
module mult_N1024_CC512 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [1:0] b;
  output [2047:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423;
  wire   [2047:0] sreg;

  DFF \sreg_reg[2045]  ( .D(c[2047]), .CLK(clk), .RST(rst), .Q(sreg[2045]) );
  DFF \sreg_reg[2044]  ( .D(c[2046]), .CLK(clk), .RST(rst), .Q(sreg[2044]) );
  DFF \sreg_reg[2043]  ( .D(c[2045]), .CLK(clk), .RST(rst), .Q(sreg[2043]) );
  DFF \sreg_reg[2042]  ( .D(c[2044]), .CLK(clk), .RST(rst), .Q(sreg[2042]) );
  DFF \sreg_reg[2041]  ( .D(c[2043]), .CLK(clk), .RST(rst), .Q(sreg[2041]) );
  DFF \sreg_reg[2040]  ( .D(c[2042]), .CLK(clk), .RST(rst), .Q(sreg[2040]) );
  DFF \sreg_reg[2039]  ( .D(c[2041]), .CLK(clk), .RST(rst), .Q(sreg[2039]) );
  DFF \sreg_reg[2038]  ( .D(c[2040]), .CLK(clk), .RST(rst), .Q(sreg[2038]) );
  DFF \sreg_reg[2037]  ( .D(c[2039]), .CLK(clk), .RST(rst), .Q(sreg[2037]) );
  DFF \sreg_reg[2036]  ( .D(c[2038]), .CLK(clk), .RST(rst), .Q(sreg[2036]) );
  DFF \sreg_reg[2035]  ( .D(c[2037]), .CLK(clk), .RST(rst), .Q(sreg[2035]) );
  DFF \sreg_reg[2034]  ( .D(c[2036]), .CLK(clk), .RST(rst), .Q(sreg[2034]) );
  DFF \sreg_reg[2033]  ( .D(c[2035]), .CLK(clk), .RST(rst), .Q(sreg[2033]) );
  DFF \sreg_reg[2032]  ( .D(c[2034]), .CLK(clk), .RST(rst), .Q(sreg[2032]) );
  DFF \sreg_reg[2031]  ( .D(c[2033]), .CLK(clk), .RST(rst), .Q(sreg[2031]) );
  DFF \sreg_reg[2030]  ( .D(c[2032]), .CLK(clk), .RST(rst), .Q(sreg[2030]) );
  DFF \sreg_reg[2029]  ( .D(c[2031]), .CLK(clk), .RST(rst), .Q(sreg[2029]) );
  DFF \sreg_reg[2028]  ( .D(c[2030]), .CLK(clk), .RST(rst), .Q(sreg[2028]) );
  DFF \sreg_reg[2027]  ( .D(c[2029]), .CLK(clk), .RST(rst), .Q(sreg[2027]) );
  DFF \sreg_reg[2026]  ( .D(c[2028]), .CLK(clk), .RST(rst), .Q(sreg[2026]) );
  DFF \sreg_reg[2025]  ( .D(c[2027]), .CLK(clk), .RST(rst), .Q(sreg[2025]) );
  DFF \sreg_reg[2024]  ( .D(c[2026]), .CLK(clk), .RST(rst), .Q(sreg[2024]) );
  DFF \sreg_reg[2023]  ( .D(c[2025]), .CLK(clk), .RST(rst), .Q(sreg[2023]) );
  DFF \sreg_reg[2022]  ( .D(c[2024]), .CLK(clk), .RST(rst), .Q(sreg[2022]) );
  DFF \sreg_reg[2021]  ( .D(c[2023]), .CLK(clk), .RST(rst), .Q(sreg[2021]) );
  DFF \sreg_reg[2020]  ( .D(c[2022]), .CLK(clk), .RST(rst), .Q(sreg[2020]) );
  DFF \sreg_reg[2019]  ( .D(c[2021]), .CLK(clk), .RST(rst), .Q(sreg[2019]) );
  DFF \sreg_reg[2018]  ( .D(c[2020]), .CLK(clk), .RST(rst), .Q(sreg[2018]) );
  DFF \sreg_reg[2017]  ( .D(c[2019]), .CLK(clk), .RST(rst), .Q(sreg[2017]) );
  DFF \sreg_reg[2016]  ( .D(c[2018]), .CLK(clk), .RST(rst), .Q(sreg[2016]) );
  DFF \sreg_reg[2015]  ( .D(c[2017]), .CLK(clk), .RST(rst), .Q(sreg[2015]) );
  DFF \sreg_reg[2014]  ( .D(c[2016]), .CLK(clk), .RST(rst), .Q(sreg[2014]) );
  DFF \sreg_reg[2013]  ( .D(c[2015]), .CLK(clk), .RST(rst), .Q(sreg[2013]) );
  DFF \sreg_reg[2012]  ( .D(c[2014]), .CLK(clk), .RST(rst), .Q(sreg[2012]) );
  DFF \sreg_reg[2011]  ( .D(c[2013]), .CLK(clk), .RST(rst), .Q(sreg[2011]) );
  DFF \sreg_reg[2010]  ( .D(c[2012]), .CLK(clk), .RST(rst), .Q(sreg[2010]) );
  DFF \sreg_reg[2009]  ( .D(c[2011]), .CLK(clk), .RST(rst), .Q(sreg[2009]) );
  DFF \sreg_reg[2008]  ( .D(c[2010]), .CLK(clk), .RST(rst), .Q(sreg[2008]) );
  DFF \sreg_reg[2007]  ( .D(c[2009]), .CLK(clk), .RST(rst), .Q(sreg[2007]) );
  DFF \sreg_reg[2006]  ( .D(c[2008]), .CLK(clk), .RST(rst), .Q(sreg[2006]) );
  DFF \sreg_reg[2005]  ( .D(c[2007]), .CLK(clk), .RST(rst), .Q(sreg[2005]) );
  DFF \sreg_reg[2004]  ( .D(c[2006]), .CLK(clk), .RST(rst), .Q(sreg[2004]) );
  DFF \sreg_reg[2003]  ( .D(c[2005]), .CLK(clk), .RST(rst), .Q(sreg[2003]) );
  DFF \sreg_reg[2002]  ( .D(c[2004]), .CLK(clk), .RST(rst), .Q(sreg[2002]) );
  DFF \sreg_reg[2001]  ( .D(c[2003]), .CLK(clk), .RST(rst), .Q(sreg[2001]) );
  DFF \sreg_reg[2000]  ( .D(c[2002]), .CLK(clk), .RST(rst), .Q(sreg[2000]) );
  DFF \sreg_reg[1999]  ( .D(c[2001]), .CLK(clk), .RST(rst), .Q(sreg[1999]) );
  DFF \sreg_reg[1998]  ( .D(c[2000]), .CLK(clk), .RST(rst), .Q(sreg[1998]) );
  DFF \sreg_reg[1997]  ( .D(c[1999]), .CLK(clk), .RST(rst), .Q(sreg[1997]) );
  DFF \sreg_reg[1996]  ( .D(c[1998]), .CLK(clk), .RST(rst), .Q(sreg[1996]) );
  DFF \sreg_reg[1995]  ( .D(c[1997]), .CLK(clk), .RST(rst), .Q(sreg[1995]) );
  DFF \sreg_reg[1994]  ( .D(c[1996]), .CLK(clk), .RST(rst), .Q(sreg[1994]) );
  DFF \sreg_reg[1993]  ( .D(c[1995]), .CLK(clk), .RST(rst), .Q(sreg[1993]) );
  DFF \sreg_reg[1992]  ( .D(c[1994]), .CLK(clk), .RST(rst), .Q(sreg[1992]) );
  DFF \sreg_reg[1991]  ( .D(c[1993]), .CLK(clk), .RST(rst), .Q(sreg[1991]) );
  DFF \sreg_reg[1990]  ( .D(c[1992]), .CLK(clk), .RST(rst), .Q(sreg[1990]) );
  DFF \sreg_reg[1989]  ( .D(c[1991]), .CLK(clk), .RST(rst), .Q(sreg[1989]) );
  DFF \sreg_reg[1988]  ( .D(c[1990]), .CLK(clk), .RST(rst), .Q(sreg[1988]) );
  DFF \sreg_reg[1987]  ( .D(c[1989]), .CLK(clk), .RST(rst), .Q(sreg[1987]) );
  DFF \sreg_reg[1986]  ( .D(c[1988]), .CLK(clk), .RST(rst), .Q(sreg[1986]) );
  DFF \sreg_reg[1985]  ( .D(c[1987]), .CLK(clk), .RST(rst), .Q(sreg[1985]) );
  DFF \sreg_reg[1984]  ( .D(c[1986]), .CLK(clk), .RST(rst), .Q(sreg[1984]) );
  DFF \sreg_reg[1983]  ( .D(c[1985]), .CLK(clk), .RST(rst), .Q(sreg[1983]) );
  DFF \sreg_reg[1982]  ( .D(c[1984]), .CLK(clk), .RST(rst), .Q(sreg[1982]) );
  DFF \sreg_reg[1981]  ( .D(c[1983]), .CLK(clk), .RST(rst), .Q(sreg[1981]) );
  DFF \sreg_reg[1980]  ( .D(c[1982]), .CLK(clk), .RST(rst), .Q(sreg[1980]) );
  DFF \sreg_reg[1979]  ( .D(c[1981]), .CLK(clk), .RST(rst), .Q(sreg[1979]) );
  DFF \sreg_reg[1978]  ( .D(c[1980]), .CLK(clk), .RST(rst), .Q(sreg[1978]) );
  DFF \sreg_reg[1977]  ( .D(c[1979]), .CLK(clk), .RST(rst), .Q(sreg[1977]) );
  DFF \sreg_reg[1976]  ( .D(c[1978]), .CLK(clk), .RST(rst), .Q(sreg[1976]) );
  DFF \sreg_reg[1975]  ( .D(c[1977]), .CLK(clk), .RST(rst), .Q(sreg[1975]) );
  DFF \sreg_reg[1974]  ( .D(c[1976]), .CLK(clk), .RST(rst), .Q(sreg[1974]) );
  DFF \sreg_reg[1973]  ( .D(c[1975]), .CLK(clk), .RST(rst), .Q(sreg[1973]) );
  DFF \sreg_reg[1972]  ( .D(c[1974]), .CLK(clk), .RST(rst), .Q(sreg[1972]) );
  DFF \sreg_reg[1971]  ( .D(c[1973]), .CLK(clk), .RST(rst), .Q(sreg[1971]) );
  DFF \sreg_reg[1970]  ( .D(c[1972]), .CLK(clk), .RST(rst), .Q(sreg[1970]) );
  DFF \sreg_reg[1969]  ( .D(c[1971]), .CLK(clk), .RST(rst), .Q(sreg[1969]) );
  DFF \sreg_reg[1968]  ( .D(c[1970]), .CLK(clk), .RST(rst), .Q(sreg[1968]) );
  DFF \sreg_reg[1967]  ( .D(c[1969]), .CLK(clk), .RST(rst), .Q(sreg[1967]) );
  DFF \sreg_reg[1966]  ( .D(c[1968]), .CLK(clk), .RST(rst), .Q(sreg[1966]) );
  DFF \sreg_reg[1965]  ( .D(c[1967]), .CLK(clk), .RST(rst), .Q(sreg[1965]) );
  DFF \sreg_reg[1964]  ( .D(c[1966]), .CLK(clk), .RST(rst), .Q(sreg[1964]) );
  DFF \sreg_reg[1963]  ( .D(c[1965]), .CLK(clk), .RST(rst), .Q(sreg[1963]) );
  DFF \sreg_reg[1962]  ( .D(c[1964]), .CLK(clk), .RST(rst), .Q(sreg[1962]) );
  DFF \sreg_reg[1961]  ( .D(c[1963]), .CLK(clk), .RST(rst), .Q(sreg[1961]) );
  DFF \sreg_reg[1960]  ( .D(c[1962]), .CLK(clk), .RST(rst), .Q(sreg[1960]) );
  DFF \sreg_reg[1959]  ( .D(c[1961]), .CLK(clk), .RST(rst), .Q(sreg[1959]) );
  DFF \sreg_reg[1958]  ( .D(c[1960]), .CLK(clk), .RST(rst), .Q(sreg[1958]) );
  DFF \sreg_reg[1957]  ( .D(c[1959]), .CLK(clk), .RST(rst), .Q(sreg[1957]) );
  DFF \sreg_reg[1956]  ( .D(c[1958]), .CLK(clk), .RST(rst), .Q(sreg[1956]) );
  DFF \sreg_reg[1955]  ( .D(c[1957]), .CLK(clk), .RST(rst), .Q(sreg[1955]) );
  DFF \sreg_reg[1954]  ( .D(c[1956]), .CLK(clk), .RST(rst), .Q(sreg[1954]) );
  DFF \sreg_reg[1953]  ( .D(c[1955]), .CLK(clk), .RST(rst), .Q(sreg[1953]) );
  DFF \sreg_reg[1952]  ( .D(c[1954]), .CLK(clk), .RST(rst), .Q(sreg[1952]) );
  DFF \sreg_reg[1951]  ( .D(c[1953]), .CLK(clk), .RST(rst), .Q(sreg[1951]) );
  DFF \sreg_reg[1950]  ( .D(c[1952]), .CLK(clk), .RST(rst), .Q(sreg[1950]) );
  DFF \sreg_reg[1949]  ( .D(c[1951]), .CLK(clk), .RST(rst), .Q(sreg[1949]) );
  DFF \sreg_reg[1948]  ( .D(c[1950]), .CLK(clk), .RST(rst), .Q(sreg[1948]) );
  DFF \sreg_reg[1947]  ( .D(c[1949]), .CLK(clk), .RST(rst), .Q(sreg[1947]) );
  DFF \sreg_reg[1946]  ( .D(c[1948]), .CLK(clk), .RST(rst), .Q(sreg[1946]) );
  DFF \sreg_reg[1945]  ( .D(c[1947]), .CLK(clk), .RST(rst), .Q(sreg[1945]) );
  DFF \sreg_reg[1944]  ( .D(c[1946]), .CLK(clk), .RST(rst), .Q(sreg[1944]) );
  DFF \sreg_reg[1943]  ( .D(c[1945]), .CLK(clk), .RST(rst), .Q(sreg[1943]) );
  DFF \sreg_reg[1942]  ( .D(c[1944]), .CLK(clk), .RST(rst), .Q(sreg[1942]) );
  DFF \sreg_reg[1941]  ( .D(c[1943]), .CLK(clk), .RST(rst), .Q(sreg[1941]) );
  DFF \sreg_reg[1940]  ( .D(c[1942]), .CLK(clk), .RST(rst), .Q(sreg[1940]) );
  DFF \sreg_reg[1939]  ( .D(c[1941]), .CLK(clk), .RST(rst), .Q(sreg[1939]) );
  DFF \sreg_reg[1938]  ( .D(c[1940]), .CLK(clk), .RST(rst), .Q(sreg[1938]) );
  DFF \sreg_reg[1937]  ( .D(c[1939]), .CLK(clk), .RST(rst), .Q(sreg[1937]) );
  DFF \sreg_reg[1936]  ( .D(c[1938]), .CLK(clk), .RST(rst), .Q(sreg[1936]) );
  DFF \sreg_reg[1935]  ( .D(c[1937]), .CLK(clk), .RST(rst), .Q(sreg[1935]) );
  DFF \sreg_reg[1934]  ( .D(c[1936]), .CLK(clk), .RST(rst), .Q(sreg[1934]) );
  DFF \sreg_reg[1933]  ( .D(c[1935]), .CLK(clk), .RST(rst), .Q(sreg[1933]) );
  DFF \sreg_reg[1932]  ( .D(c[1934]), .CLK(clk), .RST(rst), .Q(sreg[1932]) );
  DFF \sreg_reg[1931]  ( .D(c[1933]), .CLK(clk), .RST(rst), .Q(sreg[1931]) );
  DFF \sreg_reg[1930]  ( .D(c[1932]), .CLK(clk), .RST(rst), .Q(sreg[1930]) );
  DFF \sreg_reg[1929]  ( .D(c[1931]), .CLK(clk), .RST(rst), .Q(sreg[1929]) );
  DFF \sreg_reg[1928]  ( .D(c[1930]), .CLK(clk), .RST(rst), .Q(sreg[1928]) );
  DFF \sreg_reg[1927]  ( .D(c[1929]), .CLK(clk), .RST(rst), .Q(sreg[1927]) );
  DFF \sreg_reg[1926]  ( .D(c[1928]), .CLK(clk), .RST(rst), .Q(sreg[1926]) );
  DFF \sreg_reg[1925]  ( .D(c[1927]), .CLK(clk), .RST(rst), .Q(sreg[1925]) );
  DFF \sreg_reg[1924]  ( .D(c[1926]), .CLK(clk), .RST(rst), .Q(sreg[1924]) );
  DFF \sreg_reg[1923]  ( .D(c[1925]), .CLK(clk), .RST(rst), .Q(sreg[1923]) );
  DFF \sreg_reg[1922]  ( .D(c[1924]), .CLK(clk), .RST(rst), .Q(sreg[1922]) );
  DFF \sreg_reg[1921]  ( .D(c[1923]), .CLK(clk), .RST(rst), .Q(sreg[1921]) );
  DFF \sreg_reg[1920]  ( .D(c[1922]), .CLK(clk), .RST(rst), .Q(sreg[1920]) );
  DFF \sreg_reg[1919]  ( .D(c[1921]), .CLK(clk), .RST(rst), .Q(sreg[1919]) );
  DFF \sreg_reg[1918]  ( .D(c[1920]), .CLK(clk), .RST(rst), .Q(sreg[1918]) );
  DFF \sreg_reg[1917]  ( .D(c[1919]), .CLK(clk), .RST(rst), .Q(sreg[1917]) );
  DFF \sreg_reg[1916]  ( .D(c[1918]), .CLK(clk), .RST(rst), .Q(sreg[1916]) );
  DFF \sreg_reg[1915]  ( .D(c[1917]), .CLK(clk), .RST(rst), .Q(sreg[1915]) );
  DFF \sreg_reg[1914]  ( .D(c[1916]), .CLK(clk), .RST(rst), .Q(sreg[1914]) );
  DFF \sreg_reg[1913]  ( .D(c[1915]), .CLK(clk), .RST(rst), .Q(sreg[1913]) );
  DFF \sreg_reg[1912]  ( .D(c[1914]), .CLK(clk), .RST(rst), .Q(sreg[1912]) );
  DFF \sreg_reg[1911]  ( .D(c[1913]), .CLK(clk), .RST(rst), .Q(sreg[1911]) );
  DFF \sreg_reg[1910]  ( .D(c[1912]), .CLK(clk), .RST(rst), .Q(sreg[1910]) );
  DFF \sreg_reg[1909]  ( .D(c[1911]), .CLK(clk), .RST(rst), .Q(sreg[1909]) );
  DFF \sreg_reg[1908]  ( .D(c[1910]), .CLK(clk), .RST(rst), .Q(sreg[1908]) );
  DFF \sreg_reg[1907]  ( .D(c[1909]), .CLK(clk), .RST(rst), .Q(sreg[1907]) );
  DFF \sreg_reg[1906]  ( .D(c[1908]), .CLK(clk), .RST(rst), .Q(sreg[1906]) );
  DFF \sreg_reg[1905]  ( .D(c[1907]), .CLK(clk), .RST(rst), .Q(sreg[1905]) );
  DFF \sreg_reg[1904]  ( .D(c[1906]), .CLK(clk), .RST(rst), .Q(sreg[1904]) );
  DFF \sreg_reg[1903]  ( .D(c[1905]), .CLK(clk), .RST(rst), .Q(sreg[1903]) );
  DFF \sreg_reg[1902]  ( .D(c[1904]), .CLK(clk), .RST(rst), .Q(sreg[1902]) );
  DFF \sreg_reg[1901]  ( .D(c[1903]), .CLK(clk), .RST(rst), .Q(sreg[1901]) );
  DFF \sreg_reg[1900]  ( .D(c[1902]), .CLK(clk), .RST(rst), .Q(sreg[1900]) );
  DFF \sreg_reg[1899]  ( .D(c[1901]), .CLK(clk), .RST(rst), .Q(sreg[1899]) );
  DFF \sreg_reg[1898]  ( .D(c[1900]), .CLK(clk), .RST(rst), .Q(sreg[1898]) );
  DFF \sreg_reg[1897]  ( .D(c[1899]), .CLK(clk), .RST(rst), .Q(sreg[1897]) );
  DFF \sreg_reg[1896]  ( .D(c[1898]), .CLK(clk), .RST(rst), .Q(sreg[1896]) );
  DFF \sreg_reg[1895]  ( .D(c[1897]), .CLK(clk), .RST(rst), .Q(sreg[1895]) );
  DFF \sreg_reg[1894]  ( .D(c[1896]), .CLK(clk), .RST(rst), .Q(sreg[1894]) );
  DFF \sreg_reg[1893]  ( .D(c[1895]), .CLK(clk), .RST(rst), .Q(sreg[1893]) );
  DFF \sreg_reg[1892]  ( .D(c[1894]), .CLK(clk), .RST(rst), .Q(sreg[1892]) );
  DFF \sreg_reg[1891]  ( .D(c[1893]), .CLK(clk), .RST(rst), .Q(sreg[1891]) );
  DFF \sreg_reg[1890]  ( .D(c[1892]), .CLK(clk), .RST(rst), .Q(sreg[1890]) );
  DFF \sreg_reg[1889]  ( .D(c[1891]), .CLK(clk), .RST(rst), .Q(sreg[1889]) );
  DFF \sreg_reg[1888]  ( .D(c[1890]), .CLK(clk), .RST(rst), .Q(sreg[1888]) );
  DFF \sreg_reg[1887]  ( .D(c[1889]), .CLK(clk), .RST(rst), .Q(sreg[1887]) );
  DFF \sreg_reg[1886]  ( .D(c[1888]), .CLK(clk), .RST(rst), .Q(sreg[1886]) );
  DFF \sreg_reg[1885]  ( .D(c[1887]), .CLK(clk), .RST(rst), .Q(sreg[1885]) );
  DFF \sreg_reg[1884]  ( .D(c[1886]), .CLK(clk), .RST(rst), .Q(sreg[1884]) );
  DFF \sreg_reg[1883]  ( .D(c[1885]), .CLK(clk), .RST(rst), .Q(sreg[1883]) );
  DFF \sreg_reg[1882]  ( .D(c[1884]), .CLK(clk), .RST(rst), .Q(sreg[1882]) );
  DFF \sreg_reg[1881]  ( .D(c[1883]), .CLK(clk), .RST(rst), .Q(sreg[1881]) );
  DFF \sreg_reg[1880]  ( .D(c[1882]), .CLK(clk), .RST(rst), .Q(sreg[1880]) );
  DFF \sreg_reg[1879]  ( .D(c[1881]), .CLK(clk), .RST(rst), .Q(sreg[1879]) );
  DFF \sreg_reg[1878]  ( .D(c[1880]), .CLK(clk), .RST(rst), .Q(sreg[1878]) );
  DFF \sreg_reg[1877]  ( .D(c[1879]), .CLK(clk), .RST(rst), .Q(sreg[1877]) );
  DFF \sreg_reg[1876]  ( .D(c[1878]), .CLK(clk), .RST(rst), .Q(sreg[1876]) );
  DFF \sreg_reg[1875]  ( .D(c[1877]), .CLK(clk), .RST(rst), .Q(sreg[1875]) );
  DFF \sreg_reg[1874]  ( .D(c[1876]), .CLK(clk), .RST(rst), .Q(sreg[1874]) );
  DFF \sreg_reg[1873]  ( .D(c[1875]), .CLK(clk), .RST(rst), .Q(sreg[1873]) );
  DFF \sreg_reg[1872]  ( .D(c[1874]), .CLK(clk), .RST(rst), .Q(sreg[1872]) );
  DFF \sreg_reg[1871]  ( .D(c[1873]), .CLK(clk), .RST(rst), .Q(sreg[1871]) );
  DFF \sreg_reg[1870]  ( .D(c[1872]), .CLK(clk), .RST(rst), .Q(sreg[1870]) );
  DFF \sreg_reg[1869]  ( .D(c[1871]), .CLK(clk), .RST(rst), .Q(sreg[1869]) );
  DFF \sreg_reg[1868]  ( .D(c[1870]), .CLK(clk), .RST(rst), .Q(sreg[1868]) );
  DFF \sreg_reg[1867]  ( .D(c[1869]), .CLK(clk), .RST(rst), .Q(sreg[1867]) );
  DFF \sreg_reg[1866]  ( .D(c[1868]), .CLK(clk), .RST(rst), .Q(sreg[1866]) );
  DFF \sreg_reg[1865]  ( .D(c[1867]), .CLK(clk), .RST(rst), .Q(sreg[1865]) );
  DFF \sreg_reg[1864]  ( .D(c[1866]), .CLK(clk), .RST(rst), .Q(sreg[1864]) );
  DFF \sreg_reg[1863]  ( .D(c[1865]), .CLK(clk), .RST(rst), .Q(sreg[1863]) );
  DFF \sreg_reg[1862]  ( .D(c[1864]), .CLK(clk), .RST(rst), .Q(sreg[1862]) );
  DFF \sreg_reg[1861]  ( .D(c[1863]), .CLK(clk), .RST(rst), .Q(sreg[1861]) );
  DFF \sreg_reg[1860]  ( .D(c[1862]), .CLK(clk), .RST(rst), .Q(sreg[1860]) );
  DFF \sreg_reg[1859]  ( .D(c[1861]), .CLK(clk), .RST(rst), .Q(sreg[1859]) );
  DFF \sreg_reg[1858]  ( .D(c[1860]), .CLK(clk), .RST(rst), .Q(sreg[1858]) );
  DFF \sreg_reg[1857]  ( .D(c[1859]), .CLK(clk), .RST(rst), .Q(sreg[1857]) );
  DFF \sreg_reg[1856]  ( .D(c[1858]), .CLK(clk), .RST(rst), .Q(sreg[1856]) );
  DFF \sreg_reg[1855]  ( .D(c[1857]), .CLK(clk), .RST(rst), .Q(sreg[1855]) );
  DFF \sreg_reg[1854]  ( .D(c[1856]), .CLK(clk), .RST(rst), .Q(sreg[1854]) );
  DFF \sreg_reg[1853]  ( .D(c[1855]), .CLK(clk), .RST(rst), .Q(sreg[1853]) );
  DFF \sreg_reg[1852]  ( .D(c[1854]), .CLK(clk), .RST(rst), .Q(sreg[1852]) );
  DFF \sreg_reg[1851]  ( .D(c[1853]), .CLK(clk), .RST(rst), .Q(sreg[1851]) );
  DFF \sreg_reg[1850]  ( .D(c[1852]), .CLK(clk), .RST(rst), .Q(sreg[1850]) );
  DFF \sreg_reg[1849]  ( .D(c[1851]), .CLK(clk), .RST(rst), .Q(sreg[1849]) );
  DFF \sreg_reg[1848]  ( .D(c[1850]), .CLK(clk), .RST(rst), .Q(sreg[1848]) );
  DFF \sreg_reg[1847]  ( .D(c[1849]), .CLK(clk), .RST(rst), .Q(sreg[1847]) );
  DFF \sreg_reg[1846]  ( .D(c[1848]), .CLK(clk), .RST(rst), .Q(sreg[1846]) );
  DFF \sreg_reg[1845]  ( .D(c[1847]), .CLK(clk), .RST(rst), .Q(sreg[1845]) );
  DFF \sreg_reg[1844]  ( .D(c[1846]), .CLK(clk), .RST(rst), .Q(sreg[1844]) );
  DFF \sreg_reg[1843]  ( .D(c[1845]), .CLK(clk), .RST(rst), .Q(sreg[1843]) );
  DFF \sreg_reg[1842]  ( .D(c[1844]), .CLK(clk), .RST(rst), .Q(sreg[1842]) );
  DFF \sreg_reg[1841]  ( .D(c[1843]), .CLK(clk), .RST(rst), .Q(sreg[1841]) );
  DFF \sreg_reg[1840]  ( .D(c[1842]), .CLK(clk), .RST(rst), .Q(sreg[1840]) );
  DFF \sreg_reg[1839]  ( .D(c[1841]), .CLK(clk), .RST(rst), .Q(sreg[1839]) );
  DFF \sreg_reg[1838]  ( .D(c[1840]), .CLK(clk), .RST(rst), .Q(sreg[1838]) );
  DFF \sreg_reg[1837]  ( .D(c[1839]), .CLK(clk), .RST(rst), .Q(sreg[1837]) );
  DFF \sreg_reg[1836]  ( .D(c[1838]), .CLK(clk), .RST(rst), .Q(sreg[1836]) );
  DFF \sreg_reg[1835]  ( .D(c[1837]), .CLK(clk), .RST(rst), .Q(sreg[1835]) );
  DFF \sreg_reg[1834]  ( .D(c[1836]), .CLK(clk), .RST(rst), .Q(sreg[1834]) );
  DFF \sreg_reg[1833]  ( .D(c[1835]), .CLK(clk), .RST(rst), .Q(sreg[1833]) );
  DFF \sreg_reg[1832]  ( .D(c[1834]), .CLK(clk), .RST(rst), .Q(sreg[1832]) );
  DFF \sreg_reg[1831]  ( .D(c[1833]), .CLK(clk), .RST(rst), .Q(sreg[1831]) );
  DFF \sreg_reg[1830]  ( .D(c[1832]), .CLK(clk), .RST(rst), .Q(sreg[1830]) );
  DFF \sreg_reg[1829]  ( .D(c[1831]), .CLK(clk), .RST(rst), .Q(sreg[1829]) );
  DFF \sreg_reg[1828]  ( .D(c[1830]), .CLK(clk), .RST(rst), .Q(sreg[1828]) );
  DFF \sreg_reg[1827]  ( .D(c[1829]), .CLK(clk), .RST(rst), .Q(sreg[1827]) );
  DFF \sreg_reg[1826]  ( .D(c[1828]), .CLK(clk), .RST(rst), .Q(sreg[1826]) );
  DFF \sreg_reg[1825]  ( .D(c[1827]), .CLK(clk), .RST(rst), .Q(sreg[1825]) );
  DFF \sreg_reg[1824]  ( .D(c[1826]), .CLK(clk), .RST(rst), .Q(sreg[1824]) );
  DFF \sreg_reg[1823]  ( .D(c[1825]), .CLK(clk), .RST(rst), .Q(sreg[1823]) );
  DFF \sreg_reg[1822]  ( .D(c[1824]), .CLK(clk), .RST(rst), .Q(sreg[1822]) );
  DFF \sreg_reg[1821]  ( .D(c[1823]), .CLK(clk), .RST(rst), .Q(sreg[1821]) );
  DFF \sreg_reg[1820]  ( .D(c[1822]), .CLK(clk), .RST(rst), .Q(sreg[1820]) );
  DFF \sreg_reg[1819]  ( .D(c[1821]), .CLK(clk), .RST(rst), .Q(sreg[1819]) );
  DFF \sreg_reg[1818]  ( .D(c[1820]), .CLK(clk), .RST(rst), .Q(sreg[1818]) );
  DFF \sreg_reg[1817]  ( .D(c[1819]), .CLK(clk), .RST(rst), .Q(sreg[1817]) );
  DFF \sreg_reg[1816]  ( .D(c[1818]), .CLK(clk), .RST(rst), .Q(sreg[1816]) );
  DFF \sreg_reg[1815]  ( .D(c[1817]), .CLK(clk), .RST(rst), .Q(sreg[1815]) );
  DFF \sreg_reg[1814]  ( .D(c[1816]), .CLK(clk), .RST(rst), .Q(sreg[1814]) );
  DFF \sreg_reg[1813]  ( .D(c[1815]), .CLK(clk), .RST(rst), .Q(sreg[1813]) );
  DFF \sreg_reg[1812]  ( .D(c[1814]), .CLK(clk), .RST(rst), .Q(sreg[1812]) );
  DFF \sreg_reg[1811]  ( .D(c[1813]), .CLK(clk), .RST(rst), .Q(sreg[1811]) );
  DFF \sreg_reg[1810]  ( .D(c[1812]), .CLK(clk), .RST(rst), .Q(sreg[1810]) );
  DFF \sreg_reg[1809]  ( .D(c[1811]), .CLK(clk), .RST(rst), .Q(sreg[1809]) );
  DFF \sreg_reg[1808]  ( .D(c[1810]), .CLK(clk), .RST(rst), .Q(sreg[1808]) );
  DFF \sreg_reg[1807]  ( .D(c[1809]), .CLK(clk), .RST(rst), .Q(sreg[1807]) );
  DFF \sreg_reg[1806]  ( .D(c[1808]), .CLK(clk), .RST(rst), .Q(sreg[1806]) );
  DFF \sreg_reg[1805]  ( .D(c[1807]), .CLK(clk), .RST(rst), .Q(sreg[1805]) );
  DFF \sreg_reg[1804]  ( .D(c[1806]), .CLK(clk), .RST(rst), .Q(sreg[1804]) );
  DFF \sreg_reg[1803]  ( .D(c[1805]), .CLK(clk), .RST(rst), .Q(sreg[1803]) );
  DFF \sreg_reg[1802]  ( .D(c[1804]), .CLK(clk), .RST(rst), .Q(sreg[1802]) );
  DFF \sreg_reg[1801]  ( .D(c[1803]), .CLK(clk), .RST(rst), .Q(sreg[1801]) );
  DFF \sreg_reg[1800]  ( .D(c[1802]), .CLK(clk), .RST(rst), .Q(sreg[1800]) );
  DFF \sreg_reg[1799]  ( .D(c[1801]), .CLK(clk), .RST(rst), .Q(sreg[1799]) );
  DFF \sreg_reg[1798]  ( .D(c[1800]), .CLK(clk), .RST(rst), .Q(sreg[1798]) );
  DFF \sreg_reg[1797]  ( .D(c[1799]), .CLK(clk), .RST(rst), .Q(sreg[1797]) );
  DFF \sreg_reg[1796]  ( .D(c[1798]), .CLK(clk), .RST(rst), .Q(sreg[1796]) );
  DFF \sreg_reg[1795]  ( .D(c[1797]), .CLK(clk), .RST(rst), .Q(sreg[1795]) );
  DFF \sreg_reg[1794]  ( .D(c[1796]), .CLK(clk), .RST(rst), .Q(sreg[1794]) );
  DFF \sreg_reg[1793]  ( .D(c[1795]), .CLK(clk), .RST(rst), .Q(sreg[1793]) );
  DFF \sreg_reg[1792]  ( .D(c[1794]), .CLK(clk), .RST(rst), .Q(sreg[1792]) );
  DFF \sreg_reg[1791]  ( .D(c[1793]), .CLK(clk), .RST(rst), .Q(sreg[1791]) );
  DFF \sreg_reg[1790]  ( .D(c[1792]), .CLK(clk), .RST(rst), .Q(sreg[1790]) );
  DFF \sreg_reg[1789]  ( .D(c[1791]), .CLK(clk), .RST(rst), .Q(sreg[1789]) );
  DFF \sreg_reg[1788]  ( .D(c[1790]), .CLK(clk), .RST(rst), .Q(sreg[1788]) );
  DFF \sreg_reg[1787]  ( .D(c[1789]), .CLK(clk), .RST(rst), .Q(sreg[1787]) );
  DFF \sreg_reg[1786]  ( .D(c[1788]), .CLK(clk), .RST(rst), .Q(sreg[1786]) );
  DFF \sreg_reg[1785]  ( .D(c[1787]), .CLK(clk), .RST(rst), .Q(sreg[1785]) );
  DFF \sreg_reg[1784]  ( .D(c[1786]), .CLK(clk), .RST(rst), .Q(sreg[1784]) );
  DFF \sreg_reg[1783]  ( .D(c[1785]), .CLK(clk), .RST(rst), .Q(sreg[1783]) );
  DFF \sreg_reg[1782]  ( .D(c[1784]), .CLK(clk), .RST(rst), .Q(sreg[1782]) );
  DFF \sreg_reg[1781]  ( .D(c[1783]), .CLK(clk), .RST(rst), .Q(sreg[1781]) );
  DFF \sreg_reg[1780]  ( .D(c[1782]), .CLK(clk), .RST(rst), .Q(sreg[1780]) );
  DFF \sreg_reg[1779]  ( .D(c[1781]), .CLK(clk), .RST(rst), .Q(sreg[1779]) );
  DFF \sreg_reg[1778]  ( .D(c[1780]), .CLK(clk), .RST(rst), .Q(sreg[1778]) );
  DFF \sreg_reg[1777]  ( .D(c[1779]), .CLK(clk), .RST(rst), .Q(sreg[1777]) );
  DFF \sreg_reg[1776]  ( .D(c[1778]), .CLK(clk), .RST(rst), .Q(sreg[1776]) );
  DFF \sreg_reg[1775]  ( .D(c[1777]), .CLK(clk), .RST(rst), .Q(sreg[1775]) );
  DFF \sreg_reg[1774]  ( .D(c[1776]), .CLK(clk), .RST(rst), .Q(sreg[1774]) );
  DFF \sreg_reg[1773]  ( .D(c[1775]), .CLK(clk), .RST(rst), .Q(sreg[1773]) );
  DFF \sreg_reg[1772]  ( .D(c[1774]), .CLK(clk), .RST(rst), .Q(sreg[1772]) );
  DFF \sreg_reg[1771]  ( .D(c[1773]), .CLK(clk), .RST(rst), .Q(sreg[1771]) );
  DFF \sreg_reg[1770]  ( .D(c[1772]), .CLK(clk), .RST(rst), .Q(sreg[1770]) );
  DFF \sreg_reg[1769]  ( .D(c[1771]), .CLK(clk), .RST(rst), .Q(sreg[1769]) );
  DFF \sreg_reg[1768]  ( .D(c[1770]), .CLK(clk), .RST(rst), .Q(sreg[1768]) );
  DFF \sreg_reg[1767]  ( .D(c[1769]), .CLK(clk), .RST(rst), .Q(sreg[1767]) );
  DFF \sreg_reg[1766]  ( .D(c[1768]), .CLK(clk), .RST(rst), .Q(sreg[1766]) );
  DFF \sreg_reg[1765]  ( .D(c[1767]), .CLK(clk), .RST(rst), .Q(sreg[1765]) );
  DFF \sreg_reg[1764]  ( .D(c[1766]), .CLK(clk), .RST(rst), .Q(sreg[1764]) );
  DFF \sreg_reg[1763]  ( .D(c[1765]), .CLK(clk), .RST(rst), .Q(sreg[1763]) );
  DFF \sreg_reg[1762]  ( .D(c[1764]), .CLK(clk), .RST(rst), .Q(sreg[1762]) );
  DFF \sreg_reg[1761]  ( .D(c[1763]), .CLK(clk), .RST(rst), .Q(sreg[1761]) );
  DFF \sreg_reg[1760]  ( .D(c[1762]), .CLK(clk), .RST(rst), .Q(sreg[1760]) );
  DFF \sreg_reg[1759]  ( .D(c[1761]), .CLK(clk), .RST(rst), .Q(sreg[1759]) );
  DFF \sreg_reg[1758]  ( .D(c[1760]), .CLK(clk), .RST(rst), .Q(sreg[1758]) );
  DFF \sreg_reg[1757]  ( .D(c[1759]), .CLK(clk), .RST(rst), .Q(sreg[1757]) );
  DFF \sreg_reg[1756]  ( .D(c[1758]), .CLK(clk), .RST(rst), .Q(sreg[1756]) );
  DFF \sreg_reg[1755]  ( .D(c[1757]), .CLK(clk), .RST(rst), .Q(sreg[1755]) );
  DFF \sreg_reg[1754]  ( .D(c[1756]), .CLK(clk), .RST(rst), .Q(sreg[1754]) );
  DFF \sreg_reg[1753]  ( .D(c[1755]), .CLK(clk), .RST(rst), .Q(sreg[1753]) );
  DFF \sreg_reg[1752]  ( .D(c[1754]), .CLK(clk), .RST(rst), .Q(sreg[1752]) );
  DFF \sreg_reg[1751]  ( .D(c[1753]), .CLK(clk), .RST(rst), .Q(sreg[1751]) );
  DFF \sreg_reg[1750]  ( .D(c[1752]), .CLK(clk), .RST(rst), .Q(sreg[1750]) );
  DFF \sreg_reg[1749]  ( .D(c[1751]), .CLK(clk), .RST(rst), .Q(sreg[1749]) );
  DFF \sreg_reg[1748]  ( .D(c[1750]), .CLK(clk), .RST(rst), .Q(sreg[1748]) );
  DFF \sreg_reg[1747]  ( .D(c[1749]), .CLK(clk), .RST(rst), .Q(sreg[1747]) );
  DFF \sreg_reg[1746]  ( .D(c[1748]), .CLK(clk), .RST(rst), .Q(sreg[1746]) );
  DFF \sreg_reg[1745]  ( .D(c[1747]), .CLK(clk), .RST(rst), .Q(sreg[1745]) );
  DFF \sreg_reg[1744]  ( .D(c[1746]), .CLK(clk), .RST(rst), .Q(sreg[1744]) );
  DFF \sreg_reg[1743]  ( .D(c[1745]), .CLK(clk), .RST(rst), .Q(sreg[1743]) );
  DFF \sreg_reg[1742]  ( .D(c[1744]), .CLK(clk), .RST(rst), .Q(sreg[1742]) );
  DFF \sreg_reg[1741]  ( .D(c[1743]), .CLK(clk), .RST(rst), .Q(sreg[1741]) );
  DFF \sreg_reg[1740]  ( .D(c[1742]), .CLK(clk), .RST(rst), .Q(sreg[1740]) );
  DFF \sreg_reg[1739]  ( .D(c[1741]), .CLK(clk), .RST(rst), .Q(sreg[1739]) );
  DFF \sreg_reg[1738]  ( .D(c[1740]), .CLK(clk), .RST(rst), .Q(sreg[1738]) );
  DFF \sreg_reg[1737]  ( .D(c[1739]), .CLK(clk), .RST(rst), .Q(sreg[1737]) );
  DFF \sreg_reg[1736]  ( .D(c[1738]), .CLK(clk), .RST(rst), .Q(sreg[1736]) );
  DFF \sreg_reg[1735]  ( .D(c[1737]), .CLK(clk), .RST(rst), .Q(sreg[1735]) );
  DFF \sreg_reg[1734]  ( .D(c[1736]), .CLK(clk), .RST(rst), .Q(sreg[1734]) );
  DFF \sreg_reg[1733]  ( .D(c[1735]), .CLK(clk), .RST(rst), .Q(sreg[1733]) );
  DFF \sreg_reg[1732]  ( .D(c[1734]), .CLK(clk), .RST(rst), .Q(sreg[1732]) );
  DFF \sreg_reg[1731]  ( .D(c[1733]), .CLK(clk), .RST(rst), .Q(sreg[1731]) );
  DFF \sreg_reg[1730]  ( .D(c[1732]), .CLK(clk), .RST(rst), .Q(sreg[1730]) );
  DFF \sreg_reg[1729]  ( .D(c[1731]), .CLK(clk), .RST(rst), .Q(sreg[1729]) );
  DFF \sreg_reg[1728]  ( .D(c[1730]), .CLK(clk), .RST(rst), .Q(sreg[1728]) );
  DFF \sreg_reg[1727]  ( .D(c[1729]), .CLK(clk), .RST(rst), .Q(sreg[1727]) );
  DFF \sreg_reg[1726]  ( .D(c[1728]), .CLK(clk), .RST(rst), .Q(sreg[1726]) );
  DFF \sreg_reg[1725]  ( .D(c[1727]), .CLK(clk), .RST(rst), .Q(sreg[1725]) );
  DFF \sreg_reg[1724]  ( .D(c[1726]), .CLK(clk), .RST(rst), .Q(sreg[1724]) );
  DFF \sreg_reg[1723]  ( .D(c[1725]), .CLK(clk), .RST(rst), .Q(sreg[1723]) );
  DFF \sreg_reg[1722]  ( .D(c[1724]), .CLK(clk), .RST(rst), .Q(sreg[1722]) );
  DFF \sreg_reg[1721]  ( .D(c[1723]), .CLK(clk), .RST(rst), .Q(sreg[1721]) );
  DFF \sreg_reg[1720]  ( .D(c[1722]), .CLK(clk), .RST(rst), .Q(sreg[1720]) );
  DFF \sreg_reg[1719]  ( .D(c[1721]), .CLK(clk), .RST(rst), .Q(sreg[1719]) );
  DFF \sreg_reg[1718]  ( .D(c[1720]), .CLK(clk), .RST(rst), .Q(sreg[1718]) );
  DFF \sreg_reg[1717]  ( .D(c[1719]), .CLK(clk), .RST(rst), .Q(sreg[1717]) );
  DFF \sreg_reg[1716]  ( .D(c[1718]), .CLK(clk), .RST(rst), .Q(sreg[1716]) );
  DFF \sreg_reg[1715]  ( .D(c[1717]), .CLK(clk), .RST(rst), .Q(sreg[1715]) );
  DFF \sreg_reg[1714]  ( .D(c[1716]), .CLK(clk), .RST(rst), .Q(sreg[1714]) );
  DFF \sreg_reg[1713]  ( .D(c[1715]), .CLK(clk), .RST(rst), .Q(sreg[1713]) );
  DFF \sreg_reg[1712]  ( .D(c[1714]), .CLK(clk), .RST(rst), .Q(sreg[1712]) );
  DFF \sreg_reg[1711]  ( .D(c[1713]), .CLK(clk), .RST(rst), .Q(sreg[1711]) );
  DFF \sreg_reg[1710]  ( .D(c[1712]), .CLK(clk), .RST(rst), .Q(sreg[1710]) );
  DFF \sreg_reg[1709]  ( .D(c[1711]), .CLK(clk), .RST(rst), .Q(sreg[1709]) );
  DFF \sreg_reg[1708]  ( .D(c[1710]), .CLK(clk), .RST(rst), .Q(sreg[1708]) );
  DFF \sreg_reg[1707]  ( .D(c[1709]), .CLK(clk), .RST(rst), .Q(sreg[1707]) );
  DFF \sreg_reg[1706]  ( .D(c[1708]), .CLK(clk), .RST(rst), .Q(sreg[1706]) );
  DFF \sreg_reg[1705]  ( .D(c[1707]), .CLK(clk), .RST(rst), .Q(sreg[1705]) );
  DFF \sreg_reg[1704]  ( .D(c[1706]), .CLK(clk), .RST(rst), .Q(sreg[1704]) );
  DFF \sreg_reg[1703]  ( .D(c[1705]), .CLK(clk), .RST(rst), .Q(sreg[1703]) );
  DFF \sreg_reg[1702]  ( .D(c[1704]), .CLK(clk), .RST(rst), .Q(sreg[1702]) );
  DFF \sreg_reg[1701]  ( .D(c[1703]), .CLK(clk), .RST(rst), .Q(sreg[1701]) );
  DFF \sreg_reg[1700]  ( .D(c[1702]), .CLK(clk), .RST(rst), .Q(sreg[1700]) );
  DFF \sreg_reg[1699]  ( .D(c[1701]), .CLK(clk), .RST(rst), .Q(sreg[1699]) );
  DFF \sreg_reg[1698]  ( .D(c[1700]), .CLK(clk), .RST(rst), .Q(sreg[1698]) );
  DFF \sreg_reg[1697]  ( .D(c[1699]), .CLK(clk), .RST(rst), .Q(sreg[1697]) );
  DFF \sreg_reg[1696]  ( .D(c[1698]), .CLK(clk), .RST(rst), .Q(sreg[1696]) );
  DFF \sreg_reg[1695]  ( .D(c[1697]), .CLK(clk), .RST(rst), .Q(sreg[1695]) );
  DFF \sreg_reg[1694]  ( .D(c[1696]), .CLK(clk), .RST(rst), .Q(sreg[1694]) );
  DFF \sreg_reg[1693]  ( .D(c[1695]), .CLK(clk), .RST(rst), .Q(sreg[1693]) );
  DFF \sreg_reg[1692]  ( .D(c[1694]), .CLK(clk), .RST(rst), .Q(sreg[1692]) );
  DFF \sreg_reg[1691]  ( .D(c[1693]), .CLK(clk), .RST(rst), .Q(sreg[1691]) );
  DFF \sreg_reg[1690]  ( .D(c[1692]), .CLK(clk), .RST(rst), .Q(sreg[1690]) );
  DFF \sreg_reg[1689]  ( .D(c[1691]), .CLK(clk), .RST(rst), .Q(sreg[1689]) );
  DFF \sreg_reg[1688]  ( .D(c[1690]), .CLK(clk), .RST(rst), .Q(sreg[1688]) );
  DFF \sreg_reg[1687]  ( .D(c[1689]), .CLK(clk), .RST(rst), .Q(sreg[1687]) );
  DFF \sreg_reg[1686]  ( .D(c[1688]), .CLK(clk), .RST(rst), .Q(sreg[1686]) );
  DFF \sreg_reg[1685]  ( .D(c[1687]), .CLK(clk), .RST(rst), .Q(sreg[1685]) );
  DFF \sreg_reg[1684]  ( .D(c[1686]), .CLK(clk), .RST(rst), .Q(sreg[1684]) );
  DFF \sreg_reg[1683]  ( .D(c[1685]), .CLK(clk), .RST(rst), .Q(sreg[1683]) );
  DFF \sreg_reg[1682]  ( .D(c[1684]), .CLK(clk), .RST(rst), .Q(sreg[1682]) );
  DFF \sreg_reg[1681]  ( .D(c[1683]), .CLK(clk), .RST(rst), .Q(sreg[1681]) );
  DFF \sreg_reg[1680]  ( .D(c[1682]), .CLK(clk), .RST(rst), .Q(sreg[1680]) );
  DFF \sreg_reg[1679]  ( .D(c[1681]), .CLK(clk), .RST(rst), .Q(sreg[1679]) );
  DFF \sreg_reg[1678]  ( .D(c[1680]), .CLK(clk), .RST(rst), .Q(sreg[1678]) );
  DFF \sreg_reg[1677]  ( .D(c[1679]), .CLK(clk), .RST(rst), .Q(sreg[1677]) );
  DFF \sreg_reg[1676]  ( .D(c[1678]), .CLK(clk), .RST(rst), .Q(sreg[1676]) );
  DFF \sreg_reg[1675]  ( .D(c[1677]), .CLK(clk), .RST(rst), .Q(sreg[1675]) );
  DFF \sreg_reg[1674]  ( .D(c[1676]), .CLK(clk), .RST(rst), .Q(sreg[1674]) );
  DFF \sreg_reg[1673]  ( .D(c[1675]), .CLK(clk), .RST(rst), .Q(sreg[1673]) );
  DFF \sreg_reg[1672]  ( .D(c[1674]), .CLK(clk), .RST(rst), .Q(sreg[1672]) );
  DFF \sreg_reg[1671]  ( .D(c[1673]), .CLK(clk), .RST(rst), .Q(sreg[1671]) );
  DFF \sreg_reg[1670]  ( .D(c[1672]), .CLK(clk), .RST(rst), .Q(sreg[1670]) );
  DFF \sreg_reg[1669]  ( .D(c[1671]), .CLK(clk), .RST(rst), .Q(sreg[1669]) );
  DFF \sreg_reg[1668]  ( .D(c[1670]), .CLK(clk), .RST(rst), .Q(sreg[1668]) );
  DFF \sreg_reg[1667]  ( .D(c[1669]), .CLK(clk), .RST(rst), .Q(sreg[1667]) );
  DFF \sreg_reg[1666]  ( .D(c[1668]), .CLK(clk), .RST(rst), .Q(sreg[1666]) );
  DFF \sreg_reg[1665]  ( .D(c[1667]), .CLK(clk), .RST(rst), .Q(sreg[1665]) );
  DFF \sreg_reg[1664]  ( .D(c[1666]), .CLK(clk), .RST(rst), .Q(sreg[1664]) );
  DFF \sreg_reg[1663]  ( .D(c[1665]), .CLK(clk), .RST(rst), .Q(sreg[1663]) );
  DFF \sreg_reg[1662]  ( .D(c[1664]), .CLK(clk), .RST(rst), .Q(sreg[1662]) );
  DFF \sreg_reg[1661]  ( .D(c[1663]), .CLK(clk), .RST(rst), .Q(sreg[1661]) );
  DFF \sreg_reg[1660]  ( .D(c[1662]), .CLK(clk), .RST(rst), .Q(sreg[1660]) );
  DFF \sreg_reg[1659]  ( .D(c[1661]), .CLK(clk), .RST(rst), .Q(sreg[1659]) );
  DFF \sreg_reg[1658]  ( .D(c[1660]), .CLK(clk), .RST(rst), .Q(sreg[1658]) );
  DFF \sreg_reg[1657]  ( .D(c[1659]), .CLK(clk), .RST(rst), .Q(sreg[1657]) );
  DFF \sreg_reg[1656]  ( .D(c[1658]), .CLK(clk), .RST(rst), .Q(sreg[1656]) );
  DFF \sreg_reg[1655]  ( .D(c[1657]), .CLK(clk), .RST(rst), .Q(sreg[1655]) );
  DFF \sreg_reg[1654]  ( .D(c[1656]), .CLK(clk), .RST(rst), .Q(sreg[1654]) );
  DFF \sreg_reg[1653]  ( .D(c[1655]), .CLK(clk), .RST(rst), .Q(sreg[1653]) );
  DFF \sreg_reg[1652]  ( .D(c[1654]), .CLK(clk), .RST(rst), .Q(sreg[1652]) );
  DFF \sreg_reg[1651]  ( .D(c[1653]), .CLK(clk), .RST(rst), .Q(sreg[1651]) );
  DFF \sreg_reg[1650]  ( .D(c[1652]), .CLK(clk), .RST(rst), .Q(sreg[1650]) );
  DFF \sreg_reg[1649]  ( .D(c[1651]), .CLK(clk), .RST(rst), .Q(sreg[1649]) );
  DFF \sreg_reg[1648]  ( .D(c[1650]), .CLK(clk), .RST(rst), .Q(sreg[1648]) );
  DFF \sreg_reg[1647]  ( .D(c[1649]), .CLK(clk), .RST(rst), .Q(sreg[1647]) );
  DFF \sreg_reg[1646]  ( .D(c[1648]), .CLK(clk), .RST(rst), .Q(sreg[1646]) );
  DFF \sreg_reg[1645]  ( .D(c[1647]), .CLK(clk), .RST(rst), .Q(sreg[1645]) );
  DFF \sreg_reg[1644]  ( .D(c[1646]), .CLK(clk), .RST(rst), .Q(sreg[1644]) );
  DFF \sreg_reg[1643]  ( .D(c[1645]), .CLK(clk), .RST(rst), .Q(sreg[1643]) );
  DFF \sreg_reg[1642]  ( .D(c[1644]), .CLK(clk), .RST(rst), .Q(sreg[1642]) );
  DFF \sreg_reg[1641]  ( .D(c[1643]), .CLK(clk), .RST(rst), .Q(sreg[1641]) );
  DFF \sreg_reg[1640]  ( .D(c[1642]), .CLK(clk), .RST(rst), .Q(sreg[1640]) );
  DFF \sreg_reg[1639]  ( .D(c[1641]), .CLK(clk), .RST(rst), .Q(sreg[1639]) );
  DFF \sreg_reg[1638]  ( .D(c[1640]), .CLK(clk), .RST(rst), .Q(sreg[1638]) );
  DFF \sreg_reg[1637]  ( .D(c[1639]), .CLK(clk), .RST(rst), .Q(sreg[1637]) );
  DFF \sreg_reg[1636]  ( .D(c[1638]), .CLK(clk), .RST(rst), .Q(sreg[1636]) );
  DFF \sreg_reg[1635]  ( .D(c[1637]), .CLK(clk), .RST(rst), .Q(sreg[1635]) );
  DFF \sreg_reg[1634]  ( .D(c[1636]), .CLK(clk), .RST(rst), .Q(sreg[1634]) );
  DFF \sreg_reg[1633]  ( .D(c[1635]), .CLK(clk), .RST(rst), .Q(sreg[1633]) );
  DFF \sreg_reg[1632]  ( .D(c[1634]), .CLK(clk), .RST(rst), .Q(sreg[1632]) );
  DFF \sreg_reg[1631]  ( .D(c[1633]), .CLK(clk), .RST(rst), .Q(sreg[1631]) );
  DFF \sreg_reg[1630]  ( .D(c[1632]), .CLK(clk), .RST(rst), .Q(sreg[1630]) );
  DFF \sreg_reg[1629]  ( .D(c[1631]), .CLK(clk), .RST(rst), .Q(sreg[1629]) );
  DFF \sreg_reg[1628]  ( .D(c[1630]), .CLK(clk), .RST(rst), .Q(sreg[1628]) );
  DFF \sreg_reg[1627]  ( .D(c[1629]), .CLK(clk), .RST(rst), .Q(sreg[1627]) );
  DFF \sreg_reg[1626]  ( .D(c[1628]), .CLK(clk), .RST(rst), .Q(sreg[1626]) );
  DFF \sreg_reg[1625]  ( .D(c[1627]), .CLK(clk), .RST(rst), .Q(sreg[1625]) );
  DFF \sreg_reg[1624]  ( .D(c[1626]), .CLK(clk), .RST(rst), .Q(sreg[1624]) );
  DFF \sreg_reg[1623]  ( .D(c[1625]), .CLK(clk), .RST(rst), .Q(sreg[1623]) );
  DFF \sreg_reg[1622]  ( .D(c[1624]), .CLK(clk), .RST(rst), .Q(sreg[1622]) );
  DFF \sreg_reg[1621]  ( .D(c[1623]), .CLK(clk), .RST(rst), .Q(sreg[1621]) );
  DFF \sreg_reg[1620]  ( .D(c[1622]), .CLK(clk), .RST(rst), .Q(sreg[1620]) );
  DFF \sreg_reg[1619]  ( .D(c[1621]), .CLK(clk), .RST(rst), .Q(sreg[1619]) );
  DFF \sreg_reg[1618]  ( .D(c[1620]), .CLK(clk), .RST(rst), .Q(sreg[1618]) );
  DFF \sreg_reg[1617]  ( .D(c[1619]), .CLK(clk), .RST(rst), .Q(sreg[1617]) );
  DFF \sreg_reg[1616]  ( .D(c[1618]), .CLK(clk), .RST(rst), .Q(sreg[1616]) );
  DFF \sreg_reg[1615]  ( .D(c[1617]), .CLK(clk), .RST(rst), .Q(sreg[1615]) );
  DFF \sreg_reg[1614]  ( .D(c[1616]), .CLK(clk), .RST(rst), .Q(sreg[1614]) );
  DFF \sreg_reg[1613]  ( .D(c[1615]), .CLK(clk), .RST(rst), .Q(sreg[1613]) );
  DFF \sreg_reg[1612]  ( .D(c[1614]), .CLK(clk), .RST(rst), .Q(sreg[1612]) );
  DFF \sreg_reg[1611]  ( .D(c[1613]), .CLK(clk), .RST(rst), .Q(sreg[1611]) );
  DFF \sreg_reg[1610]  ( .D(c[1612]), .CLK(clk), .RST(rst), .Q(sreg[1610]) );
  DFF \sreg_reg[1609]  ( .D(c[1611]), .CLK(clk), .RST(rst), .Q(sreg[1609]) );
  DFF \sreg_reg[1608]  ( .D(c[1610]), .CLK(clk), .RST(rst), .Q(sreg[1608]) );
  DFF \sreg_reg[1607]  ( .D(c[1609]), .CLK(clk), .RST(rst), .Q(sreg[1607]) );
  DFF \sreg_reg[1606]  ( .D(c[1608]), .CLK(clk), .RST(rst), .Q(sreg[1606]) );
  DFF \sreg_reg[1605]  ( .D(c[1607]), .CLK(clk), .RST(rst), .Q(sreg[1605]) );
  DFF \sreg_reg[1604]  ( .D(c[1606]), .CLK(clk), .RST(rst), .Q(sreg[1604]) );
  DFF \sreg_reg[1603]  ( .D(c[1605]), .CLK(clk), .RST(rst), .Q(sreg[1603]) );
  DFF \sreg_reg[1602]  ( .D(c[1604]), .CLK(clk), .RST(rst), .Q(sreg[1602]) );
  DFF \sreg_reg[1601]  ( .D(c[1603]), .CLK(clk), .RST(rst), .Q(sreg[1601]) );
  DFF \sreg_reg[1600]  ( .D(c[1602]), .CLK(clk), .RST(rst), .Q(sreg[1600]) );
  DFF \sreg_reg[1599]  ( .D(c[1601]), .CLK(clk), .RST(rst), .Q(sreg[1599]) );
  DFF \sreg_reg[1598]  ( .D(c[1600]), .CLK(clk), .RST(rst), .Q(sreg[1598]) );
  DFF \sreg_reg[1597]  ( .D(c[1599]), .CLK(clk), .RST(rst), .Q(sreg[1597]) );
  DFF \sreg_reg[1596]  ( .D(c[1598]), .CLK(clk), .RST(rst), .Q(sreg[1596]) );
  DFF \sreg_reg[1595]  ( .D(c[1597]), .CLK(clk), .RST(rst), .Q(sreg[1595]) );
  DFF \sreg_reg[1594]  ( .D(c[1596]), .CLK(clk), .RST(rst), .Q(sreg[1594]) );
  DFF \sreg_reg[1593]  ( .D(c[1595]), .CLK(clk), .RST(rst), .Q(sreg[1593]) );
  DFF \sreg_reg[1592]  ( .D(c[1594]), .CLK(clk), .RST(rst), .Q(sreg[1592]) );
  DFF \sreg_reg[1591]  ( .D(c[1593]), .CLK(clk), .RST(rst), .Q(sreg[1591]) );
  DFF \sreg_reg[1590]  ( .D(c[1592]), .CLK(clk), .RST(rst), .Q(sreg[1590]) );
  DFF \sreg_reg[1589]  ( .D(c[1591]), .CLK(clk), .RST(rst), .Q(sreg[1589]) );
  DFF \sreg_reg[1588]  ( .D(c[1590]), .CLK(clk), .RST(rst), .Q(sreg[1588]) );
  DFF \sreg_reg[1587]  ( .D(c[1589]), .CLK(clk), .RST(rst), .Q(sreg[1587]) );
  DFF \sreg_reg[1586]  ( .D(c[1588]), .CLK(clk), .RST(rst), .Q(sreg[1586]) );
  DFF \sreg_reg[1585]  ( .D(c[1587]), .CLK(clk), .RST(rst), .Q(sreg[1585]) );
  DFF \sreg_reg[1584]  ( .D(c[1586]), .CLK(clk), .RST(rst), .Q(sreg[1584]) );
  DFF \sreg_reg[1583]  ( .D(c[1585]), .CLK(clk), .RST(rst), .Q(sreg[1583]) );
  DFF \sreg_reg[1582]  ( .D(c[1584]), .CLK(clk), .RST(rst), .Q(sreg[1582]) );
  DFF \sreg_reg[1581]  ( .D(c[1583]), .CLK(clk), .RST(rst), .Q(sreg[1581]) );
  DFF \sreg_reg[1580]  ( .D(c[1582]), .CLK(clk), .RST(rst), .Q(sreg[1580]) );
  DFF \sreg_reg[1579]  ( .D(c[1581]), .CLK(clk), .RST(rst), .Q(sreg[1579]) );
  DFF \sreg_reg[1578]  ( .D(c[1580]), .CLK(clk), .RST(rst), .Q(sreg[1578]) );
  DFF \sreg_reg[1577]  ( .D(c[1579]), .CLK(clk), .RST(rst), .Q(sreg[1577]) );
  DFF \sreg_reg[1576]  ( .D(c[1578]), .CLK(clk), .RST(rst), .Q(sreg[1576]) );
  DFF \sreg_reg[1575]  ( .D(c[1577]), .CLK(clk), .RST(rst), .Q(sreg[1575]) );
  DFF \sreg_reg[1574]  ( .D(c[1576]), .CLK(clk), .RST(rst), .Q(sreg[1574]) );
  DFF \sreg_reg[1573]  ( .D(c[1575]), .CLK(clk), .RST(rst), .Q(sreg[1573]) );
  DFF \sreg_reg[1572]  ( .D(c[1574]), .CLK(clk), .RST(rst), .Q(sreg[1572]) );
  DFF \sreg_reg[1571]  ( .D(c[1573]), .CLK(clk), .RST(rst), .Q(sreg[1571]) );
  DFF \sreg_reg[1570]  ( .D(c[1572]), .CLK(clk), .RST(rst), .Q(sreg[1570]) );
  DFF \sreg_reg[1569]  ( .D(c[1571]), .CLK(clk), .RST(rst), .Q(sreg[1569]) );
  DFF \sreg_reg[1568]  ( .D(c[1570]), .CLK(clk), .RST(rst), .Q(sreg[1568]) );
  DFF \sreg_reg[1567]  ( .D(c[1569]), .CLK(clk), .RST(rst), .Q(sreg[1567]) );
  DFF \sreg_reg[1566]  ( .D(c[1568]), .CLK(clk), .RST(rst), .Q(sreg[1566]) );
  DFF \sreg_reg[1565]  ( .D(c[1567]), .CLK(clk), .RST(rst), .Q(sreg[1565]) );
  DFF \sreg_reg[1564]  ( .D(c[1566]), .CLK(clk), .RST(rst), .Q(sreg[1564]) );
  DFF \sreg_reg[1563]  ( .D(c[1565]), .CLK(clk), .RST(rst), .Q(sreg[1563]) );
  DFF \sreg_reg[1562]  ( .D(c[1564]), .CLK(clk), .RST(rst), .Q(sreg[1562]) );
  DFF \sreg_reg[1561]  ( .D(c[1563]), .CLK(clk), .RST(rst), .Q(sreg[1561]) );
  DFF \sreg_reg[1560]  ( .D(c[1562]), .CLK(clk), .RST(rst), .Q(sreg[1560]) );
  DFF \sreg_reg[1559]  ( .D(c[1561]), .CLK(clk), .RST(rst), .Q(sreg[1559]) );
  DFF \sreg_reg[1558]  ( .D(c[1560]), .CLK(clk), .RST(rst), .Q(sreg[1558]) );
  DFF \sreg_reg[1557]  ( .D(c[1559]), .CLK(clk), .RST(rst), .Q(sreg[1557]) );
  DFF \sreg_reg[1556]  ( .D(c[1558]), .CLK(clk), .RST(rst), .Q(sreg[1556]) );
  DFF \sreg_reg[1555]  ( .D(c[1557]), .CLK(clk), .RST(rst), .Q(sreg[1555]) );
  DFF \sreg_reg[1554]  ( .D(c[1556]), .CLK(clk), .RST(rst), .Q(sreg[1554]) );
  DFF \sreg_reg[1553]  ( .D(c[1555]), .CLK(clk), .RST(rst), .Q(sreg[1553]) );
  DFF \sreg_reg[1552]  ( .D(c[1554]), .CLK(clk), .RST(rst), .Q(sreg[1552]) );
  DFF \sreg_reg[1551]  ( .D(c[1553]), .CLK(clk), .RST(rst), .Q(sreg[1551]) );
  DFF \sreg_reg[1550]  ( .D(c[1552]), .CLK(clk), .RST(rst), .Q(sreg[1550]) );
  DFF \sreg_reg[1549]  ( .D(c[1551]), .CLK(clk), .RST(rst), .Q(sreg[1549]) );
  DFF \sreg_reg[1548]  ( .D(c[1550]), .CLK(clk), .RST(rst), .Q(sreg[1548]) );
  DFF \sreg_reg[1547]  ( .D(c[1549]), .CLK(clk), .RST(rst), .Q(sreg[1547]) );
  DFF \sreg_reg[1546]  ( .D(c[1548]), .CLK(clk), .RST(rst), .Q(sreg[1546]) );
  DFF \sreg_reg[1545]  ( .D(c[1547]), .CLK(clk), .RST(rst), .Q(sreg[1545]) );
  DFF \sreg_reg[1544]  ( .D(c[1546]), .CLK(clk), .RST(rst), .Q(sreg[1544]) );
  DFF \sreg_reg[1543]  ( .D(c[1545]), .CLK(clk), .RST(rst), .Q(sreg[1543]) );
  DFF \sreg_reg[1542]  ( .D(c[1544]), .CLK(clk), .RST(rst), .Q(sreg[1542]) );
  DFF \sreg_reg[1541]  ( .D(c[1543]), .CLK(clk), .RST(rst), .Q(sreg[1541]) );
  DFF \sreg_reg[1540]  ( .D(c[1542]), .CLK(clk), .RST(rst), .Q(sreg[1540]) );
  DFF \sreg_reg[1539]  ( .D(c[1541]), .CLK(clk), .RST(rst), .Q(sreg[1539]) );
  DFF \sreg_reg[1538]  ( .D(c[1540]), .CLK(clk), .RST(rst), .Q(sreg[1538]) );
  DFF \sreg_reg[1537]  ( .D(c[1539]), .CLK(clk), .RST(rst), .Q(sreg[1537]) );
  DFF \sreg_reg[1536]  ( .D(c[1538]), .CLK(clk), .RST(rst), .Q(sreg[1536]) );
  DFF \sreg_reg[1535]  ( .D(c[1537]), .CLK(clk), .RST(rst), .Q(sreg[1535]) );
  DFF \sreg_reg[1534]  ( .D(c[1536]), .CLK(clk), .RST(rst), .Q(sreg[1534]) );
  DFF \sreg_reg[1533]  ( .D(c[1535]), .CLK(clk), .RST(rst), .Q(sreg[1533]) );
  DFF \sreg_reg[1532]  ( .D(c[1534]), .CLK(clk), .RST(rst), .Q(sreg[1532]) );
  DFF \sreg_reg[1531]  ( .D(c[1533]), .CLK(clk), .RST(rst), .Q(sreg[1531]) );
  DFF \sreg_reg[1530]  ( .D(c[1532]), .CLK(clk), .RST(rst), .Q(sreg[1530]) );
  DFF \sreg_reg[1529]  ( .D(c[1531]), .CLK(clk), .RST(rst), .Q(sreg[1529]) );
  DFF \sreg_reg[1528]  ( .D(c[1530]), .CLK(clk), .RST(rst), .Q(sreg[1528]) );
  DFF \sreg_reg[1527]  ( .D(c[1529]), .CLK(clk), .RST(rst), .Q(sreg[1527]) );
  DFF \sreg_reg[1526]  ( .D(c[1528]), .CLK(clk), .RST(rst), .Q(sreg[1526]) );
  DFF \sreg_reg[1525]  ( .D(c[1527]), .CLK(clk), .RST(rst), .Q(sreg[1525]) );
  DFF \sreg_reg[1524]  ( .D(c[1526]), .CLK(clk), .RST(rst), .Q(sreg[1524]) );
  DFF \sreg_reg[1523]  ( .D(c[1525]), .CLK(clk), .RST(rst), .Q(sreg[1523]) );
  DFF \sreg_reg[1522]  ( .D(c[1524]), .CLK(clk), .RST(rst), .Q(sreg[1522]) );
  DFF \sreg_reg[1521]  ( .D(c[1523]), .CLK(clk), .RST(rst), .Q(sreg[1521]) );
  DFF \sreg_reg[1520]  ( .D(c[1522]), .CLK(clk), .RST(rst), .Q(sreg[1520]) );
  DFF \sreg_reg[1519]  ( .D(c[1521]), .CLK(clk), .RST(rst), .Q(sreg[1519]) );
  DFF \sreg_reg[1518]  ( .D(c[1520]), .CLK(clk), .RST(rst), .Q(sreg[1518]) );
  DFF \sreg_reg[1517]  ( .D(c[1519]), .CLK(clk), .RST(rst), .Q(sreg[1517]) );
  DFF \sreg_reg[1516]  ( .D(c[1518]), .CLK(clk), .RST(rst), .Q(sreg[1516]) );
  DFF \sreg_reg[1515]  ( .D(c[1517]), .CLK(clk), .RST(rst), .Q(sreg[1515]) );
  DFF \sreg_reg[1514]  ( .D(c[1516]), .CLK(clk), .RST(rst), .Q(sreg[1514]) );
  DFF \sreg_reg[1513]  ( .D(c[1515]), .CLK(clk), .RST(rst), .Q(sreg[1513]) );
  DFF \sreg_reg[1512]  ( .D(c[1514]), .CLK(clk), .RST(rst), .Q(sreg[1512]) );
  DFF \sreg_reg[1511]  ( .D(c[1513]), .CLK(clk), .RST(rst), .Q(sreg[1511]) );
  DFF \sreg_reg[1510]  ( .D(c[1512]), .CLK(clk), .RST(rst), .Q(sreg[1510]) );
  DFF \sreg_reg[1509]  ( .D(c[1511]), .CLK(clk), .RST(rst), .Q(sreg[1509]) );
  DFF \sreg_reg[1508]  ( .D(c[1510]), .CLK(clk), .RST(rst), .Q(sreg[1508]) );
  DFF \sreg_reg[1507]  ( .D(c[1509]), .CLK(clk), .RST(rst), .Q(sreg[1507]) );
  DFF \sreg_reg[1506]  ( .D(c[1508]), .CLK(clk), .RST(rst), .Q(sreg[1506]) );
  DFF \sreg_reg[1505]  ( .D(c[1507]), .CLK(clk), .RST(rst), .Q(sreg[1505]) );
  DFF \sreg_reg[1504]  ( .D(c[1506]), .CLK(clk), .RST(rst), .Q(sreg[1504]) );
  DFF \sreg_reg[1503]  ( .D(c[1505]), .CLK(clk), .RST(rst), .Q(sreg[1503]) );
  DFF \sreg_reg[1502]  ( .D(c[1504]), .CLK(clk), .RST(rst), .Q(sreg[1502]) );
  DFF \sreg_reg[1501]  ( .D(c[1503]), .CLK(clk), .RST(rst), .Q(sreg[1501]) );
  DFF \sreg_reg[1500]  ( .D(c[1502]), .CLK(clk), .RST(rst), .Q(sreg[1500]) );
  DFF \sreg_reg[1499]  ( .D(c[1501]), .CLK(clk), .RST(rst), .Q(sreg[1499]) );
  DFF \sreg_reg[1498]  ( .D(c[1500]), .CLK(clk), .RST(rst), .Q(sreg[1498]) );
  DFF \sreg_reg[1497]  ( .D(c[1499]), .CLK(clk), .RST(rst), .Q(sreg[1497]) );
  DFF \sreg_reg[1496]  ( .D(c[1498]), .CLK(clk), .RST(rst), .Q(sreg[1496]) );
  DFF \sreg_reg[1495]  ( .D(c[1497]), .CLK(clk), .RST(rst), .Q(sreg[1495]) );
  DFF \sreg_reg[1494]  ( .D(c[1496]), .CLK(clk), .RST(rst), .Q(sreg[1494]) );
  DFF \sreg_reg[1493]  ( .D(c[1495]), .CLK(clk), .RST(rst), .Q(sreg[1493]) );
  DFF \sreg_reg[1492]  ( .D(c[1494]), .CLK(clk), .RST(rst), .Q(sreg[1492]) );
  DFF \sreg_reg[1491]  ( .D(c[1493]), .CLK(clk), .RST(rst), .Q(sreg[1491]) );
  DFF \sreg_reg[1490]  ( .D(c[1492]), .CLK(clk), .RST(rst), .Q(sreg[1490]) );
  DFF \sreg_reg[1489]  ( .D(c[1491]), .CLK(clk), .RST(rst), .Q(sreg[1489]) );
  DFF \sreg_reg[1488]  ( .D(c[1490]), .CLK(clk), .RST(rst), .Q(sreg[1488]) );
  DFF \sreg_reg[1487]  ( .D(c[1489]), .CLK(clk), .RST(rst), .Q(sreg[1487]) );
  DFF \sreg_reg[1486]  ( .D(c[1488]), .CLK(clk), .RST(rst), .Q(sreg[1486]) );
  DFF \sreg_reg[1485]  ( .D(c[1487]), .CLK(clk), .RST(rst), .Q(sreg[1485]) );
  DFF \sreg_reg[1484]  ( .D(c[1486]), .CLK(clk), .RST(rst), .Q(sreg[1484]) );
  DFF \sreg_reg[1483]  ( .D(c[1485]), .CLK(clk), .RST(rst), .Q(sreg[1483]) );
  DFF \sreg_reg[1482]  ( .D(c[1484]), .CLK(clk), .RST(rst), .Q(sreg[1482]) );
  DFF \sreg_reg[1481]  ( .D(c[1483]), .CLK(clk), .RST(rst), .Q(sreg[1481]) );
  DFF \sreg_reg[1480]  ( .D(c[1482]), .CLK(clk), .RST(rst), .Q(sreg[1480]) );
  DFF \sreg_reg[1479]  ( .D(c[1481]), .CLK(clk), .RST(rst), .Q(sreg[1479]) );
  DFF \sreg_reg[1478]  ( .D(c[1480]), .CLK(clk), .RST(rst), .Q(sreg[1478]) );
  DFF \sreg_reg[1477]  ( .D(c[1479]), .CLK(clk), .RST(rst), .Q(sreg[1477]) );
  DFF \sreg_reg[1476]  ( .D(c[1478]), .CLK(clk), .RST(rst), .Q(sreg[1476]) );
  DFF \sreg_reg[1475]  ( .D(c[1477]), .CLK(clk), .RST(rst), .Q(sreg[1475]) );
  DFF \sreg_reg[1474]  ( .D(c[1476]), .CLK(clk), .RST(rst), .Q(sreg[1474]) );
  DFF \sreg_reg[1473]  ( .D(c[1475]), .CLK(clk), .RST(rst), .Q(sreg[1473]) );
  DFF \sreg_reg[1472]  ( .D(c[1474]), .CLK(clk), .RST(rst), .Q(sreg[1472]) );
  DFF \sreg_reg[1471]  ( .D(c[1473]), .CLK(clk), .RST(rst), .Q(sreg[1471]) );
  DFF \sreg_reg[1470]  ( .D(c[1472]), .CLK(clk), .RST(rst), .Q(sreg[1470]) );
  DFF \sreg_reg[1469]  ( .D(c[1471]), .CLK(clk), .RST(rst), .Q(sreg[1469]) );
  DFF \sreg_reg[1468]  ( .D(c[1470]), .CLK(clk), .RST(rst), .Q(sreg[1468]) );
  DFF \sreg_reg[1467]  ( .D(c[1469]), .CLK(clk), .RST(rst), .Q(sreg[1467]) );
  DFF \sreg_reg[1466]  ( .D(c[1468]), .CLK(clk), .RST(rst), .Q(sreg[1466]) );
  DFF \sreg_reg[1465]  ( .D(c[1467]), .CLK(clk), .RST(rst), .Q(sreg[1465]) );
  DFF \sreg_reg[1464]  ( .D(c[1466]), .CLK(clk), .RST(rst), .Q(sreg[1464]) );
  DFF \sreg_reg[1463]  ( .D(c[1465]), .CLK(clk), .RST(rst), .Q(sreg[1463]) );
  DFF \sreg_reg[1462]  ( .D(c[1464]), .CLK(clk), .RST(rst), .Q(sreg[1462]) );
  DFF \sreg_reg[1461]  ( .D(c[1463]), .CLK(clk), .RST(rst), .Q(sreg[1461]) );
  DFF \sreg_reg[1460]  ( .D(c[1462]), .CLK(clk), .RST(rst), .Q(sreg[1460]) );
  DFF \sreg_reg[1459]  ( .D(c[1461]), .CLK(clk), .RST(rst), .Q(sreg[1459]) );
  DFF \sreg_reg[1458]  ( .D(c[1460]), .CLK(clk), .RST(rst), .Q(sreg[1458]) );
  DFF \sreg_reg[1457]  ( .D(c[1459]), .CLK(clk), .RST(rst), .Q(sreg[1457]) );
  DFF \sreg_reg[1456]  ( .D(c[1458]), .CLK(clk), .RST(rst), .Q(sreg[1456]) );
  DFF \sreg_reg[1455]  ( .D(c[1457]), .CLK(clk), .RST(rst), .Q(sreg[1455]) );
  DFF \sreg_reg[1454]  ( .D(c[1456]), .CLK(clk), .RST(rst), .Q(sreg[1454]) );
  DFF \sreg_reg[1453]  ( .D(c[1455]), .CLK(clk), .RST(rst), .Q(sreg[1453]) );
  DFF \sreg_reg[1452]  ( .D(c[1454]), .CLK(clk), .RST(rst), .Q(sreg[1452]) );
  DFF \sreg_reg[1451]  ( .D(c[1453]), .CLK(clk), .RST(rst), .Q(sreg[1451]) );
  DFF \sreg_reg[1450]  ( .D(c[1452]), .CLK(clk), .RST(rst), .Q(sreg[1450]) );
  DFF \sreg_reg[1449]  ( .D(c[1451]), .CLK(clk), .RST(rst), .Q(sreg[1449]) );
  DFF \sreg_reg[1448]  ( .D(c[1450]), .CLK(clk), .RST(rst), .Q(sreg[1448]) );
  DFF \sreg_reg[1447]  ( .D(c[1449]), .CLK(clk), .RST(rst), .Q(sreg[1447]) );
  DFF \sreg_reg[1446]  ( .D(c[1448]), .CLK(clk), .RST(rst), .Q(sreg[1446]) );
  DFF \sreg_reg[1445]  ( .D(c[1447]), .CLK(clk), .RST(rst), .Q(sreg[1445]) );
  DFF \sreg_reg[1444]  ( .D(c[1446]), .CLK(clk), .RST(rst), .Q(sreg[1444]) );
  DFF \sreg_reg[1443]  ( .D(c[1445]), .CLK(clk), .RST(rst), .Q(sreg[1443]) );
  DFF \sreg_reg[1442]  ( .D(c[1444]), .CLK(clk), .RST(rst), .Q(sreg[1442]) );
  DFF \sreg_reg[1441]  ( .D(c[1443]), .CLK(clk), .RST(rst), .Q(sreg[1441]) );
  DFF \sreg_reg[1440]  ( .D(c[1442]), .CLK(clk), .RST(rst), .Q(sreg[1440]) );
  DFF \sreg_reg[1439]  ( .D(c[1441]), .CLK(clk), .RST(rst), .Q(sreg[1439]) );
  DFF \sreg_reg[1438]  ( .D(c[1440]), .CLK(clk), .RST(rst), .Q(sreg[1438]) );
  DFF \sreg_reg[1437]  ( .D(c[1439]), .CLK(clk), .RST(rst), .Q(sreg[1437]) );
  DFF \sreg_reg[1436]  ( .D(c[1438]), .CLK(clk), .RST(rst), .Q(sreg[1436]) );
  DFF \sreg_reg[1435]  ( .D(c[1437]), .CLK(clk), .RST(rst), .Q(sreg[1435]) );
  DFF \sreg_reg[1434]  ( .D(c[1436]), .CLK(clk), .RST(rst), .Q(sreg[1434]) );
  DFF \sreg_reg[1433]  ( .D(c[1435]), .CLK(clk), .RST(rst), .Q(sreg[1433]) );
  DFF \sreg_reg[1432]  ( .D(c[1434]), .CLK(clk), .RST(rst), .Q(sreg[1432]) );
  DFF \sreg_reg[1431]  ( .D(c[1433]), .CLK(clk), .RST(rst), .Q(sreg[1431]) );
  DFF \sreg_reg[1430]  ( .D(c[1432]), .CLK(clk), .RST(rst), .Q(sreg[1430]) );
  DFF \sreg_reg[1429]  ( .D(c[1431]), .CLK(clk), .RST(rst), .Q(sreg[1429]) );
  DFF \sreg_reg[1428]  ( .D(c[1430]), .CLK(clk), .RST(rst), .Q(sreg[1428]) );
  DFF \sreg_reg[1427]  ( .D(c[1429]), .CLK(clk), .RST(rst), .Q(sreg[1427]) );
  DFF \sreg_reg[1426]  ( .D(c[1428]), .CLK(clk), .RST(rst), .Q(sreg[1426]) );
  DFF \sreg_reg[1425]  ( .D(c[1427]), .CLK(clk), .RST(rst), .Q(sreg[1425]) );
  DFF \sreg_reg[1424]  ( .D(c[1426]), .CLK(clk), .RST(rst), .Q(sreg[1424]) );
  DFF \sreg_reg[1423]  ( .D(c[1425]), .CLK(clk), .RST(rst), .Q(sreg[1423]) );
  DFF \sreg_reg[1422]  ( .D(c[1424]), .CLK(clk), .RST(rst), .Q(sreg[1422]) );
  DFF \sreg_reg[1421]  ( .D(c[1423]), .CLK(clk), .RST(rst), .Q(sreg[1421]) );
  DFF \sreg_reg[1420]  ( .D(c[1422]), .CLK(clk), .RST(rst), .Q(sreg[1420]) );
  DFF \sreg_reg[1419]  ( .D(c[1421]), .CLK(clk), .RST(rst), .Q(sreg[1419]) );
  DFF \sreg_reg[1418]  ( .D(c[1420]), .CLK(clk), .RST(rst), .Q(sreg[1418]) );
  DFF \sreg_reg[1417]  ( .D(c[1419]), .CLK(clk), .RST(rst), .Q(sreg[1417]) );
  DFF \sreg_reg[1416]  ( .D(c[1418]), .CLK(clk), .RST(rst), .Q(sreg[1416]) );
  DFF \sreg_reg[1415]  ( .D(c[1417]), .CLK(clk), .RST(rst), .Q(sreg[1415]) );
  DFF \sreg_reg[1414]  ( .D(c[1416]), .CLK(clk), .RST(rst), .Q(sreg[1414]) );
  DFF \sreg_reg[1413]  ( .D(c[1415]), .CLK(clk), .RST(rst), .Q(sreg[1413]) );
  DFF \sreg_reg[1412]  ( .D(c[1414]), .CLK(clk), .RST(rst), .Q(sreg[1412]) );
  DFF \sreg_reg[1411]  ( .D(c[1413]), .CLK(clk), .RST(rst), .Q(sreg[1411]) );
  DFF \sreg_reg[1410]  ( .D(c[1412]), .CLK(clk), .RST(rst), .Q(sreg[1410]) );
  DFF \sreg_reg[1409]  ( .D(c[1411]), .CLK(clk), .RST(rst), .Q(sreg[1409]) );
  DFF \sreg_reg[1408]  ( .D(c[1410]), .CLK(clk), .RST(rst), .Q(sreg[1408]) );
  DFF \sreg_reg[1407]  ( .D(c[1409]), .CLK(clk), .RST(rst), .Q(sreg[1407]) );
  DFF \sreg_reg[1406]  ( .D(c[1408]), .CLK(clk), .RST(rst), .Q(sreg[1406]) );
  DFF \sreg_reg[1405]  ( .D(c[1407]), .CLK(clk), .RST(rst), .Q(sreg[1405]) );
  DFF \sreg_reg[1404]  ( .D(c[1406]), .CLK(clk), .RST(rst), .Q(sreg[1404]) );
  DFF \sreg_reg[1403]  ( .D(c[1405]), .CLK(clk), .RST(rst), .Q(sreg[1403]) );
  DFF \sreg_reg[1402]  ( .D(c[1404]), .CLK(clk), .RST(rst), .Q(sreg[1402]) );
  DFF \sreg_reg[1401]  ( .D(c[1403]), .CLK(clk), .RST(rst), .Q(sreg[1401]) );
  DFF \sreg_reg[1400]  ( .D(c[1402]), .CLK(clk), .RST(rst), .Q(sreg[1400]) );
  DFF \sreg_reg[1399]  ( .D(c[1401]), .CLK(clk), .RST(rst), .Q(sreg[1399]) );
  DFF \sreg_reg[1398]  ( .D(c[1400]), .CLK(clk), .RST(rst), .Q(sreg[1398]) );
  DFF \sreg_reg[1397]  ( .D(c[1399]), .CLK(clk), .RST(rst), .Q(sreg[1397]) );
  DFF \sreg_reg[1396]  ( .D(c[1398]), .CLK(clk), .RST(rst), .Q(sreg[1396]) );
  DFF \sreg_reg[1395]  ( .D(c[1397]), .CLK(clk), .RST(rst), .Q(sreg[1395]) );
  DFF \sreg_reg[1394]  ( .D(c[1396]), .CLK(clk), .RST(rst), .Q(sreg[1394]) );
  DFF \sreg_reg[1393]  ( .D(c[1395]), .CLK(clk), .RST(rst), .Q(sreg[1393]) );
  DFF \sreg_reg[1392]  ( .D(c[1394]), .CLK(clk), .RST(rst), .Q(sreg[1392]) );
  DFF \sreg_reg[1391]  ( .D(c[1393]), .CLK(clk), .RST(rst), .Q(sreg[1391]) );
  DFF \sreg_reg[1390]  ( .D(c[1392]), .CLK(clk), .RST(rst), .Q(sreg[1390]) );
  DFF \sreg_reg[1389]  ( .D(c[1391]), .CLK(clk), .RST(rst), .Q(sreg[1389]) );
  DFF \sreg_reg[1388]  ( .D(c[1390]), .CLK(clk), .RST(rst), .Q(sreg[1388]) );
  DFF \sreg_reg[1387]  ( .D(c[1389]), .CLK(clk), .RST(rst), .Q(sreg[1387]) );
  DFF \sreg_reg[1386]  ( .D(c[1388]), .CLK(clk), .RST(rst), .Q(sreg[1386]) );
  DFF \sreg_reg[1385]  ( .D(c[1387]), .CLK(clk), .RST(rst), .Q(sreg[1385]) );
  DFF \sreg_reg[1384]  ( .D(c[1386]), .CLK(clk), .RST(rst), .Q(sreg[1384]) );
  DFF \sreg_reg[1383]  ( .D(c[1385]), .CLK(clk), .RST(rst), .Q(sreg[1383]) );
  DFF \sreg_reg[1382]  ( .D(c[1384]), .CLK(clk), .RST(rst), .Q(sreg[1382]) );
  DFF \sreg_reg[1381]  ( .D(c[1383]), .CLK(clk), .RST(rst), .Q(sreg[1381]) );
  DFF \sreg_reg[1380]  ( .D(c[1382]), .CLK(clk), .RST(rst), .Q(sreg[1380]) );
  DFF \sreg_reg[1379]  ( .D(c[1381]), .CLK(clk), .RST(rst), .Q(sreg[1379]) );
  DFF \sreg_reg[1378]  ( .D(c[1380]), .CLK(clk), .RST(rst), .Q(sreg[1378]) );
  DFF \sreg_reg[1377]  ( .D(c[1379]), .CLK(clk), .RST(rst), .Q(sreg[1377]) );
  DFF \sreg_reg[1376]  ( .D(c[1378]), .CLK(clk), .RST(rst), .Q(sreg[1376]) );
  DFF \sreg_reg[1375]  ( .D(c[1377]), .CLK(clk), .RST(rst), .Q(sreg[1375]) );
  DFF \sreg_reg[1374]  ( .D(c[1376]), .CLK(clk), .RST(rst), .Q(sreg[1374]) );
  DFF \sreg_reg[1373]  ( .D(c[1375]), .CLK(clk), .RST(rst), .Q(sreg[1373]) );
  DFF \sreg_reg[1372]  ( .D(c[1374]), .CLK(clk), .RST(rst), .Q(sreg[1372]) );
  DFF \sreg_reg[1371]  ( .D(c[1373]), .CLK(clk), .RST(rst), .Q(sreg[1371]) );
  DFF \sreg_reg[1370]  ( .D(c[1372]), .CLK(clk), .RST(rst), .Q(sreg[1370]) );
  DFF \sreg_reg[1369]  ( .D(c[1371]), .CLK(clk), .RST(rst), .Q(sreg[1369]) );
  DFF \sreg_reg[1368]  ( .D(c[1370]), .CLK(clk), .RST(rst), .Q(sreg[1368]) );
  DFF \sreg_reg[1367]  ( .D(c[1369]), .CLK(clk), .RST(rst), .Q(sreg[1367]) );
  DFF \sreg_reg[1366]  ( .D(c[1368]), .CLK(clk), .RST(rst), .Q(sreg[1366]) );
  DFF \sreg_reg[1365]  ( .D(c[1367]), .CLK(clk), .RST(rst), .Q(sreg[1365]) );
  DFF \sreg_reg[1364]  ( .D(c[1366]), .CLK(clk), .RST(rst), .Q(sreg[1364]) );
  DFF \sreg_reg[1363]  ( .D(c[1365]), .CLK(clk), .RST(rst), .Q(sreg[1363]) );
  DFF \sreg_reg[1362]  ( .D(c[1364]), .CLK(clk), .RST(rst), .Q(sreg[1362]) );
  DFF \sreg_reg[1361]  ( .D(c[1363]), .CLK(clk), .RST(rst), .Q(sreg[1361]) );
  DFF \sreg_reg[1360]  ( .D(c[1362]), .CLK(clk), .RST(rst), .Q(sreg[1360]) );
  DFF \sreg_reg[1359]  ( .D(c[1361]), .CLK(clk), .RST(rst), .Q(sreg[1359]) );
  DFF \sreg_reg[1358]  ( .D(c[1360]), .CLK(clk), .RST(rst), .Q(sreg[1358]) );
  DFF \sreg_reg[1357]  ( .D(c[1359]), .CLK(clk), .RST(rst), .Q(sreg[1357]) );
  DFF \sreg_reg[1356]  ( .D(c[1358]), .CLK(clk), .RST(rst), .Q(sreg[1356]) );
  DFF \sreg_reg[1355]  ( .D(c[1357]), .CLK(clk), .RST(rst), .Q(sreg[1355]) );
  DFF \sreg_reg[1354]  ( .D(c[1356]), .CLK(clk), .RST(rst), .Q(sreg[1354]) );
  DFF \sreg_reg[1353]  ( .D(c[1355]), .CLK(clk), .RST(rst), .Q(sreg[1353]) );
  DFF \sreg_reg[1352]  ( .D(c[1354]), .CLK(clk), .RST(rst), .Q(sreg[1352]) );
  DFF \sreg_reg[1351]  ( .D(c[1353]), .CLK(clk), .RST(rst), .Q(sreg[1351]) );
  DFF \sreg_reg[1350]  ( .D(c[1352]), .CLK(clk), .RST(rst), .Q(sreg[1350]) );
  DFF \sreg_reg[1349]  ( .D(c[1351]), .CLK(clk), .RST(rst), .Q(sreg[1349]) );
  DFF \sreg_reg[1348]  ( .D(c[1350]), .CLK(clk), .RST(rst), .Q(sreg[1348]) );
  DFF \sreg_reg[1347]  ( .D(c[1349]), .CLK(clk), .RST(rst), .Q(sreg[1347]) );
  DFF \sreg_reg[1346]  ( .D(c[1348]), .CLK(clk), .RST(rst), .Q(sreg[1346]) );
  DFF \sreg_reg[1345]  ( .D(c[1347]), .CLK(clk), .RST(rst), .Q(sreg[1345]) );
  DFF \sreg_reg[1344]  ( .D(c[1346]), .CLK(clk), .RST(rst), .Q(sreg[1344]) );
  DFF \sreg_reg[1343]  ( .D(c[1345]), .CLK(clk), .RST(rst), .Q(sreg[1343]) );
  DFF \sreg_reg[1342]  ( .D(c[1344]), .CLK(clk), .RST(rst), .Q(sreg[1342]) );
  DFF \sreg_reg[1341]  ( .D(c[1343]), .CLK(clk), .RST(rst), .Q(sreg[1341]) );
  DFF \sreg_reg[1340]  ( .D(c[1342]), .CLK(clk), .RST(rst), .Q(sreg[1340]) );
  DFF \sreg_reg[1339]  ( .D(c[1341]), .CLK(clk), .RST(rst), .Q(sreg[1339]) );
  DFF \sreg_reg[1338]  ( .D(c[1340]), .CLK(clk), .RST(rst), .Q(sreg[1338]) );
  DFF \sreg_reg[1337]  ( .D(c[1339]), .CLK(clk), .RST(rst), .Q(sreg[1337]) );
  DFF \sreg_reg[1336]  ( .D(c[1338]), .CLK(clk), .RST(rst), .Q(sreg[1336]) );
  DFF \sreg_reg[1335]  ( .D(c[1337]), .CLK(clk), .RST(rst), .Q(sreg[1335]) );
  DFF \sreg_reg[1334]  ( .D(c[1336]), .CLK(clk), .RST(rst), .Q(sreg[1334]) );
  DFF \sreg_reg[1333]  ( .D(c[1335]), .CLK(clk), .RST(rst), .Q(sreg[1333]) );
  DFF \sreg_reg[1332]  ( .D(c[1334]), .CLK(clk), .RST(rst), .Q(sreg[1332]) );
  DFF \sreg_reg[1331]  ( .D(c[1333]), .CLK(clk), .RST(rst), .Q(sreg[1331]) );
  DFF \sreg_reg[1330]  ( .D(c[1332]), .CLK(clk), .RST(rst), .Q(sreg[1330]) );
  DFF \sreg_reg[1329]  ( .D(c[1331]), .CLK(clk), .RST(rst), .Q(sreg[1329]) );
  DFF \sreg_reg[1328]  ( .D(c[1330]), .CLK(clk), .RST(rst), .Q(sreg[1328]) );
  DFF \sreg_reg[1327]  ( .D(c[1329]), .CLK(clk), .RST(rst), .Q(sreg[1327]) );
  DFF \sreg_reg[1326]  ( .D(c[1328]), .CLK(clk), .RST(rst), .Q(sreg[1326]) );
  DFF \sreg_reg[1325]  ( .D(c[1327]), .CLK(clk), .RST(rst), .Q(sreg[1325]) );
  DFF \sreg_reg[1324]  ( .D(c[1326]), .CLK(clk), .RST(rst), .Q(sreg[1324]) );
  DFF \sreg_reg[1323]  ( .D(c[1325]), .CLK(clk), .RST(rst), .Q(sreg[1323]) );
  DFF \sreg_reg[1322]  ( .D(c[1324]), .CLK(clk), .RST(rst), .Q(sreg[1322]) );
  DFF \sreg_reg[1321]  ( .D(c[1323]), .CLK(clk), .RST(rst), .Q(sreg[1321]) );
  DFF \sreg_reg[1320]  ( .D(c[1322]), .CLK(clk), .RST(rst), .Q(sreg[1320]) );
  DFF \sreg_reg[1319]  ( .D(c[1321]), .CLK(clk), .RST(rst), .Q(sreg[1319]) );
  DFF \sreg_reg[1318]  ( .D(c[1320]), .CLK(clk), .RST(rst), .Q(sreg[1318]) );
  DFF \sreg_reg[1317]  ( .D(c[1319]), .CLK(clk), .RST(rst), .Q(sreg[1317]) );
  DFF \sreg_reg[1316]  ( .D(c[1318]), .CLK(clk), .RST(rst), .Q(sreg[1316]) );
  DFF \sreg_reg[1315]  ( .D(c[1317]), .CLK(clk), .RST(rst), .Q(sreg[1315]) );
  DFF \sreg_reg[1314]  ( .D(c[1316]), .CLK(clk), .RST(rst), .Q(sreg[1314]) );
  DFF \sreg_reg[1313]  ( .D(c[1315]), .CLK(clk), .RST(rst), .Q(sreg[1313]) );
  DFF \sreg_reg[1312]  ( .D(c[1314]), .CLK(clk), .RST(rst), .Q(sreg[1312]) );
  DFF \sreg_reg[1311]  ( .D(c[1313]), .CLK(clk), .RST(rst), .Q(sreg[1311]) );
  DFF \sreg_reg[1310]  ( .D(c[1312]), .CLK(clk), .RST(rst), .Q(sreg[1310]) );
  DFF \sreg_reg[1309]  ( .D(c[1311]), .CLK(clk), .RST(rst), .Q(sreg[1309]) );
  DFF \sreg_reg[1308]  ( .D(c[1310]), .CLK(clk), .RST(rst), .Q(sreg[1308]) );
  DFF \sreg_reg[1307]  ( .D(c[1309]), .CLK(clk), .RST(rst), .Q(sreg[1307]) );
  DFF \sreg_reg[1306]  ( .D(c[1308]), .CLK(clk), .RST(rst), .Q(sreg[1306]) );
  DFF \sreg_reg[1305]  ( .D(c[1307]), .CLK(clk), .RST(rst), .Q(sreg[1305]) );
  DFF \sreg_reg[1304]  ( .D(c[1306]), .CLK(clk), .RST(rst), .Q(sreg[1304]) );
  DFF \sreg_reg[1303]  ( .D(c[1305]), .CLK(clk), .RST(rst), .Q(sreg[1303]) );
  DFF \sreg_reg[1302]  ( .D(c[1304]), .CLK(clk), .RST(rst), .Q(sreg[1302]) );
  DFF \sreg_reg[1301]  ( .D(c[1303]), .CLK(clk), .RST(rst), .Q(sreg[1301]) );
  DFF \sreg_reg[1300]  ( .D(c[1302]), .CLK(clk), .RST(rst), .Q(sreg[1300]) );
  DFF \sreg_reg[1299]  ( .D(c[1301]), .CLK(clk), .RST(rst), .Q(sreg[1299]) );
  DFF \sreg_reg[1298]  ( .D(c[1300]), .CLK(clk), .RST(rst), .Q(sreg[1298]) );
  DFF \sreg_reg[1297]  ( .D(c[1299]), .CLK(clk), .RST(rst), .Q(sreg[1297]) );
  DFF \sreg_reg[1296]  ( .D(c[1298]), .CLK(clk), .RST(rst), .Q(sreg[1296]) );
  DFF \sreg_reg[1295]  ( .D(c[1297]), .CLK(clk), .RST(rst), .Q(sreg[1295]) );
  DFF \sreg_reg[1294]  ( .D(c[1296]), .CLK(clk), .RST(rst), .Q(sreg[1294]) );
  DFF \sreg_reg[1293]  ( .D(c[1295]), .CLK(clk), .RST(rst), .Q(sreg[1293]) );
  DFF \sreg_reg[1292]  ( .D(c[1294]), .CLK(clk), .RST(rst), .Q(sreg[1292]) );
  DFF \sreg_reg[1291]  ( .D(c[1293]), .CLK(clk), .RST(rst), .Q(sreg[1291]) );
  DFF \sreg_reg[1290]  ( .D(c[1292]), .CLK(clk), .RST(rst), .Q(sreg[1290]) );
  DFF \sreg_reg[1289]  ( .D(c[1291]), .CLK(clk), .RST(rst), .Q(sreg[1289]) );
  DFF \sreg_reg[1288]  ( .D(c[1290]), .CLK(clk), .RST(rst), .Q(sreg[1288]) );
  DFF \sreg_reg[1287]  ( .D(c[1289]), .CLK(clk), .RST(rst), .Q(sreg[1287]) );
  DFF \sreg_reg[1286]  ( .D(c[1288]), .CLK(clk), .RST(rst), .Q(sreg[1286]) );
  DFF \sreg_reg[1285]  ( .D(c[1287]), .CLK(clk), .RST(rst), .Q(sreg[1285]) );
  DFF \sreg_reg[1284]  ( .D(c[1286]), .CLK(clk), .RST(rst), .Q(sreg[1284]) );
  DFF \sreg_reg[1283]  ( .D(c[1285]), .CLK(clk), .RST(rst), .Q(sreg[1283]) );
  DFF \sreg_reg[1282]  ( .D(c[1284]), .CLK(clk), .RST(rst), .Q(sreg[1282]) );
  DFF \sreg_reg[1281]  ( .D(c[1283]), .CLK(clk), .RST(rst), .Q(sreg[1281]) );
  DFF \sreg_reg[1280]  ( .D(c[1282]), .CLK(clk), .RST(rst), .Q(sreg[1280]) );
  DFF \sreg_reg[1279]  ( .D(c[1281]), .CLK(clk), .RST(rst), .Q(sreg[1279]) );
  DFF \sreg_reg[1278]  ( .D(c[1280]), .CLK(clk), .RST(rst), .Q(sreg[1278]) );
  DFF \sreg_reg[1277]  ( .D(c[1279]), .CLK(clk), .RST(rst), .Q(sreg[1277]) );
  DFF \sreg_reg[1276]  ( .D(c[1278]), .CLK(clk), .RST(rst), .Q(sreg[1276]) );
  DFF \sreg_reg[1275]  ( .D(c[1277]), .CLK(clk), .RST(rst), .Q(sreg[1275]) );
  DFF \sreg_reg[1274]  ( .D(c[1276]), .CLK(clk), .RST(rst), .Q(sreg[1274]) );
  DFF \sreg_reg[1273]  ( .D(c[1275]), .CLK(clk), .RST(rst), .Q(sreg[1273]) );
  DFF \sreg_reg[1272]  ( .D(c[1274]), .CLK(clk), .RST(rst), .Q(sreg[1272]) );
  DFF \sreg_reg[1271]  ( .D(c[1273]), .CLK(clk), .RST(rst), .Q(sreg[1271]) );
  DFF \sreg_reg[1270]  ( .D(c[1272]), .CLK(clk), .RST(rst), .Q(sreg[1270]) );
  DFF \sreg_reg[1269]  ( .D(c[1271]), .CLK(clk), .RST(rst), .Q(sreg[1269]) );
  DFF \sreg_reg[1268]  ( .D(c[1270]), .CLK(clk), .RST(rst), .Q(sreg[1268]) );
  DFF \sreg_reg[1267]  ( .D(c[1269]), .CLK(clk), .RST(rst), .Q(sreg[1267]) );
  DFF \sreg_reg[1266]  ( .D(c[1268]), .CLK(clk), .RST(rst), .Q(sreg[1266]) );
  DFF \sreg_reg[1265]  ( .D(c[1267]), .CLK(clk), .RST(rst), .Q(sreg[1265]) );
  DFF \sreg_reg[1264]  ( .D(c[1266]), .CLK(clk), .RST(rst), .Q(sreg[1264]) );
  DFF \sreg_reg[1263]  ( .D(c[1265]), .CLK(clk), .RST(rst), .Q(sreg[1263]) );
  DFF \sreg_reg[1262]  ( .D(c[1264]), .CLK(clk), .RST(rst), .Q(sreg[1262]) );
  DFF \sreg_reg[1261]  ( .D(c[1263]), .CLK(clk), .RST(rst), .Q(sreg[1261]) );
  DFF \sreg_reg[1260]  ( .D(c[1262]), .CLK(clk), .RST(rst), .Q(sreg[1260]) );
  DFF \sreg_reg[1259]  ( .D(c[1261]), .CLK(clk), .RST(rst), .Q(sreg[1259]) );
  DFF \sreg_reg[1258]  ( .D(c[1260]), .CLK(clk), .RST(rst), .Q(sreg[1258]) );
  DFF \sreg_reg[1257]  ( .D(c[1259]), .CLK(clk), .RST(rst), .Q(sreg[1257]) );
  DFF \sreg_reg[1256]  ( .D(c[1258]), .CLK(clk), .RST(rst), .Q(sreg[1256]) );
  DFF \sreg_reg[1255]  ( .D(c[1257]), .CLK(clk), .RST(rst), .Q(sreg[1255]) );
  DFF \sreg_reg[1254]  ( .D(c[1256]), .CLK(clk), .RST(rst), .Q(sreg[1254]) );
  DFF \sreg_reg[1253]  ( .D(c[1255]), .CLK(clk), .RST(rst), .Q(sreg[1253]) );
  DFF \sreg_reg[1252]  ( .D(c[1254]), .CLK(clk), .RST(rst), .Q(sreg[1252]) );
  DFF \sreg_reg[1251]  ( .D(c[1253]), .CLK(clk), .RST(rst), .Q(sreg[1251]) );
  DFF \sreg_reg[1250]  ( .D(c[1252]), .CLK(clk), .RST(rst), .Q(sreg[1250]) );
  DFF \sreg_reg[1249]  ( .D(c[1251]), .CLK(clk), .RST(rst), .Q(sreg[1249]) );
  DFF \sreg_reg[1248]  ( .D(c[1250]), .CLK(clk), .RST(rst), .Q(sreg[1248]) );
  DFF \sreg_reg[1247]  ( .D(c[1249]), .CLK(clk), .RST(rst), .Q(sreg[1247]) );
  DFF \sreg_reg[1246]  ( .D(c[1248]), .CLK(clk), .RST(rst), .Q(sreg[1246]) );
  DFF \sreg_reg[1245]  ( .D(c[1247]), .CLK(clk), .RST(rst), .Q(sreg[1245]) );
  DFF \sreg_reg[1244]  ( .D(c[1246]), .CLK(clk), .RST(rst), .Q(sreg[1244]) );
  DFF \sreg_reg[1243]  ( .D(c[1245]), .CLK(clk), .RST(rst), .Q(sreg[1243]) );
  DFF \sreg_reg[1242]  ( .D(c[1244]), .CLK(clk), .RST(rst), .Q(sreg[1242]) );
  DFF \sreg_reg[1241]  ( .D(c[1243]), .CLK(clk), .RST(rst), .Q(sreg[1241]) );
  DFF \sreg_reg[1240]  ( .D(c[1242]), .CLK(clk), .RST(rst), .Q(sreg[1240]) );
  DFF \sreg_reg[1239]  ( .D(c[1241]), .CLK(clk), .RST(rst), .Q(sreg[1239]) );
  DFF \sreg_reg[1238]  ( .D(c[1240]), .CLK(clk), .RST(rst), .Q(sreg[1238]) );
  DFF \sreg_reg[1237]  ( .D(c[1239]), .CLK(clk), .RST(rst), .Q(sreg[1237]) );
  DFF \sreg_reg[1236]  ( .D(c[1238]), .CLK(clk), .RST(rst), .Q(sreg[1236]) );
  DFF \sreg_reg[1235]  ( .D(c[1237]), .CLK(clk), .RST(rst), .Q(sreg[1235]) );
  DFF \sreg_reg[1234]  ( .D(c[1236]), .CLK(clk), .RST(rst), .Q(sreg[1234]) );
  DFF \sreg_reg[1233]  ( .D(c[1235]), .CLK(clk), .RST(rst), .Q(sreg[1233]) );
  DFF \sreg_reg[1232]  ( .D(c[1234]), .CLK(clk), .RST(rst), .Q(sreg[1232]) );
  DFF \sreg_reg[1231]  ( .D(c[1233]), .CLK(clk), .RST(rst), .Q(sreg[1231]) );
  DFF \sreg_reg[1230]  ( .D(c[1232]), .CLK(clk), .RST(rst), .Q(sreg[1230]) );
  DFF \sreg_reg[1229]  ( .D(c[1231]), .CLK(clk), .RST(rst), .Q(sreg[1229]) );
  DFF \sreg_reg[1228]  ( .D(c[1230]), .CLK(clk), .RST(rst), .Q(sreg[1228]) );
  DFF \sreg_reg[1227]  ( .D(c[1229]), .CLK(clk), .RST(rst), .Q(sreg[1227]) );
  DFF \sreg_reg[1226]  ( .D(c[1228]), .CLK(clk), .RST(rst), .Q(sreg[1226]) );
  DFF \sreg_reg[1225]  ( .D(c[1227]), .CLK(clk), .RST(rst), .Q(sreg[1225]) );
  DFF \sreg_reg[1224]  ( .D(c[1226]), .CLK(clk), .RST(rst), .Q(sreg[1224]) );
  DFF \sreg_reg[1223]  ( .D(c[1225]), .CLK(clk), .RST(rst), .Q(sreg[1223]) );
  DFF \sreg_reg[1222]  ( .D(c[1224]), .CLK(clk), .RST(rst), .Q(sreg[1222]) );
  DFF \sreg_reg[1221]  ( .D(c[1223]), .CLK(clk), .RST(rst), .Q(sreg[1221]) );
  DFF \sreg_reg[1220]  ( .D(c[1222]), .CLK(clk), .RST(rst), .Q(sreg[1220]) );
  DFF \sreg_reg[1219]  ( .D(c[1221]), .CLK(clk), .RST(rst), .Q(sreg[1219]) );
  DFF \sreg_reg[1218]  ( .D(c[1220]), .CLK(clk), .RST(rst), .Q(sreg[1218]) );
  DFF \sreg_reg[1217]  ( .D(c[1219]), .CLK(clk), .RST(rst), .Q(sreg[1217]) );
  DFF \sreg_reg[1216]  ( .D(c[1218]), .CLK(clk), .RST(rst), .Q(sreg[1216]) );
  DFF \sreg_reg[1215]  ( .D(c[1217]), .CLK(clk), .RST(rst), .Q(sreg[1215]) );
  DFF \sreg_reg[1214]  ( .D(c[1216]), .CLK(clk), .RST(rst), .Q(sreg[1214]) );
  DFF \sreg_reg[1213]  ( .D(c[1215]), .CLK(clk), .RST(rst), .Q(sreg[1213]) );
  DFF \sreg_reg[1212]  ( .D(c[1214]), .CLK(clk), .RST(rst), .Q(sreg[1212]) );
  DFF \sreg_reg[1211]  ( .D(c[1213]), .CLK(clk), .RST(rst), .Q(sreg[1211]) );
  DFF \sreg_reg[1210]  ( .D(c[1212]), .CLK(clk), .RST(rst), .Q(sreg[1210]) );
  DFF \sreg_reg[1209]  ( .D(c[1211]), .CLK(clk), .RST(rst), .Q(sreg[1209]) );
  DFF \sreg_reg[1208]  ( .D(c[1210]), .CLK(clk), .RST(rst), .Q(sreg[1208]) );
  DFF \sreg_reg[1207]  ( .D(c[1209]), .CLK(clk), .RST(rst), .Q(sreg[1207]) );
  DFF \sreg_reg[1206]  ( .D(c[1208]), .CLK(clk), .RST(rst), .Q(sreg[1206]) );
  DFF \sreg_reg[1205]  ( .D(c[1207]), .CLK(clk), .RST(rst), .Q(sreg[1205]) );
  DFF \sreg_reg[1204]  ( .D(c[1206]), .CLK(clk), .RST(rst), .Q(sreg[1204]) );
  DFF \sreg_reg[1203]  ( .D(c[1205]), .CLK(clk), .RST(rst), .Q(sreg[1203]) );
  DFF \sreg_reg[1202]  ( .D(c[1204]), .CLK(clk), .RST(rst), .Q(sreg[1202]) );
  DFF \sreg_reg[1201]  ( .D(c[1203]), .CLK(clk), .RST(rst), .Q(sreg[1201]) );
  DFF \sreg_reg[1200]  ( .D(c[1202]), .CLK(clk), .RST(rst), .Q(sreg[1200]) );
  DFF \sreg_reg[1199]  ( .D(c[1201]), .CLK(clk), .RST(rst), .Q(sreg[1199]) );
  DFF \sreg_reg[1198]  ( .D(c[1200]), .CLK(clk), .RST(rst), .Q(sreg[1198]) );
  DFF \sreg_reg[1197]  ( .D(c[1199]), .CLK(clk), .RST(rst), .Q(sreg[1197]) );
  DFF \sreg_reg[1196]  ( .D(c[1198]), .CLK(clk), .RST(rst), .Q(sreg[1196]) );
  DFF \sreg_reg[1195]  ( .D(c[1197]), .CLK(clk), .RST(rst), .Q(sreg[1195]) );
  DFF \sreg_reg[1194]  ( .D(c[1196]), .CLK(clk), .RST(rst), .Q(sreg[1194]) );
  DFF \sreg_reg[1193]  ( .D(c[1195]), .CLK(clk), .RST(rst), .Q(sreg[1193]) );
  DFF \sreg_reg[1192]  ( .D(c[1194]), .CLK(clk), .RST(rst), .Q(sreg[1192]) );
  DFF \sreg_reg[1191]  ( .D(c[1193]), .CLK(clk), .RST(rst), .Q(sreg[1191]) );
  DFF \sreg_reg[1190]  ( .D(c[1192]), .CLK(clk), .RST(rst), .Q(sreg[1190]) );
  DFF \sreg_reg[1189]  ( .D(c[1191]), .CLK(clk), .RST(rst), .Q(sreg[1189]) );
  DFF \sreg_reg[1188]  ( .D(c[1190]), .CLK(clk), .RST(rst), .Q(sreg[1188]) );
  DFF \sreg_reg[1187]  ( .D(c[1189]), .CLK(clk), .RST(rst), .Q(sreg[1187]) );
  DFF \sreg_reg[1186]  ( .D(c[1188]), .CLK(clk), .RST(rst), .Q(sreg[1186]) );
  DFF \sreg_reg[1185]  ( .D(c[1187]), .CLK(clk), .RST(rst), .Q(sreg[1185]) );
  DFF \sreg_reg[1184]  ( .D(c[1186]), .CLK(clk), .RST(rst), .Q(sreg[1184]) );
  DFF \sreg_reg[1183]  ( .D(c[1185]), .CLK(clk), .RST(rst), .Q(sreg[1183]) );
  DFF \sreg_reg[1182]  ( .D(c[1184]), .CLK(clk), .RST(rst), .Q(sreg[1182]) );
  DFF \sreg_reg[1181]  ( .D(c[1183]), .CLK(clk), .RST(rst), .Q(sreg[1181]) );
  DFF \sreg_reg[1180]  ( .D(c[1182]), .CLK(clk), .RST(rst), .Q(sreg[1180]) );
  DFF \sreg_reg[1179]  ( .D(c[1181]), .CLK(clk), .RST(rst), .Q(sreg[1179]) );
  DFF \sreg_reg[1178]  ( .D(c[1180]), .CLK(clk), .RST(rst), .Q(sreg[1178]) );
  DFF \sreg_reg[1177]  ( .D(c[1179]), .CLK(clk), .RST(rst), .Q(sreg[1177]) );
  DFF \sreg_reg[1176]  ( .D(c[1178]), .CLK(clk), .RST(rst), .Q(sreg[1176]) );
  DFF \sreg_reg[1175]  ( .D(c[1177]), .CLK(clk), .RST(rst), .Q(sreg[1175]) );
  DFF \sreg_reg[1174]  ( .D(c[1176]), .CLK(clk), .RST(rst), .Q(sreg[1174]) );
  DFF \sreg_reg[1173]  ( .D(c[1175]), .CLK(clk), .RST(rst), .Q(sreg[1173]) );
  DFF \sreg_reg[1172]  ( .D(c[1174]), .CLK(clk), .RST(rst), .Q(sreg[1172]) );
  DFF \sreg_reg[1171]  ( .D(c[1173]), .CLK(clk), .RST(rst), .Q(sreg[1171]) );
  DFF \sreg_reg[1170]  ( .D(c[1172]), .CLK(clk), .RST(rst), .Q(sreg[1170]) );
  DFF \sreg_reg[1169]  ( .D(c[1171]), .CLK(clk), .RST(rst), .Q(sreg[1169]) );
  DFF \sreg_reg[1168]  ( .D(c[1170]), .CLK(clk), .RST(rst), .Q(sreg[1168]) );
  DFF \sreg_reg[1167]  ( .D(c[1169]), .CLK(clk), .RST(rst), .Q(sreg[1167]) );
  DFF \sreg_reg[1166]  ( .D(c[1168]), .CLK(clk), .RST(rst), .Q(sreg[1166]) );
  DFF \sreg_reg[1165]  ( .D(c[1167]), .CLK(clk), .RST(rst), .Q(sreg[1165]) );
  DFF \sreg_reg[1164]  ( .D(c[1166]), .CLK(clk), .RST(rst), .Q(sreg[1164]) );
  DFF \sreg_reg[1163]  ( .D(c[1165]), .CLK(clk), .RST(rst), .Q(sreg[1163]) );
  DFF \sreg_reg[1162]  ( .D(c[1164]), .CLK(clk), .RST(rst), .Q(sreg[1162]) );
  DFF \sreg_reg[1161]  ( .D(c[1163]), .CLK(clk), .RST(rst), .Q(sreg[1161]) );
  DFF \sreg_reg[1160]  ( .D(c[1162]), .CLK(clk), .RST(rst), .Q(sreg[1160]) );
  DFF \sreg_reg[1159]  ( .D(c[1161]), .CLK(clk), .RST(rst), .Q(sreg[1159]) );
  DFF \sreg_reg[1158]  ( .D(c[1160]), .CLK(clk), .RST(rst), .Q(sreg[1158]) );
  DFF \sreg_reg[1157]  ( .D(c[1159]), .CLK(clk), .RST(rst), .Q(sreg[1157]) );
  DFF \sreg_reg[1156]  ( .D(c[1158]), .CLK(clk), .RST(rst), .Q(sreg[1156]) );
  DFF \sreg_reg[1155]  ( .D(c[1157]), .CLK(clk), .RST(rst), .Q(sreg[1155]) );
  DFF \sreg_reg[1154]  ( .D(c[1156]), .CLK(clk), .RST(rst), .Q(sreg[1154]) );
  DFF \sreg_reg[1153]  ( .D(c[1155]), .CLK(clk), .RST(rst), .Q(sreg[1153]) );
  DFF \sreg_reg[1152]  ( .D(c[1154]), .CLK(clk), .RST(rst), .Q(sreg[1152]) );
  DFF \sreg_reg[1151]  ( .D(c[1153]), .CLK(clk), .RST(rst), .Q(sreg[1151]) );
  DFF \sreg_reg[1150]  ( .D(c[1152]), .CLK(clk), .RST(rst), .Q(sreg[1150]) );
  DFF \sreg_reg[1149]  ( .D(c[1151]), .CLK(clk), .RST(rst), .Q(sreg[1149]) );
  DFF \sreg_reg[1148]  ( .D(c[1150]), .CLK(clk), .RST(rst), .Q(sreg[1148]) );
  DFF \sreg_reg[1147]  ( .D(c[1149]), .CLK(clk), .RST(rst), .Q(sreg[1147]) );
  DFF \sreg_reg[1146]  ( .D(c[1148]), .CLK(clk), .RST(rst), .Q(sreg[1146]) );
  DFF \sreg_reg[1145]  ( .D(c[1147]), .CLK(clk), .RST(rst), .Q(sreg[1145]) );
  DFF \sreg_reg[1144]  ( .D(c[1146]), .CLK(clk), .RST(rst), .Q(sreg[1144]) );
  DFF \sreg_reg[1143]  ( .D(c[1145]), .CLK(clk), .RST(rst), .Q(sreg[1143]) );
  DFF \sreg_reg[1142]  ( .D(c[1144]), .CLK(clk), .RST(rst), .Q(sreg[1142]) );
  DFF \sreg_reg[1141]  ( .D(c[1143]), .CLK(clk), .RST(rst), .Q(sreg[1141]) );
  DFF \sreg_reg[1140]  ( .D(c[1142]), .CLK(clk), .RST(rst), .Q(sreg[1140]) );
  DFF \sreg_reg[1139]  ( .D(c[1141]), .CLK(clk), .RST(rst), .Q(sreg[1139]) );
  DFF \sreg_reg[1138]  ( .D(c[1140]), .CLK(clk), .RST(rst), .Q(sreg[1138]) );
  DFF \sreg_reg[1137]  ( .D(c[1139]), .CLK(clk), .RST(rst), .Q(sreg[1137]) );
  DFF \sreg_reg[1136]  ( .D(c[1138]), .CLK(clk), .RST(rst), .Q(sreg[1136]) );
  DFF \sreg_reg[1135]  ( .D(c[1137]), .CLK(clk), .RST(rst), .Q(sreg[1135]) );
  DFF \sreg_reg[1134]  ( .D(c[1136]), .CLK(clk), .RST(rst), .Q(sreg[1134]) );
  DFF \sreg_reg[1133]  ( .D(c[1135]), .CLK(clk), .RST(rst), .Q(sreg[1133]) );
  DFF \sreg_reg[1132]  ( .D(c[1134]), .CLK(clk), .RST(rst), .Q(sreg[1132]) );
  DFF \sreg_reg[1131]  ( .D(c[1133]), .CLK(clk), .RST(rst), .Q(sreg[1131]) );
  DFF \sreg_reg[1130]  ( .D(c[1132]), .CLK(clk), .RST(rst), .Q(sreg[1130]) );
  DFF \sreg_reg[1129]  ( .D(c[1131]), .CLK(clk), .RST(rst), .Q(sreg[1129]) );
  DFF \sreg_reg[1128]  ( .D(c[1130]), .CLK(clk), .RST(rst), .Q(sreg[1128]) );
  DFF \sreg_reg[1127]  ( .D(c[1129]), .CLK(clk), .RST(rst), .Q(sreg[1127]) );
  DFF \sreg_reg[1126]  ( .D(c[1128]), .CLK(clk), .RST(rst), .Q(sreg[1126]) );
  DFF \sreg_reg[1125]  ( .D(c[1127]), .CLK(clk), .RST(rst), .Q(sreg[1125]) );
  DFF \sreg_reg[1124]  ( .D(c[1126]), .CLK(clk), .RST(rst), .Q(sreg[1124]) );
  DFF \sreg_reg[1123]  ( .D(c[1125]), .CLK(clk), .RST(rst), .Q(sreg[1123]) );
  DFF \sreg_reg[1122]  ( .D(c[1124]), .CLK(clk), .RST(rst), .Q(sreg[1122]) );
  DFF \sreg_reg[1121]  ( .D(c[1123]), .CLK(clk), .RST(rst), .Q(sreg[1121]) );
  DFF \sreg_reg[1120]  ( .D(c[1122]), .CLK(clk), .RST(rst), .Q(sreg[1120]) );
  DFF \sreg_reg[1119]  ( .D(c[1121]), .CLK(clk), .RST(rst), .Q(sreg[1119]) );
  DFF \sreg_reg[1118]  ( .D(c[1120]), .CLK(clk), .RST(rst), .Q(sreg[1118]) );
  DFF \sreg_reg[1117]  ( .D(c[1119]), .CLK(clk), .RST(rst), .Q(sreg[1117]) );
  DFF \sreg_reg[1116]  ( .D(c[1118]), .CLK(clk), .RST(rst), .Q(sreg[1116]) );
  DFF \sreg_reg[1115]  ( .D(c[1117]), .CLK(clk), .RST(rst), .Q(sreg[1115]) );
  DFF \sreg_reg[1114]  ( .D(c[1116]), .CLK(clk), .RST(rst), .Q(sreg[1114]) );
  DFF \sreg_reg[1113]  ( .D(c[1115]), .CLK(clk), .RST(rst), .Q(sreg[1113]) );
  DFF \sreg_reg[1112]  ( .D(c[1114]), .CLK(clk), .RST(rst), .Q(sreg[1112]) );
  DFF \sreg_reg[1111]  ( .D(c[1113]), .CLK(clk), .RST(rst), .Q(sreg[1111]) );
  DFF \sreg_reg[1110]  ( .D(c[1112]), .CLK(clk), .RST(rst), .Q(sreg[1110]) );
  DFF \sreg_reg[1109]  ( .D(c[1111]), .CLK(clk), .RST(rst), .Q(sreg[1109]) );
  DFF \sreg_reg[1108]  ( .D(c[1110]), .CLK(clk), .RST(rst), .Q(sreg[1108]) );
  DFF \sreg_reg[1107]  ( .D(c[1109]), .CLK(clk), .RST(rst), .Q(sreg[1107]) );
  DFF \sreg_reg[1106]  ( .D(c[1108]), .CLK(clk), .RST(rst), .Q(sreg[1106]) );
  DFF \sreg_reg[1105]  ( .D(c[1107]), .CLK(clk), .RST(rst), .Q(sreg[1105]) );
  DFF \sreg_reg[1104]  ( .D(c[1106]), .CLK(clk), .RST(rst), .Q(sreg[1104]) );
  DFF \sreg_reg[1103]  ( .D(c[1105]), .CLK(clk), .RST(rst), .Q(sreg[1103]) );
  DFF \sreg_reg[1102]  ( .D(c[1104]), .CLK(clk), .RST(rst), .Q(sreg[1102]) );
  DFF \sreg_reg[1101]  ( .D(c[1103]), .CLK(clk), .RST(rst), .Q(sreg[1101]) );
  DFF \sreg_reg[1100]  ( .D(c[1102]), .CLK(clk), .RST(rst), .Q(sreg[1100]) );
  DFF \sreg_reg[1099]  ( .D(c[1101]), .CLK(clk), .RST(rst), .Q(sreg[1099]) );
  DFF \sreg_reg[1098]  ( .D(c[1100]), .CLK(clk), .RST(rst), .Q(sreg[1098]) );
  DFF \sreg_reg[1097]  ( .D(c[1099]), .CLK(clk), .RST(rst), .Q(sreg[1097]) );
  DFF \sreg_reg[1096]  ( .D(c[1098]), .CLK(clk), .RST(rst), .Q(sreg[1096]) );
  DFF \sreg_reg[1095]  ( .D(c[1097]), .CLK(clk), .RST(rst), .Q(sreg[1095]) );
  DFF \sreg_reg[1094]  ( .D(c[1096]), .CLK(clk), .RST(rst), .Q(sreg[1094]) );
  DFF \sreg_reg[1093]  ( .D(c[1095]), .CLK(clk), .RST(rst), .Q(sreg[1093]) );
  DFF \sreg_reg[1092]  ( .D(c[1094]), .CLK(clk), .RST(rst), .Q(sreg[1092]) );
  DFF \sreg_reg[1091]  ( .D(c[1093]), .CLK(clk), .RST(rst), .Q(sreg[1091]) );
  DFF \sreg_reg[1090]  ( .D(c[1092]), .CLK(clk), .RST(rst), .Q(sreg[1090]) );
  DFF \sreg_reg[1089]  ( .D(c[1091]), .CLK(clk), .RST(rst), .Q(sreg[1089]) );
  DFF \sreg_reg[1088]  ( .D(c[1090]), .CLK(clk), .RST(rst), .Q(sreg[1088]) );
  DFF \sreg_reg[1087]  ( .D(c[1089]), .CLK(clk), .RST(rst), .Q(sreg[1087]) );
  DFF \sreg_reg[1086]  ( .D(c[1088]), .CLK(clk), .RST(rst), .Q(sreg[1086]) );
  DFF \sreg_reg[1085]  ( .D(c[1087]), .CLK(clk), .RST(rst), .Q(sreg[1085]) );
  DFF \sreg_reg[1084]  ( .D(c[1086]), .CLK(clk), .RST(rst), .Q(sreg[1084]) );
  DFF \sreg_reg[1083]  ( .D(c[1085]), .CLK(clk), .RST(rst), .Q(sreg[1083]) );
  DFF \sreg_reg[1082]  ( .D(c[1084]), .CLK(clk), .RST(rst), .Q(sreg[1082]) );
  DFF \sreg_reg[1081]  ( .D(c[1083]), .CLK(clk), .RST(rst), .Q(sreg[1081]) );
  DFF \sreg_reg[1080]  ( .D(c[1082]), .CLK(clk), .RST(rst), .Q(sreg[1080]) );
  DFF \sreg_reg[1079]  ( .D(c[1081]), .CLK(clk), .RST(rst), .Q(sreg[1079]) );
  DFF \sreg_reg[1078]  ( .D(c[1080]), .CLK(clk), .RST(rst), .Q(sreg[1078]) );
  DFF \sreg_reg[1077]  ( .D(c[1079]), .CLK(clk), .RST(rst), .Q(sreg[1077]) );
  DFF \sreg_reg[1076]  ( .D(c[1078]), .CLK(clk), .RST(rst), .Q(sreg[1076]) );
  DFF \sreg_reg[1075]  ( .D(c[1077]), .CLK(clk), .RST(rst), .Q(sreg[1075]) );
  DFF \sreg_reg[1074]  ( .D(c[1076]), .CLK(clk), .RST(rst), .Q(sreg[1074]) );
  DFF \sreg_reg[1073]  ( .D(c[1075]), .CLK(clk), .RST(rst), .Q(sreg[1073]) );
  DFF \sreg_reg[1072]  ( .D(c[1074]), .CLK(clk), .RST(rst), .Q(sreg[1072]) );
  DFF \sreg_reg[1071]  ( .D(c[1073]), .CLK(clk), .RST(rst), .Q(sreg[1071]) );
  DFF \sreg_reg[1070]  ( .D(c[1072]), .CLK(clk), .RST(rst), .Q(sreg[1070]) );
  DFF \sreg_reg[1069]  ( .D(c[1071]), .CLK(clk), .RST(rst), .Q(sreg[1069]) );
  DFF \sreg_reg[1068]  ( .D(c[1070]), .CLK(clk), .RST(rst), .Q(sreg[1068]) );
  DFF \sreg_reg[1067]  ( .D(c[1069]), .CLK(clk), .RST(rst), .Q(sreg[1067]) );
  DFF \sreg_reg[1066]  ( .D(c[1068]), .CLK(clk), .RST(rst), .Q(sreg[1066]) );
  DFF \sreg_reg[1065]  ( .D(c[1067]), .CLK(clk), .RST(rst), .Q(sreg[1065]) );
  DFF \sreg_reg[1064]  ( .D(c[1066]), .CLK(clk), .RST(rst), .Q(sreg[1064]) );
  DFF \sreg_reg[1063]  ( .D(c[1065]), .CLK(clk), .RST(rst), .Q(sreg[1063]) );
  DFF \sreg_reg[1062]  ( .D(c[1064]), .CLK(clk), .RST(rst), .Q(sreg[1062]) );
  DFF \sreg_reg[1061]  ( .D(c[1063]), .CLK(clk), .RST(rst), .Q(sreg[1061]) );
  DFF \sreg_reg[1060]  ( .D(c[1062]), .CLK(clk), .RST(rst), .Q(sreg[1060]) );
  DFF \sreg_reg[1059]  ( .D(c[1061]), .CLK(clk), .RST(rst), .Q(sreg[1059]) );
  DFF \sreg_reg[1058]  ( .D(c[1060]), .CLK(clk), .RST(rst), .Q(sreg[1058]) );
  DFF \sreg_reg[1057]  ( .D(c[1059]), .CLK(clk), .RST(rst), .Q(sreg[1057]) );
  DFF \sreg_reg[1056]  ( .D(c[1058]), .CLK(clk), .RST(rst), .Q(sreg[1056]) );
  DFF \sreg_reg[1055]  ( .D(c[1057]), .CLK(clk), .RST(rst), .Q(sreg[1055]) );
  DFF \sreg_reg[1054]  ( .D(c[1056]), .CLK(clk), .RST(rst), .Q(sreg[1054]) );
  DFF \sreg_reg[1053]  ( .D(c[1055]), .CLK(clk), .RST(rst), .Q(sreg[1053]) );
  DFF \sreg_reg[1052]  ( .D(c[1054]), .CLK(clk), .RST(rst), .Q(sreg[1052]) );
  DFF \sreg_reg[1051]  ( .D(c[1053]), .CLK(clk), .RST(rst), .Q(sreg[1051]) );
  DFF \sreg_reg[1050]  ( .D(c[1052]), .CLK(clk), .RST(rst), .Q(sreg[1050]) );
  DFF \sreg_reg[1049]  ( .D(c[1051]), .CLK(clk), .RST(rst), .Q(sreg[1049]) );
  DFF \sreg_reg[1048]  ( .D(c[1050]), .CLK(clk), .RST(rst), .Q(sreg[1048]) );
  DFF \sreg_reg[1047]  ( .D(c[1049]), .CLK(clk), .RST(rst), .Q(sreg[1047]) );
  DFF \sreg_reg[1046]  ( .D(c[1048]), .CLK(clk), .RST(rst), .Q(sreg[1046]) );
  DFF \sreg_reg[1045]  ( .D(c[1047]), .CLK(clk), .RST(rst), .Q(sreg[1045]) );
  DFF \sreg_reg[1044]  ( .D(c[1046]), .CLK(clk), .RST(rst), .Q(sreg[1044]) );
  DFF \sreg_reg[1043]  ( .D(c[1045]), .CLK(clk), .RST(rst), .Q(sreg[1043]) );
  DFF \sreg_reg[1042]  ( .D(c[1044]), .CLK(clk), .RST(rst), .Q(sreg[1042]) );
  DFF \sreg_reg[1041]  ( .D(c[1043]), .CLK(clk), .RST(rst), .Q(sreg[1041]) );
  DFF \sreg_reg[1040]  ( .D(c[1042]), .CLK(clk), .RST(rst), .Q(sreg[1040]) );
  DFF \sreg_reg[1039]  ( .D(c[1041]), .CLK(clk), .RST(rst), .Q(sreg[1039]) );
  DFF \sreg_reg[1038]  ( .D(c[1040]), .CLK(clk), .RST(rst), .Q(sreg[1038]) );
  DFF \sreg_reg[1037]  ( .D(c[1039]), .CLK(clk), .RST(rst), .Q(sreg[1037]) );
  DFF \sreg_reg[1036]  ( .D(c[1038]), .CLK(clk), .RST(rst), .Q(sreg[1036]) );
  DFF \sreg_reg[1035]  ( .D(c[1037]), .CLK(clk), .RST(rst), .Q(sreg[1035]) );
  DFF \sreg_reg[1034]  ( .D(c[1036]), .CLK(clk), .RST(rst), .Q(sreg[1034]) );
  DFF \sreg_reg[1033]  ( .D(c[1035]), .CLK(clk), .RST(rst), .Q(sreg[1033]) );
  DFF \sreg_reg[1032]  ( .D(c[1034]), .CLK(clk), .RST(rst), .Q(sreg[1032]) );
  DFF \sreg_reg[1031]  ( .D(c[1033]), .CLK(clk), .RST(rst), .Q(sreg[1031]) );
  DFF \sreg_reg[1030]  ( .D(c[1032]), .CLK(clk), .RST(rst), .Q(sreg[1030]) );
  DFF \sreg_reg[1029]  ( .D(c[1031]), .CLK(clk), .RST(rst), .Q(sreg[1029]) );
  DFF \sreg_reg[1028]  ( .D(c[1030]), .CLK(clk), .RST(rst), .Q(sreg[1028]) );
  DFF \sreg_reg[1027]  ( .D(c[1029]), .CLK(clk), .RST(rst), .Q(sreg[1027]) );
  DFF \sreg_reg[1026]  ( .D(c[1028]), .CLK(clk), .RST(rst), .Q(sreg[1026]) );
  DFF \sreg_reg[1025]  ( .D(c[1027]), .CLK(clk), .RST(rst), .Q(sreg[1025]) );
  DFF \sreg_reg[1024]  ( .D(c[1026]), .CLK(clk), .RST(rst), .Q(sreg[1024]) );
  DFF \sreg_reg[1023]  ( .D(c[1025]), .CLK(clk), .RST(rst), .Q(sreg[1023]) );
  DFF \sreg_reg[1022]  ( .D(c[1024]), .CLK(clk), .RST(rst), .Q(sreg[1022]) );
  DFF \sreg_reg[1021]  ( .D(c[1023]), .CLK(clk), .RST(rst), .Q(c[1021]) );
  DFF \sreg_reg[1020]  ( .D(c[1022]), .CLK(clk), .RST(rst), .Q(c[1020]) );
  DFF \sreg_reg[1019]  ( .D(c[1021]), .CLK(clk), .RST(rst), .Q(c[1019]) );
  DFF \sreg_reg[1018]  ( .D(c[1020]), .CLK(clk), .RST(rst), .Q(c[1018]) );
  DFF \sreg_reg[1017]  ( .D(c[1019]), .CLK(clk), .RST(rst), .Q(c[1017]) );
  DFF \sreg_reg[1016]  ( .D(c[1018]), .CLK(clk), .RST(rst), .Q(c[1016]) );
  DFF \sreg_reg[1015]  ( .D(c[1017]), .CLK(clk), .RST(rst), .Q(c[1015]) );
  DFF \sreg_reg[1014]  ( .D(c[1016]), .CLK(clk), .RST(rst), .Q(c[1014]) );
  DFF \sreg_reg[1013]  ( .D(c[1015]), .CLK(clk), .RST(rst), .Q(c[1013]) );
  DFF \sreg_reg[1012]  ( .D(c[1014]), .CLK(clk), .RST(rst), .Q(c[1012]) );
  DFF \sreg_reg[1011]  ( .D(c[1013]), .CLK(clk), .RST(rst), .Q(c[1011]) );
  DFF \sreg_reg[1010]  ( .D(c[1012]), .CLK(clk), .RST(rst), .Q(c[1010]) );
  DFF \sreg_reg[1009]  ( .D(c[1011]), .CLK(clk), .RST(rst), .Q(c[1009]) );
  DFF \sreg_reg[1008]  ( .D(c[1010]), .CLK(clk), .RST(rst), .Q(c[1008]) );
  DFF \sreg_reg[1007]  ( .D(c[1009]), .CLK(clk), .RST(rst), .Q(c[1007]) );
  DFF \sreg_reg[1006]  ( .D(c[1008]), .CLK(clk), .RST(rst), .Q(c[1006]) );
  DFF \sreg_reg[1005]  ( .D(c[1007]), .CLK(clk), .RST(rst), .Q(c[1005]) );
  DFF \sreg_reg[1004]  ( .D(c[1006]), .CLK(clk), .RST(rst), .Q(c[1004]) );
  DFF \sreg_reg[1003]  ( .D(c[1005]), .CLK(clk), .RST(rst), .Q(c[1003]) );
  DFF \sreg_reg[1002]  ( .D(c[1004]), .CLK(clk), .RST(rst), .Q(c[1002]) );
  DFF \sreg_reg[1001]  ( .D(c[1003]), .CLK(clk), .RST(rst), .Q(c[1001]) );
  DFF \sreg_reg[1000]  ( .D(c[1002]), .CLK(clk), .RST(rst), .Q(c[1000]) );
  DFF \sreg_reg[999]  ( .D(c[1001]), .CLK(clk), .RST(rst), .Q(c[999]) );
  DFF \sreg_reg[998]  ( .D(c[1000]), .CLK(clk), .RST(rst), .Q(c[998]) );
  DFF \sreg_reg[997]  ( .D(c[999]), .CLK(clk), .RST(rst), .Q(c[997]) );
  DFF \sreg_reg[996]  ( .D(c[998]), .CLK(clk), .RST(rst), .Q(c[996]) );
  DFF \sreg_reg[995]  ( .D(c[997]), .CLK(clk), .RST(rst), .Q(c[995]) );
  DFF \sreg_reg[994]  ( .D(c[996]), .CLK(clk), .RST(rst), .Q(c[994]) );
  DFF \sreg_reg[993]  ( .D(c[995]), .CLK(clk), .RST(rst), .Q(c[993]) );
  DFF \sreg_reg[992]  ( .D(c[994]), .CLK(clk), .RST(rst), .Q(c[992]) );
  DFF \sreg_reg[991]  ( .D(c[993]), .CLK(clk), .RST(rst), .Q(c[991]) );
  DFF \sreg_reg[990]  ( .D(c[992]), .CLK(clk), .RST(rst), .Q(c[990]) );
  DFF \sreg_reg[989]  ( .D(c[991]), .CLK(clk), .RST(rst), .Q(c[989]) );
  DFF \sreg_reg[988]  ( .D(c[990]), .CLK(clk), .RST(rst), .Q(c[988]) );
  DFF \sreg_reg[987]  ( .D(c[989]), .CLK(clk), .RST(rst), .Q(c[987]) );
  DFF \sreg_reg[986]  ( .D(c[988]), .CLK(clk), .RST(rst), .Q(c[986]) );
  DFF \sreg_reg[985]  ( .D(c[987]), .CLK(clk), .RST(rst), .Q(c[985]) );
  DFF \sreg_reg[984]  ( .D(c[986]), .CLK(clk), .RST(rst), .Q(c[984]) );
  DFF \sreg_reg[983]  ( .D(c[985]), .CLK(clk), .RST(rst), .Q(c[983]) );
  DFF \sreg_reg[982]  ( .D(c[984]), .CLK(clk), .RST(rst), .Q(c[982]) );
  DFF \sreg_reg[981]  ( .D(c[983]), .CLK(clk), .RST(rst), .Q(c[981]) );
  DFF \sreg_reg[980]  ( .D(c[982]), .CLK(clk), .RST(rst), .Q(c[980]) );
  DFF \sreg_reg[979]  ( .D(c[981]), .CLK(clk), .RST(rst), .Q(c[979]) );
  DFF \sreg_reg[978]  ( .D(c[980]), .CLK(clk), .RST(rst), .Q(c[978]) );
  DFF \sreg_reg[977]  ( .D(c[979]), .CLK(clk), .RST(rst), .Q(c[977]) );
  DFF \sreg_reg[976]  ( .D(c[978]), .CLK(clk), .RST(rst), .Q(c[976]) );
  DFF \sreg_reg[975]  ( .D(c[977]), .CLK(clk), .RST(rst), .Q(c[975]) );
  DFF \sreg_reg[974]  ( .D(c[976]), .CLK(clk), .RST(rst), .Q(c[974]) );
  DFF \sreg_reg[973]  ( .D(c[975]), .CLK(clk), .RST(rst), .Q(c[973]) );
  DFF \sreg_reg[972]  ( .D(c[974]), .CLK(clk), .RST(rst), .Q(c[972]) );
  DFF \sreg_reg[971]  ( .D(c[973]), .CLK(clk), .RST(rst), .Q(c[971]) );
  DFF \sreg_reg[970]  ( .D(c[972]), .CLK(clk), .RST(rst), .Q(c[970]) );
  DFF \sreg_reg[969]  ( .D(c[971]), .CLK(clk), .RST(rst), .Q(c[969]) );
  DFF \sreg_reg[968]  ( .D(c[970]), .CLK(clk), .RST(rst), .Q(c[968]) );
  DFF \sreg_reg[967]  ( .D(c[969]), .CLK(clk), .RST(rst), .Q(c[967]) );
  DFF \sreg_reg[966]  ( .D(c[968]), .CLK(clk), .RST(rst), .Q(c[966]) );
  DFF \sreg_reg[965]  ( .D(c[967]), .CLK(clk), .RST(rst), .Q(c[965]) );
  DFF \sreg_reg[964]  ( .D(c[966]), .CLK(clk), .RST(rst), .Q(c[964]) );
  DFF \sreg_reg[963]  ( .D(c[965]), .CLK(clk), .RST(rst), .Q(c[963]) );
  DFF \sreg_reg[962]  ( .D(c[964]), .CLK(clk), .RST(rst), .Q(c[962]) );
  DFF \sreg_reg[961]  ( .D(c[963]), .CLK(clk), .RST(rst), .Q(c[961]) );
  DFF \sreg_reg[960]  ( .D(c[962]), .CLK(clk), .RST(rst), .Q(c[960]) );
  DFF \sreg_reg[959]  ( .D(c[961]), .CLK(clk), .RST(rst), .Q(c[959]) );
  DFF \sreg_reg[958]  ( .D(c[960]), .CLK(clk), .RST(rst), .Q(c[958]) );
  DFF \sreg_reg[957]  ( .D(c[959]), .CLK(clk), .RST(rst), .Q(c[957]) );
  DFF \sreg_reg[956]  ( .D(c[958]), .CLK(clk), .RST(rst), .Q(c[956]) );
  DFF \sreg_reg[955]  ( .D(c[957]), .CLK(clk), .RST(rst), .Q(c[955]) );
  DFF \sreg_reg[954]  ( .D(c[956]), .CLK(clk), .RST(rst), .Q(c[954]) );
  DFF \sreg_reg[953]  ( .D(c[955]), .CLK(clk), .RST(rst), .Q(c[953]) );
  DFF \sreg_reg[952]  ( .D(c[954]), .CLK(clk), .RST(rst), .Q(c[952]) );
  DFF \sreg_reg[951]  ( .D(c[953]), .CLK(clk), .RST(rst), .Q(c[951]) );
  DFF \sreg_reg[950]  ( .D(c[952]), .CLK(clk), .RST(rst), .Q(c[950]) );
  DFF \sreg_reg[949]  ( .D(c[951]), .CLK(clk), .RST(rst), .Q(c[949]) );
  DFF \sreg_reg[948]  ( .D(c[950]), .CLK(clk), .RST(rst), .Q(c[948]) );
  DFF \sreg_reg[947]  ( .D(c[949]), .CLK(clk), .RST(rst), .Q(c[947]) );
  DFF \sreg_reg[946]  ( .D(c[948]), .CLK(clk), .RST(rst), .Q(c[946]) );
  DFF \sreg_reg[945]  ( .D(c[947]), .CLK(clk), .RST(rst), .Q(c[945]) );
  DFF \sreg_reg[944]  ( .D(c[946]), .CLK(clk), .RST(rst), .Q(c[944]) );
  DFF \sreg_reg[943]  ( .D(c[945]), .CLK(clk), .RST(rst), .Q(c[943]) );
  DFF \sreg_reg[942]  ( .D(c[944]), .CLK(clk), .RST(rst), .Q(c[942]) );
  DFF \sreg_reg[941]  ( .D(c[943]), .CLK(clk), .RST(rst), .Q(c[941]) );
  DFF \sreg_reg[940]  ( .D(c[942]), .CLK(clk), .RST(rst), .Q(c[940]) );
  DFF \sreg_reg[939]  ( .D(c[941]), .CLK(clk), .RST(rst), .Q(c[939]) );
  DFF \sreg_reg[938]  ( .D(c[940]), .CLK(clk), .RST(rst), .Q(c[938]) );
  DFF \sreg_reg[937]  ( .D(c[939]), .CLK(clk), .RST(rst), .Q(c[937]) );
  DFF \sreg_reg[936]  ( .D(c[938]), .CLK(clk), .RST(rst), .Q(c[936]) );
  DFF \sreg_reg[935]  ( .D(c[937]), .CLK(clk), .RST(rst), .Q(c[935]) );
  DFF \sreg_reg[934]  ( .D(c[936]), .CLK(clk), .RST(rst), .Q(c[934]) );
  DFF \sreg_reg[933]  ( .D(c[935]), .CLK(clk), .RST(rst), .Q(c[933]) );
  DFF \sreg_reg[932]  ( .D(c[934]), .CLK(clk), .RST(rst), .Q(c[932]) );
  DFF \sreg_reg[931]  ( .D(c[933]), .CLK(clk), .RST(rst), .Q(c[931]) );
  DFF \sreg_reg[930]  ( .D(c[932]), .CLK(clk), .RST(rst), .Q(c[930]) );
  DFF \sreg_reg[929]  ( .D(c[931]), .CLK(clk), .RST(rst), .Q(c[929]) );
  DFF \sreg_reg[928]  ( .D(c[930]), .CLK(clk), .RST(rst), .Q(c[928]) );
  DFF \sreg_reg[927]  ( .D(c[929]), .CLK(clk), .RST(rst), .Q(c[927]) );
  DFF \sreg_reg[926]  ( .D(c[928]), .CLK(clk), .RST(rst), .Q(c[926]) );
  DFF \sreg_reg[925]  ( .D(c[927]), .CLK(clk), .RST(rst), .Q(c[925]) );
  DFF \sreg_reg[924]  ( .D(c[926]), .CLK(clk), .RST(rst), .Q(c[924]) );
  DFF \sreg_reg[923]  ( .D(c[925]), .CLK(clk), .RST(rst), .Q(c[923]) );
  DFF \sreg_reg[922]  ( .D(c[924]), .CLK(clk), .RST(rst), .Q(c[922]) );
  DFF \sreg_reg[921]  ( .D(c[923]), .CLK(clk), .RST(rst), .Q(c[921]) );
  DFF \sreg_reg[920]  ( .D(c[922]), .CLK(clk), .RST(rst), .Q(c[920]) );
  DFF \sreg_reg[919]  ( .D(c[921]), .CLK(clk), .RST(rst), .Q(c[919]) );
  DFF \sreg_reg[918]  ( .D(c[920]), .CLK(clk), .RST(rst), .Q(c[918]) );
  DFF \sreg_reg[917]  ( .D(c[919]), .CLK(clk), .RST(rst), .Q(c[917]) );
  DFF \sreg_reg[916]  ( .D(c[918]), .CLK(clk), .RST(rst), .Q(c[916]) );
  DFF \sreg_reg[915]  ( .D(c[917]), .CLK(clk), .RST(rst), .Q(c[915]) );
  DFF \sreg_reg[914]  ( .D(c[916]), .CLK(clk), .RST(rst), .Q(c[914]) );
  DFF \sreg_reg[913]  ( .D(c[915]), .CLK(clk), .RST(rst), .Q(c[913]) );
  DFF \sreg_reg[912]  ( .D(c[914]), .CLK(clk), .RST(rst), .Q(c[912]) );
  DFF \sreg_reg[911]  ( .D(c[913]), .CLK(clk), .RST(rst), .Q(c[911]) );
  DFF \sreg_reg[910]  ( .D(c[912]), .CLK(clk), .RST(rst), .Q(c[910]) );
  DFF \sreg_reg[909]  ( .D(c[911]), .CLK(clk), .RST(rst), .Q(c[909]) );
  DFF \sreg_reg[908]  ( .D(c[910]), .CLK(clk), .RST(rst), .Q(c[908]) );
  DFF \sreg_reg[907]  ( .D(c[909]), .CLK(clk), .RST(rst), .Q(c[907]) );
  DFF \sreg_reg[906]  ( .D(c[908]), .CLK(clk), .RST(rst), .Q(c[906]) );
  DFF \sreg_reg[905]  ( .D(c[907]), .CLK(clk), .RST(rst), .Q(c[905]) );
  DFF \sreg_reg[904]  ( .D(c[906]), .CLK(clk), .RST(rst), .Q(c[904]) );
  DFF \sreg_reg[903]  ( .D(c[905]), .CLK(clk), .RST(rst), .Q(c[903]) );
  DFF \sreg_reg[902]  ( .D(c[904]), .CLK(clk), .RST(rst), .Q(c[902]) );
  DFF \sreg_reg[901]  ( .D(c[903]), .CLK(clk), .RST(rst), .Q(c[901]) );
  DFF \sreg_reg[900]  ( .D(c[902]), .CLK(clk), .RST(rst), .Q(c[900]) );
  DFF \sreg_reg[899]  ( .D(c[901]), .CLK(clk), .RST(rst), .Q(c[899]) );
  DFF \sreg_reg[898]  ( .D(c[900]), .CLK(clk), .RST(rst), .Q(c[898]) );
  DFF \sreg_reg[897]  ( .D(c[899]), .CLK(clk), .RST(rst), .Q(c[897]) );
  DFF \sreg_reg[896]  ( .D(c[898]), .CLK(clk), .RST(rst), .Q(c[896]) );
  DFF \sreg_reg[895]  ( .D(c[897]), .CLK(clk), .RST(rst), .Q(c[895]) );
  DFF \sreg_reg[894]  ( .D(c[896]), .CLK(clk), .RST(rst), .Q(c[894]) );
  DFF \sreg_reg[893]  ( .D(c[895]), .CLK(clk), .RST(rst), .Q(c[893]) );
  DFF \sreg_reg[892]  ( .D(c[894]), .CLK(clk), .RST(rst), .Q(c[892]) );
  DFF \sreg_reg[891]  ( .D(c[893]), .CLK(clk), .RST(rst), .Q(c[891]) );
  DFF \sreg_reg[890]  ( .D(c[892]), .CLK(clk), .RST(rst), .Q(c[890]) );
  DFF \sreg_reg[889]  ( .D(c[891]), .CLK(clk), .RST(rst), .Q(c[889]) );
  DFF \sreg_reg[888]  ( .D(c[890]), .CLK(clk), .RST(rst), .Q(c[888]) );
  DFF \sreg_reg[887]  ( .D(c[889]), .CLK(clk), .RST(rst), .Q(c[887]) );
  DFF \sreg_reg[886]  ( .D(c[888]), .CLK(clk), .RST(rst), .Q(c[886]) );
  DFF \sreg_reg[885]  ( .D(c[887]), .CLK(clk), .RST(rst), .Q(c[885]) );
  DFF \sreg_reg[884]  ( .D(c[886]), .CLK(clk), .RST(rst), .Q(c[884]) );
  DFF \sreg_reg[883]  ( .D(c[885]), .CLK(clk), .RST(rst), .Q(c[883]) );
  DFF \sreg_reg[882]  ( .D(c[884]), .CLK(clk), .RST(rst), .Q(c[882]) );
  DFF \sreg_reg[881]  ( .D(c[883]), .CLK(clk), .RST(rst), .Q(c[881]) );
  DFF \sreg_reg[880]  ( .D(c[882]), .CLK(clk), .RST(rst), .Q(c[880]) );
  DFF \sreg_reg[879]  ( .D(c[881]), .CLK(clk), .RST(rst), .Q(c[879]) );
  DFF \sreg_reg[878]  ( .D(c[880]), .CLK(clk), .RST(rst), .Q(c[878]) );
  DFF \sreg_reg[877]  ( .D(c[879]), .CLK(clk), .RST(rst), .Q(c[877]) );
  DFF \sreg_reg[876]  ( .D(c[878]), .CLK(clk), .RST(rst), .Q(c[876]) );
  DFF \sreg_reg[875]  ( .D(c[877]), .CLK(clk), .RST(rst), .Q(c[875]) );
  DFF \sreg_reg[874]  ( .D(c[876]), .CLK(clk), .RST(rst), .Q(c[874]) );
  DFF \sreg_reg[873]  ( .D(c[875]), .CLK(clk), .RST(rst), .Q(c[873]) );
  DFF \sreg_reg[872]  ( .D(c[874]), .CLK(clk), .RST(rst), .Q(c[872]) );
  DFF \sreg_reg[871]  ( .D(c[873]), .CLK(clk), .RST(rst), .Q(c[871]) );
  DFF \sreg_reg[870]  ( .D(c[872]), .CLK(clk), .RST(rst), .Q(c[870]) );
  DFF \sreg_reg[869]  ( .D(c[871]), .CLK(clk), .RST(rst), .Q(c[869]) );
  DFF \sreg_reg[868]  ( .D(c[870]), .CLK(clk), .RST(rst), .Q(c[868]) );
  DFF \sreg_reg[867]  ( .D(c[869]), .CLK(clk), .RST(rst), .Q(c[867]) );
  DFF \sreg_reg[866]  ( .D(c[868]), .CLK(clk), .RST(rst), .Q(c[866]) );
  DFF \sreg_reg[865]  ( .D(c[867]), .CLK(clk), .RST(rst), .Q(c[865]) );
  DFF \sreg_reg[864]  ( .D(c[866]), .CLK(clk), .RST(rst), .Q(c[864]) );
  DFF \sreg_reg[863]  ( .D(c[865]), .CLK(clk), .RST(rst), .Q(c[863]) );
  DFF \sreg_reg[862]  ( .D(c[864]), .CLK(clk), .RST(rst), .Q(c[862]) );
  DFF \sreg_reg[861]  ( .D(c[863]), .CLK(clk), .RST(rst), .Q(c[861]) );
  DFF \sreg_reg[860]  ( .D(c[862]), .CLK(clk), .RST(rst), .Q(c[860]) );
  DFF \sreg_reg[859]  ( .D(c[861]), .CLK(clk), .RST(rst), .Q(c[859]) );
  DFF \sreg_reg[858]  ( .D(c[860]), .CLK(clk), .RST(rst), .Q(c[858]) );
  DFF \sreg_reg[857]  ( .D(c[859]), .CLK(clk), .RST(rst), .Q(c[857]) );
  DFF \sreg_reg[856]  ( .D(c[858]), .CLK(clk), .RST(rst), .Q(c[856]) );
  DFF \sreg_reg[855]  ( .D(c[857]), .CLK(clk), .RST(rst), .Q(c[855]) );
  DFF \sreg_reg[854]  ( .D(c[856]), .CLK(clk), .RST(rst), .Q(c[854]) );
  DFF \sreg_reg[853]  ( .D(c[855]), .CLK(clk), .RST(rst), .Q(c[853]) );
  DFF \sreg_reg[852]  ( .D(c[854]), .CLK(clk), .RST(rst), .Q(c[852]) );
  DFF \sreg_reg[851]  ( .D(c[853]), .CLK(clk), .RST(rst), .Q(c[851]) );
  DFF \sreg_reg[850]  ( .D(c[852]), .CLK(clk), .RST(rst), .Q(c[850]) );
  DFF \sreg_reg[849]  ( .D(c[851]), .CLK(clk), .RST(rst), .Q(c[849]) );
  DFF \sreg_reg[848]  ( .D(c[850]), .CLK(clk), .RST(rst), .Q(c[848]) );
  DFF \sreg_reg[847]  ( .D(c[849]), .CLK(clk), .RST(rst), .Q(c[847]) );
  DFF \sreg_reg[846]  ( .D(c[848]), .CLK(clk), .RST(rst), .Q(c[846]) );
  DFF \sreg_reg[845]  ( .D(c[847]), .CLK(clk), .RST(rst), .Q(c[845]) );
  DFF \sreg_reg[844]  ( .D(c[846]), .CLK(clk), .RST(rst), .Q(c[844]) );
  DFF \sreg_reg[843]  ( .D(c[845]), .CLK(clk), .RST(rst), .Q(c[843]) );
  DFF \sreg_reg[842]  ( .D(c[844]), .CLK(clk), .RST(rst), .Q(c[842]) );
  DFF \sreg_reg[841]  ( .D(c[843]), .CLK(clk), .RST(rst), .Q(c[841]) );
  DFF \sreg_reg[840]  ( .D(c[842]), .CLK(clk), .RST(rst), .Q(c[840]) );
  DFF \sreg_reg[839]  ( .D(c[841]), .CLK(clk), .RST(rst), .Q(c[839]) );
  DFF \sreg_reg[838]  ( .D(c[840]), .CLK(clk), .RST(rst), .Q(c[838]) );
  DFF \sreg_reg[837]  ( .D(c[839]), .CLK(clk), .RST(rst), .Q(c[837]) );
  DFF \sreg_reg[836]  ( .D(c[838]), .CLK(clk), .RST(rst), .Q(c[836]) );
  DFF \sreg_reg[835]  ( .D(c[837]), .CLK(clk), .RST(rst), .Q(c[835]) );
  DFF \sreg_reg[834]  ( .D(c[836]), .CLK(clk), .RST(rst), .Q(c[834]) );
  DFF \sreg_reg[833]  ( .D(c[835]), .CLK(clk), .RST(rst), .Q(c[833]) );
  DFF \sreg_reg[832]  ( .D(c[834]), .CLK(clk), .RST(rst), .Q(c[832]) );
  DFF \sreg_reg[831]  ( .D(c[833]), .CLK(clk), .RST(rst), .Q(c[831]) );
  DFF \sreg_reg[830]  ( .D(c[832]), .CLK(clk), .RST(rst), .Q(c[830]) );
  DFF \sreg_reg[829]  ( .D(c[831]), .CLK(clk), .RST(rst), .Q(c[829]) );
  DFF \sreg_reg[828]  ( .D(c[830]), .CLK(clk), .RST(rst), .Q(c[828]) );
  DFF \sreg_reg[827]  ( .D(c[829]), .CLK(clk), .RST(rst), .Q(c[827]) );
  DFF \sreg_reg[826]  ( .D(c[828]), .CLK(clk), .RST(rst), .Q(c[826]) );
  DFF \sreg_reg[825]  ( .D(c[827]), .CLK(clk), .RST(rst), .Q(c[825]) );
  DFF \sreg_reg[824]  ( .D(c[826]), .CLK(clk), .RST(rst), .Q(c[824]) );
  DFF \sreg_reg[823]  ( .D(c[825]), .CLK(clk), .RST(rst), .Q(c[823]) );
  DFF \sreg_reg[822]  ( .D(c[824]), .CLK(clk), .RST(rst), .Q(c[822]) );
  DFF \sreg_reg[821]  ( .D(c[823]), .CLK(clk), .RST(rst), .Q(c[821]) );
  DFF \sreg_reg[820]  ( .D(c[822]), .CLK(clk), .RST(rst), .Q(c[820]) );
  DFF \sreg_reg[819]  ( .D(c[821]), .CLK(clk), .RST(rst), .Q(c[819]) );
  DFF \sreg_reg[818]  ( .D(c[820]), .CLK(clk), .RST(rst), .Q(c[818]) );
  DFF \sreg_reg[817]  ( .D(c[819]), .CLK(clk), .RST(rst), .Q(c[817]) );
  DFF \sreg_reg[816]  ( .D(c[818]), .CLK(clk), .RST(rst), .Q(c[816]) );
  DFF \sreg_reg[815]  ( .D(c[817]), .CLK(clk), .RST(rst), .Q(c[815]) );
  DFF \sreg_reg[814]  ( .D(c[816]), .CLK(clk), .RST(rst), .Q(c[814]) );
  DFF \sreg_reg[813]  ( .D(c[815]), .CLK(clk), .RST(rst), .Q(c[813]) );
  DFF \sreg_reg[812]  ( .D(c[814]), .CLK(clk), .RST(rst), .Q(c[812]) );
  DFF \sreg_reg[811]  ( .D(c[813]), .CLK(clk), .RST(rst), .Q(c[811]) );
  DFF \sreg_reg[810]  ( .D(c[812]), .CLK(clk), .RST(rst), .Q(c[810]) );
  DFF \sreg_reg[809]  ( .D(c[811]), .CLK(clk), .RST(rst), .Q(c[809]) );
  DFF \sreg_reg[808]  ( .D(c[810]), .CLK(clk), .RST(rst), .Q(c[808]) );
  DFF \sreg_reg[807]  ( .D(c[809]), .CLK(clk), .RST(rst), .Q(c[807]) );
  DFF \sreg_reg[806]  ( .D(c[808]), .CLK(clk), .RST(rst), .Q(c[806]) );
  DFF \sreg_reg[805]  ( .D(c[807]), .CLK(clk), .RST(rst), .Q(c[805]) );
  DFF \sreg_reg[804]  ( .D(c[806]), .CLK(clk), .RST(rst), .Q(c[804]) );
  DFF \sreg_reg[803]  ( .D(c[805]), .CLK(clk), .RST(rst), .Q(c[803]) );
  DFF \sreg_reg[802]  ( .D(c[804]), .CLK(clk), .RST(rst), .Q(c[802]) );
  DFF \sreg_reg[801]  ( .D(c[803]), .CLK(clk), .RST(rst), .Q(c[801]) );
  DFF \sreg_reg[800]  ( .D(c[802]), .CLK(clk), .RST(rst), .Q(c[800]) );
  DFF \sreg_reg[799]  ( .D(c[801]), .CLK(clk), .RST(rst), .Q(c[799]) );
  DFF \sreg_reg[798]  ( .D(c[800]), .CLK(clk), .RST(rst), .Q(c[798]) );
  DFF \sreg_reg[797]  ( .D(c[799]), .CLK(clk), .RST(rst), .Q(c[797]) );
  DFF \sreg_reg[796]  ( .D(c[798]), .CLK(clk), .RST(rst), .Q(c[796]) );
  DFF \sreg_reg[795]  ( .D(c[797]), .CLK(clk), .RST(rst), .Q(c[795]) );
  DFF \sreg_reg[794]  ( .D(c[796]), .CLK(clk), .RST(rst), .Q(c[794]) );
  DFF \sreg_reg[793]  ( .D(c[795]), .CLK(clk), .RST(rst), .Q(c[793]) );
  DFF \sreg_reg[792]  ( .D(c[794]), .CLK(clk), .RST(rst), .Q(c[792]) );
  DFF \sreg_reg[791]  ( .D(c[793]), .CLK(clk), .RST(rst), .Q(c[791]) );
  DFF \sreg_reg[790]  ( .D(c[792]), .CLK(clk), .RST(rst), .Q(c[790]) );
  DFF \sreg_reg[789]  ( .D(c[791]), .CLK(clk), .RST(rst), .Q(c[789]) );
  DFF \sreg_reg[788]  ( .D(c[790]), .CLK(clk), .RST(rst), .Q(c[788]) );
  DFF \sreg_reg[787]  ( .D(c[789]), .CLK(clk), .RST(rst), .Q(c[787]) );
  DFF \sreg_reg[786]  ( .D(c[788]), .CLK(clk), .RST(rst), .Q(c[786]) );
  DFF \sreg_reg[785]  ( .D(c[787]), .CLK(clk), .RST(rst), .Q(c[785]) );
  DFF \sreg_reg[784]  ( .D(c[786]), .CLK(clk), .RST(rst), .Q(c[784]) );
  DFF \sreg_reg[783]  ( .D(c[785]), .CLK(clk), .RST(rst), .Q(c[783]) );
  DFF \sreg_reg[782]  ( .D(c[784]), .CLK(clk), .RST(rst), .Q(c[782]) );
  DFF \sreg_reg[781]  ( .D(c[783]), .CLK(clk), .RST(rst), .Q(c[781]) );
  DFF \sreg_reg[780]  ( .D(c[782]), .CLK(clk), .RST(rst), .Q(c[780]) );
  DFF \sreg_reg[779]  ( .D(c[781]), .CLK(clk), .RST(rst), .Q(c[779]) );
  DFF \sreg_reg[778]  ( .D(c[780]), .CLK(clk), .RST(rst), .Q(c[778]) );
  DFF \sreg_reg[777]  ( .D(c[779]), .CLK(clk), .RST(rst), .Q(c[777]) );
  DFF \sreg_reg[776]  ( .D(c[778]), .CLK(clk), .RST(rst), .Q(c[776]) );
  DFF \sreg_reg[775]  ( .D(c[777]), .CLK(clk), .RST(rst), .Q(c[775]) );
  DFF \sreg_reg[774]  ( .D(c[776]), .CLK(clk), .RST(rst), .Q(c[774]) );
  DFF \sreg_reg[773]  ( .D(c[775]), .CLK(clk), .RST(rst), .Q(c[773]) );
  DFF \sreg_reg[772]  ( .D(c[774]), .CLK(clk), .RST(rst), .Q(c[772]) );
  DFF \sreg_reg[771]  ( .D(c[773]), .CLK(clk), .RST(rst), .Q(c[771]) );
  DFF \sreg_reg[770]  ( .D(c[772]), .CLK(clk), .RST(rst), .Q(c[770]) );
  DFF \sreg_reg[769]  ( .D(c[771]), .CLK(clk), .RST(rst), .Q(c[769]) );
  DFF \sreg_reg[768]  ( .D(c[770]), .CLK(clk), .RST(rst), .Q(c[768]) );
  DFF \sreg_reg[767]  ( .D(c[769]), .CLK(clk), .RST(rst), .Q(c[767]) );
  DFF \sreg_reg[766]  ( .D(c[768]), .CLK(clk), .RST(rst), .Q(c[766]) );
  DFF \sreg_reg[765]  ( .D(c[767]), .CLK(clk), .RST(rst), .Q(c[765]) );
  DFF \sreg_reg[764]  ( .D(c[766]), .CLK(clk), .RST(rst), .Q(c[764]) );
  DFF \sreg_reg[763]  ( .D(c[765]), .CLK(clk), .RST(rst), .Q(c[763]) );
  DFF \sreg_reg[762]  ( .D(c[764]), .CLK(clk), .RST(rst), .Q(c[762]) );
  DFF \sreg_reg[761]  ( .D(c[763]), .CLK(clk), .RST(rst), .Q(c[761]) );
  DFF \sreg_reg[760]  ( .D(c[762]), .CLK(clk), .RST(rst), .Q(c[760]) );
  DFF \sreg_reg[759]  ( .D(c[761]), .CLK(clk), .RST(rst), .Q(c[759]) );
  DFF \sreg_reg[758]  ( .D(c[760]), .CLK(clk), .RST(rst), .Q(c[758]) );
  DFF \sreg_reg[757]  ( .D(c[759]), .CLK(clk), .RST(rst), .Q(c[757]) );
  DFF \sreg_reg[756]  ( .D(c[758]), .CLK(clk), .RST(rst), .Q(c[756]) );
  DFF \sreg_reg[755]  ( .D(c[757]), .CLK(clk), .RST(rst), .Q(c[755]) );
  DFF \sreg_reg[754]  ( .D(c[756]), .CLK(clk), .RST(rst), .Q(c[754]) );
  DFF \sreg_reg[753]  ( .D(c[755]), .CLK(clk), .RST(rst), .Q(c[753]) );
  DFF \sreg_reg[752]  ( .D(c[754]), .CLK(clk), .RST(rst), .Q(c[752]) );
  DFF \sreg_reg[751]  ( .D(c[753]), .CLK(clk), .RST(rst), .Q(c[751]) );
  DFF \sreg_reg[750]  ( .D(c[752]), .CLK(clk), .RST(rst), .Q(c[750]) );
  DFF \sreg_reg[749]  ( .D(c[751]), .CLK(clk), .RST(rst), .Q(c[749]) );
  DFF \sreg_reg[748]  ( .D(c[750]), .CLK(clk), .RST(rst), .Q(c[748]) );
  DFF \sreg_reg[747]  ( .D(c[749]), .CLK(clk), .RST(rst), .Q(c[747]) );
  DFF \sreg_reg[746]  ( .D(c[748]), .CLK(clk), .RST(rst), .Q(c[746]) );
  DFF \sreg_reg[745]  ( .D(c[747]), .CLK(clk), .RST(rst), .Q(c[745]) );
  DFF \sreg_reg[744]  ( .D(c[746]), .CLK(clk), .RST(rst), .Q(c[744]) );
  DFF \sreg_reg[743]  ( .D(c[745]), .CLK(clk), .RST(rst), .Q(c[743]) );
  DFF \sreg_reg[742]  ( .D(c[744]), .CLK(clk), .RST(rst), .Q(c[742]) );
  DFF \sreg_reg[741]  ( .D(c[743]), .CLK(clk), .RST(rst), .Q(c[741]) );
  DFF \sreg_reg[740]  ( .D(c[742]), .CLK(clk), .RST(rst), .Q(c[740]) );
  DFF \sreg_reg[739]  ( .D(c[741]), .CLK(clk), .RST(rst), .Q(c[739]) );
  DFF \sreg_reg[738]  ( .D(c[740]), .CLK(clk), .RST(rst), .Q(c[738]) );
  DFF \sreg_reg[737]  ( .D(c[739]), .CLK(clk), .RST(rst), .Q(c[737]) );
  DFF \sreg_reg[736]  ( .D(c[738]), .CLK(clk), .RST(rst), .Q(c[736]) );
  DFF \sreg_reg[735]  ( .D(c[737]), .CLK(clk), .RST(rst), .Q(c[735]) );
  DFF \sreg_reg[734]  ( .D(c[736]), .CLK(clk), .RST(rst), .Q(c[734]) );
  DFF \sreg_reg[733]  ( .D(c[735]), .CLK(clk), .RST(rst), .Q(c[733]) );
  DFF \sreg_reg[732]  ( .D(c[734]), .CLK(clk), .RST(rst), .Q(c[732]) );
  DFF \sreg_reg[731]  ( .D(c[733]), .CLK(clk), .RST(rst), .Q(c[731]) );
  DFF \sreg_reg[730]  ( .D(c[732]), .CLK(clk), .RST(rst), .Q(c[730]) );
  DFF \sreg_reg[729]  ( .D(c[731]), .CLK(clk), .RST(rst), .Q(c[729]) );
  DFF \sreg_reg[728]  ( .D(c[730]), .CLK(clk), .RST(rst), .Q(c[728]) );
  DFF \sreg_reg[727]  ( .D(c[729]), .CLK(clk), .RST(rst), .Q(c[727]) );
  DFF \sreg_reg[726]  ( .D(c[728]), .CLK(clk), .RST(rst), .Q(c[726]) );
  DFF \sreg_reg[725]  ( .D(c[727]), .CLK(clk), .RST(rst), .Q(c[725]) );
  DFF \sreg_reg[724]  ( .D(c[726]), .CLK(clk), .RST(rst), .Q(c[724]) );
  DFF \sreg_reg[723]  ( .D(c[725]), .CLK(clk), .RST(rst), .Q(c[723]) );
  DFF \sreg_reg[722]  ( .D(c[724]), .CLK(clk), .RST(rst), .Q(c[722]) );
  DFF \sreg_reg[721]  ( .D(c[723]), .CLK(clk), .RST(rst), .Q(c[721]) );
  DFF \sreg_reg[720]  ( .D(c[722]), .CLK(clk), .RST(rst), .Q(c[720]) );
  DFF \sreg_reg[719]  ( .D(c[721]), .CLK(clk), .RST(rst), .Q(c[719]) );
  DFF \sreg_reg[718]  ( .D(c[720]), .CLK(clk), .RST(rst), .Q(c[718]) );
  DFF \sreg_reg[717]  ( .D(c[719]), .CLK(clk), .RST(rst), .Q(c[717]) );
  DFF \sreg_reg[716]  ( .D(c[718]), .CLK(clk), .RST(rst), .Q(c[716]) );
  DFF \sreg_reg[715]  ( .D(c[717]), .CLK(clk), .RST(rst), .Q(c[715]) );
  DFF \sreg_reg[714]  ( .D(c[716]), .CLK(clk), .RST(rst), .Q(c[714]) );
  DFF \sreg_reg[713]  ( .D(c[715]), .CLK(clk), .RST(rst), .Q(c[713]) );
  DFF \sreg_reg[712]  ( .D(c[714]), .CLK(clk), .RST(rst), .Q(c[712]) );
  DFF \sreg_reg[711]  ( .D(c[713]), .CLK(clk), .RST(rst), .Q(c[711]) );
  DFF \sreg_reg[710]  ( .D(c[712]), .CLK(clk), .RST(rst), .Q(c[710]) );
  DFF \sreg_reg[709]  ( .D(c[711]), .CLK(clk), .RST(rst), .Q(c[709]) );
  DFF \sreg_reg[708]  ( .D(c[710]), .CLK(clk), .RST(rst), .Q(c[708]) );
  DFF \sreg_reg[707]  ( .D(c[709]), .CLK(clk), .RST(rst), .Q(c[707]) );
  DFF \sreg_reg[706]  ( .D(c[708]), .CLK(clk), .RST(rst), .Q(c[706]) );
  DFF \sreg_reg[705]  ( .D(c[707]), .CLK(clk), .RST(rst), .Q(c[705]) );
  DFF \sreg_reg[704]  ( .D(c[706]), .CLK(clk), .RST(rst), .Q(c[704]) );
  DFF \sreg_reg[703]  ( .D(c[705]), .CLK(clk), .RST(rst), .Q(c[703]) );
  DFF \sreg_reg[702]  ( .D(c[704]), .CLK(clk), .RST(rst), .Q(c[702]) );
  DFF \sreg_reg[701]  ( .D(c[703]), .CLK(clk), .RST(rst), .Q(c[701]) );
  DFF \sreg_reg[700]  ( .D(c[702]), .CLK(clk), .RST(rst), .Q(c[700]) );
  DFF \sreg_reg[699]  ( .D(c[701]), .CLK(clk), .RST(rst), .Q(c[699]) );
  DFF \sreg_reg[698]  ( .D(c[700]), .CLK(clk), .RST(rst), .Q(c[698]) );
  DFF \sreg_reg[697]  ( .D(c[699]), .CLK(clk), .RST(rst), .Q(c[697]) );
  DFF \sreg_reg[696]  ( .D(c[698]), .CLK(clk), .RST(rst), .Q(c[696]) );
  DFF \sreg_reg[695]  ( .D(c[697]), .CLK(clk), .RST(rst), .Q(c[695]) );
  DFF \sreg_reg[694]  ( .D(c[696]), .CLK(clk), .RST(rst), .Q(c[694]) );
  DFF \sreg_reg[693]  ( .D(c[695]), .CLK(clk), .RST(rst), .Q(c[693]) );
  DFF \sreg_reg[692]  ( .D(c[694]), .CLK(clk), .RST(rst), .Q(c[692]) );
  DFF \sreg_reg[691]  ( .D(c[693]), .CLK(clk), .RST(rst), .Q(c[691]) );
  DFF \sreg_reg[690]  ( .D(c[692]), .CLK(clk), .RST(rst), .Q(c[690]) );
  DFF \sreg_reg[689]  ( .D(c[691]), .CLK(clk), .RST(rst), .Q(c[689]) );
  DFF \sreg_reg[688]  ( .D(c[690]), .CLK(clk), .RST(rst), .Q(c[688]) );
  DFF \sreg_reg[687]  ( .D(c[689]), .CLK(clk), .RST(rst), .Q(c[687]) );
  DFF \sreg_reg[686]  ( .D(c[688]), .CLK(clk), .RST(rst), .Q(c[686]) );
  DFF \sreg_reg[685]  ( .D(c[687]), .CLK(clk), .RST(rst), .Q(c[685]) );
  DFF \sreg_reg[684]  ( .D(c[686]), .CLK(clk), .RST(rst), .Q(c[684]) );
  DFF \sreg_reg[683]  ( .D(c[685]), .CLK(clk), .RST(rst), .Q(c[683]) );
  DFF \sreg_reg[682]  ( .D(c[684]), .CLK(clk), .RST(rst), .Q(c[682]) );
  DFF \sreg_reg[681]  ( .D(c[683]), .CLK(clk), .RST(rst), .Q(c[681]) );
  DFF \sreg_reg[680]  ( .D(c[682]), .CLK(clk), .RST(rst), .Q(c[680]) );
  DFF \sreg_reg[679]  ( .D(c[681]), .CLK(clk), .RST(rst), .Q(c[679]) );
  DFF \sreg_reg[678]  ( .D(c[680]), .CLK(clk), .RST(rst), .Q(c[678]) );
  DFF \sreg_reg[677]  ( .D(c[679]), .CLK(clk), .RST(rst), .Q(c[677]) );
  DFF \sreg_reg[676]  ( .D(c[678]), .CLK(clk), .RST(rst), .Q(c[676]) );
  DFF \sreg_reg[675]  ( .D(c[677]), .CLK(clk), .RST(rst), .Q(c[675]) );
  DFF \sreg_reg[674]  ( .D(c[676]), .CLK(clk), .RST(rst), .Q(c[674]) );
  DFF \sreg_reg[673]  ( .D(c[675]), .CLK(clk), .RST(rst), .Q(c[673]) );
  DFF \sreg_reg[672]  ( .D(c[674]), .CLK(clk), .RST(rst), .Q(c[672]) );
  DFF \sreg_reg[671]  ( .D(c[673]), .CLK(clk), .RST(rst), .Q(c[671]) );
  DFF \sreg_reg[670]  ( .D(c[672]), .CLK(clk), .RST(rst), .Q(c[670]) );
  DFF \sreg_reg[669]  ( .D(c[671]), .CLK(clk), .RST(rst), .Q(c[669]) );
  DFF \sreg_reg[668]  ( .D(c[670]), .CLK(clk), .RST(rst), .Q(c[668]) );
  DFF \sreg_reg[667]  ( .D(c[669]), .CLK(clk), .RST(rst), .Q(c[667]) );
  DFF \sreg_reg[666]  ( .D(c[668]), .CLK(clk), .RST(rst), .Q(c[666]) );
  DFF \sreg_reg[665]  ( .D(c[667]), .CLK(clk), .RST(rst), .Q(c[665]) );
  DFF \sreg_reg[664]  ( .D(c[666]), .CLK(clk), .RST(rst), .Q(c[664]) );
  DFF \sreg_reg[663]  ( .D(c[665]), .CLK(clk), .RST(rst), .Q(c[663]) );
  DFF \sreg_reg[662]  ( .D(c[664]), .CLK(clk), .RST(rst), .Q(c[662]) );
  DFF \sreg_reg[661]  ( .D(c[663]), .CLK(clk), .RST(rst), .Q(c[661]) );
  DFF \sreg_reg[660]  ( .D(c[662]), .CLK(clk), .RST(rst), .Q(c[660]) );
  DFF \sreg_reg[659]  ( .D(c[661]), .CLK(clk), .RST(rst), .Q(c[659]) );
  DFF \sreg_reg[658]  ( .D(c[660]), .CLK(clk), .RST(rst), .Q(c[658]) );
  DFF \sreg_reg[657]  ( .D(c[659]), .CLK(clk), .RST(rst), .Q(c[657]) );
  DFF \sreg_reg[656]  ( .D(c[658]), .CLK(clk), .RST(rst), .Q(c[656]) );
  DFF \sreg_reg[655]  ( .D(c[657]), .CLK(clk), .RST(rst), .Q(c[655]) );
  DFF \sreg_reg[654]  ( .D(c[656]), .CLK(clk), .RST(rst), .Q(c[654]) );
  DFF \sreg_reg[653]  ( .D(c[655]), .CLK(clk), .RST(rst), .Q(c[653]) );
  DFF \sreg_reg[652]  ( .D(c[654]), .CLK(clk), .RST(rst), .Q(c[652]) );
  DFF \sreg_reg[651]  ( .D(c[653]), .CLK(clk), .RST(rst), .Q(c[651]) );
  DFF \sreg_reg[650]  ( .D(c[652]), .CLK(clk), .RST(rst), .Q(c[650]) );
  DFF \sreg_reg[649]  ( .D(c[651]), .CLK(clk), .RST(rst), .Q(c[649]) );
  DFF \sreg_reg[648]  ( .D(c[650]), .CLK(clk), .RST(rst), .Q(c[648]) );
  DFF \sreg_reg[647]  ( .D(c[649]), .CLK(clk), .RST(rst), .Q(c[647]) );
  DFF \sreg_reg[646]  ( .D(c[648]), .CLK(clk), .RST(rst), .Q(c[646]) );
  DFF \sreg_reg[645]  ( .D(c[647]), .CLK(clk), .RST(rst), .Q(c[645]) );
  DFF \sreg_reg[644]  ( .D(c[646]), .CLK(clk), .RST(rst), .Q(c[644]) );
  DFF \sreg_reg[643]  ( .D(c[645]), .CLK(clk), .RST(rst), .Q(c[643]) );
  DFF \sreg_reg[642]  ( .D(c[644]), .CLK(clk), .RST(rst), .Q(c[642]) );
  DFF \sreg_reg[641]  ( .D(c[643]), .CLK(clk), .RST(rst), .Q(c[641]) );
  DFF \sreg_reg[640]  ( .D(c[642]), .CLK(clk), .RST(rst), .Q(c[640]) );
  DFF \sreg_reg[639]  ( .D(c[641]), .CLK(clk), .RST(rst), .Q(c[639]) );
  DFF \sreg_reg[638]  ( .D(c[640]), .CLK(clk), .RST(rst), .Q(c[638]) );
  DFF \sreg_reg[637]  ( .D(c[639]), .CLK(clk), .RST(rst), .Q(c[637]) );
  DFF \sreg_reg[636]  ( .D(c[638]), .CLK(clk), .RST(rst), .Q(c[636]) );
  DFF \sreg_reg[635]  ( .D(c[637]), .CLK(clk), .RST(rst), .Q(c[635]) );
  DFF \sreg_reg[634]  ( .D(c[636]), .CLK(clk), .RST(rst), .Q(c[634]) );
  DFF \sreg_reg[633]  ( .D(c[635]), .CLK(clk), .RST(rst), .Q(c[633]) );
  DFF \sreg_reg[632]  ( .D(c[634]), .CLK(clk), .RST(rst), .Q(c[632]) );
  DFF \sreg_reg[631]  ( .D(c[633]), .CLK(clk), .RST(rst), .Q(c[631]) );
  DFF \sreg_reg[630]  ( .D(c[632]), .CLK(clk), .RST(rst), .Q(c[630]) );
  DFF \sreg_reg[629]  ( .D(c[631]), .CLK(clk), .RST(rst), .Q(c[629]) );
  DFF \sreg_reg[628]  ( .D(c[630]), .CLK(clk), .RST(rst), .Q(c[628]) );
  DFF \sreg_reg[627]  ( .D(c[629]), .CLK(clk), .RST(rst), .Q(c[627]) );
  DFF \sreg_reg[626]  ( .D(c[628]), .CLK(clk), .RST(rst), .Q(c[626]) );
  DFF \sreg_reg[625]  ( .D(c[627]), .CLK(clk), .RST(rst), .Q(c[625]) );
  DFF \sreg_reg[624]  ( .D(c[626]), .CLK(clk), .RST(rst), .Q(c[624]) );
  DFF \sreg_reg[623]  ( .D(c[625]), .CLK(clk), .RST(rst), .Q(c[623]) );
  DFF \sreg_reg[622]  ( .D(c[624]), .CLK(clk), .RST(rst), .Q(c[622]) );
  DFF \sreg_reg[621]  ( .D(c[623]), .CLK(clk), .RST(rst), .Q(c[621]) );
  DFF \sreg_reg[620]  ( .D(c[622]), .CLK(clk), .RST(rst), .Q(c[620]) );
  DFF \sreg_reg[619]  ( .D(c[621]), .CLK(clk), .RST(rst), .Q(c[619]) );
  DFF \sreg_reg[618]  ( .D(c[620]), .CLK(clk), .RST(rst), .Q(c[618]) );
  DFF \sreg_reg[617]  ( .D(c[619]), .CLK(clk), .RST(rst), .Q(c[617]) );
  DFF \sreg_reg[616]  ( .D(c[618]), .CLK(clk), .RST(rst), .Q(c[616]) );
  DFF \sreg_reg[615]  ( .D(c[617]), .CLK(clk), .RST(rst), .Q(c[615]) );
  DFF \sreg_reg[614]  ( .D(c[616]), .CLK(clk), .RST(rst), .Q(c[614]) );
  DFF \sreg_reg[613]  ( .D(c[615]), .CLK(clk), .RST(rst), .Q(c[613]) );
  DFF \sreg_reg[612]  ( .D(c[614]), .CLK(clk), .RST(rst), .Q(c[612]) );
  DFF \sreg_reg[611]  ( .D(c[613]), .CLK(clk), .RST(rst), .Q(c[611]) );
  DFF \sreg_reg[610]  ( .D(c[612]), .CLK(clk), .RST(rst), .Q(c[610]) );
  DFF \sreg_reg[609]  ( .D(c[611]), .CLK(clk), .RST(rst), .Q(c[609]) );
  DFF \sreg_reg[608]  ( .D(c[610]), .CLK(clk), .RST(rst), .Q(c[608]) );
  DFF \sreg_reg[607]  ( .D(c[609]), .CLK(clk), .RST(rst), .Q(c[607]) );
  DFF \sreg_reg[606]  ( .D(c[608]), .CLK(clk), .RST(rst), .Q(c[606]) );
  DFF \sreg_reg[605]  ( .D(c[607]), .CLK(clk), .RST(rst), .Q(c[605]) );
  DFF \sreg_reg[604]  ( .D(c[606]), .CLK(clk), .RST(rst), .Q(c[604]) );
  DFF \sreg_reg[603]  ( .D(c[605]), .CLK(clk), .RST(rst), .Q(c[603]) );
  DFF \sreg_reg[602]  ( .D(c[604]), .CLK(clk), .RST(rst), .Q(c[602]) );
  DFF \sreg_reg[601]  ( .D(c[603]), .CLK(clk), .RST(rst), .Q(c[601]) );
  DFF \sreg_reg[600]  ( .D(c[602]), .CLK(clk), .RST(rst), .Q(c[600]) );
  DFF \sreg_reg[599]  ( .D(c[601]), .CLK(clk), .RST(rst), .Q(c[599]) );
  DFF \sreg_reg[598]  ( .D(c[600]), .CLK(clk), .RST(rst), .Q(c[598]) );
  DFF \sreg_reg[597]  ( .D(c[599]), .CLK(clk), .RST(rst), .Q(c[597]) );
  DFF \sreg_reg[596]  ( .D(c[598]), .CLK(clk), .RST(rst), .Q(c[596]) );
  DFF \sreg_reg[595]  ( .D(c[597]), .CLK(clk), .RST(rst), .Q(c[595]) );
  DFF \sreg_reg[594]  ( .D(c[596]), .CLK(clk), .RST(rst), .Q(c[594]) );
  DFF \sreg_reg[593]  ( .D(c[595]), .CLK(clk), .RST(rst), .Q(c[593]) );
  DFF \sreg_reg[592]  ( .D(c[594]), .CLK(clk), .RST(rst), .Q(c[592]) );
  DFF \sreg_reg[591]  ( .D(c[593]), .CLK(clk), .RST(rst), .Q(c[591]) );
  DFF \sreg_reg[590]  ( .D(c[592]), .CLK(clk), .RST(rst), .Q(c[590]) );
  DFF \sreg_reg[589]  ( .D(c[591]), .CLK(clk), .RST(rst), .Q(c[589]) );
  DFF \sreg_reg[588]  ( .D(c[590]), .CLK(clk), .RST(rst), .Q(c[588]) );
  DFF \sreg_reg[587]  ( .D(c[589]), .CLK(clk), .RST(rst), .Q(c[587]) );
  DFF \sreg_reg[586]  ( .D(c[588]), .CLK(clk), .RST(rst), .Q(c[586]) );
  DFF \sreg_reg[585]  ( .D(c[587]), .CLK(clk), .RST(rst), .Q(c[585]) );
  DFF \sreg_reg[584]  ( .D(c[586]), .CLK(clk), .RST(rst), .Q(c[584]) );
  DFF \sreg_reg[583]  ( .D(c[585]), .CLK(clk), .RST(rst), .Q(c[583]) );
  DFF \sreg_reg[582]  ( .D(c[584]), .CLK(clk), .RST(rst), .Q(c[582]) );
  DFF \sreg_reg[581]  ( .D(c[583]), .CLK(clk), .RST(rst), .Q(c[581]) );
  DFF \sreg_reg[580]  ( .D(c[582]), .CLK(clk), .RST(rst), .Q(c[580]) );
  DFF \sreg_reg[579]  ( .D(c[581]), .CLK(clk), .RST(rst), .Q(c[579]) );
  DFF \sreg_reg[578]  ( .D(c[580]), .CLK(clk), .RST(rst), .Q(c[578]) );
  DFF \sreg_reg[577]  ( .D(c[579]), .CLK(clk), .RST(rst), .Q(c[577]) );
  DFF \sreg_reg[576]  ( .D(c[578]), .CLK(clk), .RST(rst), .Q(c[576]) );
  DFF \sreg_reg[575]  ( .D(c[577]), .CLK(clk), .RST(rst), .Q(c[575]) );
  DFF \sreg_reg[574]  ( .D(c[576]), .CLK(clk), .RST(rst), .Q(c[574]) );
  DFF \sreg_reg[573]  ( .D(c[575]), .CLK(clk), .RST(rst), .Q(c[573]) );
  DFF \sreg_reg[572]  ( .D(c[574]), .CLK(clk), .RST(rst), .Q(c[572]) );
  DFF \sreg_reg[571]  ( .D(c[573]), .CLK(clk), .RST(rst), .Q(c[571]) );
  DFF \sreg_reg[570]  ( .D(c[572]), .CLK(clk), .RST(rst), .Q(c[570]) );
  DFF \sreg_reg[569]  ( .D(c[571]), .CLK(clk), .RST(rst), .Q(c[569]) );
  DFF \sreg_reg[568]  ( .D(c[570]), .CLK(clk), .RST(rst), .Q(c[568]) );
  DFF \sreg_reg[567]  ( .D(c[569]), .CLK(clk), .RST(rst), .Q(c[567]) );
  DFF \sreg_reg[566]  ( .D(c[568]), .CLK(clk), .RST(rst), .Q(c[566]) );
  DFF \sreg_reg[565]  ( .D(c[567]), .CLK(clk), .RST(rst), .Q(c[565]) );
  DFF \sreg_reg[564]  ( .D(c[566]), .CLK(clk), .RST(rst), .Q(c[564]) );
  DFF \sreg_reg[563]  ( .D(c[565]), .CLK(clk), .RST(rst), .Q(c[563]) );
  DFF \sreg_reg[562]  ( .D(c[564]), .CLK(clk), .RST(rst), .Q(c[562]) );
  DFF \sreg_reg[561]  ( .D(c[563]), .CLK(clk), .RST(rst), .Q(c[561]) );
  DFF \sreg_reg[560]  ( .D(c[562]), .CLK(clk), .RST(rst), .Q(c[560]) );
  DFF \sreg_reg[559]  ( .D(c[561]), .CLK(clk), .RST(rst), .Q(c[559]) );
  DFF \sreg_reg[558]  ( .D(c[560]), .CLK(clk), .RST(rst), .Q(c[558]) );
  DFF \sreg_reg[557]  ( .D(c[559]), .CLK(clk), .RST(rst), .Q(c[557]) );
  DFF \sreg_reg[556]  ( .D(c[558]), .CLK(clk), .RST(rst), .Q(c[556]) );
  DFF \sreg_reg[555]  ( .D(c[557]), .CLK(clk), .RST(rst), .Q(c[555]) );
  DFF \sreg_reg[554]  ( .D(c[556]), .CLK(clk), .RST(rst), .Q(c[554]) );
  DFF \sreg_reg[553]  ( .D(c[555]), .CLK(clk), .RST(rst), .Q(c[553]) );
  DFF \sreg_reg[552]  ( .D(c[554]), .CLK(clk), .RST(rst), .Q(c[552]) );
  DFF \sreg_reg[551]  ( .D(c[553]), .CLK(clk), .RST(rst), .Q(c[551]) );
  DFF \sreg_reg[550]  ( .D(c[552]), .CLK(clk), .RST(rst), .Q(c[550]) );
  DFF \sreg_reg[549]  ( .D(c[551]), .CLK(clk), .RST(rst), .Q(c[549]) );
  DFF \sreg_reg[548]  ( .D(c[550]), .CLK(clk), .RST(rst), .Q(c[548]) );
  DFF \sreg_reg[547]  ( .D(c[549]), .CLK(clk), .RST(rst), .Q(c[547]) );
  DFF \sreg_reg[546]  ( .D(c[548]), .CLK(clk), .RST(rst), .Q(c[546]) );
  DFF \sreg_reg[545]  ( .D(c[547]), .CLK(clk), .RST(rst), .Q(c[545]) );
  DFF \sreg_reg[544]  ( .D(c[546]), .CLK(clk), .RST(rst), .Q(c[544]) );
  DFF \sreg_reg[543]  ( .D(c[545]), .CLK(clk), .RST(rst), .Q(c[543]) );
  DFF \sreg_reg[542]  ( .D(c[544]), .CLK(clk), .RST(rst), .Q(c[542]) );
  DFF \sreg_reg[541]  ( .D(c[543]), .CLK(clk), .RST(rst), .Q(c[541]) );
  DFF \sreg_reg[540]  ( .D(c[542]), .CLK(clk), .RST(rst), .Q(c[540]) );
  DFF \sreg_reg[539]  ( .D(c[541]), .CLK(clk), .RST(rst), .Q(c[539]) );
  DFF \sreg_reg[538]  ( .D(c[540]), .CLK(clk), .RST(rst), .Q(c[538]) );
  DFF \sreg_reg[537]  ( .D(c[539]), .CLK(clk), .RST(rst), .Q(c[537]) );
  DFF \sreg_reg[536]  ( .D(c[538]), .CLK(clk), .RST(rst), .Q(c[536]) );
  DFF \sreg_reg[535]  ( .D(c[537]), .CLK(clk), .RST(rst), .Q(c[535]) );
  DFF \sreg_reg[534]  ( .D(c[536]), .CLK(clk), .RST(rst), .Q(c[534]) );
  DFF \sreg_reg[533]  ( .D(c[535]), .CLK(clk), .RST(rst), .Q(c[533]) );
  DFF \sreg_reg[532]  ( .D(c[534]), .CLK(clk), .RST(rst), .Q(c[532]) );
  DFF \sreg_reg[531]  ( .D(c[533]), .CLK(clk), .RST(rst), .Q(c[531]) );
  DFF \sreg_reg[530]  ( .D(c[532]), .CLK(clk), .RST(rst), .Q(c[530]) );
  DFF \sreg_reg[529]  ( .D(c[531]), .CLK(clk), .RST(rst), .Q(c[529]) );
  DFF \sreg_reg[528]  ( .D(c[530]), .CLK(clk), .RST(rst), .Q(c[528]) );
  DFF \sreg_reg[527]  ( .D(c[529]), .CLK(clk), .RST(rst), .Q(c[527]) );
  DFF \sreg_reg[526]  ( .D(c[528]), .CLK(clk), .RST(rst), .Q(c[526]) );
  DFF \sreg_reg[525]  ( .D(c[527]), .CLK(clk), .RST(rst), .Q(c[525]) );
  DFF \sreg_reg[524]  ( .D(c[526]), .CLK(clk), .RST(rst), .Q(c[524]) );
  DFF \sreg_reg[523]  ( .D(c[525]), .CLK(clk), .RST(rst), .Q(c[523]) );
  DFF \sreg_reg[522]  ( .D(c[524]), .CLK(clk), .RST(rst), .Q(c[522]) );
  DFF \sreg_reg[521]  ( .D(c[523]), .CLK(clk), .RST(rst), .Q(c[521]) );
  DFF \sreg_reg[520]  ( .D(c[522]), .CLK(clk), .RST(rst), .Q(c[520]) );
  DFF \sreg_reg[519]  ( .D(c[521]), .CLK(clk), .RST(rst), .Q(c[519]) );
  DFF \sreg_reg[518]  ( .D(c[520]), .CLK(clk), .RST(rst), .Q(c[518]) );
  DFF \sreg_reg[517]  ( .D(c[519]), .CLK(clk), .RST(rst), .Q(c[517]) );
  DFF \sreg_reg[516]  ( .D(c[518]), .CLK(clk), .RST(rst), .Q(c[516]) );
  DFF \sreg_reg[515]  ( .D(c[517]), .CLK(clk), .RST(rst), .Q(c[515]) );
  DFF \sreg_reg[514]  ( .D(c[516]), .CLK(clk), .RST(rst), .Q(c[514]) );
  DFF \sreg_reg[513]  ( .D(c[515]), .CLK(clk), .RST(rst), .Q(c[513]) );
  DFF \sreg_reg[512]  ( .D(c[514]), .CLK(clk), .RST(rst), .Q(c[512]) );
  DFF \sreg_reg[511]  ( .D(c[513]), .CLK(clk), .RST(rst), .Q(c[511]) );
  DFF \sreg_reg[510]  ( .D(c[512]), .CLK(clk), .RST(rst), .Q(c[510]) );
  DFF \sreg_reg[509]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(c[509]) );
  DFF \sreg_reg[508]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(c[508]) );
  DFF \sreg_reg[507]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(c[507]) );
  DFF \sreg_reg[506]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(c[506]) );
  DFF \sreg_reg[505]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(c[505]) );
  DFF \sreg_reg[504]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(c[504]) );
  DFF \sreg_reg[503]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(c[503]) );
  DFF \sreg_reg[502]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(c[502]) );
  DFF \sreg_reg[501]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(c[501]) );
  DFF \sreg_reg[500]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(c[500]) );
  DFF \sreg_reg[499]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(c[499]) );
  DFF \sreg_reg[498]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(c[498]) );
  DFF \sreg_reg[497]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(c[497]) );
  DFF \sreg_reg[496]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(c[496]) );
  DFF \sreg_reg[495]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(c[495]) );
  DFF \sreg_reg[494]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(c[494]) );
  DFF \sreg_reg[493]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(c[493]) );
  DFF \sreg_reg[492]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(c[492]) );
  DFF \sreg_reg[491]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(c[491]) );
  DFF \sreg_reg[490]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(c[490]) );
  DFF \sreg_reg[489]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(c[489]) );
  DFF \sreg_reg[488]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(c[488]) );
  DFF \sreg_reg[487]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(c[487]) );
  DFF \sreg_reg[486]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(c[486]) );
  DFF \sreg_reg[485]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(c[485]) );
  DFF \sreg_reg[484]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(c[484]) );
  DFF \sreg_reg[483]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(c[483]) );
  DFF \sreg_reg[482]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(c[482]) );
  DFF \sreg_reg[481]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(c[481]) );
  DFF \sreg_reg[480]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(c[480]) );
  DFF \sreg_reg[479]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(c[479]) );
  DFF \sreg_reg[478]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(c[478]) );
  DFF \sreg_reg[477]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(c[477]) );
  DFF \sreg_reg[476]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(c[476]) );
  DFF \sreg_reg[475]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(c[475]) );
  DFF \sreg_reg[474]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(c[474]) );
  DFF \sreg_reg[473]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(c[473]) );
  DFF \sreg_reg[472]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(c[472]) );
  DFF \sreg_reg[471]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(c[471]) );
  DFF \sreg_reg[470]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(c[470]) );
  DFF \sreg_reg[469]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(c[469]) );
  DFF \sreg_reg[468]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(c[468]) );
  DFF \sreg_reg[467]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(c[467]) );
  DFF \sreg_reg[466]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(c[466]) );
  DFF \sreg_reg[465]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(c[465]) );
  DFF \sreg_reg[464]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(c[464]) );
  DFF \sreg_reg[463]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(c[463]) );
  DFF \sreg_reg[462]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(c[462]) );
  DFF \sreg_reg[461]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(c[461]) );
  DFF \sreg_reg[460]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(c[460]) );
  DFF \sreg_reg[459]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(c[459]) );
  DFF \sreg_reg[458]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(c[458]) );
  DFF \sreg_reg[457]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(c[457]) );
  DFF \sreg_reg[456]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(c[456]) );
  DFF \sreg_reg[455]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(c[455]) );
  DFF \sreg_reg[454]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(c[454]) );
  DFF \sreg_reg[453]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(c[453]) );
  DFF \sreg_reg[452]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(c[452]) );
  DFF \sreg_reg[451]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(c[451]) );
  DFF \sreg_reg[450]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(c[450]) );
  DFF \sreg_reg[449]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(c[449]) );
  DFF \sreg_reg[448]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(c[448]) );
  DFF \sreg_reg[447]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(c[447]) );
  DFF \sreg_reg[446]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(c[446]) );
  DFF \sreg_reg[445]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(c[445]) );
  DFF \sreg_reg[444]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(c[444]) );
  DFF \sreg_reg[443]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(c[443]) );
  DFF \sreg_reg[442]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(c[442]) );
  DFF \sreg_reg[441]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(c[441]) );
  DFF \sreg_reg[440]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(c[440]) );
  DFF \sreg_reg[439]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(c[439]) );
  DFF \sreg_reg[438]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(c[438]) );
  DFF \sreg_reg[437]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(c[437]) );
  DFF \sreg_reg[436]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(c[436]) );
  DFF \sreg_reg[435]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(c[435]) );
  DFF \sreg_reg[434]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(c[434]) );
  DFF \sreg_reg[433]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(c[433]) );
  DFF \sreg_reg[432]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(c[432]) );
  DFF \sreg_reg[431]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(c[431]) );
  DFF \sreg_reg[430]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(c[430]) );
  DFF \sreg_reg[429]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(c[429]) );
  DFF \sreg_reg[428]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(c[428]) );
  DFF \sreg_reg[427]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(c[427]) );
  DFF \sreg_reg[426]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(c[426]) );
  DFF \sreg_reg[425]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(c[425]) );
  DFF \sreg_reg[424]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(c[424]) );
  DFF \sreg_reg[423]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(c[423]) );
  DFF \sreg_reg[422]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(c[422]) );
  DFF \sreg_reg[421]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(c[421]) );
  DFF \sreg_reg[420]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(c[420]) );
  DFF \sreg_reg[419]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(c[419]) );
  DFF \sreg_reg[418]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(c[418]) );
  DFF \sreg_reg[417]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(c[417]) );
  DFF \sreg_reg[416]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(c[416]) );
  DFF \sreg_reg[415]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(c[415]) );
  DFF \sreg_reg[414]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(c[414]) );
  DFF \sreg_reg[413]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(c[413]) );
  DFF \sreg_reg[412]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(c[412]) );
  DFF \sreg_reg[411]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(c[411]) );
  DFF \sreg_reg[410]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(c[410]) );
  DFF \sreg_reg[409]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(c[409]) );
  DFF \sreg_reg[408]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(c[408]) );
  DFF \sreg_reg[407]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(c[407]) );
  DFF \sreg_reg[406]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(c[406]) );
  DFF \sreg_reg[405]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(c[405]) );
  DFF \sreg_reg[404]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(c[404]) );
  DFF \sreg_reg[403]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(c[403]) );
  DFF \sreg_reg[402]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(c[402]) );
  DFF \sreg_reg[401]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(c[401]) );
  DFF \sreg_reg[400]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(c[400]) );
  DFF \sreg_reg[399]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(c[399]) );
  DFF \sreg_reg[398]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(c[398]) );
  DFF \sreg_reg[397]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(c[397]) );
  DFF \sreg_reg[396]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(c[396]) );
  DFF \sreg_reg[395]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(c[395]) );
  DFF \sreg_reg[394]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(c[394]) );
  DFF \sreg_reg[393]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(c[393]) );
  DFF \sreg_reg[392]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(c[392]) );
  DFF \sreg_reg[391]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(c[391]) );
  DFF \sreg_reg[390]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(c[390]) );
  DFF \sreg_reg[389]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(c[389]) );
  DFF \sreg_reg[388]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(c[388]) );
  DFF \sreg_reg[387]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(c[387]) );
  DFF \sreg_reg[386]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(c[386]) );
  DFF \sreg_reg[385]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(c[385]) );
  DFF \sreg_reg[384]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(c[384]) );
  DFF \sreg_reg[383]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(c[383]) );
  DFF \sreg_reg[382]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(c[382]) );
  DFF \sreg_reg[381]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(c[381]) );
  DFF \sreg_reg[380]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(c[380]) );
  DFF \sreg_reg[379]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(c[379]) );
  DFF \sreg_reg[378]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(c[378]) );
  DFF \sreg_reg[377]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(c[377]) );
  DFF \sreg_reg[376]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(c[376]) );
  DFF \sreg_reg[375]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(c[375]) );
  DFF \sreg_reg[374]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(c[374]) );
  DFF \sreg_reg[373]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(c[373]) );
  DFF \sreg_reg[372]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(c[372]) );
  DFF \sreg_reg[371]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(c[371]) );
  DFF \sreg_reg[370]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(c[370]) );
  DFF \sreg_reg[369]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(c[369]) );
  DFF \sreg_reg[368]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(c[368]) );
  DFF \sreg_reg[367]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(c[367]) );
  DFF \sreg_reg[366]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(c[366]) );
  DFF \sreg_reg[365]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(c[365]) );
  DFF \sreg_reg[364]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(c[364]) );
  DFF \sreg_reg[363]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(c[363]) );
  DFF \sreg_reg[362]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(c[362]) );
  DFF \sreg_reg[361]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(c[361]) );
  DFF \sreg_reg[360]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(c[360]) );
  DFF \sreg_reg[359]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(c[359]) );
  DFF \sreg_reg[358]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(c[358]) );
  DFF \sreg_reg[357]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(c[357]) );
  DFF \sreg_reg[356]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(c[356]) );
  DFF \sreg_reg[355]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(c[355]) );
  DFF \sreg_reg[354]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(c[354]) );
  DFF \sreg_reg[353]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(c[353]) );
  DFF \sreg_reg[352]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(c[352]) );
  DFF \sreg_reg[351]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(c[351]) );
  DFF \sreg_reg[350]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(c[350]) );
  DFF \sreg_reg[349]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(c[349]) );
  DFF \sreg_reg[348]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(c[348]) );
  DFF \sreg_reg[347]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(c[347]) );
  DFF \sreg_reg[346]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(c[346]) );
  DFF \sreg_reg[345]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(c[345]) );
  DFF \sreg_reg[344]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(c[344]) );
  DFF \sreg_reg[343]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(c[343]) );
  DFF \sreg_reg[342]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(c[342]) );
  DFF \sreg_reg[341]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(c[341]) );
  DFF \sreg_reg[340]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(c[340]) );
  DFF \sreg_reg[339]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(c[339]) );
  DFF \sreg_reg[338]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(c[338]) );
  DFF \sreg_reg[337]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(c[337]) );
  DFF \sreg_reg[336]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(c[336]) );
  DFF \sreg_reg[335]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(c[335]) );
  DFF \sreg_reg[334]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(c[334]) );
  DFF \sreg_reg[333]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(c[333]) );
  DFF \sreg_reg[332]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(c[332]) );
  DFF \sreg_reg[331]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(c[331]) );
  DFF \sreg_reg[330]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(c[330]) );
  DFF \sreg_reg[329]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(c[329]) );
  DFF \sreg_reg[328]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(c[328]) );
  DFF \sreg_reg[327]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(c[327]) );
  DFF \sreg_reg[326]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(c[326]) );
  DFF \sreg_reg[325]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(c[325]) );
  DFF \sreg_reg[324]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(c[324]) );
  DFF \sreg_reg[323]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(c[323]) );
  DFF \sreg_reg[322]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(c[322]) );
  DFF \sreg_reg[321]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(c[321]) );
  DFF \sreg_reg[320]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(c[320]) );
  DFF \sreg_reg[319]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(c[319]) );
  DFF \sreg_reg[318]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(c[318]) );
  DFF \sreg_reg[317]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(c[317]) );
  DFF \sreg_reg[316]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(c[316]) );
  DFF \sreg_reg[315]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(c[315]) );
  DFF \sreg_reg[314]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(c[314]) );
  DFF \sreg_reg[313]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(c[313]) );
  DFF \sreg_reg[312]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(c[312]) );
  DFF \sreg_reg[311]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(c[311]) );
  DFF \sreg_reg[310]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(c[310]) );
  DFF \sreg_reg[309]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(c[309]) );
  DFF \sreg_reg[308]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(c[308]) );
  DFF \sreg_reg[307]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(c[307]) );
  DFF \sreg_reg[306]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(c[306]) );
  DFF \sreg_reg[305]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(c[305]) );
  DFF \sreg_reg[304]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(c[304]) );
  DFF \sreg_reg[303]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(c[303]) );
  DFF \sreg_reg[302]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(c[302]) );
  DFF \sreg_reg[301]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(c[301]) );
  DFF \sreg_reg[300]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(c[300]) );
  DFF \sreg_reg[299]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(c[299]) );
  DFF \sreg_reg[298]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(c[298]) );
  DFF \sreg_reg[297]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(c[297]) );
  DFF \sreg_reg[296]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(c[296]) );
  DFF \sreg_reg[295]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(c[295]) );
  DFF \sreg_reg[294]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(c[294]) );
  DFF \sreg_reg[293]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(c[293]) );
  DFF \sreg_reg[292]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(c[292]) );
  DFF \sreg_reg[291]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(c[291]) );
  DFF \sreg_reg[290]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(c[290]) );
  DFF \sreg_reg[289]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(c[289]) );
  DFF \sreg_reg[288]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(c[288]) );
  DFF \sreg_reg[287]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(c[287]) );
  DFF \sreg_reg[286]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(c[286]) );
  DFF \sreg_reg[285]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(c[285]) );
  DFF \sreg_reg[284]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(c[284]) );
  DFF \sreg_reg[283]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(c[283]) );
  DFF \sreg_reg[282]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(c[282]) );
  DFF \sreg_reg[281]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(c[281]) );
  DFF \sreg_reg[280]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(c[280]) );
  DFF \sreg_reg[279]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(c[279]) );
  DFF \sreg_reg[278]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(c[278]) );
  DFF \sreg_reg[277]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(c[277]) );
  DFF \sreg_reg[276]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(c[276]) );
  DFF \sreg_reg[275]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(c[275]) );
  DFF \sreg_reg[274]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(c[274]) );
  DFF \sreg_reg[273]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(c[273]) );
  DFF \sreg_reg[272]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(c[272]) );
  DFF \sreg_reg[271]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(c[271]) );
  DFF \sreg_reg[270]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(c[270]) );
  DFF \sreg_reg[269]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(c[269]) );
  DFF \sreg_reg[268]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(c[268]) );
  DFF \sreg_reg[267]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(c[267]) );
  DFF \sreg_reg[266]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(c[266]) );
  DFF \sreg_reg[265]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(c[265]) );
  DFF \sreg_reg[264]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(c[264]) );
  DFF \sreg_reg[263]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(c[263]) );
  DFF \sreg_reg[262]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(c[262]) );
  DFF \sreg_reg[261]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(c[261]) );
  DFF \sreg_reg[260]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(c[260]) );
  DFF \sreg_reg[259]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(c[259]) );
  DFF \sreg_reg[258]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(c[258]) );
  DFF \sreg_reg[257]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(c[257]) );
  DFF \sreg_reg[256]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(c[256]) );
  DFF \sreg_reg[255]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(c[255]) );
  DFF \sreg_reg[254]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(c[254]) );
  DFF \sreg_reg[253]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[252]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[251]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[0]) );
  OR U5 ( .A(n4276), .B(n4275), .Z(n1) );
  NAND U6 ( .A(n4278), .B(n4277), .Z(n2) );
  NAND U7 ( .A(n1), .B(n2), .Z(n4284) );
  OR U8 ( .A(n4391), .B(n4390), .Z(n3) );
  NAND U9 ( .A(n4393), .B(n4392), .Z(n4) );
  NAND U10 ( .A(n3), .B(n4), .Z(n4399) );
  OR U11 ( .A(n4488), .B(n4487), .Z(n5) );
  NAND U12 ( .A(n4490), .B(n4489), .Z(n6) );
  NAND U13 ( .A(n5), .B(n6), .Z(n4496) );
  OR U14 ( .A(n4612), .B(n4611), .Z(n7) );
  NAND U15 ( .A(n4614), .B(n4613), .Z(n8) );
  NAND U16 ( .A(n7), .B(n8), .Z(n4621) );
  OR U17 ( .A(n4700), .B(n4699), .Z(n9) );
  NAND U18 ( .A(n4702), .B(n4701), .Z(n10) );
  NAND U19 ( .A(n9), .B(n10), .Z(n4708) );
  OR U20 ( .A(n4833), .B(n4832), .Z(n11) );
  NAND U21 ( .A(n4835), .B(n4834), .Z(n12) );
  NAND U22 ( .A(n11), .B(n12), .Z(n4841) );
  OR U23 ( .A(n4966), .B(n4965), .Z(n13) );
  NAND U24 ( .A(n4968), .B(n4967), .Z(n14) );
  NAND U25 ( .A(n13), .B(n14), .Z(n4974) );
  OR U26 ( .A(n5135), .B(n5134), .Z(n15) );
  NAND U27 ( .A(n5137), .B(n5136), .Z(n16) );
  NAND U28 ( .A(n15), .B(n16), .Z(n5143) );
  OR U29 ( .A(n5250), .B(n5249), .Z(n17) );
  NAND U30 ( .A(n5252), .B(n5251), .Z(n18) );
  NAND U31 ( .A(n17), .B(n18), .Z(n5258) );
  OR U32 ( .A(n5365), .B(n5364), .Z(n19) );
  NAND U33 ( .A(n5367), .B(n5366), .Z(n20) );
  NAND U34 ( .A(n19), .B(n20), .Z(n5373) );
  OR U35 ( .A(n5462), .B(n5461), .Z(n21) );
  NAND U36 ( .A(n5464), .B(n5463), .Z(n22) );
  NAND U37 ( .A(n21), .B(n22), .Z(n5470) );
  OR U38 ( .A(n5595), .B(n5594), .Z(n23) );
  NAND U39 ( .A(n5597), .B(n5596), .Z(n24) );
  NAND U40 ( .A(n23), .B(n24), .Z(n5603) );
  OR U41 ( .A(n5692), .B(n5691), .Z(n25) );
  NAND U42 ( .A(n5694), .B(n5693), .Z(n26) );
  NAND U43 ( .A(n25), .B(n26), .Z(n5700) );
  OR U44 ( .A(n5843), .B(n5842), .Z(n27) );
  NAND U45 ( .A(n5845), .B(n5844), .Z(n28) );
  NAND U46 ( .A(n27), .B(n28), .Z(n5851) );
  OR U47 ( .A(n5967), .B(n5966), .Z(n29) );
  NAND U48 ( .A(n5969), .B(n5968), .Z(n30) );
  NAND U49 ( .A(n29), .B(n30), .Z(n5976) );
  OR U50 ( .A(n6073), .B(n6072), .Z(n31) );
  NAND U51 ( .A(n6075), .B(n6074), .Z(n32) );
  NAND U52 ( .A(n31), .B(n32), .Z(n6081) );
  OR U53 ( .A(n6161), .B(n6160), .Z(n33) );
  NAND U54 ( .A(n6163), .B(n6162), .Z(n34) );
  NAND U55 ( .A(n33), .B(n34), .Z(n6170) );
  OR U56 ( .A(n6285), .B(n6284), .Z(n35) );
  NAND U57 ( .A(n6287), .B(n6286), .Z(n36) );
  NAND U58 ( .A(n35), .B(n36), .Z(n6293) );
  OR U59 ( .A(n6436), .B(n6435), .Z(n37) );
  NAND U60 ( .A(n6438), .B(n6437), .Z(n38) );
  NAND U61 ( .A(n37), .B(n38), .Z(n6444) );
  OR U62 ( .A(n6551), .B(n6550), .Z(n39) );
  NAND U63 ( .A(n6553), .B(n6552), .Z(n40) );
  NAND U64 ( .A(n39), .B(n40), .Z(n6559) );
  OR U65 ( .A(n6666), .B(n6665), .Z(n41) );
  NAND U66 ( .A(n6668), .B(n6667), .Z(n42) );
  NAND U67 ( .A(n41), .B(n42), .Z(n6674) );
  OR U68 ( .A(n6763), .B(n6762), .Z(n43) );
  NAND U69 ( .A(n6765), .B(n6764), .Z(n44) );
  NAND U70 ( .A(n43), .B(n44), .Z(n6771) );
  OR U71 ( .A(n6932), .B(n6931), .Z(n45) );
  NAND U72 ( .A(n6934), .B(n6933), .Z(n46) );
  NAND U73 ( .A(n45), .B(n46), .Z(n6940) );
  OR U74 ( .A(n7011), .B(n7010), .Z(n47) );
  NAND U75 ( .A(n7013), .B(n7012), .Z(n48) );
  NAND U76 ( .A(n47), .B(n48), .Z(n7019) );
  OR U77 ( .A(n7108), .B(n7107), .Z(n49) );
  NAND U78 ( .A(n7110), .B(n7109), .Z(n50) );
  NAND U79 ( .A(n49), .B(n50), .Z(n7117) );
  OR U80 ( .A(n7205), .B(n7204), .Z(n51) );
  NAND U81 ( .A(n7207), .B(n7206), .Z(n52) );
  NAND U82 ( .A(n51), .B(n52), .Z(n7213) );
  OR U83 ( .A(n7320), .B(n7319), .Z(n53) );
  NAND U84 ( .A(n7322), .B(n7321), .Z(n54) );
  NAND U85 ( .A(n53), .B(n54), .Z(n7328) );
  OR U86 ( .A(n7453), .B(n7452), .Z(n55) );
  NAND U87 ( .A(n7455), .B(n7454), .Z(n56) );
  NAND U88 ( .A(n55), .B(n56), .Z(n7462) );
  OR U89 ( .A(n7550), .B(n7549), .Z(n57) );
  NAND U90 ( .A(n7552), .B(n7551), .Z(n58) );
  NAND U91 ( .A(n57), .B(n58), .Z(n7558) );
  OR U92 ( .A(n7665), .B(n7664), .Z(n59) );
  NAND U93 ( .A(n7667), .B(n7666), .Z(n60) );
  NAND U94 ( .A(n59), .B(n60), .Z(n7673) );
  OR U95 ( .A(n7789), .B(n7788), .Z(n61) );
  NAND U96 ( .A(n7791), .B(n7790), .Z(n62) );
  NAND U97 ( .A(n61), .B(n62), .Z(n7798) );
  OR U98 ( .A(n7877), .B(n7876), .Z(n63) );
  NAND U99 ( .A(n7879), .B(n7878), .Z(n64) );
  NAND U100 ( .A(n63), .B(n64), .Z(n7885) );
  OR U101 ( .A(n7983), .B(n7982), .Z(n65) );
  NAND U102 ( .A(n7985), .B(n7984), .Z(n66) );
  NAND U103 ( .A(n65), .B(n66), .Z(n7992) );
  OR U104 ( .A(n8089), .B(n8088), .Z(n67) );
  NAND U105 ( .A(n8091), .B(n8090), .Z(n68) );
  NAND U106 ( .A(n67), .B(n68), .Z(n8097) );
  OR U107 ( .A(n8204), .B(n8203), .Z(n69) );
  NAND U108 ( .A(n8206), .B(n8205), .Z(n70) );
  NAND U109 ( .A(n69), .B(n70), .Z(n8212) );
  OR U110 ( .A(n8301), .B(n8300), .Z(n71) );
  NAND U111 ( .A(n8303), .B(n8302), .Z(n72) );
  NAND U112 ( .A(n71), .B(n72), .Z(n8309) );
  OR U113 ( .A(n8416), .B(n8415), .Z(n73) );
  NAND U114 ( .A(n8418), .B(n8417), .Z(n74) );
  NAND U115 ( .A(n73), .B(n74), .Z(n8425) );
  OR U116 ( .A(n8549), .B(n8548), .Z(n75) );
  NAND U117 ( .A(n8551), .B(n8550), .Z(n76) );
  NAND U118 ( .A(n75), .B(n76), .Z(n8557) );
  OR U119 ( .A(n8664), .B(n8663), .Z(n77) );
  NAND U120 ( .A(n8666), .B(n8665), .Z(n78) );
  NAND U121 ( .A(n77), .B(n78), .Z(n8672) );
  OR U122 ( .A(n8779), .B(n8778), .Z(n79) );
  NAND U123 ( .A(n8781), .B(n8780), .Z(n80) );
  NAND U124 ( .A(n79), .B(n80), .Z(n8787) );
  OR U125 ( .A(n8912), .B(n8911), .Z(n81) );
  NAND U126 ( .A(n8914), .B(n8913), .Z(n82) );
  NAND U127 ( .A(n81), .B(n82), .Z(n8920) );
  OR U128 ( .A(n9045), .B(n9044), .Z(n83) );
  NAND U129 ( .A(n9047), .B(n9046), .Z(n84) );
  NAND U130 ( .A(n83), .B(n84), .Z(n9053) );
  OR U131 ( .A(n9160), .B(n9159), .Z(n85) );
  NAND U132 ( .A(n9162), .B(n9161), .Z(n86) );
  NAND U133 ( .A(n85), .B(n86), .Z(n9168) );
  OR U134 ( .A(n9239), .B(n9238), .Z(n87) );
  NAND U135 ( .A(n9241), .B(n9240), .Z(n88) );
  NAND U136 ( .A(n87), .B(n88), .Z(n9247) );
  OR U137 ( .A(n9354), .B(n9353), .Z(n89) );
  NAND U138 ( .A(n9356), .B(n9355), .Z(n90) );
  NAND U139 ( .A(n89), .B(n90), .Z(n9362) );
  OR U140 ( .A(n9433), .B(n9432), .Z(n91) );
  NAND U141 ( .A(n9435), .B(n9434), .Z(n92) );
  NAND U142 ( .A(n91), .B(n92), .Z(n9441) );
  OR U143 ( .A(n9548), .B(n9547), .Z(n93) );
  NAND U144 ( .A(n9550), .B(n9549), .Z(n94) );
  NAND U145 ( .A(n93), .B(n94), .Z(n9556) );
  OR U146 ( .A(n9681), .B(n9680), .Z(n95) );
  NAND U147 ( .A(n9683), .B(n9682), .Z(n96) );
  NAND U148 ( .A(n95), .B(n96), .Z(n9689) );
  OR U149 ( .A(n9778), .B(n9777), .Z(n97) );
  NAND U150 ( .A(n9780), .B(n9779), .Z(n98) );
  NAND U151 ( .A(n97), .B(n98), .Z(n9786) );
  OR U152 ( .A(n9875), .B(n9874), .Z(n99) );
  NAND U153 ( .A(n9877), .B(n9876), .Z(n100) );
  NAND U154 ( .A(n99), .B(n100), .Z(n9883) );
  OR U155 ( .A(n9990), .B(n9989), .Z(n101) );
  NAND U156 ( .A(n9992), .B(n9991), .Z(n102) );
  NAND U157 ( .A(n101), .B(n102), .Z(n9998) );
  OR U158 ( .A(n10123), .B(n10122), .Z(n103) );
  NAND U159 ( .A(n10125), .B(n10124), .Z(n104) );
  NAND U160 ( .A(n103), .B(n104), .Z(n10131) );
  OR U161 ( .A(n10220), .B(n10219), .Z(n105) );
  NAND U162 ( .A(n10222), .B(n10221), .Z(n106) );
  NAND U163 ( .A(n105), .B(n106), .Z(n10228) );
  OR U164 ( .A(n10353), .B(n10352), .Z(n107) );
  NAND U165 ( .A(n10355), .B(n10354), .Z(n108) );
  NAND U166 ( .A(n107), .B(n108), .Z(n10361) );
  OR U167 ( .A(n10468), .B(n10467), .Z(n109) );
  NAND U168 ( .A(n10470), .B(n10469), .Z(n110) );
  NAND U169 ( .A(n109), .B(n110), .Z(n10477) );
  OR U170 ( .A(n10565), .B(n10564), .Z(n111) );
  NAND U171 ( .A(n10567), .B(n10566), .Z(n112) );
  NAND U172 ( .A(n111), .B(n112), .Z(n10573) );
  OR U173 ( .A(n10680), .B(n10679), .Z(n113) );
  NAND U174 ( .A(n10682), .B(n10681), .Z(n114) );
  NAND U175 ( .A(n113), .B(n114), .Z(n10689) );
  OR U176 ( .A(n10786), .B(n10785), .Z(n115) );
  NAND U177 ( .A(n10788), .B(n10787), .Z(n116) );
  NAND U178 ( .A(n115), .B(n116), .Z(n10794) );
  OR U179 ( .A(n10946), .B(n10945), .Z(n117) );
  NAND U180 ( .A(n10948), .B(n10947), .Z(n118) );
  NAND U181 ( .A(n117), .B(n118), .Z(n10954) );
  OR U182 ( .A(n11115), .B(n11114), .Z(n119) );
  NAND U183 ( .A(n11117), .B(n11116), .Z(n120) );
  NAND U184 ( .A(n119), .B(n120), .Z(n11123) );
  OR U185 ( .A(n11203), .B(n11202), .Z(n121) );
  NAND U186 ( .A(n11205), .B(n11204), .Z(n122) );
  NAND U187 ( .A(n121), .B(n122), .Z(n11212) );
  OR U188 ( .A(n11309), .B(n11308), .Z(n123) );
  NAND U189 ( .A(n11311), .B(n11310), .Z(n124) );
  NAND U190 ( .A(n123), .B(n124), .Z(n11317) );
  OR U191 ( .A(n11478), .B(n11477), .Z(n125) );
  NAND U192 ( .A(n11480), .B(n11479), .Z(n126) );
  NAND U193 ( .A(n125), .B(n126), .Z(n11486) );
  OR U194 ( .A(n11611), .B(n11610), .Z(n127) );
  NAND U195 ( .A(n11613), .B(n11612), .Z(n128) );
  NAND U196 ( .A(n127), .B(n128), .Z(n11619) );
  OR U197 ( .A(n11744), .B(n11743), .Z(n129) );
  NAND U198 ( .A(n11746), .B(n11745), .Z(n130) );
  NAND U199 ( .A(n129), .B(n130), .Z(n11752) );
  OR U200 ( .A(n11913), .B(n11912), .Z(n131) );
  NAND U201 ( .A(n11915), .B(n11914), .Z(n132) );
  NAND U202 ( .A(n131), .B(n132), .Z(n11921) );
  OR U203 ( .A(n12019), .B(n12018), .Z(n133) );
  NAND U204 ( .A(n12021), .B(n12020), .Z(n134) );
  NAND U205 ( .A(n133), .B(n134), .Z(n12027) );
  OR U206 ( .A(n12116), .B(n12115), .Z(n135) );
  NAND U207 ( .A(n12118), .B(n12117), .Z(n136) );
  NAND U208 ( .A(n135), .B(n136), .Z(n12125) );
  OR U209 ( .A(n12213), .B(n12212), .Z(n137) );
  NAND U210 ( .A(n12215), .B(n12214), .Z(n138) );
  NAND U211 ( .A(n137), .B(n138), .Z(n12222) );
  OR U212 ( .A(n4292), .B(n4291), .Z(n139) );
  NAND U213 ( .A(n4294), .B(n4293), .Z(n140) );
  NAND U214 ( .A(n139), .B(n140), .Z(n4300) );
  OR U215 ( .A(n4407), .B(n4406), .Z(n141) );
  NAND U216 ( .A(n4409), .B(n4408), .Z(n142) );
  NAND U217 ( .A(n141), .B(n142), .Z(n4415) );
  OR U218 ( .A(n4522), .B(n4521), .Z(n143) );
  NAND U219 ( .A(n4524), .B(n4523), .Z(n144) );
  NAND U220 ( .A(n143), .B(n144), .Z(n4530) );
  OR U221 ( .A(n4619), .B(n4618), .Z(n145) );
  NAND U222 ( .A(n4621), .B(n4620), .Z(n146) );
  NAND U223 ( .A(n145), .B(n146), .Z(n4628) );
  OR U224 ( .A(n4716), .B(n4715), .Z(n147) );
  NAND U225 ( .A(n4718), .B(n4717), .Z(n148) );
  NAND U226 ( .A(n147), .B(n148), .Z(n4724) );
  OR U227 ( .A(n4849), .B(n4848), .Z(n149) );
  NAND U228 ( .A(n4851), .B(n4850), .Z(n150) );
  NAND U229 ( .A(n149), .B(n150), .Z(n4857) );
  OR U230 ( .A(n4982), .B(n4981), .Z(n151) );
  NAND U231 ( .A(n4984), .B(n4983), .Z(n152) );
  NAND U232 ( .A(n151), .B(n152), .Z(n4990) );
  OR U233 ( .A(n5151), .B(n5150), .Z(n153) );
  NAND U234 ( .A(n5153), .B(n5152), .Z(n154) );
  NAND U235 ( .A(n153), .B(n154), .Z(n5159) );
  OR U236 ( .A(n5266), .B(n5265), .Z(n155) );
  NAND U237 ( .A(n5268), .B(n5267), .Z(n156) );
  NAND U238 ( .A(n155), .B(n156), .Z(n5274) );
  OR U239 ( .A(n5381), .B(n5380), .Z(n157) );
  NAND U240 ( .A(n5383), .B(n5382), .Z(n158) );
  NAND U241 ( .A(n157), .B(n158), .Z(n5390) );
  OR U242 ( .A(n5478), .B(n5477), .Z(n159) );
  NAND U243 ( .A(n5480), .B(n5479), .Z(n160) );
  NAND U244 ( .A(n159), .B(n160), .Z(n5486) );
  OR U245 ( .A(n5611), .B(n5610), .Z(n161) );
  NAND U246 ( .A(n5613), .B(n5612), .Z(n162) );
  NAND U247 ( .A(n161), .B(n162), .Z(n5619) );
  OR U248 ( .A(n5708), .B(n5707), .Z(n163) );
  NAND U249 ( .A(n5710), .B(n5709), .Z(n164) );
  NAND U250 ( .A(n163), .B(n164), .Z(n5716) );
  OR U251 ( .A(n5859), .B(n5858), .Z(n165) );
  NAND U252 ( .A(n5861), .B(n5860), .Z(n166) );
  NAND U253 ( .A(n165), .B(n166), .Z(n5867) );
  OR U254 ( .A(n5974), .B(n5973), .Z(n167) );
  NAND U255 ( .A(n5976), .B(n5975), .Z(n168) );
  NAND U256 ( .A(n167), .B(n168), .Z(n5982) );
  OR U257 ( .A(n6089), .B(n6088), .Z(n169) );
  NAND U258 ( .A(n6091), .B(n6090), .Z(n170) );
  NAND U259 ( .A(n169), .B(n170), .Z(n6097) );
  OR U260 ( .A(n6168), .B(n6167), .Z(n171) );
  NAND U261 ( .A(n6170), .B(n6169), .Z(n172) );
  NAND U262 ( .A(n171), .B(n172), .Z(n6176) );
  OR U263 ( .A(n6301), .B(n6300), .Z(n173) );
  NAND U264 ( .A(n6303), .B(n6302), .Z(n174) );
  NAND U265 ( .A(n173), .B(n174), .Z(n6309) );
  OR U266 ( .A(n6452), .B(n6451), .Z(n175) );
  NAND U267 ( .A(n6454), .B(n6453), .Z(n176) );
  NAND U268 ( .A(n175), .B(n176), .Z(n6460) );
  OR U269 ( .A(n6567), .B(n6566), .Z(n177) );
  NAND U270 ( .A(n6569), .B(n6568), .Z(n178) );
  NAND U271 ( .A(n177), .B(n178), .Z(n6575) );
  OR U272 ( .A(n6700), .B(n6699), .Z(n179) );
  NAND U273 ( .A(n6702), .B(n6701), .Z(n180) );
  NAND U274 ( .A(n179), .B(n180), .Z(n6709) );
  OR U275 ( .A(n6779), .B(n6778), .Z(n181) );
  NAND U276 ( .A(n6781), .B(n6780), .Z(n182) );
  NAND U277 ( .A(n181), .B(n182), .Z(n6787) );
  OR U278 ( .A(n6948), .B(n6947), .Z(n183) );
  NAND U279 ( .A(n6950), .B(n6949), .Z(n184) );
  NAND U280 ( .A(n183), .B(n184), .Z(n6956) );
  OR U281 ( .A(n7027), .B(n7026), .Z(n185) );
  NAND U282 ( .A(n7029), .B(n7028), .Z(n186) );
  NAND U283 ( .A(n185), .B(n186), .Z(n7035) );
  OR U284 ( .A(n7115), .B(n7114), .Z(n187) );
  NAND U285 ( .A(n7117), .B(n7116), .Z(n188) );
  NAND U286 ( .A(n187), .B(n188), .Z(n7124) );
  OR U287 ( .A(n7221), .B(n7220), .Z(n189) );
  NAND U288 ( .A(n7223), .B(n7222), .Z(n190) );
  NAND U289 ( .A(n189), .B(n190), .Z(n7229) );
  OR U290 ( .A(n7354), .B(n7353), .Z(n191) );
  NAND U291 ( .A(n7356), .B(n7355), .Z(n192) );
  NAND U292 ( .A(n191), .B(n192), .Z(n7362) );
  OR U293 ( .A(n7460), .B(n7459), .Z(n193) );
  NAND U294 ( .A(n7462), .B(n7461), .Z(n194) );
  NAND U295 ( .A(n193), .B(n194), .Z(n7468) );
  OR U296 ( .A(n7584), .B(n7583), .Z(n195) );
  NAND U297 ( .A(n7586), .B(n7585), .Z(n196) );
  NAND U298 ( .A(n195), .B(n196), .Z(n7593) );
  OR U299 ( .A(n7681), .B(n7680), .Z(n197) );
  NAND U300 ( .A(n7683), .B(n7682), .Z(n198) );
  NAND U301 ( .A(n197), .B(n198), .Z(n7689) );
  OR U302 ( .A(n7796), .B(n7795), .Z(n199) );
  NAND U303 ( .A(n7798), .B(n7797), .Z(n200) );
  NAND U304 ( .A(n199), .B(n200), .Z(n7805) );
  OR U305 ( .A(n7893), .B(n7892), .Z(n201) );
  NAND U306 ( .A(n7895), .B(n7894), .Z(n202) );
  NAND U307 ( .A(n201), .B(n202), .Z(n7901) );
  OR U308 ( .A(n7990), .B(n7989), .Z(n203) );
  NAND U309 ( .A(n7992), .B(n7991), .Z(n204) );
  NAND U310 ( .A(n203), .B(n204), .Z(n7998) );
  OR U311 ( .A(n8105), .B(n8104), .Z(n205) );
  NAND U312 ( .A(n8107), .B(n8106), .Z(n206) );
  NAND U313 ( .A(n205), .B(n206), .Z(n8113) );
  OR U314 ( .A(n8220), .B(n8219), .Z(n207) );
  NAND U315 ( .A(n8222), .B(n8221), .Z(n208) );
  NAND U316 ( .A(n207), .B(n208), .Z(n8228) );
  OR U317 ( .A(n8317), .B(n8316), .Z(n209) );
  NAND U318 ( .A(n8319), .B(n8318), .Z(n210) );
  NAND U319 ( .A(n209), .B(n210), .Z(n8325) );
  OR U320 ( .A(n8423), .B(n8422), .Z(n211) );
  NAND U321 ( .A(n8425), .B(n8424), .Z(n212) );
  NAND U322 ( .A(n211), .B(n212), .Z(n8432) );
  OR U323 ( .A(n8583), .B(n8582), .Z(n213) );
  NAND U324 ( .A(n8585), .B(n8584), .Z(n214) );
  NAND U325 ( .A(n213), .B(n214), .Z(n8591) );
  OR U326 ( .A(n8680), .B(n8679), .Z(n215) );
  NAND U327 ( .A(n8682), .B(n8681), .Z(n216) );
  NAND U328 ( .A(n215), .B(n216), .Z(n8688) );
  OR U329 ( .A(n8795), .B(n8794), .Z(n217) );
  NAND U330 ( .A(n8797), .B(n8796), .Z(n218) );
  NAND U331 ( .A(n217), .B(n218), .Z(n8803) );
  OR U332 ( .A(n8928), .B(n8927), .Z(n219) );
  NAND U333 ( .A(n8930), .B(n8929), .Z(n220) );
  NAND U334 ( .A(n219), .B(n220), .Z(n8936) );
  OR U335 ( .A(n9079), .B(n9078), .Z(n221) );
  NAND U336 ( .A(n9081), .B(n9080), .Z(n222) );
  NAND U337 ( .A(n221), .B(n222), .Z(n9087) );
  OR U338 ( .A(n9176), .B(n9175), .Z(n223) );
  NAND U339 ( .A(n9178), .B(n9177), .Z(n224) );
  NAND U340 ( .A(n223), .B(n224), .Z(n9185) );
  OR U341 ( .A(n9255), .B(n9254), .Z(n225) );
  NAND U342 ( .A(n9257), .B(n9256), .Z(n226) );
  NAND U343 ( .A(n225), .B(n226), .Z(n9263) );
  OR U344 ( .A(n9370), .B(n9369), .Z(n227) );
  NAND U345 ( .A(n9372), .B(n9371), .Z(n228) );
  NAND U346 ( .A(n227), .B(n228), .Z(n9378) );
  OR U347 ( .A(n9449), .B(n9448), .Z(n229) );
  NAND U348 ( .A(n9451), .B(n9450), .Z(n230) );
  NAND U349 ( .A(n229), .B(n230), .Z(n9457) );
  OR U350 ( .A(n9564), .B(n9563), .Z(n231) );
  NAND U351 ( .A(n9566), .B(n9565), .Z(n232) );
  NAND U352 ( .A(n231), .B(n232), .Z(n9572) );
  OR U353 ( .A(n9697), .B(n9696), .Z(n233) );
  NAND U354 ( .A(n9699), .B(n9698), .Z(n234) );
  NAND U355 ( .A(n233), .B(n234), .Z(n9705) );
  OR U356 ( .A(n9794), .B(n9793), .Z(n235) );
  NAND U357 ( .A(n9796), .B(n9795), .Z(n236) );
  NAND U358 ( .A(n235), .B(n236), .Z(n9802) );
  OR U359 ( .A(n9891), .B(n9890), .Z(n237) );
  NAND U360 ( .A(n9893), .B(n9892), .Z(n238) );
  NAND U361 ( .A(n237), .B(n238), .Z(n9899) );
  OR U362 ( .A(n10006), .B(n10005), .Z(n239) );
  NAND U363 ( .A(n10008), .B(n10007), .Z(n240) );
  NAND U364 ( .A(n239), .B(n240), .Z(n10014) );
  OR U365 ( .A(n10139), .B(n10138), .Z(n241) );
  NAND U366 ( .A(n10141), .B(n10140), .Z(n242) );
  NAND U367 ( .A(n241), .B(n242), .Z(n10147) );
  OR U368 ( .A(n10236), .B(n10235), .Z(n243) );
  NAND U369 ( .A(n10238), .B(n10237), .Z(n244) );
  NAND U370 ( .A(n243), .B(n244), .Z(n10244) );
  OR U371 ( .A(n10369), .B(n10368), .Z(n245) );
  NAND U372 ( .A(n10371), .B(n10370), .Z(n246) );
  NAND U373 ( .A(n245), .B(n246), .Z(n10377) );
  OR U374 ( .A(n10475), .B(n10474), .Z(n247) );
  NAND U375 ( .A(n10477), .B(n10476), .Z(n248) );
  NAND U376 ( .A(n247), .B(n248), .Z(n10484) );
  OR U377 ( .A(n10581), .B(n10580), .Z(n249) );
  NAND U378 ( .A(n10583), .B(n10582), .Z(n250) );
  NAND U379 ( .A(n249), .B(n250), .Z(n10589) );
  OR U380 ( .A(n10687), .B(n10686), .Z(n251) );
  NAND U381 ( .A(n10689), .B(n10688), .Z(n252) );
  NAND U382 ( .A(n251), .B(n252), .Z(n10696) );
  OR U383 ( .A(n10811), .B(n10810), .Z(n253) );
  NAND U384 ( .A(n10813), .B(n10812), .Z(n254) );
  NAND U385 ( .A(n253), .B(n254), .Z(n10819) );
  OR U386 ( .A(n10962), .B(n10961), .Z(n255) );
  NAND U387 ( .A(n10964), .B(n10963), .Z(n256) );
  NAND U388 ( .A(n255), .B(n256), .Z(n10970) );
  OR U389 ( .A(n11131), .B(n11130), .Z(n257) );
  NAND U390 ( .A(n11133), .B(n11132), .Z(n258) );
  NAND U391 ( .A(n257), .B(n258), .Z(n11139) );
  OR U392 ( .A(n11210), .B(n11209), .Z(n259) );
  NAND U393 ( .A(n11212), .B(n11211), .Z(n260) );
  NAND U394 ( .A(n259), .B(n260), .Z(n11218) );
  OR U395 ( .A(n11325), .B(n11324), .Z(n261) );
  NAND U396 ( .A(n11327), .B(n11326), .Z(n262) );
  NAND U397 ( .A(n261), .B(n262), .Z(n11333) );
  OR U398 ( .A(n11512), .B(n11511), .Z(n263) );
  NAND U399 ( .A(n11514), .B(n11513), .Z(n264) );
  NAND U400 ( .A(n263), .B(n264), .Z(n11520) );
  OR U401 ( .A(n11627), .B(n11626), .Z(n265) );
  NAND U402 ( .A(n11629), .B(n11628), .Z(n266) );
  NAND U403 ( .A(n265), .B(n266), .Z(n11635) );
  OR U404 ( .A(n11760), .B(n11759), .Z(n267) );
  NAND U405 ( .A(n11762), .B(n11761), .Z(n268) );
  NAND U406 ( .A(n267), .B(n268), .Z(n11768) );
  OR U407 ( .A(n11929), .B(n11928), .Z(n269) );
  NAND U408 ( .A(n11931), .B(n11930), .Z(n270) );
  NAND U409 ( .A(n269), .B(n270), .Z(n11937) );
  OR U410 ( .A(n12044), .B(n12043), .Z(n271) );
  NAND U411 ( .A(n12046), .B(n12045), .Z(n272) );
  NAND U412 ( .A(n271), .B(n272), .Z(n12052) );
  OR U413 ( .A(n12123), .B(n12122), .Z(n273) );
  NAND U414 ( .A(n12125), .B(n12124), .Z(n274) );
  NAND U415 ( .A(n273), .B(n274), .Z(n12131) );
  OR U416 ( .A(n12220), .B(n12219), .Z(n275) );
  NAND U417 ( .A(n12222), .B(n12221), .Z(n276) );
  NAND U418 ( .A(n275), .B(n276), .Z(n12228) );
  OR U419 ( .A(n4064), .B(n4063), .Z(n277) );
  NAND U420 ( .A(n4066), .B(n4065), .Z(n278) );
  NAND U421 ( .A(n277), .B(n278), .Z(n4072) );
  OR U422 ( .A(n4164), .B(n4163), .Z(n279) );
  NAND U423 ( .A(n4166), .B(n4165), .Z(n280) );
  NAND U424 ( .A(n279), .B(n280), .Z(n4173) );
  OR U425 ( .A(n4308), .B(n4307), .Z(n281) );
  NAND U426 ( .A(n4310), .B(n4309), .Z(n282) );
  NAND U427 ( .A(n281), .B(n282), .Z(n4316) );
  OR U428 ( .A(n4423), .B(n4422), .Z(n283) );
  NAND U429 ( .A(n4425), .B(n4424), .Z(n284) );
  NAND U430 ( .A(n283), .B(n284), .Z(n4432) );
  OR U431 ( .A(n4556), .B(n4555), .Z(n285) );
  NAND U432 ( .A(n4558), .B(n4557), .Z(n286) );
  NAND U433 ( .A(n285), .B(n286), .Z(n4564) );
  OR U434 ( .A(n4626), .B(n4625), .Z(n287) );
  NAND U435 ( .A(n4628), .B(n4627), .Z(n288) );
  NAND U436 ( .A(n287), .B(n288), .Z(n4635) );
  OR U437 ( .A(n4732), .B(n4731), .Z(n289) );
  NAND U438 ( .A(n4734), .B(n4733), .Z(n290) );
  NAND U439 ( .A(n289), .B(n290), .Z(n4740) );
  OR U440 ( .A(n4865), .B(n4864), .Z(n291) );
  NAND U441 ( .A(n4867), .B(n4866), .Z(n292) );
  NAND U442 ( .A(n291), .B(n292), .Z(n4873) );
  OR U443 ( .A(n4998), .B(n4997), .Z(n293) );
  NAND U444 ( .A(n5000), .B(n4999), .Z(n294) );
  NAND U445 ( .A(n293), .B(n294), .Z(n5006) );
  OR U446 ( .A(n5185), .B(n5184), .Z(n295) );
  NAND U447 ( .A(n5187), .B(n5186), .Z(n296) );
  NAND U448 ( .A(n295), .B(n296), .Z(n5193) );
  OR U449 ( .A(n5282), .B(n5281), .Z(n297) );
  NAND U450 ( .A(n5284), .B(n5283), .Z(n298) );
  NAND U451 ( .A(n297), .B(n298), .Z(n5290) );
  OR U452 ( .A(n5388), .B(n5387), .Z(n299) );
  NAND U453 ( .A(n5390), .B(n5389), .Z(n300) );
  NAND U454 ( .A(n299), .B(n300), .Z(n5397) );
  OR U455 ( .A(n5494), .B(n5493), .Z(n301) );
  NAND U456 ( .A(n5496), .B(n5495), .Z(n302) );
  NAND U457 ( .A(n301), .B(n302), .Z(n5502) );
  OR U458 ( .A(n5627), .B(n5626), .Z(n303) );
  NAND U459 ( .A(n5629), .B(n5628), .Z(n304) );
  NAND U460 ( .A(n303), .B(n304), .Z(n5635) );
  OR U461 ( .A(n5724), .B(n5723), .Z(n305) );
  NAND U462 ( .A(n5726), .B(n5725), .Z(n306) );
  NAND U463 ( .A(n305), .B(n306), .Z(n5732) );
  OR U464 ( .A(n5875), .B(n5874), .Z(n307) );
  NAND U465 ( .A(n5877), .B(n5876), .Z(n308) );
  NAND U466 ( .A(n307), .B(n308), .Z(n5883) );
  OR U467 ( .A(n5990), .B(n5989), .Z(n309) );
  NAND U468 ( .A(n5992), .B(n5991), .Z(n310) );
  NAND U469 ( .A(n309), .B(n310), .Z(n5998) );
  OR U470 ( .A(n6105), .B(n6104), .Z(n311) );
  NAND U471 ( .A(n6107), .B(n6106), .Z(n312) );
  NAND U472 ( .A(n311), .B(n312), .Z(n6113) );
  OR U473 ( .A(n6202), .B(n6201), .Z(n313) );
  NAND U474 ( .A(n6204), .B(n6203), .Z(n314) );
  NAND U475 ( .A(n313), .B(n314), .Z(n6211) );
  OR U476 ( .A(n6317), .B(n6316), .Z(n315) );
  NAND U477 ( .A(n6319), .B(n6318), .Z(n316) );
  NAND U478 ( .A(n315), .B(n316), .Z(n6325) );
  OR U479 ( .A(n6468), .B(n6467), .Z(n317) );
  NAND U480 ( .A(n6470), .B(n6469), .Z(n318) );
  NAND U481 ( .A(n317), .B(n318), .Z(n6476) );
  OR U482 ( .A(n6583), .B(n6582), .Z(n319) );
  NAND U483 ( .A(n6585), .B(n6584), .Z(n320) );
  NAND U484 ( .A(n319), .B(n320), .Z(n6591) );
  OR U485 ( .A(n6707), .B(n6706), .Z(n321) );
  NAND U486 ( .A(n6709), .B(n6708), .Z(n322) );
  NAND U487 ( .A(n321), .B(n322), .Z(n6716) );
  OR U488 ( .A(n6813), .B(n6812), .Z(n323) );
  NAND U489 ( .A(n6815), .B(n6814), .Z(n324) );
  NAND U490 ( .A(n323), .B(n324), .Z(n6821) );
  OR U491 ( .A(n6964), .B(n6963), .Z(n325) );
  NAND U492 ( .A(n6966), .B(n6965), .Z(n326) );
  NAND U493 ( .A(n325), .B(n326), .Z(n6973) );
  OR U494 ( .A(n7043), .B(n7042), .Z(n327) );
  NAND U495 ( .A(n7045), .B(n7044), .Z(n328) );
  NAND U496 ( .A(n327), .B(n328), .Z(n7051) );
  OR U497 ( .A(n7122), .B(n7121), .Z(n329) );
  NAND U498 ( .A(n7124), .B(n7123), .Z(n330) );
  NAND U499 ( .A(n329), .B(n330), .Z(n7130) );
  OR U500 ( .A(n7237), .B(n7236), .Z(n331) );
  NAND U501 ( .A(n7239), .B(n7238), .Z(n332) );
  NAND U502 ( .A(n331), .B(n332), .Z(n7245) );
  OR U503 ( .A(n7370), .B(n7369), .Z(n333) );
  NAND U504 ( .A(n7372), .B(n7371), .Z(n334) );
  NAND U505 ( .A(n333), .B(n334), .Z(n7379) );
  OR U506 ( .A(n7485), .B(n7484), .Z(n335) );
  NAND U507 ( .A(n7487), .B(n7486), .Z(n336) );
  NAND U508 ( .A(n335), .B(n336), .Z(n7494) );
  OR U509 ( .A(n7591), .B(n7590), .Z(n337) );
  NAND U510 ( .A(n7593), .B(n7592), .Z(n338) );
  NAND U511 ( .A(n337), .B(n338), .Z(n7600) );
  OR U512 ( .A(n7697), .B(n7696), .Z(n339) );
  NAND U513 ( .A(n7699), .B(n7698), .Z(n340) );
  NAND U514 ( .A(n339), .B(n340), .Z(n7705) );
  OR U515 ( .A(n7803), .B(n7802), .Z(n341) );
  NAND U516 ( .A(n7805), .B(n7804), .Z(n342) );
  NAND U517 ( .A(n341), .B(n342), .Z(n7812) );
  OR U518 ( .A(n7909), .B(n7908), .Z(n343) );
  NAND U519 ( .A(n7911), .B(n7910), .Z(n344) );
  NAND U520 ( .A(n343), .B(n344), .Z(n7917) );
  OR U521 ( .A(n8006), .B(n8005), .Z(n345) );
  NAND U522 ( .A(n8008), .B(n8007), .Z(n346) );
  NAND U523 ( .A(n345), .B(n346), .Z(n8015) );
  OR U524 ( .A(n8121), .B(n8120), .Z(n347) );
  NAND U525 ( .A(n8123), .B(n8122), .Z(n348) );
  NAND U526 ( .A(n347), .B(n348), .Z(n8129) );
  OR U527 ( .A(n8236), .B(n8235), .Z(n349) );
  NAND U528 ( .A(n8238), .B(n8237), .Z(n350) );
  NAND U529 ( .A(n349), .B(n350), .Z(n8244) );
  OR U530 ( .A(n8333), .B(n8332), .Z(n351) );
  NAND U531 ( .A(n8335), .B(n8334), .Z(n352) );
  NAND U532 ( .A(n351), .B(n352), .Z(n8341) );
  OR U533 ( .A(n8430), .B(n8429), .Z(n353) );
  NAND U534 ( .A(n8432), .B(n8431), .Z(n354) );
  NAND U535 ( .A(n353), .B(n354), .Z(n8438) );
  OR U536 ( .A(n8599), .B(n8598), .Z(n355) );
  NAND U537 ( .A(n8601), .B(n8600), .Z(n356) );
  NAND U538 ( .A(n355), .B(n356), .Z(n8607) );
  OR U539 ( .A(n8696), .B(n8695), .Z(n357) );
  NAND U540 ( .A(n8698), .B(n8697), .Z(n358) );
  NAND U541 ( .A(n357), .B(n358), .Z(n8704) );
  OR U542 ( .A(n8811), .B(n8810), .Z(n359) );
  NAND U543 ( .A(n8813), .B(n8812), .Z(n360) );
  NAND U544 ( .A(n359), .B(n360), .Z(n8820) );
  OR U545 ( .A(n8944), .B(n8943), .Z(n361) );
  NAND U546 ( .A(n8946), .B(n8945), .Z(n362) );
  NAND U547 ( .A(n361), .B(n362), .Z(n8953) );
  OR U548 ( .A(n9095), .B(n9094), .Z(n363) );
  NAND U549 ( .A(n9097), .B(n9096), .Z(n364) );
  NAND U550 ( .A(n363), .B(n364), .Z(n9103) );
  OR U551 ( .A(n9183), .B(n9182), .Z(n365) );
  NAND U552 ( .A(n9185), .B(n9184), .Z(n366) );
  NAND U553 ( .A(n365), .B(n366), .Z(n9192) );
  OR U554 ( .A(n9289), .B(n9288), .Z(n367) );
  NAND U555 ( .A(n9291), .B(n9290), .Z(n368) );
  NAND U556 ( .A(n367), .B(n368), .Z(n9297) );
  OR U557 ( .A(n9386), .B(n9385), .Z(n369) );
  NAND U558 ( .A(n9388), .B(n9387), .Z(n370) );
  NAND U559 ( .A(n369), .B(n370), .Z(n9394) );
  OR U560 ( .A(n9465), .B(n9464), .Z(n371) );
  NAND U561 ( .A(n9467), .B(n9466), .Z(n372) );
  NAND U562 ( .A(n371), .B(n372), .Z(n9473) );
  OR U563 ( .A(n9580), .B(n9579), .Z(n373) );
  NAND U564 ( .A(n9582), .B(n9581), .Z(n374) );
  NAND U565 ( .A(n373), .B(n374), .Z(n9588) );
  OR U566 ( .A(n9713), .B(n9712), .Z(n375) );
  NAND U567 ( .A(n9715), .B(n9714), .Z(n376) );
  NAND U568 ( .A(n375), .B(n376), .Z(n9721) );
  OR U569 ( .A(n9810), .B(n9809), .Z(n377) );
  NAND U570 ( .A(n9812), .B(n9811), .Z(n378) );
  NAND U571 ( .A(n377), .B(n378), .Z(n9819) );
  OR U572 ( .A(n9907), .B(n9906), .Z(n379) );
  NAND U573 ( .A(n9909), .B(n9908), .Z(n380) );
  NAND U574 ( .A(n379), .B(n380), .Z(n9915) );
  OR U575 ( .A(n10022), .B(n10021), .Z(n381) );
  NAND U576 ( .A(n10024), .B(n10023), .Z(n382) );
  NAND U577 ( .A(n381), .B(n382), .Z(n10030) );
  OR U578 ( .A(n10155), .B(n10154), .Z(n383) );
  NAND U579 ( .A(n10157), .B(n10156), .Z(n384) );
  NAND U580 ( .A(n383), .B(n384), .Z(n10163) );
  OR U581 ( .A(n10252), .B(n10251), .Z(n385) );
  NAND U582 ( .A(n10254), .B(n10253), .Z(n386) );
  NAND U583 ( .A(n385), .B(n386), .Z(n10260) );
  OR U584 ( .A(n10385), .B(n10384), .Z(n387) );
  NAND U585 ( .A(n10387), .B(n10386), .Z(n388) );
  NAND U586 ( .A(n387), .B(n388), .Z(n10393) );
  OR U587 ( .A(n10482), .B(n10481), .Z(n389) );
  NAND U588 ( .A(n10484), .B(n10483), .Z(n390) );
  NAND U589 ( .A(n389), .B(n390), .Z(n10490) );
  OR U590 ( .A(n10597), .B(n10596), .Z(n391) );
  NAND U591 ( .A(n10599), .B(n10598), .Z(n392) );
  NAND U592 ( .A(n391), .B(n392), .Z(n10605) );
  OR U593 ( .A(n10694), .B(n10693), .Z(n393) );
  NAND U594 ( .A(n10696), .B(n10695), .Z(n394) );
  NAND U595 ( .A(n393), .B(n394), .Z(n10702) );
  OR U596 ( .A(n10827), .B(n10826), .Z(n395) );
  NAND U597 ( .A(n10829), .B(n10828), .Z(n396) );
  NAND U598 ( .A(n395), .B(n396), .Z(n10835) );
  OR U599 ( .A(n10978), .B(n10977), .Z(n397) );
  NAND U600 ( .A(n10980), .B(n10979), .Z(n398) );
  NAND U601 ( .A(n397), .B(n398), .Z(n10987) );
  OR U602 ( .A(n11147), .B(n11146), .Z(n399) );
  NAND U603 ( .A(n11149), .B(n11148), .Z(n400) );
  NAND U604 ( .A(n399), .B(n400), .Z(n11155) );
  OR U605 ( .A(n11226), .B(n11225), .Z(n401) );
  NAND U606 ( .A(n11228), .B(n11227), .Z(n402) );
  NAND U607 ( .A(n401), .B(n402), .Z(n11234) );
  OR U608 ( .A(n11341), .B(n11340), .Z(n403) );
  NAND U609 ( .A(n11343), .B(n11342), .Z(n404) );
  NAND U610 ( .A(n403), .B(n404), .Z(n11349) );
  OR U611 ( .A(n11528), .B(n11527), .Z(n405) );
  NAND U612 ( .A(n11530), .B(n11529), .Z(n406) );
  NAND U613 ( .A(n405), .B(n406), .Z(n11537) );
  OR U614 ( .A(n11643), .B(n11642), .Z(n407) );
  NAND U615 ( .A(n11645), .B(n11644), .Z(n408) );
  NAND U616 ( .A(n407), .B(n408), .Z(n11651) );
  OR U617 ( .A(n11830), .B(n11829), .Z(n409) );
  NAND U618 ( .A(n11832), .B(n11831), .Z(n410) );
  NAND U619 ( .A(n409), .B(n410), .Z(n11838) );
  OR U620 ( .A(n11945), .B(n11944), .Z(n411) );
  NAND U621 ( .A(n11947), .B(n11946), .Z(n412) );
  NAND U622 ( .A(n411), .B(n412), .Z(n11953) );
  OR U623 ( .A(n12060), .B(n12059), .Z(n413) );
  NAND U624 ( .A(n12062), .B(n12061), .Z(n414) );
  NAND U625 ( .A(n413), .B(n414), .Z(n12068) );
  OR U626 ( .A(n12139), .B(n12138), .Z(n415) );
  NAND U627 ( .A(n12141), .B(n12140), .Z(n416) );
  NAND U628 ( .A(n415), .B(n416), .Z(n12147) );
  OR U629 ( .A(n12254), .B(n12253), .Z(n417) );
  NAND U630 ( .A(n12256), .B(n12255), .Z(n418) );
  NAND U631 ( .A(n417), .B(n418), .Z(n12262) );
  OR U632 ( .A(n12336), .B(n12335), .Z(n419) );
  NAND U633 ( .A(n12338), .B(n12337), .Z(n420) );
  NAND U634 ( .A(n419), .B(n420), .Z(n12344) );
  OR U635 ( .A(n4089), .B(n4088), .Z(n421) );
  NAND U636 ( .A(n4091), .B(n4090), .Z(n422) );
  NAND U637 ( .A(n421), .B(n422), .Z(n4097) );
  OR U638 ( .A(n4171), .B(n4170), .Z(n423) );
  NAND U639 ( .A(n4173), .B(n4172), .Z(n424) );
  NAND U640 ( .A(n423), .B(n424), .Z(n4179) );
  OR U641 ( .A(n4324), .B(n4323), .Z(n425) );
  NAND U642 ( .A(n4326), .B(n4325), .Z(n426) );
  NAND U643 ( .A(n425), .B(n426), .Z(n4332) );
  OR U644 ( .A(n4430), .B(n4429), .Z(n427) );
  NAND U645 ( .A(n4432), .B(n4431), .Z(n428) );
  NAND U646 ( .A(n427), .B(n428), .Z(n4439) );
  OR U647 ( .A(n4572), .B(n4571), .Z(n429) );
  NAND U648 ( .A(n4574), .B(n4573), .Z(n430) );
  NAND U649 ( .A(n429), .B(n430), .Z(n4581) );
  OR U650 ( .A(n4633), .B(n4632), .Z(n431) );
  NAND U651 ( .A(n4635), .B(n4634), .Z(n432) );
  NAND U652 ( .A(n431), .B(n432), .Z(n4641) );
  OR U653 ( .A(n4748), .B(n4747), .Z(n433) );
  NAND U654 ( .A(n4750), .B(n4749), .Z(n434) );
  NAND U655 ( .A(n433), .B(n434), .Z(n4756) );
  OR U656 ( .A(n4890), .B(n4889), .Z(n435) );
  NAND U657 ( .A(n4892), .B(n4891), .Z(n436) );
  NAND U658 ( .A(n435), .B(n436), .Z(n4899) );
  OR U659 ( .A(n5032), .B(n5031), .Z(n437) );
  NAND U660 ( .A(n5034), .B(n5033), .Z(n438) );
  NAND U661 ( .A(n437), .B(n438), .Z(n5040) );
  OR U662 ( .A(n5201), .B(n5200), .Z(n439) );
  NAND U663 ( .A(n5203), .B(n5202), .Z(n440) );
  NAND U664 ( .A(n439), .B(n440), .Z(n5209) );
  OR U665 ( .A(n5298), .B(n5297), .Z(n441) );
  NAND U666 ( .A(n5300), .B(n5299), .Z(n442) );
  NAND U667 ( .A(n441), .B(n442), .Z(n5306) );
  OR U668 ( .A(n5395), .B(n5394), .Z(n443) );
  NAND U669 ( .A(n5397), .B(n5396), .Z(n444) );
  NAND U670 ( .A(n443), .B(n444), .Z(n5404) );
  OR U671 ( .A(n5510), .B(n5509), .Z(n445) );
  NAND U672 ( .A(n5512), .B(n5511), .Z(n446) );
  NAND U673 ( .A(n445), .B(n446), .Z(n5518) );
  OR U674 ( .A(n5643), .B(n5642), .Z(n447) );
  NAND U675 ( .A(n5645), .B(n5644), .Z(n448) );
  NAND U676 ( .A(n447), .B(n448), .Z(n5652) );
  OR U677 ( .A(n5740), .B(n5739), .Z(n449) );
  NAND U678 ( .A(n5742), .B(n5741), .Z(n450) );
  NAND U679 ( .A(n449), .B(n450), .Z(n5748) );
  OR U680 ( .A(n5891), .B(n5890), .Z(n451) );
  NAND U681 ( .A(n5893), .B(n5892), .Z(n452) );
  NAND U682 ( .A(n451), .B(n452), .Z(n5899) );
  OR U683 ( .A(n6006), .B(n6005), .Z(n453) );
  NAND U684 ( .A(n6008), .B(n6007), .Z(n454) );
  NAND U685 ( .A(n453), .B(n454), .Z(n6014) );
  OR U686 ( .A(n6121), .B(n6120), .Z(n455) );
  NAND U687 ( .A(n6123), .B(n6122), .Z(n456) );
  NAND U688 ( .A(n455), .B(n456), .Z(n6130) );
  OR U689 ( .A(n6209), .B(n6208), .Z(n457) );
  NAND U690 ( .A(n6211), .B(n6210), .Z(n458) );
  NAND U691 ( .A(n457), .B(n458), .Z(n6218) );
  OR U692 ( .A(n6333), .B(n6332), .Z(n459) );
  NAND U693 ( .A(n6335), .B(n6334), .Z(n460) );
  NAND U694 ( .A(n459), .B(n460), .Z(n6341) );
  OR U695 ( .A(n6484), .B(n6483), .Z(n461) );
  NAND U696 ( .A(n6486), .B(n6485), .Z(n462) );
  NAND U697 ( .A(n461), .B(n462), .Z(n6492) );
  OR U698 ( .A(n6599), .B(n6598), .Z(n463) );
  NAND U699 ( .A(n6601), .B(n6600), .Z(n464) );
  NAND U700 ( .A(n463), .B(n464), .Z(n6607) );
  OR U701 ( .A(n6714), .B(n6713), .Z(n465) );
  NAND U702 ( .A(n6716), .B(n6715), .Z(n466) );
  NAND U703 ( .A(n465), .B(n466), .Z(n6722) );
  OR U704 ( .A(n6847), .B(n6846), .Z(n467) );
  NAND U705 ( .A(n6849), .B(n6848), .Z(n468) );
  NAND U706 ( .A(n467), .B(n468), .Z(n6855) );
  OR U707 ( .A(n6971), .B(n6970), .Z(n469) );
  NAND U708 ( .A(n6973), .B(n6972), .Z(n470) );
  NAND U709 ( .A(n469), .B(n470), .Z(n6980) );
  OR U710 ( .A(n7059), .B(n7058), .Z(n471) );
  NAND U711 ( .A(n7061), .B(n7060), .Z(n472) );
  NAND U712 ( .A(n471), .B(n472), .Z(n7068) );
  OR U713 ( .A(n7138), .B(n7137), .Z(n473) );
  NAND U714 ( .A(n7140), .B(n7139), .Z(n474) );
  NAND U715 ( .A(n473), .B(n474), .Z(n7146) );
  OR U716 ( .A(n7253), .B(n7252), .Z(n475) );
  NAND U717 ( .A(n7255), .B(n7254), .Z(n476) );
  NAND U718 ( .A(n475), .B(n476), .Z(n7261) );
  OR U719 ( .A(n7377), .B(n7376), .Z(n477) );
  NAND U720 ( .A(n7379), .B(n7378), .Z(n478) );
  NAND U721 ( .A(n477), .B(n478), .Z(n7385) );
  OR U722 ( .A(n7492), .B(n7491), .Z(n479) );
  NAND U723 ( .A(n7494), .B(n7493), .Z(n480) );
  NAND U724 ( .A(n479), .B(n480), .Z(n7501) );
  OR U725 ( .A(n7598), .B(n7597), .Z(n481) );
  NAND U726 ( .A(n7600), .B(n7599), .Z(n482) );
  NAND U727 ( .A(n481), .B(n482), .Z(n7606) );
  OR U728 ( .A(n7713), .B(n7712), .Z(n483) );
  NAND U729 ( .A(n7715), .B(n7714), .Z(n484) );
  NAND U730 ( .A(n483), .B(n484), .Z(n7721) );
  OR U731 ( .A(n7810), .B(n7809), .Z(n485) );
  NAND U732 ( .A(n7812), .B(n7811), .Z(n486) );
  NAND U733 ( .A(n485), .B(n486), .Z(n7818) );
  OR U734 ( .A(n7925), .B(n7924), .Z(n487) );
  NAND U735 ( .A(n7927), .B(n7926), .Z(n488) );
  NAND U736 ( .A(n487), .B(n488), .Z(n7933) );
  OR U737 ( .A(n8013), .B(n8012), .Z(n489) );
  NAND U738 ( .A(n8015), .B(n8014), .Z(n490) );
  NAND U739 ( .A(n489), .B(n490), .Z(n8021) );
  OR U740 ( .A(n8137), .B(n8136), .Z(n491) );
  NAND U741 ( .A(n8139), .B(n8138), .Z(n492) );
  NAND U742 ( .A(n491), .B(n492), .Z(n8145) );
  OR U743 ( .A(n8252), .B(n8251), .Z(n493) );
  NAND U744 ( .A(n8254), .B(n8253), .Z(n494) );
  NAND U745 ( .A(n493), .B(n494), .Z(n8261) );
  OR U746 ( .A(n8349), .B(n8348), .Z(n495) );
  NAND U747 ( .A(n8351), .B(n8350), .Z(n496) );
  NAND U748 ( .A(n495), .B(n496), .Z(n8357) );
  OR U749 ( .A(n8446), .B(n8445), .Z(n497) );
  NAND U750 ( .A(n8448), .B(n8447), .Z(n498) );
  NAND U751 ( .A(n497), .B(n498), .Z(n8454) );
  OR U752 ( .A(n8615), .B(n8614), .Z(n499) );
  NAND U753 ( .A(n8617), .B(n8616), .Z(n500) );
  NAND U754 ( .A(n499), .B(n500), .Z(n8623) );
  OR U755 ( .A(n8712), .B(n8711), .Z(n501) );
  NAND U756 ( .A(n8714), .B(n8713), .Z(n502) );
  NAND U757 ( .A(n501), .B(n502), .Z(n8720) );
  OR U758 ( .A(n8818), .B(n8817), .Z(n503) );
  NAND U759 ( .A(n8820), .B(n8819), .Z(n504) );
  NAND U760 ( .A(n503), .B(n504), .Z(n8826) );
  OR U761 ( .A(n8951), .B(n8950), .Z(n505) );
  NAND U762 ( .A(n8953), .B(n8952), .Z(n506) );
  NAND U763 ( .A(n505), .B(n506), .Z(n8960) );
  OR U764 ( .A(n9111), .B(n9110), .Z(n507) );
  NAND U765 ( .A(n9113), .B(n9112), .Z(n508) );
  NAND U766 ( .A(n507), .B(n508), .Z(n9120) );
  OR U767 ( .A(n9190), .B(n9189), .Z(n509) );
  NAND U768 ( .A(n9192), .B(n9191), .Z(n510) );
  NAND U769 ( .A(n509), .B(n510), .Z(n9198) );
  OR U770 ( .A(n9305), .B(n9304), .Z(n511) );
  NAND U771 ( .A(n9307), .B(n9306), .Z(n512) );
  NAND U772 ( .A(n511), .B(n512), .Z(n9313) );
  OR U773 ( .A(n9402), .B(n9401), .Z(n513) );
  NAND U774 ( .A(n9404), .B(n9403), .Z(n514) );
  NAND U775 ( .A(n513), .B(n514), .Z(n9411) );
  OR U776 ( .A(n9481), .B(n9480), .Z(n515) );
  NAND U777 ( .A(n9483), .B(n9482), .Z(n516) );
  NAND U778 ( .A(n515), .B(n516), .Z(n9489) );
  OR U779 ( .A(n9596), .B(n9595), .Z(n517) );
  NAND U780 ( .A(n9598), .B(n9597), .Z(n518) );
  NAND U781 ( .A(n517), .B(n518), .Z(n9604) );
  OR U782 ( .A(n9729), .B(n9728), .Z(n519) );
  NAND U783 ( .A(n9731), .B(n9730), .Z(n520) );
  NAND U784 ( .A(n519), .B(n520), .Z(n9738) );
  OR U785 ( .A(n9817), .B(n9816), .Z(n521) );
  NAND U786 ( .A(n9819), .B(n9818), .Z(n522) );
  NAND U787 ( .A(n521), .B(n522), .Z(n9826) );
  OR U788 ( .A(n9923), .B(n9922), .Z(n523) );
  NAND U789 ( .A(n9925), .B(n9924), .Z(n524) );
  NAND U790 ( .A(n523), .B(n524), .Z(n9931) );
  OR U791 ( .A(n10056), .B(n10055), .Z(n525) );
  NAND U792 ( .A(n10058), .B(n10057), .Z(n526) );
  NAND U793 ( .A(n525), .B(n526), .Z(n10064) );
  OR U794 ( .A(n10171), .B(n10170), .Z(n527) );
  NAND U795 ( .A(n10173), .B(n10172), .Z(n528) );
  NAND U796 ( .A(n527), .B(n528), .Z(n10179) );
  OR U797 ( .A(n10268), .B(n10267), .Z(n529) );
  NAND U798 ( .A(n10270), .B(n10269), .Z(n530) );
  NAND U799 ( .A(n529), .B(n530), .Z(n10276) );
  OR U800 ( .A(n10401), .B(n10400), .Z(n531) );
  NAND U801 ( .A(n10403), .B(n10402), .Z(n532) );
  NAND U802 ( .A(n531), .B(n532), .Z(n10409) );
  OR U803 ( .A(n10498), .B(n10497), .Z(n533) );
  NAND U804 ( .A(n10500), .B(n10499), .Z(n534) );
  NAND U805 ( .A(n533), .B(n534), .Z(n10506) );
  OR U806 ( .A(n10613), .B(n10612), .Z(n535) );
  NAND U807 ( .A(n10615), .B(n10614), .Z(n536) );
  NAND U808 ( .A(n535), .B(n536), .Z(n10622) );
  OR U809 ( .A(n10710), .B(n10709), .Z(n537) );
  NAND U810 ( .A(n10712), .B(n10711), .Z(n538) );
  NAND U811 ( .A(n537), .B(n538), .Z(n10718) );
  OR U812 ( .A(n10843), .B(n10842), .Z(n539) );
  NAND U813 ( .A(n10845), .B(n10844), .Z(n540) );
  NAND U814 ( .A(n539), .B(n540), .Z(n10851) );
  OR U815 ( .A(n10985), .B(n10984), .Z(n541) );
  NAND U816 ( .A(n10987), .B(n10986), .Z(n542) );
  NAND U817 ( .A(n541), .B(n542), .Z(n10994) );
  OR U818 ( .A(n11163), .B(n11162), .Z(n543) );
  NAND U819 ( .A(n11165), .B(n11164), .Z(n544) );
  NAND U820 ( .A(n543), .B(n544), .Z(n11172) );
  OR U821 ( .A(n11242), .B(n11241), .Z(n545) );
  NAND U822 ( .A(n11244), .B(n11243), .Z(n546) );
  NAND U823 ( .A(n545), .B(n546), .Z(n11250) );
  OR U824 ( .A(n11393), .B(n11392), .Z(n547) );
  NAND U825 ( .A(n11395), .B(n11394), .Z(n548) );
  NAND U826 ( .A(n547), .B(n548), .Z(n11401) );
  OR U827 ( .A(n11535), .B(n11534), .Z(n549) );
  NAND U828 ( .A(n11537), .B(n11536), .Z(n550) );
  NAND U829 ( .A(n549), .B(n550), .Z(n11544) );
  OR U830 ( .A(n11677), .B(n11676), .Z(n551) );
  NAND U831 ( .A(n11679), .B(n11678), .Z(n552) );
  NAND U832 ( .A(n551), .B(n552), .Z(n11685) );
  OR U833 ( .A(n11846), .B(n11845), .Z(n553) );
  NAND U834 ( .A(n11848), .B(n11847), .Z(n554) );
  NAND U835 ( .A(n553), .B(n554), .Z(n11854) );
  OR U836 ( .A(n11961), .B(n11960), .Z(n555) );
  NAND U837 ( .A(n11963), .B(n11962), .Z(n556) );
  NAND U838 ( .A(n555), .B(n556), .Z(n11969) );
  OR U839 ( .A(n12076), .B(n12075), .Z(n557) );
  NAND U840 ( .A(n12078), .B(n12077), .Z(n558) );
  NAND U841 ( .A(n557), .B(n558), .Z(n12085) );
  OR U842 ( .A(n12155), .B(n12154), .Z(n559) );
  NAND U843 ( .A(n12157), .B(n12156), .Z(n560) );
  NAND U844 ( .A(n559), .B(n560), .Z(n12163) );
  OR U845 ( .A(n12270), .B(n12269), .Z(n561) );
  NAND U846 ( .A(n12272), .B(n12271), .Z(n562) );
  NAND U847 ( .A(n561), .B(n562), .Z(n12279) );
  OR U848 ( .A(n12352), .B(n12351), .Z(n563) );
  NAND U849 ( .A(n12354), .B(n12353), .Z(n564) );
  NAND U850 ( .A(n563), .B(n564), .Z(n12360) );
  OR U851 ( .A(n4105), .B(n4104), .Z(n565) );
  NAND U852 ( .A(n4107), .B(n4106), .Z(n566) );
  NAND U853 ( .A(n565), .B(n566), .Z(n4113) );
  OR U854 ( .A(n4225), .B(n4224), .Z(n567) );
  NAND U855 ( .A(n4227), .B(n4226), .Z(n568) );
  NAND U856 ( .A(n567), .B(n568), .Z(n4233) );
  OR U857 ( .A(n4340), .B(n4339), .Z(n569) );
  NAND U858 ( .A(n4342), .B(n4341), .Z(n570) );
  NAND U859 ( .A(n569), .B(n570), .Z(n4349) );
  OR U860 ( .A(n4437), .B(n4436), .Z(n571) );
  NAND U861 ( .A(n4439), .B(n4438), .Z(n572) );
  NAND U862 ( .A(n571), .B(n572), .Z(n4445) );
  OR U863 ( .A(n4579), .B(n4578), .Z(n573) );
  NAND U864 ( .A(n4581), .B(n4580), .Z(n574) );
  NAND U865 ( .A(n573), .B(n574), .Z(n4588) );
  OR U866 ( .A(n4649), .B(n4648), .Z(n575) );
  NAND U867 ( .A(n4651), .B(n4650), .Z(n576) );
  NAND U868 ( .A(n575), .B(n576), .Z(n4657) );
  OR U869 ( .A(n4764), .B(n4763), .Z(n577) );
  NAND U870 ( .A(n4766), .B(n4765), .Z(n578) );
  NAND U871 ( .A(n577), .B(n578), .Z(n4772) );
  OR U872 ( .A(n4897), .B(n4896), .Z(n579) );
  NAND U873 ( .A(n4899), .B(n4898), .Z(n580) );
  NAND U874 ( .A(n579), .B(n580), .Z(n4906) );
  OR U875 ( .A(n5048), .B(n5047), .Z(n581) );
  NAND U876 ( .A(n5050), .B(n5049), .Z(n582) );
  NAND U877 ( .A(n581), .B(n582), .Z(n5056) );
  OR U878 ( .A(n5217), .B(n5216), .Z(n583) );
  NAND U879 ( .A(n5219), .B(n5218), .Z(n584) );
  NAND U880 ( .A(n583), .B(n584), .Z(n5226) );
  OR U881 ( .A(n5314), .B(n5313), .Z(n585) );
  NAND U882 ( .A(n5316), .B(n5315), .Z(n586) );
  NAND U883 ( .A(n585), .B(n586), .Z(n5322) );
  OR U884 ( .A(n5402), .B(n5401), .Z(n587) );
  NAND U885 ( .A(n5404), .B(n5403), .Z(n588) );
  NAND U886 ( .A(n587), .B(n588), .Z(n5411) );
  OR U887 ( .A(n5526), .B(n5525), .Z(n589) );
  NAND U888 ( .A(n5528), .B(n5527), .Z(n590) );
  NAND U889 ( .A(n589), .B(n590), .Z(n5534) );
  OR U890 ( .A(n5650), .B(n5649), .Z(n591) );
  NAND U891 ( .A(n5652), .B(n5651), .Z(n592) );
  NAND U892 ( .A(n591), .B(n592), .Z(n5659) );
  OR U893 ( .A(n5774), .B(n5773), .Z(n593) );
  NAND U894 ( .A(n5776), .B(n5775), .Z(n594) );
  NAND U895 ( .A(n593), .B(n594), .Z(n5782) );
  OR U896 ( .A(n5907), .B(n5906), .Z(n595) );
  NAND U897 ( .A(n5909), .B(n5908), .Z(n596) );
  NAND U898 ( .A(n595), .B(n596), .Z(n5915) );
  OR U899 ( .A(n6022), .B(n6021), .Z(n597) );
  NAND U900 ( .A(n6024), .B(n6023), .Z(n598) );
  NAND U901 ( .A(n597), .B(n598), .Z(n6030) );
  OR U902 ( .A(n6128), .B(n6127), .Z(n599) );
  NAND U903 ( .A(n6130), .B(n6129), .Z(n600) );
  NAND U904 ( .A(n599), .B(n600), .Z(n6137) );
  OR U905 ( .A(n6216), .B(n6215), .Z(n601) );
  NAND U906 ( .A(n6218), .B(n6217), .Z(n602) );
  NAND U907 ( .A(n601), .B(n602), .Z(n6224) );
  OR U908 ( .A(n6367), .B(n6366), .Z(n603) );
  NAND U909 ( .A(n6369), .B(n6368), .Z(n604) );
  NAND U910 ( .A(n603), .B(n604), .Z(n6375) );
  OR U911 ( .A(n6500), .B(n6499), .Z(n605) );
  NAND U912 ( .A(n6502), .B(n6501), .Z(n606) );
  NAND U913 ( .A(n605), .B(n606), .Z(n6508) );
  OR U914 ( .A(n6615), .B(n6614), .Z(n607) );
  NAND U915 ( .A(n6617), .B(n6616), .Z(n608) );
  NAND U916 ( .A(n607), .B(n608), .Z(n6623) );
  OR U917 ( .A(n6730), .B(n6729), .Z(n609) );
  NAND U918 ( .A(n6732), .B(n6731), .Z(n610) );
  NAND U919 ( .A(n609), .B(n610), .Z(n6739) );
  OR U920 ( .A(n6863), .B(n6862), .Z(n611) );
  NAND U921 ( .A(n6865), .B(n6864), .Z(n612) );
  NAND U922 ( .A(n611), .B(n612), .Z(n6871) );
  OR U923 ( .A(n6978), .B(n6977), .Z(n613) );
  NAND U924 ( .A(n6980), .B(n6979), .Z(n614) );
  NAND U925 ( .A(n613), .B(n614), .Z(n6986) );
  OR U926 ( .A(n7066), .B(n7065), .Z(n615) );
  NAND U927 ( .A(n7068), .B(n7067), .Z(n616) );
  NAND U928 ( .A(n615), .B(n616), .Z(n7075) );
  OR U929 ( .A(n7154), .B(n7153), .Z(n617) );
  NAND U930 ( .A(n7156), .B(n7155), .Z(n618) );
  NAND U931 ( .A(n617), .B(n618), .Z(n7162) );
  OR U932 ( .A(n7269), .B(n7268), .Z(n619) );
  NAND U933 ( .A(n7271), .B(n7270), .Z(n620) );
  NAND U934 ( .A(n619), .B(n620), .Z(n7277) );
  OR U935 ( .A(n7402), .B(n7401), .Z(n621) );
  NAND U936 ( .A(n7404), .B(n7403), .Z(n622) );
  NAND U937 ( .A(n621), .B(n622), .Z(n7410) );
  OR U938 ( .A(n7499), .B(n7498), .Z(n623) );
  NAND U939 ( .A(n7501), .B(n7500), .Z(n624) );
  NAND U940 ( .A(n623), .B(n624), .Z(n7508) );
  OR U941 ( .A(n7614), .B(n7613), .Z(n625) );
  NAND U942 ( .A(n7616), .B(n7615), .Z(n626) );
  NAND U943 ( .A(n625), .B(n626), .Z(n7622) );
  OR U944 ( .A(n7747), .B(n7746), .Z(n627) );
  NAND U945 ( .A(n7749), .B(n7748), .Z(n628) );
  NAND U946 ( .A(n627), .B(n628), .Z(n7755) );
  OR U947 ( .A(n7826), .B(n7825), .Z(n629) );
  NAND U948 ( .A(n7828), .B(n7827), .Z(n630) );
  NAND U949 ( .A(n629), .B(n630), .Z(n7834) );
  OR U950 ( .A(n7941), .B(n7940), .Z(n631) );
  NAND U951 ( .A(n7943), .B(n7942), .Z(n632) );
  NAND U952 ( .A(n631), .B(n632), .Z(n7949) );
  OR U953 ( .A(n8029), .B(n8028), .Z(n633) );
  NAND U954 ( .A(n8031), .B(n8030), .Z(n634) );
  NAND U955 ( .A(n633), .B(n634), .Z(n8037) );
  OR U956 ( .A(n8153), .B(n8152), .Z(n635) );
  NAND U957 ( .A(n8155), .B(n8154), .Z(n636) );
  NAND U958 ( .A(n635), .B(n636), .Z(n8161) );
  OR U959 ( .A(n8259), .B(n8258), .Z(n637) );
  NAND U960 ( .A(n8261), .B(n8260), .Z(n638) );
  NAND U961 ( .A(n637), .B(n638), .Z(n8268) );
  OR U962 ( .A(n8365), .B(n8364), .Z(n639) );
  NAND U963 ( .A(n8367), .B(n8366), .Z(n640) );
  NAND U964 ( .A(n639), .B(n640), .Z(n8373) );
  OR U965 ( .A(n8462), .B(n8461), .Z(n641) );
  NAND U966 ( .A(n8464), .B(n8463), .Z(n642) );
  NAND U967 ( .A(n641), .B(n642), .Z(n8470) );
  OR U968 ( .A(n8631), .B(n8630), .Z(n643) );
  NAND U969 ( .A(n8633), .B(n8632), .Z(n644) );
  NAND U970 ( .A(n643), .B(n644), .Z(n8640) );
  OR U971 ( .A(n8728), .B(n8727), .Z(n645) );
  NAND U972 ( .A(n8730), .B(n8729), .Z(n646) );
  NAND U973 ( .A(n645), .B(n646), .Z(n8736) );
  OR U974 ( .A(n8843), .B(n8842), .Z(n647) );
  NAND U975 ( .A(n8845), .B(n8844), .Z(n648) );
  NAND U976 ( .A(n647), .B(n648), .Z(n8851) );
  OR U977 ( .A(n8958), .B(n8957), .Z(n649) );
  NAND U978 ( .A(n8960), .B(n8959), .Z(n650) );
  NAND U979 ( .A(n649), .B(n650), .Z(n8966) );
  OR U980 ( .A(n9118), .B(n9117), .Z(n651) );
  NAND U981 ( .A(n9120), .B(n9119), .Z(n652) );
  NAND U982 ( .A(n651), .B(n652), .Z(n9127) );
  OR U983 ( .A(n9206), .B(n9205), .Z(n653) );
  NAND U984 ( .A(n9208), .B(n9207), .Z(n654) );
  NAND U985 ( .A(n653), .B(n654), .Z(n9215) );
  OR U986 ( .A(n9321), .B(n9320), .Z(n655) );
  NAND U987 ( .A(n9323), .B(n9322), .Z(n656) );
  NAND U988 ( .A(n655), .B(n656), .Z(n9330) );
  OR U989 ( .A(n9409), .B(n9408), .Z(n657) );
  NAND U990 ( .A(n9411), .B(n9410), .Z(n658) );
  NAND U991 ( .A(n657), .B(n658), .Z(n9418) );
  OR U992 ( .A(n9515), .B(n9514), .Z(n659) );
  NAND U993 ( .A(n9517), .B(n9516), .Z(n660) );
  NAND U994 ( .A(n659), .B(n660), .Z(n9523) );
  OR U995 ( .A(n9630), .B(n9629), .Z(n661) );
  NAND U996 ( .A(n9632), .B(n9631), .Z(n662) );
  NAND U997 ( .A(n661), .B(n662), .Z(n9638) );
  OR U998 ( .A(n9736), .B(n9735), .Z(n663) );
  NAND U999 ( .A(n9738), .B(n9737), .Z(n664) );
  NAND U1000 ( .A(n663), .B(n664), .Z(n9745) );
  OR U1001 ( .A(n9824), .B(n9823), .Z(n665) );
  NAND U1002 ( .A(n9826), .B(n9825), .Z(n666) );
  NAND U1003 ( .A(n665), .B(n666), .Z(n9832) );
  OR U1004 ( .A(n9939), .B(n9938), .Z(n667) );
  NAND U1005 ( .A(n9941), .B(n9940), .Z(n668) );
  NAND U1006 ( .A(n667), .B(n668), .Z(n9947) );
  OR U1007 ( .A(n10072), .B(n10071), .Z(n669) );
  NAND U1008 ( .A(n10074), .B(n10073), .Z(n670) );
  NAND U1009 ( .A(n669), .B(n670), .Z(n10080) );
  OR U1010 ( .A(n10187), .B(n10186), .Z(n671) );
  NAND U1011 ( .A(n10189), .B(n10188), .Z(n672) );
  NAND U1012 ( .A(n671), .B(n672), .Z(n10196) );
  OR U1013 ( .A(n10284), .B(n10283), .Z(n673) );
  NAND U1014 ( .A(n10286), .B(n10285), .Z(n674) );
  NAND U1015 ( .A(n673), .B(n674), .Z(n10292) );
  OR U1016 ( .A(n10417), .B(n10416), .Z(n675) );
  NAND U1017 ( .A(n10419), .B(n10418), .Z(n676) );
  NAND U1018 ( .A(n675), .B(n676), .Z(n10425) );
  OR U1019 ( .A(n10514), .B(n10513), .Z(n677) );
  NAND U1020 ( .A(n10516), .B(n10515), .Z(n678) );
  NAND U1021 ( .A(n677), .B(n678), .Z(n10522) );
  OR U1022 ( .A(n10620), .B(n10619), .Z(n679) );
  NAND U1023 ( .A(n10622), .B(n10621), .Z(n680) );
  NAND U1024 ( .A(n679), .B(n680), .Z(n10629) );
  OR U1025 ( .A(n10726), .B(n10725), .Z(n681) );
  NAND U1026 ( .A(n10728), .B(n10727), .Z(n682) );
  NAND U1027 ( .A(n681), .B(n682), .Z(n10735) );
  OR U1028 ( .A(n10868), .B(n10867), .Z(n683) );
  NAND U1029 ( .A(n10870), .B(n10869), .Z(n684) );
  NAND U1030 ( .A(n683), .B(n684), .Z(n10876) );
  OR U1031 ( .A(n10992), .B(n10991), .Z(n685) );
  NAND U1032 ( .A(n10994), .B(n10993), .Z(n686) );
  NAND U1033 ( .A(n685), .B(n686), .Z(n11000) );
  OR U1034 ( .A(n11170), .B(n11169), .Z(n687) );
  NAND U1035 ( .A(n11172), .B(n11171), .Z(n688) );
  NAND U1036 ( .A(n687), .B(n688), .Z(n11179) );
  OR U1037 ( .A(n11258), .B(n11257), .Z(n689) );
  NAND U1038 ( .A(n11260), .B(n11259), .Z(n690) );
  NAND U1039 ( .A(n689), .B(n690), .Z(n11266) );
  OR U1040 ( .A(n11418), .B(n11417), .Z(n691) );
  NAND U1041 ( .A(n11420), .B(n11419), .Z(n692) );
  NAND U1042 ( .A(n691), .B(n692), .Z(n11427) );
  OR U1043 ( .A(n11542), .B(n11541), .Z(n693) );
  NAND U1044 ( .A(n11544), .B(n11543), .Z(n694) );
  NAND U1045 ( .A(n693), .B(n694), .Z(n11550) );
  OR U1046 ( .A(n11693), .B(n11692), .Z(n695) );
  NAND U1047 ( .A(n11695), .B(n11694), .Z(n696) );
  NAND U1048 ( .A(n695), .B(n696), .Z(n11702) );
  OR U1049 ( .A(n11862), .B(n11861), .Z(n697) );
  NAND U1050 ( .A(n11864), .B(n11863), .Z(n698) );
  NAND U1051 ( .A(n697), .B(n698), .Z(n11870) );
  OR U1052 ( .A(n11977), .B(n11976), .Z(n699) );
  NAND U1053 ( .A(n11979), .B(n11978), .Z(n700) );
  NAND U1054 ( .A(n699), .B(n700), .Z(n11985) );
  OR U1055 ( .A(n12083), .B(n12082), .Z(n701) );
  NAND U1056 ( .A(n12085), .B(n12084), .Z(n702) );
  NAND U1057 ( .A(n701), .B(n702), .Z(n12092) );
  OR U1058 ( .A(n12171), .B(n12170), .Z(n703) );
  NAND U1059 ( .A(n12173), .B(n12172), .Z(n704) );
  NAND U1060 ( .A(n703), .B(n704), .Z(n12179) );
  OR U1061 ( .A(n12277), .B(n12276), .Z(n705) );
  NAND U1062 ( .A(n12279), .B(n12278), .Z(n706) );
  NAND U1063 ( .A(n705), .B(n706), .Z(n12285) );
  OR U1064 ( .A(n12368), .B(n12367), .Z(n707) );
  NAND U1065 ( .A(n12370), .B(n12369), .Z(n708) );
  NAND U1066 ( .A(n707), .B(n708), .Z(n12376) );
  OR U1067 ( .A(n4049), .B(n4050), .Z(n709) );
  NAND U1068 ( .A(n4055), .B(n4048), .Z(n710) );
  NAND U1069 ( .A(n709), .B(n710), .Z(n4057) );
  NAND U1070 ( .A(n4141), .B(sreg[1040]), .Z(n711) );
  XOR U1071 ( .A(sreg[1040]), .B(n4141), .Z(n712) );
  NANDN U1072 ( .A(n4140), .B(n712), .Z(n713) );
  NAND U1073 ( .A(n711), .B(n713), .Z(n4150) );
  OR U1074 ( .A(n4157), .B(n4156), .Z(n714) );
  NAND U1075 ( .A(n4159), .B(n4158), .Z(n715) );
  NAND U1076 ( .A(n714), .B(n715), .Z(n4166) );
  NAND U1077 ( .A(n4209), .B(sreg[1048]), .Z(n716) );
  XOR U1078 ( .A(sreg[1048]), .B(n4209), .Z(n717) );
  NANDN U1079 ( .A(n4208), .B(n717), .Z(n718) );
  NAND U1080 ( .A(n716), .B(n718), .Z(n4218) );
  OR U1081 ( .A(n4241), .B(n4240), .Z(n719) );
  NAND U1082 ( .A(n4243), .B(n4242), .Z(n720) );
  NAND U1083 ( .A(n719), .B(n720), .Z(n4249) );
  OR U1084 ( .A(n4347), .B(n4346), .Z(n721) );
  NAND U1085 ( .A(n4349), .B(n4348), .Z(n722) );
  NAND U1086 ( .A(n721), .B(n722), .Z(n4356) );
  OR U1087 ( .A(n4453), .B(n4452), .Z(n723) );
  NAND U1088 ( .A(n4455), .B(n4454), .Z(n724) );
  NAND U1089 ( .A(n723), .B(n724), .Z(n4461) );
  OR U1090 ( .A(n4586), .B(n4585), .Z(n725) );
  NAND U1091 ( .A(n4588), .B(n4587), .Z(n726) );
  NAND U1092 ( .A(n725), .B(n726), .Z(n4594) );
  OR U1093 ( .A(n4665), .B(n4664), .Z(n727) );
  NAND U1094 ( .A(n4667), .B(n4666), .Z(n728) );
  NAND U1095 ( .A(n727), .B(n728), .Z(n4673) );
  OR U1096 ( .A(n4780), .B(n4779), .Z(n729) );
  NAND U1097 ( .A(n4782), .B(n4781), .Z(n730) );
  NAND U1098 ( .A(n729), .B(n730), .Z(n4788) );
  OR U1099 ( .A(n4904), .B(n4903), .Z(n731) );
  NAND U1100 ( .A(n4906), .B(n4905), .Z(n732) );
  NAND U1101 ( .A(n731), .B(n732), .Z(n4913) );
  OR U1102 ( .A(n5064), .B(n5063), .Z(n733) );
  NAND U1103 ( .A(n5066), .B(n5065), .Z(n734) );
  NAND U1104 ( .A(n733), .B(n734), .Z(n5072) );
  OR U1105 ( .A(n5224), .B(n5223), .Z(n735) );
  NAND U1106 ( .A(n5226), .B(n5225), .Z(n736) );
  NAND U1107 ( .A(n735), .B(n736), .Z(n5233) );
  OR U1108 ( .A(n5330), .B(n5329), .Z(n737) );
  NAND U1109 ( .A(n5332), .B(n5331), .Z(n738) );
  NAND U1110 ( .A(n737), .B(n738), .Z(n5338) );
  OR U1111 ( .A(n5409), .B(n5408), .Z(n739) );
  NAND U1112 ( .A(n5411), .B(n5410), .Z(n740) );
  NAND U1113 ( .A(n739), .B(n740), .Z(n5417) );
  OR U1114 ( .A(n5560), .B(n5559), .Z(n741) );
  NAND U1115 ( .A(n5562), .B(n5561), .Z(n742) );
  NAND U1116 ( .A(n741), .B(n742), .Z(n5568) );
  OR U1117 ( .A(n5657), .B(n5656), .Z(n743) );
  NAND U1118 ( .A(n5659), .B(n5658), .Z(n744) );
  NAND U1119 ( .A(n743), .B(n744), .Z(n5665) );
  OR U1120 ( .A(n5790), .B(n5789), .Z(n745) );
  NAND U1121 ( .A(n5792), .B(n5791), .Z(n746) );
  NAND U1122 ( .A(n745), .B(n746), .Z(n5798) );
  OR U1123 ( .A(n5941), .B(n5940), .Z(n747) );
  NAND U1124 ( .A(n5943), .B(n5942), .Z(n748) );
  NAND U1125 ( .A(n747), .B(n748), .Z(n5949) );
  OR U1126 ( .A(n6038), .B(n6037), .Z(n749) );
  NAND U1127 ( .A(n6040), .B(n6039), .Z(n750) );
  NAND U1128 ( .A(n749), .B(n750), .Z(n6046) );
  OR U1129 ( .A(n6135), .B(n6134), .Z(n751) );
  NAND U1130 ( .A(n6137), .B(n6136), .Z(n752) );
  NAND U1131 ( .A(n751), .B(n752), .Z(n6143) );
  OR U1132 ( .A(n6232), .B(n6231), .Z(n753) );
  NAND U1133 ( .A(n6234), .B(n6233), .Z(n754) );
  NAND U1134 ( .A(n753), .B(n754), .Z(n6240) );
  OR U1135 ( .A(n6383), .B(n6382), .Z(n755) );
  NAND U1136 ( .A(n6385), .B(n6384), .Z(n756) );
  NAND U1137 ( .A(n755), .B(n756), .Z(n6391) );
  OR U1138 ( .A(n6516), .B(n6515), .Z(n757) );
  NAND U1139 ( .A(n6518), .B(n6517), .Z(n758) );
  NAND U1140 ( .A(n757), .B(n758), .Z(n6524) );
  OR U1141 ( .A(n6631), .B(n6630), .Z(n759) );
  NAND U1142 ( .A(n6633), .B(n6632), .Z(n760) );
  NAND U1143 ( .A(n759), .B(n760), .Z(n6639) );
  OR U1144 ( .A(n6737), .B(n6736), .Z(n761) );
  NAND U1145 ( .A(n6739), .B(n6738), .Z(n762) );
  NAND U1146 ( .A(n761), .B(n762), .Z(n6746) );
  OR U1147 ( .A(n6897), .B(n6896), .Z(n763) );
  NAND U1148 ( .A(n6899), .B(n6898), .Z(n764) );
  NAND U1149 ( .A(n763), .B(n764), .Z(n6905) );
  OR U1150 ( .A(n6994), .B(n6993), .Z(n765) );
  NAND U1151 ( .A(n6996), .B(n6995), .Z(n766) );
  NAND U1152 ( .A(n765), .B(n766), .Z(n7003) );
  OR U1153 ( .A(n7073), .B(n7072), .Z(n767) );
  NAND U1154 ( .A(n7075), .B(n7074), .Z(n768) );
  NAND U1155 ( .A(n767), .B(n768), .Z(n7081) );
  OR U1156 ( .A(n7170), .B(n7169), .Z(n769) );
  NAND U1157 ( .A(n7172), .B(n7171), .Z(n770) );
  NAND U1158 ( .A(n769), .B(n770), .Z(n7178) );
  OR U1159 ( .A(n7285), .B(n7284), .Z(n771) );
  NAND U1160 ( .A(n7287), .B(n7286), .Z(n772) );
  NAND U1161 ( .A(n771), .B(n772), .Z(n7293) );
  OR U1162 ( .A(n7418), .B(n7417), .Z(n773) );
  NAND U1163 ( .A(n7420), .B(n7419), .Z(n774) );
  NAND U1164 ( .A(n773), .B(n774), .Z(n7426) );
  OR U1165 ( .A(n7506), .B(n7505), .Z(n775) );
  NAND U1166 ( .A(n7508), .B(n7507), .Z(n776) );
  NAND U1167 ( .A(n775), .B(n776), .Z(n7514) );
  OR U1168 ( .A(n7630), .B(n7629), .Z(n777) );
  NAND U1169 ( .A(n7632), .B(n7631), .Z(n778) );
  NAND U1170 ( .A(n777), .B(n778), .Z(n7638) );
  OR U1171 ( .A(n7763), .B(n7762), .Z(n779) );
  NAND U1172 ( .A(n7765), .B(n7764), .Z(n780) );
  NAND U1173 ( .A(n779), .B(n780), .Z(n7772) );
  OR U1174 ( .A(n7842), .B(n7841), .Z(n781) );
  NAND U1175 ( .A(n7844), .B(n7843), .Z(n782) );
  NAND U1176 ( .A(n781), .B(n782), .Z(n7850) );
  OR U1177 ( .A(n7957), .B(n7956), .Z(n783) );
  NAND U1178 ( .A(n7959), .B(n7958), .Z(n784) );
  NAND U1179 ( .A(n783), .B(n784), .Z(n7965) );
  OR U1180 ( .A(n8045), .B(n8044), .Z(n785) );
  NAND U1181 ( .A(n8047), .B(n8046), .Z(n786) );
  NAND U1182 ( .A(n785), .B(n786), .Z(n8054) );
  OR U1183 ( .A(n8169), .B(n8168), .Z(n787) );
  NAND U1184 ( .A(n8171), .B(n8170), .Z(n788) );
  NAND U1185 ( .A(n787), .B(n788), .Z(n8177) );
  OR U1186 ( .A(n8266), .B(n8265), .Z(n789) );
  NAND U1187 ( .A(n8268), .B(n8267), .Z(n790) );
  NAND U1188 ( .A(n789), .B(n790), .Z(n8274) );
  OR U1189 ( .A(n8381), .B(n8380), .Z(n791) );
  NAND U1190 ( .A(n8383), .B(n8382), .Z(n792) );
  NAND U1191 ( .A(n791), .B(n792), .Z(n8389) );
  OR U1192 ( .A(n8478), .B(n8477), .Z(n793) );
  NAND U1193 ( .A(n8480), .B(n8479), .Z(n794) );
  NAND U1194 ( .A(n793), .B(n794), .Z(n8486) );
  OR U1195 ( .A(n8638), .B(n8637), .Z(n795) );
  NAND U1196 ( .A(n8640), .B(n8639), .Z(n796) );
  NAND U1197 ( .A(n795), .B(n796), .Z(n8647) );
  OR U1198 ( .A(n8744), .B(n8743), .Z(n797) );
  NAND U1199 ( .A(n8746), .B(n8745), .Z(n798) );
  NAND U1200 ( .A(n797), .B(n798), .Z(n8752) );
  OR U1201 ( .A(n8859), .B(n8858), .Z(n799) );
  NAND U1202 ( .A(n8861), .B(n8860), .Z(n800) );
  NAND U1203 ( .A(n799), .B(n800), .Z(n8867) );
  OR U1204 ( .A(n8992), .B(n8991), .Z(n801) );
  NAND U1205 ( .A(n8994), .B(n8993), .Z(n802) );
  NAND U1206 ( .A(n801), .B(n802), .Z(n9000) );
  OR U1207 ( .A(n9125), .B(n9124), .Z(n803) );
  NAND U1208 ( .A(n9127), .B(n9126), .Z(n804) );
  NAND U1209 ( .A(n803), .B(n804), .Z(n9133) );
  OR U1210 ( .A(n9213), .B(n9212), .Z(n805) );
  NAND U1211 ( .A(n9215), .B(n9214), .Z(n806) );
  NAND U1212 ( .A(n805), .B(n806), .Z(n9222) );
  OR U1213 ( .A(n9328), .B(n9327), .Z(n807) );
  NAND U1214 ( .A(n9330), .B(n9329), .Z(n808) );
  NAND U1215 ( .A(n807), .B(n808), .Z(n9337) );
  OR U1216 ( .A(n9416), .B(n9415), .Z(n809) );
  NAND U1217 ( .A(n9418), .B(n9417), .Z(n810) );
  NAND U1218 ( .A(n809), .B(n810), .Z(n9425) );
  OR U1219 ( .A(n9531), .B(n9530), .Z(n811) );
  NAND U1220 ( .A(n9533), .B(n9532), .Z(n812) );
  NAND U1221 ( .A(n811), .B(n812), .Z(n9540) );
  OR U1222 ( .A(n9646), .B(n9645), .Z(n813) );
  NAND U1223 ( .A(n9648), .B(n9647), .Z(n814) );
  NAND U1224 ( .A(n813), .B(n814), .Z(n9654) );
  OR U1225 ( .A(n9743), .B(n9742), .Z(n815) );
  NAND U1226 ( .A(n9745), .B(n9744), .Z(n816) );
  NAND U1227 ( .A(n815), .B(n816), .Z(n9751) );
  OR U1228 ( .A(n9840), .B(n9839), .Z(n817) );
  NAND U1229 ( .A(n9842), .B(n9841), .Z(n818) );
  NAND U1230 ( .A(n817), .B(n818), .Z(n9848) );
  OR U1231 ( .A(n9955), .B(n9954), .Z(n819) );
  NAND U1232 ( .A(n9957), .B(n9956), .Z(n820) );
  NAND U1233 ( .A(n819), .B(n820), .Z(n9963) );
  OR U1234 ( .A(n10088), .B(n10087), .Z(n821) );
  NAND U1235 ( .A(n10090), .B(n10089), .Z(n822) );
  NAND U1236 ( .A(n821), .B(n822), .Z(n10097) );
  OR U1237 ( .A(n10194), .B(n10193), .Z(n823) );
  NAND U1238 ( .A(n10196), .B(n10195), .Z(n824) );
  NAND U1239 ( .A(n823), .B(n824), .Z(n10203) );
  OR U1240 ( .A(n10300), .B(n10299), .Z(n825) );
  NAND U1241 ( .A(n10302), .B(n10301), .Z(n826) );
  NAND U1242 ( .A(n825), .B(n826), .Z(n10308) );
  OR U1243 ( .A(n10433), .B(n10432), .Z(n827) );
  NAND U1244 ( .A(n10435), .B(n10434), .Z(n828) );
  NAND U1245 ( .A(n827), .B(n828), .Z(n10441) );
  OR U1246 ( .A(n10530), .B(n10529), .Z(n829) );
  NAND U1247 ( .A(n10532), .B(n10531), .Z(n830) );
  NAND U1248 ( .A(n829), .B(n830), .Z(n10538) );
  OR U1249 ( .A(n10627), .B(n10626), .Z(n831) );
  NAND U1250 ( .A(n10629), .B(n10628), .Z(n832) );
  NAND U1251 ( .A(n831), .B(n832), .Z(n10635) );
  OR U1252 ( .A(n10733), .B(n10732), .Z(n833) );
  NAND U1253 ( .A(n10735), .B(n10734), .Z(n834) );
  NAND U1254 ( .A(n833), .B(n834), .Z(n10741) );
  OR U1255 ( .A(n10902), .B(n10901), .Z(n835) );
  NAND U1256 ( .A(n10904), .B(n10903), .Z(n836) );
  NAND U1257 ( .A(n835), .B(n836), .Z(n10910) );
  OR U1258 ( .A(n11062), .B(n11061), .Z(n837) );
  NAND U1259 ( .A(n11064), .B(n11063), .Z(n838) );
  NAND U1260 ( .A(n837), .B(n838), .Z(n11070) );
  OR U1261 ( .A(n11177), .B(n11176), .Z(n839) );
  NAND U1262 ( .A(n11179), .B(n11178), .Z(n840) );
  NAND U1263 ( .A(n839), .B(n840), .Z(n11185) );
  OR U1264 ( .A(n11274), .B(n11273), .Z(n841) );
  NAND U1265 ( .A(n11276), .B(n11275), .Z(n842) );
  NAND U1266 ( .A(n841), .B(n842), .Z(n11282) );
  OR U1267 ( .A(n11425), .B(n11424), .Z(n843) );
  NAND U1268 ( .A(n11427), .B(n11426), .Z(n844) );
  NAND U1269 ( .A(n843), .B(n844), .Z(n11433) );
  OR U1270 ( .A(n11576), .B(n11575), .Z(n845) );
  NAND U1271 ( .A(n11578), .B(n11577), .Z(n846) );
  NAND U1272 ( .A(n845), .B(n846), .Z(n11584) );
  OR U1273 ( .A(n11700), .B(n11699), .Z(n847) );
  NAND U1274 ( .A(n11702), .B(n11701), .Z(n848) );
  NAND U1275 ( .A(n847), .B(n848), .Z(n11708) );
  OR U1276 ( .A(n11878), .B(n11877), .Z(n849) );
  NAND U1277 ( .A(n11880), .B(n11879), .Z(n850) );
  NAND U1278 ( .A(n849), .B(n850), .Z(n11886) );
  OR U1279 ( .A(n11993), .B(n11992), .Z(n851) );
  NAND U1280 ( .A(n11995), .B(n11994), .Z(n852) );
  NAND U1281 ( .A(n851), .B(n852), .Z(n12001) );
  OR U1282 ( .A(n12090), .B(n12089), .Z(n853) );
  NAND U1283 ( .A(n12092), .B(n12091), .Z(n854) );
  NAND U1284 ( .A(n853), .B(n854), .Z(n12098) );
  OR U1285 ( .A(n12187), .B(n12186), .Z(n855) );
  NAND U1286 ( .A(n12189), .B(n12188), .Z(n856) );
  NAND U1287 ( .A(n855), .B(n856), .Z(n12195) );
  OR U1288 ( .A(n12302), .B(n12301), .Z(n857) );
  NAND U1289 ( .A(n12304), .B(n12303), .Z(n858) );
  NAND U1290 ( .A(n857), .B(n858), .Z(n12310) );
  OR U1291 ( .A(n12384), .B(n12383), .Z(n859) );
  NAND U1292 ( .A(n12386), .B(n12385), .Z(n860) );
  NAND U1293 ( .A(n859), .B(n860), .Z(n12392) );
  OR U1294 ( .A(n4121), .B(n4120), .Z(n861) );
  NAND U1295 ( .A(n4123), .B(n4122), .Z(n862) );
  NAND U1296 ( .A(n861), .B(n862), .Z(n4129) );
  NAND U1297 ( .A(n4014), .B(sreg[1025]), .Z(n863) );
  XOR U1298 ( .A(sreg[1025]), .B(n4014), .Z(n864) );
  NANDN U1299 ( .A(n4013), .B(n864), .Z(n865) );
  NAND U1300 ( .A(n863), .B(n865), .Z(n4022) );
  NAND U1301 ( .A(n4068), .B(sreg[1031]), .Z(n866) );
  XOR U1302 ( .A(sreg[1031]), .B(n4068), .Z(n867) );
  NAND U1303 ( .A(n867), .B(n4067), .Z(n868) );
  NAND U1304 ( .A(n866), .B(n868), .Z(n4076) );
  NAND U1305 ( .A(n4093), .B(sreg[1034]), .Z(n869) );
  XOR U1306 ( .A(sreg[1034]), .B(n4093), .Z(n870) );
  NANDN U1307 ( .A(n4092), .B(n870), .Z(n871) );
  NAND U1308 ( .A(n869), .B(n871), .Z(n4101) );
  XOR U1309 ( .A(n4117), .B(sreg[1037]), .Z(n872) );
  NANDN U1310 ( .A(n4118), .B(n872), .Z(n873) );
  NAND U1311 ( .A(n4117), .B(sreg[1037]), .Z(n874) );
  AND U1312 ( .A(n873), .B(n874), .Z(n4124) );
  NAND U1313 ( .A(n4161), .B(sreg[1042]), .Z(n875) );
  XOR U1314 ( .A(sreg[1042]), .B(n4161), .Z(n876) );
  NAND U1315 ( .A(n876), .B(n4160), .Z(n877) );
  NAND U1316 ( .A(n875), .B(n877), .Z(n4167) );
  NAND U1317 ( .A(n4183), .B(sreg[1045]), .Z(n878) );
  XOR U1318 ( .A(sreg[1045]), .B(n4183), .Z(n879) );
  NANDN U1319 ( .A(n4184), .B(n879), .Z(n880) );
  NAND U1320 ( .A(n878), .B(n880), .Z(n4192) );
  NAND U1321 ( .A(n4229), .B(sreg[1050]), .Z(n881) );
  XOR U1322 ( .A(sreg[1050]), .B(n4229), .Z(n882) );
  NAND U1323 ( .A(n882), .B(n4228), .Z(n883) );
  NAND U1324 ( .A(n881), .B(n883), .Z(n4237) );
  XOR U1325 ( .A(n4253), .B(sreg[1053]), .Z(n884) );
  NANDN U1326 ( .A(n4254), .B(n884), .Z(n885) );
  NAND U1327 ( .A(n4253), .B(sreg[1053]), .Z(n886) );
  AND U1328 ( .A(n885), .B(n886), .Z(n4263) );
  NAND U1329 ( .A(n4280), .B(sreg[1056]), .Z(n887) );
  XOR U1330 ( .A(sreg[1056]), .B(n4280), .Z(n888) );
  NANDN U1331 ( .A(n4279), .B(n888), .Z(n889) );
  NAND U1332 ( .A(n887), .B(n889), .Z(n4288) );
  XOR U1333 ( .A(n4304), .B(sreg[1059]), .Z(n890) );
  NANDN U1334 ( .A(n4305), .B(n890), .Z(n891) );
  NAND U1335 ( .A(n4304), .B(sreg[1059]), .Z(n892) );
  AND U1336 ( .A(n891), .B(n892), .Z(n4311) );
  NAND U1337 ( .A(n4328), .B(sreg[1062]), .Z(n893) );
  XOR U1338 ( .A(sreg[1062]), .B(n4328), .Z(n894) );
  NANDN U1339 ( .A(n4327), .B(n894), .Z(n895) );
  NAND U1340 ( .A(n893), .B(n895), .Z(n4336) );
  NAND U1341 ( .A(n4351), .B(sreg[1065]), .Z(n896) );
  XOR U1342 ( .A(sreg[1065]), .B(n4351), .Z(n897) );
  NAND U1343 ( .A(n897), .B(n4350), .Z(n898) );
  NAND U1344 ( .A(n896), .B(n898), .Z(n4360) );
  NAND U1345 ( .A(n4378), .B(sreg[1068]), .Z(n899) );
  XOR U1346 ( .A(sreg[1068]), .B(n4378), .Z(n900) );
  NANDN U1347 ( .A(n4379), .B(n900), .Z(n901) );
  NAND U1348 ( .A(n899), .B(n901), .Z(n4387) );
  XOR U1349 ( .A(n4403), .B(sreg[1071]), .Z(n902) );
  NANDN U1350 ( .A(n4404), .B(n902), .Z(n903) );
  NAND U1351 ( .A(n4403), .B(sreg[1071]), .Z(n904) );
  AND U1352 ( .A(n903), .B(n904), .Z(n4410) );
  NAND U1353 ( .A(n4427), .B(sreg[1074]), .Z(n905) );
  XOR U1354 ( .A(sreg[1074]), .B(n4427), .Z(n906) );
  NANDN U1355 ( .A(n4426), .B(n906), .Z(n907) );
  NAND U1356 ( .A(n905), .B(n907), .Z(n4433) );
  XOR U1357 ( .A(n4449), .B(sreg[1077]), .Z(n908) );
  NANDN U1358 ( .A(n4450), .B(n908), .Z(n909) );
  NAND U1359 ( .A(n4449), .B(sreg[1077]), .Z(n910) );
  AND U1360 ( .A(n909), .B(n910), .Z(n4456) );
  NAND U1361 ( .A(n4476), .B(sreg[1080]), .Z(n911) );
  XOR U1362 ( .A(sreg[1080]), .B(n4476), .Z(n912) );
  NANDN U1363 ( .A(n4475), .B(n912), .Z(n913) );
  NAND U1364 ( .A(n911), .B(n913), .Z(n4484) );
  NAND U1365 ( .A(n4500), .B(sreg[1083]), .Z(n914) );
  XOR U1366 ( .A(sreg[1083]), .B(n4500), .Z(n915) );
  NANDN U1367 ( .A(n4501), .B(n915), .Z(n916) );
  NAND U1368 ( .A(n914), .B(n916), .Z(n4509) );
  NAND U1369 ( .A(n4526), .B(sreg[1086]), .Z(n917) );
  XOR U1370 ( .A(sreg[1086]), .B(n4526), .Z(n918) );
  NANDN U1371 ( .A(n4525), .B(n918), .Z(n919) );
  NAND U1372 ( .A(n917), .B(n919), .Z(n4534) );
  XOR U1373 ( .A(n4552), .B(sreg[1089]), .Z(n920) );
  NANDN U1374 ( .A(n4553), .B(n920), .Z(n921) );
  NAND U1375 ( .A(n4552), .B(sreg[1089]), .Z(n922) );
  AND U1376 ( .A(n921), .B(n922), .Z(n4559) );
  NAND U1377 ( .A(n4576), .B(sreg[1092]), .Z(n923) );
  XOR U1378 ( .A(sreg[1092]), .B(n4576), .Z(n924) );
  NANDN U1379 ( .A(n4575), .B(n924), .Z(n925) );
  NAND U1380 ( .A(n923), .B(n925), .Z(n4582) );
  XOR U1381 ( .A(n4598), .B(sreg[1095]), .Z(n926) );
  NANDN U1382 ( .A(n4599), .B(n926), .Z(n927) );
  NAND U1383 ( .A(n4598), .B(sreg[1095]), .Z(n928) );
  AND U1384 ( .A(n927), .B(n928), .Z(n4608) );
  NAND U1385 ( .A(n4623), .B(sreg[1098]), .Z(n929) );
  XOR U1386 ( .A(sreg[1098]), .B(n4623), .Z(n930) );
  NAND U1387 ( .A(n930), .B(n4622), .Z(n931) );
  NAND U1388 ( .A(n929), .B(n931), .Z(n4629) );
  XOR U1389 ( .A(n4645), .B(sreg[1101]), .Z(n932) );
  NANDN U1390 ( .A(n4646), .B(n932), .Z(n933) );
  NAND U1391 ( .A(n4645), .B(sreg[1101]), .Z(n934) );
  AND U1392 ( .A(n933), .B(n934), .Z(n4652) );
  NAND U1393 ( .A(n4669), .B(sreg[1104]), .Z(n935) );
  XOR U1394 ( .A(sreg[1104]), .B(n4669), .Z(n936) );
  NANDN U1395 ( .A(n4668), .B(n936), .Z(n937) );
  NAND U1396 ( .A(n935), .B(n937), .Z(n4677) );
  XOR U1397 ( .A(n4696), .B(sreg[1107]), .Z(n938) );
  NANDN U1398 ( .A(n4697), .B(n938), .Z(n939) );
  NAND U1399 ( .A(n4696), .B(sreg[1107]), .Z(n940) );
  AND U1400 ( .A(n939), .B(n940), .Z(n4703) );
  NAND U1401 ( .A(n4720), .B(sreg[1110]), .Z(n941) );
  XOR U1402 ( .A(sreg[1110]), .B(n4720), .Z(n942) );
  NANDN U1403 ( .A(n4719), .B(n942), .Z(n943) );
  NAND U1404 ( .A(n941), .B(n943), .Z(n4728) );
  XOR U1405 ( .A(n4744), .B(sreg[1113]), .Z(n944) );
  NANDN U1406 ( .A(n4745), .B(n944), .Z(n945) );
  NAND U1407 ( .A(n4744), .B(sreg[1113]), .Z(n946) );
  AND U1408 ( .A(n945), .B(n946), .Z(n4751) );
  NAND U1409 ( .A(n4768), .B(sreg[1116]), .Z(n947) );
  XOR U1410 ( .A(sreg[1116]), .B(n4768), .Z(n948) );
  NANDN U1411 ( .A(n4767), .B(n948), .Z(n949) );
  NAND U1412 ( .A(n947), .B(n949), .Z(n4776) );
  XOR U1413 ( .A(n4792), .B(sreg[1119]), .Z(n950) );
  NANDN U1414 ( .A(n4793), .B(n950), .Z(n951) );
  NAND U1415 ( .A(n4792), .B(sreg[1119]), .Z(n952) );
  AND U1416 ( .A(n951), .B(n952), .Z(n4802) );
  NAND U1417 ( .A(n4820), .B(sreg[1122]), .Z(n953) );
  XOR U1418 ( .A(sreg[1122]), .B(n4820), .Z(n954) );
  NANDN U1419 ( .A(n4821), .B(n954), .Z(n955) );
  NAND U1420 ( .A(n953), .B(n955), .Z(n4829) );
  XOR U1421 ( .A(n4845), .B(sreg[1125]), .Z(n956) );
  NANDN U1422 ( .A(n4846), .B(n956), .Z(n957) );
  NAND U1423 ( .A(n4845), .B(sreg[1125]), .Z(n958) );
  AND U1424 ( .A(n957), .B(n958), .Z(n4852) );
  NAND U1425 ( .A(n4869), .B(sreg[1128]), .Z(n959) );
  XOR U1426 ( .A(sreg[1128]), .B(n4869), .Z(n960) );
  NANDN U1427 ( .A(n4868), .B(n960), .Z(n961) );
  NAND U1428 ( .A(n959), .B(n961), .Z(n4877) );
  NAND U1429 ( .A(n4894), .B(sreg[1131]), .Z(n962) );
  XOR U1430 ( .A(sreg[1131]), .B(n4894), .Z(n963) );
  NANDN U1431 ( .A(n4893), .B(n963), .Z(n964) );
  NAND U1432 ( .A(n962), .B(n964), .Z(n4900) );
  NAND U1433 ( .A(n4918), .B(sreg[1134]), .Z(n965) );
  XOR U1434 ( .A(sreg[1134]), .B(n4918), .Z(n966) );
  NAND U1435 ( .A(n966), .B(n4917), .Z(n967) );
  NAND U1436 ( .A(n965), .B(n967), .Z(n4926) );
  NAND U1437 ( .A(n4944), .B(sreg[1137]), .Z(n968) );
  XOR U1438 ( .A(sreg[1137]), .B(n4944), .Z(n969) );
  NANDN U1439 ( .A(n4945), .B(n969), .Z(n970) );
  NAND U1440 ( .A(n968), .B(n970), .Z(n4953) );
  NAND U1441 ( .A(n4970), .B(sreg[1140]), .Z(n971) );
  XOR U1442 ( .A(sreg[1140]), .B(n4970), .Z(n972) );
  NANDN U1443 ( .A(n4969), .B(n972), .Z(n973) );
  NAND U1444 ( .A(n971), .B(n973), .Z(n4978) );
  XOR U1445 ( .A(n4994), .B(sreg[1143]), .Z(n974) );
  NANDN U1446 ( .A(n4995), .B(n974), .Z(n975) );
  NAND U1447 ( .A(n4994), .B(sreg[1143]), .Z(n976) );
  AND U1448 ( .A(n975), .B(n976), .Z(n5001) );
  NAND U1449 ( .A(n5019), .B(sreg[1146]), .Z(n977) );
  XOR U1450 ( .A(sreg[1146]), .B(n5019), .Z(n978) );
  NANDN U1451 ( .A(n5020), .B(n978), .Z(n979) );
  NAND U1452 ( .A(n977), .B(n979), .Z(n5028) );
  XOR U1453 ( .A(n5044), .B(sreg[1149]), .Z(n980) );
  NANDN U1454 ( .A(n5045), .B(n980), .Z(n981) );
  NAND U1455 ( .A(n5044), .B(sreg[1149]), .Z(n982) );
  AND U1456 ( .A(n981), .B(n982), .Z(n5051) );
  NAND U1457 ( .A(n5068), .B(sreg[1152]), .Z(n983) );
  XOR U1458 ( .A(sreg[1152]), .B(n5068), .Z(n984) );
  NANDN U1459 ( .A(n5067), .B(n984), .Z(n985) );
  NAND U1460 ( .A(n983), .B(n985), .Z(n5076) );
  NAND U1461 ( .A(n5095), .B(sreg[1155]), .Z(n986) );
  XOR U1462 ( .A(sreg[1155]), .B(n5095), .Z(n987) );
  NANDN U1463 ( .A(n5096), .B(n987), .Z(n988) );
  NAND U1464 ( .A(n986), .B(n988), .Z(n5104) );
  NAND U1465 ( .A(n5122), .B(sreg[1158]), .Z(n989) );
  XOR U1466 ( .A(sreg[1158]), .B(n5122), .Z(n990) );
  NANDN U1467 ( .A(n5123), .B(n990), .Z(n991) );
  NAND U1468 ( .A(n989), .B(n991), .Z(n5131) );
  XOR U1469 ( .A(n5147), .B(sreg[1161]), .Z(n992) );
  NANDN U1470 ( .A(n5148), .B(n992), .Z(n993) );
  NAND U1471 ( .A(n5147), .B(sreg[1161]), .Z(n994) );
  AND U1472 ( .A(n993), .B(n994), .Z(n5154) );
  NAND U1473 ( .A(n5172), .B(sreg[1164]), .Z(n995) );
  XOR U1474 ( .A(sreg[1164]), .B(n5172), .Z(n996) );
  NANDN U1475 ( .A(n5173), .B(n996), .Z(n997) );
  NAND U1476 ( .A(n995), .B(n997), .Z(n5181) );
  XOR U1477 ( .A(n5197), .B(sreg[1167]), .Z(n998) );
  NANDN U1478 ( .A(n5198), .B(n998), .Z(n999) );
  NAND U1479 ( .A(n5197), .B(sreg[1167]), .Z(n1000) );
  AND U1480 ( .A(n999), .B(n1000), .Z(n5204) );
  NAND U1481 ( .A(n5221), .B(sreg[1170]), .Z(n1001) );
  XOR U1482 ( .A(sreg[1170]), .B(n5221), .Z(n1002) );
  NANDN U1483 ( .A(n5220), .B(n1002), .Z(n1003) );
  NAND U1484 ( .A(n1001), .B(n1003), .Z(n5227) );
  XOR U1485 ( .A(n5246), .B(sreg[1173]), .Z(n1004) );
  NANDN U1486 ( .A(n5247), .B(n1004), .Z(n1005) );
  NAND U1487 ( .A(n5246), .B(sreg[1173]), .Z(n1006) );
  AND U1488 ( .A(n1005), .B(n1006), .Z(n5253) );
  NAND U1489 ( .A(n5270), .B(sreg[1176]), .Z(n1007) );
  XOR U1490 ( .A(sreg[1176]), .B(n5270), .Z(n1008) );
  NANDN U1491 ( .A(n5269), .B(n1008), .Z(n1009) );
  NAND U1492 ( .A(n1007), .B(n1009), .Z(n5278) );
  XOR U1493 ( .A(n5294), .B(sreg[1179]), .Z(n1010) );
  NANDN U1494 ( .A(n5295), .B(n1010), .Z(n1011) );
  NAND U1495 ( .A(n5294), .B(sreg[1179]), .Z(n1012) );
  AND U1496 ( .A(n1011), .B(n1012), .Z(n5301) );
  NAND U1497 ( .A(n5318), .B(sreg[1182]), .Z(n1013) );
  XOR U1498 ( .A(sreg[1182]), .B(n5318), .Z(n1014) );
  NANDN U1499 ( .A(n5317), .B(n1014), .Z(n1015) );
  NAND U1500 ( .A(n1013), .B(n1015), .Z(n5326) );
  XOR U1501 ( .A(n5342), .B(sreg[1185]), .Z(n1016) );
  NANDN U1502 ( .A(n5343), .B(n1016), .Z(n1017) );
  NAND U1503 ( .A(n5342), .B(sreg[1185]), .Z(n1018) );
  AND U1504 ( .A(n1017), .B(n1018), .Z(n5352) );
  NAND U1505 ( .A(n5369), .B(sreg[1188]), .Z(n1019) );
  XOR U1506 ( .A(sreg[1188]), .B(n5369), .Z(n1020) );
  NANDN U1507 ( .A(n5368), .B(n1020), .Z(n1021) );
  NAND U1508 ( .A(n1019), .B(n1021), .Z(n5377) );
  NAND U1509 ( .A(n5392), .B(sreg[1191]), .Z(n1022) );
  XOR U1510 ( .A(sreg[1191]), .B(n5392), .Z(n1023) );
  NAND U1511 ( .A(n1023), .B(n5391), .Z(n1024) );
  NAND U1512 ( .A(n1022), .B(n1024), .Z(n5398) );
  NAND U1513 ( .A(n5413), .B(sreg[1194]), .Z(n1025) );
  XOR U1514 ( .A(sreg[1194]), .B(n5413), .Z(n1026) );
  NAND U1515 ( .A(n1026), .B(n5412), .Z(n1027) );
  NAND U1516 ( .A(n1025), .B(n1027), .Z(n5421) );
  NAND U1517 ( .A(n5440), .B(sreg[1197]), .Z(n1028) );
  XOR U1518 ( .A(sreg[1197]), .B(n5440), .Z(n1029) );
  NANDN U1519 ( .A(n5441), .B(n1029), .Z(n1030) );
  NAND U1520 ( .A(n1028), .B(n1030), .Z(n5449) );
  NAND U1521 ( .A(n5466), .B(sreg[1200]), .Z(n1031) );
  XOR U1522 ( .A(sreg[1200]), .B(n5466), .Z(n1032) );
  NANDN U1523 ( .A(n5465), .B(n1032), .Z(n1033) );
  NAND U1524 ( .A(n1031), .B(n1033), .Z(n5474) );
  XOR U1525 ( .A(n5490), .B(sreg[1203]), .Z(n1034) );
  NANDN U1526 ( .A(n5491), .B(n1034), .Z(n1035) );
  NAND U1527 ( .A(n5490), .B(sreg[1203]), .Z(n1036) );
  AND U1528 ( .A(n1035), .B(n1036), .Z(n5497) );
  NAND U1529 ( .A(n5514), .B(sreg[1206]), .Z(n1037) );
  XOR U1530 ( .A(sreg[1206]), .B(n5514), .Z(n1038) );
  NANDN U1531 ( .A(n5513), .B(n1038), .Z(n1039) );
  NAND U1532 ( .A(n1037), .B(n1039), .Z(n5522) );
  NAND U1533 ( .A(n5538), .B(sreg[1209]), .Z(n1040) );
  XOR U1534 ( .A(sreg[1209]), .B(n5538), .Z(n1041) );
  NANDN U1535 ( .A(n5539), .B(n1041), .Z(n1042) );
  NAND U1536 ( .A(n1040), .B(n1042), .Z(n5547) );
  NAND U1537 ( .A(n5564), .B(sreg[1212]), .Z(n1043) );
  XOR U1538 ( .A(sreg[1212]), .B(n5564), .Z(n1044) );
  NANDN U1539 ( .A(n5563), .B(n1044), .Z(n1045) );
  NAND U1540 ( .A(n1043), .B(n1045), .Z(n5572) );
  XOR U1541 ( .A(n5591), .B(sreg[1215]), .Z(n1046) );
  NANDN U1542 ( .A(n5592), .B(n1046), .Z(n1047) );
  NAND U1543 ( .A(n5591), .B(sreg[1215]), .Z(n1048) );
  AND U1544 ( .A(n1047), .B(n1048), .Z(n5598) );
  NAND U1545 ( .A(n5615), .B(sreg[1218]), .Z(n1049) );
  XOR U1546 ( .A(sreg[1218]), .B(n5615), .Z(n1050) );
  NANDN U1547 ( .A(n5614), .B(n1050), .Z(n1051) );
  NAND U1548 ( .A(n1049), .B(n1051), .Z(n5623) );
  XOR U1549 ( .A(n5639), .B(sreg[1221]), .Z(n1052) );
  NANDN U1550 ( .A(n5640), .B(n1052), .Z(n1053) );
  NAND U1551 ( .A(n5639), .B(sreg[1221]), .Z(n1054) );
  AND U1552 ( .A(n1053), .B(n1054), .Z(n5646) );
  NAND U1553 ( .A(n5661), .B(sreg[1224]), .Z(n1055) );
  XOR U1554 ( .A(sreg[1224]), .B(n5661), .Z(n1056) );
  NAND U1555 ( .A(n1056), .B(n5660), .Z(n1057) );
  NAND U1556 ( .A(n1055), .B(n1057), .Z(n5669) );
  XOR U1557 ( .A(n5688), .B(sreg[1227]), .Z(n1058) );
  NANDN U1558 ( .A(n5689), .B(n1058), .Z(n1059) );
  NAND U1559 ( .A(n5688), .B(sreg[1227]), .Z(n1060) );
  AND U1560 ( .A(n1059), .B(n1060), .Z(n5695) );
  NAND U1561 ( .A(n5712), .B(sreg[1230]), .Z(n1061) );
  XOR U1562 ( .A(sreg[1230]), .B(n5712), .Z(n1062) );
  NANDN U1563 ( .A(n5711), .B(n1062), .Z(n1063) );
  NAND U1564 ( .A(n1061), .B(n1063), .Z(n5720) );
  XOR U1565 ( .A(n5736), .B(sreg[1233]), .Z(n1064) );
  NANDN U1566 ( .A(n5737), .B(n1064), .Z(n1065) );
  NAND U1567 ( .A(n5736), .B(sreg[1233]), .Z(n1066) );
  AND U1568 ( .A(n1065), .B(n1066), .Z(n5743) );
  NAND U1569 ( .A(n5761), .B(sreg[1236]), .Z(n1067) );
  XOR U1570 ( .A(sreg[1236]), .B(n5761), .Z(n1068) );
  NANDN U1571 ( .A(n5762), .B(n1068), .Z(n1069) );
  NAND U1572 ( .A(n1067), .B(n1069), .Z(n5770) );
  XOR U1573 ( .A(n5786), .B(sreg[1239]), .Z(n1070) );
  NANDN U1574 ( .A(n5787), .B(n1070), .Z(n1071) );
  NAND U1575 ( .A(n5786), .B(sreg[1239]), .Z(n1072) );
  AND U1576 ( .A(n1071), .B(n1072), .Z(n5793) );
  NAND U1577 ( .A(n5811), .B(sreg[1242]), .Z(n1073) );
  XOR U1578 ( .A(sreg[1242]), .B(n5811), .Z(n1074) );
  NANDN U1579 ( .A(n5812), .B(n1074), .Z(n1075) );
  NAND U1580 ( .A(n1073), .B(n1075), .Z(n5820) );
  XOR U1581 ( .A(n5839), .B(sreg[1245]), .Z(n1076) );
  NANDN U1582 ( .A(n5840), .B(n1076), .Z(n1077) );
  NAND U1583 ( .A(n5839), .B(sreg[1245]), .Z(n1078) );
  AND U1584 ( .A(n1077), .B(n1078), .Z(n5846) );
  NAND U1585 ( .A(n5863), .B(sreg[1248]), .Z(n1079) );
  XOR U1586 ( .A(sreg[1248]), .B(n5863), .Z(n1080) );
  NANDN U1587 ( .A(n5862), .B(n1080), .Z(n1081) );
  NAND U1588 ( .A(n1079), .B(n1081), .Z(n5871) );
  XOR U1589 ( .A(n5887), .B(sreg[1251]), .Z(n1082) );
  NANDN U1590 ( .A(n5888), .B(n1082), .Z(n1083) );
  NAND U1591 ( .A(n5887), .B(sreg[1251]), .Z(n1084) );
  AND U1592 ( .A(n1083), .B(n1084), .Z(n5894) );
  NAND U1593 ( .A(n5911), .B(sreg[1254]), .Z(n1085) );
  XOR U1594 ( .A(sreg[1254]), .B(n5911), .Z(n1086) );
  NANDN U1595 ( .A(n5910), .B(n1086), .Z(n1087) );
  NAND U1596 ( .A(n1085), .B(n1087), .Z(n5919) );
  XOR U1597 ( .A(n5937), .B(sreg[1257]), .Z(n1088) );
  NANDN U1598 ( .A(n5938), .B(n1088), .Z(n1089) );
  NAND U1599 ( .A(n5937), .B(sreg[1257]), .Z(n1090) );
  AND U1600 ( .A(n1089), .B(n1090), .Z(n5944) );
  NAND U1601 ( .A(n5964), .B(sreg[1260]), .Z(n1091) );
  XOR U1602 ( .A(sreg[1260]), .B(n5964), .Z(n1092) );
  NANDN U1603 ( .A(n5963), .B(n1092), .Z(n1093) );
  NAND U1604 ( .A(n1091), .B(n1093), .Z(n5970) );
  XOR U1605 ( .A(n5986), .B(sreg[1263]), .Z(n1094) );
  NANDN U1606 ( .A(n5987), .B(n1094), .Z(n1095) );
  NAND U1607 ( .A(n5986), .B(sreg[1263]), .Z(n1096) );
  AND U1608 ( .A(n1095), .B(n1096), .Z(n5993) );
  NAND U1609 ( .A(n6010), .B(sreg[1266]), .Z(n1097) );
  XOR U1610 ( .A(sreg[1266]), .B(n6010), .Z(n1098) );
  NANDN U1611 ( .A(n6009), .B(n1098), .Z(n1099) );
  NAND U1612 ( .A(n1097), .B(n1099), .Z(n6018) );
  XOR U1613 ( .A(n6034), .B(sreg[1269]), .Z(n1100) );
  NANDN U1614 ( .A(n6035), .B(n1100), .Z(n1101) );
  NAND U1615 ( .A(n6034), .B(sreg[1269]), .Z(n1102) );
  AND U1616 ( .A(n1101), .B(n1102), .Z(n6041) );
  NAND U1617 ( .A(n6061), .B(sreg[1272]), .Z(n1103) );
  XOR U1618 ( .A(sreg[1272]), .B(n6061), .Z(n1104) );
  NANDN U1619 ( .A(n6060), .B(n1104), .Z(n1105) );
  NAND U1620 ( .A(n1103), .B(n1105), .Z(n6069) );
  XOR U1621 ( .A(n6085), .B(sreg[1275]), .Z(n1106) );
  NANDN U1622 ( .A(n6086), .B(n1106), .Z(n1107) );
  NAND U1623 ( .A(n6085), .B(sreg[1275]), .Z(n1108) );
  AND U1624 ( .A(n1107), .B(n1108), .Z(n6092) );
  NAND U1625 ( .A(n6109), .B(sreg[1278]), .Z(n1109) );
  XOR U1626 ( .A(sreg[1278]), .B(n6109), .Z(n1110) );
  NANDN U1627 ( .A(n6108), .B(n1110), .Z(n1111) );
  NAND U1628 ( .A(n1109), .B(n1111), .Z(n6117) );
  NAND U1629 ( .A(n6132), .B(sreg[1281]), .Z(n1112) );
  XOR U1630 ( .A(sreg[1281]), .B(n6132), .Z(n1113) );
  NAND U1631 ( .A(n1113), .B(n6131), .Z(n1114) );
  NAND U1632 ( .A(n1112), .B(n1114), .Z(n6138) );
  NAND U1633 ( .A(n6158), .B(sreg[1284]), .Z(n1115) );
  XOR U1634 ( .A(sreg[1284]), .B(n6158), .Z(n1116) );
  NANDN U1635 ( .A(n6157), .B(n1116), .Z(n1117) );
  NAND U1636 ( .A(n1115), .B(n1117), .Z(n6164) );
  NAND U1637 ( .A(n6180), .B(sreg[1287]), .Z(n1118) );
  XOR U1638 ( .A(sreg[1287]), .B(n6180), .Z(n1119) );
  NANDN U1639 ( .A(n6181), .B(n1119), .Z(n1120) );
  NAND U1640 ( .A(n1118), .B(n1120), .Z(n6189) );
  NAND U1641 ( .A(n6206), .B(sreg[1290]), .Z(n1121) );
  XOR U1642 ( .A(sreg[1290]), .B(n6206), .Z(n1122) );
  NANDN U1643 ( .A(n6205), .B(n1122), .Z(n1123) );
  NAND U1644 ( .A(n1121), .B(n1123), .Z(n6212) );
  XOR U1645 ( .A(n6228), .B(sreg[1293]), .Z(n1124) );
  NANDN U1646 ( .A(n6229), .B(n1124), .Z(n1125) );
  NAND U1647 ( .A(n6228), .B(sreg[1293]), .Z(n1126) );
  AND U1648 ( .A(n1125), .B(n1126), .Z(n6235) );
  NAND U1649 ( .A(n6255), .B(sreg[1296]), .Z(n1127) );
  XOR U1650 ( .A(sreg[1296]), .B(n6255), .Z(n1128) );
  NANDN U1651 ( .A(n6254), .B(n1128), .Z(n1129) );
  NAND U1652 ( .A(n1127), .B(n1129), .Z(n6263) );
  XOR U1653 ( .A(n6281), .B(sreg[1299]), .Z(n1130) );
  NANDN U1654 ( .A(n6282), .B(n1130), .Z(n1131) );
  NAND U1655 ( .A(n6281), .B(sreg[1299]), .Z(n1132) );
  AND U1656 ( .A(n1131), .B(n1132), .Z(n6288) );
  NAND U1657 ( .A(n6305), .B(sreg[1302]), .Z(n1133) );
  XOR U1658 ( .A(sreg[1302]), .B(n6305), .Z(n1134) );
  NANDN U1659 ( .A(n6304), .B(n1134), .Z(n1135) );
  NAND U1660 ( .A(n1133), .B(n1135), .Z(n6313) );
  XOR U1661 ( .A(n6329), .B(sreg[1305]), .Z(n1136) );
  NANDN U1662 ( .A(n6330), .B(n1136), .Z(n1137) );
  NAND U1663 ( .A(n6329), .B(sreg[1305]), .Z(n1138) );
  AND U1664 ( .A(n1137), .B(n1138), .Z(n6336) );
  NAND U1665 ( .A(n6354), .B(sreg[1308]), .Z(n1139) );
  XOR U1666 ( .A(sreg[1308]), .B(n6354), .Z(n1140) );
  NANDN U1667 ( .A(n6355), .B(n1140), .Z(n1141) );
  NAND U1668 ( .A(n1139), .B(n1141), .Z(n6363) );
  XOR U1669 ( .A(n6379), .B(sreg[1311]), .Z(n1142) );
  NANDN U1670 ( .A(n6380), .B(n1142), .Z(n1143) );
  NAND U1671 ( .A(n6379), .B(sreg[1311]), .Z(n1144) );
  AND U1672 ( .A(n1143), .B(n1144), .Z(n6386) );
  NAND U1673 ( .A(n6404), .B(sreg[1314]), .Z(n1145) );
  XOR U1674 ( .A(sreg[1314]), .B(n6404), .Z(n1146) );
  NANDN U1675 ( .A(n6405), .B(n1146), .Z(n1147) );
  NAND U1676 ( .A(n1145), .B(n1147), .Z(n6413) );
  XOR U1677 ( .A(n6432), .B(sreg[1317]), .Z(n1148) );
  NANDN U1678 ( .A(n6433), .B(n1148), .Z(n1149) );
  NAND U1679 ( .A(n6432), .B(sreg[1317]), .Z(n1150) );
  AND U1680 ( .A(n1149), .B(n1150), .Z(n6439) );
  NAND U1681 ( .A(n6456), .B(sreg[1320]), .Z(n1151) );
  XOR U1682 ( .A(sreg[1320]), .B(n6456), .Z(n1152) );
  NANDN U1683 ( .A(n6455), .B(n1152), .Z(n1153) );
  NAND U1684 ( .A(n1151), .B(n1153), .Z(n6464) );
  XOR U1685 ( .A(n6480), .B(sreg[1323]), .Z(n1154) );
  NANDN U1686 ( .A(n6481), .B(n1154), .Z(n1155) );
  NAND U1687 ( .A(n6480), .B(sreg[1323]), .Z(n1156) );
  AND U1688 ( .A(n1155), .B(n1156), .Z(n6487) );
  NAND U1689 ( .A(n6504), .B(sreg[1326]), .Z(n1157) );
  XOR U1690 ( .A(sreg[1326]), .B(n6504), .Z(n1158) );
  NANDN U1691 ( .A(n6503), .B(n1158), .Z(n1159) );
  NAND U1692 ( .A(n1157), .B(n1159), .Z(n6512) );
  XOR U1693 ( .A(n6528), .B(sreg[1329]), .Z(n1160) );
  NANDN U1694 ( .A(n6529), .B(n1160), .Z(n1161) );
  NAND U1695 ( .A(n6528), .B(sreg[1329]), .Z(n1162) );
  AND U1696 ( .A(n1161), .B(n1162), .Z(n6538) );
  NAND U1697 ( .A(n6555), .B(sreg[1332]), .Z(n1163) );
  XOR U1698 ( .A(sreg[1332]), .B(n6555), .Z(n1164) );
  NANDN U1699 ( .A(n6554), .B(n1164), .Z(n1165) );
  NAND U1700 ( .A(n1163), .B(n1165), .Z(n6563) );
  XOR U1701 ( .A(n6579), .B(sreg[1335]), .Z(n1166) );
  NANDN U1702 ( .A(n6580), .B(n1166), .Z(n1167) );
  NAND U1703 ( .A(n6579), .B(sreg[1335]), .Z(n1168) );
  AND U1704 ( .A(n1167), .B(n1168), .Z(n6586) );
  NAND U1705 ( .A(n6603), .B(sreg[1338]), .Z(n1169) );
  XOR U1706 ( .A(sreg[1338]), .B(n6603), .Z(n1170) );
  NANDN U1707 ( .A(n6602), .B(n1170), .Z(n1171) );
  NAND U1708 ( .A(n1169), .B(n1171), .Z(n6611) );
  XOR U1709 ( .A(n6627), .B(sreg[1341]), .Z(n1172) );
  NANDN U1710 ( .A(n6628), .B(n1172), .Z(n1173) );
  NAND U1711 ( .A(n6627), .B(sreg[1341]), .Z(n1174) );
  AND U1712 ( .A(n1173), .B(n1174), .Z(n6634) );
  NAND U1713 ( .A(n6654), .B(sreg[1344]), .Z(n1175) );
  XOR U1714 ( .A(sreg[1344]), .B(n6654), .Z(n1176) );
  NANDN U1715 ( .A(n6653), .B(n1176), .Z(n1177) );
  NAND U1716 ( .A(n1175), .B(n1177), .Z(n6662) );
  NAND U1717 ( .A(n6678), .B(sreg[1347]), .Z(n1178) );
  XOR U1718 ( .A(sreg[1347]), .B(n6678), .Z(n1179) );
  NANDN U1719 ( .A(n6679), .B(n1179), .Z(n1180) );
  NAND U1720 ( .A(n1178), .B(n1180), .Z(n6687) );
  NAND U1721 ( .A(n6704), .B(sreg[1350]), .Z(n1181) );
  XOR U1722 ( .A(sreg[1350]), .B(n6704), .Z(n1182) );
  NANDN U1723 ( .A(n6703), .B(n1182), .Z(n1183) );
  NAND U1724 ( .A(n1181), .B(n1183), .Z(n6710) );
  XOR U1725 ( .A(n6726), .B(sreg[1353]), .Z(n1184) );
  NANDN U1726 ( .A(n6727), .B(n1184), .Z(n1185) );
  NAND U1727 ( .A(n6726), .B(sreg[1353]), .Z(n1186) );
  AND U1728 ( .A(n1185), .B(n1186), .Z(n6733) );
  NAND U1729 ( .A(n6751), .B(sreg[1356]), .Z(n1187) );
  XOR U1730 ( .A(sreg[1356]), .B(n6751), .Z(n1188) );
  NAND U1731 ( .A(n1188), .B(n6750), .Z(n1189) );
  NAND U1732 ( .A(n1187), .B(n1189), .Z(n6759) );
  XOR U1733 ( .A(n6775), .B(sreg[1359]), .Z(n1190) );
  NANDN U1734 ( .A(n6776), .B(n1190), .Z(n1191) );
  NAND U1735 ( .A(n6775), .B(sreg[1359]), .Z(n1192) );
  AND U1736 ( .A(n1191), .B(n1192), .Z(n6782) );
  NAND U1737 ( .A(n6800), .B(sreg[1362]), .Z(n1193) );
  XOR U1738 ( .A(sreg[1362]), .B(n6800), .Z(n1194) );
  NANDN U1739 ( .A(n6801), .B(n1194), .Z(n1195) );
  NAND U1740 ( .A(n1193), .B(n1195), .Z(n6809) );
  NAND U1741 ( .A(n6825), .B(sreg[1365]), .Z(n1196) );
  XOR U1742 ( .A(sreg[1365]), .B(n6825), .Z(n1197) );
  NANDN U1743 ( .A(n6826), .B(n1197), .Z(n1198) );
  NAND U1744 ( .A(n1196), .B(n1198), .Z(n6834) );
  NAND U1745 ( .A(n6851), .B(sreg[1368]), .Z(n1199) );
  XOR U1746 ( .A(sreg[1368]), .B(n6851), .Z(n1200) );
  NANDN U1747 ( .A(n6850), .B(n1200), .Z(n1201) );
  NAND U1748 ( .A(n1199), .B(n1201), .Z(n6859) );
  NAND U1749 ( .A(n6875), .B(sreg[1371]), .Z(n1202) );
  XOR U1750 ( .A(sreg[1371]), .B(n6875), .Z(n1203) );
  NANDN U1751 ( .A(n6876), .B(n1203), .Z(n1204) );
  NAND U1752 ( .A(n1202), .B(n1204), .Z(n6884) );
  NAND U1753 ( .A(n6901), .B(sreg[1374]), .Z(n1205) );
  XOR U1754 ( .A(sreg[1374]), .B(n6901), .Z(n1206) );
  NANDN U1755 ( .A(n6900), .B(n1206), .Z(n1207) );
  NAND U1756 ( .A(n1205), .B(n1207), .Z(n6909) );
  XOR U1757 ( .A(n6928), .B(sreg[1377]), .Z(n1208) );
  NANDN U1758 ( .A(n6929), .B(n1208), .Z(n1209) );
  NAND U1759 ( .A(n6928), .B(sreg[1377]), .Z(n1210) );
  AND U1760 ( .A(n1209), .B(n1210), .Z(n6935) );
  NAND U1761 ( .A(n6952), .B(sreg[1380]), .Z(n1211) );
  XOR U1762 ( .A(sreg[1380]), .B(n6952), .Z(n1212) );
  NANDN U1763 ( .A(n6951), .B(n1212), .Z(n1213) );
  NAND U1764 ( .A(n1211), .B(n1213), .Z(n6960) );
  NAND U1765 ( .A(n6975), .B(sreg[1383]), .Z(n1214) );
  XOR U1766 ( .A(sreg[1383]), .B(n6975), .Z(n1215) );
  NAND U1767 ( .A(n1215), .B(n6974), .Z(n1216) );
  NAND U1768 ( .A(n1214), .B(n1216), .Z(n6981) );
  NAND U1769 ( .A(n6998), .B(sreg[1386]), .Z(n1217) );
  XOR U1770 ( .A(sreg[1386]), .B(n6998), .Z(n1218) );
  NANDN U1771 ( .A(n6997), .B(n1218), .Z(n1219) );
  NAND U1772 ( .A(n1217), .B(n1219), .Z(n7007) );
  XOR U1773 ( .A(n7023), .B(sreg[1389]), .Z(n1220) );
  NANDN U1774 ( .A(n7024), .B(n1220), .Z(n1221) );
  NAND U1775 ( .A(n7023), .B(sreg[1389]), .Z(n1222) );
  AND U1776 ( .A(n1221), .B(n1222), .Z(n7030) );
  NAND U1777 ( .A(n7047), .B(sreg[1392]), .Z(n1223) );
  XOR U1778 ( .A(sreg[1392]), .B(n7047), .Z(n1224) );
  NANDN U1779 ( .A(n7046), .B(n1224), .Z(n1225) );
  NAND U1780 ( .A(n1223), .B(n1225), .Z(n7055) );
  NAND U1781 ( .A(n7070), .B(sreg[1395]), .Z(n1226) );
  XOR U1782 ( .A(sreg[1395]), .B(n7070), .Z(n1227) );
  NAND U1783 ( .A(n1227), .B(n7069), .Z(n1228) );
  NAND U1784 ( .A(n1226), .B(n1228), .Z(n7076) );
  NAND U1785 ( .A(n7096), .B(sreg[1398]), .Z(n1229) );
  XOR U1786 ( .A(sreg[1398]), .B(n7096), .Z(n1230) );
  NANDN U1787 ( .A(n7095), .B(n1230), .Z(n1231) );
  NAND U1788 ( .A(n1229), .B(n1231), .Z(n7104) );
  NAND U1789 ( .A(n7119), .B(sreg[1401]), .Z(n1232) );
  XOR U1790 ( .A(sreg[1401]), .B(n7119), .Z(n1233) );
  NAND U1791 ( .A(n1233), .B(n7118), .Z(n1234) );
  NAND U1792 ( .A(n1232), .B(n1234), .Z(n7125) );
  NAND U1793 ( .A(n7142), .B(sreg[1404]), .Z(n1235) );
  XOR U1794 ( .A(sreg[1404]), .B(n7142), .Z(n1236) );
  NANDN U1795 ( .A(n7141), .B(n1236), .Z(n1237) );
  NAND U1796 ( .A(n1235), .B(n1237), .Z(n7150) );
  XOR U1797 ( .A(n7166), .B(sreg[1407]), .Z(n1238) );
  NANDN U1798 ( .A(n7167), .B(n1238), .Z(n1239) );
  NAND U1799 ( .A(n7166), .B(sreg[1407]), .Z(n1240) );
  AND U1800 ( .A(n1239), .B(n1240), .Z(n7173) );
  NAND U1801 ( .A(n7193), .B(sreg[1410]), .Z(n1241) );
  XOR U1802 ( .A(sreg[1410]), .B(n7193), .Z(n1242) );
  NANDN U1803 ( .A(n7192), .B(n1242), .Z(n1243) );
  NAND U1804 ( .A(n1241), .B(n1243), .Z(n7201) );
  XOR U1805 ( .A(n7217), .B(sreg[1413]), .Z(n1244) );
  NANDN U1806 ( .A(n7218), .B(n1244), .Z(n1245) );
  NAND U1807 ( .A(n7217), .B(sreg[1413]), .Z(n1246) );
  AND U1808 ( .A(n1245), .B(n1246), .Z(n7224) );
  NAND U1809 ( .A(n7241), .B(sreg[1416]), .Z(n1247) );
  XOR U1810 ( .A(sreg[1416]), .B(n7241), .Z(n1248) );
  NANDN U1811 ( .A(n7240), .B(n1248), .Z(n1249) );
  NAND U1812 ( .A(n1247), .B(n1249), .Z(n7249) );
  XOR U1813 ( .A(n7265), .B(sreg[1419]), .Z(n1250) );
  NANDN U1814 ( .A(n7266), .B(n1250), .Z(n1251) );
  NAND U1815 ( .A(n7265), .B(sreg[1419]), .Z(n1252) );
  AND U1816 ( .A(n1251), .B(n1252), .Z(n7272) );
  NAND U1817 ( .A(n7289), .B(sreg[1422]), .Z(n1253) );
  XOR U1818 ( .A(sreg[1422]), .B(n7289), .Z(n1254) );
  NANDN U1819 ( .A(n7288), .B(n1254), .Z(n1255) );
  NAND U1820 ( .A(n1253), .B(n1255), .Z(n7297) );
  XOR U1821 ( .A(n7316), .B(sreg[1425]), .Z(n1256) );
  NANDN U1822 ( .A(n7317), .B(n1256), .Z(n1257) );
  NAND U1823 ( .A(n7316), .B(sreg[1425]), .Z(n1258) );
  AND U1824 ( .A(n1257), .B(n1258), .Z(n7323) );
  NAND U1825 ( .A(n7341), .B(sreg[1428]), .Z(n1259) );
  XOR U1826 ( .A(sreg[1428]), .B(n7341), .Z(n1260) );
  NANDN U1827 ( .A(n7342), .B(n1260), .Z(n1261) );
  NAND U1828 ( .A(n1259), .B(n1261), .Z(n7350) );
  XOR U1829 ( .A(n7366), .B(sreg[1431]), .Z(n1262) );
  NANDN U1830 ( .A(n7367), .B(n1262), .Z(n1263) );
  NAND U1831 ( .A(n7366), .B(sreg[1431]), .Z(n1264) );
  AND U1832 ( .A(n1263), .B(n1264), .Z(n7373) );
  NAND U1833 ( .A(n7389), .B(sreg[1434]), .Z(n1265) );
  XOR U1834 ( .A(sreg[1434]), .B(n7389), .Z(n1266) );
  NANDN U1835 ( .A(n7390), .B(n1266), .Z(n1267) );
  NAND U1836 ( .A(n1265), .B(n1267), .Z(n7398) );
  XOR U1837 ( .A(n7414), .B(sreg[1437]), .Z(n1268) );
  NANDN U1838 ( .A(n7415), .B(n1268), .Z(n1269) );
  NAND U1839 ( .A(n7414), .B(sreg[1437]), .Z(n1270) );
  AND U1840 ( .A(n1269), .B(n1270), .Z(n7421) );
  NAND U1841 ( .A(n7441), .B(sreg[1440]), .Z(n1271) );
  XOR U1842 ( .A(sreg[1440]), .B(n7441), .Z(n1272) );
  NANDN U1843 ( .A(n7440), .B(n1272), .Z(n1273) );
  NAND U1844 ( .A(n1271), .B(n1273), .Z(n7449) );
  NAND U1845 ( .A(n7464), .B(sreg[1443]), .Z(n1274) );
  XOR U1846 ( .A(sreg[1443]), .B(n7464), .Z(n1275) );
  NAND U1847 ( .A(n1275), .B(n7463), .Z(n1276) );
  NAND U1848 ( .A(n1274), .B(n1276), .Z(n7472) );
  NAND U1849 ( .A(n7489), .B(sreg[1446]), .Z(n1277) );
  XOR U1850 ( .A(sreg[1446]), .B(n7489), .Z(n1278) );
  NANDN U1851 ( .A(n7488), .B(n1278), .Z(n1279) );
  NAND U1852 ( .A(n1277), .B(n1279), .Z(n7495) );
  NAND U1853 ( .A(n7510), .B(sreg[1449]), .Z(n1280) );
  XOR U1854 ( .A(sreg[1449]), .B(n7510), .Z(n1281) );
  NAND U1855 ( .A(n1281), .B(n7509), .Z(n1282) );
  NAND U1856 ( .A(n1280), .B(n1282), .Z(n7518) );
  NAND U1857 ( .A(n7538), .B(sreg[1452]), .Z(n1283) );
  XOR U1858 ( .A(sreg[1452]), .B(n7538), .Z(n1284) );
  NANDN U1859 ( .A(n7537), .B(n1284), .Z(n1285) );
  NAND U1860 ( .A(n1283), .B(n1285), .Z(n7546) );
  NAND U1861 ( .A(n7562), .B(sreg[1455]), .Z(n1286) );
  XOR U1862 ( .A(sreg[1455]), .B(n7562), .Z(n1287) );
  NANDN U1863 ( .A(n7563), .B(n1287), .Z(n1288) );
  NAND U1864 ( .A(n1286), .B(n1288), .Z(n7571) );
  NAND U1865 ( .A(n7588), .B(sreg[1458]), .Z(n1289) );
  XOR U1866 ( .A(sreg[1458]), .B(n7588), .Z(n1290) );
  NANDN U1867 ( .A(n7587), .B(n1290), .Z(n1291) );
  NAND U1868 ( .A(n1289), .B(n1291), .Z(n7594) );
  XOR U1869 ( .A(n7610), .B(sreg[1461]), .Z(n1292) );
  NANDN U1870 ( .A(n7611), .B(n1292), .Z(n1293) );
  NAND U1871 ( .A(n7610), .B(sreg[1461]), .Z(n1294) );
  AND U1872 ( .A(n1293), .B(n1294), .Z(n7617) );
  NAND U1873 ( .A(n7634), .B(sreg[1464]), .Z(n1295) );
  XOR U1874 ( .A(sreg[1464]), .B(n7634), .Z(n1296) );
  NANDN U1875 ( .A(n7633), .B(n1296), .Z(n1297) );
  NAND U1876 ( .A(n1295), .B(n1297), .Z(n7642) );
  XOR U1877 ( .A(n7661), .B(sreg[1467]), .Z(n1298) );
  NANDN U1878 ( .A(n7662), .B(n1298), .Z(n1299) );
  NAND U1879 ( .A(n7661), .B(sreg[1467]), .Z(n1300) );
  AND U1880 ( .A(n1299), .B(n1300), .Z(n7668) );
  NAND U1881 ( .A(n7685), .B(sreg[1470]), .Z(n1301) );
  XOR U1882 ( .A(sreg[1470]), .B(n7685), .Z(n1302) );
  NANDN U1883 ( .A(n7684), .B(n1302), .Z(n1303) );
  NAND U1884 ( .A(n1301), .B(n1303), .Z(n7693) );
  XOR U1885 ( .A(n7709), .B(sreg[1473]), .Z(n1304) );
  NANDN U1886 ( .A(n7710), .B(n1304), .Z(n1305) );
  NAND U1887 ( .A(n7709), .B(sreg[1473]), .Z(n1306) );
  AND U1888 ( .A(n1305), .B(n1306), .Z(n7716) );
  NAND U1889 ( .A(n7734), .B(sreg[1476]), .Z(n1307) );
  XOR U1890 ( .A(sreg[1476]), .B(n7734), .Z(n1308) );
  NANDN U1891 ( .A(n7735), .B(n1308), .Z(n1309) );
  NAND U1892 ( .A(n1307), .B(n1309), .Z(n7743) );
  XOR U1893 ( .A(n7759), .B(sreg[1479]), .Z(n1310) );
  NANDN U1894 ( .A(n7760), .B(n1310), .Z(n1311) );
  NAND U1895 ( .A(n7759), .B(sreg[1479]), .Z(n1312) );
  AND U1896 ( .A(n1311), .B(n1312), .Z(n7766) );
  XOR U1897 ( .A(n7785), .B(sreg[1482]), .Z(n1313) );
  NANDN U1898 ( .A(n7786), .B(n1313), .Z(n1314) );
  NAND U1899 ( .A(n7785), .B(sreg[1482]), .Z(n1315) );
  AND U1900 ( .A(n1314), .B(n1315), .Z(n7792) );
  NAND U1901 ( .A(n7807), .B(sreg[1485]), .Z(n1316) );
  XOR U1902 ( .A(sreg[1485]), .B(n7807), .Z(n1317) );
  NAND U1903 ( .A(n1317), .B(n7806), .Z(n1318) );
  NAND U1904 ( .A(n1316), .B(n1318), .Z(n7813) );
  NAND U1905 ( .A(n7830), .B(sreg[1488]), .Z(n1319) );
  XOR U1906 ( .A(sreg[1488]), .B(n7830), .Z(n1320) );
  NANDN U1907 ( .A(n7829), .B(n1320), .Z(n1321) );
  NAND U1908 ( .A(n1319), .B(n1321), .Z(n7838) );
  XOR U1909 ( .A(n7854), .B(sreg[1491]), .Z(n1322) );
  NANDN U1910 ( .A(n7855), .B(n1322), .Z(n1323) );
  NAND U1911 ( .A(n7854), .B(sreg[1491]), .Z(n1324) );
  AND U1912 ( .A(n1323), .B(n1324), .Z(n7864) );
  NAND U1913 ( .A(n7881), .B(sreg[1494]), .Z(n1325) );
  XOR U1914 ( .A(sreg[1494]), .B(n7881), .Z(n1326) );
  NANDN U1915 ( .A(n7880), .B(n1326), .Z(n1327) );
  NAND U1916 ( .A(n1325), .B(n1327), .Z(n7889) );
  XOR U1917 ( .A(n7905), .B(sreg[1497]), .Z(n1328) );
  NANDN U1918 ( .A(n7906), .B(n1328), .Z(n1329) );
  NAND U1919 ( .A(n7905), .B(sreg[1497]), .Z(n1330) );
  AND U1920 ( .A(n1329), .B(n1330), .Z(n7912) );
  NAND U1921 ( .A(n7929), .B(sreg[1500]), .Z(n1331) );
  XOR U1922 ( .A(sreg[1500]), .B(n7929), .Z(n1332) );
  NANDN U1923 ( .A(n7928), .B(n1332), .Z(n1333) );
  NAND U1924 ( .A(n1331), .B(n1333), .Z(n7937) );
  XOR U1925 ( .A(n7953), .B(sreg[1503]), .Z(n1334) );
  NANDN U1926 ( .A(n7954), .B(n1334), .Z(n1335) );
  NAND U1927 ( .A(n7953), .B(sreg[1503]), .Z(n1336) );
  AND U1928 ( .A(n1335), .B(n1336), .Z(n7960) );
  NAND U1929 ( .A(n7980), .B(sreg[1506]), .Z(n1337) );
  XOR U1930 ( .A(sreg[1506]), .B(n7980), .Z(n1338) );
  NANDN U1931 ( .A(n7979), .B(n1338), .Z(n1339) );
  NAND U1932 ( .A(n1337), .B(n1339), .Z(n7986) );
  XOR U1933 ( .A(n8002), .B(sreg[1509]), .Z(n1340) );
  NANDN U1934 ( .A(n8003), .B(n1340), .Z(n1341) );
  NAND U1935 ( .A(n8002), .B(sreg[1509]), .Z(n1342) );
  AND U1936 ( .A(n1341), .B(n1342), .Z(n8009) );
  XOR U1937 ( .A(n8025), .B(sreg[1512]), .Z(n1343) );
  NANDN U1938 ( .A(n8026), .B(n1343), .Z(n1344) );
  NAND U1939 ( .A(n8025), .B(sreg[1512]), .Z(n1345) );
  AND U1940 ( .A(n1344), .B(n1345), .Z(n8032) );
  NAND U1941 ( .A(n8049), .B(sreg[1515]), .Z(n1346) );
  XOR U1942 ( .A(sreg[1515]), .B(n8049), .Z(n1347) );
  NANDN U1943 ( .A(n8048), .B(n1347), .Z(n1348) );
  NAND U1944 ( .A(n1346), .B(n1348), .Z(n8058) );
  NAND U1945 ( .A(n8076), .B(sreg[1518]), .Z(n1349) );
  XOR U1946 ( .A(sreg[1518]), .B(n8076), .Z(n1350) );
  NANDN U1947 ( .A(n8077), .B(n1350), .Z(n1351) );
  NAND U1948 ( .A(n1349), .B(n1351), .Z(n8085) );
  XOR U1949 ( .A(n8101), .B(sreg[1521]), .Z(n1352) );
  NANDN U1950 ( .A(n8102), .B(n1352), .Z(n1353) );
  NAND U1951 ( .A(n8101), .B(sreg[1521]), .Z(n1354) );
  AND U1952 ( .A(n1353), .B(n1354), .Z(n8108) );
  NAND U1953 ( .A(n8125), .B(sreg[1524]), .Z(n1355) );
  XOR U1954 ( .A(sreg[1524]), .B(n8125), .Z(n1356) );
  NANDN U1955 ( .A(n8124), .B(n1356), .Z(n1357) );
  NAND U1956 ( .A(n1355), .B(n1357), .Z(n8133) );
  XOR U1957 ( .A(n8149), .B(sreg[1527]), .Z(n1358) );
  NANDN U1958 ( .A(n8150), .B(n1358), .Z(n1359) );
  NAND U1959 ( .A(n8149), .B(sreg[1527]), .Z(n1360) );
  AND U1960 ( .A(n1359), .B(n1360), .Z(n8156) );
  NAND U1961 ( .A(n8173), .B(sreg[1530]), .Z(n1361) );
  XOR U1962 ( .A(sreg[1530]), .B(n8173), .Z(n1362) );
  NANDN U1963 ( .A(n8172), .B(n1362), .Z(n1363) );
  NAND U1964 ( .A(n1361), .B(n1363), .Z(n8181) );
  XOR U1965 ( .A(n8200), .B(sreg[1533]), .Z(n1364) );
  NANDN U1966 ( .A(n8201), .B(n1364), .Z(n1365) );
  NAND U1967 ( .A(n8200), .B(sreg[1533]), .Z(n1366) );
  AND U1968 ( .A(n1365), .B(n1366), .Z(n8207) );
  NAND U1969 ( .A(n8224), .B(sreg[1536]), .Z(n1367) );
  XOR U1970 ( .A(sreg[1536]), .B(n8224), .Z(n1368) );
  NANDN U1971 ( .A(n8223), .B(n1368), .Z(n1369) );
  NAND U1972 ( .A(n1367), .B(n1369), .Z(n8232) );
  XOR U1973 ( .A(n8248), .B(sreg[1539]), .Z(n1370) );
  NANDN U1974 ( .A(n8249), .B(n1370), .Z(n1371) );
  NAND U1975 ( .A(n8248), .B(sreg[1539]), .Z(n1372) );
  AND U1976 ( .A(n1371), .B(n1372), .Z(n8255) );
  NAND U1977 ( .A(n8270), .B(sreg[1542]), .Z(n1373) );
  XOR U1978 ( .A(sreg[1542]), .B(n8270), .Z(n1374) );
  NAND U1979 ( .A(n1374), .B(n8269), .Z(n1375) );
  NAND U1980 ( .A(n1373), .B(n1375), .Z(n8278) );
  XOR U1981 ( .A(n8297), .B(sreg[1545]), .Z(n1376) );
  NANDN U1982 ( .A(n8298), .B(n1376), .Z(n1377) );
  NAND U1983 ( .A(n8297), .B(sreg[1545]), .Z(n1378) );
  AND U1984 ( .A(n1377), .B(n1378), .Z(n8304) );
  NAND U1985 ( .A(n8321), .B(sreg[1548]), .Z(n1379) );
  XOR U1986 ( .A(sreg[1548]), .B(n8321), .Z(n1380) );
  NANDN U1987 ( .A(n8320), .B(n1380), .Z(n1381) );
  NAND U1988 ( .A(n1379), .B(n1381), .Z(n8329) );
  XOR U1989 ( .A(n8345), .B(sreg[1551]), .Z(n1382) );
  NANDN U1990 ( .A(n8346), .B(n1382), .Z(n1383) );
  NAND U1991 ( .A(n8345), .B(sreg[1551]), .Z(n1384) );
  AND U1992 ( .A(n1383), .B(n1384), .Z(n8352) );
  NAND U1993 ( .A(n8369), .B(sreg[1554]), .Z(n1385) );
  XOR U1994 ( .A(sreg[1554]), .B(n8369), .Z(n1386) );
  NANDN U1995 ( .A(n8368), .B(n1386), .Z(n1387) );
  NAND U1996 ( .A(n1385), .B(n1387), .Z(n8377) );
  XOR U1997 ( .A(n8393), .B(sreg[1557]), .Z(n1388) );
  NANDN U1998 ( .A(n8394), .B(n1388), .Z(n1389) );
  NAND U1999 ( .A(n8393), .B(sreg[1557]), .Z(n1390) );
  AND U2000 ( .A(n1389), .B(n1390), .Z(n8403) );
  NAND U2001 ( .A(n8420), .B(sreg[1560]), .Z(n1391) );
  XOR U2002 ( .A(sreg[1560]), .B(n8420), .Z(n1392) );
  NANDN U2003 ( .A(n8419), .B(n1392), .Z(n1393) );
  NAND U2004 ( .A(n1391), .B(n1393), .Z(n8426) );
  XOR U2005 ( .A(n8442), .B(sreg[1563]), .Z(n1394) );
  NANDN U2006 ( .A(n8443), .B(n1394), .Z(n1395) );
  NAND U2007 ( .A(n8442), .B(sreg[1563]), .Z(n1396) );
  AND U2008 ( .A(n1395), .B(n1396), .Z(n8449) );
  NAND U2009 ( .A(n8466), .B(sreg[1566]), .Z(n1397) );
  XOR U2010 ( .A(sreg[1566]), .B(n8466), .Z(n1398) );
  NANDN U2011 ( .A(n8465), .B(n1398), .Z(n1399) );
  NAND U2012 ( .A(n1397), .B(n1399), .Z(n8474) );
  XOR U2013 ( .A(n8490), .B(sreg[1569]), .Z(n1400) );
  NANDN U2014 ( .A(n8491), .B(n1400), .Z(n1401) );
  NAND U2015 ( .A(n8490), .B(sreg[1569]), .Z(n1402) );
  AND U2016 ( .A(n1401), .B(n1402), .Z(n8500) );
  NAND U2017 ( .A(n8518), .B(sreg[1572]), .Z(n1403) );
  XOR U2018 ( .A(sreg[1572]), .B(n8518), .Z(n1404) );
  NANDN U2019 ( .A(n8519), .B(n1404), .Z(n1405) );
  NAND U2020 ( .A(n1403), .B(n1405), .Z(n8527) );
  XOR U2021 ( .A(n8545), .B(sreg[1575]), .Z(n1406) );
  NANDN U2022 ( .A(n8546), .B(n1406), .Z(n1407) );
  NAND U2023 ( .A(n8545), .B(sreg[1575]), .Z(n1408) );
  AND U2024 ( .A(n1407), .B(n1408), .Z(n8552) );
  NAND U2025 ( .A(n8570), .B(sreg[1578]), .Z(n1409) );
  XOR U2026 ( .A(sreg[1578]), .B(n8570), .Z(n1410) );
  NANDN U2027 ( .A(n8571), .B(n1410), .Z(n1411) );
  NAND U2028 ( .A(n1409), .B(n1411), .Z(n8579) );
  XOR U2029 ( .A(n8595), .B(sreg[1581]), .Z(n1412) );
  NANDN U2030 ( .A(n8596), .B(n1412), .Z(n1413) );
  NAND U2031 ( .A(n8595), .B(sreg[1581]), .Z(n1414) );
  AND U2032 ( .A(n1413), .B(n1414), .Z(n8602) );
  NAND U2033 ( .A(n8619), .B(sreg[1584]), .Z(n1415) );
  XOR U2034 ( .A(sreg[1584]), .B(n8619), .Z(n1416) );
  NANDN U2035 ( .A(n8618), .B(n1416), .Z(n1417) );
  NAND U2036 ( .A(n1415), .B(n1417), .Z(n8627) );
  NAND U2037 ( .A(n8642), .B(sreg[1587]), .Z(n1418) );
  XOR U2038 ( .A(sreg[1587]), .B(n8642), .Z(n1419) );
  NAND U2039 ( .A(n1419), .B(n8641), .Z(n1420) );
  NAND U2040 ( .A(n1418), .B(n1420), .Z(n8651) );
  NAND U2041 ( .A(n8668), .B(sreg[1590]), .Z(n1421) );
  XOR U2042 ( .A(sreg[1590]), .B(n8668), .Z(n1422) );
  NANDN U2043 ( .A(n8667), .B(n1422), .Z(n1423) );
  NAND U2044 ( .A(n1421), .B(n1423), .Z(n8676) );
  XOR U2045 ( .A(n8692), .B(sreg[1593]), .Z(n1424) );
  NANDN U2046 ( .A(n8693), .B(n1424), .Z(n1425) );
  NAND U2047 ( .A(n8692), .B(sreg[1593]), .Z(n1426) );
  AND U2048 ( .A(n1425), .B(n1426), .Z(n8699) );
  NAND U2049 ( .A(n8716), .B(sreg[1596]), .Z(n1427) );
  XOR U2050 ( .A(sreg[1596]), .B(n8716), .Z(n1428) );
  NANDN U2051 ( .A(n8715), .B(n1428), .Z(n1429) );
  NAND U2052 ( .A(n1427), .B(n1429), .Z(n8724) );
  XOR U2053 ( .A(n8740), .B(sreg[1599]), .Z(n1430) );
  NANDN U2054 ( .A(n8741), .B(n1430), .Z(n1431) );
  NAND U2055 ( .A(n8740), .B(sreg[1599]), .Z(n1432) );
  AND U2056 ( .A(n1431), .B(n1432), .Z(n8747) );
  NAND U2057 ( .A(n8767), .B(sreg[1602]), .Z(n1433) );
  XOR U2058 ( .A(sreg[1602]), .B(n8767), .Z(n1434) );
  NANDN U2059 ( .A(n8766), .B(n1434), .Z(n1435) );
  NAND U2060 ( .A(n1433), .B(n1435), .Z(n8775) );
  XOR U2061 ( .A(n8791), .B(sreg[1605]), .Z(n1436) );
  NANDN U2062 ( .A(n8792), .B(n1436), .Z(n1437) );
  NAND U2063 ( .A(n8791), .B(sreg[1605]), .Z(n1438) );
  AND U2064 ( .A(n1437), .B(n1438), .Z(n8798) );
  NAND U2065 ( .A(n8815), .B(sreg[1608]), .Z(n1439) );
  XOR U2066 ( .A(sreg[1608]), .B(n8815), .Z(n1440) );
  NANDN U2067 ( .A(n8814), .B(n1440), .Z(n1441) );
  NAND U2068 ( .A(n1439), .B(n1441), .Z(n8821) );
  XOR U2069 ( .A(n8839), .B(sreg[1611]), .Z(n1442) );
  NANDN U2070 ( .A(n8840), .B(n1442), .Z(n1443) );
  NAND U2071 ( .A(n8839), .B(sreg[1611]), .Z(n1444) );
  AND U2072 ( .A(n1443), .B(n1444), .Z(n8846) );
  NAND U2073 ( .A(n8863), .B(sreg[1614]), .Z(n1445) );
  XOR U2074 ( .A(sreg[1614]), .B(n8863), .Z(n1446) );
  NANDN U2075 ( .A(n8862), .B(n1446), .Z(n1447) );
  NAND U2076 ( .A(n1445), .B(n1447), .Z(n8871) );
  NAND U2077 ( .A(n8890), .B(sreg[1617]), .Z(n1448) );
  XOR U2078 ( .A(sreg[1617]), .B(n8890), .Z(n1449) );
  NANDN U2079 ( .A(n8891), .B(n1449), .Z(n1450) );
  NAND U2080 ( .A(n1448), .B(n1450), .Z(n8899) );
  NAND U2081 ( .A(n8916), .B(sreg[1620]), .Z(n1451) );
  XOR U2082 ( .A(sreg[1620]), .B(n8916), .Z(n1452) );
  NANDN U2083 ( .A(n8915), .B(n1452), .Z(n1453) );
  NAND U2084 ( .A(n1451), .B(n1453), .Z(n8924) );
  XOR U2085 ( .A(n8940), .B(sreg[1623]), .Z(n1454) );
  NANDN U2086 ( .A(n8941), .B(n1454), .Z(n1455) );
  NAND U2087 ( .A(n8940), .B(sreg[1623]), .Z(n1456) );
  AND U2088 ( .A(n1455), .B(n1456), .Z(n8947) );
  NAND U2089 ( .A(n8962), .B(sreg[1626]), .Z(n1457) );
  XOR U2090 ( .A(sreg[1626]), .B(n8962), .Z(n1458) );
  NAND U2091 ( .A(n1458), .B(n8961), .Z(n1459) );
  NAND U2092 ( .A(n1457), .B(n1459), .Z(n8970) );
  XOR U2093 ( .A(n8988), .B(sreg[1629]), .Z(n1460) );
  NANDN U2094 ( .A(n8989), .B(n1460), .Z(n1461) );
  NAND U2095 ( .A(n8988), .B(sreg[1629]), .Z(n1462) );
  AND U2096 ( .A(n1461), .B(n1462), .Z(n8995) );
  NAND U2097 ( .A(n9013), .B(sreg[1632]), .Z(n1463) );
  XOR U2098 ( .A(sreg[1632]), .B(n9013), .Z(n1464) );
  NANDN U2099 ( .A(n9014), .B(n1464), .Z(n1465) );
  NAND U2100 ( .A(n1463), .B(n1465), .Z(n9022) );
  XOR U2101 ( .A(n9041), .B(sreg[1635]), .Z(n1466) );
  NANDN U2102 ( .A(n9042), .B(n1466), .Z(n1467) );
  NAND U2103 ( .A(n9041), .B(sreg[1635]), .Z(n1468) );
  AND U2104 ( .A(n1467), .B(n1468), .Z(n9048) );
  NAND U2105 ( .A(n9066), .B(sreg[1638]), .Z(n1469) );
  XOR U2106 ( .A(sreg[1638]), .B(n9066), .Z(n1470) );
  NANDN U2107 ( .A(n9067), .B(n1470), .Z(n1471) );
  NAND U2108 ( .A(n1469), .B(n1471), .Z(n9075) );
  XOR U2109 ( .A(n9091), .B(sreg[1641]), .Z(n1472) );
  NANDN U2110 ( .A(n9092), .B(n1472), .Z(n1473) );
  NAND U2111 ( .A(n9091), .B(sreg[1641]), .Z(n1474) );
  AND U2112 ( .A(n1473), .B(n1474), .Z(n9098) );
  NAND U2113 ( .A(n9115), .B(sreg[1644]), .Z(n1475) );
  XOR U2114 ( .A(sreg[1644]), .B(n9115), .Z(n1476) );
  NANDN U2115 ( .A(n9114), .B(n1476), .Z(n1477) );
  NAND U2116 ( .A(n1475), .B(n1477), .Z(n9121) );
  XOR U2117 ( .A(n9137), .B(sreg[1647]), .Z(n1478) );
  NANDN U2118 ( .A(n9138), .B(n1478), .Z(n1479) );
  NAND U2119 ( .A(n9137), .B(sreg[1647]), .Z(n1480) );
  AND U2120 ( .A(n1479), .B(n1480), .Z(n9147) );
  NAND U2121 ( .A(n9164), .B(sreg[1650]), .Z(n1481) );
  XOR U2122 ( .A(sreg[1650]), .B(n9164), .Z(n1482) );
  NANDN U2123 ( .A(n9163), .B(n1482), .Z(n1483) );
  NAND U2124 ( .A(n1481), .B(n1483), .Z(n9172) );
  NAND U2125 ( .A(n9187), .B(sreg[1653]), .Z(n1484) );
  XOR U2126 ( .A(sreg[1653]), .B(n9187), .Z(n1485) );
  NAND U2127 ( .A(n1485), .B(n9186), .Z(n1486) );
  NAND U2128 ( .A(n1484), .B(n1486), .Z(n9193) );
  NAND U2129 ( .A(n9210), .B(sreg[1656]), .Z(n1487) );
  XOR U2130 ( .A(sreg[1656]), .B(n9210), .Z(n1488) );
  NANDN U2131 ( .A(n9209), .B(n1488), .Z(n1489) );
  NAND U2132 ( .A(n1487), .B(n1489), .Z(n9216) );
  XOR U2133 ( .A(n9235), .B(sreg[1659]), .Z(n1490) );
  NANDN U2134 ( .A(n9236), .B(n1490), .Z(n1491) );
  NAND U2135 ( .A(n9235), .B(sreg[1659]), .Z(n1492) );
  AND U2136 ( .A(n1491), .B(n1492), .Z(n9242) );
  NAND U2137 ( .A(n9259), .B(sreg[1662]), .Z(n1493) );
  XOR U2138 ( .A(sreg[1662]), .B(n9259), .Z(n1494) );
  NANDN U2139 ( .A(n9258), .B(n1494), .Z(n1495) );
  NAND U2140 ( .A(n1493), .B(n1495), .Z(n9267) );
  XOR U2141 ( .A(n9285), .B(sreg[1665]), .Z(n1496) );
  NANDN U2142 ( .A(n9286), .B(n1496), .Z(n1497) );
  NAND U2143 ( .A(n9285), .B(sreg[1665]), .Z(n1498) );
  AND U2144 ( .A(n1497), .B(n1498), .Z(n9292) );
  NAND U2145 ( .A(n9309), .B(sreg[1668]), .Z(n1499) );
  XOR U2146 ( .A(sreg[1668]), .B(n9309), .Z(n1500) );
  NANDN U2147 ( .A(n9308), .B(n1500), .Z(n1501) );
  NAND U2148 ( .A(n1499), .B(n1501), .Z(n9317) );
  NAND U2149 ( .A(n9332), .B(sreg[1671]), .Z(n1502) );
  XOR U2150 ( .A(sreg[1671]), .B(n9332), .Z(n1503) );
  NAND U2151 ( .A(n1503), .B(n9331), .Z(n1504) );
  NAND U2152 ( .A(n1502), .B(n1504), .Z(n9341) );
  NAND U2153 ( .A(n9358), .B(sreg[1674]), .Z(n1505) );
  XOR U2154 ( .A(sreg[1674]), .B(n9358), .Z(n1506) );
  NANDN U2155 ( .A(n9357), .B(n1506), .Z(n1507) );
  NAND U2156 ( .A(n1505), .B(n1507), .Z(n9366) );
  XOR U2157 ( .A(n9382), .B(sreg[1677]), .Z(n1508) );
  NANDN U2158 ( .A(n9383), .B(n1508), .Z(n1509) );
  NAND U2159 ( .A(n9382), .B(sreg[1677]), .Z(n1510) );
  AND U2160 ( .A(n1509), .B(n1510), .Z(n9389) );
  NAND U2161 ( .A(n9406), .B(sreg[1680]), .Z(n1511) );
  XOR U2162 ( .A(sreg[1680]), .B(n9406), .Z(n1512) );
  NANDN U2163 ( .A(n9405), .B(n1512), .Z(n1513) );
  NAND U2164 ( .A(n1511), .B(n1513), .Z(n9412) );
  NAND U2165 ( .A(n9430), .B(sreg[1683]), .Z(n1514) );
  XOR U2166 ( .A(sreg[1683]), .B(n9430), .Z(n1515) );
  NAND U2167 ( .A(n1515), .B(n9429), .Z(n1516) );
  NAND U2168 ( .A(n1514), .B(n1516), .Z(n9436) );
  NAND U2169 ( .A(n9453), .B(sreg[1686]), .Z(n1517) );
  XOR U2170 ( .A(sreg[1686]), .B(n9453), .Z(n1518) );
  NANDN U2171 ( .A(n9452), .B(n1518), .Z(n1519) );
  NAND U2172 ( .A(n1517), .B(n1519), .Z(n9461) );
  XOR U2173 ( .A(n9477), .B(sreg[1689]), .Z(n1520) );
  NANDN U2174 ( .A(n9478), .B(n1520), .Z(n1521) );
  NAND U2175 ( .A(n9477), .B(sreg[1689]), .Z(n1522) );
  AND U2176 ( .A(n1521), .B(n1522), .Z(n9484) );
  NAND U2177 ( .A(n9502), .B(sreg[1692]), .Z(n1523) );
  XOR U2178 ( .A(sreg[1692]), .B(n9502), .Z(n1524) );
  NANDN U2179 ( .A(n9503), .B(n1524), .Z(n1525) );
  NAND U2180 ( .A(n1523), .B(n1525), .Z(n9511) );
  XOR U2181 ( .A(n9527), .B(sreg[1695]), .Z(n1526) );
  NANDN U2182 ( .A(n9528), .B(n1526), .Z(n1527) );
  NAND U2183 ( .A(n9527), .B(sreg[1695]), .Z(n1528) );
  AND U2184 ( .A(n1527), .B(n1528), .Z(n9534) );
  NAND U2185 ( .A(n9552), .B(sreg[1698]), .Z(n1529) );
  XOR U2186 ( .A(sreg[1698]), .B(n9552), .Z(n1530) );
  NAND U2187 ( .A(n1530), .B(n9551), .Z(n1531) );
  NAND U2188 ( .A(n1529), .B(n1531), .Z(n9560) );
  XOR U2189 ( .A(n9576), .B(sreg[1701]), .Z(n1532) );
  NANDN U2190 ( .A(n9577), .B(n1532), .Z(n1533) );
  NAND U2191 ( .A(n9576), .B(sreg[1701]), .Z(n1534) );
  AND U2192 ( .A(n1533), .B(n1534), .Z(n9583) );
  NAND U2193 ( .A(n9600), .B(sreg[1704]), .Z(n1535) );
  XOR U2194 ( .A(sreg[1704]), .B(n9600), .Z(n1536) );
  NANDN U2195 ( .A(n9599), .B(n1536), .Z(n1537) );
  NAND U2196 ( .A(n1535), .B(n1537), .Z(n9608) );
  XOR U2197 ( .A(n9626), .B(sreg[1707]), .Z(n1538) );
  NANDN U2198 ( .A(n9627), .B(n1538), .Z(n1539) );
  NAND U2199 ( .A(n9626), .B(sreg[1707]), .Z(n1540) );
  AND U2200 ( .A(n1539), .B(n1540), .Z(n9633) );
  NAND U2201 ( .A(n9650), .B(sreg[1710]), .Z(n1541) );
  XOR U2202 ( .A(sreg[1710]), .B(n9650), .Z(n1542) );
  NANDN U2203 ( .A(n9649), .B(n1542), .Z(n1543) );
  NAND U2204 ( .A(n1541), .B(n1543), .Z(n9658) );
  XOR U2205 ( .A(n9677), .B(sreg[1713]), .Z(n1544) );
  NANDN U2206 ( .A(n9678), .B(n1544), .Z(n1545) );
  NAND U2207 ( .A(n9677), .B(sreg[1713]), .Z(n1546) );
  AND U2208 ( .A(n1545), .B(n1546), .Z(n9684) );
  NAND U2209 ( .A(n9701), .B(sreg[1716]), .Z(n1547) );
  XOR U2210 ( .A(sreg[1716]), .B(n9701), .Z(n1548) );
  NANDN U2211 ( .A(n9700), .B(n1548), .Z(n1549) );
  NAND U2212 ( .A(n1547), .B(n1549), .Z(n9709) );
  XOR U2213 ( .A(n9725), .B(sreg[1719]), .Z(n1550) );
  NANDN U2214 ( .A(n9726), .B(n1550), .Z(n1551) );
  NAND U2215 ( .A(n9725), .B(sreg[1719]), .Z(n1552) );
  AND U2216 ( .A(n1551), .B(n1552), .Z(n9732) );
  NAND U2217 ( .A(n9747), .B(sreg[1722]), .Z(n1553) );
  XOR U2218 ( .A(sreg[1722]), .B(n9747), .Z(n1554) );
  NAND U2219 ( .A(n1554), .B(n9746), .Z(n1555) );
  NAND U2220 ( .A(n1553), .B(n1555), .Z(n9755) );
  XOR U2221 ( .A(n9774), .B(sreg[1725]), .Z(n1556) );
  NANDN U2222 ( .A(n9775), .B(n1556), .Z(n1557) );
  NAND U2223 ( .A(n9774), .B(sreg[1725]), .Z(n1558) );
  AND U2224 ( .A(n1557), .B(n1558), .Z(n9781) );
  NAND U2225 ( .A(n9798), .B(sreg[1728]), .Z(n1559) );
  XOR U2226 ( .A(sreg[1728]), .B(n9798), .Z(n1560) );
  NANDN U2227 ( .A(n9797), .B(n1560), .Z(n1561) );
  NAND U2228 ( .A(n1559), .B(n1561), .Z(n9806) );
  NAND U2229 ( .A(n9821), .B(sreg[1731]), .Z(n1562) );
  XOR U2230 ( .A(sreg[1731]), .B(n9821), .Z(n1563) );
  NAND U2231 ( .A(n1563), .B(n9820), .Z(n1564) );
  NAND U2232 ( .A(n1562), .B(n1564), .Z(n9827) );
  NAND U2233 ( .A(n9844), .B(sreg[1734]), .Z(n1565) );
  XOR U2234 ( .A(sreg[1734]), .B(n9844), .Z(n1566) );
  NANDN U2235 ( .A(n9843), .B(n1566), .Z(n1567) );
  NAND U2236 ( .A(n1565), .B(n1567), .Z(n9852) );
  XOR U2237 ( .A(n9871), .B(sreg[1737]), .Z(n1568) );
  NANDN U2238 ( .A(n9872), .B(n1568), .Z(n1569) );
  NAND U2239 ( .A(n9871), .B(sreg[1737]), .Z(n1570) );
  AND U2240 ( .A(n1569), .B(n1570), .Z(n9878) );
  NAND U2241 ( .A(n9895), .B(sreg[1740]), .Z(n1571) );
  XOR U2242 ( .A(sreg[1740]), .B(n9895), .Z(n1572) );
  NANDN U2243 ( .A(n9894), .B(n1572), .Z(n1573) );
  NAND U2244 ( .A(n1571), .B(n1573), .Z(n9903) );
  XOR U2245 ( .A(n9919), .B(sreg[1743]), .Z(n1574) );
  NANDN U2246 ( .A(n9920), .B(n1574), .Z(n1575) );
  NAND U2247 ( .A(n9919), .B(sreg[1743]), .Z(n1576) );
  AND U2248 ( .A(n1575), .B(n1576), .Z(n9926) );
  NAND U2249 ( .A(n9943), .B(sreg[1746]), .Z(n1577) );
  XOR U2250 ( .A(sreg[1746]), .B(n9943), .Z(n1578) );
  NANDN U2251 ( .A(n9942), .B(n1578), .Z(n1579) );
  NAND U2252 ( .A(n1577), .B(n1579), .Z(n9951) );
  XOR U2253 ( .A(n9967), .B(sreg[1749]), .Z(n1580) );
  NANDN U2254 ( .A(n9968), .B(n1580), .Z(n1581) );
  NAND U2255 ( .A(n9967), .B(sreg[1749]), .Z(n1582) );
  AND U2256 ( .A(n1581), .B(n1582), .Z(n9977) );
  NAND U2257 ( .A(n9994), .B(sreg[1752]), .Z(n1583) );
  XOR U2258 ( .A(sreg[1752]), .B(n9994), .Z(n1584) );
  NANDN U2259 ( .A(n9993), .B(n1584), .Z(n1585) );
  NAND U2260 ( .A(n1583), .B(n1585), .Z(n10002) );
  XOR U2261 ( .A(n10018), .B(sreg[1755]), .Z(n1586) );
  NANDN U2262 ( .A(n10019), .B(n1586), .Z(n1587) );
  NAND U2263 ( .A(n10018), .B(sreg[1755]), .Z(n1588) );
  AND U2264 ( .A(n1587), .B(n1588), .Z(n10025) );
  NAND U2265 ( .A(n10043), .B(sreg[1758]), .Z(n1589) );
  XOR U2266 ( .A(sreg[1758]), .B(n10043), .Z(n1590) );
  NANDN U2267 ( .A(n10044), .B(n1590), .Z(n1591) );
  NAND U2268 ( .A(n1589), .B(n1591), .Z(n10052) );
  XOR U2269 ( .A(n10068), .B(sreg[1761]), .Z(n1592) );
  NANDN U2270 ( .A(n10069), .B(n1592), .Z(n1593) );
  NAND U2271 ( .A(n10068), .B(sreg[1761]), .Z(n1594) );
  AND U2272 ( .A(n1593), .B(n1594), .Z(n10075) );
  NAND U2273 ( .A(n10092), .B(sreg[1764]), .Z(n1595) );
  XOR U2274 ( .A(sreg[1764]), .B(n10092), .Z(n1596) );
  NANDN U2275 ( .A(n10091), .B(n1596), .Z(n1597) );
  NAND U2276 ( .A(n1595), .B(n1597), .Z(n10101) );
  XOR U2277 ( .A(n10119), .B(sreg[1767]), .Z(n1598) );
  NANDN U2278 ( .A(n10120), .B(n1598), .Z(n1599) );
  NAND U2279 ( .A(n10119), .B(sreg[1767]), .Z(n1600) );
  AND U2280 ( .A(n1599), .B(n1600), .Z(n10126) );
  NAND U2281 ( .A(n10143), .B(sreg[1770]), .Z(n1601) );
  XOR U2282 ( .A(sreg[1770]), .B(n10143), .Z(n1602) );
  NANDN U2283 ( .A(n10142), .B(n1602), .Z(n1603) );
  NAND U2284 ( .A(n1601), .B(n1603), .Z(n10151) );
  XOR U2285 ( .A(n10167), .B(sreg[1773]), .Z(n1604) );
  NANDN U2286 ( .A(n10168), .B(n1604), .Z(n1605) );
  NAND U2287 ( .A(n10167), .B(sreg[1773]), .Z(n1606) );
  AND U2288 ( .A(n1605), .B(n1606), .Z(n10174) );
  NAND U2289 ( .A(n10191), .B(sreg[1776]), .Z(n1607) );
  XOR U2290 ( .A(sreg[1776]), .B(n10191), .Z(n1608) );
  NANDN U2291 ( .A(n10190), .B(n1608), .Z(n1609) );
  NAND U2292 ( .A(n1607), .B(n1609), .Z(n10197) );
  XOR U2293 ( .A(n10216), .B(sreg[1779]), .Z(n1610) );
  NANDN U2294 ( .A(n10217), .B(n1610), .Z(n1611) );
  NAND U2295 ( .A(n10216), .B(sreg[1779]), .Z(n1612) );
  AND U2296 ( .A(n1611), .B(n1612), .Z(n10223) );
  NAND U2297 ( .A(n10240), .B(sreg[1782]), .Z(n1613) );
  XOR U2298 ( .A(sreg[1782]), .B(n10240), .Z(n1614) );
  NANDN U2299 ( .A(n10239), .B(n1614), .Z(n1615) );
  NAND U2300 ( .A(n1613), .B(n1615), .Z(n10248) );
  XOR U2301 ( .A(n10264), .B(sreg[1785]), .Z(n1616) );
  NANDN U2302 ( .A(n10265), .B(n1616), .Z(n1617) );
  NAND U2303 ( .A(n10264), .B(sreg[1785]), .Z(n1618) );
  AND U2304 ( .A(n1617), .B(n1618), .Z(n10271) );
  NAND U2305 ( .A(n10288), .B(sreg[1788]), .Z(n1619) );
  XOR U2306 ( .A(sreg[1788]), .B(n10288), .Z(n1620) );
  NANDN U2307 ( .A(n10287), .B(n1620), .Z(n1621) );
  NAND U2308 ( .A(n1619), .B(n1621), .Z(n10296) );
  XOR U2309 ( .A(n10312), .B(sreg[1791]), .Z(n1622) );
  NANDN U2310 ( .A(n10313), .B(n1622), .Z(n1623) );
  NAND U2311 ( .A(n10312), .B(sreg[1791]), .Z(n1624) );
  AND U2312 ( .A(n1623), .B(n1624), .Z(n10322) );
  NAND U2313 ( .A(n10340), .B(sreg[1794]), .Z(n1625) );
  XOR U2314 ( .A(sreg[1794]), .B(n10340), .Z(n1626) );
  NANDN U2315 ( .A(n10341), .B(n1626), .Z(n1627) );
  NAND U2316 ( .A(n1625), .B(n1627), .Z(n10349) );
  XOR U2317 ( .A(n10365), .B(sreg[1797]), .Z(n1628) );
  NANDN U2318 ( .A(n10366), .B(n1628), .Z(n1629) );
  NAND U2319 ( .A(n10365), .B(sreg[1797]), .Z(n1630) );
  AND U2320 ( .A(n1629), .B(n1630), .Z(n10372) );
  NAND U2321 ( .A(n10389), .B(sreg[1800]), .Z(n1631) );
  XOR U2322 ( .A(sreg[1800]), .B(n10389), .Z(n1632) );
  NANDN U2323 ( .A(n10388), .B(n1632), .Z(n1633) );
  NAND U2324 ( .A(n1631), .B(n1633), .Z(n10397) );
  XOR U2325 ( .A(n10413), .B(sreg[1803]), .Z(n1634) );
  NANDN U2326 ( .A(n10414), .B(n1634), .Z(n1635) );
  NAND U2327 ( .A(n10413), .B(sreg[1803]), .Z(n1636) );
  AND U2328 ( .A(n1635), .B(n1636), .Z(n10420) );
  NAND U2329 ( .A(n10437), .B(sreg[1806]), .Z(n1637) );
  XOR U2330 ( .A(sreg[1806]), .B(n10437), .Z(n1638) );
  NANDN U2331 ( .A(n10436), .B(n1638), .Z(n1639) );
  NAND U2332 ( .A(n1637), .B(n1639), .Z(n10445) );
  XOR U2333 ( .A(n10464), .B(sreg[1809]), .Z(n1640) );
  NANDN U2334 ( .A(n10465), .B(n1640), .Z(n1641) );
  NAND U2335 ( .A(n10464), .B(sreg[1809]), .Z(n1642) );
  AND U2336 ( .A(n1641), .B(n1642), .Z(n10471) );
  NAND U2337 ( .A(n10486), .B(sreg[1812]), .Z(n1643) );
  XOR U2338 ( .A(sreg[1812]), .B(n10486), .Z(n1644) );
  NAND U2339 ( .A(n1644), .B(n10485), .Z(n1645) );
  NAND U2340 ( .A(n1643), .B(n1645), .Z(n10494) );
  XOR U2341 ( .A(n10510), .B(sreg[1815]), .Z(n1646) );
  NANDN U2342 ( .A(n10511), .B(n1646), .Z(n1647) );
  NAND U2343 ( .A(n10510), .B(sreg[1815]), .Z(n1648) );
  AND U2344 ( .A(n1647), .B(n1648), .Z(n10517) );
  NAND U2345 ( .A(n10534), .B(sreg[1818]), .Z(n1649) );
  XOR U2346 ( .A(sreg[1818]), .B(n10534), .Z(n1650) );
  NANDN U2347 ( .A(n10533), .B(n1650), .Z(n1651) );
  NAND U2348 ( .A(n1649), .B(n1651), .Z(n10542) );
  XOR U2349 ( .A(n10561), .B(sreg[1821]), .Z(n1652) );
  NANDN U2350 ( .A(n10562), .B(n1652), .Z(n1653) );
  NAND U2351 ( .A(n10561), .B(sreg[1821]), .Z(n1654) );
  AND U2352 ( .A(n1653), .B(n1654), .Z(n10568) );
  NAND U2353 ( .A(n10585), .B(sreg[1824]), .Z(n1655) );
  XOR U2354 ( .A(sreg[1824]), .B(n10585), .Z(n1656) );
  NANDN U2355 ( .A(n10584), .B(n1656), .Z(n1657) );
  NAND U2356 ( .A(n1655), .B(n1657), .Z(n10593) );
  XOR U2357 ( .A(n10609), .B(sreg[1827]), .Z(n1658) );
  NANDN U2358 ( .A(n10610), .B(n1658), .Z(n1659) );
  NAND U2359 ( .A(n10609), .B(sreg[1827]), .Z(n1660) );
  AND U2360 ( .A(n1659), .B(n1660), .Z(n10616) );
  NAND U2361 ( .A(n10631), .B(sreg[1830]), .Z(n1661) );
  XOR U2362 ( .A(sreg[1830]), .B(n10631), .Z(n1662) );
  NAND U2363 ( .A(n1662), .B(n10630), .Z(n1663) );
  NAND U2364 ( .A(n1661), .B(n1663), .Z(n10639) );
  XOR U2365 ( .A(n10657), .B(sreg[1833]), .Z(n1664) );
  NANDN U2366 ( .A(n10658), .B(n1664), .Z(n1665) );
  NAND U2367 ( .A(n10657), .B(sreg[1833]), .Z(n1666) );
  AND U2368 ( .A(n1665), .B(n1666), .Z(n10667) );
  NAND U2369 ( .A(n10684), .B(sreg[1836]), .Z(n1667) );
  XOR U2370 ( .A(sreg[1836]), .B(n10684), .Z(n1668) );
  NANDN U2371 ( .A(n10683), .B(n1668), .Z(n1669) );
  NAND U2372 ( .A(n1667), .B(n1669), .Z(n10690) );
  XOR U2373 ( .A(n10706), .B(sreg[1839]), .Z(n1670) );
  NANDN U2374 ( .A(n10707), .B(n1670), .Z(n1671) );
  NAND U2375 ( .A(n10706), .B(sreg[1839]), .Z(n1672) );
  AND U2376 ( .A(n1671), .B(n1672), .Z(n10713) );
  NAND U2377 ( .A(n10730), .B(sreg[1842]), .Z(n1673) );
  XOR U2378 ( .A(sreg[1842]), .B(n10730), .Z(n1674) );
  NANDN U2379 ( .A(n10729), .B(n1674), .Z(n1675) );
  NAND U2380 ( .A(n1673), .B(n1675), .Z(n10736) );
  XOR U2381 ( .A(n10754), .B(sreg[1845]), .Z(n1676) );
  NANDN U2382 ( .A(n10755), .B(n1676), .Z(n1677) );
  NAND U2383 ( .A(n10754), .B(sreg[1845]), .Z(n1678) );
  AND U2384 ( .A(n1677), .B(n1678), .Z(n10764) );
  XOR U2385 ( .A(n10782), .B(sreg[1848]), .Z(n1679) );
  NANDN U2386 ( .A(n10783), .B(n1679), .Z(n1680) );
  NAND U2387 ( .A(n10782), .B(sreg[1848]), .Z(n1681) );
  AND U2388 ( .A(n1680), .B(n1681), .Z(n10789) );
  XOR U2389 ( .A(n10807), .B(sreg[1851]), .Z(n1682) );
  NANDN U2390 ( .A(n10808), .B(n1682), .Z(n1683) );
  NAND U2391 ( .A(n10807), .B(sreg[1851]), .Z(n1684) );
  AND U2392 ( .A(n1683), .B(n1684), .Z(n10814) );
  NAND U2393 ( .A(n10831), .B(sreg[1854]), .Z(n1685) );
  XOR U2394 ( .A(sreg[1854]), .B(n10831), .Z(n1686) );
  NANDN U2395 ( .A(n10830), .B(n1686), .Z(n1687) );
  NAND U2396 ( .A(n1685), .B(n1687), .Z(n10839) );
  NAND U2397 ( .A(n10855), .B(sreg[1857]), .Z(n1688) );
  XOR U2398 ( .A(sreg[1857]), .B(n10855), .Z(n1689) );
  NANDN U2399 ( .A(n10856), .B(n1689), .Z(n1690) );
  NAND U2400 ( .A(n1688), .B(n1690), .Z(n10864) );
  NAND U2401 ( .A(n10880), .B(sreg[1860]), .Z(n1691) );
  XOR U2402 ( .A(sreg[1860]), .B(n10880), .Z(n1692) );
  NANDN U2403 ( .A(n10881), .B(n1692), .Z(n1693) );
  NAND U2404 ( .A(n1691), .B(n1693), .Z(n10889) );
  NAND U2405 ( .A(n10906), .B(sreg[1863]), .Z(n1694) );
  XOR U2406 ( .A(sreg[1863]), .B(n10906), .Z(n1695) );
  NANDN U2407 ( .A(n10905), .B(n1695), .Z(n1696) );
  NAND U2408 ( .A(n1694), .B(n1696), .Z(n10914) );
  NAND U2409 ( .A(n10934), .B(sreg[1866]), .Z(n1697) );
  XOR U2410 ( .A(sreg[1866]), .B(n10934), .Z(n1698) );
  NANDN U2411 ( .A(n10933), .B(n1698), .Z(n1699) );
  NAND U2412 ( .A(n1697), .B(n1699), .Z(n10942) );
  XOR U2413 ( .A(n10958), .B(sreg[1869]), .Z(n1700) );
  NANDN U2414 ( .A(n10959), .B(n1700), .Z(n1701) );
  NAND U2415 ( .A(n10958), .B(sreg[1869]), .Z(n1702) );
  AND U2416 ( .A(n1701), .B(n1702), .Z(n10965) );
  NAND U2417 ( .A(n10982), .B(sreg[1872]), .Z(n1703) );
  XOR U2418 ( .A(sreg[1872]), .B(n10982), .Z(n1704) );
  NANDN U2419 ( .A(n10981), .B(n1704), .Z(n1705) );
  NAND U2420 ( .A(n1703), .B(n1705), .Z(n10988) );
  NAND U2421 ( .A(n11004), .B(sreg[1875]), .Z(n1706) );
  XOR U2422 ( .A(sreg[1875]), .B(n11004), .Z(n1707) );
  NANDN U2423 ( .A(n11005), .B(n1707), .Z(n1708) );
  NAND U2424 ( .A(n1706), .B(n1708), .Z(n11013) );
  NAND U2425 ( .A(n11031), .B(sreg[1878]), .Z(n1709) );
  XOR U2426 ( .A(sreg[1878]), .B(n11031), .Z(n1710) );
  NANDN U2427 ( .A(n11032), .B(n1710), .Z(n1711) );
  NAND U2428 ( .A(n1709), .B(n1711), .Z(n11040) );
  XOR U2429 ( .A(n11058), .B(sreg[1881]), .Z(n1712) );
  NANDN U2430 ( .A(n11059), .B(n1712), .Z(n1713) );
  NAND U2431 ( .A(n11058), .B(sreg[1881]), .Z(n1714) );
  AND U2432 ( .A(n1713), .B(n1714), .Z(n11065) );
  NAND U2433 ( .A(n11083), .B(sreg[1884]), .Z(n1715) );
  XOR U2434 ( .A(sreg[1884]), .B(n11083), .Z(n1716) );
  NANDN U2435 ( .A(n11084), .B(n1716), .Z(n1717) );
  NAND U2436 ( .A(n1715), .B(n1717), .Z(n11092) );
  XOR U2437 ( .A(n11111), .B(sreg[1887]), .Z(n1718) );
  NANDN U2438 ( .A(n11112), .B(n1718), .Z(n1719) );
  NAND U2439 ( .A(n11111), .B(sreg[1887]), .Z(n1720) );
  AND U2440 ( .A(n1719), .B(n1720), .Z(n11118) );
  NAND U2441 ( .A(n11135), .B(sreg[1890]), .Z(n1721) );
  XOR U2442 ( .A(sreg[1890]), .B(n11135), .Z(n1722) );
  NANDN U2443 ( .A(n11134), .B(n1722), .Z(n1723) );
  NAND U2444 ( .A(n1721), .B(n1723), .Z(n11143) );
  XOR U2445 ( .A(n11159), .B(sreg[1893]), .Z(n1724) );
  NANDN U2446 ( .A(n11160), .B(n1724), .Z(n1725) );
  NAND U2447 ( .A(n11159), .B(sreg[1893]), .Z(n1726) );
  AND U2448 ( .A(n1725), .B(n1726), .Z(n11166) );
  NAND U2449 ( .A(n11181), .B(sreg[1896]), .Z(n1727) );
  XOR U2450 ( .A(sreg[1896]), .B(n11181), .Z(n1728) );
  NAND U2451 ( .A(n1728), .B(n11180), .Z(n1729) );
  NAND U2452 ( .A(n1727), .B(n1729), .Z(n11189) );
  NAND U2453 ( .A(n11207), .B(sreg[1899]), .Z(n1730) );
  XOR U2454 ( .A(sreg[1899]), .B(n11207), .Z(n1731) );
  NAND U2455 ( .A(n1731), .B(n11206), .Z(n1732) );
  NAND U2456 ( .A(n1730), .B(n1732), .Z(n11213) );
  NAND U2457 ( .A(n11230), .B(sreg[1902]), .Z(n1733) );
  XOR U2458 ( .A(sreg[1902]), .B(n11230), .Z(n1734) );
  NANDN U2459 ( .A(n11229), .B(n1734), .Z(n1735) );
  NAND U2460 ( .A(n1733), .B(n1735), .Z(n11238) );
  XOR U2461 ( .A(n11254), .B(sreg[1905]), .Z(n1736) );
  NANDN U2462 ( .A(n11255), .B(n1736), .Z(n1737) );
  NAND U2463 ( .A(n11254), .B(sreg[1905]), .Z(n1738) );
  AND U2464 ( .A(n1737), .B(n1738), .Z(n11261) );
  NAND U2465 ( .A(n11278), .B(sreg[1908]), .Z(n1739) );
  XOR U2466 ( .A(sreg[1908]), .B(n11278), .Z(n1740) );
  NANDN U2467 ( .A(n11277), .B(n1740), .Z(n1741) );
  NAND U2468 ( .A(n1739), .B(n1741), .Z(n11286) );
  XOR U2469 ( .A(n11305), .B(sreg[1911]), .Z(n1742) );
  NANDN U2470 ( .A(n11306), .B(n1742), .Z(n1743) );
  NAND U2471 ( .A(n11305), .B(sreg[1911]), .Z(n1744) );
  AND U2472 ( .A(n1743), .B(n1744), .Z(n11312) );
  NAND U2473 ( .A(n11329), .B(sreg[1914]), .Z(n1745) );
  XOR U2474 ( .A(sreg[1914]), .B(n11329), .Z(n1746) );
  NANDN U2475 ( .A(n11328), .B(n1746), .Z(n1747) );
  NAND U2476 ( .A(n1745), .B(n1747), .Z(n11337) );
  NAND U2477 ( .A(n11353), .B(sreg[1917]), .Z(n1748) );
  XOR U2478 ( .A(sreg[1917]), .B(n11353), .Z(n1749) );
  NANDN U2479 ( .A(n11354), .B(n1749), .Z(n1750) );
  NAND U2480 ( .A(n1748), .B(n1750), .Z(n11362) );
  NAND U2481 ( .A(n11380), .B(sreg[1920]), .Z(n1751) );
  XOR U2482 ( .A(sreg[1920]), .B(n11380), .Z(n1752) );
  NANDN U2483 ( .A(n11381), .B(n1752), .Z(n1753) );
  NAND U2484 ( .A(n1751), .B(n1753), .Z(n11389) );
  NAND U2485 ( .A(n11405), .B(sreg[1923]), .Z(n1754) );
  XOR U2486 ( .A(sreg[1923]), .B(n11405), .Z(n1755) );
  NANDN U2487 ( .A(n11406), .B(n1755), .Z(n1756) );
  NAND U2488 ( .A(n1754), .B(n1756), .Z(n11414) );
  NAND U2489 ( .A(n11429), .B(sreg[1926]), .Z(n1757) );
  XOR U2490 ( .A(sreg[1926]), .B(n11429), .Z(n1758) );
  NAND U2491 ( .A(n1758), .B(n11428), .Z(n1759) );
  NAND U2492 ( .A(n1757), .B(n1759), .Z(n11437) );
  XOR U2493 ( .A(n11455), .B(sreg[1929]), .Z(n1760) );
  NANDN U2494 ( .A(n11456), .B(n1760), .Z(n1761) );
  NAND U2495 ( .A(n11455), .B(sreg[1929]), .Z(n1762) );
  AND U2496 ( .A(n1761), .B(n1762), .Z(n11465) );
  NAND U2497 ( .A(n11482), .B(sreg[1932]), .Z(n1763) );
  XOR U2498 ( .A(sreg[1932]), .B(n11482), .Z(n1764) );
  NANDN U2499 ( .A(n11481), .B(n1764), .Z(n1765) );
  NAND U2500 ( .A(n1763), .B(n1765), .Z(n11490) );
  XOR U2501 ( .A(n11508), .B(sreg[1935]), .Z(n1766) );
  NANDN U2502 ( .A(n11509), .B(n1766), .Z(n1767) );
  NAND U2503 ( .A(n11508), .B(sreg[1935]), .Z(n1768) );
  AND U2504 ( .A(n1767), .B(n1768), .Z(n11515) );
  NAND U2505 ( .A(n11532), .B(sreg[1938]), .Z(n1769) );
  XOR U2506 ( .A(sreg[1938]), .B(n11532), .Z(n1770) );
  NANDN U2507 ( .A(n11531), .B(n1770), .Z(n1771) );
  NAND U2508 ( .A(n1769), .B(n1771), .Z(n11538) );
  NAND U2509 ( .A(n11554), .B(sreg[1941]), .Z(n1772) );
  XOR U2510 ( .A(sreg[1941]), .B(n11554), .Z(n1773) );
  NANDN U2511 ( .A(n11555), .B(n1773), .Z(n1774) );
  NAND U2512 ( .A(n1772), .B(n1774), .Z(n11563) );
  NAND U2513 ( .A(n11580), .B(sreg[1944]), .Z(n1775) );
  XOR U2514 ( .A(sreg[1944]), .B(n11580), .Z(n1776) );
  NANDN U2515 ( .A(n11579), .B(n1776), .Z(n1777) );
  NAND U2516 ( .A(n1775), .B(n1777), .Z(n11588) );
  XOR U2517 ( .A(n11607), .B(sreg[1947]), .Z(n1778) );
  NANDN U2518 ( .A(n11608), .B(n1778), .Z(n1779) );
  NAND U2519 ( .A(n11607), .B(sreg[1947]), .Z(n1780) );
  AND U2520 ( .A(n1779), .B(n1780), .Z(n11614) );
  NAND U2521 ( .A(n11631), .B(sreg[1950]), .Z(n1781) );
  XOR U2522 ( .A(sreg[1950]), .B(n11631), .Z(n1782) );
  NANDN U2523 ( .A(n11630), .B(n1782), .Z(n1783) );
  NAND U2524 ( .A(n1781), .B(n1783), .Z(n11639) );
  NAND U2525 ( .A(n11655), .B(sreg[1953]), .Z(n1784) );
  XOR U2526 ( .A(sreg[1953]), .B(n11655), .Z(n1785) );
  NANDN U2527 ( .A(n11656), .B(n1785), .Z(n1786) );
  NAND U2528 ( .A(n1784), .B(n1786), .Z(n11664) );
  NAND U2529 ( .A(n11681), .B(sreg[1956]), .Z(n1787) );
  XOR U2530 ( .A(sreg[1956]), .B(n11681), .Z(n1788) );
  NANDN U2531 ( .A(n11680), .B(n1788), .Z(n1789) );
  NAND U2532 ( .A(n1787), .B(n1789), .Z(n11689) );
  NAND U2533 ( .A(n11704), .B(sreg[1959]), .Z(n1790) );
  XOR U2534 ( .A(sreg[1959]), .B(n11704), .Z(n1791) );
  NAND U2535 ( .A(n1791), .B(n11703), .Z(n1792) );
  NAND U2536 ( .A(n1790), .B(n1792), .Z(n11712) );
  NAND U2537 ( .A(n11732), .B(sreg[1962]), .Z(n1793) );
  XOR U2538 ( .A(sreg[1962]), .B(n11732), .Z(n1794) );
  NANDN U2539 ( .A(n11731), .B(n1794), .Z(n1795) );
  NAND U2540 ( .A(n1793), .B(n1795), .Z(n11740) );
  XOR U2541 ( .A(n11756), .B(sreg[1965]), .Z(n1796) );
  NANDN U2542 ( .A(n11757), .B(n1796), .Z(n1797) );
  NAND U2543 ( .A(n11756), .B(sreg[1965]), .Z(n1798) );
  AND U2544 ( .A(n1797), .B(n1798), .Z(n11763) );
  NAND U2545 ( .A(n11781), .B(sreg[1968]), .Z(n1799) );
  XOR U2546 ( .A(sreg[1968]), .B(n11781), .Z(n1800) );
  NANDN U2547 ( .A(n11782), .B(n1800), .Z(n1801) );
  NAND U2548 ( .A(n1799), .B(n1801), .Z(n11790) );
  NAND U2549 ( .A(n11808), .B(sreg[1971]), .Z(n1802) );
  XOR U2550 ( .A(sreg[1971]), .B(n11808), .Z(n1803) );
  NANDN U2551 ( .A(n11809), .B(n1803), .Z(n1804) );
  NAND U2552 ( .A(n1802), .B(n1804), .Z(n11817) );
  NAND U2553 ( .A(n11834), .B(sreg[1974]), .Z(n1805) );
  XOR U2554 ( .A(sreg[1974]), .B(n11834), .Z(n1806) );
  NANDN U2555 ( .A(n11833), .B(n1806), .Z(n1807) );
  NAND U2556 ( .A(n1805), .B(n1807), .Z(n11842) );
  XOR U2557 ( .A(n11858), .B(sreg[1977]), .Z(n1808) );
  NANDN U2558 ( .A(n11859), .B(n1808), .Z(n1809) );
  NAND U2559 ( .A(n11858), .B(sreg[1977]), .Z(n1810) );
  AND U2560 ( .A(n1809), .B(n1810), .Z(n11865) );
  NAND U2561 ( .A(n11882), .B(sreg[1980]), .Z(n1811) );
  XOR U2562 ( .A(sreg[1980]), .B(n11882), .Z(n1812) );
  NANDN U2563 ( .A(n11881), .B(n1812), .Z(n1813) );
  NAND U2564 ( .A(n1811), .B(n1813), .Z(n11890) );
  XOR U2565 ( .A(n11909), .B(sreg[1983]), .Z(n1814) );
  NANDN U2566 ( .A(n11910), .B(n1814), .Z(n1815) );
  NAND U2567 ( .A(n11909), .B(sreg[1983]), .Z(n1816) );
  AND U2568 ( .A(n1815), .B(n1816), .Z(n11916) );
  NAND U2569 ( .A(n11933), .B(sreg[1986]), .Z(n1817) );
  XOR U2570 ( .A(sreg[1986]), .B(n11933), .Z(n1818) );
  NANDN U2571 ( .A(n11932), .B(n1818), .Z(n1819) );
  NAND U2572 ( .A(n1817), .B(n1819), .Z(n11941) );
  XOR U2573 ( .A(n11957), .B(sreg[1989]), .Z(n1820) );
  NANDN U2574 ( .A(n11958), .B(n1820), .Z(n1821) );
  NAND U2575 ( .A(n11957), .B(sreg[1989]), .Z(n1822) );
  AND U2576 ( .A(n1821), .B(n1822), .Z(n11964) );
  NAND U2577 ( .A(n11981), .B(sreg[1992]), .Z(n1823) );
  XOR U2578 ( .A(sreg[1992]), .B(n11981), .Z(n1824) );
  NANDN U2579 ( .A(n11980), .B(n1824), .Z(n1825) );
  NAND U2580 ( .A(n1823), .B(n1825), .Z(n11989) );
  XOR U2581 ( .A(n12005), .B(sreg[1995]), .Z(n1826) );
  NANDN U2582 ( .A(n12006), .B(n1826), .Z(n1827) );
  NAND U2583 ( .A(n12005), .B(sreg[1995]), .Z(n1828) );
  AND U2584 ( .A(n1827), .B(n1828), .Z(n12015) );
  NAND U2585 ( .A(n12031), .B(sreg[1998]), .Z(n1829) );
  XOR U2586 ( .A(sreg[1998]), .B(n12031), .Z(n1830) );
  NANDN U2587 ( .A(n12032), .B(n1830), .Z(n1831) );
  NAND U2588 ( .A(n1829), .B(n1831), .Z(n12040) );
  XOR U2589 ( .A(n12056), .B(sreg[2001]), .Z(n1832) );
  NANDN U2590 ( .A(n12057), .B(n1832), .Z(n1833) );
  NAND U2591 ( .A(n12056), .B(sreg[2001]), .Z(n1834) );
  AND U2592 ( .A(n1833), .B(n1834), .Z(n12063) );
  NAND U2593 ( .A(n12080), .B(sreg[2004]), .Z(n1835) );
  XOR U2594 ( .A(sreg[2004]), .B(n12080), .Z(n1836) );
  NANDN U2595 ( .A(n12079), .B(n1836), .Z(n1837) );
  NAND U2596 ( .A(n1835), .B(n1837), .Z(n12086) );
  XOR U2597 ( .A(n12102), .B(sreg[2007]), .Z(n1838) );
  NANDN U2598 ( .A(n12103), .B(n1838), .Z(n1839) );
  NAND U2599 ( .A(n12102), .B(sreg[2007]), .Z(n1840) );
  AND U2600 ( .A(n1839), .B(n1840), .Z(n12112) );
  NAND U2601 ( .A(n12127), .B(sreg[2010]), .Z(n1841) );
  XOR U2602 ( .A(sreg[2010]), .B(n12127), .Z(n1842) );
  NAND U2603 ( .A(n1842), .B(n12126), .Z(n1843) );
  NAND U2604 ( .A(n1841), .B(n1843), .Z(n12135) );
  XOR U2605 ( .A(n12151), .B(sreg[2013]), .Z(n1844) );
  NANDN U2606 ( .A(n12152), .B(n1844), .Z(n1845) );
  NAND U2607 ( .A(n12151), .B(sreg[2013]), .Z(n1846) );
  AND U2608 ( .A(n1845), .B(n1846), .Z(n12158) );
  NAND U2609 ( .A(n12175), .B(sreg[2016]), .Z(n1847) );
  XOR U2610 ( .A(sreg[2016]), .B(n12175), .Z(n1848) );
  NANDN U2611 ( .A(n12174), .B(n1848), .Z(n1849) );
  NAND U2612 ( .A(n1847), .B(n1849), .Z(n12183) );
  XOR U2613 ( .A(n12199), .B(sreg[2019]), .Z(n1850) );
  NANDN U2614 ( .A(n12200), .B(n1850), .Z(n1851) );
  NAND U2615 ( .A(n12199), .B(sreg[2019]), .Z(n1852) );
  AND U2616 ( .A(n1851), .B(n1852), .Z(n12209) );
  NAND U2617 ( .A(n12224), .B(sreg[2022]), .Z(n1853) );
  XOR U2618 ( .A(sreg[2022]), .B(n12224), .Z(n1854) );
  NAND U2619 ( .A(n1854), .B(n12223), .Z(n1855) );
  NAND U2620 ( .A(n1853), .B(n1855), .Z(n12232) );
  XOR U2621 ( .A(n12250), .B(sreg[2025]), .Z(n1856) );
  NANDN U2622 ( .A(n12251), .B(n1856), .Z(n1857) );
  NAND U2623 ( .A(n12250), .B(sreg[2025]), .Z(n1858) );
  AND U2624 ( .A(n1857), .B(n1858), .Z(n12257) );
  NAND U2625 ( .A(n12274), .B(sreg[2028]), .Z(n1859) );
  XOR U2626 ( .A(sreg[2028]), .B(n12274), .Z(n1860) );
  NANDN U2627 ( .A(n12273), .B(n1860), .Z(n1861) );
  NAND U2628 ( .A(n1859), .B(n1861), .Z(n12280) );
  XOR U2629 ( .A(n12298), .B(sreg[2031]), .Z(n1862) );
  NANDN U2630 ( .A(n12299), .B(n1862), .Z(n1863) );
  NAND U2631 ( .A(n12298), .B(sreg[2031]), .Z(n1864) );
  AND U2632 ( .A(n1863), .B(n1864), .Z(n12305) );
  NAND U2633 ( .A(n12323), .B(sreg[2034]), .Z(n1865) );
  XOR U2634 ( .A(sreg[2034]), .B(n12323), .Z(n1866) );
  NANDN U2635 ( .A(n12324), .B(n1866), .Z(n1867) );
  NAND U2636 ( .A(n1865), .B(n1867), .Z(n12332) );
  XOR U2637 ( .A(n12348), .B(sreg[2037]), .Z(n1868) );
  NANDN U2638 ( .A(n12349), .B(n1868), .Z(n1869) );
  NAND U2639 ( .A(n12348), .B(sreg[2037]), .Z(n1870) );
  AND U2640 ( .A(n1869), .B(n1870), .Z(n12355) );
  NAND U2641 ( .A(n12372), .B(sreg[2040]), .Z(n1871) );
  XOR U2642 ( .A(sreg[2040]), .B(n12372), .Z(n1872) );
  NANDN U2643 ( .A(n12371), .B(n1872), .Z(n1873) );
  NAND U2644 ( .A(n1871), .B(n1873), .Z(n12380) );
  NAND U2645 ( .A(n12396), .B(sreg[2043]), .Z(n1874) );
  XOR U2646 ( .A(sreg[2043]), .B(n12396), .Z(n1875) );
  NANDN U2647 ( .A(n12397), .B(n1875), .Z(n1876) );
  NAND U2648 ( .A(n1874), .B(n1876), .Z(n12407) );
  NAND U2649 ( .A(n4022), .B(sreg[1026]), .Z(n1877) );
  XOR U2650 ( .A(sreg[1026]), .B(n4022), .Z(n1878) );
  NANDN U2651 ( .A(n4023), .B(n1878), .Z(n1879) );
  NAND U2652 ( .A(n1877), .B(n1879), .Z(n4025) );
  XOR U2653 ( .A(n4052), .B(sreg[1029]), .Z(n1880) );
  NANDN U2654 ( .A(n4051), .B(n1880), .Z(n1881) );
  NAND U2655 ( .A(n4052), .B(sreg[1029]), .Z(n1882) );
  AND U2656 ( .A(n1881), .B(n1882), .Z(n4060) );
  NAND U2657 ( .A(n4076), .B(sreg[1032]), .Z(n1883) );
  XOR U2658 ( .A(sreg[1032]), .B(n4076), .Z(n1884) );
  NANDN U2659 ( .A(n4077), .B(n1884), .Z(n1885) );
  NAND U2660 ( .A(n1883), .B(n1885), .Z(n4085) );
  XOR U2661 ( .A(n4101), .B(sreg[1035]), .Z(n1886) );
  NANDN U2662 ( .A(n4102), .B(n1886), .Z(n1887) );
  NAND U2663 ( .A(n4101), .B(sreg[1035]), .Z(n1888) );
  AND U2664 ( .A(n1887), .B(n1888), .Z(n4108) );
  NAND U2665 ( .A(n4125), .B(sreg[1038]), .Z(n1889) );
  XOR U2666 ( .A(sreg[1038]), .B(n4125), .Z(n1890) );
  NANDN U2667 ( .A(n4124), .B(n1890), .Z(n1891) );
  NAND U2668 ( .A(n1889), .B(n1891), .Z(n4133) );
  NAND U2669 ( .A(n4168), .B(sreg[1043]), .Z(n1892) );
  XOR U2670 ( .A(sreg[1043]), .B(n4168), .Z(n1893) );
  NAND U2671 ( .A(n1893), .B(n4167), .Z(n1894) );
  NAND U2672 ( .A(n1892), .B(n1894), .Z(n4174) );
  XOR U2673 ( .A(n4192), .B(sreg[1046]), .Z(n1895) );
  NANDN U2674 ( .A(n4193), .B(n1895), .Z(n1896) );
  NAND U2675 ( .A(n4192), .B(sreg[1046]), .Z(n1897) );
  AND U2676 ( .A(n1896), .B(n1897), .Z(n4201) );
  XOR U2677 ( .A(n4237), .B(sreg[1051]), .Z(n1898) );
  NANDN U2678 ( .A(n4238), .B(n1898), .Z(n1899) );
  NAND U2679 ( .A(n4237), .B(sreg[1051]), .Z(n1900) );
  AND U2680 ( .A(n1899), .B(n1900), .Z(n4244) );
  NAND U2681 ( .A(n4264), .B(sreg[1054]), .Z(n1901) );
  XOR U2682 ( .A(sreg[1054]), .B(n4264), .Z(n1902) );
  NANDN U2683 ( .A(n4263), .B(n1902), .Z(n1903) );
  NAND U2684 ( .A(n1901), .B(n1903), .Z(n4272) );
  XOR U2685 ( .A(n4288), .B(sreg[1057]), .Z(n1904) );
  NANDN U2686 ( .A(n4289), .B(n1904), .Z(n1905) );
  NAND U2687 ( .A(n4288), .B(sreg[1057]), .Z(n1906) );
  AND U2688 ( .A(n1905), .B(n1906), .Z(n4295) );
  NAND U2689 ( .A(n4312), .B(sreg[1060]), .Z(n1907) );
  XOR U2690 ( .A(sreg[1060]), .B(n4312), .Z(n1908) );
  NANDN U2691 ( .A(n4311), .B(n1908), .Z(n1909) );
  NAND U2692 ( .A(n1907), .B(n1909), .Z(n4320) );
  XOR U2693 ( .A(n4336), .B(sreg[1063]), .Z(n1910) );
  NANDN U2694 ( .A(n4337), .B(n1910), .Z(n1911) );
  NAND U2695 ( .A(n4336), .B(sreg[1063]), .Z(n1912) );
  AND U2696 ( .A(n1911), .B(n1912), .Z(n4343) );
  NAND U2697 ( .A(n4361), .B(sreg[1066]), .Z(n1913) );
  XOR U2698 ( .A(sreg[1066]), .B(n4361), .Z(n1914) );
  NAND U2699 ( .A(n1914), .B(n4360), .Z(n1915) );
  NAND U2700 ( .A(n1913), .B(n1915), .Z(n4369) );
  XOR U2701 ( .A(n4387), .B(sreg[1069]), .Z(n1916) );
  NANDN U2702 ( .A(n4388), .B(n1916), .Z(n1917) );
  NAND U2703 ( .A(n4387), .B(sreg[1069]), .Z(n1918) );
  AND U2704 ( .A(n1917), .B(n1918), .Z(n4394) );
  NAND U2705 ( .A(n4411), .B(sreg[1072]), .Z(n1919) );
  XOR U2706 ( .A(sreg[1072]), .B(n4411), .Z(n1920) );
  NANDN U2707 ( .A(n4410), .B(n1920), .Z(n1921) );
  NAND U2708 ( .A(n1919), .B(n1921), .Z(n4419) );
  NAND U2709 ( .A(n4434), .B(sreg[1075]), .Z(n1922) );
  XOR U2710 ( .A(sreg[1075]), .B(n4434), .Z(n1923) );
  NAND U2711 ( .A(n1923), .B(n4433), .Z(n1924) );
  NAND U2712 ( .A(n1922), .B(n1924), .Z(n4440) );
  NAND U2713 ( .A(n4457), .B(sreg[1078]), .Z(n1925) );
  XOR U2714 ( .A(sreg[1078]), .B(n4457), .Z(n1926) );
  NANDN U2715 ( .A(n4456), .B(n1926), .Z(n1927) );
  NAND U2716 ( .A(n1925), .B(n1927), .Z(n4465) );
  XOR U2717 ( .A(n4484), .B(sreg[1081]), .Z(n1928) );
  NANDN U2718 ( .A(n4485), .B(n1928), .Z(n1929) );
  NAND U2719 ( .A(n4484), .B(sreg[1081]), .Z(n1930) );
  AND U2720 ( .A(n1929), .B(n1930), .Z(n4491) );
  NAND U2721 ( .A(n4509), .B(sreg[1084]), .Z(n1931) );
  XOR U2722 ( .A(sreg[1084]), .B(n4509), .Z(n1932) );
  NANDN U2723 ( .A(n4510), .B(n1932), .Z(n1933) );
  NAND U2724 ( .A(n1931), .B(n1933), .Z(n4518) );
  NAND U2725 ( .A(n4534), .B(sreg[1087]), .Z(n1934) );
  XOR U2726 ( .A(sreg[1087]), .B(n4534), .Z(n1935) );
  NANDN U2727 ( .A(n4535), .B(n1935), .Z(n1936) );
  NAND U2728 ( .A(n1934), .B(n1936), .Z(n4543) );
  NAND U2729 ( .A(n4560), .B(sreg[1090]), .Z(n1937) );
  XOR U2730 ( .A(sreg[1090]), .B(n4560), .Z(n1938) );
  NANDN U2731 ( .A(n4559), .B(n1938), .Z(n1939) );
  NAND U2732 ( .A(n1937), .B(n1939), .Z(n4568) );
  NAND U2733 ( .A(n4583), .B(sreg[1093]), .Z(n1940) );
  XOR U2734 ( .A(sreg[1093]), .B(n4583), .Z(n1941) );
  NAND U2735 ( .A(n1941), .B(n4582), .Z(n1942) );
  NAND U2736 ( .A(n1940), .B(n1942), .Z(n4589) );
  NAND U2737 ( .A(n4609), .B(sreg[1096]), .Z(n1943) );
  XOR U2738 ( .A(sreg[1096]), .B(n4609), .Z(n1944) );
  NANDN U2739 ( .A(n4608), .B(n1944), .Z(n1945) );
  NAND U2740 ( .A(n1943), .B(n1945), .Z(n4615) );
  NAND U2741 ( .A(n4630), .B(sreg[1099]), .Z(n1946) );
  XOR U2742 ( .A(sreg[1099]), .B(n4630), .Z(n1947) );
  NAND U2743 ( .A(n1947), .B(n4629), .Z(n1948) );
  NAND U2744 ( .A(n1946), .B(n1948), .Z(n4636) );
  NAND U2745 ( .A(n4653), .B(sreg[1102]), .Z(n1949) );
  XOR U2746 ( .A(sreg[1102]), .B(n4653), .Z(n1950) );
  NANDN U2747 ( .A(n4652), .B(n1950), .Z(n1951) );
  NAND U2748 ( .A(n1949), .B(n1951), .Z(n4661) );
  XOR U2749 ( .A(n4677), .B(sreg[1105]), .Z(n1952) );
  NANDN U2750 ( .A(n4678), .B(n1952), .Z(n1953) );
  NAND U2751 ( .A(n4677), .B(sreg[1105]), .Z(n1954) );
  AND U2752 ( .A(n1953), .B(n1954), .Z(n4687) );
  NAND U2753 ( .A(n4704), .B(sreg[1108]), .Z(n1955) );
  XOR U2754 ( .A(sreg[1108]), .B(n4704), .Z(n1956) );
  NANDN U2755 ( .A(n4703), .B(n1956), .Z(n1957) );
  NAND U2756 ( .A(n1955), .B(n1957), .Z(n4712) );
  XOR U2757 ( .A(n4728), .B(sreg[1111]), .Z(n1958) );
  NANDN U2758 ( .A(n4729), .B(n1958), .Z(n1959) );
  NAND U2759 ( .A(n4728), .B(sreg[1111]), .Z(n1960) );
  AND U2760 ( .A(n1959), .B(n1960), .Z(n4735) );
  NAND U2761 ( .A(n4752), .B(sreg[1114]), .Z(n1961) );
  XOR U2762 ( .A(sreg[1114]), .B(n4752), .Z(n1962) );
  NANDN U2763 ( .A(n4751), .B(n1962), .Z(n1963) );
  NAND U2764 ( .A(n1961), .B(n1963), .Z(n4760) );
  XOR U2765 ( .A(n4776), .B(sreg[1117]), .Z(n1964) );
  NANDN U2766 ( .A(n4777), .B(n1964), .Z(n1965) );
  NAND U2767 ( .A(n4776), .B(sreg[1117]), .Z(n1966) );
  AND U2768 ( .A(n1965), .B(n1966), .Z(n4783) );
  NAND U2769 ( .A(n4803), .B(sreg[1120]), .Z(n1967) );
  XOR U2770 ( .A(sreg[1120]), .B(n4803), .Z(n1968) );
  NANDN U2771 ( .A(n4802), .B(n1968), .Z(n1969) );
  NAND U2772 ( .A(n1967), .B(n1969), .Z(n4811) );
  XOR U2773 ( .A(n4829), .B(sreg[1123]), .Z(n1970) );
  NANDN U2774 ( .A(n4830), .B(n1970), .Z(n1971) );
  NAND U2775 ( .A(n4829), .B(sreg[1123]), .Z(n1972) );
  AND U2776 ( .A(n1971), .B(n1972), .Z(n4836) );
  NAND U2777 ( .A(n4853), .B(sreg[1126]), .Z(n1973) );
  XOR U2778 ( .A(sreg[1126]), .B(n4853), .Z(n1974) );
  NANDN U2779 ( .A(n4852), .B(n1974), .Z(n1975) );
  NAND U2780 ( .A(n1973), .B(n1975), .Z(n4861) );
  NAND U2781 ( .A(n4877), .B(sreg[1129]), .Z(n1976) );
  XOR U2782 ( .A(sreg[1129]), .B(n4877), .Z(n1977) );
  NANDN U2783 ( .A(n4878), .B(n1977), .Z(n1978) );
  NAND U2784 ( .A(n1976), .B(n1978), .Z(n4886) );
  NAND U2785 ( .A(n4901), .B(sreg[1132]), .Z(n1979) );
  XOR U2786 ( .A(sreg[1132]), .B(n4901), .Z(n1980) );
  NAND U2787 ( .A(n1980), .B(n4900), .Z(n1981) );
  NAND U2788 ( .A(n1979), .B(n1981), .Z(n4907) );
  NAND U2789 ( .A(n4926), .B(sreg[1135]), .Z(n1982) );
  XOR U2790 ( .A(sreg[1135]), .B(n4926), .Z(n1983) );
  NANDN U2791 ( .A(n4927), .B(n1983), .Z(n1984) );
  NAND U2792 ( .A(n1982), .B(n1984), .Z(n4935) );
  NAND U2793 ( .A(n4953), .B(sreg[1138]), .Z(n1985) );
  XOR U2794 ( .A(sreg[1138]), .B(n4953), .Z(n1986) );
  NANDN U2795 ( .A(n4954), .B(n1986), .Z(n1987) );
  NAND U2796 ( .A(n1985), .B(n1987), .Z(n4962) );
  XOR U2797 ( .A(n4978), .B(sreg[1141]), .Z(n1988) );
  NANDN U2798 ( .A(n4979), .B(n1988), .Z(n1989) );
  NAND U2799 ( .A(n4978), .B(sreg[1141]), .Z(n1990) );
  AND U2800 ( .A(n1989), .B(n1990), .Z(n4985) );
  NAND U2801 ( .A(n5002), .B(sreg[1144]), .Z(n1991) );
  XOR U2802 ( .A(sreg[1144]), .B(n5002), .Z(n1992) );
  NANDN U2803 ( .A(n5001), .B(n1992), .Z(n1993) );
  NAND U2804 ( .A(n1991), .B(n1993), .Z(n5010) );
  XOR U2805 ( .A(n5028), .B(sreg[1147]), .Z(n1994) );
  NANDN U2806 ( .A(n5029), .B(n1994), .Z(n1995) );
  NAND U2807 ( .A(n5028), .B(sreg[1147]), .Z(n1996) );
  AND U2808 ( .A(n1995), .B(n1996), .Z(n5035) );
  NAND U2809 ( .A(n5052), .B(sreg[1150]), .Z(n1997) );
  XOR U2810 ( .A(sreg[1150]), .B(n5052), .Z(n1998) );
  NANDN U2811 ( .A(n5051), .B(n1998), .Z(n1999) );
  NAND U2812 ( .A(n1997), .B(n1999), .Z(n5060) );
  XOR U2813 ( .A(n5076), .B(sreg[1153]), .Z(n2000) );
  NANDN U2814 ( .A(n5077), .B(n2000), .Z(n2001) );
  NAND U2815 ( .A(n5076), .B(sreg[1153]), .Z(n2002) );
  AND U2816 ( .A(n2001), .B(n2002), .Z(n5086) );
  NAND U2817 ( .A(n5104), .B(sreg[1156]), .Z(n2003) );
  XOR U2818 ( .A(sreg[1156]), .B(n5104), .Z(n2004) );
  NANDN U2819 ( .A(n5105), .B(n2004), .Z(n2005) );
  NAND U2820 ( .A(n2003), .B(n2005), .Z(n5113) );
  XOR U2821 ( .A(n5131), .B(sreg[1159]), .Z(n2006) );
  NANDN U2822 ( .A(n5132), .B(n2006), .Z(n2007) );
  NAND U2823 ( .A(n5131), .B(sreg[1159]), .Z(n2008) );
  AND U2824 ( .A(n2007), .B(n2008), .Z(n5138) );
  NAND U2825 ( .A(n5155), .B(sreg[1162]), .Z(n2009) );
  XOR U2826 ( .A(sreg[1162]), .B(n5155), .Z(n2010) );
  NANDN U2827 ( .A(n5154), .B(n2010), .Z(n2011) );
  NAND U2828 ( .A(n2009), .B(n2011), .Z(n5163) );
  XOR U2829 ( .A(n5181), .B(sreg[1165]), .Z(n2012) );
  NANDN U2830 ( .A(n5182), .B(n2012), .Z(n2013) );
  NAND U2831 ( .A(n5181), .B(sreg[1165]), .Z(n2014) );
  AND U2832 ( .A(n2013), .B(n2014), .Z(n5188) );
  NAND U2833 ( .A(n5205), .B(sreg[1168]), .Z(n2015) );
  XOR U2834 ( .A(sreg[1168]), .B(n5205), .Z(n2016) );
  NANDN U2835 ( .A(n5204), .B(n2016), .Z(n2017) );
  NAND U2836 ( .A(n2015), .B(n2017), .Z(n5213) );
  NAND U2837 ( .A(n5228), .B(sreg[1171]), .Z(n2018) );
  XOR U2838 ( .A(sreg[1171]), .B(n5228), .Z(n2019) );
  NAND U2839 ( .A(n2019), .B(n5227), .Z(n2020) );
  NAND U2840 ( .A(n2018), .B(n2020), .Z(n5237) );
  NAND U2841 ( .A(n5254), .B(sreg[1174]), .Z(n2021) );
  XOR U2842 ( .A(sreg[1174]), .B(n5254), .Z(n2022) );
  NANDN U2843 ( .A(n5253), .B(n2022), .Z(n2023) );
  NAND U2844 ( .A(n2021), .B(n2023), .Z(n5262) );
  XOR U2845 ( .A(n5278), .B(sreg[1177]), .Z(n2024) );
  NANDN U2846 ( .A(n5279), .B(n2024), .Z(n2025) );
  NAND U2847 ( .A(n5278), .B(sreg[1177]), .Z(n2026) );
  AND U2848 ( .A(n2025), .B(n2026), .Z(n5285) );
  NAND U2849 ( .A(n5302), .B(sreg[1180]), .Z(n2027) );
  XOR U2850 ( .A(sreg[1180]), .B(n5302), .Z(n2028) );
  NANDN U2851 ( .A(n5301), .B(n2028), .Z(n2029) );
  NAND U2852 ( .A(n2027), .B(n2029), .Z(n5310) );
  XOR U2853 ( .A(n5326), .B(sreg[1183]), .Z(n2030) );
  NANDN U2854 ( .A(n5327), .B(n2030), .Z(n2031) );
  NAND U2855 ( .A(n5326), .B(sreg[1183]), .Z(n2032) );
  AND U2856 ( .A(n2031), .B(n2032), .Z(n5333) );
  NAND U2857 ( .A(n5353), .B(sreg[1186]), .Z(n2033) );
  XOR U2858 ( .A(sreg[1186]), .B(n5353), .Z(n2034) );
  NANDN U2859 ( .A(n5352), .B(n2034), .Z(n2035) );
  NAND U2860 ( .A(n2033), .B(n2035), .Z(n5361) );
  XOR U2861 ( .A(n5377), .B(sreg[1189]), .Z(n2036) );
  NANDN U2862 ( .A(n5378), .B(n2036), .Z(n2037) );
  NAND U2863 ( .A(n5377), .B(sreg[1189]), .Z(n2038) );
  AND U2864 ( .A(n2037), .B(n2038), .Z(n5384) );
  NAND U2865 ( .A(n5399), .B(sreg[1192]), .Z(n2039) );
  XOR U2866 ( .A(sreg[1192]), .B(n5399), .Z(n2040) );
  NAND U2867 ( .A(n2040), .B(n5398), .Z(n2041) );
  NAND U2868 ( .A(n2039), .B(n2041), .Z(n5405) );
  XOR U2869 ( .A(n5421), .B(sreg[1195]), .Z(n2042) );
  NANDN U2870 ( .A(n5422), .B(n2042), .Z(n2043) );
  NAND U2871 ( .A(n5421), .B(sreg[1195]), .Z(n2044) );
  AND U2872 ( .A(n2043), .B(n2044), .Z(n5431) );
  NAND U2873 ( .A(n5449), .B(sreg[1198]), .Z(n2045) );
  XOR U2874 ( .A(sreg[1198]), .B(n5449), .Z(n2046) );
  NANDN U2875 ( .A(n5450), .B(n2046), .Z(n2047) );
  NAND U2876 ( .A(n2045), .B(n2047), .Z(n5458) );
  XOR U2877 ( .A(n5474), .B(sreg[1201]), .Z(n2048) );
  NANDN U2878 ( .A(n5475), .B(n2048), .Z(n2049) );
  NAND U2879 ( .A(n5474), .B(sreg[1201]), .Z(n2050) );
  AND U2880 ( .A(n2049), .B(n2050), .Z(n5481) );
  NAND U2881 ( .A(n5498), .B(sreg[1204]), .Z(n2051) );
  XOR U2882 ( .A(sreg[1204]), .B(n5498), .Z(n2052) );
  NANDN U2883 ( .A(n5497), .B(n2052), .Z(n2053) );
  NAND U2884 ( .A(n2051), .B(n2053), .Z(n5506) );
  XOR U2885 ( .A(n5522), .B(sreg[1207]), .Z(n2054) );
  NANDN U2886 ( .A(n5523), .B(n2054), .Z(n2055) );
  NAND U2887 ( .A(n5522), .B(sreg[1207]), .Z(n2056) );
  AND U2888 ( .A(n2055), .B(n2056), .Z(n5529) );
  NAND U2889 ( .A(n5547), .B(sreg[1210]), .Z(n2057) );
  XOR U2890 ( .A(sreg[1210]), .B(n5547), .Z(n2058) );
  NANDN U2891 ( .A(n5548), .B(n2058), .Z(n2059) );
  NAND U2892 ( .A(n2057), .B(n2059), .Z(n5556) );
  XOR U2893 ( .A(n5572), .B(sreg[1213]), .Z(n2060) );
  NANDN U2894 ( .A(n5573), .B(n2060), .Z(n2061) );
  NAND U2895 ( .A(n5572), .B(sreg[1213]), .Z(n2062) );
  AND U2896 ( .A(n2061), .B(n2062), .Z(n5582) );
  NAND U2897 ( .A(n5599), .B(sreg[1216]), .Z(n2063) );
  XOR U2898 ( .A(sreg[1216]), .B(n5599), .Z(n2064) );
  NANDN U2899 ( .A(n5598), .B(n2064), .Z(n2065) );
  NAND U2900 ( .A(n2063), .B(n2065), .Z(n5607) );
  XOR U2901 ( .A(n5623), .B(sreg[1219]), .Z(n2066) );
  NANDN U2902 ( .A(n5624), .B(n2066), .Z(n2067) );
  NAND U2903 ( .A(n5623), .B(sreg[1219]), .Z(n2068) );
  AND U2904 ( .A(n2067), .B(n2068), .Z(n5630) );
  NAND U2905 ( .A(n5647), .B(sreg[1222]), .Z(n2069) );
  XOR U2906 ( .A(sreg[1222]), .B(n5647), .Z(n2070) );
  NANDN U2907 ( .A(n5646), .B(n2070), .Z(n2071) );
  NAND U2908 ( .A(n2069), .B(n2071), .Z(n5653) );
  XOR U2909 ( .A(n5669), .B(sreg[1225]), .Z(n2072) );
  NANDN U2910 ( .A(n5670), .B(n2072), .Z(n2073) );
  NAND U2911 ( .A(n5669), .B(sreg[1225]), .Z(n2074) );
  AND U2912 ( .A(n2073), .B(n2074), .Z(n5679) );
  NAND U2913 ( .A(n5696), .B(sreg[1228]), .Z(n2075) );
  XOR U2914 ( .A(sreg[1228]), .B(n5696), .Z(n2076) );
  NANDN U2915 ( .A(n5695), .B(n2076), .Z(n2077) );
  NAND U2916 ( .A(n2075), .B(n2077), .Z(n5704) );
  XOR U2917 ( .A(n5720), .B(sreg[1231]), .Z(n2078) );
  NANDN U2918 ( .A(n5721), .B(n2078), .Z(n2079) );
  NAND U2919 ( .A(n5720), .B(sreg[1231]), .Z(n2080) );
  AND U2920 ( .A(n2079), .B(n2080), .Z(n5727) );
  NAND U2921 ( .A(n5744), .B(sreg[1234]), .Z(n2081) );
  XOR U2922 ( .A(sreg[1234]), .B(n5744), .Z(n2082) );
  NANDN U2923 ( .A(n5743), .B(n2082), .Z(n2083) );
  NAND U2924 ( .A(n2081), .B(n2083), .Z(n5752) );
  XOR U2925 ( .A(n5770), .B(sreg[1237]), .Z(n2084) );
  NANDN U2926 ( .A(n5771), .B(n2084), .Z(n2085) );
  NAND U2927 ( .A(n5770), .B(sreg[1237]), .Z(n2086) );
  AND U2928 ( .A(n2085), .B(n2086), .Z(n5777) );
  NAND U2929 ( .A(n5794), .B(sreg[1240]), .Z(n2087) );
  XOR U2930 ( .A(sreg[1240]), .B(n5794), .Z(n2088) );
  NANDN U2931 ( .A(n5793), .B(n2088), .Z(n2089) );
  NAND U2932 ( .A(n2087), .B(n2089), .Z(n5802) );
  XOR U2933 ( .A(n5820), .B(sreg[1243]), .Z(n2090) );
  NANDN U2934 ( .A(n5821), .B(n2090), .Z(n2091) );
  NAND U2935 ( .A(n5820), .B(sreg[1243]), .Z(n2092) );
  AND U2936 ( .A(n2091), .B(n2092), .Z(n5830) );
  NAND U2937 ( .A(n5847), .B(sreg[1246]), .Z(n2093) );
  XOR U2938 ( .A(sreg[1246]), .B(n5847), .Z(n2094) );
  NANDN U2939 ( .A(n5846), .B(n2094), .Z(n2095) );
  NAND U2940 ( .A(n2093), .B(n2095), .Z(n5855) );
  XOR U2941 ( .A(n5871), .B(sreg[1249]), .Z(n2096) );
  NANDN U2942 ( .A(n5872), .B(n2096), .Z(n2097) );
  NAND U2943 ( .A(n5871), .B(sreg[1249]), .Z(n2098) );
  AND U2944 ( .A(n2097), .B(n2098), .Z(n5878) );
  NAND U2945 ( .A(n5895), .B(sreg[1252]), .Z(n2099) );
  XOR U2946 ( .A(sreg[1252]), .B(n5895), .Z(n2100) );
  NANDN U2947 ( .A(n5894), .B(n2100), .Z(n2101) );
  NAND U2948 ( .A(n2099), .B(n2101), .Z(n5903) );
  NAND U2949 ( .A(n5919), .B(sreg[1255]), .Z(n2102) );
  XOR U2950 ( .A(sreg[1255]), .B(n5919), .Z(n2103) );
  NANDN U2951 ( .A(n5920), .B(n2103), .Z(n2104) );
  NAND U2952 ( .A(n2102), .B(n2104), .Z(n5928) );
  NAND U2953 ( .A(n5945), .B(sreg[1258]), .Z(n2105) );
  XOR U2954 ( .A(sreg[1258]), .B(n5945), .Z(n2106) );
  NANDN U2955 ( .A(n5944), .B(n2106), .Z(n2107) );
  NAND U2956 ( .A(n2105), .B(n2107), .Z(n5953) );
  NAND U2957 ( .A(n5971), .B(sreg[1261]), .Z(n2108) );
  XOR U2958 ( .A(sreg[1261]), .B(n5971), .Z(n2109) );
  NAND U2959 ( .A(n2109), .B(n5970), .Z(n2110) );
  NAND U2960 ( .A(n2108), .B(n2110), .Z(n5977) );
  NAND U2961 ( .A(n5994), .B(sreg[1264]), .Z(n2111) );
  XOR U2962 ( .A(sreg[1264]), .B(n5994), .Z(n2112) );
  NANDN U2963 ( .A(n5993), .B(n2112), .Z(n2113) );
  NAND U2964 ( .A(n2111), .B(n2113), .Z(n6002) );
  XOR U2965 ( .A(n6018), .B(sreg[1267]), .Z(n2114) );
  NANDN U2966 ( .A(n6019), .B(n2114), .Z(n2115) );
  NAND U2967 ( .A(n6018), .B(sreg[1267]), .Z(n2116) );
  AND U2968 ( .A(n2115), .B(n2116), .Z(n6025) );
  NAND U2969 ( .A(n6042), .B(sreg[1270]), .Z(n2117) );
  XOR U2970 ( .A(sreg[1270]), .B(n6042), .Z(n2118) );
  NANDN U2971 ( .A(n6041), .B(n2118), .Z(n2119) );
  NAND U2972 ( .A(n2117), .B(n2119), .Z(n6050) );
  XOR U2973 ( .A(n6069), .B(sreg[1273]), .Z(n2120) );
  NANDN U2974 ( .A(n6070), .B(n2120), .Z(n2121) );
  NAND U2975 ( .A(n6069), .B(sreg[1273]), .Z(n2122) );
  AND U2976 ( .A(n2121), .B(n2122), .Z(n6076) );
  NAND U2977 ( .A(n6093), .B(sreg[1276]), .Z(n2123) );
  XOR U2978 ( .A(sreg[1276]), .B(n6093), .Z(n2124) );
  NANDN U2979 ( .A(n6092), .B(n2124), .Z(n2125) );
  NAND U2980 ( .A(n2123), .B(n2125), .Z(n6101) );
  XOR U2981 ( .A(n6117), .B(sreg[1279]), .Z(n2126) );
  NANDN U2982 ( .A(n6118), .B(n2126), .Z(n2127) );
  NAND U2983 ( .A(n6117), .B(sreg[1279]), .Z(n2128) );
  AND U2984 ( .A(n2127), .B(n2128), .Z(n6124) );
  NAND U2985 ( .A(n6139), .B(sreg[1282]), .Z(n2129) );
  XOR U2986 ( .A(sreg[1282]), .B(n6139), .Z(n2130) );
  NAND U2987 ( .A(n2130), .B(n6138), .Z(n2131) );
  NAND U2988 ( .A(n2129), .B(n2131), .Z(n6147) );
  NAND U2989 ( .A(n6165), .B(sreg[1285]), .Z(n2132) );
  XOR U2990 ( .A(sreg[1285]), .B(n6165), .Z(n2133) );
  NAND U2991 ( .A(n2133), .B(n6164), .Z(n2134) );
  NAND U2992 ( .A(n2132), .B(n2134), .Z(n6171) );
  NAND U2993 ( .A(n6189), .B(sreg[1288]), .Z(n2135) );
  XOR U2994 ( .A(sreg[1288]), .B(n6189), .Z(n2136) );
  NANDN U2995 ( .A(n6190), .B(n2136), .Z(n2137) );
  NAND U2996 ( .A(n2135), .B(n2137), .Z(n6198) );
  NAND U2997 ( .A(n6213), .B(sreg[1291]), .Z(n2138) );
  XOR U2998 ( .A(sreg[1291]), .B(n6213), .Z(n2139) );
  NAND U2999 ( .A(n2139), .B(n6212), .Z(n2140) );
  NAND U3000 ( .A(n2138), .B(n2140), .Z(n6219) );
  NAND U3001 ( .A(n6236), .B(sreg[1294]), .Z(n2141) );
  XOR U3002 ( .A(sreg[1294]), .B(n6236), .Z(n2142) );
  NANDN U3003 ( .A(n6235), .B(n2142), .Z(n2143) );
  NAND U3004 ( .A(n2141), .B(n2143), .Z(n6244) );
  NAND U3005 ( .A(n6263), .B(sreg[1297]), .Z(n2144) );
  XOR U3006 ( .A(sreg[1297]), .B(n6263), .Z(n2145) );
  NANDN U3007 ( .A(n6264), .B(n2145), .Z(n2146) );
  NAND U3008 ( .A(n2144), .B(n2146), .Z(n6272) );
  NAND U3009 ( .A(n6289), .B(sreg[1300]), .Z(n2147) );
  XOR U3010 ( .A(sreg[1300]), .B(n6289), .Z(n2148) );
  NANDN U3011 ( .A(n6288), .B(n2148), .Z(n2149) );
  NAND U3012 ( .A(n2147), .B(n2149), .Z(n6297) );
  XOR U3013 ( .A(n6313), .B(sreg[1303]), .Z(n2150) );
  NANDN U3014 ( .A(n6314), .B(n2150), .Z(n2151) );
  NAND U3015 ( .A(n6313), .B(sreg[1303]), .Z(n2152) );
  AND U3016 ( .A(n2151), .B(n2152), .Z(n6320) );
  NAND U3017 ( .A(n6337), .B(sreg[1306]), .Z(n2153) );
  XOR U3018 ( .A(sreg[1306]), .B(n6337), .Z(n2154) );
  NANDN U3019 ( .A(n6336), .B(n2154), .Z(n2155) );
  NAND U3020 ( .A(n2153), .B(n2155), .Z(n6345) );
  XOR U3021 ( .A(n6363), .B(sreg[1309]), .Z(n2156) );
  NANDN U3022 ( .A(n6364), .B(n2156), .Z(n2157) );
  NAND U3023 ( .A(n6363), .B(sreg[1309]), .Z(n2158) );
  AND U3024 ( .A(n2157), .B(n2158), .Z(n6370) );
  NAND U3025 ( .A(n6387), .B(sreg[1312]), .Z(n2159) );
  XOR U3026 ( .A(sreg[1312]), .B(n6387), .Z(n2160) );
  NANDN U3027 ( .A(n6386), .B(n2160), .Z(n2161) );
  NAND U3028 ( .A(n2159), .B(n2161), .Z(n6395) );
  XOR U3029 ( .A(n6413), .B(sreg[1315]), .Z(n2162) );
  NANDN U3030 ( .A(n6414), .B(n2162), .Z(n2163) );
  NAND U3031 ( .A(n6413), .B(sreg[1315]), .Z(n2164) );
  AND U3032 ( .A(n2163), .B(n2164), .Z(n6423) );
  NAND U3033 ( .A(n6440), .B(sreg[1318]), .Z(n2165) );
  XOR U3034 ( .A(sreg[1318]), .B(n6440), .Z(n2166) );
  NANDN U3035 ( .A(n6439), .B(n2166), .Z(n2167) );
  NAND U3036 ( .A(n2165), .B(n2167), .Z(n6448) );
  XOR U3037 ( .A(n6464), .B(sreg[1321]), .Z(n2168) );
  NANDN U3038 ( .A(n6465), .B(n2168), .Z(n2169) );
  NAND U3039 ( .A(n6464), .B(sreg[1321]), .Z(n2170) );
  AND U3040 ( .A(n2169), .B(n2170), .Z(n6471) );
  NAND U3041 ( .A(n6488), .B(sreg[1324]), .Z(n2171) );
  XOR U3042 ( .A(sreg[1324]), .B(n6488), .Z(n2172) );
  NANDN U3043 ( .A(n6487), .B(n2172), .Z(n2173) );
  NAND U3044 ( .A(n2171), .B(n2173), .Z(n6496) );
  XOR U3045 ( .A(n6512), .B(sreg[1327]), .Z(n2174) );
  NANDN U3046 ( .A(n6513), .B(n2174), .Z(n2175) );
  NAND U3047 ( .A(n6512), .B(sreg[1327]), .Z(n2176) );
  AND U3048 ( .A(n2175), .B(n2176), .Z(n6519) );
  NAND U3049 ( .A(n6539), .B(sreg[1330]), .Z(n2177) );
  XOR U3050 ( .A(sreg[1330]), .B(n6539), .Z(n2178) );
  NANDN U3051 ( .A(n6538), .B(n2178), .Z(n2179) );
  NAND U3052 ( .A(n2177), .B(n2179), .Z(n6547) );
  XOR U3053 ( .A(n6563), .B(sreg[1333]), .Z(n2180) );
  NANDN U3054 ( .A(n6564), .B(n2180), .Z(n2181) );
  NAND U3055 ( .A(n6563), .B(sreg[1333]), .Z(n2182) );
  AND U3056 ( .A(n2181), .B(n2182), .Z(n6570) );
  NAND U3057 ( .A(n6587), .B(sreg[1336]), .Z(n2183) );
  XOR U3058 ( .A(sreg[1336]), .B(n6587), .Z(n2184) );
  NANDN U3059 ( .A(n6586), .B(n2184), .Z(n2185) );
  NAND U3060 ( .A(n2183), .B(n2185), .Z(n6595) );
  XOR U3061 ( .A(n6611), .B(sreg[1339]), .Z(n2186) );
  NANDN U3062 ( .A(n6612), .B(n2186), .Z(n2187) );
  NAND U3063 ( .A(n6611), .B(sreg[1339]), .Z(n2188) );
  AND U3064 ( .A(n2187), .B(n2188), .Z(n6618) );
  NAND U3065 ( .A(n6635), .B(sreg[1342]), .Z(n2189) );
  XOR U3066 ( .A(sreg[1342]), .B(n6635), .Z(n2190) );
  NANDN U3067 ( .A(n6634), .B(n2190), .Z(n2191) );
  NAND U3068 ( .A(n2189), .B(n2191), .Z(n6643) );
  XOR U3069 ( .A(n6662), .B(sreg[1345]), .Z(n2192) );
  NANDN U3070 ( .A(n6663), .B(n2192), .Z(n2193) );
  NAND U3071 ( .A(n6662), .B(sreg[1345]), .Z(n2194) );
  AND U3072 ( .A(n2193), .B(n2194), .Z(n6669) );
  NAND U3073 ( .A(n6687), .B(sreg[1348]), .Z(n2195) );
  XOR U3074 ( .A(sreg[1348]), .B(n6687), .Z(n2196) );
  NANDN U3075 ( .A(n6688), .B(n2196), .Z(n2197) );
  NAND U3076 ( .A(n2195), .B(n2197), .Z(n6696) );
  NAND U3077 ( .A(n6711), .B(sreg[1351]), .Z(n2198) );
  XOR U3078 ( .A(sreg[1351]), .B(n6711), .Z(n2199) );
  NAND U3079 ( .A(n2199), .B(n6710), .Z(n2200) );
  NAND U3080 ( .A(n2198), .B(n2200), .Z(n6717) );
  NAND U3081 ( .A(n6734), .B(sreg[1354]), .Z(n2201) );
  XOR U3082 ( .A(sreg[1354]), .B(n6734), .Z(n2202) );
  NANDN U3083 ( .A(n6733), .B(n2202), .Z(n2203) );
  NAND U3084 ( .A(n2201), .B(n2203), .Z(n6740) );
  XOR U3085 ( .A(n6759), .B(sreg[1357]), .Z(n2204) );
  NANDN U3086 ( .A(n6760), .B(n2204), .Z(n2205) );
  NAND U3087 ( .A(n6759), .B(sreg[1357]), .Z(n2206) );
  AND U3088 ( .A(n2205), .B(n2206), .Z(n6766) );
  NAND U3089 ( .A(n6783), .B(sreg[1360]), .Z(n2207) );
  XOR U3090 ( .A(sreg[1360]), .B(n6783), .Z(n2208) );
  NANDN U3091 ( .A(n6782), .B(n2208), .Z(n2209) );
  NAND U3092 ( .A(n2207), .B(n2209), .Z(n6791) );
  XOR U3093 ( .A(n6809), .B(sreg[1363]), .Z(n2210) );
  NANDN U3094 ( .A(n6810), .B(n2210), .Z(n2211) );
  NAND U3095 ( .A(n6809), .B(sreg[1363]), .Z(n2212) );
  AND U3096 ( .A(n2211), .B(n2212), .Z(n6816) );
  NAND U3097 ( .A(n6834), .B(sreg[1366]), .Z(n2213) );
  XOR U3098 ( .A(sreg[1366]), .B(n6834), .Z(n2214) );
  NANDN U3099 ( .A(n6835), .B(n2214), .Z(n2215) );
  NAND U3100 ( .A(n2213), .B(n2215), .Z(n6843) );
  XOR U3101 ( .A(n6859), .B(sreg[1369]), .Z(n2216) );
  NANDN U3102 ( .A(n6860), .B(n2216), .Z(n2217) );
  NAND U3103 ( .A(n6859), .B(sreg[1369]), .Z(n2218) );
  AND U3104 ( .A(n2217), .B(n2218), .Z(n6866) );
  NAND U3105 ( .A(n6884), .B(sreg[1372]), .Z(n2219) );
  XOR U3106 ( .A(sreg[1372]), .B(n6884), .Z(n2220) );
  NANDN U3107 ( .A(n6885), .B(n2220), .Z(n2221) );
  NAND U3108 ( .A(n2219), .B(n2221), .Z(n6893) );
  XOR U3109 ( .A(n6909), .B(sreg[1375]), .Z(n2222) );
  NANDN U3110 ( .A(n6910), .B(n2222), .Z(n2223) );
  NAND U3111 ( .A(n6909), .B(sreg[1375]), .Z(n2224) );
  AND U3112 ( .A(n2223), .B(n2224), .Z(n6919) );
  NAND U3113 ( .A(n6936), .B(sreg[1378]), .Z(n2225) );
  XOR U3114 ( .A(sreg[1378]), .B(n6936), .Z(n2226) );
  NANDN U3115 ( .A(n6935), .B(n2226), .Z(n2227) );
  NAND U3116 ( .A(n2225), .B(n2227), .Z(n6944) );
  XOR U3117 ( .A(n6960), .B(sreg[1381]), .Z(n2228) );
  NANDN U3118 ( .A(n6961), .B(n2228), .Z(n2229) );
  NAND U3119 ( .A(n6960), .B(sreg[1381]), .Z(n2230) );
  AND U3120 ( .A(n2229), .B(n2230), .Z(n6967) );
  NAND U3121 ( .A(n6982), .B(sreg[1384]), .Z(n2231) );
  XOR U3122 ( .A(sreg[1384]), .B(n6982), .Z(n2232) );
  NAND U3123 ( .A(n2232), .B(n6981), .Z(n2233) );
  NAND U3124 ( .A(n2231), .B(n2233), .Z(n6990) );
  NAND U3125 ( .A(n7008), .B(sreg[1387]), .Z(n2234) );
  XOR U3126 ( .A(sreg[1387]), .B(n7008), .Z(n2235) );
  NAND U3127 ( .A(n2235), .B(n7007), .Z(n2236) );
  NAND U3128 ( .A(n2234), .B(n2236), .Z(n7014) );
  NAND U3129 ( .A(n7031), .B(sreg[1390]), .Z(n2237) );
  XOR U3130 ( .A(sreg[1390]), .B(n7031), .Z(n2238) );
  NANDN U3131 ( .A(n7030), .B(n2238), .Z(n2239) );
  NAND U3132 ( .A(n2237), .B(n2239), .Z(n7039) );
  XOR U3133 ( .A(n7055), .B(sreg[1393]), .Z(n2240) );
  NANDN U3134 ( .A(n7056), .B(n2240), .Z(n2241) );
  NAND U3135 ( .A(n7055), .B(sreg[1393]), .Z(n2242) );
  AND U3136 ( .A(n2241), .B(n2242), .Z(n7062) );
  NAND U3137 ( .A(n7077), .B(sreg[1396]), .Z(n2243) );
  XOR U3138 ( .A(sreg[1396]), .B(n7077), .Z(n2244) );
  NAND U3139 ( .A(n2244), .B(n7076), .Z(n2245) );
  NAND U3140 ( .A(n2243), .B(n2245), .Z(n7085) );
  XOR U3141 ( .A(n7104), .B(sreg[1399]), .Z(n2246) );
  NANDN U3142 ( .A(n7105), .B(n2246), .Z(n2247) );
  NAND U3143 ( .A(n7104), .B(sreg[1399]), .Z(n2248) );
  AND U3144 ( .A(n2247), .B(n2248), .Z(n7111) );
  NAND U3145 ( .A(n7126), .B(sreg[1402]), .Z(n2249) );
  XOR U3146 ( .A(sreg[1402]), .B(n7126), .Z(n2250) );
  NAND U3147 ( .A(n2250), .B(n7125), .Z(n2251) );
  NAND U3148 ( .A(n2249), .B(n2251), .Z(n7134) );
  XOR U3149 ( .A(n7150), .B(sreg[1405]), .Z(n2252) );
  NANDN U3150 ( .A(n7151), .B(n2252), .Z(n2253) );
  NAND U3151 ( .A(n7150), .B(sreg[1405]), .Z(n2254) );
  AND U3152 ( .A(n2253), .B(n2254), .Z(n7157) );
  NAND U3153 ( .A(n7174), .B(sreg[1408]), .Z(n2255) );
  XOR U3154 ( .A(sreg[1408]), .B(n7174), .Z(n2256) );
  NANDN U3155 ( .A(n7173), .B(n2256), .Z(n2257) );
  NAND U3156 ( .A(n2255), .B(n2257), .Z(n7182) );
  XOR U3157 ( .A(n7201), .B(sreg[1411]), .Z(n2258) );
  NANDN U3158 ( .A(n7202), .B(n2258), .Z(n2259) );
  NAND U3159 ( .A(n7201), .B(sreg[1411]), .Z(n2260) );
  AND U3160 ( .A(n2259), .B(n2260), .Z(n7208) );
  NAND U3161 ( .A(n7225), .B(sreg[1414]), .Z(n2261) );
  XOR U3162 ( .A(sreg[1414]), .B(n7225), .Z(n2262) );
  NANDN U3163 ( .A(n7224), .B(n2262), .Z(n2263) );
  NAND U3164 ( .A(n2261), .B(n2263), .Z(n7233) );
  XOR U3165 ( .A(n7249), .B(sreg[1417]), .Z(n2264) );
  NANDN U3166 ( .A(n7250), .B(n2264), .Z(n2265) );
  NAND U3167 ( .A(n7249), .B(sreg[1417]), .Z(n2266) );
  AND U3168 ( .A(n2265), .B(n2266), .Z(n7256) );
  NAND U3169 ( .A(n7273), .B(sreg[1420]), .Z(n2267) );
  XOR U3170 ( .A(sreg[1420]), .B(n7273), .Z(n2268) );
  NANDN U3171 ( .A(n7272), .B(n2268), .Z(n2269) );
  NAND U3172 ( .A(n2267), .B(n2269), .Z(n7281) );
  XOR U3173 ( .A(n7297), .B(sreg[1423]), .Z(n2270) );
  NANDN U3174 ( .A(n7298), .B(n2270), .Z(n2271) );
  NAND U3175 ( .A(n7297), .B(sreg[1423]), .Z(n2272) );
  AND U3176 ( .A(n2271), .B(n2272), .Z(n7307) );
  NAND U3177 ( .A(n7324), .B(sreg[1426]), .Z(n2273) );
  XOR U3178 ( .A(sreg[1426]), .B(n7324), .Z(n2274) );
  NANDN U3179 ( .A(n7323), .B(n2274), .Z(n2275) );
  NAND U3180 ( .A(n2273), .B(n2275), .Z(n7332) );
  XOR U3181 ( .A(n7350), .B(sreg[1429]), .Z(n2276) );
  NANDN U3182 ( .A(n7351), .B(n2276), .Z(n2277) );
  NAND U3183 ( .A(n7350), .B(sreg[1429]), .Z(n2278) );
  AND U3184 ( .A(n2277), .B(n2278), .Z(n7357) );
  NAND U3185 ( .A(n7374), .B(sreg[1432]), .Z(n2279) );
  XOR U3186 ( .A(sreg[1432]), .B(n7374), .Z(n2280) );
  NANDN U3187 ( .A(n7373), .B(n2280), .Z(n2281) );
  NAND U3188 ( .A(n2279), .B(n2281), .Z(n7380) );
  XOR U3189 ( .A(n7398), .B(sreg[1435]), .Z(n2282) );
  NANDN U3190 ( .A(n7399), .B(n2282), .Z(n2283) );
  NAND U3191 ( .A(n7398), .B(sreg[1435]), .Z(n2284) );
  AND U3192 ( .A(n2283), .B(n2284), .Z(n7405) );
  NAND U3193 ( .A(n7422), .B(sreg[1438]), .Z(n2285) );
  XOR U3194 ( .A(sreg[1438]), .B(n7422), .Z(n2286) );
  NANDN U3195 ( .A(n7421), .B(n2286), .Z(n2287) );
  NAND U3196 ( .A(n2285), .B(n2287), .Z(n7430) );
  XOR U3197 ( .A(n7449), .B(sreg[1441]), .Z(n2288) );
  NANDN U3198 ( .A(n7450), .B(n2288), .Z(n2289) );
  NAND U3199 ( .A(n7449), .B(sreg[1441]), .Z(n2290) );
  AND U3200 ( .A(n2289), .B(n2290), .Z(n7456) );
  NAND U3201 ( .A(n7472), .B(sreg[1444]), .Z(n2291) );
  XOR U3202 ( .A(sreg[1444]), .B(n7472), .Z(n2292) );
  NANDN U3203 ( .A(n7473), .B(n2292), .Z(n2293) );
  NAND U3204 ( .A(n2291), .B(n2293), .Z(n7481) );
  NAND U3205 ( .A(n7496), .B(sreg[1447]), .Z(n2294) );
  XOR U3206 ( .A(sreg[1447]), .B(n7496), .Z(n2295) );
  NAND U3207 ( .A(n2295), .B(n7495), .Z(n2296) );
  NAND U3208 ( .A(n2294), .B(n2296), .Z(n7502) );
  NAND U3209 ( .A(n7518), .B(sreg[1450]), .Z(n2297) );
  XOR U3210 ( .A(sreg[1450]), .B(n7518), .Z(n2298) );
  NANDN U3211 ( .A(n7519), .B(n2298), .Z(n2299) );
  NAND U3212 ( .A(n2297), .B(n2299), .Z(n7527) );
  XOR U3213 ( .A(n7546), .B(sreg[1453]), .Z(n2300) );
  NANDN U3214 ( .A(n7547), .B(n2300), .Z(n2301) );
  NAND U3215 ( .A(n7546), .B(sreg[1453]), .Z(n2302) );
  AND U3216 ( .A(n2301), .B(n2302), .Z(n7553) );
  NAND U3217 ( .A(n7571), .B(sreg[1456]), .Z(n2303) );
  XOR U3218 ( .A(sreg[1456]), .B(n7571), .Z(n2304) );
  NANDN U3219 ( .A(n7572), .B(n2304), .Z(n2305) );
  NAND U3220 ( .A(n2303), .B(n2305), .Z(n7580) );
  NAND U3221 ( .A(n7595), .B(sreg[1459]), .Z(n2306) );
  XOR U3222 ( .A(sreg[1459]), .B(n7595), .Z(n2307) );
  NAND U3223 ( .A(n2307), .B(n7594), .Z(n2308) );
  NAND U3224 ( .A(n2306), .B(n2308), .Z(n7601) );
  NAND U3225 ( .A(n7618), .B(sreg[1462]), .Z(n2309) );
  XOR U3226 ( .A(sreg[1462]), .B(n7618), .Z(n2310) );
  NANDN U3227 ( .A(n7617), .B(n2310), .Z(n2311) );
  NAND U3228 ( .A(n2309), .B(n2311), .Z(n7626) );
  XOR U3229 ( .A(n7642), .B(sreg[1465]), .Z(n2312) );
  NANDN U3230 ( .A(n7643), .B(n2312), .Z(n2313) );
  NAND U3231 ( .A(n7642), .B(sreg[1465]), .Z(n2314) );
  AND U3232 ( .A(n2313), .B(n2314), .Z(n7652) );
  NAND U3233 ( .A(n7669), .B(sreg[1468]), .Z(n2315) );
  XOR U3234 ( .A(sreg[1468]), .B(n7669), .Z(n2316) );
  NANDN U3235 ( .A(n7668), .B(n2316), .Z(n2317) );
  NAND U3236 ( .A(n2315), .B(n2317), .Z(n7677) );
  XOR U3237 ( .A(n7693), .B(sreg[1471]), .Z(n2318) );
  NANDN U3238 ( .A(n7694), .B(n2318), .Z(n2319) );
  NAND U3239 ( .A(n7693), .B(sreg[1471]), .Z(n2320) );
  AND U3240 ( .A(n2319), .B(n2320), .Z(n7700) );
  NAND U3241 ( .A(n7717), .B(sreg[1474]), .Z(n2321) );
  XOR U3242 ( .A(sreg[1474]), .B(n7717), .Z(n2322) );
  NANDN U3243 ( .A(n7716), .B(n2322), .Z(n2323) );
  NAND U3244 ( .A(n2321), .B(n2323), .Z(n7725) );
  XOR U3245 ( .A(n7743), .B(sreg[1477]), .Z(n2324) );
  NANDN U3246 ( .A(n7744), .B(n2324), .Z(n2325) );
  NAND U3247 ( .A(n7743), .B(sreg[1477]), .Z(n2326) );
  AND U3248 ( .A(n2325), .B(n2326), .Z(n7750) );
  NAND U3249 ( .A(n7767), .B(sreg[1480]), .Z(n2327) );
  XOR U3250 ( .A(sreg[1480]), .B(n7767), .Z(n2328) );
  NANDN U3251 ( .A(n7766), .B(n2328), .Z(n2329) );
  NAND U3252 ( .A(n2327), .B(n2329), .Z(n7776) );
  NAND U3253 ( .A(n7793), .B(sreg[1483]), .Z(n2330) );
  XOR U3254 ( .A(sreg[1483]), .B(n7793), .Z(n2331) );
  NANDN U3255 ( .A(n7792), .B(n2331), .Z(n2332) );
  NAND U3256 ( .A(n2330), .B(n2332), .Z(n7799) );
  NAND U3257 ( .A(n7814), .B(sreg[1486]), .Z(n2333) );
  XOR U3258 ( .A(sreg[1486]), .B(n7814), .Z(n2334) );
  NAND U3259 ( .A(n2334), .B(n7813), .Z(n2335) );
  NAND U3260 ( .A(n2333), .B(n2335), .Z(n7822) );
  XOR U3261 ( .A(n7838), .B(sreg[1489]), .Z(n2336) );
  NANDN U3262 ( .A(n7839), .B(n2336), .Z(n2337) );
  NAND U3263 ( .A(n7838), .B(sreg[1489]), .Z(n2338) );
  AND U3264 ( .A(n2337), .B(n2338), .Z(n7845) );
  NAND U3265 ( .A(n7865), .B(sreg[1492]), .Z(n2339) );
  XOR U3266 ( .A(sreg[1492]), .B(n7865), .Z(n2340) );
  NANDN U3267 ( .A(n7864), .B(n2340), .Z(n2341) );
  NAND U3268 ( .A(n2339), .B(n2341), .Z(n7873) );
  XOR U3269 ( .A(n7889), .B(sreg[1495]), .Z(n2342) );
  NANDN U3270 ( .A(n7890), .B(n2342), .Z(n2343) );
  NAND U3271 ( .A(n7889), .B(sreg[1495]), .Z(n2344) );
  AND U3272 ( .A(n2343), .B(n2344), .Z(n7896) );
  NAND U3273 ( .A(n7913), .B(sreg[1498]), .Z(n2345) );
  XOR U3274 ( .A(sreg[1498]), .B(n7913), .Z(n2346) );
  NANDN U3275 ( .A(n7912), .B(n2346), .Z(n2347) );
  NAND U3276 ( .A(n2345), .B(n2347), .Z(n7921) );
  XOR U3277 ( .A(n7937), .B(sreg[1501]), .Z(n2348) );
  NANDN U3278 ( .A(n7938), .B(n2348), .Z(n2349) );
  NAND U3279 ( .A(n7937), .B(sreg[1501]), .Z(n2350) );
  AND U3280 ( .A(n2349), .B(n2350), .Z(n7944) );
  NAND U3281 ( .A(n7961), .B(sreg[1504]), .Z(n2351) );
  XOR U3282 ( .A(sreg[1504]), .B(n7961), .Z(n2352) );
  NANDN U3283 ( .A(n7960), .B(n2352), .Z(n2353) );
  NAND U3284 ( .A(n2351), .B(n2353), .Z(n7969) );
  NAND U3285 ( .A(n7987), .B(sreg[1507]), .Z(n2354) );
  XOR U3286 ( .A(sreg[1507]), .B(n7987), .Z(n2355) );
  NAND U3287 ( .A(n2355), .B(n7986), .Z(n2356) );
  NAND U3288 ( .A(n2354), .B(n2356), .Z(n7993) );
  NAND U3289 ( .A(n8010), .B(sreg[1510]), .Z(n2357) );
  XOR U3290 ( .A(sreg[1510]), .B(n8010), .Z(n2358) );
  NANDN U3291 ( .A(n8009), .B(n2358), .Z(n2359) );
  NAND U3292 ( .A(n2357), .B(n2359), .Z(n8016) );
  NAND U3293 ( .A(n8033), .B(sreg[1513]), .Z(n2360) );
  XOR U3294 ( .A(sreg[1513]), .B(n8033), .Z(n2361) );
  NANDN U3295 ( .A(n8032), .B(n2361), .Z(n2362) );
  NAND U3296 ( .A(n2360), .B(n2362), .Z(n8041) );
  NAND U3297 ( .A(n8059), .B(sreg[1516]), .Z(n2363) );
  XOR U3298 ( .A(sreg[1516]), .B(n8059), .Z(n2364) );
  NAND U3299 ( .A(n2364), .B(n8058), .Z(n2365) );
  NAND U3300 ( .A(n2363), .B(n2365), .Z(n8067) );
  XOR U3301 ( .A(n8085), .B(sreg[1519]), .Z(n2366) );
  NANDN U3302 ( .A(n8086), .B(n2366), .Z(n2367) );
  NAND U3303 ( .A(n8085), .B(sreg[1519]), .Z(n2368) );
  AND U3304 ( .A(n2367), .B(n2368), .Z(n8092) );
  NAND U3305 ( .A(n8109), .B(sreg[1522]), .Z(n2369) );
  XOR U3306 ( .A(sreg[1522]), .B(n8109), .Z(n2370) );
  NANDN U3307 ( .A(n8108), .B(n2370), .Z(n2371) );
  NAND U3308 ( .A(n2369), .B(n2371), .Z(n8117) );
  XOR U3309 ( .A(n8133), .B(sreg[1525]), .Z(n2372) );
  NANDN U3310 ( .A(n8134), .B(n2372), .Z(n2373) );
  NAND U3311 ( .A(n8133), .B(sreg[1525]), .Z(n2374) );
  AND U3312 ( .A(n2373), .B(n2374), .Z(n8140) );
  NAND U3313 ( .A(n8157), .B(sreg[1528]), .Z(n2375) );
  XOR U3314 ( .A(sreg[1528]), .B(n8157), .Z(n2376) );
  NANDN U3315 ( .A(n8156), .B(n2376), .Z(n2377) );
  NAND U3316 ( .A(n2375), .B(n2377), .Z(n8165) );
  XOR U3317 ( .A(n8181), .B(sreg[1531]), .Z(n2378) );
  NANDN U3318 ( .A(n8182), .B(n2378), .Z(n2379) );
  NAND U3319 ( .A(n8181), .B(sreg[1531]), .Z(n2380) );
  AND U3320 ( .A(n2379), .B(n2380), .Z(n8191) );
  NAND U3321 ( .A(n8208), .B(sreg[1534]), .Z(n2381) );
  XOR U3322 ( .A(sreg[1534]), .B(n8208), .Z(n2382) );
  NANDN U3323 ( .A(n8207), .B(n2382), .Z(n2383) );
  NAND U3324 ( .A(n2381), .B(n2383), .Z(n8216) );
  XOR U3325 ( .A(n8232), .B(sreg[1537]), .Z(n2384) );
  NANDN U3326 ( .A(n8233), .B(n2384), .Z(n2385) );
  NAND U3327 ( .A(n8232), .B(sreg[1537]), .Z(n2386) );
  AND U3328 ( .A(n2385), .B(n2386), .Z(n8239) );
  NAND U3329 ( .A(n8256), .B(sreg[1540]), .Z(n2387) );
  XOR U3330 ( .A(sreg[1540]), .B(n8256), .Z(n2388) );
  NANDN U3331 ( .A(n8255), .B(n2388), .Z(n2389) );
  NAND U3332 ( .A(n2387), .B(n2389), .Z(n8262) );
  XOR U3333 ( .A(n8278), .B(sreg[1543]), .Z(n2390) );
  NANDN U3334 ( .A(n8279), .B(n2390), .Z(n2391) );
  NAND U3335 ( .A(n8278), .B(sreg[1543]), .Z(n2392) );
  AND U3336 ( .A(n2391), .B(n2392), .Z(n8288) );
  NAND U3337 ( .A(n8305), .B(sreg[1546]), .Z(n2393) );
  XOR U3338 ( .A(sreg[1546]), .B(n8305), .Z(n2394) );
  NANDN U3339 ( .A(n8304), .B(n2394), .Z(n2395) );
  NAND U3340 ( .A(n2393), .B(n2395), .Z(n8313) );
  XOR U3341 ( .A(n8329), .B(sreg[1549]), .Z(n2396) );
  NANDN U3342 ( .A(n8330), .B(n2396), .Z(n2397) );
  NAND U3343 ( .A(n8329), .B(sreg[1549]), .Z(n2398) );
  AND U3344 ( .A(n2397), .B(n2398), .Z(n8336) );
  NAND U3345 ( .A(n8353), .B(sreg[1552]), .Z(n2399) );
  XOR U3346 ( .A(sreg[1552]), .B(n8353), .Z(n2400) );
  NANDN U3347 ( .A(n8352), .B(n2400), .Z(n2401) );
  NAND U3348 ( .A(n2399), .B(n2401), .Z(n8361) );
  XOR U3349 ( .A(n8377), .B(sreg[1555]), .Z(n2402) );
  NANDN U3350 ( .A(n8378), .B(n2402), .Z(n2403) );
  NAND U3351 ( .A(n8377), .B(sreg[1555]), .Z(n2404) );
  AND U3352 ( .A(n2403), .B(n2404), .Z(n8384) );
  NAND U3353 ( .A(n8404), .B(sreg[1558]), .Z(n2405) );
  XOR U3354 ( .A(sreg[1558]), .B(n8404), .Z(n2406) );
  NANDN U3355 ( .A(n8403), .B(n2406), .Z(n2407) );
  NAND U3356 ( .A(n2405), .B(n2407), .Z(n8412) );
  NAND U3357 ( .A(n8427), .B(sreg[1561]), .Z(n2408) );
  XOR U3358 ( .A(sreg[1561]), .B(n8427), .Z(n2409) );
  NAND U3359 ( .A(n2409), .B(n8426), .Z(n2410) );
  NAND U3360 ( .A(n2408), .B(n2410), .Z(n8433) );
  NAND U3361 ( .A(n8450), .B(sreg[1564]), .Z(n2411) );
  XOR U3362 ( .A(sreg[1564]), .B(n8450), .Z(n2412) );
  NANDN U3363 ( .A(n8449), .B(n2412), .Z(n2413) );
  NAND U3364 ( .A(n2411), .B(n2413), .Z(n8458) );
  XOR U3365 ( .A(n8474), .B(sreg[1567]), .Z(n2414) );
  NANDN U3366 ( .A(n8475), .B(n2414), .Z(n2415) );
  NAND U3367 ( .A(n8474), .B(sreg[1567]), .Z(n2416) );
  AND U3368 ( .A(n2415), .B(n2416), .Z(n8481) );
  NAND U3369 ( .A(n8501), .B(sreg[1570]), .Z(n2417) );
  XOR U3370 ( .A(sreg[1570]), .B(n8501), .Z(n2418) );
  NANDN U3371 ( .A(n8500), .B(n2418), .Z(n2419) );
  NAND U3372 ( .A(n2417), .B(n2419), .Z(n8509) );
  NAND U3373 ( .A(n8527), .B(sreg[1573]), .Z(n2420) );
  XOR U3374 ( .A(sreg[1573]), .B(n8527), .Z(n2421) );
  NANDN U3375 ( .A(n8528), .B(n2421), .Z(n2422) );
  NAND U3376 ( .A(n2420), .B(n2422), .Z(n8536) );
  NAND U3377 ( .A(n8553), .B(sreg[1576]), .Z(n2423) );
  XOR U3378 ( .A(sreg[1576]), .B(n8553), .Z(n2424) );
  NANDN U3379 ( .A(n8552), .B(n2424), .Z(n2425) );
  NAND U3380 ( .A(n2423), .B(n2425), .Z(n8561) );
  XOR U3381 ( .A(n8579), .B(sreg[1579]), .Z(n2426) );
  NANDN U3382 ( .A(n8580), .B(n2426), .Z(n2427) );
  NAND U3383 ( .A(n8579), .B(sreg[1579]), .Z(n2428) );
  AND U3384 ( .A(n2427), .B(n2428), .Z(n8586) );
  NAND U3385 ( .A(n8603), .B(sreg[1582]), .Z(n2429) );
  XOR U3386 ( .A(sreg[1582]), .B(n8603), .Z(n2430) );
  NANDN U3387 ( .A(n8602), .B(n2430), .Z(n2431) );
  NAND U3388 ( .A(n2429), .B(n2431), .Z(n8611) );
  XOR U3389 ( .A(n8627), .B(sreg[1585]), .Z(n2432) );
  NANDN U3390 ( .A(n8628), .B(n2432), .Z(n2433) );
  NAND U3391 ( .A(n8627), .B(sreg[1585]), .Z(n2434) );
  AND U3392 ( .A(n2433), .B(n2434), .Z(n8634) );
  NAND U3393 ( .A(n8652), .B(sreg[1588]), .Z(n2435) );
  XOR U3394 ( .A(sreg[1588]), .B(n8652), .Z(n2436) );
  NAND U3395 ( .A(n2436), .B(n8651), .Z(n2437) );
  NAND U3396 ( .A(n2435), .B(n2437), .Z(n8660) );
  XOR U3397 ( .A(n8676), .B(sreg[1591]), .Z(n2438) );
  NANDN U3398 ( .A(n8677), .B(n2438), .Z(n2439) );
  NAND U3399 ( .A(n8676), .B(sreg[1591]), .Z(n2440) );
  AND U3400 ( .A(n2439), .B(n2440), .Z(n8683) );
  NAND U3401 ( .A(n8700), .B(sreg[1594]), .Z(n2441) );
  XOR U3402 ( .A(sreg[1594]), .B(n8700), .Z(n2442) );
  NANDN U3403 ( .A(n8699), .B(n2442), .Z(n2443) );
  NAND U3404 ( .A(n2441), .B(n2443), .Z(n8708) );
  XOR U3405 ( .A(n8724), .B(sreg[1597]), .Z(n2444) );
  NANDN U3406 ( .A(n8725), .B(n2444), .Z(n2445) );
  NAND U3407 ( .A(n8724), .B(sreg[1597]), .Z(n2446) );
  AND U3408 ( .A(n2445), .B(n2446), .Z(n8731) );
  NAND U3409 ( .A(n8748), .B(sreg[1600]), .Z(n2447) );
  XOR U3410 ( .A(sreg[1600]), .B(n8748), .Z(n2448) );
  NANDN U3411 ( .A(n8747), .B(n2448), .Z(n2449) );
  NAND U3412 ( .A(n2447), .B(n2449), .Z(n8756) );
  XOR U3413 ( .A(n8775), .B(sreg[1603]), .Z(n2450) );
  NANDN U3414 ( .A(n8776), .B(n2450), .Z(n2451) );
  NAND U3415 ( .A(n8775), .B(sreg[1603]), .Z(n2452) );
  AND U3416 ( .A(n2451), .B(n2452), .Z(n8782) );
  NAND U3417 ( .A(n8799), .B(sreg[1606]), .Z(n2453) );
  XOR U3418 ( .A(sreg[1606]), .B(n8799), .Z(n2454) );
  NANDN U3419 ( .A(n8798), .B(n2454), .Z(n2455) );
  NAND U3420 ( .A(n2453), .B(n2455), .Z(n8807) );
  NAND U3421 ( .A(n8822), .B(sreg[1609]), .Z(n2456) );
  XOR U3422 ( .A(sreg[1609]), .B(n8822), .Z(n2457) );
  NAND U3423 ( .A(n2457), .B(n8821), .Z(n2458) );
  NAND U3424 ( .A(n2456), .B(n2458), .Z(n8830) );
  NAND U3425 ( .A(n8847), .B(sreg[1612]), .Z(n2459) );
  XOR U3426 ( .A(sreg[1612]), .B(n8847), .Z(n2460) );
  NANDN U3427 ( .A(n8846), .B(n2460), .Z(n2461) );
  NAND U3428 ( .A(n2459), .B(n2461), .Z(n8855) );
  XOR U3429 ( .A(n8871), .B(sreg[1615]), .Z(n2462) );
  NANDN U3430 ( .A(n8872), .B(n2462), .Z(n2463) );
  NAND U3431 ( .A(n8871), .B(sreg[1615]), .Z(n2464) );
  AND U3432 ( .A(n2463), .B(n2464), .Z(n8881) );
  NAND U3433 ( .A(n8899), .B(sreg[1618]), .Z(n2465) );
  XOR U3434 ( .A(sreg[1618]), .B(n8899), .Z(n2466) );
  NANDN U3435 ( .A(n8900), .B(n2466), .Z(n2467) );
  NAND U3436 ( .A(n2465), .B(n2467), .Z(n8908) );
  XOR U3437 ( .A(n8924), .B(sreg[1621]), .Z(n2468) );
  NANDN U3438 ( .A(n8925), .B(n2468), .Z(n2469) );
  NAND U3439 ( .A(n8924), .B(sreg[1621]), .Z(n2470) );
  AND U3440 ( .A(n2469), .B(n2470), .Z(n8931) );
  NAND U3441 ( .A(n8948), .B(sreg[1624]), .Z(n2471) );
  XOR U3442 ( .A(sreg[1624]), .B(n8948), .Z(n2472) );
  NANDN U3443 ( .A(n8947), .B(n2472), .Z(n2473) );
  NAND U3444 ( .A(n2471), .B(n2473), .Z(n8954) );
  NAND U3445 ( .A(n8970), .B(sreg[1627]), .Z(n2474) );
  XOR U3446 ( .A(sreg[1627]), .B(n8970), .Z(n2475) );
  NANDN U3447 ( .A(n8971), .B(n2475), .Z(n2476) );
  NAND U3448 ( .A(n2474), .B(n2476), .Z(n8979) );
  NAND U3449 ( .A(n8996), .B(sreg[1630]), .Z(n2477) );
  XOR U3450 ( .A(sreg[1630]), .B(n8996), .Z(n2478) );
  NANDN U3451 ( .A(n8995), .B(n2478), .Z(n2479) );
  NAND U3452 ( .A(n2477), .B(n2479), .Z(n9004) );
  XOR U3453 ( .A(n9022), .B(sreg[1633]), .Z(n2480) );
  NANDN U3454 ( .A(n9023), .B(n2480), .Z(n2481) );
  NAND U3455 ( .A(n9022), .B(sreg[1633]), .Z(n2482) );
  AND U3456 ( .A(n2481), .B(n2482), .Z(n9032) );
  NAND U3457 ( .A(n9049), .B(sreg[1636]), .Z(n2483) );
  XOR U3458 ( .A(sreg[1636]), .B(n9049), .Z(n2484) );
  NANDN U3459 ( .A(n9048), .B(n2484), .Z(n2485) );
  NAND U3460 ( .A(n2483), .B(n2485), .Z(n9057) );
  XOR U3461 ( .A(n9075), .B(sreg[1639]), .Z(n2486) );
  NANDN U3462 ( .A(n9076), .B(n2486), .Z(n2487) );
  NAND U3463 ( .A(n9075), .B(sreg[1639]), .Z(n2488) );
  AND U3464 ( .A(n2487), .B(n2488), .Z(n9082) );
  NAND U3465 ( .A(n9099), .B(sreg[1642]), .Z(n2489) );
  XOR U3466 ( .A(sreg[1642]), .B(n9099), .Z(n2490) );
  NANDN U3467 ( .A(n9098), .B(n2490), .Z(n2491) );
  NAND U3468 ( .A(n2489), .B(n2491), .Z(n9107) );
  NAND U3469 ( .A(n9122), .B(sreg[1645]), .Z(n2492) );
  XOR U3470 ( .A(sreg[1645]), .B(n9122), .Z(n2493) );
  NAND U3471 ( .A(n2493), .B(n9121), .Z(n2494) );
  NAND U3472 ( .A(n2492), .B(n2494), .Z(n9128) );
  NAND U3473 ( .A(n9148), .B(sreg[1648]), .Z(n2495) );
  XOR U3474 ( .A(sreg[1648]), .B(n9148), .Z(n2496) );
  NANDN U3475 ( .A(n9147), .B(n2496), .Z(n2497) );
  NAND U3476 ( .A(n2495), .B(n2497), .Z(n9156) );
  XOR U3477 ( .A(n9172), .B(sreg[1651]), .Z(n2498) );
  NANDN U3478 ( .A(n9173), .B(n2498), .Z(n2499) );
  NAND U3479 ( .A(n9172), .B(sreg[1651]), .Z(n2500) );
  AND U3480 ( .A(n2499), .B(n2500), .Z(n9179) );
  NAND U3481 ( .A(n9194), .B(sreg[1654]), .Z(n2501) );
  XOR U3482 ( .A(sreg[1654]), .B(n9194), .Z(n2502) );
  NAND U3483 ( .A(n2502), .B(n9193), .Z(n2503) );
  NAND U3484 ( .A(n2501), .B(n2503), .Z(n9202) );
  NAND U3485 ( .A(n9217), .B(sreg[1657]), .Z(n2504) );
  XOR U3486 ( .A(sreg[1657]), .B(n9217), .Z(n2505) );
  NAND U3487 ( .A(n2505), .B(n9216), .Z(n2506) );
  NAND U3488 ( .A(n2504), .B(n2506), .Z(n9226) );
  NAND U3489 ( .A(n9243), .B(sreg[1660]), .Z(n2507) );
  XOR U3490 ( .A(sreg[1660]), .B(n9243), .Z(n2508) );
  NANDN U3491 ( .A(n9242), .B(n2508), .Z(n2509) );
  NAND U3492 ( .A(n2507), .B(n2509), .Z(n9251) );
  NAND U3493 ( .A(n9267), .B(sreg[1663]), .Z(n2510) );
  XOR U3494 ( .A(sreg[1663]), .B(n9267), .Z(n2511) );
  NANDN U3495 ( .A(n9268), .B(n2511), .Z(n2512) );
  NAND U3496 ( .A(n2510), .B(n2512), .Z(n9276) );
  NAND U3497 ( .A(n9293), .B(sreg[1666]), .Z(n2513) );
  XOR U3498 ( .A(sreg[1666]), .B(n9293), .Z(n2514) );
  NANDN U3499 ( .A(n9292), .B(n2514), .Z(n2515) );
  NAND U3500 ( .A(n2513), .B(n2515), .Z(n9301) );
  XOR U3501 ( .A(n9317), .B(sreg[1669]), .Z(n2516) );
  NANDN U3502 ( .A(n9318), .B(n2516), .Z(n2517) );
  NAND U3503 ( .A(n9317), .B(sreg[1669]), .Z(n2518) );
  AND U3504 ( .A(n2517), .B(n2518), .Z(n9324) );
  NAND U3505 ( .A(n9342), .B(sreg[1672]), .Z(n2519) );
  XOR U3506 ( .A(sreg[1672]), .B(n9342), .Z(n2520) );
  NAND U3507 ( .A(n2520), .B(n9341), .Z(n2521) );
  NAND U3508 ( .A(n2519), .B(n2521), .Z(n9350) );
  XOR U3509 ( .A(n9366), .B(sreg[1675]), .Z(n2522) );
  NANDN U3510 ( .A(n9367), .B(n2522), .Z(n2523) );
  NAND U3511 ( .A(n9366), .B(sreg[1675]), .Z(n2524) );
  AND U3512 ( .A(n2523), .B(n2524), .Z(n9373) );
  NAND U3513 ( .A(n9390), .B(sreg[1678]), .Z(n2525) );
  XOR U3514 ( .A(sreg[1678]), .B(n9390), .Z(n2526) );
  NANDN U3515 ( .A(n9389), .B(n2526), .Z(n2527) );
  NAND U3516 ( .A(n2525), .B(n2527), .Z(n9398) );
  NAND U3517 ( .A(n9413), .B(sreg[1681]), .Z(n2528) );
  XOR U3518 ( .A(sreg[1681]), .B(n9413), .Z(n2529) );
  NAND U3519 ( .A(n2529), .B(n9412), .Z(n2530) );
  NAND U3520 ( .A(n2528), .B(n2530), .Z(n9419) );
  NAND U3521 ( .A(n9437), .B(sreg[1684]), .Z(n2531) );
  XOR U3522 ( .A(sreg[1684]), .B(n9437), .Z(n2532) );
  NAND U3523 ( .A(n2532), .B(n9436), .Z(n2533) );
  NAND U3524 ( .A(n2531), .B(n2533), .Z(n9445) );
  XOR U3525 ( .A(n9461), .B(sreg[1687]), .Z(n2534) );
  NANDN U3526 ( .A(n9462), .B(n2534), .Z(n2535) );
  NAND U3527 ( .A(n9461), .B(sreg[1687]), .Z(n2536) );
  AND U3528 ( .A(n2535), .B(n2536), .Z(n9468) );
  NAND U3529 ( .A(n9485), .B(sreg[1690]), .Z(n2537) );
  XOR U3530 ( .A(sreg[1690]), .B(n9485), .Z(n2538) );
  NANDN U3531 ( .A(n9484), .B(n2538), .Z(n2539) );
  NAND U3532 ( .A(n2537), .B(n2539), .Z(n9493) );
  XOR U3533 ( .A(n9511), .B(sreg[1693]), .Z(n2540) );
  NANDN U3534 ( .A(n9512), .B(n2540), .Z(n2541) );
  NAND U3535 ( .A(n9511), .B(sreg[1693]), .Z(n2542) );
  AND U3536 ( .A(n2541), .B(n2542), .Z(n9518) );
  NAND U3537 ( .A(n9535), .B(sreg[1696]), .Z(n2543) );
  XOR U3538 ( .A(sreg[1696]), .B(n9535), .Z(n2544) );
  NANDN U3539 ( .A(n9534), .B(n2544), .Z(n2545) );
  NAND U3540 ( .A(n2543), .B(n2545), .Z(n9544) );
  XOR U3541 ( .A(n9560), .B(sreg[1699]), .Z(n2546) );
  NANDN U3542 ( .A(n9561), .B(n2546), .Z(n2547) );
  NAND U3543 ( .A(n9560), .B(sreg[1699]), .Z(n2548) );
  AND U3544 ( .A(n2547), .B(n2548), .Z(n9567) );
  NAND U3545 ( .A(n9584), .B(sreg[1702]), .Z(n2549) );
  XOR U3546 ( .A(sreg[1702]), .B(n9584), .Z(n2550) );
  NANDN U3547 ( .A(n9583), .B(n2550), .Z(n2551) );
  NAND U3548 ( .A(n2549), .B(n2551), .Z(n9592) );
  NAND U3549 ( .A(n9608), .B(sreg[1705]), .Z(n2552) );
  XOR U3550 ( .A(sreg[1705]), .B(n9608), .Z(n2553) );
  NANDN U3551 ( .A(n9609), .B(n2553), .Z(n2554) );
  NAND U3552 ( .A(n2552), .B(n2554), .Z(n9617) );
  NAND U3553 ( .A(n9634), .B(sreg[1708]), .Z(n2555) );
  XOR U3554 ( .A(sreg[1708]), .B(n9634), .Z(n2556) );
  NANDN U3555 ( .A(n9633), .B(n2556), .Z(n2557) );
  NAND U3556 ( .A(n2555), .B(n2557), .Z(n9642) );
  XOR U3557 ( .A(n9658), .B(sreg[1711]), .Z(n2558) );
  NANDN U3558 ( .A(n9659), .B(n2558), .Z(n2559) );
  NAND U3559 ( .A(n9658), .B(sreg[1711]), .Z(n2560) );
  AND U3560 ( .A(n2559), .B(n2560), .Z(n9668) );
  NAND U3561 ( .A(n9685), .B(sreg[1714]), .Z(n2561) );
  XOR U3562 ( .A(sreg[1714]), .B(n9685), .Z(n2562) );
  NANDN U3563 ( .A(n9684), .B(n2562), .Z(n2563) );
  NAND U3564 ( .A(n2561), .B(n2563), .Z(n9693) );
  XOR U3565 ( .A(n9709), .B(sreg[1717]), .Z(n2564) );
  NANDN U3566 ( .A(n9710), .B(n2564), .Z(n2565) );
  NAND U3567 ( .A(n9709), .B(sreg[1717]), .Z(n2566) );
  AND U3568 ( .A(n2565), .B(n2566), .Z(n9716) );
  NAND U3569 ( .A(n9733), .B(sreg[1720]), .Z(n2567) );
  XOR U3570 ( .A(sreg[1720]), .B(n9733), .Z(n2568) );
  NANDN U3571 ( .A(n9732), .B(n2568), .Z(n2569) );
  NAND U3572 ( .A(n2567), .B(n2569), .Z(n9739) );
  XOR U3573 ( .A(n9755), .B(sreg[1723]), .Z(n2570) );
  NANDN U3574 ( .A(n9756), .B(n2570), .Z(n2571) );
  NAND U3575 ( .A(n9755), .B(sreg[1723]), .Z(n2572) );
  AND U3576 ( .A(n2571), .B(n2572), .Z(n9765) );
  NAND U3577 ( .A(n9782), .B(sreg[1726]), .Z(n2573) );
  XOR U3578 ( .A(sreg[1726]), .B(n9782), .Z(n2574) );
  NANDN U3579 ( .A(n9781), .B(n2574), .Z(n2575) );
  NAND U3580 ( .A(n2573), .B(n2575), .Z(n9790) );
  XOR U3581 ( .A(n9806), .B(sreg[1729]), .Z(n2576) );
  NANDN U3582 ( .A(n9807), .B(n2576), .Z(n2577) );
  NAND U3583 ( .A(n9806), .B(sreg[1729]), .Z(n2578) );
  AND U3584 ( .A(n2577), .B(n2578), .Z(n9813) );
  NAND U3585 ( .A(n9828), .B(sreg[1732]), .Z(n2579) );
  XOR U3586 ( .A(sreg[1732]), .B(n9828), .Z(n2580) );
  NAND U3587 ( .A(n2580), .B(n9827), .Z(n2581) );
  NAND U3588 ( .A(n2579), .B(n2581), .Z(n9836) );
  XOR U3589 ( .A(n9852), .B(sreg[1735]), .Z(n2582) );
  NANDN U3590 ( .A(n9853), .B(n2582), .Z(n2583) );
  NAND U3591 ( .A(n9852), .B(sreg[1735]), .Z(n2584) );
  AND U3592 ( .A(n2583), .B(n2584), .Z(n9862) );
  NAND U3593 ( .A(n9879), .B(sreg[1738]), .Z(n2585) );
  XOR U3594 ( .A(sreg[1738]), .B(n9879), .Z(n2586) );
  NANDN U3595 ( .A(n9878), .B(n2586), .Z(n2587) );
  NAND U3596 ( .A(n2585), .B(n2587), .Z(n9887) );
  XOR U3597 ( .A(n9903), .B(sreg[1741]), .Z(n2588) );
  NANDN U3598 ( .A(n9904), .B(n2588), .Z(n2589) );
  NAND U3599 ( .A(n9903), .B(sreg[1741]), .Z(n2590) );
  AND U3600 ( .A(n2589), .B(n2590), .Z(n9910) );
  NAND U3601 ( .A(n9927), .B(sreg[1744]), .Z(n2591) );
  XOR U3602 ( .A(sreg[1744]), .B(n9927), .Z(n2592) );
  NANDN U3603 ( .A(n9926), .B(n2592), .Z(n2593) );
  NAND U3604 ( .A(n2591), .B(n2593), .Z(n9935) );
  XOR U3605 ( .A(n9951), .B(sreg[1747]), .Z(n2594) );
  NANDN U3606 ( .A(n9952), .B(n2594), .Z(n2595) );
  NAND U3607 ( .A(n9951), .B(sreg[1747]), .Z(n2596) );
  AND U3608 ( .A(n2595), .B(n2596), .Z(n9958) );
  NAND U3609 ( .A(n9978), .B(sreg[1750]), .Z(n2597) );
  XOR U3610 ( .A(sreg[1750]), .B(n9978), .Z(n2598) );
  NANDN U3611 ( .A(n9977), .B(n2598), .Z(n2599) );
  NAND U3612 ( .A(n2597), .B(n2599), .Z(n9986) );
  XOR U3613 ( .A(n10002), .B(sreg[1753]), .Z(n2600) );
  NANDN U3614 ( .A(n10003), .B(n2600), .Z(n2601) );
  NAND U3615 ( .A(n10002), .B(sreg[1753]), .Z(n2602) );
  AND U3616 ( .A(n2601), .B(n2602), .Z(n10009) );
  NAND U3617 ( .A(n10026), .B(sreg[1756]), .Z(n2603) );
  XOR U3618 ( .A(sreg[1756]), .B(n10026), .Z(n2604) );
  NANDN U3619 ( .A(n10025), .B(n2604), .Z(n2605) );
  NAND U3620 ( .A(n2603), .B(n2605), .Z(n10034) );
  XOR U3621 ( .A(n10052), .B(sreg[1759]), .Z(n2606) );
  NANDN U3622 ( .A(n10053), .B(n2606), .Z(n2607) );
  NAND U3623 ( .A(n10052), .B(sreg[1759]), .Z(n2608) );
  AND U3624 ( .A(n2607), .B(n2608), .Z(n10059) );
  NAND U3625 ( .A(n10076), .B(sreg[1762]), .Z(n2609) );
  XOR U3626 ( .A(sreg[1762]), .B(n10076), .Z(n2610) );
  NANDN U3627 ( .A(n10075), .B(n2610), .Z(n2611) );
  NAND U3628 ( .A(n2609), .B(n2611), .Z(n10084) );
  NAND U3629 ( .A(n10102), .B(sreg[1765]), .Z(n2612) );
  XOR U3630 ( .A(sreg[1765]), .B(n10102), .Z(n2613) );
  NAND U3631 ( .A(n2613), .B(n10101), .Z(n2614) );
  NAND U3632 ( .A(n2612), .B(n2614), .Z(n10110) );
  NAND U3633 ( .A(n10127), .B(sreg[1768]), .Z(n2615) );
  XOR U3634 ( .A(sreg[1768]), .B(n10127), .Z(n2616) );
  NANDN U3635 ( .A(n10126), .B(n2616), .Z(n2617) );
  NAND U3636 ( .A(n2615), .B(n2617), .Z(n10135) );
  XOR U3637 ( .A(n10151), .B(sreg[1771]), .Z(n2618) );
  NANDN U3638 ( .A(n10152), .B(n2618), .Z(n2619) );
  NAND U3639 ( .A(n10151), .B(sreg[1771]), .Z(n2620) );
  AND U3640 ( .A(n2619), .B(n2620), .Z(n10158) );
  NAND U3641 ( .A(n10175), .B(sreg[1774]), .Z(n2621) );
  XOR U3642 ( .A(sreg[1774]), .B(n10175), .Z(n2622) );
  NANDN U3643 ( .A(n10174), .B(n2622), .Z(n2623) );
  NAND U3644 ( .A(n2621), .B(n2623), .Z(n10183) );
  NAND U3645 ( .A(n10198), .B(sreg[1777]), .Z(n2624) );
  XOR U3646 ( .A(sreg[1777]), .B(n10198), .Z(n2625) );
  NAND U3647 ( .A(n2625), .B(n10197), .Z(n2626) );
  NAND U3648 ( .A(n2624), .B(n2626), .Z(n10207) );
  NAND U3649 ( .A(n10224), .B(sreg[1780]), .Z(n2627) );
  XOR U3650 ( .A(sreg[1780]), .B(n10224), .Z(n2628) );
  NANDN U3651 ( .A(n10223), .B(n2628), .Z(n2629) );
  NAND U3652 ( .A(n2627), .B(n2629), .Z(n10232) );
  XOR U3653 ( .A(n10248), .B(sreg[1783]), .Z(n2630) );
  NANDN U3654 ( .A(n10249), .B(n2630), .Z(n2631) );
  NAND U3655 ( .A(n10248), .B(sreg[1783]), .Z(n2632) );
  AND U3656 ( .A(n2631), .B(n2632), .Z(n10255) );
  NAND U3657 ( .A(n10272), .B(sreg[1786]), .Z(n2633) );
  XOR U3658 ( .A(sreg[1786]), .B(n10272), .Z(n2634) );
  NANDN U3659 ( .A(n10271), .B(n2634), .Z(n2635) );
  NAND U3660 ( .A(n2633), .B(n2635), .Z(n10280) );
  XOR U3661 ( .A(n10296), .B(sreg[1789]), .Z(n2636) );
  NANDN U3662 ( .A(n10297), .B(n2636), .Z(n2637) );
  NAND U3663 ( .A(n10296), .B(sreg[1789]), .Z(n2638) );
  AND U3664 ( .A(n2637), .B(n2638), .Z(n10303) );
  NAND U3665 ( .A(n10323), .B(sreg[1792]), .Z(n2639) );
  XOR U3666 ( .A(sreg[1792]), .B(n10323), .Z(n2640) );
  NANDN U3667 ( .A(n10322), .B(n2640), .Z(n2641) );
  NAND U3668 ( .A(n2639), .B(n2641), .Z(n10331) );
  XOR U3669 ( .A(n10349), .B(sreg[1795]), .Z(n2642) );
  NANDN U3670 ( .A(n10350), .B(n2642), .Z(n2643) );
  NAND U3671 ( .A(n10349), .B(sreg[1795]), .Z(n2644) );
  AND U3672 ( .A(n2643), .B(n2644), .Z(n10356) );
  NAND U3673 ( .A(n10373), .B(sreg[1798]), .Z(n2645) );
  XOR U3674 ( .A(sreg[1798]), .B(n10373), .Z(n2646) );
  NANDN U3675 ( .A(n10372), .B(n2646), .Z(n2647) );
  NAND U3676 ( .A(n2645), .B(n2647), .Z(n10381) );
  XOR U3677 ( .A(n10397), .B(sreg[1801]), .Z(n2648) );
  NANDN U3678 ( .A(n10398), .B(n2648), .Z(n2649) );
  NAND U3679 ( .A(n10397), .B(sreg[1801]), .Z(n2650) );
  AND U3680 ( .A(n2649), .B(n2650), .Z(n10404) );
  NAND U3681 ( .A(n10421), .B(sreg[1804]), .Z(n2651) );
  XOR U3682 ( .A(sreg[1804]), .B(n10421), .Z(n2652) );
  NANDN U3683 ( .A(n10420), .B(n2652), .Z(n2653) );
  NAND U3684 ( .A(n2651), .B(n2653), .Z(n10429) );
  XOR U3685 ( .A(n10445), .B(sreg[1807]), .Z(n2654) );
  NANDN U3686 ( .A(n10446), .B(n2654), .Z(n2655) );
  NAND U3687 ( .A(n10445), .B(sreg[1807]), .Z(n2656) );
  AND U3688 ( .A(n2655), .B(n2656), .Z(n10455) );
  NAND U3689 ( .A(n10472), .B(sreg[1810]), .Z(n2657) );
  XOR U3690 ( .A(sreg[1810]), .B(n10472), .Z(n2658) );
  NANDN U3691 ( .A(n10471), .B(n2658), .Z(n2659) );
  NAND U3692 ( .A(n2657), .B(n2659), .Z(n10478) );
  XOR U3693 ( .A(n10494), .B(sreg[1813]), .Z(n2660) );
  NANDN U3694 ( .A(n10495), .B(n2660), .Z(n2661) );
  NAND U3695 ( .A(n10494), .B(sreg[1813]), .Z(n2662) );
  AND U3696 ( .A(n2661), .B(n2662), .Z(n10501) );
  NAND U3697 ( .A(n10518), .B(sreg[1816]), .Z(n2663) );
  XOR U3698 ( .A(sreg[1816]), .B(n10518), .Z(n2664) );
  NANDN U3699 ( .A(n10517), .B(n2664), .Z(n2665) );
  NAND U3700 ( .A(n2663), .B(n2665), .Z(n10526) );
  XOR U3701 ( .A(n10542), .B(sreg[1819]), .Z(n2666) );
  NANDN U3702 ( .A(n10543), .B(n2666), .Z(n2667) );
  NAND U3703 ( .A(n10542), .B(sreg[1819]), .Z(n2668) );
  AND U3704 ( .A(n2667), .B(n2668), .Z(n10552) );
  NAND U3705 ( .A(n10569), .B(sreg[1822]), .Z(n2669) );
  XOR U3706 ( .A(sreg[1822]), .B(n10569), .Z(n2670) );
  NANDN U3707 ( .A(n10568), .B(n2670), .Z(n2671) );
  NAND U3708 ( .A(n2669), .B(n2671), .Z(n10577) );
  XOR U3709 ( .A(n10593), .B(sreg[1825]), .Z(n2672) );
  NANDN U3710 ( .A(n10594), .B(n2672), .Z(n2673) );
  NAND U3711 ( .A(n10593), .B(sreg[1825]), .Z(n2674) );
  AND U3712 ( .A(n2673), .B(n2674), .Z(n10600) );
  NAND U3713 ( .A(n10617), .B(sreg[1828]), .Z(n2675) );
  XOR U3714 ( .A(sreg[1828]), .B(n10617), .Z(n2676) );
  NANDN U3715 ( .A(n10616), .B(n2676), .Z(n2677) );
  NAND U3716 ( .A(n2675), .B(n2677), .Z(n10623) );
  NAND U3717 ( .A(n10639), .B(sreg[1831]), .Z(n2678) );
  XOR U3718 ( .A(sreg[1831]), .B(n10639), .Z(n2679) );
  NANDN U3719 ( .A(n10640), .B(n2679), .Z(n2680) );
  NAND U3720 ( .A(n2678), .B(n2680), .Z(n10648) );
  NAND U3721 ( .A(n10668), .B(sreg[1834]), .Z(n2681) );
  XOR U3722 ( .A(sreg[1834]), .B(n10668), .Z(n2682) );
  NANDN U3723 ( .A(n10667), .B(n2682), .Z(n2683) );
  NAND U3724 ( .A(n2681), .B(n2683), .Z(n10676) );
  NAND U3725 ( .A(n10691), .B(sreg[1837]), .Z(n2684) );
  XOR U3726 ( .A(sreg[1837]), .B(n10691), .Z(n2685) );
  NAND U3727 ( .A(n2685), .B(n10690), .Z(n2686) );
  NAND U3728 ( .A(n2684), .B(n2686), .Z(n10697) );
  NAND U3729 ( .A(n10714), .B(sreg[1840]), .Z(n2687) );
  XOR U3730 ( .A(sreg[1840]), .B(n10714), .Z(n2688) );
  NANDN U3731 ( .A(n10713), .B(n2688), .Z(n2689) );
  NAND U3732 ( .A(n2687), .B(n2689), .Z(n10722) );
  NAND U3733 ( .A(n10737), .B(sreg[1843]), .Z(n2690) );
  XOR U3734 ( .A(sreg[1843]), .B(n10737), .Z(n2691) );
  NAND U3735 ( .A(n2691), .B(n10736), .Z(n2692) );
  NAND U3736 ( .A(n2690), .B(n2692), .Z(n10745) );
  NAND U3737 ( .A(n10765), .B(sreg[1846]), .Z(n2693) );
  XOR U3738 ( .A(sreg[1846]), .B(n10765), .Z(n2694) );
  NANDN U3739 ( .A(n10764), .B(n2694), .Z(n2695) );
  NAND U3740 ( .A(n2693), .B(n2695), .Z(n10773) );
  NAND U3741 ( .A(n10790), .B(sreg[1849]), .Z(n2696) );
  XOR U3742 ( .A(sreg[1849]), .B(n10790), .Z(n2697) );
  NANDN U3743 ( .A(n10789), .B(n2697), .Z(n2698) );
  NAND U3744 ( .A(n2696), .B(n2698), .Z(n10798) );
  NAND U3745 ( .A(n10815), .B(sreg[1852]), .Z(n2699) );
  XOR U3746 ( .A(sreg[1852]), .B(n10815), .Z(n2700) );
  NANDN U3747 ( .A(n10814), .B(n2700), .Z(n2701) );
  NAND U3748 ( .A(n2699), .B(n2701), .Z(n10823) );
  XOR U3749 ( .A(n10839), .B(sreg[1855]), .Z(n2702) );
  NANDN U3750 ( .A(n10840), .B(n2702), .Z(n2703) );
  NAND U3751 ( .A(n10839), .B(sreg[1855]), .Z(n2704) );
  AND U3752 ( .A(n2703), .B(n2704), .Z(n10846) );
  XOR U3753 ( .A(n10864), .B(sreg[1858]), .Z(n2705) );
  NANDN U3754 ( .A(n10865), .B(n2705), .Z(n2706) );
  NAND U3755 ( .A(n10864), .B(sreg[1858]), .Z(n2707) );
  AND U3756 ( .A(n2706), .B(n2707), .Z(n10871) );
  NAND U3757 ( .A(n10889), .B(sreg[1861]), .Z(n2708) );
  XOR U3758 ( .A(sreg[1861]), .B(n10889), .Z(n2709) );
  NANDN U3759 ( .A(n10890), .B(n2709), .Z(n2710) );
  NAND U3760 ( .A(n2708), .B(n2710), .Z(n10898) );
  NAND U3761 ( .A(n10914), .B(sreg[1864]), .Z(n2711) );
  XOR U3762 ( .A(sreg[1864]), .B(n10914), .Z(n2712) );
  NANDN U3763 ( .A(n10915), .B(n2712), .Z(n2713) );
  NAND U3764 ( .A(n2711), .B(n2713), .Z(n10923) );
  XOR U3765 ( .A(n10942), .B(sreg[1867]), .Z(n2714) );
  NANDN U3766 ( .A(n10943), .B(n2714), .Z(n2715) );
  NAND U3767 ( .A(n10942), .B(sreg[1867]), .Z(n2716) );
  AND U3768 ( .A(n2715), .B(n2716), .Z(n10949) );
  NAND U3769 ( .A(n10966), .B(sreg[1870]), .Z(n2717) );
  XOR U3770 ( .A(sreg[1870]), .B(n10966), .Z(n2718) );
  NANDN U3771 ( .A(n10965), .B(n2718), .Z(n2719) );
  NAND U3772 ( .A(n2717), .B(n2719), .Z(n10974) );
  NAND U3773 ( .A(n10989), .B(sreg[1873]), .Z(n2720) );
  XOR U3774 ( .A(sreg[1873]), .B(n10989), .Z(n2721) );
  NAND U3775 ( .A(n2721), .B(n10988), .Z(n2722) );
  NAND U3776 ( .A(n2720), .B(n2722), .Z(n10995) );
  NAND U3777 ( .A(n11013), .B(sreg[1876]), .Z(n2723) );
  XOR U3778 ( .A(sreg[1876]), .B(n11013), .Z(n2724) );
  NANDN U3779 ( .A(n11014), .B(n2724), .Z(n2725) );
  NAND U3780 ( .A(n2723), .B(n2725), .Z(n11022) );
  NAND U3781 ( .A(n11040), .B(sreg[1879]), .Z(n2726) );
  XOR U3782 ( .A(sreg[1879]), .B(n11040), .Z(n2727) );
  NANDN U3783 ( .A(n11041), .B(n2727), .Z(n2728) );
  NAND U3784 ( .A(n2726), .B(n2728), .Z(n11049) );
  NAND U3785 ( .A(n11066), .B(sreg[1882]), .Z(n2729) );
  XOR U3786 ( .A(sreg[1882]), .B(n11066), .Z(n2730) );
  NANDN U3787 ( .A(n11065), .B(n2730), .Z(n2731) );
  NAND U3788 ( .A(n2729), .B(n2731), .Z(n11074) );
  XOR U3789 ( .A(n11092), .B(sreg[1885]), .Z(n2732) );
  NANDN U3790 ( .A(n11093), .B(n2732), .Z(n2733) );
  NAND U3791 ( .A(n11092), .B(sreg[1885]), .Z(n2734) );
  AND U3792 ( .A(n2733), .B(n2734), .Z(n11102) );
  NAND U3793 ( .A(n11119), .B(sreg[1888]), .Z(n2735) );
  XOR U3794 ( .A(sreg[1888]), .B(n11119), .Z(n2736) );
  NANDN U3795 ( .A(n11118), .B(n2736), .Z(n2737) );
  NAND U3796 ( .A(n2735), .B(n2737), .Z(n11127) );
  XOR U3797 ( .A(n11143), .B(sreg[1891]), .Z(n2738) );
  NANDN U3798 ( .A(n11144), .B(n2738), .Z(n2739) );
  NAND U3799 ( .A(n11143), .B(sreg[1891]), .Z(n2740) );
  AND U3800 ( .A(n2739), .B(n2740), .Z(n11150) );
  NAND U3801 ( .A(n11167), .B(sreg[1894]), .Z(n2741) );
  XOR U3802 ( .A(sreg[1894]), .B(n11167), .Z(n2742) );
  NANDN U3803 ( .A(n11166), .B(n2742), .Z(n2743) );
  NAND U3804 ( .A(n2741), .B(n2743), .Z(n11173) );
  XOR U3805 ( .A(n11189), .B(sreg[1897]), .Z(n2744) );
  NANDN U3806 ( .A(n11190), .B(n2744), .Z(n2745) );
  NAND U3807 ( .A(n11189), .B(sreg[1897]), .Z(n2746) );
  AND U3808 ( .A(n2745), .B(n2746), .Z(n11199) );
  NAND U3809 ( .A(n11214), .B(sreg[1900]), .Z(n2747) );
  XOR U3810 ( .A(sreg[1900]), .B(n11214), .Z(n2748) );
  NAND U3811 ( .A(n2748), .B(n11213), .Z(n2749) );
  NAND U3812 ( .A(n2747), .B(n2749), .Z(n11222) );
  XOR U3813 ( .A(n11238), .B(sreg[1903]), .Z(n2750) );
  NANDN U3814 ( .A(n11239), .B(n2750), .Z(n2751) );
  NAND U3815 ( .A(n11238), .B(sreg[1903]), .Z(n2752) );
  AND U3816 ( .A(n2751), .B(n2752), .Z(n11245) );
  NAND U3817 ( .A(n11262), .B(sreg[1906]), .Z(n2753) );
  XOR U3818 ( .A(sreg[1906]), .B(n11262), .Z(n2754) );
  NANDN U3819 ( .A(n11261), .B(n2754), .Z(n2755) );
  NAND U3820 ( .A(n2753), .B(n2755), .Z(n11270) );
  XOR U3821 ( .A(n11286), .B(sreg[1909]), .Z(n2756) );
  NANDN U3822 ( .A(n11287), .B(n2756), .Z(n2757) );
  NAND U3823 ( .A(n11286), .B(sreg[1909]), .Z(n2758) );
  AND U3824 ( .A(n2757), .B(n2758), .Z(n11296) );
  NAND U3825 ( .A(n11313), .B(sreg[1912]), .Z(n2759) );
  XOR U3826 ( .A(sreg[1912]), .B(n11313), .Z(n2760) );
  NANDN U3827 ( .A(n11312), .B(n2760), .Z(n2761) );
  NAND U3828 ( .A(n2759), .B(n2761), .Z(n11321) );
  XOR U3829 ( .A(n11337), .B(sreg[1915]), .Z(n2762) );
  NANDN U3830 ( .A(n11338), .B(n2762), .Z(n2763) );
  NAND U3831 ( .A(n11337), .B(sreg[1915]), .Z(n2764) );
  AND U3832 ( .A(n2763), .B(n2764), .Z(n11344) );
  NAND U3833 ( .A(n11362), .B(sreg[1918]), .Z(n2765) );
  XOR U3834 ( .A(sreg[1918]), .B(n11362), .Z(n2766) );
  NANDN U3835 ( .A(n11363), .B(n2766), .Z(n2767) );
  NAND U3836 ( .A(n2765), .B(n2767), .Z(n11371) );
  XOR U3837 ( .A(n11389), .B(sreg[1921]), .Z(n2768) );
  NANDN U3838 ( .A(n11390), .B(n2768), .Z(n2769) );
  NAND U3839 ( .A(n11389), .B(sreg[1921]), .Z(n2770) );
  AND U3840 ( .A(n2769), .B(n2770), .Z(n11396) );
  XOR U3841 ( .A(n11414), .B(sreg[1924]), .Z(n2771) );
  NANDN U3842 ( .A(n11415), .B(n2771), .Z(n2772) );
  NAND U3843 ( .A(n11414), .B(sreg[1924]), .Z(n2773) );
  AND U3844 ( .A(n2772), .B(n2773), .Z(n11421) );
  NAND U3845 ( .A(n11437), .B(sreg[1927]), .Z(n2774) );
  XOR U3846 ( .A(sreg[1927]), .B(n11437), .Z(n2775) );
  NANDN U3847 ( .A(n11438), .B(n2775), .Z(n2776) );
  NAND U3848 ( .A(n2774), .B(n2776), .Z(n11446) );
  NAND U3849 ( .A(n11466), .B(sreg[1930]), .Z(n2777) );
  XOR U3850 ( .A(sreg[1930]), .B(n11466), .Z(n2778) );
  NANDN U3851 ( .A(n11465), .B(n2778), .Z(n2779) );
  NAND U3852 ( .A(n2777), .B(n2779), .Z(n11474) );
  NAND U3853 ( .A(n11490), .B(sreg[1933]), .Z(n2780) );
  XOR U3854 ( .A(sreg[1933]), .B(n11490), .Z(n2781) );
  NANDN U3855 ( .A(n11491), .B(n2781), .Z(n2782) );
  NAND U3856 ( .A(n2780), .B(n2782), .Z(n11499) );
  NAND U3857 ( .A(n11516), .B(sreg[1936]), .Z(n2783) );
  XOR U3858 ( .A(sreg[1936]), .B(n11516), .Z(n2784) );
  NANDN U3859 ( .A(n11515), .B(n2784), .Z(n2785) );
  NAND U3860 ( .A(n2783), .B(n2785), .Z(n11524) );
  NAND U3861 ( .A(n11539), .B(sreg[1939]), .Z(n2786) );
  XOR U3862 ( .A(sreg[1939]), .B(n11539), .Z(n2787) );
  NAND U3863 ( .A(n2787), .B(n11538), .Z(n2788) );
  NAND U3864 ( .A(n2786), .B(n2788), .Z(n11545) );
  NAND U3865 ( .A(n11563), .B(sreg[1942]), .Z(n2789) );
  XOR U3866 ( .A(sreg[1942]), .B(n11563), .Z(n2790) );
  NANDN U3867 ( .A(n11564), .B(n2790), .Z(n2791) );
  NAND U3868 ( .A(n2789), .B(n2791), .Z(n11572) );
  XOR U3869 ( .A(n11588), .B(sreg[1945]), .Z(n2792) );
  NANDN U3870 ( .A(n11589), .B(n2792), .Z(n2793) );
  NAND U3871 ( .A(n11588), .B(sreg[1945]), .Z(n2794) );
  AND U3872 ( .A(n2793), .B(n2794), .Z(n11598) );
  NAND U3873 ( .A(n11615), .B(sreg[1948]), .Z(n2795) );
  XOR U3874 ( .A(sreg[1948]), .B(n11615), .Z(n2796) );
  NANDN U3875 ( .A(n11614), .B(n2796), .Z(n2797) );
  NAND U3876 ( .A(n2795), .B(n2797), .Z(n11623) );
  XOR U3877 ( .A(n11639), .B(sreg[1951]), .Z(n2798) );
  NANDN U3878 ( .A(n11640), .B(n2798), .Z(n2799) );
  NAND U3879 ( .A(n11639), .B(sreg[1951]), .Z(n2800) );
  AND U3880 ( .A(n2799), .B(n2800), .Z(n11646) );
  NAND U3881 ( .A(n11664), .B(sreg[1954]), .Z(n2801) );
  XOR U3882 ( .A(sreg[1954]), .B(n11664), .Z(n2802) );
  NANDN U3883 ( .A(n11665), .B(n2802), .Z(n2803) );
  NAND U3884 ( .A(n2801), .B(n2803), .Z(n11673) );
  XOR U3885 ( .A(n11689), .B(sreg[1957]), .Z(n2804) );
  NANDN U3886 ( .A(n11690), .B(n2804), .Z(n2805) );
  NAND U3887 ( .A(n11689), .B(sreg[1957]), .Z(n2806) );
  AND U3888 ( .A(n2805), .B(n2806), .Z(n11696) );
  NAND U3889 ( .A(n11712), .B(sreg[1960]), .Z(n2807) );
  XOR U3890 ( .A(sreg[1960]), .B(n11712), .Z(n2808) );
  NANDN U3891 ( .A(n11713), .B(n2808), .Z(n2809) );
  NAND U3892 ( .A(n2807), .B(n2809), .Z(n11721) );
  XOR U3893 ( .A(n11740), .B(sreg[1963]), .Z(n2810) );
  NANDN U3894 ( .A(n11741), .B(n2810), .Z(n2811) );
  NAND U3895 ( .A(n11740), .B(sreg[1963]), .Z(n2812) );
  AND U3896 ( .A(n2811), .B(n2812), .Z(n11747) );
  NAND U3897 ( .A(n11764), .B(sreg[1966]), .Z(n2813) );
  XOR U3898 ( .A(sreg[1966]), .B(n11764), .Z(n2814) );
  NANDN U3899 ( .A(n11763), .B(n2814), .Z(n2815) );
  NAND U3900 ( .A(n2813), .B(n2815), .Z(n11772) );
  NAND U3901 ( .A(n11790), .B(sreg[1969]), .Z(n2816) );
  XOR U3902 ( .A(sreg[1969]), .B(n11790), .Z(n2817) );
  NANDN U3903 ( .A(n11791), .B(n2817), .Z(n2818) );
  NAND U3904 ( .A(n2816), .B(n2818), .Z(n11799) );
  NAND U3905 ( .A(n11817), .B(sreg[1972]), .Z(n2819) );
  XOR U3906 ( .A(sreg[1972]), .B(n11817), .Z(n2820) );
  NANDN U3907 ( .A(n11818), .B(n2820), .Z(n2821) );
  NAND U3908 ( .A(n2819), .B(n2821), .Z(n11826) );
  XOR U3909 ( .A(n11842), .B(sreg[1975]), .Z(n2822) );
  NANDN U3910 ( .A(n11843), .B(n2822), .Z(n2823) );
  NAND U3911 ( .A(n11842), .B(sreg[1975]), .Z(n2824) );
  AND U3912 ( .A(n2823), .B(n2824), .Z(n11849) );
  NAND U3913 ( .A(n11866), .B(sreg[1978]), .Z(n2825) );
  XOR U3914 ( .A(sreg[1978]), .B(n11866), .Z(n2826) );
  NANDN U3915 ( .A(n11865), .B(n2826), .Z(n2827) );
  NAND U3916 ( .A(n2825), .B(n2827), .Z(n11874) );
  XOR U3917 ( .A(n11890), .B(sreg[1981]), .Z(n2828) );
  NANDN U3918 ( .A(n11891), .B(n2828), .Z(n2829) );
  NAND U3919 ( .A(n11890), .B(sreg[1981]), .Z(n2830) );
  AND U3920 ( .A(n2829), .B(n2830), .Z(n11900) );
  NAND U3921 ( .A(n11917), .B(sreg[1984]), .Z(n2831) );
  XOR U3922 ( .A(sreg[1984]), .B(n11917), .Z(n2832) );
  NANDN U3923 ( .A(n11916), .B(n2832), .Z(n2833) );
  NAND U3924 ( .A(n2831), .B(n2833), .Z(n11925) );
  XOR U3925 ( .A(n11941), .B(sreg[1987]), .Z(n2834) );
  NANDN U3926 ( .A(n11942), .B(n2834), .Z(n2835) );
  NAND U3927 ( .A(n11941), .B(sreg[1987]), .Z(n2836) );
  AND U3928 ( .A(n2835), .B(n2836), .Z(n11948) );
  NAND U3929 ( .A(n11965), .B(sreg[1990]), .Z(n2837) );
  XOR U3930 ( .A(sreg[1990]), .B(n11965), .Z(n2838) );
  NANDN U3931 ( .A(n11964), .B(n2838), .Z(n2839) );
  NAND U3932 ( .A(n2837), .B(n2839), .Z(n11973) );
  XOR U3933 ( .A(n11989), .B(sreg[1993]), .Z(n2840) );
  NANDN U3934 ( .A(n11990), .B(n2840), .Z(n2841) );
  NAND U3935 ( .A(n11989), .B(sreg[1993]), .Z(n2842) );
  AND U3936 ( .A(n2841), .B(n2842), .Z(n11996) );
  NAND U3937 ( .A(n12016), .B(sreg[1996]), .Z(n2843) );
  XOR U3938 ( .A(sreg[1996]), .B(n12016), .Z(n2844) );
  NANDN U3939 ( .A(n12015), .B(n2844), .Z(n2845) );
  NAND U3940 ( .A(n2843), .B(n2845), .Z(n12022) );
  XOR U3941 ( .A(n12040), .B(sreg[1999]), .Z(n2846) );
  NANDN U3942 ( .A(n12041), .B(n2846), .Z(n2847) );
  NAND U3943 ( .A(n12040), .B(sreg[1999]), .Z(n2848) );
  AND U3944 ( .A(n2847), .B(n2848), .Z(n12047) );
  NAND U3945 ( .A(n12064), .B(sreg[2002]), .Z(n2849) );
  XOR U3946 ( .A(sreg[2002]), .B(n12064), .Z(n2850) );
  NANDN U3947 ( .A(n12063), .B(n2850), .Z(n2851) );
  NAND U3948 ( .A(n2849), .B(n2851), .Z(n12072) );
  NAND U3949 ( .A(n12087), .B(sreg[2005]), .Z(n2852) );
  XOR U3950 ( .A(sreg[2005]), .B(n12087), .Z(n2853) );
  NAND U3951 ( .A(n2853), .B(n12086), .Z(n2854) );
  NAND U3952 ( .A(n2852), .B(n2854), .Z(n12093) );
  NAND U3953 ( .A(n12113), .B(sreg[2008]), .Z(n2855) );
  XOR U3954 ( .A(sreg[2008]), .B(n12113), .Z(n2856) );
  NANDN U3955 ( .A(n12112), .B(n2856), .Z(n2857) );
  NAND U3956 ( .A(n2855), .B(n2857), .Z(n12119) );
  XOR U3957 ( .A(n12135), .B(sreg[2011]), .Z(n2858) );
  NANDN U3958 ( .A(n12136), .B(n2858), .Z(n2859) );
  NAND U3959 ( .A(n12135), .B(sreg[2011]), .Z(n2860) );
  AND U3960 ( .A(n2859), .B(n2860), .Z(n12142) );
  NAND U3961 ( .A(n12159), .B(sreg[2014]), .Z(n2861) );
  XOR U3962 ( .A(sreg[2014]), .B(n12159), .Z(n2862) );
  NANDN U3963 ( .A(n12158), .B(n2862), .Z(n2863) );
  NAND U3964 ( .A(n2861), .B(n2863), .Z(n12167) );
  XOR U3965 ( .A(n12183), .B(sreg[2017]), .Z(n2864) );
  NANDN U3966 ( .A(n12184), .B(n2864), .Z(n2865) );
  NAND U3967 ( .A(n12183), .B(sreg[2017]), .Z(n2866) );
  AND U3968 ( .A(n2865), .B(n2866), .Z(n12190) );
  NAND U3969 ( .A(n12210), .B(sreg[2020]), .Z(n2867) );
  XOR U3970 ( .A(sreg[2020]), .B(n12210), .Z(n2868) );
  NANDN U3971 ( .A(n12209), .B(n2868), .Z(n2869) );
  NAND U3972 ( .A(n2867), .B(n2869), .Z(n12216) );
  NAND U3973 ( .A(n12232), .B(sreg[2023]), .Z(n2870) );
  XOR U3974 ( .A(sreg[2023]), .B(n12232), .Z(n2871) );
  NANDN U3975 ( .A(n12233), .B(n2871), .Z(n2872) );
  NAND U3976 ( .A(n2870), .B(n2872), .Z(n12241) );
  NAND U3977 ( .A(n12258), .B(sreg[2026]), .Z(n2873) );
  XOR U3978 ( .A(sreg[2026]), .B(n12258), .Z(n2874) );
  NANDN U3979 ( .A(n12257), .B(n2874), .Z(n2875) );
  NAND U3980 ( .A(n2873), .B(n2875), .Z(n12266) );
  NAND U3981 ( .A(n12281), .B(sreg[2029]), .Z(n2876) );
  XOR U3982 ( .A(sreg[2029]), .B(n12281), .Z(n2877) );
  NAND U3983 ( .A(n2877), .B(n12280), .Z(n2878) );
  NAND U3984 ( .A(n2876), .B(n2878), .Z(n12289) );
  NAND U3985 ( .A(n12306), .B(sreg[2032]), .Z(n2879) );
  XOR U3986 ( .A(sreg[2032]), .B(n12306), .Z(n2880) );
  NANDN U3987 ( .A(n12305), .B(n2880), .Z(n2881) );
  NAND U3988 ( .A(n2879), .B(n2881), .Z(n12314) );
  XOR U3989 ( .A(n12332), .B(sreg[2035]), .Z(n2882) );
  NANDN U3990 ( .A(n12333), .B(n2882), .Z(n2883) );
  NAND U3991 ( .A(n12332), .B(sreg[2035]), .Z(n2884) );
  AND U3992 ( .A(n2883), .B(n2884), .Z(n12339) );
  NAND U3993 ( .A(n12356), .B(sreg[2038]), .Z(n2885) );
  XOR U3994 ( .A(sreg[2038]), .B(n12356), .Z(n2886) );
  NANDN U3995 ( .A(n12355), .B(n2886), .Z(n2887) );
  NAND U3996 ( .A(n2885), .B(n2887), .Z(n12364) );
  XOR U3997 ( .A(n12380), .B(sreg[2041]), .Z(n2888) );
  NANDN U3998 ( .A(n12381), .B(n2888), .Z(n2889) );
  NAND U3999 ( .A(n12380), .B(sreg[2041]), .Z(n2890) );
  AND U4000 ( .A(n2889), .B(n2890), .Z(n12387) );
  NAND U4001 ( .A(n12408), .B(n12407), .Z(n2891) );
  XOR U4002 ( .A(n12407), .B(n12408), .Z(n2892) );
  NAND U4003 ( .A(n2892), .B(sreg[2044]), .Z(n2893) );
  NAND U4004 ( .A(n2891), .B(n2893), .Z(n12415) );
  OR U4005 ( .A(n4137), .B(n4136), .Z(n2894) );
  NAND U4006 ( .A(n4139), .B(n4138), .Z(n2895) );
  NAND U4007 ( .A(n2894), .B(n2895), .Z(n4146) );
  OR U4008 ( .A(n4205), .B(n4204), .Z(n2896) );
  NAND U4009 ( .A(n4207), .B(n4206), .Z(n2897) );
  NAND U4010 ( .A(n2896), .B(n2897), .Z(n4214) );
  NAND U4011 ( .A(n4026), .B(n4025), .Z(n2898) );
  XOR U4012 ( .A(n4025), .B(n4026), .Z(n2899) );
  NAND U4013 ( .A(n2899), .B(sreg[1027]), .Z(n2900) );
  NAND U4014 ( .A(n2898), .B(n2900), .Z(n4043) );
  XOR U4015 ( .A(n4061), .B(n4060), .Z(n2901) );
  NANDN U4016 ( .A(sreg[1030]), .B(n2901), .Z(n2902) );
  NAND U4017 ( .A(n4061), .B(n4060), .Z(n2903) );
  AND U4018 ( .A(n2902), .B(n2903), .Z(n4067) );
  XOR U4019 ( .A(n4085), .B(sreg[1033]), .Z(n2904) );
  NANDN U4020 ( .A(n4086), .B(n2904), .Z(n2905) );
  NAND U4021 ( .A(n4085), .B(sreg[1033]), .Z(n2906) );
  AND U4022 ( .A(n2905), .B(n2906), .Z(n4092) );
  NAND U4023 ( .A(n4109), .B(sreg[1036]), .Z(n2907) );
  XOR U4024 ( .A(sreg[1036]), .B(n4109), .Z(n2908) );
  NANDN U4025 ( .A(n4108), .B(n2908), .Z(n2909) );
  NAND U4026 ( .A(n2907), .B(n2909), .Z(n4117) );
  XOR U4027 ( .A(n4133), .B(sreg[1039]), .Z(n2910) );
  NANDN U4028 ( .A(n4134), .B(n2910), .Z(n2911) );
  NAND U4029 ( .A(n4133), .B(sreg[1039]), .Z(n2912) );
  AND U4030 ( .A(n2911), .B(n2912), .Z(n4140) );
  NAND U4031 ( .A(n4175), .B(sreg[1044]), .Z(n2913) );
  XOR U4032 ( .A(sreg[1044]), .B(n4175), .Z(n2914) );
  NAND U4033 ( .A(n2914), .B(n4174), .Z(n2915) );
  NAND U4034 ( .A(n2913), .B(n2915), .Z(n4183) );
  NAND U4035 ( .A(n4202), .B(n4201), .Z(n2916) );
  XOR U4036 ( .A(n4201), .B(n4202), .Z(n2917) );
  NANDN U4037 ( .A(sreg[1047]), .B(n2917), .Z(n2918) );
  NAND U4038 ( .A(n2916), .B(n2918), .Z(n4208) );
  NAND U4039 ( .A(n4245), .B(sreg[1052]), .Z(n2919) );
  XOR U4040 ( .A(sreg[1052]), .B(n4245), .Z(n2920) );
  NANDN U4041 ( .A(n4244), .B(n2920), .Z(n2921) );
  NAND U4042 ( .A(n2919), .B(n2921), .Z(n4253) );
  XOR U4043 ( .A(n4272), .B(sreg[1055]), .Z(n2922) );
  NANDN U4044 ( .A(n4273), .B(n2922), .Z(n2923) );
  NAND U4045 ( .A(n4272), .B(sreg[1055]), .Z(n2924) );
  AND U4046 ( .A(n2923), .B(n2924), .Z(n4279) );
  NAND U4047 ( .A(n4296), .B(sreg[1058]), .Z(n2925) );
  XOR U4048 ( .A(sreg[1058]), .B(n4296), .Z(n2926) );
  NANDN U4049 ( .A(n4295), .B(n2926), .Z(n2927) );
  NAND U4050 ( .A(n2925), .B(n2927), .Z(n4304) );
  XOR U4051 ( .A(n4320), .B(sreg[1061]), .Z(n2928) );
  NANDN U4052 ( .A(n4321), .B(n2928), .Z(n2929) );
  NAND U4053 ( .A(n4320), .B(sreg[1061]), .Z(n2930) );
  AND U4054 ( .A(n2929), .B(n2930), .Z(n4327) );
  NAND U4055 ( .A(n4344), .B(sreg[1064]), .Z(n2931) );
  XOR U4056 ( .A(sreg[1064]), .B(n4344), .Z(n2932) );
  NANDN U4057 ( .A(n4343), .B(n2932), .Z(n2933) );
  NAND U4058 ( .A(n2931), .B(n2933), .Z(n4350) );
  NAND U4059 ( .A(n4369), .B(sreg[1067]), .Z(n2934) );
  XOR U4060 ( .A(sreg[1067]), .B(n4369), .Z(n2935) );
  NANDN U4061 ( .A(n4370), .B(n2935), .Z(n2936) );
  NAND U4062 ( .A(n2934), .B(n2936), .Z(n4378) );
  NAND U4063 ( .A(n4395), .B(sreg[1070]), .Z(n2937) );
  XOR U4064 ( .A(sreg[1070]), .B(n4395), .Z(n2938) );
  NANDN U4065 ( .A(n4394), .B(n2938), .Z(n2939) );
  NAND U4066 ( .A(n2937), .B(n2939), .Z(n4403) );
  XOR U4067 ( .A(n4419), .B(sreg[1073]), .Z(n2940) );
  NANDN U4068 ( .A(n4420), .B(n2940), .Z(n2941) );
  NAND U4069 ( .A(n4419), .B(sreg[1073]), .Z(n2942) );
  AND U4070 ( .A(n2941), .B(n2942), .Z(n4426) );
  NAND U4071 ( .A(n4441), .B(sreg[1076]), .Z(n2943) );
  XOR U4072 ( .A(sreg[1076]), .B(n4441), .Z(n2944) );
  NAND U4073 ( .A(n2944), .B(n4440), .Z(n2945) );
  NAND U4074 ( .A(n2943), .B(n2945), .Z(n4449) );
  XOR U4075 ( .A(n4465), .B(sreg[1079]), .Z(n2946) );
  NANDN U4076 ( .A(n4466), .B(n2946), .Z(n2947) );
  NAND U4077 ( .A(n4465), .B(sreg[1079]), .Z(n2948) );
  AND U4078 ( .A(n2947), .B(n2948), .Z(n4475) );
  NAND U4079 ( .A(n4492), .B(sreg[1082]), .Z(n2949) );
  XOR U4080 ( .A(sreg[1082]), .B(n4492), .Z(n2950) );
  NANDN U4081 ( .A(n4491), .B(n2950), .Z(n2951) );
  NAND U4082 ( .A(n2949), .B(n2951), .Z(n4500) );
  XOR U4083 ( .A(n4518), .B(sreg[1085]), .Z(n2952) );
  NANDN U4084 ( .A(n4519), .B(n2952), .Z(n2953) );
  NAND U4085 ( .A(n4518), .B(sreg[1085]), .Z(n2954) );
  AND U4086 ( .A(n2953), .B(n2954), .Z(n4525) );
  NAND U4087 ( .A(n4543), .B(sreg[1088]), .Z(n2955) );
  XOR U4088 ( .A(sreg[1088]), .B(n4543), .Z(n2956) );
  NANDN U4089 ( .A(n4544), .B(n2956), .Z(n2957) );
  NAND U4090 ( .A(n2955), .B(n2957), .Z(n4552) );
  XOR U4091 ( .A(n4568), .B(sreg[1091]), .Z(n2958) );
  NANDN U4092 ( .A(n4569), .B(n2958), .Z(n2959) );
  NAND U4093 ( .A(n4568), .B(sreg[1091]), .Z(n2960) );
  AND U4094 ( .A(n2959), .B(n2960), .Z(n4575) );
  NAND U4095 ( .A(n4590), .B(sreg[1094]), .Z(n2961) );
  XOR U4096 ( .A(sreg[1094]), .B(n4590), .Z(n2962) );
  NAND U4097 ( .A(n2962), .B(n4589), .Z(n2963) );
  NAND U4098 ( .A(n2961), .B(n2963), .Z(n4598) );
  NAND U4099 ( .A(n4616), .B(sreg[1097]), .Z(n2964) );
  XOR U4100 ( .A(sreg[1097]), .B(n4616), .Z(n2965) );
  NAND U4101 ( .A(n2965), .B(n4615), .Z(n2966) );
  NAND U4102 ( .A(n2964), .B(n2966), .Z(n4622) );
  NAND U4103 ( .A(n4637), .B(sreg[1100]), .Z(n2967) );
  XOR U4104 ( .A(sreg[1100]), .B(n4637), .Z(n2968) );
  NAND U4105 ( .A(n2968), .B(n4636), .Z(n2969) );
  NAND U4106 ( .A(n2967), .B(n2969), .Z(n4645) );
  XOR U4107 ( .A(n4661), .B(sreg[1103]), .Z(n2970) );
  NANDN U4108 ( .A(n4662), .B(n2970), .Z(n2971) );
  NAND U4109 ( .A(n4661), .B(sreg[1103]), .Z(n2972) );
  AND U4110 ( .A(n2971), .B(n2972), .Z(n4668) );
  NAND U4111 ( .A(n4688), .B(sreg[1106]), .Z(n2973) );
  XOR U4112 ( .A(sreg[1106]), .B(n4688), .Z(n2974) );
  NANDN U4113 ( .A(n4687), .B(n2974), .Z(n2975) );
  NAND U4114 ( .A(n2973), .B(n2975), .Z(n4696) );
  XOR U4115 ( .A(n4712), .B(sreg[1109]), .Z(n2976) );
  NANDN U4116 ( .A(n4713), .B(n2976), .Z(n2977) );
  NAND U4117 ( .A(n4712), .B(sreg[1109]), .Z(n2978) );
  AND U4118 ( .A(n2977), .B(n2978), .Z(n4719) );
  NAND U4119 ( .A(n4736), .B(sreg[1112]), .Z(n2979) );
  XOR U4120 ( .A(sreg[1112]), .B(n4736), .Z(n2980) );
  NANDN U4121 ( .A(n4735), .B(n2980), .Z(n2981) );
  NAND U4122 ( .A(n2979), .B(n2981), .Z(n4744) );
  XOR U4123 ( .A(n4760), .B(sreg[1115]), .Z(n2982) );
  NANDN U4124 ( .A(n4761), .B(n2982), .Z(n2983) );
  NAND U4125 ( .A(n4760), .B(sreg[1115]), .Z(n2984) );
  AND U4126 ( .A(n2983), .B(n2984), .Z(n4767) );
  NAND U4127 ( .A(n4784), .B(sreg[1118]), .Z(n2985) );
  XOR U4128 ( .A(sreg[1118]), .B(n4784), .Z(n2986) );
  NANDN U4129 ( .A(n4783), .B(n2986), .Z(n2987) );
  NAND U4130 ( .A(n2985), .B(n2987), .Z(n4792) );
  NAND U4131 ( .A(n4811), .B(sreg[1121]), .Z(n2988) );
  XOR U4132 ( .A(sreg[1121]), .B(n4811), .Z(n2989) );
  NANDN U4133 ( .A(n4812), .B(n2989), .Z(n2990) );
  NAND U4134 ( .A(n2988), .B(n2990), .Z(n4820) );
  NAND U4135 ( .A(n4837), .B(sreg[1124]), .Z(n2991) );
  XOR U4136 ( .A(sreg[1124]), .B(n4837), .Z(n2992) );
  NANDN U4137 ( .A(n4836), .B(n2992), .Z(n2993) );
  NAND U4138 ( .A(n2991), .B(n2993), .Z(n4845) );
  XOR U4139 ( .A(n4861), .B(sreg[1127]), .Z(n2994) );
  NANDN U4140 ( .A(n4862), .B(n2994), .Z(n2995) );
  NAND U4141 ( .A(n4861), .B(sreg[1127]), .Z(n2996) );
  AND U4142 ( .A(n2995), .B(n2996), .Z(n4868) );
  XOR U4143 ( .A(n4886), .B(sreg[1130]), .Z(n2997) );
  NANDN U4144 ( .A(n4887), .B(n2997), .Z(n2998) );
  NAND U4145 ( .A(n4886), .B(sreg[1130]), .Z(n2999) );
  AND U4146 ( .A(n2998), .B(n2999), .Z(n4893) );
  NAND U4147 ( .A(n4908), .B(sreg[1133]), .Z(n3000) );
  XOR U4148 ( .A(sreg[1133]), .B(n4908), .Z(n3001) );
  NAND U4149 ( .A(n3001), .B(n4907), .Z(n3002) );
  NAND U4150 ( .A(n3000), .B(n3002), .Z(n4917) );
  NAND U4151 ( .A(n4935), .B(sreg[1136]), .Z(n3003) );
  XOR U4152 ( .A(sreg[1136]), .B(n4935), .Z(n3004) );
  NANDN U4153 ( .A(n4936), .B(n3004), .Z(n3005) );
  NAND U4154 ( .A(n3003), .B(n3005), .Z(n4944) );
  XOR U4155 ( .A(n4962), .B(sreg[1139]), .Z(n3006) );
  NANDN U4156 ( .A(n4963), .B(n3006), .Z(n3007) );
  NAND U4157 ( .A(n4962), .B(sreg[1139]), .Z(n3008) );
  AND U4158 ( .A(n3007), .B(n3008), .Z(n4969) );
  NAND U4159 ( .A(n4986), .B(sreg[1142]), .Z(n3009) );
  XOR U4160 ( .A(sreg[1142]), .B(n4986), .Z(n3010) );
  NANDN U4161 ( .A(n4985), .B(n3010), .Z(n3011) );
  NAND U4162 ( .A(n3009), .B(n3011), .Z(n4994) );
  NAND U4163 ( .A(n5010), .B(sreg[1145]), .Z(n3012) );
  XOR U4164 ( .A(sreg[1145]), .B(n5010), .Z(n3013) );
  NANDN U4165 ( .A(n5011), .B(n3013), .Z(n3014) );
  NAND U4166 ( .A(n3012), .B(n3014), .Z(n5019) );
  NAND U4167 ( .A(n5036), .B(sreg[1148]), .Z(n3015) );
  XOR U4168 ( .A(sreg[1148]), .B(n5036), .Z(n3016) );
  NANDN U4169 ( .A(n5035), .B(n3016), .Z(n3017) );
  NAND U4170 ( .A(n3015), .B(n3017), .Z(n5044) );
  XOR U4171 ( .A(n5060), .B(sreg[1151]), .Z(n3018) );
  NANDN U4172 ( .A(n5061), .B(n3018), .Z(n3019) );
  NAND U4173 ( .A(n5060), .B(sreg[1151]), .Z(n3020) );
  AND U4174 ( .A(n3019), .B(n3020), .Z(n5067) );
  NAND U4175 ( .A(n5087), .B(sreg[1154]), .Z(n3021) );
  XOR U4176 ( .A(sreg[1154]), .B(n5087), .Z(n3022) );
  NANDN U4177 ( .A(n5086), .B(n3022), .Z(n3023) );
  NAND U4178 ( .A(n3021), .B(n3023), .Z(n5095) );
  NAND U4179 ( .A(n5113), .B(sreg[1157]), .Z(n3024) );
  XOR U4180 ( .A(sreg[1157]), .B(n5113), .Z(n3025) );
  NANDN U4181 ( .A(n5114), .B(n3025), .Z(n3026) );
  NAND U4182 ( .A(n3024), .B(n3026), .Z(n5122) );
  NAND U4183 ( .A(n5139), .B(sreg[1160]), .Z(n3027) );
  XOR U4184 ( .A(sreg[1160]), .B(n5139), .Z(n3028) );
  NANDN U4185 ( .A(n5138), .B(n3028), .Z(n3029) );
  NAND U4186 ( .A(n3027), .B(n3029), .Z(n5147) );
  NAND U4187 ( .A(n5163), .B(sreg[1163]), .Z(n3030) );
  XOR U4188 ( .A(sreg[1163]), .B(n5163), .Z(n3031) );
  NANDN U4189 ( .A(n5164), .B(n3031), .Z(n3032) );
  NAND U4190 ( .A(n3030), .B(n3032), .Z(n5172) );
  NAND U4191 ( .A(n5189), .B(sreg[1166]), .Z(n3033) );
  XOR U4192 ( .A(sreg[1166]), .B(n5189), .Z(n3034) );
  NANDN U4193 ( .A(n5188), .B(n3034), .Z(n3035) );
  NAND U4194 ( .A(n3033), .B(n3035), .Z(n5197) );
  XOR U4195 ( .A(n5213), .B(sreg[1169]), .Z(n3036) );
  NANDN U4196 ( .A(n5214), .B(n3036), .Z(n3037) );
  NAND U4197 ( .A(n5213), .B(sreg[1169]), .Z(n3038) );
  AND U4198 ( .A(n3037), .B(n3038), .Z(n5220) );
  NAND U4199 ( .A(n5238), .B(sreg[1172]), .Z(n3039) );
  XOR U4200 ( .A(sreg[1172]), .B(n5238), .Z(n3040) );
  NAND U4201 ( .A(n3040), .B(n5237), .Z(n3041) );
  NAND U4202 ( .A(n3039), .B(n3041), .Z(n5246) );
  XOR U4203 ( .A(n5262), .B(sreg[1175]), .Z(n3042) );
  NANDN U4204 ( .A(n5263), .B(n3042), .Z(n3043) );
  NAND U4205 ( .A(n5262), .B(sreg[1175]), .Z(n3044) );
  AND U4206 ( .A(n3043), .B(n3044), .Z(n5269) );
  NAND U4207 ( .A(n5286), .B(sreg[1178]), .Z(n3045) );
  XOR U4208 ( .A(sreg[1178]), .B(n5286), .Z(n3046) );
  NANDN U4209 ( .A(n5285), .B(n3046), .Z(n3047) );
  NAND U4210 ( .A(n3045), .B(n3047), .Z(n5294) );
  XOR U4211 ( .A(n5310), .B(sreg[1181]), .Z(n3048) );
  NANDN U4212 ( .A(n5311), .B(n3048), .Z(n3049) );
  NAND U4213 ( .A(n5310), .B(sreg[1181]), .Z(n3050) );
  AND U4214 ( .A(n3049), .B(n3050), .Z(n5317) );
  NAND U4215 ( .A(n5334), .B(sreg[1184]), .Z(n3051) );
  XOR U4216 ( .A(sreg[1184]), .B(n5334), .Z(n3052) );
  NANDN U4217 ( .A(n5333), .B(n3052), .Z(n3053) );
  NAND U4218 ( .A(n3051), .B(n3053), .Z(n5342) );
  XOR U4219 ( .A(n5361), .B(sreg[1187]), .Z(n3054) );
  NANDN U4220 ( .A(n5362), .B(n3054), .Z(n3055) );
  NAND U4221 ( .A(n5361), .B(sreg[1187]), .Z(n3056) );
  AND U4222 ( .A(n3055), .B(n3056), .Z(n5368) );
  NAND U4223 ( .A(n5385), .B(sreg[1190]), .Z(n3057) );
  XOR U4224 ( .A(sreg[1190]), .B(n5385), .Z(n3058) );
  NANDN U4225 ( .A(n5384), .B(n3058), .Z(n3059) );
  NAND U4226 ( .A(n3057), .B(n3059), .Z(n5391) );
  NAND U4227 ( .A(n5406), .B(sreg[1193]), .Z(n3060) );
  XOR U4228 ( .A(sreg[1193]), .B(n5406), .Z(n3061) );
  NAND U4229 ( .A(n3061), .B(n5405), .Z(n3062) );
  NAND U4230 ( .A(n3060), .B(n3062), .Z(n5412) );
  NAND U4231 ( .A(n5432), .B(sreg[1196]), .Z(n3063) );
  XOR U4232 ( .A(sreg[1196]), .B(n5432), .Z(n3064) );
  NANDN U4233 ( .A(n5431), .B(n3064), .Z(n3065) );
  NAND U4234 ( .A(n3063), .B(n3065), .Z(n5440) );
  XOR U4235 ( .A(n5458), .B(sreg[1199]), .Z(n3066) );
  NANDN U4236 ( .A(n5459), .B(n3066), .Z(n3067) );
  NAND U4237 ( .A(n5458), .B(sreg[1199]), .Z(n3068) );
  AND U4238 ( .A(n3067), .B(n3068), .Z(n5465) );
  NAND U4239 ( .A(n5482), .B(sreg[1202]), .Z(n3069) );
  XOR U4240 ( .A(sreg[1202]), .B(n5482), .Z(n3070) );
  NANDN U4241 ( .A(n5481), .B(n3070), .Z(n3071) );
  NAND U4242 ( .A(n3069), .B(n3071), .Z(n5490) );
  XOR U4243 ( .A(n5506), .B(sreg[1205]), .Z(n3072) );
  NANDN U4244 ( .A(n5507), .B(n3072), .Z(n3073) );
  NAND U4245 ( .A(n5506), .B(sreg[1205]), .Z(n3074) );
  AND U4246 ( .A(n3073), .B(n3074), .Z(n5513) );
  NAND U4247 ( .A(n5530), .B(sreg[1208]), .Z(n3075) );
  XOR U4248 ( .A(sreg[1208]), .B(n5530), .Z(n3076) );
  NANDN U4249 ( .A(n5529), .B(n3076), .Z(n3077) );
  NAND U4250 ( .A(n3075), .B(n3077), .Z(n5538) );
  XOR U4251 ( .A(n5556), .B(sreg[1211]), .Z(n3078) );
  NANDN U4252 ( .A(n5557), .B(n3078), .Z(n3079) );
  NAND U4253 ( .A(n5556), .B(sreg[1211]), .Z(n3080) );
  AND U4254 ( .A(n3079), .B(n3080), .Z(n5563) );
  NAND U4255 ( .A(n5583), .B(sreg[1214]), .Z(n3081) );
  XOR U4256 ( .A(sreg[1214]), .B(n5583), .Z(n3082) );
  NANDN U4257 ( .A(n5582), .B(n3082), .Z(n3083) );
  NAND U4258 ( .A(n3081), .B(n3083), .Z(n5591) );
  XOR U4259 ( .A(n5607), .B(sreg[1217]), .Z(n3084) );
  NANDN U4260 ( .A(n5608), .B(n3084), .Z(n3085) );
  NAND U4261 ( .A(n5607), .B(sreg[1217]), .Z(n3086) );
  AND U4262 ( .A(n3085), .B(n3086), .Z(n5614) );
  NAND U4263 ( .A(n5631), .B(sreg[1220]), .Z(n3087) );
  XOR U4264 ( .A(sreg[1220]), .B(n5631), .Z(n3088) );
  NANDN U4265 ( .A(n5630), .B(n3088), .Z(n3089) );
  NAND U4266 ( .A(n3087), .B(n3089), .Z(n5639) );
  NAND U4267 ( .A(n5654), .B(sreg[1223]), .Z(n3090) );
  XOR U4268 ( .A(sreg[1223]), .B(n5654), .Z(n3091) );
  NAND U4269 ( .A(n3091), .B(n5653), .Z(n3092) );
  NAND U4270 ( .A(n3090), .B(n3092), .Z(n5660) );
  NAND U4271 ( .A(n5680), .B(sreg[1226]), .Z(n3093) );
  XOR U4272 ( .A(sreg[1226]), .B(n5680), .Z(n3094) );
  NANDN U4273 ( .A(n5679), .B(n3094), .Z(n3095) );
  NAND U4274 ( .A(n3093), .B(n3095), .Z(n5688) );
  XOR U4275 ( .A(n5704), .B(sreg[1229]), .Z(n3096) );
  NANDN U4276 ( .A(n5705), .B(n3096), .Z(n3097) );
  NAND U4277 ( .A(n5704), .B(sreg[1229]), .Z(n3098) );
  AND U4278 ( .A(n3097), .B(n3098), .Z(n5711) );
  NAND U4279 ( .A(n5728), .B(sreg[1232]), .Z(n3099) );
  XOR U4280 ( .A(sreg[1232]), .B(n5728), .Z(n3100) );
  NANDN U4281 ( .A(n5727), .B(n3100), .Z(n3101) );
  NAND U4282 ( .A(n3099), .B(n3101), .Z(n5736) );
  NAND U4283 ( .A(n5752), .B(sreg[1235]), .Z(n3102) );
  XOR U4284 ( .A(sreg[1235]), .B(n5752), .Z(n3103) );
  NANDN U4285 ( .A(n5753), .B(n3103), .Z(n3104) );
  NAND U4286 ( .A(n3102), .B(n3104), .Z(n5761) );
  NAND U4287 ( .A(n5778), .B(sreg[1238]), .Z(n3105) );
  XOR U4288 ( .A(sreg[1238]), .B(n5778), .Z(n3106) );
  NANDN U4289 ( .A(n5777), .B(n3106), .Z(n3107) );
  NAND U4290 ( .A(n3105), .B(n3107), .Z(n5786) );
  NAND U4291 ( .A(n5802), .B(sreg[1241]), .Z(n3108) );
  XOR U4292 ( .A(sreg[1241]), .B(n5802), .Z(n3109) );
  NANDN U4293 ( .A(n5803), .B(n3109), .Z(n3110) );
  NAND U4294 ( .A(n3108), .B(n3110), .Z(n5811) );
  NAND U4295 ( .A(n5831), .B(sreg[1244]), .Z(n3111) );
  XOR U4296 ( .A(sreg[1244]), .B(n5831), .Z(n3112) );
  NANDN U4297 ( .A(n5830), .B(n3112), .Z(n3113) );
  NAND U4298 ( .A(n3111), .B(n3113), .Z(n5839) );
  XOR U4299 ( .A(n5855), .B(sreg[1247]), .Z(n3114) );
  NANDN U4300 ( .A(n5856), .B(n3114), .Z(n3115) );
  NAND U4301 ( .A(n5855), .B(sreg[1247]), .Z(n3116) );
  AND U4302 ( .A(n3115), .B(n3116), .Z(n5862) );
  NAND U4303 ( .A(n5879), .B(sreg[1250]), .Z(n3117) );
  XOR U4304 ( .A(sreg[1250]), .B(n5879), .Z(n3118) );
  NANDN U4305 ( .A(n5878), .B(n3118), .Z(n3119) );
  NAND U4306 ( .A(n3117), .B(n3119), .Z(n5887) );
  XOR U4307 ( .A(n5903), .B(sreg[1253]), .Z(n3120) );
  NANDN U4308 ( .A(n5904), .B(n3120), .Z(n3121) );
  NAND U4309 ( .A(n5903), .B(sreg[1253]), .Z(n3122) );
  AND U4310 ( .A(n3121), .B(n3122), .Z(n5910) );
  NAND U4311 ( .A(n5928), .B(sreg[1256]), .Z(n3123) );
  XOR U4312 ( .A(sreg[1256]), .B(n5928), .Z(n3124) );
  NANDN U4313 ( .A(n5929), .B(n3124), .Z(n3125) );
  NAND U4314 ( .A(n3123), .B(n3125), .Z(n5937) );
  XOR U4315 ( .A(n5953), .B(sreg[1259]), .Z(n3126) );
  NANDN U4316 ( .A(n5954), .B(n3126), .Z(n3127) );
  NAND U4317 ( .A(n5953), .B(sreg[1259]), .Z(n3128) );
  AND U4318 ( .A(n3127), .B(n3128), .Z(n5963) );
  NAND U4319 ( .A(n5978), .B(sreg[1262]), .Z(n3129) );
  XOR U4320 ( .A(sreg[1262]), .B(n5978), .Z(n3130) );
  NAND U4321 ( .A(n3130), .B(n5977), .Z(n3131) );
  NAND U4322 ( .A(n3129), .B(n3131), .Z(n5986) );
  XOR U4323 ( .A(n6002), .B(sreg[1265]), .Z(n3132) );
  NANDN U4324 ( .A(n6003), .B(n3132), .Z(n3133) );
  NAND U4325 ( .A(n6002), .B(sreg[1265]), .Z(n3134) );
  AND U4326 ( .A(n3133), .B(n3134), .Z(n6009) );
  NAND U4327 ( .A(n6026), .B(sreg[1268]), .Z(n3135) );
  XOR U4328 ( .A(sreg[1268]), .B(n6026), .Z(n3136) );
  NANDN U4329 ( .A(n6025), .B(n3136), .Z(n3137) );
  NAND U4330 ( .A(n3135), .B(n3137), .Z(n6034) );
  XOR U4331 ( .A(n6050), .B(sreg[1271]), .Z(n3138) );
  NANDN U4332 ( .A(n6051), .B(n3138), .Z(n3139) );
  NAND U4333 ( .A(n6050), .B(sreg[1271]), .Z(n3140) );
  AND U4334 ( .A(n3139), .B(n3140), .Z(n6060) );
  NAND U4335 ( .A(n6077), .B(sreg[1274]), .Z(n3141) );
  XOR U4336 ( .A(sreg[1274]), .B(n6077), .Z(n3142) );
  NANDN U4337 ( .A(n6076), .B(n3142), .Z(n3143) );
  NAND U4338 ( .A(n3141), .B(n3143), .Z(n6085) );
  XOR U4339 ( .A(n6101), .B(sreg[1277]), .Z(n3144) );
  NANDN U4340 ( .A(n6102), .B(n3144), .Z(n3145) );
  NAND U4341 ( .A(n6101), .B(sreg[1277]), .Z(n3146) );
  AND U4342 ( .A(n3145), .B(n3146), .Z(n6108) );
  NAND U4343 ( .A(n6125), .B(sreg[1280]), .Z(n3147) );
  XOR U4344 ( .A(sreg[1280]), .B(n6125), .Z(n3148) );
  NANDN U4345 ( .A(n6124), .B(n3148), .Z(n3149) );
  NAND U4346 ( .A(n3147), .B(n3149), .Z(n6131) );
  XOR U4347 ( .A(n6147), .B(sreg[1283]), .Z(n3150) );
  NANDN U4348 ( .A(n6148), .B(n3150), .Z(n3151) );
  NAND U4349 ( .A(n6147), .B(sreg[1283]), .Z(n3152) );
  AND U4350 ( .A(n3151), .B(n3152), .Z(n6157) );
  NAND U4351 ( .A(n6172), .B(sreg[1286]), .Z(n3153) );
  XOR U4352 ( .A(sreg[1286]), .B(n6172), .Z(n3154) );
  NAND U4353 ( .A(n3154), .B(n6171), .Z(n3155) );
  NAND U4354 ( .A(n3153), .B(n3155), .Z(n6180) );
  XOR U4355 ( .A(n6198), .B(sreg[1289]), .Z(n3156) );
  NANDN U4356 ( .A(n6199), .B(n3156), .Z(n3157) );
  NAND U4357 ( .A(n6198), .B(sreg[1289]), .Z(n3158) );
  AND U4358 ( .A(n3157), .B(n3158), .Z(n6205) );
  NAND U4359 ( .A(n6220), .B(sreg[1292]), .Z(n3159) );
  XOR U4360 ( .A(sreg[1292]), .B(n6220), .Z(n3160) );
  NAND U4361 ( .A(n3160), .B(n6219), .Z(n3161) );
  NAND U4362 ( .A(n3159), .B(n3161), .Z(n6228) );
  XOR U4363 ( .A(n6244), .B(sreg[1295]), .Z(n3162) );
  NANDN U4364 ( .A(n6245), .B(n3162), .Z(n3163) );
  NAND U4365 ( .A(n6244), .B(sreg[1295]), .Z(n3164) );
  AND U4366 ( .A(n3163), .B(n3164), .Z(n6254) );
  NAND U4367 ( .A(n6272), .B(sreg[1298]), .Z(n3165) );
  XOR U4368 ( .A(sreg[1298]), .B(n6272), .Z(n3166) );
  NANDN U4369 ( .A(n6273), .B(n3166), .Z(n3167) );
  NAND U4370 ( .A(n3165), .B(n3167), .Z(n6281) );
  XOR U4371 ( .A(n6297), .B(sreg[1301]), .Z(n3168) );
  NANDN U4372 ( .A(n6298), .B(n3168), .Z(n3169) );
  NAND U4373 ( .A(n6297), .B(sreg[1301]), .Z(n3170) );
  AND U4374 ( .A(n3169), .B(n3170), .Z(n6304) );
  NAND U4375 ( .A(n6321), .B(sreg[1304]), .Z(n3171) );
  XOR U4376 ( .A(sreg[1304]), .B(n6321), .Z(n3172) );
  NANDN U4377 ( .A(n6320), .B(n3172), .Z(n3173) );
  NAND U4378 ( .A(n3171), .B(n3173), .Z(n6329) );
  NAND U4379 ( .A(n6345), .B(sreg[1307]), .Z(n3174) );
  XOR U4380 ( .A(sreg[1307]), .B(n6345), .Z(n3175) );
  NANDN U4381 ( .A(n6346), .B(n3175), .Z(n3176) );
  NAND U4382 ( .A(n3174), .B(n3176), .Z(n6354) );
  NAND U4383 ( .A(n6371), .B(sreg[1310]), .Z(n3177) );
  XOR U4384 ( .A(sreg[1310]), .B(n6371), .Z(n3178) );
  NANDN U4385 ( .A(n6370), .B(n3178), .Z(n3179) );
  NAND U4386 ( .A(n3177), .B(n3179), .Z(n6379) );
  NAND U4387 ( .A(n6395), .B(sreg[1313]), .Z(n3180) );
  XOR U4388 ( .A(sreg[1313]), .B(n6395), .Z(n3181) );
  NANDN U4389 ( .A(n6396), .B(n3181), .Z(n3182) );
  NAND U4390 ( .A(n3180), .B(n3182), .Z(n6404) );
  NAND U4391 ( .A(n6424), .B(sreg[1316]), .Z(n3183) );
  XOR U4392 ( .A(sreg[1316]), .B(n6424), .Z(n3184) );
  NANDN U4393 ( .A(n6423), .B(n3184), .Z(n3185) );
  NAND U4394 ( .A(n3183), .B(n3185), .Z(n6432) );
  XOR U4395 ( .A(n6448), .B(sreg[1319]), .Z(n3186) );
  NANDN U4396 ( .A(n6449), .B(n3186), .Z(n3187) );
  NAND U4397 ( .A(n6448), .B(sreg[1319]), .Z(n3188) );
  AND U4398 ( .A(n3187), .B(n3188), .Z(n6455) );
  NAND U4399 ( .A(n6472), .B(sreg[1322]), .Z(n3189) );
  XOR U4400 ( .A(sreg[1322]), .B(n6472), .Z(n3190) );
  NANDN U4401 ( .A(n6471), .B(n3190), .Z(n3191) );
  NAND U4402 ( .A(n3189), .B(n3191), .Z(n6480) );
  XOR U4403 ( .A(n6496), .B(sreg[1325]), .Z(n3192) );
  NANDN U4404 ( .A(n6497), .B(n3192), .Z(n3193) );
  NAND U4405 ( .A(n6496), .B(sreg[1325]), .Z(n3194) );
  AND U4406 ( .A(n3193), .B(n3194), .Z(n6503) );
  NAND U4407 ( .A(n6520), .B(sreg[1328]), .Z(n3195) );
  XOR U4408 ( .A(sreg[1328]), .B(n6520), .Z(n3196) );
  NANDN U4409 ( .A(n6519), .B(n3196), .Z(n3197) );
  NAND U4410 ( .A(n3195), .B(n3197), .Z(n6528) );
  XOR U4411 ( .A(n6547), .B(sreg[1331]), .Z(n3198) );
  NANDN U4412 ( .A(n6548), .B(n3198), .Z(n3199) );
  NAND U4413 ( .A(n6547), .B(sreg[1331]), .Z(n3200) );
  AND U4414 ( .A(n3199), .B(n3200), .Z(n6554) );
  NAND U4415 ( .A(n6571), .B(sreg[1334]), .Z(n3201) );
  XOR U4416 ( .A(sreg[1334]), .B(n6571), .Z(n3202) );
  NANDN U4417 ( .A(n6570), .B(n3202), .Z(n3203) );
  NAND U4418 ( .A(n3201), .B(n3203), .Z(n6579) );
  XOR U4419 ( .A(n6595), .B(sreg[1337]), .Z(n3204) );
  NANDN U4420 ( .A(n6596), .B(n3204), .Z(n3205) );
  NAND U4421 ( .A(n6595), .B(sreg[1337]), .Z(n3206) );
  AND U4422 ( .A(n3205), .B(n3206), .Z(n6602) );
  NAND U4423 ( .A(n6619), .B(sreg[1340]), .Z(n3207) );
  XOR U4424 ( .A(sreg[1340]), .B(n6619), .Z(n3208) );
  NANDN U4425 ( .A(n6618), .B(n3208), .Z(n3209) );
  NAND U4426 ( .A(n3207), .B(n3209), .Z(n6627) );
  XOR U4427 ( .A(n6643), .B(sreg[1343]), .Z(n3210) );
  NANDN U4428 ( .A(n6644), .B(n3210), .Z(n3211) );
  NAND U4429 ( .A(n6643), .B(sreg[1343]), .Z(n3212) );
  AND U4430 ( .A(n3211), .B(n3212), .Z(n6653) );
  NAND U4431 ( .A(n6670), .B(sreg[1346]), .Z(n3213) );
  XOR U4432 ( .A(sreg[1346]), .B(n6670), .Z(n3214) );
  NANDN U4433 ( .A(n6669), .B(n3214), .Z(n3215) );
  NAND U4434 ( .A(n3213), .B(n3215), .Z(n6678) );
  XOR U4435 ( .A(n6696), .B(sreg[1349]), .Z(n3216) );
  NANDN U4436 ( .A(n6697), .B(n3216), .Z(n3217) );
  NAND U4437 ( .A(n6696), .B(sreg[1349]), .Z(n3218) );
  AND U4438 ( .A(n3217), .B(n3218), .Z(n6703) );
  NAND U4439 ( .A(n6718), .B(sreg[1352]), .Z(n3219) );
  XOR U4440 ( .A(sreg[1352]), .B(n6718), .Z(n3220) );
  NAND U4441 ( .A(n3220), .B(n6717), .Z(n3221) );
  NAND U4442 ( .A(n3219), .B(n3221), .Z(n6726) );
  NAND U4443 ( .A(n6741), .B(sreg[1355]), .Z(n3222) );
  XOR U4444 ( .A(sreg[1355]), .B(n6741), .Z(n3223) );
  NAND U4445 ( .A(n3223), .B(n6740), .Z(n3224) );
  NAND U4446 ( .A(n3222), .B(n3224), .Z(n6750) );
  NAND U4447 ( .A(n6767), .B(sreg[1358]), .Z(n3225) );
  XOR U4448 ( .A(sreg[1358]), .B(n6767), .Z(n3226) );
  NANDN U4449 ( .A(n6766), .B(n3226), .Z(n3227) );
  NAND U4450 ( .A(n3225), .B(n3227), .Z(n6775) );
  NAND U4451 ( .A(n6791), .B(sreg[1361]), .Z(n3228) );
  XOR U4452 ( .A(sreg[1361]), .B(n6791), .Z(n3229) );
  NANDN U4453 ( .A(n6792), .B(n3229), .Z(n3230) );
  NAND U4454 ( .A(n3228), .B(n3230), .Z(n6800) );
  NAND U4455 ( .A(n6817), .B(sreg[1364]), .Z(n3231) );
  XOR U4456 ( .A(sreg[1364]), .B(n6817), .Z(n3232) );
  NANDN U4457 ( .A(n6816), .B(n3232), .Z(n3233) );
  NAND U4458 ( .A(n3231), .B(n3233), .Z(n6825) );
  XOR U4459 ( .A(n6843), .B(sreg[1367]), .Z(n3234) );
  NANDN U4460 ( .A(n6844), .B(n3234), .Z(n3235) );
  NAND U4461 ( .A(n6843), .B(sreg[1367]), .Z(n3236) );
  AND U4462 ( .A(n3235), .B(n3236), .Z(n6850) );
  NAND U4463 ( .A(n6867), .B(sreg[1370]), .Z(n3237) );
  XOR U4464 ( .A(sreg[1370]), .B(n6867), .Z(n3238) );
  NANDN U4465 ( .A(n6866), .B(n3238), .Z(n3239) );
  NAND U4466 ( .A(n3237), .B(n3239), .Z(n6875) );
  XOR U4467 ( .A(n6893), .B(sreg[1373]), .Z(n3240) );
  NANDN U4468 ( .A(n6894), .B(n3240), .Z(n3241) );
  NAND U4469 ( .A(n6893), .B(sreg[1373]), .Z(n3242) );
  AND U4470 ( .A(n3241), .B(n3242), .Z(n6900) );
  NAND U4471 ( .A(n6920), .B(sreg[1376]), .Z(n3243) );
  XOR U4472 ( .A(sreg[1376]), .B(n6920), .Z(n3244) );
  NANDN U4473 ( .A(n6919), .B(n3244), .Z(n3245) );
  NAND U4474 ( .A(n3243), .B(n3245), .Z(n6928) );
  XOR U4475 ( .A(n6944), .B(sreg[1379]), .Z(n3246) );
  NANDN U4476 ( .A(n6945), .B(n3246), .Z(n3247) );
  NAND U4477 ( .A(n6944), .B(sreg[1379]), .Z(n3248) );
  AND U4478 ( .A(n3247), .B(n3248), .Z(n6951) );
  NAND U4479 ( .A(n6968), .B(sreg[1382]), .Z(n3249) );
  XOR U4480 ( .A(sreg[1382]), .B(n6968), .Z(n3250) );
  NANDN U4481 ( .A(n6967), .B(n3250), .Z(n3251) );
  NAND U4482 ( .A(n3249), .B(n3251), .Z(n6974) );
  XOR U4483 ( .A(n6990), .B(sreg[1385]), .Z(n3252) );
  NANDN U4484 ( .A(n6991), .B(n3252), .Z(n3253) );
  NAND U4485 ( .A(n6990), .B(sreg[1385]), .Z(n3254) );
  AND U4486 ( .A(n3253), .B(n3254), .Z(n6997) );
  NAND U4487 ( .A(n7015), .B(sreg[1388]), .Z(n3255) );
  XOR U4488 ( .A(sreg[1388]), .B(n7015), .Z(n3256) );
  NAND U4489 ( .A(n3256), .B(n7014), .Z(n3257) );
  NAND U4490 ( .A(n3255), .B(n3257), .Z(n7023) );
  XOR U4491 ( .A(n7039), .B(sreg[1391]), .Z(n3258) );
  NANDN U4492 ( .A(n7040), .B(n3258), .Z(n3259) );
  NAND U4493 ( .A(n7039), .B(sreg[1391]), .Z(n3260) );
  AND U4494 ( .A(n3259), .B(n3260), .Z(n7046) );
  NAND U4495 ( .A(n7063), .B(sreg[1394]), .Z(n3261) );
  XOR U4496 ( .A(sreg[1394]), .B(n7063), .Z(n3262) );
  NANDN U4497 ( .A(n7062), .B(n3262), .Z(n3263) );
  NAND U4498 ( .A(n3261), .B(n3263), .Z(n7069) );
  XOR U4499 ( .A(n7085), .B(sreg[1397]), .Z(n3264) );
  NANDN U4500 ( .A(n7086), .B(n3264), .Z(n3265) );
  NAND U4501 ( .A(n7085), .B(sreg[1397]), .Z(n3266) );
  AND U4502 ( .A(n3265), .B(n3266), .Z(n7095) );
  NAND U4503 ( .A(n7112), .B(sreg[1400]), .Z(n3267) );
  XOR U4504 ( .A(sreg[1400]), .B(n7112), .Z(n3268) );
  NANDN U4505 ( .A(n7111), .B(n3268), .Z(n3269) );
  NAND U4506 ( .A(n3267), .B(n3269), .Z(n7118) );
  XOR U4507 ( .A(n7134), .B(sreg[1403]), .Z(n3270) );
  NANDN U4508 ( .A(n7135), .B(n3270), .Z(n3271) );
  NAND U4509 ( .A(n7134), .B(sreg[1403]), .Z(n3272) );
  AND U4510 ( .A(n3271), .B(n3272), .Z(n7141) );
  NAND U4511 ( .A(n7158), .B(sreg[1406]), .Z(n3273) );
  XOR U4512 ( .A(sreg[1406]), .B(n7158), .Z(n3274) );
  NANDN U4513 ( .A(n7157), .B(n3274), .Z(n3275) );
  NAND U4514 ( .A(n3273), .B(n3275), .Z(n7166) );
  XOR U4515 ( .A(n7182), .B(sreg[1409]), .Z(n3276) );
  NANDN U4516 ( .A(n7183), .B(n3276), .Z(n3277) );
  NAND U4517 ( .A(n7182), .B(sreg[1409]), .Z(n3278) );
  AND U4518 ( .A(n3277), .B(n3278), .Z(n7192) );
  NAND U4519 ( .A(n7209), .B(sreg[1412]), .Z(n3279) );
  XOR U4520 ( .A(sreg[1412]), .B(n7209), .Z(n3280) );
  NANDN U4521 ( .A(n7208), .B(n3280), .Z(n3281) );
  NAND U4522 ( .A(n3279), .B(n3281), .Z(n7217) );
  XOR U4523 ( .A(n7233), .B(sreg[1415]), .Z(n3282) );
  NANDN U4524 ( .A(n7234), .B(n3282), .Z(n3283) );
  NAND U4525 ( .A(n7233), .B(sreg[1415]), .Z(n3284) );
  AND U4526 ( .A(n3283), .B(n3284), .Z(n7240) );
  NAND U4527 ( .A(n7257), .B(sreg[1418]), .Z(n3285) );
  XOR U4528 ( .A(sreg[1418]), .B(n7257), .Z(n3286) );
  NANDN U4529 ( .A(n7256), .B(n3286), .Z(n3287) );
  NAND U4530 ( .A(n3285), .B(n3287), .Z(n7265) );
  XOR U4531 ( .A(n7281), .B(sreg[1421]), .Z(n3288) );
  NANDN U4532 ( .A(n7282), .B(n3288), .Z(n3289) );
  NAND U4533 ( .A(n7281), .B(sreg[1421]), .Z(n3290) );
  AND U4534 ( .A(n3289), .B(n3290), .Z(n7288) );
  NAND U4535 ( .A(n7308), .B(sreg[1424]), .Z(n3291) );
  XOR U4536 ( .A(sreg[1424]), .B(n7308), .Z(n3292) );
  NANDN U4537 ( .A(n7307), .B(n3292), .Z(n3293) );
  NAND U4538 ( .A(n3291), .B(n3293), .Z(n7316) );
  NAND U4539 ( .A(n7332), .B(sreg[1427]), .Z(n3294) );
  XOR U4540 ( .A(sreg[1427]), .B(n7332), .Z(n3295) );
  NANDN U4541 ( .A(n7333), .B(n3295), .Z(n3296) );
  NAND U4542 ( .A(n3294), .B(n3296), .Z(n7341) );
  NAND U4543 ( .A(n7358), .B(sreg[1430]), .Z(n3297) );
  XOR U4544 ( .A(sreg[1430]), .B(n7358), .Z(n3298) );
  NANDN U4545 ( .A(n7357), .B(n3298), .Z(n3299) );
  NAND U4546 ( .A(n3297), .B(n3299), .Z(n7366) );
  NAND U4547 ( .A(n7381), .B(sreg[1433]), .Z(n3300) );
  XOR U4548 ( .A(sreg[1433]), .B(n7381), .Z(n3301) );
  NAND U4549 ( .A(n3301), .B(n7380), .Z(n3302) );
  NAND U4550 ( .A(n3300), .B(n3302), .Z(n7389) );
  NAND U4551 ( .A(n7406), .B(sreg[1436]), .Z(n3303) );
  XOR U4552 ( .A(sreg[1436]), .B(n7406), .Z(n3304) );
  NANDN U4553 ( .A(n7405), .B(n3304), .Z(n3305) );
  NAND U4554 ( .A(n3303), .B(n3305), .Z(n7414) );
  XOR U4555 ( .A(n7430), .B(sreg[1439]), .Z(n3306) );
  NANDN U4556 ( .A(n7431), .B(n3306), .Z(n3307) );
  NAND U4557 ( .A(n7430), .B(sreg[1439]), .Z(n3308) );
  AND U4558 ( .A(n3307), .B(n3308), .Z(n7440) );
  NAND U4559 ( .A(n7457), .B(sreg[1442]), .Z(n3309) );
  XOR U4560 ( .A(sreg[1442]), .B(n7457), .Z(n3310) );
  NANDN U4561 ( .A(n7456), .B(n3310), .Z(n3311) );
  NAND U4562 ( .A(n3309), .B(n3311), .Z(n7463) );
  XOR U4563 ( .A(n7481), .B(sreg[1445]), .Z(n3312) );
  NANDN U4564 ( .A(n7482), .B(n3312), .Z(n3313) );
  NAND U4565 ( .A(n7481), .B(sreg[1445]), .Z(n3314) );
  AND U4566 ( .A(n3313), .B(n3314), .Z(n7488) );
  NAND U4567 ( .A(n7503), .B(sreg[1448]), .Z(n3315) );
  XOR U4568 ( .A(sreg[1448]), .B(n7503), .Z(n3316) );
  NAND U4569 ( .A(n3316), .B(n7502), .Z(n3317) );
  NAND U4570 ( .A(n3315), .B(n3317), .Z(n7509) );
  XOR U4571 ( .A(n7527), .B(sreg[1451]), .Z(n3318) );
  NANDN U4572 ( .A(n7528), .B(n3318), .Z(n3319) );
  NAND U4573 ( .A(n7527), .B(sreg[1451]), .Z(n3320) );
  AND U4574 ( .A(n3319), .B(n3320), .Z(n7537) );
  NAND U4575 ( .A(n7554), .B(sreg[1454]), .Z(n3321) );
  XOR U4576 ( .A(sreg[1454]), .B(n7554), .Z(n3322) );
  NANDN U4577 ( .A(n7553), .B(n3322), .Z(n3323) );
  NAND U4578 ( .A(n3321), .B(n3323), .Z(n7562) );
  XOR U4579 ( .A(n7580), .B(sreg[1457]), .Z(n3324) );
  NANDN U4580 ( .A(n7581), .B(n3324), .Z(n3325) );
  NAND U4581 ( .A(n7580), .B(sreg[1457]), .Z(n3326) );
  AND U4582 ( .A(n3325), .B(n3326), .Z(n7587) );
  NAND U4583 ( .A(n7602), .B(sreg[1460]), .Z(n3327) );
  XOR U4584 ( .A(sreg[1460]), .B(n7602), .Z(n3328) );
  NAND U4585 ( .A(n3328), .B(n7601), .Z(n3329) );
  NAND U4586 ( .A(n3327), .B(n3329), .Z(n7610) );
  XOR U4587 ( .A(n7626), .B(sreg[1463]), .Z(n3330) );
  NANDN U4588 ( .A(n7627), .B(n3330), .Z(n3331) );
  NAND U4589 ( .A(n7626), .B(sreg[1463]), .Z(n3332) );
  AND U4590 ( .A(n3331), .B(n3332), .Z(n7633) );
  NAND U4591 ( .A(n7653), .B(sreg[1466]), .Z(n3333) );
  XOR U4592 ( .A(sreg[1466]), .B(n7653), .Z(n3334) );
  NANDN U4593 ( .A(n7652), .B(n3334), .Z(n3335) );
  NAND U4594 ( .A(n3333), .B(n3335), .Z(n7661) );
  XOR U4595 ( .A(n7677), .B(sreg[1469]), .Z(n3336) );
  NANDN U4596 ( .A(n7678), .B(n3336), .Z(n3337) );
  NAND U4597 ( .A(n7677), .B(sreg[1469]), .Z(n3338) );
  AND U4598 ( .A(n3337), .B(n3338), .Z(n7684) );
  NAND U4599 ( .A(n7701), .B(sreg[1472]), .Z(n3339) );
  XOR U4600 ( .A(sreg[1472]), .B(n7701), .Z(n3340) );
  NANDN U4601 ( .A(n7700), .B(n3340), .Z(n3341) );
  NAND U4602 ( .A(n3339), .B(n3341), .Z(n7709) );
  NAND U4603 ( .A(n7725), .B(sreg[1475]), .Z(n3342) );
  XOR U4604 ( .A(sreg[1475]), .B(n7725), .Z(n3343) );
  NANDN U4605 ( .A(n7726), .B(n3343), .Z(n3344) );
  NAND U4606 ( .A(n3342), .B(n3344), .Z(n7734) );
  NAND U4607 ( .A(n7751), .B(sreg[1478]), .Z(n3345) );
  XOR U4608 ( .A(sreg[1478]), .B(n7751), .Z(n3346) );
  NANDN U4609 ( .A(n7750), .B(n3346), .Z(n3347) );
  NAND U4610 ( .A(n3345), .B(n3347), .Z(n7759) );
  NAND U4611 ( .A(n7777), .B(sreg[1481]), .Z(n3348) );
  XOR U4612 ( .A(sreg[1481]), .B(n7777), .Z(n3349) );
  NAND U4613 ( .A(n3349), .B(n7776), .Z(n3350) );
  NAND U4614 ( .A(n3348), .B(n3350), .Z(n7785) );
  NAND U4615 ( .A(n7800), .B(sreg[1484]), .Z(n3351) );
  XOR U4616 ( .A(sreg[1484]), .B(n7800), .Z(n3352) );
  NAND U4617 ( .A(n3352), .B(n7799), .Z(n3353) );
  NAND U4618 ( .A(n3351), .B(n3353), .Z(n7806) );
  XOR U4619 ( .A(n7822), .B(sreg[1487]), .Z(n3354) );
  NANDN U4620 ( .A(n7823), .B(n3354), .Z(n3355) );
  NAND U4621 ( .A(n7822), .B(sreg[1487]), .Z(n3356) );
  AND U4622 ( .A(n3355), .B(n3356), .Z(n7829) );
  NAND U4623 ( .A(n7846), .B(sreg[1490]), .Z(n3357) );
  XOR U4624 ( .A(sreg[1490]), .B(n7846), .Z(n3358) );
  NANDN U4625 ( .A(n7845), .B(n3358), .Z(n3359) );
  NAND U4626 ( .A(n3357), .B(n3359), .Z(n7854) );
  XOR U4627 ( .A(n7873), .B(sreg[1493]), .Z(n3360) );
  NANDN U4628 ( .A(n7874), .B(n3360), .Z(n3361) );
  NAND U4629 ( .A(n7873), .B(sreg[1493]), .Z(n3362) );
  AND U4630 ( .A(n3361), .B(n3362), .Z(n7880) );
  NAND U4631 ( .A(n7897), .B(sreg[1496]), .Z(n3363) );
  XOR U4632 ( .A(sreg[1496]), .B(n7897), .Z(n3364) );
  NANDN U4633 ( .A(n7896), .B(n3364), .Z(n3365) );
  NAND U4634 ( .A(n3363), .B(n3365), .Z(n7905) );
  XOR U4635 ( .A(n7921), .B(sreg[1499]), .Z(n3366) );
  NANDN U4636 ( .A(n7922), .B(n3366), .Z(n3367) );
  NAND U4637 ( .A(n7921), .B(sreg[1499]), .Z(n3368) );
  AND U4638 ( .A(n3367), .B(n3368), .Z(n7928) );
  NAND U4639 ( .A(n7945), .B(sreg[1502]), .Z(n3369) );
  XOR U4640 ( .A(sreg[1502]), .B(n7945), .Z(n3370) );
  NANDN U4641 ( .A(n7944), .B(n3370), .Z(n3371) );
  NAND U4642 ( .A(n3369), .B(n3371), .Z(n7953) );
  XOR U4643 ( .A(n7969), .B(sreg[1505]), .Z(n3372) );
  NANDN U4644 ( .A(n7970), .B(n3372), .Z(n3373) );
  NAND U4645 ( .A(n7969), .B(sreg[1505]), .Z(n3374) );
  AND U4646 ( .A(n3373), .B(n3374), .Z(n7979) );
  NAND U4647 ( .A(n7994), .B(sreg[1508]), .Z(n3375) );
  XOR U4648 ( .A(sreg[1508]), .B(n7994), .Z(n3376) );
  NAND U4649 ( .A(n3376), .B(n7993), .Z(n3377) );
  NAND U4650 ( .A(n3375), .B(n3377), .Z(n8002) );
  NAND U4651 ( .A(n8017), .B(sreg[1511]), .Z(n3378) );
  XOR U4652 ( .A(sreg[1511]), .B(n8017), .Z(n3379) );
  NAND U4653 ( .A(n3379), .B(n8016), .Z(n3380) );
  NAND U4654 ( .A(n3378), .B(n3380), .Z(n8025) );
  XOR U4655 ( .A(n8041), .B(sreg[1514]), .Z(n3381) );
  NANDN U4656 ( .A(n8042), .B(n3381), .Z(n3382) );
  NAND U4657 ( .A(n8041), .B(sreg[1514]), .Z(n3383) );
  AND U4658 ( .A(n3382), .B(n3383), .Z(n8048) );
  NAND U4659 ( .A(n8067), .B(sreg[1517]), .Z(n3384) );
  XOR U4660 ( .A(sreg[1517]), .B(n8067), .Z(n3385) );
  NANDN U4661 ( .A(n8068), .B(n3385), .Z(n3386) );
  NAND U4662 ( .A(n3384), .B(n3386), .Z(n8076) );
  NAND U4663 ( .A(n8093), .B(sreg[1520]), .Z(n3387) );
  XOR U4664 ( .A(sreg[1520]), .B(n8093), .Z(n3388) );
  NANDN U4665 ( .A(n8092), .B(n3388), .Z(n3389) );
  NAND U4666 ( .A(n3387), .B(n3389), .Z(n8101) );
  XOR U4667 ( .A(n8117), .B(sreg[1523]), .Z(n3390) );
  NANDN U4668 ( .A(n8118), .B(n3390), .Z(n3391) );
  NAND U4669 ( .A(n8117), .B(sreg[1523]), .Z(n3392) );
  AND U4670 ( .A(n3391), .B(n3392), .Z(n8124) );
  NAND U4671 ( .A(n8141), .B(sreg[1526]), .Z(n3393) );
  XOR U4672 ( .A(sreg[1526]), .B(n8141), .Z(n3394) );
  NANDN U4673 ( .A(n8140), .B(n3394), .Z(n3395) );
  NAND U4674 ( .A(n3393), .B(n3395), .Z(n8149) );
  XOR U4675 ( .A(n8165), .B(sreg[1529]), .Z(n3396) );
  NANDN U4676 ( .A(n8166), .B(n3396), .Z(n3397) );
  NAND U4677 ( .A(n8165), .B(sreg[1529]), .Z(n3398) );
  AND U4678 ( .A(n3397), .B(n3398), .Z(n8172) );
  NAND U4679 ( .A(n8192), .B(sreg[1532]), .Z(n3399) );
  XOR U4680 ( .A(sreg[1532]), .B(n8192), .Z(n3400) );
  NANDN U4681 ( .A(n8191), .B(n3400), .Z(n3401) );
  NAND U4682 ( .A(n3399), .B(n3401), .Z(n8200) );
  XOR U4683 ( .A(n8216), .B(sreg[1535]), .Z(n3402) );
  NANDN U4684 ( .A(n8217), .B(n3402), .Z(n3403) );
  NAND U4685 ( .A(n8216), .B(sreg[1535]), .Z(n3404) );
  AND U4686 ( .A(n3403), .B(n3404), .Z(n8223) );
  NAND U4687 ( .A(n8240), .B(sreg[1538]), .Z(n3405) );
  XOR U4688 ( .A(sreg[1538]), .B(n8240), .Z(n3406) );
  NANDN U4689 ( .A(n8239), .B(n3406), .Z(n3407) );
  NAND U4690 ( .A(n3405), .B(n3407), .Z(n8248) );
  NAND U4691 ( .A(n8263), .B(sreg[1541]), .Z(n3408) );
  XOR U4692 ( .A(sreg[1541]), .B(n8263), .Z(n3409) );
  NAND U4693 ( .A(n3409), .B(n8262), .Z(n3410) );
  NAND U4694 ( .A(n3408), .B(n3410), .Z(n8269) );
  NAND U4695 ( .A(n8289), .B(sreg[1544]), .Z(n3411) );
  XOR U4696 ( .A(sreg[1544]), .B(n8289), .Z(n3412) );
  NANDN U4697 ( .A(n8288), .B(n3412), .Z(n3413) );
  NAND U4698 ( .A(n3411), .B(n3413), .Z(n8297) );
  XOR U4699 ( .A(n8313), .B(sreg[1547]), .Z(n3414) );
  NANDN U4700 ( .A(n8314), .B(n3414), .Z(n3415) );
  NAND U4701 ( .A(n8313), .B(sreg[1547]), .Z(n3416) );
  AND U4702 ( .A(n3415), .B(n3416), .Z(n8320) );
  NAND U4703 ( .A(n8337), .B(sreg[1550]), .Z(n3417) );
  XOR U4704 ( .A(sreg[1550]), .B(n8337), .Z(n3418) );
  NANDN U4705 ( .A(n8336), .B(n3418), .Z(n3419) );
  NAND U4706 ( .A(n3417), .B(n3419), .Z(n8345) );
  XOR U4707 ( .A(n8361), .B(sreg[1553]), .Z(n3420) );
  NANDN U4708 ( .A(n8362), .B(n3420), .Z(n3421) );
  NAND U4709 ( .A(n8361), .B(sreg[1553]), .Z(n3422) );
  AND U4710 ( .A(n3421), .B(n3422), .Z(n8368) );
  NAND U4711 ( .A(n8385), .B(sreg[1556]), .Z(n3423) );
  XOR U4712 ( .A(sreg[1556]), .B(n8385), .Z(n3424) );
  NANDN U4713 ( .A(n8384), .B(n3424), .Z(n3425) );
  NAND U4714 ( .A(n3423), .B(n3425), .Z(n8393) );
  XOR U4715 ( .A(n8412), .B(sreg[1559]), .Z(n3426) );
  NANDN U4716 ( .A(n8413), .B(n3426), .Z(n3427) );
  NAND U4717 ( .A(n8412), .B(sreg[1559]), .Z(n3428) );
  AND U4718 ( .A(n3427), .B(n3428), .Z(n8419) );
  NAND U4719 ( .A(n8434), .B(sreg[1562]), .Z(n3429) );
  XOR U4720 ( .A(sreg[1562]), .B(n8434), .Z(n3430) );
  NAND U4721 ( .A(n3430), .B(n8433), .Z(n3431) );
  NAND U4722 ( .A(n3429), .B(n3431), .Z(n8442) );
  XOR U4723 ( .A(n8458), .B(sreg[1565]), .Z(n3432) );
  NANDN U4724 ( .A(n8459), .B(n3432), .Z(n3433) );
  NAND U4725 ( .A(n8458), .B(sreg[1565]), .Z(n3434) );
  AND U4726 ( .A(n3433), .B(n3434), .Z(n8465) );
  NAND U4727 ( .A(n8482), .B(sreg[1568]), .Z(n3435) );
  XOR U4728 ( .A(sreg[1568]), .B(n8482), .Z(n3436) );
  NANDN U4729 ( .A(n8481), .B(n3436), .Z(n3437) );
  NAND U4730 ( .A(n3435), .B(n3437), .Z(n8490) );
  NAND U4731 ( .A(n8509), .B(sreg[1571]), .Z(n3438) );
  XOR U4732 ( .A(sreg[1571]), .B(n8509), .Z(n3439) );
  NANDN U4733 ( .A(n8510), .B(n3439), .Z(n3440) );
  NAND U4734 ( .A(n3438), .B(n3440), .Z(n8518) );
  NAND U4735 ( .A(n8536), .B(sreg[1574]), .Z(n3441) );
  XOR U4736 ( .A(sreg[1574]), .B(n8536), .Z(n3442) );
  NANDN U4737 ( .A(n8537), .B(n3442), .Z(n3443) );
  NAND U4738 ( .A(n3441), .B(n3443), .Z(n8545) );
  NAND U4739 ( .A(n8561), .B(sreg[1577]), .Z(n3444) );
  XOR U4740 ( .A(sreg[1577]), .B(n8561), .Z(n3445) );
  NANDN U4741 ( .A(n8562), .B(n3445), .Z(n3446) );
  NAND U4742 ( .A(n3444), .B(n3446), .Z(n8570) );
  NAND U4743 ( .A(n8587), .B(sreg[1580]), .Z(n3447) );
  XOR U4744 ( .A(sreg[1580]), .B(n8587), .Z(n3448) );
  NANDN U4745 ( .A(n8586), .B(n3448), .Z(n3449) );
  NAND U4746 ( .A(n3447), .B(n3449), .Z(n8595) );
  XOR U4747 ( .A(n8611), .B(sreg[1583]), .Z(n3450) );
  NANDN U4748 ( .A(n8612), .B(n3450), .Z(n3451) );
  NAND U4749 ( .A(n8611), .B(sreg[1583]), .Z(n3452) );
  AND U4750 ( .A(n3451), .B(n3452), .Z(n8618) );
  NAND U4751 ( .A(n8635), .B(sreg[1586]), .Z(n3453) );
  XOR U4752 ( .A(sreg[1586]), .B(n8635), .Z(n3454) );
  NANDN U4753 ( .A(n8634), .B(n3454), .Z(n3455) );
  NAND U4754 ( .A(n3453), .B(n3455), .Z(n8641) );
  XOR U4755 ( .A(n8660), .B(sreg[1589]), .Z(n3456) );
  NANDN U4756 ( .A(n8661), .B(n3456), .Z(n3457) );
  NAND U4757 ( .A(n8660), .B(sreg[1589]), .Z(n3458) );
  AND U4758 ( .A(n3457), .B(n3458), .Z(n8667) );
  NAND U4759 ( .A(n8684), .B(sreg[1592]), .Z(n3459) );
  XOR U4760 ( .A(sreg[1592]), .B(n8684), .Z(n3460) );
  NANDN U4761 ( .A(n8683), .B(n3460), .Z(n3461) );
  NAND U4762 ( .A(n3459), .B(n3461), .Z(n8692) );
  XOR U4763 ( .A(n8708), .B(sreg[1595]), .Z(n3462) );
  NANDN U4764 ( .A(n8709), .B(n3462), .Z(n3463) );
  NAND U4765 ( .A(n8708), .B(sreg[1595]), .Z(n3464) );
  AND U4766 ( .A(n3463), .B(n3464), .Z(n8715) );
  NAND U4767 ( .A(n8732), .B(sreg[1598]), .Z(n3465) );
  XOR U4768 ( .A(sreg[1598]), .B(n8732), .Z(n3466) );
  NANDN U4769 ( .A(n8731), .B(n3466), .Z(n3467) );
  NAND U4770 ( .A(n3465), .B(n3467), .Z(n8740) );
  XOR U4771 ( .A(n8756), .B(sreg[1601]), .Z(n3468) );
  NANDN U4772 ( .A(n8757), .B(n3468), .Z(n3469) );
  NAND U4773 ( .A(n8756), .B(sreg[1601]), .Z(n3470) );
  AND U4774 ( .A(n3469), .B(n3470), .Z(n8766) );
  NAND U4775 ( .A(n8783), .B(sreg[1604]), .Z(n3471) );
  XOR U4776 ( .A(sreg[1604]), .B(n8783), .Z(n3472) );
  NANDN U4777 ( .A(n8782), .B(n3472), .Z(n3473) );
  NAND U4778 ( .A(n3471), .B(n3473), .Z(n8791) );
  XOR U4779 ( .A(n8807), .B(sreg[1607]), .Z(n3474) );
  NANDN U4780 ( .A(n8808), .B(n3474), .Z(n3475) );
  NAND U4781 ( .A(n8807), .B(sreg[1607]), .Z(n3476) );
  AND U4782 ( .A(n3475), .B(n3476), .Z(n8814) );
  NAND U4783 ( .A(n8830), .B(sreg[1610]), .Z(n3477) );
  XOR U4784 ( .A(sreg[1610]), .B(n8830), .Z(n3478) );
  NANDN U4785 ( .A(n8831), .B(n3478), .Z(n3479) );
  NAND U4786 ( .A(n3477), .B(n3479), .Z(n8839) );
  XOR U4787 ( .A(n8855), .B(sreg[1613]), .Z(n3480) );
  NANDN U4788 ( .A(n8856), .B(n3480), .Z(n3481) );
  NAND U4789 ( .A(n8855), .B(sreg[1613]), .Z(n3482) );
  AND U4790 ( .A(n3481), .B(n3482), .Z(n8862) );
  NAND U4791 ( .A(n8882), .B(sreg[1616]), .Z(n3483) );
  XOR U4792 ( .A(sreg[1616]), .B(n8882), .Z(n3484) );
  NANDN U4793 ( .A(n8881), .B(n3484), .Z(n3485) );
  NAND U4794 ( .A(n3483), .B(n3485), .Z(n8890) );
  XOR U4795 ( .A(n8908), .B(sreg[1619]), .Z(n3486) );
  NANDN U4796 ( .A(n8909), .B(n3486), .Z(n3487) );
  NAND U4797 ( .A(n8908), .B(sreg[1619]), .Z(n3488) );
  AND U4798 ( .A(n3487), .B(n3488), .Z(n8915) );
  NAND U4799 ( .A(n8932), .B(sreg[1622]), .Z(n3489) );
  XOR U4800 ( .A(sreg[1622]), .B(n8932), .Z(n3490) );
  NANDN U4801 ( .A(n8931), .B(n3490), .Z(n3491) );
  NAND U4802 ( .A(n3489), .B(n3491), .Z(n8940) );
  NAND U4803 ( .A(n8955), .B(sreg[1625]), .Z(n3492) );
  XOR U4804 ( .A(sreg[1625]), .B(n8955), .Z(n3493) );
  NAND U4805 ( .A(n3493), .B(n8954), .Z(n3494) );
  NAND U4806 ( .A(n3492), .B(n3494), .Z(n8961) );
  NAND U4807 ( .A(n8979), .B(sreg[1628]), .Z(n3495) );
  XOR U4808 ( .A(sreg[1628]), .B(n8979), .Z(n3496) );
  NANDN U4809 ( .A(n8980), .B(n3496), .Z(n3497) );
  NAND U4810 ( .A(n3495), .B(n3497), .Z(n8988) );
  NAND U4811 ( .A(n9004), .B(sreg[1631]), .Z(n3498) );
  XOR U4812 ( .A(sreg[1631]), .B(n9004), .Z(n3499) );
  NANDN U4813 ( .A(n9005), .B(n3499), .Z(n3500) );
  NAND U4814 ( .A(n3498), .B(n3500), .Z(n9013) );
  NAND U4815 ( .A(n9033), .B(sreg[1634]), .Z(n3501) );
  XOR U4816 ( .A(sreg[1634]), .B(n9033), .Z(n3502) );
  NANDN U4817 ( .A(n9032), .B(n3502), .Z(n3503) );
  NAND U4818 ( .A(n3501), .B(n3503), .Z(n9041) );
  NAND U4819 ( .A(n9057), .B(sreg[1637]), .Z(n3504) );
  XOR U4820 ( .A(sreg[1637]), .B(n9057), .Z(n3505) );
  NANDN U4821 ( .A(n9058), .B(n3505), .Z(n3506) );
  NAND U4822 ( .A(n3504), .B(n3506), .Z(n9066) );
  NAND U4823 ( .A(n9083), .B(sreg[1640]), .Z(n3507) );
  XOR U4824 ( .A(sreg[1640]), .B(n9083), .Z(n3508) );
  NANDN U4825 ( .A(n9082), .B(n3508), .Z(n3509) );
  NAND U4826 ( .A(n3507), .B(n3509), .Z(n9091) );
  XOR U4827 ( .A(n9107), .B(sreg[1643]), .Z(n3510) );
  NANDN U4828 ( .A(n9108), .B(n3510), .Z(n3511) );
  NAND U4829 ( .A(n9107), .B(sreg[1643]), .Z(n3512) );
  AND U4830 ( .A(n3511), .B(n3512), .Z(n9114) );
  NAND U4831 ( .A(n9129), .B(sreg[1646]), .Z(n3513) );
  XOR U4832 ( .A(sreg[1646]), .B(n9129), .Z(n3514) );
  NAND U4833 ( .A(n3514), .B(n9128), .Z(n3515) );
  NAND U4834 ( .A(n3513), .B(n3515), .Z(n9137) );
  XOR U4835 ( .A(n9156), .B(sreg[1649]), .Z(n3516) );
  NANDN U4836 ( .A(n9157), .B(n3516), .Z(n3517) );
  NAND U4837 ( .A(n9156), .B(sreg[1649]), .Z(n3518) );
  AND U4838 ( .A(n3517), .B(n3518), .Z(n9163) );
  NAND U4839 ( .A(n9180), .B(sreg[1652]), .Z(n3519) );
  XOR U4840 ( .A(sreg[1652]), .B(n9180), .Z(n3520) );
  NANDN U4841 ( .A(n9179), .B(n3520), .Z(n3521) );
  NAND U4842 ( .A(n3519), .B(n3521), .Z(n9186) );
  XOR U4843 ( .A(n9202), .B(sreg[1655]), .Z(n3522) );
  NANDN U4844 ( .A(n9203), .B(n3522), .Z(n3523) );
  NAND U4845 ( .A(n9202), .B(sreg[1655]), .Z(n3524) );
  AND U4846 ( .A(n3523), .B(n3524), .Z(n9209) );
  NAND U4847 ( .A(n9227), .B(sreg[1658]), .Z(n3525) );
  XOR U4848 ( .A(sreg[1658]), .B(n9227), .Z(n3526) );
  NAND U4849 ( .A(n3526), .B(n9226), .Z(n3527) );
  NAND U4850 ( .A(n3525), .B(n3527), .Z(n9235) );
  XOR U4851 ( .A(n9251), .B(sreg[1661]), .Z(n3528) );
  NANDN U4852 ( .A(n9252), .B(n3528), .Z(n3529) );
  NAND U4853 ( .A(n9251), .B(sreg[1661]), .Z(n3530) );
  AND U4854 ( .A(n3529), .B(n3530), .Z(n9258) );
  NAND U4855 ( .A(n9276), .B(sreg[1664]), .Z(n3531) );
  XOR U4856 ( .A(sreg[1664]), .B(n9276), .Z(n3532) );
  NANDN U4857 ( .A(n9277), .B(n3532), .Z(n3533) );
  NAND U4858 ( .A(n3531), .B(n3533), .Z(n9285) );
  XOR U4859 ( .A(n9301), .B(sreg[1667]), .Z(n3534) );
  NANDN U4860 ( .A(n9302), .B(n3534), .Z(n3535) );
  NAND U4861 ( .A(n9301), .B(sreg[1667]), .Z(n3536) );
  AND U4862 ( .A(n3535), .B(n3536), .Z(n9308) );
  NAND U4863 ( .A(n9325), .B(sreg[1670]), .Z(n3537) );
  XOR U4864 ( .A(sreg[1670]), .B(n9325), .Z(n3538) );
  NANDN U4865 ( .A(n9324), .B(n3538), .Z(n3539) );
  NAND U4866 ( .A(n3537), .B(n3539), .Z(n9331) );
  XOR U4867 ( .A(n9350), .B(sreg[1673]), .Z(n3540) );
  NANDN U4868 ( .A(n9351), .B(n3540), .Z(n3541) );
  NAND U4869 ( .A(n9350), .B(sreg[1673]), .Z(n3542) );
  AND U4870 ( .A(n3541), .B(n3542), .Z(n9357) );
  NAND U4871 ( .A(n9374), .B(sreg[1676]), .Z(n3543) );
  XOR U4872 ( .A(sreg[1676]), .B(n9374), .Z(n3544) );
  NANDN U4873 ( .A(n9373), .B(n3544), .Z(n3545) );
  NAND U4874 ( .A(n3543), .B(n3545), .Z(n9382) );
  XOR U4875 ( .A(n9398), .B(sreg[1679]), .Z(n3546) );
  NANDN U4876 ( .A(n9399), .B(n3546), .Z(n3547) );
  NAND U4877 ( .A(n9398), .B(sreg[1679]), .Z(n3548) );
  AND U4878 ( .A(n3547), .B(n3548), .Z(n9405) );
  NAND U4879 ( .A(n9420), .B(sreg[1682]), .Z(n3549) );
  XOR U4880 ( .A(sreg[1682]), .B(n9420), .Z(n3550) );
  NAND U4881 ( .A(n3550), .B(n9419), .Z(n3551) );
  NAND U4882 ( .A(n3549), .B(n3551), .Z(n9429) );
  XOR U4883 ( .A(n9445), .B(sreg[1685]), .Z(n3552) );
  NANDN U4884 ( .A(n9446), .B(n3552), .Z(n3553) );
  NAND U4885 ( .A(n9445), .B(sreg[1685]), .Z(n3554) );
  AND U4886 ( .A(n3553), .B(n3554), .Z(n9452) );
  NAND U4887 ( .A(n9469), .B(sreg[1688]), .Z(n3555) );
  XOR U4888 ( .A(sreg[1688]), .B(n9469), .Z(n3556) );
  NANDN U4889 ( .A(n9468), .B(n3556), .Z(n3557) );
  NAND U4890 ( .A(n3555), .B(n3557), .Z(n9477) );
  NAND U4891 ( .A(n9493), .B(sreg[1691]), .Z(n3558) );
  XOR U4892 ( .A(sreg[1691]), .B(n9493), .Z(n3559) );
  NANDN U4893 ( .A(n9494), .B(n3559), .Z(n3560) );
  NAND U4894 ( .A(n3558), .B(n3560), .Z(n9502) );
  NAND U4895 ( .A(n9519), .B(sreg[1694]), .Z(n3561) );
  XOR U4896 ( .A(sreg[1694]), .B(n9519), .Z(n3562) );
  NANDN U4897 ( .A(n9518), .B(n3562), .Z(n3563) );
  NAND U4898 ( .A(n3561), .B(n3563), .Z(n9527) );
  NAND U4899 ( .A(n9545), .B(sreg[1697]), .Z(n3564) );
  XOR U4900 ( .A(sreg[1697]), .B(n9545), .Z(n3565) );
  NAND U4901 ( .A(n3565), .B(n9544), .Z(n3566) );
  NAND U4902 ( .A(n3564), .B(n3566), .Z(n9551) );
  NAND U4903 ( .A(n9568), .B(sreg[1700]), .Z(n3567) );
  XOR U4904 ( .A(sreg[1700]), .B(n9568), .Z(n3568) );
  NANDN U4905 ( .A(n9567), .B(n3568), .Z(n3569) );
  NAND U4906 ( .A(n3567), .B(n3569), .Z(n9576) );
  XOR U4907 ( .A(n9592), .B(sreg[1703]), .Z(n3570) );
  NANDN U4908 ( .A(n9593), .B(n3570), .Z(n3571) );
  NAND U4909 ( .A(n9592), .B(sreg[1703]), .Z(n3572) );
  AND U4910 ( .A(n3571), .B(n3572), .Z(n9599) );
  NAND U4911 ( .A(n9617), .B(sreg[1706]), .Z(n3573) );
  XOR U4912 ( .A(sreg[1706]), .B(n9617), .Z(n3574) );
  NANDN U4913 ( .A(n9618), .B(n3574), .Z(n3575) );
  NAND U4914 ( .A(n3573), .B(n3575), .Z(n9626) );
  XOR U4915 ( .A(n9642), .B(sreg[1709]), .Z(n3576) );
  NANDN U4916 ( .A(n9643), .B(n3576), .Z(n3577) );
  NAND U4917 ( .A(n9642), .B(sreg[1709]), .Z(n3578) );
  AND U4918 ( .A(n3577), .B(n3578), .Z(n9649) );
  NAND U4919 ( .A(n9669), .B(sreg[1712]), .Z(n3579) );
  XOR U4920 ( .A(sreg[1712]), .B(n9669), .Z(n3580) );
  NANDN U4921 ( .A(n9668), .B(n3580), .Z(n3581) );
  NAND U4922 ( .A(n3579), .B(n3581), .Z(n9677) );
  XOR U4923 ( .A(n9693), .B(sreg[1715]), .Z(n3582) );
  NANDN U4924 ( .A(n9694), .B(n3582), .Z(n3583) );
  NAND U4925 ( .A(n9693), .B(sreg[1715]), .Z(n3584) );
  AND U4926 ( .A(n3583), .B(n3584), .Z(n9700) );
  NAND U4927 ( .A(n9717), .B(sreg[1718]), .Z(n3585) );
  XOR U4928 ( .A(sreg[1718]), .B(n9717), .Z(n3586) );
  NANDN U4929 ( .A(n9716), .B(n3586), .Z(n3587) );
  NAND U4930 ( .A(n3585), .B(n3587), .Z(n9725) );
  NAND U4931 ( .A(n9740), .B(sreg[1721]), .Z(n3588) );
  XOR U4932 ( .A(sreg[1721]), .B(n9740), .Z(n3589) );
  NAND U4933 ( .A(n3589), .B(n9739), .Z(n3590) );
  NAND U4934 ( .A(n3588), .B(n3590), .Z(n9746) );
  NAND U4935 ( .A(n9766), .B(sreg[1724]), .Z(n3591) );
  XOR U4936 ( .A(sreg[1724]), .B(n9766), .Z(n3592) );
  NANDN U4937 ( .A(n9765), .B(n3592), .Z(n3593) );
  NAND U4938 ( .A(n3591), .B(n3593), .Z(n9774) );
  XOR U4939 ( .A(n9790), .B(sreg[1727]), .Z(n3594) );
  NANDN U4940 ( .A(n9791), .B(n3594), .Z(n3595) );
  NAND U4941 ( .A(n9790), .B(sreg[1727]), .Z(n3596) );
  AND U4942 ( .A(n3595), .B(n3596), .Z(n9797) );
  NAND U4943 ( .A(n9814), .B(sreg[1730]), .Z(n3597) );
  XOR U4944 ( .A(sreg[1730]), .B(n9814), .Z(n3598) );
  NANDN U4945 ( .A(n9813), .B(n3598), .Z(n3599) );
  NAND U4946 ( .A(n3597), .B(n3599), .Z(n9820) );
  XOR U4947 ( .A(n9836), .B(sreg[1733]), .Z(n3600) );
  NANDN U4948 ( .A(n9837), .B(n3600), .Z(n3601) );
  NAND U4949 ( .A(n9836), .B(sreg[1733]), .Z(n3602) );
  AND U4950 ( .A(n3601), .B(n3602), .Z(n9843) );
  NAND U4951 ( .A(n9863), .B(sreg[1736]), .Z(n3603) );
  XOR U4952 ( .A(sreg[1736]), .B(n9863), .Z(n3604) );
  NANDN U4953 ( .A(n9862), .B(n3604), .Z(n3605) );
  NAND U4954 ( .A(n3603), .B(n3605), .Z(n9871) );
  XOR U4955 ( .A(n9887), .B(sreg[1739]), .Z(n3606) );
  NANDN U4956 ( .A(n9888), .B(n3606), .Z(n3607) );
  NAND U4957 ( .A(n9887), .B(sreg[1739]), .Z(n3608) );
  AND U4958 ( .A(n3607), .B(n3608), .Z(n9894) );
  NAND U4959 ( .A(n9911), .B(sreg[1742]), .Z(n3609) );
  XOR U4960 ( .A(sreg[1742]), .B(n9911), .Z(n3610) );
  NANDN U4961 ( .A(n9910), .B(n3610), .Z(n3611) );
  NAND U4962 ( .A(n3609), .B(n3611), .Z(n9919) );
  XOR U4963 ( .A(n9935), .B(sreg[1745]), .Z(n3612) );
  NANDN U4964 ( .A(n9936), .B(n3612), .Z(n3613) );
  NAND U4965 ( .A(n9935), .B(sreg[1745]), .Z(n3614) );
  AND U4966 ( .A(n3613), .B(n3614), .Z(n9942) );
  NAND U4967 ( .A(n9959), .B(sreg[1748]), .Z(n3615) );
  XOR U4968 ( .A(sreg[1748]), .B(n9959), .Z(n3616) );
  NANDN U4969 ( .A(n9958), .B(n3616), .Z(n3617) );
  NAND U4970 ( .A(n3615), .B(n3617), .Z(n9967) );
  XOR U4971 ( .A(n9986), .B(sreg[1751]), .Z(n3618) );
  NANDN U4972 ( .A(n9987), .B(n3618), .Z(n3619) );
  NAND U4973 ( .A(n9986), .B(sreg[1751]), .Z(n3620) );
  AND U4974 ( .A(n3619), .B(n3620), .Z(n9993) );
  NAND U4975 ( .A(n10010), .B(sreg[1754]), .Z(n3621) );
  XOR U4976 ( .A(sreg[1754]), .B(n10010), .Z(n3622) );
  NANDN U4977 ( .A(n10009), .B(n3622), .Z(n3623) );
  NAND U4978 ( .A(n3621), .B(n3623), .Z(n10018) );
  NAND U4979 ( .A(n10034), .B(sreg[1757]), .Z(n3624) );
  XOR U4980 ( .A(sreg[1757]), .B(n10034), .Z(n3625) );
  NANDN U4981 ( .A(n10035), .B(n3625), .Z(n3626) );
  NAND U4982 ( .A(n3624), .B(n3626), .Z(n10043) );
  NAND U4983 ( .A(n10060), .B(sreg[1760]), .Z(n3627) );
  XOR U4984 ( .A(sreg[1760]), .B(n10060), .Z(n3628) );
  NANDN U4985 ( .A(n10059), .B(n3628), .Z(n3629) );
  NAND U4986 ( .A(n3627), .B(n3629), .Z(n10068) );
  XOR U4987 ( .A(n10084), .B(sreg[1763]), .Z(n3630) );
  NANDN U4988 ( .A(n10085), .B(n3630), .Z(n3631) );
  NAND U4989 ( .A(n10084), .B(sreg[1763]), .Z(n3632) );
  AND U4990 ( .A(n3631), .B(n3632), .Z(n10091) );
  NAND U4991 ( .A(n10110), .B(sreg[1766]), .Z(n3633) );
  XOR U4992 ( .A(sreg[1766]), .B(n10110), .Z(n3634) );
  NANDN U4993 ( .A(n10111), .B(n3634), .Z(n3635) );
  NAND U4994 ( .A(n3633), .B(n3635), .Z(n10119) );
  XOR U4995 ( .A(n10135), .B(sreg[1769]), .Z(n3636) );
  NANDN U4996 ( .A(n10136), .B(n3636), .Z(n3637) );
  NAND U4997 ( .A(n10135), .B(sreg[1769]), .Z(n3638) );
  AND U4998 ( .A(n3637), .B(n3638), .Z(n10142) );
  NAND U4999 ( .A(n10159), .B(sreg[1772]), .Z(n3639) );
  XOR U5000 ( .A(sreg[1772]), .B(n10159), .Z(n3640) );
  NANDN U5001 ( .A(n10158), .B(n3640), .Z(n3641) );
  NAND U5002 ( .A(n3639), .B(n3641), .Z(n10167) );
  XOR U5003 ( .A(n10183), .B(sreg[1775]), .Z(n3642) );
  NANDN U5004 ( .A(n10184), .B(n3642), .Z(n3643) );
  NAND U5005 ( .A(n10183), .B(sreg[1775]), .Z(n3644) );
  AND U5006 ( .A(n3643), .B(n3644), .Z(n10190) );
  NAND U5007 ( .A(n10208), .B(sreg[1778]), .Z(n3645) );
  XOR U5008 ( .A(sreg[1778]), .B(n10208), .Z(n3646) );
  NAND U5009 ( .A(n3646), .B(n10207), .Z(n3647) );
  NAND U5010 ( .A(n3645), .B(n3647), .Z(n10216) );
  XOR U5011 ( .A(n10232), .B(sreg[1781]), .Z(n3648) );
  NANDN U5012 ( .A(n10233), .B(n3648), .Z(n3649) );
  NAND U5013 ( .A(n10232), .B(sreg[1781]), .Z(n3650) );
  AND U5014 ( .A(n3649), .B(n3650), .Z(n10239) );
  NAND U5015 ( .A(n10256), .B(sreg[1784]), .Z(n3651) );
  XOR U5016 ( .A(sreg[1784]), .B(n10256), .Z(n3652) );
  NANDN U5017 ( .A(n10255), .B(n3652), .Z(n3653) );
  NAND U5018 ( .A(n3651), .B(n3653), .Z(n10264) );
  XOR U5019 ( .A(n10280), .B(sreg[1787]), .Z(n3654) );
  NANDN U5020 ( .A(n10281), .B(n3654), .Z(n3655) );
  NAND U5021 ( .A(n10280), .B(sreg[1787]), .Z(n3656) );
  AND U5022 ( .A(n3655), .B(n3656), .Z(n10287) );
  NAND U5023 ( .A(n10304), .B(sreg[1790]), .Z(n3657) );
  XOR U5024 ( .A(sreg[1790]), .B(n10304), .Z(n3658) );
  NANDN U5025 ( .A(n10303), .B(n3658), .Z(n3659) );
  NAND U5026 ( .A(n3657), .B(n3659), .Z(n10312) );
  NAND U5027 ( .A(n10331), .B(sreg[1793]), .Z(n3660) );
  XOR U5028 ( .A(sreg[1793]), .B(n10331), .Z(n3661) );
  NANDN U5029 ( .A(n10332), .B(n3661), .Z(n3662) );
  NAND U5030 ( .A(n3660), .B(n3662), .Z(n10340) );
  NAND U5031 ( .A(n10357), .B(sreg[1796]), .Z(n3663) );
  XOR U5032 ( .A(sreg[1796]), .B(n10357), .Z(n3664) );
  NANDN U5033 ( .A(n10356), .B(n3664), .Z(n3665) );
  NAND U5034 ( .A(n3663), .B(n3665), .Z(n10365) );
  XOR U5035 ( .A(n10381), .B(sreg[1799]), .Z(n3666) );
  NANDN U5036 ( .A(n10382), .B(n3666), .Z(n3667) );
  NAND U5037 ( .A(n10381), .B(sreg[1799]), .Z(n3668) );
  AND U5038 ( .A(n3667), .B(n3668), .Z(n10388) );
  NAND U5039 ( .A(n10405), .B(sreg[1802]), .Z(n3669) );
  XOR U5040 ( .A(sreg[1802]), .B(n10405), .Z(n3670) );
  NANDN U5041 ( .A(n10404), .B(n3670), .Z(n3671) );
  NAND U5042 ( .A(n3669), .B(n3671), .Z(n10413) );
  XOR U5043 ( .A(n10429), .B(sreg[1805]), .Z(n3672) );
  NANDN U5044 ( .A(n10430), .B(n3672), .Z(n3673) );
  NAND U5045 ( .A(n10429), .B(sreg[1805]), .Z(n3674) );
  AND U5046 ( .A(n3673), .B(n3674), .Z(n10436) );
  NAND U5047 ( .A(n10456), .B(sreg[1808]), .Z(n3675) );
  XOR U5048 ( .A(sreg[1808]), .B(n10456), .Z(n3676) );
  NANDN U5049 ( .A(n10455), .B(n3676), .Z(n3677) );
  NAND U5050 ( .A(n3675), .B(n3677), .Z(n10464) );
  NAND U5051 ( .A(n10479), .B(sreg[1811]), .Z(n3678) );
  XOR U5052 ( .A(sreg[1811]), .B(n10479), .Z(n3679) );
  NAND U5053 ( .A(n3679), .B(n10478), .Z(n3680) );
  NAND U5054 ( .A(n3678), .B(n3680), .Z(n10485) );
  NAND U5055 ( .A(n10502), .B(sreg[1814]), .Z(n3681) );
  XOR U5056 ( .A(sreg[1814]), .B(n10502), .Z(n3682) );
  NANDN U5057 ( .A(n10501), .B(n3682), .Z(n3683) );
  NAND U5058 ( .A(n3681), .B(n3683), .Z(n10510) );
  XOR U5059 ( .A(n10526), .B(sreg[1817]), .Z(n3684) );
  NANDN U5060 ( .A(n10527), .B(n3684), .Z(n3685) );
  NAND U5061 ( .A(n10526), .B(sreg[1817]), .Z(n3686) );
  AND U5062 ( .A(n3685), .B(n3686), .Z(n10533) );
  NAND U5063 ( .A(n10553), .B(sreg[1820]), .Z(n3687) );
  XOR U5064 ( .A(sreg[1820]), .B(n10553), .Z(n3688) );
  NANDN U5065 ( .A(n10552), .B(n3688), .Z(n3689) );
  NAND U5066 ( .A(n3687), .B(n3689), .Z(n10561) );
  XOR U5067 ( .A(n10577), .B(sreg[1823]), .Z(n3690) );
  NANDN U5068 ( .A(n10578), .B(n3690), .Z(n3691) );
  NAND U5069 ( .A(n10577), .B(sreg[1823]), .Z(n3692) );
  AND U5070 ( .A(n3691), .B(n3692), .Z(n10584) );
  NAND U5071 ( .A(n10601), .B(sreg[1826]), .Z(n3693) );
  XOR U5072 ( .A(sreg[1826]), .B(n10601), .Z(n3694) );
  NANDN U5073 ( .A(n10600), .B(n3694), .Z(n3695) );
  NAND U5074 ( .A(n3693), .B(n3695), .Z(n10609) );
  NAND U5075 ( .A(n10624), .B(sreg[1829]), .Z(n3696) );
  XOR U5076 ( .A(sreg[1829]), .B(n10624), .Z(n3697) );
  NAND U5077 ( .A(n3697), .B(n10623), .Z(n3698) );
  NAND U5078 ( .A(n3696), .B(n3698), .Z(n10630) );
  NAND U5079 ( .A(n10648), .B(sreg[1832]), .Z(n3699) );
  XOR U5080 ( .A(sreg[1832]), .B(n10648), .Z(n3700) );
  NANDN U5081 ( .A(n10649), .B(n3700), .Z(n3701) );
  NAND U5082 ( .A(n3699), .B(n3701), .Z(n10657) );
  XOR U5083 ( .A(n10676), .B(sreg[1835]), .Z(n3702) );
  NANDN U5084 ( .A(n10677), .B(n3702), .Z(n3703) );
  NAND U5085 ( .A(n10676), .B(sreg[1835]), .Z(n3704) );
  AND U5086 ( .A(n3703), .B(n3704), .Z(n10683) );
  NAND U5087 ( .A(n10698), .B(sreg[1838]), .Z(n3705) );
  XOR U5088 ( .A(sreg[1838]), .B(n10698), .Z(n3706) );
  NAND U5089 ( .A(n3706), .B(n10697), .Z(n3707) );
  NAND U5090 ( .A(n3705), .B(n3707), .Z(n10706) );
  XOR U5091 ( .A(n10722), .B(sreg[1841]), .Z(n3708) );
  NANDN U5092 ( .A(n10723), .B(n3708), .Z(n3709) );
  NAND U5093 ( .A(n10722), .B(sreg[1841]), .Z(n3710) );
  AND U5094 ( .A(n3709), .B(n3710), .Z(n10729) );
  NAND U5095 ( .A(n10745), .B(sreg[1844]), .Z(n3711) );
  XOR U5096 ( .A(sreg[1844]), .B(n10745), .Z(n3712) );
  NANDN U5097 ( .A(n10746), .B(n3712), .Z(n3713) );
  NAND U5098 ( .A(n3711), .B(n3713), .Z(n10754) );
  NAND U5099 ( .A(n10773), .B(sreg[1847]), .Z(n3714) );
  XOR U5100 ( .A(sreg[1847]), .B(n10773), .Z(n3715) );
  NANDN U5101 ( .A(n10774), .B(n3715), .Z(n3716) );
  NAND U5102 ( .A(n3714), .B(n3716), .Z(n10782) );
  NAND U5103 ( .A(n10798), .B(sreg[1850]), .Z(n3717) );
  XOR U5104 ( .A(sreg[1850]), .B(n10798), .Z(n3718) );
  NANDN U5105 ( .A(n10799), .B(n3718), .Z(n3719) );
  NAND U5106 ( .A(n3717), .B(n3719), .Z(n10807) );
  XOR U5107 ( .A(n10823), .B(sreg[1853]), .Z(n3720) );
  NANDN U5108 ( .A(n10824), .B(n3720), .Z(n3721) );
  NAND U5109 ( .A(n10823), .B(sreg[1853]), .Z(n3722) );
  AND U5110 ( .A(n3721), .B(n3722), .Z(n10830) );
  NAND U5111 ( .A(n10847), .B(sreg[1856]), .Z(n3723) );
  XOR U5112 ( .A(sreg[1856]), .B(n10847), .Z(n3724) );
  NANDN U5113 ( .A(n10846), .B(n3724), .Z(n3725) );
  NAND U5114 ( .A(n3723), .B(n3725), .Z(n10855) );
  NAND U5115 ( .A(n10872), .B(sreg[1859]), .Z(n3726) );
  XOR U5116 ( .A(sreg[1859]), .B(n10872), .Z(n3727) );
  NANDN U5117 ( .A(n10871), .B(n3727), .Z(n3728) );
  NAND U5118 ( .A(n3726), .B(n3728), .Z(n10880) );
  XOR U5119 ( .A(n10898), .B(sreg[1862]), .Z(n3729) );
  NANDN U5120 ( .A(n10899), .B(n3729), .Z(n3730) );
  NAND U5121 ( .A(n10898), .B(sreg[1862]), .Z(n3731) );
  AND U5122 ( .A(n3730), .B(n3731), .Z(n10905) );
  XOR U5123 ( .A(n10923), .B(sreg[1865]), .Z(n3732) );
  NANDN U5124 ( .A(n10924), .B(n3732), .Z(n3733) );
  NAND U5125 ( .A(n10923), .B(sreg[1865]), .Z(n3734) );
  AND U5126 ( .A(n3733), .B(n3734), .Z(n10933) );
  NAND U5127 ( .A(n10950), .B(sreg[1868]), .Z(n3735) );
  XOR U5128 ( .A(sreg[1868]), .B(n10950), .Z(n3736) );
  NANDN U5129 ( .A(n10949), .B(n3736), .Z(n3737) );
  NAND U5130 ( .A(n3735), .B(n3737), .Z(n10958) );
  XOR U5131 ( .A(n10974), .B(sreg[1871]), .Z(n3738) );
  NANDN U5132 ( .A(n10975), .B(n3738), .Z(n3739) );
  NAND U5133 ( .A(n10974), .B(sreg[1871]), .Z(n3740) );
  AND U5134 ( .A(n3739), .B(n3740), .Z(n10981) );
  NAND U5135 ( .A(n10996), .B(sreg[1874]), .Z(n3741) );
  XOR U5136 ( .A(sreg[1874]), .B(n10996), .Z(n3742) );
  NAND U5137 ( .A(n3742), .B(n10995), .Z(n3743) );
  NAND U5138 ( .A(n3741), .B(n3743), .Z(n11004) );
  NAND U5139 ( .A(n11022), .B(sreg[1877]), .Z(n3744) );
  XOR U5140 ( .A(sreg[1877]), .B(n11022), .Z(n3745) );
  NANDN U5141 ( .A(n11023), .B(n3745), .Z(n3746) );
  NAND U5142 ( .A(n3744), .B(n3746), .Z(n11031) );
  NAND U5143 ( .A(n11049), .B(sreg[1880]), .Z(n3747) );
  XOR U5144 ( .A(sreg[1880]), .B(n11049), .Z(n3748) );
  NANDN U5145 ( .A(n11050), .B(n3748), .Z(n3749) );
  NAND U5146 ( .A(n3747), .B(n3749), .Z(n11058) );
  NAND U5147 ( .A(n11074), .B(sreg[1883]), .Z(n3750) );
  XOR U5148 ( .A(sreg[1883]), .B(n11074), .Z(n3751) );
  NANDN U5149 ( .A(n11075), .B(n3751), .Z(n3752) );
  NAND U5150 ( .A(n3750), .B(n3752), .Z(n11083) );
  NAND U5151 ( .A(n11103), .B(sreg[1886]), .Z(n3753) );
  XOR U5152 ( .A(sreg[1886]), .B(n11103), .Z(n3754) );
  NANDN U5153 ( .A(n11102), .B(n3754), .Z(n3755) );
  NAND U5154 ( .A(n3753), .B(n3755), .Z(n11111) );
  XOR U5155 ( .A(n11127), .B(sreg[1889]), .Z(n3756) );
  NANDN U5156 ( .A(n11128), .B(n3756), .Z(n3757) );
  NAND U5157 ( .A(n11127), .B(sreg[1889]), .Z(n3758) );
  AND U5158 ( .A(n3757), .B(n3758), .Z(n11134) );
  NAND U5159 ( .A(n11151), .B(sreg[1892]), .Z(n3759) );
  XOR U5160 ( .A(sreg[1892]), .B(n11151), .Z(n3760) );
  NANDN U5161 ( .A(n11150), .B(n3760), .Z(n3761) );
  NAND U5162 ( .A(n3759), .B(n3761), .Z(n11159) );
  NAND U5163 ( .A(n11174), .B(sreg[1895]), .Z(n3762) );
  XOR U5164 ( .A(sreg[1895]), .B(n11174), .Z(n3763) );
  NAND U5165 ( .A(n3763), .B(n11173), .Z(n3764) );
  NAND U5166 ( .A(n3762), .B(n3764), .Z(n11180) );
  NAND U5167 ( .A(n11200), .B(sreg[1898]), .Z(n3765) );
  XOR U5168 ( .A(sreg[1898]), .B(n11200), .Z(n3766) );
  NANDN U5169 ( .A(n11199), .B(n3766), .Z(n3767) );
  NAND U5170 ( .A(n3765), .B(n3767), .Z(n11206) );
  XOR U5171 ( .A(n11222), .B(sreg[1901]), .Z(n3768) );
  NANDN U5172 ( .A(n11223), .B(n3768), .Z(n3769) );
  NAND U5173 ( .A(n11222), .B(sreg[1901]), .Z(n3770) );
  AND U5174 ( .A(n3769), .B(n3770), .Z(n11229) );
  NAND U5175 ( .A(n11246), .B(sreg[1904]), .Z(n3771) );
  XOR U5176 ( .A(sreg[1904]), .B(n11246), .Z(n3772) );
  NANDN U5177 ( .A(n11245), .B(n3772), .Z(n3773) );
  NAND U5178 ( .A(n3771), .B(n3773), .Z(n11254) );
  XOR U5179 ( .A(n11270), .B(sreg[1907]), .Z(n3774) );
  NANDN U5180 ( .A(n11271), .B(n3774), .Z(n3775) );
  NAND U5181 ( .A(n11270), .B(sreg[1907]), .Z(n3776) );
  AND U5182 ( .A(n3775), .B(n3776), .Z(n11277) );
  NAND U5183 ( .A(n11297), .B(sreg[1910]), .Z(n3777) );
  XOR U5184 ( .A(sreg[1910]), .B(n11297), .Z(n3778) );
  NANDN U5185 ( .A(n11296), .B(n3778), .Z(n3779) );
  NAND U5186 ( .A(n3777), .B(n3779), .Z(n11305) );
  XOR U5187 ( .A(n11321), .B(sreg[1913]), .Z(n3780) );
  NANDN U5188 ( .A(n11322), .B(n3780), .Z(n3781) );
  NAND U5189 ( .A(n11321), .B(sreg[1913]), .Z(n3782) );
  AND U5190 ( .A(n3781), .B(n3782), .Z(n11328) );
  NAND U5191 ( .A(n11345), .B(sreg[1916]), .Z(n3783) );
  XOR U5192 ( .A(sreg[1916]), .B(n11345), .Z(n3784) );
  NANDN U5193 ( .A(n11344), .B(n3784), .Z(n3785) );
  NAND U5194 ( .A(n3783), .B(n3785), .Z(n11353) );
  NAND U5195 ( .A(n11371), .B(sreg[1919]), .Z(n3786) );
  XOR U5196 ( .A(sreg[1919]), .B(n11371), .Z(n3787) );
  NANDN U5197 ( .A(n11372), .B(n3787), .Z(n3788) );
  NAND U5198 ( .A(n3786), .B(n3788), .Z(n11380) );
  NAND U5199 ( .A(n11397), .B(sreg[1922]), .Z(n3789) );
  XOR U5200 ( .A(sreg[1922]), .B(n11397), .Z(n3790) );
  NANDN U5201 ( .A(n11396), .B(n3790), .Z(n3791) );
  NAND U5202 ( .A(n3789), .B(n3791), .Z(n11405) );
  NAND U5203 ( .A(n11422), .B(sreg[1925]), .Z(n3792) );
  XOR U5204 ( .A(sreg[1925]), .B(n11422), .Z(n3793) );
  NANDN U5205 ( .A(n11421), .B(n3793), .Z(n3794) );
  NAND U5206 ( .A(n3792), .B(n3794), .Z(n11428) );
  NAND U5207 ( .A(n11446), .B(sreg[1928]), .Z(n3795) );
  XOR U5208 ( .A(sreg[1928]), .B(n11446), .Z(n3796) );
  NANDN U5209 ( .A(n11447), .B(n3796), .Z(n3797) );
  NAND U5210 ( .A(n3795), .B(n3797), .Z(n11455) );
  XOR U5211 ( .A(n11474), .B(sreg[1931]), .Z(n3798) );
  NANDN U5212 ( .A(n11475), .B(n3798), .Z(n3799) );
  NAND U5213 ( .A(n11474), .B(sreg[1931]), .Z(n3800) );
  AND U5214 ( .A(n3799), .B(n3800), .Z(n11481) );
  NAND U5215 ( .A(n11499), .B(sreg[1934]), .Z(n3801) );
  XOR U5216 ( .A(sreg[1934]), .B(n11499), .Z(n3802) );
  NANDN U5217 ( .A(n11500), .B(n3802), .Z(n3803) );
  NAND U5218 ( .A(n3801), .B(n3803), .Z(n11508) );
  XOR U5219 ( .A(n11524), .B(sreg[1937]), .Z(n3804) );
  NANDN U5220 ( .A(n11525), .B(n3804), .Z(n3805) );
  NAND U5221 ( .A(n11524), .B(sreg[1937]), .Z(n3806) );
  AND U5222 ( .A(n3805), .B(n3806), .Z(n11531) );
  NAND U5223 ( .A(n11546), .B(sreg[1940]), .Z(n3807) );
  XOR U5224 ( .A(sreg[1940]), .B(n11546), .Z(n3808) );
  NAND U5225 ( .A(n3808), .B(n11545), .Z(n3809) );
  NAND U5226 ( .A(n3807), .B(n3809), .Z(n11554) );
  XOR U5227 ( .A(n11572), .B(sreg[1943]), .Z(n3810) );
  NANDN U5228 ( .A(n11573), .B(n3810), .Z(n3811) );
  NAND U5229 ( .A(n11572), .B(sreg[1943]), .Z(n3812) );
  AND U5230 ( .A(n3811), .B(n3812), .Z(n11579) );
  NAND U5231 ( .A(n11599), .B(sreg[1946]), .Z(n3813) );
  XOR U5232 ( .A(sreg[1946]), .B(n11599), .Z(n3814) );
  NANDN U5233 ( .A(n11598), .B(n3814), .Z(n3815) );
  NAND U5234 ( .A(n3813), .B(n3815), .Z(n11607) );
  XOR U5235 ( .A(n11623), .B(sreg[1949]), .Z(n3816) );
  NANDN U5236 ( .A(n11624), .B(n3816), .Z(n3817) );
  NAND U5237 ( .A(n11623), .B(sreg[1949]), .Z(n3818) );
  AND U5238 ( .A(n3817), .B(n3818), .Z(n11630) );
  NAND U5239 ( .A(n11647), .B(sreg[1952]), .Z(n3819) );
  XOR U5240 ( .A(sreg[1952]), .B(n11647), .Z(n3820) );
  NANDN U5241 ( .A(n11646), .B(n3820), .Z(n3821) );
  NAND U5242 ( .A(n3819), .B(n3821), .Z(n11655) );
  XOR U5243 ( .A(n11673), .B(sreg[1955]), .Z(n3822) );
  NANDN U5244 ( .A(n11674), .B(n3822), .Z(n3823) );
  NAND U5245 ( .A(n11673), .B(sreg[1955]), .Z(n3824) );
  AND U5246 ( .A(n3823), .B(n3824), .Z(n11680) );
  NAND U5247 ( .A(n11697), .B(sreg[1958]), .Z(n3825) );
  XOR U5248 ( .A(sreg[1958]), .B(n11697), .Z(n3826) );
  NANDN U5249 ( .A(n11696), .B(n3826), .Z(n3827) );
  NAND U5250 ( .A(n3825), .B(n3827), .Z(n11703) );
  XOR U5251 ( .A(n11721), .B(sreg[1961]), .Z(n3828) );
  NANDN U5252 ( .A(n11722), .B(n3828), .Z(n3829) );
  NAND U5253 ( .A(n11721), .B(sreg[1961]), .Z(n3830) );
  AND U5254 ( .A(n3829), .B(n3830), .Z(n11731) );
  NAND U5255 ( .A(n11748), .B(sreg[1964]), .Z(n3831) );
  XOR U5256 ( .A(sreg[1964]), .B(n11748), .Z(n3832) );
  NANDN U5257 ( .A(n11747), .B(n3832), .Z(n3833) );
  NAND U5258 ( .A(n3831), .B(n3833), .Z(n11756) );
  NAND U5259 ( .A(n11772), .B(sreg[1967]), .Z(n3834) );
  XOR U5260 ( .A(sreg[1967]), .B(n11772), .Z(n3835) );
  NANDN U5261 ( .A(n11773), .B(n3835), .Z(n3836) );
  NAND U5262 ( .A(n3834), .B(n3836), .Z(n11781) );
  NAND U5263 ( .A(n11799), .B(sreg[1970]), .Z(n3837) );
  XOR U5264 ( .A(sreg[1970]), .B(n11799), .Z(n3838) );
  NANDN U5265 ( .A(n11800), .B(n3838), .Z(n3839) );
  NAND U5266 ( .A(n3837), .B(n3839), .Z(n11808) );
  XOR U5267 ( .A(n11826), .B(sreg[1973]), .Z(n3840) );
  NANDN U5268 ( .A(n11827), .B(n3840), .Z(n3841) );
  NAND U5269 ( .A(n11826), .B(sreg[1973]), .Z(n3842) );
  AND U5270 ( .A(n3841), .B(n3842), .Z(n11833) );
  NAND U5271 ( .A(n11850), .B(sreg[1976]), .Z(n3843) );
  XOR U5272 ( .A(sreg[1976]), .B(n11850), .Z(n3844) );
  NANDN U5273 ( .A(n11849), .B(n3844), .Z(n3845) );
  NAND U5274 ( .A(n3843), .B(n3845), .Z(n11858) );
  XOR U5275 ( .A(n11874), .B(sreg[1979]), .Z(n3846) );
  NANDN U5276 ( .A(n11875), .B(n3846), .Z(n3847) );
  NAND U5277 ( .A(n11874), .B(sreg[1979]), .Z(n3848) );
  AND U5278 ( .A(n3847), .B(n3848), .Z(n11881) );
  NAND U5279 ( .A(n11901), .B(sreg[1982]), .Z(n3849) );
  XOR U5280 ( .A(sreg[1982]), .B(n11901), .Z(n3850) );
  NANDN U5281 ( .A(n11900), .B(n3850), .Z(n3851) );
  NAND U5282 ( .A(n3849), .B(n3851), .Z(n11909) );
  XOR U5283 ( .A(n11925), .B(sreg[1985]), .Z(n3852) );
  NANDN U5284 ( .A(n11926), .B(n3852), .Z(n3853) );
  NAND U5285 ( .A(n11925), .B(sreg[1985]), .Z(n3854) );
  AND U5286 ( .A(n3853), .B(n3854), .Z(n11932) );
  NAND U5287 ( .A(n11949), .B(sreg[1988]), .Z(n3855) );
  XOR U5288 ( .A(sreg[1988]), .B(n11949), .Z(n3856) );
  NANDN U5289 ( .A(n11948), .B(n3856), .Z(n3857) );
  NAND U5290 ( .A(n3855), .B(n3857), .Z(n11957) );
  XOR U5291 ( .A(n11973), .B(sreg[1991]), .Z(n3858) );
  NANDN U5292 ( .A(n11974), .B(n3858), .Z(n3859) );
  NAND U5293 ( .A(n11973), .B(sreg[1991]), .Z(n3860) );
  AND U5294 ( .A(n3859), .B(n3860), .Z(n11980) );
  NAND U5295 ( .A(n11997), .B(sreg[1994]), .Z(n3861) );
  XOR U5296 ( .A(sreg[1994]), .B(n11997), .Z(n3862) );
  NANDN U5297 ( .A(n11996), .B(n3862), .Z(n3863) );
  NAND U5298 ( .A(n3861), .B(n3863), .Z(n12005) );
  NAND U5299 ( .A(n12023), .B(sreg[1997]), .Z(n3864) );
  XOR U5300 ( .A(sreg[1997]), .B(n12023), .Z(n3865) );
  NAND U5301 ( .A(n3865), .B(n12022), .Z(n3866) );
  NAND U5302 ( .A(n3864), .B(n3866), .Z(n12031) );
  NAND U5303 ( .A(n12048), .B(sreg[2000]), .Z(n3867) );
  XOR U5304 ( .A(sreg[2000]), .B(n12048), .Z(n3868) );
  NANDN U5305 ( .A(n12047), .B(n3868), .Z(n3869) );
  NAND U5306 ( .A(n3867), .B(n3869), .Z(n12056) );
  XOR U5307 ( .A(n12072), .B(sreg[2003]), .Z(n3870) );
  NANDN U5308 ( .A(n12073), .B(n3870), .Z(n3871) );
  NAND U5309 ( .A(n12072), .B(sreg[2003]), .Z(n3872) );
  AND U5310 ( .A(n3871), .B(n3872), .Z(n12079) );
  NAND U5311 ( .A(n12094), .B(sreg[2006]), .Z(n3873) );
  XOR U5312 ( .A(sreg[2006]), .B(n12094), .Z(n3874) );
  NAND U5313 ( .A(n3874), .B(n12093), .Z(n3875) );
  NAND U5314 ( .A(n3873), .B(n3875), .Z(n12102) );
  NAND U5315 ( .A(n12120), .B(sreg[2009]), .Z(n3876) );
  XOR U5316 ( .A(sreg[2009]), .B(n12120), .Z(n3877) );
  NAND U5317 ( .A(n3877), .B(n12119), .Z(n3878) );
  NAND U5318 ( .A(n3876), .B(n3878), .Z(n12126) );
  NAND U5319 ( .A(n12143), .B(sreg[2012]), .Z(n3879) );
  XOR U5320 ( .A(sreg[2012]), .B(n12143), .Z(n3880) );
  NANDN U5321 ( .A(n12142), .B(n3880), .Z(n3881) );
  NAND U5322 ( .A(n3879), .B(n3881), .Z(n12151) );
  XOR U5323 ( .A(n12167), .B(sreg[2015]), .Z(n3882) );
  NANDN U5324 ( .A(n12168), .B(n3882), .Z(n3883) );
  NAND U5325 ( .A(n12167), .B(sreg[2015]), .Z(n3884) );
  AND U5326 ( .A(n3883), .B(n3884), .Z(n12174) );
  NAND U5327 ( .A(n12191), .B(sreg[2018]), .Z(n3885) );
  XOR U5328 ( .A(sreg[2018]), .B(n12191), .Z(n3886) );
  NANDN U5329 ( .A(n12190), .B(n3886), .Z(n3887) );
  NAND U5330 ( .A(n3885), .B(n3887), .Z(n12199) );
  NAND U5331 ( .A(n12217), .B(sreg[2021]), .Z(n3888) );
  XOR U5332 ( .A(sreg[2021]), .B(n12217), .Z(n3889) );
  NAND U5333 ( .A(n3889), .B(n12216), .Z(n3890) );
  NAND U5334 ( .A(n3888), .B(n3890), .Z(n12223) );
  NAND U5335 ( .A(n12241), .B(sreg[2024]), .Z(n3891) );
  XOR U5336 ( .A(sreg[2024]), .B(n12241), .Z(n3892) );
  NANDN U5337 ( .A(n12242), .B(n3892), .Z(n3893) );
  NAND U5338 ( .A(n3891), .B(n3893), .Z(n12250) );
  XOR U5339 ( .A(n12266), .B(sreg[2027]), .Z(n3894) );
  NANDN U5340 ( .A(n12267), .B(n3894), .Z(n3895) );
  NAND U5341 ( .A(n12266), .B(sreg[2027]), .Z(n3896) );
  AND U5342 ( .A(n3895), .B(n3896), .Z(n12273) );
  NAND U5343 ( .A(n12289), .B(sreg[2030]), .Z(n3897) );
  XOR U5344 ( .A(sreg[2030]), .B(n12289), .Z(n3898) );
  NANDN U5345 ( .A(n12290), .B(n3898), .Z(n3899) );
  NAND U5346 ( .A(n3897), .B(n3899), .Z(n12298) );
  NAND U5347 ( .A(n12314), .B(sreg[2033]), .Z(n3900) );
  XOR U5348 ( .A(sreg[2033]), .B(n12314), .Z(n3901) );
  NANDN U5349 ( .A(n12315), .B(n3901), .Z(n3902) );
  NAND U5350 ( .A(n3900), .B(n3902), .Z(n12323) );
  NAND U5351 ( .A(n12340), .B(sreg[2036]), .Z(n3903) );
  XOR U5352 ( .A(sreg[2036]), .B(n12340), .Z(n3904) );
  NANDN U5353 ( .A(n12339), .B(n3904), .Z(n3905) );
  NAND U5354 ( .A(n3903), .B(n3905), .Z(n12348) );
  XOR U5355 ( .A(n12364), .B(sreg[2039]), .Z(n3906) );
  NANDN U5356 ( .A(n12365), .B(n3906), .Z(n3907) );
  NAND U5357 ( .A(n12364), .B(sreg[2039]), .Z(n3908) );
  AND U5358 ( .A(n3907), .B(n3908), .Z(n12371) );
  NAND U5359 ( .A(n12388), .B(sreg[2042]), .Z(n3909) );
  XOR U5360 ( .A(sreg[2042]), .B(n12388), .Z(n3910) );
  NANDN U5361 ( .A(n12387), .B(n3910), .Z(n3911) );
  NAND U5362 ( .A(n3909), .B(n3911), .Z(n12396) );
  NAND U5363 ( .A(n12416), .B(n12415), .Z(n3912) );
  XOR U5364 ( .A(n12415), .B(n12416), .Z(n3913) );
  NAND U5365 ( .A(n3913), .B(sreg[2045]), .Z(n3914) );
  NAND U5366 ( .A(n3912), .B(n3914), .Z(n12420) );
  IV U5367 ( .A(b[0]), .Z(n3915) );
  IV U5368 ( .A(b[0]), .Z(n3916) );
  IV U5369 ( .A(b[0]), .Z(n3917) );
  IV U5370 ( .A(b[0]), .Z(n3918) );
  IV U5371 ( .A(b[0]), .Z(n3919) );
  IV U5372 ( .A(b[0]), .Z(n3920) );
  IV U5373 ( .A(b[0]), .Z(n3921) );
  IV U5374 ( .A(b[0]), .Z(n3922) );
  IV U5375 ( .A(b[0]), .Z(n3923) );
  IV U5376 ( .A(b[0]), .Z(n3924) );
  IV U5377 ( .A(b[0]), .Z(n3925) );
  IV U5378 ( .A(b[0]), .Z(n3926) );
  IV U5379 ( .A(b[0]), .Z(n3927) );
  IV U5380 ( .A(b[0]), .Z(n3928) );
  IV U5381 ( .A(b[0]), .Z(n3929) );
  IV U5382 ( .A(b[0]), .Z(n3930) );
  IV U5383 ( .A(b[0]), .Z(n3931) );
  IV U5384 ( .A(b[0]), .Z(n3932) );
  IV U5385 ( .A(b[0]), .Z(n3933) );
  IV U5386 ( .A(b[0]), .Z(n3934) );
  IV U5387 ( .A(b[0]), .Z(n3935) );
  IV U5388 ( .A(b[0]), .Z(n3936) );
  IV U5389 ( .A(b[0]), .Z(n3937) );
  IV U5390 ( .A(b[0]), .Z(n3938) );
  IV U5391 ( .A(b[0]), .Z(n3939) );
  IV U5392 ( .A(b[0]), .Z(n3940) );
  IV U5393 ( .A(b[0]), .Z(n3941) );
  IV U5394 ( .A(b[0]), .Z(n3942) );
  IV U5395 ( .A(b[0]), .Z(n3943) );
  IV U5396 ( .A(b[0]), .Z(n3944) );
  IV U5397 ( .A(b[0]), .Z(n3945) );
  IV U5398 ( .A(b[0]), .Z(n3946) );
  IV U5399 ( .A(b[0]), .Z(n3947) );
  IV U5400 ( .A(b[0]), .Z(n3948) );
  IV U5401 ( .A(b[0]), .Z(n3949) );
  IV U5402 ( .A(b[0]), .Z(n3950) );
  IV U5403 ( .A(b[0]), .Z(n3951) );
  IV U5404 ( .A(b[0]), .Z(n3952) );
  IV U5405 ( .A(b[0]), .Z(n3953) );
  IV U5406 ( .A(b[0]), .Z(n3954) );
  IV U5407 ( .A(b[0]), .Z(n3955) );
  IV U5408 ( .A(b[0]), .Z(n3956) );
  IV U5409 ( .A(b[0]), .Z(n3957) );
  IV U5410 ( .A(b[0]), .Z(n3958) );
  IV U5411 ( .A(b[0]), .Z(n3959) );
  IV U5412 ( .A(b[0]), .Z(n3960) );
  IV U5413 ( .A(b[0]), .Z(n3961) );
  IV U5414 ( .A(b[0]), .Z(n3962) );
  IV U5415 ( .A(b[0]), .Z(n3963) );
  IV U5416 ( .A(b[0]), .Z(n3964) );
  IV U5417 ( .A(b[0]), .Z(n3965) );
  IV U5418 ( .A(b[0]), .Z(n3966) );
  IV U5419 ( .A(b[0]), .Z(n3967) );
  IV U5420 ( .A(b[0]), .Z(n3968) );
  IV U5421 ( .A(b[0]), .Z(n3969) );
  IV U5422 ( .A(b[0]), .Z(n3970) );
  IV U5423 ( .A(b[0]), .Z(n3971) );
  IV U5424 ( .A(b[0]), .Z(n3972) );
  IV U5425 ( .A(b[0]), .Z(n3973) );
  IV U5426 ( .A(b[0]), .Z(n3974) );
  IV U5427 ( .A(b[0]), .Z(n3975) );
  IV U5428 ( .A(b[0]), .Z(n3976) );
  IV U5429 ( .A(b[0]), .Z(n3977) );
  IV U5430 ( .A(b[0]), .Z(n3978) );
  IV U5431 ( .A(b[0]), .Z(n3979) );
  IV U5432 ( .A(b[0]), .Z(n3980) );
  IV U5433 ( .A(b[0]), .Z(n3981) );
  IV U5434 ( .A(b[0]), .Z(n3982) );
  IV U5435 ( .A(b[0]), .Z(n3983) );
  IV U5436 ( .A(b[0]), .Z(n3984) );
  IV U5437 ( .A(b[0]), .Z(n3985) );
  IV U5438 ( .A(b[0]), .Z(n3986) );
  IV U5439 ( .A(b[0]), .Z(n3987) );
  NANDN U5440 ( .A(n3915), .B(a[0]), .Z(n3988) );
  XNOR U5441 ( .A(sreg[1022]), .B(n3988), .Z(c[1022]) );
  NAND U5442 ( .A(b[1]), .B(a[0]), .Z(n3996) );
  NANDN U5443 ( .A(n3915), .B(a[1]), .Z(n3995) );
  XOR U5444 ( .A(n3996), .B(n3995), .Z(n3990) );
  XNOR U5445 ( .A(sreg[1023]), .B(n3990), .Z(n3992) );
  NANDN U5446 ( .A(n3988), .B(sreg[1022]), .Z(n3991) );
  XOR U5447 ( .A(n3992), .B(n3991), .Z(c[1023]) );
  AND U5448 ( .A(a[2]), .B(b[0]), .Z(n4008) );
  AND U5449 ( .A(a[1]), .B(n3988), .Z(n3989) );
  NAND U5450 ( .A(n3989), .B(b[1]), .Z(n3997) );
  XNOR U5451 ( .A(n4008), .B(n3997), .Z(n4002) );
  XNOR U5452 ( .A(sreg[1024]), .B(n4002), .Z(n4004) );
  NAND U5453 ( .A(sreg[1023]), .B(n3990), .Z(n3994) );
  OR U5454 ( .A(n3992), .B(n3991), .Z(n3993) );
  AND U5455 ( .A(n3994), .B(n3993), .Z(n4003) );
  XOR U5456 ( .A(n4004), .B(n4003), .Z(c[1024]) );
  OR U5457 ( .A(n3996), .B(n3995), .Z(n3999) );
  NANDN U5458 ( .A(n3997), .B(n4008), .Z(n3998) );
  NAND U5459 ( .A(n3999), .B(n3998), .Z(n4009) );
  ANDN U5460 ( .B(a[3]), .A(n3915), .Z(n4001) );
  NAND U5461 ( .A(b[1]), .B(a[2]), .Z(n4000) );
  XNOR U5462 ( .A(n4001), .B(n4000), .Z(n4010) );
  XOR U5463 ( .A(n4009), .B(n4010), .Z(n4014) );
  NAND U5464 ( .A(sreg[1024]), .B(n4002), .Z(n4006) );
  OR U5465 ( .A(n4004), .B(n4003), .Z(n4005) );
  AND U5466 ( .A(n4006), .B(n4005), .Z(n4013) );
  XNOR U5467 ( .A(n4013), .B(sreg[1025]), .Z(n4007) );
  XOR U5468 ( .A(n4014), .B(n4007), .Z(c[1025]) );
  NAND U5469 ( .A(b[1]), .B(a[3]), .Z(n4018) );
  AND U5470 ( .A(a[4]), .B(b[0]), .Z(n4028) );
  NANDN U5471 ( .A(n4018), .B(n4008), .Z(n4012) );
  NAND U5472 ( .A(n4010), .B(n4009), .Z(n4011) );
  NAND U5473 ( .A(n4012), .B(n4011), .Z(n4016) );
  XOR U5474 ( .A(n4028), .B(n4016), .Z(n4017) );
  XOR U5475 ( .A(n4018), .B(n4017), .Z(n4023) );
  XOR U5476 ( .A(n4022), .B(sreg[1026]), .Z(n4015) );
  XNOR U5477 ( .A(n4023), .B(n4015), .Z(c[1026]) );
  NAND U5478 ( .A(n4016), .B(n4028), .Z(n4020) );
  NANDN U5479 ( .A(n4018), .B(n4017), .Z(n4019) );
  NAND U5480 ( .A(n4020), .B(n4019), .Z(n4030) );
  ANDN U5481 ( .B(a[5]), .A(n3915), .Z(n4036) );
  NAND U5482 ( .A(b[1]), .B(a[4]), .Z(n4021) );
  XNOR U5483 ( .A(n4036), .B(n4021), .Z(n4031) );
  XOR U5484 ( .A(n4030), .B(n4031), .Z(n4026) );
  XOR U5485 ( .A(n4025), .B(sreg[1027]), .Z(n4024) );
  XOR U5486 ( .A(n4026), .B(n4024), .Z(c[1027]) );
  ANDN U5487 ( .B(a[6]), .A(n3915), .Z(n4048) );
  NAND U5488 ( .A(b[1]), .B(a[5]), .Z(n4027) );
  XOR U5489 ( .A(n4048), .B(n4027), .Z(n4039) );
  AND U5490 ( .A(a[5]), .B(b[1]), .Z(n4029) );
  NAND U5491 ( .A(n4029), .B(n4028), .Z(n4033) );
  NAND U5492 ( .A(n4031), .B(n4030), .Z(n4032) );
  NAND U5493 ( .A(n4033), .B(n4032), .Z(n4038) );
  XNOR U5494 ( .A(n4039), .B(n4038), .Z(n4042) );
  XNOR U5495 ( .A(sreg[1028]), .B(n4042), .Z(n4044) );
  XNOR U5496 ( .A(n4043), .B(n4044), .Z(c[1028]) );
  ANDN U5497 ( .B(a[7]), .A(n3915), .Z(n4035) );
  NAND U5498 ( .A(b[1]), .B(a[6]), .Z(n4034) );
  XOR U5499 ( .A(n4035), .B(n4034), .Z(n4050) );
  AND U5500 ( .A(a[6]), .B(b[1]), .Z(n4037) );
  NAND U5501 ( .A(n4037), .B(n4036), .Z(n4041) );
  NANDN U5502 ( .A(n4039), .B(n4038), .Z(n4040) );
  AND U5503 ( .A(n4041), .B(n4040), .Z(n4049) );
  XOR U5504 ( .A(n4050), .B(n4049), .Z(n4052) );
  NAND U5505 ( .A(sreg[1028]), .B(n4042), .Z(n4046) );
  NANDN U5506 ( .A(n4044), .B(n4043), .Z(n4045) );
  AND U5507 ( .A(n4046), .B(n4045), .Z(n4051) );
  XNOR U5508 ( .A(n4051), .B(sreg[1029]), .Z(n4047) );
  XOR U5509 ( .A(n4052), .B(n4047), .Z(c[1029]) );
  AND U5510 ( .A(a[7]), .B(b[1]), .Z(n4055) );
  NAND U5511 ( .A(b[0]), .B(a[8]), .Z(n4054) );
  XOR U5512 ( .A(n4055), .B(n4054), .Z(n4056) );
  XOR U5513 ( .A(n4057), .B(n4056), .Z(n4061) );
  XOR U5514 ( .A(sreg[1030]), .B(n4060), .Z(n4053) );
  XOR U5515 ( .A(n4061), .B(n4053), .Z(c[1030]) );
  NANDN U5516 ( .A(n4055), .B(n4054), .Z(n4059) );
  OR U5517 ( .A(n4057), .B(n4056), .Z(n4058) );
  NAND U5518 ( .A(n4059), .B(n4058), .Z(n4066) );
  ANDN U5519 ( .B(a[9]), .A(n3916), .Z(n4064) );
  AND U5520 ( .A(b[1]), .B(a[8]), .Z(n4063) );
  XOR U5521 ( .A(n4064), .B(n4063), .Z(n4065) );
  XNOR U5522 ( .A(n4066), .B(n4065), .Z(n4068) );
  XNOR U5523 ( .A(sreg[1031]), .B(n4067), .Z(n4062) );
  XNOR U5524 ( .A(n4068), .B(n4062), .Z(c[1031]) );
  NAND U5525 ( .A(b[0]), .B(a[10]), .Z(n4071) );
  NAND U5526 ( .A(a[9]), .B(b[1]), .Z(n4070) );
  XNOR U5527 ( .A(n4071), .B(n4070), .Z(n4073) );
  XNOR U5528 ( .A(n4072), .B(n4073), .Z(n4077) );
  XOR U5529 ( .A(n4076), .B(sreg[1032]), .Z(n4069) );
  XNOR U5530 ( .A(n4077), .B(n4069), .Z(c[1032]) );
  NAND U5531 ( .A(n4071), .B(n4070), .Z(n4075) );
  NANDN U5532 ( .A(n4073), .B(n4072), .Z(n4074) );
  NAND U5533 ( .A(n4075), .B(n4074), .Z(n4081) );
  NAND U5534 ( .A(b[0]), .B(a[11]), .Z(n4080) );
  NAND U5535 ( .A(a[10]), .B(b[1]), .Z(n4079) );
  XNOR U5536 ( .A(n4080), .B(n4079), .Z(n4082) );
  XNOR U5537 ( .A(n4081), .B(n4082), .Z(n4086) );
  XOR U5538 ( .A(n4085), .B(sreg[1033]), .Z(n4078) );
  XNOR U5539 ( .A(n4086), .B(n4078), .Z(c[1033]) );
  NAND U5540 ( .A(n4080), .B(n4079), .Z(n4084) );
  NANDN U5541 ( .A(n4082), .B(n4081), .Z(n4083) );
  NAND U5542 ( .A(n4084), .B(n4083), .Z(n4091) );
  ANDN U5543 ( .B(a[12]), .A(n3916), .Z(n4089) );
  AND U5544 ( .A(b[1]), .B(a[11]), .Z(n4088) );
  XOR U5545 ( .A(n4089), .B(n4088), .Z(n4090) );
  XNOR U5546 ( .A(n4091), .B(n4090), .Z(n4093) );
  XOR U5547 ( .A(sreg[1034]), .B(n4092), .Z(n4087) );
  XNOR U5548 ( .A(n4093), .B(n4087), .Z(c[1034]) );
  NAND U5549 ( .A(b[0]), .B(a[13]), .Z(n4096) );
  NAND U5550 ( .A(a[12]), .B(b[1]), .Z(n4095) );
  XNOR U5551 ( .A(n4096), .B(n4095), .Z(n4098) );
  XNOR U5552 ( .A(n4097), .B(n4098), .Z(n4102) );
  XOR U5553 ( .A(n4101), .B(sreg[1035]), .Z(n4094) );
  XNOR U5554 ( .A(n4102), .B(n4094), .Z(c[1035]) );
  NAND U5555 ( .A(n4096), .B(n4095), .Z(n4100) );
  NANDN U5556 ( .A(n4098), .B(n4097), .Z(n4099) );
  NAND U5557 ( .A(n4100), .B(n4099), .Z(n4107) );
  ANDN U5558 ( .B(a[14]), .A(n3916), .Z(n4105) );
  AND U5559 ( .A(b[1]), .B(a[13]), .Z(n4104) );
  XOR U5560 ( .A(n4105), .B(n4104), .Z(n4106) );
  XNOR U5561 ( .A(n4107), .B(n4106), .Z(n4109) );
  XOR U5562 ( .A(sreg[1036]), .B(n4108), .Z(n4103) );
  XNOR U5563 ( .A(n4109), .B(n4103), .Z(c[1036]) );
  NAND U5564 ( .A(b[0]), .B(a[15]), .Z(n4112) );
  NAND U5565 ( .A(a[14]), .B(b[1]), .Z(n4111) );
  XNOR U5566 ( .A(n4112), .B(n4111), .Z(n4114) );
  XNOR U5567 ( .A(n4113), .B(n4114), .Z(n4118) );
  XOR U5568 ( .A(n4117), .B(sreg[1037]), .Z(n4110) );
  XNOR U5569 ( .A(n4118), .B(n4110), .Z(c[1037]) );
  NAND U5570 ( .A(n4112), .B(n4111), .Z(n4116) );
  NANDN U5571 ( .A(n4114), .B(n4113), .Z(n4115) );
  NAND U5572 ( .A(n4116), .B(n4115), .Z(n4123) );
  ANDN U5573 ( .B(a[16]), .A(n3916), .Z(n4121) );
  AND U5574 ( .A(b[1]), .B(a[15]), .Z(n4120) );
  XOR U5575 ( .A(n4121), .B(n4120), .Z(n4122) );
  XNOR U5576 ( .A(n4123), .B(n4122), .Z(n4125) );
  XOR U5577 ( .A(sreg[1038]), .B(n4124), .Z(n4119) );
  XNOR U5578 ( .A(n4125), .B(n4119), .Z(c[1038]) );
  NAND U5579 ( .A(b[0]), .B(a[17]), .Z(n4128) );
  NAND U5580 ( .A(a[16]), .B(b[1]), .Z(n4127) );
  XNOR U5581 ( .A(n4128), .B(n4127), .Z(n4130) );
  XNOR U5582 ( .A(n4129), .B(n4130), .Z(n4134) );
  XOR U5583 ( .A(n4133), .B(sreg[1039]), .Z(n4126) );
  XNOR U5584 ( .A(n4134), .B(n4126), .Z(c[1039]) );
  NAND U5585 ( .A(n4128), .B(n4127), .Z(n4132) );
  NANDN U5586 ( .A(n4130), .B(n4129), .Z(n4131) );
  NAND U5587 ( .A(n4132), .B(n4131), .Z(n4139) );
  ANDN U5588 ( .B(a[18]), .A(n3916), .Z(n4137) );
  AND U5589 ( .A(b[1]), .B(a[17]), .Z(n4136) );
  XOR U5590 ( .A(n4137), .B(n4136), .Z(n4138) );
  XNOR U5591 ( .A(n4139), .B(n4138), .Z(n4141) );
  XOR U5592 ( .A(sreg[1040]), .B(n4140), .Z(n4135) );
  XNOR U5593 ( .A(n4141), .B(n4135), .Z(c[1040]) );
  ANDN U5594 ( .B(a[19]), .A(n3916), .Z(n4144) );
  AND U5595 ( .A(b[1]), .B(a[18]), .Z(n4143) );
  XOR U5596 ( .A(n4144), .B(n4143), .Z(n4145) );
  XOR U5597 ( .A(n4146), .B(n4145), .Z(n4152) );
  IV U5598 ( .A(n4150), .Z(n4149) );
  XOR U5599 ( .A(n4149), .B(sreg[1041]), .Z(n4142) );
  XOR U5600 ( .A(n4152), .B(n4142), .Z(c[1041]) );
  OR U5601 ( .A(n4144), .B(n4143), .Z(n4148) );
  NAND U5602 ( .A(n4146), .B(n4145), .Z(n4147) );
  NAND U5603 ( .A(n4148), .B(n4147), .Z(n4159) );
  ANDN U5604 ( .B(a[20]), .A(n3916), .Z(n4157) );
  AND U5605 ( .A(b[1]), .B(a[19]), .Z(n4156) );
  XOR U5606 ( .A(n4157), .B(n4156), .Z(n4158) );
  XNOR U5607 ( .A(n4159), .B(n4158), .Z(n4161) );
  NANDN U5608 ( .A(n4149), .B(sreg[1041]), .Z(n4154) );
  OR U5609 ( .A(sreg[1041]), .B(n4150), .Z(n4151) );
  NANDN U5610 ( .A(n4152), .B(n4151), .Z(n4153) );
  NAND U5611 ( .A(n4154), .B(n4153), .Z(n4160) );
  XNOR U5612 ( .A(sreg[1042]), .B(n4160), .Z(n4155) );
  XNOR U5613 ( .A(n4161), .B(n4155), .Z(c[1042]) );
  ANDN U5614 ( .B(a[21]), .A(n3917), .Z(n4164) );
  AND U5615 ( .A(b[1]), .B(a[20]), .Z(n4163) );
  XOR U5616 ( .A(n4164), .B(n4163), .Z(n4165) );
  XNOR U5617 ( .A(n4166), .B(n4165), .Z(n4168) );
  XNOR U5618 ( .A(sreg[1043]), .B(n4167), .Z(n4162) );
  XNOR U5619 ( .A(n4168), .B(n4162), .Z(c[1043]) );
  ANDN U5620 ( .B(a[22]), .A(n3917), .Z(n4171) );
  AND U5621 ( .A(b[1]), .B(a[21]), .Z(n4170) );
  XOR U5622 ( .A(n4171), .B(n4170), .Z(n4172) );
  XNOR U5623 ( .A(n4173), .B(n4172), .Z(n4175) );
  XNOR U5624 ( .A(sreg[1044]), .B(n4174), .Z(n4169) );
  XNOR U5625 ( .A(n4175), .B(n4169), .Z(c[1044]) );
  NAND U5626 ( .A(b[0]), .B(a[23]), .Z(n4178) );
  NAND U5627 ( .A(a[22]), .B(b[1]), .Z(n4177) );
  XNOR U5628 ( .A(n4178), .B(n4177), .Z(n4180) );
  XNOR U5629 ( .A(n4179), .B(n4180), .Z(n4184) );
  XOR U5630 ( .A(n4183), .B(sreg[1045]), .Z(n4176) );
  XNOR U5631 ( .A(n4184), .B(n4176), .Z(c[1045]) );
  NAND U5632 ( .A(n4178), .B(n4177), .Z(n4182) );
  NANDN U5633 ( .A(n4180), .B(n4179), .Z(n4181) );
  NAND U5634 ( .A(n4182), .B(n4181), .Z(n4189) );
  ANDN U5635 ( .B(a[24]), .A(n3917), .Z(n4187) );
  AND U5636 ( .A(b[1]), .B(a[23]), .Z(n4186) );
  XOR U5637 ( .A(n4187), .B(n4186), .Z(n4188) );
  XOR U5638 ( .A(n4189), .B(n4188), .Z(n4193) );
  XNOR U5639 ( .A(n4192), .B(sreg[1046]), .Z(n4185) );
  XOR U5640 ( .A(n4193), .B(n4185), .Z(c[1046]) );
  OR U5641 ( .A(n4187), .B(n4186), .Z(n4191) );
  NAND U5642 ( .A(n4189), .B(n4188), .Z(n4190) );
  NAND U5643 ( .A(n4191), .B(n4190), .Z(n4197) );
  NAND U5644 ( .A(b[0]), .B(a[25]), .Z(n4196) );
  NAND U5645 ( .A(a[24]), .B(b[1]), .Z(n4195) );
  XNOR U5646 ( .A(n4196), .B(n4195), .Z(n4198) );
  XNOR U5647 ( .A(n4197), .B(n4198), .Z(n4202) );
  XNOR U5648 ( .A(n4201), .B(sreg[1047]), .Z(n4194) );
  XNOR U5649 ( .A(n4202), .B(n4194), .Z(c[1047]) );
  NAND U5650 ( .A(n4196), .B(n4195), .Z(n4200) );
  NANDN U5651 ( .A(n4198), .B(n4197), .Z(n4199) );
  NAND U5652 ( .A(n4200), .B(n4199), .Z(n4207) );
  ANDN U5653 ( .B(a[26]), .A(n3917), .Z(n4205) );
  AND U5654 ( .A(b[1]), .B(a[25]), .Z(n4204) );
  XOR U5655 ( .A(n4205), .B(n4204), .Z(n4206) );
  XNOR U5656 ( .A(n4207), .B(n4206), .Z(n4209) );
  XOR U5657 ( .A(sreg[1048]), .B(n4208), .Z(n4203) );
  XNOR U5658 ( .A(n4209), .B(n4203), .Z(c[1048]) );
  ANDN U5659 ( .B(a[27]), .A(n3917), .Z(n4212) );
  AND U5660 ( .A(b[1]), .B(a[26]), .Z(n4211) );
  XOR U5661 ( .A(n4212), .B(n4211), .Z(n4213) );
  XOR U5662 ( .A(n4214), .B(n4213), .Z(n4220) );
  IV U5663 ( .A(n4218), .Z(n4217) );
  XOR U5664 ( .A(n4217), .B(sreg[1049]), .Z(n4210) );
  XOR U5665 ( .A(n4220), .B(n4210), .Z(c[1049]) );
  OR U5666 ( .A(n4212), .B(n4211), .Z(n4216) );
  NAND U5667 ( .A(n4214), .B(n4213), .Z(n4215) );
  NAND U5668 ( .A(n4216), .B(n4215), .Z(n4227) );
  ANDN U5669 ( .B(a[28]), .A(n3917), .Z(n4225) );
  AND U5670 ( .A(b[1]), .B(a[27]), .Z(n4224) );
  XOR U5671 ( .A(n4225), .B(n4224), .Z(n4226) );
  XNOR U5672 ( .A(n4227), .B(n4226), .Z(n4229) );
  NANDN U5673 ( .A(n4217), .B(sreg[1049]), .Z(n4222) );
  OR U5674 ( .A(sreg[1049]), .B(n4218), .Z(n4219) );
  NANDN U5675 ( .A(n4220), .B(n4219), .Z(n4221) );
  NAND U5676 ( .A(n4222), .B(n4221), .Z(n4228) );
  XNOR U5677 ( .A(sreg[1050]), .B(n4228), .Z(n4223) );
  XNOR U5678 ( .A(n4229), .B(n4223), .Z(c[1050]) );
  NAND U5679 ( .A(b[0]), .B(a[29]), .Z(n4232) );
  NAND U5680 ( .A(a[28]), .B(b[1]), .Z(n4231) );
  XNOR U5681 ( .A(n4232), .B(n4231), .Z(n4234) );
  XNOR U5682 ( .A(n4233), .B(n4234), .Z(n4238) );
  XOR U5683 ( .A(n4237), .B(sreg[1051]), .Z(n4230) );
  XNOR U5684 ( .A(n4238), .B(n4230), .Z(c[1051]) );
  NAND U5685 ( .A(n4232), .B(n4231), .Z(n4236) );
  NANDN U5686 ( .A(n4234), .B(n4233), .Z(n4235) );
  NAND U5687 ( .A(n4236), .B(n4235), .Z(n4243) );
  ANDN U5688 ( .B(a[30]), .A(n3917), .Z(n4241) );
  AND U5689 ( .A(b[1]), .B(a[29]), .Z(n4240) );
  XOR U5690 ( .A(n4241), .B(n4240), .Z(n4242) );
  XNOR U5691 ( .A(n4243), .B(n4242), .Z(n4245) );
  XOR U5692 ( .A(sreg[1052]), .B(n4244), .Z(n4239) );
  XNOR U5693 ( .A(n4245), .B(n4239), .Z(c[1052]) );
  NAND U5694 ( .A(b[0]), .B(a[31]), .Z(n4248) );
  NAND U5695 ( .A(a[30]), .B(b[1]), .Z(n4247) );
  XNOR U5696 ( .A(n4248), .B(n4247), .Z(n4250) );
  XNOR U5697 ( .A(n4249), .B(n4250), .Z(n4254) );
  XOR U5698 ( .A(n4253), .B(sreg[1053]), .Z(n4246) );
  XNOR U5699 ( .A(n4254), .B(n4246), .Z(c[1053]) );
  NAND U5700 ( .A(n4248), .B(n4247), .Z(n4252) );
  NANDN U5701 ( .A(n4250), .B(n4249), .Z(n4251) );
  NAND U5702 ( .A(n4252), .B(n4251), .Z(n4259) );
  ANDN U5703 ( .B(a[32]), .A(n3918), .Z(n4257) );
  AND U5704 ( .A(b[1]), .B(a[31]), .Z(n4256) );
  XOR U5705 ( .A(n4257), .B(n4256), .Z(n4258) );
  XNOR U5706 ( .A(n4259), .B(n4258), .Z(n4264) );
  XOR U5707 ( .A(sreg[1054]), .B(n4263), .Z(n4255) );
  XNOR U5708 ( .A(n4264), .B(n4255), .Z(c[1054]) );
  OR U5709 ( .A(n4257), .B(n4256), .Z(n4262) );
  IV U5710 ( .A(n4258), .Z(n4260) );
  NANDN U5711 ( .A(n4260), .B(n4259), .Z(n4261) );
  NAND U5712 ( .A(n4262), .B(n4261), .Z(n4268) );
  NAND U5713 ( .A(b[0]), .B(a[33]), .Z(n4267) );
  NAND U5714 ( .A(a[32]), .B(b[1]), .Z(n4266) );
  XNOR U5715 ( .A(n4267), .B(n4266), .Z(n4269) );
  XNOR U5716 ( .A(n4268), .B(n4269), .Z(n4273) );
  XOR U5717 ( .A(n4272), .B(sreg[1055]), .Z(n4265) );
  XNOR U5718 ( .A(n4273), .B(n4265), .Z(c[1055]) );
  NAND U5719 ( .A(n4267), .B(n4266), .Z(n4271) );
  NANDN U5720 ( .A(n4269), .B(n4268), .Z(n4270) );
  NAND U5721 ( .A(n4271), .B(n4270), .Z(n4278) );
  ANDN U5722 ( .B(a[34]), .A(n3918), .Z(n4276) );
  AND U5723 ( .A(b[1]), .B(a[33]), .Z(n4275) );
  XOR U5724 ( .A(n4276), .B(n4275), .Z(n4277) );
  XNOR U5725 ( .A(n4278), .B(n4277), .Z(n4280) );
  XOR U5726 ( .A(sreg[1056]), .B(n4279), .Z(n4274) );
  XNOR U5727 ( .A(n4280), .B(n4274), .Z(c[1056]) );
  NAND U5728 ( .A(b[0]), .B(a[35]), .Z(n4283) );
  NAND U5729 ( .A(a[34]), .B(b[1]), .Z(n4282) );
  XNOR U5730 ( .A(n4283), .B(n4282), .Z(n4285) );
  XNOR U5731 ( .A(n4284), .B(n4285), .Z(n4289) );
  XOR U5732 ( .A(n4288), .B(sreg[1057]), .Z(n4281) );
  XNOR U5733 ( .A(n4289), .B(n4281), .Z(c[1057]) );
  NAND U5734 ( .A(n4283), .B(n4282), .Z(n4287) );
  NANDN U5735 ( .A(n4285), .B(n4284), .Z(n4286) );
  NAND U5736 ( .A(n4287), .B(n4286), .Z(n4294) );
  ANDN U5737 ( .B(a[36]), .A(n3918), .Z(n4292) );
  AND U5738 ( .A(b[1]), .B(a[35]), .Z(n4291) );
  XOR U5739 ( .A(n4292), .B(n4291), .Z(n4293) );
  XNOR U5740 ( .A(n4294), .B(n4293), .Z(n4296) );
  XOR U5741 ( .A(sreg[1058]), .B(n4295), .Z(n4290) );
  XNOR U5742 ( .A(n4296), .B(n4290), .Z(c[1058]) );
  NAND U5743 ( .A(b[0]), .B(a[37]), .Z(n4299) );
  NAND U5744 ( .A(a[36]), .B(b[1]), .Z(n4298) );
  XNOR U5745 ( .A(n4299), .B(n4298), .Z(n4301) );
  XNOR U5746 ( .A(n4300), .B(n4301), .Z(n4305) );
  XOR U5747 ( .A(n4304), .B(sreg[1059]), .Z(n4297) );
  XNOR U5748 ( .A(n4305), .B(n4297), .Z(c[1059]) );
  NAND U5749 ( .A(n4299), .B(n4298), .Z(n4303) );
  NANDN U5750 ( .A(n4301), .B(n4300), .Z(n4302) );
  NAND U5751 ( .A(n4303), .B(n4302), .Z(n4310) );
  ANDN U5752 ( .B(a[38]), .A(n3918), .Z(n4308) );
  AND U5753 ( .A(b[1]), .B(a[37]), .Z(n4307) );
  XOR U5754 ( .A(n4308), .B(n4307), .Z(n4309) );
  XNOR U5755 ( .A(n4310), .B(n4309), .Z(n4312) );
  XOR U5756 ( .A(sreg[1060]), .B(n4311), .Z(n4306) );
  XNOR U5757 ( .A(n4312), .B(n4306), .Z(c[1060]) );
  NAND U5758 ( .A(b[0]), .B(a[39]), .Z(n4315) );
  NAND U5759 ( .A(a[38]), .B(b[1]), .Z(n4314) );
  XNOR U5760 ( .A(n4315), .B(n4314), .Z(n4317) );
  XNOR U5761 ( .A(n4316), .B(n4317), .Z(n4321) );
  XOR U5762 ( .A(n4320), .B(sreg[1061]), .Z(n4313) );
  XNOR U5763 ( .A(n4321), .B(n4313), .Z(c[1061]) );
  NAND U5764 ( .A(n4315), .B(n4314), .Z(n4319) );
  NANDN U5765 ( .A(n4317), .B(n4316), .Z(n4318) );
  NAND U5766 ( .A(n4319), .B(n4318), .Z(n4326) );
  ANDN U5767 ( .B(a[40]), .A(n3918), .Z(n4324) );
  AND U5768 ( .A(b[1]), .B(a[39]), .Z(n4323) );
  XOR U5769 ( .A(n4324), .B(n4323), .Z(n4325) );
  XNOR U5770 ( .A(n4326), .B(n4325), .Z(n4328) );
  XOR U5771 ( .A(sreg[1062]), .B(n4327), .Z(n4322) );
  XNOR U5772 ( .A(n4328), .B(n4322), .Z(c[1062]) );
  NAND U5773 ( .A(b[0]), .B(a[41]), .Z(n4331) );
  NAND U5774 ( .A(a[40]), .B(b[1]), .Z(n4330) );
  XNOR U5775 ( .A(n4331), .B(n4330), .Z(n4333) );
  XNOR U5776 ( .A(n4332), .B(n4333), .Z(n4337) );
  XOR U5777 ( .A(n4336), .B(sreg[1063]), .Z(n4329) );
  XNOR U5778 ( .A(n4337), .B(n4329), .Z(c[1063]) );
  NAND U5779 ( .A(n4331), .B(n4330), .Z(n4335) );
  NANDN U5780 ( .A(n4333), .B(n4332), .Z(n4334) );
  NAND U5781 ( .A(n4335), .B(n4334), .Z(n4342) );
  ANDN U5782 ( .B(a[42]), .A(n3918), .Z(n4340) );
  AND U5783 ( .A(b[1]), .B(a[41]), .Z(n4339) );
  XOR U5784 ( .A(n4340), .B(n4339), .Z(n4341) );
  XNOR U5785 ( .A(n4342), .B(n4341), .Z(n4344) );
  XOR U5786 ( .A(sreg[1064]), .B(n4343), .Z(n4338) );
  XNOR U5787 ( .A(n4344), .B(n4338), .Z(c[1064]) );
  ANDN U5788 ( .B(a[43]), .A(n3918), .Z(n4347) );
  AND U5789 ( .A(b[1]), .B(a[42]), .Z(n4346) );
  XOR U5790 ( .A(n4347), .B(n4346), .Z(n4348) );
  XNOR U5791 ( .A(n4349), .B(n4348), .Z(n4351) );
  XNOR U5792 ( .A(sreg[1065]), .B(n4350), .Z(n4345) );
  XNOR U5793 ( .A(n4351), .B(n4345), .Z(c[1065]) );
  ANDN U5794 ( .B(a[44]), .A(n3919), .Z(n4354) );
  AND U5795 ( .A(b[1]), .B(a[43]), .Z(n4353) );
  XOR U5796 ( .A(n4354), .B(n4353), .Z(n4355) );
  XNOR U5797 ( .A(n4356), .B(n4355), .Z(n4361) );
  XNOR U5798 ( .A(sreg[1066]), .B(n4360), .Z(n4352) );
  XNOR U5799 ( .A(n4361), .B(n4352), .Z(c[1066]) );
  OR U5800 ( .A(n4354), .B(n4353), .Z(n4359) );
  IV U5801 ( .A(n4355), .Z(n4357) );
  NANDN U5802 ( .A(n4357), .B(n4356), .Z(n4358) );
  NAND U5803 ( .A(n4359), .B(n4358), .Z(n4365) );
  NAND U5804 ( .A(b[0]), .B(a[45]), .Z(n4364) );
  NAND U5805 ( .A(a[44]), .B(b[1]), .Z(n4363) );
  XNOR U5806 ( .A(n4364), .B(n4363), .Z(n4366) );
  XNOR U5807 ( .A(n4365), .B(n4366), .Z(n4370) );
  XOR U5808 ( .A(n4369), .B(sreg[1067]), .Z(n4362) );
  XNOR U5809 ( .A(n4370), .B(n4362), .Z(c[1067]) );
  NAND U5810 ( .A(n4364), .B(n4363), .Z(n4368) );
  NANDN U5811 ( .A(n4366), .B(n4365), .Z(n4367) );
  NAND U5812 ( .A(n4368), .B(n4367), .Z(n4374) );
  NAND U5813 ( .A(b[0]), .B(a[46]), .Z(n4373) );
  NAND U5814 ( .A(a[45]), .B(b[1]), .Z(n4372) );
  XNOR U5815 ( .A(n4373), .B(n4372), .Z(n4375) );
  XNOR U5816 ( .A(n4374), .B(n4375), .Z(n4379) );
  XOR U5817 ( .A(n4378), .B(sreg[1068]), .Z(n4371) );
  XNOR U5818 ( .A(n4379), .B(n4371), .Z(c[1068]) );
  NAND U5819 ( .A(n4373), .B(n4372), .Z(n4377) );
  NANDN U5820 ( .A(n4375), .B(n4374), .Z(n4376) );
  NAND U5821 ( .A(n4377), .B(n4376), .Z(n4383) );
  NAND U5822 ( .A(b[0]), .B(a[47]), .Z(n4382) );
  NAND U5823 ( .A(a[46]), .B(b[1]), .Z(n4381) );
  XNOR U5824 ( .A(n4382), .B(n4381), .Z(n4384) );
  XNOR U5825 ( .A(n4383), .B(n4384), .Z(n4388) );
  XOR U5826 ( .A(n4387), .B(sreg[1069]), .Z(n4380) );
  XNOR U5827 ( .A(n4388), .B(n4380), .Z(c[1069]) );
  NAND U5828 ( .A(n4382), .B(n4381), .Z(n4386) );
  NANDN U5829 ( .A(n4384), .B(n4383), .Z(n4385) );
  NAND U5830 ( .A(n4386), .B(n4385), .Z(n4393) );
  ANDN U5831 ( .B(a[48]), .A(n3919), .Z(n4391) );
  AND U5832 ( .A(b[1]), .B(a[47]), .Z(n4390) );
  XOR U5833 ( .A(n4391), .B(n4390), .Z(n4392) );
  XNOR U5834 ( .A(n4393), .B(n4392), .Z(n4395) );
  XOR U5835 ( .A(sreg[1070]), .B(n4394), .Z(n4389) );
  XNOR U5836 ( .A(n4395), .B(n4389), .Z(c[1070]) );
  NAND U5837 ( .A(b[0]), .B(a[49]), .Z(n4398) );
  NAND U5838 ( .A(a[48]), .B(b[1]), .Z(n4397) );
  XNOR U5839 ( .A(n4398), .B(n4397), .Z(n4400) );
  XNOR U5840 ( .A(n4399), .B(n4400), .Z(n4404) );
  XOR U5841 ( .A(n4403), .B(sreg[1071]), .Z(n4396) );
  XNOR U5842 ( .A(n4404), .B(n4396), .Z(c[1071]) );
  NAND U5843 ( .A(n4398), .B(n4397), .Z(n4402) );
  NANDN U5844 ( .A(n4400), .B(n4399), .Z(n4401) );
  NAND U5845 ( .A(n4402), .B(n4401), .Z(n4409) );
  ANDN U5846 ( .B(a[50]), .A(n3919), .Z(n4407) );
  AND U5847 ( .A(b[1]), .B(a[49]), .Z(n4406) );
  XOR U5848 ( .A(n4407), .B(n4406), .Z(n4408) );
  XNOR U5849 ( .A(n4409), .B(n4408), .Z(n4411) );
  XOR U5850 ( .A(sreg[1072]), .B(n4410), .Z(n4405) );
  XNOR U5851 ( .A(n4411), .B(n4405), .Z(c[1072]) );
  NAND U5852 ( .A(b[0]), .B(a[51]), .Z(n4414) );
  NAND U5853 ( .A(a[50]), .B(b[1]), .Z(n4413) );
  XNOR U5854 ( .A(n4414), .B(n4413), .Z(n4416) );
  XNOR U5855 ( .A(n4415), .B(n4416), .Z(n4420) );
  XOR U5856 ( .A(n4419), .B(sreg[1073]), .Z(n4412) );
  XNOR U5857 ( .A(n4420), .B(n4412), .Z(c[1073]) );
  NAND U5858 ( .A(n4414), .B(n4413), .Z(n4418) );
  NANDN U5859 ( .A(n4416), .B(n4415), .Z(n4417) );
  NAND U5860 ( .A(n4418), .B(n4417), .Z(n4425) );
  ANDN U5861 ( .B(a[52]), .A(n3919), .Z(n4423) );
  AND U5862 ( .A(b[1]), .B(a[51]), .Z(n4422) );
  XOR U5863 ( .A(n4423), .B(n4422), .Z(n4424) );
  XNOR U5864 ( .A(n4425), .B(n4424), .Z(n4427) );
  XOR U5865 ( .A(sreg[1074]), .B(n4426), .Z(n4421) );
  XNOR U5866 ( .A(n4427), .B(n4421), .Z(c[1074]) );
  ANDN U5867 ( .B(a[53]), .A(n3919), .Z(n4430) );
  AND U5868 ( .A(b[1]), .B(a[52]), .Z(n4429) );
  XOR U5869 ( .A(n4430), .B(n4429), .Z(n4431) );
  XNOR U5870 ( .A(n4432), .B(n4431), .Z(n4434) );
  XNOR U5871 ( .A(sreg[1075]), .B(n4433), .Z(n4428) );
  XNOR U5872 ( .A(n4434), .B(n4428), .Z(c[1075]) );
  ANDN U5873 ( .B(a[54]), .A(n3919), .Z(n4437) );
  AND U5874 ( .A(b[1]), .B(a[53]), .Z(n4436) );
  XOR U5875 ( .A(n4437), .B(n4436), .Z(n4438) );
  XNOR U5876 ( .A(n4439), .B(n4438), .Z(n4441) );
  XNOR U5877 ( .A(sreg[1076]), .B(n4440), .Z(n4435) );
  XNOR U5878 ( .A(n4441), .B(n4435), .Z(c[1076]) );
  NAND U5879 ( .A(b[0]), .B(a[55]), .Z(n4444) );
  NAND U5880 ( .A(a[54]), .B(b[1]), .Z(n4443) );
  XNOR U5881 ( .A(n4444), .B(n4443), .Z(n4446) );
  XNOR U5882 ( .A(n4445), .B(n4446), .Z(n4450) );
  XOR U5883 ( .A(n4449), .B(sreg[1077]), .Z(n4442) );
  XNOR U5884 ( .A(n4450), .B(n4442), .Z(c[1077]) );
  NAND U5885 ( .A(n4444), .B(n4443), .Z(n4448) );
  NANDN U5886 ( .A(n4446), .B(n4445), .Z(n4447) );
  NAND U5887 ( .A(n4448), .B(n4447), .Z(n4455) );
  ANDN U5888 ( .B(a[56]), .A(n3919), .Z(n4453) );
  AND U5889 ( .A(b[1]), .B(a[55]), .Z(n4452) );
  XOR U5890 ( .A(n4453), .B(n4452), .Z(n4454) );
  XNOR U5891 ( .A(n4455), .B(n4454), .Z(n4457) );
  XOR U5892 ( .A(sreg[1078]), .B(n4456), .Z(n4451) );
  XNOR U5893 ( .A(n4457), .B(n4451), .Z(c[1078]) );
  NAND U5894 ( .A(b[0]), .B(a[57]), .Z(n4460) );
  NAND U5895 ( .A(a[56]), .B(b[1]), .Z(n4459) );
  XNOR U5896 ( .A(n4460), .B(n4459), .Z(n4462) );
  XNOR U5897 ( .A(n4461), .B(n4462), .Z(n4466) );
  XOR U5898 ( .A(n4465), .B(sreg[1079]), .Z(n4458) );
  XNOR U5899 ( .A(n4466), .B(n4458), .Z(c[1079]) );
  NAND U5900 ( .A(n4460), .B(n4459), .Z(n4464) );
  NANDN U5901 ( .A(n4462), .B(n4461), .Z(n4463) );
  NAND U5902 ( .A(n4464), .B(n4463), .Z(n4471) );
  ANDN U5903 ( .B(a[58]), .A(n3920), .Z(n4469) );
  AND U5904 ( .A(b[1]), .B(a[57]), .Z(n4468) );
  XOR U5905 ( .A(n4469), .B(n4468), .Z(n4470) );
  XNOR U5906 ( .A(n4471), .B(n4470), .Z(n4476) );
  XOR U5907 ( .A(sreg[1080]), .B(n4475), .Z(n4467) );
  XNOR U5908 ( .A(n4476), .B(n4467), .Z(c[1080]) );
  OR U5909 ( .A(n4469), .B(n4468), .Z(n4474) );
  IV U5910 ( .A(n4470), .Z(n4472) );
  NANDN U5911 ( .A(n4472), .B(n4471), .Z(n4473) );
  NAND U5912 ( .A(n4474), .B(n4473), .Z(n4480) );
  NAND U5913 ( .A(b[0]), .B(a[59]), .Z(n4479) );
  NAND U5914 ( .A(a[58]), .B(b[1]), .Z(n4478) );
  XNOR U5915 ( .A(n4479), .B(n4478), .Z(n4481) );
  XNOR U5916 ( .A(n4480), .B(n4481), .Z(n4485) );
  XOR U5917 ( .A(n4484), .B(sreg[1081]), .Z(n4477) );
  XNOR U5918 ( .A(n4485), .B(n4477), .Z(c[1081]) );
  NAND U5919 ( .A(n4479), .B(n4478), .Z(n4483) );
  NANDN U5920 ( .A(n4481), .B(n4480), .Z(n4482) );
  NAND U5921 ( .A(n4483), .B(n4482), .Z(n4490) );
  ANDN U5922 ( .B(a[60]), .A(n3920), .Z(n4488) );
  AND U5923 ( .A(b[1]), .B(a[59]), .Z(n4487) );
  XOR U5924 ( .A(n4488), .B(n4487), .Z(n4489) );
  XNOR U5925 ( .A(n4490), .B(n4489), .Z(n4492) );
  XOR U5926 ( .A(sreg[1082]), .B(n4491), .Z(n4486) );
  XNOR U5927 ( .A(n4492), .B(n4486), .Z(c[1082]) );
  NAND U5928 ( .A(b[0]), .B(a[61]), .Z(n4495) );
  NAND U5929 ( .A(a[60]), .B(b[1]), .Z(n4494) );
  XNOR U5930 ( .A(n4495), .B(n4494), .Z(n4497) );
  XNOR U5931 ( .A(n4496), .B(n4497), .Z(n4501) );
  XOR U5932 ( .A(n4500), .B(sreg[1083]), .Z(n4493) );
  XNOR U5933 ( .A(n4501), .B(n4493), .Z(c[1083]) );
  NAND U5934 ( .A(n4495), .B(n4494), .Z(n4499) );
  NANDN U5935 ( .A(n4497), .B(n4496), .Z(n4498) );
  NAND U5936 ( .A(n4499), .B(n4498), .Z(n4505) );
  NAND U5937 ( .A(b[0]), .B(a[62]), .Z(n4504) );
  NAND U5938 ( .A(a[61]), .B(b[1]), .Z(n4503) );
  XNOR U5939 ( .A(n4504), .B(n4503), .Z(n4506) );
  XNOR U5940 ( .A(n4505), .B(n4506), .Z(n4510) );
  XOR U5941 ( .A(n4509), .B(sreg[1084]), .Z(n4502) );
  XNOR U5942 ( .A(n4510), .B(n4502), .Z(c[1084]) );
  NAND U5943 ( .A(n4504), .B(n4503), .Z(n4508) );
  NANDN U5944 ( .A(n4506), .B(n4505), .Z(n4507) );
  NAND U5945 ( .A(n4508), .B(n4507), .Z(n4514) );
  NAND U5946 ( .A(b[0]), .B(a[63]), .Z(n4513) );
  NAND U5947 ( .A(a[62]), .B(b[1]), .Z(n4512) );
  XNOR U5948 ( .A(n4513), .B(n4512), .Z(n4515) );
  XNOR U5949 ( .A(n4514), .B(n4515), .Z(n4519) );
  XOR U5950 ( .A(n4518), .B(sreg[1085]), .Z(n4511) );
  XNOR U5951 ( .A(n4519), .B(n4511), .Z(c[1085]) );
  NAND U5952 ( .A(n4513), .B(n4512), .Z(n4517) );
  NANDN U5953 ( .A(n4515), .B(n4514), .Z(n4516) );
  NAND U5954 ( .A(n4517), .B(n4516), .Z(n4524) );
  ANDN U5955 ( .B(a[64]), .A(n3920), .Z(n4522) );
  AND U5956 ( .A(b[1]), .B(a[63]), .Z(n4521) );
  XOR U5957 ( .A(n4522), .B(n4521), .Z(n4523) );
  XNOR U5958 ( .A(n4524), .B(n4523), .Z(n4526) );
  XOR U5959 ( .A(sreg[1086]), .B(n4525), .Z(n4520) );
  XNOR U5960 ( .A(n4526), .B(n4520), .Z(c[1086]) );
  NAND U5961 ( .A(b[0]), .B(a[65]), .Z(n4529) );
  NAND U5962 ( .A(a[64]), .B(b[1]), .Z(n4528) );
  XNOR U5963 ( .A(n4529), .B(n4528), .Z(n4531) );
  XNOR U5964 ( .A(n4530), .B(n4531), .Z(n4535) );
  XOR U5965 ( .A(n4534), .B(sreg[1087]), .Z(n4527) );
  XNOR U5966 ( .A(n4535), .B(n4527), .Z(c[1087]) );
  NAND U5967 ( .A(n4529), .B(n4528), .Z(n4533) );
  NANDN U5968 ( .A(n4531), .B(n4530), .Z(n4532) );
  NAND U5969 ( .A(n4533), .B(n4532), .Z(n4539) );
  NAND U5970 ( .A(b[0]), .B(a[66]), .Z(n4538) );
  NAND U5971 ( .A(a[65]), .B(b[1]), .Z(n4537) );
  XNOR U5972 ( .A(n4538), .B(n4537), .Z(n4540) );
  XNOR U5973 ( .A(n4539), .B(n4540), .Z(n4544) );
  XOR U5974 ( .A(n4543), .B(sreg[1088]), .Z(n4536) );
  XNOR U5975 ( .A(n4544), .B(n4536), .Z(c[1088]) );
  NAND U5976 ( .A(n4538), .B(n4537), .Z(n4542) );
  NANDN U5977 ( .A(n4540), .B(n4539), .Z(n4541) );
  NAND U5978 ( .A(n4542), .B(n4541), .Z(n4548) );
  NAND U5979 ( .A(b[0]), .B(a[67]), .Z(n4547) );
  NAND U5980 ( .A(a[66]), .B(b[1]), .Z(n4546) );
  XNOR U5981 ( .A(n4547), .B(n4546), .Z(n4549) );
  XNOR U5982 ( .A(n4548), .B(n4549), .Z(n4553) );
  XOR U5983 ( .A(n4552), .B(sreg[1089]), .Z(n4545) );
  XNOR U5984 ( .A(n4553), .B(n4545), .Z(c[1089]) );
  NAND U5985 ( .A(n4547), .B(n4546), .Z(n4551) );
  NANDN U5986 ( .A(n4549), .B(n4548), .Z(n4550) );
  NAND U5987 ( .A(n4551), .B(n4550), .Z(n4558) );
  ANDN U5988 ( .B(a[68]), .A(n3920), .Z(n4556) );
  AND U5989 ( .A(b[1]), .B(a[67]), .Z(n4555) );
  XOR U5990 ( .A(n4556), .B(n4555), .Z(n4557) );
  XNOR U5991 ( .A(n4558), .B(n4557), .Z(n4560) );
  XOR U5992 ( .A(sreg[1090]), .B(n4559), .Z(n4554) );
  XNOR U5993 ( .A(n4560), .B(n4554), .Z(c[1090]) );
  NAND U5994 ( .A(b[0]), .B(a[69]), .Z(n4563) );
  NAND U5995 ( .A(a[68]), .B(b[1]), .Z(n4562) );
  XNOR U5996 ( .A(n4563), .B(n4562), .Z(n4565) );
  XNOR U5997 ( .A(n4564), .B(n4565), .Z(n4569) );
  XOR U5998 ( .A(n4568), .B(sreg[1091]), .Z(n4561) );
  XNOR U5999 ( .A(n4569), .B(n4561), .Z(c[1091]) );
  NAND U6000 ( .A(n4563), .B(n4562), .Z(n4567) );
  NANDN U6001 ( .A(n4565), .B(n4564), .Z(n4566) );
  NAND U6002 ( .A(n4567), .B(n4566), .Z(n4574) );
  ANDN U6003 ( .B(a[70]), .A(n3920), .Z(n4572) );
  AND U6004 ( .A(b[1]), .B(a[69]), .Z(n4571) );
  XOR U6005 ( .A(n4572), .B(n4571), .Z(n4573) );
  XNOR U6006 ( .A(n4574), .B(n4573), .Z(n4576) );
  XOR U6007 ( .A(sreg[1092]), .B(n4575), .Z(n4570) );
  XNOR U6008 ( .A(n4576), .B(n4570), .Z(c[1092]) );
  ANDN U6009 ( .B(a[71]), .A(n3920), .Z(n4579) );
  AND U6010 ( .A(b[1]), .B(a[70]), .Z(n4578) );
  XOR U6011 ( .A(n4579), .B(n4578), .Z(n4580) );
  XNOR U6012 ( .A(n4581), .B(n4580), .Z(n4583) );
  XNOR U6013 ( .A(sreg[1093]), .B(n4582), .Z(n4577) );
  XNOR U6014 ( .A(n4583), .B(n4577), .Z(c[1093]) );
  ANDN U6015 ( .B(a[72]), .A(n3920), .Z(n4586) );
  AND U6016 ( .A(b[1]), .B(a[71]), .Z(n4585) );
  XOR U6017 ( .A(n4586), .B(n4585), .Z(n4587) );
  XNOR U6018 ( .A(n4588), .B(n4587), .Z(n4590) );
  XNOR U6019 ( .A(sreg[1094]), .B(n4589), .Z(n4584) );
  XNOR U6020 ( .A(n4590), .B(n4584), .Z(c[1094]) );
  NAND U6021 ( .A(b[0]), .B(a[73]), .Z(n4593) );
  NAND U6022 ( .A(a[72]), .B(b[1]), .Z(n4592) );
  XNOR U6023 ( .A(n4593), .B(n4592), .Z(n4595) );
  XNOR U6024 ( .A(n4594), .B(n4595), .Z(n4599) );
  XOR U6025 ( .A(n4598), .B(sreg[1095]), .Z(n4591) );
  XNOR U6026 ( .A(n4599), .B(n4591), .Z(c[1095]) );
  NAND U6027 ( .A(n4593), .B(n4592), .Z(n4597) );
  NANDN U6028 ( .A(n4595), .B(n4594), .Z(n4596) );
  NAND U6029 ( .A(n4597), .B(n4596), .Z(n4604) );
  ANDN U6030 ( .B(a[74]), .A(n3921), .Z(n4602) );
  AND U6031 ( .A(b[1]), .B(a[73]), .Z(n4601) );
  XOR U6032 ( .A(n4602), .B(n4601), .Z(n4603) );
  XNOR U6033 ( .A(n4604), .B(n4603), .Z(n4609) );
  XOR U6034 ( .A(sreg[1096]), .B(n4608), .Z(n4600) );
  XNOR U6035 ( .A(n4609), .B(n4600), .Z(c[1096]) );
  OR U6036 ( .A(n4602), .B(n4601), .Z(n4607) );
  IV U6037 ( .A(n4603), .Z(n4605) );
  NANDN U6038 ( .A(n4605), .B(n4604), .Z(n4606) );
  NAND U6039 ( .A(n4607), .B(n4606), .Z(n4614) );
  ANDN U6040 ( .B(a[75]), .A(n3921), .Z(n4612) );
  AND U6041 ( .A(b[1]), .B(a[74]), .Z(n4611) );
  XOR U6042 ( .A(n4612), .B(n4611), .Z(n4613) );
  XNOR U6043 ( .A(n4614), .B(n4613), .Z(n4616) );
  XNOR U6044 ( .A(sreg[1097]), .B(n4615), .Z(n4610) );
  XNOR U6045 ( .A(n4616), .B(n4610), .Z(c[1097]) );
  ANDN U6046 ( .B(a[76]), .A(n3921), .Z(n4619) );
  AND U6047 ( .A(b[1]), .B(a[75]), .Z(n4618) );
  XOR U6048 ( .A(n4619), .B(n4618), .Z(n4620) );
  XNOR U6049 ( .A(n4621), .B(n4620), .Z(n4623) );
  XNOR U6050 ( .A(sreg[1098]), .B(n4622), .Z(n4617) );
  XNOR U6051 ( .A(n4623), .B(n4617), .Z(c[1098]) );
  ANDN U6052 ( .B(a[77]), .A(n3921), .Z(n4626) );
  AND U6053 ( .A(b[1]), .B(a[76]), .Z(n4625) );
  XOR U6054 ( .A(n4626), .B(n4625), .Z(n4627) );
  XNOR U6055 ( .A(n4628), .B(n4627), .Z(n4630) );
  XNOR U6056 ( .A(sreg[1099]), .B(n4629), .Z(n4624) );
  XNOR U6057 ( .A(n4630), .B(n4624), .Z(c[1099]) );
  ANDN U6058 ( .B(a[78]), .A(n3921), .Z(n4633) );
  AND U6059 ( .A(b[1]), .B(a[77]), .Z(n4632) );
  XOR U6060 ( .A(n4633), .B(n4632), .Z(n4634) );
  XNOR U6061 ( .A(n4635), .B(n4634), .Z(n4637) );
  XNOR U6062 ( .A(sreg[1100]), .B(n4636), .Z(n4631) );
  XNOR U6063 ( .A(n4637), .B(n4631), .Z(c[1100]) );
  NAND U6064 ( .A(b[0]), .B(a[79]), .Z(n4640) );
  NAND U6065 ( .A(a[78]), .B(b[1]), .Z(n4639) );
  XNOR U6066 ( .A(n4640), .B(n4639), .Z(n4642) );
  XNOR U6067 ( .A(n4641), .B(n4642), .Z(n4646) );
  XOR U6068 ( .A(n4645), .B(sreg[1101]), .Z(n4638) );
  XNOR U6069 ( .A(n4646), .B(n4638), .Z(c[1101]) );
  NAND U6070 ( .A(n4640), .B(n4639), .Z(n4644) );
  NANDN U6071 ( .A(n4642), .B(n4641), .Z(n4643) );
  NAND U6072 ( .A(n4644), .B(n4643), .Z(n4651) );
  ANDN U6073 ( .B(a[80]), .A(n3921), .Z(n4649) );
  AND U6074 ( .A(b[1]), .B(a[79]), .Z(n4648) );
  XOR U6075 ( .A(n4649), .B(n4648), .Z(n4650) );
  XNOR U6076 ( .A(n4651), .B(n4650), .Z(n4653) );
  XOR U6077 ( .A(sreg[1102]), .B(n4652), .Z(n4647) );
  XNOR U6078 ( .A(n4653), .B(n4647), .Z(c[1102]) );
  NAND U6079 ( .A(b[0]), .B(a[81]), .Z(n4656) );
  NAND U6080 ( .A(a[80]), .B(b[1]), .Z(n4655) );
  XNOR U6081 ( .A(n4656), .B(n4655), .Z(n4658) );
  XNOR U6082 ( .A(n4657), .B(n4658), .Z(n4662) );
  XOR U6083 ( .A(n4661), .B(sreg[1103]), .Z(n4654) );
  XNOR U6084 ( .A(n4662), .B(n4654), .Z(c[1103]) );
  NAND U6085 ( .A(n4656), .B(n4655), .Z(n4660) );
  NANDN U6086 ( .A(n4658), .B(n4657), .Z(n4659) );
  NAND U6087 ( .A(n4660), .B(n4659), .Z(n4667) );
  ANDN U6088 ( .B(a[82]), .A(n3921), .Z(n4665) );
  AND U6089 ( .A(b[1]), .B(a[81]), .Z(n4664) );
  XOR U6090 ( .A(n4665), .B(n4664), .Z(n4666) );
  XNOR U6091 ( .A(n4667), .B(n4666), .Z(n4669) );
  XOR U6092 ( .A(sreg[1104]), .B(n4668), .Z(n4663) );
  XNOR U6093 ( .A(n4669), .B(n4663), .Z(c[1104]) );
  NAND U6094 ( .A(b[0]), .B(a[83]), .Z(n4672) );
  NAND U6095 ( .A(a[82]), .B(b[1]), .Z(n4671) );
  XNOR U6096 ( .A(n4672), .B(n4671), .Z(n4674) );
  XNOR U6097 ( .A(n4673), .B(n4674), .Z(n4678) );
  XOR U6098 ( .A(n4677), .B(sreg[1105]), .Z(n4670) );
  XNOR U6099 ( .A(n4678), .B(n4670), .Z(c[1105]) );
  NAND U6100 ( .A(n4672), .B(n4671), .Z(n4676) );
  NANDN U6101 ( .A(n4674), .B(n4673), .Z(n4675) );
  NAND U6102 ( .A(n4676), .B(n4675), .Z(n4683) );
  ANDN U6103 ( .B(a[84]), .A(n3922), .Z(n4681) );
  AND U6104 ( .A(b[1]), .B(a[83]), .Z(n4680) );
  XOR U6105 ( .A(n4681), .B(n4680), .Z(n4682) );
  XNOR U6106 ( .A(n4683), .B(n4682), .Z(n4688) );
  XOR U6107 ( .A(sreg[1106]), .B(n4687), .Z(n4679) );
  XNOR U6108 ( .A(n4688), .B(n4679), .Z(c[1106]) );
  OR U6109 ( .A(n4681), .B(n4680), .Z(n4686) );
  IV U6110 ( .A(n4682), .Z(n4684) );
  NANDN U6111 ( .A(n4684), .B(n4683), .Z(n4685) );
  NAND U6112 ( .A(n4686), .B(n4685), .Z(n4692) );
  NAND U6113 ( .A(b[0]), .B(a[85]), .Z(n4691) );
  NAND U6114 ( .A(a[84]), .B(b[1]), .Z(n4690) );
  XNOR U6115 ( .A(n4691), .B(n4690), .Z(n4693) );
  XNOR U6116 ( .A(n4692), .B(n4693), .Z(n4697) );
  XOR U6117 ( .A(n4696), .B(sreg[1107]), .Z(n4689) );
  XNOR U6118 ( .A(n4697), .B(n4689), .Z(c[1107]) );
  NAND U6119 ( .A(n4691), .B(n4690), .Z(n4695) );
  NANDN U6120 ( .A(n4693), .B(n4692), .Z(n4694) );
  NAND U6121 ( .A(n4695), .B(n4694), .Z(n4702) );
  ANDN U6122 ( .B(a[86]), .A(n3922), .Z(n4700) );
  AND U6123 ( .A(b[1]), .B(a[85]), .Z(n4699) );
  XOR U6124 ( .A(n4700), .B(n4699), .Z(n4701) );
  XNOR U6125 ( .A(n4702), .B(n4701), .Z(n4704) );
  XOR U6126 ( .A(sreg[1108]), .B(n4703), .Z(n4698) );
  XNOR U6127 ( .A(n4704), .B(n4698), .Z(c[1108]) );
  NAND U6128 ( .A(b[0]), .B(a[87]), .Z(n4707) );
  NAND U6129 ( .A(a[86]), .B(b[1]), .Z(n4706) );
  XNOR U6130 ( .A(n4707), .B(n4706), .Z(n4709) );
  XNOR U6131 ( .A(n4708), .B(n4709), .Z(n4713) );
  XOR U6132 ( .A(n4712), .B(sreg[1109]), .Z(n4705) );
  XNOR U6133 ( .A(n4713), .B(n4705), .Z(c[1109]) );
  NAND U6134 ( .A(n4707), .B(n4706), .Z(n4711) );
  NANDN U6135 ( .A(n4709), .B(n4708), .Z(n4710) );
  NAND U6136 ( .A(n4711), .B(n4710), .Z(n4718) );
  ANDN U6137 ( .B(a[88]), .A(n3922), .Z(n4716) );
  AND U6138 ( .A(b[1]), .B(a[87]), .Z(n4715) );
  XOR U6139 ( .A(n4716), .B(n4715), .Z(n4717) );
  XNOR U6140 ( .A(n4718), .B(n4717), .Z(n4720) );
  XOR U6141 ( .A(sreg[1110]), .B(n4719), .Z(n4714) );
  XNOR U6142 ( .A(n4720), .B(n4714), .Z(c[1110]) );
  NAND U6143 ( .A(b[0]), .B(a[89]), .Z(n4723) );
  NAND U6144 ( .A(a[88]), .B(b[1]), .Z(n4722) );
  XNOR U6145 ( .A(n4723), .B(n4722), .Z(n4725) );
  XNOR U6146 ( .A(n4724), .B(n4725), .Z(n4729) );
  XOR U6147 ( .A(n4728), .B(sreg[1111]), .Z(n4721) );
  XNOR U6148 ( .A(n4729), .B(n4721), .Z(c[1111]) );
  NAND U6149 ( .A(n4723), .B(n4722), .Z(n4727) );
  NANDN U6150 ( .A(n4725), .B(n4724), .Z(n4726) );
  NAND U6151 ( .A(n4727), .B(n4726), .Z(n4734) );
  ANDN U6152 ( .B(a[90]), .A(n3922), .Z(n4732) );
  AND U6153 ( .A(b[1]), .B(a[89]), .Z(n4731) );
  XOR U6154 ( .A(n4732), .B(n4731), .Z(n4733) );
  XNOR U6155 ( .A(n4734), .B(n4733), .Z(n4736) );
  XOR U6156 ( .A(sreg[1112]), .B(n4735), .Z(n4730) );
  XNOR U6157 ( .A(n4736), .B(n4730), .Z(c[1112]) );
  NAND U6158 ( .A(b[0]), .B(a[91]), .Z(n4739) );
  NAND U6159 ( .A(a[90]), .B(b[1]), .Z(n4738) );
  XNOR U6160 ( .A(n4739), .B(n4738), .Z(n4741) );
  XNOR U6161 ( .A(n4740), .B(n4741), .Z(n4745) );
  XOR U6162 ( .A(n4744), .B(sreg[1113]), .Z(n4737) );
  XNOR U6163 ( .A(n4745), .B(n4737), .Z(c[1113]) );
  NAND U6164 ( .A(n4739), .B(n4738), .Z(n4743) );
  NANDN U6165 ( .A(n4741), .B(n4740), .Z(n4742) );
  NAND U6166 ( .A(n4743), .B(n4742), .Z(n4750) );
  ANDN U6167 ( .B(a[92]), .A(n3922), .Z(n4748) );
  AND U6168 ( .A(b[1]), .B(a[91]), .Z(n4747) );
  XOR U6169 ( .A(n4748), .B(n4747), .Z(n4749) );
  XNOR U6170 ( .A(n4750), .B(n4749), .Z(n4752) );
  XOR U6171 ( .A(sreg[1114]), .B(n4751), .Z(n4746) );
  XNOR U6172 ( .A(n4752), .B(n4746), .Z(c[1114]) );
  NAND U6173 ( .A(b[0]), .B(a[93]), .Z(n4755) );
  NAND U6174 ( .A(a[92]), .B(b[1]), .Z(n4754) );
  XNOR U6175 ( .A(n4755), .B(n4754), .Z(n4757) );
  XNOR U6176 ( .A(n4756), .B(n4757), .Z(n4761) );
  XOR U6177 ( .A(n4760), .B(sreg[1115]), .Z(n4753) );
  XNOR U6178 ( .A(n4761), .B(n4753), .Z(c[1115]) );
  NAND U6179 ( .A(n4755), .B(n4754), .Z(n4759) );
  NANDN U6180 ( .A(n4757), .B(n4756), .Z(n4758) );
  NAND U6181 ( .A(n4759), .B(n4758), .Z(n4766) );
  ANDN U6182 ( .B(a[94]), .A(n3922), .Z(n4764) );
  AND U6183 ( .A(b[1]), .B(a[93]), .Z(n4763) );
  XOR U6184 ( .A(n4764), .B(n4763), .Z(n4765) );
  XNOR U6185 ( .A(n4766), .B(n4765), .Z(n4768) );
  XOR U6186 ( .A(sreg[1116]), .B(n4767), .Z(n4762) );
  XNOR U6187 ( .A(n4768), .B(n4762), .Z(c[1116]) );
  NAND U6188 ( .A(b[0]), .B(a[95]), .Z(n4771) );
  NAND U6189 ( .A(a[94]), .B(b[1]), .Z(n4770) );
  XNOR U6190 ( .A(n4771), .B(n4770), .Z(n4773) );
  XNOR U6191 ( .A(n4772), .B(n4773), .Z(n4777) );
  XOR U6192 ( .A(n4776), .B(sreg[1117]), .Z(n4769) );
  XNOR U6193 ( .A(n4777), .B(n4769), .Z(c[1117]) );
  NAND U6194 ( .A(n4771), .B(n4770), .Z(n4775) );
  NANDN U6195 ( .A(n4773), .B(n4772), .Z(n4774) );
  NAND U6196 ( .A(n4775), .B(n4774), .Z(n4782) );
  ANDN U6197 ( .B(a[96]), .A(n3922), .Z(n4780) );
  AND U6198 ( .A(b[1]), .B(a[95]), .Z(n4779) );
  XOR U6199 ( .A(n4780), .B(n4779), .Z(n4781) );
  XNOR U6200 ( .A(n4782), .B(n4781), .Z(n4784) );
  XOR U6201 ( .A(sreg[1118]), .B(n4783), .Z(n4778) );
  XNOR U6202 ( .A(n4784), .B(n4778), .Z(c[1118]) );
  NAND U6203 ( .A(b[0]), .B(a[97]), .Z(n4787) );
  NAND U6204 ( .A(a[96]), .B(b[1]), .Z(n4786) );
  XNOR U6205 ( .A(n4787), .B(n4786), .Z(n4789) );
  XNOR U6206 ( .A(n4788), .B(n4789), .Z(n4793) );
  XOR U6207 ( .A(n4792), .B(sreg[1119]), .Z(n4785) );
  XNOR U6208 ( .A(n4793), .B(n4785), .Z(c[1119]) );
  NAND U6209 ( .A(n4787), .B(n4786), .Z(n4791) );
  NANDN U6210 ( .A(n4789), .B(n4788), .Z(n4790) );
  NAND U6211 ( .A(n4791), .B(n4790), .Z(n4798) );
  ANDN U6212 ( .B(a[98]), .A(n3923), .Z(n4796) );
  AND U6213 ( .A(b[1]), .B(a[97]), .Z(n4795) );
  XOR U6214 ( .A(n4796), .B(n4795), .Z(n4797) );
  XNOR U6215 ( .A(n4798), .B(n4797), .Z(n4803) );
  XOR U6216 ( .A(sreg[1120]), .B(n4802), .Z(n4794) );
  XNOR U6217 ( .A(n4803), .B(n4794), .Z(c[1120]) );
  OR U6218 ( .A(n4796), .B(n4795), .Z(n4801) );
  IV U6219 ( .A(n4797), .Z(n4799) );
  NANDN U6220 ( .A(n4799), .B(n4798), .Z(n4800) );
  NAND U6221 ( .A(n4801), .B(n4800), .Z(n4807) );
  NAND U6222 ( .A(b[0]), .B(a[99]), .Z(n4806) );
  NAND U6223 ( .A(a[98]), .B(b[1]), .Z(n4805) );
  XNOR U6224 ( .A(n4806), .B(n4805), .Z(n4808) );
  XNOR U6225 ( .A(n4807), .B(n4808), .Z(n4812) );
  XOR U6226 ( .A(n4811), .B(sreg[1121]), .Z(n4804) );
  XNOR U6227 ( .A(n4812), .B(n4804), .Z(c[1121]) );
  NAND U6228 ( .A(n4806), .B(n4805), .Z(n4810) );
  NANDN U6229 ( .A(n4808), .B(n4807), .Z(n4809) );
  NAND U6230 ( .A(n4810), .B(n4809), .Z(n4816) );
  NAND U6231 ( .A(b[0]), .B(a[100]), .Z(n4815) );
  NAND U6232 ( .A(a[99]), .B(b[1]), .Z(n4814) );
  XNOR U6233 ( .A(n4815), .B(n4814), .Z(n4817) );
  XNOR U6234 ( .A(n4816), .B(n4817), .Z(n4821) );
  XOR U6235 ( .A(n4820), .B(sreg[1122]), .Z(n4813) );
  XNOR U6236 ( .A(n4821), .B(n4813), .Z(c[1122]) );
  NAND U6237 ( .A(n4815), .B(n4814), .Z(n4819) );
  NANDN U6238 ( .A(n4817), .B(n4816), .Z(n4818) );
  NAND U6239 ( .A(n4819), .B(n4818), .Z(n4825) );
  NAND U6240 ( .A(b[0]), .B(a[101]), .Z(n4824) );
  NAND U6241 ( .A(a[100]), .B(b[1]), .Z(n4823) );
  XNOR U6242 ( .A(n4824), .B(n4823), .Z(n4826) );
  XNOR U6243 ( .A(n4825), .B(n4826), .Z(n4830) );
  XOR U6244 ( .A(n4829), .B(sreg[1123]), .Z(n4822) );
  XNOR U6245 ( .A(n4830), .B(n4822), .Z(c[1123]) );
  NAND U6246 ( .A(n4824), .B(n4823), .Z(n4828) );
  NANDN U6247 ( .A(n4826), .B(n4825), .Z(n4827) );
  NAND U6248 ( .A(n4828), .B(n4827), .Z(n4835) );
  ANDN U6249 ( .B(a[102]), .A(n3923), .Z(n4833) );
  AND U6250 ( .A(b[1]), .B(a[101]), .Z(n4832) );
  XOR U6251 ( .A(n4833), .B(n4832), .Z(n4834) );
  XNOR U6252 ( .A(n4835), .B(n4834), .Z(n4837) );
  XOR U6253 ( .A(sreg[1124]), .B(n4836), .Z(n4831) );
  XNOR U6254 ( .A(n4837), .B(n4831), .Z(c[1124]) );
  NAND U6255 ( .A(b[0]), .B(a[103]), .Z(n4840) );
  NAND U6256 ( .A(a[102]), .B(b[1]), .Z(n4839) );
  XNOR U6257 ( .A(n4840), .B(n4839), .Z(n4842) );
  XNOR U6258 ( .A(n4841), .B(n4842), .Z(n4846) );
  XOR U6259 ( .A(n4845), .B(sreg[1125]), .Z(n4838) );
  XNOR U6260 ( .A(n4846), .B(n4838), .Z(c[1125]) );
  NAND U6261 ( .A(n4840), .B(n4839), .Z(n4844) );
  NANDN U6262 ( .A(n4842), .B(n4841), .Z(n4843) );
  NAND U6263 ( .A(n4844), .B(n4843), .Z(n4851) );
  ANDN U6264 ( .B(a[104]), .A(n3923), .Z(n4849) );
  AND U6265 ( .A(b[1]), .B(a[103]), .Z(n4848) );
  XOR U6266 ( .A(n4849), .B(n4848), .Z(n4850) );
  XNOR U6267 ( .A(n4851), .B(n4850), .Z(n4853) );
  XOR U6268 ( .A(sreg[1126]), .B(n4852), .Z(n4847) );
  XNOR U6269 ( .A(n4853), .B(n4847), .Z(c[1126]) );
  NAND U6270 ( .A(b[0]), .B(a[105]), .Z(n4856) );
  NAND U6271 ( .A(a[104]), .B(b[1]), .Z(n4855) );
  XNOR U6272 ( .A(n4856), .B(n4855), .Z(n4858) );
  XNOR U6273 ( .A(n4857), .B(n4858), .Z(n4862) );
  XOR U6274 ( .A(n4861), .B(sreg[1127]), .Z(n4854) );
  XNOR U6275 ( .A(n4862), .B(n4854), .Z(c[1127]) );
  NAND U6276 ( .A(n4856), .B(n4855), .Z(n4860) );
  NANDN U6277 ( .A(n4858), .B(n4857), .Z(n4859) );
  NAND U6278 ( .A(n4860), .B(n4859), .Z(n4867) );
  ANDN U6279 ( .B(a[106]), .A(n3923), .Z(n4865) );
  AND U6280 ( .A(b[1]), .B(a[105]), .Z(n4864) );
  XOR U6281 ( .A(n4865), .B(n4864), .Z(n4866) );
  XNOR U6282 ( .A(n4867), .B(n4866), .Z(n4869) );
  XOR U6283 ( .A(sreg[1128]), .B(n4868), .Z(n4863) );
  XNOR U6284 ( .A(n4869), .B(n4863), .Z(c[1128]) );
  NAND U6285 ( .A(b[0]), .B(a[107]), .Z(n4872) );
  NAND U6286 ( .A(a[106]), .B(b[1]), .Z(n4871) );
  XNOR U6287 ( .A(n4872), .B(n4871), .Z(n4874) );
  XNOR U6288 ( .A(n4873), .B(n4874), .Z(n4878) );
  XOR U6289 ( .A(n4877), .B(sreg[1129]), .Z(n4870) );
  XNOR U6290 ( .A(n4878), .B(n4870), .Z(c[1129]) );
  NAND U6291 ( .A(n4872), .B(n4871), .Z(n4876) );
  NANDN U6292 ( .A(n4874), .B(n4873), .Z(n4875) );
  NAND U6293 ( .A(n4876), .B(n4875), .Z(n4882) );
  NAND U6294 ( .A(b[0]), .B(a[108]), .Z(n4881) );
  NAND U6295 ( .A(a[107]), .B(b[1]), .Z(n4880) );
  XNOR U6296 ( .A(n4881), .B(n4880), .Z(n4883) );
  XNOR U6297 ( .A(n4882), .B(n4883), .Z(n4887) );
  XOR U6298 ( .A(n4886), .B(sreg[1130]), .Z(n4879) );
  XNOR U6299 ( .A(n4887), .B(n4879), .Z(c[1130]) );
  NAND U6300 ( .A(n4881), .B(n4880), .Z(n4885) );
  NANDN U6301 ( .A(n4883), .B(n4882), .Z(n4884) );
  NAND U6302 ( .A(n4885), .B(n4884), .Z(n4892) );
  ANDN U6303 ( .B(a[109]), .A(n3923), .Z(n4890) );
  AND U6304 ( .A(b[1]), .B(a[108]), .Z(n4889) );
  XOR U6305 ( .A(n4890), .B(n4889), .Z(n4891) );
  XNOR U6306 ( .A(n4892), .B(n4891), .Z(n4894) );
  XOR U6307 ( .A(sreg[1131]), .B(n4893), .Z(n4888) );
  XNOR U6308 ( .A(n4894), .B(n4888), .Z(c[1131]) );
  ANDN U6309 ( .B(a[110]), .A(n3923), .Z(n4897) );
  AND U6310 ( .A(b[1]), .B(a[109]), .Z(n4896) );
  XOR U6311 ( .A(n4897), .B(n4896), .Z(n4898) );
  XNOR U6312 ( .A(n4899), .B(n4898), .Z(n4901) );
  XNOR U6313 ( .A(sreg[1132]), .B(n4900), .Z(n4895) );
  XNOR U6314 ( .A(n4901), .B(n4895), .Z(c[1132]) );
  ANDN U6315 ( .B(a[111]), .A(n3923), .Z(n4904) );
  AND U6316 ( .A(b[1]), .B(a[110]), .Z(n4903) );
  XOR U6317 ( .A(n4904), .B(n4903), .Z(n4905) );
  XNOR U6318 ( .A(n4906), .B(n4905), .Z(n4908) );
  XNOR U6319 ( .A(sreg[1133]), .B(n4907), .Z(n4902) );
  XNOR U6320 ( .A(n4908), .B(n4902), .Z(c[1133]) );
  ANDN U6321 ( .B(a[112]), .A(n3924), .Z(n4911) );
  AND U6322 ( .A(b[1]), .B(a[111]), .Z(n4910) );
  XOR U6323 ( .A(n4911), .B(n4910), .Z(n4912) );
  XNOR U6324 ( .A(n4913), .B(n4912), .Z(n4918) );
  XNOR U6325 ( .A(sreg[1134]), .B(n4917), .Z(n4909) );
  XNOR U6326 ( .A(n4918), .B(n4909), .Z(c[1134]) );
  OR U6327 ( .A(n4911), .B(n4910), .Z(n4916) );
  IV U6328 ( .A(n4912), .Z(n4914) );
  NANDN U6329 ( .A(n4914), .B(n4913), .Z(n4915) );
  NAND U6330 ( .A(n4916), .B(n4915), .Z(n4922) );
  NAND U6331 ( .A(b[0]), .B(a[113]), .Z(n4921) );
  NAND U6332 ( .A(a[112]), .B(b[1]), .Z(n4920) );
  XNOR U6333 ( .A(n4921), .B(n4920), .Z(n4923) );
  XNOR U6334 ( .A(n4922), .B(n4923), .Z(n4927) );
  XOR U6335 ( .A(n4926), .B(sreg[1135]), .Z(n4919) );
  XNOR U6336 ( .A(n4927), .B(n4919), .Z(c[1135]) );
  NAND U6337 ( .A(n4921), .B(n4920), .Z(n4925) );
  NANDN U6338 ( .A(n4923), .B(n4922), .Z(n4924) );
  NAND U6339 ( .A(n4925), .B(n4924), .Z(n4931) );
  NAND U6340 ( .A(b[0]), .B(a[114]), .Z(n4930) );
  NAND U6341 ( .A(a[113]), .B(b[1]), .Z(n4929) );
  XNOR U6342 ( .A(n4930), .B(n4929), .Z(n4932) );
  XNOR U6343 ( .A(n4931), .B(n4932), .Z(n4936) );
  XOR U6344 ( .A(n4935), .B(sreg[1136]), .Z(n4928) );
  XNOR U6345 ( .A(n4936), .B(n4928), .Z(c[1136]) );
  NAND U6346 ( .A(n4930), .B(n4929), .Z(n4934) );
  NANDN U6347 ( .A(n4932), .B(n4931), .Z(n4933) );
  NAND U6348 ( .A(n4934), .B(n4933), .Z(n4940) );
  NAND U6349 ( .A(b[0]), .B(a[115]), .Z(n4939) );
  NAND U6350 ( .A(a[114]), .B(b[1]), .Z(n4938) );
  XNOR U6351 ( .A(n4939), .B(n4938), .Z(n4941) );
  XNOR U6352 ( .A(n4940), .B(n4941), .Z(n4945) );
  XOR U6353 ( .A(n4944), .B(sreg[1137]), .Z(n4937) );
  XNOR U6354 ( .A(n4945), .B(n4937), .Z(c[1137]) );
  NAND U6355 ( .A(n4939), .B(n4938), .Z(n4943) );
  NANDN U6356 ( .A(n4941), .B(n4940), .Z(n4942) );
  NAND U6357 ( .A(n4943), .B(n4942), .Z(n4949) );
  NAND U6358 ( .A(b[0]), .B(a[116]), .Z(n4948) );
  NAND U6359 ( .A(a[115]), .B(b[1]), .Z(n4947) );
  XNOR U6360 ( .A(n4948), .B(n4947), .Z(n4950) );
  XNOR U6361 ( .A(n4949), .B(n4950), .Z(n4954) );
  XOR U6362 ( .A(n4953), .B(sreg[1138]), .Z(n4946) );
  XNOR U6363 ( .A(n4954), .B(n4946), .Z(c[1138]) );
  NAND U6364 ( .A(n4948), .B(n4947), .Z(n4952) );
  NANDN U6365 ( .A(n4950), .B(n4949), .Z(n4951) );
  NAND U6366 ( .A(n4952), .B(n4951), .Z(n4958) );
  NAND U6367 ( .A(b[0]), .B(a[117]), .Z(n4957) );
  NAND U6368 ( .A(a[116]), .B(b[1]), .Z(n4956) );
  XNOR U6369 ( .A(n4957), .B(n4956), .Z(n4959) );
  XNOR U6370 ( .A(n4958), .B(n4959), .Z(n4963) );
  XOR U6371 ( .A(n4962), .B(sreg[1139]), .Z(n4955) );
  XNOR U6372 ( .A(n4963), .B(n4955), .Z(c[1139]) );
  NAND U6373 ( .A(n4957), .B(n4956), .Z(n4961) );
  NANDN U6374 ( .A(n4959), .B(n4958), .Z(n4960) );
  NAND U6375 ( .A(n4961), .B(n4960), .Z(n4968) );
  ANDN U6376 ( .B(a[118]), .A(n3924), .Z(n4966) );
  AND U6377 ( .A(b[1]), .B(a[117]), .Z(n4965) );
  XOR U6378 ( .A(n4966), .B(n4965), .Z(n4967) );
  XNOR U6379 ( .A(n4968), .B(n4967), .Z(n4970) );
  XOR U6380 ( .A(sreg[1140]), .B(n4969), .Z(n4964) );
  XNOR U6381 ( .A(n4970), .B(n4964), .Z(c[1140]) );
  NAND U6382 ( .A(b[0]), .B(a[119]), .Z(n4973) );
  NAND U6383 ( .A(a[118]), .B(b[1]), .Z(n4972) );
  XNOR U6384 ( .A(n4973), .B(n4972), .Z(n4975) );
  XNOR U6385 ( .A(n4974), .B(n4975), .Z(n4979) );
  XOR U6386 ( .A(n4978), .B(sreg[1141]), .Z(n4971) );
  XNOR U6387 ( .A(n4979), .B(n4971), .Z(c[1141]) );
  NAND U6388 ( .A(n4973), .B(n4972), .Z(n4977) );
  NANDN U6389 ( .A(n4975), .B(n4974), .Z(n4976) );
  NAND U6390 ( .A(n4977), .B(n4976), .Z(n4984) );
  ANDN U6391 ( .B(a[120]), .A(n3924), .Z(n4982) );
  AND U6392 ( .A(b[1]), .B(a[119]), .Z(n4981) );
  XOR U6393 ( .A(n4982), .B(n4981), .Z(n4983) );
  XNOR U6394 ( .A(n4984), .B(n4983), .Z(n4986) );
  XOR U6395 ( .A(sreg[1142]), .B(n4985), .Z(n4980) );
  XNOR U6396 ( .A(n4986), .B(n4980), .Z(c[1142]) );
  NAND U6397 ( .A(b[0]), .B(a[121]), .Z(n4989) );
  NAND U6398 ( .A(a[120]), .B(b[1]), .Z(n4988) );
  XNOR U6399 ( .A(n4989), .B(n4988), .Z(n4991) );
  XNOR U6400 ( .A(n4990), .B(n4991), .Z(n4995) );
  XOR U6401 ( .A(n4994), .B(sreg[1143]), .Z(n4987) );
  XNOR U6402 ( .A(n4995), .B(n4987), .Z(c[1143]) );
  NAND U6403 ( .A(n4989), .B(n4988), .Z(n4993) );
  NANDN U6404 ( .A(n4991), .B(n4990), .Z(n4992) );
  NAND U6405 ( .A(n4993), .B(n4992), .Z(n5000) );
  ANDN U6406 ( .B(a[122]), .A(n3924), .Z(n4998) );
  AND U6407 ( .A(b[1]), .B(a[121]), .Z(n4997) );
  XOR U6408 ( .A(n4998), .B(n4997), .Z(n4999) );
  XNOR U6409 ( .A(n5000), .B(n4999), .Z(n5002) );
  XOR U6410 ( .A(sreg[1144]), .B(n5001), .Z(n4996) );
  XNOR U6411 ( .A(n5002), .B(n4996), .Z(c[1144]) );
  NAND U6412 ( .A(b[0]), .B(a[123]), .Z(n5005) );
  NAND U6413 ( .A(a[122]), .B(b[1]), .Z(n5004) );
  XNOR U6414 ( .A(n5005), .B(n5004), .Z(n5007) );
  XNOR U6415 ( .A(n5006), .B(n5007), .Z(n5011) );
  XOR U6416 ( .A(n5010), .B(sreg[1145]), .Z(n5003) );
  XNOR U6417 ( .A(n5011), .B(n5003), .Z(c[1145]) );
  NAND U6418 ( .A(n5005), .B(n5004), .Z(n5009) );
  NANDN U6419 ( .A(n5007), .B(n5006), .Z(n5008) );
  NAND U6420 ( .A(n5009), .B(n5008), .Z(n5015) );
  NAND U6421 ( .A(b[0]), .B(a[124]), .Z(n5014) );
  NAND U6422 ( .A(a[123]), .B(b[1]), .Z(n5013) );
  XNOR U6423 ( .A(n5014), .B(n5013), .Z(n5016) );
  XNOR U6424 ( .A(n5015), .B(n5016), .Z(n5020) );
  XOR U6425 ( .A(n5019), .B(sreg[1146]), .Z(n5012) );
  XNOR U6426 ( .A(n5020), .B(n5012), .Z(c[1146]) );
  NAND U6427 ( .A(n5014), .B(n5013), .Z(n5018) );
  NANDN U6428 ( .A(n5016), .B(n5015), .Z(n5017) );
  NAND U6429 ( .A(n5018), .B(n5017), .Z(n5024) );
  NAND U6430 ( .A(b[0]), .B(a[125]), .Z(n5023) );
  NAND U6431 ( .A(a[124]), .B(b[1]), .Z(n5022) );
  XNOR U6432 ( .A(n5023), .B(n5022), .Z(n5025) );
  XNOR U6433 ( .A(n5024), .B(n5025), .Z(n5029) );
  XOR U6434 ( .A(n5028), .B(sreg[1147]), .Z(n5021) );
  XNOR U6435 ( .A(n5029), .B(n5021), .Z(c[1147]) );
  NAND U6436 ( .A(n5023), .B(n5022), .Z(n5027) );
  NANDN U6437 ( .A(n5025), .B(n5024), .Z(n5026) );
  NAND U6438 ( .A(n5027), .B(n5026), .Z(n5034) );
  ANDN U6439 ( .B(a[126]), .A(n3924), .Z(n5032) );
  AND U6440 ( .A(b[1]), .B(a[125]), .Z(n5031) );
  XOR U6441 ( .A(n5032), .B(n5031), .Z(n5033) );
  XNOR U6442 ( .A(n5034), .B(n5033), .Z(n5036) );
  XOR U6443 ( .A(sreg[1148]), .B(n5035), .Z(n5030) );
  XNOR U6444 ( .A(n5036), .B(n5030), .Z(c[1148]) );
  NAND U6445 ( .A(b[0]), .B(a[127]), .Z(n5039) );
  NAND U6446 ( .A(a[126]), .B(b[1]), .Z(n5038) );
  XNOR U6447 ( .A(n5039), .B(n5038), .Z(n5041) );
  XNOR U6448 ( .A(n5040), .B(n5041), .Z(n5045) );
  XOR U6449 ( .A(n5044), .B(sreg[1149]), .Z(n5037) );
  XNOR U6450 ( .A(n5045), .B(n5037), .Z(c[1149]) );
  NAND U6451 ( .A(n5039), .B(n5038), .Z(n5043) );
  NANDN U6452 ( .A(n5041), .B(n5040), .Z(n5042) );
  NAND U6453 ( .A(n5043), .B(n5042), .Z(n5050) );
  ANDN U6454 ( .B(a[128]), .A(n3924), .Z(n5048) );
  AND U6455 ( .A(b[1]), .B(a[127]), .Z(n5047) );
  XOR U6456 ( .A(n5048), .B(n5047), .Z(n5049) );
  XNOR U6457 ( .A(n5050), .B(n5049), .Z(n5052) );
  XOR U6458 ( .A(sreg[1150]), .B(n5051), .Z(n5046) );
  XNOR U6459 ( .A(n5052), .B(n5046), .Z(c[1150]) );
  NAND U6460 ( .A(b[0]), .B(a[129]), .Z(n5055) );
  NAND U6461 ( .A(a[128]), .B(b[1]), .Z(n5054) );
  XNOR U6462 ( .A(n5055), .B(n5054), .Z(n5057) );
  XNOR U6463 ( .A(n5056), .B(n5057), .Z(n5061) );
  XOR U6464 ( .A(n5060), .B(sreg[1151]), .Z(n5053) );
  XNOR U6465 ( .A(n5061), .B(n5053), .Z(c[1151]) );
  NAND U6466 ( .A(n5055), .B(n5054), .Z(n5059) );
  NANDN U6467 ( .A(n5057), .B(n5056), .Z(n5058) );
  NAND U6468 ( .A(n5059), .B(n5058), .Z(n5066) );
  ANDN U6469 ( .B(a[130]), .A(n3924), .Z(n5064) );
  AND U6470 ( .A(b[1]), .B(a[129]), .Z(n5063) );
  XOR U6471 ( .A(n5064), .B(n5063), .Z(n5065) );
  XNOR U6472 ( .A(n5066), .B(n5065), .Z(n5068) );
  XOR U6473 ( .A(sreg[1152]), .B(n5067), .Z(n5062) );
  XNOR U6474 ( .A(n5068), .B(n5062), .Z(c[1152]) );
  NAND U6475 ( .A(b[0]), .B(a[131]), .Z(n5071) );
  NAND U6476 ( .A(a[130]), .B(b[1]), .Z(n5070) );
  XNOR U6477 ( .A(n5071), .B(n5070), .Z(n5073) );
  XNOR U6478 ( .A(n5072), .B(n5073), .Z(n5077) );
  XOR U6479 ( .A(n5076), .B(sreg[1153]), .Z(n5069) );
  XNOR U6480 ( .A(n5077), .B(n5069), .Z(c[1153]) );
  NAND U6481 ( .A(n5071), .B(n5070), .Z(n5075) );
  NANDN U6482 ( .A(n5073), .B(n5072), .Z(n5074) );
  NAND U6483 ( .A(n5075), .B(n5074), .Z(n5082) );
  ANDN U6484 ( .B(a[132]), .A(n3925), .Z(n5080) );
  AND U6485 ( .A(b[1]), .B(a[131]), .Z(n5079) );
  XOR U6486 ( .A(n5080), .B(n5079), .Z(n5081) );
  XNOR U6487 ( .A(n5082), .B(n5081), .Z(n5087) );
  XOR U6488 ( .A(sreg[1154]), .B(n5086), .Z(n5078) );
  XNOR U6489 ( .A(n5087), .B(n5078), .Z(c[1154]) );
  OR U6490 ( .A(n5080), .B(n5079), .Z(n5085) );
  IV U6491 ( .A(n5081), .Z(n5083) );
  NANDN U6492 ( .A(n5083), .B(n5082), .Z(n5084) );
  NAND U6493 ( .A(n5085), .B(n5084), .Z(n5091) );
  NAND U6494 ( .A(b[0]), .B(a[133]), .Z(n5090) );
  NAND U6495 ( .A(a[132]), .B(b[1]), .Z(n5089) );
  XNOR U6496 ( .A(n5090), .B(n5089), .Z(n5092) );
  XNOR U6497 ( .A(n5091), .B(n5092), .Z(n5096) );
  XOR U6498 ( .A(n5095), .B(sreg[1155]), .Z(n5088) );
  XNOR U6499 ( .A(n5096), .B(n5088), .Z(c[1155]) );
  NAND U6500 ( .A(n5090), .B(n5089), .Z(n5094) );
  NANDN U6501 ( .A(n5092), .B(n5091), .Z(n5093) );
  NAND U6502 ( .A(n5094), .B(n5093), .Z(n5100) );
  NAND U6503 ( .A(b[0]), .B(a[134]), .Z(n5099) );
  NAND U6504 ( .A(a[133]), .B(b[1]), .Z(n5098) );
  XNOR U6505 ( .A(n5099), .B(n5098), .Z(n5101) );
  XNOR U6506 ( .A(n5100), .B(n5101), .Z(n5105) );
  XOR U6507 ( .A(n5104), .B(sreg[1156]), .Z(n5097) );
  XNOR U6508 ( .A(n5105), .B(n5097), .Z(c[1156]) );
  NAND U6509 ( .A(n5099), .B(n5098), .Z(n5103) );
  NANDN U6510 ( .A(n5101), .B(n5100), .Z(n5102) );
  NAND U6511 ( .A(n5103), .B(n5102), .Z(n5109) );
  NAND U6512 ( .A(b[0]), .B(a[135]), .Z(n5108) );
  NAND U6513 ( .A(a[134]), .B(b[1]), .Z(n5107) );
  XNOR U6514 ( .A(n5108), .B(n5107), .Z(n5110) );
  XNOR U6515 ( .A(n5109), .B(n5110), .Z(n5114) );
  XOR U6516 ( .A(n5113), .B(sreg[1157]), .Z(n5106) );
  XNOR U6517 ( .A(n5114), .B(n5106), .Z(c[1157]) );
  NAND U6518 ( .A(n5108), .B(n5107), .Z(n5112) );
  NANDN U6519 ( .A(n5110), .B(n5109), .Z(n5111) );
  NAND U6520 ( .A(n5112), .B(n5111), .Z(n5118) );
  NAND U6521 ( .A(b[0]), .B(a[136]), .Z(n5117) );
  NAND U6522 ( .A(a[135]), .B(b[1]), .Z(n5116) );
  XNOR U6523 ( .A(n5117), .B(n5116), .Z(n5119) );
  XNOR U6524 ( .A(n5118), .B(n5119), .Z(n5123) );
  XOR U6525 ( .A(n5122), .B(sreg[1158]), .Z(n5115) );
  XNOR U6526 ( .A(n5123), .B(n5115), .Z(c[1158]) );
  NAND U6527 ( .A(n5117), .B(n5116), .Z(n5121) );
  NANDN U6528 ( .A(n5119), .B(n5118), .Z(n5120) );
  NAND U6529 ( .A(n5121), .B(n5120), .Z(n5127) );
  NAND U6530 ( .A(b[0]), .B(a[137]), .Z(n5126) );
  NAND U6531 ( .A(a[136]), .B(b[1]), .Z(n5125) );
  XNOR U6532 ( .A(n5126), .B(n5125), .Z(n5128) );
  XNOR U6533 ( .A(n5127), .B(n5128), .Z(n5132) );
  XOR U6534 ( .A(n5131), .B(sreg[1159]), .Z(n5124) );
  XNOR U6535 ( .A(n5132), .B(n5124), .Z(c[1159]) );
  NAND U6536 ( .A(n5126), .B(n5125), .Z(n5130) );
  NANDN U6537 ( .A(n5128), .B(n5127), .Z(n5129) );
  NAND U6538 ( .A(n5130), .B(n5129), .Z(n5137) );
  ANDN U6539 ( .B(a[138]), .A(n3925), .Z(n5135) );
  AND U6540 ( .A(b[1]), .B(a[137]), .Z(n5134) );
  XOR U6541 ( .A(n5135), .B(n5134), .Z(n5136) );
  XNOR U6542 ( .A(n5137), .B(n5136), .Z(n5139) );
  XOR U6543 ( .A(sreg[1160]), .B(n5138), .Z(n5133) );
  XNOR U6544 ( .A(n5139), .B(n5133), .Z(c[1160]) );
  NAND U6545 ( .A(b[0]), .B(a[139]), .Z(n5142) );
  NAND U6546 ( .A(a[138]), .B(b[1]), .Z(n5141) );
  XNOR U6547 ( .A(n5142), .B(n5141), .Z(n5144) );
  XNOR U6548 ( .A(n5143), .B(n5144), .Z(n5148) );
  XOR U6549 ( .A(n5147), .B(sreg[1161]), .Z(n5140) );
  XNOR U6550 ( .A(n5148), .B(n5140), .Z(c[1161]) );
  NAND U6551 ( .A(n5142), .B(n5141), .Z(n5146) );
  NANDN U6552 ( .A(n5144), .B(n5143), .Z(n5145) );
  NAND U6553 ( .A(n5146), .B(n5145), .Z(n5153) );
  ANDN U6554 ( .B(a[140]), .A(n3925), .Z(n5151) );
  AND U6555 ( .A(b[1]), .B(a[139]), .Z(n5150) );
  XOR U6556 ( .A(n5151), .B(n5150), .Z(n5152) );
  XNOR U6557 ( .A(n5153), .B(n5152), .Z(n5155) );
  XOR U6558 ( .A(sreg[1162]), .B(n5154), .Z(n5149) );
  XNOR U6559 ( .A(n5155), .B(n5149), .Z(c[1162]) );
  NAND U6560 ( .A(b[0]), .B(a[141]), .Z(n5158) );
  NAND U6561 ( .A(a[140]), .B(b[1]), .Z(n5157) );
  XNOR U6562 ( .A(n5158), .B(n5157), .Z(n5160) );
  XNOR U6563 ( .A(n5159), .B(n5160), .Z(n5164) );
  XOR U6564 ( .A(n5163), .B(sreg[1163]), .Z(n5156) );
  XNOR U6565 ( .A(n5164), .B(n5156), .Z(c[1163]) );
  NAND U6566 ( .A(n5158), .B(n5157), .Z(n5162) );
  NANDN U6567 ( .A(n5160), .B(n5159), .Z(n5161) );
  NAND U6568 ( .A(n5162), .B(n5161), .Z(n5168) );
  NAND U6569 ( .A(b[0]), .B(a[142]), .Z(n5167) );
  NAND U6570 ( .A(a[141]), .B(b[1]), .Z(n5166) );
  XNOR U6571 ( .A(n5167), .B(n5166), .Z(n5169) );
  XNOR U6572 ( .A(n5168), .B(n5169), .Z(n5173) );
  XOR U6573 ( .A(n5172), .B(sreg[1164]), .Z(n5165) );
  XNOR U6574 ( .A(n5173), .B(n5165), .Z(c[1164]) );
  NAND U6575 ( .A(n5167), .B(n5166), .Z(n5171) );
  NANDN U6576 ( .A(n5169), .B(n5168), .Z(n5170) );
  NAND U6577 ( .A(n5171), .B(n5170), .Z(n5177) );
  NAND U6578 ( .A(b[0]), .B(a[143]), .Z(n5176) );
  NAND U6579 ( .A(a[142]), .B(b[1]), .Z(n5175) );
  XNOR U6580 ( .A(n5176), .B(n5175), .Z(n5178) );
  XNOR U6581 ( .A(n5177), .B(n5178), .Z(n5182) );
  XOR U6582 ( .A(n5181), .B(sreg[1165]), .Z(n5174) );
  XNOR U6583 ( .A(n5182), .B(n5174), .Z(c[1165]) );
  NAND U6584 ( .A(n5176), .B(n5175), .Z(n5180) );
  NANDN U6585 ( .A(n5178), .B(n5177), .Z(n5179) );
  NAND U6586 ( .A(n5180), .B(n5179), .Z(n5187) );
  ANDN U6587 ( .B(a[144]), .A(n3925), .Z(n5185) );
  AND U6588 ( .A(b[1]), .B(a[143]), .Z(n5184) );
  XOR U6589 ( .A(n5185), .B(n5184), .Z(n5186) );
  XNOR U6590 ( .A(n5187), .B(n5186), .Z(n5189) );
  XOR U6591 ( .A(sreg[1166]), .B(n5188), .Z(n5183) );
  XNOR U6592 ( .A(n5189), .B(n5183), .Z(c[1166]) );
  NAND U6593 ( .A(b[0]), .B(a[145]), .Z(n5192) );
  NAND U6594 ( .A(a[144]), .B(b[1]), .Z(n5191) );
  XNOR U6595 ( .A(n5192), .B(n5191), .Z(n5194) );
  XNOR U6596 ( .A(n5193), .B(n5194), .Z(n5198) );
  XOR U6597 ( .A(n5197), .B(sreg[1167]), .Z(n5190) );
  XNOR U6598 ( .A(n5198), .B(n5190), .Z(c[1167]) );
  NAND U6599 ( .A(n5192), .B(n5191), .Z(n5196) );
  NANDN U6600 ( .A(n5194), .B(n5193), .Z(n5195) );
  NAND U6601 ( .A(n5196), .B(n5195), .Z(n5203) );
  ANDN U6602 ( .B(a[146]), .A(n3925), .Z(n5201) );
  AND U6603 ( .A(b[1]), .B(a[145]), .Z(n5200) );
  XOR U6604 ( .A(n5201), .B(n5200), .Z(n5202) );
  XNOR U6605 ( .A(n5203), .B(n5202), .Z(n5205) );
  XOR U6606 ( .A(sreg[1168]), .B(n5204), .Z(n5199) );
  XNOR U6607 ( .A(n5205), .B(n5199), .Z(c[1168]) );
  NAND U6608 ( .A(b[0]), .B(a[147]), .Z(n5208) );
  NAND U6609 ( .A(a[146]), .B(b[1]), .Z(n5207) );
  XNOR U6610 ( .A(n5208), .B(n5207), .Z(n5210) );
  XNOR U6611 ( .A(n5209), .B(n5210), .Z(n5214) );
  XOR U6612 ( .A(n5213), .B(sreg[1169]), .Z(n5206) );
  XNOR U6613 ( .A(n5214), .B(n5206), .Z(c[1169]) );
  NAND U6614 ( .A(n5208), .B(n5207), .Z(n5212) );
  NANDN U6615 ( .A(n5210), .B(n5209), .Z(n5211) );
  NAND U6616 ( .A(n5212), .B(n5211), .Z(n5219) );
  ANDN U6617 ( .B(a[148]), .A(n3925), .Z(n5217) );
  AND U6618 ( .A(b[1]), .B(a[147]), .Z(n5216) );
  XOR U6619 ( .A(n5217), .B(n5216), .Z(n5218) );
  XNOR U6620 ( .A(n5219), .B(n5218), .Z(n5221) );
  XOR U6621 ( .A(sreg[1170]), .B(n5220), .Z(n5215) );
  XNOR U6622 ( .A(n5221), .B(n5215), .Z(c[1170]) );
  ANDN U6623 ( .B(a[149]), .A(n3925), .Z(n5224) );
  AND U6624 ( .A(b[1]), .B(a[148]), .Z(n5223) );
  XOR U6625 ( .A(n5224), .B(n5223), .Z(n5225) );
  XNOR U6626 ( .A(n5226), .B(n5225), .Z(n5228) );
  XNOR U6627 ( .A(sreg[1171]), .B(n5227), .Z(n5222) );
  XNOR U6628 ( .A(n5228), .B(n5222), .Z(c[1171]) );
  ANDN U6629 ( .B(a[150]), .A(n3926), .Z(n5231) );
  AND U6630 ( .A(b[1]), .B(a[149]), .Z(n5230) );
  XOR U6631 ( .A(n5231), .B(n5230), .Z(n5232) );
  XNOR U6632 ( .A(n5233), .B(n5232), .Z(n5238) );
  XNOR U6633 ( .A(sreg[1172]), .B(n5237), .Z(n5229) );
  XNOR U6634 ( .A(n5238), .B(n5229), .Z(c[1172]) );
  OR U6635 ( .A(n5231), .B(n5230), .Z(n5236) );
  IV U6636 ( .A(n5232), .Z(n5234) );
  NANDN U6637 ( .A(n5234), .B(n5233), .Z(n5235) );
  NAND U6638 ( .A(n5236), .B(n5235), .Z(n5242) );
  NAND U6639 ( .A(b[0]), .B(a[151]), .Z(n5241) );
  NAND U6640 ( .A(a[150]), .B(b[1]), .Z(n5240) );
  XNOR U6641 ( .A(n5241), .B(n5240), .Z(n5243) );
  XNOR U6642 ( .A(n5242), .B(n5243), .Z(n5247) );
  XOR U6643 ( .A(n5246), .B(sreg[1173]), .Z(n5239) );
  XNOR U6644 ( .A(n5247), .B(n5239), .Z(c[1173]) );
  NAND U6645 ( .A(n5241), .B(n5240), .Z(n5245) );
  NANDN U6646 ( .A(n5243), .B(n5242), .Z(n5244) );
  NAND U6647 ( .A(n5245), .B(n5244), .Z(n5252) );
  ANDN U6648 ( .B(a[152]), .A(n3926), .Z(n5250) );
  AND U6649 ( .A(b[1]), .B(a[151]), .Z(n5249) );
  XOR U6650 ( .A(n5250), .B(n5249), .Z(n5251) );
  XNOR U6651 ( .A(n5252), .B(n5251), .Z(n5254) );
  XOR U6652 ( .A(sreg[1174]), .B(n5253), .Z(n5248) );
  XNOR U6653 ( .A(n5254), .B(n5248), .Z(c[1174]) );
  NAND U6654 ( .A(b[0]), .B(a[153]), .Z(n5257) );
  NAND U6655 ( .A(a[152]), .B(b[1]), .Z(n5256) );
  XNOR U6656 ( .A(n5257), .B(n5256), .Z(n5259) );
  XNOR U6657 ( .A(n5258), .B(n5259), .Z(n5263) );
  XOR U6658 ( .A(n5262), .B(sreg[1175]), .Z(n5255) );
  XNOR U6659 ( .A(n5263), .B(n5255), .Z(c[1175]) );
  NAND U6660 ( .A(n5257), .B(n5256), .Z(n5261) );
  NANDN U6661 ( .A(n5259), .B(n5258), .Z(n5260) );
  NAND U6662 ( .A(n5261), .B(n5260), .Z(n5268) );
  ANDN U6663 ( .B(a[154]), .A(n3926), .Z(n5266) );
  AND U6664 ( .A(b[1]), .B(a[153]), .Z(n5265) );
  XOR U6665 ( .A(n5266), .B(n5265), .Z(n5267) );
  XNOR U6666 ( .A(n5268), .B(n5267), .Z(n5270) );
  XOR U6667 ( .A(sreg[1176]), .B(n5269), .Z(n5264) );
  XNOR U6668 ( .A(n5270), .B(n5264), .Z(c[1176]) );
  NAND U6669 ( .A(b[0]), .B(a[155]), .Z(n5273) );
  NAND U6670 ( .A(a[154]), .B(b[1]), .Z(n5272) );
  XNOR U6671 ( .A(n5273), .B(n5272), .Z(n5275) );
  XNOR U6672 ( .A(n5274), .B(n5275), .Z(n5279) );
  XOR U6673 ( .A(n5278), .B(sreg[1177]), .Z(n5271) );
  XNOR U6674 ( .A(n5279), .B(n5271), .Z(c[1177]) );
  NAND U6675 ( .A(n5273), .B(n5272), .Z(n5277) );
  NANDN U6676 ( .A(n5275), .B(n5274), .Z(n5276) );
  NAND U6677 ( .A(n5277), .B(n5276), .Z(n5284) );
  ANDN U6678 ( .B(a[156]), .A(n3926), .Z(n5282) );
  AND U6679 ( .A(b[1]), .B(a[155]), .Z(n5281) );
  XOR U6680 ( .A(n5282), .B(n5281), .Z(n5283) );
  XNOR U6681 ( .A(n5284), .B(n5283), .Z(n5286) );
  XOR U6682 ( .A(sreg[1178]), .B(n5285), .Z(n5280) );
  XNOR U6683 ( .A(n5286), .B(n5280), .Z(c[1178]) );
  NAND U6684 ( .A(b[0]), .B(a[157]), .Z(n5289) );
  NAND U6685 ( .A(a[156]), .B(b[1]), .Z(n5288) );
  XNOR U6686 ( .A(n5289), .B(n5288), .Z(n5291) );
  XNOR U6687 ( .A(n5290), .B(n5291), .Z(n5295) );
  XOR U6688 ( .A(n5294), .B(sreg[1179]), .Z(n5287) );
  XNOR U6689 ( .A(n5295), .B(n5287), .Z(c[1179]) );
  NAND U6690 ( .A(n5289), .B(n5288), .Z(n5293) );
  NANDN U6691 ( .A(n5291), .B(n5290), .Z(n5292) );
  NAND U6692 ( .A(n5293), .B(n5292), .Z(n5300) );
  ANDN U6693 ( .B(a[158]), .A(n3926), .Z(n5298) );
  AND U6694 ( .A(b[1]), .B(a[157]), .Z(n5297) );
  XOR U6695 ( .A(n5298), .B(n5297), .Z(n5299) );
  XNOR U6696 ( .A(n5300), .B(n5299), .Z(n5302) );
  XOR U6697 ( .A(sreg[1180]), .B(n5301), .Z(n5296) );
  XNOR U6698 ( .A(n5302), .B(n5296), .Z(c[1180]) );
  NAND U6699 ( .A(b[0]), .B(a[159]), .Z(n5305) );
  NAND U6700 ( .A(a[158]), .B(b[1]), .Z(n5304) );
  XNOR U6701 ( .A(n5305), .B(n5304), .Z(n5307) );
  XNOR U6702 ( .A(n5306), .B(n5307), .Z(n5311) );
  XOR U6703 ( .A(n5310), .B(sreg[1181]), .Z(n5303) );
  XNOR U6704 ( .A(n5311), .B(n5303), .Z(c[1181]) );
  NAND U6705 ( .A(n5305), .B(n5304), .Z(n5309) );
  NANDN U6706 ( .A(n5307), .B(n5306), .Z(n5308) );
  NAND U6707 ( .A(n5309), .B(n5308), .Z(n5316) );
  ANDN U6708 ( .B(a[160]), .A(n3926), .Z(n5314) );
  AND U6709 ( .A(b[1]), .B(a[159]), .Z(n5313) );
  XOR U6710 ( .A(n5314), .B(n5313), .Z(n5315) );
  XNOR U6711 ( .A(n5316), .B(n5315), .Z(n5318) );
  XOR U6712 ( .A(sreg[1182]), .B(n5317), .Z(n5312) );
  XNOR U6713 ( .A(n5318), .B(n5312), .Z(c[1182]) );
  NAND U6714 ( .A(b[0]), .B(a[161]), .Z(n5321) );
  NAND U6715 ( .A(a[160]), .B(b[1]), .Z(n5320) );
  XNOR U6716 ( .A(n5321), .B(n5320), .Z(n5323) );
  XNOR U6717 ( .A(n5322), .B(n5323), .Z(n5327) );
  XOR U6718 ( .A(n5326), .B(sreg[1183]), .Z(n5319) );
  XNOR U6719 ( .A(n5327), .B(n5319), .Z(c[1183]) );
  NAND U6720 ( .A(n5321), .B(n5320), .Z(n5325) );
  NANDN U6721 ( .A(n5323), .B(n5322), .Z(n5324) );
  NAND U6722 ( .A(n5325), .B(n5324), .Z(n5332) );
  ANDN U6723 ( .B(a[162]), .A(n3926), .Z(n5330) );
  AND U6724 ( .A(b[1]), .B(a[161]), .Z(n5329) );
  XOR U6725 ( .A(n5330), .B(n5329), .Z(n5331) );
  XNOR U6726 ( .A(n5332), .B(n5331), .Z(n5334) );
  XOR U6727 ( .A(sreg[1184]), .B(n5333), .Z(n5328) );
  XNOR U6728 ( .A(n5334), .B(n5328), .Z(c[1184]) );
  NAND U6729 ( .A(b[0]), .B(a[163]), .Z(n5337) );
  NAND U6730 ( .A(a[162]), .B(b[1]), .Z(n5336) );
  XNOR U6731 ( .A(n5337), .B(n5336), .Z(n5339) );
  XNOR U6732 ( .A(n5338), .B(n5339), .Z(n5343) );
  XOR U6733 ( .A(n5342), .B(sreg[1185]), .Z(n5335) );
  XNOR U6734 ( .A(n5343), .B(n5335), .Z(c[1185]) );
  NAND U6735 ( .A(n5337), .B(n5336), .Z(n5341) );
  NANDN U6736 ( .A(n5339), .B(n5338), .Z(n5340) );
  NAND U6737 ( .A(n5341), .B(n5340), .Z(n5348) );
  ANDN U6738 ( .B(a[164]), .A(n3927), .Z(n5346) );
  AND U6739 ( .A(b[1]), .B(a[163]), .Z(n5345) );
  XOR U6740 ( .A(n5346), .B(n5345), .Z(n5347) );
  XNOR U6741 ( .A(n5348), .B(n5347), .Z(n5353) );
  XOR U6742 ( .A(sreg[1186]), .B(n5352), .Z(n5344) );
  XNOR U6743 ( .A(n5353), .B(n5344), .Z(c[1186]) );
  OR U6744 ( .A(n5346), .B(n5345), .Z(n5351) );
  IV U6745 ( .A(n5347), .Z(n5349) );
  NANDN U6746 ( .A(n5349), .B(n5348), .Z(n5350) );
  NAND U6747 ( .A(n5351), .B(n5350), .Z(n5357) );
  NAND U6748 ( .A(b[0]), .B(a[165]), .Z(n5356) );
  NAND U6749 ( .A(a[164]), .B(b[1]), .Z(n5355) );
  XNOR U6750 ( .A(n5356), .B(n5355), .Z(n5358) );
  XNOR U6751 ( .A(n5357), .B(n5358), .Z(n5362) );
  XOR U6752 ( .A(n5361), .B(sreg[1187]), .Z(n5354) );
  XNOR U6753 ( .A(n5362), .B(n5354), .Z(c[1187]) );
  NAND U6754 ( .A(n5356), .B(n5355), .Z(n5360) );
  NANDN U6755 ( .A(n5358), .B(n5357), .Z(n5359) );
  NAND U6756 ( .A(n5360), .B(n5359), .Z(n5367) );
  ANDN U6757 ( .B(a[166]), .A(n3927), .Z(n5365) );
  AND U6758 ( .A(b[1]), .B(a[165]), .Z(n5364) );
  XOR U6759 ( .A(n5365), .B(n5364), .Z(n5366) );
  XNOR U6760 ( .A(n5367), .B(n5366), .Z(n5369) );
  XOR U6761 ( .A(sreg[1188]), .B(n5368), .Z(n5363) );
  XNOR U6762 ( .A(n5369), .B(n5363), .Z(c[1188]) );
  NAND U6763 ( .A(b[0]), .B(a[167]), .Z(n5372) );
  NAND U6764 ( .A(a[166]), .B(b[1]), .Z(n5371) );
  XNOR U6765 ( .A(n5372), .B(n5371), .Z(n5374) );
  XNOR U6766 ( .A(n5373), .B(n5374), .Z(n5378) );
  XOR U6767 ( .A(n5377), .B(sreg[1189]), .Z(n5370) );
  XNOR U6768 ( .A(n5378), .B(n5370), .Z(c[1189]) );
  NAND U6769 ( .A(n5372), .B(n5371), .Z(n5376) );
  NANDN U6770 ( .A(n5374), .B(n5373), .Z(n5375) );
  NAND U6771 ( .A(n5376), .B(n5375), .Z(n5383) );
  ANDN U6772 ( .B(a[168]), .A(n3927), .Z(n5381) );
  AND U6773 ( .A(b[1]), .B(a[167]), .Z(n5380) );
  XOR U6774 ( .A(n5381), .B(n5380), .Z(n5382) );
  XNOR U6775 ( .A(n5383), .B(n5382), .Z(n5385) );
  XOR U6776 ( .A(sreg[1190]), .B(n5384), .Z(n5379) );
  XNOR U6777 ( .A(n5385), .B(n5379), .Z(c[1190]) );
  ANDN U6778 ( .B(a[169]), .A(n3927), .Z(n5388) );
  AND U6779 ( .A(b[1]), .B(a[168]), .Z(n5387) );
  XOR U6780 ( .A(n5388), .B(n5387), .Z(n5389) );
  XNOR U6781 ( .A(n5390), .B(n5389), .Z(n5392) );
  XNOR U6782 ( .A(sreg[1191]), .B(n5391), .Z(n5386) );
  XNOR U6783 ( .A(n5392), .B(n5386), .Z(c[1191]) );
  ANDN U6784 ( .B(a[170]), .A(n3927), .Z(n5395) );
  AND U6785 ( .A(b[1]), .B(a[169]), .Z(n5394) );
  XOR U6786 ( .A(n5395), .B(n5394), .Z(n5396) );
  XNOR U6787 ( .A(n5397), .B(n5396), .Z(n5399) );
  XNOR U6788 ( .A(sreg[1192]), .B(n5398), .Z(n5393) );
  XNOR U6789 ( .A(n5399), .B(n5393), .Z(c[1192]) );
  ANDN U6790 ( .B(a[171]), .A(n3927), .Z(n5402) );
  AND U6791 ( .A(b[1]), .B(a[170]), .Z(n5401) );
  XOR U6792 ( .A(n5402), .B(n5401), .Z(n5403) );
  XNOR U6793 ( .A(n5404), .B(n5403), .Z(n5406) );
  XNOR U6794 ( .A(sreg[1193]), .B(n5405), .Z(n5400) );
  XNOR U6795 ( .A(n5406), .B(n5400), .Z(c[1193]) );
  ANDN U6796 ( .B(a[172]), .A(n3927), .Z(n5409) );
  AND U6797 ( .A(b[1]), .B(a[171]), .Z(n5408) );
  XOR U6798 ( .A(n5409), .B(n5408), .Z(n5410) );
  XNOR U6799 ( .A(n5411), .B(n5410), .Z(n5413) );
  XNOR U6800 ( .A(sreg[1194]), .B(n5412), .Z(n5407) );
  XNOR U6801 ( .A(n5413), .B(n5407), .Z(c[1194]) );
  NAND U6802 ( .A(b[0]), .B(a[173]), .Z(n5416) );
  NAND U6803 ( .A(a[172]), .B(b[1]), .Z(n5415) );
  XNOR U6804 ( .A(n5416), .B(n5415), .Z(n5418) );
  XNOR U6805 ( .A(n5417), .B(n5418), .Z(n5422) );
  XOR U6806 ( .A(n5421), .B(sreg[1195]), .Z(n5414) );
  XNOR U6807 ( .A(n5422), .B(n5414), .Z(c[1195]) );
  NAND U6808 ( .A(n5416), .B(n5415), .Z(n5420) );
  NANDN U6809 ( .A(n5418), .B(n5417), .Z(n5419) );
  NAND U6810 ( .A(n5420), .B(n5419), .Z(n5427) );
  ANDN U6811 ( .B(a[174]), .A(n3928), .Z(n5425) );
  AND U6812 ( .A(b[1]), .B(a[173]), .Z(n5424) );
  XOR U6813 ( .A(n5425), .B(n5424), .Z(n5426) );
  XNOR U6814 ( .A(n5427), .B(n5426), .Z(n5432) );
  XOR U6815 ( .A(sreg[1196]), .B(n5431), .Z(n5423) );
  XNOR U6816 ( .A(n5432), .B(n5423), .Z(c[1196]) );
  OR U6817 ( .A(n5425), .B(n5424), .Z(n5430) );
  IV U6818 ( .A(n5426), .Z(n5428) );
  NANDN U6819 ( .A(n5428), .B(n5427), .Z(n5429) );
  NAND U6820 ( .A(n5430), .B(n5429), .Z(n5436) );
  NAND U6821 ( .A(b[0]), .B(a[175]), .Z(n5435) );
  NAND U6822 ( .A(a[174]), .B(b[1]), .Z(n5434) );
  XNOR U6823 ( .A(n5435), .B(n5434), .Z(n5437) );
  XNOR U6824 ( .A(n5436), .B(n5437), .Z(n5441) );
  XOR U6825 ( .A(n5440), .B(sreg[1197]), .Z(n5433) );
  XNOR U6826 ( .A(n5441), .B(n5433), .Z(c[1197]) );
  NAND U6827 ( .A(n5435), .B(n5434), .Z(n5439) );
  NANDN U6828 ( .A(n5437), .B(n5436), .Z(n5438) );
  NAND U6829 ( .A(n5439), .B(n5438), .Z(n5445) );
  NAND U6830 ( .A(b[0]), .B(a[176]), .Z(n5444) );
  NAND U6831 ( .A(a[175]), .B(b[1]), .Z(n5443) );
  XNOR U6832 ( .A(n5444), .B(n5443), .Z(n5446) );
  XNOR U6833 ( .A(n5445), .B(n5446), .Z(n5450) );
  XOR U6834 ( .A(n5449), .B(sreg[1198]), .Z(n5442) );
  XNOR U6835 ( .A(n5450), .B(n5442), .Z(c[1198]) );
  NAND U6836 ( .A(n5444), .B(n5443), .Z(n5448) );
  NANDN U6837 ( .A(n5446), .B(n5445), .Z(n5447) );
  NAND U6838 ( .A(n5448), .B(n5447), .Z(n5454) );
  NAND U6839 ( .A(b[0]), .B(a[177]), .Z(n5453) );
  NAND U6840 ( .A(a[176]), .B(b[1]), .Z(n5452) );
  XNOR U6841 ( .A(n5453), .B(n5452), .Z(n5455) );
  XNOR U6842 ( .A(n5454), .B(n5455), .Z(n5459) );
  XOR U6843 ( .A(n5458), .B(sreg[1199]), .Z(n5451) );
  XNOR U6844 ( .A(n5459), .B(n5451), .Z(c[1199]) );
  NAND U6845 ( .A(n5453), .B(n5452), .Z(n5457) );
  NANDN U6846 ( .A(n5455), .B(n5454), .Z(n5456) );
  NAND U6847 ( .A(n5457), .B(n5456), .Z(n5464) );
  ANDN U6848 ( .B(a[178]), .A(n3928), .Z(n5462) );
  AND U6849 ( .A(b[1]), .B(a[177]), .Z(n5461) );
  XOR U6850 ( .A(n5462), .B(n5461), .Z(n5463) );
  XNOR U6851 ( .A(n5464), .B(n5463), .Z(n5466) );
  XOR U6852 ( .A(sreg[1200]), .B(n5465), .Z(n5460) );
  XNOR U6853 ( .A(n5466), .B(n5460), .Z(c[1200]) );
  NAND U6854 ( .A(b[0]), .B(a[179]), .Z(n5469) );
  NAND U6855 ( .A(a[178]), .B(b[1]), .Z(n5468) );
  XNOR U6856 ( .A(n5469), .B(n5468), .Z(n5471) );
  XNOR U6857 ( .A(n5470), .B(n5471), .Z(n5475) );
  XOR U6858 ( .A(n5474), .B(sreg[1201]), .Z(n5467) );
  XNOR U6859 ( .A(n5475), .B(n5467), .Z(c[1201]) );
  NAND U6860 ( .A(n5469), .B(n5468), .Z(n5473) );
  NANDN U6861 ( .A(n5471), .B(n5470), .Z(n5472) );
  NAND U6862 ( .A(n5473), .B(n5472), .Z(n5480) );
  ANDN U6863 ( .B(a[180]), .A(n3928), .Z(n5478) );
  AND U6864 ( .A(b[1]), .B(a[179]), .Z(n5477) );
  XOR U6865 ( .A(n5478), .B(n5477), .Z(n5479) );
  XNOR U6866 ( .A(n5480), .B(n5479), .Z(n5482) );
  XOR U6867 ( .A(sreg[1202]), .B(n5481), .Z(n5476) );
  XNOR U6868 ( .A(n5482), .B(n5476), .Z(c[1202]) );
  NAND U6869 ( .A(b[0]), .B(a[181]), .Z(n5485) );
  NAND U6870 ( .A(a[180]), .B(b[1]), .Z(n5484) );
  XNOR U6871 ( .A(n5485), .B(n5484), .Z(n5487) );
  XNOR U6872 ( .A(n5486), .B(n5487), .Z(n5491) );
  XOR U6873 ( .A(n5490), .B(sreg[1203]), .Z(n5483) );
  XNOR U6874 ( .A(n5491), .B(n5483), .Z(c[1203]) );
  NAND U6875 ( .A(n5485), .B(n5484), .Z(n5489) );
  NANDN U6876 ( .A(n5487), .B(n5486), .Z(n5488) );
  NAND U6877 ( .A(n5489), .B(n5488), .Z(n5496) );
  ANDN U6878 ( .B(a[182]), .A(n3928), .Z(n5494) );
  AND U6879 ( .A(b[1]), .B(a[181]), .Z(n5493) );
  XOR U6880 ( .A(n5494), .B(n5493), .Z(n5495) );
  XNOR U6881 ( .A(n5496), .B(n5495), .Z(n5498) );
  XOR U6882 ( .A(sreg[1204]), .B(n5497), .Z(n5492) );
  XNOR U6883 ( .A(n5498), .B(n5492), .Z(c[1204]) );
  NAND U6884 ( .A(b[0]), .B(a[183]), .Z(n5501) );
  NAND U6885 ( .A(a[182]), .B(b[1]), .Z(n5500) );
  XNOR U6886 ( .A(n5501), .B(n5500), .Z(n5503) );
  XNOR U6887 ( .A(n5502), .B(n5503), .Z(n5507) );
  XOR U6888 ( .A(n5506), .B(sreg[1205]), .Z(n5499) );
  XNOR U6889 ( .A(n5507), .B(n5499), .Z(c[1205]) );
  NAND U6890 ( .A(n5501), .B(n5500), .Z(n5505) );
  NANDN U6891 ( .A(n5503), .B(n5502), .Z(n5504) );
  NAND U6892 ( .A(n5505), .B(n5504), .Z(n5512) );
  ANDN U6893 ( .B(a[184]), .A(n3928), .Z(n5510) );
  AND U6894 ( .A(b[1]), .B(a[183]), .Z(n5509) );
  XOR U6895 ( .A(n5510), .B(n5509), .Z(n5511) );
  XNOR U6896 ( .A(n5512), .B(n5511), .Z(n5514) );
  XOR U6897 ( .A(sreg[1206]), .B(n5513), .Z(n5508) );
  XNOR U6898 ( .A(n5514), .B(n5508), .Z(c[1206]) );
  NAND U6899 ( .A(b[0]), .B(a[185]), .Z(n5517) );
  NAND U6900 ( .A(a[184]), .B(b[1]), .Z(n5516) );
  XNOR U6901 ( .A(n5517), .B(n5516), .Z(n5519) );
  XNOR U6902 ( .A(n5518), .B(n5519), .Z(n5523) );
  XOR U6903 ( .A(n5522), .B(sreg[1207]), .Z(n5515) );
  XNOR U6904 ( .A(n5523), .B(n5515), .Z(c[1207]) );
  NAND U6905 ( .A(n5517), .B(n5516), .Z(n5521) );
  NANDN U6906 ( .A(n5519), .B(n5518), .Z(n5520) );
  NAND U6907 ( .A(n5521), .B(n5520), .Z(n5528) );
  ANDN U6908 ( .B(a[186]), .A(n3928), .Z(n5526) );
  AND U6909 ( .A(b[1]), .B(a[185]), .Z(n5525) );
  XOR U6910 ( .A(n5526), .B(n5525), .Z(n5527) );
  XNOR U6911 ( .A(n5528), .B(n5527), .Z(n5530) );
  XOR U6912 ( .A(sreg[1208]), .B(n5529), .Z(n5524) );
  XNOR U6913 ( .A(n5530), .B(n5524), .Z(c[1208]) );
  NAND U6914 ( .A(b[0]), .B(a[187]), .Z(n5533) );
  NAND U6915 ( .A(a[186]), .B(b[1]), .Z(n5532) );
  XNOR U6916 ( .A(n5533), .B(n5532), .Z(n5535) );
  XNOR U6917 ( .A(n5534), .B(n5535), .Z(n5539) );
  XOR U6918 ( .A(n5538), .B(sreg[1209]), .Z(n5531) );
  XNOR U6919 ( .A(n5539), .B(n5531), .Z(c[1209]) );
  NAND U6920 ( .A(n5533), .B(n5532), .Z(n5537) );
  NANDN U6921 ( .A(n5535), .B(n5534), .Z(n5536) );
  NAND U6922 ( .A(n5537), .B(n5536), .Z(n5543) );
  NAND U6923 ( .A(b[0]), .B(a[188]), .Z(n5542) );
  NAND U6924 ( .A(a[187]), .B(b[1]), .Z(n5541) );
  XNOR U6925 ( .A(n5542), .B(n5541), .Z(n5544) );
  XNOR U6926 ( .A(n5543), .B(n5544), .Z(n5548) );
  XOR U6927 ( .A(n5547), .B(sreg[1210]), .Z(n5540) );
  XNOR U6928 ( .A(n5548), .B(n5540), .Z(c[1210]) );
  NAND U6929 ( .A(n5542), .B(n5541), .Z(n5546) );
  NANDN U6930 ( .A(n5544), .B(n5543), .Z(n5545) );
  NAND U6931 ( .A(n5546), .B(n5545), .Z(n5552) );
  NAND U6932 ( .A(b[0]), .B(a[189]), .Z(n5551) );
  NAND U6933 ( .A(a[188]), .B(b[1]), .Z(n5550) );
  XNOR U6934 ( .A(n5551), .B(n5550), .Z(n5553) );
  XNOR U6935 ( .A(n5552), .B(n5553), .Z(n5557) );
  XOR U6936 ( .A(n5556), .B(sreg[1211]), .Z(n5549) );
  XNOR U6937 ( .A(n5557), .B(n5549), .Z(c[1211]) );
  NAND U6938 ( .A(n5551), .B(n5550), .Z(n5555) );
  NANDN U6939 ( .A(n5553), .B(n5552), .Z(n5554) );
  NAND U6940 ( .A(n5555), .B(n5554), .Z(n5562) );
  ANDN U6941 ( .B(a[190]), .A(n3928), .Z(n5560) );
  AND U6942 ( .A(b[1]), .B(a[189]), .Z(n5559) );
  XOR U6943 ( .A(n5560), .B(n5559), .Z(n5561) );
  XNOR U6944 ( .A(n5562), .B(n5561), .Z(n5564) );
  XOR U6945 ( .A(sreg[1212]), .B(n5563), .Z(n5558) );
  XNOR U6946 ( .A(n5564), .B(n5558), .Z(c[1212]) );
  NAND U6947 ( .A(b[0]), .B(a[191]), .Z(n5567) );
  NAND U6948 ( .A(a[190]), .B(b[1]), .Z(n5566) );
  XNOR U6949 ( .A(n5567), .B(n5566), .Z(n5569) );
  XNOR U6950 ( .A(n5568), .B(n5569), .Z(n5573) );
  XOR U6951 ( .A(n5572), .B(sreg[1213]), .Z(n5565) );
  XNOR U6952 ( .A(n5573), .B(n5565), .Z(c[1213]) );
  NAND U6953 ( .A(n5567), .B(n5566), .Z(n5571) );
  NANDN U6954 ( .A(n5569), .B(n5568), .Z(n5570) );
  NAND U6955 ( .A(n5571), .B(n5570), .Z(n5578) );
  ANDN U6956 ( .B(a[192]), .A(n3929), .Z(n5576) );
  AND U6957 ( .A(b[1]), .B(a[191]), .Z(n5575) );
  XOR U6958 ( .A(n5576), .B(n5575), .Z(n5577) );
  XNOR U6959 ( .A(n5578), .B(n5577), .Z(n5583) );
  XOR U6960 ( .A(sreg[1214]), .B(n5582), .Z(n5574) );
  XNOR U6961 ( .A(n5583), .B(n5574), .Z(c[1214]) );
  OR U6962 ( .A(n5576), .B(n5575), .Z(n5581) );
  IV U6963 ( .A(n5577), .Z(n5579) );
  NANDN U6964 ( .A(n5579), .B(n5578), .Z(n5580) );
  NAND U6965 ( .A(n5581), .B(n5580), .Z(n5587) );
  NAND U6966 ( .A(b[0]), .B(a[193]), .Z(n5586) );
  NAND U6967 ( .A(a[192]), .B(b[1]), .Z(n5585) );
  XNOR U6968 ( .A(n5586), .B(n5585), .Z(n5588) );
  XNOR U6969 ( .A(n5587), .B(n5588), .Z(n5592) );
  XOR U6970 ( .A(n5591), .B(sreg[1215]), .Z(n5584) );
  XNOR U6971 ( .A(n5592), .B(n5584), .Z(c[1215]) );
  NAND U6972 ( .A(n5586), .B(n5585), .Z(n5590) );
  NANDN U6973 ( .A(n5588), .B(n5587), .Z(n5589) );
  NAND U6974 ( .A(n5590), .B(n5589), .Z(n5597) );
  ANDN U6975 ( .B(a[194]), .A(n3929), .Z(n5595) );
  AND U6976 ( .A(b[1]), .B(a[193]), .Z(n5594) );
  XOR U6977 ( .A(n5595), .B(n5594), .Z(n5596) );
  XNOR U6978 ( .A(n5597), .B(n5596), .Z(n5599) );
  XOR U6979 ( .A(sreg[1216]), .B(n5598), .Z(n5593) );
  XNOR U6980 ( .A(n5599), .B(n5593), .Z(c[1216]) );
  NAND U6981 ( .A(b[0]), .B(a[195]), .Z(n5602) );
  NAND U6982 ( .A(a[194]), .B(b[1]), .Z(n5601) );
  XNOR U6983 ( .A(n5602), .B(n5601), .Z(n5604) );
  XNOR U6984 ( .A(n5603), .B(n5604), .Z(n5608) );
  XOR U6985 ( .A(n5607), .B(sreg[1217]), .Z(n5600) );
  XNOR U6986 ( .A(n5608), .B(n5600), .Z(c[1217]) );
  NAND U6987 ( .A(n5602), .B(n5601), .Z(n5606) );
  NANDN U6988 ( .A(n5604), .B(n5603), .Z(n5605) );
  NAND U6989 ( .A(n5606), .B(n5605), .Z(n5613) );
  ANDN U6990 ( .B(a[196]), .A(n3929), .Z(n5611) );
  AND U6991 ( .A(b[1]), .B(a[195]), .Z(n5610) );
  XOR U6992 ( .A(n5611), .B(n5610), .Z(n5612) );
  XNOR U6993 ( .A(n5613), .B(n5612), .Z(n5615) );
  XOR U6994 ( .A(sreg[1218]), .B(n5614), .Z(n5609) );
  XNOR U6995 ( .A(n5615), .B(n5609), .Z(c[1218]) );
  NAND U6996 ( .A(b[0]), .B(a[197]), .Z(n5618) );
  NAND U6997 ( .A(a[196]), .B(b[1]), .Z(n5617) );
  XNOR U6998 ( .A(n5618), .B(n5617), .Z(n5620) );
  XNOR U6999 ( .A(n5619), .B(n5620), .Z(n5624) );
  XOR U7000 ( .A(n5623), .B(sreg[1219]), .Z(n5616) );
  XNOR U7001 ( .A(n5624), .B(n5616), .Z(c[1219]) );
  NAND U7002 ( .A(n5618), .B(n5617), .Z(n5622) );
  NANDN U7003 ( .A(n5620), .B(n5619), .Z(n5621) );
  NAND U7004 ( .A(n5622), .B(n5621), .Z(n5629) );
  ANDN U7005 ( .B(a[198]), .A(n3929), .Z(n5627) );
  AND U7006 ( .A(b[1]), .B(a[197]), .Z(n5626) );
  XOR U7007 ( .A(n5627), .B(n5626), .Z(n5628) );
  XNOR U7008 ( .A(n5629), .B(n5628), .Z(n5631) );
  XOR U7009 ( .A(sreg[1220]), .B(n5630), .Z(n5625) );
  XNOR U7010 ( .A(n5631), .B(n5625), .Z(c[1220]) );
  NAND U7011 ( .A(b[0]), .B(a[199]), .Z(n5634) );
  NAND U7012 ( .A(a[198]), .B(b[1]), .Z(n5633) );
  XNOR U7013 ( .A(n5634), .B(n5633), .Z(n5636) );
  XNOR U7014 ( .A(n5635), .B(n5636), .Z(n5640) );
  XOR U7015 ( .A(n5639), .B(sreg[1221]), .Z(n5632) );
  XNOR U7016 ( .A(n5640), .B(n5632), .Z(c[1221]) );
  NAND U7017 ( .A(n5634), .B(n5633), .Z(n5638) );
  NANDN U7018 ( .A(n5636), .B(n5635), .Z(n5637) );
  NAND U7019 ( .A(n5638), .B(n5637), .Z(n5645) );
  ANDN U7020 ( .B(a[200]), .A(n3929), .Z(n5643) );
  AND U7021 ( .A(b[1]), .B(a[199]), .Z(n5642) );
  XOR U7022 ( .A(n5643), .B(n5642), .Z(n5644) );
  XNOR U7023 ( .A(n5645), .B(n5644), .Z(n5647) );
  XOR U7024 ( .A(sreg[1222]), .B(n5646), .Z(n5641) );
  XNOR U7025 ( .A(n5647), .B(n5641), .Z(c[1222]) );
  ANDN U7026 ( .B(a[201]), .A(n3929), .Z(n5650) );
  AND U7027 ( .A(b[1]), .B(a[200]), .Z(n5649) );
  XOR U7028 ( .A(n5650), .B(n5649), .Z(n5651) );
  XNOR U7029 ( .A(n5652), .B(n5651), .Z(n5654) );
  XNOR U7030 ( .A(sreg[1223]), .B(n5653), .Z(n5648) );
  XNOR U7031 ( .A(n5654), .B(n5648), .Z(c[1223]) );
  ANDN U7032 ( .B(a[202]), .A(n3929), .Z(n5657) );
  AND U7033 ( .A(b[1]), .B(a[201]), .Z(n5656) );
  XOR U7034 ( .A(n5657), .B(n5656), .Z(n5658) );
  XNOR U7035 ( .A(n5659), .B(n5658), .Z(n5661) );
  XNOR U7036 ( .A(sreg[1224]), .B(n5660), .Z(n5655) );
  XNOR U7037 ( .A(n5661), .B(n5655), .Z(c[1224]) );
  NAND U7038 ( .A(b[0]), .B(a[203]), .Z(n5664) );
  NAND U7039 ( .A(a[202]), .B(b[1]), .Z(n5663) );
  XNOR U7040 ( .A(n5664), .B(n5663), .Z(n5666) );
  XNOR U7041 ( .A(n5665), .B(n5666), .Z(n5670) );
  XOR U7042 ( .A(n5669), .B(sreg[1225]), .Z(n5662) );
  XNOR U7043 ( .A(n5670), .B(n5662), .Z(c[1225]) );
  NAND U7044 ( .A(n5664), .B(n5663), .Z(n5668) );
  NANDN U7045 ( .A(n5666), .B(n5665), .Z(n5667) );
  NAND U7046 ( .A(n5668), .B(n5667), .Z(n5675) );
  ANDN U7047 ( .B(a[204]), .A(n3930), .Z(n5673) );
  AND U7048 ( .A(b[1]), .B(a[203]), .Z(n5672) );
  XOR U7049 ( .A(n5673), .B(n5672), .Z(n5674) );
  XNOR U7050 ( .A(n5675), .B(n5674), .Z(n5680) );
  XOR U7051 ( .A(sreg[1226]), .B(n5679), .Z(n5671) );
  XNOR U7052 ( .A(n5680), .B(n5671), .Z(c[1226]) );
  OR U7053 ( .A(n5673), .B(n5672), .Z(n5678) );
  IV U7054 ( .A(n5674), .Z(n5676) );
  NANDN U7055 ( .A(n5676), .B(n5675), .Z(n5677) );
  NAND U7056 ( .A(n5678), .B(n5677), .Z(n5684) );
  NAND U7057 ( .A(b[0]), .B(a[205]), .Z(n5683) );
  NAND U7058 ( .A(a[204]), .B(b[1]), .Z(n5682) );
  XNOR U7059 ( .A(n5683), .B(n5682), .Z(n5685) );
  XNOR U7060 ( .A(n5684), .B(n5685), .Z(n5689) );
  XOR U7061 ( .A(n5688), .B(sreg[1227]), .Z(n5681) );
  XNOR U7062 ( .A(n5689), .B(n5681), .Z(c[1227]) );
  NAND U7063 ( .A(n5683), .B(n5682), .Z(n5687) );
  NANDN U7064 ( .A(n5685), .B(n5684), .Z(n5686) );
  NAND U7065 ( .A(n5687), .B(n5686), .Z(n5694) );
  ANDN U7066 ( .B(a[206]), .A(n3930), .Z(n5692) );
  AND U7067 ( .A(b[1]), .B(a[205]), .Z(n5691) );
  XOR U7068 ( .A(n5692), .B(n5691), .Z(n5693) );
  XNOR U7069 ( .A(n5694), .B(n5693), .Z(n5696) );
  XOR U7070 ( .A(sreg[1228]), .B(n5695), .Z(n5690) );
  XNOR U7071 ( .A(n5696), .B(n5690), .Z(c[1228]) );
  NAND U7072 ( .A(b[0]), .B(a[207]), .Z(n5699) );
  NAND U7073 ( .A(a[206]), .B(b[1]), .Z(n5698) );
  XNOR U7074 ( .A(n5699), .B(n5698), .Z(n5701) );
  XNOR U7075 ( .A(n5700), .B(n5701), .Z(n5705) );
  XOR U7076 ( .A(n5704), .B(sreg[1229]), .Z(n5697) );
  XNOR U7077 ( .A(n5705), .B(n5697), .Z(c[1229]) );
  NAND U7078 ( .A(n5699), .B(n5698), .Z(n5703) );
  NANDN U7079 ( .A(n5701), .B(n5700), .Z(n5702) );
  NAND U7080 ( .A(n5703), .B(n5702), .Z(n5710) );
  ANDN U7081 ( .B(a[208]), .A(n3930), .Z(n5708) );
  AND U7082 ( .A(b[1]), .B(a[207]), .Z(n5707) );
  XOR U7083 ( .A(n5708), .B(n5707), .Z(n5709) );
  XNOR U7084 ( .A(n5710), .B(n5709), .Z(n5712) );
  XOR U7085 ( .A(sreg[1230]), .B(n5711), .Z(n5706) );
  XNOR U7086 ( .A(n5712), .B(n5706), .Z(c[1230]) );
  NAND U7087 ( .A(b[0]), .B(a[209]), .Z(n5715) );
  NAND U7088 ( .A(a[208]), .B(b[1]), .Z(n5714) );
  XNOR U7089 ( .A(n5715), .B(n5714), .Z(n5717) );
  XNOR U7090 ( .A(n5716), .B(n5717), .Z(n5721) );
  XOR U7091 ( .A(n5720), .B(sreg[1231]), .Z(n5713) );
  XNOR U7092 ( .A(n5721), .B(n5713), .Z(c[1231]) );
  NAND U7093 ( .A(n5715), .B(n5714), .Z(n5719) );
  NANDN U7094 ( .A(n5717), .B(n5716), .Z(n5718) );
  NAND U7095 ( .A(n5719), .B(n5718), .Z(n5726) );
  ANDN U7096 ( .B(a[210]), .A(n3930), .Z(n5724) );
  AND U7097 ( .A(b[1]), .B(a[209]), .Z(n5723) );
  XOR U7098 ( .A(n5724), .B(n5723), .Z(n5725) );
  XNOR U7099 ( .A(n5726), .B(n5725), .Z(n5728) );
  XOR U7100 ( .A(sreg[1232]), .B(n5727), .Z(n5722) );
  XNOR U7101 ( .A(n5728), .B(n5722), .Z(c[1232]) );
  NAND U7102 ( .A(b[0]), .B(a[211]), .Z(n5731) );
  NAND U7103 ( .A(a[210]), .B(b[1]), .Z(n5730) );
  XNOR U7104 ( .A(n5731), .B(n5730), .Z(n5733) );
  XNOR U7105 ( .A(n5732), .B(n5733), .Z(n5737) );
  XOR U7106 ( .A(n5736), .B(sreg[1233]), .Z(n5729) );
  XNOR U7107 ( .A(n5737), .B(n5729), .Z(c[1233]) );
  NAND U7108 ( .A(n5731), .B(n5730), .Z(n5735) );
  NANDN U7109 ( .A(n5733), .B(n5732), .Z(n5734) );
  NAND U7110 ( .A(n5735), .B(n5734), .Z(n5742) );
  ANDN U7111 ( .B(a[212]), .A(n3930), .Z(n5740) );
  AND U7112 ( .A(b[1]), .B(a[211]), .Z(n5739) );
  XOR U7113 ( .A(n5740), .B(n5739), .Z(n5741) );
  XNOR U7114 ( .A(n5742), .B(n5741), .Z(n5744) );
  XOR U7115 ( .A(sreg[1234]), .B(n5743), .Z(n5738) );
  XNOR U7116 ( .A(n5744), .B(n5738), .Z(c[1234]) );
  NAND U7117 ( .A(b[0]), .B(a[213]), .Z(n5747) );
  NAND U7118 ( .A(a[212]), .B(b[1]), .Z(n5746) );
  XNOR U7119 ( .A(n5747), .B(n5746), .Z(n5749) );
  XNOR U7120 ( .A(n5748), .B(n5749), .Z(n5753) );
  XOR U7121 ( .A(n5752), .B(sreg[1235]), .Z(n5745) );
  XNOR U7122 ( .A(n5753), .B(n5745), .Z(c[1235]) );
  NAND U7123 ( .A(n5747), .B(n5746), .Z(n5751) );
  NANDN U7124 ( .A(n5749), .B(n5748), .Z(n5750) );
  NAND U7125 ( .A(n5751), .B(n5750), .Z(n5757) );
  NAND U7126 ( .A(b[0]), .B(a[214]), .Z(n5756) );
  NAND U7127 ( .A(a[213]), .B(b[1]), .Z(n5755) );
  XNOR U7128 ( .A(n5756), .B(n5755), .Z(n5758) );
  XNOR U7129 ( .A(n5757), .B(n5758), .Z(n5762) );
  XOR U7130 ( .A(n5761), .B(sreg[1236]), .Z(n5754) );
  XNOR U7131 ( .A(n5762), .B(n5754), .Z(c[1236]) );
  NAND U7132 ( .A(n5756), .B(n5755), .Z(n5760) );
  NANDN U7133 ( .A(n5758), .B(n5757), .Z(n5759) );
  NAND U7134 ( .A(n5760), .B(n5759), .Z(n5766) );
  NAND U7135 ( .A(b[0]), .B(a[215]), .Z(n5765) );
  NAND U7136 ( .A(a[214]), .B(b[1]), .Z(n5764) );
  XNOR U7137 ( .A(n5765), .B(n5764), .Z(n5767) );
  XNOR U7138 ( .A(n5766), .B(n5767), .Z(n5771) );
  XOR U7139 ( .A(n5770), .B(sreg[1237]), .Z(n5763) );
  XNOR U7140 ( .A(n5771), .B(n5763), .Z(c[1237]) );
  NAND U7141 ( .A(n5765), .B(n5764), .Z(n5769) );
  NANDN U7142 ( .A(n5767), .B(n5766), .Z(n5768) );
  NAND U7143 ( .A(n5769), .B(n5768), .Z(n5776) );
  ANDN U7144 ( .B(a[216]), .A(n3930), .Z(n5774) );
  AND U7145 ( .A(b[1]), .B(a[215]), .Z(n5773) );
  XOR U7146 ( .A(n5774), .B(n5773), .Z(n5775) );
  XNOR U7147 ( .A(n5776), .B(n5775), .Z(n5778) );
  XOR U7148 ( .A(sreg[1238]), .B(n5777), .Z(n5772) );
  XNOR U7149 ( .A(n5778), .B(n5772), .Z(c[1238]) );
  NAND U7150 ( .A(b[0]), .B(a[217]), .Z(n5781) );
  NAND U7151 ( .A(a[216]), .B(b[1]), .Z(n5780) );
  XNOR U7152 ( .A(n5781), .B(n5780), .Z(n5783) );
  XNOR U7153 ( .A(n5782), .B(n5783), .Z(n5787) );
  XOR U7154 ( .A(n5786), .B(sreg[1239]), .Z(n5779) );
  XNOR U7155 ( .A(n5787), .B(n5779), .Z(c[1239]) );
  NAND U7156 ( .A(n5781), .B(n5780), .Z(n5785) );
  NANDN U7157 ( .A(n5783), .B(n5782), .Z(n5784) );
  NAND U7158 ( .A(n5785), .B(n5784), .Z(n5792) );
  ANDN U7159 ( .B(a[218]), .A(n3930), .Z(n5790) );
  AND U7160 ( .A(b[1]), .B(a[217]), .Z(n5789) );
  XOR U7161 ( .A(n5790), .B(n5789), .Z(n5791) );
  XNOR U7162 ( .A(n5792), .B(n5791), .Z(n5794) );
  XOR U7163 ( .A(sreg[1240]), .B(n5793), .Z(n5788) );
  XNOR U7164 ( .A(n5794), .B(n5788), .Z(c[1240]) );
  NAND U7165 ( .A(b[0]), .B(a[219]), .Z(n5797) );
  NAND U7166 ( .A(a[218]), .B(b[1]), .Z(n5796) );
  XNOR U7167 ( .A(n5797), .B(n5796), .Z(n5799) );
  XNOR U7168 ( .A(n5798), .B(n5799), .Z(n5803) );
  XOR U7169 ( .A(n5802), .B(sreg[1241]), .Z(n5795) );
  XNOR U7170 ( .A(n5803), .B(n5795), .Z(c[1241]) );
  NAND U7171 ( .A(n5797), .B(n5796), .Z(n5801) );
  NANDN U7172 ( .A(n5799), .B(n5798), .Z(n5800) );
  NAND U7173 ( .A(n5801), .B(n5800), .Z(n5807) );
  NAND U7174 ( .A(b[0]), .B(a[220]), .Z(n5806) );
  NAND U7175 ( .A(a[219]), .B(b[1]), .Z(n5805) );
  XNOR U7176 ( .A(n5806), .B(n5805), .Z(n5808) );
  XNOR U7177 ( .A(n5807), .B(n5808), .Z(n5812) );
  XOR U7178 ( .A(n5811), .B(sreg[1242]), .Z(n5804) );
  XNOR U7179 ( .A(n5812), .B(n5804), .Z(c[1242]) );
  NAND U7180 ( .A(n5806), .B(n5805), .Z(n5810) );
  NANDN U7181 ( .A(n5808), .B(n5807), .Z(n5809) );
  NAND U7182 ( .A(n5810), .B(n5809), .Z(n5816) );
  NAND U7183 ( .A(b[0]), .B(a[221]), .Z(n5815) );
  NAND U7184 ( .A(a[220]), .B(b[1]), .Z(n5814) );
  XNOR U7185 ( .A(n5815), .B(n5814), .Z(n5817) );
  XNOR U7186 ( .A(n5816), .B(n5817), .Z(n5821) );
  XOR U7187 ( .A(n5820), .B(sreg[1243]), .Z(n5813) );
  XNOR U7188 ( .A(n5821), .B(n5813), .Z(c[1243]) );
  NAND U7189 ( .A(n5815), .B(n5814), .Z(n5819) );
  NANDN U7190 ( .A(n5817), .B(n5816), .Z(n5818) );
  NAND U7191 ( .A(n5819), .B(n5818), .Z(n5826) );
  ANDN U7192 ( .B(a[222]), .A(n3931), .Z(n5824) );
  AND U7193 ( .A(b[1]), .B(a[221]), .Z(n5823) );
  XOR U7194 ( .A(n5824), .B(n5823), .Z(n5825) );
  XNOR U7195 ( .A(n5826), .B(n5825), .Z(n5831) );
  XOR U7196 ( .A(sreg[1244]), .B(n5830), .Z(n5822) );
  XNOR U7197 ( .A(n5831), .B(n5822), .Z(c[1244]) );
  OR U7198 ( .A(n5824), .B(n5823), .Z(n5829) );
  IV U7199 ( .A(n5825), .Z(n5827) );
  NANDN U7200 ( .A(n5827), .B(n5826), .Z(n5828) );
  NAND U7201 ( .A(n5829), .B(n5828), .Z(n5835) );
  NAND U7202 ( .A(b[0]), .B(a[223]), .Z(n5834) );
  NAND U7203 ( .A(a[222]), .B(b[1]), .Z(n5833) );
  XNOR U7204 ( .A(n5834), .B(n5833), .Z(n5836) );
  XNOR U7205 ( .A(n5835), .B(n5836), .Z(n5840) );
  XOR U7206 ( .A(n5839), .B(sreg[1245]), .Z(n5832) );
  XNOR U7207 ( .A(n5840), .B(n5832), .Z(c[1245]) );
  NAND U7208 ( .A(n5834), .B(n5833), .Z(n5838) );
  NANDN U7209 ( .A(n5836), .B(n5835), .Z(n5837) );
  NAND U7210 ( .A(n5838), .B(n5837), .Z(n5845) );
  ANDN U7211 ( .B(a[224]), .A(n3931), .Z(n5843) );
  AND U7212 ( .A(b[1]), .B(a[223]), .Z(n5842) );
  XOR U7213 ( .A(n5843), .B(n5842), .Z(n5844) );
  XNOR U7214 ( .A(n5845), .B(n5844), .Z(n5847) );
  XOR U7215 ( .A(sreg[1246]), .B(n5846), .Z(n5841) );
  XNOR U7216 ( .A(n5847), .B(n5841), .Z(c[1246]) );
  NAND U7217 ( .A(b[0]), .B(a[225]), .Z(n5850) );
  NAND U7218 ( .A(a[224]), .B(b[1]), .Z(n5849) );
  XNOR U7219 ( .A(n5850), .B(n5849), .Z(n5852) );
  XNOR U7220 ( .A(n5851), .B(n5852), .Z(n5856) );
  XOR U7221 ( .A(n5855), .B(sreg[1247]), .Z(n5848) );
  XNOR U7222 ( .A(n5856), .B(n5848), .Z(c[1247]) );
  NAND U7223 ( .A(n5850), .B(n5849), .Z(n5854) );
  NANDN U7224 ( .A(n5852), .B(n5851), .Z(n5853) );
  NAND U7225 ( .A(n5854), .B(n5853), .Z(n5861) );
  ANDN U7226 ( .B(a[226]), .A(n3931), .Z(n5859) );
  AND U7227 ( .A(b[1]), .B(a[225]), .Z(n5858) );
  XOR U7228 ( .A(n5859), .B(n5858), .Z(n5860) );
  XNOR U7229 ( .A(n5861), .B(n5860), .Z(n5863) );
  XOR U7230 ( .A(sreg[1248]), .B(n5862), .Z(n5857) );
  XNOR U7231 ( .A(n5863), .B(n5857), .Z(c[1248]) );
  NAND U7232 ( .A(b[0]), .B(a[227]), .Z(n5866) );
  NAND U7233 ( .A(a[226]), .B(b[1]), .Z(n5865) );
  XNOR U7234 ( .A(n5866), .B(n5865), .Z(n5868) );
  XNOR U7235 ( .A(n5867), .B(n5868), .Z(n5872) );
  XOR U7236 ( .A(n5871), .B(sreg[1249]), .Z(n5864) );
  XNOR U7237 ( .A(n5872), .B(n5864), .Z(c[1249]) );
  NAND U7238 ( .A(n5866), .B(n5865), .Z(n5870) );
  NANDN U7239 ( .A(n5868), .B(n5867), .Z(n5869) );
  NAND U7240 ( .A(n5870), .B(n5869), .Z(n5877) );
  ANDN U7241 ( .B(a[228]), .A(n3931), .Z(n5875) );
  AND U7242 ( .A(b[1]), .B(a[227]), .Z(n5874) );
  XOR U7243 ( .A(n5875), .B(n5874), .Z(n5876) );
  XNOR U7244 ( .A(n5877), .B(n5876), .Z(n5879) );
  XOR U7245 ( .A(sreg[1250]), .B(n5878), .Z(n5873) );
  XNOR U7246 ( .A(n5879), .B(n5873), .Z(c[1250]) );
  NAND U7247 ( .A(b[0]), .B(a[229]), .Z(n5882) );
  NAND U7248 ( .A(a[228]), .B(b[1]), .Z(n5881) );
  XNOR U7249 ( .A(n5882), .B(n5881), .Z(n5884) );
  XNOR U7250 ( .A(n5883), .B(n5884), .Z(n5888) );
  XOR U7251 ( .A(n5887), .B(sreg[1251]), .Z(n5880) );
  XNOR U7252 ( .A(n5888), .B(n5880), .Z(c[1251]) );
  NAND U7253 ( .A(n5882), .B(n5881), .Z(n5886) );
  NANDN U7254 ( .A(n5884), .B(n5883), .Z(n5885) );
  NAND U7255 ( .A(n5886), .B(n5885), .Z(n5893) );
  ANDN U7256 ( .B(a[230]), .A(n3931), .Z(n5891) );
  AND U7257 ( .A(b[1]), .B(a[229]), .Z(n5890) );
  XOR U7258 ( .A(n5891), .B(n5890), .Z(n5892) );
  XNOR U7259 ( .A(n5893), .B(n5892), .Z(n5895) );
  XOR U7260 ( .A(sreg[1252]), .B(n5894), .Z(n5889) );
  XNOR U7261 ( .A(n5895), .B(n5889), .Z(c[1252]) );
  NAND U7262 ( .A(b[0]), .B(a[231]), .Z(n5898) );
  NAND U7263 ( .A(a[230]), .B(b[1]), .Z(n5897) );
  XNOR U7264 ( .A(n5898), .B(n5897), .Z(n5900) );
  XNOR U7265 ( .A(n5899), .B(n5900), .Z(n5904) );
  XOR U7266 ( .A(n5903), .B(sreg[1253]), .Z(n5896) );
  XNOR U7267 ( .A(n5904), .B(n5896), .Z(c[1253]) );
  NAND U7268 ( .A(n5898), .B(n5897), .Z(n5902) );
  NANDN U7269 ( .A(n5900), .B(n5899), .Z(n5901) );
  NAND U7270 ( .A(n5902), .B(n5901), .Z(n5909) );
  ANDN U7271 ( .B(a[232]), .A(n3931), .Z(n5907) );
  AND U7272 ( .A(b[1]), .B(a[231]), .Z(n5906) );
  XOR U7273 ( .A(n5907), .B(n5906), .Z(n5908) );
  XNOR U7274 ( .A(n5909), .B(n5908), .Z(n5911) );
  XOR U7275 ( .A(sreg[1254]), .B(n5910), .Z(n5905) );
  XNOR U7276 ( .A(n5911), .B(n5905), .Z(c[1254]) );
  NAND U7277 ( .A(b[0]), .B(a[233]), .Z(n5914) );
  NAND U7278 ( .A(a[232]), .B(b[1]), .Z(n5913) );
  XNOR U7279 ( .A(n5914), .B(n5913), .Z(n5916) );
  XNOR U7280 ( .A(n5915), .B(n5916), .Z(n5920) );
  XOR U7281 ( .A(n5919), .B(sreg[1255]), .Z(n5912) );
  XNOR U7282 ( .A(n5920), .B(n5912), .Z(c[1255]) );
  NAND U7283 ( .A(n5914), .B(n5913), .Z(n5918) );
  NANDN U7284 ( .A(n5916), .B(n5915), .Z(n5917) );
  NAND U7285 ( .A(n5918), .B(n5917), .Z(n5924) );
  NAND U7286 ( .A(b[0]), .B(a[234]), .Z(n5923) );
  NAND U7287 ( .A(a[233]), .B(b[1]), .Z(n5922) );
  XNOR U7288 ( .A(n5923), .B(n5922), .Z(n5925) );
  XNOR U7289 ( .A(n5924), .B(n5925), .Z(n5929) );
  XOR U7290 ( .A(n5928), .B(sreg[1256]), .Z(n5921) );
  XNOR U7291 ( .A(n5929), .B(n5921), .Z(c[1256]) );
  NAND U7292 ( .A(n5923), .B(n5922), .Z(n5927) );
  NANDN U7293 ( .A(n5925), .B(n5924), .Z(n5926) );
  NAND U7294 ( .A(n5927), .B(n5926), .Z(n5933) );
  NAND U7295 ( .A(b[0]), .B(a[235]), .Z(n5932) );
  NAND U7296 ( .A(a[234]), .B(b[1]), .Z(n5931) );
  XNOR U7297 ( .A(n5932), .B(n5931), .Z(n5934) );
  XNOR U7298 ( .A(n5933), .B(n5934), .Z(n5938) );
  XOR U7299 ( .A(n5937), .B(sreg[1257]), .Z(n5930) );
  XNOR U7300 ( .A(n5938), .B(n5930), .Z(c[1257]) );
  NAND U7301 ( .A(n5932), .B(n5931), .Z(n5936) );
  NANDN U7302 ( .A(n5934), .B(n5933), .Z(n5935) );
  NAND U7303 ( .A(n5936), .B(n5935), .Z(n5943) );
  ANDN U7304 ( .B(a[236]), .A(n3931), .Z(n5941) );
  AND U7305 ( .A(b[1]), .B(a[235]), .Z(n5940) );
  XOR U7306 ( .A(n5941), .B(n5940), .Z(n5942) );
  XNOR U7307 ( .A(n5943), .B(n5942), .Z(n5945) );
  XOR U7308 ( .A(sreg[1258]), .B(n5944), .Z(n5939) );
  XNOR U7309 ( .A(n5945), .B(n5939), .Z(c[1258]) );
  NAND U7310 ( .A(b[0]), .B(a[237]), .Z(n5948) );
  NAND U7311 ( .A(a[236]), .B(b[1]), .Z(n5947) );
  XNOR U7312 ( .A(n5948), .B(n5947), .Z(n5950) );
  XNOR U7313 ( .A(n5949), .B(n5950), .Z(n5954) );
  XOR U7314 ( .A(n5953), .B(sreg[1259]), .Z(n5946) );
  XNOR U7315 ( .A(n5954), .B(n5946), .Z(c[1259]) );
  NAND U7316 ( .A(n5948), .B(n5947), .Z(n5952) );
  NANDN U7317 ( .A(n5950), .B(n5949), .Z(n5951) );
  NAND U7318 ( .A(n5952), .B(n5951), .Z(n5959) );
  ANDN U7319 ( .B(a[238]), .A(n3932), .Z(n5957) );
  AND U7320 ( .A(b[1]), .B(a[237]), .Z(n5956) );
  XOR U7321 ( .A(n5957), .B(n5956), .Z(n5958) );
  XNOR U7322 ( .A(n5959), .B(n5958), .Z(n5964) );
  XOR U7323 ( .A(sreg[1260]), .B(n5963), .Z(n5955) );
  XNOR U7324 ( .A(n5964), .B(n5955), .Z(c[1260]) );
  OR U7325 ( .A(n5957), .B(n5956), .Z(n5962) );
  IV U7326 ( .A(n5958), .Z(n5960) );
  NANDN U7327 ( .A(n5960), .B(n5959), .Z(n5961) );
  NAND U7328 ( .A(n5962), .B(n5961), .Z(n5969) );
  ANDN U7329 ( .B(a[239]), .A(n3932), .Z(n5967) );
  AND U7330 ( .A(b[1]), .B(a[238]), .Z(n5966) );
  XOR U7331 ( .A(n5967), .B(n5966), .Z(n5968) );
  XNOR U7332 ( .A(n5969), .B(n5968), .Z(n5971) );
  XNOR U7333 ( .A(sreg[1261]), .B(n5970), .Z(n5965) );
  XNOR U7334 ( .A(n5971), .B(n5965), .Z(c[1261]) );
  ANDN U7335 ( .B(a[240]), .A(n3932), .Z(n5974) );
  AND U7336 ( .A(b[1]), .B(a[239]), .Z(n5973) );
  XOR U7337 ( .A(n5974), .B(n5973), .Z(n5975) );
  XNOR U7338 ( .A(n5976), .B(n5975), .Z(n5978) );
  XNOR U7339 ( .A(sreg[1262]), .B(n5977), .Z(n5972) );
  XNOR U7340 ( .A(n5978), .B(n5972), .Z(c[1262]) );
  NAND U7341 ( .A(b[0]), .B(a[241]), .Z(n5981) );
  NAND U7342 ( .A(a[240]), .B(b[1]), .Z(n5980) );
  XNOR U7343 ( .A(n5981), .B(n5980), .Z(n5983) );
  XNOR U7344 ( .A(n5982), .B(n5983), .Z(n5987) );
  XOR U7345 ( .A(n5986), .B(sreg[1263]), .Z(n5979) );
  XNOR U7346 ( .A(n5987), .B(n5979), .Z(c[1263]) );
  NAND U7347 ( .A(n5981), .B(n5980), .Z(n5985) );
  NANDN U7348 ( .A(n5983), .B(n5982), .Z(n5984) );
  NAND U7349 ( .A(n5985), .B(n5984), .Z(n5992) );
  ANDN U7350 ( .B(a[242]), .A(n3932), .Z(n5990) );
  AND U7351 ( .A(b[1]), .B(a[241]), .Z(n5989) );
  XOR U7352 ( .A(n5990), .B(n5989), .Z(n5991) );
  XNOR U7353 ( .A(n5992), .B(n5991), .Z(n5994) );
  XOR U7354 ( .A(sreg[1264]), .B(n5993), .Z(n5988) );
  XNOR U7355 ( .A(n5994), .B(n5988), .Z(c[1264]) );
  NAND U7356 ( .A(b[0]), .B(a[243]), .Z(n5997) );
  NAND U7357 ( .A(a[242]), .B(b[1]), .Z(n5996) );
  XNOR U7358 ( .A(n5997), .B(n5996), .Z(n5999) );
  XNOR U7359 ( .A(n5998), .B(n5999), .Z(n6003) );
  XOR U7360 ( .A(n6002), .B(sreg[1265]), .Z(n5995) );
  XNOR U7361 ( .A(n6003), .B(n5995), .Z(c[1265]) );
  NAND U7362 ( .A(n5997), .B(n5996), .Z(n6001) );
  NANDN U7363 ( .A(n5999), .B(n5998), .Z(n6000) );
  NAND U7364 ( .A(n6001), .B(n6000), .Z(n6008) );
  ANDN U7365 ( .B(a[244]), .A(n3932), .Z(n6006) );
  AND U7366 ( .A(b[1]), .B(a[243]), .Z(n6005) );
  XOR U7367 ( .A(n6006), .B(n6005), .Z(n6007) );
  XNOR U7368 ( .A(n6008), .B(n6007), .Z(n6010) );
  XOR U7369 ( .A(sreg[1266]), .B(n6009), .Z(n6004) );
  XNOR U7370 ( .A(n6010), .B(n6004), .Z(c[1266]) );
  NAND U7371 ( .A(b[0]), .B(a[245]), .Z(n6013) );
  NAND U7372 ( .A(a[244]), .B(b[1]), .Z(n6012) );
  XNOR U7373 ( .A(n6013), .B(n6012), .Z(n6015) );
  XNOR U7374 ( .A(n6014), .B(n6015), .Z(n6019) );
  XOR U7375 ( .A(n6018), .B(sreg[1267]), .Z(n6011) );
  XNOR U7376 ( .A(n6019), .B(n6011), .Z(c[1267]) );
  NAND U7377 ( .A(n6013), .B(n6012), .Z(n6017) );
  NANDN U7378 ( .A(n6015), .B(n6014), .Z(n6016) );
  NAND U7379 ( .A(n6017), .B(n6016), .Z(n6024) );
  ANDN U7380 ( .B(a[246]), .A(n3932), .Z(n6022) );
  AND U7381 ( .A(b[1]), .B(a[245]), .Z(n6021) );
  XOR U7382 ( .A(n6022), .B(n6021), .Z(n6023) );
  XNOR U7383 ( .A(n6024), .B(n6023), .Z(n6026) );
  XOR U7384 ( .A(sreg[1268]), .B(n6025), .Z(n6020) );
  XNOR U7385 ( .A(n6026), .B(n6020), .Z(c[1268]) );
  NAND U7386 ( .A(b[0]), .B(a[247]), .Z(n6029) );
  NAND U7387 ( .A(a[246]), .B(b[1]), .Z(n6028) );
  XNOR U7388 ( .A(n6029), .B(n6028), .Z(n6031) );
  XNOR U7389 ( .A(n6030), .B(n6031), .Z(n6035) );
  XOR U7390 ( .A(n6034), .B(sreg[1269]), .Z(n6027) );
  XNOR U7391 ( .A(n6035), .B(n6027), .Z(c[1269]) );
  NAND U7392 ( .A(n6029), .B(n6028), .Z(n6033) );
  NANDN U7393 ( .A(n6031), .B(n6030), .Z(n6032) );
  NAND U7394 ( .A(n6033), .B(n6032), .Z(n6040) );
  ANDN U7395 ( .B(a[248]), .A(n3932), .Z(n6038) );
  AND U7396 ( .A(b[1]), .B(a[247]), .Z(n6037) );
  XOR U7397 ( .A(n6038), .B(n6037), .Z(n6039) );
  XNOR U7398 ( .A(n6040), .B(n6039), .Z(n6042) );
  XOR U7399 ( .A(sreg[1270]), .B(n6041), .Z(n6036) );
  XNOR U7400 ( .A(n6042), .B(n6036), .Z(c[1270]) );
  NAND U7401 ( .A(b[0]), .B(a[249]), .Z(n6045) );
  NAND U7402 ( .A(a[248]), .B(b[1]), .Z(n6044) );
  XNOR U7403 ( .A(n6045), .B(n6044), .Z(n6047) );
  XNOR U7404 ( .A(n6046), .B(n6047), .Z(n6051) );
  XOR U7405 ( .A(n6050), .B(sreg[1271]), .Z(n6043) );
  XNOR U7406 ( .A(n6051), .B(n6043), .Z(c[1271]) );
  NAND U7407 ( .A(n6045), .B(n6044), .Z(n6049) );
  NANDN U7408 ( .A(n6047), .B(n6046), .Z(n6048) );
  NAND U7409 ( .A(n6049), .B(n6048), .Z(n6056) );
  ANDN U7410 ( .B(a[250]), .A(n3933), .Z(n6054) );
  AND U7411 ( .A(b[1]), .B(a[249]), .Z(n6053) );
  XOR U7412 ( .A(n6054), .B(n6053), .Z(n6055) );
  XNOR U7413 ( .A(n6056), .B(n6055), .Z(n6061) );
  XOR U7414 ( .A(sreg[1272]), .B(n6060), .Z(n6052) );
  XNOR U7415 ( .A(n6061), .B(n6052), .Z(c[1272]) );
  OR U7416 ( .A(n6054), .B(n6053), .Z(n6059) );
  IV U7417 ( .A(n6055), .Z(n6057) );
  NANDN U7418 ( .A(n6057), .B(n6056), .Z(n6058) );
  NAND U7419 ( .A(n6059), .B(n6058), .Z(n6065) );
  NAND U7420 ( .A(b[0]), .B(a[251]), .Z(n6064) );
  NAND U7421 ( .A(a[250]), .B(b[1]), .Z(n6063) );
  XNOR U7422 ( .A(n6064), .B(n6063), .Z(n6066) );
  XNOR U7423 ( .A(n6065), .B(n6066), .Z(n6070) );
  XOR U7424 ( .A(n6069), .B(sreg[1273]), .Z(n6062) );
  XNOR U7425 ( .A(n6070), .B(n6062), .Z(c[1273]) );
  NAND U7426 ( .A(n6064), .B(n6063), .Z(n6068) );
  NANDN U7427 ( .A(n6066), .B(n6065), .Z(n6067) );
  NAND U7428 ( .A(n6068), .B(n6067), .Z(n6075) );
  ANDN U7429 ( .B(a[252]), .A(n3933), .Z(n6073) );
  AND U7430 ( .A(b[1]), .B(a[251]), .Z(n6072) );
  XOR U7431 ( .A(n6073), .B(n6072), .Z(n6074) );
  XNOR U7432 ( .A(n6075), .B(n6074), .Z(n6077) );
  XOR U7433 ( .A(sreg[1274]), .B(n6076), .Z(n6071) );
  XNOR U7434 ( .A(n6077), .B(n6071), .Z(c[1274]) );
  NAND U7435 ( .A(b[0]), .B(a[253]), .Z(n6080) );
  NAND U7436 ( .A(a[252]), .B(b[1]), .Z(n6079) );
  XNOR U7437 ( .A(n6080), .B(n6079), .Z(n6082) );
  XNOR U7438 ( .A(n6081), .B(n6082), .Z(n6086) );
  XOR U7439 ( .A(n6085), .B(sreg[1275]), .Z(n6078) );
  XNOR U7440 ( .A(n6086), .B(n6078), .Z(c[1275]) );
  NAND U7441 ( .A(n6080), .B(n6079), .Z(n6084) );
  NANDN U7442 ( .A(n6082), .B(n6081), .Z(n6083) );
  NAND U7443 ( .A(n6084), .B(n6083), .Z(n6091) );
  ANDN U7444 ( .B(a[254]), .A(n3933), .Z(n6089) );
  AND U7445 ( .A(b[1]), .B(a[253]), .Z(n6088) );
  XOR U7446 ( .A(n6089), .B(n6088), .Z(n6090) );
  XNOR U7447 ( .A(n6091), .B(n6090), .Z(n6093) );
  XOR U7448 ( .A(sreg[1276]), .B(n6092), .Z(n6087) );
  XNOR U7449 ( .A(n6093), .B(n6087), .Z(c[1276]) );
  NAND U7450 ( .A(b[0]), .B(a[255]), .Z(n6096) );
  NAND U7451 ( .A(a[254]), .B(b[1]), .Z(n6095) );
  XNOR U7452 ( .A(n6096), .B(n6095), .Z(n6098) );
  XNOR U7453 ( .A(n6097), .B(n6098), .Z(n6102) );
  XOR U7454 ( .A(n6101), .B(sreg[1277]), .Z(n6094) );
  XNOR U7455 ( .A(n6102), .B(n6094), .Z(c[1277]) );
  NAND U7456 ( .A(n6096), .B(n6095), .Z(n6100) );
  NANDN U7457 ( .A(n6098), .B(n6097), .Z(n6099) );
  NAND U7458 ( .A(n6100), .B(n6099), .Z(n6107) );
  ANDN U7459 ( .B(a[256]), .A(n3933), .Z(n6105) );
  AND U7460 ( .A(b[1]), .B(a[255]), .Z(n6104) );
  XOR U7461 ( .A(n6105), .B(n6104), .Z(n6106) );
  XNOR U7462 ( .A(n6107), .B(n6106), .Z(n6109) );
  XOR U7463 ( .A(sreg[1278]), .B(n6108), .Z(n6103) );
  XNOR U7464 ( .A(n6109), .B(n6103), .Z(c[1278]) );
  NAND U7465 ( .A(b[0]), .B(a[257]), .Z(n6112) );
  NAND U7466 ( .A(a[256]), .B(b[1]), .Z(n6111) );
  XNOR U7467 ( .A(n6112), .B(n6111), .Z(n6114) );
  XNOR U7468 ( .A(n6113), .B(n6114), .Z(n6118) );
  XOR U7469 ( .A(n6117), .B(sreg[1279]), .Z(n6110) );
  XNOR U7470 ( .A(n6118), .B(n6110), .Z(c[1279]) );
  NAND U7471 ( .A(n6112), .B(n6111), .Z(n6116) );
  NANDN U7472 ( .A(n6114), .B(n6113), .Z(n6115) );
  NAND U7473 ( .A(n6116), .B(n6115), .Z(n6123) );
  ANDN U7474 ( .B(a[258]), .A(n3933), .Z(n6121) );
  AND U7475 ( .A(b[1]), .B(a[257]), .Z(n6120) );
  XOR U7476 ( .A(n6121), .B(n6120), .Z(n6122) );
  XNOR U7477 ( .A(n6123), .B(n6122), .Z(n6125) );
  XOR U7478 ( .A(sreg[1280]), .B(n6124), .Z(n6119) );
  XNOR U7479 ( .A(n6125), .B(n6119), .Z(c[1280]) );
  ANDN U7480 ( .B(a[259]), .A(n3933), .Z(n6128) );
  AND U7481 ( .A(b[1]), .B(a[258]), .Z(n6127) );
  XOR U7482 ( .A(n6128), .B(n6127), .Z(n6129) );
  XNOR U7483 ( .A(n6130), .B(n6129), .Z(n6132) );
  XNOR U7484 ( .A(sreg[1281]), .B(n6131), .Z(n6126) );
  XNOR U7485 ( .A(n6132), .B(n6126), .Z(c[1281]) );
  ANDN U7486 ( .B(a[260]), .A(n3933), .Z(n6135) );
  AND U7487 ( .A(b[1]), .B(a[259]), .Z(n6134) );
  XOR U7488 ( .A(n6135), .B(n6134), .Z(n6136) );
  XNOR U7489 ( .A(n6137), .B(n6136), .Z(n6139) );
  XNOR U7490 ( .A(sreg[1282]), .B(n6138), .Z(n6133) );
  XNOR U7491 ( .A(n6139), .B(n6133), .Z(c[1282]) );
  NAND U7492 ( .A(b[0]), .B(a[261]), .Z(n6142) );
  NAND U7493 ( .A(a[260]), .B(b[1]), .Z(n6141) );
  XNOR U7494 ( .A(n6142), .B(n6141), .Z(n6144) );
  XNOR U7495 ( .A(n6143), .B(n6144), .Z(n6148) );
  XOR U7496 ( .A(n6147), .B(sreg[1283]), .Z(n6140) );
  XNOR U7497 ( .A(n6148), .B(n6140), .Z(c[1283]) );
  NAND U7498 ( .A(n6142), .B(n6141), .Z(n6146) );
  NANDN U7499 ( .A(n6144), .B(n6143), .Z(n6145) );
  NAND U7500 ( .A(n6146), .B(n6145), .Z(n6153) );
  ANDN U7501 ( .B(a[262]), .A(n3934), .Z(n6151) );
  AND U7502 ( .A(b[1]), .B(a[261]), .Z(n6150) );
  XOR U7503 ( .A(n6151), .B(n6150), .Z(n6152) );
  XNOR U7504 ( .A(n6153), .B(n6152), .Z(n6158) );
  XOR U7505 ( .A(sreg[1284]), .B(n6157), .Z(n6149) );
  XNOR U7506 ( .A(n6158), .B(n6149), .Z(c[1284]) );
  OR U7507 ( .A(n6151), .B(n6150), .Z(n6156) );
  IV U7508 ( .A(n6152), .Z(n6154) );
  NANDN U7509 ( .A(n6154), .B(n6153), .Z(n6155) );
  NAND U7510 ( .A(n6156), .B(n6155), .Z(n6163) );
  ANDN U7511 ( .B(a[263]), .A(n3934), .Z(n6161) );
  AND U7512 ( .A(b[1]), .B(a[262]), .Z(n6160) );
  XOR U7513 ( .A(n6161), .B(n6160), .Z(n6162) );
  XNOR U7514 ( .A(n6163), .B(n6162), .Z(n6165) );
  XNOR U7515 ( .A(sreg[1285]), .B(n6164), .Z(n6159) );
  XNOR U7516 ( .A(n6165), .B(n6159), .Z(c[1285]) );
  ANDN U7517 ( .B(a[264]), .A(n3934), .Z(n6168) );
  AND U7518 ( .A(b[1]), .B(a[263]), .Z(n6167) );
  XOR U7519 ( .A(n6168), .B(n6167), .Z(n6169) );
  XNOR U7520 ( .A(n6170), .B(n6169), .Z(n6172) );
  XNOR U7521 ( .A(sreg[1286]), .B(n6171), .Z(n6166) );
  XNOR U7522 ( .A(n6172), .B(n6166), .Z(c[1286]) );
  NAND U7523 ( .A(b[0]), .B(a[265]), .Z(n6175) );
  NAND U7524 ( .A(a[264]), .B(b[1]), .Z(n6174) );
  XNOR U7525 ( .A(n6175), .B(n6174), .Z(n6177) );
  XNOR U7526 ( .A(n6176), .B(n6177), .Z(n6181) );
  XOR U7527 ( .A(n6180), .B(sreg[1287]), .Z(n6173) );
  XNOR U7528 ( .A(n6181), .B(n6173), .Z(c[1287]) );
  NAND U7529 ( .A(n6175), .B(n6174), .Z(n6179) );
  NANDN U7530 ( .A(n6177), .B(n6176), .Z(n6178) );
  NAND U7531 ( .A(n6179), .B(n6178), .Z(n6185) );
  NAND U7532 ( .A(b[0]), .B(a[266]), .Z(n6184) );
  NAND U7533 ( .A(a[265]), .B(b[1]), .Z(n6183) );
  XNOR U7534 ( .A(n6184), .B(n6183), .Z(n6186) );
  XNOR U7535 ( .A(n6185), .B(n6186), .Z(n6190) );
  XOR U7536 ( .A(n6189), .B(sreg[1288]), .Z(n6182) );
  XNOR U7537 ( .A(n6190), .B(n6182), .Z(c[1288]) );
  NAND U7538 ( .A(n6184), .B(n6183), .Z(n6188) );
  NANDN U7539 ( .A(n6186), .B(n6185), .Z(n6187) );
  NAND U7540 ( .A(n6188), .B(n6187), .Z(n6194) );
  NAND U7541 ( .A(b[0]), .B(a[267]), .Z(n6193) );
  NAND U7542 ( .A(a[266]), .B(b[1]), .Z(n6192) );
  XNOR U7543 ( .A(n6193), .B(n6192), .Z(n6195) );
  XNOR U7544 ( .A(n6194), .B(n6195), .Z(n6199) );
  XOR U7545 ( .A(n6198), .B(sreg[1289]), .Z(n6191) );
  XNOR U7546 ( .A(n6199), .B(n6191), .Z(c[1289]) );
  NAND U7547 ( .A(n6193), .B(n6192), .Z(n6197) );
  NANDN U7548 ( .A(n6195), .B(n6194), .Z(n6196) );
  NAND U7549 ( .A(n6197), .B(n6196), .Z(n6204) );
  ANDN U7550 ( .B(a[268]), .A(n3934), .Z(n6202) );
  AND U7551 ( .A(b[1]), .B(a[267]), .Z(n6201) );
  XOR U7552 ( .A(n6202), .B(n6201), .Z(n6203) );
  XNOR U7553 ( .A(n6204), .B(n6203), .Z(n6206) );
  XOR U7554 ( .A(sreg[1290]), .B(n6205), .Z(n6200) );
  XNOR U7555 ( .A(n6206), .B(n6200), .Z(c[1290]) );
  ANDN U7556 ( .B(a[269]), .A(n3934), .Z(n6209) );
  AND U7557 ( .A(b[1]), .B(a[268]), .Z(n6208) );
  XOR U7558 ( .A(n6209), .B(n6208), .Z(n6210) );
  XNOR U7559 ( .A(n6211), .B(n6210), .Z(n6213) );
  XNOR U7560 ( .A(sreg[1291]), .B(n6212), .Z(n6207) );
  XNOR U7561 ( .A(n6213), .B(n6207), .Z(c[1291]) );
  ANDN U7562 ( .B(a[270]), .A(n3934), .Z(n6216) );
  AND U7563 ( .A(b[1]), .B(a[269]), .Z(n6215) );
  XOR U7564 ( .A(n6216), .B(n6215), .Z(n6217) );
  XNOR U7565 ( .A(n6218), .B(n6217), .Z(n6220) );
  XNOR U7566 ( .A(sreg[1292]), .B(n6219), .Z(n6214) );
  XNOR U7567 ( .A(n6220), .B(n6214), .Z(c[1292]) );
  NAND U7568 ( .A(b[0]), .B(a[271]), .Z(n6223) );
  NAND U7569 ( .A(a[270]), .B(b[1]), .Z(n6222) );
  XNOR U7570 ( .A(n6223), .B(n6222), .Z(n6225) );
  XNOR U7571 ( .A(n6224), .B(n6225), .Z(n6229) );
  XOR U7572 ( .A(n6228), .B(sreg[1293]), .Z(n6221) );
  XNOR U7573 ( .A(n6229), .B(n6221), .Z(c[1293]) );
  NAND U7574 ( .A(n6223), .B(n6222), .Z(n6227) );
  NANDN U7575 ( .A(n6225), .B(n6224), .Z(n6226) );
  NAND U7576 ( .A(n6227), .B(n6226), .Z(n6234) );
  ANDN U7577 ( .B(a[272]), .A(n3934), .Z(n6232) );
  AND U7578 ( .A(b[1]), .B(a[271]), .Z(n6231) );
  XOR U7579 ( .A(n6232), .B(n6231), .Z(n6233) );
  XNOR U7580 ( .A(n6234), .B(n6233), .Z(n6236) );
  XOR U7581 ( .A(sreg[1294]), .B(n6235), .Z(n6230) );
  XNOR U7582 ( .A(n6236), .B(n6230), .Z(c[1294]) );
  NAND U7583 ( .A(b[0]), .B(a[273]), .Z(n6239) );
  NAND U7584 ( .A(a[272]), .B(b[1]), .Z(n6238) );
  XNOR U7585 ( .A(n6239), .B(n6238), .Z(n6241) );
  XNOR U7586 ( .A(n6240), .B(n6241), .Z(n6245) );
  XOR U7587 ( .A(n6244), .B(sreg[1295]), .Z(n6237) );
  XNOR U7588 ( .A(n6245), .B(n6237), .Z(c[1295]) );
  NAND U7589 ( .A(n6239), .B(n6238), .Z(n6243) );
  NANDN U7590 ( .A(n6241), .B(n6240), .Z(n6242) );
  NAND U7591 ( .A(n6243), .B(n6242), .Z(n6250) );
  ANDN U7592 ( .B(a[274]), .A(n3935), .Z(n6248) );
  AND U7593 ( .A(b[1]), .B(a[273]), .Z(n6247) );
  XOR U7594 ( .A(n6248), .B(n6247), .Z(n6249) );
  XNOR U7595 ( .A(n6250), .B(n6249), .Z(n6255) );
  XOR U7596 ( .A(sreg[1296]), .B(n6254), .Z(n6246) );
  XNOR U7597 ( .A(n6255), .B(n6246), .Z(c[1296]) );
  OR U7598 ( .A(n6248), .B(n6247), .Z(n6253) );
  IV U7599 ( .A(n6249), .Z(n6251) );
  NANDN U7600 ( .A(n6251), .B(n6250), .Z(n6252) );
  NAND U7601 ( .A(n6253), .B(n6252), .Z(n6259) );
  NAND U7602 ( .A(b[0]), .B(a[275]), .Z(n6258) );
  NAND U7603 ( .A(a[274]), .B(b[1]), .Z(n6257) );
  XNOR U7604 ( .A(n6258), .B(n6257), .Z(n6260) );
  XNOR U7605 ( .A(n6259), .B(n6260), .Z(n6264) );
  XOR U7606 ( .A(n6263), .B(sreg[1297]), .Z(n6256) );
  XNOR U7607 ( .A(n6264), .B(n6256), .Z(c[1297]) );
  NAND U7608 ( .A(n6258), .B(n6257), .Z(n6262) );
  NANDN U7609 ( .A(n6260), .B(n6259), .Z(n6261) );
  NAND U7610 ( .A(n6262), .B(n6261), .Z(n6268) );
  NAND U7611 ( .A(b[0]), .B(a[276]), .Z(n6267) );
  NAND U7612 ( .A(a[275]), .B(b[1]), .Z(n6266) );
  XNOR U7613 ( .A(n6267), .B(n6266), .Z(n6269) );
  XNOR U7614 ( .A(n6268), .B(n6269), .Z(n6273) );
  XOR U7615 ( .A(n6272), .B(sreg[1298]), .Z(n6265) );
  XNOR U7616 ( .A(n6273), .B(n6265), .Z(c[1298]) );
  NAND U7617 ( .A(n6267), .B(n6266), .Z(n6271) );
  NANDN U7618 ( .A(n6269), .B(n6268), .Z(n6270) );
  NAND U7619 ( .A(n6271), .B(n6270), .Z(n6277) );
  NAND U7620 ( .A(b[0]), .B(a[277]), .Z(n6276) );
  NAND U7621 ( .A(a[276]), .B(b[1]), .Z(n6275) );
  XNOR U7622 ( .A(n6276), .B(n6275), .Z(n6278) );
  XNOR U7623 ( .A(n6277), .B(n6278), .Z(n6282) );
  XOR U7624 ( .A(n6281), .B(sreg[1299]), .Z(n6274) );
  XNOR U7625 ( .A(n6282), .B(n6274), .Z(c[1299]) );
  NAND U7626 ( .A(n6276), .B(n6275), .Z(n6280) );
  NANDN U7627 ( .A(n6278), .B(n6277), .Z(n6279) );
  NAND U7628 ( .A(n6280), .B(n6279), .Z(n6287) );
  ANDN U7629 ( .B(a[278]), .A(n3935), .Z(n6285) );
  AND U7630 ( .A(b[1]), .B(a[277]), .Z(n6284) );
  XOR U7631 ( .A(n6285), .B(n6284), .Z(n6286) );
  XNOR U7632 ( .A(n6287), .B(n6286), .Z(n6289) );
  XOR U7633 ( .A(sreg[1300]), .B(n6288), .Z(n6283) );
  XNOR U7634 ( .A(n6289), .B(n6283), .Z(c[1300]) );
  NAND U7635 ( .A(b[0]), .B(a[279]), .Z(n6292) );
  NAND U7636 ( .A(a[278]), .B(b[1]), .Z(n6291) );
  XNOR U7637 ( .A(n6292), .B(n6291), .Z(n6294) );
  XNOR U7638 ( .A(n6293), .B(n6294), .Z(n6298) );
  XOR U7639 ( .A(n6297), .B(sreg[1301]), .Z(n6290) );
  XNOR U7640 ( .A(n6298), .B(n6290), .Z(c[1301]) );
  NAND U7641 ( .A(n6292), .B(n6291), .Z(n6296) );
  NANDN U7642 ( .A(n6294), .B(n6293), .Z(n6295) );
  NAND U7643 ( .A(n6296), .B(n6295), .Z(n6303) );
  ANDN U7644 ( .B(a[280]), .A(n3935), .Z(n6301) );
  AND U7645 ( .A(b[1]), .B(a[279]), .Z(n6300) );
  XOR U7646 ( .A(n6301), .B(n6300), .Z(n6302) );
  XNOR U7647 ( .A(n6303), .B(n6302), .Z(n6305) );
  XOR U7648 ( .A(sreg[1302]), .B(n6304), .Z(n6299) );
  XNOR U7649 ( .A(n6305), .B(n6299), .Z(c[1302]) );
  NAND U7650 ( .A(b[0]), .B(a[281]), .Z(n6308) );
  NAND U7651 ( .A(a[280]), .B(b[1]), .Z(n6307) );
  XNOR U7652 ( .A(n6308), .B(n6307), .Z(n6310) );
  XNOR U7653 ( .A(n6309), .B(n6310), .Z(n6314) );
  XOR U7654 ( .A(n6313), .B(sreg[1303]), .Z(n6306) );
  XNOR U7655 ( .A(n6314), .B(n6306), .Z(c[1303]) );
  NAND U7656 ( .A(n6308), .B(n6307), .Z(n6312) );
  NANDN U7657 ( .A(n6310), .B(n6309), .Z(n6311) );
  NAND U7658 ( .A(n6312), .B(n6311), .Z(n6319) );
  ANDN U7659 ( .B(a[282]), .A(n3935), .Z(n6317) );
  AND U7660 ( .A(b[1]), .B(a[281]), .Z(n6316) );
  XOR U7661 ( .A(n6317), .B(n6316), .Z(n6318) );
  XNOR U7662 ( .A(n6319), .B(n6318), .Z(n6321) );
  XOR U7663 ( .A(sreg[1304]), .B(n6320), .Z(n6315) );
  XNOR U7664 ( .A(n6321), .B(n6315), .Z(c[1304]) );
  NAND U7665 ( .A(b[0]), .B(a[283]), .Z(n6324) );
  NAND U7666 ( .A(a[282]), .B(b[1]), .Z(n6323) );
  XNOR U7667 ( .A(n6324), .B(n6323), .Z(n6326) );
  XNOR U7668 ( .A(n6325), .B(n6326), .Z(n6330) );
  XOR U7669 ( .A(n6329), .B(sreg[1305]), .Z(n6322) );
  XNOR U7670 ( .A(n6330), .B(n6322), .Z(c[1305]) );
  NAND U7671 ( .A(n6324), .B(n6323), .Z(n6328) );
  NANDN U7672 ( .A(n6326), .B(n6325), .Z(n6327) );
  NAND U7673 ( .A(n6328), .B(n6327), .Z(n6335) );
  ANDN U7674 ( .B(a[284]), .A(n3935), .Z(n6333) );
  AND U7675 ( .A(b[1]), .B(a[283]), .Z(n6332) );
  XOR U7676 ( .A(n6333), .B(n6332), .Z(n6334) );
  XNOR U7677 ( .A(n6335), .B(n6334), .Z(n6337) );
  XOR U7678 ( .A(sreg[1306]), .B(n6336), .Z(n6331) );
  XNOR U7679 ( .A(n6337), .B(n6331), .Z(c[1306]) );
  NAND U7680 ( .A(b[0]), .B(a[285]), .Z(n6340) );
  NAND U7681 ( .A(a[284]), .B(b[1]), .Z(n6339) );
  XNOR U7682 ( .A(n6340), .B(n6339), .Z(n6342) );
  XNOR U7683 ( .A(n6341), .B(n6342), .Z(n6346) );
  XOR U7684 ( .A(n6345), .B(sreg[1307]), .Z(n6338) );
  XNOR U7685 ( .A(n6346), .B(n6338), .Z(c[1307]) );
  NAND U7686 ( .A(n6340), .B(n6339), .Z(n6344) );
  NANDN U7687 ( .A(n6342), .B(n6341), .Z(n6343) );
  NAND U7688 ( .A(n6344), .B(n6343), .Z(n6350) );
  NAND U7689 ( .A(b[0]), .B(a[286]), .Z(n6349) );
  NAND U7690 ( .A(a[285]), .B(b[1]), .Z(n6348) );
  XNOR U7691 ( .A(n6349), .B(n6348), .Z(n6351) );
  XNOR U7692 ( .A(n6350), .B(n6351), .Z(n6355) );
  XOR U7693 ( .A(n6354), .B(sreg[1308]), .Z(n6347) );
  XNOR U7694 ( .A(n6355), .B(n6347), .Z(c[1308]) );
  NAND U7695 ( .A(n6349), .B(n6348), .Z(n6353) );
  NANDN U7696 ( .A(n6351), .B(n6350), .Z(n6352) );
  NAND U7697 ( .A(n6353), .B(n6352), .Z(n6359) );
  NAND U7698 ( .A(b[0]), .B(a[287]), .Z(n6358) );
  NAND U7699 ( .A(a[286]), .B(b[1]), .Z(n6357) );
  XNOR U7700 ( .A(n6358), .B(n6357), .Z(n6360) );
  XNOR U7701 ( .A(n6359), .B(n6360), .Z(n6364) );
  XOR U7702 ( .A(n6363), .B(sreg[1309]), .Z(n6356) );
  XNOR U7703 ( .A(n6364), .B(n6356), .Z(c[1309]) );
  NAND U7704 ( .A(n6358), .B(n6357), .Z(n6362) );
  NANDN U7705 ( .A(n6360), .B(n6359), .Z(n6361) );
  NAND U7706 ( .A(n6362), .B(n6361), .Z(n6369) );
  ANDN U7707 ( .B(a[288]), .A(n3935), .Z(n6367) );
  AND U7708 ( .A(b[1]), .B(a[287]), .Z(n6366) );
  XOR U7709 ( .A(n6367), .B(n6366), .Z(n6368) );
  XNOR U7710 ( .A(n6369), .B(n6368), .Z(n6371) );
  XOR U7711 ( .A(sreg[1310]), .B(n6370), .Z(n6365) );
  XNOR U7712 ( .A(n6371), .B(n6365), .Z(c[1310]) );
  NAND U7713 ( .A(b[0]), .B(a[289]), .Z(n6374) );
  NAND U7714 ( .A(a[288]), .B(b[1]), .Z(n6373) );
  XNOR U7715 ( .A(n6374), .B(n6373), .Z(n6376) );
  XNOR U7716 ( .A(n6375), .B(n6376), .Z(n6380) );
  XOR U7717 ( .A(n6379), .B(sreg[1311]), .Z(n6372) );
  XNOR U7718 ( .A(n6380), .B(n6372), .Z(c[1311]) );
  NAND U7719 ( .A(n6374), .B(n6373), .Z(n6378) );
  NANDN U7720 ( .A(n6376), .B(n6375), .Z(n6377) );
  NAND U7721 ( .A(n6378), .B(n6377), .Z(n6385) );
  ANDN U7722 ( .B(a[290]), .A(n3935), .Z(n6383) );
  AND U7723 ( .A(b[1]), .B(a[289]), .Z(n6382) );
  XOR U7724 ( .A(n6383), .B(n6382), .Z(n6384) );
  XNOR U7725 ( .A(n6385), .B(n6384), .Z(n6387) );
  XOR U7726 ( .A(sreg[1312]), .B(n6386), .Z(n6381) );
  XNOR U7727 ( .A(n6387), .B(n6381), .Z(c[1312]) );
  NAND U7728 ( .A(b[0]), .B(a[291]), .Z(n6390) );
  NAND U7729 ( .A(a[290]), .B(b[1]), .Z(n6389) );
  XNOR U7730 ( .A(n6390), .B(n6389), .Z(n6392) );
  XNOR U7731 ( .A(n6391), .B(n6392), .Z(n6396) );
  XOR U7732 ( .A(n6395), .B(sreg[1313]), .Z(n6388) );
  XNOR U7733 ( .A(n6396), .B(n6388), .Z(c[1313]) );
  NAND U7734 ( .A(n6390), .B(n6389), .Z(n6394) );
  NANDN U7735 ( .A(n6392), .B(n6391), .Z(n6393) );
  NAND U7736 ( .A(n6394), .B(n6393), .Z(n6400) );
  NAND U7737 ( .A(b[0]), .B(a[292]), .Z(n6399) );
  NAND U7738 ( .A(a[291]), .B(b[1]), .Z(n6398) );
  XNOR U7739 ( .A(n6399), .B(n6398), .Z(n6401) );
  XNOR U7740 ( .A(n6400), .B(n6401), .Z(n6405) );
  XOR U7741 ( .A(n6404), .B(sreg[1314]), .Z(n6397) );
  XNOR U7742 ( .A(n6405), .B(n6397), .Z(c[1314]) );
  NAND U7743 ( .A(n6399), .B(n6398), .Z(n6403) );
  NANDN U7744 ( .A(n6401), .B(n6400), .Z(n6402) );
  NAND U7745 ( .A(n6403), .B(n6402), .Z(n6409) );
  NAND U7746 ( .A(b[0]), .B(a[293]), .Z(n6408) );
  NAND U7747 ( .A(a[292]), .B(b[1]), .Z(n6407) );
  XNOR U7748 ( .A(n6408), .B(n6407), .Z(n6410) );
  XNOR U7749 ( .A(n6409), .B(n6410), .Z(n6414) );
  XOR U7750 ( .A(n6413), .B(sreg[1315]), .Z(n6406) );
  XNOR U7751 ( .A(n6414), .B(n6406), .Z(c[1315]) );
  NAND U7752 ( .A(n6408), .B(n6407), .Z(n6412) );
  NANDN U7753 ( .A(n6410), .B(n6409), .Z(n6411) );
  NAND U7754 ( .A(n6412), .B(n6411), .Z(n6419) );
  ANDN U7755 ( .B(a[294]), .A(n3936), .Z(n6417) );
  AND U7756 ( .A(b[1]), .B(a[293]), .Z(n6416) );
  XOR U7757 ( .A(n6417), .B(n6416), .Z(n6418) );
  XNOR U7758 ( .A(n6419), .B(n6418), .Z(n6424) );
  XOR U7759 ( .A(sreg[1316]), .B(n6423), .Z(n6415) );
  XNOR U7760 ( .A(n6424), .B(n6415), .Z(c[1316]) );
  OR U7761 ( .A(n6417), .B(n6416), .Z(n6422) );
  IV U7762 ( .A(n6418), .Z(n6420) );
  NANDN U7763 ( .A(n6420), .B(n6419), .Z(n6421) );
  NAND U7764 ( .A(n6422), .B(n6421), .Z(n6428) );
  NAND U7765 ( .A(b[0]), .B(a[295]), .Z(n6427) );
  NAND U7766 ( .A(a[294]), .B(b[1]), .Z(n6426) );
  XNOR U7767 ( .A(n6427), .B(n6426), .Z(n6429) );
  XNOR U7768 ( .A(n6428), .B(n6429), .Z(n6433) );
  XOR U7769 ( .A(n6432), .B(sreg[1317]), .Z(n6425) );
  XNOR U7770 ( .A(n6433), .B(n6425), .Z(c[1317]) );
  NAND U7771 ( .A(n6427), .B(n6426), .Z(n6431) );
  NANDN U7772 ( .A(n6429), .B(n6428), .Z(n6430) );
  NAND U7773 ( .A(n6431), .B(n6430), .Z(n6438) );
  ANDN U7774 ( .B(a[296]), .A(n3936), .Z(n6436) );
  AND U7775 ( .A(b[1]), .B(a[295]), .Z(n6435) );
  XOR U7776 ( .A(n6436), .B(n6435), .Z(n6437) );
  XNOR U7777 ( .A(n6438), .B(n6437), .Z(n6440) );
  XOR U7778 ( .A(sreg[1318]), .B(n6439), .Z(n6434) );
  XNOR U7779 ( .A(n6440), .B(n6434), .Z(c[1318]) );
  NAND U7780 ( .A(b[0]), .B(a[297]), .Z(n6443) );
  NAND U7781 ( .A(a[296]), .B(b[1]), .Z(n6442) );
  XNOR U7782 ( .A(n6443), .B(n6442), .Z(n6445) );
  XNOR U7783 ( .A(n6444), .B(n6445), .Z(n6449) );
  XOR U7784 ( .A(n6448), .B(sreg[1319]), .Z(n6441) );
  XNOR U7785 ( .A(n6449), .B(n6441), .Z(c[1319]) );
  NAND U7786 ( .A(n6443), .B(n6442), .Z(n6447) );
  NANDN U7787 ( .A(n6445), .B(n6444), .Z(n6446) );
  NAND U7788 ( .A(n6447), .B(n6446), .Z(n6454) );
  ANDN U7789 ( .B(a[298]), .A(n3936), .Z(n6452) );
  AND U7790 ( .A(b[1]), .B(a[297]), .Z(n6451) );
  XOR U7791 ( .A(n6452), .B(n6451), .Z(n6453) );
  XNOR U7792 ( .A(n6454), .B(n6453), .Z(n6456) );
  XOR U7793 ( .A(sreg[1320]), .B(n6455), .Z(n6450) );
  XNOR U7794 ( .A(n6456), .B(n6450), .Z(c[1320]) );
  NAND U7795 ( .A(b[0]), .B(a[299]), .Z(n6459) );
  NAND U7796 ( .A(a[298]), .B(b[1]), .Z(n6458) );
  XNOR U7797 ( .A(n6459), .B(n6458), .Z(n6461) );
  XNOR U7798 ( .A(n6460), .B(n6461), .Z(n6465) );
  XOR U7799 ( .A(n6464), .B(sreg[1321]), .Z(n6457) );
  XNOR U7800 ( .A(n6465), .B(n6457), .Z(c[1321]) );
  NAND U7801 ( .A(n6459), .B(n6458), .Z(n6463) );
  NANDN U7802 ( .A(n6461), .B(n6460), .Z(n6462) );
  NAND U7803 ( .A(n6463), .B(n6462), .Z(n6470) );
  ANDN U7804 ( .B(a[300]), .A(n3936), .Z(n6468) );
  AND U7805 ( .A(b[1]), .B(a[299]), .Z(n6467) );
  XOR U7806 ( .A(n6468), .B(n6467), .Z(n6469) );
  XNOR U7807 ( .A(n6470), .B(n6469), .Z(n6472) );
  XOR U7808 ( .A(sreg[1322]), .B(n6471), .Z(n6466) );
  XNOR U7809 ( .A(n6472), .B(n6466), .Z(c[1322]) );
  NAND U7810 ( .A(b[0]), .B(a[301]), .Z(n6475) );
  NAND U7811 ( .A(a[300]), .B(b[1]), .Z(n6474) );
  XNOR U7812 ( .A(n6475), .B(n6474), .Z(n6477) );
  XNOR U7813 ( .A(n6476), .B(n6477), .Z(n6481) );
  XOR U7814 ( .A(n6480), .B(sreg[1323]), .Z(n6473) );
  XNOR U7815 ( .A(n6481), .B(n6473), .Z(c[1323]) );
  NAND U7816 ( .A(n6475), .B(n6474), .Z(n6479) );
  NANDN U7817 ( .A(n6477), .B(n6476), .Z(n6478) );
  NAND U7818 ( .A(n6479), .B(n6478), .Z(n6486) );
  ANDN U7819 ( .B(a[302]), .A(n3936), .Z(n6484) );
  AND U7820 ( .A(b[1]), .B(a[301]), .Z(n6483) );
  XOR U7821 ( .A(n6484), .B(n6483), .Z(n6485) );
  XNOR U7822 ( .A(n6486), .B(n6485), .Z(n6488) );
  XOR U7823 ( .A(sreg[1324]), .B(n6487), .Z(n6482) );
  XNOR U7824 ( .A(n6488), .B(n6482), .Z(c[1324]) );
  NAND U7825 ( .A(b[0]), .B(a[303]), .Z(n6491) );
  NAND U7826 ( .A(a[302]), .B(b[1]), .Z(n6490) );
  XNOR U7827 ( .A(n6491), .B(n6490), .Z(n6493) );
  XNOR U7828 ( .A(n6492), .B(n6493), .Z(n6497) );
  XOR U7829 ( .A(n6496), .B(sreg[1325]), .Z(n6489) );
  XNOR U7830 ( .A(n6497), .B(n6489), .Z(c[1325]) );
  NAND U7831 ( .A(n6491), .B(n6490), .Z(n6495) );
  NANDN U7832 ( .A(n6493), .B(n6492), .Z(n6494) );
  NAND U7833 ( .A(n6495), .B(n6494), .Z(n6502) );
  ANDN U7834 ( .B(a[304]), .A(n3936), .Z(n6500) );
  AND U7835 ( .A(b[1]), .B(a[303]), .Z(n6499) );
  XOR U7836 ( .A(n6500), .B(n6499), .Z(n6501) );
  XNOR U7837 ( .A(n6502), .B(n6501), .Z(n6504) );
  XOR U7838 ( .A(sreg[1326]), .B(n6503), .Z(n6498) );
  XNOR U7839 ( .A(n6504), .B(n6498), .Z(c[1326]) );
  NAND U7840 ( .A(b[0]), .B(a[305]), .Z(n6507) );
  NAND U7841 ( .A(a[304]), .B(b[1]), .Z(n6506) );
  XNOR U7842 ( .A(n6507), .B(n6506), .Z(n6509) );
  XNOR U7843 ( .A(n6508), .B(n6509), .Z(n6513) );
  XOR U7844 ( .A(n6512), .B(sreg[1327]), .Z(n6505) );
  XNOR U7845 ( .A(n6513), .B(n6505), .Z(c[1327]) );
  NAND U7846 ( .A(n6507), .B(n6506), .Z(n6511) );
  NANDN U7847 ( .A(n6509), .B(n6508), .Z(n6510) );
  NAND U7848 ( .A(n6511), .B(n6510), .Z(n6518) );
  ANDN U7849 ( .B(a[306]), .A(n3936), .Z(n6516) );
  AND U7850 ( .A(b[1]), .B(a[305]), .Z(n6515) );
  XOR U7851 ( .A(n6516), .B(n6515), .Z(n6517) );
  XNOR U7852 ( .A(n6518), .B(n6517), .Z(n6520) );
  XOR U7853 ( .A(sreg[1328]), .B(n6519), .Z(n6514) );
  XNOR U7854 ( .A(n6520), .B(n6514), .Z(c[1328]) );
  NAND U7855 ( .A(b[0]), .B(a[307]), .Z(n6523) );
  NAND U7856 ( .A(a[306]), .B(b[1]), .Z(n6522) );
  XNOR U7857 ( .A(n6523), .B(n6522), .Z(n6525) );
  XNOR U7858 ( .A(n6524), .B(n6525), .Z(n6529) );
  XOR U7859 ( .A(n6528), .B(sreg[1329]), .Z(n6521) );
  XNOR U7860 ( .A(n6529), .B(n6521), .Z(c[1329]) );
  NAND U7861 ( .A(n6523), .B(n6522), .Z(n6527) );
  NANDN U7862 ( .A(n6525), .B(n6524), .Z(n6526) );
  NAND U7863 ( .A(n6527), .B(n6526), .Z(n6534) );
  ANDN U7864 ( .B(a[308]), .A(n3937), .Z(n6532) );
  AND U7865 ( .A(b[1]), .B(a[307]), .Z(n6531) );
  XOR U7866 ( .A(n6532), .B(n6531), .Z(n6533) );
  XNOR U7867 ( .A(n6534), .B(n6533), .Z(n6539) );
  XOR U7868 ( .A(sreg[1330]), .B(n6538), .Z(n6530) );
  XNOR U7869 ( .A(n6539), .B(n6530), .Z(c[1330]) );
  OR U7870 ( .A(n6532), .B(n6531), .Z(n6537) );
  IV U7871 ( .A(n6533), .Z(n6535) );
  NANDN U7872 ( .A(n6535), .B(n6534), .Z(n6536) );
  NAND U7873 ( .A(n6537), .B(n6536), .Z(n6543) );
  NAND U7874 ( .A(b[0]), .B(a[309]), .Z(n6542) );
  NAND U7875 ( .A(a[308]), .B(b[1]), .Z(n6541) );
  XNOR U7876 ( .A(n6542), .B(n6541), .Z(n6544) );
  XNOR U7877 ( .A(n6543), .B(n6544), .Z(n6548) );
  XOR U7878 ( .A(n6547), .B(sreg[1331]), .Z(n6540) );
  XNOR U7879 ( .A(n6548), .B(n6540), .Z(c[1331]) );
  NAND U7880 ( .A(n6542), .B(n6541), .Z(n6546) );
  NANDN U7881 ( .A(n6544), .B(n6543), .Z(n6545) );
  NAND U7882 ( .A(n6546), .B(n6545), .Z(n6553) );
  ANDN U7883 ( .B(a[310]), .A(n3937), .Z(n6551) );
  AND U7884 ( .A(b[1]), .B(a[309]), .Z(n6550) );
  XOR U7885 ( .A(n6551), .B(n6550), .Z(n6552) );
  XNOR U7886 ( .A(n6553), .B(n6552), .Z(n6555) );
  XOR U7887 ( .A(sreg[1332]), .B(n6554), .Z(n6549) );
  XNOR U7888 ( .A(n6555), .B(n6549), .Z(c[1332]) );
  NAND U7889 ( .A(b[0]), .B(a[311]), .Z(n6558) );
  NAND U7890 ( .A(a[310]), .B(b[1]), .Z(n6557) );
  XNOR U7891 ( .A(n6558), .B(n6557), .Z(n6560) );
  XNOR U7892 ( .A(n6559), .B(n6560), .Z(n6564) );
  XOR U7893 ( .A(n6563), .B(sreg[1333]), .Z(n6556) );
  XNOR U7894 ( .A(n6564), .B(n6556), .Z(c[1333]) );
  NAND U7895 ( .A(n6558), .B(n6557), .Z(n6562) );
  NANDN U7896 ( .A(n6560), .B(n6559), .Z(n6561) );
  NAND U7897 ( .A(n6562), .B(n6561), .Z(n6569) );
  ANDN U7898 ( .B(a[312]), .A(n3937), .Z(n6567) );
  AND U7899 ( .A(b[1]), .B(a[311]), .Z(n6566) );
  XOR U7900 ( .A(n6567), .B(n6566), .Z(n6568) );
  XNOR U7901 ( .A(n6569), .B(n6568), .Z(n6571) );
  XOR U7902 ( .A(sreg[1334]), .B(n6570), .Z(n6565) );
  XNOR U7903 ( .A(n6571), .B(n6565), .Z(c[1334]) );
  NAND U7904 ( .A(b[0]), .B(a[313]), .Z(n6574) );
  NAND U7905 ( .A(a[312]), .B(b[1]), .Z(n6573) );
  XNOR U7906 ( .A(n6574), .B(n6573), .Z(n6576) );
  XNOR U7907 ( .A(n6575), .B(n6576), .Z(n6580) );
  XOR U7908 ( .A(n6579), .B(sreg[1335]), .Z(n6572) );
  XNOR U7909 ( .A(n6580), .B(n6572), .Z(c[1335]) );
  NAND U7910 ( .A(n6574), .B(n6573), .Z(n6578) );
  NANDN U7911 ( .A(n6576), .B(n6575), .Z(n6577) );
  NAND U7912 ( .A(n6578), .B(n6577), .Z(n6585) );
  ANDN U7913 ( .B(a[314]), .A(n3937), .Z(n6583) );
  AND U7914 ( .A(b[1]), .B(a[313]), .Z(n6582) );
  XOR U7915 ( .A(n6583), .B(n6582), .Z(n6584) );
  XNOR U7916 ( .A(n6585), .B(n6584), .Z(n6587) );
  XOR U7917 ( .A(sreg[1336]), .B(n6586), .Z(n6581) );
  XNOR U7918 ( .A(n6587), .B(n6581), .Z(c[1336]) );
  NAND U7919 ( .A(b[0]), .B(a[315]), .Z(n6590) );
  NAND U7920 ( .A(a[314]), .B(b[1]), .Z(n6589) );
  XNOR U7921 ( .A(n6590), .B(n6589), .Z(n6592) );
  XNOR U7922 ( .A(n6591), .B(n6592), .Z(n6596) );
  XOR U7923 ( .A(n6595), .B(sreg[1337]), .Z(n6588) );
  XNOR U7924 ( .A(n6596), .B(n6588), .Z(c[1337]) );
  NAND U7925 ( .A(n6590), .B(n6589), .Z(n6594) );
  NANDN U7926 ( .A(n6592), .B(n6591), .Z(n6593) );
  NAND U7927 ( .A(n6594), .B(n6593), .Z(n6601) );
  ANDN U7928 ( .B(a[316]), .A(n3937), .Z(n6599) );
  AND U7929 ( .A(b[1]), .B(a[315]), .Z(n6598) );
  XOR U7930 ( .A(n6599), .B(n6598), .Z(n6600) );
  XNOR U7931 ( .A(n6601), .B(n6600), .Z(n6603) );
  XOR U7932 ( .A(sreg[1338]), .B(n6602), .Z(n6597) );
  XNOR U7933 ( .A(n6603), .B(n6597), .Z(c[1338]) );
  NAND U7934 ( .A(b[0]), .B(a[317]), .Z(n6606) );
  NAND U7935 ( .A(a[316]), .B(b[1]), .Z(n6605) );
  XNOR U7936 ( .A(n6606), .B(n6605), .Z(n6608) );
  XNOR U7937 ( .A(n6607), .B(n6608), .Z(n6612) );
  XOR U7938 ( .A(n6611), .B(sreg[1339]), .Z(n6604) );
  XNOR U7939 ( .A(n6612), .B(n6604), .Z(c[1339]) );
  NAND U7940 ( .A(n6606), .B(n6605), .Z(n6610) );
  NANDN U7941 ( .A(n6608), .B(n6607), .Z(n6609) );
  NAND U7942 ( .A(n6610), .B(n6609), .Z(n6617) );
  ANDN U7943 ( .B(a[318]), .A(n3937), .Z(n6615) );
  AND U7944 ( .A(b[1]), .B(a[317]), .Z(n6614) );
  XOR U7945 ( .A(n6615), .B(n6614), .Z(n6616) );
  XNOR U7946 ( .A(n6617), .B(n6616), .Z(n6619) );
  XOR U7947 ( .A(sreg[1340]), .B(n6618), .Z(n6613) );
  XNOR U7948 ( .A(n6619), .B(n6613), .Z(c[1340]) );
  NAND U7949 ( .A(b[0]), .B(a[319]), .Z(n6622) );
  NAND U7950 ( .A(a[318]), .B(b[1]), .Z(n6621) );
  XNOR U7951 ( .A(n6622), .B(n6621), .Z(n6624) );
  XNOR U7952 ( .A(n6623), .B(n6624), .Z(n6628) );
  XOR U7953 ( .A(n6627), .B(sreg[1341]), .Z(n6620) );
  XNOR U7954 ( .A(n6628), .B(n6620), .Z(c[1341]) );
  NAND U7955 ( .A(n6622), .B(n6621), .Z(n6626) );
  NANDN U7956 ( .A(n6624), .B(n6623), .Z(n6625) );
  NAND U7957 ( .A(n6626), .B(n6625), .Z(n6633) );
  ANDN U7958 ( .B(a[320]), .A(n3937), .Z(n6631) );
  AND U7959 ( .A(b[1]), .B(a[319]), .Z(n6630) );
  XOR U7960 ( .A(n6631), .B(n6630), .Z(n6632) );
  XNOR U7961 ( .A(n6633), .B(n6632), .Z(n6635) );
  XOR U7962 ( .A(sreg[1342]), .B(n6634), .Z(n6629) );
  XNOR U7963 ( .A(n6635), .B(n6629), .Z(c[1342]) );
  NAND U7964 ( .A(b[0]), .B(a[321]), .Z(n6638) );
  NAND U7965 ( .A(a[320]), .B(b[1]), .Z(n6637) );
  XNOR U7966 ( .A(n6638), .B(n6637), .Z(n6640) );
  XNOR U7967 ( .A(n6639), .B(n6640), .Z(n6644) );
  XOR U7968 ( .A(n6643), .B(sreg[1343]), .Z(n6636) );
  XNOR U7969 ( .A(n6644), .B(n6636), .Z(c[1343]) );
  NAND U7970 ( .A(n6638), .B(n6637), .Z(n6642) );
  NANDN U7971 ( .A(n6640), .B(n6639), .Z(n6641) );
  NAND U7972 ( .A(n6642), .B(n6641), .Z(n6649) );
  ANDN U7973 ( .B(a[322]), .A(n3938), .Z(n6647) );
  AND U7974 ( .A(b[1]), .B(a[321]), .Z(n6646) );
  XOR U7975 ( .A(n6647), .B(n6646), .Z(n6648) );
  XNOR U7976 ( .A(n6649), .B(n6648), .Z(n6654) );
  XOR U7977 ( .A(sreg[1344]), .B(n6653), .Z(n6645) );
  XNOR U7978 ( .A(n6654), .B(n6645), .Z(c[1344]) );
  OR U7979 ( .A(n6647), .B(n6646), .Z(n6652) );
  IV U7980 ( .A(n6648), .Z(n6650) );
  NANDN U7981 ( .A(n6650), .B(n6649), .Z(n6651) );
  NAND U7982 ( .A(n6652), .B(n6651), .Z(n6658) );
  NAND U7983 ( .A(b[0]), .B(a[323]), .Z(n6657) );
  NAND U7984 ( .A(a[322]), .B(b[1]), .Z(n6656) );
  XNOR U7985 ( .A(n6657), .B(n6656), .Z(n6659) );
  XNOR U7986 ( .A(n6658), .B(n6659), .Z(n6663) );
  XOR U7987 ( .A(n6662), .B(sreg[1345]), .Z(n6655) );
  XNOR U7988 ( .A(n6663), .B(n6655), .Z(c[1345]) );
  NAND U7989 ( .A(n6657), .B(n6656), .Z(n6661) );
  NANDN U7990 ( .A(n6659), .B(n6658), .Z(n6660) );
  NAND U7991 ( .A(n6661), .B(n6660), .Z(n6668) );
  ANDN U7992 ( .B(a[324]), .A(n3938), .Z(n6666) );
  AND U7993 ( .A(b[1]), .B(a[323]), .Z(n6665) );
  XOR U7994 ( .A(n6666), .B(n6665), .Z(n6667) );
  XNOR U7995 ( .A(n6668), .B(n6667), .Z(n6670) );
  XOR U7996 ( .A(sreg[1346]), .B(n6669), .Z(n6664) );
  XNOR U7997 ( .A(n6670), .B(n6664), .Z(c[1346]) );
  NAND U7998 ( .A(b[0]), .B(a[325]), .Z(n6673) );
  NAND U7999 ( .A(a[324]), .B(b[1]), .Z(n6672) );
  XNOR U8000 ( .A(n6673), .B(n6672), .Z(n6675) );
  XNOR U8001 ( .A(n6674), .B(n6675), .Z(n6679) );
  XOR U8002 ( .A(n6678), .B(sreg[1347]), .Z(n6671) );
  XNOR U8003 ( .A(n6679), .B(n6671), .Z(c[1347]) );
  NAND U8004 ( .A(n6673), .B(n6672), .Z(n6677) );
  NANDN U8005 ( .A(n6675), .B(n6674), .Z(n6676) );
  NAND U8006 ( .A(n6677), .B(n6676), .Z(n6683) );
  NAND U8007 ( .A(b[0]), .B(a[326]), .Z(n6682) );
  NAND U8008 ( .A(a[325]), .B(b[1]), .Z(n6681) );
  XNOR U8009 ( .A(n6682), .B(n6681), .Z(n6684) );
  XNOR U8010 ( .A(n6683), .B(n6684), .Z(n6688) );
  XOR U8011 ( .A(n6687), .B(sreg[1348]), .Z(n6680) );
  XNOR U8012 ( .A(n6688), .B(n6680), .Z(c[1348]) );
  NAND U8013 ( .A(n6682), .B(n6681), .Z(n6686) );
  NANDN U8014 ( .A(n6684), .B(n6683), .Z(n6685) );
  NAND U8015 ( .A(n6686), .B(n6685), .Z(n6692) );
  NAND U8016 ( .A(b[0]), .B(a[327]), .Z(n6691) );
  NAND U8017 ( .A(a[326]), .B(b[1]), .Z(n6690) );
  XNOR U8018 ( .A(n6691), .B(n6690), .Z(n6693) );
  XNOR U8019 ( .A(n6692), .B(n6693), .Z(n6697) );
  XOR U8020 ( .A(n6696), .B(sreg[1349]), .Z(n6689) );
  XNOR U8021 ( .A(n6697), .B(n6689), .Z(c[1349]) );
  NAND U8022 ( .A(n6691), .B(n6690), .Z(n6695) );
  NANDN U8023 ( .A(n6693), .B(n6692), .Z(n6694) );
  NAND U8024 ( .A(n6695), .B(n6694), .Z(n6702) );
  ANDN U8025 ( .B(a[328]), .A(n3938), .Z(n6700) );
  AND U8026 ( .A(b[1]), .B(a[327]), .Z(n6699) );
  XOR U8027 ( .A(n6700), .B(n6699), .Z(n6701) );
  XNOR U8028 ( .A(n6702), .B(n6701), .Z(n6704) );
  XOR U8029 ( .A(sreg[1350]), .B(n6703), .Z(n6698) );
  XNOR U8030 ( .A(n6704), .B(n6698), .Z(c[1350]) );
  ANDN U8031 ( .B(a[329]), .A(n3938), .Z(n6707) );
  AND U8032 ( .A(b[1]), .B(a[328]), .Z(n6706) );
  XOR U8033 ( .A(n6707), .B(n6706), .Z(n6708) );
  XNOR U8034 ( .A(n6709), .B(n6708), .Z(n6711) );
  XNOR U8035 ( .A(sreg[1351]), .B(n6710), .Z(n6705) );
  XNOR U8036 ( .A(n6711), .B(n6705), .Z(c[1351]) );
  ANDN U8037 ( .B(a[330]), .A(n3938), .Z(n6714) );
  AND U8038 ( .A(b[1]), .B(a[329]), .Z(n6713) );
  XOR U8039 ( .A(n6714), .B(n6713), .Z(n6715) );
  XNOR U8040 ( .A(n6716), .B(n6715), .Z(n6718) );
  XNOR U8041 ( .A(sreg[1352]), .B(n6717), .Z(n6712) );
  XNOR U8042 ( .A(n6718), .B(n6712), .Z(c[1352]) );
  NAND U8043 ( .A(b[0]), .B(a[331]), .Z(n6721) );
  NAND U8044 ( .A(a[330]), .B(b[1]), .Z(n6720) );
  XNOR U8045 ( .A(n6721), .B(n6720), .Z(n6723) );
  XNOR U8046 ( .A(n6722), .B(n6723), .Z(n6727) );
  XOR U8047 ( .A(n6726), .B(sreg[1353]), .Z(n6719) );
  XNOR U8048 ( .A(n6727), .B(n6719), .Z(c[1353]) );
  NAND U8049 ( .A(n6721), .B(n6720), .Z(n6725) );
  NANDN U8050 ( .A(n6723), .B(n6722), .Z(n6724) );
  NAND U8051 ( .A(n6725), .B(n6724), .Z(n6732) );
  ANDN U8052 ( .B(a[332]), .A(n3938), .Z(n6730) );
  AND U8053 ( .A(b[1]), .B(a[331]), .Z(n6729) );
  XOR U8054 ( .A(n6730), .B(n6729), .Z(n6731) );
  XNOR U8055 ( .A(n6732), .B(n6731), .Z(n6734) );
  XOR U8056 ( .A(sreg[1354]), .B(n6733), .Z(n6728) );
  XNOR U8057 ( .A(n6734), .B(n6728), .Z(c[1354]) );
  ANDN U8058 ( .B(a[333]), .A(n3938), .Z(n6737) );
  AND U8059 ( .A(b[1]), .B(a[332]), .Z(n6736) );
  XOR U8060 ( .A(n6737), .B(n6736), .Z(n6738) );
  XNOR U8061 ( .A(n6739), .B(n6738), .Z(n6741) );
  XNOR U8062 ( .A(sreg[1355]), .B(n6740), .Z(n6735) );
  XNOR U8063 ( .A(n6741), .B(n6735), .Z(c[1355]) );
  ANDN U8064 ( .B(a[334]), .A(n3939), .Z(n6744) );
  AND U8065 ( .A(b[1]), .B(a[333]), .Z(n6743) );
  XOR U8066 ( .A(n6744), .B(n6743), .Z(n6745) );
  XNOR U8067 ( .A(n6746), .B(n6745), .Z(n6751) );
  XNOR U8068 ( .A(sreg[1356]), .B(n6750), .Z(n6742) );
  XNOR U8069 ( .A(n6751), .B(n6742), .Z(c[1356]) );
  OR U8070 ( .A(n6744), .B(n6743), .Z(n6749) );
  IV U8071 ( .A(n6745), .Z(n6747) );
  NANDN U8072 ( .A(n6747), .B(n6746), .Z(n6748) );
  NAND U8073 ( .A(n6749), .B(n6748), .Z(n6755) );
  NAND U8074 ( .A(b[0]), .B(a[335]), .Z(n6754) );
  NAND U8075 ( .A(a[334]), .B(b[1]), .Z(n6753) );
  XNOR U8076 ( .A(n6754), .B(n6753), .Z(n6756) );
  XNOR U8077 ( .A(n6755), .B(n6756), .Z(n6760) );
  XOR U8078 ( .A(n6759), .B(sreg[1357]), .Z(n6752) );
  XNOR U8079 ( .A(n6760), .B(n6752), .Z(c[1357]) );
  NAND U8080 ( .A(n6754), .B(n6753), .Z(n6758) );
  NANDN U8081 ( .A(n6756), .B(n6755), .Z(n6757) );
  NAND U8082 ( .A(n6758), .B(n6757), .Z(n6765) );
  ANDN U8083 ( .B(a[336]), .A(n3939), .Z(n6763) );
  AND U8084 ( .A(b[1]), .B(a[335]), .Z(n6762) );
  XOR U8085 ( .A(n6763), .B(n6762), .Z(n6764) );
  XNOR U8086 ( .A(n6765), .B(n6764), .Z(n6767) );
  XOR U8087 ( .A(sreg[1358]), .B(n6766), .Z(n6761) );
  XNOR U8088 ( .A(n6767), .B(n6761), .Z(c[1358]) );
  NAND U8089 ( .A(b[0]), .B(a[337]), .Z(n6770) );
  NAND U8090 ( .A(a[336]), .B(b[1]), .Z(n6769) );
  XNOR U8091 ( .A(n6770), .B(n6769), .Z(n6772) );
  XNOR U8092 ( .A(n6771), .B(n6772), .Z(n6776) );
  XOR U8093 ( .A(n6775), .B(sreg[1359]), .Z(n6768) );
  XNOR U8094 ( .A(n6776), .B(n6768), .Z(c[1359]) );
  NAND U8095 ( .A(n6770), .B(n6769), .Z(n6774) );
  NANDN U8096 ( .A(n6772), .B(n6771), .Z(n6773) );
  NAND U8097 ( .A(n6774), .B(n6773), .Z(n6781) );
  ANDN U8098 ( .B(a[338]), .A(n3939), .Z(n6779) );
  AND U8099 ( .A(b[1]), .B(a[337]), .Z(n6778) );
  XOR U8100 ( .A(n6779), .B(n6778), .Z(n6780) );
  XNOR U8101 ( .A(n6781), .B(n6780), .Z(n6783) );
  XOR U8102 ( .A(sreg[1360]), .B(n6782), .Z(n6777) );
  XNOR U8103 ( .A(n6783), .B(n6777), .Z(c[1360]) );
  NAND U8104 ( .A(b[0]), .B(a[339]), .Z(n6786) );
  NAND U8105 ( .A(a[338]), .B(b[1]), .Z(n6785) );
  XNOR U8106 ( .A(n6786), .B(n6785), .Z(n6788) );
  XNOR U8107 ( .A(n6787), .B(n6788), .Z(n6792) );
  XOR U8108 ( .A(n6791), .B(sreg[1361]), .Z(n6784) );
  XNOR U8109 ( .A(n6792), .B(n6784), .Z(c[1361]) );
  NAND U8110 ( .A(n6786), .B(n6785), .Z(n6790) );
  NANDN U8111 ( .A(n6788), .B(n6787), .Z(n6789) );
  NAND U8112 ( .A(n6790), .B(n6789), .Z(n6796) );
  NAND U8113 ( .A(b[0]), .B(a[340]), .Z(n6795) );
  NAND U8114 ( .A(a[339]), .B(b[1]), .Z(n6794) );
  XNOR U8115 ( .A(n6795), .B(n6794), .Z(n6797) );
  XNOR U8116 ( .A(n6796), .B(n6797), .Z(n6801) );
  XOR U8117 ( .A(n6800), .B(sreg[1362]), .Z(n6793) );
  XNOR U8118 ( .A(n6801), .B(n6793), .Z(c[1362]) );
  NAND U8119 ( .A(n6795), .B(n6794), .Z(n6799) );
  NANDN U8120 ( .A(n6797), .B(n6796), .Z(n6798) );
  NAND U8121 ( .A(n6799), .B(n6798), .Z(n6805) );
  NAND U8122 ( .A(b[0]), .B(a[341]), .Z(n6804) );
  NAND U8123 ( .A(a[340]), .B(b[1]), .Z(n6803) );
  XNOR U8124 ( .A(n6804), .B(n6803), .Z(n6806) );
  XNOR U8125 ( .A(n6805), .B(n6806), .Z(n6810) );
  XOR U8126 ( .A(n6809), .B(sreg[1363]), .Z(n6802) );
  XNOR U8127 ( .A(n6810), .B(n6802), .Z(c[1363]) );
  NAND U8128 ( .A(n6804), .B(n6803), .Z(n6808) );
  NANDN U8129 ( .A(n6806), .B(n6805), .Z(n6807) );
  NAND U8130 ( .A(n6808), .B(n6807), .Z(n6815) );
  ANDN U8131 ( .B(a[342]), .A(n3939), .Z(n6813) );
  AND U8132 ( .A(b[1]), .B(a[341]), .Z(n6812) );
  XOR U8133 ( .A(n6813), .B(n6812), .Z(n6814) );
  XNOR U8134 ( .A(n6815), .B(n6814), .Z(n6817) );
  XOR U8135 ( .A(sreg[1364]), .B(n6816), .Z(n6811) );
  XNOR U8136 ( .A(n6817), .B(n6811), .Z(c[1364]) );
  NAND U8137 ( .A(b[0]), .B(a[343]), .Z(n6820) );
  NAND U8138 ( .A(a[342]), .B(b[1]), .Z(n6819) );
  XNOR U8139 ( .A(n6820), .B(n6819), .Z(n6822) );
  XNOR U8140 ( .A(n6821), .B(n6822), .Z(n6826) );
  XOR U8141 ( .A(n6825), .B(sreg[1365]), .Z(n6818) );
  XNOR U8142 ( .A(n6826), .B(n6818), .Z(c[1365]) );
  NAND U8143 ( .A(n6820), .B(n6819), .Z(n6824) );
  NANDN U8144 ( .A(n6822), .B(n6821), .Z(n6823) );
  NAND U8145 ( .A(n6824), .B(n6823), .Z(n6830) );
  NAND U8146 ( .A(b[0]), .B(a[344]), .Z(n6829) );
  NAND U8147 ( .A(a[343]), .B(b[1]), .Z(n6828) );
  XNOR U8148 ( .A(n6829), .B(n6828), .Z(n6831) );
  XNOR U8149 ( .A(n6830), .B(n6831), .Z(n6835) );
  XOR U8150 ( .A(n6834), .B(sreg[1366]), .Z(n6827) );
  XNOR U8151 ( .A(n6835), .B(n6827), .Z(c[1366]) );
  NAND U8152 ( .A(n6829), .B(n6828), .Z(n6833) );
  NANDN U8153 ( .A(n6831), .B(n6830), .Z(n6832) );
  NAND U8154 ( .A(n6833), .B(n6832), .Z(n6839) );
  NAND U8155 ( .A(b[0]), .B(a[345]), .Z(n6838) );
  NAND U8156 ( .A(a[344]), .B(b[1]), .Z(n6837) );
  XNOR U8157 ( .A(n6838), .B(n6837), .Z(n6840) );
  XNOR U8158 ( .A(n6839), .B(n6840), .Z(n6844) );
  XOR U8159 ( .A(n6843), .B(sreg[1367]), .Z(n6836) );
  XNOR U8160 ( .A(n6844), .B(n6836), .Z(c[1367]) );
  NAND U8161 ( .A(n6838), .B(n6837), .Z(n6842) );
  NANDN U8162 ( .A(n6840), .B(n6839), .Z(n6841) );
  NAND U8163 ( .A(n6842), .B(n6841), .Z(n6849) );
  ANDN U8164 ( .B(a[346]), .A(n3939), .Z(n6847) );
  AND U8165 ( .A(b[1]), .B(a[345]), .Z(n6846) );
  XOR U8166 ( .A(n6847), .B(n6846), .Z(n6848) );
  XNOR U8167 ( .A(n6849), .B(n6848), .Z(n6851) );
  XOR U8168 ( .A(sreg[1368]), .B(n6850), .Z(n6845) );
  XNOR U8169 ( .A(n6851), .B(n6845), .Z(c[1368]) );
  NAND U8170 ( .A(b[0]), .B(a[347]), .Z(n6854) );
  NAND U8171 ( .A(a[346]), .B(b[1]), .Z(n6853) );
  XNOR U8172 ( .A(n6854), .B(n6853), .Z(n6856) );
  XNOR U8173 ( .A(n6855), .B(n6856), .Z(n6860) );
  XOR U8174 ( .A(n6859), .B(sreg[1369]), .Z(n6852) );
  XNOR U8175 ( .A(n6860), .B(n6852), .Z(c[1369]) );
  NAND U8176 ( .A(n6854), .B(n6853), .Z(n6858) );
  NANDN U8177 ( .A(n6856), .B(n6855), .Z(n6857) );
  NAND U8178 ( .A(n6858), .B(n6857), .Z(n6865) );
  ANDN U8179 ( .B(a[348]), .A(n3939), .Z(n6863) );
  AND U8180 ( .A(b[1]), .B(a[347]), .Z(n6862) );
  XOR U8181 ( .A(n6863), .B(n6862), .Z(n6864) );
  XNOR U8182 ( .A(n6865), .B(n6864), .Z(n6867) );
  XOR U8183 ( .A(sreg[1370]), .B(n6866), .Z(n6861) );
  XNOR U8184 ( .A(n6867), .B(n6861), .Z(c[1370]) );
  NAND U8185 ( .A(b[0]), .B(a[349]), .Z(n6870) );
  NAND U8186 ( .A(a[348]), .B(b[1]), .Z(n6869) );
  XNOR U8187 ( .A(n6870), .B(n6869), .Z(n6872) );
  XNOR U8188 ( .A(n6871), .B(n6872), .Z(n6876) );
  XOR U8189 ( .A(n6875), .B(sreg[1371]), .Z(n6868) );
  XNOR U8190 ( .A(n6876), .B(n6868), .Z(c[1371]) );
  NAND U8191 ( .A(n6870), .B(n6869), .Z(n6874) );
  NANDN U8192 ( .A(n6872), .B(n6871), .Z(n6873) );
  NAND U8193 ( .A(n6874), .B(n6873), .Z(n6880) );
  NAND U8194 ( .A(b[0]), .B(a[350]), .Z(n6879) );
  NAND U8195 ( .A(a[349]), .B(b[1]), .Z(n6878) );
  XNOR U8196 ( .A(n6879), .B(n6878), .Z(n6881) );
  XNOR U8197 ( .A(n6880), .B(n6881), .Z(n6885) );
  XOR U8198 ( .A(n6884), .B(sreg[1372]), .Z(n6877) );
  XNOR U8199 ( .A(n6885), .B(n6877), .Z(c[1372]) );
  NAND U8200 ( .A(n6879), .B(n6878), .Z(n6883) );
  NANDN U8201 ( .A(n6881), .B(n6880), .Z(n6882) );
  NAND U8202 ( .A(n6883), .B(n6882), .Z(n6889) );
  NAND U8203 ( .A(b[0]), .B(a[351]), .Z(n6888) );
  NAND U8204 ( .A(a[350]), .B(b[1]), .Z(n6887) );
  XNOR U8205 ( .A(n6888), .B(n6887), .Z(n6890) );
  XNOR U8206 ( .A(n6889), .B(n6890), .Z(n6894) );
  XOR U8207 ( .A(n6893), .B(sreg[1373]), .Z(n6886) );
  XNOR U8208 ( .A(n6894), .B(n6886), .Z(c[1373]) );
  NAND U8209 ( .A(n6888), .B(n6887), .Z(n6892) );
  NANDN U8210 ( .A(n6890), .B(n6889), .Z(n6891) );
  NAND U8211 ( .A(n6892), .B(n6891), .Z(n6899) );
  ANDN U8212 ( .B(a[352]), .A(n3939), .Z(n6897) );
  AND U8213 ( .A(b[1]), .B(a[351]), .Z(n6896) );
  XOR U8214 ( .A(n6897), .B(n6896), .Z(n6898) );
  XNOR U8215 ( .A(n6899), .B(n6898), .Z(n6901) );
  XOR U8216 ( .A(sreg[1374]), .B(n6900), .Z(n6895) );
  XNOR U8217 ( .A(n6901), .B(n6895), .Z(c[1374]) );
  NAND U8218 ( .A(b[0]), .B(a[353]), .Z(n6904) );
  NAND U8219 ( .A(a[352]), .B(b[1]), .Z(n6903) );
  XNOR U8220 ( .A(n6904), .B(n6903), .Z(n6906) );
  XNOR U8221 ( .A(n6905), .B(n6906), .Z(n6910) );
  XOR U8222 ( .A(n6909), .B(sreg[1375]), .Z(n6902) );
  XNOR U8223 ( .A(n6910), .B(n6902), .Z(c[1375]) );
  NAND U8224 ( .A(n6904), .B(n6903), .Z(n6908) );
  NANDN U8225 ( .A(n6906), .B(n6905), .Z(n6907) );
  NAND U8226 ( .A(n6908), .B(n6907), .Z(n6915) );
  ANDN U8227 ( .B(a[354]), .A(n3940), .Z(n6913) );
  AND U8228 ( .A(b[1]), .B(a[353]), .Z(n6912) );
  XOR U8229 ( .A(n6913), .B(n6912), .Z(n6914) );
  XNOR U8230 ( .A(n6915), .B(n6914), .Z(n6920) );
  XOR U8231 ( .A(sreg[1376]), .B(n6919), .Z(n6911) );
  XNOR U8232 ( .A(n6920), .B(n6911), .Z(c[1376]) );
  OR U8233 ( .A(n6913), .B(n6912), .Z(n6918) );
  IV U8234 ( .A(n6914), .Z(n6916) );
  NANDN U8235 ( .A(n6916), .B(n6915), .Z(n6917) );
  NAND U8236 ( .A(n6918), .B(n6917), .Z(n6924) );
  NAND U8237 ( .A(b[0]), .B(a[355]), .Z(n6923) );
  NAND U8238 ( .A(a[354]), .B(b[1]), .Z(n6922) );
  XNOR U8239 ( .A(n6923), .B(n6922), .Z(n6925) );
  XNOR U8240 ( .A(n6924), .B(n6925), .Z(n6929) );
  XOR U8241 ( .A(n6928), .B(sreg[1377]), .Z(n6921) );
  XNOR U8242 ( .A(n6929), .B(n6921), .Z(c[1377]) );
  NAND U8243 ( .A(n6923), .B(n6922), .Z(n6927) );
  NANDN U8244 ( .A(n6925), .B(n6924), .Z(n6926) );
  NAND U8245 ( .A(n6927), .B(n6926), .Z(n6934) );
  ANDN U8246 ( .B(a[356]), .A(n3940), .Z(n6932) );
  AND U8247 ( .A(b[1]), .B(a[355]), .Z(n6931) );
  XOR U8248 ( .A(n6932), .B(n6931), .Z(n6933) );
  XNOR U8249 ( .A(n6934), .B(n6933), .Z(n6936) );
  XOR U8250 ( .A(sreg[1378]), .B(n6935), .Z(n6930) );
  XNOR U8251 ( .A(n6936), .B(n6930), .Z(c[1378]) );
  NAND U8252 ( .A(b[0]), .B(a[357]), .Z(n6939) );
  NAND U8253 ( .A(a[356]), .B(b[1]), .Z(n6938) );
  XNOR U8254 ( .A(n6939), .B(n6938), .Z(n6941) );
  XNOR U8255 ( .A(n6940), .B(n6941), .Z(n6945) );
  XOR U8256 ( .A(n6944), .B(sreg[1379]), .Z(n6937) );
  XNOR U8257 ( .A(n6945), .B(n6937), .Z(c[1379]) );
  NAND U8258 ( .A(n6939), .B(n6938), .Z(n6943) );
  NANDN U8259 ( .A(n6941), .B(n6940), .Z(n6942) );
  NAND U8260 ( .A(n6943), .B(n6942), .Z(n6950) );
  ANDN U8261 ( .B(a[358]), .A(n3940), .Z(n6948) );
  AND U8262 ( .A(b[1]), .B(a[357]), .Z(n6947) );
  XOR U8263 ( .A(n6948), .B(n6947), .Z(n6949) );
  XNOR U8264 ( .A(n6950), .B(n6949), .Z(n6952) );
  XOR U8265 ( .A(sreg[1380]), .B(n6951), .Z(n6946) );
  XNOR U8266 ( .A(n6952), .B(n6946), .Z(c[1380]) );
  NAND U8267 ( .A(b[0]), .B(a[359]), .Z(n6955) );
  NAND U8268 ( .A(a[358]), .B(b[1]), .Z(n6954) );
  XNOR U8269 ( .A(n6955), .B(n6954), .Z(n6957) );
  XNOR U8270 ( .A(n6956), .B(n6957), .Z(n6961) );
  XOR U8271 ( .A(n6960), .B(sreg[1381]), .Z(n6953) );
  XNOR U8272 ( .A(n6961), .B(n6953), .Z(c[1381]) );
  NAND U8273 ( .A(n6955), .B(n6954), .Z(n6959) );
  NANDN U8274 ( .A(n6957), .B(n6956), .Z(n6958) );
  NAND U8275 ( .A(n6959), .B(n6958), .Z(n6966) );
  ANDN U8276 ( .B(a[360]), .A(n3940), .Z(n6964) );
  AND U8277 ( .A(b[1]), .B(a[359]), .Z(n6963) );
  XOR U8278 ( .A(n6964), .B(n6963), .Z(n6965) );
  XNOR U8279 ( .A(n6966), .B(n6965), .Z(n6968) );
  XOR U8280 ( .A(sreg[1382]), .B(n6967), .Z(n6962) );
  XNOR U8281 ( .A(n6968), .B(n6962), .Z(c[1382]) );
  ANDN U8282 ( .B(a[361]), .A(n3940), .Z(n6971) );
  AND U8283 ( .A(b[1]), .B(a[360]), .Z(n6970) );
  XOR U8284 ( .A(n6971), .B(n6970), .Z(n6972) );
  XNOR U8285 ( .A(n6973), .B(n6972), .Z(n6975) );
  XNOR U8286 ( .A(sreg[1383]), .B(n6974), .Z(n6969) );
  XNOR U8287 ( .A(n6975), .B(n6969), .Z(c[1383]) );
  ANDN U8288 ( .B(a[362]), .A(n3940), .Z(n6978) );
  AND U8289 ( .A(b[1]), .B(a[361]), .Z(n6977) );
  XOR U8290 ( .A(n6978), .B(n6977), .Z(n6979) );
  XNOR U8291 ( .A(n6980), .B(n6979), .Z(n6982) );
  XNOR U8292 ( .A(sreg[1384]), .B(n6981), .Z(n6976) );
  XNOR U8293 ( .A(n6982), .B(n6976), .Z(c[1384]) );
  NAND U8294 ( .A(b[0]), .B(a[363]), .Z(n6985) );
  NAND U8295 ( .A(a[362]), .B(b[1]), .Z(n6984) );
  XNOR U8296 ( .A(n6985), .B(n6984), .Z(n6987) );
  XNOR U8297 ( .A(n6986), .B(n6987), .Z(n6991) );
  XOR U8298 ( .A(n6990), .B(sreg[1385]), .Z(n6983) );
  XNOR U8299 ( .A(n6991), .B(n6983), .Z(c[1385]) );
  NAND U8300 ( .A(n6985), .B(n6984), .Z(n6989) );
  NANDN U8301 ( .A(n6987), .B(n6986), .Z(n6988) );
  NAND U8302 ( .A(n6989), .B(n6988), .Z(n6996) );
  ANDN U8303 ( .B(a[364]), .A(n3940), .Z(n6994) );
  AND U8304 ( .A(b[1]), .B(a[363]), .Z(n6993) );
  XOR U8305 ( .A(n6994), .B(n6993), .Z(n6995) );
  XNOR U8306 ( .A(n6996), .B(n6995), .Z(n6998) );
  XOR U8307 ( .A(sreg[1386]), .B(n6997), .Z(n6992) );
  XNOR U8308 ( .A(n6998), .B(n6992), .Z(c[1386]) );
  ANDN U8309 ( .B(a[365]), .A(n3941), .Z(n7001) );
  AND U8310 ( .A(b[1]), .B(a[364]), .Z(n7000) );
  XOR U8311 ( .A(n7001), .B(n7000), .Z(n7002) );
  XNOR U8312 ( .A(n7003), .B(n7002), .Z(n7008) );
  XNOR U8313 ( .A(sreg[1387]), .B(n7007), .Z(n6999) );
  XNOR U8314 ( .A(n7008), .B(n6999), .Z(c[1387]) );
  OR U8315 ( .A(n7001), .B(n7000), .Z(n7006) );
  IV U8316 ( .A(n7002), .Z(n7004) );
  NANDN U8317 ( .A(n7004), .B(n7003), .Z(n7005) );
  NAND U8318 ( .A(n7006), .B(n7005), .Z(n7013) );
  ANDN U8319 ( .B(a[366]), .A(n3941), .Z(n7011) );
  AND U8320 ( .A(b[1]), .B(a[365]), .Z(n7010) );
  XOR U8321 ( .A(n7011), .B(n7010), .Z(n7012) );
  XNOR U8322 ( .A(n7013), .B(n7012), .Z(n7015) );
  XNOR U8323 ( .A(sreg[1388]), .B(n7014), .Z(n7009) );
  XNOR U8324 ( .A(n7015), .B(n7009), .Z(c[1388]) );
  NAND U8325 ( .A(b[0]), .B(a[367]), .Z(n7018) );
  NAND U8326 ( .A(a[366]), .B(b[1]), .Z(n7017) );
  XNOR U8327 ( .A(n7018), .B(n7017), .Z(n7020) );
  XNOR U8328 ( .A(n7019), .B(n7020), .Z(n7024) );
  XOR U8329 ( .A(n7023), .B(sreg[1389]), .Z(n7016) );
  XNOR U8330 ( .A(n7024), .B(n7016), .Z(c[1389]) );
  NAND U8331 ( .A(n7018), .B(n7017), .Z(n7022) );
  NANDN U8332 ( .A(n7020), .B(n7019), .Z(n7021) );
  NAND U8333 ( .A(n7022), .B(n7021), .Z(n7029) );
  ANDN U8334 ( .B(a[368]), .A(n3941), .Z(n7027) );
  AND U8335 ( .A(b[1]), .B(a[367]), .Z(n7026) );
  XOR U8336 ( .A(n7027), .B(n7026), .Z(n7028) );
  XNOR U8337 ( .A(n7029), .B(n7028), .Z(n7031) );
  XOR U8338 ( .A(sreg[1390]), .B(n7030), .Z(n7025) );
  XNOR U8339 ( .A(n7031), .B(n7025), .Z(c[1390]) );
  NAND U8340 ( .A(b[0]), .B(a[369]), .Z(n7034) );
  NAND U8341 ( .A(a[368]), .B(b[1]), .Z(n7033) );
  XNOR U8342 ( .A(n7034), .B(n7033), .Z(n7036) );
  XNOR U8343 ( .A(n7035), .B(n7036), .Z(n7040) );
  XOR U8344 ( .A(n7039), .B(sreg[1391]), .Z(n7032) );
  XNOR U8345 ( .A(n7040), .B(n7032), .Z(c[1391]) );
  NAND U8346 ( .A(n7034), .B(n7033), .Z(n7038) );
  NANDN U8347 ( .A(n7036), .B(n7035), .Z(n7037) );
  NAND U8348 ( .A(n7038), .B(n7037), .Z(n7045) );
  ANDN U8349 ( .B(a[370]), .A(n3941), .Z(n7043) );
  AND U8350 ( .A(b[1]), .B(a[369]), .Z(n7042) );
  XOR U8351 ( .A(n7043), .B(n7042), .Z(n7044) );
  XNOR U8352 ( .A(n7045), .B(n7044), .Z(n7047) );
  XOR U8353 ( .A(sreg[1392]), .B(n7046), .Z(n7041) );
  XNOR U8354 ( .A(n7047), .B(n7041), .Z(c[1392]) );
  NAND U8355 ( .A(b[0]), .B(a[371]), .Z(n7050) );
  NAND U8356 ( .A(a[370]), .B(b[1]), .Z(n7049) );
  XNOR U8357 ( .A(n7050), .B(n7049), .Z(n7052) );
  XNOR U8358 ( .A(n7051), .B(n7052), .Z(n7056) );
  XOR U8359 ( .A(n7055), .B(sreg[1393]), .Z(n7048) );
  XNOR U8360 ( .A(n7056), .B(n7048), .Z(c[1393]) );
  NAND U8361 ( .A(n7050), .B(n7049), .Z(n7054) );
  NANDN U8362 ( .A(n7052), .B(n7051), .Z(n7053) );
  NAND U8363 ( .A(n7054), .B(n7053), .Z(n7061) );
  ANDN U8364 ( .B(a[372]), .A(n3941), .Z(n7059) );
  AND U8365 ( .A(b[1]), .B(a[371]), .Z(n7058) );
  XOR U8366 ( .A(n7059), .B(n7058), .Z(n7060) );
  XNOR U8367 ( .A(n7061), .B(n7060), .Z(n7063) );
  XOR U8368 ( .A(sreg[1394]), .B(n7062), .Z(n7057) );
  XNOR U8369 ( .A(n7063), .B(n7057), .Z(c[1394]) );
  ANDN U8370 ( .B(a[373]), .A(n3941), .Z(n7066) );
  AND U8371 ( .A(b[1]), .B(a[372]), .Z(n7065) );
  XOR U8372 ( .A(n7066), .B(n7065), .Z(n7067) );
  XNOR U8373 ( .A(n7068), .B(n7067), .Z(n7070) );
  XNOR U8374 ( .A(sreg[1395]), .B(n7069), .Z(n7064) );
  XNOR U8375 ( .A(n7070), .B(n7064), .Z(c[1395]) );
  ANDN U8376 ( .B(a[374]), .A(n3941), .Z(n7073) );
  AND U8377 ( .A(b[1]), .B(a[373]), .Z(n7072) );
  XOR U8378 ( .A(n7073), .B(n7072), .Z(n7074) );
  XNOR U8379 ( .A(n7075), .B(n7074), .Z(n7077) );
  XNOR U8380 ( .A(sreg[1396]), .B(n7076), .Z(n7071) );
  XNOR U8381 ( .A(n7077), .B(n7071), .Z(c[1396]) );
  NAND U8382 ( .A(b[0]), .B(a[375]), .Z(n7080) );
  NAND U8383 ( .A(a[374]), .B(b[1]), .Z(n7079) );
  XNOR U8384 ( .A(n7080), .B(n7079), .Z(n7082) );
  XNOR U8385 ( .A(n7081), .B(n7082), .Z(n7086) );
  XOR U8386 ( .A(n7085), .B(sreg[1397]), .Z(n7078) );
  XNOR U8387 ( .A(n7086), .B(n7078), .Z(c[1397]) );
  NAND U8388 ( .A(n7080), .B(n7079), .Z(n7084) );
  NANDN U8389 ( .A(n7082), .B(n7081), .Z(n7083) );
  NAND U8390 ( .A(n7084), .B(n7083), .Z(n7091) );
  ANDN U8391 ( .B(a[376]), .A(n3942), .Z(n7089) );
  AND U8392 ( .A(b[1]), .B(a[375]), .Z(n7088) );
  XOR U8393 ( .A(n7089), .B(n7088), .Z(n7090) );
  XNOR U8394 ( .A(n7091), .B(n7090), .Z(n7096) );
  XOR U8395 ( .A(sreg[1398]), .B(n7095), .Z(n7087) );
  XNOR U8396 ( .A(n7096), .B(n7087), .Z(c[1398]) );
  OR U8397 ( .A(n7089), .B(n7088), .Z(n7094) );
  IV U8398 ( .A(n7090), .Z(n7092) );
  NANDN U8399 ( .A(n7092), .B(n7091), .Z(n7093) );
  NAND U8400 ( .A(n7094), .B(n7093), .Z(n7100) );
  NAND U8401 ( .A(b[0]), .B(a[377]), .Z(n7099) );
  NAND U8402 ( .A(a[376]), .B(b[1]), .Z(n7098) );
  XNOR U8403 ( .A(n7099), .B(n7098), .Z(n7101) );
  XNOR U8404 ( .A(n7100), .B(n7101), .Z(n7105) );
  XOR U8405 ( .A(n7104), .B(sreg[1399]), .Z(n7097) );
  XNOR U8406 ( .A(n7105), .B(n7097), .Z(c[1399]) );
  NAND U8407 ( .A(n7099), .B(n7098), .Z(n7103) );
  NANDN U8408 ( .A(n7101), .B(n7100), .Z(n7102) );
  NAND U8409 ( .A(n7103), .B(n7102), .Z(n7110) );
  ANDN U8410 ( .B(a[378]), .A(n3942), .Z(n7108) );
  AND U8411 ( .A(b[1]), .B(a[377]), .Z(n7107) );
  XOR U8412 ( .A(n7108), .B(n7107), .Z(n7109) );
  XNOR U8413 ( .A(n7110), .B(n7109), .Z(n7112) );
  XOR U8414 ( .A(sreg[1400]), .B(n7111), .Z(n7106) );
  XNOR U8415 ( .A(n7112), .B(n7106), .Z(c[1400]) );
  ANDN U8416 ( .B(a[379]), .A(n3942), .Z(n7115) );
  AND U8417 ( .A(b[1]), .B(a[378]), .Z(n7114) );
  XOR U8418 ( .A(n7115), .B(n7114), .Z(n7116) );
  XNOR U8419 ( .A(n7117), .B(n7116), .Z(n7119) );
  XNOR U8420 ( .A(sreg[1401]), .B(n7118), .Z(n7113) );
  XNOR U8421 ( .A(n7119), .B(n7113), .Z(c[1401]) );
  ANDN U8422 ( .B(a[380]), .A(n3942), .Z(n7122) );
  AND U8423 ( .A(b[1]), .B(a[379]), .Z(n7121) );
  XOR U8424 ( .A(n7122), .B(n7121), .Z(n7123) );
  XNOR U8425 ( .A(n7124), .B(n7123), .Z(n7126) );
  XNOR U8426 ( .A(sreg[1402]), .B(n7125), .Z(n7120) );
  XNOR U8427 ( .A(n7126), .B(n7120), .Z(c[1402]) );
  NAND U8428 ( .A(b[0]), .B(a[381]), .Z(n7129) );
  NAND U8429 ( .A(a[380]), .B(b[1]), .Z(n7128) );
  XNOR U8430 ( .A(n7129), .B(n7128), .Z(n7131) );
  XNOR U8431 ( .A(n7130), .B(n7131), .Z(n7135) );
  XOR U8432 ( .A(n7134), .B(sreg[1403]), .Z(n7127) );
  XNOR U8433 ( .A(n7135), .B(n7127), .Z(c[1403]) );
  NAND U8434 ( .A(n7129), .B(n7128), .Z(n7133) );
  NANDN U8435 ( .A(n7131), .B(n7130), .Z(n7132) );
  NAND U8436 ( .A(n7133), .B(n7132), .Z(n7140) );
  ANDN U8437 ( .B(a[382]), .A(n3942), .Z(n7138) );
  AND U8438 ( .A(b[1]), .B(a[381]), .Z(n7137) );
  XOR U8439 ( .A(n7138), .B(n7137), .Z(n7139) );
  XNOR U8440 ( .A(n7140), .B(n7139), .Z(n7142) );
  XOR U8441 ( .A(sreg[1404]), .B(n7141), .Z(n7136) );
  XNOR U8442 ( .A(n7142), .B(n7136), .Z(c[1404]) );
  NAND U8443 ( .A(b[0]), .B(a[383]), .Z(n7145) );
  NAND U8444 ( .A(a[382]), .B(b[1]), .Z(n7144) );
  XNOR U8445 ( .A(n7145), .B(n7144), .Z(n7147) );
  XNOR U8446 ( .A(n7146), .B(n7147), .Z(n7151) );
  XOR U8447 ( .A(n7150), .B(sreg[1405]), .Z(n7143) );
  XNOR U8448 ( .A(n7151), .B(n7143), .Z(c[1405]) );
  NAND U8449 ( .A(n7145), .B(n7144), .Z(n7149) );
  NANDN U8450 ( .A(n7147), .B(n7146), .Z(n7148) );
  NAND U8451 ( .A(n7149), .B(n7148), .Z(n7156) );
  ANDN U8452 ( .B(a[384]), .A(n3942), .Z(n7154) );
  AND U8453 ( .A(b[1]), .B(a[383]), .Z(n7153) );
  XOR U8454 ( .A(n7154), .B(n7153), .Z(n7155) );
  XNOR U8455 ( .A(n7156), .B(n7155), .Z(n7158) );
  XOR U8456 ( .A(sreg[1406]), .B(n7157), .Z(n7152) );
  XNOR U8457 ( .A(n7158), .B(n7152), .Z(c[1406]) );
  NAND U8458 ( .A(b[0]), .B(a[385]), .Z(n7161) );
  NAND U8459 ( .A(a[384]), .B(b[1]), .Z(n7160) );
  XNOR U8460 ( .A(n7161), .B(n7160), .Z(n7163) );
  XNOR U8461 ( .A(n7162), .B(n7163), .Z(n7167) );
  XOR U8462 ( .A(n7166), .B(sreg[1407]), .Z(n7159) );
  XNOR U8463 ( .A(n7167), .B(n7159), .Z(c[1407]) );
  NAND U8464 ( .A(n7161), .B(n7160), .Z(n7165) );
  NANDN U8465 ( .A(n7163), .B(n7162), .Z(n7164) );
  NAND U8466 ( .A(n7165), .B(n7164), .Z(n7172) );
  ANDN U8467 ( .B(a[386]), .A(n3942), .Z(n7170) );
  AND U8468 ( .A(b[1]), .B(a[385]), .Z(n7169) );
  XOR U8469 ( .A(n7170), .B(n7169), .Z(n7171) );
  XNOR U8470 ( .A(n7172), .B(n7171), .Z(n7174) );
  XOR U8471 ( .A(sreg[1408]), .B(n7173), .Z(n7168) );
  XNOR U8472 ( .A(n7174), .B(n7168), .Z(c[1408]) );
  NAND U8473 ( .A(b[0]), .B(a[387]), .Z(n7177) );
  NAND U8474 ( .A(a[386]), .B(b[1]), .Z(n7176) );
  XNOR U8475 ( .A(n7177), .B(n7176), .Z(n7179) );
  XNOR U8476 ( .A(n7178), .B(n7179), .Z(n7183) );
  XOR U8477 ( .A(n7182), .B(sreg[1409]), .Z(n7175) );
  XNOR U8478 ( .A(n7183), .B(n7175), .Z(c[1409]) );
  NAND U8479 ( .A(n7177), .B(n7176), .Z(n7181) );
  NANDN U8480 ( .A(n7179), .B(n7178), .Z(n7180) );
  NAND U8481 ( .A(n7181), .B(n7180), .Z(n7188) );
  ANDN U8482 ( .B(a[388]), .A(n3943), .Z(n7186) );
  AND U8483 ( .A(b[1]), .B(a[387]), .Z(n7185) );
  XOR U8484 ( .A(n7186), .B(n7185), .Z(n7187) );
  XNOR U8485 ( .A(n7188), .B(n7187), .Z(n7193) );
  XOR U8486 ( .A(sreg[1410]), .B(n7192), .Z(n7184) );
  XNOR U8487 ( .A(n7193), .B(n7184), .Z(c[1410]) );
  OR U8488 ( .A(n7186), .B(n7185), .Z(n7191) );
  IV U8489 ( .A(n7187), .Z(n7189) );
  NANDN U8490 ( .A(n7189), .B(n7188), .Z(n7190) );
  NAND U8491 ( .A(n7191), .B(n7190), .Z(n7197) );
  NAND U8492 ( .A(b[0]), .B(a[389]), .Z(n7196) );
  NAND U8493 ( .A(a[388]), .B(b[1]), .Z(n7195) );
  XNOR U8494 ( .A(n7196), .B(n7195), .Z(n7198) );
  XNOR U8495 ( .A(n7197), .B(n7198), .Z(n7202) );
  XOR U8496 ( .A(n7201), .B(sreg[1411]), .Z(n7194) );
  XNOR U8497 ( .A(n7202), .B(n7194), .Z(c[1411]) );
  NAND U8498 ( .A(n7196), .B(n7195), .Z(n7200) );
  NANDN U8499 ( .A(n7198), .B(n7197), .Z(n7199) );
  NAND U8500 ( .A(n7200), .B(n7199), .Z(n7207) );
  ANDN U8501 ( .B(a[390]), .A(n3943), .Z(n7205) );
  AND U8502 ( .A(b[1]), .B(a[389]), .Z(n7204) );
  XOR U8503 ( .A(n7205), .B(n7204), .Z(n7206) );
  XNOR U8504 ( .A(n7207), .B(n7206), .Z(n7209) );
  XOR U8505 ( .A(sreg[1412]), .B(n7208), .Z(n7203) );
  XNOR U8506 ( .A(n7209), .B(n7203), .Z(c[1412]) );
  NAND U8507 ( .A(b[0]), .B(a[391]), .Z(n7212) );
  NAND U8508 ( .A(a[390]), .B(b[1]), .Z(n7211) );
  XNOR U8509 ( .A(n7212), .B(n7211), .Z(n7214) );
  XNOR U8510 ( .A(n7213), .B(n7214), .Z(n7218) );
  XOR U8511 ( .A(n7217), .B(sreg[1413]), .Z(n7210) );
  XNOR U8512 ( .A(n7218), .B(n7210), .Z(c[1413]) );
  NAND U8513 ( .A(n7212), .B(n7211), .Z(n7216) );
  NANDN U8514 ( .A(n7214), .B(n7213), .Z(n7215) );
  NAND U8515 ( .A(n7216), .B(n7215), .Z(n7223) );
  ANDN U8516 ( .B(a[392]), .A(n3943), .Z(n7221) );
  AND U8517 ( .A(b[1]), .B(a[391]), .Z(n7220) );
  XOR U8518 ( .A(n7221), .B(n7220), .Z(n7222) );
  XNOR U8519 ( .A(n7223), .B(n7222), .Z(n7225) );
  XOR U8520 ( .A(sreg[1414]), .B(n7224), .Z(n7219) );
  XNOR U8521 ( .A(n7225), .B(n7219), .Z(c[1414]) );
  NAND U8522 ( .A(b[0]), .B(a[393]), .Z(n7228) );
  NAND U8523 ( .A(a[392]), .B(b[1]), .Z(n7227) );
  XNOR U8524 ( .A(n7228), .B(n7227), .Z(n7230) );
  XNOR U8525 ( .A(n7229), .B(n7230), .Z(n7234) );
  XOR U8526 ( .A(n7233), .B(sreg[1415]), .Z(n7226) );
  XNOR U8527 ( .A(n7234), .B(n7226), .Z(c[1415]) );
  NAND U8528 ( .A(n7228), .B(n7227), .Z(n7232) );
  NANDN U8529 ( .A(n7230), .B(n7229), .Z(n7231) );
  NAND U8530 ( .A(n7232), .B(n7231), .Z(n7239) );
  ANDN U8531 ( .B(a[394]), .A(n3943), .Z(n7237) );
  AND U8532 ( .A(b[1]), .B(a[393]), .Z(n7236) );
  XOR U8533 ( .A(n7237), .B(n7236), .Z(n7238) );
  XNOR U8534 ( .A(n7239), .B(n7238), .Z(n7241) );
  XOR U8535 ( .A(sreg[1416]), .B(n7240), .Z(n7235) );
  XNOR U8536 ( .A(n7241), .B(n7235), .Z(c[1416]) );
  NAND U8537 ( .A(b[0]), .B(a[395]), .Z(n7244) );
  NAND U8538 ( .A(a[394]), .B(b[1]), .Z(n7243) );
  XNOR U8539 ( .A(n7244), .B(n7243), .Z(n7246) );
  XNOR U8540 ( .A(n7245), .B(n7246), .Z(n7250) );
  XOR U8541 ( .A(n7249), .B(sreg[1417]), .Z(n7242) );
  XNOR U8542 ( .A(n7250), .B(n7242), .Z(c[1417]) );
  NAND U8543 ( .A(n7244), .B(n7243), .Z(n7248) );
  NANDN U8544 ( .A(n7246), .B(n7245), .Z(n7247) );
  NAND U8545 ( .A(n7248), .B(n7247), .Z(n7255) );
  ANDN U8546 ( .B(a[396]), .A(n3943), .Z(n7253) );
  AND U8547 ( .A(b[1]), .B(a[395]), .Z(n7252) );
  XOR U8548 ( .A(n7253), .B(n7252), .Z(n7254) );
  XNOR U8549 ( .A(n7255), .B(n7254), .Z(n7257) );
  XOR U8550 ( .A(sreg[1418]), .B(n7256), .Z(n7251) );
  XNOR U8551 ( .A(n7257), .B(n7251), .Z(c[1418]) );
  NAND U8552 ( .A(b[0]), .B(a[397]), .Z(n7260) );
  NAND U8553 ( .A(a[396]), .B(b[1]), .Z(n7259) );
  XNOR U8554 ( .A(n7260), .B(n7259), .Z(n7262) );
  XNOR U8555 ( .A(n7261), .B(n7262), .Z(n7266) );
  XOR U8556 ( .A(n7265), .B(sreg[1419]), .Z(n7258) );
  XNOR U8557 ( .A(n7266), .B(n7258), .Z(c[1419]) );
  NAND U8558 ( .A(n7260), .B(n7259), .Z(n7264) );
  NANDN U8559 ( .A(n7262), .B(n7261), .Z(n7263) );
  NAND U8560 ( .A(n7264), .B(n7263), .Z(n7271) );
  ANDN U8561 ( .B(a[398]), .A(n3943), .Z(n7269) );
  AND U8562 ( .A(b[1]), .B(a[397]), .Z(n7268) );
  XOR U8563 ( .A(n7269), .B(n7268), .Z(n7270) );
  XNOR U8564 ( .A(n7271), .B(n7270), .Z(n7273) );
  XOR U8565 ( .A(sreg[1420]), .B(n7272), .Z(n7267) );
  XNOR U8566 ( .A(n7273), .B(n7267), .Z(c[1420]) );
  NAND U8567 ( .A(b[0]), .B(a[399]), .Z(n7276) );
  NAND U8568 ( .A(a[398]), .B(b[1]), .Z(n7275) );
  XNOR U8569 ( .A(n7276), .B(n7275), .Z(n7278) );
  XNOR U8570 ( .A(n7277), .B(n7278), .Z(n7282) );
  XOR U8571 ( .A(n7281), .B(sreg[1421]), .Z(n7274) );
  XNOR U8572 ( .A(n7282), .B(n7274), .Z(c[1421]) );
  NAND U8573 ( .A(n7276), .B(n7275), .Z(n7280) );
  NANDN U8574 ( .A(n7278), .B(n7277), .Z(n7279) );
  NAND U8575 ( .A(n7280), .B(n7279), .Z(n7287) );
  ANDN U8576 ( .B(a[400]), .A(n3943), .Z(n7285) );
  AND U8577 ( .A(b[1]), .B(a[399]), .Z(n7284) );
  XOR U8578 ( .A(n7285), .B(n7284), .Z(n7286) );
  XNOR U8579 ( .A(n7287), .B(n7286), .Z(n7289) );
  XOR U8580 ( .A(sreg[1422]), .B(n7288), .Z(n7283) );
  XNOR U8581 ( .A(n7289), .B(n7283), .Z(c[1422]) );
  NAND U8582 ( .A(b[0]), .B(a[401]), .Z(n7292) );
  NAND U8583 ( .A(a[400]), .B(b[1]), .Z(n7291) );
  XNOR U8584 ( .A(n7292), .B(n7291), .Z(n7294) );
  XNOR U8585 ( .A(n7293), .B(n7294), .Z(n7298) );
  XOR U8586 ( .A(n7297), .B(sreg[1423]), .Z(n7290) );
  XNOR U8587 ( .A(n7298), .B(n7290), .Z(c[1423]) );
  NAND U8588 ( .A(n7292), .B(n7291), .Z(n7296) );
  NANDN U8589 ( .A(n7294), .B(n7293), .Z(n7295) );
  NAND U8590 ( .A(n7296), .B(n7295), .Z(n7303) );
  ANDN U8591 ( .B(a[402]), .A(n3944), .Z(n7301) );
  AND U8592 ( .A(b[1]), .B(a[401]), .Z(n7300) );
  XOR U8593 ( .A(n7301), .B(n7300), .Z(n7302) );
  XNOR U8594 ( .A(n7303), .B(n7302), .Z(n7308) );
  XOR U8595 ( .A(sreg[1424]), .B(n7307), .Z(n7299) );
  XNOR U8596 ( .A(n7308), .B(n7299), .Z(c[1424]) );
  OR U8597 ( .A(n7301), .B(n7300), .Z(n7306) );
  IV U8598 ( .A(n7302), .Z(n7304) );
  NANDN U8599 ( .A(n7304), .B(n7303), .Z(n7305) );
  NAND U8600 ( .A(n7306), .B(n7305), .Z(n7312) );
  NAND U8601 ( .A(b[0]), .B(a[403]), .Z(n7311) );
  NAND U8602 ( .A(a[402]), .B(b[1]), .Z(n7310) );
  XNOR U8603 ( .A(n7311), .B(n7310), .Z(n7313) );
  XNOR U8604 ( .A(n7312), .B(n7313), .Z(n7317) );
  XOR U8605 ( .A(n7316), .B(sreg[1425]), .Z(n7309) );
  XNOR U8606 ( .A(n7317), .B(n7309), .Z(c[1425]) );
  NAND U8607 ( .A(n7311), .B(n7310), .Z(n7315) );
  NANDN U8608 ( .A(n7313), .B(n7312), .Z(n7314) );
  NAND U8609 ( .A(n7315), .B(n7314), .Z(n7322) );
  ANDN U8610 ( .B(a[404]), .A(n3944), .Z(n7320) );
  AND U8611 ( .A(b[1]), .B(a[403]), .Z(n7319) );
  XOR U8612 ( .A(n7320), .B(n7319), .Z(n7321) );
  XNOR U8613 ( .A(n7322), .B(n7321), .Z(n7324) );
  XOR U8614 ( .A(sreg[1426]), .B(n7323), .Z(n7318) );
  XNOR U8615 ( .A(n7324), .B(n7318), .Z(c[1426]) );
  NAND U8616 ( .A(b[0]), .B(a[405]), .Z(n7327) );
  NAND U8617 ( .A(a[404]), .B(b[1]), .Z(n7326) );
  XNOR U8618 ( .A(n7327), .B(n7326), .Z(n7329) );
  XNOR U8619 ( .A(n7328), .B(n7329), .Z(n7333) );
  XOR U8620 ( .A(n7332), .B(sreg[1427]), .Z(n7325) );
  XNOR U8621 ( .A(n7333), .B(n7325), .Z(c[1427]) );
  NAND U8622 ( .A(n7327), .B(n7326), .Z(n7331) );
  NANDN U8623 ( .A(n7329), .B(n7328), .Z(n7330) );
  NAND U8624 ( .A(n7331), .B(n7330), .Z(n7337) );
  NAND U8625 ( .A(b[0]), .B(a[406]), .Z(n7336) );
  NAND U8626 ( .A(a[405]), .B(b[1]), .Z(n7335) );
  XNOR U8627 ( .A(n7336), .B(n7335), .Z(n7338) );
  XNOR U8628 ( .A(n7337), .B(n7338), .Z(n7342) );
  XOR U8629 ( .A(n7341), .B(sreg[1428]), .Z(n7334) );
  XNOR U8630 ( .A(n7342), .B(n7334), .Z(c[1428]) );
  NAND U8631 ( .A(n7336), .B(n7335), .Z(n7340) );
  NANDN U8632 ( .A(n7338), .B(n7337), .Z(n7339) );
  NAND U8633 ( .A(n7340), .B(n7339), .Z(n7346) );
  NAND U8634 ( .A(b[0]), .B(a[407]), .Z(n7345) );
  NAND U8635 ( .A(a[406]), .B(b[1]), .Z(n7344) );
  XNOR U8636 ( .A(n7345), .B(n7344), .Z(n7347) );
  XNOR U8637 ( .A(n7346), .B(n7347), .Z(n7351) );
  XOR U8638 ( .A(n7350), .B(sreg[1429]), .Z(n7343) );
  XNOR U8639 ( .A(n7351), .B(n7343), .Z(c[1429]) );
  NAND U8640 ( .A(n7345), .B(n7344), .Z(n7349) );
  NANDN U8641 ( .A(n7347), .B(n7346), .Z(n7348) );
  NAND U8642 ( .A(n7349), .B(n7348), .Z(n7356) );
  ANDN U8643 ( .B(a[408]), .A(n3944), .Z(n7354) );
  AND U8644 ( .A(b[1]), .B(a[407]), .Z(n7353) );
  XOR U8645 ( .A(n7354), .B(n7353), .Z(n7355) );
  XNOR U8646 ( .A(n7356), .B(n7355), .Z(n7358) );
  XOR U8647 ( .A(sreg[1430]), .B(n7357), .Z(n7352) );
  XNOR U8648 ( .A(n7358), .B(n7352), .Z(c[1430]) );
  NAND U8649 ( .A(b[0]), .B(a[409]), .Z(n7361) );
  NAND U8650 ( .A(a[408]), .B(b[1]), .Z(n7360) );
  XNOR U8651 ( .A(n7361), .B(n7360), .Z(n7363) );
  XNOR U8652 ( .A(n7362), .B(n7363), .Z(n7367) );
  XOR U8653 ( .A(n7366), .B(sreg[1431]), .Z(n7359) );
  XNOR U8654 ( .A(n7367), .B(n7359), .Z(c[1431]) );
  NAND U8655 ( .A(n7361), .B(n7360), .Z(n7365) );
  NANDN U8656 ( .A(n7363), .B(n7362), .Z(n7364) );
  NAND U8657 ( .A(n7365), .B(n7364), .Z(n7372) );
  ANDN U8658 ( .B(a[410]), .A(n3944), .Z(n7370) );
  AND U8659 ( .A(b[1]), .B(a[409]), .Z(n7369) );
  XOR U8660 ( .A(n7370), .B(n7369), .Z(n7371) );
  XNOR U8661 ( .A(n7372), .B(n7371), .Z(n7374) );
  XOR U8662 ( .A(sreg[1432]), .B(n7373), .Z(n7368) );
  XNOR U8663 ( .A(n7374), .B(n7368), .Z(c[1432]) );
  ANDN U8664 ( .B(a[411]), .A(n3944), .Z(n7377) );
  AND U8665 ( .A(b[1]), .B(a[410]), .Z(n7376) );
  XOR U8666 ( .A(n7377), .B(n7376), .Z(n7378) );
  XNOR U8667 ( .A(n7379), .B(n7378), .Z(n7381) );
  XNOR U8668 ( .A(sreg[1433]), .B(n7380), .Z(n7375) );
  XNOR U8669 ( .A(n7381), .B(n7375), .Z(c[1433]) );
  NAND U8670 ( .A(b[0]), .B(a[412]), .Z(n7384) );
  NAND U8671 ( .A(a[411]), .B(b[1]), .Z(n7383) );
  XNOR U8672 ( .A(n7384), .B(n7383), .Z(n7386) );
  XNOR U8673 ( .A(n7385), .B(n7386), .Z(n7390) );
  XOR U8674 ( .A(n7389), .B(sreg[1434]), .Z(n7382) );
  XNOR U8675 ( .A(n7390), .B(n7382), .Z(c[1434]) );
  NAND U8676 ( .A(n7384), .B(n7383), .Z(n7388) );
  NANDN U8677 ( .A(n7386), .B(n7385), .Z(n7387) );
  NAND U8678 ( .A(n7388), .B(n7387), .Z(n7394) );
  NAND U8679 ( .A(b[0]), .B(a[413]), .Z(n7393) );
  NAND U8680 ( .A(a[412]), .B(b[1]), .Z(n7392) );
  XNOR U8681 ( .A(n7393), .B(n7392), .Z(n7395) );
  XNOR U8682 ( .A(n7394), .B(n7395), .Z(n7399) );
  XOR U8683 ( .A(n7398), .B(sreg[1435]), .Z(n7391) );
  XNOR U8684 ( .A(n7399), .B(n7391), .Z(c[1435]) );
  NAND U8685 ( .A(n7393), .B(n7392), .Z(n7397) );
  NANDN U8686 ( .A(n7395), .B(n7394), .Z(n7396) );
  NAND U8687 ( .A(n7397), .B(n7396), .Z(n7404) );
  ANDN U8688 ( .B(a[414]), .A(n3944), .Z(n7402) );
  AND U8689 ( .A(b[1]), .B(a[413]), .Z(n7401) );
  XOR U8690 ( .A(n7402), .B(n7401), .Z(n7403) );
  XNOR U8691 ( .A(n7404), .B(n7403), .Z(n7406) );
  XOR U8692 ( .A(sreg[1436]), .B(n7405), .Z(n7400) );
  XNOR U8693 ( .A(n7406), .B(n7400), .Z(c[1436]) );
  NAND U8694 ( .A(b[0]), .B(a[415]), .Z(n7409) );
  NAND U8695 ( .A(a[414]), .B(b[1]), .Z(n7408) );
  XNOR U8696 ( .A(n7409), .B(n7408), .Z(n7411) );
  XNOR U8697 ( .A(n7410), .B(n7411), .Z(n7415) );
  XOR U8698 ( .A(n7414), .B(sreg[1437]), .Z(n7407) );
  XNOR U8699 ( .A(n7415), .B(n7407), .Z(c[1437]) );
  NAND U8700 ( .A(n7409), .B(n7408), .Z(n7413) );
  NANDN U8701 ( .A(n7411), .B(n7410), .Z(n7412) );
  NAND U8702 ( .A(n7413), .B(n7412), .Z(n7420) );
  ANDN U8703 ( .B(a[416]), .A(n3944), .Z(n7418) );
  AND U8704 ( .A(b[1]), .B(a[415]), .Z(n7417) );
  XOR U8705 ( .A(n7418), .B(n7417), .Z(n7419) );
  XNOR U8706 ( .A(n7420), .B(n7419), .Z(n7422) );
  XOR U8707 ( .A(sreg[1438]), .B(n7421), .Z(n7416) );
  XNOR U8708 ( .A(n7422), .B(n7416), .Z(c[1438]) );
  NAND U8709 ( .A(b[0]), .B(a[417]), .Z(n7425) );
  NAND U8710 ( .A(a[416]), .B(b[1]), .Z(n7424) );
  XNOR U8711 ( .A(n7425), .B(n7424), .Z(n7427) );
  XNOR U8712 ( .A(n7426), .B(n7427), .Z(n7431) );
  XOR U8713 ( .A(n7430), .B(sreg[1439]), .Z(n7423) );
  XNOR U8714 ( .A(n7431), .B(n7423), .Z(c[1439]) );
  NAND U8715 ( .A(n7425), .B(n7424), .Z(n7429) );
  NANDN U8716 ( .A(n7427), .B(n7426), .Z(n7428) );
  NAND U8717 ( .A(n7429), .B(n7428), .Z(n7436) );
  ANDN U8718 ( .B(a[418]), .A(n3945), .Z(n7434) );
  AND U8719 ( .A(b[1]), .B(a[417]), .Z(n7433) );
  XOR U8720 ( .A(n7434), .B(n7433), .Z(n7435) );
  XNOR U8721 ( .A(n7436), .B(n7435), .Z(n7441) );
  XOR U8722 ( .A(sreg[1440]), .B(n7440), .Z(n7432) );
  XNOR U8723 ( .A(n7441), .B(n7432), .Z(c[1440]) );
  OR U8724 ( .A(n7434), .B(n7433), .Z(n7439) );
  IV U8725 ( .A(n7435), .Z(n7437) );
  NANDN U8726 ( .A(n7437), .B(n7436), .Z(n7438) );
  NAND U8727 ( .A(n7439), .B(n7438), .Z(n7445) );
  NAND U8728 ( .A(b[0]), .B(a[419]), .Z(n7444) );
  NAND U8729 ( .A(a[418]), .B(b[1]), .Z(n7443) );
  XNOR U8730 ( .A(n7444), .B(n7443), .Z(n7446) );
  XNOR U8731 ( .A(n7445), .B(n7446), .Z(n7450) );
  XOR U8732 ( .A(n7449), .B(sreg[1441]), .Z(n7442) );
  XNOR U8733 ( .A(n7450), .B(n7442), .Z(c[1441]) );
  NAND U8734 ( .A(n7444), .B(n7443), .Z(n7448) );
  NANDN U8735 ( .A(n7446), .B(n7445), .Z(n7447) );
  NAND U8736 ( .A(n7448), .B(n7447), .Z(n7455) );
  ANDN U8737 ( .B(a[420]), .A(n3945), .Z(n7453) );
  AND U8738 ( .A(b[1]), .B(a[419]), .Z(n7452) );
  XOR U8739 ( .A(n7453), .B(n7452), .Z(n7454) );
  XNOR U8740 ( .A(n7455), .B(n7454), .Z(n7457) );
  XOR U8741 ( .A(sreg[1442]), .B(n7456), .Z(n7451) );
  XNOR U8742 ( .A(n7457), .B(n7451), .Z(c[1442]) );
  ANDN U8743 ( .B(a[421]), .A(n3945), .Z(n7460) );
  AND U8744 ( .A(b[1]), .B(a[420]), .Z(n7459) );
  XOR U8745 ( .A(n7460), .B(n7459), .Z(n7461) );
  XNOR U8746 ( .A(n7462), .B(n7461), .Z(n7464) );
  XNOR U8747 ( .A(sreg[1443]), .B(n7463), .Z(n7458) );
  XNOR U8748 ( .A(n7464), .B(n7458), .Z(c[1443]) );
  NAND U8749 ( .A(b[0]), .B(a[422]), .Z(n7467) );
  NAND U8750 ( .A(a[421]), .B(b[1]), .Z(n7466) );
  XNOR U8751 ( .A(n7467), .B(n7466), .Z(n7469) );
  XNOR U8752 ( .A(n7468), .B(n7469), .Z(n7473) );
  XOR U8753 ( .A(n7472), .B(sreg[1444]), .Z(n7465) );
  XNOR U8754 ( .A(n7473), .B(n7465), .Z(c[1444]) );
  NAND U8755 ( .A(n7467), .B(n7466), .Z(n7471) );
  NANDN U8756 ( .A(n7469), .B(n7468), .Z(n7470) );
  NAND U8757 ( .A(n7471), .B(n7470), .Z(n7477) );
  NAND U8758 ( .A(b[0]), .B(a[423]), .Z(n7476) );
  NAND U8759 ( .A(a[422]), .B(b[1]), .Z(n7475) );
  XNOR U8760 ( .A(n7476), .B(n7475), .Z(n7478) );
  XNOR U8761 ( .A(n7477), .B(n7478), .Z(n7482) );
  XOR U8762 ( .A(n7481), .B(sreg[1445]), .Z(n7474) );
  XNOR U8763 ( .A(n7482), .B(n7474), .Z(c[1445]) );
  NAND U8764 ( .A(n7476), .B(n7475), .Z(n7480) );
  NANDN U8765 ( .A(n7478), .B(n7477), .Z(n7479) );
  NAND U8766 ( .A(n7480), .B(n7479), .Z(n7487) );
  ANDN U8767 ( .B(a[424]), .A(n3945), .Z(n7485) );
  AND U8768 ( .A(b[1]), .B(a[423]), .Z(n7484) );
  XOR U8769 ( .A(n7485), .B(n7484), .Z(n7486) );
  XNOR U8770 ( .A(n7487), .B(n7486), .Z(n7489) );
  XOR U8771 ( .A(sreg[1446]), .B(n7488), .Z(n7483) );
  XNOR U8772 ( .A(n7489), .B(n7483), .Z(c[1446]) );
  ANDN U8773 ( .B(a[425]), .A(n3945), .Z(n7492) );
  AND U8774 ( .A(b[1]), .B(a[424]), .Z(n7491) );
  XOR U8775 ( .A(n7492), .B(n7491), .Z(n7493) );
  XNOR U8776 ( .A(n7494), .B(n7493), .Z(n7496) );
  XNOR U8777 ( .A(sreg[1447]), .B(n7495), .Z(n7490) );
  XNOR U8778 ( .A(n7496), .B(n7490), .Z(c[1447]) );
  ANDN U8779 ( .B(a[426]), .A(n3945), .Z(n7499) );
  AND U8780 ( .A(b[1]), .B(a[425]), .Z(n7498) );
  XOR U8781 ( .A(n7499), .B(n7498), .Z(n7500) );
  XNOR U8782 ( .A(n7501), .B(n7500), .Z(n7503) );
  XNOR U8783 ( .A(sreg[1448]), .B(n7502), .Z(n7497) );
  XNOR U8784 ( .A(n7503), .B(n7497), .Z(c[1448]) );
  ANDN U8785 ( .B(a[427]), .A(n3945), .Z(n7506) );
  AND U8786 ( .A(b[1]), .B(a[426]), .Z(n7505) );
  XOR U8787 ( .A(n7506), .B(n7505), .Z(n7507) );
  XNOR U8788 ( .A(n7508), .B(n7507), .Z(n7510) );
  XNOR U8789 ( .A(sreg[1449]), .B(n7509), .Z(n7504) );
  XNOR U8790 ( .A(n7510), .B(n7504), .Z(c[1449]) );
  NAND U8791 ( .A(b[0]), .B(a[428]), .Z(n7513) );
  NAND U8792 ( .A(a[427]), .B(b[1]), .Z(n7512) );
  XNOR U8793 ( .A(n7513), .B(n7512), .Z(n7515) );
  XNOR U8794 ( .A(n7514), .B(n7515), .Z(n7519) );
  XOR U8795 ( .A(n7518), .B(sreg[1450]), .Z(n7511) );
  XNOR U8796 ( .A(n7519), .B(n7511), .Z(c[1450]) );
  NAND U8797 ( .A(n7513), .B(n7512), .Z(n7517) );
  NANDN U8798 ( .A(n7515), .B(n7514), .Z(n7516) );
  NAND U8799 ( .A(n7517), .B(n7516), .Z(n7523) );
  NAND U8800 ( .A(b[0]), .B(a[429]), .Z(n7522) );
  NAND U8801 ( .A(a[428]), .B(b[1]), .Z(n7521) );
  XNOR U8802 ( .A(n7522), .B(n7521), .Z(n7524) );
  XNOR U8803 ( .A(n7523), .B(n7524), .Z(n7528) );
  XOR U8804 ( .A(n7527), .B(sreg[1451]), .Z(n7520) );
  XNOR U8805 ( .A(n7528), .B(n7520), .Z(c[1451]) );
  NAND U8806 ( .A(n7522), .B(n7521), .Z(n7526) );
  NANDN U8807 ( .A(n7524), .B(n7523), .Z(n7525) );
  NAND U8808 ( .A(n7526), .B(n7525), .Z(n7533) );
  ANDN U8809 ( .B(a[430]), .A(n3946), .Z(n7531) );
  AND U8810 ( .A(b[1]), .B(a[429]), .Z(n7530) );
  XOR U8811 ( .A(n7531), .B(n7530), .Z(n7532) );
  XNOR U8812 ( .A(n7533), .B(n7532), .Z(n7538) );
  XOR U8813 ( .A(sreg[1452]), .B(n7537), .Z(n7529) );
  XNOR U8814 ( .A(n7538), .B(n7529), .Z(c[1452]) );
  OR U8815 ( .A(n7531), .B(n7530), .Z(n7536) );
  IV U8816 ( .A(n7532), .Z(n7534) );
  NANDN U8817 ( .A(n7534), .B(n7533), .Z(n7535) );
  NAND U8818 ( .A(n7536), .B(n7535), .Z(n7542) );
  NAND U8819 ( .A(b[0]), .B(a[431]), .Z(n7541) );
  NAND U8820 ( .A(a[430]), .B(b[1]), .Z(n7540) );
  XNOR U8821 ( .A(n7541), .B(n7540), .Z(n7543) );
  XNOR U8822 ( .A(n7542), .B(n7543), .Z(n7547) );
  XOR U8823 ( .A(n7546), .B(sreg[1453]), .Z(n7539) );
  XNOR U8824 ( .A(n7547), .B(n7539), .Z(c[1453]) );
  NAND U8825 ( .A(n7541), .B(n7540), .Z(n7545) );
  NANDN U8826 ( .A(n7543), .B(n7542), .Z(n7544) );
  NAND U8827 ( .A(n7545), .B(n7544), .Z(n7552) );
  ANDN U8828 ( .B(a[432]), .A(n3946), .Z(n7550) );
  AND U8829 ( .A(b[1]), .B(a[431]), .Z(n7549) );
  XOR U8830 ( .A(n7550), .B(n7549), .Z(n7551) );
  XNOR U8831 ( .A(n7552), .B(n7551), .Z(n7554) );
  XOR U8832 ( .A(sreg[1454]), .B(n7553), .Z(n7548) );
  XNOR U8833 ( .A(n7554), .B(n7548), .Z(c[1454]) );
  NAND U8834 ( .A(b[0]), .B(a[433]), .Z(n7557) );
  NAND U8835 ( .A(a[432]), .B(b[1]), .Z(n7556) );
  XNOR U8836 ( .A(n7557), .B(n7556), .Z(n7559) );
  XNOR U8837 ( .A(n7558), .B(n7559), .Z(n7563) );
  XOR U8838 ( .A(n7562), .B(sreg[1455]), .Z(n7555) );
  XNOR U8839 ( .A(n7563), .B(n7555), .Z(c[1455]) );
  NAND U8840 ( .A(n7557), .B(n7556), .Z(n7561) );
  NANDN U8841 ( .A(n7559), .B(n7558), .Z(n7560) );
  NAND U8842 ( .A(n7561), .B(n7560), .Z(n7567) );
  NAND U8843 ( .A(b[0]), .B(a[434]), .Z(n7566) );
  NAND U8844 ( .A(a[433]), .B(b[1]), .Z(n7565) );
  XNOR U8845 ( .A(n7566), .B(n7565), .Z(n7568) );
  XNOR U8846 ( .A(n7567), .B(n7568), .Z(n7572) );
  XOR U8847 ( .A(n7571), .B(sreg[1456]), .Z(n7564) );
  XNOR U8848 ( .A(n7572), .B(n7564), .Z(c[1456]) );
  NAND U8849 ( .A(n7566), .B(n7565), .Z(n7570) );
  NANDN U8850 ( .A(n7568), .B(n7567), .Z(n7569) );
  NAND U8851 ( .A(n7570), .B(n7569), .Z(n7576) );
  NAND U8852 ( .A(b[0]), .B(a[435]), .Z(n7575) );
  NAND U8853 ( .A(a[434]), .B(b[1]), .Z(n7574) );
  XNOR U8854 ( .A(n7575), .B(n7574), .Z(n7577) );
  XNOR U8855 ( .A(n7576), .B(n7577), .Z(n7581) );
  XOR U8856 ( .A(n7580), .B(sreg[1457]), .Z(n7573) );
  XNOR U8857 ( .A(n7581), .B(n7573), .Z(c[1457]) );
  NAND U8858 ( .A(n7575), .B(n7574), .Z(n7579) );
  NANDN U8859 ( .A(n7577), .B(n7576), .Z(n7578) );
  NAND U8860 ( .A(n7579), .B(n7578), .Z(n7586) );
  ANDN U8861 ( .B(a[436]), .A(n3946), .Z(n7584) );
  AND U8862 ( .A(b[1]), .B(a[435]), .Z(n7583) );
  XOR U8863 ( .A(n7584), .B(n7583), .Z(n7585) );
  XNOR U8864 ( .A(n7586), .B(n7585), .Z(n7588) );
  XOR U8865 ( .A(sreg[1458]), .B(n7587), .Z(n7582) );
  XNOR U8866 ( .A(n7588), .B(n7582), .Z(c[1458]) );
  ANDN U8867 ( .B(a[437]), .A(n3946), .Z(n7591) );
  AND U8868 ( .A(b[1]), .B(a[436]), .Z(n7590) );
  XOR U8869 ( .A(n7591), .B(n7590), .Z(n7592) );
  XNOR U8870 ( .A(n7593), .B(n7592), .Z(n7595) );
  XNOR U8871 ( .A(sreg[1459]), .B(n7594), .Z(n7589) );
  XNOR U8872 ( .A(n7595), .B(n7589), .Z(c[1459]) );
  ANDN U8873 ( .B(a[438]), .A(n3946), .Z(n7598) );
  AND U8874 ( .A(b[1]), .B(a[437]), .Z(n7597) );
  XOR U8875 ( .A(n7598), .B(n7597), .Z(n7599) );
  XNOR U8876 ( .A(n7600), .B(n7599), .Z(n7602) );
  XNOR U8877 ( .A(sreg[1460]), .B(n7601), .Z(n7596) );
  XNOR U8878 ( .A(n7602), .B(n7596), .Z(c[1460]) );
  NAND U8879 ( .A(b[0]), .B(a[439]), .Z(n7605) );
  NAND U8880 ( .A(a[438]), .B(b[1]), .Z(n7604) );
  XNOR U8881 ( .A(n7605), .B(n7604), .Z(n7607) );
  XNOR U8882 ( .A(n7606), .B(n7607), .Z(n7611) );
  XOR U8883 ( .A(n7610), .B(sreg[1461]), .Z(n7603) );
  XNOR U8884 ( .A(n7611), .B(n7603), .Z(c[1461]) );
  NAND U8885 ( .A(n7605), .B(n7604), .Z(n7609) );
  NANDN U8886 ( .A(n7607), .B(n7606), .Z(n7608) );
  NAND U8887 ( .A(n7609), .B(n7608), .Z(n7616) );
  ANDN U8888 ( .B(a[440]), .A(n3946), .Z(n7614) );
  AND U8889 ( .A(b[1]), .B(a[439]), .Z(n7613) );
  XOR U8890 ( .A(n7614), .B(n7613), .Z(n7615) );
  XNOR U8891 ( .A(n7616), .B(n7615), .Z(n7618) );
  XOR U8892 ( .A(sreg[1462]), .B(n7617), .Z(n7612) );
  XNOR U8893 ( .A(n7618), .B(n7612), .Z(c[1462]) );
  NAND U8894 ( .A(b[0]), .B(a[441]), .Z(n7621) );
  NAND U8895 ( .A(a[440]), .B(b[1]), .Z(n7620) );
  XNOR U8896 ( .A(n7621), .B(n7620), .Z(n7623) );
  XNOR U8897 ( .A(n7622), .B(n7623), .Z(n7627) );
  XOR U8898 ( .A(n7626), .B(sreg[1463]), .Z(n7619) );
  XNOR U8899 ( .A(n7627), .B(n7619), .Z(c[1463]) );
  NAND U8900 ( .A(n7621), .B(n7620), .Z(n7625) );
  NANDN U8901 ( .A(n7623), .B(n7622), .Z(n7624) );
  NAND U8902 ( .A(n7625), .B(n7624), .Z(n7632) );
  ANDN U8903 ( .B(a[442]), .A(n3946), .Z(n7630) );
  AND U8904 ( .A(b[1]), .B(a[441]), .Z(n7629) );
  XOR U8905 ( .A(n7630), .B(n7629), .Z(n7631) );
  XNOR U8906 ( .A(n7632), .B(n7631), .Z(n7634) );
  XOR U8907 ( .A(sreg[1464]), .B(n7633), .Z(n7628) );
  XNOR U8908 ( .A(n7634), .B(n7628), .Z(c[1464]) );
  NAND U8909 ( .A(b[0]), .B(a[443]), .Z(n7637) );
  NAND U8910 ( .A(a[442]), .B(b[1]), .Z(n7636) );
  XNOR U8911 ( .A(n7637), .B(n7636), .Z(n7639) );
  XNOR U8912 ( .A(n7638), .B(n7639), .Z(n7643) );
  XOR U8913 ( .A(n7642), .B(sreg[1465]), .Z(n7635) );
  XNOR U8914 ( .A(n7643), .B(n7635), .Z(c[1465]) );
  NAND U8915 ( .A(n7637), .B(n7636), .Z(n7641) );
  NANDN U8916 ( .A(n7639), .B(n7638), .Z(n7640) );
  NAND U8917 ( .A(n7641), .B(n7640), .Z(n7648) );
  ANDN U8918 ( .B(a[444]), .A(n3947), .Z(n7646) );
  AND U8919 ( .A(b[1]), .B(a[443]), .Z(n7645) );
  XOR U8920 ( .A(n7646), .B(n7645), .Z(n7647) );
  XNOR U8921 ( .A(n7648), .B(n7647), .Z(n7653) );
  XOR U8922 ( .A(sreg[1466]), .B(n7652), .Z(n7644) );
  XNOR U8923 ( .A(n7653), .B(n7644), .Z(c[1466]) );
  OR U8924 ( .A(n7646), .B(n7645), .Z(n7651) );
  IV U8925 ( .A(n7647), .Z(n7649) );
  NANDN U8926 ( .A(n7649), .B(n7648), .Z(n7650) );
  NAND U8927 ( .A(n7651), .B(n7650), .Z(n7657) );
  NAND U8928 ( .A(b[0]), .B(a[445]), .Z(n7656) );
  NAND U8929 ( .A(a[444]), .B(b[1]), .Z(n7655) );
  XNOR U8930 ( .A(n7656), .B(n7655), .Z(n7658) );
  XNOR U8931 ( .A(n7657), .B(n7658), .Z(n7662) );
  XOR U8932 ( .A(n7661), .B(sreg[1467]), .Z(n7654) );
  XNOR U8933 ( .A(n7662), .B(n7654), .Z(c[1467]) );
  NAND U8934 ( .A(n7656), .B(n7655), .Z(n7660) );
  NANDN U8935 ( .A(n7658), .B(n7657), .Z(n7659) );
  NAND U8936 ( .A(n7660), .B(n7659), .Z(n7667) );
  ANDN U8937 ( .B(a[446]), .A(n3947), .Z(n7665) );
  AND U8938 ( .A(b[1]), .B(a[445]), .Z(n7664) );
  XOR U8939 ( .A(n7665), .B(n7664), .Z(n7666) );
  XNOR U8940 ( .A(n7667), .B(n7666), .Z(n7669) );
  XOR U8941 ( .A(sreg[1468]), .B(n7668), .Z(n7663) );
  XNOR U8942 ( .A(n7669), .B(n7663), .Z(c[1468]) );
  NAND U8943 ( .A(b[0]), .B(a[447]), .Z(n7672) );
  NAND U8944 ( .A(a[446]), .B(b[1]), .Z(n7671) );
  XNOR U8945 ( .A(n7672), .B(n7671), .Z(n7674) );
  XNOR U8946 ( .A(n7673), .B(n7674), .Z(n7678) );
  XOR U8947 ( .A(n7677), .B(sreg[1469]), .Z(n7670) );
  XNOR U8948 ( .A(n7678), .B(n7670), .Z(c[1469]) );
  NAND U8949 ( .A(n7672), .B(n7671), .Z(n7676) );
  NANDN U8950 ( .A(n7674), .B(n7673), .Z(n7675) );
  NAND U8951 ( .A(n7676), .B(n7675), .Z(n7683) );
  ANDN U8952 ( .B(a[448]), .A(n3947), .Z(n7681) );
  AND U8953 ( .A(b[1]), .B(a[447]), .Z(n7680) );
  XOR U8954 ( .A(n7681), .B(n7680), .Z(n7682) );
  XNOR U8955 ( .A(n7683), .B(n7682), .Z(n7685) );
  XOR U8956 ( .A(sreg[1470]), .B(n7684), .Z(n7679) );
  XNOR U8957 ( .A(n7685), .B(n7679), .Z(c[1470]) );
  NAND U8958 ( .A(b[0]), .B(a[449]), .Z(n7688) );
  NAND U8959 ( .A(a[448]), .B(b[1]), .Z(n7687) );
  XNOR U8960 ( .A(n7688), .B(n7687), .Z(n7690) );
  XNOR U8961 ( .A(n7689), .B(n7690), .Z(n7694) );
  XOR U8962 ( .A(n7693), .B(sreg[1471]), .Z(n7686) );
  XNOR U8963 ( .A(n7694), .B(n7686), .Z(c[1471]) );
  NAND U8964 ( .A(n7688), .B(n7687), .Z(n7692) );
  NANDN U8965 ( .A(n7690), .B(n7689), .Z(n7691) );
  NAND U8966 ( .A(n7692), .B(n7691), .Z(n7699) );
  ANDN U8967 ( .B(a[450]), .A(n3947), .Z(n7697) );
  AND U8968 ( .A(b[1]), .B(a[449]), .Z(n7696) );
  XOR U8969 ( .A(n7697), .B(n7696), .Z(n7698) );
  XNOR U8970 ( .A(n7699), .B(n7698), .Z(n7701) );
  XOR U8971 ( .A(sreg[1472]), .B(n7700), .Z(n7695) );
  XNOR U8972 ( .A(n7701), .B(n7695), .Z(c[1472]) );
  NAND U8973 ( .A(b[0]), .B(a[451]), .Z(n7704) );
  NAND U8974 ( .A(a[450]), .B(b[1]), .Z(n7703) );
  XNOR U8975 ( .A(n7704), .B(n7703), .Z(n7706) );
  XNOR U8976 ( .A(n7705), .B(n7706), .Z(n7710) );
  XOR U8977 ( .A(n7709), .B(sreg[1473]), .Z(n7702) );
  XNOR U8978 ( .A(n7710), .B(n7702), .Z(c[1473]) );
  NAND U8979 ( .A(n7704), .B(n7703), .Z(n7708) );
  NANDN U8980 ( .A(n7706), .B(n7705), .Z(n7707) );
  NAND U8981 ( .A(n7708), .B(n7707), .Z(n7715) );
  ANDN U8982 ( .B(a[452]), .A(n3947), .Z(n7713) );
  AND U8983 ( .A(b[1]), .B(a[451]), .Z(n7712) );
  XOR U8984 ( .A(n7713), .B(n7712), .Z(n7714) );
  XNOR U8985 ( .A(n7715), .B(n7714), .Z(n7717) );
  XOR U8986 ( .A(sreg[1474]), .B(n7716), .Z(n7711) );
  XNOR U8987 ( .A(n7717), .B(n7711), .Z(c[1474]) );
  NAND U8988 ( .A(b[0]), .B(a[453]), .Z(n7720) );
  NAND U8989 ( .A(a[452]), .B(b[1]), .Z(n7719) );
  XNOR U8990 ( .A(n7720), .B(n7719), .Z(n7722) );
  XNOR U8991 ( .A(n7721), .B(n7722), .Z(n7726) );
  XOR U8992 ( .A(n7725), .B(sreg[1475]), .Z(n7718) );
  XNOR U8993 ( .A(n7726), .B(n7718), .Z(c[1475]) );
  NAND U8994 ( .A(n7720), .B(n7719), .Z(n7724) );
  NANDN U8995 ( .A(n7722), .B(n7721), .Z(n7723) );
  NAND U8996 ( .A(n7724), .B(n7723), .Z(n7730) );
  NAND U8997 ( .A(b[0]), .B(a[454]), .Z(n7729) );
  NAND U8998 ( .A(a[453]), .B(b[1]), .Z(n7728) );
  XNOR U8999 ( .A(n7729), .B(n7728), .Z(n7731) );
  XNOR U9000 ( .A(n7730), .B(n7731), .Z(n7735) );
  XOR U9001 ( .A(n7734), .B(sreg[1476]), .Z(n7727) );
  XNOR U9002 ( .A(n7735), .B(n7727), .Z(c[1476]) );
  NAND U9003 ( .A(n7729), .B(n7728), .Z(n7733) );
  NANDN U9004 ( .A(n7731), .B(n7730), .Z(n7732) );
  NAND U9005 ( .A(n7733), .B(n7732), .Z(n7739) );
  NAND U9006 ( .A(b[0]), .B(a[455]), .Z(n7738) );
  NAND U9007 ( .A(a[454]), .B(b[1]), .Z(n7737) );
  XNOR U9008 ( .A(n7738), .B(n7737), .Z(n7740) );
  XNOR U9009 ( .A(n7739), .B(n7740), .Z(n7744) );
  XOR U9010 ( .A(n7743), .B(sreg[1477]), .Z(n7736) );
  XNOR U9011 ( .A(n7744), .B(n7736), .Z(c[1477]) );
  NAND U9012 ( .A(n7738), .B(n7737), .Z(n7742) );
  NANDN U9013 ( .A(n7740), .B(n7739), .Z(n7741) );
  NAND U9014 ( .A(n7742), .B(n7741), .Z(n7749) );
  ANDN U9015 ( .B(a[456]), .A(n3947), .Z(n7747) );
  AND U9016 ( .A(b[1]), .B(a[455]), .Z(n7746) );
  XOR U9017 ( .A(n7747), .B(n7746), .Z(n7748) );
  XNOR U9018 ( .A(n7749), .B(n7748), .Z(n7751) );
  XOR U9019 ( .A(sreg[1478]), .B(n7750), .Z(n7745) );
  XNOR U9020 ( .A(n7751), .B(n7745), .Z(c[1478]) );
  NAND U9021 ( .A(b[0]), .B(a[457]), .Z(n7754) );
  NAND U9022 ( .A(a[456]), .B(b[1]), .Z(n7753) );
  XNOR U9023 ( .A(n7754), .B(n7753), .Z(n7756) );
  XNOR U9024 ( .A(n7755), .B(n7756), .Z(n7760) );
  XOR U9025 ( .A(n7759), .B(sreg[1479]), .Z(n7752) );
  XNOR U9026 ( .A(n7760), .B(n7752), .Z(c[1479]) );
  NAND U9027 ( .A(n7754), .B(n7753), .Z(n7758) );
  NANDN U9028 ( .A(n7756), .B(n7755), .Z(n7757) );
  NAND U9029 ( .A(n7758), .B(n7757), .Z(n7765) );
  ANDN U9030 ( .B(a[458]), .A(n3947), .Z(n7763) );
  AND U9031 ( .A(b[1]), .B(a[457]), .Z(n7762) );
  XOR U9032 ( .A(n7763), .B(n7762), .Z(n7764) );
  XNOR U9033 ( .A(n7765), .B(n7764), .Z(n7767) );
  XOR U9034 ( .A(sreg[1480]), .B(n7766), .Z(n7761) );
  XNOR U9035 ( .A(n7767), .B(n7761), .Z(c[1480]) );
  ANDN U9036 ( .B(a[459]), .A(n3948), .Z(n7770) );
  AND U9037 ( .A(b[1]), .B(a[458]), .Z(n7769) );
  XOR U9038 ( .A(n7770), .B(n7769), .Z(n7771) );
  XNOR U9039 ( .A(n7772), .B(n7771), .Z(n7777) );
  XNOR U9040 ( .A(sreg[1481]), .B(n7776), .Z(n7768) );
  XNOR U9041 ( .A(n7777), .B(n7768), .Z(c[1481]) );
  OR U9042 ( .A(n7770), .B(n7769), .Z(n7775) );
  IV U9043 ( .A(n7771), .Z(n7773) );
  NANDN U9044 ( .A(n7773), .B(n7772), .Z(n7774) );
  NAND U9045 ( .A(n7775), .B(n7774), .Z(n7781) );
  NAND U9046 ( .A(b[0]), .B(a[460]), .Z(n7780) );
  NAND U9047 ( .A(a[459]), .B(b[1]), .Z(n7779) );
  XNOR U9048 ( .A(n7780), .B(n7779), .Z(n7782) );
  XNOR U9049 ( .A(n7781), .B(n7782), .Z(n7786) );
  XOR U9050 ( .A(n7785), .B(sreg[1482]), .Z(n7778) );
  XNOR U9051 ( .A(n7786), .B(n7778), .Z(c[1482]) );
  NAND U9052 ( .A(n7780), .B(n7779), .Z(n7784) );
  NANDN U9053 ( .A(n7782), .B(n7781), .Z(n7783) );
  NAND U9054 ( .A(n7784), .B(n7783), .Z(n7791) );
  ANDN U9055 ( .B(a[461]), .A(n3948), .Z(n7789) );
  AND U9056 ( .A(b[1]), .B(a[460]), .Z(n7788) );
  XOR U9057 ( .A(n7789), .B(n7788), .Z(n7790) );
  XNOR U9058 ( .A(n7791), .B(n7790), .Z(n7793) );
  XOR U9059 ( .A(sreg[1483]), .B(n7792), .Z(n7787) );
  XNOR U9060 ( .A(n7793), .B(n7787), .Z(c[1483]) );
  ANDN U9061 ( .B(a[462]), .A(n3948), .Z(n7796) );
  AND U9062 ( .A(b[1]), .B(a[461]), .Z(n7795) );
  XOR U9063 ( .A(n7796), .B(n7795), .Z(n7797) );
  XNOR U9064 ( .A(n7798), .B(n7797), .Z(n7800) );
  XNOR U9065 ( .A(sreg[1484]), .B(n7799), .Z(n7794) );
  XNOR U9066 ( .A(n7800), .B(n7794), .Z(c[1484]) );
  ANDN U9067 ( .B(a[463]), .A(n3948), .Z(n7803) );
  AND U9068 ( .A(b[1]), .B(a[462]), .Z(n7802) );
  XOR U9069 ( .A(n7803), .B(n7802), .Z(n7804) );
  XNOR U9070 ( .A(n7805), .B(n7804), .Z(n7807) );
  XNOR U9071 ( .A(sreg[1485]), .B(n7806), .Z(n7801) );
  XNOR U9072 ( .A(n7807), .B(n7801), .Z(c[1485]) );
  ANDN U9073 ( .B(a[464]), .A(n3948), .Z(n7810) );
  AND U9074 ( .A(b[1]), .B(a[463]), .Z(n7809) );
  XOR U9075 ( .A(n7810), .B(n7809), .Z(n7811) );
  XNOR U9076 ( .A(n7812), .B(n7811), .Z(n7814) );
  XNOR U9077 ( .A(sreg[1486]), .B(n7813), .Z(n7808) );
  XNOR U9078 ( .A(n7814), .B(n7808), .Z(c[1486]) );
  NAND U9079 ( .A(b[0]), .B(a[465]), .Z(n7817) );
  NAND U9080 ( .A(a[464]), .B(b[1]), .Z(n7816) );
  XNOR U9081 ( .A(n7817), .B(n7816), .Z(n7819) );
  XNOR U9082 ( .A(n7818), .B(n7819), .Z(n7823) );
  XOR U9083 ( .A(n7822), .B(sreg[1487]), .Z(n7815) );
  XNOR U9084 ( .A(n7823), .B(n7815), .Z(c[1487]) );
  NAND U9085 ( .A(n7817), .B(n7816), .Z(n7821) );
  NANDN U9086 ( .A(n7819), .B(n7818), .Z(n7820) );
  NAND U9087 ( .A(n7821), .B(n7820), .Z(n7828) );
  ANDN U9088 ( .B(a[466]), .A(n3948), .Z(n7826) );
  AND U9089 ( .A(b[1]), .B(a[465]), .Z(n7825) );
  XOR U9090 ( .A(n7826), .B(n7825), .Z(n7827) );
  XNOR U9091 ( .A(n7828), .B(n7827), .Z(n7830) );
  XOR U9092 ( .A(sreg[1488]), .B(n7829), .Z(n7824) );
  XNOR U9093 ( .A(n7830), .B(n7824), .Z(c[1488]) );
  NAND U9094 ( .A(b[0]), .B(a[467]), .Z(n7833) );
  NAND U9095 ( .A(a[466]), .B(b[1]), .Z(n7832) );
  XNOR U9096 ( .A(n7833), .B(n7832), .Z(n7835) );
  XNOR U9097 ( .A(n7834), .B(n7835), .Z(n7839) );
  XOR U9098 ( .A(n7838), .B(sreg[1489]), .Z(n7831) );
  XNOR U9099 ( .A(n7839), .B(n7831), .Z(c[1489]) );
  NAND U9100 ( .A(n7833), .B(n7832), .Z(n7837) );
  NANDN U9101 ( .A(n7835), .B(n7834), .Z(n7836) );
  NAND U9102 ( .A(n7837), .B(n7836), .Z(n7844) );
  ANDN U9103 ( .B(a[468]), .A(n3948), .Z(n7842) );
  AND U9104 ( .A(b[1]), .B(a[467]), .Z(n7841) );
  XOR U9105 ( .A(n7842), .B(n7841), .Z(n7843) );
  XNOR U9106 ( .A(n7844), .B(n7843), .Z(n7846) );
  XOR U9107 ( .A(sreg[1490]), .B(n7845), .Z(n7840) );
  XNOR U9108 ( .A(n7846), .B(n7840), .Z(c[1490]) );
  NAND U9109 ( .A(b[0]), .B(a[469]), .Z(n7849) );
  NAND U9110 ( .A(a[468]), .B(b[1]), .Z(n7848) );
  XNOR U9111 ( .A(n7849), .B(n7848), .Z(n7851) );
  XNOR U9112 ( .A(n7850), .B(n7851), .Z(n7855) );
  XOR U9113 ( .A(n7854), .B(sreg[1491]), .Z(n7847) );
  XNOR U9114 ( .A(n7855), .B(n7847), .Z(c[1491]) );
  NAND U9115 ( .A(n7849), .B(n7848), .Z(n7853) );
  NANDN U9116 ( .A(n7851), .B(n7850), .Z(n7852) );
  NAND U9117 ( .A(n7853), .B(n7852), .Z(n7860) );
  ANDN U9118 ( .B(a[470]), .A(n3949), .Z(n7858) );
  AND U9119 ( .A(b[1]), .B(a[469]), .Z(n7857) );
  XOR U9120 ( .A(n7858), .B(n7857), .Z(n7859) );
  XNOR U9121 ( .A(n7860), .B(n7859), .Z(n7865) );
  XOR U9122 ( .A(sreg[1492]), .B(n7864), .Z(n7856) );
  XNOR U9123 ( .A(n7865), .B(n7856), .Z(c[1492]) );
  OR U9124 ( .A(n7858), .B(n7857), .Z(n7863) );
  IV U9125 ( .A(n7859), .Z(n7861) );
  NANDN U9126 ( .A(n7861), .B(n7860), .Z(n7862) );
  NAND U9127 ( .A(n7863), .B(n7862), .Z(n7869) );
  NAND U9128 ( .A(b[0]), .B(a[471]), .Z(n7868) );
  NAND U9129 ( .A(a[470]), .B(b[1]), .Z(n7867) );
  XNOR U9130 ( .A(n7868), .B(n7867), .Z(n7870) );
  XNOR U9131 ( .A(n7869), .B(n7870), .Z(n7874) );
  XOR U9132 ( .A(n7873), .B(sreg[1493]), .Z(n7866) );
  XNOR U9133 ( .A(n7874), .B(n7866), .Z(c[1493]) );
  NAND U9134 ( .A(n7868), .B(n7867), .Z(n7872) );
  NANDN U9135 ( .A(n7870), .B(n7869), .Z(n7871) );
  NAND U9136 ( .A(n7872), .B(n7871), .Z(n7879) );
  ANDN U9137 ( .B(a[472]), .A(n3949), .Z(n7877) );
  AND U9138 ( .A(b[1]), .B(a[471]), .Z(n7876) );
  XOR U9139 ( .A(n7877), .B(n7876), .Z(n7878) );
  XNOR U9140 ( .A(n7879), .B(n7878), .Z(n7881) );
  XOR U9141 ( .A(sreg[1494]), .B(n7880), .Z(n7875) );
  XNOR U9142 ( .A(n7881), .B(n7875), .Z(c[1494]) );
  NAND U9143 ( .A(b[0]), .B(a[473]), .Z(n7884) );
  NAND U9144 ( .A(a[472]), .B(b[1]), .Z(n7883) );
  XNOR U9145 ( .A(n7884), .B(n7883), .Z(n7886) );
  XNOR U9146 ( .A(n7885), .B(n7886), .Z(n7890) );
  XOR U9147 ( .A(n7889), .B(sreg[1495]), .Z(n7882) );
  XNOR U9148 ( .A(n7890), .B(n7882), .Z(c[1495]) );
  NAND U9149 ( .A(n7884), .B(n7883), .Z(n7888) );
  NANDN U9150 ( .A(n7886), .B(n7885), .Z(n7887) );
  NAND U9151 ( .A(n7888), .B(n7887), .Z(n7895) );
  ANDN U9152 ( .B(a[474]), .A(n3949), .Z(n7893) );
  AND U9153 ( .A(b[1]), .B(a[473]), .Z(n7892) );
  XOR U9154 ( .A(n7893), .B(n7892), .Z(n7894) );
  XNOR U9155 ( .A(n7895), .B(n7894), .Z(n7897) );
  XOR U9156 ( .A(sreg[1496]), .B(n7896), .Z(n7891) );
  XNOR U9157 ( .A(n7897), .B(n7891), .Z(c[1496]) );
  NAND U9158 ( .A(b[0]), .B(a[475]), .Z(n7900) );
  NAND U9159 ( .A(a[474]), .B(b[1]), .Z(n7899) );
  XNOR U9160 ( .A(n7900), .B(n7899), .Z(n7902) );
  XNOR U9161 ( .A(n7901), .B(n7902), .Z(n7906) );
  XOR U9162 ( .A(n7905), .B(sreg[1497]), .Z(n7898) );
  XNOR U9163 ( .A(n7906), .B(n7898), .Z(c[1497]) );
  NAND U9164 ( .A(n7900), .B(n7899), .Z(n7904) );
  NANDN U9165 ( .A(n7902), .B(n7901), .Z(n7903) );
  NAND U9166 ( .A(n7904), .B(n7903), .Z(n7911) );
  ANDN U9167 ( .B(a[476]), .A(n3949), .Z(n7909) );
  AND U9168 ( .A(b[1]), .B(a[475]), .Z(n7908) );
  XOR U9169 ( .A(n7909), .B(n7908), .Z(n7910) );
  XNOR U9170 ( .A(n7911), .B(n7910), .Z(n7913) );
  XOR U9171 ( .A(sreg[1498]), .B(n7912), .Z(n7907) );
  XNOR U9172 ( .A(n7913), .B(n7907), .Z(c[1498]) );
  NAND U9173 ( .A(b[0]), .B(a[477]), .Z(n7916) );
  NAND U9174 ( .A(a[476]), .B(b[1]), .Z(n7915) );
  XNOR U9175 ( .A(n7916), .B(n7915), .Z(n7918) );
  XNOR U9176 ( .A(n7917), .B(n7918), .Z(n7922) );
  XOR U9177 ( .A(n7921), .B(sreg[1499]), .Z(n7914) );
  XNOR U9178 ( .A(n7922), .B(n7914), .Z(c[1499]) );
  NAND U9179 ( .A(n7916), .B(n7915), .Z(n7920) );
  NANDN U9180 ( .A(n7918), .B(n7917), .Z(n7919) );
  NAND U9181 ( .A(n7920), .B(n7919), .Z(n7927) );
  ANDN U9182 ( .B(a[478]), .A(n3949), .Z(n7925) );
  AND U9183 ( .A(b[1]), .B(a[477]), .Z(n7924) );
  XOR U9184 ( .A(n7925), .B(n7924), .Z(n7926) );
  XNOR U9185 ( .A(n7927), .B(n7926), .Z(n7929) );
  XOR U9186 ( .A(sreg[1500]), .B(n7928), .Z(n7923) );
  XNOR U9187 ( .A(n7929), .B(n7923), .Z(c[1500]) );
  NAND U9188 ( .A(b[0]), .B(a[479]), .Z(n7932) );
  NAND U9189 ( .A(a[478]), .B(b[1]), .Z(n7931) );
  XNOR U9190 ( .A(n7932), .B(n7931), .Z(n7934) );
  XNOR U9191 ( .A(n7933), .B(n7934), .Z(n7938) );
  XOR U9192 ( .A(n7937), .B(sreg[1501]), .Z(n7930) );
  XNOR U9193 ( .A(n7938), .B(n7930), .Z(c[1501]) );
  NAND U9194 ( .A(n7932), .B(n7931), .Z(n7936) );
  NANDN U9195 ( .A(n7934), .B(n7933), .Z(n7935) );
  NAND U9196 ( .A(n7936), .B(n7935), .Z(n7943) );
  ANDN U9197 ( .B(a[480]), .A(n3949), .Z(n7941) );
  AND U9198 ( .A(b[1]), .B(a[479]), .Z(n7940) );
  XOR U9199 ( .A(n7941), .B(n7940), .Z(n7942) );
  XNOR U9200 ( .A(n7943), .B(n7942), .Z(n7945) );
  XOR U9201 ( .A(sreg[1502]), .B(n7944), .Z(n7939) );
  XNOR U9202 ( .A(n7945), .B(n7939), .Z(c[1502]) );
  NAND U9203 ( .A(b[0]), .B(a[481]), .Z(n7948) );
  NAND U9204 ( .A(a[480]), .B(b[1]), .Z(n7947) );
  XNOR U9205 ( .A(n7948), .B(n7947), .Z(n7950) );
  XNOR U9206 ( .A(n7949), .B(n7950), .Z(n7954) );
  XOR U9207 ( .A(n7953), .B(sreg[1503]), .Z(n7946) );
  XNOR U9208 ( .A(n7954), .B(n7946), .Z(c[1503]) );
  NAND U9209 ( .A(n7948), .B(n7947), .Z(n7952) );
  NANDN U9210 ( .A(n7950), .B(n7949), .Z(n7951) );
  NAND U9211 ( .A(n7952), .B(n7951), .Z(n7959) );
  ANDN U9212 ( .B(a[482]), .A(n3949), .Z(n7957) );
  AND U9213 ( .A(b[1]), .B(a[481]), .Z(n7956) );
  XOR U9214 ( .A(n7957), .B(n7956), .Z(n7958) );
  XNOR U9215 ( .A(n7959), .B(n7958), .Z(n7961) );
  XOR U9216 ( .A(sreg[1504]), .B(n7960), .Z(n7955) );
  XNOR U9217 ( .A(n7961), .B(n7955), .Z(c[1504]) );
  NAND U9218 ( .A(b[0]), .B(a[483]), .Z(n7964) );
  NAND U9219 ( .A(a[482]), .B(b[1]), .Z(n7963) );
  XNOR U9220 ( .A(n7964), .B(n7963), .Z(n7966) );
  XNOR U9221 ( .A(n7965), .B(n7966), .Z(n7970) );
  XOR U9222 ( .A(n7969), .B(sreg[1505]), .Z(n7962) );
  XNOR U9223 ( .A(n7970), .B(n7962), .Z(c[1505]) );
  NAND U9224 ( .A(n7964), .B(n7963), .Z(n7968) );
  NANDN U9225 ( .A(n7966), .B(n7965), .Z(n7967) );
  NAND U9226 ( .A(n7968), .B(n7967), .Z(n7975) );
  ANDN U9227 ( .B(a[484]), .A(n3950), .Z(n7973) );
  AND U9228 ( .A(b[1]), .B(a[483]), .Z(n7972) );
  XOR U9229 ( .A(n7973), .B(n7972), .Z(n7974) );
  XNOR U9230 ( .A(n7975), .B(n7974), .Z(n7980) );
  XOR U9231 ( .A(sreg[1506]), .B(n7979), .Z(n7971) );
  XNOR U9232 ( .A(n7980), .B(n7971), .Z(c[1506]) );
  OR U9233 ( .A(n7973), .B(n7972), .Z(n7978) );
  IV U9234 ( .A(n7974), .Z(n7976) );
  NANDN U9235 ( .A(n7976), .B(n7975), .Z(n7977) );
  NAND U9236 ( .A(n7978), .B(n7977), .Z(n7985) );
  ANDN U9237 ( .B(a[485]), .A(n3950), .Z(n7983) );
  AND U9238 ( .A(b[1]), .B(a[484]), .Z(n7982) );
  XOR U9239 ( .A(n7983), .B(n7982), .Z(n7984) );
  XNOR U9240 ( .A(n7985), .B(n7984), .Z(n7987) );
  XNOR U9241 ( .A(sreg[1507]), .B(n7986), .Z(n7981) );
  XNOR U9242 ( .A(n7987), .B(n7981), .Z(c[1507]) );
  ANDN U9243 ( .B(a[486]), .A(n3950), .Z(n7990) );
  AND U9244 ( .A(b[1]), .B(a[485]), .Z(n7989) );
  XOR U9245 ( .A(n7990), .B(n7989), .Z(n7991) );
  XNOR U9246 ( .A(n7992), .B(n7991), .Z(n7994) );
  XNOR U9247 ( .A(sreg[1508]), .B(n7993), .Z(n7988) );
  XNOR U9248 ( .A(n7994), .B(n7988), .Z(c[1508]) );
  NAND U9249 ( .A(b[0]), .B(a[487]), .Z(n7997) );
  NAND U9250 ( .A(a[486]), .B(b[1]), .Z(n7996) );
  XNOR U9251 ( .A(n7997), .B(n7996), .Z(n7999) );
  XNOR U9252 ( .A(n7998), .B(n7999), .Z(n8003) );
  XOR U9253 ( .A(n8002), .B(sreg[1509]), .Z(n7995) );
  XNOR U9254 ( .A(n8003), .B(n7995), .Z(c[1509]) );
  NAND U9255 ( .A(n7997), .B(n7996), .Z(n8001) );
  NANDN U9256 ( .A(n7999), .B(n7998), .Z(n8000) );
  NAND U9257 ( .A(n8001), .B(n8000), .Z(n8008) );
  ANDN U9258 ( .B(a[488]), .A(n3950), .Z(n8006) );
  AND U9259 ( .A(b[1]), .B(a[487]), .Z(n8005) );
  XOR U9260 ( .A(n8006), .B(n8005), .Z(n8007) );
  XNOR U9261 ( .A(n8008), .B(n8007), .Z(n8010) );
  XOR U9262 ( .A(sreg[1510]), .B(n8009), .Z(n8004) );
  XNOR U9263 ( .A(n8010), .B(n8004), .Z(c[1510]) );
  ANDN U9264 ( .B(a[489]), .A(n3950), .Z(n8013) );
  AND U9265 ( .A(b[1]), .B(a[488]), .Z(n8012) );
  XOR U9266 ( .A(n8013), .B(n8012), .Z(n8014) );
  XNOR U9267 ( .A(n8015), .B(n8014), .Z(n8017) );
  XNOR U9268 ( .A(sreg[1511]), .B(n8016), .Z(n8011) );
  XNOR U9269 ( .A(n8017), .B(n8011), .Z(c[1511]) );
  NAND U9270 ( .A(b[0]), .B(a[490]), .Z(n8020) );
  NAND U9271 ( .A(a[489]), .B(b[1]), .Z(n8019) );
  XNOR U9272 ( .A(n8020), .B(n8019), .Z(n8022) );
  XNOR U9273 ( .A(n8021), .B(n8022), .Z(n8026) );
  XOR U9274 ( .A(n8025), .B(sreg[1512]), .Z(n8018) );
  XNOR U9275 ( .A(n8026), .B(n8018), .Z(c[1512]) );
  NAND U9276 ( .A(n8020), .B(n8019), .Z(n8024) );
  NANDN U9277 ( .A(n8022), .B(n8021), .Z(n8023) );
  NAND U9278 ( .A(n8024), .B(n8023), .Z(n8031) );
  ANDN U9279 ( .B(a[491]), .A(n3950), .Z(n8029) );
  AND U9280 ( .A(b[1]), .B(a[490]), .Z(n8028) );
  XOR U9281 ( .A(n8029), .B(n8028), .Z(n8030) );
  XNOR U9282 ( .A(n8031), .B(n8030), .Z(n8033) );
  XOR U9283 ( .A(sreg[1513]), .B(n8032), .Z(n8027) );
  XNOR U9284 ( .A(n8033), .B(n8027), .Z(c[1513]) );
  NAND U9285 ( .A(b[0]), .B(a[492]), .Z(n8036) );
  NAND U9286 ( .A(a[491]), .B(b[1]), .Z(n8035) );
  XNOR U9287 ( .A(n8036), .B(n8035), .Z(n8038) );
  XNOR U9288 ( .A(n8037), .B(n8038), .Z(n8042) );
  XOR U9289 ( .A(n8041), .B(sreg[1514]), .Z(n8034) );
  XNOR U9290 ( .A(n8042), .B(n8034), .Z(c[1514]) );
  NAND U9291 ( .A(n8036), .B(n8035), .Z(n8040) );
  NANDN U9292 ( .A(n8038), .B(n8037), .Z(n8039) );
  NAND U9293 ( .A(n8040), .B(n8039), .Z(n8047) );
  ANDN U9294 ( .B(a[493]), .A(n3950), .Z(n8045) );
  AND U9295 ( .A(b[1]), .B(a[492]), .Z(n8044) );
  XOR U9296 ( .A(n8045), .B(n8044), .Z(n8046) );
  XNOR U9297 ( .A(n8047), .B(n8046), .Z(n8049) );
  XOR U9298 ( .A(sreg[1515]), .B(n8048), .Z(n8043) );
  XNOR U9299 ( .A(n8049), .B(n8043), .Z(c[1515]) );
  ANDN U9300 ( .B(a[494]), .A(n3951), .Z(n8052) );
  AND U9301 ( .A(b[1]), .B(a[493]), .Z(n8051) );
  XOR U9302 ( .A(n8052), .B(n8051), .Z(n8053) );
  XNOR U9303 ( .A(n8054), .B(n8053), .Z(n8059) );
  XNOR U9304 ( .A(sreg[1516]), .B(n8058), .Z(n8050) );
  XNOR U9305 ( .A(n8059), .B(n8050), .Z(c[1516]) );
  OR U9306 ( .A(n8052), .B(n8051), .Z(n8057) );
  IV U9307 ( .A(n8053), .Z(n8055) );
  NANDN U9308 ( .A(n8055), .B(n8054), .Z(n8056) );
  NAND U9309 ( .A(n8057), .B(n8056), .Z(n8063) );
  NAND U9310 ( .A(b[0]), .B(a[495]), .Z(n8062) );
  NAND U9311 ( .A(a[494]), .B(b[1]), .Z(n8061) );
  XNOR U9312 ( .A(n8062), .B(n8061), .Z(n8064) );
  XNOR U9313 ( .A(n8063), .B(n8064), .Z(n8068) );
  XOR U9314 ( .A(n8067), .B(sreg[1517]), .Z(n8060) );
  XNOR U9315 ( .A(n8068), .B(n8060), .Z(c[1517]) );
  NAND U9316 ( .A(n8062), .B(n8061), .Z(n8066) );
  NANDN U9317 ( .A(n8064), .B(n8063), .Z(n8065) );
  NAND U9318 ( .A(n8066), .B(n8065), .Z(n8072) );
  NAND U9319 ( .A(b[0]), .B(a[496]), .Z(n8071) );
  NAND U9320 ( .A(a[495]), .B(b[1]), .Z(n8070) );
  XNOR U9321 ( .A(n8071), .B(n8070), .Z(n8073) );
  XNOR U9322 ( .A(n8072), .B(n8073), .Z(n8077) );
  XOR U9323 ( .A(n8076), .B(sreg[1518]), .Z(n8069) );
  XNOR U9324 ( .A(n8077), .B(n8069), .Z(c[1518]) );
  NAND U9325 ( .A(n8071), .B(n8070), .Z(n8075) );
  NANDN U9326 ( .A(n8073), .B(n8072), .Z(n8074) );
  NAND U9327 ( .A(n8075), .B(n8074), .Z(n8081) );
  NAND U9328 ( .A(b[0]), .B(a[497]), .Z(n8080) );
  NAND U9329 ( .A(a[496]), .B(b[1]), .Z(n8079) );
  XNOR U9330 ( .A(n8080), .B(n8079), .Z(n8082) );
  XNOR U9331 ( .A(n8081), .B(n8082), .Z(n8086) );
  XOR U9332 ( .A(n8085), .B(sreg[1519]), .Z(n8078) );
  XNOR U9333 ( .A(n8086), .B(n8078), .Z(c[1519]) );
  NAND U9334 ( .A(n8080), .B(n8079), .Z(n8084) );
  NANDN U9335 ( .A(n8082), .B(n8081), .Z(n8083) );
  NAND U9336 ( .A(n8084), .B(n8083), .Z(n8091) );
  ANDN U9337 ( .B(a[498]), .A(n3951), .Z(n8089) );
  AND U9338 ( .A(b[1]), .B(a[497]), .Z(n8088) );
  XOR U9339 ( .A(n8089), .B(n8088), .Z(n8090) );
  XNOR U9340 ( .A(n8091), .B(n8090), .Z(n8093) );
  XOR U9341 ( .A(sreg[1520]), .B(n8092), .Z(n8087) );
  XNOR U9342 ( .A(n8093), .B(n8087), .Z(c[1520]) );
  NAND U9343 ( .A(b[0]), .B(a[499]), .Z(n8096) );
  NAND U9344 ( .A(a[498]), .B(b[1]), .Z(n8095) );
  XNOR U9345 ( .A(n8096), .B(n8095), .Z(n8098) );
  XNOR U9346 ( .A(n8097), .B(n8098), .Z(n8102) );
  XOR U9347 ( .A(n8101), .B(sreg[1521]), .Z(n8094) );
  XNOR U9348 ( .A(n8102), .B(n8094), .Z(c[1521]) );
  NAND U9349 ( .A(n8096), .B(n8095), .Z(n8100) );
  NANDN U9350 ( .A(n8098), .B(n8097), .Z(n8099) );
  NAND U9351 ( .A(n8100), .B(n8099), .Z(n8107) );
  ANDN U9352 ( .B(a[500]), .A(n3951), .Z(n8105) );
  AND U9353 ( .A(b[1]), .B(a[499]), .Z(n8104) );
  XOR U9354 ( .A(n8105), .B(n8104), .Z(n8106) );
  XNOR U9355 ( .A(n8107), .B(n8106), .Z(n8109) );
  XOR U9356 ( .A(sreg[1522]), .B(n8108), .Z(n8103) );
  XNOR U9357 ( .A(n8109), .B(n8103), .Z(c[1522]) );
  NAND U9358 ( .A(b[0]), .B(a[501]), .Z(n8112) );
  NAND U9359 ( .A(a[500]), .B(b[1]), .Z(n8111) );
  XNOR U9360 ( .A(n8112), .B(n8111), .Z(n8114) );
  XNOR U9361 ( .A(n8113), .B(n8114), .Z(n8118) );
  XOR U9362 ( .A(n8117), .B(sreg[1523]), .Z(n8110) );
  XNOR U9363 ( .A(n8118), .B(n8110), .Z(c[1523]) );
  NAND U9364 ( .A(n8112), .B(n8111), .Z(n8116) );
  NANDN U9365 ( .A(n8114), .B(n8113), .Z(n8115) );
  NAND U9366 ( .A(n8116), .B(n8115), .Z(n8123) );
  ANDN U9367 ( .B(a[502]), .A(n3951), .Z(n8121) );
  AND U9368 ( .A(b[1]), .B(a[501]), .Z(n8120) );
  XOR U9369 ( .A(n8121), .B(n8120), .Z(n8122) );
  XNOR U9370 ( .A(n8123), .B(n8122), .Z(n8125) );
  XOR U9371 ( .A(sreg[1524]), .B(n8124), .Z(n8119) );
  XNOR U9372 ( .A(n8125), .B(n8119), .Z(c[1524]) );
  NAND U9373 ( .A(b[0]), .B(a[503]), .Z(n8128) );
  NAND U9374 ( .A(a[502]), .B(b[1]), .Z(n8127) );
  XNOR U9375 ( .A(n8128), .B(n8127), .Z(n8130) );
  XNOR U9376 ( .A(n8129), .B(n8130), .Z(n8134) );
  XOR U9377 ( .A(n8133), .B(sreg[1525]), .Z(n8126) );
  XNOR U9378 ( .A(n8134), .B(n8126), .Z(c[1525]) );
  NAND U9379 ( .A(n8128), .B(n8127), .Z(n8132) );
  NANDN U9380 ( .A(n8130), .B(n8129), .Z(n8131) );
  NAND U9381 ( .A(n8132), .B(n8131), .Z(n8139) );
  ANDN U9382 ( .B(a[504]), .A(n3951), .Z(n8137) );
  AND U9383 ( .A(b[1]), .B(a[503]), .Z(n8136) );
  XOR U9384 ( .A(n8137), .B(n8136), .Z(n8138) );
  XNOR U9385 ( .A(n8139), .B(n8138), .Z(n8141) );
  XOR U9386 ( .A(sreg[1526]), .B(n8140), .Z(n8135) );
  XNOR U9387 ( .A(n8141), .B(n8135), .Z(c[1526]) );
  NAND U9388 ( .A(b[0]), .B(a[505]), .Z(n8144) );
  NAND U9389 ( .A(a[504]), .B(b[1]), .Z(n8143) );
  XNOR U9390 ( .A(n8144), .B(n8143), .Z(n8146) );
  XNOR U9391 ( .A(n8145), .B(n8146), .Z(n8150) );
  XOR U9392 ( .A(n8149), .B(sreg[1527]), .Z(n8142) );
  XNOR U9393 ( .A(n8150), .B(n8142), .Z(c[1527]) );
  NAND U9394 ( .A(n8144), .B(n8143), .Z(n8148) );
  NANDN U9395 ( .A(n8146), .B(n8145), .Z(n8147) );
  NAND U9396 ( .A(n8148), .B(n8147), .Z(n8155) );
  ANDN U9397 ( .B(a[506]), .A(n3951), .Z(n8153) );
  AND U9398 ( .A(b[1]), .B(a[505]), .Z(n8152) );
  XOR U9399 ( .A(n8153), .B(n8152), .Z(n8154) );
  XNOR U9400 ( .A(n8155), .B(n8154), .Z(n8157) );
  XOR U9401 ( .A(sreg[1528]), .B(n8156), .Z(n8151) );
  XNOR U9402 ( .A(n8157), .B(n8151), .Z(c[1528]) );
  NAND U9403 ( .A(b[0]), .B(a[507]), .Z(n8160) );
  NAND U9404 ( .A(a[506]), .B(b[1]), .Z(n8159) );
  XNOR U9405 ( .A(n8160), .B(n8159), .Z(n8162) );
  XNOR U9406 ( .A(n8161), .B(n8162), .Z(n8166) );
  XOR U9407 ( .A(n8165), .B(sreg[1529]), .Z(n8158) );
  XNOR U9408 ( .A(n8166), .B(n8158), .Z(c[1529]) );
  NAND U9409 ( .A(n8160), .B(n8159), .Z(n8164) );
  NANDN U9410 ( .A(n8162), .B(n8161), .Z(n8163) );
  NAND U9411 ( .A(n8164), .B(n8163), .Z(n8171) );
  ANDN U9412 ( .B(a[508]), .A(n3951), .Z(n8169) );
  AND U9413 ( .A(b[1]), .B(a[507]), .Z(n8168) );
  XOR U9414 ( .A(n8169), .B(n8168), .Z(n8170) );
  XNOR U9415 ( .A(n8171), .B(n8170), .Z(n8173) );
  XOR U9416 ( .A(sreg[1530]), .B(n8172), .Z(n8167) );
  XNOR U9417 ( .A(n8173), .B(n8167), .Z(c[1530]) );
  NAND U9418 ( .A(b[0]), .B(a[509]), .Z(n8176) );
  NAND U9419 ( .A(a[508]), .B(b[1]), .Z(n8175) );
  XNOR U9420 ( .A(n8176), .B(n8175), .Z(n8178) );
  XNOR U9421 ( .A(n8177), .B(n8178), .Z(n8182) );
  XOR U9422 ( .A(n8181), .B(sreg[1531]), .Z(n8174) );
  XNOR U9423 ( .A(n8182), .B(n8174), .Z(c[1531]) );
  NAND U9424 ( .A(n8176), .B(n8175), .Z(n8180) );
  NANDN U9425 ( .A(n8178), .B(n8177), .Z(n8179) );
  NAND U9426 ( .A(n8180), .B(n8179), .Z(n8187) );
  ANDN U9427 ( .B(a[510]), .A(n3952), .Z(n8185) );
  AND U9428 ( .A(b[1]), .B(a[509]), .Z(n8184) );
  XOR U9429 ( .A(n8185), .B(n8184), .Z(n8186) );
  XNOR U9430 ( .A(n8187), .B(n8186), .Z(n8192) );
  XOR U9431 ( .A(sreg[1532]), .B(n8191), .Z(n8183) );
  XNOR U9432 ( .A(n8192), .B(n8183), .Z(c[1532]) );
  OR U9433 ( .A(n8185), .B(n8184), .Z(n8190) );
  IV U9434 ( .A(n8186), .Z(n8188) );
  NANDN U9435 ( .A(n8188), .B(n8187), .Z(n8189) );
  NAND U9436 ( .A(n8190), .B(n8189), .Z(n8196) );
  NAND U9437 ( .A(b[0]), .B(a[511]), .Z(n8195) );
  NAND U9438 ( .A(a[510]), .B(b[1]), .Z(n8194) );
  XNOR U9439 ( .A(n8195), .B(n8194), .Z(n8197) );
  XNOR U9440 ( .A(n8196), .B(n8197), .Z(n8201) );
  XOR U9441 ( .A(n8200), .B(sreg[1533]), .Z(n8193) );
  XNOR U9442 ( .A(n8201), .B(n8193), .Z(c[1533]) );
  NAND U9443 ( .A(n8195), .B(n8194), .Z(n8199) );
  NANDN U9444 ( .A(n8197), .B(n8196), .Z(n8198) );
  NAND U9445 ( .A(n8199), .B(n8198), .Z(n8206) );
  ANDN U9446 ( .B(a[512]), .A(n3952), .Z(n8204) );
  AND U9447 ( .A(b[1]), .B(a[511]), .Z(n8203) );
  XOR U9448 ( .A(n8204), .B(n8203), .Z(n8205) );
  XNOR U9449 ( .A(n8206), .B(n8205), .Z(n8208) );
  XOR U9450 ( .A(sreg[1534]), .B(n8207), .Z(n8202) );
  XNOR U9451 ( .A(n8208), .B(n8202), .Z(c[1534]) );
  NAND U9452 ( .A(b[0]), .B(a[513]), .Z(n8211) );
  NAND U9453 ( .A(a[512]), .B(b[1]), .Z(n8210) );
  XNOR U9454 ( .A(n8211), .B(n8210), .Z(n8213) );
  XNOR U9455 ( .A(n8212), .B(n8213), .Z(n8217) );
  XOR U9456 ( .A(n8216), .B(sreg[1535]), .Z(n8209) );
  XNOR U9457 ( .A(n8217), .B(n8209), .Z(c[1535]) );
  NAND U9458 ( .A(n8211), .B(n8210), .Z(n8215) );
  NANDN U9459 ( .A(n8213), .B(n8212), .Z(n8214) );
  NAND U9460 ( .A(n8215), .B(n8214), .Z(n8222) );
  ANDN U9461 ( .B(a[514]), .A(n3952), .Z(n8220) );
  AND U9462 ( .A(b[1]), .B(a[513]), .Z(n8219) );
  XOR U9463 ( .A(n8220), .B(n8219), .Z(n8221) );
  XNOR U9464 ( .A(n8222), .B(n8221), .Z(n8224) );
  XOR U9465 ( .A(sreg[1536]), .B(n8223), .Z(n8218) );
  XNOR U9466 ( .A(n8224), .B(n8218), .Z(c[1536]) );
  NAND U9467 ( .A(b[0]), .B(a[515]), .Z(n8227) );
  NAND U9468 ( .A(a[514]), .B(b[1]), .Z(n8226) );
  XNOR U9469 ( .A(n8227), .B(n8226), .Z(n8229) );
  XNOR U9470 ( .A(n8228), .B(n8229), .Z(n8233) );
  XOR U9471 ( .A(n8232), .B(sreg[1537]), .Z(n8225) );
  XNOR U9472 ( .A(n8233), .B(n8225), .Z(c[1537]) );
  NAND U9473 ( .A(n8227), .B(n8226), .Z(n8231) );
  NANDN U9474 ( .A(n8229), .B(n8228), .Z(n8230) );
  NAND U9475 ( .A(n8231), .B(n8230), .Z(n8238) );
  ANDN U9476 ( .B(a[516]), .A(n3952), .Z(n8236) );
  AND U9477 ( .A(b[1]), .B(a[515]), .Z(n8235) );
  XOR U9478 ( .A(n8236), .B(n8235), .Z(n8237) );
  XNOR U9479 ( .A(n8238), .B(n8237), .Z(n8240) );
  XOR U9480 ( .A(sreg[1538]), .B(n8239), .Z(n8234) );
  XNOR U9481 ( .A(n8240), .B(n8234), .Z(c[1538]) );
  NAND U9482 ( .A(b[0]), .B(a[517]), .Z(n8243) );
  NAND U9483 ( .A(a[516]), .B(b[1]), .Z(n8242) );
  XNOR U9484 ( .A(n8243), .B(n8242), .Z(n8245) );
  XNOR U9485 ( .A(n8244), .B(n8245), .Z(n8249) );
  XOR U9486 ( .A(n8248), .B(sreg[1539]), .Z(n8241) );
  XNOR U9487 ( .A(n8249), .B(n8241), .Z(c[1539]) );
  NAND U9488 ( .A(n8243), .B(n8242), .Z(n8247) );
  NANDN U9489 ( .A(n8245), .B(n8244), .Z(n8246) );
  NAND U9490 ( .A(n8247), .B(n8246), .Z(n8254) );
  ANDN U9491 ( .B(a[518]), .A(n3952), .Z(n8252) );
  AND U9492 ( .A(b[1]), .B(a[517]), .Z(n8251) );
  XOR U9493 ( .A(n8252), .B(n8251), .Z(n8253) );
  XNOR U9494 ( .A(n8254), .B(n8253), .Z(n8256) );
  XOR U9495 ( .A(sreg[1540]), .B(n8255), .Z(n8250) );
  XNOR U9496 ( .A(n8256), .B(n8250), .Z(c[1540]) );
  ANDN U9497 ( .B(a[519]), .A(n3952), .Z(n8259) );
  AND U9498 ( .A(b[1]), .B(a[518]), .Z(n8258) );
  XOR U9499 ( .A(n8259), .B(n8258), .Z(n8260) );
  XNOR U9500 ( .A(n8261), .B(n8260), .Z(n8263) );
  XNOR U9501 ( .A(sreg[1541]), .B(n8262), .Z(n8257) );
  XNOR U9502 ( .A(n8263), .B(n8257), .Z(c[1541]) );
  ANDN U9503 ( .B(a[520]), .A(n3952), .Z(n8266) );
  AND U9504 ( .A(b[1]), .B(a[519]), .Z(n8265) );
  XOR U9505 ( .A(n8266), .B(n8265), .Z(n8267) );
  XNOR U9506 ( .A(n8268), .B(n8267), .Z(n8270) );
  XNOR U9507 ( .A(sreg[1542]), .B(n8269), .Z(n8264) );
  XNOR U9508 ( .A(n8270), .B(n8264), .Z(c[1542]) );
  NAND U9509 ( .A(b[0]), .B(a[521]), .Z(n8273) );
  NAND U9510 ( .A(a[520]), .B(b[1]), .Z(n8272) );
  XNOR U9511 ( .A(n8273), .B(n8272), .Z(n8275) );
  XNOR U9512 ( .A(n8274), .B(n8275), .Z(n8279) );
  XOR U9513 ( .A(n8278), .B(sreg[1543]), .Z(n8271) );
  XNOR U9514 ( .A(n8279), .B(n8271), .Z(c[1543]) );
  NAND U9515 ( .A(n8273), .B(n8272), .Z(n8277) );
  NANDN U9516 ( .A(n8275), .B(n8274), .Z(n8276) );
  NAND U9517 ( .A(n8277), .B(n8276), .Z(n8284) );
  ANDN U9518 ( .B(a[522]), .A(n3953), .Z(n8282) );
  AND U9519 ( .A(b[1]), .B(a[521]), .Z(n8281) );
  XOR U9520 ( .A(n8282), .B(n8281), .Z(n8283) );
  XNOR U9521 ( .A(n8284), .B(n8283), .Z(n8289) );
  XOR U9522 ( .A(sreg[1544]), .B(n8288), .Z(n8280) );
  XNOR U9523 ( .A(n8289), .B(n8280), .Z(c[1544]) );
  OR U9524 ( .A(n8282), .B(n8281), .Z(n8287) );
  IV U9525 ( .A(n8283), .Z(n8285) );
  NANDN U9526 ( .A(n8285), .B(n8284), .Z(n8286) );
  NAND U9527 ( .A(n8287), .B(n8286), .Z(n8293) );
  NAND U9528 ( .A(b[0]), .B(a[523]), .Z(n8292) );
  NAND U9529 ( .A(a[522]), .B(b[1]), .Z(n8291) );
  XNOR U9530 ( .A(n8292), .B(n8291), .Z(n8294) );
  XNOR U9531 ( .A(n8293), .B(n8294), .Z(n8298) );
  XOR U9532 ( .A(n8297), .B(sreg[1545]), .Z(n8290) );
  XNOR U9533 ( .A(n8298), .B(n8290), .Z(c[1545]) );
  NAND U9534 ( .A(n8292), .B(n8291), .Z(n8296) );
  NANDN U9535 ( .A(n8294), .B(n8293), .Z(n8295) );
  NAND U9536 ( .A(n8296), .B(n8295), .Z(n8303) );
  ANDN U9537 ( .B(a[524]), .A(n3953), .Z(n8301) );
  AND U9538 ( .A(b[1]), .B(a[523]), .Z(n8300) );
  XOR U9539 ( .A(n8301), .B(n8300), .Z(n8302) );
  XNOR U9540 ( .A(n8303), .B(n8302), .Z(n8305) );
  XOR U9541 ( .A(sreg[1546]), .B(n8304), .Z(n8299) );
  XNOR U9542 ( .A(n8305), .B(n8299), .Z(c[1546]) );
  NAND U9543 ( .A(b[0]), .B(a[525]), .Z(n8308) );
  NAND U9544 ( .A(a[524]), .B(b[1]), .Z(n8307) );
  XNOR U9545 ( .A(n8308), .B(n8307), .Z(n8310) );
  XNOR U9546 ( .A(n8309), .B(n8310), .Z(n8314) );
  XOR U9547 ( .A(n8313), .B(sreg[1547]), .Z(n8306) );
  XNOR U9548 ( .A(n8314), .B(n8306), .Z(c[1547]) );
  NAND U9549 ( .A(n8308), .B(n8307), .Z(n8312) );
  NANDN U9550 ( .A(n8310), .B(n8309), .Z(n8311) );
  NAND U9551 ( .A(n8312), .B(n8311), .Z(n8319) );
  ANDN U9552 ( .B(a[526]), .A(n3953), .Z(n8317) );
  AND U9553 ( .A(b[1]), .B(a[525]), .Z(n8316) );
  XOR U9554 ( .A(n8317), .B(n8316), .Z(n8318) );
  XNOR U9555 ( .A(n8319), .B(n8318), .Z(n8321) );
  XOR U9556 ( .A(sreg[1548]), .B(n8320), .Z(n8315) );
  XNOR U9557 ( .A(n8321), .B(n8315), .Z(c[1548]) );
  NAND U9558 ( .A(b[0]), .B(a[527]), .Z(n8324) );
  NAND U9559 ( .A(a[526]), .B(b[1]), .Z(n8323) );
  XNOR U9560 ( .A(n8324), .B(n8323), .Z(n8326) );
  XNOR U9561 ( .A(n8325), .B(n8326), .Z(n8330) );
  XOR U9562 ( .A(n8329), .B(sreg[1549]), .Z(n8322) );
  XNOR U9563 ( .A(n8330), .B(n8322), .Z(c[1549]) );
  NAND U9564 ( .A(n8324), .B(n8323), .Z(n8328) );
  NANDN U9565 ( .A(n8326), .B(n8325), .Z(n8327) );
  NAND U9566 ( .A(n8328), .B(n8327), .Z(n8335) );
  ANDN U9567 ( .B(a[528]), .A(n3953), .Z(n8333) );
  AND U9568 ( .A(b[1]), .B(a[527]), .Z(n8332) );
  XOR U9569 ( .A(n8333), .B(n8332), .Z(n8334) );
  XNOR U9570 ( .A(n8335), .B(n8334), .Z(n8337) );
  XOR U9571 ( .A(sreg[1550]), .B(n8336), .Z(n8331) );
  XNOR U9572 ( .A(n8337), .B(n8331), .Z(c[1550]) );
  NAND U9573 ( .A(b[0]), .B(a[529]), .Z(n8340) );
  NAND U9574 ( .A(a[528]), .B(b[1]), .Z(n8339) );
  XNOR U9575 ( .A(n8340), .B(n8339), .Z(n8342) );
  XNOR U9576 ( .A(n8341), .B(n8342), .Z(n8346) );
  XOR U9577 ( .A(n8345), .B(sreg[1551]), .Z(n8338) );
  XNOR U9578 ( .A(n8346), .B(n8338), .Z(c[1551]) );
  NAND U9579 ( .A(n8340), .B(n8339), .Z(n8344) );
  NANDN U9580 ( .A(n8342), .B(n8341), .Z(n8343) );
  NAND U9581 ( .A(n8344), .B(n8343), .Z(n8351) );
  ANDN U9582 ( .B(a[530]), .A(n3953), .Z(n8349) );
  AND U9583 ( .A(b[1]), .B(a[529]), .Z(n8348) );
  XOR U9584 ( .A(n8349), .B(n8348), .Z(n8350) );
  XNOR U9585 ( .A(n8351), .B(n8350), .Z(n8353) );
  XOR U9586 ( .A(sreg[1552]), .B(n8352), .Z(n8347) );
  XNOR U9587 ( .A(n8353), .B(n8347), .Z(c[1552]) );
  NAND U9588 ( .A(b[0]), .B(a[531]), .Z(n8356) );
  NAND U9589 ( .A(a[530]), .B(b[1]), .Z(n8355) );
  XNOR U9590 ( .A(n8356), .B(n8355), .Z(n8358) );
  XNOR U9591 ( .A(n8357), .B(n8358), .Z(n8362) );
  XOR U9592 ( .A(n8361), .B(sreg[1553]), .Z(n8354) );
  XNOR U9593 ( .A(n8362), .B(n8354), .Z(c[1553]) );
  NAND U9594 ( .A(n8356), .B(n8355), .Z(n8360) );
  NANDN U9595 ( .A(n8358), .B(n8357), .Z(n8359) );
  NAND U9596 ( .A(n8360), .B(n8359), .Z(n8367) );
  ANDN U9597 ( .B(a[532]), .A(n3953), .Z(n8365) );
  AND U9598 ( .A(b[1]), .B(a[531]), .Z(n8364) );
  XOR U9599 ( .A(n8365), .B(n8364), .Z(n8366) );
  XNOR U9600 ( .A(n8367), .B(n8366), .Z(n8369) );
  XOR U9601 ( .A(sreg[1554]), .B(n8368), .Z(n8363) );
  XNOR U9602 ( .A(n8369), .B(n8363), .Z(c[1554]) );
  NAND U9603 ( .A(b[0]), .B(a[533]), .Z(n8372) );
  NAND U9604 ( .A(a[532]), .B(b[1]), .Z(n8371) );
  XNOR U9605 ( .A(n8372), .B(n8371), .Z(n8374) );
  XNOR U9606 ( .A(n8373), .B(n8374), .Z(n8378) );
  XOR U9607 ( .A(n8377), .B(sreg[1555]), .Z(n8370) );
  XNOR U9608 ( .A(n8378), .B(n8370), .Z(c[1555]) );
  NAND U9609 ( .A(n8372), .B(n8371), .Z(n8376) );
  NANDN U9610 ( .A(n8374), .B(n8373), .Z(n8375) );
  NAND U9611 ( .A(n8376), .B(n8375), .Z(n8383) );
  ANDN U9612 ( .B(a[534]), .A(n3953), .Z(n8381) );
  AND U9613 ( .A(b[1]), .B(a[533]), .Z(n8380) );
  XOR U9614 ( .A(n8381), .B(n8380), .Z(n8382) );
  XNOR U9615 ( .A(n8383), .B(n8382), .Z(n8385) );
  XOR U9616 ( .A(sreg[1556]), .B(n8384), .Z(n8379) );
  XNOR U9617 ( .A(n8385), .B(n8379), .Z(c[1556]) );
  NAND U9618 ( .A(b[0]), .B(a[535]), .Z(n8388) );
  NAND U9619 ( .A(a[534]), .B(b[1]), .Z(n8387) );
  XNOR U9620 ( .A(n8388), .B(n8387), .Z(n8390) );
  XNOR U9621 ( .A(n8389), .B(n8390), .Z(n8394) );
  XOR U9622 ( .A(n8393), .B(sreg[1557]), .Z(n8386) );
  XNOR U9623 ( .A(n8394), .B(n8386), .Z(c[1557]) );
  NAND U9624 ( .A(n8388), .B(n8387), .Z(n8392) );
  NANDN U9625 ( .A(n8390), .B(n8389), .Z(n8391) );
  NAND U9626 ( .A(n8392), .B(n8391), .Z(n8399) );
  ANDN U9627 ( .B(a[536]), .A(n3954), .Z(n8397) );
  AND U9628 ( .A(b[1]), .B(a[535]), .Z(n8396) );
  XOR U9629 ( .A(n8397), .B(n8396), .Z(n8398) );
  XNOR U9630 ( .A(n8399), .B(n8398), .Z(n8404) );
  XOR U9631 ( .A(sreg[1558]), .B(n8403), .Z(n8395) );
  XNOR U9632 ( .A(n8404), .B(n8395), .Z(c[1558]) );
  OR U9633 ( .A(n8397), .B(n8396), .Z(n8402) );
  IV U9634 ( .A(n8398), .Z(n8400) );
  NANDN U9635 ( .A(n8400), .B(n8399), .Z(n8401) );
  NAND U9636 ( .A(n8402), .B(n8401), .Z(n8408) );
  NAND U9637 ( .A(b[0]), .B(a[537]), .Z(n8407) );
  NAND U9638 ( .A(a[536]), .B(b[1]), .Z(n8406) );
  XNOR U9639 ( .A(n8407), .B(n8406), .Z(n8409) );
  XNOR U9640 ( .A(n8408), .B(n8409), .Z(n8413) );
  XOR U9641 ( .A(n8412), .B(sreg[1559]), .Z(n8405) );
  XNOR U9642 ( .A(n8413), .B(n8405), .Z(c[1559]) );
  NAND U9643 ( .A(n8407), .B(n8406), .Z(n8411) );
  NANDN U9644 ( .A(n8409), .B(n8408), .Z(n8410) );
  NAND U9645 ( .A(n8411), .B(n8410), .Z(n8418) );
  ANDN U9646 ( .B(a[538]), .A(n3954), .Z(n8416) );
  AND U9647 ( .A(b[1]), .B(a[537]), .Z(n8415) );
  XOR U9648 ( .A(n8416), .B(n8415), .Z(n8417) );
  XNOR U9649 ( .A(n8418), .B(n8417), .Z(n8420) );
  XOR U9650 ( .A(sreg[1560]), .B(n8419), .Z(n8414) );
  XNOR U9651 ( .A(n8420), .B(n8414), .Z(c[1560]) );
  ANDN U9652 ( .B(a[539]), .A(n3954), .Z(n8423) );
  AND U9653 ( .A(b[1]), .B(a[538]), .Z(n8422) );
  XOR U9654 ( .A(n8423), .B(n8422), .Z(n8424) );
  XNOR U9655 ( .A(n8425), .B(n8424), .Z(n8427) );
  XNOR U9656 ( .A(sreg[1561]), .B(n8426), .Z(n8421) );
  XNOR U9657 ( .A(n8427), .B(n8421), .Z(c[1561]) );
  ANDN U9658 ( .B(a[540]), .A(n3954), .Z(n8430) );
  AND U9659 ( .A(b[1]), .B(a[539]), .Z(n8429) );
  XOR U9660 ( .A(n8430), .B(n8429), .Z(n8431) );
  XNOR U9661 ( .A(n8432), .B(n8431), .Z(n8434) );
  XNOR U9662 ( .A(sreg[1562]), .B(n8433), .Z(n8428) );
  XNOR U9663 ( .A(n8434), .B(n8428), .Z(c[1562]) );
  NAND U9664 ( .A(b[0]), .B(a[541]), .Z(n8437) );
  NAND U9665 ( .A(a[540]), .B(b[1]), .Z(n8436) );
  XNOR U9666 ( .A(n8437), .B(n8436), .Z(n8439) );
  XNOR U9667 ( .A(n8438), .B(n8439), .Z(n8443) );
  XOR U9668 ( .A(n8442), .B(sreg[1563]), .Z(n8435) );
  XNOR U9669 ( .A(n8443), .B(n8435), .Z(c[1563]) );
  NAND U9670 ( .A(n8437), .B(n8436), .Z(n8441) );
  NANDN U9671 ( .A(n8439), .B(n8438), .Z(n8440) );
  NAND U9672 ( .A(n8441), .B(n8440), .Z(n8448) );
  ANDN U9673 ( .B(a[542]), .A(n3954), .Z(n8446) );
  AND U9674 ( .A(b[1]), .B(a[541]), .Z(n8445) );
  XOR U9675 ( .A(n8446), .B(n8445), .Z(n8447) );
  XNOR U9676 ( .A(n8448), .B(n8447), .Z(n8450) );
  XOR U9677 ( .A(sreg[1564]), .B(n8449), .Z(n8444) );
  XNOR U9678 ( .A(n8450), .B(n8444), .Z(c[1564]) );
  NAND U9679 ( .A(b[0]), .B(a[543]), .Z(n8453) );
  NAND U9680 ( .A(a[542]), .B(b[1]), .Z(n8452) );
  XNOR U9681 ( .A(n8453), .B(n8452), .Z(n8455) );
  XNOR U9682 ( .A(n8454), .B(n8455), .Z(n8459) );
  XOR U9683 ( .A(n8458), .B(sreg[1565]), .Z(n8451) );
  XNOR U9684 ( .A(n8459), .B(n8451), .Z(c[1565]) );
  NAND U9685 ( .A(n8453), .B(n8452), .Z(n8457) );
  NANDN U9686 ( .A(n8455), .B(n8454), .Z(n8456) );
  NAND U9687 ( .A(n8457), .B(n8456), .Z(n8464) );
  ANDN U9688 ( .B(a[544]), .A(n3954), .Z(n8462) );
  AND U9689 ( .A(b[1]), .B(a[543]), .Z(n8461) );
  XOR U9690 ( .A(n8462), .B(n8461), .Z(n8463) );
  XNOR U9691 ( .A(n8464), .B(n8463), .Z(n8466) );
  XOR U9692 ( .A(sreg[1566]), .B(n8465), .Z(n8460) );
  XNOR U9693 ( .A(n8466), .B(n8460), .Z(c[1566]) );
  NAND U9694 ( .A(b[0]), .B(a[545]), .Z(n8469) );
  NAND U9695 ( .A(a[544]), .B(b[1]), .Z(n8468) );
  XNOR U9696 ( .A(n8469), .B(n8468), .Z(n8471) );
  XNOR U9697 ( .A(n8470), .B(n8471), .Z(n8475) );
  XOR U9698 ( .A(n8474), .B(sreg[1567]), .Z(n8467) );
  XNOR U9699 ( .A(n8475), .B(n8467), .Z(c[1567]) );
  NAND U9700 ( .A(n8469), .B(n8468), .Z(n8473) );
  NANDN U9701 ( .A(n8471), .B(n8470), .Z(n8472) );
  NAND U9702 ( .A(n8473), .B(n8472), .Z(n8480) );
  ANDN U9703 ( .B(a[546]), .A(n3954), .Z(n8478) );
  AND U9704 ( .A(b[1]), .B(a[545]), .Z(n8477) );
  XOR U9705 ( .A(n8478), .B(n8477), .Z(n8479) );
  XNOR U9706 ( .A(n8480), .B(n8479), .Z(n8482) );
  XOR U9707 ( .A(sreg[1568]), .B(n8481), .Z(n8476) );
  XNOR U9708 ( .A(n8482), .B(n8476), .Z(c[1568]) );
  NAND U9709 ( .A(b[0]), .B(a[547]), .Z(n8485) );
  NAND U9710 ( .A(a[546]), .B(b[1]), .Z(n8484) );
  XNOR U9711 ( .A(n8485), .B(n8484), .Z(n8487) );
  XNOR U9712 ( .A(n8486), .B(n8487), .Z(n8491) );
  XOR U9713 ( .A(n8490), .B(sreg[1569]), .Z(n8483) );
  XNOR U9714 ( .A(n8491), .B(n8483), .Z(c[1569]) );
  NAND U9715 ( .A(n8485), .B(n8484), .Z(n8489) );
  NANDN U9716 ( .A(n8487), .B(n8486), .Z(n8488) );
  NAND U9717 ( .A(n8489), .B(n8488), .Z(n8496) );
  ANDN U9718 ( .B(a[548]), .A(n3955), .Z(n8494) );
  AND U9719 ( .A(b[1]), .B(a[547]), .Z(n8493) );
  XOR U9720 ( .A(n8494), .B(n8493), .Z(n8495) );
  XNOR U9721 ( .A(n8496), .B(n8495), .Z(n8501) );
  XOR U9722 ( .A(sreg[1570]), .B(n8500), .Z(n8492) );
  XNOR U9723 ( .A(n8501), .B(n8492), .Z(c[1570]) );
  OR U9724 ( .A(n8494), .B(n8493), .Z(n8499) );
  IV U9725 ( .A(n8495), .Z(n8497) );
  NANDN U9726 ( .A(n8497), .B(n8496), .Z(n8498) );
  NAND U9727 ( .A(n8499), .B(n8498), .Z(n8505) );
  NAND U9728 ( .A(b[0]), .B(a[549]), .Z(n8504) );
  NAND U9729 ( .A(a[548]), .B(b[1]), .Z(n8503) );
  XNOR U9730 ( .A(n8504), .B(n8503), .Z(n8506) );
  XNOR U9731 ( .A(n8505), .B(n8506), .Z(n8510) );
  XOR U9732 ( .A(n8509), .B(sreg[1571]), .Z(n8502) );
  XNOR U9733 ( .A(n8510), .B(n8502), .Z(c[1571]) );
  NAND U9734 ( .A(n8504), .B(n8503), .Z(n8508) );
  NANDN U9735 ( .A(n8506), .B(n8505), .Z(n8507) );
  NAND U9736 ( .A(n8508), .B(n8507), .Z(n8514) );
  NAND U9737 ( .A(b[0]), .B(a[550]), .Z(n8513) );
  NAND U9738 ( .A(a[549]), .B(b[1]), .Z(n8512) );
  XNOR U9739 ( .A(n8513), .B(n8512), .Z(n8515) );
  XNOR U9740 ( .A(n8514), .B(n8515), .Z(n8519) );
  XOR U9741 ( .A(n8518), .B(sreg[1572]), .Z(n8511) );
  XNOR U9742 ( .A(n8519), .B(n8511), .Z(c[1572]) );
  NAND U9743 ( .A(n8513), .B(n8512), .Z(n8517) );
  NANDN U9744 ( .A(n8515), .B(n8514), .Z(n8516) );
  NAND U9745 ( .A(n8517), .B(n8516), .Z(n8523) );
  NAND U9746 ( .A(b[0]), .B(a[551]), .Z(n8522) );
  NAND U9747 ( .A(a[550]), .B(b[1]), .Z(n8521) );
  XNOR U9748 ( .A(n8522), .B(n8521), .Z(n8524) );
  XNOR U9749 ( .A(n8523), .B(n8524), .Z(n8528) );
  XOR U9750 ( .A(n8527), .B(sreg[1573]), .Z(n8520) );
  XNOR U9751 ( .A(n8528), .B(n8520), .Z(c[1573]) );
  NAND U9752 ( .A(n8522), .B(n8521), .Z(n8526) );
  NANDN U9753 ( .A(n8524), .B(n8523), .Z(n8525) );
  NAND U9754 ( .A(n8526), .B(n8525), .Z(n8532) );
  NAND U9755 ( .A(b[0]), .B(a[552]), .Z(n8531) );
  NAND U9756 ( .A(a[551]), .B(b[1]), .Z(n8530) );
  XNOR U9757 ( .A(n8531), .B(n8530), .Z(n8533) );
  XNOR U9758 ( .A(n8532), .B(n8533), .Z(n8537) );
  XOR U9759 ( .A(n8536), .B(sreg[1574]), .Z(n8529) );
  XNOR U9760 ( .A(n8537), .B(n8529), .Z(c[1574]) );
  NAND U9761 ( .A(n8531), .B(n8530), .Z(n8535) );
  NANDN U9762 ( .A(n8533), .B(n8532), .Z(n8534) );
  NAND U9763 ( .A(n8535), .B(n8534), .Z(n8541) );
  NAND U9764 ( .A(b[0]), .B(a[553]), .Z(n8540) );
  NAND U9765 ( .A(a[552]), .B(b[1]), .Z(n8539) );
  XNOR U9766 ( .A(n8540), .B(n8539), .Z(n8542) );
  XNOR U9767 ( .A(n8541), .B(n8542), .Z(n8546) );
  XOR U9768 ( .A(n8545), .B(sreg[1575]), .Z(n8538) );
  XNOR U9769 ( .A(n8546), .B(n8538), .Z(c[1575]) );
  NAND U9770 ( .A(n8540), .B(n8539), .Z(n8544) );
  NANDN U9771 ( .A(n8542), .B(n8541), .Z(n8543) );
  NAND U9772 ( .A(n8544), .B(n8543), .Z(n8551) );
  ANDN U9773 ( .B(a[554]), .A(n3955), .Z(n8549) );
  AND U9774 ( .A(b[1]), .B(a[553]), .Z(n8548) );
  XOR U9775 ( .A(n8549), .B(n8548), .Z(n8550) );
  XNOR U9776 ( .A(n8551), .B(n8550), .Z(n8553) );
  XOR U9777 ( .A(sreg[1576]), .B(n8552), .Z(n8547) );
  XNOR U9778 ( .A(n8553), .B(n8547), .Z(c[1576]) );
  NAND U9779 ( .A(b[0]), .B(a[555]), .Z(n8556) );
  NAND U9780 ( .A(a[554]), .B(b[1]), .Z(n8555) );
  XNOR U9781 ( .A(n8556), .B(n8555), .Z(n8558) );
  XNOR U9782 ( .A(n8557), .B(n8558), .Z(n8562) );
  XOR U9783 ( .A(n8561), .B(sreg[1577]), .Z(n8554) );
  XNOR U9784 ( .A(n8562), .B(n8554), .Z(c[1577]) );
  NAND U9785 ( .A(n8556), .B(n8555), .Z(n8560) );
  NANDN U9786 ( .A(n8558), .B(n8557), .Z(n8559) );
  NAND U9787 ( .A(n8560), .B(n8559), .Z(n8566) );
  NAND U9788 ( .A(b[0]), .B(a[556]), .Z(n8565) );
  NAND U9789 ( .A(a[555]), .B(b[1]), .Z(n8564) );
  XNOR U9790 ( .A(n8565), .B(n8564), .Z(n8567) );
  XNOR U9791 ( .A(n8566), .B(n8567), .Z(n8571) );
  XOR U9792 ( .A(n8570), .B(sreg[1578]), .Z(n8563) );
  XNOR U9793 ( .A(n8571), .B(n8563), .Z(c[1578]) );
  NAND U9794 ( .A(n8565), .B(n8564), .Z(n8569) );
  NANDN U9795 ( .A(n8567), .B(n8566), .Z(n8568) );
  NAND U9796 ( .A(n8569), .B(n8568), .Z(n8575) );
  NAND U9797 ( .A(b[0]), .B(a[557]), .Z(n8574) );
  NAND U9798 ( .A(a[556]), .B(b[1]), .Z(n8573) );
  XNOR U9799 ( .A(n8574), .B(n8573), .Z(n8576) );
  XNOR U9800 ( .A(n8575), .B(n8576), .Z(n8580) );
  XOR U9801 ( .A(n8579), .B(sreg[1579]), .Z(n8572) );
  XNOR U9802 ( .A(n8580), .B(n8572), .Z(c[1579]) );
  NAND U9803 ( .A(n8574), .B(n8573), .Z(n8578) );
  NANDN U9804 ( .A(n8576), .B(n8575), .Z(n8577) );
  NAND U9805 ( .A(n8578), .B(n8577), .Z(n8585) );
  ANDN U9806 ( .B(a[558]), .A(n3955), .Z(n8583) );
  AND U9807 ( .A(b[1]), .B(a[557]), .Z(n8582) );
  XOR U9808 ( .A(n8583), .B(n8582), .Z(n8584) );
  XNOR U9809 ( .A(n8585), .B(n8584), .Z(n8587) );
  XOR U9810 ( .A(sreg[1580]), .B(n8586), .Z(n8581) );
  XNOR U9811 ( .A(n8587), .B(n8581), .Z(c[1580]) );
  NAND U9812 ( .A(b[0]), .B(a[559]), .Z(n8590) );
  NAND U9813 ( .A(a[558]), .B(b[1]), .Z(n8589) );
  XNOR U9814 ( .A(n8590), .B(n8589), .Z(n8592) );
  XNOR U9815 ( .A(n8591), .B(n8592), .Z(n8596) );
  XOR U9816 ( .A(n8595), .B(sreg[1581]), .Z(n8588) );
  XNOR U9817 ( .A(n8596), .B(n8588), .Z(c[1581]) );
  NAND U9818 ( .A(n8590), .B(n8589), .Z(n8594) );
  NANDN U9819 ( .A(n8592), .B(n8591), .Z(n8593) );
  NAND U9820 ( .A(n8594), .B(n8593), .Z(n8601) );
  ANDN U9821 ( .B(a[560]), .A(n3955), .Z(n8599) );
  AND U9822 ( .A(b[1]), .B(a[559]), .Z(n8598) );
  XOR U9823 ( .A(n8599), .B(n8598), .Z(n8600) );
  XNOR U9824 ( .A(n8601), .B(n8600), .Z(n8603) );
  XOR U9825 ( .A(sreg[1582]), .B(n8602), .Z(n8597) );
  XNOR U9826 ( .A(n8603), .B(n8597), .Z(c[1582]) );
  NAND U9827 ( .A(b[0]), .B(a[561]), .Z(n8606) );
  NAND U9828 ( .A(a[560]), .B(b[1]), .Z(n8605) );
  XNOR U9829 ( .A(n8606), .B(n8605), .Z(n8608) );
  XNOR U9830 ( .A(n8607), .B(n8608), .Z(n8612) );
  XOR U9831 ( .A(n8611), .B(sreg[1583]), .Z(n8604) );
  XNOR U9832 ( .A(n8612), .B(n8604), .Z(c[1583]) );
  NAND U9833 ( .A(n8606), .B(n8605), .Z(n8610) );
  NANDN U9834 ( .A(n8608), .B(n8607), .Z(n8609) );
  NAND U9835 ( .A(n8610), .B(n8609), .Z(n8617) );
  ANDN U9836 ( .B(a[562]), .A(n3955), .Z(n8615) );
  AND U9837 ( .A(b[1]), .B(a[561]), .Z(n8614) );
  XOR U9838 ( .A(n8615), .B(n8614), .Z(n8616) );
  XNOR U9839 ( .A(n8617), .B(n8616), .Z(n8619) );
  XOR U9840 ( .A(sreg[1584]), .B(n8618), .Z(n8613) );
  XNOR U9841 ( .A(n8619), .B(n8613), .Z(c[1584]) );
  NAND U9842 ( .A(b[0]), .B(a[563]), .Z(n8622) );
  NAND U9843 ( .A(a[562]), .B(b[1]), .Z(n8621) );
  XNOR U9844 ( .A(n8622), .B(n8621), .Z(n8624) );
  XNOR U9845 ( .A(n8623), .B(n8624), .Z(n8628) );
  XOR U9846 ( .A(n8627), .B(sreg[1585]), .Z(n8620) );
  XNOR U9847 ( .A(n8628), .B(n8620), .Z(c[1585]) );
  NAND U9848 ( .A(n8622), .B(n8621), .Z(n8626) );
  NANDN U9849 ( .A(n8624), .B(n8623), .Z(n8625) );
  NAND U9850 ( .A(n8626), .B(n8625), .Z(n8633) );
  ANDN U9851 ( .B(a[564]), .A(n3955), .Z(n8631) );
  AND U9852 ( .A(b[1]), .B(a[563]), .Z(n8630) );
  XOR U9853 ( .A(n8631), .B(n8630), .Z(n8632) );
  XNOR U9854 ( .A(n8633), .B(n8632), .Z(n8635) );
  XOR U9855 ( .A(sreg[1586]), .B(n8634), .Z(n8629) );
  XNOR U9856 ( .A(n8635), .B(n8629), .Z(c[1586]) );
  ANDN U9857 ( .B(a[565]), .A(n3955), .Z(n8638) );
  AND U9858 ( .A(b[1]), .B(a[564]), .Z(n8637) );
  XOR U9859 ( .A(n8638), .B(n8637), .Z(n8639) );
  XNOR U9860 ( .A(n8640), .B(n8639), .Z(n8642) );
  XNOR U9861 ( .A(sreg[1587]), .B(n8641), .Z(n8636) );
  XNOR U9862 ( .A(n8642), .B(n8636), .Z(c[1587]) );
  ANDN U9863 ( .B(a[566]), .A(n3956), .Z(n8645) );
  AND U9864 ( .A(b[1]), .B(a[565]), .Z(n8644) );
  XOR U9865 ( .A(n8645), .B(n8644), .Z(n8646) );
  XNOR U9866 ( .A(n8647), .B(n8646), .Z(n8652) );
  XNOR U9867 ( .A(sreg[1588]), .B(n8651), .Z(n8643) );
  XNOR U9868 ( .A(n8652), .B(n8643), .Z(c[1588]) );
  OR U9869 ( .A(n8645), .B(n8644), .Z(n8650) );
  IV U9870 ( .A(n8646), .Z(n8648) );
  NANDN U9871 ( .A(n8648), .B(n8647), .Z(n8649) );
  NAND U9872 ( .A(n8650), .B(n8649), .Z(n8656) );
  NAND U9873 ( .A(b[0]), .B(a[567]), .Z(n8655) );
  NAND U9874 ( .A(a[566]), .B(b[1]), .Z(n8654) );
  XNOR U9875 ( .A(n8655), .B(n8654), .Z(n8657) );
  XNOR U9876 ( .A(n8656), .B(n8657), .Z(n8661) );
  XOR U9877 ( .A(n8660), .B(sreg[1589]), .Z(n8653) );
  XNOR U9878 ( .A(n8661), .B(n8653), .Z(c[1589]) );
  NAND U9879 ( .A(n8655), .B(n8654), .Z(n8659) );
  NANDN U9880 ( .A(n8657), .B(n8656), .Z(n8658) );
  NAND U9881 ( .A(n8659), .B(n8658), .Z(n8666) );
  ANDN U9882 ( .B(a[568]), .A(n3956), .Z(n8664) );
  AND U9883 ( .A(b[1]), .B(a[567]), .Z(n8663) );
  XOR U9884 ( .A(n8664), .B(n8663), .Z(n8665) );
  XNOR U9885 ( .A(n8666), .B(n8665), .Z(n8668) );
  XOR U9886 ( .A(sreg[1590]), .B(n8667), .Z(n8662) );
  XNOR U9887 ( .A(n8668), .B(n8662), .Z(c[1590]) );
  NAND U9888 ( .A(b[0]), .B(a[569]), .Z(n8671) );
  NAND U9889 ( .A(a[568]), .B(b[1]), .Z(n8670) );
  XNOR U9890 ( .A(n8671), .B(n8670), .Z(n8673) );
  XNOR U9891 ( .A(n8672), .B(n8673), .Z(n8677) );
  XOR U9892 ( .A(n8676), .B(sreg[1591]), .Z(n8669) );
  XNOR U9893 ( .A(n8677), .B(n8669), .Z(c[1591]) );
  NAND U9894 ( .A(n8671), .B(n8670), .Z(n8675) );
  NANDN U9895 ( .A(n8673), .B(n8672), .Z(n8674) );
  NAND U9896 ( .A(n8675), .B(n8674), .Z(n8682) );
  ANDN U9897 ( .B(a[570]), .A(n3956), .Z(n8680) );
  AND U9898 ( .A(b[1]), .B(a[569]), .Z(n8679) );
  XOR U9899 ( .A(n8680), .B(n8679), .Z(n8681) );
  XNOR U9900 ( .A(n8682), .B(n8681), .Z(n8684) );
  XOR U9901 ( .A(sreg[1592]), .B(n8683), .Z(n8678) );
  XNOR U9902 ( .A(n8684), .B(n8678), .Z(c[1592]) );
  NAND U9903 ( .A(b[0]), .B(a[571]), .Z(n8687) );
  NAND U9904 ( .A(a[570]), .B(b[1]), .Z(n8686) );
  XNOR U9905 ( .A(n8687), .B(n8686), .Z(n8689) );
  XNOR U9906 ( .A(n8688), .B(n8689), .Z(n8693) );
  XOR U9907 ( .A(n8692), .B(sreg[1593]), .Z(n8685) );
  XNOR U9908 ( .A(n8693), .B(n8685), .Z(c[1593]) );
  NAND U9909 ( .A(n8687), .B(n8686), .Z(n8691) );
  NANDN U9910 ( .A(n8689), .B(n8688), .Z(n8690) );
  NAND U9911 ( .A(n8691), .B(n8690), .Z(n8698) );
  ANDN U9912 ( .B(a[572]), .A(n3956), .Z(n8696) );
  AND U9913 ( .A(b[1]), .B(a[571]), .Z(n8695) );
  XOR U9914 ( .A(n8696), .B(n8695), .Z(n8697) );
  XNOR U9915 ( .A(n8698), .B(n8697), .Z(n8700) );
  XOR U9916 ( .A(sreg[1594]), .B(n8699), .Z(n8694) );
  XNOR U9917 ( .A(n8700), .B(n8694), .Z(c[1594]) );
  NAND U9918 ( .A(b[0]), .B(a[573]), .Z(n8703) );
  NAND U9919 ( .A(a[572]), .B(b[1]), .Z(n8702) );
  XNOR U9920 ( .A(n8703), .B(n8702), .Z(n8705) );
  XNOR U9921 ( .A(n8704), .B(n8705), .Z(n8709) );
  XOR U9922 ( .A(n8708), .B(sreg[1595]), .Z(n8701) );
  XNOR U9923 ( .A(n8709), .B(n8701), .Z(c[1595]) );
  NAND U9924 ( .A(n8703), .B(n8702), .Z(n8707) );
  NANDN U9925 ( .A(n8705), .B(n8704), .Z(n8706) );
  NAND U9926 ( .A(n8707), .B(n8706), .Z(n8714) );
  ANDN U9927 ( .B(a[574]), .A(n3956), .Z(n8712) );
  AND U9928 ( .A(b[1]), .B(a[573]), .Z(n8711) );
  XOR U9929 ( .A(n8712), .B(n8711), .Z(n8713) );
  XNOR U9930 ( .A(n8714), .B(n8713), .Z(n8716) );
  XOR U9931 ( .A(sreg[1596]), .B(n8715), .Z(n8710) );
  XNOR U9932 ( .A(n8716), .B(n8710), .Z(c[1596]) );
  NAND U9933 ( .A(b[0]), .B(a[575]), .Z(n8719) );
  NAND U9934 ( .A(a[574]), .B(b[1]), .Z(n8718) );
  XNOR U9935 ( .A(n8719), .B(n8718), .Z(n8721) );
  XNOR U9936 ( .A(n8720), .B(n8721), .Z(n8725) );
  XOR U9937 ( .A(n8724), .B(sreg[1597]), .Z(n8717) );
  XNOR U9938 ( .A(n8725), .B(n8717), .Z(c[1597]) );
  NAND U9939 ( .A(n8719), .B(n8718), .Z(n8723) );
  NANDN U9940 ( .A(n8721), .B(n8720), .Z(n8722) );
  NAND U9941 ( .A(n8723), .B(n8722), .Z(n8730) );
  ANDN U9942 ( .B(a[576]), .A(n3956), .Z(n8728) );
  AND U9943 ( .A(b[1]), .B(a[575]), .Z(n8727) );
  XOR U9944 ( .A(n8728), .B(n8727), .Z(n8729) );
  XNOR U9945 ( .A(n8730), .B(n8729), .Z(n8732) );
  XOR U9946 ( .A(sreg[1598]), .B(n8731), .Z(n8726) );
  XNOR U9947 ( .A(n8732), .B(n8726), .Z(c[1598]) );
  NAND U9948 ( .A(b[0]), .B(a[577]), .Z(n8735) );
  NAND U9949 ( .A(a[576]), .B(b[1]), .Z(n8734) );
  XNOR U9950 ( .A(n8735), .B(n8734), .Z(n8737) );
  XNOR U9951 ( .A(n8736), .B(n8737), .Z(n8741) );
  XOR U9952 ( .A(n8740), .B(sreg[1599]), .Z(n8733) );
  XNOR U9953 ( .A(n8741), .B(n8733), .Z(c[1599]) );
  NAND U9954 ( .A(n8735), .B(n8734), .Z(n8739) );
  NANDN U9955 ( .A(n8737), .B(n8736), .Z(n8738) );
  NAND U9956 ( .A(n8739), .B(n8738), .Z(n8746) );
  ANDN U9957 ( .B(a[578]), .A(n3956), .Z(n8744) );
  AND U9958 ( .A(b[1]), .B(a[577]), .Z(n8743) );
  XOR U9959 ( .A(n8744), .B(n8743), .Z(n8745) );
  XNOR U9960 ( .A(n8746), .B(n8745), .Z(n8748) );
  XOR U9961 ( .A(sreg[1600]), .B(n8747), .Z(n8742) );
  XNOR U9962 ( .A(n8748), .B(n8742), .Z(c[1600]) );
  NAND U9963 ( .A(b[0]), .B(a[579]), .Z(n8751) );
  NAND U9964 ( .A(a[578]), .B(b[1]), .Z(n8750) );
  XNOR U9965 ( .A(n8751), .B(n8750), .Z(n8753) );
  XNOR U9966 ( .A(n8752), .B(n8753), .Z(n8757) );
  XOR U9967 ( .A(n8756), .B(sreg[1601]), .Z(n8749) );
  XNOR U9968 ( .A(n8757), .B(n8749), .Z(c[1601]) );
  NAND U9969 ( .A(n8751), .B(n8750), .Z(n8755) );
  NANDN U9970 ( .A(n8753), .B(n8752), .Z(n8754) );
  NAND U9971 ( .A(n8755), .B(n8754), .Z(n8762) );
  ANDN U9972 ( .B(a[580]), .A(n3957), .Z(n8760) );
  AND U9973 ( .A(b[1]), .B(a[579]), .Z(n8759) );
  XOR U9974 ( .A(n8760), .B(n8759), .Z(n8761) );
  XNOR U9975 ( .A(n8762), .B(n8761), .Z(n8767) );
  XOR U9976 ( .A(sreg[1602]), .B(n8766), .Z(n8758) );
  XNOR U9977 ( .A(n8767), .B(n8758), .Z(c[1602]) );
  OR U9978 ( .A(n8760), .B(n8759), .Z(n8765) );
  IV U9979 ( .A(n8761), .Z(n8763) );
  NANDN U9980 ( .A(n8763), .B(n8762), .Z(n8764) );
  NAND U9981 ( .A(n8765), .B(n8764), .Z(n8771) );
  NAND U9982 ( .A(b[0]), .B(a[581]), .Z(n8770) );
  NAND U9983 ( .A(a[580]), .B(b[1]), .Z(n8769) );
  XNOR U9984 ( .A(n8770), .B(n8769), .Z(n8772) );
  XNOR U9985 ( .A(n8771), .B(n8772), .Z(n8776) );
  XOR U9986 ( .A(n8775), .B(sreg[1603]), .Z(n8768) );
  XNOR U9987 ( .A(n8776), .B(n8768), .Z(c[1603]) );
  NAND U9988 ( .A(n8770), .B(n8769), .Z(n8774) );
  NANDN U9989 ( .A(n8772), .B(n8771), .Z(n8773) );
  NAND U9990 ( .A(n8774), .B(n8773), .Z(n8781) );
  ANDN U9991 ( .B(a[582]), .A(n3957), .Z(n8779) );
  AND U9992 ( .A(b[1]), .B(a[581]), .Z(n8778) );
  XOR U9993 ( .A(n8779), .B(n8778), .Z(n8780) );
  XNOR U9994 ( .A(n8781), .B(n8780), .Z(n8783) );
  XOR U9995 ( .A(sreg[1604]), .B(n8782), .Z(n8777) );
  XNOR U9996 ( .A(n8783), .B(n8777), .Z(c[1604]) );
  NAND U9997 ( .A(b[0]), .B(a[583]), .Z(n8786) );
  NAND U9998 ( .A(a[582]), .B(b[1]), .Z(n8785) );
  XNOR U9999 ( .A(n8786), .B(n8785), .Z(n8788) );
  XNOR U10000 ( .A(n8787), .B(n8788), .Z(n8792) );
  XOR U10001 ( .A(n8791), .B(sreg[1605]), .Z(n8784) );
  XNOR U10002 ( .A(n8792), .B(n8784), .Z(c[1605]) );
  NAND U10003 ( .A(n8786), .B(n8785), .Z(n8790) );
  NANDN U10004 ( .A(n8788), .B(n8787), .Z(n8789) );
  NAND U10005 ( .A(n8790), .B(n8789), .Z(n8797) );
  ANDN U10006 ( .B(a[584]), .A(n3957), .Z(n8795) );
  AND U10007 ( .A(b[1]), .B(a[583]), .Z(n8794) );
  XOR U10008 ( .A(n8795), .B(n8794), .Z(n8796) );
  XNOR U10009 ( .A(n8797), .B(n8796), .Z(n8799) );
  XOR U10010 ( .A(sreg[1606]), .B(n8798), .Z(n8793) );
  XNOR U10011 ( .A(n8799), .B(n8793), .Z(c[1606]) );
  NAND U10012 ( .A(b[0]), .B(a[585]), .Z(n8802) );
  NAND U10013 ( .A(a[584]), .B(b[1]), .Z(n8801) );
  XNOR U10014 ( .A(n8802), .B(n8801), .Z(n8804) );
  XNOR U10015 ( .A(n8803), .B(n8804), .Z(n8808) );
  XOR U10016 ( .A(n8807), .B(sreg[1607]), .Z(n8800) );
  XNOR U10017 ( .A(n8808), .B(n8800), .Z(c[1607]) );
  NAND U10018 ( .A(n8802), .B(n8801), .Z(n8806) );
  NANDN U10019 ( .A(n8804), .B(n8803), .Z(n8805) );
  NAND U10020 ( .A(n8806), .B(n8805), .Z(n8813) );
  ANDN U10021 ( .B(a[586]), .A(n3957), .Z(n8811) );
  AND U10022 ( .A(b[1]), .B(a[585]), .Z(n8810) );
  XOR U10023 ( .A(n8811), .B(n8810), .Z(n8812) );
  XNOR U10024 ( .A(n8813), .B(n8812), .Z(n8815) );
  XOR U10025 ( .A(sreg[1608]), .B(n8814), .Z(n8809) );
  XNOR U10026 ( .A(n8815), .B(n8809), .Z(c[1608]) );
  ANDN U10027 ( .B(a[587]), .A(n3957), .Z(n8818) );
  AND U10028 ( .A(b[1]), .B(a[586]), .Z(n8817) );
  XOR U10029 ( .A(n8818), .B(n8817), .Z(n8819) );
  XNOR U10030 ( .A(n8820), .B(n8819), .Z(n8822) );
  XNOR U10031 ( .A(sreg[1609]), .B(n8821), .Z(n8816) );
  XNOR U10032 ( .A(n8822), .B(n8816), .Z(c[1609]) );
  NAND U10033 ( .A(b[0]), .B(a[588]), .Z(n8825) );
  NAND U10034 ( .A(a[587]), .B(b[1]), .Z(n8824) );
  XNOR U10035 ( .A(n8825), .B(n8824), .Z(n8827) );
  XNOR U10036 ( .A(n8826), .B(n8827), .Z(n8831) );
  XOR U10037 ( .A(n8830), .B(sreg[1610]), .Z(n8823) );
  XNOR U10038 ( .A(n8831), .B(n8823), .Z(c[1610]) );
  NAND U10039 ( .A(n8825), .B(n8824), .Z(n8829) );
  NANDN U10040 ( .A(n8827), .B(n8826), .Z(n8828) );
  NAND U10041 ( .A(n8829), .B(n8828), .Z(n8835) );
  NAND U10042 ( .A(b[0]), .B(a[589]), .Z(n8834) );
  NAND U10043 ( .A(a[588]), .B(b[1]), .Z(n8833) );
  XNOR U10044 ( .A(n8834), .B(n8833), .Z(n8836) );
  XNOR U10045 ( .A(n8835), .B(n8836), .Z(n8840) );
  XOR U10046 ( .A(n8839), .B(sreg[1611]), .Z(n8832) );
  XNOR U10047 ( .A(n8840), .B(n8832), .Z(c[1611]) );
  NAND U10048 ( .A(n8834), .B(n8833), .Z(n8838) );
  NANDN U10049 ( .A(n8836), .B(n8835), .Z(n8837) );
  NAND U10050 ( .A(n8838), .B(n8837), .Z(n8845) );
  ANDN U10051 ( .B(a[590]), .A(n3957), .Z(n8843) );
  AND U10052 ( .A(b[1]), .B(a[589]), .Z(n8842) );
  XOR U10053 ( .A(n8843), .B(n8842), .Z(n8844) );
  XNOR U10054 ( .A(n8845), .B(n8844), .Z(n8847) );
  XOR U10055 ( .A(sreg[1612]), .B(n8846), .Z(n8841) );
  XNOR U10056 ( .A(n8847), .B(n8841), .Z(c[1612]) );
  NAND U10057 ( .A(b[0]), .B(a[591]), .Z(n8850) );
  NAND U10058 ( .A(a[590]), .B(b[1]), .Z(n8849) );
  XNOR U10059 ( .A(n8850), .B(n8849), .Z(n8852) );
  XNOR U10060 ( .A(n8851), .B(n8852), .Z(n8856) );
  XOR U10061 ( .A(n8855), .B(sreg[1613]), .Z(n8848) );
  XNOR U10062 ( .A(n8856), .B(n8848), .Z(c[1613]) );
  NAND U10063 ( .A(n8850), .B(n8849), .Z(n8854) );
  NANDN U10064 ( .A(n8852), .B(n8851), .Z(n8853) );
  NAND U10065 ( .A(n8854), .B(n8853), .Z(n8861) );
  ANDN U10066 ( .B(a[592]), .A(n3957), .Z(n8859) );
  AND U10067 ( .A(b[1]), .B(a[591]), .Z(n8858) );
  XOR U10068 ( .A(n8859), .B(n8858), .Z(n8860) );
  XNOR U10069 ( .A(n8861), .B(n8860), .Z(n8863) );
  XOR U10070 ( .A(sreg[1614]), .B(n8862), .Z(n8857) );
  XNOR U10071 ( .A(n8863), .B(n8857), .Z(c[1614]) );
  NAND U10072 ( .A(b[0]), .B(a[593]), .Z(n8866) );
  NAND U10073 ( .A(a[592]), .B(b[1]), .Z(n8865) );
  XNOR U10074 ( .A(n8866), .B(n8865), .Z(n8868) );
  XNOR U10075 ( .A(n8867), .B(n8868), .Z(n8872) );
  XOR U10076 ( .A(n8871), .B(sreg[1615]), .Z(n8864) );
  XNOR U10077 ( .A(n8872), .B(n8864), .Z(c[1615]) );
  NAND U10078 ( .A(n8866), .B(n8865), .Z(n8870) );
  NANDN U10079 ( .A(n8868), .B(n8867), .Z(n8869) );
  NAND U10080 ( .A(n8870), .B(n8869), .Z(n8877) );
  ANDN U10081 ( .B(a[594]), .A(n3958), .Z(n8875) );
  AND U10082 ( .A(b[1]), .B(a[593]), .Z(n8874) );
  XOR U10083 ( .A(n8875), .B(n8874), .Z(n8876) );
  XNOR U10084 ( .A(n8877), .B(n8876), .Z(n8882) );
  XOR U10085 ( .A(sreg[1616]), .B(n8881), .Z(n8873) );
  XNOR U10086 ( .A(n8882), .B(n8873), .Z(c[1616]) );
  OR U10087 ( .A(n8875), .B(n8874), .Z(n8880) );
  IV U10088 ( .A(n8876), .Z(n8878) );
  NANDN U10089 ( .A(n8878), .B(n8877), .Z(n8879) );
  NAND U10090 ( .A(n8880), .B(n8879), .Z(n8886) );
  NAND U10091 ( .A(b[0]), .B(a[595]), .Z(n8885) );
  NAND U10092 ( .A(a[594]), .B(b[1]), .Z(n8884) );
  XNOR U10093 ( .A(n8885), .B(n8884), .Z(n8887) );
  XNOR U10094 ( .A(n8886), .B(n8887), .Z(n8891) );
  XOR U10095 ( .A(n8890), .B(sreg[1617]), .Z(n8883) );
  XNOR U10096 ( .A(n8891), .B(n8883), .Z(c[1617]) );
  NAND U10097 ( .A(n8885), .B(n8884), .Z(n8889) );
  NANDN U10098 ( .A(n8887), .B(n8886), .Z(n8888) );
  NAND U10099 ( .A(n8889), .B(n8888), .Z(n8895) );
  NAND U10100 ( .A(b[0]), .B(a[596]), .Z(n8894) );
  NAND U10101 ( .A(a[595]), .B(b[1]), .Z(n8893) );
  XNOR U10102 ( .A(n8894), .B(n8893), .Z(n8896) );
  XNOR U10103 ( .A(n8895), .B(n8896), .Z(n8900) );
  XOR U10104 ( .A(n8899), .B(sreg[1618]), .Z(n8892) );
  XNOR U10105 ( .A(n8900), .B(n8892), .Z(c[1618]) );
  NAND U10106 ( .A(n8894), .B(n8893), .Z(n8898) );
  NANDN U10107 ( .A(n8896), .B(n8895), .Z(n8897) );
  NAND U10108 ( .A(n8898), .B(n8897), .Z(n8904) );
  NAND U10109 ( .A(b[0]), .B(a[597]), .Z(n8903) );
  NAND U10110 ( .A(a[596]), .B(b[1]), .Z(n8902) );
  XNOR U10111 ( .A(n8903), .B(n8902), .Z(n8905) );
  XNOR U10112 ( .A(n8904), .B(n8905), .Z(n8909) );
  XOR U10113 ( .A(n8908), .B(sreg[1619]), .Z(n8901) );
  XNOR U10114 ( .A(n8909), .B(n8901), .Z(c[1619]) );
  NAND U10115 ( .A(n8903), .B(n8902), .Z(n8907) );
  NANDN U10116 ( .A(n8905), .B(n8904), .Z(n8906) );
  NAND U10117 ( .A(n8907), .B(n8906), .Z(n8914) );
  ANDN U10118 ( .B(a[598]), .A(n3958), .Z(n8912) );
  AND U10119 ( .A(b[1]), .B(a[597]), .Z(n8911) );
  XOR U10120 ( .A(n8912), .B(n8911), .Z(n8913) );
  XNOR U10121 ( .A(n8914), .B(n8913), .Z(n8916) );
  XOR U10122 ( .A(sreg[1620]), .B(n8915), .Z(n8910) );
  XNOR U10123 ( .A(n8916), .B(n8910), .Z(c[1620]) );
  NAND U10124 ( .A(b[0]), .B(a[599]), .Z(n8919) );
  NAND U10125 ( .A(a[598]), .B(b[1]), .Z(n8918) );
  XNOR U10126 ( .A(n8919), .B(n8918), .Z(n8921) );
  XNOR U10127 ( .A(n8920), .B(n8921), .Z(n8925) );
  XOR U10128 ( .A(n8924), .B(sreg[1621]), .Z(n8917) );
  XNOR U10129 ( .A(n8925), .B(n8917), .Z(c[1621]) );
  NAND U10130 ( .A(n8919), .B(n8918), .Z(n8923) );
  NANDN U10131 ( .A(n8921), .B(n8920), .Z(n8922) );
  NAND U10132 ( .A(n8923), .B(n8922), .Z(n8930) );
  ANDN U10133 ( .B(a[600]), .A(n3958), .Z(n8928) );
  AND U10134 ( .A(b[1]), .B(a[599]), .Z(n8927) );
  XOR U10135 ( .A(n8928), .B(n8927), .Z(n8929) );
  XNOR U10136 ( .A(n8930), .B(n8929), .Z(n8932) );
  XOR U10137 ( .A(sreg[1622]), .B(n8931), .Z(n8926) );
  XNOR U10138 ( .A(n8932), .B(n8926), .Z(c[1622]) );
  NAND U10139 ( .A(b[0]), .B(a[601]), .Z(n8935) );
  NAND U10140 ( .A(a[600]), .B(b[1]), .Z(n8934) );
  XNOR U10141 ( .A(n8935), .B(n8934), .Z(n8937) );
  XNOR U10142 ( .A(n8936), .B(n8937), .Z(n8941) );
  XOR U10143 ( .A(n8940), .B(sreg[1623]), .Z(n8933) );
  XNOR U10144 ( .A(n8941), .B(n8933), .Z(c[1623]) );
  NAND U10145 ( .A(n8935), .B(n8934), .Z(n8939) );
  NANDN U10146 ( .A(n8937), .B(n8936), .Z(n8938) );
  NAND U10147 ( .A(n8939), .B(n8938), .Z(n8946) );
  ANDN U10148 ( .B(a[602]), .A(n3958), .Z(n8944) );
  AND U10149 ( .A(b[1]), .B(a[601]), .Z(n8943) );
  XOR U10150 ( .A(n8944), .B(n8943), .Z(n8945) );
  XNOR U10151 ( .A(n8946), .B(n8945), .Z(n8948) );
  XOR U10152 ( .A(sreg[1624]), .B(n8947), .Z(n8942) );
  XNOR U10153 ( .A(n8948), .B(n8942), .Z(c[1624]) );
  ANDN U10154 ( .B(a[603]), .A(n3958), .Z(n8951) );
  AND U10155 ( .A(b[1]), .B(a[602]), .Z(n8950) );
  XOR U10156 ( .A(n8951), .B(n8950), .Z(n8952) );
  XNOR U10157 ( .A(n8953), .B(n8952), .Z(n8955) );
  XNOR U10158 ( .A(sreg[1625]), .B(n8954), .Z(n8949) );
  XNOR U10159 ( .A(n8955), .B(n8949), .Z(c[1625]) );
  ANDN U10160 ( .B(a[604]), .A(n3958), .Z(n8958) );
  AND U10161 ( .A(b[1]), .B(a[603]), .Z(n8957) );
  XOR U10162 ( .A(n8958), .B(n8957), .Z(n8959) );
  XNOR U10163 ( .A(n8960), .B(n8959), .Z(n8962) );
  XNOR U10164 ( .A(sreg[1626]), .B(n8961), .Z(n8956) );
  XNOR U10165 ( .A(n8962), .B(n8956), .Z(c[1626]) );
  NAND U10166 ( .A(b[0]), .B(a[605]), .Z(n8965) );
  NAND U10167 ( .A(a[604]), .B(b[1]), .Z(n8964) );
  XNOR U10168 ( .A(n8965), .B(n8964), .Z(n8967) );
  XNOR U10169 ( .A(n8966), .B(n8967), .Z(n8971) );
  XOR U10170 ( .A(n8970), .B(sreg[1627]), .Z(n8963) );
  XNOR U10171 ( .A(n8971), .B(n8963), .Z(c[1627]) );
  NAND U10172 ( .A(n8965), .B(n8964), .Z(n8969) );
  NANDN U10173 ( .A(n8967), .B(n8966), .Z(n8968) );
  NAND U10174 ( .A(n8969), .B(n8968), .Z(n8975) );
  NAND U10175 ( .A(b[0]), .B(a[606]), .Z(n8974) );
  NAND U10176 ( .A(a[605]), .B(b[1]), .Z(n8973) );
  XNOR U10177 ( .A(n8974), .B(n8973), .Z(n8976) );
  XNOR U10178 ( .A(n8975), .B(n8976), .Z(n8980) );
  XOR U10179 ( .A(n8979), .B(sreg[1628]), .Z(n8972) );
  XNOR U10180 ( .A(n8980), .B(n8972), .Z(c[1628]) );
  NAND U10181 ( .A(n8974), .B(n8973), .Z(n8978) );
  NANDN U10182 ( .A(n8976), .B(n8975), .Z(n8977) );
  NAND U10183 ( .A(n8978), .B(n8977), .Z(n8984) );
  NAND U10184 ( .A(b[0]), .B(a[607]), .Z(n8983) );
  NAND U10185 ( .A(a[606]), .B(b[1]), .Z(n8982) );
  XNOR U10186 ( .A(n8983), .B(n8982), .Z(n8985) );
  XNOR U10187 ( .A(n8984), .B(n8985), .Z(n8989) );
  XOR U10188 ( .A(n8988), .B(sreg[1629]), .Z(n8981) );
  XNOR U10189 ( .A(n8989), .B(n8981), .Z(c[1629]) );
  NAND U10190 ( .A(n8983), .B(n8982), .Z(n8987) );
  NANDN U10191 ( .A(n8985), .B(n8984), .Z(n8986) );
  NAND U10192 ( .A(n8987), .B(n8986), .Z(n8994) );
  ANDN U10193 ( .B(a[608]), .A(n3958), .Z(n8992) );
  AND U10194 ( .A(b[1]), .B(a[607]), .Z(n8991) );
  XOR U10195 ( .A(n8992), .B(n8991), .Z(n8993) );
  XNOR U10196 ( .A(n8994), .B(n8993), .Z(n8996) );
  XOR U10197 ( .A(sreg[1630]), .B(n8995), .Z(n8990) );
  XNOR U10198 ( .A(n8996), .B(n8990), .Z(c[1630]) );
  NAND U10199 ( .A(b[0]), .B(a[609]), .Z(n8999) );
  NAND U10200 ( .A(a[608]), .B(b[1]), .Z(n8998) );
  XNOR U10201 ( .A(n8999), .B(n8998), .Z(n9001) );
  XNOR U10202 ( .A(n9000), .B(n9001), .Z(n9005) );
  XOR U10203 ( .A(n9004), .B(sreg[1631]), .Z(n8997) );
  XNOR U10204 ( .A(n9005), .B(n8997), .Z(c[1631]) );
  NAND U10205 ( .A(n8999), .B(n8998), .Z(n9003) );
  NANDN U10206 ( .A(n9001), .B(n9000), .Z(n9002) );
  NAND U10207 ( .A(n9003), .B(n9002), .Z(n9009) );
  NAND U10208 ( .A(b[0]), .B(a[610]), .Z(n9008) );
  NAND U10209 ( .A(a[609]), .B(b[1]), .Z(n9007) );
  XNOR U10210 ( .A(n9008), .B(n9007), .Z(n9010) );
  XNOR U10211 ( .A(n9009), .B(n9010), .Z(n9014) );
  XOR U10212 ( .A(n9013), .B(sreg[1632]), .Z(n9006) );
  XNOR U10213 ( .A(n9014), .B(n9006), .Z(c[1632]) );
  NAND U10214 ( .A(n9008), .B(n9007), .Z(n9012) );
  NANDN U10215 ( .A(n9010), .B(n9009), .Z(n9011) );
  NAND U10216 ( .A(n9012), .B(n9011), .Z(n9018) );
  NAND U10217 ( .A(b[0]), .B(a[611]), .Z(n9017) );
  NAND U10218 ( .A(a[610]), .B(b[1]), .Z(n9016) );
  XNOR U10219 ( .A(n9017), .B(n9016), .Z(n9019) );
  XNOR U10220 ( .A(n9018), .B(n9019), .Z(n9023) );
  XOR U10221 ( .A(n9022), .B(sreg[1633]), .Z(n9015) );
  XNOR U10222 ( .A(n9023), .B(n9015), .Z(c[1633]) );
  NAND U10223 ( .A(n9017), .B(n9016), .Z(n9021) );
  NANDN U10224 ( .A(n9019), .B(n9018), .Z(n9020) );
  NAND U10225 ( .A(n9021), .B(n9020), .Z(n9028) );
  ANDN U10226 ( .B(a[612]), .A(n3959), .Z(n9026) );
  AND U10227 ( .A(b[1]), .B(a[611]), .Z(n9025) );
  XOR U10228 ( .A(n9026), .B(n9025), .Z(n9027) );
  XNOR U10229 ( .A(n9028), .B(n9027), .Z(n9033) );
  XOR U10230 ( .A(sreg[1634]), .B(n9032), .Z(n9024) );
  XNOR U10231 ( .A(n9033), .B(n9024), .Z(c[1634]) );
  OR U10232 ( .A(n9026), .B(n9025), .Z(n9031) );
  IV U10233 ( .A(n9027), .Z(n9029) );
  NANDN U10234 ( .A(n9029), .B(n9028), .Z(n9030) );
  NAND U10235 ( .A(n9031), .B(n9030), .Z(n9037) );
  NAND U10236 ( .A(b[0]), .B(a[613]), .Z(n9036) );
  NAND U10237 ( .A(a[612]), .B(b[1]), .Z(n9035) );
  XNOR U10238 ( .A(n9036), .B(n9035), .Z(n9038) );
  XNOR U10239 ( .A(n9037), .B(n9038), .Z(n9042) );
  XOR U10240 ( .A(n9041), .B(sreg[1635]), .Z(n9034) );
  XNOR U10241 ( .A(n9042), .B(n9034), .Z(c[1635]) );
  NAND U10242 ( .A(n9036), .B(n9035), .Z(n9040) );
  NANDN U10243 ( .A(n9038), .B(n9037), .Z(n9039) );
  NAND U10244 ( .A(n9040), .B(n9039), .Z(n9047) );
  ANDN U10245 ( .B(a[614]), .A(n3959), .Z(n9045) );
  AND U10246 ( .A(b[1]), .B(a[613]), .Z(n9044) );
  XOR U10247 ( .A(n9045), .B(n9044), .Z(n9046) );
  XNOR U10248 ( .A(n9047), .B(n9046), .Z(n9049) );
  XOR U10249 ( .A(sreg[1636]), .B(n9048), .Z(n9043) );
  XNOR U10250 ( .A(n9049), .B(n9043), .Z(c[1636]) );
  NAND U10251 ( .A(b[0]), .B(a[615]), .Z(n9052) );
  NAND U10252 ( .A(a[614]), .B(b[1]), .Z(n9051) );
  XNOR U10253 ( .A(n9052), .B(n9051), .Z(n9054) );
  XNOR U10254 ( .A(n9053), .B(n9054), .Z(n9058) );
  XOR U10255 ( .A(n9057), .B(sreg[1637]), .Z(n9050) );
  XNOR U10256 ( .A(n9058), .B(n9050), .Z(c[1637]) );
  NAND U10257 ( .A(n9052), .B(n9051), .Z(n9056) );
  NANDN U10258 ( .A(n9054), .B(n9053), .Z(n9055) );
  NAND U10259 ( .A(n9056), .B(n9055), .Z(n9062) );
  NAND U10260 ( .A(b[0]), .B(a[616]), .Z(n9061) );
  NAND U10261 ( .A(a[615]), .B(b[1]), .Z(n9060) );
  XNOR U10262 ( .A(n9061), .B(n9060), .Z(n9063) );
  XNOR U10263 ( .A(n9062), .B(n9063), .Z(n9067) );
  XOR U10264 ( .A(n9066), .B(sreg[1638]), .Z(n9059) );
  XNOR U10265 ( .A(n9067), .B(n9059), .Z(c[1638]) );
  NAND U10266 ( .A(n9061), .B(n9060), .Z(n9065) );
  NANDN U10267 ( .A(n9063), .B(n9062), .Z(n9064) );
  NAND U10268 ( .A(n9065), .B(n9064), .Z(n9071) );
  NAND U10269 ( .A(b[0]), .B(a[617]), .Z(n9070) );
  NAND U10270 ( .A(a[616]), .B(b[1]), .Z(n9069) );
  XNOR U10271 ( .A(n9070), .B(n9069), .Z(n9072) );
  XNOR U10272 ( .A(n9071), .B(n9072), .Z(n9076) );
  XOR U10273 ( .A(n9075), .B(sreg[1639]), .Z(n9068) );
  XNOR U10274 ( .A(n9076), .B(n9068), .Z(c[1639]) );
  NAND U10275 ( .A(n9070), .B(n9069), .Z(n9074) );
  NANDN U10276 ( .A(n9072), .B(n9071), .Z(n9073) );
  NAND U10277 ( .A(n9074), .B(n9073), .Z(n9081) );
  ANDN U10278 ( .B(a[618]), .A(n3959), .Z(n9079) );
  AND U10279 ( .A(b[1]), .B(a[617]), .Z(n9078) );
  XOR U10280 ( .A(n9079), .B(n9078), .Z(n9080) );
  XNOR U10281 ( .A(n9081), .B(n9080), .Z(n9083) );
  XOR U10282 ( .A(sreg[1640]), .B(n9082), .Z(n9077) );
  XNOR U10283 ( .A(n9083), .B(n9077), .Z(c[1640]) );
  NAND U10284 ( .A(b[0]), .B(a[619]), .Z(n9086) );
  NAND U10285 ( .A(a[618]), .B(b[1]), .Z(n9085) );
  XNOR U10286 ( .A(n9086), .B(n9085), .Z(n9088) );
  XNOR U10287 ( .A(n9087), .B(n9088), .Z(n9092) );
  XOR U10288 ( .A(n9091), .B(sreg[1641]), .Z(n9084) );
  XNOR U10289 ( .A(n9092), .B(n9084), .Z(c[1641]) );
  NAND U10290 ( .A(n9086), .B(n9085), .Z(n9090) );
  NANDN U10291 ( .A(n9088), .B(n9087), .Z(n9089) );
  NAND U10292 ( .A(n9090), .B(n9089), .Z(n9097) );
  ANDN U10293 ( .B(a[620]), .A(n3959), .Z(n9095) );
  AND U10294 ( .A(b[1]), .B(a[619]), .Z(n9094) );
  XOR U10295 ( .A(n9095), .B(n9094), .Z(n9096) );
  XNOR U10296 ( .A(n9097), .B(n9096), .Z(n9099) );
  XOR U10297 ( .A(sreg[1642]), .B(n9098), .Z(n9093) );
  XNOR U10298 ( .A(n9099), .B(n9093), .Z(c[1642]) );
  NAND U10299 ( .A(b[0]), .B(a[621]), .Z(n9102) );
  NAND U10300 ( .A(a[620]), .B(b[1]), .Z(n9101) );
  XNOR U10301 ( .A(n9102), .B(n9101), .Z(n9104) );
  XNOR U10302 ( .A(n9103), .B(n9104), .Z(n9108) );
  XOR U10303 ( .A(n9107), .B(sreg[1643]), .Z(n9100) );
  XNOR U10304 ( .A(n9108), .B(n9100), .Z(c[1643]) );
  NAND U10305 ( .A(n9102), .B(n9101), .Z(n9106) );
  NANDN U10306 ( .A(n9104), .B(n9103), .Z(n9105) );
  NAND U10307 ( .A(n9106), .B(n9105), .Z(n9113) );
  ANDN U10308 ( .B(a[622]), .A(n3959), .Z(n9111) );
  AND U10309 ( .A(b[1]), .B(a[621]), .Z(n9110) );
  XOR U10310 ( .A(n9111), .B(n9110), .Z(n9112) );
  XNOR U10311 ( .A(n9113), .B(n9112), .Z(n9115) );
  XOR U10312 ( .A(sreg[1644]), .B(n9114), .Z(n9109) );
  XNOR U10313 ( .A(n9115), .B(n9109), .Z(c[1644]) );
  ANDN U10314 ( .B(a[623]), .A(n3959), .Z(n9118) );
  AND U10315 ( .A(b[1]), .B(a[622]), .Z(n9117) );
  XOR U10316 ( .A(n9118), .B(n9117), .Z(n9119) );
  XNOR U10317 ( .A(n9120), .B(n9119), .Z(n9122) );
  XNOR U10318 ( .A(sreg[1645]), .B(n9121), .Z(n9116) );
  XNOR U10319 ( .A(n9122), .B(n9116), .Z(c[1645]) );
  ANDN U10320 ( .B(a[624]), .A(n3959), .Z(n9125) );
  AND U10321 ( .A(b[1]), .B(a[623]), .Z(n9124) );
  XOR U10322 ( .A(n9125), .B(n9124), .Z(n9126) );
  XNOR U10323 ( .A(n9127), .B(n9126), .Z(n9129) );
  XNOR U10324 ( .A(sreg[1646]), .B(n9128), .Z(n9123) );
  XNOR U10325 ( .A(n9129), .B(n9123), .Z(c[1646]) );
  NAND U10326 ( .A(b[0]), .B(a[625]), .Z(n9132) );
  NAND U10327 ( .A(a[624]), .B(b[1]), .Z(n9131) );
  XNOR U10328 ( .A(n9132), .B(n9131), .Z(n9134) );
  XNOR U10329 ( .A(n9133), .B(n9134), .Z(n9138) );
  XOR U10330 ( .A(n9137), .B(sreg[1647]), .Z(n9130) );
  XNOR U10331 ( .A(n9138), .B(n9130), .Z(c[1647]) );
  NAND U10332 ( .A(n9132), .B(n9131), .Z(n9136) );
  NANDN U10333 ( .A(n9134), .B(n9133), .Z(n9135) );
  NAND U10334 ( .A(n9136), .B(n9135), .Z(n9143) );
  ANDN U10335 ( .B(a[626]), .A(n3960), .Z(n9141) );
  AND U10336 ( .A(b[1]), .B(a[625]), .Z(n9140) );
  XOR U10337 ( .A(n9141), .B(n9140), .Z(n9142) );
  XNOR U10338 ( .A(n9143), .B(n9142), .Z(n9148) );
  XOR U10339 ( .A(sreg[1648]), .B(n9147), .Z(n9139) );
  XNOR U10340 ( .A(n9148), .B(n9139), .Z(c[1648]) );
  OR U10341 ( .A(n9141), .B(n9140), .Z(n9146) );
  IV U10342 ( .A(n9142), .Z(n9144) );
  NANDN U10343 ( .A(n9144), .B(n9143), .Z(n9145) );
  NAND U10344 ( .A(n9146), .B(n9145), .Z(n9152) );
  NAND U10345 ( .A(b[0]), .B(a[627]), .Z(n9151) );
  NAND U10346 ( .A(a[626]), .B(b[1]), .Z(n9150) );
  XNOR U10347 ( .A(n9151), .B(n9150), .Z(n9153) );
  XNOR U10348 ( .A(n9152), .B(n9153), .Z(n9157) );
  XOR U10349 ( .A(n9156), .B(sreg[1649]), .Z(n9149) );
  XNOR U10350 ( .A(n9157), .B(n9149), .Z(c[1649]) );
  NAND U10351 ( .A(n9151), .B(n9150), .Z(n9155) );
  NANDN U10352 ( .A(n9153), .B(n9152), .Z(n9154) );
  NAND U10353 ( .A(n9155), .B(n9154), .Z(n9162) );
  ANDN U10354 ( .B(a[628]), .A(n3960), .Z(n9160) );
  AND U10355 ( .A(b[1]), .B(a[627]), .Z(n9159) );
  XOR U10356 ( .A(n9160), .B(n9159), .Z(n9161) );
  XNOR U10357 ( .A(n9162), .B(n9161), .Z(n9164) );
  XOR U10358 ( .A(sreg[1650]), .B(n9163), .Z(n9158) );
  XNOR U10359 ( .A(n9164), .B(n9158), .Z(c[1650]) );
  NAND U10360 ( .A(b[0]), .B(a[629]), .Z(n9167) );
  NAND U10361 ( .A(a[628]), .B(b[1]), .Z(n9166) );
  XNOR U10362 ( .A(n9167), .B(n9166), .Z(n9169) );
  XNOR U10363 ( .A(n9168), .B(n9169), .Z(n9173) );
  XOR U10364 ( .A(n9172), .B(sreg[1651]), .Z(n9165) );
  XNOR U10365 ( .A(n9173), .B(n9165), .Z(c[1651]) );
  NAND U10366 ( .A(n9167), .B(n9166), .Z(n9171) );
  NANDN U10367 ( .A(n9169), .B(n9168), .Z(n9170) );
  NAND U10368 ( .A(n9171), .B(n9170), .Z(n9178) );
  ANDN U10369 ( .B(a[630]), .A(n3960), .Z(n9176) );
  AND U10370 ( .A(b[1]), .B(a[629]), .Z(n9175) );
  XOR U10371 ( .A(n9176), .B(n9175), .Z(n9177) );
  XNOR U10372 ( .A(n9178), .B(n9177), .Z(n9180) );
  XOR U10373 ( .A(sreg[1652]), .B(n9179), .Z(n9174) );
  XNOR U10374 ( .A(n9180), .B(n9174), .Z(c[1652]) );
  ANDN U10375 ( .B(a[631]), .A(n3960), .Z(n9183) );
  AND U10376 ( .A(b[1]), .B(a[630]), .Z(n9182) );
  XOR U10377 ( .A(n9183), .B(n9182), .Z(n9184) );
  XNOR U10378 ( .A(n9185), .B(n9184), .Z(n9187) );
  XNOR U10379 ( .A(sreg[1653]), .B(n9186), .Z(n9181) );
  XNOR U10380 ( .A(n9187), .B(n9181), .Z(c[1653]) );
  ANDN U10381 ( .B(a[632]), .A(n3960), .Z(n9190) );
  AND U10382 ( .A(b[1]), .B(a[631]), .Z(n9189) );
  XOR U10383 ( .A(n9190), .B(n9189), .Z(n9191) );
  XNOR U10384 ( .A(n9192), .B(n9191), .Z(n9194) );
  XNOR U10385 ( .A(sreg[1654]), .B(n9193), .Z(n9188) );
  XNOR U10386 ( .A(n9194), .B(n9188), .Z(c[1654]) );
  NAND U10387 ( .A(b[0]), .B(a[633]), .Z(n9197) );
  NAND U10388 ( .A(a[632]), .B(b[1]), .Z(n9196) );
  XNOR U10389 ( .A(n9197), .B(n9196), .Z(n9199) );
  XNOR U10390 ( .A(n9198), .B(n9199), .Z(n9203) );
  XOR U10391 ( .A(n9202), .B(sreg[1655]), .Z(n9195) );
  XNOR U10392 ( .A(n9203), .B(n9195), .Z(c[1655]) );
  NAND U10393 ( .A(n9197), .B(n9196), .Z(n9201) );
  NANDN U10394 ( .A(n9199), .B(n9198), .Z(n9200) );
  NAND U10395 ( .A(n9201), .B(n9200), .Z(n9208) );
  ANDN U10396 ( .B(a[634]), .A(n3960), .Z(n9206) );
  AND U10397 ( .A(b[1]), .B(a[633]), .Z(n9205) );
  XOR U10398 ( .A(n9206), .B(n9205), .Z(n9207) );
  XNOR U10399 ( .A(n9208), .B(n9207), .Z(n9210) );
  XOR U10400 ( .A(sreg[1656]), .B(n9209), .Z(n9204) );
  XNOR U10401 ( .A(n9210), .B(n9204), .Z(c[1656]) );
  ANDN U10402 ( .B(a[635]), .A(n3960), .Z(n9213) );
  AND U10403 ( .A(b[1]), .B(a[634]), .Z(n9212) );
  XOR U10404 ( .A(n9213), .B(n9212), .Z(n9214) );
  XNOR U10405 ( .A(n9215), .B(n9214), .Z(n9217) );
  XNOR U10406 ( .A(sreg[1657]), .B(n9216), .Z(n9211) );
  XNOR U10407 ( .A(n9217), .B(n9211), .Z(c[1657]) );
  ANDN U10408 ( .B(a[636]), .A(n3961), .Z(n9220) );
  AND U10409 ( .A(b[1]), .B(a[635]), .Z(n9219) );
  XOR U10410 ( .A(n9220), .B(n9219), .Z(n9221) );
  XNOR U10411 ( .A(n9222), .B(n9221), .Z(n9227) );
  XNOR U10412 ( .A(sreg[1658]), .B(n9226), .Z(n9218) );
  XNOR U10413 ( .A(n9227), .B(n9218), .Z(c[1658]) );
  OR U10414 ( .A(n9220), .B(n9219), .Z(n9225) );
  IV U10415 ( .A(n9221), .Z(n9223) );
  NANDN U10416 ( .A(n9223), .B(n9222), .Z(n9224) );
  NAND U10417 ( .A(n9225), .B(n9224), .Z(n9231) );
  NAND U10418 ( .A(b[0]), .B(a[637]), .Z(n9230) );
  NAND U10419 ( .A(a[636]), .B(b[1]), .Z(n9229) );
  XNOR U10420 ( .A(n9230), .B(n9229), .Z(n9232) );
  XNOR U10421 ( .A(n9231), .B(n9232), .Z(n9236) );
  XOR U10422 ( .A(n9235), .B(sreg[1659]), .Z(n9228) );
  XNOR U10423 ( .A(n9236), .B(n9228), .Z(c[1659]) );
  NAND U10424 ( .A(n9230), .B(n9229), .Z(n9234) );
  NANDN U10425 ( .A(n9232), .B(n9231), .Z(n9233) );
  NAND U10426 ( .A(n9234), .B(n9233), .Z(n9241) );
  ANDN U10427 ( .B(a[638]), .A(n3961), .Z(n9239) );
  AND U10428 ( .A(b[1]), .B(a[637]), .Z(n9238) );
  XOR U10429 ( .A(n9239), .B(n9238), .Z(n9240) );
  XNOR U10430 ( .A(n9241), .B(n9240), .Z(n9243) );
  XOR U10431 ( .A(sreg[1660]), .B(n9242), .Z(n9237) );
  XNOR U10432 ( .A(n9243), .B(n9237), .Z(c[1660]) );
  NAND U10433 ( .A(b[0]), .B(a[639]), .Z(n9246) );
  NAND U10434 ( .A(a[638]), .B(b[1]), .Z(n9245) );
  XNOR U10435 ( .A(n9246), .B(n9245), .Z(n9248) );
  XNOR U10436 ( .A(n9247), .B(n9248), .Z(n9252) );
  XOR U10437 ( .A(n9251), .B(sreg[1661]), .Z(n9244) );
  XNOR U10438 ( .A(n9252), .B(n9244), .Z(c[1661]) );
  NAND U10439 ( .A(n9246), .B(n9245), .Z(n9250) );
  NANDN U10440 ( .A(n9248), .B(n9247), .Z(n9249) );
  NAND U10441 ( .A(n9250), .B(n9249), .Z(n9257) );
  ANDN U10442 ( .B(a[640]), .A(n3961), .Z(n9255) );
  AND U10443 ( .A(b[1]), .B(a[639]), .Z(n9254) );
  XOR U10444 ( .A(n9255), .B(n9254), .Z(n9256) );
  XNOR U10445 ( .A(n9257), .B(n9256), .Z(n9259) );
  XOR U10446 ( .A(sreg[1662]), .B(n9258), .Z(n9253) );
  XNOR U10447 ( .A(n9259), .B(n9253), .Z(c[1662]) );
  NAND U10448 ( .A(b[0]), .B(a[641]), .Z(n9262) );
  NAND U10449 ( .A(a[640]), .B(b[1]), .Z(n9261) );
  XNOR U10450 ( .A(n9262), .B(n9261), .Z(n9264) );
  XNOR U10451 ( .A(n9263), .B(n9264), .Z(n9268) );
  XOR U10452 ( .A(n9267), .B(sreg[1663]), .Z(n9260) );
  XNOR U10453 ( .A(n9268), .B(n9260), .Z(c[1663]) );
  NAND U10454 ( .A(n9262), .B(n9261), .Z(n9266) );
  NANDN U10455 ( .A(n9264), .B(n9263), .Z(n9265) );
  NAND U10456 ( .A(n9266), .B(n9265), .Z(n9272) );
  NAND U10457 ( .A(b[0]), .B(a[642]), .Z(n9271) );
  NAND U10458 ( .A(a[641]), .B(b[1]), .Z(n9270) );
  XNOR U10459 ( .A(n9271), .B(n9270), .Z(n9273) );
  XNOR U10460 ( .A(n9272), .B(n9273), .Z(n9277) );
  XOR U10461 ( .A(n9276), .B(sreg[1664]), .Z(n9269) );
  XNOR U10462 ( .A(n9277), .B(n9269), .Z(c[1664]) );
  NAND U10463 ( .A(n9271), .B(n9270), .Z(n9275) );
  NANDN U10464 ( .A(n9273), .B(n9272), .Z(n9274) );
  NAND U10465 ( .A(n9275), .B(n9274), .Z(n9281) );
  NAND U10466 ( .A(b[0]), .B(a[643]), .Z(n9280) );
  NAND U10467 ( .A(a[642]), .B(b[1]), .Z(n9279) );
  XNOR U10468 ( .A(n9280), .B(n9279), .Z(n9282) );
  XNOR U10469 ( .A(n9281), .B(n9282), .Z(n9286) );
  XOR U10470 ( .A(n9285), .B(sreg[1665]), .Z(n9278) );
  XNOR U10471 ( .A(n9286), .B(n9278), .Z(c[1665]) );
  NAND U10472 ( .A(n9280), .B(n9279), .Z(n9284) );
  NANDN U10473 ( .A(n9282), .B(n9281), .Z(n9283) );
  NAND U10474 ( .A(n9284), .B(n9283), .Z(n9291) );
  ANDN U10475 ( .B(a[644]), .A(n3961), .Z(n9289) );
  AND U10476 ( .A(b[1]), .B(a[643]), .Z(n9288) );
  XOR U10477 ( .A(n9289), .B(n9288), .Z(n9290) );
  XNOR U10478 ( .A(n9291), .B(n9290), .Z(n9293) );
  XOR U10479 ( .A(sreg[1666]), .B(n9292), .Z(n9287) );
  XNOR U10480 ( .A(n9293), .B(n9287), .Z(c[1666]) );
  NAND U10481 ( .A(b[0]), .B(a[645]), .Z(n9296) );
  NAND U10482 ( .A(a[644]), .B(b[1]), .Z(n9295) );
  XNOR U10483 ( .A(n9296), .B(n9295), .Z(n9298) );
  XNOR U10484 ( .A(n9297), .B(n9298), .Z(n9302) );
  XOR U10485 ( .A(n9301), .B(sreg[1667]), .Z(n9294) );
  XNOR U10486 ( .A(n9302), .B(n9294), .Z(c[1667]) );
  NAND U10487 ( .A(n9296), .B(n9295), .Z(n9300) );
  NANDN U10488 ( .A(n9298), .B(n9297), .Z(n9299) );
  NAND U10489 ( .A(n9300), .B(n9299), .Z(n9307) );
  ANDN U10490 ( .B(a[646]), .A(n3961), .Z(n9305) );
  AND U10491 ( .A(b[1]), .B(a[645]), .Z(n9304) );
  XOR U10492 ( .A(n9305), .B(n9304), .Z(n9306) );
  XNOR U10493 ( .A(n9307), .B(n9306), .Z(n9309) );
  XOR U10494 ( .A(sreg[1668]), .B(n9308), .Z(n9303) );
  XNOR U10495 ( .A(n9309), .B(n9303), .Z(c[1668]) );
  NAND U10496 ( .A(b[0]), .B(a[647]), .Z(n9312) );
  NAND U10497 ( .A(a[646]), .B(b[1]), .Z(n9311) );
  XNOR U10498 ( .A(n9312), .B(n9311), .Z(n9314) );
  XNOR U10499 ( .A(n9313), .B(n9314), .Z(n9318) );
  XOR U10500 ( .A(n9317), .B(sreg[1669]), .Z(n9310) );
  XNOR U10501 ( .A(n9318), .B(n9310), .Z(c[1669]) );
  NAND U10502 ( .A(n9312), .B(n9311), .Z(n9316) );
  NANDN U10503 ( .A(n9314), .B(n9313), .Z(n9315) );
  NAND U10504 ( .A(n9316), .B(n9315), .Z(n9323) );
  ANDN U10505 ( .B(a[648]), .A(n3961), .Z(n9321) );
  AND U10506 ( .A(b[1]), .B(a[647]), .Z(n9320) );
  XOR U10507 ( .A(n9321), .B(n9320), .Z(n9322) );
  XNOR U10508 ( .A(n9323), .B(n9322), .Z(n9325) );
  XOR U10509 ( .A(sreg[1670]), .B(n9324), .Z(n9319) );
  XNOR U10510 ( .A(n9325), .B(n9319), .Z(c[1670]) );
  ANDN U10511 ( .B(a[649]), .A(n3961), .Z(n9328) );
  AND U10512 ( .A(b[1]), .B(a[648]), .Z(n9327) );
  XOR U10513 ( .A(n9328), .B(n9327), .Z(n9329) );
  XNOR U10514 ( .A(n9330), .B(n9329), .Z(n9332) );
  XNOR U10515 ( .A(sreg[1671]), .B(n9331), .Z(n9326) );
  XNOR U10516 ( .A(n9332), .B(n9326), .Z(c[1671]) );
  ANDN U10517 ( .B(a[650]), .A(n3962), .Z(n9335) );
  AND U10518 ( .A(b[1]), .B(a[649]), .Z(n9334) );
  XOR U10519 ( .A(n9335), .B(n9334), .Z(n9336) );
  XNOR U10520 ( .A(n9337), .B(n9336), .Z(n9342) );
  XNOR U10521 ( .A(sreg[1672]), .B(n9341), .Z(n9333) );
  XNOR U10522 ( .A(n9342), .B(n9333), .Z(c[1672]) );
  OR U10523 ( .A(n9335), .B(n9334), .Z(n9340) );
  IV U10524 ( .A(n9336), .Z(n9338) );
  NANDN U10525 ( .A(n9338), .B(n9337), .Z(n9339) );
  NAND U10526 ( .A(n9340), .B(n9339), .Z(n9346) );
  NAND U10527 ( .A(b[0]), .B(a[651]), .Z(n9345) );
  NAND U10528 ( .A(a[650]), .B(b[1]), .Z(n9344) );
  XNOR U10529 ( .A(n9345), .B(n9344), .Z(n9347) );
  XNOR U10530 ( .A(n9346), .B(n9347), .Z(n9351) );
  XOR U10531 ( .A(n9350), .B(sreg[1673]), .Z(n9343) );
  XNOR U10532 ( .A(n9351), .B(n9343), .Z(c[1673]) );
  NAND U10533 ( .A(n9345), .B(n9344), .Z(n9349) );
  NANDN U10534 ( .A(n9347), .B(n9346), .Z(n9348) );
  NAND U10535 ( .A(n9349), .B(n9348), .Z(n9356) );
  ANDN U10536 ( .B(a[652]), .A(n3962), .Z(n9354) );
  AND U10537 ( .A(b[1]), .B(a[651]), .Z(n9353) );
  XOR U10538 ( .A(n9354), .B(n9353), .Z(n9355) );
  XNOR U10539 ( .A(n9356), .B(n9355), .Z(n9358) );
  XOR U10540 ( .A(sreg[1674]), .B(n9357), .Z(n9352) );
  XNOR U10541 ( .A(n9358), .B(n9352), .Z(c[1674]) );
  NAND U10542 ( .A(b[0]), .B(a[653]), .Z(n9361) );
  NAND U10543 ( .A(a[652]), .B(b[1]), .Z(n9360) );
  XNOR U10544 ( .A(n9361), .B(n9360), .Z(n9363) );
  XNOR U10545 ( .A(n9362), .B(n9363), .Z(n9367) );
  XOR U10546 ( .A(n9366), .B(sreg[1675]), .Z(n9359) );
  XNOR U10547 ( .A(n9367), .B(n9359), .Z(c[1675]) );
  NAND U10548 ( .A(n9361), .B(n9360), .Z(n9365) );
  NANDN U10549 ( .A(n9363), .B(n9362), .Z(n9364) );
  NAND U10550 ( .A(n9365), .B(n9364), .Z(n9372) );
  ANDN U10551 ( .B(a[654]), .A(n3962), .Z(n9370) );
  AND U10552 ( .A(b[1]), .B(a[653]), .Z(n9369) );
  XOR U10553 ( .A(n9370), .B(n9369), .Z(n9371) );
  XNOR U10554 ( .A(n9372), .B(n9371), .Z(n9374) );
  XOR U10555 ( .A(sreg[1676]), .B(n9373), .Z(n9368) );
  XNOR U10556 ( .A(n9374), .B(n9368), .Z(c[1676]) );
  NAND U10557 ( .A(b[0]), .B(a[655]), .Z(n9377) );
  NAND U10558 ( .A(a[654]), .B(b[1]), .Z(n9376) );
  XNOR U10559 ( .A(n9377), .B(n9376), .Z(n9379) );
  XNOR U10560 ( .A(n9378), .B(n9379), .Z(n9383) );
  XOR U10561 ( .A(n9382), .B(sreg[1677]), .Z(n9375) );
  XNOR U10562 ( .A(n9383), .B(n9375), .Z(c[1677]) );
  NAND U10563 ( .A(n9377), .B(n9376), .Z(n9381) );
  NANDN U10564 ( .A(n9379), .B(n9378), .Z(n9380) );
  NAND U10565 ( .A(n9381), .B(n9380), .Z(n9388) );
  ANDN U10566 ( .B(a[656]), .A(n3962), .Z(n9386) );
  AND U10567 ( .A(b[1]), .B(a[655]), .Z(n9385) );
  XOR U10568 ( .A(n9386), .B(n9385), .Z(n9387) );
  XNOR U10569 ( .A(n9388), .B(n9387), .Z(n9390) );
  XOR U10570 ( .A(sreg[1678]), .B(n9389), .Z(n9384) );
  XNOR U10571 ( .A(n9390), .B(n9384), .Z(c[1678]) );
  NAND U10572 ( .A(b[0]), .B(a[657]), .Z(n9393) );
  NAND U10573 ( .A(a[656]), .B(b[1]), .Z(n9392) );
  XNOR U10574 ( .A(n9393), .B(n9392), .Z(n9395) );
  XNOR U10575 ( .A(n9394), .B(n9395), .Z(n9399) );
  XOR U10576 ( .A(n9398), .B(sreg[1679]), .Z(n9391) );
  XNOR U10577 ( .A(n9399), .B(n9391), .Z(c[1679]) );
  NAND U10578 ( .A(n9393), .B(n9392), .Z(n9397) );
  NANDN U10579 ( .A(n9395), .B(n9394), .Z(n9396) );
  NAND U10580 ( .A(n9397), .B(n9396), .Z(n9404) );
  ANDN U10581 ( .B(a[658]), .A(n3962), .Z(n9402) );
  AND U10582 ( .A(b[1]), .B(a[657]), .Z(n9401) );
  XOR U10583 ( .A(n9402), .B(n9401), .Z(n9403) );
  XNOR U10584 ( .A(n9404), .B(n9403), .Z(n9406) );
  XOR U10585 ( .A(sreg[1680]), .B(n9405), .Z(n9400) );
  XNOR U10586 ( .A(n9406), .B(n9400), .Z(c[1680]) );
  ANDN U10587 ( .B(a[659]), .A(n3962), .Z(n9409) );
  AND U10588 ( .A(b[1]), .B(a[658]), .Z(n9408) );
  XOR U10589 ( .A(n9409), .B(n9408), .Z(n9410) );
  XNOR U10590 ( .A(n9411), .B(n9410), .Z(n9413) );
  XNOR U10591 ( .A(sreg[1681]), .B(n9412), .Z(n9407) );
  XNOR U10592 ( .A(n9413), .B(n9407), .Z(c[1681]) );
  ANDN U10593 ( .B(a[660]), .A(n3962), .Z(n9416) );
  AND U10594 ( .A(b[1]), .B(a[659]), .Z(n9415) );
  XOR U10595 ( .A(n9416), .B(n9415), .Z(n9417) );
  XNOR U10596 ( .A(n9418), .B(n9417), .Z(n9420) );
  XNOR U10597 ( .A(sreg[1682]), .B(n9419), .Z(n9414) );
  XNOR U10598 ( .A(n9420), .B(n9414), .Z(c[1682]) );
  ANDN U10599 ( .B(a[661]), .A(n3963), .Z(n9423) );
  AND U10600 ( .A(b[1]), .B(a[660]), .Z(n9422) );
  XOR U10601 ( .A(n9423), .B(n9422), .Z(n9424) );
  XNOR U10602 ( .A(n9425), .B(n9424), .Z(n9430) );
  XNOR U10603 ( .A(sreg[1683]), .B(n9429), .Z(n9421) );
  XNOR U10604 ( .A(n9430), .B(n9421), .Z(c[1683]) );
  OR U10605 ( .A(n9423), .B(n9422), .Z(n9428) );
  IV U10606 ( .A(n9424), .Z(n9426) );
  NANDN U10607 ( .A(n9426), .B(n9425), .Z(n9427) );
  NAND U10608 ( .A(n9428), .B(n9427), .Z(n9435) );
  ANDN U10609 ( .B(a[662]), .A(n3963), .Z(n9433) );
  AND U10610 ( .A(b[1]), .B(a[661]), .Z(n9432) );
  XOR U10611 ( .A(n9433), .B(n9432), .Z(n9434) );
  XNOR U10612 ( .A(n9435), .B(n9434), .Z(n9437) );
  XNOR U10613 ( .A(sreg[1684]), .B(n9436), .Z(n9431) );
  XNOR U10614 ( .A(n9437), .B(n9431), .Z(c[1684]) );
  NAND U10615 ( .A(b[0]), .B(a[663]), .Z(n9440) );
  NAND U10616 ( .A(a[662]), .B(b[1]), .Z(n9439) );
  XNOR U10617 ( .A(n9440), .B(n9439), .Z(n9442) );
  XNOR U10618 ( .A(n9441), .B(n9442), .Z(n9446) );
  XOR U10619 ( .A(n9445), .B(sreg[1685]), .Z(n9438) );
  XNOR U10620 ( .A(n9446), .B(n9438), .Z(c[1685]) );
  NAND U10621 ( .A(n9440), .B(n9439), .Z(n9444) );
  NANDN U10622 ( .A(n9442), .B(n9441), .Z(n9443) );
  NAND U10623 ( .A(n9444), .B(n9443), .Z(n9451) );
  ANDN U10624 ( .B(a[664]), .A(n3963), .Z(n9449) );
  AND U10625 ( .A(b[1]), .B(a[663]), .Z(n9448) );
  XOR U10626 ( .A(n9449), .B(n9448), .Z(n9450) );
  XNOR U10627 ( .A(n9451), .B(n9450), .Z(n9453) );
  XOR U10628 ( .A(sreg[1686]), .B(n9452), .Z(n9447) );
  XNOR U10629 ( .A(n9453), .B(n9447), .Z(c[1686]) );
  NAND U10630 ( .A(b[0]), .B(a[665]), .Z(n9456) );
  NAND U10631 ( .A(a[664]), .B(b[1]), .Z(n9455) );
  XNOR U10632 ( .A(n9456), .B(n9455), .Z(n9458) );
  XNOR U10633 ( .A(n9457), .B(n9458), .Z(n9462) );
  XOR U10634 ( .A(n9461), .B(sreg[1687]), .Z(n9454) );
  XNOR U10635 ( .A(n9462), .B(n9454), .Z(c[1687]) );
  NAND U10636 ( .A(n9456), .B(n9455), .Z(n9460) );
  NANDN U10637 ( .A(n9458), .B(n9457), .Z(n9459) );
  NAND U10638 ( .A(n9460), .B(n9459), .Z(n9467) );
  ANDN U10639 ( .B(a[666]), .A(n3963), .Z(n9465) );
  AND U10640 ( .A(b[1]), .B(a[665]), .Z(n9464) );
  XOR U10641 ( .A(n9465), .B(n9464), .Z(n9466) );
  XNOR U10642 ( .A(n9467), .B(n9466), .Z(n9469) );
  XOR U10643 ( .A(sreg[1688]), .B(n9468), .Z(n9463) );
  XNOR U10644 ( .A(n9469), .B(n9463), .Z(c[1688]) );
  NAND U10645 ( .A(b[0]), .B(a[667]), .Z(n9472) );
  NAND U10646 ( .A(a[666]), .B(b[1]), .Z(n9471) );
  XNOR U10647 ( .A(n9472), .B(n9471), .Z(n9474) );
  XNOR U10648 ( .A(n9473), .B(n9474), .Z(n9478) );
  XOR U10649 ( .A(n9477), .B(sreg[1689]), .Z(n9470) );
  XNOR U10650 ( .A(n9478), .B(n9470), .Z(c[1689]) );
  NAND U10651 ( .A(n9472), .B(n9471), .Z(n9476) );
  NANDN U10652 ( .A(n9474), .B(n9473), .Z(n9475) );
  NAND U10653 ( .A(n9476), .B(n9475), .Z(n9483) );
  ANDN U10654 ( .B(a[668]), .A(n3963), .Z(n9481) );
  AND U10655 ( .A(b[1]), .B(a[667]), .Z(n9480) );
  XOR U10656 ( .A(n9481), .B(n9480), .Z(n9482) );
  XNOR U10657 ( .A(n9483), .B(n9482), .Z(n9485) );
  XOR U10658 ( .A(sreg[1690]), .B(n9484), .Z(n9479) );
  XNOR U10659 ( .A(n9485), .B(n9479), .Z(c[1690]) );
  NAND U10660 ( .A(b[0]), .B(a[669]), .Z(n9488) );
  NAND U10661 ( .A(a[668]), .B(b[1]), .Z(n9487) );
  XNOR U10662 ( .A(n9488), .B(n9487), .Z(n9490) );
  XNOR U10663 ( .A(n9489), .B(n9490), .Z(n9494) );
  XOR U10664 ( .A(n9493), .B(sreg[1691]), .Z(n9486) );
  XNOR U10665 ( .A(n9494), .B(n9486), .Z(c[1691]) );
  NAND U10666 ( .A(n9488), .B(n9487), .Z(n9492) );
  NANDN U10667 ( .A(n9490), .B(n9489), .Z(n9491) );
  NAND U10668 ( .A(n9492), .B(n9491), .Z(n9498) );
  NAND U10669 ( .A(b[0]), .B(a[670]), .Z(n9497) );
  NAND U10670 ( .A(a[669]), .B(b[1]), .Z(n9496) );
  XNOR U10671 ( .A(n9497), .B(n9496), .Z(n9499) );
  XNOR U10672 ( .A(n9498), .B(n9499), .Z(n9503) );
  XOR U10673 ( .A(n9502), .B(sreg[1692]), .Z(n9495) );
  XNOR U10674 ( .A(n9503), .B(n9495), .Z(c[1692]) );
  NAND U10675 ( .A(n9497), .B(n9496), .Z(n9501) );
  NANDN U10676 ( .A(n9499), .B(n9498), .Z(n9500) );
  NAND U10677 ( .A(n9501), .B(n9500), .Z(n9507) );
  NAND U10678 ( .A(b[0]), .B(a[671]), .Z(n9506) );
  NAND U10679 ( .A(a[670]), .B(b[1]), .Z(n9505) );
  XNOR U10680 ( .A(n9506), .B(n9505), .Z(n9508) );
  XNOR U10681 ( .A(n9507), .B(n9508), .Z(n9512) );
  XOR U10682 ( .A(n9511), .B(sreg[1693]), .Z(n9504) );
  XNOR U10683 ( .A(n9512), .B(n9504), .Z(c[1693]) );
  NAND U10684 ( .A(n9506), .B(n9505), .Z(n9510) );
  NANDN U10685 ( .A(n9508), .B(n9507), .Z(n9509) );
  NAND U10686 ( .A(n9510), .B(n9509), .Z(n9517) );
  ANDN U10687 ( .B(a[672]), .A(n3963), .Z(n9515) );
  AND U10688 ( .A(b[1]), .B(a[671]), .Z(n9514) );
  XOR U10689 ( .A(n9515), .B(n9514), .Z(n9516) );
  XNOR U10690 ( .A(n9517), .B(n9516), .Z(n9519) );
  XOR U10691 ( .A(sreg[1694]), .B(n9518), .Z(n9513) );
  XNOR U10692 ( .A(n9519), .B(n9513), .Z(c[1694]) );
  NAND U10693 ( .A(b[0]), .B(a[673]), .Z(n9522) );
  NAND U10694 ( .A(a[672]), .B(b[1]), .Z(n9521) );
  XNOR U10695 ( .A(n9522), .B(n9521), .Z(n9524) );
  XNOR U10696 ( .A(n9523), .B(n9524), .Z(n9528) );
  XOR U10697 ( .A(n9527), .B(sreg[1695]), .Z(n9520) );
  XNOR U10698 ( .A(n9528), .B(n9520), .Z(c[1695]) );
  NAND U10699 ( .A(n9522), .B(n9521), .Z(n9526) );
  NANDN U10700 ( .A(n9524), .B(n9523), .Z(n9525) );
  NAND U10701 ( .A(n9526), .B(n9525), .Z(n9533) );
  ANDN U10702 ( .B(a[674]), .A(n3963), .Z(n9531) );
  AND U10703 ( .A(b[1]), .B(a[673]), .Z(n9530) );
  XOR U10704 ( .A(n9531), .B(n9530), .Z(n9532) );
  XNOR U10705 ( .A(n9533), .B(n9532), .Z(n9535) );
  XOR U10706 ( .A(sreg[1696]), .B(n9534), .Z(n9529) );
  XNOR U10707 ( .A(n9535), .B(n9529), .Z(c[1696]) );
  ANDN U10708 ( .B(a[675]), .A(n3964), .Z(n9538) );
  AND U10709 ( .A(b[1]), .B(a[674]), .Z(n9537) );
  XOR U10710 ( .A(n9538), .B(n9537), .Z(n9539) );
  XNOR U10711 ( .A(n9540), .B(n9539), .Z(n9545) );
  XNOR U10712 ( .A(sreg[1697]), .B(n9544), .Z(n9536) );
  XNOR U10713 ( .A(n9545), .B(n9536), .Z(c[1697]) );
  OR U10714 ( .A(n9538), .B(n9537), .Z(n9543) );
  IV U10715 ( .A(n9539), .Z(n9541) );
  NANDN U10716 ( .A(n9541), .B(n9540), .Z(n9542) );
  NAND U10717 ( .A(n9543), .B(n9542), .Z(n9550) );
  ANDN U10718 ( .B(a[676]), .A(n3964), .Z(n9548) );
  AND U10719 ( .A(b[1]), .B(a[675]), .Z(n9547) );
  XOR U10720 ( .A(n9548), .B(n9547), .Z(n9549) );
  XNOR U10721 ( .A(n9550), .B(n9549), .Z(n9552) );
  XNOR U10722 ( .A(sreg[1698]), .B(n9551), .Z(n9546) );
  XNOR U10723 ( .A(n9552), .B(n9546), .Z(c[1698]) );
  NAND U10724 ( .A(b[0]), .B(a[677]), .Z(n9555) );
  NAND U10725 ( .A(a[676]), .B(b[1]), .Z(n9554) );
  XNOR U10726 ( .A(n9555), .B(n9554), .Z(n9557) );
  XNOR U10727 ( .A(n9556), .B(n9557), .Z(n9561) );
  XOR U10728 ( .A(n9560), .B(sreg[1699]), .Z(n9553) );
  XNOR U10729 ( .A(n9561), .B(n9553), .Z(c[1699]) );
  NAND U10730 ( .A(n9555), .B(n9554), .Z(n9559) );
  NANDN U10731 ( .A(n9557), .B(n9556), .Z(n9558) );
  NAND U10732 ( .A(n9559), .B(n9558), .Z(n9566) );
  ANDN U10733 ( .B(a[678]), .A(n3964), .Z(n9564) );
  AND U10734 ( .A(b[1]), .B(a[677]), .Z(n9563) );
  XOR U10735 ( .A(n9564), .B(n9563), .Z(n9565) );
  XNOR U10736 ( .A(n9566), .B(n9565), .Z(n9568) );
  XOR U10737 ( .A(sreg[1700]), .B(n9567), .Z(n9562) );
  XNOR U10738 ( .A(n9568), .B(n9562), .Z(c[1700]) );
  NAND U10739 ( .A(b[0]), .B(a[679]), .Z(n9571) );
  NAND U10740 ( .A(a[678]), .B(b[1]), .Z(n9570) );
  XNOR U10741 ( .A(n9571), .B(n9570), .Z(n9573) );
  XNOR U10742 ( .A(n9572), .B(n9573), .Z(n9577) );
  XOR U10743 ( .A(n9576), .B(sreg[1701]), .Z(n9569) );
  XNOR U10744 ( .A(n9577), .B(n9569), .Z(c[1701]) );
  NAND U10745 ( .A(n9571), .B(n9570), .Z(n9575) );
  NANDN U10746 ( .A(n9573), .B(n9572), .Z(n9574) );
  NAND U10747 ( .A(n9575), .B(n9574), .Z(n9582) );
  ANDN U10748 ( .B(a[680]), .A(n3964), .Z(n9580) );
  AND U10749 ( .A(b[1]), .B(a[679]), .Z(n9579) );
  XOR U10750 ( .A(n9580), .B(n9579), .Z(n9581) );
  XNOR U10751 ( .A(n9582), .B(n9581), .Z(n9584) );
  XOR U10752 ( .A(sreg[1702]), .B(n9583), .Z(n9578) );
  XNOR U10753 ( .A(n9584), .B(n9578), .Z(c[1702]) );
  NAND U10754 ( .A(b[0]), .B(a[681]), .Z(n9587) );
  NAND U10755 ( .A(a[680]), .B(b[1]), .Z(n9586) );
  XNOR U10756 ( .A(n9587), .B(n9586), .Z(n9589) );
  XNOR U10757 ( .A(n9588), .B(n9589), .Z(n9593) );
  XOR U10758 ( .A(n9592), .B(sreg[1703]), .Z(n9585) );
  XNOR U10759 ( .A(n9593), .B(n9585), .Z(c[1703]) );
  NAND U10760 ( .A(n9587), .B(n9586), .Z(n9591) );
  NANDN U10761 ( .A(n9589), .B(n9588), .Z(n9590) );
  NAND U10762 ( .A(n9591), .B(n9590), .Z(n9598) );
  ANDN U10763 ( .B(a[682]), .A(n3964), .Z(n9596) );
  AND U10764 ( .A(b[1]), .B(a[681]), .Z(n9595) );
  XOR U10765 ( .A(n9596), .B(n9595), .Z(n9597) );
  XNOR U10766 ( .A(n9598), .B(n9597), .Z(n9600) );
  XOR U10767 ( .A(sreg[1704]), .B(n9599), .Z(n9594) );
  XNOR U10768 ( .A(n9600), .B(n9594), .Z(c[1704]) );
  NAND U10769 ( .A(b[0]), .B(a[683]), .Z(n9603) );
  NAND U10770 ( .A(a[682]), .B(b[1]), .Z(n9602) );
  XNOR U10771 ( .A(n9603), .B(n9602), .Z(n9605) );
  XNOR U10772 ( .A(n9604), .B(n9605), .Z(n9609) );
  XOR U10773 ( .A(n9608), .B(sreg[1705]), .Z(n9601) );
  XNOR U10774 ( .A(n9609), .B(n9601), .Z(c[1705]) );
  NAND U10775 ( .A(n9603), .B(n9602), .Z(n9607) );
  NANDN U10776 ( .A(n9605), .B(n9604), .Z(n9606) );
  NAND U10777 ( .A(n9607), .B(n9606), .Z(n9613) );
  NAND U10778 ( .A(b[0]), .B(a[684]), .Z(n9612) );
  NAND U10779 ( .A(a[683]), .B(b[1]), .Z(n9611) );
  XNOR U10780 ( .A(n9612), .B(n9611), .Z(n9614) );
  XNOR U10781 ( .A(n9613), .B(n9614), .Z(n9618) );
  XOR U10782 ( .A(n9617), .B(sreg[1706]), .Z(n9610) );
  XNOR U10783 ( .A(n9618), .B(n9610), .Z(c[1706]) );
  NAND U10784 ( .A(n9612), .B(n9611), .Z(n9616) );
  NANDN U10785 ( .A(n9614), .B(n9613), .Z(n9615) );
  NAND U10786 ( .A(n9616), .B(n9615), .Z(n9622) );
  NAND U10787 ( .A(b[0]), .B(a[685]), .Z(n9621) );
  NAND U10788 ( .A(a[684]), .B(b[1]), .Z(n9620) );
  XNOR U10789 ( .A(n9621), .B(n9620), .Z(n9623) );
  XNOR U10790 ( .A(n9622), .B(n9623), .Z(n9627) );
  XOR U10791 ( .A(n9626), .B(sreg[1707]), .Z(n9619) );
  XNOR U10792 ( .A(n9627), .B(n9619), .Z(c[1707]) );
  NAND U10793 ( .A(n9621), .B(n9620), .Z(n9625) );
  NANDN U10794 ( .A(n9623), .B(n9622), .Z(n9624) );
  NAND U10795 ( .A(n9625), .B(n9624), .Z(n9632) );
  ANDN U10796 ( .B(a[686]), .A(n3964), .Z(n9630) );
  AND U10797 ( .A(b[1]), .B(a[685]), .Z(n9629) );
  XOR U10798 ( .A(n9630), .B(n9629), .Z(n9631) );
  XNOR U10799 ( .A(n9632), .B(n9631), .Z(n9634) );
  XOR U10800 ( .A(sreg[1708]), .B(n9633), .Z(n9628) );
  XNOR U10801 ( .A(n9634), .B(n9628), .Z(c[1708]) );
  NAND U10802 ( .A(b[0]), .B(a[687]), .Z(n9637) );
  NAND U10803 ( .A(a[686]), .B(b[1]), .Z(n9636) );
  XNOR U10804 ( .A(n9637), .B(n9636), .Z(n9639) );
  XNOR U10805 ( .A(n9638), .B(n9639), .Z(n9643) );
  XOR U10806 ( .A(n9642), .B(sreg[1709]), .Z(n9635) );
  XNOR U10807 ( .A(n9643), .B(n9635), .Z(c[1709]) );
  NAND U10808 ( .A(n9637), .B(n9636), .Z(n9641) );
  NANDN U10809 ( .A(n9639), .B(n9638), .Z(n9640) );
  NAND U10810 ( .A(n9641), .B(n9640), .Z(n9648) );
  ANDN U10811 ( .B(a[688]), .A(n3964), .Z(n9646) );
  AND U10812 ( .A(b[1]), .B(a[687]), .Z(n9645) );
  XOR U10813 ( .A(n9646), .B(n9645), .Z(n9647) );
  XNOR U10814 ( .A(n9648), .B(n9647), .Z(n9650) );
  XOR U10815 ( .A(sreg[1710]), .B(n9649), .Z(n9644) );
  XNOR U10816 ( .A(n9650), .B(n9644), .Z(c[1710]) );
  NAND U10817 ( .A(b[0]), .B(a[689]), .Z(n9653) );
  NAND U10818 ( .A(a[688]), .B(b[1]), .Z(n9652) );
  XNOR U10819 ( .A(n9653), .B(n9652), .Z(n9655) );
  XNOR U10820 ( .A(n9654), .B(n9655), .Z(n9659) );
  XOR U10821 ( .A(n9658), .B(sreg[1711]), .Z(n9651) );
  XNOR U10822 ( .A(n9659), .B(n9651), .Z(c[1711]) );
  NAND U10823 ( .A(n9653), .B(n9652), .Z(n9657) );
  NANDN U10824 ( .A(n9655), .B(n9654), .Z(n9656) );
  NAND U10825 ( .A(n9657), .B(n9656), .Z(n9664) );
  ANDN U10826 ( .B(a[690]), .A(n3965), .Z(n9662) );
  AND U10827 ( .A(b[1]), .B(a[689]), .Z(n9661) );
  XOR U10828 ( .A(n9662), .B(n9661), .Z(n9663) );
  XNOR U10829 ( .A(n9664), .B(n9663), .Z(n9669) );
  XOR U10830 ( .A(sreg[1712]), .B(n9668), .Z(n9660) );
  XNOR U10831 ( .A(n9669), .B(n9660), .Z(c[1712]) );
  OR U10832 ( .A(n9662), .B(n9661), .Z(n9667) );
  IV U10833 ( .A(n9663), .Z(n9665) );
  NANDN U10834 ( .A(n9665), .B(n9664), .Z(n9666) );
  NAND U10835 ( .A(n9667), .B(n9666), .Z(n9673) );
  NAND U10836 ( .A(b[0]), .B(a[691]), .Z(n9672) );
  NAND U10837 ( .A(a[690]), .B(b[1]), .Z(n9671) );
  XNOR U10838 ( .A(n9672), .B(n9671), .Z(n9674) );
  XNOR U10839 ( .A(n9673), .B(n9674), .Z(n9678) );
  XOR U10840 ( .A(n9677), .B(sreg[1713]), .Z(n9670) );
  XNOR U10841 ( .A(n9678), .B(n9670), .Z(c[1713]) );
  NAND U10842 ( .A(n9672), .B(n9671), .Z(n9676) );
  NANDN U10843 ( .A(n9674), .B(n9673), .Z(n9675) );
  NAND U10844 ( .A(n9676), .B(n9675), .Z(n9683) );
  ANDN U10845 ( .B(a[692]), .A(n3965), .Z(n9681) );
  AND U10846 ( .A(b[1]), .B(a[691]), .Z(n9680) );
  XOR U10847 ( .A(n9681), .B(n9680), .Z(n9682) );
  XNOR U10848 ( .A(n9683), .B(n9682), .Z(n9685) );
  XOR U10849 ( .A(sreg[1714]), .B(n9684), .Z(n9679) );
  XNOR U10850 ( .A(n9685), .B(n9679), .Z(c[1714]) );
  NAND U10851 ( .A(b[0]), .B(a[693]), .Z(n9688) );
  NAND U10852 ( .A(a[692]), .B(b[1]), .Z(n9687) );
  XNOR U10853 ( .A(n9688), .B(n9687), .Z(n9690) );
  XNOR U10854 ( .A(n9689), .B(n9690), .Z(n9694) );
  XOR U10855 ( .A(n9693), .B(sreg[1715]), .Z(n9686) );
  XNOR U10856 ( .A(n9694), .B(n9686), .Z(c[1715]) );
  NAND U10857 ( .A(n9688), .B(n9687), .Z(n9692) );
  NANDN U10858 ( .A(n9690), .B(n9689), .Z(n9691) );
  NAND U10859 ( .A(n9692), .B(n9691), .Z(n9699) );
  ANDN U10860 ( .B(a[694]), .A(n3965), .Z(n9697) );
  AND U10861 ( .A(b[1]), .B(a[693]), .Z(n9696) );
  XOR U10862 ( .A(n9697), .B(n9696), .Z(n9698) );
  XNOR U10863 ( .A(n9699), .B(n9698), .Z(n9701) );
  XOR U10864 ( .A(sreg[1716]), .B(n9700), .Z(n9695) );
  XNOR U10865 ( .A(n9701), .B(n9695), .Z(c[1716]) );
  NAND U10866 ( .A(b[0]), .B(a[695]), .Z(n9704) );
  NAND U10867 ( .A(a[694]), .B(b[1]), .Z(n9703) );
  XNOR U10868 ( .A(n9704), .B(n9703), .Z(n9706) );
  XNOR U10869 ( .A(n9705), .B(n9706), .Z(n9710) );
  XOR U10870 ( .A(n9709), .B(sreg[1717]), .Z(n9702) );
  XNOR U10871 ( .A(n9710), .B(n9702), .Z(c[1717]) );
  NAND U10872 ( .A(n9704), .B(n9703), .Z(n9708) );
  NANDN U10873 ( .A(n9706), .B(n9705), .Z(n9707) );
  NAND U10874 ( .A(n9708), .B(n9707), .Z(n9715) );
  ANDN U10875 ( .B(a[696]), .A(n3965), .Z(n9713) );
  AND U10876 ( .A(b[1]), .B(a[695]), .Z(n9712) );
  XOR U10877 ( .A(n9713), .B(n9712), .Z(n9714) );
  XNOR U10878 ( .A(n9715), .B(n9714), .Z(n9717) );
  XOR U10879 ( .A(sreg[1718]), .B(n9716), .Z(n9711) );
  XNOR U10880 ( .A(n9717), .B(n9711), .Z(c[1718]) );
  NAND U10881 ( .A(b[0]), .B(a[697]), .Z(n9720) );
  NAND U10882 ( .A(a[696]), .B(b[1]), .Z(n9719) );
  XNOR U10883 ( .A(n9720), .B(n9719), .Z(n9722) );
  XNOR U10884 ( .A(n9721), .B(n9722), .Z(n9726) );
  XOR U10885 ( .A(n9725), .B(sreg[1719]), .Z(n9718) );
  XNOR U10886 ( .A(n9726), .B(n9718), .Z(c[1719]) );
  NAND U10887 ( .A(n9720), .B(n9719), .Z(n9724) );
  NANDN U10888 ( .A(n9722), .B(n9721), .Z(n9723) );
  NAND U10889 ( .A(n9724), .B(n9723), .Z(n9731) );
  ANDN U10890 ( .B(a[698]), .A(n3965), .Z(n9729) );
  AND U10891 ( .A(b[1]), .B(a[697]), .Z(n9728) );
  XOR U10892 ( .A(n9729), .B(n9728), .Z(n9730) );
  XNOR U10893 ( .A(n9731), .B(n9730), .Z(n9733) );
  XOR U10894 ( .A(sreg[1720]), .B(n9732), .Z(n9727) );
  XNOR U10895 ( .A(n9733), .B(n9727), .Z(c[1720]) );
  ANDN U10896 ( .B(a[699]), .A(n3965), .Z(n9736) );
  AND U10897 ( .A(b[1]), .B(a[698]), .Z(n9735) );
  XOR U10898 ( .A(n9736), .B(n9735), .Z(n9737) );
  XNOR U10899 ( .A(n9738), .B(n9737), .Z(n9740) );
  XNOR U10900 ( .A(sreg[1721]), .B(n9739), .Z(n9734) );
  XNOR U10901 ( .A(n9740), .B(n9734), .Z(c[1721]) );
  ANDN U10902 ( .B(a[700]), .A(n3965), .Z(n9743) );
  AND U10903 ( .A(b[1]), .B(a[699]), .Z(n9742) );
  XOR U10904 ( .A(n9743), .B(n9742), .Z(n9744) );
  XNOR U10905 ( .A(n9745), .B(n9744), .Z(n9747) );
  XNOR U10906 ( .A(sreg[1722]), .B(n9746), .Z(n9741) );
  XNOR U10907 ( .A(n9747), .B(n9741), .Z(c[1722]) );
  NAND U10908 ( .A(b[0]), .B(a[701]), .Z(n9750) );
  NAND U10909 ( .A(a[700]), .B(b[1]), .Z(n9749) );
  XNOR U10910 ( .A(n9750), .B(n9749), .Z(n9752) );
  XNOR U10911 ( .A(n9751), .B(n9752), .Z(n9756) );
  XOR U10912 ( .A(n9755), .B(sreg[1723]), .Z(n9748) );
  XNOR U10913 ( .A(n9756), .B(n9748), .Z(c[1723]) );
  NAND U10914 ( .A(n9750), .B(n9749), .Z(n9754) );
  NANDN U10915 ( .A(n9752), .B(n9751), .Z(n9753) );
  NAND U10916 ( .A(n9754), .B(n9753), .Z(n9761) );
  ANDN U10917 ( .B(a[702]), .A(n3966), .Z(n9759) );
  AND U10918 ( .A(b[1]), .B(a[701]), .Z(n9758) );
  XOR U10919 ( .A(n9759), .B(n9758), .Z(n9760) );
  XNOR U10920 ( .A(n9761), .B(n9760), .Z(n9766) );
  XOR U10921 ( .A(sreg[1724]), .B(n9765), .Z(n9757) );
  XNOR U10922 ( .A(n9766), .B(n9757), .Z(c[1724]) );
  OR U10923 ( .A(n9759), .B(n9758), .Z(n9764) );
  IV U10924 ( .A(n9760), .Z(n9762) );
  NANDN U10925 ( .A(n9762), .B(n9761), .Z(n9763) );
  NAND U10926 ( .A(n9764), .B(n9763), .Z(n9770) );
  NAND U10927 ( .A(b[0]), .B(a[703]), .Z(n9769) );
  NAND U10928 ( .A(a[702]), .B(b[1]), .Z(n9768) );
  XNOR U10929 ( .A(n9769), .B(n9768), .Z(n9771) );
  XNOR U10930 ( .A(n9770), .B(n9771), .Z(n9775) );
  XOR U10931 ( .A(n9774), .B(sreg[1725]), .Z(n9767) );
  XNOR U10932 ( .A(n9775), .B(n9767), .Z(c[1725]) );
  NAND U10933 ( .A(n9769), .B(n9768), .Z(n9773) );
  NANDN U10934 ( .A(n9771), .B(n9770), .Z(n9772) );
  NAND U10935 ( .A(n9773), .B(n9772), .Z(n9780) );
  ANDN U10936 ( .B(a[704]), .A(n3966), .Z(n9778) );
  AND U10937 ( .A(b[1]), .B(a[703]), .Z(n9777) );
  XOR U10938 ( .A(n9778), .B(n9777), .Z(n9779) );
  XNOR U10939 ( .A(n9780), .B(n9779), .Z(n9782) );
  XOR U10940 ( .A(sreg[1726]), .B(n9781), .Z(n9776) );
  XNOR U10941 ( .A(n9782), .B(n9776), .Z(c[1726]) );
  NAND U10942 ( .A(b[0]), .B(a[705]), .Z(n9785) );
  NAND U10943 ( .A(a[704]), .B(b[1]), .Z(n9784) );
  XNOR U10944 ( .A(n9785), .B(n9784), .Z(n9787) );
  XNOR U10945 ( .A(n9786), .B(n9787), .Z(n9791) );
  XOR U10946 ( .A(n9790), .B(sreg[1727]), .Z(n9783) );
  XNOR U10947 ( .A(n9791), .B(n9783), .Z(c[1727]) );
  NAND U10948 ( .A(n9785), .B(n9784), .Z(n9789) );
  NANDN U10949 ( .A(n9787), .B(n9786), .Z(n9788) );
  NAND U10950 ( .A(n9789), .B(n9788), .Z(n9796) );
  ANDN U10951 ( .B(a[706]), .A(n3966), .Z(n9794) );
  AND U10952 ( .A(b[1]), .B(a[705]), .Z(n9793) );
  XOR U10953 ( .A(n9794), .B(n9793), .Z(n9795) );
  XNOR U10954 ( .A(n9796), .B(n9795), .Z(n9798) );
  XOR U10955 ( .A(sreg[1728]), .B(n9797), .Z(n9792) );
  XNOR U10956 ( .A(n9798), .B(n9792), .Z(c[1728]) );
  NAND U10957 ( .A(b[0]), .B(a[707]), .Z(n9801) );
  NAND U10958 ( .A(a[706]), .B(b[1]), .Z(n9800) );
  XNOR U10959 ( .A(n9801), .B(n9800), .Z(n9803) );
  XNOR U10960 ( .A(n9802), .B(n9803), .Z(n9807) );
  XOR U10961 ( .A(n9806), .B(sreg[1729]), .Z(n9799) );
  XNOR U10962 ( .A(n9807), .B(n9799), .Z(c[1729]) );
  NAND U10963 ( .A(n9801), .B(n9800), .Z(n9805) );
  NANDN U10964 ( .A(n9803), .B(n9802), .Z(n9804) );
  NAND U10965 ( .A(n9805), .B(n9804), .Z(n9812) );
  ANDN U10966 ( .B(a[708]), .A(n3966), .Z(n9810) );
  AND U10967 ( .A(b[1]), .B(a[707]), .Z(n9809) );
  XOR U10968 ( .A(n9810), .B(n9809), .Z(n9811) );
  XNOR U10969 ( .A(n9812), .B(n9811), .Z(n9814) );
  XOR U10970 ( .A(sreg[1730]), .B(n9813), .Z(n9808) );
  XNOR U10971 ( .A(n9814), .B(n9808), .Z(c[1730]) );
  ANDN U10972 ( .B(a[709]), .A(n3966), .Z(n9817) );
  AND U10973 ( .A(b[1]), .B(a[708]), .Z(n9816) );
  XOR U10974 ( .A(n9817), .B(n9816), .Z(n9818) );
  XNOR U10975 ( .A(n9819), .B(n9818), .Z(n9821) );
  XNOR U10976 ( .A(sreg[1731]), .B(n9820), .Z(n9815) );
  XNOR U10977 ( .A(n9821), .B(n9815), .Z(c[1731]) );
  ANDN U10978 ( .B(a[710]), .A(n3966), .Z(n9824) );
  AND U10979 ( .A(b[1]), .B(a[709]), .Z(n9823) );
  XOR U10980 ( .A(n9824), .B(n9823), .Z(n9825) );
  XNOR U10981 ( .A(n9826), .B(n9825), .Z(n9828) );
  XNOR U10982 ( .A(sreg[1732]), .B(n9827), .Z(n9822) );
  XNOR U10983 ( .A(n9828), .B(n9822), .Z(c[1732]) );
  NAND U10984 ( .A(b[0]), .B(a[711]), .Z(n9831) );
  NAND U10985 ( .A(a[710]), .B(b[1]), .Z(n9830) );
  XNOR U10986 ( .A(n9831), .B(n9830), .Z(n9833) );
  XNOR U10987 ( .A(n9832), .B(n9833), .Z(n9837) );
  XOR U10988 ( .A(n9836), .B(sreg[1733]), .Z(n9829) );
  XNOR U10989 ( .A(n9837), .B(n9829), .Z(c[1733]) );
  NAND U10990 ( .A(n9831), .B(n9830), .Z(n9835) );
  NANDN U10991 ( .A(n9833), .B(n9832), .Z(n9834) );
  NAND U10992 ( .A(n9835), .B(n9834), .Z(n9842) );
  ANDN U10993 ( .B(a[712]), .A(n3966), .Z(n9840) );
  AND U10994 ( .A(b[1]), .B(a[711]), .Z(n9839) );
  XOR U10995 ( .A(n9840), .B(n9839), .Z(n9841) );
  XNOR U10996 ( .A(n9842), .B(n9841), .Z(n9844) );
  XOR U10997 ( .A(sreg[1734]), .B(n9843), .Z(n9838) );
  XNOR U10998 ( .A(n9844), .B(n9838), .Z(c[1734]) );
  NAND U10999 ( .A(b[0]), .B(a[713]), .Z(n9847) );
  NAND U11000 ( .A(a[712]), .B(b[1]), .Z(n9846) );
  XNOR U11001 ( .A(n9847), .B(n9846), .Z(n9849) );
  XNOR U11002 ( .A(n9848), .B(n9849), .Z(n9853) );
  XOR U11003 ( .A(n9852), .B(sreg[1735]), .Z(n9845) );
  XNOR U11004 ( .A(n9853), .B(n9845), .Z(c[1735]) );
  NAND U11005 ( .A(n9847), .B(n9846), .Z(n9851) );
  NANDN U11006 ( .A(n9849), .B(n9848), .Z(n9850) );
  NAND U11007 ( .A(n9851), .B(n9850), .Z(n9858) );
  ANDN U11008 ( .B(a[714]), .A(n3967), .Z(n9856) );
  AND U11009 ( .A(b[1]), .B(a[713]), .Z(n9855) );
  XOR U11010 ( .A(n9856), .B(n9855), .Z(n9857) );
  XNOR U11011 ( .A(n9858), .B(n9857), .Z(n9863) );
  XOR U11012 ( .A(sreg[1736]), .B(n9862), .Z(n9854) );
  XNOR U11013 ( .A(n9863), .B(n9854), .Z(c[1736]) );
  OR U11014 ( .A(n9856), .B(n9855), .Z(n9861) );
  IV U11015 ( .A(n9857), .Z(n9859) );
  NANDN U11016 ( .A(n9859), .B(n9858), .Z(n9860) );
  NAND U11017 ( .A(n9861), .B(n9860), .Z(n9867) );
  NAND U11018 ( .A(b[0]), .B(a[715]), .Z(n9866) );
  NAND U11019 ( .A(a[714]), .B(b[1]), .Z(n9865) );
  XNOR U11020 ( .A(n9866), .B(n9865), .Z(n9868) );
  XNOR U11021 ( .A(n9867), .B(n9868), .Z(n9872) );
  XOR U11022 ( .A(n9871), .B(sreg[1737]), .Z(n9864) );
  XNOR U11023 ( .A(n9872), .B(n9864), .Z(c[1737]) );
  NAND U11024 ( .A(n9866), .B(n9865), .Z(n9870) );
  NANDN U11025 ( .A(n9868), .B(n9867), .Z(n9869) );
  NAND U11026 ( .A(n9870), .B(n9869), .Z(n9877) );
  ANDN U11027 ( .B(a[716]), .A(n3967), .Z(n9875) );
  AND U11028 ( .A(b[1]), .B(a[715]), .Z(n9874) );
  XOR U11029 ( .A(n9875), .B(n9874), .Z(n9876) );
  XNOR U11030 ( .A(n9877), .B(n9876), .Z(n9879) );
  XOR U11031 ( .A(sreg[1738]), .B(n9878), .Z(n9873) );
  XNOR U11032 ( .A(n9879), .B(n9873), .Z(c[1738]) );
  NAND U11033 ( .A(b[0]), .B(a[717]), .Z(n9882) );
  NAND U11034 ( .A(a[716]), .B(b[1]), .Z(n9881) );
  XNOR U11035 ( .A(n9882), .B(n9881), .Z(n9884) );
  XNOR U11036 ( .A(n9883), .B(n9884), .Z(n9888) );
  XOR U11037 ( .A(n9887), .B(sreg[1739]), .Z(n9880) );
  XNOR U11038 ( .A(n9888), .B(n9880), .Z(c[1739]) );
  NAND U11039 ( .A(n9882), .B(n9881), .Z(n9886) );
  NANDN U11040 ( .A(n9884), .B(n9883), .Z(n9885) );
  NAND U11041 ( .A(n9886), .B(n9885), .Z(n9893) );
  ANDN U11042 ( .B(a[718]), .A(n3967), .Z(n9891) );
  AND U11043 ( .A(b[1]), .B(a[717]), .Z(n9890) );
  XOR U11044 ( .A(n9891), .B(n9890), .Z(n9892) );
  XNOR U11045 ( .A(n9893), .B(n9892), .Z(n9895) );
  XOR U11046 ( .A(sreg[1740]), .B(n9894), .Z(n9889) );
  XNOR U11047 ( .A(n9895), .B(n9889), .Z(c[1740]) );
  NAND U11048 ( .A(b[0]), .B(a[719]), .Z(n9898) );
  NAND U11049 ( .A(a[718]), .B(b[1]), .Z(n9897) );
  XNOR U11050 ( .A(n9898), .B(n9897), .Z(n9900) );
  XNOR U11051 ( .A(n9899), .B(n9900), .Z(n9904) );
  XOR U11052 ( .A(n9903), .B(sreg[1741]), .Z(n9896) );
  XNOR U11053 ( .A(n9904), .B(n9896), .Z(c[1741]) );
  NAND U11054 ( .A(n9898), .B(n9897), .Z(n9902) );
  NANDN U11055 ( .A(n9900), .B(n9899), .Z(n9901) );
  NAND U11056 ( .A(n9902), .B(n9901), .Z(n9909) );
  ANDN U11057 ( .B(a[720]), .A(n3967), .Z(n9907) );
  AND U11058 ( .A(b[1]), .B(a[719]), .Z(n9906) );
  XOR U11059 ( .A(n9907), .B(n9906), .Z(n9908) );
  XNOR U11060 ( .A(n9909), .B(n9908), .Z(n9911) );
  XOR U11061 ( .A(sreg[1742]), .B(n9910), .Z(n9905) );
  XNOR U11062 ( .A(n9911), .B(n9905), .Z(c[1742]) );
  NAND U11063 ( .A(b[0]), .B(a[721]), .Z(n9914) );
  NAND U11064 ( .A(a[720]), .B(b[1]), .Z(n9913) );
  XNOR U11065 ( .A(n9914), .B(n9913), .Z(n9916) );
  XNOR U11066 ( .A(n9915), .B(n9916), .Z(n9920) );
  XOR U11067 ( .A(n9919), .B(sreg[1743]), .Z(n9912) );
  XNOR U11068 ( .A(n9920), .B(n9912), .Z(c[1743]) );
  NAND U11069 ( .A(n9914), .B(n9913), .Z(n9918) );
  NANDN U11070 ( .A(n9916), .B(n9915), .Z(n9917) );
  NAND U11071 ( .A(n9918), .B(n9917), .Z(n9925) );
  ANDN U11072 ( .B(a[722]), .A(n3967), .Z(n9923) );
  AND U11073 ( .A(b[1]), .B(a[721]), .Z(n9922) );
  XOR U11074 ( .A(n9923), .B(n9922), .Z(n9924) );
  XNOR U11075 ( .A(n9925), .B(n9924), .Z(n9927) );
  XOR U11076 ( .A(sreg[1744]), .B(n9926), .Z(n9921) );
  XNOR U11077 ( .A(n9927), .B(n9921), .Z(c[1744]) );
  NAND U11078 ( .A(b[0]), .B(a[723]), .Z(n9930) );
  NAND U11079 ( .A(a[722]), .B(b[1]), .Z(n9929) );
  XNOR U11080 ( .A(n9930), .B(n9929), .Z(n9932) );
  XNOR U11081 ( .A(n9931), .B(n9932), .Z(n9936) );
  XOR U11082 ( .A(n9935), .B(sreg[1745]), .Z(n9928) );
  XNOR U11083 ( .A(n9936), .B(n9928), .Z(c[1745]) );
  NAND U11084 ( .A(n9930), .B(n9929), .Z(n9934) );
  NANDN U11085 ( .A(n9932), .B(n9931), .Z(n9933) );
  NAND U11086 ( .A(n9934), .B(n9933), .Z(n9941) );
  ANDN U11087 ( .B(a[724]), .A(n3967), .Z(n9939) );
  AND U11088 ( .A(b[1]), .B(a[723]), .Z(n9938) );
  XOR U11089 ( .A(n9939), .B(n9938), .Z(n9940) );
  XNOR U11090 ( .A(n9941), .B(n9940), .Z(n9943) );
  XOR U11091 ( .A(sreg[1746]), .B(n9942), .Z(n9937) );
  XNOR U11092 ( .A(n9943), .B(n9937), .Z(c[1746]) );
  NAND U11093 ( .A(b[0]), .B(a[725]), .Z(n9946) );
  NAND U11094 ( .A(a[724]), .B(b[1]), .Z(n9945) );
  XNOR U11095 ( .A(n9946), .B(n9945), .Z(n9948) );
  XNOR U11096 ( .A(n9947), .B(n9948), .Z(n9952) );
  XOR U11097 ( .A(n9951), .B(sreg[1747]), .Z(n9944) );
  XNOR U11098 ( .A(n9952), .B(n9944), .Z(c[1747]) );
  NAND U11099 ( .A(n9946), .B(n9945), .Z(n9950) );
  NANDN U11100 ( .A(n9948), .B(n9947), .Z(n9949) );
  NAND U11101 ( .A(n9950), .B(n9949), .Z(n9957) );
  ANDN U11102 ( .B(a[726]), .A(n3967), .Z(n9955) );
  AND U11103 ( .A(b[1]), .B(a[725]), .Z(n9954) );
  XOR U11104 ( .A(n9955), .B(n9954), .Z(n9956) );
  XNOR U11105 ( .A(n9957), .B(n9956), .Z(n9959) );
  XOR U11106 ( .A(sreg[1748]), .B(n9958), .Z(n9953) );
  XNOR U11107 ( .A(n9959), .B(n9953), .Z(c[1748]) );
  NAND U11108 ( .A(b[0]), .B(a[727]), .Z(n9962) );
  NAND U11109 ( .A(a[726]), .B(b[1]), .Z(n9961) );
  XNOR U11110 ( .A(n9962), .B(n9961), .Z(n9964) );
  XNOR U11111 ( .A(n9963), .B(n9964), .Z(n9968) );
  XOR U11112 ( .A(n9967), .B(sreg[1749]), .Z(n9960) );
  XNOR U11113 ( .A(n9968), .B(n9960), .Z(c[1749]) );
  NAND U11114 ( .A(n9962), .B(n9961), .Z(n9966) );
  NANDN U11115 ( .A(n9964), .B(n9963), .Z(n9965) );
  NAND U11116 ( .A(n9966), .B(n9965), .Z(n9973) );
  ANDN U11117 ( .B(a[728]), .A(n3968), .Z(n9971) );
  AND U11118 ( .A(b[1]), .B(a[727]), .Z(n9970) );
  XOR U11119 ( .A(n9971), .B(n9970), .Z(n9972) );
  XNOR U11120 ( .A(n9973), .B(n9972), .Z(n9978) );
  XOR U11121 ( .A(sreg[1750]), .B(n9977), .Z(n9969) );
  XNOR U11122 ( .A(n9978), .B(n9969), .Z(c[1750]) );
  OR U11123 ( .A(n9971), .B(n9970), .Z(n9976) );
  IV U11124 ( .A(n9972), .Z(n9974) );
  NANDN U11125 ( .A(n9974), .B(n9973), .Z(n9975) );
  NAND U11126 ( .A(n9976), .B(n9975), .Z(n9982) );
  NAND U11127 ( .A(b[0]), .B(a[729]), .Z(n9981) );
  NAND U11128 ( .A(a[728]), .B(b[1]), .Z(n9980) );
  XNOR U11129 ( .A(n9981), .B(n9980), .Z(n9983) );
  XNOR U11130 ( .A(n9982), .B(n9983), .Z(n9987) );
  XOR U11131 ( .A(n9986), .B(sreg[1751]), .Z(n9979) );
  XNOR U11132 ( .A(n9987), .B(n9979), .Z(c[1751]) );
  NAND U11133 ( .A(n9981), .B(n9980), .Z(n9985) );
  NANDN U11134 ( .A(n9983), .B(n9982), .Z(n9984) );
  NAND U11135 ( .A(n9985), .B(n9984), .Z(n9992) );
  ANDN U11136 ( .B(a[730]), .A(n3968), .Z(n9990) );
  AND U11137 ( .A(b[1]), .B(a[729]), .Z(n9989) );
  XOR U11138 ( .A(n9990), .B(n9989), .Z(n9991) );
  XNOR U11139 ( .A(n9992), .B(n9991), .Z(n9994) );
  XOR U11140 ( .A(sreg[1752]), .B(n9993), .Z(n9988) );
  XNOR U11141 ( .A(n9994), .B(n9988), .Z(c[1752]) );
  NAND U11142 ( .A(b[0]), .B(a[731]), .Z(n9997) );
  NAND U11143 ( .A(a[730]), .B(b[1]), .Z(n9996) );
  XNOR U11144 ( .A(n9997), .B(n9996), .Z(n9999) );
  XNOR U11145 ( .A(n9998), .B(n9999), .Z(n10003) );
  XOR U11146 ( .A(n10002), .B(sreg[1753]), .Z(n9995) );
  XNOR U11147 ( .A(n10003), .B(n9995), .Z(c[1753]) );
  NAND U11148 ( .A(n9997), .B(n9996), .Z(n10001) );
  NANDN U11149 ( .A(n9999), .B(n9998), .Z(n10000) );
  NAND U11150 ( .A(n10001), .B(n10000), .Z(n10008) );
  ANDN U11151 ( .B(a[732]), .A(n3968), .Z(n10006) );
  AND U11152 ( .A(b[1]), .B(a[731]), .Z(n10005) );
  XOR U11153 ( .A(n10006), .B(n10005), .Z(n10007) );
  XNOR U11154 ( .A(n10008), .B(n10007), .Z(n10010) );
  XOR U11155 ( .A(sreg[1754]), .B(n10009), .Z(n10004) );
  XNOR U11156 ( .A(n10010), .B(n10004), .Z(c[1754]) );
  NAND U11157 ( .A(b[0]), .B(a[733]), .Z(n10013) );
  NAND U11158 ( .A(a[732]), .B(b[1]), .Z(n10012) );
  XNOR U11159 ( .A(n10013), .B(n10012), .Z(n10015) );
  XNOR U11160 ( .A(n10014), .B(n10015), .Z(n10019) );
  XOR U11161 ( .A(n10018), .B(sreg[1755]), .Z(n10011) );
  XNOR U11162 ( .A(n10019), .B(n10011), .Z(c[1755]) );
  NAND U11163 ( .A(n10013), .B(n10012), .Z(n10017) );
  NANDN U11164 ( .A(n10015), .B(n10014), .Z(n10016) );
  NAND U11165 ( .A(n10017), .B(n10016), .Z(n10024) );
  ANDN U11166 ( .B(a[734]), .A(n3968), .Z(n10022) );
  AND U11167 ( .A(b[1]), .B(a[733]), .Z(n10021) );
  XOR U11168 ( .A(n10022), .B(n10021), .Z(n10023) );
  XNOR U11169 ( .A(n10024), .B(n10023), .Z(n10026) );
  XOR U11170 ( .A(sreg[1756]), .B(n10025), .Z(n10020) );
  XNOR U11171 ( .A(n10026), .B(n10020), .Z(c[1756]) );
  NAND U11172 ( .A(b[0]), .B(a[735]), .Z(n10029) );
  NAND U11173 ( .A(a[734]), .B(b[1]), .Z(n10028) );
  XNOR U11174 ( .A(n10029), .B(n10028), .Z(n10031) );
  XNOR U11175 ( .A(n10030), .B(n10031), .Z(n10035) );
  XOR U11176 ( .A(n10034), .B(sreg[1757]), .Z(n10027) );
  XNOR U11177 ( .A(n10035), .B(n10027), .Z(c[1757]) );
  NAND U11178 ( .A(n10029), .B(n10028), .Z(n10033) );
  NANDN U11179 ( .A(n10031), .B(n10030), .Z(n10032) );
  NAND U11180 ( .A(n10033), .B(n10032), .Z(n10039) );
  NAND U11181 ( .A(b[0]), .B(a[736]), .Z(n10038) );
  NAND U11182 ( .A(a[735]), .B(b[1]), .Z(n10037) );
  XNOR U11183 ( .A(n10038), .B(n10037), .Z(n10040) );
  XNOR U11184 ( .A(n10039), .B(n10040), .Z(n10044) );
  XOR U11185 ( .A(n10043), .B(sreg[1758]), .Z(n10036) );
  XNOR U11186 ( .A(n10044), .B(n10036), .Z(c[1758]) );
  NAND U11187 ( .A(n10038), .B(n10037), .Z(n10042) );
  NANDN U11188 ( .A(n10040), .B(n10039), .Z(n10041) );
  NAND U11189 ( .A(n10042), .B(n10041), .Z(n10048) );
  NAND U11190 ( .A(b[0]), .B(a[737]), .Z(n10047) );
  NAND U11191 ( .A(a[736]), .B(b[1]), .Z(n10046) );
  XNOR U11192 ( .A(n10047), .B(n10046), .Z(n10049) );
  XNOR U11193 ( .A(n10048), .B(n10049), .Z(n10053) );
  XOR U11194 ( .A(n10052), .B(sreg[1759]), .Z(n10045) );
  XNOR U11195 ( .A(n10053), .B(n10045), .Z(c[1759]) );
  NAND U11196 ( .A(n10047), .B(n10046), .Z(n10051) );
  NANDN U11197 ( .A(n10049), .B(n10048), .Z(n10050) );
  NAND U11198 ( .A(n10051), .B(n10050), .Z(n10058) );
  ANDN U11199 ( .B(a[738]), .A(n3968), .Z(n10056) );
  AND U11200 ( .A(b[1]), .B(a[737]), .Z(n10055) );
  XOR U11201 ( .A(n10056), .B(n10055), .Z(n10057) );
  XNOR U11202 ( .A(n10058), .B(n10057), .Z(n10060) );
  XOR U11203 ( .A(sreg[1760]), .B(n10059), .Z(n10054) );
  XNOR U11204 ( .A(n10060), .B(n10054), .Z(c[1760]) );
  NAND U11205 ( .A(b[0]), .B(a[739]), .Z(n10063) );
  NAND U11206 ( .A(a[738]), .B(b[1]), .Z(n10062) );
  XNOR U11207 ( .A(n10063), .B(n10062), .Z(n10065) );
  XNOR U11208 ( .A(n10064), .B(n10065), .Z(n10069) );
  XOR U11209 ( .A(n10068), .B(sreg[1761]), .Z(n10061) );
  XNOR U11210 ( .A(n10069), .B(n10061), .Z(c[1761]) );
  NAND U11211 ( .A(n10063), .B(n10062), .Z(n10067) );
  NANDN U11212 ( .A(n10065), .B(n10064), .Z(n10066) );
  NAND U11213 ( .A(n10067), .B(n10066), .Z(n10074) );
  ANDN U11214 ( .B(a[740]), .A(n3968), .Z(n10072) );
  AND U11215 ( .A(b[1]), .B(a[739]), .Z(n10071) );
  XOR U11216 ( .A(n10072), .B(n10071), .Z(n10073) );
  XNOR U11217 ( .A(n10074), .B(n10073), .Z(n10076) );
  XOR U11218 ( .A(sreg[1762]), .B(n10075), .Z(n10070) );
  XNOR U11219 ( .A(n10076), .B(n10070), .Z(c[1762]) );
  NAND U11220 ( .A(b[0]), .B(a[741]), .Z(n10079) );
  NAND U11221 ( .A(a[740]), .B(b[1]), .Z(n10078) );
  XNOR U11222 ( .A(n10079), .B(n10078), .Z(n10081) );
  XNOR U11223 ( .A(n10080), .B(n10081), .Z(n10085) );
  XOR U11224 ( .A(n10084), .B(sreg[1763]), .Z(n10077) );
  XNOR U11225 ( .A(n10085), .B(n10077), .Z(c[1763]) );
  NAND U11226 ( .A(n10079), .B(n10078), .Z(n10083) );
  NANDN U11227 ( .A(n10081), .B(n10080), .Z(n10082) );
  NAND U11228 ( .A(n10083), .B(n10082), .Z(n10090) );
  ANDN U11229 ( .B(a[742]), .A(n3968), .Z(n10088) );
  AND U11230 ( .A(b[1]), .B(a[741]), .Z(n10087) );
  XOR U11231 ( .A(n10088), .B(n10087), .Z(n10089) );
  XNOR U11232 ( .A(n10090), .B(n10089), .Z(n10092) );
  XOR U11233 ( .A(sreg[1764]), .B(n10091), .Z(n10086) );
  XNOR U11234 ( .A(n10092), .B(n10086), .Z(c[1764]) );
  ANDN U11235 ( .B(a[743]), .A(n3969), .Z(n10095) );
  AND U11236 ( .A(b[1]), .B(a[742]), .Z(n10094) );
  XOR U11237 ( .A(n10095), .B(n10094), .Z(n10096) );
  XNOR U11238 ( .A(n10097), .B(n10096), .Z(n10102) );
  XNOR U11239 ( .A(sreg[1765]), .B(n10101), .Z(n10093) );
  XNOR U11240 ( .A(n10102), .B(n10093), .Z(c[1765]) );
  OR U11241 ( .A(n10095), .B(n10094), .Z(n10100) );
  IV U11242 ( .A(n10096), .Z(n10098) );
  NANDN U11243 ( .A(n10098), .B(n10097), .Z(n10099) );
  NAND U11244 ( .A(n10100), .B(n10099), .Z(n10106) );
  NAND U11245 ( .A(b[0]), .B(a[744]), .Z(n10105) );
  NAND U11246 ( .A(a[743]), .B(b[1]), .Z(n10104) );
  XNOR U11247 ( .A(n10105), .B(n10104), .Z(n10107) );
  XNOR U11248 ( .A(n10106), .B(n10107), .Z(n10111) );
  XOR U11249 ( .A(n10110), .B(sreg[1766]), .Z(n10103) );
  XNOR U11250 ( .A(n10111), .B(n10103), .Z(c[1766]) );
  NAND U11251 ( .A(n10105), .B(n10104), .Z(n10109) );
  NANDN U11252 ( .A(n10107), .B(n10106), .Z(n10108) );
  NAND U11253 ( .A(n10109), .B(n10108), .Z(n10115) );
  NAND U11254 ( .A(b[0]), .B(a[745]), .Z(n10114) );
  NAND U11255 ( .A(a[744]), .B(b[1]), .Z(n10113) );
  XNOR U11256 ( .A(n10114), .B(n10113), .Z(n10116) );
  XNOR U11257 ( .A(n10115), .B(n10116), .Z(n10120) );
  XOR U11258 ( .A(n10119), .B(sreg[1767]), .Z(n10112) );
  XNOR U11259 ( .A(n10120), .B(n10112), .Z(c[1767]) );
  NAND U11260 ( .A(n10114), .B(n10113), .Z(n10118) );
  NANDN U11261 ( .A(n10116), .B(n10115), .Z(n10117) );
  NAND U11262 ( .A(n10118), .B(n10117), .Z(n10125) );
  ANDN U11263 ( .B(a[746]), .A(n3969), .Z(n10123) );
  AND U11264 ( .A(b[1]), .B(a[745]), .Z(n10122) );
  XOR U11265 ( .A(n10123), .B(n10122), .Z(n10124) );
  XNOR U11266 ( .A(n10125), .B(n10124), .Z(n10127) );
  XOR U11267 ( .A(sreg[1768]), .B(n10126), .Z(n10121) );
  XNOR U11268 ( .A(n10127), .B(n10121), .Z(c[1768]) );
  NAND U11269 ( .A(b[0]), .B(a[747]), .Z(n10130) );
  NAND U11270 ( .A(a[746]), .B(b[1]), .Z(n10129) );
  XNOR U11271 ( .A(n10130), .B(n10129), .Z(n10132) );
  XNOR U11272 ( .A(n10131), .B(n10132), .Z(n10136) );
  XOR U11273 ( .A(n10135), .B(sreg[1769]), .Z(n10128) );
  XNOR U11274 ( .A(n10136), .B(n10128), .Z(c[1769]) );
  NAND U11275 ( .A(n10130), .B(n10129), .Z(n10134) );
  NANDN U11276 ( .A(n10132), .B(n10131), .Z(n10133) );
  NAND U11277 ( .A(n10134), .B(n10133), .Z(n10141) );
  ANDN U11278 ( .B(a[748]), .A(n3969), .Z(n10139) );
  AND U11279 ( .A(b[1]), .B(a[747]), .Z(n10138) );
  XOR U11280 ( .A(n10139), .B(n10138), .Z(n10140) );
  XNOR U11281 ( .A(n10141), .B(n10140), .Z(n10143) );
  XOR U11282 ( .A(sreg[1770]), .B(n10142), .Z(n10137) );
  XNOR U11283 ( .A(n10143), .B(n10137), .Z(c[1770]) );
  NAND U11284 ( .A(b[0]), .B(a[749]), .Z(n10146) );
  NAND U11285 ( .A(a[748]), .B(b[1]), .Z(n10145) );
  XNOR U11286 ( .A(n10146), .B(n10145), .Z(n10148) );
  XNOR U11287 ( .A(n10147), .B(n10148), .Z(n10152) );
  XOR U11288 ( .A(n10151), .B(sreg[1771]), .Z(n10144) );
  XNOR U11289 ( .A(n10152), .B(n10144), .Z(c[1771]) );
  NAND U11290 ( .A(n10146), .B(n10145), .Z(n10150) );
  NANDN U11291 ( .A(n10148), .B(n10147), .Z(n10149) );
  NAND U11292 ( .A(n10150), .B(n10149), .Z(n10157) );
  ANDN U11293 ( .B(a[750]), .A(n3969), .Z(n10155) );
  AND U11294 ( .A(b[1]), .B(a[749]), .Z(n10154) );
  XOR U11295 ( .A(n10155), .B(n10154), .Z(n10156) );
  XNOR U11296 ( .A(n10157), .B(n10156), .Z(n10159) );
  XOR U11297 ( .A(sreg[1772]), .B(n10158), .Z(n10153) );
  XNOR U11298 ( .A(n10159), .B(n10153), .Z(c[1772]) );
  NAND U11299 ( .A(b[0]), .B(a[751]), .Z(n10162) );
  NAND U11300 ( .A(a[750]), .B(b[1]), .Z(n10161) );
  XNOR U11301 ( .A(n10162), .B(n10161), .Z(n10164) );
  XNOR U11302 ( .A(n10163), .B(n10164), .Z(n10168) );
  XOR U11303 ( .A(n10167), .B(sreg[1773]), .Z(n10160) );
  XNOR U11304 ( .A(n10168), .B(n10160), .Z(c[1773]) );
  NAND U11305 ( .A(n10162), .B(n10161), .Z(n10166) );
  NANDN U11306 ( .A(n10164), .B(n10163), .Z(n10165) );
  NAND U11307 ( .A(n10166), .B(n10165), .Z(n10173) );
  ANDN U11308 ( .B(a[752]), .A(n3969), .Z(n10171) );
  AND U11309 ( .A(b[1]), .B(a[751]), .Z(n10170) );
  XOR U11310 ( .A(n10171), .B(n10170), .Z(n10172) );
  XNOR U11311 ( .A(n10173), .B(n10172), .Z(n10175) );
  XOR U11312 ( .A(sreg[1774]), .B(n10174), .Z(n10169) );
  XNOR U11313 ( .A(n10175), .B(n10169), .Z(c[1774]) );
  NAND U11314 ( .A(b[0]), .B(a[753]), .Z(n10178) );
  NAND U11315 ( .A(a[752]), .B(b[1]), .Z(n10177) );
  XNOR U11316 ( .A(n10178), .B(n10177), .Z(n10180) );
  XNOR U11317 ( .A(n10179), .B(n10180), .Z(n10184) );
  XOR U11318 ( .A(n10183), .B(sreg[1775]), .Z(n10176) );
  XNOR U11319 ( .A(n10184), .B(n10176), .Z(c[1775]) );
  NAND U11320 ( .A(n10178), .B(n10177), .Z(n10182) );
  NANDN U11321 ( .A(n10180), .B(n10179), .Z(n10181) );
  NAND U11322 ( .A(n10182), .B(n10181), .Z(n10189) );
  ANDN U11323 ( .B(a[754]), .A(n3969), .Z(n10187) );
  AND U11324 ( .A(b[1]), .B(a[753]), .Z(n10186) );
  XOR U11325 ( .A(n10187), .B(n10186), .Z(n10188) );
  XNOR U11326 ( .A(n10189), .B(n10188), .Z(n10191) );
  XOR U11327 ( .A(sreg[1776]), .B(n10190), .Z(n10185) );
  XNOR U11328 ( .A(n10191), .B(n10185), .Z(c[1776]) );
  ANDN U11329 ( .B(a[755]), .A(n3969), .Z(n10194) );
  AND U11330 ( .A(b[1]), .B(a[754]), .Z(n10193) );
  XOR U11331 ( .A(n10194), .B(n10193), .Z(n10195) );
  XNOR U11332 ( .A(n10196), .B(n10195), .Z(n10198) );
  XNOR U11333 ( .A(sreg[1777]), .B(n10197), .Z(n10192) );
  XNOR U11334 ( .A(n10198), .B(n10192), .Z(c[1777]) );
  ANDN U11335 ( .B(a[756]), .A(n3970), .Z(n10201) );
  AND U11336 ( .A(b[1]), .B(a[755]), .Z(n10200) );
  XOR U11337 ( .A(n10201), .B(n10200), .Z(n10202) );
  XNOR U11338 ( .A(n10203), .B(n10202), .Z(n10208) );
  XNOR U11339 ( .A(sreg[1778]), .B(n10207), .Z(n10199) );
  XNOR U11340 ( .A(n10208), .B(n10199), .Z(c[1778]) );
  OR U11341 ( .A(n10201), .B(n10200), .Z(n10206) );
  IV U11342 ( .A(n10202), .Z(n10204) );
  NANDN U11343 ( .A(n10204), .B(n10203), .Z(n10205) );
  NAND U11344 ( .A(n10206), .B(n10205), .Z(n10212) );
  NAND U11345 ( .A(b[0]), .B(a[757]), .Z(n10211) );
  NAND U11346 ( .A(a[756]), .B(b[1]), .Z(n10210) );
  XNOR U11347 ( .A(n10211), .B(n10210), .Z(n10213) );
  XNOR U11348 ( .A(n10212), .B(n10213), .Z(n10217) );
  XOR U11349 ( .A(n10216), .B(sreg[1779]), .Z(n10209) );
  XNOR U11350 ( .A(n10217), .B(n10209), .Z(c[1779]) );
  NAND U11351 ( .A(n10211), .B(n10210), .Z(n10215) );
  NANDN U11352 ( .A(n10213), .B(n10212), .Z(n10214) );
  NAND U11353 ( .A(n10215), .B(n10214), .Z(n10222) );
  ANDN U11354 ( .B(a[758]), .A(n3970), .Z(n10220) );
  AND U11355 ( .A(b[1]), .B(a[757]), .Z(n10219) );
  XOR U11356 ( .A(n10220), .B(n10219), .Z(n10221) );
  XNOR U11357 ( .A(n10222), .B(n10221), .Z(n10224) );
  XOR U11358 ( .A(sreg[1780]), .B(n10223), .Z(n10218) );
  XNOR U11359 ( .A(n10224), .B(n10218), .Z(c[1780]) );
  NAND U11360 ( .A(b[0]), .B(a[759]), .Z(n10227) );
  NAND U11361 ( .A(a[758]), .B(b[1]), .Z(n10226) );
  XNOR U11362 ( .A(n10227), .B(n10226), .Z(n10229) );
  XNOR U11363 ( .A(n10228), .B(n10229), .Z(n10233) );
  XOR U11364 ( .A(n10232), .B(sreg[1781]), .Z(n10225) );
  XNOR U11365 ( .A(n10233), .B(n10225), .Z(c[1781]) );
  NAND U11366 ( .A(n10227), .B(n10226), .Z(n10231) );
  NANDN U11367 ( .A(n10229), .B(n10228), .Z(n10230) );
  NAND U11368 ( .A(n10231), .B(n10230), .Z(n10238) );
  ANDN U11369 ( .B(a[760]), .A(n3970), .Z(n10236) );
  AND U11370 ( .A(b[1]), .B(a[759]), .Z(n10235) );
  XOR U11371 ( .A(n10236), .B(n10235), .Z(n10237) );
  XNOR U11372 ( .A(n10238), .B(n10237), .Z(n10240) );
  XOR U11373 ( .A(sreg[1782]), .B(n10239), .Z(n10234) );
  XNOR U11374 ( .A(n10240), .B(n10234), .Z(c[1782]) );
  NAND U11375 ( .A(b[0]), .B(a[761]), .Z(n10243) );
  NAND U11376 ( .A(a[760]), .B(b[1]), .Z(n10242) );
  XNOR U11377 ( .A(n10243), .B(n10242), .Z(n10245) );
  XNOR U11378 ( .A(n10244), .B(n10245), .Z(n10249) );
  XOR U11379 ( .A(n10248), .B(sreg[1783]), .Z(n10241) );
  XNOR U11380 ( .A(n10249), .B(n10241), .Z(c[1783]) );
  NAND U11381 ( .A(n10243), .B(n10242), .Z(n10247) );
  NANDN U11382 ( .A(n10245), .B(n10244), .Z(n10246) );
  NAND U11383 ( .A(n10247), .B(n10246), .Z(n10254) );
  ANDN U11384 ( .B(a[762]), .A(n3970), .Z(n10252) );
  AND U11385 ( .A(b[1]), .B(a[761]), .Z(n10251) );
  XOR U11386 ( .A(n10252), .B(n10251), .Z(n10253) );
  XNOR U11387 ( .A(n10254), .B(n10253), .Z(n10256) );
  XOR U11388 ( .A(sreg[1784]), .B(n10255), .Z(n10250) );
  XNOR U11389 ( .A(n10256), .B(n10250), .Z(c[1784]) );
  NAND U11390 ( .A(b[0]), .B(a[763]), .Z(n10259) );
  NAND U11391 ( .A(a[762]), .B(b[1]), .Z(n10258) );
  XNOR U11392 ( .A(n10259), .B(n10258), .Z(n10261) );
  XNOR U11393 ( .A(n10260), .B(n10261), .Z(n10265) );
  XOR U11394 ( .A(n10264), .B(sreg[1785]), .Z(n10257) );
  XNOR U11395 ( .A(n10265), .B(n10257), .Z(c[1785]) );
  NAND U11396 ( .A(n10259), .B(n10258), .Z(n10263) );
  NANDN U11397 ( .A(n10261), .B(n10260), .Z(n10262) );
  NAND U11398 ( .A(n10263), .B(n10262), .Z(n10270) );
  ANDN U11399 ( .B(a[764]), .A(n3970), .Z(n10268) );
  AND U11400 ( .A(b[1]), .B(a[763]), .Z(n10267) );
  XOR U11401 ( .A(n10268), .B(n10267), .Z(n10269) );
  XNOR U11402 ( .A(n10270), .B(n10269), .Z(n10272) );
  XOR U11403 ( .A(sreg[1786]), .B(n10271), .Z(n10266) );
  XNOR U11404 ( .A(n10272), .B(n10266), .Z(c[1786]) );
  NAND U11405 ( .A(b[0]), .B(a[765]), .Z(n10275) );
  NAND U11406 ( .A(a[764]), .B(b[1]), .Z(n10274) );
  XNOR U11407 ( .A(n10275), .B(n10274), .Z(n10277) );
  XNOR U11408 ( .A(n10276), .B(n10277), .Z(n10281) );
  XOR U11409 ( .A(n10280), .B(sreg[1787]), .Z(n10273) );
  XNOR U11410 ( .A(n10281), .B(n10273), .Z(c[1787]) );
  NAND U11411 ( .A(n10275), .B(n10274), .Z(n10279) );
  NANDN U11412 ( .A(n10277), .B(n10276), .Z(n10278) );
  NAND U11413 ( .A(n10279), .B(n10278), .Z(n10286) );
  ANDN U11414 ( .B(a[766]), .A(n3970), .Z(n10284) );
  AND U11415 ( .A(b[1]), .B(a[765]), .Z(n10283) );
  XOR U11416 ( .A(n10284), .B(n10283), .Z(n10285) );
  XNOR U11417 ( .A(n10286), .B(n10285), .Z(n10288) );
  XOR U11418 ( .A(sreg[1788]), .B(n10287), .Z(n10282) );
  XNOR U11419 ( .A(n10288), .B(n10282), .Z(c[1788]) );
  NAND U11420 ( .A(b[0]), .B(a[767]), .Z(n10291) );
  NAND U11421 ( .A(a[766]), .B(b[1]), .Z(n10290) );
  XNOR U11422 ( .A(n10291), .B(n10290), .Z(n10293) );
  XNOR U11423 ( .A(n10292), .B(n10293), .Z(n10297) );
  XOR U11424 ( .A(n10296), .B(sreg[1789]), .Z(n10289) );
  XNOR U11425 ( .A(n10297), .B(n10289), .Z(c[1789]) );
  NAND U11426 ( .A(n10291), .B(n10290), .Z(n10295) );
  NANDN U11427 ( .A(n10293), .B(n10292), .Z(n10294) );
  NAND U11428 ( .A(n10295), .B(n10294), .Z(n10302) );
  ANDN U11429 ( .B(a[768]), .A(n3970), .Z(n10300) );
  AND U11430 ( .A(b[1]), .B(a[767]), .Z(n10299) );
  XOR U11431 ( .A(n10300), .B(n10299), .Z(n10301) );
  XNOR U11432 ( .A(n10302), .B(n10301), .Z(n10304) );
  XOR U11433 ( .A(sreg[1790]), .B(n10303), .Z(n10298) );
  XNOR U11434 ( .A(n10304), .B(n10298), .Z(c[1790]) );
  NAND U11435 ( .A(b[0]), .B(a[769]), .Z(n10307) );
  NAND U11436 ( .A(a[768]), .B(b[1]), .Z(n10306) );
  XNOR U11437 ( .A(n10307), .B(n10306), .Z(n10309) );
  XNOR U11438 ( .A(n10308), .B(n10309), .Z(n10313) );
  XOR U11439 ( .A(n10312), .B(sreg[1791]), .Z(n10305) );
  XNOR U11440 ( .A(n10313), .B(n10305), .Z(c[1791]) );
  NAND U11441 ( .A(n10307), .B(n10306), .Z(n10311) );
  NANDN U11442 ( .A(n10309), .B(n10308), .Z(n10310) );
  NAND U11443 ( .A(n10311), .B(n10310), .Z(n10318) );
  ANDN U11444 ( .B(a[770]), .A(n3971), .Z(n10316) );
  AND U11445 ( .A(b[1]), .B(a[769]), .Z(n10315) );
  XOR U11446 ( .A(n10316), .B(n10315), .Z(n10317) );
  XNOR U11447 ( .A(n10318), .B(n10317), .Z(n10323) );
  XOR U11448 ( .A(sreg[1792]), .B(n10322), .Z(n10314) );
  XNOR U11449 ( .A(n10323), .B(n10314), .Z(c[1792]) );
  OR U11450 ( .A(n10316), .B(n10315), .Z(n10321) );
  IV U11451 ( .A(n10317), .Z(n10319) );
  NANDN U11452 ( .A(n10319), .B(n10318), .Z(n10320) );
  NAND U11453 ( .A(n10321), .B(n10320), .Z(n10327) );
  NAND U11454 ( .A(b[0]), .B(a[771]), .Z(n10326) );
  NAND U11455 ( .A(a[770]), .B(b[1]), .Z(n10325) );
  XNOR U11456 ( .A(n10326), .B(n10325), .Z(n10328) );
  XNOR U11457 ( .A(n10327), .B(n10328), .Z(n10332) );
  XOR U11458 ( .A(n10331), .B(sreg[1793]), .Z(n10324) );
  XNOR U11459 ( .A(n10332), .B(n10324), .Z(c[1793]) );
  NAND U11460 ( .A(n10326), .B(n10325), .Z(n10330) );
  NANDN U11461 ( .A(n10328), .B(n10327), .Z(n10329) );
  NAND U11462 ( .A(n10330), .B(n10329), .Z(n10336) );
  NAND U11463 ( .A(b[0]), .B(a[772]), .Z(n10335) );
  NAND U11464 ( .A(a[771]), .B(b[1]), .Z(n10334) );
  XNOR U11465 ( .A(n10335), .B(n10334), .Z(n10337) );
  XNOR U11466 ( .A(n10336), .B(n10337), .Z(n10341) );
  XOR U11467 ( .A(n10340), .B(sreg[1794]), .Z(n10333) );
  XNOR U11468 ( .A(n10341), .B(n10333), .Z(c[1794]) );
  NAND U11469 ( .A(n10335), .B(n10334), .Z(n10339) );
  NANDN U11470 ( .A(n10337), .B(n10336), .Z(n10338) );
  NAND U11471 ( .A(n10339), .B(n10338), .Z(n10345) );
  NAND U11472 ( .A(b[0]), .B(a[773]), .Z(n10344) );
  NAND U11473 ( .A(a[772]), .B(b[1]), .Z(n10343) );
  XNOR U11474 ( .A(n10344), .B(n10343), .Z(n10346) );
  XNOR U11475 ( .A(n10345), .B(n10346), .Z(n10350) );
  XOR U11476 ( .A(n10349), .B(sreg[1795]), .Z(n10342) );
  XNOR U11477 ( .A(n10350), .B(n10342), .Z(c[1795]) );
  NAND U11478 ( .A(n10344), .B(n10343), .Z(n10348) );
  NANDN U11479 ( .A(n10346), .B(n10345), .Z(n10347) );
  NAND U11480 ( .A(n10348), .B(n10347), .Z(n10355) );
  ANDN U11481 ( .B(a[774]), .A(n3971), .Z(n10353) );
  AND U11482 ( .A(b[1]), .B(a[773]), .Z(n10352) );
  XOR U11483 ( .A(n10353), .B(n10352), .Z(n10354) );
  XNOR U11484 ( .A(n10355), .B(n10354), .Z(n10357) );
  XOR U11485 ( .A(sreg[1796]), .B(n10356), .Z(n10351) );
  XNOR U11486 ( .A(n10357), .B(n10351), .Z(c[1796]) );
  NAND U11487 ( .A(b[0]), .B(a[775]), .Z(n10360) );
  NAND U11488 ( .A(a[774]), .B(b[1]), .Z(n10359) );
  XNOR U11489 ( .A(n10360), .B(n10359), .Z(n10362) );
  XNOR U11490 ( .A(n10361), .B(n10362), .Z(n10366) );
  XOR U11491 ( .A(n10365), .B(sreg[1797]), .Z(n10358) );
  XNOR U11492 ( .A(n10366), .B(n10358), .Z(c[1797]) );
  NAND U11493 ( .A(n10360), .B(n10359), .Z(n10364) );
  NANDN U11494 ( .A(n10362), .B(n10361), .Z(n10363) );
  NAND U11495 ( .A(n10364), .B(n10363), .Z(n10371) );
  ANDN U11496 ( .B(a[776]), .A(n3971), .Z(n10369) );
  AND U11497 ( .A(b[1]), .B(a[775]), .Z(n10368) );
  XOR U11498 ( .A(n10369), .B(n10368), .Z(n10370) );
  XNOR U11499 ( .A(n10371), .B(n10370), .Z(n10373) );
  XOR U11500 ( .A(sreg[1798]), .B(n10372), .Z(n10367) );
  XNOR U11501 ( .A(n10373), .B(n10367), .Z(c[1798]) );
  NAND U11502 ( .A(b[0]), .B(a[777]), .Z(n10376) );
  NAND U11503 ( .A(a[776]), .B(b[1]), .Z(n10375) );
  XNOR U11504 ( .A(n10376), .B(n10375), .Z(n10378) );
  XNOR U11505 ( .A(n10377), .B(n10378), .Z(n10382) );
  XOR U11506 ( .A(n10381), .B(sreg[1799]), .Z(n10374) );
  XNOR U11507 ( .A(n10382), .B(n10374), .Z(c[1799]) );
  NAND U11508 ( .A(n10376), .B(n10375), .Z(n10380) );
  NANDN U11509 ( .A(n10378), .B(n10377), .Z(n10379) );
  NAND U11510 ( .A(n10380), .B(n10379), .Z(n10387) );
  ANDN U11511 ( .B(a[778]), .A(n3971), .Z(n10385) );
  AND U11512 ( .A(b[1]), .B(a[777]), .Z(n10384) );
  XOR U11513 ( .A(n10385), .B(n10384), .Z(n10386) );
  XNOR U11514 ( .A(n10387), .B(n10386), .Z(n10389) );
  XOR U11515 ( .A(sreg[1800]), .B(n10388), .Z(n10383) );
  XNOR U11516 ( .A(n10389), .B(n10383), .Z(c[1800]) );
  NAND U11517 ( .A(b[0]), .B(a[779]), .Z(n10392) );
  NAND U11518 ( .A(a[778]), .B(b[1]), .Z(n10391) );
  XNOR U11519 ( .A(n10392), .B(n10391), .Z(n10394) );
  XNOR U11520 ( .A(n10393), .B(n10394), .Z(n10398) );
  XOR U11521 ( .A(n10397), .B(sreg[1801]), .Z(n10390) );
  XNOR U11522 ( .A(n10398), .B(n10390), .Z(c[1801]) );
  NAND U11523 ( .A(n10392), .B(n10391), .Z(n10396) );
  NANDN U11524 ( .A(n10394), .B(n10393), .Z(n10395) );
  NAND U11525 ( .A(n10396), .B(n10395), .Z(n10403) );
  ANDN U11526 ( .B(a[780]), .A(n3971), .Z(n10401) );
  AND U11527 ( .A(b[1]), .B(a[779]), .Z(n10400) );
  XOR U11528 ( .A(n10401), .B(n10400), .Z(n10402) );
  XNOR U11529 ( .A(n10403), .B(n10402), .Z(n10405) );
  XOR U11530 ( .A(sreg[1802]), .B(n10404), .Z(n10399) );
  XNOR U11531 ( .A(n10405), .B(n10399), .Z(c[1802]) );
  NAND U11532 ( .A(b[0]), .B(a[781]), .Z(n10408) );
  NAND U11533 ( .A(a[780]), .B(b[1]), .Z(n10407) );
  XNOR U11534 ( .A(n10408), .B(n10407), .Z(n10410) );
  XNOR U11535 ( .A(n10409), .B(n10410), .Z(n10414) );
  XOR U11536 ( .A(n10413), .B(sreg[1803]), .Z(n10406) );
  XNOR U11537 ( .A(n10414), .B(n10406), .Z(c[1803]) );
  NAND U11538 ( .A(n10408), .B(n10407), .Z(n10412) );
  NANDN U11539 ( .A(n10410), .B(n10409), .Z(n10411) );
  NAND U11540 ( .A(n10412), .B(n10411), .Z(n10419) );
  ANDN U11541 ( .B(a[782]), .A(n3971), .Z(n10417) );
  AND U11542 ( .A(b[1]), .B(a[781]), .Z(n10416) );
  XOR U11543 ( .A(n10417), .B(n10416), .Z(n10418) );
  XNOR U11544 ( .A(n10419), .B(n10418), .Z(n10421) );
  XOR U11545 ( .A(sreg[1804]), .B(n10420), .Z(n10415) );
  XNOR U11546 ( .A(n10421), .B(n10415), .Z(c[1804]) );
  NAND U11547 ( .A(b[0]), .B(a[783]), .Z(n10424) );
  NAND U11548 ( .A(a[782]), .B(b[1]), .Z(n10423) );
  XNOR U11549 ( .A(n10424), .B(n10423), .Z(n10426) );
  XNOR U11550 ( .A(n10425), .B(n10426), .Z(n10430) );
  XOR U11551 ( .A(n10429), .B(sreg[1805]), .Z(n10422) );
  XNOR U11552 ( .A(n10430), .B(n10422), .Z(c[1805]) );
  NAND U11553 ( .A(n10424), .B(n10423), .Z(n10428) );
  NANDN U11554 ( .A(n10426), .B(n10425), .Z(n10427) );
  NAND U11555 ( .A(n10428), .B(n10427), .Z(n10435) );
  ANDN U11556 ( .B(a[784]), .A(n3971), .Z(n10433) );
  AND U11557 ( .A(b[1]), .B(a[783]), .Z(n10432) );
  XOR U11558 ( .A(n10433), .B(n10432), .Z(n10434) );
  XNOR U11559 ( .A(n10435), .B(n10434), .Z(n10437) );
  XOR U11560 ( .A(sreg[1806]), .B(n10436), .Z(n10431) );
  XNOR U11561 ( .A(n10437), .B(n10431), .Z(c[1806]) );
  NAND U11562 ( .A(b[0]), .B(a[785]), .Z(n10440) );
  NAND U11563 ( .A(a[784]), .B(b[1]), .Z(n10439) );
  XNOR U11564 ( .A(n10440), .B(n10439), .Z(n10442) );
  XNOR U11565 ( .A(n10441), .B(n10442), .Z(n10446) );
  XOR U11566 ( .A(n10445), .B(sreg[1807]), .Z(n10438) );
  XNOR U11567 ( .A(n10446), .B(n10438), .Z(c[1807]) );
  NAND U11568 ( .A(n10440), .B(n10439), .Z(n10444) );
  NANDN U11569 ( .A(n10442), .B(n10441), .Z(n10443) );
  NAND U11570 ( .A(n10444), .B(n10443), .Z(n10451) );
  ANDN U11571 ( .B(a[786]), .A(n3972), .Z(n10449) );
  AND U11572 ( .A(b[1]), .B(a[785]), .Z(n10448) );
  XOR U11573 ( .A(n10449), .B(n10448), .Z(n10450) );
  XNOR U11574 ( .A(n10451), .B(n10450), .Z(n10456) );
  XOR U11575 ( .A(sreg[1808]), .B(n10455), .Z(n10447) );
  XNOR U11576 ( .A(n10456), .B(n10447), .Z(c[1808]) );
  OR U11577 ( .A(n10449), .B(n10448), .Z(n10454) );
  IV U11578 ( .A(n10450), .Z(n10452) );
  NANDN U11579 ( .A(n10452), .B(n10451), .Z(n10453) );
  NAND U11580 ( .A(n10454), .B(n10453), .Z(n10460) );
  NAND U11581 ( .A(b[0]), .B(a[787]), .Z(n10459) );
  NAND U11582 ( .A(a[786]), .B(b[1]), .Z(n10458) );
  XNOR U11583 ( .A(n10459), .B(n10458), .Z(n10461) );
  XNOR U11584 ( .A(n10460), .B(n10461), .Z(n10465) );
  XOR U11585 ( .A(n10464), .B(sreg[1809]), .Z(n10457) );
  XNOR U11586 ( .A(n10465), .B(n10457), .Z(c[1809]) );
  NAND U11587 ( .A(n10459), .B(n10458), .Z(n10463) );
  NANDN U11588 ( .A(n10461), .B(n10460), .Z(n10462) );
  NAND U11589 ( .A(n10463), .B(n10462), .Z(n10470) );
  ANDN U11590 ( .B(a[788]), .A(n3972), .Z(n10468) );
  AND U11591 ( .A(b[1]), .B(a[787]), .Z(n10467) );
  XOR U11592 ( .A(n10468), .B(n10467), .Z(n10469) );
  XNOR U11593 ( .A(n10470), .B(n10469), .Z(n10472) );
  XOR U11594 ( .A(sreg[1810]), .B(n10471), .Z(n10466) );
  XNOR U11595 ( .A(n10472), .B(n10466), .Z(c[1810]) );
  ANDN U11596 ( .B(a[789]), .A(n3972), .Z(n10475) );
  AND U11597 ( .A(b[1]), .B(a[788]), .Z(n10474) );
  XOR U11598 ( .A(n10475), .B(n10474), .Z(n10476) );
  XNOR U11599 ( .A(n10477), .B(n10476), .Z(n10479) );
  XNOR U11600 ( .A(sreg[1811]), .B(n10478), .Z(n10473) );
  XNOR U11601 ( .A(n10479), .B(n10473), .Z(c[1811]) );
  ANDN U11602 ( .B(a[790]), .A(n3972), .Z(n10482) );
  AND U11603 ( .A(b[1]), .B(a[789]), .Z(n10481) );
  XOR U11604 ( .A(n10482), .B(n10481), .Z(n10483) );
  XNOR U11605 ( .A(n10484), .B(n10483), .Z(n10486) );
  XNOR U11606 ( .A(sreg[1812]), .B(n10485), .Z(n10480) );
  XNOR U11607 ( .A(n10486), .B(n10480), .Z(c[1812]) );
  NAND U11608 ( .A(b[0]), .B(a[791]), .Z(n10489) );
  NAND U11609 ( .A(a[790]), .B(b[1]), .Z(n10488) );
  XNOR U11610 ( .A(n10489), .B(n10488), .Z(n10491) );
  XNOR U11611 ( .A(n10490), .B(n10491), .Z(n10495) );
  XOR U11612 ( .A(n10494), .B(sreg[1813]), .Z(n10487) );
  XNOR U11613 ( .A(n10495), .B(n10487), .Z(c[1813]) );
  NAND U11614 ( .A(n10489), .B(n10488), .Z(n10493) );
  NANDN U11615 ( .A(n10491), .B(n10490), .Z(n10492) );
  NAND U11616 ( .A(n10493), .B(n10492), .Z(n10500) );
  ANDN U11617 ( .B(a[792]), .A(n3972), .Z(n10498) );
  AND U11618 ( .A(b[1]), .B(a[791]), .Z(n10497) );
  XOR U11619 ( .A(n10498), .B(n10497), .Z(n10499) );
  XNOR U11620 ( .A(n10500), .B(n10499), .Z(n10502) );
  XOR U11621 ( .A(sreg[1814]), .B(n10501), .Z(n10496) );
  XNOR U11622 ( .A(n10502), .B(n10496), .Z(c[1814]) );
  NAND U11623 ( .A(b[0]), .B(a[793]), .Z(n10505) );
  NAND U11624 ( .A(a[792]), .B(b[1]), .Z(n10504) );
  XNOR U11625 ( .A(n10505), .B(n10504), .Z(n10507) );
  XNOR U11626 ( .A(n10506), .B(n10507), .Z(n10511) );
  XOR U11627 ( .A(n10510), .B(sreg[1815]), .Z(n10503) );
  XNOR U11628 ( .A(n10511), .B(n10503), .Z(c[1815]) );
  NAND U11629 ( .A(n10505), .B(n10504), .Z(n10509) );
  NANDN U11630 ( .A(n10507), .B(n10506), .Z(n10508) );
  NAND U11631 ( .A(n10509), .B(n10508), .Z(n10516) );
  ANDN U11632 ( .B(a[794]), .A(n3972), .Z(n10514) );
  AND U11633 ( .A(b[1]), .B(a[793]), .Z(n10513) );
  XOR U11634 ( .A(n10514), .B(n10513), .Z(n10515) );
  XNOR U11635 ( .A(n10516), .B(n10515), .Z(n10518) );
  XOR U11636 ( .A(sreg[1816]), .B(n10517), .Z(n10512) );
  XNOR U11637 ( .A(n10518), .B(n10512), .Z(c[1816]) );
  NAND U11638 ( .A(b[0]), .B(a[795]), .Z(n10521) );
  NAND U11639 ( .A(a[794]), .B(b[1]), .Z(n10520) );
  XNOR U11640 ( .A(n10521), .B(n10520), .Z(n10523) );
  XNOR U11641 ( .A(n10522), .B(n10523), .Z(n10527) );
  XOR U11642 ( .A(n10526), .B(sreg[1817]), .Z(n10519) );
  XNOR U11643 ( .A(n10527), .B(n10519), .Z(c[1817]) );
  NAND U11644 ( .A(n10521), .B(n10520), .Z(n10525) );
  NANDN U11645 ( .A(n10523), .B(n10522), .Z(n10524) );
  NAND U11646 ( .A(n10525), .B(n10524), .Z(n10532) );
  ANDN U11647 ( .B(a[796]), .A(n3972), .Z(n10530) );
  AND U11648 ( .A(b[1]), .B(a[795]), .Z(n10529) );
  XOR U11649 ( .A(n10530), .B(n10529), .Z(n10531) );
  XNOR U11650 ( .A(n10532), .B(n10531), .Z(n10534) );
  XOR U11651 ( .A(sreg[1818]), .B(n10533), .Z(n10528) );
  XNOR U11652 ( .A(n10534), .B(n10528), .Z(c[1818]) );
  NAND U11653 ( .A(b[0]), .B(a[797]), .Z(n10537) );
  NAND U11654 ( .A(a[796]), .B(b[1]), .Z(n10536) );
  XNOR U11655 ( .A(n10537), .B(n10536), .Z(n10539) );
  XNOR U11656 ( .A(n10538), .B(n10539), .Z(n10543) );
  XOR U11657 ( .A(n10542), .B(sreg[1819]), .Z(n10535) );
  XNOR U11658 ( .A(n10543), .B(n10535), .Z(c[1819]) );
  NAND U11659 ( .A(n10537), .B(n10536), .Z(n10541) );
  NANDN U11660 ( .A(n10539), .B(n10538), .Z(n10540) );
  NAND U11661 ( .A(n10541), .B(n10540), .Z(n10548) );
  ANDN U11662 ( .B(a[798]), .A(n3973), .Z(n10546) );
  AND U11663 ( .A(b[1]), .B(a[797]), .Z(n10545) );
  XOR U11664 ( .A(n10546), .B(n10545), .Z(n10547) );
  XNOR U11665 ( .A(n10548), .B(n10547), .Z(n10553) );
  XOR U11666 ( .A(sreg[1820]), .B(n10552), .Z(n10544) );
  XNOR U11667 ( .A(n10553), .B(n10544), .Z(c[1820]) );
  OR U11668 ( .A(n10546), .B(n10545), .Z(n10551) );
  IV U11669 ( .A(n10547), .Z(n10549) );
  NANDN U11670 ( .A(n10549), .B(n10548), .Z(n10550) );
  NAND U11671 ( .A(n10551), .B(n10550), .Z(n10557) );
  NAND U11672 ( .A(b[0]), .B(a[799]), .Z(n10556) );
  NAND U11673 ( .A(a[798]), .B(b[1]), .Z(n10555) );
  XNOR U11674 ( .A(n10556), .B(n10555), .Z(n10558) );
  XNOR U11675 ( .A(n10557), .B(n10558), .Z(n10562) );
  XOR U11676 ( .A(n10561), .B(sreg[1821]), .Z(n10554) );
  XNOR U11677 ( .A(n10562), .B(n10554), .Z(c[1821]) );
  NAND U11678 ( .A(n10556), .B(n10555), .Z(n10560) );
  NANDN U11679 ( .A(n10558), .B(n10557), .Z(n10559) );
  NAND U11680 ( .A(n10560), .B(n10559), .Z(n10567) );
  ANDN U11681 ( .B(a[800]), .A(n3973), .Z(n10565) );
  AND U11682 ( .A(b[1]), .B(a[799]), .Z(n10564) );
  XOR U11683 ( .A(n10565), .B(n10564), .Z(n10566) );
  XNOR U11684 ( .A(n10567), .B(n10566), .Z(n10569) );
  XOR U11685 ( .A(sreg[1822]), .B(n10568), .Z(n10563) );
  XNOR U11686 ( .A(n10569), .B(n10563), .Z(c[1822]) );
  NAND U11687 ( .A(b[0]), .B(a[801]), .Z(n10572) );
  NAND U11688 ( .A(a[800]), .B(b[1]), .Z(n10571) );
  XNOR U11689 ( .A(n10572), .B(n10571), .Z(n10574) );
  XNOR U11690 ( .A(n10573), .B(n10574), .Z(n10578) );
  XOR U11691 ( .A(n10577), .B(sreg[1823]), .Z(n10570) );
  XNOR U11692 ( .A(n10578), .B(n10570), .Z(c[1823]) );
  NAND U11693 ( .A(n10572), .B(n10571), .Z(n10576) );
  NANDN U11694 ( .A(n10574), .B(n10573), .Z(n10575) );
  NAND U11695 ( .A(n10576), .B(n10575), .Z(n10583) );
  ANDN U11696 ( .B(a[802]), .A(n3973), .Z(n10581) );
  AND U11697 ( .A(b[1]), .B(a[801]), .Z(n10580) );
  XOR U11698 ( .A(n10581), .B(n10580), .Z(n10582) );
  XNOR U11699 ( .A(n10583), .B(n10582), .Z(n10585) );
  XOR U11700 ( .A(sreg[1824]), .B(n10584), .Z(n10579) );
  XNOR U11701 ( .A(n10585), .B(n10579), .Z(c[1824]) );
  NAND U11702 ( .A(b[0]), .B(a[803]), .Z(n10588) );
  NAND U11703 ( .A(a[802]), .B(b[1]), .Z(n10587) );
  XNOR U11704 ( .A(n10588), .B(n10587), .Z(n10590) );
  XNOR U11705 ( .A(n10589), .B(n10590), .Z(n10594) );
  XOR U11706 ( .A(n10593), .B(sreg[1825]), .Z(n10586) );
  XNOR U11707 ( .A(n10594), .B(n10586), .Z(c[1825]) );
  NAND U11708 ( .A(n10588), .B(n10587), .Z(n10592) );
  NANDN U11709 ( .A(n10590), .B(n10589), .Z(n10591) );
  NAND U11710 ( .A(n10592), .B(n10591), .Z(n10599) );
  ANDN U11711 ( .B(a[804]), .A(n3973), .Z(n10597) );
  AND U11712 ( .A(b[1]), .B(a[803]), .Z(n10596) );
  XOR U11713 ( .A(n10597), .B(n10596), .Z(n10598) );
  XNOR U11714 ( .A(n10599), .B(n10598), .Z(n10601) );
  XOR U11715 ( .A(sreg[1826]), .B(n10600), .Z(n10595) );
  XNOR U11716 ( .A(n10601), .B(n10595), .Z(c[1826]) );
  NAND U11717 ( .A(b[0]), .B(a[805]), .Z(n10604) );
  NAND U11718 ( .A(a[804]), .B(b[1]), .Z(n10603) );
  XNOR U11719 ( .A(n10604), .B(n10603), .Z(n10606) );
  XNOR U11720 ( .A(n10605), .B(n10606), .Z(n10610) );
  XOR U11721 ( .A(n10609), .B(sreg[1827]), .Z(n10602) );
  XNOR U11722 ( .A(n10610), .B(n10602), .Z(c[1827]) );
  NAND U11723 ( .A(n10604), .B(n10603), .Z(n10608) );
  NANDN U11724 ( .A(n10606), .B(n10605), .Z(n10607) );
  NAND U11725 ( .A(n10608), .B(n10607), .Z(n10615) );
  ANDN U11726 ( .B(a[806]), .A(n3973), .Z(n10613) );
  AND U11727 ( .A(b[1]), .B(a[805]), .Z(n10612) );
  XOR U11728 ( .A(n10613), .B(n10612), .Z(n10614) );
  XNOR U11729 ( .A(n10615), .B(n10614), .Z(n10617) );
  XOR U11730 ( .A(sreg[1828]), .B(n10616), .Z(n10611) );
  XNOR U11731 ( .A(n10617), .B(n10611), .Z(c[1828]) );
  ANDN U11732 ( .B(a[807]), .A(n3973), .Z(n10620) );
  AND U11733 ( .A(b[1]), .B(a[806]), .Z(n10619) );
  XOR U11734 ( .A(n10620), .B(n10619), .Z(n10621) );
  XNOR U11735 ( .A(n10622), .B(n10621), .Z(n10624) );
  XNOR U11736 ( .A(sreg[1829]), .B(n10623), .Z(n10618) );
  XNOR U11737 ( .A(n10624), .B(n10618), .Z(c[1829]) );
  ANDN U11738 ( .B(a[808]), .A(n3973), .Z(n10627) );
  AND U11739 ( .A(b[1]), .B(a[807]), .Z(n10626) );
  XOR U11740 ( .A(n10627), .B(n10626), .Z(n10628) );
  XNOR U11741 ( .A(n10629), .B(n10628), .Z(n10631) );
  XNOR U11742 ( .A(sreg[1830]), .B(n10630), .Z(n10625) );
  XNOR U11743 ( .A(n10631), .B(n10625), .Z(c[1830]) );
  NAND U11744 ( .A(b[0]), .B(a[809]), .Z(n10634) );
  NAND U11745 ( .A(a[808]), .B(b[1]), .Z(n10633) );
  XNOR U11746 ( .A(n10634), .B(n10633), .Z(n10636) );
  XNOR U11747 ( .A(n10635), .B(n10636), .Z(n10640) );
  XOR U11748 ( .A(n10639), .B(sreg[1831]), .Z(n10632) );
  XNOR U11749 ( .A(n10640), .B(n10632), .Z(c[1831]) );
  NAND U11750 ( .A(n10634), .B(n10633), .Z(n10638) );
  NANDN U11751 ( .A(n10636), .B(n10635), .Z(n10637) );
  NAND U11752 ( .A(n10638), .B(n10637), .Z(n10644) );
  NAND U11753 ( .A(b[0]), .B(a[810]), .Z(n10643) );
  NAND U11754 ( .A(a[809]), .B(b[1]), .Z(n10642) );
  XNOR U11755 ( .A(n10643), .B(n10642), .Z(n10645) );
  XNOR U11756 ( .A(n10644), .B(n10645), .Z(n10649) );
  XOR U11757 ( .A(n10648), .B(sreg[1832]), .Z(n10641) );
  XNOR U11758 ( .A(n10649), .B(n10641), .Z(c[1832]) );
  NAND U11759 ( .A(n10643), .B(n10642), .Z(n10647) );
  NANDN U11760 ( .A(n10645), .B(n10644), .Z(n10646) );
  NAND U11761 ( .A(n10647), .B(n10646), .Z(n10653) );
  NAND U11762 ( .A(b[0]), .B(a[811]), .Z(n10652) );
  NAND U11763 ( .A(a[810]), .B(b[1]), .Z(n10651) );
  XNOR U11764 ( .A(n10652), .B(n10651), .Z(n10654) );
  XNOR U11765 ( .A(n10653), .B(n10654), .Z(n10658) );
  XOR U11766 ( .A(n10657), .B(sreg[1833]), .Z(n10650) );
  XNOR U11767 ( .A(n10658), .B(n10650), .Z(c[1833]) );
  NAND U11768 ( .A(n10652), .B(n10651), .Z(n10656) );
  NANDN U11769 ( .A(n10654), .B(n10653), .Z(n10655) );
  NAND U11770 ( .A(n10656), .B(n10655), .Z(n10663) );
  ANDN U11771 ( .B(a[812]), .A(n3974), .Z(n10661) );
  AND U11772 ( .A(b[1]), .B(a[811]), .Z(n10660) );
  XOR U11773 ( .A(n10661), .B(n10660), .Z(n10662) );
  XNOR U11774 ( .A(n10663), .B(n10662), .Z(n10668) );
  XOR U11775 ( .A(sreg[1834]), .B(n10667), .Z(n10659) );
  XNOR U11776 ( .A(n10668), .B(n10659), .Z(c[1834]) );
  OR U11777 ( .A(n10661), .B(n10660), .Z(n10666) );
  IV U11778 ( .A(n10662), .Z(n10664) );
  NANDN U11779 ( .A(n10664), .B(n10663), .Z(n10665) );
  NAND U11780 ( .A(n10666), .B(n10665), .Z(n10672) );
  NAND U11781 ( .A(b[0]), .B(a[813]), .Z(n10671) );
  NAND U11782 ( .A(a[812]), .B(b[1]), .Z(n10670) );
  XNOR U11783 ( .A(n10671), .B(n10670), .Z(n10673) );
  XNOR U11784 ( .A(n10672), .B(n10673), .Z(n10677) );
  XOR U11785 ( .A(n10676), .B(sreg[1835]), .Z(n10669) );
  XNOR U11786 ( .A(n10677), .B(n10669), .Z(c[1835]) );
  NAND U11787 ( .A(n10671), .B(n10670), .Z(n10675) );
  NANDN U11788 ( .A(n10673), .B(n10672), .Z(n10674) );
  NAND U11789 ( .A(n10675), .B(n10674), .Z(n10682) );
  ANDN U11790 ( .B(a[814]), .A(n3974), .Z(n10680) );
  AND U11791 ( .A(b[1]), .B(a[813]), .Z(n10679) );
  XOR U11792 ( .A(n10680), .B(n10679), .Z(n10681) );
  XNOR U11793 ( .A(n10682), .B(n10681), .Z(n10684) );
  XOR U11794 ( .A(sreg[1836]), .B(n10683), .Z(n10678) );
  XNOR U11795 ( .A(n10684), .B(n10678), .Z(c[1836]) );
  ANDN U11796 ( .B(a[815]), .A(n3974), .Z(n10687) );
  AND U11797 ( .A(b[1]), .B(a[814]), .Z(n10686) );
  XOR U11798 ( .A(n10687), .B(n10686), .Z(n10688) );
  XNOR U11799 ( .A(n10689), .B(n10688), .Z(n10691) );
  XNOR U11800 ( .A(sreg[1837]), .B(n10690), .Z(n10685) );
  XNOR U11801 ( .A(n10691), .B(n10685), .Z(c[1837]) );
  ANDN U11802 ( .B(a[816]), .A(n3974), .Z(n10694) );
  AND U11803 ( .A(b[1]), .B(a[815]), .Z(n10693) );
  XOR U11804 ( .A(n10694), .B(n10693), .Z(n10695) );
  XNOR U11805 ( .A(n10696), .B(n10695), .Z(n10698) );
  XNOR U11806 ( .A(sreg[1838]), .B(n10697), .Z(n10692) );
  XNOR U11807 ( .A(n10698), .B(n10692), .Z(c[1838]) );
  NAND U11808 ( .A(b[0]), .B(a[817]), .Z(n10701) );
  NAND U11809 ( .A(a[816]), .B(b[1]), .Z(n10700) );
  XNOR U11810 ( .A(n10701), .B(n10700), .Z(n10703) );
  XNOR U11811 ( .A(n10702), .B(n10703), .Z(n10707) );
  XOR U11812 ( .A(n10706), .B(sreg[1839]), .Z(n10699) );
  XNOR U11813 ( .A(n10707), .B(n10699), .Z(c[1839]) );
  NAND U11814 ( .A(n10701), .B(n10700), .Z(n10705) );
  NANDN U11815 ( .A(n10703), .B(n10702), .Z(n10704) );
  NAND U11816 ( .A(n10705), .B(n10704), .Z(n10712) );
  ANDN U11817 ( .B(a[818]), .A(n3974), .Z(n10710) );
  AND U11818 ( .A(b[1]), .B(a[817]), .Z(n10709) );
  XOR U11819 ( .A(n10710), .B(n10709), .Z(n10711) );
  XNOR U11820 ( .A(n10712), .B(n10711), .Z(n10714) );
  XOR U11821 ( .A(sreg[1840]), .B(n10713), .Z(n10708) );
  XNOR U11822 ( .A(n10714), .B(n10708), .Z(c[1840]) );
  NAND U11823 ( .A(b[0]), .B(a[819]), .Z(n10717) );
  NAND U11824 ( .A(a[818]), .B(b[1]), .Z(n10716) );
  XNOR U11825 ( .A(n10717), .B(n10716), .Z(n10719) );
  XNOR U11826 ( .A(n10718), .B(n10719), .Z(n10723) );
  XOR U11827 ( .A(n10722), .B(sreg[1841]), .Z(n10715) );
  XNOR U11828 ( .A(n10723), .B(n10715), .Z(c[1841]) );
  NAND U11829 ( .A(n10717), .B(n10716), .Z(n10721) );
  NANDN U11830 ( .A(n10719), .B(n10718), .Z(n10720) );
  NAND U11831 ( .A(n10721), .B(n10720), .Z(n10728) );
  ANDN U11832 ( .B(a[820]), .A(n3974), .Z(n10726) );
  AND U11833 ( .A(b[1]), .B(a[819]), .Z(n10725) );
  XOR U11834 ( .A(n10726), .B(n10725), .Z(n10727) );
  XNOR U11835 ( .A(n10728), .B(n10727), .Z(n10730) );
  XOR U11836 ( .A(sreg[1842]), .B(n10729), .Z(n10724) );
  XNOR U11837 ( .A(n10730), .B(n10724), .Z(c[1842]) );
  ANDN U11838 ( .B(a[821]), .A(n3974), .Z(n10733) );
  AND U11839 ( .A(b[1]), .B(a[820]), .Z(n10732) );
  XOR U11840 ( .A(n10733), .B(n10732), .Z(n10734) );
  XNOR U11841 ( .A(n10735), .B(n10734), .Z(n10737) );
  XNOR U11842 ( .A(sreg[1843]), .B(n10736), .Z(n10731) );
  XNOR U11843 ( .A(n10737), .B(n10731), .Z(c[1843]) );
  NAND U11844 ( .A(b[0]), .B(a[822]), .Z(n10740) );
  NAND U11845 ( .A(a[821]), .B(b[1]), .Z(n10739) );
  XNOR U11846 ( .A(n10740), .B(n10739), .Z(n10742) );
  XNOR U11847 ( .A(n10741), .B(n10742), .Z(n10746) );
  XOR U11848 ( .A(n10745), .B(sreg[1844]), .Z(n10738) );
  XNOR U11849 ( .A(n10746), .B(n10738), .Z(c[1844]) );
  NAND U11850 ( .A(n10740), .B(n10739), .Z(n10744) );
  NANDN U11851 ( .A(n10742), .B(n10741), .Z(n10743) );
  NAND U11852 ( .A(n10744), .B(n10743), .Z(n10750) );
  NAND U11853 ( .A(b[0]), .B(a[823]), .Z(n10749) );
  NAND U11854 ( .A(a[822]), .B(b[1]), .Z(n10748) );
  XNOR U11855 ( .A(n10749), .B(n10748), .Z(n10751) );
  XNOR U11856 ( .A(n10750), .B(n10751), .Z(n10755) );
  XOR U11857 ( .A(n10754), .B(sreg[1845]), .Z(n10747) );
  XNOR U11858 ( .A(n10755), .B(n10747), .Z(c[1845]) );
  NAND U11859 ( .A(n10749), .B(n10748), .Z(n10753) );
  NANDN U11860 ( .A(n10751), .B(n10750), .Z(n10752) );
  NAND U11861 ( .A(n10753), .B(n10752), .Z(n10760) );
  ANDN U11862 ( .B(a[824]), .A(n3975), .Z(n10758) );
  AND U11863 ( .A(b[1]), .B(a[823]), .Z(n10757) );
  XOR U11864 ( .A(n10758), .B(n10757), .Z(n10759) );
  XNOR U11865 ( .A(n10760), .B(n10759), .Z(n10765) );
  XOR U11866 ( .A(sreg[1846]), .B(n10764), .Z(n10756) );
  XNOR U11867 ( .A(n10765), .B(n10756), .Z(c[1846]) );
  OR U11868 ( .A(n10758), .B(n10757), .Z(n10763) );
  IV U11869 ( .A(n10759), .Z(n10761) );
  NANDN U11870 ( .A(n10761), .B(n10760), .Z(n10762) );
  NAND U11871 ( .A(n10763), .B(n10762), .Z(n10769) );
  NAND U11872 ( .A(b[0]), .B(a[825]), .Z(n10768) );
  NAND U11873 ( .A(a[824]), .B(b[1]), .Z(n10767) );
  XNOR U11874 ( .A(n10768), .B(n10767), .Z(n10770) );
  XNOR U11875 ( .A(n10769), .B(n10770), .Z(n10774) );
  XOR U11876 ( .A(n10773), .B(sreg[1847]), .Z(n10766) );
  XNOR U11877 ( .A(n10774), .B(n10766), .Z(c[1847]) );
  NAND U11878 ( .A(n10768), .B(n10767), .Z(n10772) );
  NANDN U11879 ( .A(n10770), .B(n10769), .Z(n10771) );
  NAND U11880 ( .A(n10772), .B(n10771), .Z(n10778) );
  NAND U11881 ( .A(b[0]), .B(a[826]), .Z(n10777) );
  NAND U11882 ( .A(a[825]), .B(b[1]), .Z(n10776) );
  XNOR U11883 ( .A(n10777), .B(n10776), .Z(n10779) );
  XNOR U11884 ( .A(n10778), .B(n10779), .Z(n10783) );
  XOR U11885 ( .A(n10782), .B(sreg[1848]), .Z(n10775) );
  XNOR U11886 ( .A(n10783), .B(n10775), .Z(c[1848]) );
  NAND U11887 ( .A(n10777), .B(n10776), .Z(n10781) );
  NANDN U11888 ( .A(n10779), .B(n10778), .Z(n10780) );
  NAND U11889 ( .A(n10781), .B(n10780), .Z(n10788) );
  ANDN U11890 ( .B(a[827]), .A(n3975), .Z(n10786) );
  AND U11891 ( .A(b[1]), .B(a[826]), .Z(n10785) );
  XOR U11892 ( .A(n10786), .B(n10785), .Z(n10787) );
  XNOR U11893 ( .A(n10788), .B(n10787), .Z(n10790) );
  XOR U11894 ( .A(sreg[1849]), .B(n10789), .Z(n10784) );
  XNOR U11895 ( .A(n10790), .B(n10784), .Z(c[1849]) );
  NAND U11896 ( .A(b[0]), .B(a[828]), .Z(n10793) );
  NAND U11897 ( .A(a[827]), .B(b[1]), .Z(n10792) );
  XNOR U11898 ( .A(n10793), .B(n10792), .Z(n10795) );
  XNOR U11899 ( .A(n10794), .B(n10795), .Z(n10799) );
  XOR U11900 ( .A(n10798), .B(sreg[1850]), .Z(n10791) );
  XNOR U11901 ( .A(n10799), .B(n10791), .Z(c[1850]) );
  NAND U11902 ( .A(n10793), .B(n10792), .Z(n10797) );
  NANDN U11903 ( .A(n10795), .B(n10794), .Z(n10796) );
  NAND U11904 ( .A(n10797), .B(n10796), .Z(n10803) );
  NAND U11905 ( .A(b[0]), .B(a[829]), .Z(n10802) );
  NAND U11906 ( .A(a[828]), .B(b[1]), .Z(n10801) );
  XNOR U11907 ( .A(n10802), .B(n10801), .Z(n10804) );
  XNOR U11908 ( .A(n10803), .B(n10804), .Z(n10808) );
  XOR U11909 ( .A(n10807), .B(sreg[1851]), .Z(n10800) );
  XNOR U11910 ( .A(n10808), .B(n10800), .Z(c[1851]) );
  NAND U11911 ( .A(n10802), .B(n10801), .Z(n10806) );
  NANDN U11912 ( .A(n10804), .B(n10803), .Z(n10805) );
  NAND U11913 ( .A(n10806), .B(n10805), .Z(n10813) );
  ANDN U11914 ( .B(a[830]), .A(n3975), .Z(n10811) );
  AND U11915 ( .A(b[1]), .B(a[829]), .Z(n10810) );
  XOR U11916 ( .A(n10811), .B(n10810), .Z(n10812) );
  XNOR U11917 ( .A(n10813), .B(n10812), .Z(n10815) );
  XOR U11918 ( .A(sreg[1852]), .B(n10814), .Z(n10809) );
  XNOR U11919 ( .A(n10815), .B(n10809), .Z(c[1852]) );
  NAND U11920 ( .A(b[0]), .B(a[831]), .Z(n10818) );
  NAND U11921 ( .A(a[830]), .B(b[1]), .Z(n10817) );
  XNOR U11922 ( .A(n10818), .B(n10817), .Z(n10820) );
  XNOR U11923 ( .A(n10819), .B(n10820), .Z(n10824) );
  XOR U11924 ( .A(n10823), .B(sreg[1853]), .Z(n10816) );
  XNOR U11925 ( .A(n10824), .B(n10816), .Z(c[1853]) );
  NAND U11926 ( .A(n10818), .B(n10817), .Z(n10822) );
  NANDN U11927 ( .A(n10820), .B(n10819), .Z(n10821) );
  NAND U11928 ( .A(n10822), .B(n10821), .Z(n10829) );
  ANDN U11929 ( .B(a[832]), .A(n3975), .Z(n10827) );
  AND U11930 ( .A(b[1]), .B(a[831]), .Z(n10826) );
  XOR U11931 ( .A(n10827), .B(n10826), .Z(n10828) );
  XNOR U11932 ( .A(n10829), .B(n10828), .Z(n10831) );
  XOR U11933 ( .A(sreg[1854]), .B(n10830), .Z(n10825) );
  XNOR U11934 ( .A(n10831), .B(n10825), .Z(c[1854]) );
  NAND U11935 ( .A(b[0]), .B(a[833]), .Z(n10834) );
  NAND U11936 ( .A(a[832]), .B(b[1]), .Z(n10833) );
  XNOR U11937 ( .A(n10834), .B(n10833), .Z(n10836) );
  XNOR U11938 ( .A(n10835), .B(n10836), .Z(n10840) );
  XOR U11939 ( .A(n10839), .B(sreg[1855]), .Z(n10832) );
  XNOR U11940 ( .A(n10840), .B(n10832), .Z(c[1855]) );
  NAND U11941 ( .A(n10834), .B(n10833), .Z(n10838) );
  NANDN U11942 ( .A(n10836), .B(n10835), .Z(n10837) );
  NAND U11943 ( .A(n10838), .B(n10837), .Z(n10845) );
  ANDN U11944 ( .B(a[834]), .A(n3975), .Z(n10843) );
  AND U11945 ( .A(b[1]), .B(a[833]), .Z(n10842) );
  XOR U11946 ( .A(n10843), .B(n10842), .Z(n10844) );
  XNOR U11947 ( .A(n10845), .B(n10844), .Z(n10847) );
  XOR U11948 ( .A(sreg[1856]), .B(n10846), .Z(n10841) );
  XNOR U11949 ( .A(n10847), .B(n10841), .Z(c[1856]) );
  NAND U11950 ( .A(b[0]), .B(a[835]), .Z(n10850) );
  NAND U11951 ( .A(a[834]), .B(b[1]), .Z(n10849) );
  XNOR U11952 ( .A(n10850), .B(n10849), .Z(n10852) );
  XNOR U11953 ( .A(n10851), .B(n10852), .Z(n10856) );
  XOR U11954 ( .A(n10855), .B(sreg[1857]), .Z(n10848) );
  XNOR U11955 ( .A(n10856), .B(n10848), .Z(c[1857]) );
  NAND U11956 ( .A(n10850), .B(n10849), .Z(n10854) );
  NANDN U11957 ( .A(n10852), .B(n10851), .Z(n10853) );
  NAND U11958 ( .A(n10854), .B(n10853), .Z(n10860) );
  NAND U11959 ( .A(b[0]), .B(a[836]), .Z(n10859) );
  NAND U11960 ( .A(a[835]), .B(b[1]), .Z(n10858) );
  XNOR U11961 ( .A(n10859), .B(n10858), .Z(n10861) );
  XNOR U11962 ( .A(n10860), .B(n10861), .Z(n10865) );
  XOR U11963 ( .A(n10864), .B(sreg[1858]), .Z(n10857) );
  XNOR U11964 ( .A(n10865), .B(n10857), .Z(c[1858]) );
  NAND U11965 ( .A(n10859), .B(n10858), .Z(n10863) );
  NANDN U11966 ( .A(n10861), .B(n10860), .Z(n10862) );
  NAND U11967 ( .A(n10863), .B(n10862), .Z(n10870) );
  ANDN U11968 ( .B(a[837]), .A(n3975), .Z(n10868) );
  AND U11969 ( .A(b[1]), .B(a[836]), .Z(n10867) );
  XOR U11970 ( .A(n10868), .B(n10867), .Z(n10869) );
  XNOR U11971 ( .A(n10870), .B(n10869), .Z(n10872) );
  XOR U11972 ( .A(sreg[1859]), .B(n10871), .Z(n10866) );
  XNOR U11973 ( .A(n10872), .B(n10866), .Z(c[1859]) );
  NAND U11974 ( .A(b[0]), .B(a[838]), .Z(n10875) );
  NAND U11975 ( .A(a[837]), .B(b[1]), .Z(n10874) );
  XNOR U11976 ( .A(n10875), .B(n10874), .Z(n10877) );
  XNOR U11977 ( .A(n10876), .B(n10877), .Z(n10881) );
  XOR U11978 ( .A(n10880), .B(sreg[1860]), .Z(n10873) );
  XNOR U11979 ( .A(n10881), .B(n10873), .Z(c[1860]) );
  NAND U11980 ( .A(n10875), .B(n10874), .Z(n10879) );
  NANDN U11981 ( .A(n10877), .B(n10876), .Z(n10878) );
  NAND U11982 ( .A(n10879), .B(n10878), .Z(n10885) );
  NAND U11983 ( .A(b[0]), .B(a[839]), .Z(n10884) );
  NAND U11984 ( .A(a[838]), .B(b[1]), .Z(n10883) );
  XNOR U11985 ( .A(n10884), .B(n10883), .Z(n10886) );
  XNOR U11986 ( .A(n10885), .B(n10886), .Z(n10890) );
  XOR U11987 ( .A(n10889), .B(sreg[1861]), .Z(n10882) );
  XNOR U11988 ( .A(n10890), .B(n10882), .Z(c[1861]) );
  NAND U11989 ( .A(n10884), .B(n10883), .Z(n10888) );
  NANDN U11990 ( .A(n10886), .B(n10885), .Z(n10887) );
  NAND U11991 ( .A(n10888), .B(n10887), .Z(n10894) );
  NAND U11992 ( .A(b[0]), .B(a[840]), .Z(n10893) );
  NAND U11993 ( .A(a[839]), .B(b[1]), .Z(n10892) );
  XNOR U11994 ( .A(n10893), .B(n10892), .Z(n10895) );
  XNOR U11995 ( .A(n10894), .B(n10895), .Z(n10899) );
  XOR U11996 ( .A(n10898), .B(sreg[1862]), .Z(n10891) );
  XNOR U11997 ( .A(n10899), .B(n10891), .Z(c[1862]) );
  NAND U11998 ( .A(n10893), .B(n10892), .Z(n10897) );
  NANDN U11999 ( .A(n10895), .B(n10894), .Z(n10896) );
  NAND U12000 ( .A(n10897), .B(n10896), .Z(n10904) );
  ANDN U12001 ( .B(a[841]), .A(n3975), .Z(n10902) );
  AND U12002 ( .A(b[1]), .B(a[840]), .Z(n10901) );
  XOR U12003 ( .A(n10902), .B(n10901), .Z(n10903) );
  XNOR U12004 ( .A(n10904), .B(n10903), .Z(n10906) );
  XOR U12005 ( .A(sreg[1863]), .B(n10905), .Z(n10900) );
  XNOR U12006 ( .A(n10906), .B(n10900), .Z(c[1863]) );
  NAND U12007 ( .A(b[0]), .B(a[842]), .Z(n10909) );
  NAND U12008 ( .A(a[841]), .B(b[1]), .Z(n10908) );
  XNOR U12009 ( .A(n10909), .B(n10908), .Z(n10911) );
  XNOR U12010 ( .A(n10910), .B(n10911), .Z(n10915) );
  XOR U12011 ( .A(n10914), .B(sreg[1864]), .Z(n10907) );
  XNOR U12012 ( .A(n10915), .B(n10907), .Z(c[1864]) );
  NAND U12013 ( .A(n10909), .B(n10908), .Z(n10913) );
  NANDN U12014 ( .A(n10911), .B(n10910), .Z(n10912) );
  NAND U12015 ( .A(n10913), .B(n10912), .Z(n10919) );
  NAND U12016 ( .A(b[0]), .B(a[843]), .Z(n10918) );
  NAND U12017 ( .A(a[842]), .B(b[1]), .Z(n10917) );
  XNOR U12018 ( .A(n10918), .B(n10917), .Z(n10920) );
  XNOR U12019 ( .A(n10919), .B(n10920), .Z(n10924) );
  XOR U12020 ( .A(n10923), .B(sreg[1865]), .Z(n10916) );
  XNOR U12021 ( .A(n10924), .B(n10916), .Z(c[1865]) );
  NAND U12022 ( .A(n10918), .B(n10917), .Z(n10922) );
  NANDN U12023 ( .A(n10920), .B(n10919), .Z(n10921) );
  NAND U12024 ( .A(n10922), .B(n10921), .Z(n10929) );
  ANDN U12025 ( .B(a[844]), .A(n3976), .Z(n10927) );
  AND U12026 ( .A(b[1]), .B(a[843]), .Z(n10926) );
  XOR U12027 ( .A(n10927), .B(n10926), .Z(n10928) );
  XNOR U12028 ( .A(n10929), .B(n10928), .Z(n10934) );
  XOR U12029 ( .A(sreg[1866]), .B(n10933), .Z(n10925) );
  XNOR U12030 ( .A(n10934), .B(n10925), .Z(c[1866]) );
  OR U12031 ( .A(n10927), .B(n10926), .Z(n10932) );
  IV U12032 ( .A(n10928), .Z(n10930) );
  NANDN U12033 ( .A(n10930), .B(n10929), .Z(n10931) );
  NAND U12034 ( .A(n10932), .B(n10931), .Z(n10938) );
  NAND U12035 ( .A(b[0]), .B(a[845]), .Z(n10937) );
  NAND U12036 ( .A(a[844]), .B(b[1]), .Z(n10936) );
  XNOR U12037 ( .A(n10937), .B(n10936), .Z(n10939) );
  XNOR U12038 ( .A(n10938), .B(n10939), .Z(n10943) );
  XOR U12039 ( .A(n10942), .B(sreg[1867]), .Z(n10935) );
  XNOR U12040 ( .A(n10943), .B(n10935), .Z(c[1867]) );
  NAND U12041 ( .A(n10937), .B(n10936), .Z(n10941) );
  NANDN U12042 ( .A(n10939), .B(n10938), .Z(n10940) );
  NAND U12043 ( .A(n10941), .B(n10940), .Z(n10948) );
  ANDN U12044 ( .B(a[846]), .A(n3976), .Z(n10946) );
  AND U12045 ( .A(b[1]), .B(a[845]), .Z(n10945) );
  XOR U12046 ( .A(n10946), .B(n10945), .Z(n10947) );
  XNOR U12047 ( .A(n10948), .B(n10947), .Z(n10950) );
  XOR U12048 ( .A(sreg[1868]), .B(n10949), .Z(n10944) );
  XNOR U12049 ( .A(n10950), .B(n10944), .Z(c[1868]) );
  NAND U12050 ( .A(b[0]), .B(a[847]), .Z(n10953) );
  NAND U12051 ( .A(a[846]), .B(b[1]), .Z(n10952) );
  XNOR U12052 ( .A(n10953), .B(n10952), .Z(n10955) );
  XNOR U12053 ( .A(n10954), .B(n10955), .Z(n10959) );
  XOR U12054 ( .A(n10958), .B(sreg[1869]), .Z(n10951) );
  XNOR U12055 ( .A(n10959), .B(n10951), .Z(c[1869]) );
  NAND U12056 ( .A(n10953), .B(n10952), .Z(n10957) );
  NANDN U12057 ( .A(n10955), .B(n10954), .Z(n10956) );
  NAND U12058 ( .A(n10957), .B(n10956), .Z(n10964) );
  ANDN U12059 ( .B(a[848]), .A(n3976), .Z(n10962) );
  AND U12060 ( .A(b[1]), .B(a[847]), .Z(n10961) );
  XOR U12061 ( .A(n10962), .B(n10961), .Z(n10963) );
  XNOR U12062 ( .A(n10964), .B(n10963), .Z(n10966) );
  XOR U12063 ( .A(sreg[1870]), .B(n10965), .Z(n10960) );
  XNOR U12064 ( .A(n10966), .B(n10960), .Z(c[1870]) );
  NAND U12065 ( .A(b[0]), .B(a[849]), .Z(n10969) );
  NAND U12066 ( .A(a[848]), .B(b[1]), .Z(n10968) );
  XNOR U12067 ( .A(n10969), .B(n10968), .Z(n10971) );
  XNOR U12068 ( .A(n10970), .B(n10971), .Z(n10975) );
  XOR U12069 ( .A(n10974), .B(sreg[1871]), .Z(n10967) );
  XNOR U12070 ( .A(n10975), .B(n10967), .Z(c[1871]) );
  NAND U12071 ( .A(n10969), .B(n10968), .Z(n10973) );
  NANDN U12072 ( .A(n10971), .B(n10970), .Z(n10972) );
  NAND U12073 ( .A(n10973), .B(n10972), .Z(n10980) );
  ANDN U12074 ( .B(a[850]), .A(n3976), .Z(n10978) );
  AND U12075 ( .A(b[1]), .B(a[849]), .Z(n10977) );
  XOR U12076 ( .A(n10978), .B(n10977), .Z(n10979) );
  XNOR U12077 ( .A(n10980), .B(n10979), .Z(n10982) );
  XOR U12078 ( .A(sreg[1872]), .B(n10981), .Z(n10976) );
  XNOR U12079 ( .A(n10982), .B(n10976), .Z(c[1872]) );
  ANDN U12080 ( .B(a[851]), .A(n3976), .Z(n10985) );
  AND U12081 ( .A(b[1]), .B(a[850]), .Z(n10984) );
  XOR U12082 ( .A(n10985), .B(n10984), .Z(n10986) );
  XNOR U12083 ( .A(n10987), .B(n10986), .Z(n10989) );
  XNOR U12084 ( .A(sreg[1873]), .B(n10988), .Z(n10983) );
  XNOR U12085 ( .A(n10989), .B(n10983), .Z(c[1873]) );
  ANDN U12086 ( .B(a[852]), .A(n3976), .Z(n10992) );
  AND U12087 ( .A(b[1]), .B(a[851]), .Z(n10991) );
  XOR U12088 ( .A(n10992), .B(n10991), .Z(n10993) );
  XNOR U12089 ( .A(n10994), .B(n10993), .Z(n10996) );
  XNOR U12090 ( .A(sreg[1874]), .B(n10995), .Z(n10990) );
  XNOR U12091 ( .A(n10996), .B(n10990), .Z(c[1874]) );
  NAND U12092 ( .A(b[0]), .B(a[853]), .Z(n10999) );
  NAND U12093 ( .A(a[852]), .B(b[1]), .Z(n10998) );
  XNOR U12094 ( .A(n10999), .B(n10998), .Z(n11001) );
  XNOR U12095 ( .A(n11000), .B(n11001), .Z(n11005) );
  XOR U12096 ( .A(n11004), .B(sreg[1875]), .Z(n10997) );
  XNOR U12097 ( .A(n11005), .B(n10997), .Z(c[1875]) );
  NAND U12098 ( .A(n10999), .B(n10998), .Z(n11003) );
  NANDN U12099 ( .A(n11001), .B(n11000), .Z(n11002) );
  NAND U12100 ( .A(n11003), .B(n11002), .Z(n11009) );
  NAND U12101 ( .A(b[0]), .B(a[854]), .Z(n11008) );
  NAND U12102 ( .A(a[853]), .B(b[1]), .Z(n11007) );
  XNOR U12103 ( .A(n11008), .B(n11007), .Z(n11010) );
  XNOR U12104 ( .A(n11009), .B(n11010), .Z(n11014) );
  XOR U12105 ( .A(n11013), .B(sreg[1876]), .Z(n11006) );
  XNOR U12106 ( .A(n11014), .B(n11006), .Z(c[1876]) );
  NAND U12107 ( .A(n11008), .B(n11007), .Z(n11012) );
  NANDN U12108 ( .A(n11010), .B(n11009), .Z(n11011) );
  NAND U12109 ( .A(n11012), .B(n11011), .Z(n11018) );
  NAND U12110 ( .A(b[0]), .B(a[855]), .Z(n11017) );
  NAND U12111 ( .A(a[854]), .B(b[1]), .Z(n11016) );
  XNOR U12112 ( .A(n11017), .B(n11016), .Z(n11019) );
  XNOR U12113 ( .A(n11018), .B(n11019), .Z(n11023) );
  XOR U12114 ( .A(n11022), .B(sreg[1877]), .Z(n11015) );
  XNOR U12115 ( .A(n11023), .B(n11015), .Z(c[1877]) );
  NAND U12116 ( .A(n11017), .B(n11016), .Z(n11021) );
  NANDN U12117 ( .A(n11019), .B(n11018), .Z(n11020) );
  NAND U12118 ( .A(n11021), .B(n11020), .Z(n11027) );
  NAND U12119 ( .A(b[0]), .B(a[856]), .Z(n11026) );
  NAND U12120 ( .A(a[855]), .B(b[1]), .Z(n11025) );
  XNOR U12121 ( .A(n11026), .B(n11025), .Z(n11028) );
  XNOR U12122 ( .A(n11027), .B(n11028), .Z(n11032) );
  XOR U12123 ( .A(n11031), .B(sreg[1878]), .Z(n11024) );
  XNOR U12124 ( .A(n11032), .B(n11024), .Z(c[1878]) );
  NAND U12125 ( .A(n11026), .B(n11025), .Z(n11030) );
  NANDN U12126 ( .A(n11028), .B(n11027), .Z(n11029) );
  NAND U12127 ( .A(n11030), .B(n11029), .Z(n11036) );
  NAND U12128 ( .A(b[0]), .B(a[857]), .Z(n11035) );
  NAND U12129 ( .A(a[856]), .B(b[1]), .Z(n11034) );
  XNOR U12130 ( .A(n11035), .B(n11034), .Z(n11037) );
  XNOR U12131 ( .A(n11036), .B(n11037), .Z(n11041) );
  XOR U12132 ( .A(n11040), .B(sreg[1879]), .Z(n11033) );
  XNOR U12133 ( .A(n11041), .B(n11033), .Z(c[1879]) );
  NAND U12134 ( .A(n11035), .B(n11034), .Z(n11039) );
  NANDN U12135 ( .A(n11037), .B(n11036), .Z(n11038) );
  NAND U12136 ( .A(n11039), .B(n11038), .Z(n11045) );
  NAND U12137 ( .A(b[0]), .B(a[858]), .Z(n11044) );
  NAND U12138 ( .A(a[857]), .B(b[1]), .Z(n11043) );
  XNOR U12139 ( .A(n11044), .B(n11043), .Z(n11046) );
  XNOR U12140 ( .A(n11045), .B(n11046), .Z(n11050) );
  XOR U12141 ( .A(n11049), .B(sreg[1880]), .Z(n11042) );
  XNOR U12142 ( .A(n11050), .B(n11042), .Z(c[1880]) );
  NAND U12143 ( .A(n11044), .B(n11043), .Z(n11048) );
  NANDN U12144 ( .A(n11046), .B(n11045), .Z(n11047) );
  NAND U12145 ( .A(n11048), .B(n11047), .Z(n11054) );
  NAND U12146 ( .A(b[0]), .B(a[859]), .Z(n11053) );
  NAND U12147 ( .A(a[858]), .B(b[1]), .Z(n11052) );
  XNOR U12148 ( .A(n11053), .B(n11052), .Z(n11055) );
  XNOR U12149 ( .A(n11054), .B(n11055), .Z(n11059) );
  XOR U12150 ( .A(n11058), .B(sreg[1881]), .Z(n11051) );
  XNOR U12151 ( .A(n11059), .B(n11051), .Z(c[1881]) );
  NAND U12152 ( .A(n11053), .B(n11052), .Z(n11057) );
  NANDN U12153 ( .A(n11055), .B(n11054), .Z(n11056) );
  NAND U12154 ( .A(n11057), .B(n11056), .Z(n11064) );
  ANDN U12155 ( .B(a[860]), .A(n3976), .Z(n11062) );
  AND U12156 ( .A(b[1]), .B(a[859]), .Z(n11061) );
  XOR U12157 ( .A(n11062), .B(n11061), .Z(n11063) );
  XNOR U12158 ( .A(n11064), .B(n11063), .Z(n11066) );
  XOR U12159 ( .A(sreg[1882]), .B(n11065), .Z(n11060) );
  XNOR U12160 ( .A(n11066), .B(n11060), .Z(c[1882]) );
  NAND U12161 ( .A(b[0]), .B(a[861]), .Z(n11069) );
  NAND U12162 ( .A(a[860]), .B(b[1]), .Z(n11068) );
  XNOR U12163 ( .A(n11069), .B(n11068), .Z(n11071) );
  XNOR U12164 ( .A(n11070), .B(n11071), .Z(n11075) );
  XOR U12165 ( .A(n11074), .B(sreg[1883]), .Z(n11067) );
  XNOR U12166 ( .A(n11075), .B(n11067), .Z(c[1883]) );
  NAND U12167 ( .A(n11069), .B(n11068), .Z(n11073) );
  NANDN U12168 ( .A(n11071), .B(n11070), .Z(n11072) );
  NAND U12169 ( .A(n11073), .B(n11072), .Z(n11079) );
  NAND U12170 ( .A(b[0]), .B(a[862]), .Z(n11078) );
  NAND U12171 ( .A(a[861]), .B(b[1]), .Z(n11077) );
  XNOR U12172 ( .A(n11078), .B(n11077), .Z(n11080) );
  XNOR U12173 ( .A(n11079), .B(n11080), .Z(n11084) );
  XOR U12174 ( .A(n11083), .B(sreg[1884]), .Z(n11076) );
  XNOR U12175 ( .A(n11084), .B(n11076), .Z(c[1884]) );
  NAND U12176 ( .A(n11078), .B(n11077), .Z(n11082) );
  NANDN U12177 ( .A(n11080), .B(n11079), .Z(n11081) );
  NAND U12178 ( .A(n11082), .B(n11081), .Z(n11088) );
  NAND U12179 ( .A(b[0]), .B(a[863]), .Z(n11087) );
  NAND U12180 ( .A(a[862]), .B(b[1]), .Z(n11086) );
  XNOR U12181 ( .A(n11087), .B(n11086), .Z(n11089) );
  XNOR U12182 ( .A(n11088), .B(n11089), .Z(n11093) );
  XOR U12183 ( .A(n11092), .B(sreg[1885]), .Z(n11085) );
  XNOR U12184 ( .A(n11093), .B(n11085), .Z(c[1885]) );
  NAND U12185 ( .A(n11087), .B(n11086), .Z(n11091) );
  NANDN U12186 ( .A(n11089), .B(n11088), .Z(n11090) );
  NAND U12187 ( .A(n11091), .B(n11090), .Z(n11098) );
  ANDN U12188 ( .B(a[864]), .A(n3977), .Z(n11096) );
  AND U12189 ( .A(b[1]), .B(a[863]), .Z(n11095) );
  XOR U12190 ( .A(n11096), .B(n11095), .Z(n11097) );
  XNOR U12191 ( .A(n11098), .B(n11097), .Z(n11103) );
  XOR U12192 ( .A(sreg[1886]), .B(n11102), .Z(n11094) );
  XNOR U12193 ( .A(n11103), .B(n11094), .Z(c[1886]) );
  OR U12194 ( .A(n11096), .B(n11095), .Z(n11101) );
  IV U12195 ( .A(n11097), .Z(n11099) );
  NANDN U12196 ( .A(n11099), .B(n11098), .Z(n11100) );
  NAND U12197 ( .A(n11101), .B(n11100), .Z(n11107) );
  NAND U12198 ( .A(b[0]), .B(a[865]), .Z(n11106) );
  NAND U12199 ( .A(a[864]), .B(b[1]), .Z(n11105) );
  XNOR U12200 ( .A(n11106), .B(n11105), .Z(n11108) );
  XNOR U12201 ( .A(n11107), .B(n11108), .Z(n11112) );
  XOR U12202 ( .A(n11111), .B(sreg[1887]), .Z(n11104) );
  XNOR U12203 ( .A(n11112), .B(n11104), .Z(c[1887]) );
  NAND U12204 ( .A(n11106), .B(n11105), .Z(n11110) );
  NANDN U12205 ( .A(n11108), .B(n11107), .Z(n11109) );
  NAND U12206 ( .A(n11110), .B(n11109), .Z(n11117) );
  ANDN U12207 ( .B(a[866]), .A(n3977), .Z(n11115) );
  AND U12208 ( .A(b[1]), .B(a[865]), .Z(n11114) );
  XOR U12209 ( .A(n11115), .B(n11114), .Z(n11116) );
  XNOR U12210 ( .A(n11117), .B(n11116), .Z(n11119) );
  XOR U12211 ( .A(sreg[1888]), .B(n11118), .Z(n11113) );
  XNOR U12212 ( .A(n11119), .B(n11113), .Z(c[1888]) );
  NAND U12213 ( .A(b[0]), .B(a[867]), .Z(n11122) );
  NAND U12214 ( .A(a[866]), .B(b[1]), .Z(n11121) );
  XNOR U12215 ( .A(n11122), .B(n11121), .Z(n11124) );
  XNOR U12216 ( .A(n11123), .B(n11124), .Z(n11128) );
  XOR U12217 ( .A(n11127), .B(sreg[1889]), .Z(n11120) );
  XNOR U12218 ( .A(n11128), .B(n11120), .Z(c[1889]) );
  NAND U12219 ( .A(n11122), .B(n11121), .Z(n11126) );
  NANDN U12220 ( .A(n11124), .B(n11123), .Z(n11125) );
  NAND U12221 ( .A(n11126), .B(n11125), .Z(n11133) );
  ANDN U12222 ( .B(a[868]), .A(n3977), .Z(n11131) );
  AND U12223 ( .A(b[1]), .B(a[867]), .Z(n11130) );
  XOR U12224 ( .A(n11131), .B(n11130), .Z(n11132) );
  XNOR U12225 ( .A(n11133), .B(n11132), .Z(n11135) );
  XOR U12226 ( .A(sreg[1890]), .B(n11134), .Z(n11129) );
  XNOR U12227 ( .A(n11135), .B(n11129), .Z(c[1890]) );
  NAND U12228 ( .A(b[0]), .B(a[869]), .Z(n11138) );
  NAND U12229 ( .A(a[868]), .B(b[1]), .Z(n11137) );
  XNOR U12230 ( .A(n11138), .B(n11137), .Z(n11140) );
  XNOR U12231 ( .A(n11139), .B(n11140), .Z(n11144) );
  XOR U12232 ( .A(n11143), .B(sreg[1891]), .Z(n11136) );
  XNOR U12233 ( .A(n11144), .B(n11136), .Z(c[1891]) );
  NAND U12234 ( .A(n11138), .B(n11137), .Z(n11142) );
  NANDN U12235 ( .A(n11140), .B(n11139), .Z(n11141) );
  NAND U12236 ( .A(n11142), .B(n11141), .Z(n11149) );
  ANDN U12237 ( .B(a[870]), .A(n3977), .Z(n11147) );
  AND U12238 ( .A(b[1]), .B(a[869]), .Z(n11146) );
  XOR U12239 ( .A(n11147), .B(n11146), .Z(n11148) );
  XNOR U12240 ( .A(n11149), .B(n11148), .Z(n11151) );
  XOR U12241 ( .A(sreg[1892]), .B(n11150), .Z(n11145) );
  XNOR U12242 ( .A(n11151), .B(n11145), .Z(c[1892]) );
  NAND U12243 ( .A(b[0]), .B(a[871]), .Z(n11154) );
  NAND U12244 ( .A(a[870]), .B(b[1]), .Z(n11153) );
  XNOR U12245 ( .A(n11154), .B(n11153), .Z(n11156) );
  XNOR U12246 ( .A(n11155), .B(n11156), .Z(n11160) );
  XOR U12247 ( .A(n11159), .B(sreg[1893]), .Z(n11152) );
  XNOR U12248 ( .A(n11160), .B(n11152), .Z(c[1893]) );
  NAND U12249 ( .A(n11154), .B(n11153), .Z(n11158) );
  NANDN U12250 ( .A(n11156), .B(n11155), .Z(n11157) );
  NAND U12251 ( .A(n11158), .B(n11157), .Z(n11165) );
  ANDN U12252 ( .B(a[872]), .A(n3977), .Z(n11163) );
  AND U12253 ( .A(b[1]), .B(a[871]), .Z(n11162) );
  XOR U12254 ( .A(n11163), .B(n11162), .Z(n11164) );
  XNOR U12255 ( .A(n11165), .B(n11164), .Z(n11167) );
  XOR U12256 ( .A(sreg[1894]), .B(n11166), .Z(n11161) );
  XNOR U12257 ( .A(n11167), .B(n11161), .Z(c[1894]) );
  ANDN U12258 ( .B(a[873]), .A(n3977), .Z(n11170) );
  AND U12259 ( .A(b[1]), .B(a[872]), .Z(n11169) );
  XOR U12260 ( .A(n11170), .B(n11169), .Z(n11171) );
  XNOR U12261 ( .A(n11172), .B(n11171), .Z(n11174) );
  XNOR U12262 ( .A(sreg[1895]), .B(n11173), .Z(n11168) );
  XNOR U12263 ( .A(n11174), .B(n11168), .Z(c[1895]) );
  ANDN U12264 ( .B(a[874]), .A(n3977), .Z(n11177) );
  AND U12265 ( .A(b[1]), .B(a[873]), .Z(n11176) );
  XOR U12266 ( .A(n11177), .B(n11176), .Z(n11178) );
  XNOR U12267 ( .A(n11179), .B(n11178), .Z(n11181) );
  XNOR U12268 ( .A(sreg[1896]), .B(n11180), .Z(n11175) );
  XNOR U12269 ( .A(n11181), .B(n11175), .Z(c[1896]) );
  NAND U12270 ( .A(b[0]), .B(a[875]), .Z(n11184) );
  NAND U12271 ( .A(a[874]), .B(b[1]), .Z(n11183) );
  XNOR U12272 ( .A(n11184), .B(n11183), .Z(n11186) );
  XNOR U12273 ( .A(n11185), .B(n11186), .Z(n11190) );
  XOR U12274 ( .A(n11189), .B(sreg[1897]), .Z(n11182) );
  XNOR U12275 ( .A(n11190), .B(n11182), .Z(c[1897]) );
  NAND U12276 ( .A(n11184), .B(n11183), .Z(n11188) );
  NANDN U12277 ( .A(n11186), .B(n11185), .Z(n11187) );
  NAND U12278 ( .A(n11188), .B(n11187), .Z(n11195) );
  ANDN U12279 ( .B(a[876]), .A(n3978), .Z(n11193) );
  AND U12280 ( .A(b[1]), .B(a[875]), .Z(n11192) );
  XOR U12281 ( .A(n11193), .B(n11192), .Z(n11194) );
  XNOR U12282 ( .A(n11195), .B(n11194), .Z(n11200) );
  XOR U12283 ( .A(sreg[1898]), .B(n11199), .Z(n11191) );
  XNOR U12284 ( .A(n11200), .B(n11191), .Z(c[1898]) );
  OR U12285 ( .A(n11193), .B(n11192), .Z(n11198) );
  IV U12286 ( .A(n11194), .Z(n11196) );
  NANDN U12287 ( .A(n11196), .B(n11195), .Z(n11197) );
  NAND U12288 ( .A(n11198), .B(n11197), .Z(n11205) );
  ANDN U12289 ( .B(a[877]), .A(n3978), .Z(n11203) );
  AND U12290 ( .A(b[1]), .B(a[876]), .Z(n11202) );
  XOR U12291 ( .A(n11203), .B(n11202), .Z(n11204) );
  XNOR U12292 ( .A(n11205), .B(n11204), .Z(n11207) );
  XNOR U12293 ( .A(sreg[1899]), .B(n11206), .Z(n11201) );
  XNOR U12294 ( .A(n11207), .B(n11201), .Z(c[1899]) );
  ANDN U12295 ( .B(a[878]), .A(n3978), .Z(n11210) );
  AND U12296 ( .A(b[1]), .B(a[877]), .Z(n11209) );
  XOR U12297 ( .A(n11210), .B(n11209), .Z(n11211) );
  XNOR U12298 ( .A(n11212), .B(n11211), .Z(n11214) );
  XNOR U12299 ( .A(sreg[1900]), .B(n11213), .Z(n11208) );
  XNOR U12300 ( .A(n11214), .B(n11208), .Z(c[1900]) );
  NAND U12301 ( .A(b[0]), .B(a[879]), .Z(n11217) );
  NAND U12302 ( .A(a[878]), .B(b[1]), .Z(n11216) );
  XNOR U12303 ( .A(n11217), .B(n11216), .Z(n11219) );
  XNOR U12304 ( .A(n11218), .B(n11219), .Z(n11223) );
  XOR U12305 ( .A(n11222), .B(sreg[1901]), .Z(n11215) );
  XNOR U12306 ( .A(n11223), .B(n11215), .Z(c[1901]) );
  NAND U12307 ( .A(n11217), .B(n11216), .Z(n11221) );
  NANDN U12308 ( .A(n11219), .B(n11218), .Z(n11220) );
  NAND U12309 ( .A(n11221), .B(n11220), .Z(n11228) );
  ANDN U12310 ( .B(a[880]), .A(n3978), .Z(n11226) );
  AND U12311 ( .A(b[1]), .B(a[879]), .Z(n11225) );
  XOR U12312 ( .A(n11226), .B(n11225), .Z(n11227) );
  XNOR U12313 ( .A(n11228), .B(n11227), .Z(n11230) );
  XOR U12314 ( .A(sreg[1902]), .B(n11229), .Z(n11224) );
  XNOR U12315 ( .A(n11230), .B(n11224), .Z(c[1902]) );
  NAND U12316 ( .A(b[0]), .B(a[881]), .Z(n11233) );
  NAND U12317 ( .A(a[880]), .B(b[1]), .Z(n11232) );
  XNOR U12318 ( .A(n11233), .B(n11232), .Z(n11235) );
  XNOR U12319 ( .A(n11234), .B(n11235), .Z(n11239) );
  XOR U12320 ( .A(n11238), .B(sreg[1903]), .Z(n11231) );
  XNOR U12321 ( .A(n11239), .B(n11231), .Z(c[1903]) );
  NAND U12322 ( .A(n11233), .B(n11232), .Z(n11237) );
  NANDN U12323 ( .A(n11235), .B(n11234), .Z(n11236) );
  NAND U12324 ( .A(n11237), .B(n11236), .Z(n11244) );
  ANDN U12325 ( .B(a[882]), .A(n3978), .Z(n11242) );
  AND U12326 ( .A(b[1]), .B(a[881]), .Z(n11241) );
  XOR U12327 ( .A(n11242), .B(n11241), .Z(n11243) );
  XNOR U12328 ( .A(n11244), .B(n11243), .Z(n11246) );
  XOR U12329 ( .A(sreg[1904]), .B(n11245), .Z(n11240) );
  XNOR U12330 ( .A(n11246), .B(n11240), .Z(c[1904]) );
  NAND U12331 ( .A(b[0]), .B(a[883]), .Z(n11249) );
  NAND U12332 ( .A(a[882]), .B(b[1]), .Z(n11248) );
  XNOR U12333 ( .A(n11249), .B(n11248), .Z(n11251) );
  XNOR U12334 ( .A(n11250), .B(n11251), .Z(n11255) );
  XOR U12335 ( .A(n11254), .B(sreg[1905]), .Z(n11247) );
  XNOR U12336 ( .A(n11255), .B(n11247), .Z(c[1905]) );
  NAND U12337 ( .A(n11249), .B(n11248), .Z(n11253) );
  NANDN U12338 ( .A(n11251), .B(n11250), .Z(n11252) );
  NAND U12339 ( .A(n11253), .B(n11252), .Z(n11260) );
  ANDN U12340 ( .B(a[884]), .A(n3978), .Z(n11258) );
  AND U12341 ( .A(b[1]), .B(a[883]), .Z(n11257) );
  XOR U12342 ( .A(n11258), .B(n11257), .Z(n11259) );
  XNOR U12343 ( .A(n11260), .B(n11259), .Z(n11262) );
  XOR U12344 ( .A(sreg[1906]), .B(n11261), .Z(n11256) );
  XNOR U12345 ( .A(n11262), .B(n11256), .Z(c[1906]) );
  NAND U12346 ( .A(b[0]), .B(a[885]), .Z(n11265) );
  NAND U12347 ( .A(a[884]), .B(b[1]), .Z(n11264) );
  XNOR U12348 ( .A(n11265), .B(n11264), .Z(n11267) );
  XNOR U12349 ( .A(n11266), .B(n11267), .Z(n11271) );
  XOR U12350 ( .A(n11270), .B(sreg[1907]), .Z(n11263) );
  XNOR U12351 ( .A(n11271), .B(n11263), .Z(c[1907]) );
  NAND U12352 ( .A(n11265), .B(n11264), .Z(n11269) );
  NANDN U12353 ( .A(n11267), .B(n11266), .Z(n11268) );
  NAND U12354 ( .A(n11269), .B(n11268), .Z(n11276) );
  ANDN U12355 ( .B(a[886]), .A(n3978), .Z(n11274) );
  AND U12356 ( .A(b[1]), .B(a[885]), .Z(n11273) );
  XOR U12357 ( .A(n11274), .B(n11273), .Z(n11275) );
  XNOR U12358 ( .A(n11276), .B(n11275), .Z(n11278) );
  XOR U12359 ( .A(sreg[1908]), .B(n11277), .Z(n11272) );
  XNOR U12360 ( .A(n11278), .B(n11272), .Z(c[1908]) );
  NAND U12361 ( .A(b[0]), .B(a[887]), .Z(n11281) );
  NAND U12362 ( .A(a[886]), .B(b[1]), .Z(n11280) );
  XNOR U12363 ( .A(n11281), .B(n11280), .Z(n11283) );
  XNOR U12364 ( .A(n11282), .B(n11283), .Z(n11287) );
  XOR U12365 ( .A(n11286), .B(sreg[1909]), .Z(n11279) );
  XNOR U12366 ( .A(n11287), .B(n11279), .Z(c[1909]) );
  NAND U12367 ( .A(n11281), .B(n11280), .Z(n11285) );
  NANDN U12368 ( .A(n11283), .B(n11282), .Z(n11284) );
  NAND U12369 ( .A(n11285), .B(n11284), .Z(n11292) );
  ANDN U12370 ( .B(a[888]), .A(n3979), .Z(n11290) );
  AND U12371 ( .A(b[1]), .B(a[887]), .Z(n11289) );
  XOR U12372 ( .A(n11290), .B(n11289), .Z(n11291) );
  XNOR U12373 ( .A(n11292), .B(n11291), .Z(n11297) );
  XOR U12374 ( .A(sreg[1910]), .B(n11296), .Z(n11288) );
  XNOR U12375 ( .A(n11297), .B(n11288), .Z(c[1910]) );
  OR U12376 ( .A(n11290), .B(n11289), .Z(n11295) );
  IV U12377 ( .A(n11291), .Z(n11293) );
  NANDN U12378 ( .A(n11293), .B(n11292), .Z(n11294) );
  NAND U12379 ( .A(n11295), .B(n11294), .Z(n11301) );
  NAND U12380 ( .A(b[0]), .B(a[889]), .Z(n11300) );
  NAND U12381 ( .A(a[888]), .B(b[1]), .Z(n11299) );
  XNOR U12382 ( .A(n11300), .B(n11299), .Z(n11302) );
  XNOR U12383 ( .A(n11301), .B(n11302), .Z(n11306) );
  XOR U12384 ( .A(n11305), .B(sreg[1911]), .Z(n11298) );
  XNOR U12385 ( .A(n11306), .B(n11298), .Z(c[1911]) );
  NAND U12386 ( .A(n11300), .B(n11299), .Z(n11304) );
  NANDN U12387 ( .A(n11302), .B(n11301), .Z(n11303) );
  NAND U12388 ( .A(n11304), .B(n11303), .Z(n11311) );
  ANDN U12389 ( .B(a[890]), .A(n3979), .Z(n11309) );
  AND U12390 ( .A(b[1]), .B(a[889]), .Z(n11308) );
  XOR U12391 ( .A(n11309), .B(n11308), .Z(n11310) );
  XNOR U12392 ( .A(n11311), .B(n11310), .Z(n11313) );
  XOR U12393 ( .A(sreg[1912]), .B(n11312), .Z(n11307) );
  XNOR U12394 ( .A(n11313), .B(n11307), .Z(c[1912]) );
  NAND U12395 ( .A(b[0]), .B(a[891]), .Z(n11316) );
  NAND U12396 ( .A(a[890]), .B(b[1]), .Z(n11315) );
  XNOR U12397 ( .A(n11316), .B(n11315), .Z(n11318) );
  XNOR U12398 ( .A(n11317), .B(n11318), .Z(n11322) );
  XOR U12399 ( .A(n11321), .B(sreg[1913]), .Z(n11314) );
  XNOR U12400 ( .A(n11322), .B(n11314), .Z(c[1913]) );
  NAND U12401 ( .A(n11316), .B(n11315), .Z(n11320) );
  NANDN U12402 ( .A(n11318), .B(n11317), .Z(n11319) );
  NAND U12403 ( .A(n11320), .B(n11319), .Z(n11327) );
  ANDN U12404 ( .B(a[892]), .A(n3979), .Z(n11325) );
  AND U12405 ( .A(b[1]), .B(a[891]), .Z(n11324) );
  XOR U12406 ( .A(n11325), .B(n11324), .Z(n11326) );
  XNOR U12407 ( .A(n11327), .B(n11326), .Z(n11329) );
  XOR U12408 ( .A(sreg[1914]), .B(n11328), .Z(n11323) );
  XNOR U12409 ( .A(n11329), .B(n11323), .Z(c[1914]) );
  NAND U12410 ( .A(b[0]), .B(a[893]), .Z(n11332) );
  NAND U12411 ( .A(a[892]), .B(b[1]), .Z(n11331) );
  XNOR U12412 ( .A(n11332), .B(n11331), .Z(n11334) );
  XNOR U12413 ( .A(n11333), .B(n11334), .Z(n11338) );
  XOR U12414 ( .A(n11337), .B(sreg[1915]), .Z(n11330) );
  XNOR U12415 ( .A(n11338), .B(n11330), .Z(c[1915]) );
  NAND U12416 ( .A(n11332), .B(n11331), .Z(n11336) );
  NANDN U12417 ( .A(n11334), .B(n11333), .Z(n11335) );
  NAND U12418 ( .A(n11336), .B(n11335), .Z(n11343) );
  ANDN U12419 ( .B(a[894]), .A(n3979), .Z(n11341) );
  AND U12420 ( .A(b[1]), .B(a[893]), .Z(n11340) );
  XOR U12421 ( .A(n11341), .B(n11340), .Z(n11342) );
  XNOR U12422 ( .A(n11343), .B(n11342), .Z(n11345) );
  XOR U12423 ( .A(sreg[1916]), .B(n11344), .Z(n11339) );
  XNOR U12424 ( .A(n11345), .B(n11339), .Z(c[1916]) );
  NAND U12425 ( .A(b[0]), .B(a[895]), .Z(n11348) );
  NAND U12426 ( .A(a[894]), .B(b[1]), .Z(n11347) );
  XNOR U12427 ( .A(n11348), .B(n11347), .Z(n11350) );
  XNOR U12428 ( .A(n11349), .B(n11350), .Z(n11354) );
  XOR U12429 ( .A(n11353), .B(sreg[1917]), .Z(n11346) );
  XNOR U12430 ( .A(n11354), .B(n11346), .Z(c[1917]) );
  NAND U12431 ( .A(n11348), .B(n11347), .Z(n11352) );
  NANDN U12432 ( .A(n11350), .B(n11349), .Z(n11351) );
  NAND U12433 ( .A(n11352), .B(n11351), .Z(n11358) );
  NAND U12434 ( .A(b[0]), .B(a[896]), .Z(n11357) );
  NAND U12435 ( .A(a[895]), .B(b[1]), .Z(n11356) );
  XNOR U12436 ( .A(n11357), .B(n11356), .Z(n11359) );
  XNOR U12437 ( .A(n11358), .B(n11359), .Z(n11363) );
  XOR U12438 ( .A(n11362), .B(sreg[1918]), .Z(n11355) );
  XNOR U12439 ( .A(n11363), .B(n11355), .Z(c[1918]) );
  NAND U12440 ( .A(n11357), .B(n11356), .Z(n11361) );
  NANDN U12441 ( .A(n11359), .B(n11358), .Z(n11360) );
  NAND U12442 ( .A(n11361), .B(n11360), .Z(n11367) );
  NAND U12443 ( .A(b[0]), .B(a[897]), .Z(n11366) );
  NAND U12444 ( .A(a[896]), .B(b[1]), .Z(n11365) );
  XNOR U12445 ( .A(n11366), .B(n11365), .Z(n11368) );
  XNOR U12446 ( .A(n11367), .B(n11368), .Z(n11372) );
  XOR U12447 ( .A(n11371), .B(sreg[1919]), .Z(n11364) );
  XNOR U12448 ( .A(n11372), .B(n11364), .Z(c[1919]) );
  NAND U12449 ( .A(n11366), .B(n11365), .Z(n11370) );
  NANDN U12450 ( .A(n11368), .B(n11367), .Z(n11369) );
  NAND U12451 ( .A(n11370), .B(n11369), .Z(n11376) );
  NAND U12452 ( .A(b[0]), .B(a[898]), .Z(n11375) );
  NAND U12453 ( .A(a[897]), .B(b[1]), .Z(n11374) );
  XNOR U12454 ( .A(n11375), .B(n11374), .Z(n11377) );
  XNOR U12455 ( .A(n11376), .B(n11377), .Z(n11381) );
  XOR U12456 ( .A(n11380), .B(sreg[1920]), .Z(n11373) );
  XNOR U12457 ( .A(n11381), .B(n11373), .Z(c[1920]) );
  NAND U12458 ( .A(n11375), .B(n11374), .Z(n11379) );
  NANDN U12459 ( .A(n11377), .B(n11376), .Z(n11378) );
  NAND U12460 ( .A(n11379), .B(n11378), .Z(n11385) );
  NAND U12461 ( .A(b[0]), .B(a[899]), .Z(n11384) );
  NAND U12462 ( .A(a[898]), .B(b[1]), .Z(n11383) );
  XNOR U12463 ( .A(n11384), .B(n11383), .Z(n11386) );
  XNOR U12464 ( .A(n11385), .B(n11386), .Z(n11390) );
  XOR U12465 ( .A(n11389), .B(sreg[1921]), .Z(n11382) );
  XNOR U12466 ( .A(n11390), .B(n11382), .Z(c[1921]) );
  NAND U12467 ( .A(n11384), .B(n11383), .Z(n11388) );
  NANDN U12468 ( .A(n11386), .B(n11385), .Z(n11387) );
  NAND U12469 ( .A(n11388), .B(n11387), .Z(n11395) );
  ANDN U12470 ( .B(a[900]), .A(n3979), .Z(n11393) );
  AND U12471 ( .A(b[1]), .B(a[899]), .Z(n11392) );
  XOR U12472 ( .A(n11393), .B(n11392), .Z(n11394) );
  XNOR U12473 ( .A(n11395), .B(n11394), .Z(n11397) );
  XOR U12474 ( .A(sreg[1922]), .B(n11396), .Z(n11391) );
  XNOR U12475 ( .A(n11397), .B(n11391), .Z(c[1922]) );
  NAND U12476 ( .A(b[0]), .B(a[901]), .Z(n11400) );
  NAND U12477 ( .A(a[900]), .B(b[1]), .Z(n11399) );
  XNOR U12478 ( .A(n11400), .B(n11399), .Z(n11402) );
  XNOR U12479 ( .A(n11401), .B(n11402), .Z(n11406) );
  XOR U12480 ( .A(n11405), .B(sreg[1923]), .Z(n11398) );
  XNOR U12481 ( .A(n11406), .B(n11398), .Z(c[1923]) );
  NAND U12482 ( .A(n11400), .B(n11399), .Z(n11404) );
  NANDN U12483 ( .A(n11402), .B(n11401), .Z(n11403) );
  NAND U12484 ( .A(n11404), .B(n11403), .Z(n11410) );
  NAND U12485 ( .A(b[0]), .B(a[902]), .Z(n11409) );
  NAND U12486 ( .A(a[901]), .B(b[1]), .Z(n11408) );
  XNOR U12487 ( .A(n11409), .B(n11408), .Z(n11411) );
  XNOR U12488 ( .A(n11410), .B(n11411), .Z(n11415) );
  XOR U12489 ( .A(n11414), .B(sreg[1924]), .Z(n11407) );
  XNOR U12490 ( .A(n11415), .B(n11407), .Z(c[1924]) );
  NAND U12491 ( .A(n11409), .B(n11408), .Z(n11413) );
  NANDN U12492 ( .A(n11411), .B(n11410), .Z(n11412) );
  NAND U12493 ( .A(n11413), .B(n11412), .Z(n11420) );
  ANDN U12494 ( .B(a[903]), .A(n3979), .Z(n11418) );
  AND U12495 ( .A(b[1]), .B(a[902]), .Z(n11417) );
  XOR U12496 ( .A(n11418), .B(n11417), .Z(n11419) );
  XNOR U12497 ( .A(n11420), .B(n11419), .Z(n11422) );
  XOR U12498 ( .A(sreg[1925]), .B(n11421), .Z(n11416) );
  XNOR U12499 ( .A(n11422), .B(n11416), .Z(c[1925]) );
  ANDN U12500 ( .B(a[904]), .A(n3979), .Z(n11425) );
  AND U12501 ( .A(b[1]), .B(a[903]), .Z(n11424) );
  XOR U12502 ( .A(n11425), .B(n11424), .Z(n11426) );
  XNOR U12503 ( .A(n11427), .B(n11426), .Z(n11429) );
  XNOR U12504 ( .A(sreg[1926]), .B(n11428), .Z(n11423) );
  XNOR U12505 ( .A(n11429), .B(n11423), .Z(c[1926]) );
  NAND U12506 ( .A(b[0]), .B(a[905]), .Z(n11432) );
  NAND U12507 ( .A(a[904]), .B(b[1]), .Z(n11431) );
  XNOR U12508 ( .A(n11432), .B(n11431), .Z(n11434) );
  XNOR U12509 ( .A(n11433), .B(n11434), .Z(n11438) );
  XOR U12510 ( .A(n11437), .B(sreg[1927]), .Z(n11430) );
  XNOR U12511 ( .A(n11438), .B(n11430), .Z(c[1927]) );
  NAND U12512 ( .A(n11432), .B(n11431), .Z(n11436) );
  NANDN U12513 ( .A(n11434), .B(n11433), .Z(n11435) );
  NAND U12514 ( .A(n11436), .B(n11435), .Z(n11442) );
  NAND U12515 ( .A(b[0]), .B(a[906]), .Z(n11441) );
  NAND U12516 ( .A(a[905]), .B(b[1]), .Z(n11440) );
  XNOR U12517 ( .A(n11441), .B(n11440), .Z(n11443) );
  XNOR U12518 ( .A(n11442), .B(n11443), .Z(n11447) );
  XOR U12519 ( .A(n11446), .B(sreg[1928]), .Z(n11439) );
  XNOR U12520 ( .A(n11447), .B(n11439), .Z(c[1928]) );
  NAND U12521 ( .A(n11441), .B(n11440), .Z(n11445) );
  NANDN U12522 ( .A(n11443), .B(n11442), .Z(n11444) );
  NAND U12523 ( .A(n11445), .B(n11444), .Z(n11451) );
  NAND U12524 ( .A(b[0]), .B(a[907]), .Z(n11450) );
  NAND U12525 ( .A(a[906]), .B(b[1]), .Z(n11449) );
  XNOR U12526 ( .A(n11450), .B(n11449), .Z(n11452) );
  XNOR U12527 ( .A(n11451), .B(n11452), .Z(n11456) );
  XOR U12528 ( .A(n11455), .B(sreg[1929]), .Z(n11448) );
  XNOR U12529 ( .A(n11456), .B(n11448), .Z(c[1929]) );
  NAND U12530 ( .A(n11450), .B(n11449), .Z(n11454) );
  NANDN U12531 ( .A(n11452), .B(n11451), .Z(n11453) );
  NAND U12532 ( .A(n11454), .B(n11453), .Z(n11461) );
  ANDN U12533 ( .B(a[908]), .A(n3980), .Z(n11459) );
  AND U12534 ( .A(b[1]), .B(a[907]), .Z(n11458) );
  XOR U12535 ( .A(n11459), .B(n11458), .Z(n11460) );
  XNOR U12536 ( .A(n11461), .B(n11460), .Z(n11466) );
  XOR U12537 ( .A(sreg[1930]), .B(n11465), .Z(n11457) );
  XNOR U12538 ( .A(n11466), .B(n11457), .Z(c[1930]) );
  OR U12539 ( .A(n11459), .B(n11458), .Z(n11464) );
  IV U12540 ( .A(n11460), .Z(n11462) );
  NANDN U12541 ( .A(n11462), .B(n11461), .Z(n11463) );
  NAND U12542 ( .A(n11464), .B(n11463), .Z(n11470) );
  NAND U12543 ( .A(b[0]), .B(a[909]), .Z(n11469) );
  NAND U12544 ( .A(a[908]), .B(b[1]), .Z(n11468) );
  XNOR U12545 ( .A(n11469), .B(n11468), .Z(n11471) );
  XNOR U12546 ( .A(n11470), .B(n11471), .Z(n11475) );
  XOR U12547 ( .A(n11474), .B(sreg[1931]), .Z(n11467) );
  XNOR U12548 ( .A(n11475), .B(n11467), .Z(c[1931]) );
  NAND U12549 ( .A(n11469), .B(n11468), .Z(n11473) );
  NANDN U12550 ( .A(n11471), .B(n11470), .Z(n11472) );
  NAND U12551 ( .A(n11473), .B(n11472), .Z(n11480) );
  ANDN U12552 ( .B(a[910]), .A(n3980), .Z(n11478) );
  AND U12553 ( .A(b[1]), .B(a[909]), .Z(n11477) );
  XOR U12554 ( .A(n11478), .B(n11477), .Z(n11479) );
  XNOR U12555 ( .A(n11480), .B(n11479), .Z(n11482) );
  XOR U12556 ( .A(sreg[1932]), .B(n11481), .Z(n11476) );
  XNOR U12557 ( .A(n11482), .B(n11476), .Z(c[1932]) );
  NAND U12558 ( .A(b[0]), .B(a[911]), .Z(n11485) );
  NAND U12559 ( .A(a[910]), .B(b[1]), .Z(n11484) );
  XNOR U12560 ( .A(n11485), .B(n11484), .Z(n11487) );
  XNOR U12561 ( .A(n11486), .B(n11487), .Z(n11491) );
  XOR U12562 ( .A(n11490), .B(sreg[1933]), .Z(n11483) );
  XNOR U12563 ( .A(n11491), .B(n11483), .Z(c[1933]) );
  NAND U12564 ( .A(n11485), .B(n11484), .Z(n11489) );
  NANDN U12565 ( .A(n11487), .B(n11486), .Z(n11488) );
  NAND U12566 ( .A(n11489), .B(n11488), .Z(n11495) );
  NAND U12567 ( .A(b[0]), .B(a[912]), .Z(n11494) );
  NAND U12568 ( .A(a[911]), .B(b[1]), .Z(n11493) );
  XNOR U12569 ( .A(n11494), .B(n11493), .Z(n11496) );
  XNOR U12570 ( .A(n11495), .B(n11496), .Z(n11500) );
  XOR U12571 ( .A(n11499), .B(sreg[1934]), .Z(n11492) );
  XNOR U12572 ( .A(n11500), .B(n11492), .Z(c[1934]) );
  NAND U12573 ( .A(n11494), .B(n11493), .Z(n11498) );
  NANDN U12574 ( .A(n11496), .B(n11495), .Z(n11497) );
  NAND U12575 ( .A(n11498), .B(n11497), .Z(n11504) );
  NAND U12576 ( .A(b[0]), .B(a[913]), .Z(n11503) );
  NAND U12577 ( .A(a[912]), .B(b[1]), .Z(n11502) );
  XNOR U12578 ( .A(n11503), .B(n11502), .Z(n11505) );
  XNOR U12579 ( .A(n11504), .B(n11505), .Z(n11509) );
  XOR U12580 ( .A(n11508), .B(sreg[1935]), .Z(n11501) );
  XNOR U12581 ( .A(n11509), .B(n11501), .Z(c[1935]) );
  NAND U12582 ( .A(n11503), .B(n11502), .Z(n11507) );
  NANDN U12583 ( .A(n11505), .B(n11504), .Z(n11506) );
  NAND U12584 ( .A(n11507), .B(n11506), .Z(n11514) );
  ANDN U12585 ( .B(a[914]), .A(n3980), .Z(n11512) );
  AND U12586 ( .A(b[1]), .B(a[913]), .Z(n11511) );
  XOR U12587 ( .A(n11512), .B(n11511), .Z(n11513) );
  XNOR U12588 ( .A(n11514), .B(n11513), .Z(n11516) );
  XOR U12589 ( .A(sreg[1936]), .B(n11515), .Z(n11510) );
  XNOR U12590 ( .A(n11516), .B(n11510), .Z(c[1936]) );
  NAND U12591 ( .A(b[0]), .B(a[915]), .Z(n11519) );
  NAND U12592 ( .A(a[914]), .B(b[1]), .Z(n11518) );
  XNOR U12593 ( .A(n11519), .B(n11518), .Z(n11521) );
  XNOR U12594 ( .A(n11520), .B(n11521), .Z(n11525) );
  XOR U12595 ( .A(n11524), .B(sreg[1937]), .Z(n11517) );
  XNOR U12596 ( .A(n11525), .B(n11517), .Z(c[1937]) );
  NAND U12597 ( .A(n11519), .B(n11518), .Z(n11523) );
  NANDN U12598 ( .A(n11521), .B(n11520), .Z(n11522) );
  NAND U12599 ( .A(n11523), .B(n11522), .Z(n11530) );
  ANDN U12600 ( .B(a[916]), .A(n3980), .Z(n11528) );
  AND U12601 ( .A(b[1]), .B(a[915]), .Z(n11527) );
  XOR U12602 ( .A(n11528), .B(n11527), .Z(n11529) );
  XNOR U12603 ( .A(n11530), .B(n11529), .Z(n11532) );
  XOR U12604 ( .A(sreg[1938]), .B(n11531), .Z(n11526) );
  XNOR U12605 ( .A(n11532), .B(n11526), .Z(c[1938]) );
  ANDN U12606 ( .B(a[917]), .A(n3980), .Z(n11535) );
  AND U12607 ( .A(b[1]), .B(a[916]), .Z(n11534) );
  XOR U12608 ( .A(n11535), .B(n11534), .Z(n11536) );
  XNOR U12609 ( .A(n11537), .B(n11536), .Z(n11539) );
  XNOR U12610 ( .A(sreg[1939]), .B(n11538), .Z(n11533) );
  XNOR U12611 ( .A(n11539), .B(n11533), .Z(c[1939]) );
  ANDN U12612 ( .B(a[918]), .A(n3980), .Z(n11542) );
  AND U12613 ( .A(b[1]), .B(a[917]), .Z(n11541) );
  XOR U12614 ( .A(n11542), .B(n11541), .Z(n11543) );
  XNOR U12615 ( .A(n11544), .B(n11543), .Z(n11546) );
  XNOR U12616 ( .A(sreg[1940]), .B(n11545), .Z(n11540) );
  XNOR U12617 ( .A(n11546), .B(n11540), .Z(c[1940]) );
  NAND U12618 ( .A(b[0]), .B(a[919]), .Z(n11549) );
  NAND U12619 ( .A(a[918]), .B(b[1]), .Z(n11548) );
  XNOR U12620 ( .A(n11549), .B(n11548), .Z(n11551) );
  XNOR U12621 ( .A(n11550), .B(n11551), .Z(n11555) );
  XOR U12622 ( .A(n11554), .B(sreg[1941]), .Z(n11547) );
  XNOR U12623 ( .A(n11555), .B(n11547), .Z(c[1941]) );
  NAND U12624 ( .A(n11549), .B(n11548), .Z(n11553) );
  NANDN U12625 ( .A(n11551), .B(n11550), .Z(n11552) );
  NAND U12626 ( .A(n11553), .B(n11552), .Z(n11559) );
  NAND U12627 ( .A(b[0]), .B(a[920]), .Z(n11558) );
  NAND U12628 ( .A(a[919]), .B(b[1]), .Z(n11557) );
  XNOR U12629 ( .A(n11558), .B(n11557), .Z(n11560) );
  XNOR U12630 ( .A(n11559), .B(n11560), .Z(n11564) );
  XOR U12631 ( .A(n11563), .B(sreg[1942]), .Z(n11556) );
  XNOR U12632 ( .A(n11564), .B(n11556), .Z(c[1942]) );
  NAND U12633 ( .A(n11558), .B(n11557), .Z(n11562) );
  NANDN U12634 ( .A(n11560), .B(n11559), .Z(n11561) );
  NAND U12635 ( .A(n11562), .B(n11561), .Z(n11568) );
  NAND U12636 ( .A(b[0]), .B(a[921]), .Z(n11567) );
  NAND U12637 ( .A(a[920]), .B(b[1]), .Z(n11566) );
  XNOR U12638 ( .A(n11567), .B(n11566), .Z(n11569) );
  XNOR U12639 ( .A(n11568), .B(n11569), .Z(n11573) );
  XOR U12640 ( .A(n11572), .B(sreg[1943]), .Z(n11565) );
  XNOR U12641 ( .A(n11573), .B(n11565), .Z(c[1943]) );
  NAND U12642 ( .A(n11567), .B(n11566), .Z(n11571) );
  NANDN U12643 ( .A(n11569), .B(n11568), .Z(n11570) );
  NAND U12644 ( .A(n11571), .B(n11570), .Z(n11578) );
  ANDN U12645 ( .B(a[922]), .A(n3980), .Z(n11576) );
  AND U12646 ( .A(b[1]), .B(a[921]), .Z(n11575) );
  XOR U12647 ( .A(n11576), .B(n11575), .Z(n11577) );
  XNOR U12648 ( .A(n11578), .B(n11577), .Z(n11580) );
  XOR U12649 ( .A(sreg[1944]), .B(n11579), .Z(n11574) );
  XNOR U12650 ( .A(n11580), .B(n11574), .Z(c[1944]) );
  NAND U12651 ( .A(b[0]), .B(a[923]), .Z(n11583) );
  NAND U12652 ( .A(a[922]), .B(b[1]), .Z(n11582) );
  XNOR U12653 ( .A(n11583), .B(n11582), .Z(n11585) );
  XNOR U12654 ( .A(n11584), .B(n11585), .Z(n11589) );
  XOR U12655 ( .A(n11588), .B(sreg[1945]), .Z(n11581) );
  XNOR U12656 ( .A(n11589), .B(n11581), .Z(c[1945]) );
  NAND U12657 ( .A(n11583), .B(n11582), .Z(n11587) );
  NANDN U12658 ( .A(n11585), .B(n11584), .Z(n11586) );
  NAND U12659 ( .A(n11587), .B(n11586), .Z(n11594) );
  ANDN U12660 ( .B(a[924]), .A(n3981), .Z(n11592) );
  AND U12661 ( .A(b[1]), .B(a[923]), .Z(n11591) );
  XOR U12662 ( .A(n11592), .B(n11591), .Z(n11593) );
  XNOR U12663 ( .A(n11594), .B(n11593), .Z(n11599) );
  XOR U12664 ( .A(sreg[1946]), .B(n11598), .Z(n11590) );
  XNOR U12665 ( .A(n11599), .B(n11590), .Z(c[1946]) );
  OR U12666 ( .A(n11592), .B(n11591), .Z(n11597) );
  IV U12667 ( .A(n11593), .Z(n11595) );
  NANDN U12668 ( .A(n11595), .B(n11594), .Z(n11596) );
  NAND U12669 ( .A(n11597), .B(n11596), .Z(n11603) );
  NAND U12670 ( .A(b[0]), .B(a[925]), .Z(n11602) );
  NAND U12671 ( .A(a[924]), .B(b[1]), .Z(n11601) );
  XNOR U12672 ( .A(n11602), .B(n11601), .Z(n11604) );
  XNOR U12673 ( .A(n11603), .B(n11604), .Z(n11608) );
  XOR U12674 ( .A(n11607), .B(sreg[1947]), .Z(n11600) );
  XNOR U12675 ( .A(n11608), .B(n11600), .Z(c[1947]) );
  NAND U12676 ( .A(n11602), .B(n11601), .Z(n11606) );
  NANDN U12677 ( .A(n11604), .B(n11603), .Z(n11605) );
  NAND U12678 ( .A(n11606), .B(n11605), .Z(n11613) );
  ANDN U12679 ( .B(a[926]), .A(n3981), .Z(n11611) );
  AND U12680 ( .A(b[1]), .B(a[925]), .Z(n11610) );
  XOR U12681 ( .A(n11611), .B(n11610), .Z(n11612) );
  XNOR U12682 ( .A(n11613), .B(n11612), .Z(n11615) );
  XOR U12683 ( .A(sreg[1948]), .B(n11614), .Z(n11609) );
  XNOR U12684 ( .A(n11615), .B(n11609), .Z(c[1948]) );
  NAND U12685 ( .A(b[0]), .B(a[927]), .Z(n11618) );
  NAND U12686 ( .A(a[926]), .B(b[1]), .Z(n11617) );
  XNOR U12687 ( .A(n11618), .B(n11617), .Z(n11620) );
  XNOR U12688 ( .A(n11619), .B(n11620), .Z(n11624) );
  XOR U12689 ( .A(n11623), .B(sreg[1949]), .Z(n11616) );
  XNOR U12690 ( .A(n11624), .B(n11616), .Z(c[1949]) );
  NAND U12691 ( .A(n11618), .B(n11617), .Z(n11622) );
  NANDN U12692 ( .A(n11620), .B(n11619), .Z(n11621) );
  NAND U12693 ( .A(n11622), .B(n11621), .Z(n11629) );
  ANDN U12694 ( .B(a[928]), .A(n3981), .Z(n11627) );
  AND U12695 ( .A(b[1]), .B(a[927]), .Z(n11626) );
  XOR U12696 ( .A(n11627), .B(n11626), .Z(n11628) );
  XNOR U12697 ( .A(n11629), .B(n11628), .Z(n11631) );
  XOR U12698 ( .A(sreg[1950]), .B(n11630), .Z(n11625) );
  XNOR U12699 ( .A(n11631), .B(n11625), .Z(c[1950]) );
  NAND U12700 ( .A(b[0]), .B(a[929]), .Z(n11634) );
  NAND U12701 ( .A(a[928]), .B(b[1]), .Z(n11633) );
  XNOR U12702 ( .A(n11634), .B(n11633), .Z(n11636) );
  XNOR U12703 ( .A(n11635), .B(n11636), .Z(n11640) );
  XOR U12704 ( .A(n11639), .B(sreg[1951]), .Z(n11632) );
  XNOR U12705 ( .A(n11640), .B(n11632), .Z(c[1951]) );
  NAND U12706 ( .A(n11634), .B(n11633), .Z(n11638) );
  NANDN U12707 ( .A(n11636), .B(n11635), .Z(n11637) );
  NAND U12708 ( .A(n11638), .B(n11637), .Z(n11645) );
  ANDN U12709 ( .B(a[930]), .A(n3981), .Z(n11643) );
  AND U12710 ( .A(b[1]), .B(a[929]), .Z(n11642) );
  XOR U12711 ( .A(n11643), .B(n11642), .Z(n11644) );
  XNOR U12712 ( .A(n11645), .B(n11644), .Z(n11647) );
  XOR U12713 ( .A(sreg[1952]), .B(n11646), .Z(n11641) );
  XNOR U12714 ( .A(n11647), .B(n11641), .Z(c[1952]) );
  NAND U12715 ( .A(b[0]), .B(a[931]), .Z(n11650) );
  NAND U12716 ( .A(a[930]), .B(b[1]), .Z(n11649) );
  XNOR U12717 ( .A(n11650), .B(n11649), .Z(n11652) );
  XNOR U12718 ( .A(n11651), .B(n11652), .Z(n11656) );
  XOR U12719 ( .A(n11655), .B(sreg[1953]), .Z(n11648) );
  XNOR U12720 ( .A(n11656), .B(n11648), .Z(c[1953]) );
  NAND U12721 ( .A(n11650), .B(n11649), .Z(n11654) );
  NANDN U12722 ( .A(n11652), .B(n11651), .Z(n11653) );
  NAND U12723 ( .A(n11654), .B(n11653), .Z(n11660) );
  NAND U12724 ( .A(b[0]), .B(a[932]), .Z(n11659) );
  NAND U12725 ( .A(a[931]), .B(b[1]), .Z(n11658) );
  XNOR U12726 ( .A(n11659), .B(n11658), .Z(n11661) );
  XNOR U12727 ( .A(n11660), .B(n11661), .Z(n11665) );
  XOR U12728 ( .A(n11664), .B(sreg[1954]), .Z(n11657) );
  XNOR U12729 ( .A(n11665), .B(n11657), .Z(c[1954]) );
  NAND U12730 ( .A(n11659), .B(n11658), .Z(n11663) );
  NANDN U12731 ( .A(n11661), .B(n11660), .Z(n11662) );
  NAND U12732 ( .A(n11663), .B(n11662), .Z(n11669) );
  NAND U12733 ( .A(b[0]), .B(a[933]), .Z(n11668) );
  NAND U12734 ( .A(a[932]), .B(b[1]), .Z(n11667) );
  XNOR U12735 ( .A(n11668), .B(n11667), .Z(n11670) );
  XNOR U12736 ( .A(n11669), .B(n11670), .Z(n11674) );
  XOR U12737 ( .A(n11673), .B(sreg[1955]), .Z(n11666) );
  XNOR U12738 ( .A(n11674), .B(n11666), .Z(c[1955]) );
  NAND U12739 ( .A(n11668), .B(n11667), .Z(n11672) );
  NANDN U12740 ( .A(n11670), .B(n11669), .Z(n11671) );
  NAND U12741 ( .A(n11672), .B(n11671), .Z(n11679) );
  ANDN U12742 ( .B(a[934]), .A(n3981), .Z(n11677) );
  AND U12743 ( .A(b[1]), .B(a[933]), .Z(n11676) );
  XOR U12744 ( .A(n11677), .B(n11676), .Z(n11678) );
  XNOR U12745 ( .A(n11679), .B(n11678), .Z(n11681) );
  XOR U12746 ( .A(sreg[1956]), .B(n11680), .Z(n11675) );
  XNOR U12747 ( .A(n11681), .B(n11675), .Z(c[1956]) );
  NAND U12748 ( .A(b[0]), .B(a[935]), .Z(n11684) );
  NAND U12749 ( .A(a[934]), .B(b[1]), .Z(n11683) );
  XNOR U12750 ( .A(n11684), .B(n11683), .Z(n11686) );
  XNOR U12751 ( .A(n11685), .B(n11686), .Z(n11690) );
  XOR U12752 ( .A(n11689), .B(sreg[1957]), .Z(n11682) );
  XNOR U12753 ( .A(n11690), .B(n11682), .Z(c[1957]) );
  NAND U12754 ( .A(n11684), .B(n11683), .Z(n11688) );
  NANDN U12755 ( .A(n11686), .B(n11685), .Z(n11687) );
  NAND U12756 ( .A(n11688), .B(n11687), .Z(n11695) );
  ANDN U12757 ( .B(a[936]), .A(n3981), .Z(n11693) );
  AND U12758 ( .A(b[1]), .B(a[935]), .Z(n11692) );
  XOR U12759 ( .A(n11693), .B(n11692), .Z(n11694) );
  XNOR U12760 ( .A(n11695), .B(n11694), .Z(n11697) );
  XOR U12761 ( .A(sreg[1958]), .B(n11696), .Z(n11691) );
  XNOR U12762 ( .A(n11697), .B(n11691), .Z(c[1958]) );
  ANDN U12763 ( .B(a[937]), .A(n3981), .Z(n11700) );
  AND U12764 ( .A(b[1]), .B(a[936]), .Z(n11699) );
  XOR U12765 ( .A(n11700), .B(n11699), .Z(n11701) );
  XNOR U12766 ( .A(n11702), .B(n11701), .Z(n11704) );
  XNOR U12767 ( .A(sreg[1959]), .B(n11703), .Z(n11698) );
  XNOR U12768 ( .A(n11704), .B(n11698), .Z(c[1959]) );
  NAND U12769 ( .A(b[0]), .B(a[938]), .Z(n11707) );
  NAND U12770 ( .A(a[937]), .B(b[1]), .Z(n11706) );
  XNOR U12771 ( .A(n11707), .B(n11706), .Z(n11709) );
  XNOR U12772 ( .A(n11708), .B(n11709), .Z(n11713) );
  XOR U12773 ( .A(n11712), .B(sreg[1960]), .Z(n11705) );
  XNOR U12774 ( .A(n11713), .B(n11705), .Z(c[1960]) );
  NAND U12775 ( .A(n11707), .B(n11706), .Z(n11711) );
  NANDN U12776 ( .A(n11709), .B(n11708), .Z(n11710) );
  NAND U12777 ( .A(n11711), .B(n11710), .Z(n11717) );
  NAND U12778 ( .A(b[0]), .B(a[939]), .Z(n11716) );
  NAND U12779 ( .A(a[938]), .B(b[1]), .Z(n11715) );
  XNOR U12780 ( .A(n11716), .B(n11715), .Z(n11718) );
  XNOR U12781 ( .A(n11717), .B(n11718), .Z(n11722) );
  XOR U12782 ( .A(n11721), .B(sreg[1961]), .Z(n11714) );
  XNOR U12783 ( .A(n11722), .B(n11714), .Z(c[1961]) );
  NAND U12784 ( .A(n11716), .B(n11715), .Z(n11720) );
  NANDN U12785 ( .A(n11718), .B(n11717), .Z(n11719) );
  NAND U12786 ( .A(n11720), .B(n11719), .Z(n11727) );
  ANDN U12787 ( .B(a[940]), .A(n3982), .Z(n11725) );
  AND U12788 ( .A(b[1]), .B(a[939]), .Z(n11724) );
  XOR U12789 ( .A(n11725), .B(n11724), .Z(n11726) );
  XNOR U12790 ( .A(n11727), .B(n11726), .Z(n11732) );
  XOR U12791 ( .A(sreg[1962]), .B(n11731), .Z(n11723) );
  XNOR U12792 ( .A(n11732), .B(n11723), .Z(c[1962]) );
  OR U12793 ( .A(n11725), .B(n11724), .Z(n11730) );
  IV U12794 ( .A(n11726), .Z(n11728) );
  NANDN U12795 ( .A(n11728), .B(n11727), .Z(n11729) );
  NAND U12796 ( .A(n11730), .B(n11729), .Z(n11736) );
  NAND U12797 ( .A(b[0]), .B(a[941]), .Z(n11735) );
  NAND U12798 ( .A(a[940]), .B(b[1]), .Z(n11734) );
  XNOR U12799 ( .A(n11735), .B(n11734), .Z(n11737) );
  XNOR U12800 ( .A(n11736), .B(n11737), .Z(n11741) );
  XOR U12801 ( .A(n11740), .B(sreg[1963]), .Z(n11733) );
  XNOR U12802 ( .A(n11741), .B(n11733), .Z(c[1963]) );
  NAND U12803 ( .A(n11735), .B(n11734), .Z(n11739) );
  NANDN U12804 ( .A(n11737), .B(n11736), .Z(n11738) );
  NAND U12805 ( .A(n11739), .B(n11738), .Z(n11746) );
  ANDN U12806 ( .B(a[942]), .A(n3982), .Z(n11744) );
  AND U12807 ( .A(b[1]), .B(a[941]), .Z(n11743) );
  XOR U12808 ( .A(n11744), .B(n11743), .Z(n11745) );
  XNOR U12809 ( .A(n11746), .B(n11745), .Z(n11748) );
  XOR U12810 ( .A(sreg[1964]), .B(n11747), .Z(n11742) );
  XNOR U12811 ( .A(n11748), .B(n11742), .Z(c[1964]) );
  NAND U12812 ( .A(b[0]), .B(a[943]), .Z(n11751) );
  NAND U12813 ( .A(a[942]), .B(b[1]), .Z(n11750) );
  XNOR U12814 ( .A(n11751), .B(n11750), .Z(n11753) );
  XNOR U12815 ( .A(n11752), .B(n11753), .Z(n11757) );
  XOR U12816 ( .A(n11756), .B(sreg[1965]), .Z(n11749) );
  XNOR U12817 ( .A(n11757), .B(n11749), .Z(c[1965]) );
  NAND U12818 ( .A(n11751), .B(n11750), .Z(n11755) );
  NANDN U12819 ( .A(n11753), .B(n11752), .Z(n11754) );
  NAND U12820 ( .A(n11755), .B(n11754), .Z(n11762) );
  ANDN U12821 ( .B(a[944]), .A(n3982), .Z(n11760) );
  AND U12822 ( .A(b[1]), .B(a[943]), .Z(n11759) );
  XOR U12823 ( .A(n11760), .B(n11759), .Z(n11761) );
  XNOR U12824 ( .A(n11762), .B(n11761), .Z(n11764) );
  XOR U12825 ( .A(sreg[1966]), .B(n11763), .Z(n11758) );
  XNOR U12826 ( .A(n11764), .B(n11758), .Z(c[1966]) );
  NAND U12827 ( .A(b[0]), .B(a[945]), .Z(n11767) );
  NAND U12828 ( .A(a[944]), .B(b[1]), .Z(n11766) );
  XNOR U12829 ( .A(n11767), .B(n11766), .Z(n11769) );
  XNOR U12830 ( .A(n11768), .B(n11769), .Z(n11773) );
  XOR U12831 ( .A(n11772), .B(sreg[1967]), .Z(n11765) );
  XNOR U12832 ( .A(n11773), .B(n11765), .Z(c[1967]) );
  NAND U12833 ( .A(n11767), .B(n11766), .Z(n11771) );
  NANDN U12834 ( .A(n11769), .B(n11768), .Z(n11770) );
  NAND U12835 ( .A(n11771), .B(n11770), .Z(n11777) );
  NAND U12836 ( .A(b[0]), .B(a[946]), .Z(n11776) );
  NAND U12837 ( .A(a[945]), .B(b[1]), .Z(n11775) );
  XNOR U12838 ( .A(n11776), .B(n11775), .Z(n11778) );
  XNOR U12839 ( .A(n11777), .B(n11778), .Z(n11782) );
  XOR U12840 ( .A(n11781), .B(sreg[1968]), .Z(n11774) );
  XNOR U12841 ( .A(n11782), .B(n11774), .Z(c[1968]) );
  NAND U12842 ( .A(n11776), .B(n11775), .Z(n11780) );
  NANDN U12843 ( .A(n11778), .B(n11777), .Z(n11779) );
  NAND U12844 ( .A(n11780), .B(n11779), .Z(n11786) );
  NAND U12845 ( .A(b[0]), .B(a[947]), .Z(n11785) );
  NAND U12846 ( .A(a[946]), .B(b[1]), .Z(n11784) );
  XNOR U12847 ( .A(n11785), .B(n11784), .Z(n11787) );
  XNOR U12848 ( .A(n11786), .B(n11787), .Z(n11791) );
  XOR U12849 ( .A(n11790), .B(sreg[1969]), .Z(n11783) );
  XNOR U12850 ( .A(n11791), .B(n11783), .Z(c[1969]) );
  NAND U12851 ( .A(n11785), .B(n11784), .Z(n11789) );
  NANDN U12852 ( .A(n11787), .B(n11786), .Z(n11788) );
  NAND U12853 ( .A(n11789), .B(n11788), .Z(n11795) );
  NAND U12854 ( .A(b[0]), .B(a[948]), .Z(n11794) );
  NAND U12855 ( .A(a[947]), .B(b[1]), .Z(n11793) );
  XNOR U12856 ( .A(n11794), .B(n11793), .Z(n11796) );
  XNOR U12857 ( .A(n11795), .B(n11796), .Z(n11800) );
  XOR U12858 ( .A(n11799), .B(sreg[1970]), .Z(n11792) );
  XNOR U12859 ( .A(n11800), .B(n11792), .Z(c[1970]) );
  NAND U12860 ( .A(n11794), .B(n11793), .Z(n11798) );
  NANDN U12861 ( .A(n11796), .B(n11795), .Z(n11797) );
  NAND U12862 ( .A(n11798), .B(n11797), .Z(n11804) );
  NAND U12863 ( .A(b[0]), .B(a[949]), .Z(n11803) );
  NAND U12864 ( .A(a[948]), .B(b[1]), .Z(n11802) );
  XNOR U12865 ( .A(n11803), .B(n11802), .Z(n11805) );
  XNOR U12866 ( .A(n11804), .B(n11805), .Z(n11809) );
  XOR U12867 ( .A(n11808), .B(sreg[1971]), .Z(n11801) );
  XNOR U12868 ( .A(n11809), .B(n11801), .Z(c[1971]) );
  NAND U12869 ( .A(n11803), .B(n11802), .Z(n11807) );
  NANDN U12870 ( .A(n11805), .B(n11804), .Z(n11806) );
  NAND U12871 ( .A(n11807), .B(n11806), .Z(n11813) );
  NAND U12872 ( .A(b[0]), .B(a[950]), .Z(n11812) );
  NAND U12873 ( .A(a[949]), .B(b[1]), .Z(n11811) );
  XNOR U12874 ( .A(n11812), .B(n11811), .Z(n11814) );
  XNOR U12875 ( .A(n11813), .B(n11814), .Z(n11818) );
  XOR U12876 ( .A(n11817), .B(sreg[1972]), .Z(n11810) );
  XNOR U12877 ( .A(n11818), .B(n11810), .Z(c[1972]) );
  NAND U12878 ( .A(n11812), .B(n11811), .Z(n11816) );
  NANDN U12879 ( .A(n11814), .B(n11813), .Z(n11815) );
  NAND U12880 ( .A(n11816), .B(n11815), .Z(n11822) );
  NAND U12881 ( .A(b[0]), .B(a[951]), .Z(n11821) );
  NAND U12882 ( .A(a[950]), .B(b[1]), .Z(n11820) );
  XNOR U12883 ( .A(n11821), .B(n11820), .Z(n11823) );
  XNOR U12884 ( .A(n11822), .B(n11823), .Z(n11827) );
  XOR U12885 ( .A(n11826), .B(sreg[1973]), .Z(n11819) );
  XNOR U12886 ( .A(n11827), .B(n11819), .Z(c[1973]) );
  NAND U12887 ( .A(n11821), .B(n11820), .Z(n11825) );
  NANDN U12888 ( .A(n11823), .B(n11822), .Z(n11824) );
  NAND U12889 ( .A(n11825), .B(n11824), .Z(n11832) );
  ANDN U12890 ( .B(a[952]), .A(n3982), .Z(n11830) );
  AND U12891 ( .A(b[1]), .B(a[951]), .Z(n11829) );
  XOR U12892 ( .A(n11830), .B(n11829), .Z(n11831) );
  XNOR U12893 ( .A(n11832), .B(n11831), .Z(n11834) );
  XOR U12894 ( .A(sreg[1974]), .B(n11833), .Z(n11828) );
  XNOR U12895 ( .A(n11834), .B(n11828), .Z(c[1974]) );
  NAND U12896 ( .A(b[0]), .B(a[953]), .Z(n11837) );
  NAND U12897 ( .A(a[952]), .B(b[1]), .Z(n11836) );
  XNOR U12898 ( .A(n11837), .B(n11836), .Z(n11839) );
  XNOR U12899 ( .A(n11838), .B(n11839), .Z(n11843) );
  XOR U12900 ( .A(n11842), .B(sreg[1975]), .Z(n11835) );
  XNOR U12901 ( .A(n11843), .B(n11835), .Z(c[1975]) );
  NAND U12902 ( .A(n11837), .B(n11836), .Z(n11841) );
  NANDN U12903 ( .A(n11839), .B(n11838), .Z(n11840) );
  NAND U12904 ( .A(n11841), .B(n11840), .Z(n11848) );
  ANDN U12905 ( .B(a[954]), .A(n3982), .Z(n11846) );
  AND U12906 ( .A(b[1]), .B(a[953]), .Z(n11845) );
  XOR U12907 ( .A(n11846), .B(n11845), .Z(n11847) );
  XNOR U12908 ( .A(n11848), .B(n11847), .Z(n11850) );
  XOR U12909 ( .A(sreg[1976]), .B(n11849), .Z(n11844) );
  XNOR U12910 ( .A(n11850), .B(n11844), .Z(c[1976]) );
  NAND U12911 ( .A(b[0]), .B(a[955]), .Z(n11853) );
  NAND U12912 ( .A(a[954]), .B(b[1]), .Z(n11852) );
  XNOR U12913 ( .A(n11853), .B(n11852), .Z(n11855) );
  XNOR U12914 ( .A(n11854), .B(n11855), .Z(n11859) );
  XOR U12915 ( .A(n11858), .B(sreg[1977]), .Z(n11851) );
  XNOR U12916 ( .A(n11859), .B(n11851), .Z(c[1977]) );
  NAND U12917 ( .A(n11853), .B(n11852), .Z(n11857) );
  NANDN U12918 ( .A(n11855), .B(n11854), .Z(n11856) );
  NAND U12919 ( .A(n11857), .B(n11856), .Z(n11864) );
  ANDN U12920 ( .B(a[956]), .A(n3982), .Z(n11862) );
  AND U12921 ( .A(b[1]), .B(a[955]), .Z(n11861) );
  XOR U12922 ( .A(n11862), .B(n11861), .Z(n11863) );
  XNOR U12923 ( .A(n11864), .B(n11863), .Z(n11866) );
  XOR U12924 ( .A(sreg[1978]), .B(n11865), .Z(n11860) );
  XNOR U12925 ( .A(n11866), .B(n11860), .Z(c[1978]) );
  NAND U12926 ( .A(b[0]), .B(a[957]), .Z(n11869) );
  NAND U12927 ( .A(a[956]), .B(b[1]), .Z(n11868) );
  XNOR U12928 ( .A(n11869), .B(n11868), .Z(n11871) );
  XNOR U12929 ( .A(n11870), .B(n11871), .Z(n11875) );
  XOR U12930 ( .A(n11874), .B(sreg[1979]), .Z(n11867) );
  XNOR U12931 ( .A(n11875), .B(n11867), .Z(c[1979]) );
  NAND U12932 ( .A(n11869), .B(n11868), .Z(n11873) );
  NANDN U12933 ( .A(n11871), .B(n11870), .Z(n11872) );
  NAND U12934 ( .A(n11873), .B(n11872), .Z(n11880) );
  ANDN U12935 ( .B(a[958]), .A(n3982), .Z(n11878) );
  AND U12936 ( .A(b[1]), .B(a[957]), .Z(n11877) );
  XOR U12937 ( .A(n11878), .B(n11877), .Z(n11879) );
  XNOR U12938 ( .A(n11880), .B(n11879), .Z(n11882) );
  XOR U12939 ( .A(sreg[1980]), .B(n11881), .Z(n11876) );
  XNOR U12940 ( .A(n11882), .B(n11876), .Z(c[1980]) );
  NAND U12941 ( .A(b[0]), .B(a[959]), .Z(n11885) );
  NAND U12942 ( .A(a[958]), .B(b[1]), .Z(n11884) );
  XNOR U12943 ( .A(n11885), .B(n11884), .Z(n11887) );
  XNOR U12944 ( .A(n11886), .B(n11887), .Z(n11891) );
  XOR U12945 ( .A(n11890), .B(sreg[1981]), .Z(n11883) );
  XNOR U12946 ( .A(n11891), .B(n11883), .Z(c[1981]) );
  NAND U12947 ( .A(n11885), .B(n11884), .Z(n11889) );
  NANDN U12948 ( .A(n11887), .B(n11886), .Z(n11888) );
  NAND U12949 ( .A(n11889), .B(n11888), .Z(n11896) );
  ANDN U12950 ( .B(a[960]), .A(n3983), .Z(n11894) );
  AND U12951 ( .A(b[1]), .B(a[959]), .Z(n11893) );
  XOR U12952 ( .A(n11894), .B(n11893), .Z(n11895) );
  XNOR U12953 ( .A(n11896), .B(n11895), .Z(n11901) );
  XOR U12954 ( .A(sreg[1982]), .B(n11900), .Z(n11892) );
  XNOR U12955 ( .A(n11901), .B(n11892), .Z(c[1982]) );
  OR U12956 ( .A(n11894), .B(n11893), .Z(n11899) );
  IV U12957 ( .A(n11895), .Z(n11897) );
  NANDN U12958 ( .A(n11897), .B(n11896), .Z(n11898) );
  NAND U12959 ( .A(n11899), .B(n11898), .Z(n11905) );
  NAND U12960 ( .A(b[0]), .B(a[961]), .Z(n11904) );
  NAND U12961 ( .A(a[960]), .B(b[1]), .Z(n11903) );
  XNOR U12962 ( .A(n11904), .B(n11903), .Z(n11906) );
  XNOR U12963 ( .A(n11905), .B(n11906), .Z(n11910) );
  XOR U12964 ( .A(n11909), .B(sreg[1983]), .Z(n11902) );
  XNOR U12965 ( .A(n11910), .B(n11902), .Z(c[1983]) );
  NAND U12966 ( .A(n11904), .B(n11903), .Z(n11908) );
  NANDN U12967 ( .A(n11906), .B(n11905), .Z(n11907) );
  NAND U12968 ( .A(n11908), .B(n11907), .Z(n11915) );
  ANDN U12969 ( .B(a[962]), .A(n3983), .Z(n11913) );
  AND U12970 ( .A(b[1]), .B(a[961]), .Z(n11912) );
  XOR U12971 ( .A(n11913), .B(n11912), .Z(n11914) );
  XNOR U12972 ( .A(n11915), .B(n11914), .Z(n11917) );
  XOR U12973 ( .A(sreg[1984]), .B(n11916), .Z(n11911) );
  XNOR U12974 ( .A(n11917), .B(n11911), .Z(c[1984]) );
  NAND U12975 ( .A(b[0]), .B(a[963]), .Z(n11920) );
  NAND U12976 ( .A(a[962]), .B(b[1]), .Z(n11919) );
  XNOR U12977 ( .A(n11920), .B(n11919), .Z(n11922) );
  XNOR U12978 ( .A(n11921), .B(n11922), .Z(n11926) );
  XOR U12979 ( .A(n11925), .B(sreg[1985]), .Z(n11918) );
  XNOR U12980 ( .A(n11926), .B(n11918), .Z(c[1985]) );
  NAND U12981 ( .A(n11920), .B(n11919), .Z(n11924) );
  NANDN U12982 ( .A(n11922), .B(n11921), .Z(n11923) );
  NAND U12983 ( .A(n11924), .B(n11923), .Z(n11931) );
  ANDN U12984 ( .B(a[964]), .A(n3983), .Z(n11929) );
  AND U12985 ( .A(b[1]), .B(a[963]), .Z(n11928) );
  XOR U12986 ( .A(n11929), .B(n11928), .Z(n11930) );
  XNOR U12987 ( .A(n11931), .B(n11930), .Z(n11933) );
  XOR U12988 ( .A(sreg[1986]), .B(n11932), .Z(n11927) );
  XNOR U12989 ( .A(n11933), .B(n11927), .Z(c[1986]) );
  NAND U12990 ( .A(b[0]), .B(a[965]), .Z(n11936) );
  NAND U12991 ( .A(a[964]), .B(b[1]), .Z(n11935) );
  XNOR U12992 ( .A(n11936), .B(n11935), .Z(n11938) );
  XNOR U12993 ( .A(n11937), .B(n11938), .Z(n11942) );
  XOR U12994 ( .A(n11941), .B(sreg[1987]), .Z(n11934) );
  XNOR U12995 ( .A(n11942), .B(n11934), .Z(c[1987]) );
  NAND U12996 ( .A(n11936), .B(n11935), .Z(n11940) );
  NANDN U12997 ( .A(n11938), .B(n11937), .Z(n11939) );
  NAND U12998 ( .A(n11940), .B(n11939), .Z(n11947) );
  ANDN U12999 ( .B(a[966]), .A(n3983), .Z(n11945) );
  AND U13000 ( .A(b[1]), .B(a[965]), .Z(n11944) );
  XOR U13001 ( .A(n11945), .B(n11944), .Z(n11946) );
  XNOR U13002 ( .A(n11947), .B(n11946), .Z(n11949) );
  XOR U13003 ( .A(sreg[1988]), .B(n11948), .Z(n11943) );
  XNOR U13004 ( .A(n11949), .B(n11943), .Z(c[1988]) );
  NAND U13005 ( .A(b[0]), .B(a[967]), .Z(n11952) );
  NAND U13006 ( .A(a[966]), .B(b[1]), .Z(n11951) );
  XNOR U13007 ( .A(n11952), .B(n11951), .Z(n11954) );
  XNOR U13008 ( .A(n11953), .B(n11954), .Z(n11958) );
  XOR U13009 ( .A(n11957), .B(sreg[1989]), .Z(n11950) );
  XNOR U13010 ( .A(n11958), .B(n11950), .Z(c[1989]) );
  NAND U13011 ( .A(n11952), .B(n11951), .Z(n11956) );
  NANDN U13012 ( .A(n11954), .B(n11953), .Z(n11955) );
  NAND U13013 ( .A(n11956), .B(n11955), .Z(n11963) );
  ANDN U13014 ( .B(a[968]), .A(n3983), .Z(n11961) );
  AND U13015 ( .A(b[1]), .B(a[967]), .Z(n11960) );
  XOR U13016 ( .A(n11961), .B(n11960), .Z(n11962) );
  XNOR U13017 ( .A(n11963), .B(n11962), .Z(n11965) );
  XOR U13018 ( .A(sreg[1990]), .B(n11964), .Z(n11959) );
  XNOR U13019 ( .A(n11965), .B(n11959), .Z(c[1990]) );
  NAND U13020 ( .A(b[0]), .B(a[969]), .Z(n11968) );
  NAND U13021 ( .A(a[968]), .B(b[1]), .Z(n11967) );
  XNOR U13022 ( .A(n11968), .B(n11967), .Z(n11970) );
  XNOR U13023 ( .A(n11969), .B(n11970), .Z(n11974) );
  XOR U13024 ( .A(n11973), .B(sreg[1991]), .Z(n11966) );
  XNOR U13025 ( .A(n11974), .B(n11966), .Z(c[1991]) );
  NAND U13026 ( .A(n11968), .B(n11967), .Z(n11972) );
  NANDN U13027 ( .A(n11970), .B(n11969), .Z(n11971) );
  NAND U13028 ( .A(n11972), .B(n11971), .Z(n11979) );
  ANDN U13029 ( .B(a[970]), .A(n3983), .Z(n11977) );
  AND U13030 ( .A(b[1]), .B(a[969]), .Z(n11976) );
  XOR U13031 ( .A(n11977), .B(n11976), .Z(n11978) );
  XNOR U13032 ( .A(n11979), .B(n11978), .Z(n11981) );
  XOR U13033 ( .A(sreg[1992]), .B(n11980), .Z(n11975) );
  XNOR U13034 ( .A(n11981), .B(n11975), .Z(c[1992]) );
  NAND U13035 ( .A(b[0]), .B(a[971]), .Z(n11984) );
  NAND U13036 ( .A(a[970]), .B(b[1]), .Z(n11983) );
  XNOR U13037 ( .A(n11984), .B(n11983), .Z(n11986) );
  XNOR U13038 ( .A(n11985), .B(n11986), .Z(n11990) );
  XOR U13039 ( .A(n11989), .B(sreg[1993]), .Z(n11982) );
  XNOR U13040 ( .A(n11990), .B(n11982), .Z(c[1993]) );
  NAND U13041 ( .A(n11984), .B(n11983), .Z(n11988) );
  NANDN U13042 ( .A(n11986), .B(n11985), .Z(n11987) );
  NAND U13043 ( .A(n11988), .B(n11987), .Z(n11995) );
  ANDN U13044 ( .B(a[972]), .A(n3983), .Z(n11993) );
  AND U13045 ( .A(b[1]), .B(a[971]), .Z(n11992) );
  XOR U13046 ( .A(n11993), .B(n11992), .Z(n11994) );
  XNOR U13047 ( .A(n11995), .B(n11994), .Z(n11997) );
  XOR U13048 ( .A(sreg[1994]), .B(n11996), .Z(n11991) );
  XNOR U13049 ( .A(n11997), .B(n11991), .Z(c[1994]) );
  NAND U13050 ( .A(b[0]), .B(a[973]), .Z(n12000) );
  NAND U13051 ( .A(a[972]), .B(b[1]), .Z(n11999) );
  XNOR U13052 ( .A(n12000), .B(n11999), .Z(n12002) );
  XNOR U13053 ( .A(n12001), .B(n12002), .Z(n12006) );
  XOR U13054 ( .A(n12005), .B(sreg[1995]), .Z(n11998) );
  XNOR U13055 ( .A(n12006), .B(n11998), .Z(c[1995]) );
  NAND U13056 ( .A(n12000), .B(n11999), .Z(n12004) );
  NANDN U13057 ( .A(n12002), .B(n12001), .Z(n12003) );
  NAND U13058 ( .A(n12004), .B(n12003), .Z(n12011) );
  ANDN U13059 ( .B(a[974]), .A(n3984), .Z(n12009) );
  AND U13060 ( .A(b[1]), .B(a[973]), .Z(n12008) );
  XOR U13061 ( .A(n12009), .B(n12008), .Z(n12010) );
  XNOR U13062 ( .A(n12011), .B(n12010), .Z(n12016) );
  XOR U13063 ( .A(sreg[1996]), .B(n12015), .Z(n12007) );
  XNOR U13064 ( .A(n12016), .B(n12007), .Z(c[1996]) );
  OR U13065 ( .A(n12009), .B(n12008), .Z(n12014) );
  IV U13066 ( .A(n12010), .Z(n12012) );
  NANDN U13067 ( .A(n12012), .B(n12011), .Z(n12013) );
  NAND U13068 ( .A(n12014), .B(n12013), .Z(n12021) );
  ANDN U13069 ( .B(a[975]), .A(n3984), .Z(n12019) );
  AND U13070 ( .A(b[1]), .B(a[974]), .Z(n12018) );
  XOR U13071 ( .A(n12019), .B(n12018), .Z(n12020) );
  XNOR U13072 ( .A(n12021), .B(n12020), .Z(n12023) );
  XNOR U13073 ( .A(sreg[1997]), .B(n12022), .Z(n12017) );
  XNOR U13074 ( .A(n12023), .B(n12017), .Z(c[1997]) );
  NAND U13075 ( .A(b[0]), .B(a[976]), .Z(n12026) );
  NAND U13076 ( .A(a[975]), .B(b[1]), .Z(n12025) );
  XNOR U13077 ( .A(n12026), .B(n12025), .Z(n12028) );
  XNOR U13078 ( .A(n12027), .B(n12028), .Z(n12032) );
  XOR U13079 ( .A(n12031), .B(sreg[1998]), .Z(n12024) );
  XNOR U13080 ( .A(n12032), .B(n12024), .Z(c[1998]) );
  NAND U13081 ( .A(n12026), .B(n12025), .Z(n12030) );
  NANDN U13082 ( .A(n12028), .B(n12027), .Z(n12029) );
  NAND U13083 ( .A(n12030), .B(n12029), .Z(n12036) );
  NAND U13084 ( .A(b[0]), .B(a[977]), .Z(n12035) );
  NAND U13085 ( .A(a[976]), .B(b[1]), .Z(n12034) );
  XNOR U13086 ( .A(n12035), .B(n12034), .Z(n12037) );
  XNOR U13087 ( .A(n12036), .B(n12037), .Z(n12041) );
  XOR U13088 ( .A(n12040), .B(sreg[1999]), .Z(n12033) );
  XNOR U13089 ( .A(n12041), .B(n12033), .Z(c[1999]) );
  NAND U13090 ( .A(n12035), .B(n12034), .Z(n12039) );
  NANDN U13091 ( .A(n12037), .B(n12036), .Z(n12038) );
  NAND U13092 ( .A(n12039), .B(n12038), .Z(n12046) );
  ANDN U13093 ( .B(a[978]), .A(n3984), .Z(n12044) );
  AND U13094 ( .A(b[1]), .B(a[977]), .Z(n12043) );
  XOR U13095 ( .A(n12044), .B(n12043), .Z(n12045) );
  XNOR U13096 ( .A(n12046), .B(n12045), .Z(n12048) );
  XOR U13097 ( .A(sreg[2000]), .B(n12047), .Z(n12042) );
  XNOR U13098 ( .A(n12048), .B(n12042), .Z(c[2000]) );
  NAND U13099 ( .A(b[0]), .B(a[979]), .Z(n12051) );
  NAND U13100 ( .A(a[978]), .B(b[1]), .Z(n12050) );
  XNOR U13101 ( .A(n12051), .B(n12050), .Z(n12053) );
  XNOR U13102 ( .A(n12052), .B(n12053), .Z(n12057) );
  XOR U13103 ( .A(n12056), .B(sreg[2001]), .Z(n12049) );
  XNOR U13104 ( .A(n12057), .B(n12049), .Z(c[2001]) );
  NAND U13105 ( .A(n12051), .B(n12050), .Z(n12055) );
  NANDN U13106 ( .A(n12053), .B(n12052), .Z(n12054) );
  NAND U13107 ( .A(n12055), .B(n12054), .Z(n12062) );
  ANDN U13108 ( .B(a[980]), .A(n3984), .Z(n12060) );
  AND U13109 ( .A(b[1]), .B(a[979]), .Z(n12059) );
  XOR U13110 ( .A(n12060), .B(n12059), .Z(n12061) );
  XNOR U13111 ( .A(n12062), .B(n12061), .Z(n12064) );
  XOR U13112 ( .A(sreg[2002]), .B(n12063), .Z(n12058) );
  XNOR U13113 ( .A(n12064), .B(n12058), .Z(c[2002]) );
  NAND U13114 ( .A(b[0]), .B(a[981]), .Z(n12067) );
  NAND U13115 ( .A(a[980]), .B(b[1]), .Z(n12066) );
  XNOR U13116 ( .A(n12067), .B(n12066), .Z(n12069) );
  XNOR U13117 ( .A(n12068), .B(n12069), .Z(n12073) );
  XOR U13118 ( .A(n12072), .B(sreg[2003]), .Z(n12065) );
  XNOR U13119 ( .A(n12073), .B(n12065), .Z(c[2003]) );
  NAND U13120 ( .A(n12067), .B(n12066), .Z(n12071) );
  NANDN U13121 ( .A(n12069), .B(n12068), .Z(n12070) );
  NAND U13122 ( .A(n12071), .B(n12070), .Z(n12078) );
  ANDN U13123 ( .B(a[982]), .A(n3984), .Z(n12076) );
  AND U13124 ( .A(b[1]), .B(a[981]), .Z(n12075) );
  XOR U13125 ( .A(n12076), .B(n12075), .Z(n12077) );
  XNOR U13126 ( .A(n12078), .B(n12077), .Z(n12080) );
  XOR U13127 ( .A(sreg[2004]), .B(n12079), .Z(n12074) );
  XNOR U13128 ( .A(n12080), .B(n12074), .Z(c[2004]) );
  ANDN U13129 ( .B(a[983]), .A(n3984), .Z(n12083) );
  AND U13130 ( .A(b[1]), .B(a[982]), .Z(n12082) );
  XOR U13131 ( .A(n12083), .B(n12082), .Z(n12084) );
  XNOR U13132 ( .A(n12085), .B(n12084), .Z(n12087) );
  XNOR U13133 ( .A(sreg[2005]), .B(n12086), .Z(n12081) );
  XNOR U13134 ( .A(n12087), .B(n12081), .Z(c[2005]) );
  ANDN U13135 ( .B(a[984]), .A(n3984), .Z(n12090) );
  AND U13136 ( .A(b[1]), .B(a[983]), .Z(n12089) );
  XOR U13137 ( .A(n12090), .B(n12089), .Z(n12091) );
  XNOR U13138 ( .A(n12092), .B(n12091), .Z(n12094) );
  XNOR U13139 ( .A(sreg[2006]), .B(n12093), .Z(n12088) );
  XNOR U13140 ( .A(n12094), .B(n12088), .Z(c[2006]) );
  NAND U13141 ( .A(b[0]), .B(a[985]), .Z(n12097) );
  NAND U13142 ( .A(a[984]), .B(b[1]), .Z(n12096) );
  XNOR U13143 ( .A(n12097), .B(n12096), .Z(n12099) );
  XNOR U13144 ( .A(n12098), .B(n12099), .Z(n12103) );
  XOR U13145 ( .A(n12102), .B(sreg[2007]), .Z(n12095) );
  XNOR U13146 ( .A(n12103), .B(n12095), .Z(c[2007]) );
  NAND U13147 ( .A(n12097), .B(n12096), .Z(n12101) );
  NANDN U13148 ( .A(n12099), .B(n12098), .Z(n12100) );
  NAND U13149 ( .A(n12101), .B(n12100), .Z(n12108) );
  ANDN U13150 ( .B(a[986]), .A(n3985), .Z(n12106) );
  AND U13151 ( .A(b[1]), .B(a[985]), .Z(n12105) );
  XOR U13152 ( .A(n12106), .B(n12105), .Z(n12107) );
  XNOR U13153 ( .A(n12108), .B(n12107), .Z(n12113) );
  XOR U13154 ( .A(sreg[2008]), .B(n12112), .Z(n12104) );
  XNOR U13155 ( .A(n12113), .B(n12104), .Z(c[2008]) );
  OR U13156 ( .A(n12106), .B(n12105), .Z(n12111) );
  IV U13157 ( .A(n12107), .Z(n12109) );
  NANDN U13158 ( .A(n12109), .B(n12108), .Z(n12110) );
  NAND U13159 ( .A(n12111), .B(n12110), .Z(n12118) );
  ANDN U13160 ( .B(a[987]), .A(n3985), .Z(n12116) );
  AND U13161 ( .A(b[1]), .B(a[986]), .Z(n12115) );
  XOR U13162 ( .A(n12116), .B(n12115), .Z(n12117) );
  XNOR U13163 ( .A(n12118), .B(n12117), .Z(n12120) );
  XNOR U13164 ( .A(sreg[2009]), .B(n12119), .Z(n12114) );
  XNOR U13165 ( .A(n12120), .B(n12114), .Z(c[2009]) );
  ANDN U13166 ( .B(a[988]), .A(n3985), .Z(n12123) );
  AND U13167 ( .A(b[1]), .B(a[987]), .Z(n12122) );
  XOR U13168 ( .A(n12123), .B(n12122), .Z(n12124) );
  XNOR U13169 ( .A(n12125), .B(n12124), .Z(n12127) );
  XNOR U13170 ( .A(sreg[2010]), .B(n12126), .Z(n12121) );
  XNOR U13171 ( .A(n12127), .B(n12121), .Z(c[2010]) );
  NAND U13172 ( .A(b[0]), .B(a[989]), .Z(n12130) );
  NAND U13173 ( .A(a[988]), .B(b[1]), .Z(n12129) );
  XNOR U13174 ( .A(n12130), .B(n12129), .Z(n12132) );
  XNOR U13175 ( .A(n12131), .B(n12132), .Z(n12136) );
  XOR U13176 ( .A(n12135), .B(sreg[2011]), .Z(n12128) );
  XNOR U13177 ( .A(n12136), .B(n12128), .Z(c[2011]) );
  NAND U13178 ( .A(n12130), .B(n12129), .Z(n12134) );
  NANDN U13179 ( .A(n12132), .B(n12131), .Z(n12133) );
  NAND U13180 ( .A(n12134), .B(n12133), .Z(n12141) );
  ANDN U13181 ( .B(a[990]), .A(n3985), .Z(n12139) );
  AND U13182 ( .A(b[1]), .B(a[989]), .Z(n12138) );
  XOR U13183 ( .A(n12139), .B(n12138), .Z(n12140) );
  XNOR U13184 ( .A(n12141), .B(n12140), .Z(n12143) );
  XOR U13185 ( .A(sreg[2012]), .B(n12142), .Z(n12137) );
  XNOR U13186 ( .A(n12143), .B(n12137), .Z(c[2012]) );
  NAND U13187 ( .A(b[0]), .B(a[991]), .Z(n12146) );
  NAND U13188 ( .A(a[990]), .B(b[1]), .Z(n12145) );
  XNOR U13189 ( .A(n12146), .B(n12145), .Z(n12148) );
  XNOR U13190 ( .A(n12147), .B(n12148), .Z(n12152) );
  XOR U13191 ( .A(n12151), .B(sreg[2013]), .Z(n12144) );
  XNOR U13192 ( .A(n12152), .B(n12144), .Z(c[2013]) );
  NAND U13193 ( .A(n12146), .B(n12145), .Z(n12150) );
  NANDN U13194 ( .A(n12148), .B(n12147), .Z(n12149) );
  NAND U13195 ( .A(n12150), .B(n12149), .Z(n12157) );
  ANDN U13196 ( .B(a[992]), .A(n3985), .Z(n12155) );
  AND U13197 ( .A(b[1]), .B(a[991]), .Z(n12154) );
  XOR U13198 ( .A(n12155), .B(n12154), .Z(n12156) );
  XNOR U13199 ( .A(n12157), .B(n12156), .Z(n12159) );
  XOR U13200 ( .A(sreg[2014]), .B(n12158), .Z(n12153) );
  XNOR U13201 ( .A(n12159), .B(n12153), .Z(c[2014]) );
  NAND U13202 ( .A(b[0]), .B(a[993]), .Z(n12162) );
  NAND U13203 ( .A(a[992]), .B(b[1]), .Z(n12161) );
  XNOR U13204 ( .A(n12162), .B(n12161), .Z(n12164) );
  XNOR U13205 ( .A(n12163), .B(n12164), .Z(n12168) );
  XOR U13206 ( .A(n12167), .B(sreg[2015]), .Z(n12160) );
  XNOR U13207 ( .A(n12168), .B(n12160), .Z(c[2015]) );
  NAND U13208 ( .A(n12162), .B(n12161), .Z(n12166) );
  NANDN U13209 ( .A(n12164), .B(n12163), .Z(n12165) );
  NAND U13210 ( .A(n12166), .B(n12165), .Z(n12173) );
  ANDN U13211 ( .B(a[994]), .A(n3985), .Z(n12171) );
  AND U13212 ( .A(b[1]), .B(a[993]), .Z(n12170) );
  XOR U13213 ( .A(n12171), .B(n12170), .Z(n12172) );
  XNOR U13214 ( .A(n12173), .B(n12172), .Z(n12175) );
  XOR U13215 ( .A(sreg[2016]), .B(n12174), .Z(n12169) );
  XNOR U13216 ( .A(n12175), .B(n12169), .Z(c[2016]) );
  NAND U13217 ( .A(b[0]), .B(a[995]), .Z(n12178) );
  NAND U13218 ( .A(a[994]), .B(b[1]), .Z(n12177) );
  XNOR U13219 ( .A(n12178), .B(n12177), .Z(n12180) );
  XNOR U13220 ( .A(n12179), .B(n12180), .Z(n12184) );
  XOR U13221 ( .A(n12183), .B(sreg[2017]), .Z(n12176) );
  XNOR U13222 ( .A(n12184), .B(n12176), .Z(c[2017]) );
  NAND U13223 ( .A(n12178), .B(n12177), .Z(n12182) );
  NANDN U13224 ( .A(n12180), .B(n12179), .Z(n12181) );
  NAND U13225 ( .A(n12182), .B(n12181), .Z(n12189) );
  ANDN U13226 ( .B(a[996]), .A(n3985), .Z(n12187) );
  AND U13227 ( .A(b[1]), .B(a[995]), .Z(n12186) );
  XOR U13228 ( .A(n12187), .B(n12186), .Z(n12188) );
  XNOR U13229 ( .A(n12189), .B(n12188), .Z(n12191) );
  XOR U13230 ( .A(sreg[2018]), .B(n12190), .Z(n12185) );
  XNOR U13231 ( .A(n12191), .B(n12185), .Z(c[2018]) );
  NAND U13232 ( .A(b[0]), .B(a[997]), .Z(n12194) );
  NAND U13233 ( .A(a[996]), .B(b[1]), .Z(n12193) );
  XNOR U13234 ( .A(n12194), .B(n12193), .Z(n12196) );
  XNOR U13235 ( .A(n12195), .B(n12196), .Z(n12200) );
  XOR U13236 ( .A(n12199), .B(sreg[2019]), .Z(n12192) );
  XNOR U13237 ( .A(n12200), .B(n12192), .Z(c[2019]) );
  NAND U13238 ( .A(n12194), .B(n12193), .Z(n12198) );
  NANDN U13239 ( .A(n12196), .B(n12195), .Z(n12197) );
  NAND U13240 ( .A(n12198), .B(n12197), .Z(n12205) );
  ANDN U13241 ( .B(a[998]), .A(n3986), .Z(n12203) );
  AND U13242 ( .A(b[1]), .B(a[997]), .Z(n12202) );
  XOR U13243 ( .A(n12203), .B(n12202), .Z(n12204) );
  XNOR U13244 ( .A(n12205), .B(n12204), .Z(n12210) );
  XOR U13245 ( .A(sreg[2020]), .B(n12209), .Z(n12201) );
  XNOR U13246 ( .A(n12210), .B(n12201), .Z(c[2020]) );
  OR U13247 ( .A(n12203), .B(n12202), .Z(n12208) );
  IV U13248 ( .A(n12204), .Z(n12206) );
  NANDN U13249 ( .A(n12206), .B(n12205), .Z(n12207) );
  NAND U13250 ( .A(n12208), .B(n12207), .Z(n12215) );
  ANDN U13251 ( .B(a[999]), .A(n3986), .Z(n12213) );
  AND U13252 ( .A(b[1]), .B(a[998]), .Z(n12212) );
  XOR U13253 ( .A(n12213), .B(n12212), .Z(n12214) );
  XNOR U13254 ( .A(n12215), .B(n12214), .Z(n12217) );
  XNOR U13255 ( .A(sreg[2021]), .B(n12216), .Z(n12211) );
  XNOR U13256 ( .A(n12217), .B(n12211), .Z(c[2021]) );
  ANDN U13257 ( .B(a[1000]), .A(n3986), .Z(n12220) );
  AND U13258 ( .A(b[1]), .B(a[999]), .Z(n12219) );
  XOR U13259 ( .A(n12220), .B(n12219), .Z(n12221) );
  XNOR U13260 ( .A(n12222), .B(n12221), .Z(n12224) );
  XNOR U13261 ( .A(sreg[2022]), .B(n12223), .Z(n12218) );
  XNOR U13262 ( .A(n12224), .B(n12218), .Z(c[2022]) );
  NAND U13263 ( .A(b[0]), .B(a[1001]), .Z(n12227) );
  NAND U13264 ( .A(a[1000]), .B(b[1]), .Z(n12226) );
  XNOR U13265 ( .A(n12227), .B(n12226), .Z(n12229) );
  XNOR U13266 ( .A(n12228), .B(n12229), .Z(n12233) );
  XOR U13267 ( .A(n12232), .B(sreg[2023]), .Z(n12225) );
  XNOR U13268 ( .A(n12233), .B(n12225), .Z(c[2023]) );
  NAND U13269 ( .A(n12227), .B(n12226), .Z(n12231) );
  NANDN U13270 ( .A(n12229), .B(n12228), .Z(n12230) );
  NAND U13271 ( .A(n12231), .B(n12230), .Z(n12237) );
  NAND U13272 ( .A(b[0]), .B(a[1002]), .Z(n12236) );
  NAND U13273 ( .A(a[1001]), .B(b[1]), .Z(n12235) );
  XNOR U13274 ( .A(n12236), .B(n12235), .Z(n12238) );
  XNOR U13275 ( .A(n12237), .B(n12238), .Z(n12242) );
  XOR U13276 ( .A(n12241), .B(sreg[2024]), .Z(n12234) );
  XNOR U13277 ( .A(n12242), .B(n12234), .Z(c[2024]) );
  NAND U13278 ( .A(n12236), .B(n12235), .Z(n12240) );
  NANDN U13279 ( .A(n12238), .B(n12237), .Z(n12239) );
  NAND U13280 ( .A(n12240), .B(n12239), .Z(n12246) );
  NAND U13281 ( .A(b[0]), .B(a[1003]), .Z(n12245) );
  NAND U13282 ( .A(a[1002]), .B(b[1]), .Z(n12244) );
  XNOR U13283 ( .A(n12245), .B(n12244), .Z(n12247) );
  XNOR U13284 ( .A(n12246), .B(n12247), .Z(n12251) );
  XOR U13285 ( .A(n12250), .B(sreg[2025]), .Z(n12243) );
  XNOR U13286 ( .A(n12251), .B(n12243), .Z(c[2025]) );
  NAND U13287 ( .A(n12245), .B(n12244), .Z(n12249) );
  NANDN U13288 ( .A(n12247), .B(n12246), .Z(n12248) );
  NAND U13289 ( .A(n12249), .B(n12248), .Z(n12256) );
  ANDN U13290 ( .B(a[1004]), .A(n3986), .Z(n12254) );
  AND U13291 ( .A(b[1]), .B(a[1003]), .Z(n12253) );
  XOR U13292 ( .A(n12254), .B(n12253), .Z(n12255) );
  XNOR U13293 ( .A(n12256), .B(n12255), .Z(n12258) );
  XOR U13294 ( .A(sreg[2026]), .B(n12257), .Z(n12252) );
  XNOR U13295 ( .A(n12258), .B(n12252), .Z(c[2026]) );
  NAND U13296 ( .A(b[0]), .B(a[1005]), .Z(n12261) );
  NAND U13297 ( .A(a[1004]), .B(b[1]), .Z(n12260) );
  XNOR U13298 ( .A(n12261), .B(n12260), .Z(n12263) );
  XNOR U13299 ( .A(n12262), .B(n12263), .Z(n12267) );
  XOR U13300 ( .A(n12266), .B(sreg[2027]), .Z(n12259) );
  XNOR U13301 ( .A(n12267), .B(n12259), .Z(c[2027]) );
  NAND U13302 ( .A(n12261), .B(n12260), .Z(n12265) );
  NANDN U13303 ( .A(n12263), .B(n12262), .Z(n12264) );
  NAND U13304 ( .A(n12265), .B(n12264), .Z(n12272) );
  ANDN U13305 ( .B(a[1006]), .A(n3986), .Z(n12270) );
  AND U13306 ( .A(b[1]), .B(a[1005]), .Z(n12269) );
  XOR U13307 ( .A(n12270), .B(n12269), .Z(n12271) );
  XNOR U13308 ( .A(n12272), .B(n12271), .Z(n12274) );
  XOR U13309 ( .A(sreg[2028]), .B(n12273), .Z(n12268) );
  XNOR U13310 ( .A(n12274), .B(n12268), .Z(c[2028]) );
  ANDN U13311 ( .B(a[1007]), .A(n3986), .Z(n12277) );
  AND U13312 ( .A(b[1]), .B(a[1006]), .Z(n12276) );
  XOR U13313 ( .A(n12277), .B(n12276), .Z(n12278) );
  XNOR U13314 ( .A(n12279), .B(n12278), .Z(n12281) );
  XNOR U13315 ( .A(sreg[2029]), .B(n12280), .Z(n12275) );
  XNOR U13316 ( .A(n12281), .B(n12275), .Z(c[2029]) );
  NAND U13317 ( .A(b[0]), .B(a[1008]), .Z(n12284) );
  NAND U13318 ( .A(a[1007]), .B(b[1]), .Z(n12283) );
  XNOR U13319 ( .A(n12284), .B(n12283), .Z(n12286) );
  XNOR U13320 ( .A(n12285), .B(n12286), .Z(n12290) );
  XOR U13321 ( .A(n12289), .B(sreg[2030]), .Z(n12282) );
  XNOR U13322 ( .A(n12290), .B(n12282), .Z(c[2030]) );
  NAND U13323 ( .A(n12284), .B(n12283), .Z(n12288) );
  NANDN U13324 ( .A(n12286), .B(n12285), .Z(n12287) );
  NAND U13325 ( .A(n12288), .B(n12287), .Z(n12294) );
  NAND U13326 ( .A(b[0]), .B(a[1009]), .Z(n12293) );
  NAND U13327 ( .A(a[1008]), .B(b[1]), .Z(n12292) );
  XNOR U13328 ( .A(n12293), .B(n12292), .Z(n12295) );
  XNOR U13329 ( .A(n12294), .B(n12295), .Z(n12299) );
  XOR U13330 ( .A(n12298), .B(sreg[2031]), .Z(n12291) );
  XNOR U13331 ( .A(n12299), .B(n12291), .Z(c[2031]) );
  NAND U13332 ( .A(n12293), .B(n12292), .Z(n12297) );
  NANDN U13333 ( .A(n12295), .B(n12294), .Z(n12296) );
  NAND U13334 ( .A(n12297), .B(n12296), .Z(n12304) );
  ANDN U13335 ( .B(a[1010]), .A(n3986), .Z(n12302) );
  AND U13336 ( .A(b[1]), .B(a[1009]), .Z(n12301) );
  XOR U13337 ( .A(n12302), .B(n12301), .Z(n12303) );
  XNOR U13338 ( .A(n12304), .B(n12303), .Z(n12306) );
  XOR U13339 ( .A(sreg[2032]), .B(n12305), .Z(n12300) );
  XNOR U13340 ( .A(n12306), .B(n12300), .Z(c[2032]) );
  NAND U13341 ( .A(b[0]), .B(a[1011]), .Z(n12309) );
  NAND U13342 ( .A(a[1010]), .B(b[1]), .Z(n12308) );
  XNOR U13343 ( .A(n12309), .B(n12308), .Z(n12311) );
  XNOR U13344 ( .A(n12310), .B(n12311), .Z(n12315) );
  XOR U13345 ( .A(n12314), .B(sreg[2033]), .Z(n12307) );
  XNOR U13346 ( .A(n12315), .B(n12307), .Z(c[2033]) );
  NAND U13347 ( .A(n12309), .B(n12308), .Z(n12313) );
  NANDN U13348 ( .A(n12311), .B(n12310), .Z(n12312) );
  NAND U13349 ( .A(n12313), .B(n12312), .Z(n12319) );
  NAND U13350 ( .A(b[0]), .B(a[1012]), .Z(n12318) );
  NAND U13351 ( .A(a[1011]), .B(b[1]), .Z(n12317) );
  XNOR U13352 ( .A(n12318), .B(n12317), .Z(n12320) );
  XNOR U13353 ( .A(n12319), .B(n12320), .Z(n12324) );
  XOR U13354 ( .A(n12323), .B(sreg[2034]), .Z(n12316) );
  XNOR U13355 ( .A(n12324), .B(n12316), .Z(c[2034]) );
  NAND U13356 ( .A(n12318), .B(n12317), .Z(n12322) );
  NANDN U13357 ( .A(n12320), .B(n12319), .Z(n12321) );
  NAND U13358 ( .A(n12322), .B(n12321), .Z(n12328) );
  NAND U13359 ( .A(b[0]), .B(a[1013]), .Z(n12327) );
  NAND U13360 ( .A(a[1012]), .B(b[1]), .Z(n12326) );
  XNOR U13361 ( .A(n12327), .B(n12326), .Z(n12329) );
  XNOR U13362 ( .A(n12328), .B(n12329), .Z(n12333) );
  XOR U13363 ( .A(n12332), .B(sreg[2035]), .Z(n12325) );
  XNOR U13364 ( .A(n12333), .B(n12325), .Z(c[2035]) );
  NAND U13365 ( .A(n12327), .B(n12326), .Z(n12331) );
  NANDN U13366 ( .A(n12329), .B(n12328), .Z(n12330) );
  NAND U13367 ( .A(n12331), .B(n12330), .Z(n12338) );
  ANDN U13368 ( .B(a[1014]), .A(n3987), .Z(n12336) );
  AND U13369 ( .A(b[1]), .B(a[1013]), .Z(n12335) );
  XOR U13370 ( .A(n12336), .B(n12335), .Z(n12337) );
  XNOR U13371 ( .A(n12338), .B(n12337), .Z(n12340) );
  XOR U13372 ( .A(sreg[2036]), .B(n12339), .Z(n12334) );
  XNOR U13373 ( .A(n12340), .B(n12334), .Z(c[2036]) );
  NAND U13374 ( .A(b[0]), .B(a[1015]), .Z(n12343) );
  NAND U13375 ( .A(a[1014]), .B(b[1]), .Z(n12342) );
  XNOR U13376 ( .A(n12343), .B(n12342), .Z(n12345) );
  XNOR U13377 ( .A(n12344), .B(n12345), .Z(n12349) );
  XOR U13378 ( .A(n12348), .B(sreg[2037]), .Z(n12341) );
  XNOR U13379 ( .A(n12349), .B(n12341), .Z(c[2037]) );
  NAND U13380 ( .A(n12343), .B(n12342), .Z(n12347) );
  NANDN U13381 ( .A(n12345), .B(n12344), .Z(n12346) );
  NAND U13382 ( .A(n12347), .B(n12346), .Z(n12354) );
  ANDN U13383 ( .B(a[1016]), .A(n3987), .Z(n12352) );
  AND U13384 ( .A(b[1]), .B(a[1015]), .Z(n12351) );
  XOR U13385 ( .A(n12352), .B(n12351), .Z(n12353) );
  XNOR U13386 ( .A(n12354), .B(n12353), .Z(n12356) );
  XOR U13387 ( .A(sreg[2038]), .B(n12355), .Z(n12350) );
  XNOR U13388 ( .A(n12356), .B(n12350), .Z(c[2038]) );
  NAND U13389 ( .A(b[0]), .B(a[1017]), .Z(n12359) );
  NAND U13390 ( .A(a[1016]), .B(b[1]), .Z(n12358) );
  XNOR U13391 ( .A(n12359), .B(n12358), .Z(n12361) );
  XNOR U13392 ( .A(n12360), .B(n12361), .Z(n12365) );
  XOR U13393 ( .A(n12364), .B(sreg[2039]), .Z(n12357) );
  XNOR U13394 ( .A(n12365), .B(n12357), .Z(c[2039]) );
  NAND U13395 ( .A(n12359), .B(n12358), .Z(n12363) );
  NANDN U13396 ( .A(n12361), .B(n12360), .Z(n12362) );
  NAND U13397 ( .A(n12363), .B(n12362), .Z(n12370) );
  ANDN U13398 ( .B(a[1018]), .A(n3987), .Z(n12368) );
  AND U13399 ( .A(b[1]), .B(a[1017]), .Z(n12367) );
  XOR U13400 ( .A(n12368), .B(n12367), .Z(n12369) );
  XNOR U13401 ( .A(n12370), .B(n12369), .Z(n12372) );
  XOR U13402 ( .A(sreg[2040]), .B(n12371), .Z(n12366) );
  XNOR U13403 ( .A(n12372), .B(n12366), .Z(c[2040]) );
  NAND U13404 ( .A(b[0]), .B(a[1019]), .Z(n12375) );
  NAND U13405 ( .A(a[1018]), .B(b[1]), .Z(n12374) );
  XNOR U13406 ( .A(n12375), .B(n12374), .Z(n12377) );
  XNOR U13407 ( .A(n12376), .B(n12377), .Z(n12381) );
  XOR U13408 ( .A(n12380), .B(sreg[2041]), .Z(n12373) );
  XNOR U13409 ( .A(n12381), .B(n12373), .Z(c[2041]) );
  NAND U13410 ( .A(n12375), .B(n12374), .Z(n12379) );
  NANDN U13411 ( .A(n12377), .B(n12376), .Z(n12378) );
  NAND U13412 ( .A(n12379), .B(n12378), .Z(n12386) );
  ANDN U13413 ( .B(a[1020]), .A(n3987), .Z(n12384) );
  AND U13414 ( .A(b[1]), .B(a[1019]), .Z(n12383) );
  XOR U13415 ( .A(n12384), .B(n12383), .Z(n12385) );
  XNOR U13416 ( .A(n12386), .B(n12385), .Z(n12388) );
  XOR U13417 ( .A(sreg[2042]), .B(n12387), .Z(n12382) );
  XNOR U13418 ( .A(n12388), .B(n12382), .Z(c[2042]) );
  NAND U13419 ( .A(b[0]), .B(a[1021]), .Z(n12391) );
  NAND U13420 ( .A(a[1020]), .B(b[1]), .Z(n12390) );
  XNOR U13421 ( .A(n12391), .B(n12390), .Z(n12393) );
  XNOR U13422 ( .A(n12392), .B(n12393), .Z(n12397) );
  XOR U13423 ( .A(n12396), .B(sreg[2043]), .Z(n12389) );
  XNOR U13424 ( .A(n12397), .B(n12389), .Z(c[2043]) );
  NAND U13425 ( .A(n12391), .B(n12390), .Z(n12395) );
  NANDN U13426 ( .A(n12393), .B(n12392), .Z(n12394) );
  NAND U13427 ( .A(n12395), .B(n12394), .Z(n12402) );
  ANDN U13428 ( .B(a[1022]), .A(n3987), .Z(n12399) );
  IV U13429 ( .A(n12399), .Z(n12410) );
  AND U13430 ( .A(a[1021]), .B(b[1]), .Z(n12400) );
  XNOR U13431 ( .A(n12410), .B(n12400), .Z(n12401) );
  XNOR U13432 ( .A(n12402), .B(n12401), .Z(n12408) );
  XOR U13433 ( .A(n12407), .B(sreg[2044]), .Z(n12398) );
  XOR U13434 ( .A(n12408), .B(n12398), .Z(c[2044]) );
  OR U13435 ( .A(n12400), .B(n12399), .Z(n12404) );
  NAND U13436 ( .A(n12402), .B(n12401), .Z(n12403) );
  NAND U13437 ( .A(n12404), .B(n12403), .Z(n12412) );
  ANDN U13438 ( .B(a[1023]), .A(n3987), .Z(n12406) );
  NAND U13439 ( .A(b[1]), .B(a[1022]), .Z(n12405) );
  XOR U13440 ( .A(n12406), .B(n12405), .Z(n12411) );
  XOR U13441 ( .A(n12412), .B(n12411), .Z(n12416) );
  XOR U13442 ( .A(n12415), .B(sreg[2045]), .Z(n12409) );
  XOR U13443 ( .A(n12416), .B(n12409), .Z(c[2045]) );
  AND U13444 ( .A(a[1023]), .B(b[1]), .Z(n12419) );
  NANDN U13445 ( .A(n12410), .B(n12419), .Z(n12414) );
  OR U13446 ( .A(n12412), .B(n12411), .Z(n12413) );
  NAND U13447 ( .A(n12414), .B(n12413), .Z(n12421) );
  XOR U13448 ( .A(n12419), .B(n12420), .Z(n12417) );
  XOR U13449 ( .A(n12421), .B(n12417), .Z(c[2046]) );
  XOR U13450 ( .A(n12421), .B(n12420), .Z(n12418) );
  NANDN U13451 ( .A(n12419), .B(n12418), .Z(n12423) );
  OR U13452 ( .A(n12421), .B(n12420), .Z(n12422) );
  AND U13453 ( .A(n12423), .B(n12422), .Z(c[2047]) );
endmodule

