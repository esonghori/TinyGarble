
module SubBytes_0 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042;

  XNOR U2962 ( .A(n2145), .B(n2148), .Z(n2168) );
  XNOR U2963 ( .A(x[103]), .B(x[98]), .Z(n3465) );
  XOR U2964 ( .A(n3655), .B(n3654), .Z(n1987) );
  XNOR U2965 ( .A(z[10]), .B(n3656), .Z(n1988) );
  XNOR U2966 ( .A(n1987), .B(n1988), .Z(z[9]) );
  ANDN U2967 ( .B(n3589), .A(n3597), .Z(n1989) );
  XNOR U2968 ( .A(n3350), .B(n3354), .Z(n1990) );
  XNOR U2969 ( .A(n1989), .B(n1990), .Z(n3377) );
  ANDN U2970 ( .B(n3774), .A(n3782), .Z(n1991) );
  XNOR U2971 ( .A(n2471), .B(n2475), .Z(n1992) );
  XNOR U2972 ( .A(n1991), .B(n1992), .Z(n2498) );
  ANDN U2973 ( .B(n3421), .A(n3764), .Z(n1993) );
  XNOR U2974 ( .A(n2046), .B(n2050), .Z(n1994) );
  XNOR U2975 ( .A(n1993), .B(n1994), .Z(n2073) );
  ANDN U2976 ( .B(n3931), .A(n3939), .Z(n1995) );
  XNOR U2977 ( .A(n2839), .B(n2843), .Z(n1996) );
  XNOR U2978 ( .A(n1995), .B(n1996), .Z(n2866) );
  ANDN U2979 ( .B(n3523), .A(n3531), .Z(n1997) );
  XNOR U2980 ( .A(n3258), .B(n3262), .Z(n1998) );
  XNOR U2981 ( .A(n1997), .B(n1998), .Z(n3285) );
  ANDN U2982 ( .B(n3694), .A(n3702), .Z(n1999) );
  XNOR U2983 ( .A(n2287), .B(n2291), .Z(n2000) );
  XNOR U2984 ( .A(n1999), .B(n2000), .Z(n2314) );
  ANDN U2985 ( .B(n3729), .A(n3737), .Z(n2001) );
  XNOR U2986 ( .A(n2379), .B(n2383), .Z(n2002) );
  XNOR U2987 ( .A(n2001), .B(n2002), .Z(n2406) );
  ANDN U2988 ( .B(n3894), .A(n3902), .Z(n2003) );
  XNOR U2989 ( .A(n2747), .B(n2751), .Z(n2004) );
  XNOR U2990 ( .A(n2003), .B(n2004), .Z(n2774) );
  ANDN U2991 ( .B(n3488), .A(n3496), .Z(n2005) );
  XNOR U2992 ( .A(n3166), .B(n3170), .Z(n2006) );
  XNOR U2993 ( .A(n2005), .B(n2006), .Z(n3193) );
  ANDN U2994 ( .B(n3845), .A(n3853), .Z(n2007) );
  XNOR U2995 ( .A(n2655), .B(n2659), .Z(n2008) );
  XNOR U2996 ( .A(n2007), .B(n2008), .Z(n2682) );
  ANDN U2997 ( .B(n3659), .A(n3667), .Z(n2009) );
  XNOR U2998 ( .A(n2195), .B(n2199), .Z(n2010) );
  XNOR U2999 ( .A(n2009), .B(n2010), .Z(n2222) );
  XNOR U3000 ( .A(n3567), .B(n2116), .Z(n2167) );
  XOR U3001 ( .A(n3623), .B(n3637), .Z(n3581) );
  ANDN U3002 ( .B(n3809), .A(n3818), .Z(n2011) );
  XNOR U3003 ( .A(n2563), .B(n2567), .Z(n2012) );
  XNOR U3004 ( .A(n2011), .B(n2012), .Z(n2590) );
  NAND U3005 ( .A(n2942), .B(n2963), .Z(n2013) );
  OR U3006 ( .A(n2989), .B(n2963), .Z(n2014) );
  NAND U3007 ( .A(n2013), .B(n2014), .Z(n2015) );
  XNOR U3008 ( .A(n2978), .B(n2015), .Z(n2016) );
  XOR U3009 ( .A(n2932), .B(n2919), .Z(n2017) );
  XNOR U3010 ( .A(n2016), .B(n2017), .Z(n2957) );
  XNOR U3011 ( .A(n3471), .B(n3463), .Z(n3444) );
  NAND U3012 ( .A(n3029), .B(n3050), .Z(n2018) );
  OR U3013 ( .A(n3076), .B(n3050), .Z(n2019) );
  NAND U3014 ( .A(n2018), .B(n2019), .Z(n2020) );
  XNOR U3015 ( .A(n3065), .B(n2020), .Z(n2021) );
  XOR U3016 ( .A(n3019), .B(n3006), .Z(n2022) );
  XNOR U3017 ( .A(n2021), .B(n2022), .Z(n3044) );
  XOR U3018 ( .A(x[98]), .B(n3084), .Z(n2023) );
  XNOR U3019 ( .A(n3083), .B(n2023), .Z(n3430) );
  IV U3020 ( .A(x[4]), .Z(n2024) );
  IV U3021 ( .A(x[0]), .Z(n2109) );
  XOR U3022 ( .A(n2109), .B(x[6]), .Z(n2025) );
  XOR U3023 ( .A(n2025), .B(x[5]), .Z(n2049) );
  IV U3024 ( .A(n2049), .Z(n3867) );
  XOR U3025 ( .A(n2024), .B(n3867), .Z(n2098) );
  XOR U3026 ( .A(x[1]), .B(x[3]), .Z(n2026) );
  XOR U3027 ( .A(x[7]), .B(n2024), .Z(n2084) );
  XNOR U3028 ( .A(n2026), .B(n2084), .Z(n2063) );
  IV U3029 ( .A(n2063), .Z(n2041) );
  XOR U3030 ( .A(n2026), .B(n2025), .Z(n2027) );
  XOR U3031 ( .A(x[2]), .B(n2027), .Z(n3421) );
  XOR U3032 ( .A(n3421), .B(n2049), .Z(n2081) );
  XOR U3033 ( .A(n2041), .B(n2081), .Z(n2094) );
  IV U3034 ( .A(x[2]), .Z(n2037) );
  XOR U3035 ( .A(x[4]), .B(n2037), .Z(n2086) );
  NOR U3036 ( .A(n2094), .B(n2086), .Z(n2029) );
  XOR U3037 ( .A(x[7]), .B(n3867), .Z(n3764) );
  XOR U3038 ( .A(n3421), .B(n3764), .Z(n2028) );
  XNOR U3039 ( .A(n2029), .B(n2028), .Z(n2030) );
  XNOR U3040 ( .A(n2109), .B(n3421), .Z(n2093) );
  NOR U3041 ( .A(n2084), .B(n2093), .Z(n2039) );
  XNOR U3042 ( .A(n2030), .B(n2039), .Z(n2051) );
  IV U3043 ( .A(x[1]), .Z(n3866) );
  XNOR U3044 ( .A(n3866), .B(x[2]), .Z(n2031) );
  XNOR U3045 ( .A(n3764), .B(n2031), .Z(n2083) );
  ANDN U3046 ( .B(n2083), .A(x[0]), .Z(n2032) );
  XNOR U3047 ( .A(n2084), .B(n2031), .Z(n2088) );
  NANDN U3048 ( .A(n2041), .B(n2088), .Z(n2042) );
  XOR U3049 ( .A(n2032), .B(n2042), .Z(n2034) );
  OR U3050 ( .A(n2083), .B(n2063), .Z(n2033) );
  NAND U3051 ( .A(n2034), .B(n2033), .Z(n2035) );
  XOR U3052 ( .A(n2051), .B(n2035), .Z(n2036) );
  XOR U3053 ( .A(n2098), .B(n2036), .Z(n2077) );
  XNOR U3054 ( .A(n2041), .B(x[0]), .Z(n2064) );
  XNOR U3055 ( .A(n3867), .B(n2064), .Z(n2111) );
  IV U3056 ( .A(x[7]), .Z(n2040) );
  XOR U3057 ( .A(n2040), .B(n2037), .Z(n2103) );
  NANDN U3058 ( .A(n2111), .B(n2103), .Z(n2038) );
  XOR U3059 ( .A(n2039), .B(n2038), .Z(n2046) );
  XOR U3060 ( .A(n3866), .B(n2040), .Z(n3765) );
  NAND U3061 ( .A(n2081), .B(n3765), .Z(n2050) );
  ANDN U3062 ( .B(n2098), .A(n2109), .Z(n2044) );
  XNOR U3063 ( .A(n2042), .B(n2041), .Z(n2043) );
  XNOR U3064 ( .A(n2044), .B(n2043), .Z(n2045) );
  XNOR U3065 ( .A(n2046), .B(n2045), .Z(n2048) );
  XNOR U3066 ( .A(x[2]), .B(n3764), .Z(n2047) );
  XNOR U3067 ( .A(n2048), .B(n2047), .Z(n2078) );
  IV U3068 ( .A(n2078), .Z(n2070) );
  AND U3069 ( .A(n2073), .B(n2070), .Z(n2066) );
  XOR U3070 ( .A(n2077), .B(n2066), .Z(n2054) );
  ANDN U3071 ( .B(n2049), .A(x[1]), .Z(n2053) );
  XNOR U3072 ( .A(n2051), .B(n2050), .Z(n2052) );
  XNOR U3073 ( .A(n2053), .B(n2052), .Z(n2072) );
  ANDN U3074 ( .B(n2054), .A(n2072), .Z(n2061) );
  IV U3075 ( .A(n2073), .Z(n2058) );
  NANDN U3076 ( .A(n2058), .B(n2072), .Z(n2055) );
  NANDN U3077 ( .A(n2061), .B(n2055), .Z(n2085) );
  NANDN U3078 ( .A(n2073), .B(n2070), .Z(n2056) );
  NAND U3079 ( .A(n2056), .B(n2072), .Z(n2060) );
  XNOR U3080 ( .A(n2070), .B(n2077), .Z(n2057) );
  NANDN U3081 ( .A(n2058), .B(n2057), .Z(n2059) );
  AND U3082 ( .A(n2060), .B(n2059), .Z(n2110) );
  OR U3083 ( .A(n2085), .B(n2110), .Z(n2062) );
  ANDN U3084 ( .B(n2062), .A(n2061), .Z(n2089) );
  NANDN U3085 ( .A(n2089), .B(n2063), .Z(n3863) );
  NANDN U3086 ( .A(n2085), .B(n2064), .Z(n2065) );
  XOR U3087 ( .A(n3863), .B(n2065), .Z(n2097) );
  NANDN U3088 ( .A(n2070), .B(n2077), .Z(n2069) );
  XNOR U3089 ( .A(n2066), .B(n2072), .Z(n2067) );
  NANDN U3090 ( .A(n2077), .B(n2067), .Z(n2068) );
  AND U3091 ( .A(n2069), .B(n2068), .Z(n3869) );
  NANDN U3092 ( .A(n2070), .B(n2073), .Z(n2071) );
  NAND U3093 ( .A(n2077), .B(n2071), .Z(n2076) );
  XNOR U3094 ( .A(n2073), .B(n2072), .Z(n2074) );
  NANDN U3095 ( .A(n2078), .B(n2074), .Z(n2075) );
  NAND U3096 ( .A(n2076), .B(n2075), .Z(n3763) );
  IV U3097 ( .A(n3763), .Z(n3420) );
  NANDN U3098 ( .A(n3869), .B(n3420), .Z(n2080) );
  NANDN U3099 ( .A(n2078), .B(n2077), .Z(n2079) );
  NAND U3100 ( .A(n2080), .B(n2079), .Z(n3766) );
  NANDN U3101 ( .A(n3766), .B(n2081), .Z(n3423) );
  NANDN U3102 ( .A(n3869), .B(n3867), .Z(n2082) );
  XNOR U3103 ( .A(n3423), .B(n2082), .Z(n2099) );
  XOR U3104 ( .A(n2097), .B(n2099), .Z(z[2]) );
  NOR U3105 ( .A(n2085), .B(n2083), .Z(n2091) );
  XOR U3106 ( .A(n3420), .B(n2110), .Z(n2092) );
  NANDN U3107 ( .A(n2084), .B(n2092), .Z(n2105) );
  XOR U3108 ( .A(n2085), .B(n3869), .Z(n2112) );
  XNOR U3109 ( .A(n2092), .B(n2112), .Z(n2095) );
  OR U3110 ( .A(n2086), .B(n2095), .Z(n2087) );
  XNOR U3111 ( .A(n2105), .B(n2087), .Z(n3862) );
  NANDN U3112 ( .A(n2089), .B(n2088), .Z(n2100) );
  XNOR U3113 ( .A(n3862), .B(n2100), .Z(n2090) );
  XOR U3114 ( .A(n2091), .B(n2090), .Z(n3771) );
  NANDN U3115 ( .A(n2093), .B(n2092), .Z(n3424) );
  OR U3116 ( .A(n2095), .B(n2094), .Z(n2096) );
  XOR U3117 ( .A(n3424), .B(n2096), .Z(n2106) );
  XOR U3118 ( .A(n2106), .B(n2097), .Z(n3427) );
  XOR U3119 ( .A(n3771), .B(n3427), .Z(n3927) );
  ANDN U3120 ( .B(n2110), .A(n2098), .Z(n2102) );
  XNOR U3121 ( .A(n2100), .B(n2099), .Z(n2101) );
  XNOR U3122 ( .A(n2102), .B(n2101), .Z(n2108) );
  NAND U3123 ( .A(n2103), .B(n2112), .Z(n2104) );
  XNOR U3124 ( .A(n2105), .B(n2104), .Z(n3767) );
  XOR U3125 ( .A(n2106), .B(n3767), .Z(n2107) );
  XOR U3126 ( .A(n2108), .B(n2107), .Z(n3770) );
  XNOR U3127 ( .A(n3927), .B(n3770), .Z(z[1]) );
  ANDN U3128 ( .B(n2110), .A(n2109), .Z(n3865) );
  ANDN U3129 ( .B(n2112), .A(n2111), .Z(n3426) );
  XNOR U3130 ( .A(n3424), .B(z[1]), .Z(n2113) );
  XNOR U3131 ( .A(n3426), .B(n2113), .Z(n2114) );
  XOR U3132 ( .A(n3863), .B(n2114), .Z(n2115) );
  XOR U3133 ( .A(n3865), .B(n2115), .Z(z[7]) );
  IV U3134 ( .A(x[9]), .Z(n3575) );
  IV U3135 ( .A(x[8]), .Z(n3638) );
  XNOR U3136 ( .A(x[14]), .B(n3638), .Z(n2121) );
  XOR U3137 ( .A(x[13]), .B(n2121), .Z(n3631) );
  ANDN U3138 ( .B(n3575), .A(n3631), .Z(n2118) );
  XNOR U3139 ( .A(x[12]), .B(x[15]), .Z(n3567) );
  XOR U3140 ( .A(x[11]), .B(x[9]), .Z(n2116) );
  XNOR U3141 ( .A(x[10]), .B(n2116), .Z(n2142) );
  XNOR U3142 ( .A(x[14]), .B(n2142), .Z(n3580) );
  NANDN U3143 ( .A(n3567), .B(n3580), .Z(n2120) );
  IV U3144 ( .A(x[12]), .Z(n2123) );
  XOR U3145 ( .A(x[10]), .B(n2123), .Z(n3569) );
  XOR U3146 ( .A(n3638), .B(n2167), .Z(n2171) );
  IV U3147 ( .A(n3631), .Z(n2161) );
  XOR U3148 ( .A(n2171), .B(n2161), .Z(n3625) );
  XNOR U3149 ( .A(n3580), .B(n3625), .Z(n3583) );
  OR U3150 ( .A(n3569), .B(n3583), .Z(n2117) );
  XOR U3151 ( .A(n2120), .B(n2117), .Z(n2137) );
  XNOR U3152 ( .A(n2118), .B(n2137), .Z(n2145) );
  IV U3153 ( .A(x[10]), .Z(n2124) );
  IV U3154 ( .A(x[15]), .Z(n3574) );
  XOR U3155 ( .A(n2124), .B(n3574), .Z(n3646) );
  NAND U3156 ( .A(n3625), .B(n3646), .Z(n2119) );
  XNOR U3157 ( .A(n2120), .B(n2119), .Z(n2128) );
  XOR U3158 ( .A(x[15]), .B(n3631), .Z(n3565) );
  XNOR U3159 ( .A(n2142), .B(n2121), .Z(n3624) );
  NAND U3160 ( .A(n3565), .B(n3624), .Z(n2122) );
  XOR U3161 ( .A(n2128), .B(n2122), .Z(n2148) );
  XNOR U3162 ( .A(n2123), .B(n2161), .Z(n3561) );
  NOR U3163 ( .A(n3638), .B(n3561), .Z(n2130) );
  XNOR U3164 ( .A(n2124), .B(x[9]), .Z(n2131) );
  XOR U3165 ( .A(n3567), .B(n2131), .Z(n3558) );
  NANDN U3166 ( .A(n3558), .B(n2167), .Z(n2132) );
  XNOR U3167 ( .A(n2132), .B(n3565), .Z(n2126) );
  XNOR U3168 ( .A(n2124), .B(n2171), .Z(n2125) );
  XNOR U3169 ( .A(n2126), .B(n2125), .Z(n2127) );
  XOR U3170 ( .A(n2128), .B(n2127), .Z(n2129) );
  XNOR U3171 ( .A(n2130), .B(n2129), .Z(n2157) );
  IV U3172 ( .A(n2157), .Z(n2147) );
  NANDN U3173 ( .A(n2168), .B(n2147), .Z(n2141) );
  XNOR U3174 ( .A(n2131), .B(n3565), .Z(n3566) );
  ANDN U3175 ( .B(n3566), .A(x[8]), .Z(n2133) );
  XOR U3176 ( .A(n2133), .B(n2132), .Z(n2135) );
  OR U3177 ( .A(n2167), .B(n3566), .Z(n2134) );
  NAND U3178 ( .A(n2135), .B(n2134), .Z(n2136) );
  XOR U3179 ( .A(n3624), .B(n2136), .Z(n2139) );
  XOR U3180 ( .A(n3567), .B(n2137), .Z(n2138) );
  XNOR U3181 ( .A(n2139), .B(n2138), .Z(n2158) );
  IV U3182 ( .A(n2158), .Z(n2154) );
  NANDN U3183 ( .A(n2154), .B(n2168), .Z(n2140) );
  NAND U3184 ( .A(n2141), .B(n2140), .Z(n2150) );
  XOR U3185 ( .A(x[13]), .B(n2142), .Z(n2153) );
  NANDN U3186 ( .A(n2153), .B(n3575), .Z(n2144) );
  NANDN U3187 ( .A(n3574), .B(n2153), .Z(n2143) );
  AND U3188 ( .A(n2144), .B(n2143), .Z(n2149) );
  XOR U3189 ( .A(n2149), .B(n2145), .Z(n2166) );
  IV U3190 ( .A(n2166), .Z(n2151) );
  ANDN U3191 ( .B(n2151), .A(n2154), .Z(n2146) );
  XOR U3192 ( .A(n2150), .B(n2146), .Z(n2164) );
  OR U3193 ( .A(n2164), .B(n2147), .Z(n3564) );
  XOR U3194 ( .A(n2149), .B(n2148), .Z(n2163) );
  NANDN U3195 ( .A(n2157), .B(n2163), .Z(n2156) );
  XNOR U3196 ( .A(n2151), .B(n2150), .Z(n2152) );
  XNOR U3197 ( .A(n2156), .B(n2152), .Z(n2165) );
  ANDN U3198 ( .B(n2154), .A(n2165), .Z(n2160) );
  XOR U3199 ( .A(n3564), .B(n2160), .Z(n3577) );
  OR U3200 ( .A(n3577), .B(n2153), .Z(n3628) );
  ANDN U3201 ( .B(n2154), .A(n2166), .Z(n2155) );
  XNOR U3202 ( .A(n2156), .B(n2155), .Z(n2169) );
  XNOR U3203 ( .A(n2158), .B(n2157), .Z(n2159) );
  NANDN U3204 ( .A(n2169), .B(n2159), .Z(n3563) );
  XOR U3205 ( .A(n3563), .B(n2160), .Z(n3633) );
  OR U3206 ( .A(n3633), .B(n2161), .Z(n2162) );
  XNOR U3207 ( .A(n3628), .B(n2162), .Z(n3585) );
  OR U3208 ( .A(n2164), .B(n2163), .Z(n3559) );
  NOR U3209 ( .A(n2166), .B(n2165), .Z(n2170) );
  XOR U3210 ( .A(n3559), .B(n2170), .Z(n3557) );
  ANDN U3211 ( .B(n2167), .A(n3557), .Z(n3640) );
  OR U3212 ( .A(n2169), .B(n2168), .Z(n3560) );
  XOR U3213 ( .A(n3560), .B(n2170), .Z(n3568) );
  OR U3214 ( .A(n3568), .B(n2171), .Z(n2172) );
  XOR U3215 ( .A(n3640), .B(n2172), .Z(n3650) );
  XNOR U3216 ( .A(n3585), .B(n3650), .Z(z[10]) );
  IV U3217 ( .A(x[20]), .Z(n2173) );
  IV U3218 ( .A(x[16]), .Z(n2258) );
  XOR U3219 ( .A(n2258), .B(x[22]), .Z(n2174) );
  XOR U3220 ( .A(n2174), .B(x[21]), .Z(n2198) );
  IV U3221 ( .A(n2198), .Z(n3682) );
  XOR U3222 ( .A(n2173), .B(n3682), .Z(n2247) );
  XOR U3223 ( .A(x[17]), .B(x[19]), .Z(n2175) );
  XOR U3224 ( .A(x[23]), .B(n2173), .Z(n2233) );
  XNOR U3225 ( .A(n2175), .B(n2233), .Z(n2212) );
  IV U3226 ( .A(n2212), .Z(n2190) );
  XOR U3227 ( .A(n2175), .B(n2174), .Z(n2176) );
  XOR U3228 ( .A(x[18]), .B(n2176), .Z(n3659) );
  XOR U3229 ( .A(n3659), .B(n2198), .Z(n2230) );
  XOR U3230 ( .A(n2190), .B(n2230), .Z(n2243) );
  IV U3231 ( .A(x[18]), .Z(n2186) );
  XOR U3232 ( .A(x[20]), .B(n2186), .Z(n2235) );
  NOR U3233 ( .A(n2243), .B(n2235), .Z(n2178) );
  XOR U3234 ( .A(x[23]), .B(n3682), .Z(n3667) );
  XOR U3235 ( .A(n3659), .B(n3667), .Z(n2177) );
  XNOR U3236 ( .A(n2178), .B(n2177), .Z(n2179) );
  XNOR U3237 ( .A(n2258), .B(n3659), .Z(n2242) );
  NOR U3238 ( .A(n2233), .B(n2242), .Z(n2188) );
  XNOR U3239 ( .A(n2179), .B(n2188), .Z(n2200) );
  IV U3240 ( .A(x[17]), .Z(n3681) );
  XNOR U3241 ( .A(n3681), .B(x[18]), .Z(n2180) );
  XNOR U3242 ( .A(n3667), .B(n2180), .Z(n2232) );
  ANDN U3243 ( .B(n2232), .A(x[16]), .Z(n2181) );
  XNOR U3244 ( .A(n2233), .B(n2180), .Z(n2237) );
  NANDN U3245 ( .A(n2190), .B(n2237), .Z(n2191) );
  XOR U3246 ( .A(n2181), .B(n2191), .Z(n2183) );
  OR U3247 ( .A(n2232), .B(n2212), .Z(n2182) );
  NAND U3248 ( .A(n2183), .B(n2182), .Z(n2184) );
  XOR U3249 ( .A(n2200), .B(n2184), .Z(n2185) );
  XOR U3250 ( .A(n2247), .B(n2185), .Z(n2226) );
  XNOR U3251 ( .A(n2190), .B(x[16]), .Z(n2213) );
  XNOR U3252 ( .A(n3682), .B(n2213), .Z(n2260) );
  IV U3253 ( .A(x[23]), .Z(n2189) );
  XOR U3254 ( .A(n2189), .B(n2186), .Z(n2252) );
  NANDN U3255 ( .A(n2260), .B(n2252), .Z(n2187) );
  XOR U3256 ( .A(n2188), .B(n2187), .Z(n2195) );
  XOR U3257 ( .A(n3681), .B(n2189), .Z(n3668) );
  NAND U3258 ( .A(n2230), .B(n3668), .Z(n2199) );
  ANDN U3259 ( .B(n2247), .A(n2258), .Z(n2193) );
  XNOR U3260 ( .A(n2191), .B(n2190), .Z(n2192) );
  XNOR U3261 ( .A(n2193), .B(n2192), .Z(n2194) );
  XNOR U3262 ( .A(n2195), .B(n2194), .Z(n2197) );
  XNOR U3263 ( .A(x[18]), .B(n3667), .Z(n2196) );
  XNOR U3264 ( .A(n2197), .B(n2196), .Z(n2227) );
  IV U3265 ( .A(n2227), .Z(n2219) );
  AND U3266 ( .A(n2222), .B(n2219), .Z(n2215) );
  XOR U3267 ( .A(n2226), .B(n2215), .Z(n2203) );
  ANDN U3268 ( .B(n2198), .A(x[17]), .Z(n2202) );
  XNOR U3269 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U3270 ( .A(n2202), .B(n2201), .Z(n2221) );
  ANDN U3271 ( .B(n2203), .A(n2221), .Z(n2210) );
  IV U3272 ( .A(n2222), .Z(n2207) );
  NANDN U3273 ( .A(n2207), .B(n2221), .Z(n2204) );
  NANDN U3274 ( .A(n2210), .B(n2204), .Z(n2234) );
  NANDN U3275 ( .A(n2222), .B(n2219), .Z(n2205) );
  NAND U3276 ( .A(n2205), .B(n2221), .Z(n2209) );
  XNOR U3277 ( .A(n2219), .B(n2226), .Z(n2206) );
  NANDN U3278 ( .A(n2207), .B(n2206), .Z(n2208) );
  AND U3279 ( .A(n2209), .B(n2208), .Z(n2259) );
  OR U3280 ( .A(n2234), .B(n2259), .Z(n2211) );
  ANDN U3281 ( .B(n2211), .A(n2210), .Z(n2238) );
  NANDN U3282 ( .A(n2238), .B(n2212), .Z(n3678) );
  NANDN U3283 ( .A(n2234), .B(n2213), .Z(n2214) );
  XOR U3284 ( .A(n3678), .B(n2214), .Z(n2246) );
  NANDN U3285 ( .A(n2219), .B(n2226), .Z(n2218) );
  XNOR U3286 ( .A(n2215), .B(n2221), .Z(n2216) );
  NANDN U3287 ( .A(n2226), .B(n2216), .Z(n2217) );
  AND U3288 ( .A(n2218), .B(n2217), .Z(n3684) );
  NANDN U3289 ( .A(n2219), .B(n2222), .Z(n2220) );
  NAND U3290 ( .A(n2226), .B(n2220), .Z(n2225) );
  XNOR U3291 ( .A(n2222), .B(n2221), .Z(n2223) );
  NANDN U3292 ( .A(n2227), .B(n2223), .Z(n2224) );
  NAND U3293 ( .A(n2225), .B(n2224), .Z(n3666) );
  IV U3294 ( .A(n3666), .Z(n3658) );
  NANDN U3295 ( .A(n3684), .B(n3658), .Z(n2229) );
  NANDN U3296 ( .A(n2227), .B(n2226), .Z(n2228) );
  NAND U3297 ( .A(n2229), .B(n2228), .Z(n3669) );
  NANDN U3298 ( .A(n3669), .B(n2230), .Z(n3661) );
  NANDN U3299 ( .A(n3684), .B(n3682), .Z(n2231) );
  XNOR U3300 ( .A(n3661), .B(n2231), .Z(n2248) );
  XOR U3301 ( .A(n2246), .B(n2248), .Z(z[18]) );
  NOR U3302 ( .A(n2234), .B(n2232), .Z(n2240) );
  XOR U3303 ( .A(n3658), .B(n2259), .Z(n2241) );
  NANDN U3304 ( .A(n2233), .B(n2241), .Z(n2254) );
  XOR U3305 ( .A(n2234), .B(n3684), .Z(n2261) );
  XNOR U3306 ( .A(n2241), .B(n2261), .Z(n2244) );
  OR U3307 ( .A(n2235), .B(n2244), .Z(n2236) );
  XNOR U3308 ( .A(n2254), .B(n2236), .Z(n3677) );
  NANDN U3309 ( .A(n2238), .B(n2237), .Z(n2249) );
  XNOR U3310 ( .A(n3677), .B(n2249), .Z(n2239) );
  XOR U3311 ( .A(n2240), .B(n2239), .Z(n3674) );
  NANDN U3312 ( .A(n2242), .B(n2241), .Z(n3662) );
  OR U3313 ( .A(n2244), .B(n2243), .Z(n2245) );
  XOR U3314 ( .A(n3662), .B(n2245), .Z(n2255) );
  XOR U3315 ( .A(n2255), .B(n2246), .Z(n3665) );
  XOR U3316 ( .A(n3674), .B(n3665), .Z(n3692) );
  ANDN U3317 ( .B(n2259), .A(n2247), .Z(n2251) );
  XNOR U3318 ( .A(n2249), .B(n2248), .Z(n2250) );
  XNOR U3319 ( .A(n2251), .B(n2250), .Z(n2257) );
  NAND U3320 ( .A(n2252), .B(n2261), .Z(n2253) );
  XNOR U3321 ( .A(n2254), .B(n2253), .Z(n3670) );
  XOR U3322 ( .A(n2255), .B(n3670), .Z(n2256) );
  XOR U3323 ( .A(n2257), .B(n2256), .Z(n3673) );
  XNOR U3324 ( .A(n3692), .B(n3673), .Z(z[17]) );
  ANDN U3325 ( .B(n2259), .A(n2258), .Z(n3680) );
  ANDN U3326 ( .B(n2261), .A(n2260), .Z(n3664) );
  XNOR U3327 ( .A(n3662), .B(z[17]), .Z(n2262) );
  XNOR U3328 ( .A(n3664), .B(n2262), .Z(n2263) );
  XOR U3329 ( .A(n3678), .B(n2263), .Z(n2264) );
  XOR U3330 ( .A(n3680), .B(n2264), .Z(z[23]) );
  IV U3331 ( .A(x[28]), .Z(n2265) );
  IV U3332 ( .A(x[24]), .Z(n2350) );
  XOR U3333 ( .A(n2350), .B(x[30]), .Z(n2266) );
  XOR U3334 ( .A(n2266), .B(x[29]), .Z(n2290) );
  IV U3335 ( .A(n2290), .Z(n3717) );
  XOR U3336 ( .A(n2265), .B(n3717), .Z(n2339) );
  XOR U3337 ( .A(x[25]), .B(x[27]), .Z(n2267) );
  XOR U3338 ( .A(x[31]), .B(n2265), .Z(n2325) );
  XNOR U3339 ( .A(n2267), .B(n2325), .Z(n2304) );
  IV U3340 ( .A(n2304), .Z(n2282) );
  XOR U3341 ( .A(n2267), .B(n2266), .Z(n2268) );
  XOR U3342 ( .A(x[26]), .B(n2268), .Z(n3694) );
  XOR U3343 ( .A(n3694), .B(n2290), .Z(n2322) );
  XOR U3344 ( .A(n2282), .B(n2322), .Z(n2335) );
  IV U3345 ( .A(x[26]), .Z(n2278) );
  XOR U3346 ( .A(x[28]), .B(n2278), .Z(n2327) );
  NOR U3347 ( .A(n2335), .B(n2327), .Z(n2270) );
  XOR U3348 ( .A(x[31]), .B(n3717), .Z(n3702) );
  XOR U3349 ( .A(n3694), .B(n3702), .Z(n2269) );
  XNOR U3350 ( .A(n2270), .B(n2269), .Z(n2271) );
  XNOR U3351 ( .A(n2350), .B(n3694), .Z(n2334) );
  NOR U3352 ( .A(n2325), .B(n2334), .Z(n2280) );
  XNOR U3353 ( .A(n2271), .B(n2280), .Z(n2292) );
  IV U3354 ( .A(x[25]), .Z(n3716) );
  XNOR U3355 ( .A(n3716), .B(x[26]), .Z(n2272) );
  XNOR U3356 ( .A(n3702), .B(n2272), .Z(n2324) );
  ANDN U3357 ( .B(n2324), .A(x[24]), .Z(n2273) );
  XNOR U3358 ( .A(n2325), .B(n2272), .Z(n2329) );
  NANDN U3359 ( .A(n2282), .B(n2329), .Z(n2283) );
  XOR U3360 ( .A(n2273), .B(n2283), .Z(n2275) );
  OR U3361 ( .A(n2324), .B(n2304), .Z(n2274) );
  NAND U3362 ( .A(n2275), .B(n2274), .Z(n2276) );
  XOR U3363 ( .A(n2292), .B(n2276), .Z(n2277) );
  XOR U3364 ( .A(n2339), .B(n2277), .Z(n2318) );
  XNOR U3365 ( .A(n2282), .B(x[24]), .Z(n2305) );
  XNOR U3366 ( .A(n3717), .B(n2305), .Z(n2352) );
  IV U3367 ( .A(x[31]), .Z(n2281) );
  XOR U3368 ( .A(n2281), .B(n2278), .Z(n2344) );
  NANDN U3369 ( .A(n2352), .B(n2344), .Z(n2279) );
  XOR U3370 ( .A(n2280), .B(n2279), .Z(n2287) );
  XOR U3371 ( .A(n3716), .B(n2281), .Z(n3703) );
  NAND U3372 ( .A(n2322), .B(n3703), .Z(n2291) );
  ANDN U3373 ( .B(n2339), .A(n2350), .Z(n2285) );
  XNOR U3374 ( .A(n2283), .B(n2282), .Z(n2284) );
  XNOR U3375 ( .A(n2285), .B(n2284), .Z(n2286) );
  XNOR U3376 ( .A(n2287), .B(n2286), .Z(n2289) );
  XNOR U3377 ( .A(x[26]), .B(n3702), .Z(n2288) );
  XNOR U3378 ( .A(n2289), .B(n2288), .Z(n2319) );
  IV U3379 ( .A(n2319), .Z(n2311) );
  AND U3380 ( .A(n2314), .B(n2311), .Z(n2307) );
  XOR U3381 ( .A(n2318), .B(n2307), .Z(n2295) );
  ANDN U3382 ( .B(n2290), .A(x[25]), .Z(n2294) );
  XNOR U3383 ( .A(n2292), .B(n2291), .Z(n2293) );
  XNOR U3384 ( .A(n2294), .B(n2293), .Z(n2313) );
  ANDN U3385 ( .B(n2295), .A(n2313), .Z(n2302) );
  IV U3386 ( .A(n2314), .Z(n2299) );
  NANDN U3387 ( .A(n2299), .B(n2313), .Z(n2296) );
  NANDN U3388 ( .A(n2302), .B(n2296), .Z(n2326) );
  NANDN U3389 ( .A(n2314), .B(n2311), .Z(n2297) );
  NAND U3390 ( .A(n2297), .B(n2313), .Z(n2301) );
  XNOR U3391 ( .A(n2311), .B(n2318), .Z(n2298) );
  NANDN U3392 ( .A(n2299), .B(n2298), .Z(n2300) );
  AND U3393 ( .A(n2301), .B(n2300), .Z(n2351) );
  OR U3394 ( .A(n2326), .B(n2351), .Z(n2303) );
  ANDN U3395 ( .B(n2303), .A(n2302), .Z(n2330) );
  NANDN U3396 ( .A(n2330), .B(n2304), .Z(n3713) );
  NANDN U3397 ( .A(n2326), .B(n2305), .Z(n2306) );
  XOR U3398 ( .A(n3713), .B(n2306), .Z(n2338) );
  NANDN U3399 ( .A(n2311), .B(n2318), .Z(n2310) );
  XNOR U3400 ( .A(n2307), .B(n2313), .Z(n2308) );
  NANDN U3401 ( .A(n2318), .B(n2308), .Z(n2309) );
  AND U3402 ( .A(n2310), .B(n2309), .Z(n3719) );
  NANDN U3403 ( .A(n2311), .B(n2314), .Z(n2312) );
  NAND U3404 ( .A(n2318), .B(n2312), .Z(n2317) );
  XNOR U3405 ( .A(n2314), .B(n2313), .Z(n2315) );
  NANDN U3406 ( .A(n2319), .B(n2315), .Z(n2316) );
  NAND U3407 ( .A(n2317), .B(n2316), .Z(n3701) );
  IV U3408 ( .A(n3701), .Z(n3693) );
  NANDN U3409 ( .A(n3719), .B(n3693), .Z(n2321) );
  NANDN U3410 ( .A(n2319), .B(n2318), .Z(n2320) );
  NAND U3411 ( .A(n2321), .B(n2320), .Z(n3704) );
  NANDN U3412 ( .A(n3704), .B(n2322), .Z(n3696) );
  NANDN U3413 ( .A(n3719), .B(n3717), .Z(n2323) );
  XNOR U3414 ( .A(n3696), .B(n2323), .Z(n2340) );
  XOR U3415 ( .A(n2338), .B(n2340), .Z(z[26]) );
  NOR U3416 ( .A(n2326), .B(n2324), .Z(n2332) );
  XOR U3417 ( .A(n3693), .B(n2351), .Z(n2333) );
  NANDN U3418 ( .A(n2325), .B(n2333), .Z(n2346) );
  XOR U3419 ( .A(n2326), .B(n3719), .Z(n2353) );
  XNOR U3420 ( .A(n2333), .B(n2353), .Z(n2336) );
  OR U3421 ( .A(n2327), .B(n2336), .Z(n2328) );
  XNOR U3422 ( .A(n2346), .B(n2328), .Z(n3712) );
  NANDN U3423 ( .A(n2330), .B(n2329), .Z(n2341) );
  XNOR U3424 ( .A(n3712), .B(n2341), .Z(n2331) );
  XOR U3425 ( .A(n2332), .B(n2331), .Z(n3709) );
  NANDN U3426 ( .A(n2334), .B(n2333), .Z(n3697) );
  OR U3427 ( .A(n2336), .B(n2335), .Z(n2337) );
  XOR U3428 ( .A(n3697), .B(n2337), .Z(n2347) );
  XOR U3429 ( .A(n2347), .B(n2338), .Z(n3700) );
  XOR U3430 ( .A(n3709), .B(n3700), .Z(n3727) );
  ANDN U3431 ( .B(n2351), .A(n2339), .Z(n2343) );
  XNOR U3432 ( .A(n2341), .B(n2340), .Z(n2342) );
  XNOR U3433 ( .A(n2343), .B(n2342), .Z(n2349) );
  NAND U3434 ( .A(n2344), .B(n2353), .Z(n2345) );
  XNOR U3435 ( .A(n2346), .B(n2345), .Z(n3705) );
  XOR U3436 ( .A(n2347), .B(n3705), .Z(n2348) );
  XOR U3437 ( .A(n2349), .B(n2348), .Z(n3708) );
  XNOR U3438 ( .A(n3727), .B(n3708), .Z(z[25]) );
  ANDN U3439 ( .B(n2351), .A(n2350), .Z(n3715) );
  ANDN U3440 ( .B(n2353), .A(n2352), .Z(n3699) );
  XNOR U3441 ( .A(n3697), .B(z[25]), .Z(n2354) );
  XNOR U3442 ( .A(n3699), .B(n2354), .Z(n2355) );
  XOR U3443 ( .A(n3713), .B(n2355), .Z(n2356) );
  XOR U3444 ( .A(n3715), .B(n2356), .Z(z[31]) );
  IV U3445 ( .A(x[36]), .Z(n2357) );
  IV U3446 ( .A(x[32]), .Z(n2442) );
  XOR U3447 ( .A(n2442), .B(x[38]), .Z(n2358) );
  XOR U3448 ( .A(n2358), .B(x[37]), .Z(n2382) );
  IV U3449 ( .A(n2382), .Z(n3752) );
  XOR U3450 ( .A(n2357), .B(n3752), .Z(n2431) );
  XOR U3451 ( .A(x[33]), .B(x[35]), .Z(n2359) );
  XOR U3452 ( .A(x[39]), .B(n2357), .Z(n2417) );
  XNOR U3453 ( .A(n2359), .B(n2417), .Z(n2396) );
  IV U3454 ( .A(n2396), .Z(n2374) );
  XOR U3455 ( .A(n2359), .B(n2358), .Z(n2360) );
  XOR U3456 ( .A(x[34]), .B(n2360), .Z(n3729) );
  XOR U3457 ( .A(n3729), .B(n2382), .Z(n2414) );
  XOR U3458 ( .A(n2374), .B(n2414), .Z(n2427) );
  IV U3459 ( .A(x[34]), .Z(n2370) );
  XOR U3460 ( .A(x[36]), .B(n2370), .Z(n2419) );
  NOR U3461 ( .A(n2427), .B(n2419), .Z(n2362) );
  XOR U3462 ( .A(x[39]), .B(n3752), .Z(n3737) );
  XOR U3463 ( .A(n3729), .B(n3737), .Z(n2361) );
  XNOR U3464 ( .A(n2362), .B(n2361), .Z(n2363) );
  XNOR U3465 ( .A(n2442), .B(n3729), .Z(n2426) );
  NOR U3466 ( .A(n2417), .B(n2426), .Z(n2372) );
  XNOR U3467 ( .A(n2363), .B(n2372), .Z(n2384) );
  IV U3468 ( .A(x[33]), .Z(n3751) );
  XNOR U3469 ( .A(n3751), .B(x[34]), .Z(n2364) );
  XNOR U3470 ( .A(n3737), .B(n2364), .Z(n2416) );
  ANDN U3471 ( .B(n2416), .A(x[32]), .Z(n2365) );
  XNOR U3472 ( .A(n2417), .B(n2364), .Z(n2421) );
  NANDN U3473 ( .A(n2374), .B(n2421), .Z(n2375) );
  XOR U3474 ( .A(n2365), .B(n2375), .Z(n2367) );
  OR U3475 ( .A(n2416), .B(n2396), .Z(n2366) );
  NAND U3476 ( .A(n2367), .B(n2366), .Z(n2368) );
  XOR U3477 ( .A(n2384), .B(n2368), .Z(n2369) );
  XOR U3478 ( .A(n2431), .B(n2369), .Z(n2410) );
  XNOR U3479 ( .A(n2374), .B(x[32]), .Z(n2397) );
  XNOR U3480 ( .A(n3752), .B(n2397), .Z(n2444) );
  IV U3481 ( .A(x[39]), .Z(n2373) );
  XOR U3482 ( .A(n2373), .B(n2370), .Z(n2436) );
  NANDN U3483 ( .A(n2444), .B(n2436), .Z(n2371) );
  XOR U3484 ( .A(n2372), .B(n2371), .Z(n2379) );
  XOR U3485 ( .A(n3751), .B(n2373), .Z(n3738) );
  NAND U3486 ( .A(n2414), .B(n3738), .Z(n2383) );
  ANDN U3487 ( .B(n2431), .A(n2442), .Z(n2377) );
  XNOR U3488 ( .A(n2375), .B(n2374), .Z(n2376) );
  XNOR U3489 ( .A(n2377), .B(n2376), .Z(n2378) );
  XNOR U3490 ( .A(n2379), .B(n2378), .Z(n2381) );
  XNOR U3491 ( .A(x[34]), .B(n3737), .Z(n2380) );
  XNOR U3492 ( .A(n2381), .B(n2380), .Z(n2411) );
  IV U3493 ( .A(n2411), .Z(n2403) );
  AND U3494 ( .A(n2406), .B(n2403), .Z(n2399) );
  XOR U3495 ( .A(n2410), .B(n2399), .Z(n2387) );
  ANDN U3496 ( .B(n2382), .A(x[33]), .Z(n2386) );
  XNOR U3497 ( .A(n2384), .B(n2383), .Z(n2385) );
  XNOR U3498 ( .A(n2386), .B(n2385), .Z(n2405) );
  ANDN U3499 ( .B(n2387), .A(n2405), .Z(n2394) );
  IV U3500 ( .A(n2406), .Z(n2391) );
  NANDN U3501 ( .A(n2391), .B(n2405), .Z(n2388) );
  NANDN U3502 ( .A(n2394), .B(n2388), .Z(n2418) );
  NANDN U3503 ( .A(n2406), .B(n2403), .Z(n2389) );
  NAND U3504 ( .A(n2389), .B(n2405), .Z(n2393) );
  XNOR U3505 ( .A(n2403), .B(n2410), .Z(n2390) );
  NANDN U3506 ( .A(n2391), .B(n2390), .Z(n2392) );
  AND U3507 ( .A(n2393), .B(n2392), .Z(n2443) );
  OR U3508 ( .A(n2418), .B(n2443), .Z(n2395) );
  ANDN U3509 ( .B(n2395), .A(n2394), .Z(n2422) );
  NANDN U3510 ( .A(n2422), .B(n2396), .Z(n3748) );
  NANDN U3511 ( .A(n2418), .B(n2397), .Z(n2398) );
  XOR U3512 ( .A(n3748), .B(n2398), .Z(n2430) );
  NANDN U3513 ( .A(n2403), .B(n2410), .Z(n2402) );
  XNOR U3514 ( .A(n2399), .B(n2405), .Z(n2400) );
  NANDN U3515 ( .A(n2410), .B(n2400), .Z(n2401) );
  AND U3516 ( .A(n2402), .B(n2401), .Z(n3754) );
  NANDN U3517 ( .A(n2403), .B(n2406), .Z(n2404) );
  NAND U3518 ( .A(n2410), .B(n2404), .Z(n2409) );
  XNOR U3519 ( .A(n2406), .B(n2405), .Z(n2407) );
  NANDN U3520 ( .A(n2411), .B(n2407), .Z(n2408) );
  NAND U3521 ( .A(n2409), .B(n2408), .Z(n3736) );
  IV U3522 ( .A(n3736), .Z(n3728) );
  NANDN U3523 ( .A(n3754), .B(n3728), .Z(n2413) );
  NANDN U3524 ( .A(n2411), .B(n2410), .Z(n2412) );
  NAND U3525 ( .A(n2413), .B(n2412), .Z(n3739) );
  NANDN U3526 ( .A(n3739), .B(n2414), .Z(n3731) );
  NANDN U3527 ( .A(n3754), .B(n3752), .Z(n2415) );
  XNOR U3528 ( .A(n3731), .B(n2415), .Z(n2432) );
  XOR U3529 ( .A(n2430), .B(n2432), .Z(z[34]) );
  NOR U3530 ( .A(n2418), .B(n2416), .Z(n2424) );
  XOR U3531 ( .A(n3728), .B(n2443), .Z(n2425) );
  NANDN U3532 ( .A(n2417), .B(n2425), .Z(n2438) );
  XOR U3533 ( .A(n2418), .B(n3754), .Z(n2445) );
  XNOR U3534 ( .A(n2425), .B(n2445), .Z(n2428) );
  OR U3535 ( .A(n2419), .B(n2428), .Z(n2420) );
  XNOR U3536 ( .A(n2438), .B(n2420), .Z(n3747) );
  NANDN U3537 ( .A(n2422), .B(n2421), .Z(n2433) );
  XNOR U3538 ( .A(n3747), .B(n2433), .Z(n2423) );
  XOR U3539 ( .A(n2424), .B(n2423), .Z(n3744) );
  NANDN U3540 ( .A(n2426), .B(n2425), .Z(n3732) );
  OR U3541 ( .A(n2428), .B(n2427), .Z(n2429) );
  XOR U3542 ( .A(n3732), .B(n2429), .Z(n2439) );
  XOR U3543 ( .A(n2439), .B(n2430), .Z(n3735) );
  XOR U3544 ( .A(n3744), .B(n3735), .Z(n3762) );
  ANDN U3545 ( .B(n2443), .A(n2431), .Z(n2435) );
  XNOR U3546 ( .A(n2433), .B(n2432), .Z(n2434) );
  XNOR U3547 ( .A(n2435), .B(n2434), .Z(n2441) );
  NAND U3548 ( .A(n2436), .B(n2445), .Z(n2437) );
  XNOR U3549 ( .A(n2438), .B(n2437), .Z(n3740) );
  XOR U3550 ( .A(n2439), .B(n3740), .Z(n2440) );
  XOR U3551 ( .A(n2441), .B(n2440), .Z(n3743) );
  XNOR U3552 ( .A(n3762), .B(n3743), .Z(z[33]) );
  ANDN U3553 ( .B(n2443), .A(n2442), .Z(n3750) );
  ANDN U3554 ( .B(n2445), .A(n2444), .Z(n3734) );
  XNOR U3555 ( .A(n3732), .B(z[33]), .Z(n2446) );
  XNOR U3556 ( .A(n3734), .B(n2446), .Z(n2447) );
  XOR U3557 ( .A(n3748), .B(n2447), .Z(n2448) );
  XOR U3558 ( .A(n3750), .B(n2448), .Z(z[39]) );
  IV U3559 ( .A(x[44]), .Z(n2449) );
  IV U3560 ( .A(x[40]), .Z(n2534) );
  XOR U3561 ( .A(n2534), .B(x[46]), .Z(n2450) );
  XOR U3562 ( .A(n2450), .B(x[45]), .Z(n2474) );
  IV U3563 ( .A(n2474), .Z(n3797) );
  XOR U3564 ( .A(n2449), .B(n3797), .Z(n2523) );
  XOR U3565 ( .A(x[41]), .B(x[43]), .Z(n2451) );
  XOR U3566 ( .A(x[47]), .B(n2449), .Z(n2509) );
  XNOR U3567 ( .A(n2451), .B(n2509), .Z(n2488) );
  IV U3568 ( .A(n2488), .Z(n2466) );
  XOR U3569 ( .A(n2451), .B(n2450), .Z(n2452) );
  XOR U3570 ( .A(x[42]), .B(n2452), .Z(n3774) );
  XOR U3571 ( .A(n3774), .B(n2474), .Z(n2506) );
  XOR U3572 ( .A(n2466), .B(n2506), .Z(n2519) );
  IV U3573 ( .A(x[42]), .Z(n2462) );
  XOR U3574 ( .A(x[44]), .B(n2462), .Z(n2511) );
  NOR U3575 ( .A(n2519), .B(n2511), .Z(n2454) );
  XOR U3576 ( .A(x[47]), .B(n3797), .Z(n3782) );
  XOR U3577 ( .A(n3774), .B(n3782), .Z(n2453) );
  XNOR U3578 ( .A(n2454), .B(n2453), .Z(n2455) );
  XNOR U3579 ( .A(n2534), .B(n3774), .Z(n2518) );
  NOR U3580 ( .A(n2509), .B(n2518), .Z(n2464) );
  XNOR U3581 ( .A(n2455), .B(n2464), .Z(n2476) );
  IV U3582 ( .A(x[41]), .Z(n3796) );
  XNOR U3583 ( .A(n3796), .B(x[42]), .Z(n2456) );
  XNOR U3584 ( .A(n3782), .B(n2456), .Z(n2508) );
  ANDN U3585 ( .B(n2508), .A(x[40]), .Z(n2457) );
  XNOR U3586 ( .A(n2509), .B(n2456), .Z(n2513) );
  NANDN U3587 ( .A(n2466), .B(n2513), .Z(n2467) );
  XOR U3588 ( .A(n2457), .B(n2467), .Z(n2459) );
  OR U3589 ( .A(n2508), .B(n2488), .Z(n2458) );
  NAND U3590 ( .A(n2459), .B(n2458), .Z(n2460) );
  XOR U3591 ( .A(n2476), .B(n2460), .Z(n2461) );
  XOR U3592 ( .A(n2523), .B(n2461), .Z(n2502) );
  XNOR U3593 ( .A(n2466), .B(x[40]), .Z(n2489) );
  XNOR U3594 ( .A(n3797), .B(n2489), .Z(n2536) );
  IV U3595 ( .A(x[47]), .Z(n2465) );
  XOR U3596 ( .A(n2465), .B(n2462), .Z(n2528) );
  NANDN U3597 ( .A(n2536), .B(n2528), .Z(n2463) );
  XOR U3598 ( .A(n2464), .B(n2463), .Z(n2471) );
  XOR U3599 ( .A(n3796), .B(n2465), .Z(n3783) );
  NAND U3600 ( .A(n2506), .B(n3783), .Z(n2475) );
  ANDN U3601 ( .B(n2523), .A(n2534), .Z(n2469) );
  XNOR U3602 ( .A(n2467), .B(n2466), .Z(n2468) );
  XNOR U3603 ( .A(n2469), .B(n2468), .Z(n2470) );
  XNOR U3604 ( .A(n2471), .B(n2470), .Z(n2473) );
  XNOR U3605 ( .A(x[42]), .B(n3782), .Z(n2472) );
  XNOR U3606 ( .A(n2473), .B(n2472), .Z(n2503) );
  IV U3607 ( .A(n2503), .Z(n2495) );
  AND U3608 ( .A(n2498), .B(n2495), .Z(n2491) );
  XOR U3609 ( .A(n2502), .B(n2491), .Z(n2479) );
  ANDN U3610 ( .B(n2474), .A(x[41]), .Z(n2478) );
  XNOR U3611 ( .A(n2476), .B(n2475), .Z(n2477) );
  XNOR U3612 ( .A(n2478), .B(n2477), .Z(n2497) );
  ANDN U3613 ( .B(n2479), .A(n2497), .Z(n2486) );
  IV U3614 ( .A(n2498), .Z(n2483) );
  NANDN U3615 ( .A(n2483), .B(n2497), .Z(n2480) );
  NANDN U3616 ( .A(n2486), .B(n2480), .Z(n2510) );
  NANDN U3617 ( .A(n2498), .B(n2495), .Z(n2481) );
  NAND U3618 ( .A(n2481), .B(n2497), .Z(n2485) );
  XNOR U3619 ( .A(n2495), .B(n2502), .Z(n2482) );
  NANDN U3620 ( .A(n2483), .B(n2482), .Z(n2484) );
  AND U3621 ( .A(n2485), .B(n2484), .Z(n2535) );
  OR U3622 ( .A(n2510), .B(n2535), .Z(n2487) );
  ANDN U3623 ( .B(n2487), .A(n2486), .Z(n2514) );
  NANDN U3624 ( .A(n2514), .B(n2488), .Z(n3793) );
  NANDN U3625 ( .A(n2510), .B(n2489), .Z(n2490) );
  XOR U3626 ( .A(n3793), .B(n2490), .Z(n2522) );
  NANDN U3627 ( .A(n2495), .B(n2502), .Z(n2494) );
  XNOR U3628 ( .A(n2491), .B(n2497), .Z(n2492) );
  NANDN U3629 ( .A(n2502), .B(n2492), .Z(n2493) );
  AND U3630 ( .A(n2494), .B(n2493), .Z(n3799) );
  NANDN U3631 ( .A(n2495), .B(n2498), .Z(n2496) );
  NAND U3632 ( .A(n2502), .B(n2496), .Z(n2501) );
  XNOR U3633 ( .A(n2498), .B(n2497), .Z(n2499) );
  NANDN U3634 ( .A(n2503), .B(n2499), .Z(n2500) );
  NAND U3635 ( .A(n2501), .B(n2500), .Z(n3781) );
  IV U3636 ( .A(n3781), .Z(n3773) );
  NANDN U3637 ( .A(n3799), .B(n3773), .Z(n2505) );
  NANDN U3638 ( .A(n2503), .B(n2502), .Z(n2504) );
  NAND U3639 ( .A(n2505), .B(n2504), .Z(n3784) );
  NANDN U3640 ( .A(n3784), .B(n2506), .Z(n3776) );
  NANDN U3641 ( .A(n3799), .B(n3797), .Z(n2507) );
  XNOR U3642 ( .A(n3776), .B(n2507), .Z(n2524) );
  XOR U3643 ( .A(n2522), .B(n2524), .Z(z[42]) );
  NOR U3644 ( .A(n2510), .B(n2508), .Z(n2516) );
  XOR U3645 ( .A(n3773), .B(n2535), .Z(n2517) );
  NANDN U3646 ( .A(n2509), .B(n2517), .Z(n2530) );
  XOR U3647 ( .A(n2510), .B(n3799), .Z(n2537) );
  XNOR U3648 ( .A(n2517), .B(n2537), .Z(n2520) );
  OR U3649 ( .A(n2511), .B(n2520), .Z(n2512) );
  XNOR U3650 ( .A(n2530), .B(n2512), .Z(n3792) );
  NANDN U3651 ( .A(n2514), .B(n2513), .Z(n2525) );
  XNOR U3652 ( .A(n3792), .B(n2525), .Z(n2515) );
  XOR U3653 ( .A(n2516), .B(n2515), .Z(n3789) );
  NANDN U3654 ( .A(n2518), .B(n2517), .Z(n3777) );
  OR U3655 ( .A(n2520), .B(n2519), .Z(n2521) );
  XOR U3656 ( .A(n3777), .B(n2521), .Z(n2531) );
  XOR U3657 ( .A(n2531), .B(n2522), .Z(n3780) );
  XOR U3658 ( .A(n3789), .B(n3780), .Z(n3807) );
  ANDN U3659 ( .B(n2535), .A(n2523), .Z(n2527) );
  XNOR U3660 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3661 ( .A(n2527), .B(n2526), .Z(n2533) );
  NAND U3662 ( .A(n2528), .B(n2537), .Z(n2529) );
  XNOR U3663 ( .A(n2530), .B(n2529), .Z(n3785) );
  XOR U3664 ( .A(n2531), .B(n3785), .Z(n2532) );
  XOR U3665 ( .A(n2533), .B(n2532), .Z(n3788) );
  XNOR U3666 ( .A(n3807), .B(n3788), .Z(z[41]) );
  ANDN U3667 ( .B(n2535), .A(n2534), .Z(n3795) );
  ANDN U3668 ( .B(n2537), .A(n2536), .Z(n3779) );
  XNOR U3669 ( .A(n3777), .B(z[41]), .Z(n2538) );
  XNOR U3670 ( .A(n3779), .B(n2538), .Z(n2539) );
  XOR U3671 ( .A(n3793), .B(n2539), .Z(n2540) );
  XOR U3672 ( .A(n3795), .B(n2540), .Z(z[47]) );
  IV U3673 ( .A(x[52]), .Z(n2541) );
  IV U3674 ( .A(x[48]), .Z(n2626) );
  XOR U3675 ( .A(n2626), .B(x[54]), .Z(n2542) );
  XOR U3676 ( .A(n2542), .B(x[53]), .Z(n2566) );
  IV U3677 ( .A(n2566), .Z(n3833) );
  XOR U3678 ( .A(n2541), .B(n3833), .Z(n2615) );
  XOR U3679 ( .A(x[49]), .B(x[51]), .Z(n2543) );
  XOR U3680 ( .A(x[55]), .B(n2541), .Z(n2601) );
  XNOR U3681 ( .A(n2543), .B(n2601), .Z(n2580) );
  IV U3682 ( .A(n2580), .Z(n2558) );
  XOR U3683 ( .A(n2543), .B(n2542), .Z(n2544) );
  XOR U3684 ( .A(x[50]), .B(n2544), .Z(n3809) );
  XOR U3685 ( .A(n3809), .B(n2566), .Z(n2598) );
  XOR U3686 ( .A(n2558), .B(n2598), .Z(n2611) );
  IV U3687 ( .A(x[50]), .Z(n2554) );
  XOR U3688 ( .A(x[52]), .B(n2554), .Z(n2603) );
  NOR U3689 ( .A(n2611), .B(n2603), .Z(n2546) );
  XOR U3690 ( .A(x[55]), .B(n3833), .Z(n3818) );
  XOR U3691 ( .A(n3809), .B(n3818), .Z(n2545) );
  XNOR U3692 ( .A(n2546), .B(n2545), .Z(n2547) );
  XNOR U3693 ( .A(n2626), .B(n3809), .Z(n2610) );
  NOR U3694 ( .A(n2601), .B(n2610), .Z(n2556) );
  XNOR U3695 ( .A(n2547), .B(n2556), .Z(n2568) );
  IV U3696 ( .A(x[49]), .Z(n3832) );
  XNOR U3697 ( .A(n3832), .B(x[50]), .Z(n2548) );
  XNOR U3698 ( .A(n3818), .B(n2548), .Z(n2600) );
  ANDN U3699 ( .B(n2600), .A(x[48]), .Z(n2549) );
  XNOR U3700 ( .A(n2601), .B(n2548), .Z(n2605) );
  NANDN U3701 ( .A(n2558), .B(n2605), .Z(n2559) );
  XOR U3702 ( .A(n2549), .B(n2559), .Z(n2551) );
  OR U3703 ( .A(n2600), .B(n2580), .Z(n2550) );
  NAND U3704 ( .A(n2551), .B(n2550), .Z(n2552) );
  XOR U3705 ( .A(n2568), .B(n2552), .Z(n2553) );
  XOR U3706 ( .A(n2615), .B(n2553), .Z(n2594) );
  XNOR U3707 ( .A(n2558), .B(x[48]), .Z(n2581) );
  XNOR U3708 ( .A(n3833), .B(n2581), .Z(n2628) );
  IV U3709 ( .A(x[55]), .Z(n2557) );
  XOR U3710 ( .A(n2557), .B(n2554), .Z(n2620) );
  NANDN U3711 ( .A(n2628), .B(n2620), .Z(n2555) );
  XOR U3712 ( .A(n2556), .B(n2555), .Z(n2563) );
  XOR U3713 ( .A(n3832), .B(n2557), .Z(n3819) );
  NAND U3714 ( .A(n2598), .B(n3819), .Z(n2567) );
  ANDN U3715 ( .B(n2615), .A(n2626), .Z(n2561) );
  XNOR U3716 ( .A(n2559), .B(n2558), .Z(n2560) );
  XNOR U3717 ( .A(n2561), .B(n2560), .Z(n2562) );
  XNOR U3718 ( .A(n2563), .B(n2562), .Z(n2565) );
  XNOR U3719 ( .A(x[50]), .B(n3818), .Z(n2564) );
  XNOR U3720 ( .A(n2565), .B(n2564), .Z(n2595) );
  IV U3721 ( .A(n2595), .Z(n2587) );
  AND U3722 ( .A(n2590), .B(n2587), .Z(n2583) );
  XOR U3723 ( .A(n2594), .B(n2583), .Z(n2571) );
  ANDN U3724 ( .B(n2566), .A(x[49]), .Z(n2570) );
  XNOR U3725 ( .A(n2568), .B(n2567), .Z(n2569) );
  XNOR U3726 ( .A(n2570), .B(n2569), .Z(n2589) );
  ANDN U3727 ( .B(n2571), .A(n2589), .Z(n2578) );
  IV U3728 ( .A(n2590), .Z(n2575) );
  NANDN U3729 ( .A(n2575), .B(n2589), .Z(n2572) );
  NANDN U3730 ( .A(n2578), .B(n2572), .Z(n2602) );
  NANDN U3731 ( .A(n2590), .B(n2587), .Z(n2573) );
  NAND U3732 ( .A(n2573), .B(n2589), .Z(n2577) );
  XNOR U3733 ( .A(n2587), .B(n2594), .Z(n2574) );
  NANDN U3734 ( .A(n2575), .B(n2574), .Z(n2576) );
  AND U3735 ( .A(n2577), .B(n2576), .Z(n2627) );
  OR U3736 ( .A(n2602), .B(n2627), .Z(n2579) );
  ANDN U3737 ( .B(n2579), .A(n2578), .Z(n2606) );
  NANDN U3738 ( .A(n2606), .B(n2580), .Z(n3829) );
  NANDN U3739 ( .A(n2602), .B(n2581), .Z(n2582) );
  XOR U3740 ( .A(n3829), .B(n2582), .Z(n2614) );
  NANDN U3741 ( .A(n2587), .B(n2594), .Z(n2586) );
  XNOR U3742 ( .A(n2583), .B(n2589), .Z(n2584) );
  NANDN U3743 ( .A(n2594), .B(n2584), .Z(n2585) );
  AND U3744 ( .A(n2586), .B(n2585), .Z(n3835) );
  NANDN U3745 ( .A(n2587), .B(n2590), .Z(n2588) );
  NAND U3746 ( .A(n2594), .B(n2588), .Z(n2593) );
  XNOR U3747 ( .A(n2590), .B(n2589), .Z(n2591) );
  NANDN U3748 ( .A(n2595), .B(n2591), .Z(n2592) );
  NAND U3749 ( .A(n2593), .B(n2592), .Z(n3817) );
  IV U3750 ( .A(n3817), .Z(n3808) );
  NANDN U3751 ( .A(n3835), .B(n3808), .Z(n2597) );
  NANDN U3752 ( .A(n2595), .B(n2594), .Z(n2596) );
  NAND U3753 ( .A(n2597), .B(n2596), .Z(n3820) );
  NANDN U3754 ( .A(n3820), .B(n2598), .Z(n3811) );
  NANDN U3755 ( .A(n3835), .B(n3833), .Z(n2599) );
  XNOR U3756 ( .A(n3811), .B(n2599), .Z(n2616) );
  XOR U3757 ( .A(n2614), .B(n2616), .Z(z[50]) );
  NOR U3758 ( .A(n2602), .B(n2600), .Z(n2608) );
  XOR U3759 ( .A(n3808), .B(n2627), .Z(n2609) );
  NANDN U3760 ( .A(n2601), .B(n2609), .Z(n2622) );
  XOR U3761 ( .A(n2602), .B(n3835), .Z(n2629) );
  XNOR U3762 ( .A(n2609), .B(n2629), .Z(n2612) );
  OR U3763 ( .A(n2603), .B(n2612), .Z(n2604) );
  XNOR U3764 ( .A(n2622), .B(n2604), .Z(n3828) );
  NANDN U3765 ( .A(n2606), .B(n2605), .Z(n2617) );
  XNOR U3766 ( .A(n3828), .B(n2617), .Z(n2607) );
  XOR U3767 ( .A(n2608), .B(n2607), .Z(n3825) );
  NANDN U3768 ( .A(n2610), .B(n2609), .Z(n3812) );
  OR U3769 ( .A(n2612), .B(n2611), .Z(n2613) );
  XOR U3770 ( .A(n3812), .B(n2613), .Z(n2623) );
  XOR U3771 ( .A(n2623), .B(n2614), .Z(n3815) );
  XOR U3772 ( .A(n3825), .B(n3815), .Z(n3843) );
  ANDN U3773 ( .B(n2627), .A(n2615), .Z(n2619) );
  XNOR U3774 ( .A(n2617), .B(n2616), .Z(n2618) );
  XNOR U3775 ( .A(n2619), .B(n2618), .Z(n2625) );
  NAND U3776 ( .A(n2620), .B(n2629), .Z(n2621) );
  XNOR U3777 ( .A(n2622), .B(n2621), .Z(n3821) );
  XOR U3778 ( .A(n2623), .B(n3821), .Z(n2624) );
  XOR U3779 ( .A(n2625), .B(n2624), .Z(n3824) );
  XNOR U3780 ( .A(n3843), .B(n3824), .Z(z[49]) );
  ANDN U3781 ( .B(n2627), .A(n2626), .Z(n3831) );
  ANDN U3782 ( .B(n2629), .A(n2628), .Z(n3814) );
  XNOR U3783 ( .A(n3812), .B(z[49]), .Z(n2630) );
  XNOR U3784 ( .A(n3814), .B(n2630), .Z(n2631) );
  XOR U3785 ( .A(n3829), .B(n2631), .Z(n2632) );
  XOR U3786 ( .A(n3831), .B(n2632), .Z(z[55]) );
  IV U3787 ( .A(x[60]), .Z(n2633) );
  IV U3788 ( .A(x[56]), .Z(n2718) );
  XOR U3789 ( .A(n2718), .B(x[62]), .Z(n2634) );
  XOR U3790 ( .A(n2634), .B(x[61]), .Z(n2658) );
  IV U3791 ( .A(n2658), .Z(n3882) );
  XOR U3792 ( .A(n2633), .B(n3882), .Z(n2707) );
  XOR U3793 ( .A(x[57]), .B(x[59]), .Z(n2635) );
  XOR U3794 ( .A(x[63]), .B(n2633), .Z(n2693) );
  XNOR U3795 ( .A(n2635), .B(n2693), .Z(n2672) );
  IV U3796 ( .A(n2672), .Z(n2650) );
  XOR U3797 ( .A(n2635), .B(n2634), .Z(n2636) );
  XOR U3798 ( .A(x[58]), .B(n2636), .Z(n3845) );
  XOR U3799 ( .A(n3845), .B(n2658), .Z(n2690) );
  XOR U3800 ( .A(n2650), .B(n2690), .Z(n2703) );
  IV U3801 ( .A(x[58]), .Z(n2646) );
  XOR U3802 ( .A(x[60]), .B(n2646), .Z(n2695) );
  NOR U3803 ( .A(n2703), .B(n2695), .Z(n2638) );
  XOR U3804 ( .A(x[63]), .B(n3882), .Z(n3853) );
  XOR U3805 ( .A(n3845), .B(n3853), .Z(n2637) );
  XNOR U3806 ( .A(n2638), .B(n2637), .Z(n2639) );
  XNOR U3807 ( .A(n2718), .B(n3845), .Z(n2702) );
  NOR U3808 ( .A(n2693), .B(n2702), .Z(n2648) );
  XNOR U3809 ( .A(n2639), .B(n2648), .Z(n2660) );
  IV U3810 ( .A(x[57]), .Z(n3881) );
  XNOR U3811 ( .A(n3881), .B(x[58]), .Z(n2640) );
  XNOR U3812 ( .A(n3853), .B(n2640), .Z(n2692) );
  ANDN U3813 ( .B(n2692), .A(x[56]), .Z(n2641) );
  XNOR U3814 ( .A(n2693), .B(n2640), .Z(n2697) );
  NANDN U3815 ( .A(n2650), .B(n2697), .Z(n2651) );
  XOR U3816 ( .A(n2641), .B(n2651), .Z(n2643) );
  OR U3817 ( .A(n2692), .B(n2672), .Z(n2642) );
  NAND U3818 ( .A(n2643), .B(n2642), .Z(n2644) );
  XOR U3819 ( .A(n2660), .B(n2644), .Z(n2645) );
  XOR U3820 ( .A(n2707), .B(n2645), .Z(n2686) );
  XNOR U3821 ( .A(n2650), .B(x[56]), .Z(n2673) );
  XNOR U3822 ( .A(n3882), .B(n2673), .Z(n2720) );
  IV U3823 ( .A(x[63]), .Z(n2649) );
  XOR U3824 ( .A(n2649), .B(n2646), .Z(n2712) );
  NANDN U3825 ( .A(n2720), .B(n2712), .Z(n2647) );
  XOR U3826 ( .A(n2648), .B(n2647), .Z(n2655) );
  XOR U3827 ( .A(n3881), .B(n2649), .Z(n3854) );
  NAND U3828 ( .A(n2690), .B(n3854), .Z(n2659) );
  ANDN U3829 ( .B(n2707), .A(n2718), .Z(n2653) );
  XNOR U3830 ( .A(n2651), .B(n2650), .Z(n2652) );
  XNOR U3831 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3832 ( .A(n2655), .B(n2654), .Z(n2657) );
  XNOR U3833 ( .A(x[58]), .B(n3853), .Z(n2656) );
  XNOR U3834 ( .A(n2657), .B(n2656), .Z(n2687) );
  IV U3835 ( .A(n2687), .Z(n2679) );
  AND U3836 ( .A(n2682), .B(n2679), .Z(n2675) );
  XOR U3837 ( .A(n2686), .B(n2675), .Z(n2663) );
  ANDN U3838 ( .B(n2658), .A(x[57]), .Z(n2662) );
  XNOR U3839 ( .A(n2660), .B(n2659), .Z(n2661) );
  XNOR U3840 ( .A(n2662), .B(n2661), .Z(n2681) );
  ANDN U3841 ( .B(n2663), .A(n2681), .Z(n2670) );
  IV U3842 ( .A(n2682), .Z(n2667) );
  NANDN U3843 ( .A(n2667), .B(n2681), .Z(n2664) );
  NANDN U3844 ( .A(n2670), .B(n2664), .Z(n2694) );
  NANDN U3845 ( .A(n2682), .B(n2679), .Z(n2665) );
  NAND U3846 ( .A(n2665), .B(n2681), .Z(n2669) );
  XNOR U3847 ( .A(n2679), .B(n2686), .Z(n2666) );
  NANDN U3848 ( .A(n2667), .B(n2666), .Z(n2668) );
  AND U3849 ( .A(n2669), .B(n2668), .Z(n2719) );
  OR U3850 ( .A(n2694), .B(n2719), .Z(n2671) );
  ANDN U3851 ( .B(n2671), .A(n2670), .Z(n2698) );
  NANDN U3852 ( .A(n2698), .B(n2672), .Z(n3878) );
  NANDN U3853 ( .A(n2694), .B(n2673), .Z(n2674) );
  XOR U3854 ( .A(n3878), .B(n2674), .Z(n2706) );
  NANDN U3855 ( .A(n2679), .B(n2686), .Z(n2678) );
  XNOR U3856 ( .A(n2675), .B(n2681), .Z(n2676) );
  NANDN U3857 ( .A(n2686), .B(n2676), .Z(n2677) );
  AND U3858 ( .A(n2678), .B(n2677), .Z(n3884) );
  NANDN U3859 ( .A(n2679), .B(n2682), .Z(n2680) );
  NAND U3860 ( .A(n2686), .B(n2680), .Z(n2685) );
  XNOR U3861 ( .A(n2682), .B(n2681), .Z(n2683) );
  NANDN U3862 ( .A(n2687), .B(n2683), .Z(n2684) );
  NAND U3863 ( .A(n2685), .B(n2684), .Z(n3852) );
  IV U3864 ( .A(n3852), .Z(n3844) );
  NANDN U3865 ( .A(n3884), .B(n3844), .Z(n2689) );
  NANDN U3866 ( .A(n2687), .B(n2686), .Z(n2688) );
  NAND U3867 ( .A(n2689), .B(n2688), .Z(n3855) );
  NANDN U3868 ( .A(n3855), .B(n2690), .Z(n3847) );
  NANDN U3869 ( .A(n3884), .B(n3882), .Z(n2691) );
  XNOR U3870 ( .A(n3847), .B(n2691), .Z(n2708) );
  XOR U3871 ( .A(n2706), .B(n2708), .Z(z[58]) );
  NOR U3872 ( .A(n2694), .B(n2692), .Z(n2700) );
  XOR U3873 ( .A(n3844), .B(n2719), .Z(n2701) );
  NANDN U3874 ( .A(n2693), .B(n2701), .Z(n2714) );
  XOR U3875 ( .A(n2694), .B(n3884), .Z(n2721) );
  XNOR U3876 ( .A(n2701), .B(n2721), .Z(n2704) );
  OR U3877 ( .A(n2695), .B(n2704), .Z(n2696) );
  XNOR U3878 ( .A(n2714), .B(n2696), .Z(n3877) );
  NANDN U3879 ( .A(n2698), .B(n2697), .Z(n2709) );
  XNOR U3880 ( .A(n3877), .B(n2709), .Z(n2699) );
  XOR U3881 ( .A(n2700), .B(n2699), .Z(n3860) );
  NANDN U3882 ( .A(n2702), .B(n2701), .Z(n3848) );
  OR U3883 ( .A(n2704), .B(n2703), .Z(n2705) );
  XOR U3884 ( .A(n3848), .B(n2705), .Z(n2715) );
  XOR U3885 ( .A(n2715), .B(n2706), .Z(n3851) );
  XOR U3886 ( .A(n3860), .B(n3851), .Z(n3892) );
  ANDN U3887 ( .B(n2719), .A(n2707), .Z(n2711) );
  XNOR U3888 ( .A(n2709), .B(n2708), .Z(n2710) );
  XNOR U3889 ( .A(n2711), .B(n2710), .Z(n2717) );
  NAND U3890 ( .A(n2712), .B(n2721), .Z(n2713) );
  XNOR U3891 ( .A(n2714), .B(n2713), .Z(n3856) );
  XOR U3892 ( .A(n2715), .B(n3856), .Z(n2716) );
  XOR U3893 ( .A(n2717), .B(n2716), .Z(n3859) );
  XNOR U3894 ( .A(n3892), .B(n3859), .Z(z[57]) );
  ANDN U3895 ( .B(n2719), .A(n2718), .Z(n3880) );
  ANDN U3896 ( .B(n2721), .A(n2720), .Z(n3850) );
  XNOR U3897 ( .A(n3848), .B(z[57]), .Z(n2722) );
  XNOR U3898 ( .A(n3850), .B(n2722), .Z(n2723) );
  XOR U3899 ( .A(n3878), .B(n2723), .Z(n2724) );
  XOR U3900 ( .A(n3880), .B(n2724), .Z(z[63]) );
  IV U3901 ( .A(x[68]), .Z(n2725) );
  IV U3902 ( .A(x[64]), .Z(n2810) );
  XOR U3903 ( .A(n2810), .B(x[70]), .Z(n2726) );
  XOR U3904 ( .A(n2726), .B(x[69]), .Z(n2750) );
  IV U3905 ( .A(n2750), .Z(n3917) );
  XOR U3906 ( .A(n2725), .B(n3917), .Z(n2799) );
  XOR U3907 ( .A(x[65]), .B(x[67]), .Z(n2727) );
  XOR U3908 ( .A(x[71]), .B(n2725), .Z(n2785) );
  XNOR U3909 ( .A(n2727), .B(n2785), .Z(n2764) );
  IV U3910 ( .A(n2764), .Z(n2742) );
  XOR U3911 ( .A(n2727), .B(n2726), .Z(n2728) );
  XOR U3912 ( .A(x[66]), .B(n2728), .Z(n3894) );
  XOR U3913 ( .A(n3894), .B(n2750), .Z(n2782) );
  XOR U3914 ( .A(n2742), .B(n2782), .Z(n2795) );
  IV U3915 ( .A(x[66]), .Z(n2738) );
  XOR U3916 ( .A(x[68]), .B(n2738), .Z(n2787) );
  NOR U3917 ( .A(n2795), .B(n2787), .Z(n2730) );
  XOR U3918 ( .A(x[71]), .B(n3917), .Z(n3902) );
  XOR U3919 ( .A(n3894), .B(n3902), .Z(n2729) );
  XNOR U3920 ( .A(n2730), .B(n2729), .Z(n2731) );
  XNOR U3921 ( .A(n2810), .B(n3894), .Z(n2794) );
  NOR U3922 ( .A(n2785), .B(n2794), .Z(n2740) );
  XNOR U3923 ( .A(n2731), .B(n2740), .Z(n2752) );
  IV U3924 ( .A(x[65]), .Z(n3916) );
  XNOR U3925 ( .A(n3916), .B(x[66]), .Z(n2732) );
  XNOR U3926 ( .A(n3902), .B(n2732), .Z(n2784) );
  ANDN U3927 ( .B(n2784), .A(x[64]), .Z(n2733) );
  XNOR U3928 ( .A(n2785), .B(n2732), .Z(n2789) );
  NANDN U3929 ( .A(n2742), .B(n2789), .Z(n2743) );
  XOR U3930 ( .A(n2733), .B(n2743), .Z(n2735) );
  OR U3931 ( .A(n2784), .B(n2764), .Z(n2734) );
  NAND U3932 ( .A(n2735), .B(n2734), .Z(n2736) );
  XOR U3933 ( .A(n2752), .B(n2736), .Z(n2737) );
  XOR U3934 ( .A(n2799), .B(n2737), .Z(n2778) );
  XNOR U3935 ( .A(n2742), .B(x[64]), .Z(n2765) );
  XNOR U3936 ( .A(n3917), .B(n2765), .Z(n2812) );
  IV U3937 ( .A(x[71]), .Z(n2741) );
  XOR U3938 ( .A(n2741), .B(n2738), .Z(n2804) );
  NANDN U3939 ( .A(n2812), .B(n2804), .Z(n2739) );
  XOR U3940 ( .A(n2740), .B(n2739), .Z(n2747) );
  XOR U3941 ( .A(n3916), .B(n2741), .Z(n3903) );
  NAND U3942 ( .A(n2782), .B(n3903), .Z(n2751) );
  ANDN U3943 ( .B(n2799), .A(n2810), .Z(n2745) );
  XNOR U3944 ( .A(n2743), .B(n2742), .Z(n2744) );
  XNOR U3945 ( .A(n2745), .B(n2744), .Z(n2746) );
  XNOR U3946 ( .A(n2747), .B(n2746), .Z(n2749) );
  XNOR U3947 ( .A(x[66]), .B(n3902), .Z(n2748) );
  XNOR U3948 ( .A(n2749), .B(n2748), .Z(n2779) );
  IV U3949 ( .A(n2779), .Z(n2771) );
  AND U3950 ( .A(n2774), .B(n2771), .Z(n2767) );
  XOR U3951 ( .A(n2778), .B(n2767), .Z(n2755) );
  ANDN U3952 ( .B(n2750), .A(x[65]), .Z(n2754) );
  XNOR U3953 ( .A(n2752), .B(n2751), .Z(n2753) );
  XNOR U3954 ( .A(n2754), .B(n2753), .Z(n2773) );
  ANDN U3955 ( .B(n2755), .A(n2773), .Z(n2762) );
  IV U3956 ( .A(n2774), .Z(n2759) );
  NANDN U3957 ( .A(n2759), .B(n2773), .Z(n2756) );
  NANDN U3958 ( .A(n2762), .B(n2756), .Z(n2786) );
  NANDN U3959 ( .A(n2774), .B(n2771), .Z(n2757) );
  NAND U3960 ( .A(n2757), .B(n2773), .Z(n2761) );
  XNOR U3961 ( .A(n2771), .B(n2778), .Z(n2758) );
  NANDN U3962 ( .A(n2759), .B(n2758), .Z(n2760) );
  AND U3963 ( .A(n2761), .B(n2760), .Z(n2811) );
  OR U3964 ( .A(n2786), .B(n2811), .Z(n2763) );
  ANDN U3965 ( .B(n2763), .A(n2762), .Z(n2790) );
  NANDN U3966 ( .A(n2790), .B(n2764), .Z(n3913) );
  NANDN U3967 ( .A(n2786), .B(n2765), .Z(n2766) );
  XOR U3968 ( .A(n3913), .B(n2766), .Z(n2798) );
  NANDN U3969 ( .A(n2771), .B(n2778), .Z(n2770) );
  XNOR U3970 ( .A(n2767), .B(n2773), .Z(n2768) );
  NANDN U3971 ( .A(n2778), .B(n2768), .Z(n2769) );
  AND U3972 ( .A(n2770), .B(n2769), .Z(n3919) );
  NANDN U3973 ( .A(n2771), .B(n2774), .Z(n2772) );
  NAND U3974 ( .A(n2778), .B(n2772), .Z(n2777) );
  XNOR U3975 ( .A(n2774), .B(n2773), .Z(n2775) );
  NANDN U3976 ( .A(n2779), .B(n2775), .Z(n2776) );
  NAND U3977 ( .A(n2777), .B(n2776), .Z(n3901) );
  IV U3978 ( .A(n3901), .Z(n3893) );
  NANDN U3979 ( .A(n3919), .B(n3893), .Z(n2781) );
  NANDN U3980 ( .A(n2779), .B(n2778), .Z(n2780) );
  NAND U3981 ( .A(n2781), .B(n2780), .Z(n3904) );
  NANDN U3982 ( .A(n3904), .B(n2782), .Z(n3896) );
  NANDN U3983 ( .A(n3919), .B(n3917), .Z(n2783) );
  XNOR U3984 ( .A(n3896), .B(n2783), .Z(n2800) );
  XOR U3985 ( .A(n2798), .B(n2800), .Z(z[66]) );
  NOR U3986 ( .A(n2786), .B(n2784), .Z(n2792) );
  XOR U3987 ( .A(n3893), .B(n2811), .Z(n2793) );
  NANDN U3988 ( .A(n2785), .B(n2793), .Z(n2806) );
  XOR U3989 ( .A(n2786), .B(n3919), .Z(n2813) );
  XNOR U3990 ( .A(n2793), .B(n2813), .Z(n2796) );
  OR U3991 ( .A(n2787), .B(n2796), .Z(n2788) );
  XNOR U3992 ( .A(n2806), .B(n2788), .Z(n3912) );
  NANDN U3993 ( .A(n2790), .B(n2789), .Z(n2801) );
  XNOR U3994 ( .A(n3912), .B(n2801), .Z(n2791) );
  XOR U3995 ( .A(n2792), .B(n2791), .Z(n3909) );
  NANDN U3996 ( .A(n2794), .B(n2793), .Z(n3897) );
  OR U3997 ( .A(n2796), .B(n2795), .Z(n2797) );
  XOR U3998 ( .A(n3897), .B(n2797), .Z(n2807) );
  XOR U3999 ( .A(n2807), .B(n2798), .Z(n3900) );
  XOR U4000 ( .A(n3909), .B(n3900), .Z(n3929) );
  ANDN U4001 ( .B(n2811), .A(n2799), .Z(n2803) );
  XNOR U4002 ( .A(n2801), .B(n2800), .Z(n2802) );
  XNOR U4003 ( .A(n2803), .B(n2802), .Z(n2809) );
  NAND U4004 ( .A(n2804), .B(n2813), .Z(n2805) );
  XNOR U4005 ( .A(n2806), .B(n2805), .Z(n3905) );
  XOR U4006 ( .A(n2807), .B(n3905), .Z(n2808) );
  XOR U4007 ( .A(n2809), .B(n2808), .Z(n3908) );
  XNOR U4008 ( .A(n3929), .B(n3908), .Z(z[65]) );
  ANDN U4009 ( .B(n2811), .A(n2810), .Z(n3915) );
  ANDN U4010 ( .B(n2813), .A(n2812), .Z(n3899) );
  XNOR U4011 ( .A(n3897), .B(z[65]), .Z(n2814) );
  XNOR U4012 ( .A(n3899), .B(n2814), .Z(n2815) );
  XOR U4013 ( .A(n3913), .B(n2815), .Z(n2816) );
  XOR U4014 ( .A(n3915), .B(n2816), .Z(z[71]) );
  IV U4015 ( .A(x[76]), .Z(n2817) );
  IV U4016 ( .A(x[72]), .Z(n2902) );
  XOR U4017 ( .A(n2902), .B(x[78]), .Z(n2818) );
  XOR U4018 ( .A(n2818), .B(x[77]), .Z(n2842) );
  IV U4019 ( .A(n2842), .Z(n3954) );
  XOR U4020 ( .A(n2817), .B(n3954), .Z(n2891) );
  XOR U4021 ( .A(x[73]), .B(x[75]), .Z(n2819) );
  XOR U4022 ( .A(x[79]), .B(n2817), .Z(n2877) );
  XNOR U4023 ( .A(n2819), .B(n2877), .Z(n2856) );
  IV U4024 ( .A(n2856), .Z(n2834) );
  XOR U4025 ( .A(n2819), .B(n2818), .Z(n2820) );
  XOR U4026 ( .A(x[74]), .B(n2820), .Z(n3931) );
  XOR U4027 ( .A(n3931), .B(n2842), .Z(n2874) );
  XOR U4028 ( .A(n2834), .B(n2874), .Z(n2887) );
  IV U4029 ( .A(x[74]), .Z(n2830) );
  XOR U4030 ( .A(x[76]), .B(n2830), .Z(n2879) );
  NOR U4031 ( .A(n2887), .B(n2879), .Z(n2822) );
  XOR U4032 ( .A(x[79]), .B(n3954), .Z(n3939) );
  XOR U4033 ( .A(n3931), .B(n3939), .Z(n2821) );
  XNOR U4034 ( .A(n2822), .B(n2821), .Z(n2823) );
  XNOR U4035 ( .A(n2902), .B(n3931), .Z(n2886) );
  NOR U4036 ( .A(n2877), .B(n2886), .Z(n2832) );
  XNOR U4037 ( .A(n2823), .B(n2832), .Z(n2844) );
  IV U4038 ( .A(x[73]), .Z(n3953) );
  XNOR U4039 ( .A(n3953), .B(x[74]), .Z(n2824) );
  XNOR U4040 ( .A(n3939), .B(n2824), .Z(n2876) );
  ANDN U4041 ( .B(n2876), .A(x[72]), .Z(n2825) );
  XNOR U4042 ( .A(n2877), .B(n2824), .Z(n2881) );
  NANDN U4043 ( .A(n2834), .B(n2881), .Z(n2835) );
  XOR U4044 ( .A(n2825), .B(n2835), .Z(n2827) );
  OR U4045 ( .A(n2876), .B(n2856), .Z(n2826) );
  NAND U4046 ( .A(n2827), .B(n2826), .Z(n2828) );
  XOR U4047 ( .A(n2844), .B(n2828), .Z(n2829) );
  XOR U4048 ( .A(n2891), .B(n2829), .Z(n2870) );
  XNOR U4049 ( .A(n2834), .B(x[72]), .Z(n2857) );
  XNOR U4050 ( .A(n3954), .B(n2857), .Z(n2904) );
  IV U4051 ( .A(x[79]), .Z(n2833) );
  XOR U4052 ( .A(n2833), .B(n2830), .Z(n2896) );
  NANDN U4053 ( .A(n2904), .B(n2896), .Z(n2831) );
  XOR U4054 ( .A(n2832), .B(n2831), .Z(n2839) );
  XOR U4055 ( .A(n3953), .B(n2833), .Z(n3940) );
  NAND U4056 ( .A(n2874), .B(n3940), .Z(n2843) );
  ANDN U4057 ( .B(n2891), .A(n2902), .Z(n2837) );
  XNOR U4058 ( .A(n2835), .B(n2834), .Z(n2836) );
  XNOR U4059 ( .A(n2837), .B(n2836), .Z(n2838) );
  XNOR U4060 ( .A(n2839), .B(n2838), .Z(n2841) );
  XNOR U4061 ( .A(x[74]), .B(n3939), .Z(n2840) );
  XNOR U4062 ( .A(n2841), .B(n2840), .Z(n2871) );
  IV U4063 ( .A(n2871), .Z(n2863) );
  AND U4064 ( .A(n2866), .B(n2863), .Z(n2859) );
  XOR U4065 ( .A(n2870), .B(n2859), .Z(n2847) );
  ANDN U4066 ( .B(n2842), .A(x[73]), .Z(n2846) );
  XNOR U4067 ( .A(n2844), .B(n2843), .Z(n2845) );
  XNOR U4068 ( .A(n2846), .B(n2845), .Z(n2865) );
  ANDN U4069 ( .B(n2847), .A(n2865), .Z(n2854) );
  IV U4070 ( .A(n2866), .Z(n2851) );
  NANDN U4071 ( .A(n2851), .B(n2865), .Z(n2848) );
  NANDN U4072 ( .A(n2854), .B(n2848), .Z(n2878) );
  NANDN U4073 ( .A(n2866), .B(n2863), .Z(n2849) );
  NAND U4074 ( .A(n2849), .B(n2865), .Z(n2853) );
  XNOR U4075 ( .A(n2863), .B(n2870), .Z(n2850) );
  NANDN U4076 ( .A(n2851), .B(n2850), .Z(n2852) );
  AND U4077 ( .A(n2853), .B(n2852), .Z(n2903) );
  OR U4078 ( .A(n2878), .B(n2903), .Z(n2855) );
  ANDN U4079 ( .B(n2855), .A(n2854), .Z(n2882) );
  NANDN U4080 ( .A(n2882), .B(n2856), .Z(n3950) );
  NANDN U4081 ( .A(n2878), .B(n2857), .Z(n2858) );
  XOR U4082 ( .A(n3950), .B(n2858), .Z(n2890) );
  NANDN U4083 ( .A(n2863), .B(n2870), .Z(n2862) );
  XNOR U4084 ( .A(n2859), .B(n2865), .Z(n2860) );
  NANDN U4085 ( .A(n2870), .B(n2860), .Z(n2861) );
  AND U4086 ( .A(n2862), .B(n2861), .Z(n3956) );
  NANDN U4087 ( .A(n2863), .B(n2866), .Z(n2864) );
  NAND U4088 ( .A(n2870), .B(n2864), .Z(n2869) );
  XNOR U4089 ( .A(n2866), .B(n2865), .Z(n2867) );
  NANDN U4090 ( .A(n2871), .B(n2867), .Z(n2868) );
  NAND U4091 ( .A(n2869), .B(n2868), .Z(n3938) );
  IV U4092 ( .A(n3938), .Z(n3930) );
  NANDN U4093 ( .A(n3956), .B(n3930), .Z(n2873) );
  NANDN U4094 ( .A(n2871), .B(n2870), .Z(n2872) );
  NAND U4095 ( .A(n2873), .B(n2872), .Z(n3941) );
  NANDN U4096 ( .A(n3941), .B(n2874), .Z(n3933) );
  NANDN U4097 ( .A(n3956), .B(n3954), .Z(n2875) );
  XNOR U4098 ( .A(n3933), .B(n2875), .Z(n2892) );
  XOR U4099 ( .A(n2890), .B(n2892), .Z(z[74]) );
  NOR U4100 ( .A(n2878), .B(n2876), .Z(n2884) );
  XOR U4101 ( .A(n3930), .B(n2903), .Z(n2885) );
  NANDN U4102 ( .A(n2877), .B(n2885), .Z(n2898) );
  XOR U4103 ( .A(n2878), .B(n3956), .Z(n2905) );
  XNOR U4104 ( .A(n2885), .B(n2905), .Z(n2888) );
  OR U4105 ( .A(n2879), .B(n2888), .Z(n2880) );
  XNOR U4106 ( .A(n2898), .B(n2880), .Z(n3949) );
  NANDN U4107 ( .A(n2882), .B(n2881), .Z(n2893) );
  XNOR U4108 ( .A(n3949), .B(n2893), .Z(n2883) );
  XOR U4109 ( .A(n2884), .B(n2883), .Z(n3946) );
  NANDN U4110 ( .A(n2886), .B(n2885), .Z(n3934) );
  OR U4111 ( .A(n2888), .B(n2887), .Z(n2889) );
  XOR U4112 ( .A(n3934), .B(n2889), .Z(n2899) );
  XOR U4113 ( .A(n2899), .B(n2890), .Z(n3937) );
  XOR U4114 ( .A(n3946), .B(n3937), .Z(n3964) );
  ANDN U4115 ( .B(n2903), .A(n2891), .Z(n2895) );
  XNOR U4116 ( .A(n2893), .B(n2892), .Z(n2894) );
  XNOR U4117 ( .A(n2895), .B(n2894), .Z(n2901) );
  NAND U4118 ( .A(n2896), .B(n2905), .Z(n2897) );
  XNOR U4119 ( .A(n2898), .B(n2897), .Z(n3942) );
  XOR U4120 ( .A(n2899), .B(n3942), .Z(n2900) );
  XOR U4121 ( .A(n2901), .B(n2900), .Z(n3945) );
  XNOR U4122 ( .A(n3964), .B(n3945), .Z(z[73]) );
  ANDN U4123 ( .B(n2903), .A(n2902), .Z(n3952) );
  ANDN U4124 ( .B(n2905), .A(n2904), .Z(n3936) );
  XNOR U4125 ( .A(n3934), .B(z[73]), .Z(n2906) );
  XNOR U4126 ( .A(n3936), .B(n2906), .Z(n2907) );
  XOR U4127 ( .A(n3950), .B(n2907), .Z(n2908) );
  XOR U4128 ( .A(n3952), .B(n2908), .Z(z[79]) );
  XOR U4129 ( .A(x[80]), .B(x[86]), .Z(n2909) );
  XOR U4130 ( .A(n2909), .B(x[85]), .Z(n3989) );
  IV U4131 ( .A(n3989), .Z(n2912) );
  XOR U4132 ( .A(x[84]), .B(n2912), .Z(n2978) );
  XNOR U4133 ( .A(x[87]), .B(n2912), .Z(n3974) );
  IV U4134 ( .A(x[81]), .Z(n3988) );
  IV U4135 ( .A(x[82]), .Z(n2916) );
  XOR U4136 ( .A(n3988), .B(n2916), .Z(n2920) );
  XOR U4137 ( .A(n3974), .B(n2920), .Z(n2963) );
  XOR U4138 ( .A(n3988), .B(x[83]), .Z(n2910) );
  IV U4139 ( .A(x[87]), .Z(n2925) );
  XOR U4140 ( .A(x[84]), .B(n2925), .Z(n2964) );
  XOR U4141 ( .A(n2910), .B(n2964), .Z(n2942) );
  IV U4142 ( .A(x[80]), .Z(n2989) );
  XOR U4143 ( .A(n2910), .B(n2909), .Z(n2911) );
  XOR U4144 ( .A(x[82]), .B(n2911), .Z(n3966) );
  XOR U4145 ( .A(n3966), .B(n2912), .Z(n2961) );
  XNOR U4146 ( .A(n2942), .B(n2961), .Z(n2974) );
  XOR U4147 ( .A(x[84]), .B(n2916), .Z(n2966) );
  NOR U4148 ( .A(n2974), .B(n2966), .Z(n2914) );
  XOR U4149 ( .A(n3966), .B(n3974), .Z(n2913) );
  XNOR U4150 ( .A(n2914), .B(n2913), .Z(n2915) );
  XNOR U4151 ( .A(n2989), .B(n3966), .Z(n2973) );
  NOR U4152 ( .A(n2964), .B(n2973), .Z(n2918) );
  XNOR U4153 ( .A(n2915), .B(n2918), .Z(n2932) );
  XOR U4154 ( .A(n2964), .B(n2920), .Z(n2968) );
  NANDN U4155 ( .A(n2968), .B(n2942), .Z(n2919) );
  IV U4156 ( .A(n2957), .Z(n2950) );
  XNOR U4157 ( .A(n2942), .B(n2989), .Z(n2943) );
  XNOR U4158 ( .A(n3989), .B(n2943), .Z(n2991) );
  XOR U4159 ( .A(x[87]), .B(n2916), .Z(n2983) );
  OR U4160 ( .A(n2991), .B(n2983), .Z(n2917) );
  XOR U4161 ( .A(n2918), .B(n2917), .Z(n2928) );
  XOR U4162 ( .A(n2919), .B(n2928), .Z(n2922) );
  XNOR U4163 ( .A(x[83]), .B(n2920), .Z(n2921) );
  XNOR U4164 ( .A(n2922), .B(n2921), .Z(n2924) );
  NANDN U4165 ( .A(x[80]), .B(n2978), .Z(n2923) );
  XNOR U4166 ( .A(n2924), .B(n2923), .Z(n2951) );
  ANDN U4167 ( .B(n3966), .A(n3974), .Z(n2926) );
  XOR U4168 ( .A(n3988), .B(n2925), .Z(n3975) );
  NAND U4169 ( .A(n2961), .B(n3975), .Z(n2930) );
  XOR U4170 ( .A(n2926), .B(n2930), .Z(n2927) );
  XNOR U4171 ( .A(n2928), .B(n2927), .Z(n2937) );
  IV U4172 ( .A(n2937), .Z(n2953) );
  AND U4173 ( .A(n2951), .B(n2953), .Z(n2945) );
  XNOR U4174 ( .A(n2950), .B(n2945), .Z(n2933) );
  ANDN U4175 ( .B(n3988), .A(n3989), .Z(n2929) );
  XOR U4176 ( .A(n2930), .B(n2929), .Z(n2931) );
  XOR U4177 ( .A(n2932), .B(n2931), .Z(n2952) );
  ANDN U4178 ( .B(n2933), .A(n2952), .Z(n2940) );
  NANDN U4179 ( .A(n2937), .B(n2952), .Z(n2934) );
  NANDN U4180 ( .A(n2940), .B(n2934), .Z(n2965) );
  NANDN U4181 ( .A(n2953), .B(n2951), .Z(n2935) );
  NAND U4182 ( .A(n2935), .B(n2952), .Z(n2939) );
  XNOR U4183 ( .A(n2951), .B(n2957), .Z(n2936) );
  NANDN U4184 ( .A(n2937), .B(n2936), .Z(n2938) );
  AND U4185 ( .A(n2939), .B(n2938), .Z(n2990) );
  OR U4186 ( .A(n2965), .B(n2990), .Z(n2941) );
  ANDN U4187 ( .B(n2941), .A(n2940), .Z(n2969) );
  NANDN U4188 ( .A(n2969), .B(n2942), .Z(n3985) );
  NANDN U4189 ( .A(n2965), .B(n2943), .Z(n2944) );
  XOR U4190 ( .A(n3985), .B(n2944), .Z(n2977) );
  NANDN U4191 ( .A(n2951), .B(n2957), .Z(n2948) );
  XNOR U4192 ( .A(n2945), .B(n2952), .Z(n2946) );
  NANDN U4193 ( .A(n2957), .B(n2946), .Z(n2947) );
  AND U4194 ( .A(n2948), .B(n2947), .Z(n3991) );
  NANDN U4195 ( .A(n2951), .B(n2953), .Z(n2949) );
  NANDN U4196 ( .A(n2950), .B(n2949), .Z(n2956) );
  IV U4197 ( .A(n2951), .Z(n2958) );
  XNOR U4198 ( .A(n2953), .B(n2952), .Z(n2954) );
  NANDN U4199 ( .A(n2958), .B(n2954), .Z(n2955) );
  NAND U4200 ( .A(n2956), .B(n2955), .Z(n3973) );
  IV U4201 ( .A(n3973), .Z(n3965) );
  NANDN U4202 ( .A(n3991), .B(n3965), .Z(n2960) );
  NANDN U4203 ( .A(n2958), .B(n2957), .Z(n2959) );
  NAND U4204 ( .A(n2960), .B(n2959), .Z(n3976) );
  NANDN U4205 ( .A(n3976), .B(n2961), .Z(n3968) );
  NANDN U4206 ( .A(n3991), .B(n3989), .Z(n2962) );
  XNOR U4207 ( .A(n3968), .B(n2962), .Z(n2979) );
  XOR U4208 ( .A(n2977), .B(n2979), .Z(z[82]) );
  ANDN U4209 ( .B(n2963), .A(n2965), .Z(n2971) );
  XOR U4210 ( .A(n3965), .B(n2990), .Z(n2972) );
  NANDN U4211 ( .A(n2964), .B(n2972), .Z(n2985) );
  XOR U4212 ( .A(n2965), .B(n3991), .Z(n2992) );
  XNOR U4213 ( .A(n2972), .B(n2992), .Z(n2975) );
  OR U4214 ( .A(n2966), .B(n2975), .Z(n2967) );
  XNOR U4215 ( .A(n2985), .B(n2967), .Z(n3984) );
  OR U4216 ( .A(n2969), .B(n2968), .Z(n2980) );
  XNOR U4217 ( .A(n3984), .B(n2980), .Z(n2970) );
  XOR U4218 ( .A(n2971), .B(n2970), .Z(n3981) );
  NANDN U4219 ( .A(n2973), .B(n2972), .Z(n3969) );
  OR U4220 ( .A(n2975), .B(n2974), .Z(n2976) );
  XOR U4221 ( .A(n3969), .B(n2976), .Z(n2986) );
  XOR U4222 ( .A(n2986), .B(n2977), .Z(n3972) );
  XOR U4223 ( .A(n3981), .B(n3972), .Z(n3999) );
  ANDN U4224 ( .B(n2990), .A(n2978), .Z(n2982) );
  XNOR U4225 ( .A(n2980), .B(n2979), .Z(n2981) );
  XNOR U4226 ( .A(n2982), .B(n2981), .Z(n2988) );
  NANDN U4227 ( .A(n2983), .B(n2992), .Z(n2984) );
  XNOR U4228 ( .A(n2985), .B(n2984), .Z(n3977) );
  XOR U4229 ( .A(n2986), .B(n3977), .Z(n2987) );
  XOR U4230 ( .A(n2988), .B(n2987), .Z(n3980) );
  XNOR U4231 ( .A(n3999), .B(n3980), .Z(z[81]) );
  ANDN U4232 ( .B(n2990), .A(n2989), .Z(n3987) );
  ANDN U4233 ( .B(n2992), .A(n2991), .Z(n3971) );
  XNOR U4234 ( .A(n3969), .B(z[81]), .Z(n2993) );
  XNOR U4235 ( .A(n3971), .B(n2993), .Z(n2994) );
  XOR U4236 ( .A(n3985), .B(n2994), .Z(n2995) );
  XOR U4237 ( .A(n3987), .B(n2995), .Z(z[87]) );
  XOR U4238 ( .A(x[88]), .B(x[94]), .Z(n2996) );
  XOR U4239 ( .A(n2996), .B(x[93]), .Z(n4026) );
  IV U4240 ( .A(n4026), .Z(n2999) );
  XOR U4241 ( .A(x[92]), .B(n2999), .Z(n3065) );
  XNOR U4242 ( .A(x[95]), .B(n2999), .Z(n4011) );
  IV U4243 ( .A(x[89]), .Z(n4025) );
  IV U4244 ( .A(x[90]), .Z(n3003) );
  XOR U4245 ( .A(n4025), .B(n3003), .Z(n3007) );
  XOR U4246 ( .A(n4011), .B(n3007), .Z(n3050) );
  XOR U4247 ( .A(n4025), .B(x[91]), .Z(n2997) );
  IV U4248 ( .A(x[95]), .Z(n3012) );
  XOR U4249 ( .A(x[92]), .B(n3012), .Z(n3051) );
  XOR U4250 ( .A(n2997), .B(n3051), .Z(n3029) );
  IV U4251 ( .A(x[88]), .Z(n3076) );
  XOR U4252 ( .A(n2997), .B(n2996), .Z(n2998) );
  XOR U4253 ( .A(x[90]), .B(n2998), .Z(n4001) );
  XOR U4254 ( .A(n4001), .B(n2999), .Z(n3048) );
  XNOR U4255 ( .A(n3029), .B(n3048), .Z(n3061) );
  XOR U4256 ( .A(x[92]), .B(n3003), .Z(n3053) );
  NOR U4257 ( .A(n3061), .B(n3053), .Z(n3001) );
  XOR U4258 ( .A(n4001), .B(n4011), .Z(n3000) );
  XNOR U4259 ( .A(n3001), .B(n3000), .Z(n3002) );
  XNOR U4260 ( .A(n3076), .B(n4001), .Z(n3060) );
  NOR U4261 ( .A(n3051), .B(n3060), .Z(n3005) );
  XNOR U4262 ( .A(n3002), .B(n3005), .Z(n3019) );
  XOR U4263 ( .A(n3051), .B(n3007), .Z(n3055) );
  NANDN U4264 ( .A(n3055), .B(n3029), .Z(n3006) );
  IV U4265 ( .A(n3044), .Z(n3037) );
  XNOR U4266 ( .A(n3029), .B(n3076), .Z(n3030) );
  XNOR U4267 ( .A(n4026), .B(n3030), .Z(n3078) );
  XOR U4268 ( .A(x[95]), .B(n3003), .Z(n3070) );
  OR U4269 ( .A(n3078), .B(n3070), .Z(n3004) );
  XOR U4270 ( .A(n3005), .B(n3004), .Z(n3015) );
  XOR U4271 ( .A(n3006), .B(n3015), .Z(n3009) );
  XNOR U4272 ( .A(x[91]), .B(n3007), .Z(n3008) );
  XNOR U4273 ( .A(n3009), .B(n3008), .Z(n3011) );
  NANDN U4274 ( .A(x[88]), .B(n3065), .Z(n3010) );
  XNOR U4275 ( .A(n3011), .B(n3010), .Z(n3038) );
  ANDN U4276 ( .B(n4001), .A(n4011), .Z(n3013) );
  XOR U4277 ( .A(n4025), .B(n3012), .Z(n4012) );
  NAND U4278 ( .A(n3048), .B(n4012), .Z(n3017) );
  XOR U4279 ( .A(n3013), .B(n3017), .Z(n3014) );
  XNOR U4280 ( .A(n3015), .B(n3014), .Z(n3024) );
  IV U4281 ( .A(n3024), .Z(n3040) );
  AND U4282 ( .A(n3038), .B(n3040), .Z(n3032) );
  XNOR U4283 ( .A(n3037), .B(n3032), .Z(n3020) );
  ANDN U4284 ( .B(n4025), .A(n4026), .Z(n3016) );
  XOR U4285 ( .A(n3017), .B(n3016), .Z(n3018) );
  XOR U4286 ( .A(n3019), .B(n3018), .Z(n3039) );
  ANDN U4287 ( .B(n3020), .A(n3039), .Z(n3027) );
  NANDN U4288 ( .A(n3024), .B(n3039), .Z(n3021) );
  NANDN U4289 ( .A(n3027), .B(n3021), .Z(n3052) );
  NANDN U4290 ( .A(n3040), .B(n3038), .Z(n3022) );
  NAND U4291 ( .A(n3022), .B(n3039), .Z(n3026) );
  XNOR U4292 ( .A(n3038), .B(n3044), .Z(n3023) );
  NANDN U4293 ( .A(n3024), .B(n3023), .Z(n3025) );
  AND U4294 ( .A(n3026), .B(n3025), .Z(n3077) );
  OR U4295 ( .A(n3052), .B(n3077), .Z(n3028) );
  ANDN U4296 ( .B(n3028), .A(n3027), .Z(n3056) );
  NANDN U4297 ( .A(n3056), .B(n3029), .Z(n4022) );
  NANDN U4298 ( .A(n3052), .B(n3030), .Z(n3031) );
  XOR U4299 ( .A(n4022), .B(n3031), .Z(n3064) );
  NANDN U4300 ( .A(n3038), .B(n3044), .Z(n3035) );
  XNOR U4301 ( .A(n3032), .B(n3039), .Z(n3033) );
  NANDN U4302 ( .A(n3044), .B(n3033), .Z(n3034) );
  AND U4303 ( .A(n3035), .B(n3034), .Z(n4028) );
  NANDN U4304 ( .A(n3038), .B(n3040), .Z(n3036) );
  NANDN U4305 ( .A(n3037), .B(n3036), .Z(n3043) );
  IV U4306 ( .A(n3038), .Z(n3045) );
  XNOR U4307 ( .A(n3040), .B(n3039), .Z(n3041) );
  NANDN U4308 ( .A(n3045), .B(n3041), .Z(n3042) );
  NAND U4309 ( .A(n3043), .B(n3042), .Z(n4010) );
  IV U4310 ( .A(n4010), .Z(n4000) );
  NANDN U4311 ( .A(n4028), .B(n4000), .Z(n3047) );
  NANDN U4312 ( .A(n3045), .B(n3044), .Z(n3046) );
  NAND U4313 ( .A(n3047), .B(n3046), .Z(n4013) );
  NANDN U4314 ( .A(n4013), .B(n3048), .Z(n4003) );
  NANDN U4315 ( .A(n4028), .B(n4026), .Z(n3049) );
  XNOR U4316 ( .A(n4003), .B(n3049), .Z(n3066) );
  XOR U4317 ( .A(n3064), .B(n3066), .Z(z[90]) );
  ANDN U4318 ( .B(n3050), .A(n3052), .Z(n3058) );
  XOR U4319 ( .A(n4000), .B(n3077), .Z(n3059) );
  NANDN U4320 ( .A(n3051), .B(n3059), .Z(n3072) );
  XOR U4321 ( .A(n3052), .B(n4028), .Z(n3079) );
  XNOR U4322 ( .A(n3059), .B(n3079), .Z(n3062) );
  OR U4323 ( .A(n3053), .B(n3062), .Z(n3054) );
  XNOR U4324 ( .A(n3072), .B(n3054), .Z(n4021) );
  OR U4325 ( .A(n3056), .B(n3055), .Z(n3067) );
  XNOR U4326 ( .A(n4021), .B(n3067), .Z(n3057) );
  XOR U4327 ( .A(n3058), .B(n3057), .Z(n4018) );
  NANDN U4328 ( .A(n3060), .B(n3059), .Z(n4004) );
  OR U4329 ( .A(n3062), .B(n3061), .Z(n3063) );
  XOR U4330 ( .A(n4004), .B(n3063), .Z(n3073) );
  XOR U4331 ( .A(n3073), .B(n3064), .Z(n4007) );
  XOR U4332 ( .A(n4018), .B(n4007), .Z(n4036) );
  ANDN U4333 ( .B(n3077), .A(n3065), .Z(n3069) );
  XNOR U4334 ( .A(n3067), .B(n3066), .Z(n3068) );
  XNOR U4335 ( .A(n3069), .B(n3068), .Z(n3075) );
  NANDN U4336 ( .A(n3070), .B(n3079), .Z(n3071) );
  XNOR U4337 ( .A(n3072), .B(n3071), .Z(n4014) );
  XOR U4338 ( .A(n3073), .B(n4014), .Z(n3074) );
  XOR U4339 ( .A(n3075), .B(n3074), .Z(n4017) );
  XNOR U4340 ( .A(n4036), .B(n4017), .Z(z[89]) );
  ANDN U4341 ( .B(n3077), .A(n3076), .Z(n4024) );
  ANDN U4342 ( .B(n3079), .A(n3078), .Z(n4006) );
  XNOR U4343 ( .A(n4004), .B(z[89]), .Z(n3080) );
  XNOR U4344 ( .A(n4006), .B(n3080), .Z(n3081) );
  XOR U4345 ( .A(n4022), .B(n3081), .Z(n3082) );
  XOR U4346 ( .A(n4024), .B(n3082), .Z(z[95]) );
  IV U4347 ( .A(x[97]), .Z(n3436) );
  IV U4348 ( .A(x[96]), .Z(n3105) );
  XNOR U4349 ( .A(n3105), .B(x[102]), .Z(n3083) );
  XNOR U4350 ( .A(x[101]), .B(n3083), .Z(n3437) );
  IV U4351 ( .A(n3437), .Z(n3085) );
  ANDN U4352 ( .B(n3436), .A(n3085), .Z(n3091) );
  XOR U4353 ( .A(x[97]), .B(x[103]), .Z(n3434) );
  XOR U4354 ( .A(x[97]), .B(x[99]), .Z(n3084) );
  XOR U4355 ( .A(n3430), .B(n3437), .Z(n3142) );
  NAND U4356 ( .A(n3434), .B(n3142), .Z(n3094) );
  XNOR U4357 ( .A(x[103]), .B(x[100]), .Z(n3443) );
  IV U4358 ( .A(n3443), .Z(n3088) );
  XOR U4359 ( .A(n3084), .B(n3088), .Z(n3108) );
  IV U4360 ( .A(n3108), .Z(n3124) );
  XOR U4361 ( .A(n3124), .B(n3142), .Z(n3459) );
  IV U4362 ( .A(x[100]), .Z(n3097) );
  XOR U4363 ( .A(x[98]), .B(n3097), .Z(n3445) );
  NOR U4364 ( .A(n3459), .B(n3445), .Z(n3087) );
  XOR U4365 ( .A(x[103]), .B(n3085), .Z(n3462) );
  XOR U4366 ( .A(n3430), .B(n3462), .Z(n3086) );
  XNOR U4367 ( .A(n3087), .B(n3086), .Z(n3089) );
  XNOR U4368 ( .A(n3105), .B(n3430), .Z(n3429) );
  ANDN U4369 ( .B(n3088), .A(n3429), .Z(n3093) );
  XNOR U4370 ( .A(n3089), .B(n3093), .Z(n3113) );
  XNOR U4371 ( .A(n3094), .B(n3113), .Z(n3090) );
  XNOR U4372 ( .A(n3091), .B(n3090), .Z(n3128) );
  NANDN U4373 ( .A(n3462), .B(n3430), .Z(n3096) );
  XOR U4374 ( .A(x[96]), .B(n3124), .Z(n3125) );
  XNOR U4375 ( .A(n3437), .B(n3125), .Z(n3428) );
  OR U4376 ( .A(n3465), .B(n3428), .Z(n3092) );
  XOR U4377 ( .A(n3093), .B(n3092), .Z(n3101) );
  XNOR U4378 ( .A(n3101), .B(n3094), .Z(n3095) );
  XNOR U4379 ( .A(n3096), .B(n3095), .Z(n3119) );
  XOR U4380 ( .A(x[98]), .B(n3436), .Z(n3104) );
  XNOR U4381 ( .A(n3443), .B(n3104), .Z(n3454) );
  OR U4382 ( .A(n3454), .B(n3124), .Z(n3106) );
  XOR U4383 ( .A(n3097), .B(n3437), .Z(n3472) );
  NOR U4384 ( .A(n3105), .B(n3472), .Z(n3099) );
  XNOR U4385 ( .A(x[98]), .B(n3108), .Z(n3098) );
  XNOR U4386 ( .A(n3099), .B(n3098), .Z(n3100) );
  XNOR U4387 ( .A(n3106), .B(n3100), .Z(n3103) );
  XOR U4388 ( .A(n3101), .B(n3462), .Z(n3102) );
  XNOR U4389 ( .A(n3103), .B(n3102), .Z(n3131) );
  IV U4390 ( .A(n3131), .Z(n3134) );
  NANDN U4391 ( .A(n3119), .B(n3134), .Z(n3136) );
  XNOR U4392 ( .A(n3462), .B(n3104), .Z(n3452) );
  ANDN U4393 ( .B(n3105), .A(n3452), .Z(n3107) );
  XOR U4394 ( .A(n3107), .B(n3106), .Z(n3110) );
  NANDN U4395 ( .A(n3108), .B(n3452), .Z(n3109) );
  NAND U4396 ( .A(n3110), .B(n3109), .Z(n3111) );
  XNOR U4397 ( .A(n3111), .B(n3472), .Z(n3112) );
  XOR U4398 ( .A(n3113), .B(n3112), .Z(n3139) );
  IV U4399 ( .A(n3139), .Z(n3135) );
  XNOR U4400 ( .A(n3136), .B(n3135), .Z(n3114) );
  NANDN U4401 ( .A(n3128), .B(n3114), .Z(n3116) );
  IV U4402 ( .A(n3128), .Z(n3137) );
  ANDN U4403 ( .B(n3119), .A(n3137), .Z(n3115) );
  ANDN U4404 ( .B(n3116), .A(n3115), .Z(n3451) );
  IV U4405 ( .A(n3119), .Z(n3129) );
  NANDN U4406 ( .A(n3129), .B(n3134), .Z(n3117) );
  NANDN U4407 ( .A(n3137), .B(n3117), .Z(n3121) );
  XNOR U4408 ( .A(n3134), .B(n3139), .Z(n3118) );
  NANDN U4409 ( .A(n3119), .B(n3118), .Z(n3120) );
  NAND U4410 ( .A(n3121), .B(n3120), .Z(n3471) );
  OR U4411 ( .A(n3451), .B(n3471), .Z(n3123) );
  NANDN U4412 ( .A(n3137), .B(n3129), .Z(n3122) );
  NAND U4413 ( .A(n3123), .B(n3122), .Z(n3453) );
  OR U4414 ( .A(n3453), .B(n3124), .Z(n3448) );
  OR U4415 ( .A(n3451), .B(n3125), .Z(n3126) );
  XNOR U4416 ( .A(n3448), .B(n3126), .Z(n3461) );
  NANDN U4417 ( .A(n3134), .B(n3129), .Z(n3127) );
  NANDN U4418 ( .A(n3135), .B(n3127), .Z(n3133) );
  XNOR U4419 ( .A(n3129), .B(n3128), .Z(n3130) );
  NANDN U4420 ( .A(n3131), .B(n3130), .Z(n3132) );
  AND U4421 ( .A(n3133), .B(n3132), .Z(n3463) );
  NANDN U4422 ( .A(n3135), .B(n3134), .Z(n3141) );
  XOR U4423 ( .A(n3137), .B(n3136), .Z(n3138) );
  NANDN U4424 ( .A(n3139), .B(n3138), .Z(n3140) );
  AND U4425 ( .A(n3141), .B(n3140), .Z(n3438) );
  XNOR U4426 ( .A(n3463), .B(n3438), .Z(n3435) );
  NANDN U4427 ( .A(n3435), .B(n3142), .Z(n3432) );
  ANDN U4428 ( .B(n3438), .A(n3437), .Z(n3143) );
  XNOR U4429 ( .A(n3432), .B(n3143), .Z(n3480) );
  XOR U4430 ( .A(n3461), .B(n3480), .Z(z[98]) );
  IV U4431 ( .A(x[108]), .Z(n3144) );
  IV U4432 ( .A(x[104]), .Z(n3229) );
  XOR U4433 ( .A(n3229), .B(x[110]), .Z(n3145) );
  XOR U4434 ( .A(n3145), .B(x[109]), .Z(n3169) );
  IV U4435 ( .A(n3169), .Z(n3511) );
  XOR U4436 ( .A(n3144), .B(n3511), .Z(n3218) );
  XOR U4437 ( .A(x[105]), .B(x[107]), .Z(n3146) );
  XOR U4438 ( .A(x[111]), .B(n3144), .Z(n3204) );
  XNOR U4439 ( .A(n3146), .B(n3204), .Z(n3183) );
  IV U4440 ( .A(n3183), .Z(n3161) );
  XOR U4441 ( .A(n3146), .B(n3145), .Z(n3147) );
  XOR U4442 ( .A(x[106]), .B(n3147), .Z(n3488) );
  XOR U4443 ( .A(n3488), .B(n3169), .Z(n3201) );
  XOR U4444 ( .A(n3161), .B(n3201), .Z(n3214) );
  IV U4445 ( .A(x[106]), .Z(n3157) );
  XOR U4446 ( .A(x[108]), .B(n3157), .Z(n3206) );
  NOR U4447 ( .A(n3214), .B(n3206), .Z(n3149) );
  XOR U4448 ( .A(x[111]), .B(n3511), .Z(n3496) );
  XOR U4449 ( .A(n3488), .B(n3496), .Z(n3148) );
  XNOR U4450 ( .A(n3149), .B(n3148), .Z(n3150) );
  XNOR U4451 ( .A(n3229), .B(n3488), .Z(n3213) );
  NOR U4452 ( .A(n3204), .B(n3213), .Z(n3159) );
  XNOR U4453 ( .A(n3150), .B(n3159), .Z(n3171) );
  IV U4454 ( .A(x[105]), .Z(n3510) );
  XNOR U4455 ( .A(n3510), .B(x[106]), .Z(n3151) );
  XNOR U4456 ( .A(n3496), .B(n3151), .Z(n3203) );
  ANDN U4457 ( .B(n3203), .A(x[104]), .Z(n3152) );
  XNOR U4458 ( .A(n3204), .B(n3151), .Z(n3208) );
  NANDN U4459 ( .A(n3161), .B(n3208), .Z(n3162) );
  XOR U4460 ( .A(n3152), .B(n3162), .Z(n3154) );
  OR U4461 ( .A(n3203), .B(n3183), .Z(n3153) );
  NAND U4462 ( .A(n3154), .B(n3153), .Z(n3155) );
  XOR U4463 ( .A(n3171), .B(n3155), .Z(n3156) );
  XOR U4464 ( .A(n3218), .B(n3156), .Z(n3197) );
  XNOR U4465 ( .A(n3161), .B(x[104]), .Z(n3184) );
  XNOR U4466 ( .A(n3511), .B(n3184), .Z(n3231) );
  IV U4467 ( .A(x[111]), .Z(n3160) );
  XOR U4468 ( .A(n3160), .B(n3157), .Z(n3223) );
  NANDN U4469 ( .A(n3231), .B(n3223), .Z(n3158) );
  XOR U4470 ( .A(n3159), .B(n3158), .Z(n3166) );
  XOR U4471 ( .A(n3510), .B(n3160), .Z(n3497) );
  NAND U4472 ( .A(n3201), .B(n3497), .Z(n3170) );
  ANDN U4473 ( .B(n3218), .A(n3229), .Z(n3164) );
  XNOR U4474 ( .A(n3162), .B(n3161), .Z(n3163) );
  XNOR U4475 ( .A(n3164), .B(n3163), .Z(n3165) );
  XNOR U4476 ( .A(n3166), .B(n3165), .Z(n3168) );
  XNOR U4477 ( .A(x[106]), .B(n3496), .Z(n3167) );
  XNOR U4478 ( .A(n3168), .B(n3167), .Z(n3198) );
  IV U4479 ( .A(n3198), .Z(n3190) );
  AND U4480 ( .A(n3193), .B(n3190), .Z(n3186) );
  XOR U4481 ( .A(n3197), .B(n3186), .Z(n3174) );
  ANDN U4482 ( .B(n3169), .A(x[105]), .Z(n3173) );
  XNOR U4483 ( .A(n3171), .B(n3170), .Z(n3172) );
  XNOR U4484 ( .A(n3173), .B(n3172), .Z(n3192) );
  ANDN U4485 ( .B(n3174), .A(n3192), .Z(n3181) );
  IV U4486 ( .A(n3193), .Z(n3178) );
  NANDN U4487 ( .A(n3178), .B(n3192), .Z(n3175) );
  NANDN U4488 ( .A(n3181), .B(n3175), .Z(n3205) );
  NANDN U4489 ( .A(n3193), .B(n3190), .Z(n3176) );
  NAND U4490 ( .A(n3176), .B(n3192), .Z(n3180) );
  XNOR U4491 ( .A(n3190), .B(n3197), .Z(n3177) );
  NANDN U4492 ( .A(n3178), .B(n3177), .Z(n3179) );
  AND U4493 ( .A(n3180), .B(n3179), .Z(n3230) );
  OR U4494 ( .A(n3205), .B(n3230), .Z(n3182) );
  ANDN U4495 ( .B(n3182), .A(n3181), .Z(n3209) );
  NANDN U4496 ( .A(n3209), .B(n3183), .Z(n3507) );
  NANDN U4497 ( .A(n3205), .B(n3184), .Z(n3185) );
  XOR U4498 ( .A(n3507), .B(n3185), .Z(n3217) );
  NANDN U4499 ( .A(n3190), .B(n3197), .Z(n3189) );
  XNOR U4500 ( .A(n3186), .B(n3192), .Z(n3187) );
  NANDN U4501 ( .A(n3197), .B(n3187), .Z(n3188) );
  AND U4502 ( .A(n3189), .B(n3188), .Z(n3513) );
  NANDN U4503 ( .A(n3190), .B(n3193), .Z(n3191) );
  NAND U4504 ( .A(n3197), .B(n3191), .Z(n3196) );
  XNOR U4505 ( .A(n3193), .B(n3192), .Z(n3194) );
  NANDN U4506 ( .A(n3198), .B(n3194), .Z(n3195) );
  NAND U4507 ( .A(n3196), .B(n3195), .Z(n3495) );
  IV U4508 ( .A(n3495), .Z(n3487) );
  NANDN U4509 ( .A(n3513), .B(n3487), .Z(n3200) );
  NANDN U4510 ( .A(n3198), .B(n3197), .Z(n3199) );
  NAND U4511 ( .A(n3200), .B(n3199), .Z(n3498) );
  NANDN U4512 ( .A(n3498), .B(n3201), .Z(n3490) );
  NANDN U4513 ( .A(n3513), .B(n3511), .Z(n3202) );
  XNOR U4514 ( .A(n3490), .B(n3202), .Z(n3219) );
  XOR U4515 ( .A(n3217), .B(n3219), .Z(z[106]) );
  NOR U4516 ( .A(n3205), .B(n3203), .Z(n3211) );
  XOR U4517 ( .A(n3487), .B(n3230), .Z(n3212) );
  NANDN U4518 ( .A(n3204), .B(n3212), .Z(n3225) );
  XOR U4519 ( .A(n3205), .B(n3513), .Z(n3232) );
  XNOR U4520 ( .A(n3212), .B(n3232), .Z(n3215) );
  OR U4521 ( .A(n3206), .B(n3215), .Z(n3207) );
  XNOR U4522 ( .A(n3225), .B(n3207), .Z(n3506) );
  NANDN U4523 ( .A(n3209), .B(n3208), .Z(n3220) );
  XNOR U4524 ( .A(n3506), .B(n3220), .Z(n3210) );
  XOR U4525 ( .A(n3211), .B(n3210), .Z(n3503) );
  NANDN U4526 ( .A(n3213), .B(n3212), .Z(n3491) );
  OR U4527 ( .A(n3215), .B(n3214), .Z(n3216) );
  XOR U4528 ( .A(n3491), .B(n3216), .Z(n3226) );
  XOR U4529 ( .A(n3226), .B(n3217), .Z(n3494) );
  XOR U4530 ( .A(n3503), .B(n3494), .Z(n3521) );
  ANDN U4531 ( .B(n3230), .A(n3218), .Z(n3222) );
  XNOR U4532 ( .A(n3220), .B(n3219), .Z(n3221) );
  XNOR U4533 ( .A(n3222), .B(n3221), .Z(n3228) );
  NAND U4534 ( .A(n3223), .B(n3232), .Z(n3224) );
  XNOR U4535 ( .A(n3225), .B(n3224), .Z(n3499) );
  XOR U4536 ( .A(n3226), .B(n3499), .Z(n3227) );
  XOR U4537 ( .A(n3228), .B(n3227), .Z(n3502) );
  XNOR U4538 ( .A(n3521), .B(n3502), .Z(z[105]) );
  ANDN U4539 ( .B(n3230), .A(n3229), .Z(n3509) );
  ANDN U4540 ( .B(n3232), .A(n3231), .Z(n3493) );
  XNOR U4541 ( .A(n3491), .B(z[105]), .Z(n3233) );
  XNOR U4542 ( .A(n3493), .B(n3233), .Z(n3234) );
  XOR U4543 ( .A(n3507), .B(n3234), .Z(n3235) );
  XOR U4544 ( .A(n3509), .B(n3235), .Z(z[111]) );
  IV U4545 ( .A(x[116]), .Z(n3236) );
  IV U4546 ( .A(x[112]), .Z(n3321) );
  XOR U4547 ( .A(n3321), .B(x[118]), .Z(n3237) );
  XOR U4548 ( .A(n3237), .B(x[117]), .Z(n3261) );
  IV U4549 ( .A(n3261), .Z(n3546) );
  XOR U4550 ( .A(n3236), .B(n3546), .Z(n3310) );
  XOR U4551 ( .A(x[113]), .B(x[115]), .Z(n3238) );
  XOR U4552 ( .A(x[119]), .B(n3236), .Z(n3296) );
  XNOR U4553 ( .A(n3238), .B(n3296), .Z(n3275) );
  IV U4554 ( .A(n3275), .Z(n3253) );
  XOR U4555 ( .A(n3238), .B(n3237), .Z(n3239) );
  XOR U4556 ( .A(x[114]), .B(n3239), .Z(n3523) );
  XOR U4557 ( .A(n3523), .B(n3261), .Z(n3293) );
  XOR U4558 ( .A(n3253), .B(n3293), .Z(n3306) );
  IV U4559 ( .A(x[114]), .Z(n3249) );
  XOR U4560 ( .A(x[116]), .B(n3249), .Z(n3298) );
  NOR U4561 ( .A(n3306), .B(n3298), .Z(n3241) );
  XOR U4562 ( .A(x[119]), .B(n3546), .Z(n3531) );
  XOR U4563 ( .A(n3523), .B(n3531), .Z(n3240) );
  XNOR U4564 ( .A(n3241), .B(n3240), .Z(n3242) );
  XNOR U4565 ( .A(n3321), .B(n3523), .Z(n3305) );
  NOR U4566 ( .A(n3296), .B(n3305), .Z(n3251) );
  XNOR U4567 ( .A(n3242), .B(n3251), .Z(n3263) );
  IV U4568 ( .A(x[113]), .Z(n3545) );
  XNOR U4569 ( .A(n3545), .B(x[114]), .Z(n3243) );
  XNOR U4570 ( .A(n3531), .B(n3243), .Z(n3295) );
  ANDN U4571 ( .B(n3295), .A(x[112]), .Z(n3244) );
  XNOR U4572 ( .A(n3296), .B(n3243), .Z(n3300) );
  NANDN U4573 ( .A(n3253), .B(n3300), .Z(n3254) );
  XOR U4574 ( .A(n3244), .B(n3254), .Z(n3246) );
  OR U4575 ( .A(n3295), .B(n3275), .Z(n3245) );
  NAND U4576 ( .A(n3246), .B(n3245), .Z(n3247) );
  XOR U4577 ( .A(n3263), .B(n3247), .Z(n3248) );
  XOR U4578 ( .A(n3310), .B(n3248), .Z(n3289) );
  XNOR U4579 ( .A(n3253), .B(x[112]), .Z(n3276) );
  XNOR U4580 ( .A(n3546), .B(n3276), .Z(n3323) );
  IV U4581 ( .A(x[119]), .Z(n3252) );
  XOR U4582 ( .A(n3252), .B(n3249), .Z(n3315) );
  NANDN U4583 ( .A(n3323), .B(n3315), .Z(n3250) );
  XOR U4584 ( .A(n3251), .B(n3250), .Z(n3258) );
  XOR U4585 ( .A(n3545), .B(n3252), .Z(n3532) );
  NAND U4586 ( .A(n3293), .B(n3532), .Z(n3262) );
  ANDN U4587 ( .B(n3310), .A(n3321), .Z(n3256) );
  XNOR U4588 ( .A(n3254), .B(n3253), .Z(n3255) );
  XNOR U4589 ( .A(n3256), .B(n3255), .Z(n3257) );
  XNOR U4590 ( .A(n3258), .B(n3257), .Z(n3260) );
  XNOR U4591 ( .A(x[114]), .B(n3531), .Z(n3259) );
  XNOR U4592 ( .A(n3260), .B(n3259), .Z(n3290) );
  IV U4593 ( .A(n3290), .Z(n3282) );
  AND U4594 ( .A(n3285), .B(n3282), .Z(n3278) );
  XOR U4595 ( .A(n3289), .B(n3278), .Z(n3266) );
  ANDN U4596 ( .B(n3261), .A(x[113]), .Z(n3265) );
  XNOR U4597 ( .A(n3263), .B(n3262), .Z(n3264) );
  XNOR U4598 ( .A(n3265), .B(n3264), .Z(n3284) );
  ANDN U4599 ( .B(n3266), .A(n3284), .Z(n3273) );
  IV U4600 ( .A(n3285), .Z(n3270) );
  NANDN U4601 ( .A(n3270), .B(n3284), .Z(n3267) );
  NANDN U4602 ( .A(n3273), .B(n3267), .Z(n3297) );
  NANDN U4603 ( .A(n3285), .B(n3282), .Z(n3268) );
  NAND U4604 ( .A(n3268), .B(n3284), .Z(n3272) );
  XNOR U4605 ( .A(n3282), .B(n3289), .Z(n3269) );
  NANDN U4606 ( .A(n3270), .B(n3269), .Z(n3271) );
  AND U4607 ( .A(n3272), .B(n3271), .Z(n3322) );
  OR U4608 ( .A(n3297), .B(n3322), .Z(n3274) );
  ANDN U4609 ( .B(n3274), .A(n3273), .Z(n3301) );
  NANDN U4610 ( .A(n3301), .B(n3275), .Z(n3542) );
  NANDN U4611 ( .A(n3297), .B(n3276), .Z(n3277) );
  XOR U4612 ( .A(n3542), .B(n3277), .Z(n3309) );
  NANDN U4613 ( .A(n3282), .B(n3289), .Z(n3281) );
  XNOR U4614 ( .A(n3278), .B(n3284), .Z(n3279) );
  NANDN U4615 ( .A(n3289), .B(n3279), .Z(n3280) );
  AND U4616 ( .A(n3281), .B(n3280), .Z(n3548) );
  NANDN U4617 ( .A(n3282), .B(n3285), .Z(n3283) );
  NAND U4618 ( .A(n3289), .B(n3283), .Z(n3288) );
  XNOR U4619 ( .A(n3285), .B(n3284), .Z(n3286) );
  NANDN U4620 ( .A(n3290), .B(n3286), .Z(n3287) );
  NAND U4621 ( .A(n3288), .B(n3287), .Z(n3530) );
  IV U4622 ( .A(n3530), .Z(n3522) );
  NANDN U4623 ( .A(n3548), .B(n3522), .Z(n3292) );
  NANDN U4624 ( .A(n3290), .B(n3289), .Z(n3291) );
  NAND U4625 ( .A(n3292), .B(n3291), .Z(n3533) );
  NANDN U4626 ( .A(n3533), .B(n3293), .Z(n3525) );
  NANDN U4627 ( .A(n3548), .B(n3546), .Z(n3294) );
  XNOR U4628 ( .A(n3525), .B(n3294), .Z(n3311) );
  XOR U4629 ( .A(n3309), .B(n3311), .Z(z[114]) );
  NOR U4630 ( .A(n3297), .B(n3295), .Z(n3303) );
  XOR U4631 ( .A(n3522), .B(n3322), .Z(n3304) );
  NANDN U4632 ( .A(n3296), .B(n3304), .Z(n3317) );
  XOR U4633 ( .A(n3297), .B(n3548), .Z(n3324) );
  XNOR U4634 ( .A(n3304), .B(n3324), .Z(n3307) );
  OR U4635 ( .A(n3298), .B(n3307), .Z(n3299) );
  XNOR U4636 ( .A(n3317), .B(n3299), .Z(n3541) );
  NANDN U4637 ( .A(n3301), .B(n3300), .Z(n3312) );
  XNOR U4638 ( .A(n3541), .B(n3312), .Z(n3302) );
  XOR U4639 ( .A(n3303), .B(n3302), .Z(n3538) );
  NANDN U4640 ( .A(n3305), .B(n3304), .Z(n3526) );
  OR U4641 ( .A(n3307), .B(n3306), .Z(n3308) );
  XOR U4642 ( .A(n3526), .B(n3308), .Z(n3318) );
  XOR U4643 ( .A(n3318), .B(n3309), .Z(n3529) );
  XOR U4644 ( .A(n3538), .B(n3529), .Z(n3556) );
  ANDN U4645 ( .B(n3322), .A(n3310), .Z(n3314) );
  XNOR U4646 ( .A(n3312), .B(n3311), .Z(n3313) );
  XNOR U4647 ( .A(n3314), .B(n3313), .Z(n3320) );
  NAND U4648 ( .A(n3315), .B(n3324), .Z(n3316) );
  XNOR U4649 ( .A(n3317), .B(n3316), .Z(n3534) );
  XOR U4650 ( .A(n3318), .B(n3534), .Z(n3319) );
  XOR U4651 ( .A(n3320), .B(n3319), .Z(n3537) );
  XNOR U4652 ( .A(n3556), .B(n3537), .Z(z[113]) );
  ANDN U4653 ( .B(n3322), .A(n3321), .Z(n3544) );
  ANDN U4654 ( .B(n3324), .A(n3323), .Z(n3528) );
  XNOR U4655 ( .A(n3526), .B(z[113]), .Z(n3325) );
  XNOR U4656 ( .A(n3528), .B(n3325), .Z(n3326) );
  XOR U4657 ( .A(n3542), .B(n3326), .Z(n3327) );
  XOR U4658 ( .A(n3544), .B(n3327), .Z(z[119]) );
  IV U4659 ( .A(x[124]), .Z(n3328) );
  IV U4660 ( .A(x[120]), .Z(n3413) );
  XOR U4661 ( .A(n3413), .B(x[126]), .Z(n3329) );
  XOR U4662 ( .A(n3329), .B(x[125]), .Z(n3353) );
  IV U4663 ( .A(n3353), .Z(n3612) );
  XOR U4664 ( .A(n3328), .B(n3612), .Z(n3402) );
  XOR U4665 ( .A(x[121]), .B(x[123]), .Z(n3330) );
  XOR U4666 ( .A(x[127]), .B(n3328), .Z(n3388) );
  XNOR U4667 ( .A(n3330), .B(n3388), .Z(n3367) );
  IV U4668 ( .A(n3367), .Z(n3345) );
  XOR U4669 ( .A(n3330), .B(n3329), .Z(n3331) );
  XOR U4670 ( .A(x[122]), .B(n3331), .Z(n3589) );
  XOR U4671 ( .A(n3589), .B(n3353), .Z(n3385) );
  XOR U4672 ( .A(n3345), .B(n3385), .Z(n3398) );
  IV U4673 ( .A(x[122]), .Z(n3341) );
  XOR U4674 ( .A(x[124]), .B(n3341), .Z(n3390) );
  NOR U4675 ( .A(n3398), .B(n3390), .Z(n3333) );
  XOR U4676 ( .A(x[127]), .B(n3612), .Z(n3597) );
  XOR U4677 ( .A(n3589), .B(n3597), .Z(n3332) );
  XNOR U4678 ( .A(n3333), .B(n3332), .Z(n3334) );
  XNOR U4679 ( .A(n3413), .B(n3589), .Z(n3397) );
  NOR U4680 ( .A(n3388), .B(n3397), .Z(n3343) );
  XNOR U4681 ( .A(n3334), .B(n3343), .Z(n3355) );
  IV U4682 ( .A(x[121]), .Z(n3611) );
  XNOR U4683 ( .A(n3611), .B(x[122]), .Z(n3335) );
  XNOR U4684 ( .A(n3597), .B(n3335), .Z(n3387) );
  ANDN U4685 ( .B(n3387), .A(x[120]), .Z(n3336) );
  XNOR U4686 ( .A(n3388), .B(n3335), .Z(n3392) );
  NANDN U4687 ( .A(n3345), .B(n3392), .Z(n3346) );
  XOR U4688 ( .A(n3336), .B(n3346), .Z(n3338) );
  OR U4689 ( .A(n3387), .B(n3367), .Z(n3337) );
  NAND U4690 ( .A(n3338), .B(n3337), .Z(n3339) );
  XOR U4691 ( .A(n3355), .B(n3339), .Z(n3340) );
  XOR U4692 ( .A(n3402), .B(n3340), .Z(n3381) );
  XNOR U4693 ( .A(n3345), .B(x[120]), .Z(n3368) );
  XNOR U4694 ( .A(n3612), .B(n3368), .Z(n3415) );
  IV U4695 ( .A(x[127]), .Z(n3344) );
  XOR U4696 ( .A(n3344), .B(n3341), .Z(n3407) );
  NANDN U4697 ( .A(n3415), .B(n3407), .Z(n3342) );
  XOR U4698 ( .A(n3343), .B(n3342), .Z(n3350) );
  XOR U4699 ( .A(n3611), .B(n3344), .Z(n3598) );
  NAND U4700 ( .A(n3385), .B(n3598), .Z(n3354) );
  ANDN U4701 ( .B(n3402), .A(n3413), .Z(n3348) );
  XNOR U4702 ( .A(n3346), .B(n3345), .Z(n3347) );
  XNOR U4703 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4704 ( .A(n3350), .B(n3349), .Z(n3352) );
  XNOR U4705 ( .A(x[122]), .B(n3597), .Z(n3351) );
  XNOR U4706 ( .A(n3352), .B(n3351), .Z(n3382) );
  IV U4707 ( .A(n3382), .Z(n3374) );
  AND U4708 ( .A(n3377), .B(n3374), .Z(n3370) );
  XOR U4709 ( .A(n3381), .B(n3370), .Z(n3358) );
  ANDN U4710 ( .B(n3353), .A(x[121]), .Z(n3357) );
  XNOR U4711 ( .A(n3355), .B(n3354), .Z(n3356) );
  XNOR U4712 ( .A(n3357), .B(n3356), .Z(n3376) );
  ANDN U4713 ( .B(n3358), .A(n3376), .Z(n3365) );
  IV U4714 ( .A(n3377), .Z(n3362) );
  NANDN U4715 ( .A(n3362), .B(n3376), .Z(n3359) );
  NANDN U4716 ( .A(n3365), .B(n3359), .Z(n3389) );
  NANDN U4717 ( .A(n3377), .B(n3374), .Z(n3360) );
  NAND U4718 ( .A(n3360), .B(n3376), .Z(n3364) );
  XNOR U4719 ( .A(n3374), .B(n3381), .Z(n3361) );
  NANDN U4720 ( .A(n3362), .B(n3361), .Z(n3363) );
  AND U4721 ( .A(n3364), .B(n3363), .Z(n3414) );
  OR U4722 ( .A(n3389), .B(n3414), .Z(n3366) );
  ANDN U4723 ( .B(n3366), .A(n3365), .Z(n3393) );
  NANDN U4724 ( .A(n3393), .B(n3367), .Z(n3608) );
  NANDN U4725 ( .A(n3389), .B(n3368), .Z(n3369) );
  XOR U4726 ( .A(n3608), .B(n3369), .Z(n3401) );
  NANDN U4727 ( .A(n3374), .B(n3381), .Z(n3373) );
  XNOR U4728 ( .A(n3370), .B(n3376), .Z(n3371) );
  NANDN U4729 ( .A(n3381), .B(n3371), .Z(n3372) );
  AND U4730 ( .A(n3373), .B(n3372), .Z(n3614) );
  NANDN U4731 ( .A(n3374), .B(n3377), .Z(n3375) );
  NAND U4732 ( .A(n3381), .B(n3375), .Z(n3380) );
  XNOR U4733 ( .A(n3377), .B(n3376), .Z(n3378) );
  NANDN U4734 ( .A(n3382), .B(n3378), .Z(n3379) );
  NAND U4735 ( .A(n3380), .B(n3379), .Z(n3596) );
  IV U4736 ( .A(n3596), .Z(n3588) );
  NANDN U4737 ( .A(n3614), .B(n3588), .Z(n3384) );
  NANDN U4738 ( .A(n3382), .B(n3381), .Z(n3383) );
  NAND U4739 ( .A(n3384), .B(n3383), .Z(n3599) );
  NANDN U4740 ( .A(n3599), .B(n3385), .Z(n3591) );
  NANDN U4741 ( .A(n3614), .B(n3612), .Z(n3386) );
  XNOR U4742 ( .A(n3591), .B(n3386), .Z(n3403) );
  XOR U4743 ( .A(n3401), .B(n3403), .Z(z[122]) );
  NOR U4744 ( .A(n3389), .B(n3387), .Z(n3395) );
  XOR U4745 ( .A(n3588), .B(n3414), .Z(n3396) );
  NANDN U4746 ( .A(n3388), .B(n3396), .Z(n3409) );
  XOR U4747 ( .A(n3389), .B(n3614), .Z(n3416) );
  XNOR U4748 ( .A(n3396), .B(n3416), .Z(n3399) );
  OR U4749 ( .A(n3390), .B(n3399), .Z(n3391) );
  XNOR U4750 ( .A(n3409), .B(n3391), .Z(n3607) );
  NANDN U4751 ( .A(n3393), .B(n3392), .Z(n3404) );
  XNOR U4752 ( .A(n3607), .B(n3404), .Z(n3394) );
  XOR U4753 ( .A(n3395), .B(n3394), .Z(n3604) );
  NANDN U4754 ( .A(n3397), .B(n3396), .Z(n3592) );
  OR U4755 ( .A(n3399), .B(n3398), .Z(n3400) );
  XOR U4756 ( .A(n3592), .B(n3400), .Z(n3410) );
  XOR U4757 ( .A(n3410), .B(n3401), .Z(n3595) );
  XOR U4758 ( .A(n3604), .B(n3595), .Z(n3622) );
  ANDN U4759 ( .B(n3414), .A(n3402), .Z(n3406) );
  XNOR U4760 ( .A(n3404), .B(n3403), .Z(n3405) );
  XNOR U4761 ( .A(n3406), .B(n3405), .Z(n3412) );
  NAND U4762 ( .A(n3407), .B(n3416), .Z(n3408) );
  XNOR U4763 ( .A(n3409), .B(n3408), .Z(n3600) );
  XOR U4764 ( .A(n3410), .B(n3600), .Z(n3411) );
  XOR U4765 ( .A(n3412), .B(n3411), .Z(n3603) );
  XNOR U4766 ( .A(n3622), .B(n3603), .Z(z[121]) );
  ANDN U4767 ( .B(n3414), .A(n3413), .Z(n3610) );
  ANDN U4768 ( .B(n3416), .A(n3415), .Z(n3594) );
  XNOR U4769 ( .A(n3592), .B(z[121]), .Z(n3417) );
  XNOR U4770 ( .A(n3594), .B(n3417), .Z(n3418) );
  XOR U4771 ( .A(n3608), .B(n3418), .Z(n3419) );
  XOR U4772 ( .A(n3610), .B(n3419), .Z(z[127]) );
  NANDN U4773 ( .A(n3421), .B(n3420), .Z(n3422) );
  XNOR U4774 ( .A(n3423), .B(n3422), .Z(n3873) );
  XNOR U4775 ( .A(n3424), .B(n3873), .Z(n3425) );
  XOR U4776 ( .A(n3426), .B(n3425), .Z(n3816) );
  XOR U4777 ( .A(n3816), .B(n3427), .Z(z[0]) );
  XNOR U4778 ( .A(n3438), .B(n3451), .Z(n3464) );
  ANDN U4779 ( .B(n3464), .A(n3428), .Z(n3485) );
  NANDN U4780 ( .A(n3429), .B(n3444), .Z(n3483) );
  NANDN U4781 ( .A(n3430), .B(n3463), .Z(n3431) );
  XNOR U4782 ( .A(n3432), .B(n3431), .Z(n3442) );
  XNOR U4783 ( .A(n3483), .B(n3442), .Z(n3433) );
  XOR U4784 ( .A(n3485), .B(n3433), .Z(n4038) );
  XNOR U4785 ( .A(n4038), .B(z[98]), .Z(z[100]) );
  NANDN U4786 ( .A(n3435), .B(n3434), .Z(n3468) );
  XOR U4787 ( .A(n3437), .B(n3436), .Z(n3439) );
  NAND U4788 ( .A(n3439), .B(n3438), .Z(n3440) );
  XOR U4789 ( .A(n3468), .B(n3440), .Z(n3441) );
  XNOR U4790 ( .A(n3442), .B(n3441), .Z(n3450) );
  NANDN U4791 ( .A(n3443), .B(n3444), .Z(n3467) );
  XNOR U4792 ( .A(n3444), .B(n3464), .Z(n3458) );
  OR U4793 ( .A(n3458), .B(n3445), .Z(n3446) );
  XNOR U4794 ( .A(n3467), .B(n3446), .Z(n3455) );
  NANDN U4795 ( .A(n3471), .B(x[96]), .Z(n3447) );
  XNOR U4796 ( .A(n3448), .B(n3447), .Z(n3482) );
  XNOR U4797 ( .A(n3455), .B(n3482), .Z(n3449) );
  XOR U4798 ( .A(n3450), .B(n3449), .Z(z[101]) );
  ANDN U4799 ( .B(n3452), .A(n3451), .Z(n3457) );
  OR U4800 ( .A(n3454), .B(n3453), .Z(n3477) );
  XNOR U4801 ( .A(n3477), .B(n3455), .Z(n3456) );
  XOR U4802 ( .A(n3457), .B(n3456), .Z(n4039) );
  OR U4803 ( .A(n3459), .B(n3458), .Z(n3460) );
  XOR U4804 ( .A(n3483), .B(n3460), .Z(n3474) );
  XOR U4805 ( .A(n3474), .B(n3461), .Z(n4037) );
  XNOR U4806 ( .A(n4039), .B(n4037), .Z(n3481) );
  AND U4807 ( .A(n3463), .B(n3462), .Z(n3470) );
  NANDN U4808 ( .A(n3465), .B(n3464), .Z(n3466) );
  XNOR U4809 ( .A(n3467), .B(n3466), .Z(n3473) );
  XNOR U4810 ( .A(n3473), .B(n3468), .Z(n3469) );
  XOR U4811 ( .A(n3470), .B(n3469), .Z(n4042) );
  XNOR U4812 ( .A(n3481), .B(n4042), .Z(z[102]) );
  ANDN U4813 ( .B(n3472), .A(n3471), .Z(n3476) );
  XOR U4814 ( .A(n3474), .B(n3473), .Z(n3475) );
  XNOR U4815 ( .A(n3476), .B(n3475), .Z(n3478) );
  XNOR U4816 ( .A(n3478), .B(n3477), .Z(n3479) );
  XNOR U4817 ( .A(n3480), .B(n3479), .Z(n4040) );
  XNOR U4818 ( .A(n4040), .B(n3481), .Z(z[97]) );
  XNOR U4819 ( .A(n3483), .B(n3482), .Z(n3484) );
  XNOR U4820 ( .A(n3485), .B(n3484), .Z(n3486) );
  XOR U4821 ( .A(n3486), .B(z[97]), .Z(z[103]) );
  NANDN U4822 ( .A(n3488), .B(n3487), .Z(n3489) );
  XNOR U4823 ( .A(n3490), .B(n3489), .Z(n3517) );
  XNOR U4824 ( .A(n3491), .B(n3517), .Z(n3492) );
  XOR U4825 ( .A(n3493), .B(n3492), .Z(n3505) );
  XOR U4826 ( .A(n3505), .B(n3494), .Z(z[104]) );
  ANDN U4827 ( .B(n3496), .A(n3495), .Z(n3501) );
  NANDN U4828 ( .A(n3498), .B(n3497), .Z(n3515) );
  XNOR U4829 ( .A(n3499), .B(n3515), .Z(n3500) );
  XOR U4830 ( .A(n3501), .B(n3500), .Z(n3520) );
  XOR U4831 ( .A(n3503), .B(n3502), .Z(n3504) );
  XOR U4832 ( .A(n3520), .B(n3504), .Z(z[107]) );
  XNOR U4833 ( .A(n3505), .B(z[106]), .Z(z[108]) );
  XNOR U4834 ( .A(n3507), .B(n3506), .Z(n3508) );
  XNOR U4835 ( .A(n3509), .B(n3508), .Z(n3519) );
  XNOR U4836 ( .A(n3511), .B(n3510), .Z(n3512) );
  NANDN U4837 ( .A(n3513), .B(n3512), .Z(n3514) );
  XOR U4838 ( .A(n3515), .B(n3514), .Z(n3516) );
  XNOR U4839 ( .A(n3517), .B(n3516), .Z(n3518) );
  XNOR U4840 ( .A(n3519), .B(n3518), .Z(z[109]) );
  XNOR U4841 ( .A(n3521), .B(n3520), .Z(z[110]) );
  NANDN U4842 ( .A(n3523), .B(n3522), .Z(n3524) );
  XNOR U4843 ( .A(n3525), .B(n3524), .Z(n3552) );
  XNOR U4844 ( .A(n3526), .B(n3552), .Z(n3527) );
  XOR U4845 ( .A(n3528), .B(n3527), .Z(n3540) );
  XOR U4846 ( .A(n3540), .B(n3529), .Z(z[112]) );
  ANDN U4847 ( .B(n3531), .A(n3530), .Z(n3536) );
  NANDN U4848 ( .A(n3533), .B(n3532), .Z(n3550) );
  XNOR U4849 ( .A(n3534), .B(n3550), .Z(n3535) );
  XOR U4850 ( .A(n3536), .B(n3535), .Z(n3555) );
  XOR U4851 ( .A(n3538), .B(n3537), .Z(n3539) );
  XOR U4852 ( .A(n3555), .B(n3539), .Z(z[115]) );
  XNOR U4853 ( .A(n3540), .B(z[114]), .Z(z[116]) );
  XNOR U4854 ( .A(n3542), .B(n3541), .Z(n3543) );
  XNOR U4855 ( .A(n3544), .B(n3543), .Z(n3554) );
  XNOR U4856 ( .A(n3546), .B(n3545), .Z(n3547) );
  NANDN U4857 ( .A(n3548), .B(n3547), .Z(n3549) );
  XOR U4858 ( .A(n3550), .B(n3549), .Z(n3551) );
  XNOR U4859 ( .A(n3552), .B(n3551), .Z(n3553) );
  XNOR U4860 ( .A(n3554), .B(n3553), .Z(z[117]) );
  XNOR U4861 ( .A(n3556), .B(n3555), .Z(z[118]) );
  NOR U4862 ( .A(n3558), .B(n3557), .Z(n3571) );
  XNOR U4863 ( .A(n3560), .B(n3559), .Z(n3637) );
  OR U4864 ( .A(n3561), .B(n3637), .Z(n3562) );
  XOR U4865 ( .A(n3571), .B(n3562), .Z(n3656) );
  XNOR U4866 ( .A(n3564), .B(n3563), .Z(n3623) );
  ANDN U4867 ( .B(n3565), .A(n3623), .Z(n3579) );
  NOR U4868 ( .A(n3566), .B(n3568), .Z(n3573) );
  NANDN U4869 ( .A(n3567), .B(n3581), .Z(n3649) );
  XOR U4870 ( .A(n3633), .B(n3568), .Z(n3647) );
  XNOR U4871 ( .A(n3581), .B(n3647), .Z(n3582) );
  OR U4872 ( .A(n3582), .B(n3569), .Z(n3570) );
  XNOR U4873 ( .A(n3649), .B(n3570), .Z(n3643) );
  XOR U4874 ( .A(n3571), .B(n3643), .Z(n3572) );
  XOR U4875 ( .A(n3573), .B(n3572), .Z(n3655) );
  XOR U4876 ( .A(n3575), .B(n3574), .Z(n3576) );
  NANDN U4877 ( .A(n3577), .B(n3576), .Z(n3635) );
  XNOR U4878 ( .A(n3655), .B(n3635), .Z(n3578) );
  XOR U4879 ( .A(n3579), .B(n3578), .Z(n3652) );
  XOR U4880 ( .A(n3656), .B(n3652), .Z(n3587) );
  NAND U4881 ( .A(n3581), .B(n3580), .Z(n3627) );
  OR U4882 ( .A(n3583), .B(n3582), .Z(n3584) );
  XNOR U4883 ( .A(n3627), .B(n3584), .Z(n3651) );
  XNOR U4884 ( .A(n3651), .B(n3585), .Z(n3586) );
  XOR U4885 ( .A(n3587), .B(n3586), .Z(z[11]) );
  NANDN U4886 ( .A(n3589), .B(n3588), .Z(n3590) );
  XNOR U4887 ( .A(n3591), .B(n3590), .Z(n3618) );
  XNOR U4888 ( .A(n3592), .B(n3618), .Z(n3593) );
  XOR U4889 ( .A(n3594), .B(n3593), .Z(n3606) );
  XOR U4890 ( .A(n3606), .B(n3595), .Z(z[120]) );
  ANDN U4891 ( .B(n3597), .A(n3596), .Z(n3602) );
  NANDN U4892 ( .A(n3599), .B(n3598), .Z(n3616) );
  XNOR U4893 ( .A(n3600), .B(n3616), .Z(n3601) );
  XOR U4894 ( .A(n3602), .B(n3601), .Z(n3621) );
  XOR U4895 ( .A(n3604), .B(n3603), .Z(n3605) );
  XOR U4896 ( .A(n3621), .B(n3605), .Z(z[123]) );
  XNOR U4897 ( .A(n3606), .B(z[122]), .Z(z[124]) );
  XNOR U4898 ( .A(n3608), .B(n3607), .Z(n3609) );
  XNOR U4899 ( .A(n3610), .B(n3609), .Z(n3620) );
  XNOR U4900 ( .A(n3612), .B(n3611), .Z(n3613) );
  NANDN U4901 ( .A(n3614), .B(n3613), .Z(n3615) );
  XOR U4902 ( .A(n3616), .B(n3615), .Z(n3617) );
  XNOR U4903 ( .A(n3618), .B(n3617), .Z(n3619) );
  XNOR U4904 ( .A(n3620), .B(n3619), .Z(z[125]) );
  XNOR U4905 ( .A(n3622), .B(n3621), .Z(z[126]) );
  ANDN U4906 ( .B(n3624), .A(n3623), .Z(n3630) );
  NAND U4907 ( .A(n3647), .B(n3625), .Z(n3626) );
  XNOR U4908 ( .A(n3627), .B(n3626), .Z(n3639) );
  XNOR U4909 ( .A(n3628), .B(n3639), .Z(n3629) );
  XOR U4910 ( .A(n3630), .B(n3629), .Z(n4008) );
  XNOR U4911 ( .A(n4008), .B(z[10]), .Z(z[12]) );
  XOR U4912 ( .A(x[9]), .B(n3631), .Z(n3632) );
  NANDN U4913 ( .A(n3633), .B(n3632), .Z(n3634) );
  XOR U4914 ( .A(n3635), .B(n3634), .Z(n3636) );
  XNOR U4915 ( .A(n4008), .B(n3636), .Z(n3645) );
  NOR U4916 ( .A(n3638), .B(n3637), .Z(n3642) );
  XOR U4917 ( .A(n3640), .B(n3639), .Z(n3641) );
  XOR U4918 ( .A(n3642), .B(n3641), .Z(n3657) );
  XNOR U4919 ( .A(n3643), .B(n3657), .Z(n3644) );
  XOR U4920 ( .A(n3645), .B(n3644), .Z(z[13]) );
  AND U4921 ( .A(n3647), .B(n3646), .Z(n3648) );
  XNOR U4922 ( .A(n3649), .B(n3648), .Z(n3654) );
  XNOR U4923 ( .A(n3651), .B(n3650), .Z(n4009) );
  XNOR U4924 ( .A(n3652), .B(n4009), .Z(n3653) );
  XOR U4925 ( .A(n3654), .B(n3653), .Z(z[14]) );
  XNOR U4926 ( .A(n3657), .B(z[9]), .Z(z[15]) );
  NANDN U4927 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U4928 ( .A(n3661), .B(n3660), .Z(n3688) );
  XNOR U4929 ( .A(n3662), .B(n3688), .Z(n3663) );
  XOR U4930 ( .A(n3664), .B(n3663), .Z(n3676) );
  XOR U4931 ( .A(n3676), .B(n3665), .Z(z[16]) );
  ANDN U4932 ( .B(n3667), .A(n3666), .Z(n3672) );
  NANDN U4933 ( .A(n3669), .B(n3668), .Z(n3686) );
  XNOR U4934 ( .A(n3670), .B(n3686), .Z(n3671) );
  XOR U4935 ( .A(n3672), .B(n3671), .Z(n3691) );
  XOR U4936 ( .A(n3674), .B(n3673), .Z(n3675) );
  XOR U4937 ( .A(n3691), .B(n3675), .Z(z[19]) );
  XNOR U4938 ( .A(n3676), .B(z[18]), .Z(z[20]) );
  XNOR U4939 ( .A(n3678), .B(n3677), .Z(n3679) );
  XNOR U4940 ( .A(n3680), .B(n3679), .Z(n3690) );
  XNOR U4941 ( .A(n3682), .B(n3681), .Z(n3683) );
  NANDN U4942 ( .A(n3684), .B(n3683), .Z(n3685) );
  XOR U4943 ( .A(n3686), .B(n3685), .Z(n3687) );
  XNOR U4944 ( .A(n3688), .B(n3687), .Z(n3689) );
  XNOR U4945 ( .A(n3690), .B(n3689), .Z(z[21]) );
  XNOR U4946 ( .A(n3692), .B(n3691), .Z(z[22]) );
  NANDN U4947 ( .A(n3694), .B(n3693), .Z(n3695) );
  XNOR U4948 ( .A(n3696), .B(n3695), .Z(n3723) );
  XNOR U4949 ( .A(n3697), .B(n3723), .Z(n3698) );
  XOR U4950 ( .A(n3699), .B(n3698), .Z(n3711) );
  XOR U4951 ( .A(n3711), .B(n3700), .Z(z[24]) );
  ANDN U4952 ( .B(n3702), .A(n3701), .Z(n3707) );
  NANDN U4953 ( .A(n3704), .B(n3703), .Z(n3721) );
  XNOR U4954 ( .A(n3705), .B(n3721), .Z(n3706) );
  XOR U4955 ( .A(n3707), .B(n3706), .Z(n3726) );
  XOR U4956 ( .A(n3709), .B(n3708), .Z(n3710) );
  XOR U4957 ( .A(n3726), .B(n3710), .Z(z[27]) );
  XNOR U4958 ( .A(n3711), .B(z[26]), .Z(z[28]) );
  XNOR U4959 ( .A(n3713), .B(n3712), .Z(n3714) );
  XNOR U4960 ( .A(n3715), .B(n3714), .Z(n3725) );
  XNOR U4961 ( .A(n3717), .B(n3716), .Z(n3718) );
  NANDN U4962 ( .A(n3719), .B(n3718), .Z(n3720) );
  XOR U4963 ( .A(n3721), .B(n3720), .Z(n3722) );
  XNOR U4964 ( .A(n3723), .B(n3722), .Z(n3724) );
  XNOR U4965 ( .A(n3725), .B(n3724), .Z(z[29]) );
  XNOR U4966 ( .A(n3727), .B(n3726), .Z(z[30]) );
  NANDN U4967 ( .A(n3729), .B(n3728), .Z(n3730) );
  XNOR U4968 ( .A(n3731), .B(n3730), .Z(n3758) );
  XNOR U4969 ( .A(n3732), .B(n3758), .Z(n3733) );
  XOR U4970 ( .A(n3734), .B(n3733), .Z(n3746) );
  XOR U4971 ( .A(n3746), .B(n3735), .Z(z[32]) );
  ANDN U4972 ( .B(n3737), .A(n3736), .Z(n3742) );
  NANDN U4973 ( .A(n3739), .B(n3738), .Z(n3756) );
  XNOR U4974 ( .A(n3740), .B(n3756), .Z(n3741) );
  XOR U4975 ( .A(n3742), .B(n3741), .Z(n3761) );
  XOR U4976 ( .A(n3744), .B(n3743), .Z(n3745) );
  XOR U4977 ( .A(n3761), .B(n3745), .Z(z[35]) );
  XNOR U4978 ( .A(n3746), .B(z[34]), .Z(z[36]) );
  XNOR U4979 ( .A(n3748), .B(n3747), .Z(n3749) );
  XNOR U4980 ( .A(n3750), .B(n3749), .Z(n3760) );
  XNOR U4981 ( .A(n3752), .B(n3751), .Z(n3753) );
  NANDN U4982 ( .A(n3754), .B(n3753), .Z(n3755) );
  XOR U4983 ( .A(n3756), .B(n3755), .Z(n3757) );
  XNOR U4984 ( .A(n3758), .B(n3757), .Z(n3759) );
  XNOR U4985 ( .A(n3760), .B(n3759), .Z(z[37]) );
  XNOR U4986 ( .A(n3762), .B(n3761), .Z(z[38]) );
  ANDN U4987 ( .B(n3764), .A(n3763), .Z(n3769) );
  NANDN U4988 ( .A(n3766), .B(n3765), .Z(n3871) );
  XNOR U4989 ( .A(n3767), .B(n3871), .Z(n3768) );
  XOR U4990 ( .A(n3769), .B(n3768), .Z(n3926) );
  XOR U4991 ( .A(n3771), .B(n3770), .Z(n3772) );
  XOR U4992 ( .A(n3926), .B(n3772), .Z(z[3]) );
  NANDN U4993 ( .A(n3774), .B(n3773), .Z(n3775) );
  XNOR U4994 ( .A(n3776), .B(n3775), .Z(n3803) );
  XNOR U4995 ( .A(n3777), .B(n3803), .Z(n3778) );
  XOR U4996 ( .A(n3779), .B(n3778), .Z(n3791) );
  XOR U4997 ( .A(n3791), .B(n3780), .Z(z[40]) );
  ANDN U4998 ( .B(n3782), .A(n3781), .Z(n3787) );
  NANDN U4999 ( .A(n3784), .B(n3783), .Z(n3801) );
  XNOR U5000 ( .A(n3785), .B(n3801), .Z(n3786) );
  XOR U5001 ( .A(n3787), .B(n3786), .Z(n3806) );
  XOR U5002 ( .A(n3789), .B(n3788), .Z(n3790) );
  XOR U5003 ( .A(n3806), .B(n3790), .Z(z[43]) );
  XNOR U5004 ( .A(n3791), .B(z[42]), .Z(z[44]) );
  XNOR U5005 ( .A(n3793), .B(n3792), .Z(n3794) );
  XNOR U5006 ( .A(n3795), .B(n3794), .Z(n3805) );
  XNOR U5007 ( .A(n3797), .B(n3796), .Z(n3798) );
  NANDN U5008 ( .A(n3799), .B(n3798), .Z(n3800) );
  XOR U5009 ( .A(n3801), .B(n3800), .Z(n3802) );
  XNOR U5010 ( .A(n3803), .B(n3802), .Z(n3804) );
  XNOR U5011 ( .A(n3805), .B(n3804), .Z(z[45]) );
  XNOR U5012 ( .A(n3807), .B(n3806), .Z(z[46]) );
  NANDN U5013 ( .A(n3809), .B(n3808), .Z(n3810) );
  XNOR U5014 ( .A(n3811), .B(n3810), .Z(n3839) );
  XNOR U5015 ( .A(n3812), .B(n3839), .Z(n3813) );
  XOR U5016 ( .A(n3814), .B(n3813), .Z(n3827) );
  XOR U5017 ( .A(n3827), .B(n3815), .Z(z[48]) );
  XNOR U5018 ( .A(n3816), .B(z[2]), .Z(z[4]) );
  ANDN U5019 ( .B(n3818), .A(n3817), .Z(n3823) );
  NANDN U5020 ( .A(n3820), .B(n3819), .Z(n3837) );
  XNOR U5021 ( .A(n3821), .B(n3837), .Z(n3822) );
  XOR U5022 ( .A(n3823), .B(n3822), .Z(n3842) );
  XOR U5023 ( .A(n3825), .B(n3824), .Z(n3826) );
  XOR U5024 ( .A(n3842), .B(n3826), .Z(z[51]) );
  XNOR U5025 ( .A(n3827), .B(z[50]), .Z(z[52]) );
  XNOR U5026 ( .A(n3829), .B(n3828), .Z(n3830) );
  XNOR U5027 ( .A(n3831), .B(n3830), .Z(n3841) );
  XNOR U5028 ( .A(n3833), .B(n3832), .Z(n3834) );
  NANDN U5029 ( .A(n3835), .B(n3834), .Z(n3836) );
  XOR U5030 ( .A(n3837), .B(n3836), .Z(n3838) );
  XNOR U5031 ( .A(n3839), .B(n3838), .Z(n3840) );
  XNOR U5032 ( .A(n3841), .B(n3840), .Z(z[53]) );
  XNOR U5033 ( .A(n3843), .B(n3842), .Z(z[54]) );
  NANDN U5034 ( .A(n3845), .B(n3844), .Z(n3846) );
  XNOR U5035 ( .A(n3847), .B(n3846), .Z(n3888) );
  XNOR U5036 ( .A(n3848), .B(n3888), .Z(n3849) );
  XOR U5037 ( .A(n3850), .B(n3849), .Z(n3876) );
  XOR U5038 ( .A(n3876), .B(n3851), .Z(z[56]) );
  ANDN U5039 ( .B(n3853), .A(n3852), .Z(n3858) );
  NANDN U5040 ( .A(n3855), .B(n3854), .Z(n3886) );
  XNOR U5041 ( .A(n3856), .B(n3886), .Z(n3857) );
  XOR U5042 ( .A(n3858), .B(n3857), .Z(n3891) );
  XOR U5043 ( .A(n3860), .B(n3859), .Z(n3861) );
  XOR U5044 ( .A(n3891), .B(n3861), .Z(z[59]) );
  XNOR U5045 ( .A(n3863), .B(n3862), .Z(n3864) );
  XNOR U5046 ( .A(n3865), .B(n3864), .Z(n3875) );
  XNOR U5047 ( .A(n3867), .B(n3866), .Z(n3868) );
  NANDN U5048 ( .A(n3869), .B(n3868), .Z(n3870) );
  XOR U5049 ( .A(n3871), .B(n3870), .Z(n3872) );
  XNOR U5050 ( .A(n3873), .B(n3872), .Z(n3874) );
  XNOR U5051 ( .A(n3875), .B(n3874), .Z(z[5]) );
  XNOR U5052 ( .A(n3876), .B(z[58]), .Z(z[60]) );
  XNOR U5053 ( .A(n3878), .B(n3877), .Z(n3879) );
  XNOR U5054 ( .A(n3880), .B(n3879), .Z(n3890) );
  XNOR U5055 ( .A(n3882), .B(n3881), .Z(n3883) );
  NANDN U5056 ( .A(n3884), .B(n3883), .Z(n3885) );
  XOR U5057 ( .A(n3886), .B(n3885), .Z(n3887) );
  XNOR U5058 ( .A(n3888), .B(n3887), .Z(n3889) );
  XNOR U5059 ( .A(n3890), .B(n3889), .Z(z[61]) );
  XNOR U5060 ( .A(n3892), .B(n3891), .Z(z[62]) );
  NANDN U5061 ( .A(n3894), .B(n3893), .Z(n3895) );
  XNOR U5062 ( .A(n3896), .B(n3895), .Z(n3923) );
  XNOR U5063 ( .A(n3897), .B(n3923), .Z(n3898) );
  XOR U5064 ( .A(n3899), .B(n3898), .Z(n3911) );
  XOR U5065 ( .A(n3911), .B(n3900), .Z(z[64]) );
  ANDN U5066 ( .B(n3902), .A(n3901), .Z(n3907) );
  NANDN U5067 ( .A(n3904), .B(n3903), .Z(n3921) );
  XNOR U5068 ( .A(n3905), .B(n3921), .Z(n3906) );
  XOR U5069 ( .A(n3907), .B(n3906), .Z(n3928) );
  XOR U5070 ( .A(n3909), .B(n3908), .Z(n3910) );
  XOR U5071 ( .A(n3928), .B(n3910), .Z(z[67]) );
  XNOR U5072 ( .A(n3911), .B(z[66]), .Z(z[68]) );
  XNOR U5073 ( .A(n3913), .B(n3912), .Z(n3914) );
  XNOR U5074 ( .A(n3915), .B(n3914), .Z(n3925) );
  XNOR U5075 ( .A(n3917), .B(n3916), .Z(n3918) );
  NANDN U5076 ( .A(n3919), .B(n3918), .Z(n3920) );
  XOR U5077 ( .A(n3921), .B(n3920), .Z(n3922) );
  XNOR U5078 ( .A(n3923), .B(n3922), .Z(n3924) );
  XNOR U5079 ( .A(n3925), .B(n3924), .Z(z[69]) );
  XNOR U5080 ( .A(n3927), .B(n3926), .Z(z[6]) );
  XNOR U5081 ( .A(n3929), .B(n3928), .Z(z[70]) );
  NANDN U5082 ( .A(n3931), .B(n3930), .Z(n3932) );
  XNOR U5083 ( .A(n3933), .B(n3932), .Z(n3960) );
  XNOR U5084 ( .A(n3934), .B(n3960), .Z(n3935) );
  XOR U5085 ( .A(n3936), .B(n3935), .Z(n3948) );
  XOR U5086 ( .A(n3948), .B(n3937), .Z(z[72]) );
  ANDN U5087 ( .B(n3939), .A(n3938), .Z(n3944) );
  NANDN U5088 ( .A(n3941), .B(n3940), .Z(n3958) );
  XNOR U5089 ( .A(n3942), .B(n3958), .Z(n3943) );
  XOR U5090 ( .A(n3944), .B(n3943), .Z(n3963) );
  XOR U5091 ( .A(n3946), .B(n3945), .Z(n3947) );
  XOR U5092 ( .A(n3963), .B(n3947), .Z(z[75]) );
  XNOR U5093 ( .A(n3948), .B(z[74]), .Z(z[76]) );
  XNOR U5094 ( .A(n3950), .B(n3949), .Z(n3951) );
  XNOR U5095 ( .A(n3952), .B(n3951), .Z(n3962) );
  XNOR U5096 ( .A(n3954), .B(n3953), .Z(n3955) );
  NANDN U5097 ( .A(n3956), .B(n3955), .Z(n3957) );
  XOR U5098 ( .A(n3958), .B(n3957), .Z(n3959) );
  XNOR U5099 ( .A(n3960), .B(n3959), .Z(n3961) );
  XNOR U5100 ( .A(n3962), .B(n3961), .Z(z[77]) );
  XNOR U5101 ( .A(n3964), .B(n3963), .Z(z[78]) );
  NANDN U5102 ( .A(n3966), .B(n3965), .Z(n3967) );
  XNOR U5103 ( .A(n3968), .B(n3967), .Z(n3995) );
  XNOR U5104 ( .A(n3969), .B(n3995), .Z(n3970) );
  XOR U5105 ( .A(n3971), .B(n3970), .Z(n3983) );
  XOR U5106 ( .A(n3983), .B(n3972), .Z(z[80]) );
  ANDN U5107 ( .B(n3974), .A(n3973), .Z(n3979) );
  NANDN U5108 ( .A(n3976), .B(n3975), .Z(n3993) );
  XNOR U5109 ( .A(n3977), .B(n3993), .Z(n3978) );
  XOR U5110 ( .A(n3979), .B(n3978), .Z(n3998) );
  XOR U5111 ( .A(n3981), .B(n3980), .Z(n3982) );
  XOR U5112 ( .A(n3998), .B(n3982), .Z(z[83]) );
  XNOR U5113 ( .A(n3983), .B(z[82]), .Z(z[84]) );
  XNOR U5114 ( .A(n3985), .B(n3984), .Z(n3986) );
  XNOR U5115 ( .A(n3987), .B(n3986), .Z(n3997) );
  XNOR U5116 ( .A(n3989), .B(n3988), .Z(n3990) );
  NANDN U5117 ( .A(n3991), .B(n3990), .Z(n3992) );
  XOR U5118 ( .A(n3993), .B(n3992), .Z(n3994) );
  XNOR U5119 ( .A(n3995), .B(n3994), .Z(n3996) );
  XNOR U5120 ( .A(n3997), .B(n3996), .Z(z[85]) );
  XNOR U5121 ( .A(n3999), .B(n3998), .Z(z[86]) );
  NANDN U5122 ( .A(n4001), .B(n4000), .Z(n4002) );
  XNOR U5123 ( .A(n4003), .B(n4002), .Z(n4032) );
  XNOR U5124 ( .A(n4004), .B(n4032), .Z(n4005) );
  XOR U5125 ( .A(n4006), .B(n4005), .Z(n4020) );
  XOR U5126 ( .A(n4020), .B(n4007), .Z(z[88]) );
  XNOR U5127 ( .A(n4009), .B(n4008), .Z(z[8]) );
  ANDN U5128 ( .B(n4011), .A(n4010), .Z(n4016) );
  NANDN U5129 ( .A(n4013), .B(n4012), .Z(n4030) );
  XNOR U5130 ( .A(n4014), .B(n4030), .Z(n4015) );
  XOR U5131 ( .A(n4016), .B(n4015), .Z(n4035) );
  XOR U5132 ( .A(n4018), .B(n4017), .Z(n4019) );
  XOR U5133 ( .A(n4035), .B(n4019), .Z(z[91]) );
  XNOR U5134 ( .A(n4020), .B(z[90]), .Z(z[92]) );
  XNOR U5135 ( .A(n4022), .B(n4021), .Z(n4023) );
  XNOR U5136 ( .A(n4024), .B(n4023), .Z(n4034) );
  XNOR U5137 ( .A(n4026), .B(n4025), .Z(n4027) );
  NANDN U5138 ( .A(n4028), .B(n4027), .Z(n4029) );
  XOR U5139 ( .A(n4030), .B(n4029), .Z(n4031) );
  XNOR U5140 ( .A(n4032), .B(n4031), .Z(n4033) );
  XNOR U5141 ( .A(n4034), .B(n4033), .Z(z[93]) );
  XNOR U5142 ( .A(n4036), .B(n4035), .Z(z[94]) );
  XNOR U5143 ( .A(n4038), .B(n4037), .Z(z[96]) );
  XOR U5144 ( .A(n4040), .B(n4039), .Z(n4041) );
  XOR U5145 ( .A(n4042), .B(n4041), .Z(z[99]) );
endmodule


module SubBytes_1 ( x, z );
  input [127:0] x;
  output [127:0] z;
  wire   n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
         n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
         n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
         n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
         n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036,
         n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
         n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
         n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
         n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076,
         n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
         n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
         n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
         n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
         n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
         n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
         n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
         n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
         n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
         n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
         n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
         n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196,
         n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
         n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
         n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
         n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236,
         n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
         n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
         n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
         n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276,
         n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
         n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
         n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
         n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
         n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
         n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
         n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
         n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356,
         n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
         n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
         n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
         n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396,
         n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
         n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436,
         n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
         n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
         n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
         n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
         n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
         n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
         n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
         n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516,
         n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
         n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
         n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
         n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
         n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
         n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
         n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
         n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
         n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
         n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
         n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906,
         n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916,
         n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
         n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936,
         n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
         n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976,
         n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986,
         n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996,
         n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042;

  XNOR U2962 ( .A(x[103]), .B(x[98]), .Z(n3465) );
  XOR U2963 ( .A(n3623), .B(n3637), .Z(n3581) );
  XNOR U2964 ( .A(n2145), .B(n2148), .Z(n2168) );
  ANDN U2965 ( .B(n3729), .A(n3737), .Z(n1987) );
  XNOR U2966 ( .A(n2379), .B(n2383), .Z(n1988) );
  XNOR U2967 ( .A(n1987), .B(n1988), .Z(n2406) );
  ANDN U2968 ( .B(n3931), .A(n3939), .Z(n1989) );
  XNOR U2969 ( .A(n2839), .B(n2843), .Z(n1990) );
  XNOR U2970 ( .A(n1989), .B(n1990), .Z(n2866) );
  ANDN U2971 ( .B(n3523), .A(n3531), .Z(n1991) );
  XNOR U2972 ( .A(n3258), .B(n3262), .Z(n1992) );
  XNOR U2973 ( .A(n1991), .B(n1992), .Z(n3285) );
  ANDN U2974 ( .B(n3694), .A(n3702), .Z(n1993) );
  XNOR U2975 ( .A(n2287), .B(n2291), .Z(n1994) );
  XNOR U2976 ( .A(n1993), .B(n1994), .Z(n2314) );
  ANDN U2977 ( .B(n3894), .A(n3902), .Z(n1995) );
  XNOR U2978 ( .A(n2747), .B(n2751), .Z(n1996) );
  XNOR U2979 ( .A(n1995), .B(n1996), .Z(n2774) );
  ANDN U2980 ( .B(n3488), .A(n3496), .Z(n1997) );
  XNOR U2981 ( .A(n3166), .B(n3170), .Z(n1998) );
  XNOR U2982 ( .A(n1997), .B(n1998), .Z(n3193) );
  ANDN U2983 ( .B(n3659), .A(n3667), .Z(n1999) );
  XNOR U2984 ( .A(n2195), .B(n2199), .Z(n2000) );
  XNOR U2985 ( .A(n1999), .B(n2000), .Z(n2222) );
  ANDN U2986 ( .B(n3845), .A(n3853), .Z(n2001) );
  XNOR U2987 ( .A(n2655), .B(n2659), .Z(n2002) );
  XNOR U2988 ( .A(n2001), .B(n2002), .Z(n2682) );
  XNOR U2989 ( .A(n3567), .B(n2116), .Z(n2167) );
  ANDN U2990 ( .B(n3809), .A(n3818), .Z(n2003) );
  XNOR U2991 ( .A(n2563), .B(n2567), .Z(n2004) );
  XNOR U2992 ( .A(n2003), .B(n2004), .Z(n2590) );
  ANDN U2993 ( .B(n3421), .A(n3764), .Z(n2005) );
  XNOR U2994 ( .A(n2046), .B(n2050), .Z(n2006) );
  XNOR U2995 ( .A(n2005), .B(n2006), .Z(n2073) );
  ANDN U2996 ( .B(n3774), .A(n3782), .Z(n2007) );
  XNOR U2997 ( .A(n2471), .B(n2475), .Z(n2008) );
  XNOR U2998 ( .A(n2007), .B(n2008), .Z(n2498) );
  ANDN U2999 ( .B(n3589), .A(n3597), .Z(n2009) );
  XNOR U3000 ( .A(n3350), .B(n3354), .Z(n2010) );
  XNOR U3001 ( .A(n2009), .B(n2010), .Z(n3377) );
  XOR U3002 ( .A(x[98]), .B(n3084), .Z(n2011) );
  XNOR U3003 ( .A(n3083), .B(n2011), .Z(n3430) );
  XNOR U3004 ( .A(n3471), .B(n3463), .Z(n3444) );
  NAND U3005 ( .A(n3029), .B(n3050), .Z(n2012) );
  OR U3006 ( .A(n3076), .B(n3050), .Z(n2013) );
  NAND U3007 ( .A(n2012), .B(n2013), .Z(n2014) );
  XNOR U3008 ( .A(n3065), .B(n2014), .Z(n2015) );
  XOR U3009 ( .A(n3019), .B(n3006), .Z(n2016) );
  XNOR U3010 ( .A(n2015), .B(n2016), .Z(n3044) );
  NAND U3011 ( .A(n2942), .B(n2963), .Z(n2017) );
  OR U3012 ( .A(n2989), .B(n2963), .Z(n2018) );
  NAND U3013 ( .A(n2017), .B(n2018), .Z(n2019) );
  XNOR U3014 ( .A(n2978), .B(n2019), .Z(n2020) );
  XOR U3015 ( .A(n2932), .B(n2919), .Z(n2021) );
  XNOR U3016 ( .A(n2020), .B(n2021), .Z(n2957) );
  XOR U3017 ( .A(n3655), .B(n3654), .Z(n2022) );
  XNOR U3018 ( .A(z[10]), .B(n3656), .Z(n2023) );
  XNOR U3019 ( .A(n2022), .B(n2023), .Z(z[9]) );
  IV U3020 ( .A(x[4]), .Z(n2024) );
  IV U3021 ( .A(x[0]), .Z(n2109) );
  XOR U3022 ( .A(n2109), .B(x[6]), .Z(n2025) );
  XOR U3023 ( .A(n2025), .B(x[5]), .Z(n2049) );
  IV U3024 ( .A(n2049), .Z(n3867) );
  XOR U3025 ( .A(n2024), .B(n3867), .Z(n2098) );
  XOR U3026 ( .A(x[1]), .B(x[3]), .Z(n2026) );
  XOR U3027 ( .A(x[7]), .B(n2024), .Z(n2084) );
  XNOR U3028 ( .A(n2026), .B(n2084), .Z(n2063) );
  IV U3029 ( .A(n2063), .Z(n2041) );
  XOR U3030 ( .A(n2026), .B(n2025), .Z(n2027) );
  XOR U3031 ( .A(x[2]), .B(n2027), .Z(n3421) );
  XOR U3032 ( .A(n3421), .B(n2049), .Z(n2081) );
  XOR U3033 ( .A(n2041), .B(n2081), .Z(n2094) );
  IV U3034 ( .A(x[2]), .Z(n2037) );
  XOR U3035 ( .A(x[4]), .B(n2037), .Z(n2086) );
  NOR U3036 ( .A(n2094), .B(n2086), .Z(n2029) );
  XOR U3037 ( .A(x[7]), .B(n3867), .Z(n3764) );
  XOR U3038 ( .A(n3421), .B(n3764), .Z(n2028) );
  XNOR U3039 ( .A(n2029), .B(n2028), .Z(n2030) );
  XNOR U3040 ( .A(n2109), .B(n3421), .Z(n2093) );
  NOR U3041 ( .A(n2084), .B(n2093), .Z(n2039) );
  XNOR U3042 ( .A(n2030), .B(n2039), .Z(n2051) );
  IV U3043 ( .A(x[1]), .Z(n3866) );
  XNOR U3044 ( .A(n3866), .B(x[2]), .Z(n2031) );
  XNOR U3045 ( .A(n3764), .B(n2031), .Z(n2083) );
  ANDN U3046 ( .B(n2083), .A(x[0]), .Z(n2032) );
  XNOR U3047 ( .A(n2084), .B(n2031), .Z(n2088) );
  NANDN U3048 ( .A(n2041), .B(n2088), .Z(n2042) );
  XOR U3049 ( .A(n2032), .B(n2042), .Z(n2034) );
  OR U3050 ( .A(n2083), .B(n2063), .Z(n2033) );
  NAND U3051 ( .A(n2034), .B(n2033), .Z(n2035) );
  XOR U3052 ( .A(n2051), .B(n2035), .Z(n2036) );
  XOR U3053 ( .A(n2098), .B(n2036), .Z(n2077) );
  XNOR U3054 ( .A(n2041), .B(x[0]), .Z(n2064) );
  XNOR U3055 ( .A(n3867), .B(n2064), .Z(n2111) );
  IV U3056 ( .A(x[7]), .Z(n2040) );
  XOR U3057 ( .A(n2040), .B(n2037), .Z(n2103) );
  NANDN U3058 ( .A(n2111), .B(n2103), .Z(n2038) );
  XOR U3059 ( .A(n2039), .B(n2038), .Z(n2046) );
  XOR U3060 ( .A(n3866), .B(n2040), .Z(n3765) );
  NAND U3061 ( .A(n2081), .B(n3765), .Z(n2050) );
  ANDN U3062 ( .B(n2098), .A(n2109), .Z(n2044) );
  XNOR U3063 ( .A(n2042), .B(n2041), .Z(n2043) );
  XNOR U3064 ( .A(n2044), .B(n2043), .Z(n2045) );
  XNOR U3065 ( .A(n2046), .B(n2045), .Z(n2048) );
  XNOR U3066 ( .A(x[2]), .B(n3764), .Z(n2047) );
  XNOR U3067 ( .A(n2048), .B(n2047), .Z(n2078) );
  IV U3068 ( .A(n2078), .Z(n2070) );
  AND U3069 ( .A(n2073), .B(n2070), .Z(n2066) );
  XOR U3070 ( .A(n2077), .B(n2066), .Z(n2054) );
  ANDN U3071 ( .B(n2049), .A(x[1]), .Z(n2053) );
  XNOR U3072 ( .A(n2051), .B(n2050), .Z(n2052) );
  XNOR U3073 ( .A(n2053), .B(n2052), .Z(n2072) );
  ANDN U3074 ( .B(n2054), .A(n2072), .Z(n2061) );
  IV U3075 ( .A(n2073), .Z(n2058) );
  NANDN U3076 ( .A(n2058), .B(n2072), .Z(n2055) );
  NANDN U3077 ( .A(n2061), .B(n2055), .Z(n2085) );
  NANDN U3078 ( .A(n2073), .B(n2070), .Z(n2056) );
  NAND U3079 ( .A(n2056), .B(n2072), .Z(n2060) );
  XNOR U3080 ( .A(n2070), .B(n2077), .Z(n2057) );
  NANDN U3081 ( .A(n2058), .B(n2057), .Z(n2059) );
  AND U3082 ( .A(n2060), .B(n2059), .Z(n2110) );
  OR U3083 ( .A(n2085), .B(n2110), .Z(n2062) );
  ANDN U3084 ( .B(n2062), .A(n2061), .Z(n2089) );
  NANDN U3085 ( .A(n2089), .B(n2063), .Z(n3863) );
  NANDN U3086 ( .A(n2085), .B(n2064), .Z(n2065) );
  XOR U3087 ( .A(n3863), .B(n2065), .Z(n2097) );
  NANDN U3088 ( .A(n2070), .B(n2077), .Z(n2069) );
  XNOR U3089 ( .A(n2066), .B(n2072), .Z(n2067) );
  NANDN U3090 ( .A(n2077), .B(n2067), .Z(n2068) );
  AND U3091 ( .A(n2069), .B(n2068), .Z(n3869) );
  NANDN U3092 ( .A(n2070), .B(n2073), .Z(n2071) );
  NAND U3093 ( .A(n2077), .B(n2071), .Z(n2076) );
  XNOR U3094 ( .A(n2073), .B(n2072), .Z(n2074) );
  NANDN U3095 ( .A(n2078), .B(n2074), .Z(n2075) );
  NAND U3096 ( .A(n2076), .B(n2075), .Z(n3763) );
  IV U3097 ( .A(n3763), .Z(n3420) );
  NANDN U3098 ( .A(n3869), .B(n3420), .Z(n2080) );
  NANDN U3099 ( .A(n2078), .B(n2077), .Z(n2079) );
  NAND U3100 ( .A(n2080), .B(n2079), .Z(n3766) );
  NANDN U3101 ( .A(n3766), .B(n2081), .Z(n3423) );
  NANDN U3102 ( .A(n3869), .B(n3867), .Z(n2082) );
  XNOR U3103 ( .A(n3423), .B(n2082), .Z(n2099) );
  XOR U3104 ( .A(n2097), .B(n2099), .Z(z[2]) );
  NOR U3105 ( .A(n2085), .B(n2083), .Z(n2091) );
  XOR U3106 ( .A(n3420), .B(n2110), .Z(n2092) );
  NANDN U3107 ( .A(n2084), .B(n2092), .Z(n2105) );
  XOR U3108 ( .A(n2085), .B(n3869), .Z(n2112) );
  XNOR U3109 ( .A(n2092), .B(n2112), .Z(n2095) );
  OR U3110 ( .A(n2086), .B(n2095), .Z(n2087) );
  XNOR U3111 ( .A(n2105), .B(n2087), .Z(n3862) );
  NANDN U3112 ( .A(n2089), .B(n2088), .Z(n2100) );
  XNOR U3113 ( .A(n3862), .B(n2100), .Z(n2090) );
  XOR U3114 ( .A(n2091), .B(n2090), .Z(n3771) );
  NANDN U3115 ( .A(n2093), .B(n2092), .Z(n3424) );
  OR U3116 ( .A(n2095), .B(n2094), .Z(n2096) );
  XOR U3117 ( .A(n3424), .B(n2096), .Z(n2106) );
  XOR U3118 ( .A(n2106), .B(n2097), .Z(n3427) );
  XOR U3119 ( .A(n3771), .B(n3427), .Z(n3927) );
  ANDN U3120 ( .B(n2110), .A(n2098), .Z(n2102) );
  XNOR U3121 ( .A(n2100), .B(n2099), .Z(n2101) );
  XNOR U3122 ( .A(n2102), .B(n2101), .Z(n2108) );
  NAND U3123 ( .A(n2103), .B(n2112), .Z(n2104) );
  XNOR U3124 ( .A(n2105), .B(n2104), .Z(n3767) );
  XOR U3125 ( .A(n2106), .B(n3767), .Z(n2107) );
  XOR U3126 ( .A(n2108), .B(n2107), .Z(n3770) );
  XNOR U3127 ( .A(n3927), .B(n3770), .Z(z[1]) );
  ANDN U3128 ( .B(n2110), .A(n2109), .Z(n3865) );
  ANDN U3129 ( .B(n2112), .A(n2111), .Z(n3426) );
  XNOR U3130 ( .A(n3424), .B(z[1]), .Z(n2113) );
  XNOR U3131 ( .A(n3426), .B(n2113), .Z(n2114) );
  XOR U3132 ( .A(n3863), .B(n2114), .Z(n2115) );
  XOR U3133 ( .A(n3865), .B(n2115), .Z(z[7]) );
  IV U3134 ( .A(x[9]), .Z(n3575) );
  IV U3135 ( .A(x[8]), .Z(n3638) );
  XNOR U3136 ( .A(x[14]), .B(n3638), .Z(n2121) );
  XOR U3137 ( .A(x[13]), .B(n2121), .Z(n3631) );
  ANDN U3138 ( .B(n3575), .A(n3631), .Z(n2118) );
  XNOR U3139 ( .A(x[12]), .B(x[15]), .Z(n3567) );
  XOR U3140 ( .A(x[11]), .B(x[9]), .Z(n2116) );
  XNOR U3141 ( .A(x[10]), .B(n2116), .Z(n2142) );
  XNOR U3142 ( .A(x[14]), .B(n2142), .Z(n3580) );
  NANDN U3143 ( .A(n3567), .B(n3580), .Z(n2120) );
  IV U3144 ( .A(x[12]), .Z(n2123) );
  XOR U3145 ( .A(x[10]), .B(n2123), .Z(n3569) );
  XOR U3146 ( .A(n3638), .B(n2167), .Z(n2171) );
  IV U3147 ( .A(n3631), .Z(n2161) );
  XOR U3148 ( .A(n2171), .B(n2161), .Z(n3625) );
  XNOR U3149 ( .A(n3580), .B(n3625), .Z(n3583) );
  OR U3150 ( .A(n3569), .B(n3583), .Z(n2117) );
  XOR U3151 ( .A(n2120), .B(n2117), .Z(n2137) );
  XNOR U3152 ( .A(n2118), .B(n2137), .Z(n2145) );
  IV U3153 ( .A(x[10]), .Z(n2124) );
  IV U3154 ( .A(x[15]), .Z(n3574) );
  XOR U3155 ( .A(n2124), .B(n3574), .Z(n3646) );
  NAND U3156 ( .A(n3625), .B(n3646), .Z(n2119) );
  XNOR U3157 ( .A(n2120), .B(n2119), .Z(n2128) );
  XOR U3158 ( .A(x[15]), .B(n3631), .Z(n3565) );
  XNOR U3159 ( .A(n2142), .B(n2121), .Z(n3624) );
  NAND U3160 ( .A(n3565), .B(n3624), .Z(n2122) );
  XOR U3161 ( .A(n2128), .B(n2122), .Z(n2148) );
  XNOR U3162 ( .A(n2123), .B(n2161), .Z(n3561) );
  NOR U3163 ( .A(n3638), .B(n3561), .Z(n2130) );
  XNOR U3164 ( .A(n2124), .B(x[9]), .Z(n2131) );
  XOR U3165 ( .A(n3567), .B(n2131), .Z(n3558) );
  NANDN U3166 ( .A(n3558), .B(n2167), .Z(n2132) );
  XNOR U3167 ( .A(n2132), .B(n3565), .Z(n2126) );
  XNOR U3168 ( .A(n2124), .B(n2171), .Z(n2125) );
  XNOR U3169 ( .A(n2126), .B(n2125), .Z(n2127) );
  XOR U3170 ( .A(n2128), .B(n2127), .Z(n2129) );
  XNOR U3171 ( .A(n2130), .B(n2129), .Z(n2157) );
  IV U3172 ( .A(n2157), .Z(n2147) );
  NANDN U3173 ( .A(n2168), .B(n2147), .Z(n2141) );
  XNOR U3174 ( .A(n2131), .B(n3565), .Z(n3566) );
  ANDN U3175 ( .B(n3566), .A(x[8]), .Z(n2133) );
  XOR U3176 ( .A(n2133), .B(n2132), .Z(n2135) );
  OR U3177 ( .A(n2167), .B(n3566), .Z(n2134) );
  NAND U3178 ( .A(n2135), .B(n2134), .Z(n2136) );
  XOR U3179 ( .A(n3624), .B(n2136), .Z(n2139) );
  XOR U3180 ( .A(n3567), .B(n2137), .Z(n2138) );
  XNOR U3181 ( .A(n2139), .B(n2138), .Z(n2158) );
  IV U3182 ( .A(n2158), .Z(n2154) );
  NANDN U3183 ( .A(n2154), .B(n2168), .Z(n2140) );
  NAND U3184 ( .A(n2141), .B(n2140), .Z(n2150) );
  XOR U3185 ( .A(x[13]), .B(n2142), .Z(n2153) );
  NANDN U3186 ( .A(n2153), .B(n3575), .Z(n2144) );
  NANDN U3187 ( .A(n3574), .B(n2153), .Z(n2143) );
  AND U3188 ( .A(n2144), .B(n2143), .Z(n2149) );
  XOR U3189 ( .A(n2149), .B(n2145), .Z(n2166) );
  IV U3190 ( .A(n2166), .Z(n2151) );
  ANDN U3191 ( .B(n2151), .A(n2154), .Z(n2146) );
  XOR U3192 ( .A(n2150), .B(n2146), .Z(n2164) );
  OR U3193 ( .A(n2164), .B(n2147), .Z(n3564) );
  XOR U3194 ( .A(n2149), .B(n2148), .Z(n2163) );
  NANDN U3195 ( .A(n2157), .B(n2163), .Z(n2156) );
  XNOR U3196 ( .A(n2151), .B(n2150), .Z(n2152) );
  XNOR U3197 ( .A(n2156), .B(n2152), .Z(n2165) );
  ANDN U3198 ( .B(n2154), .A(n2165), .Z(n2160) );
  XOR U3199 ( .A(n3564), .B(n2160), .Z(n3577) );
  OR U3200 ( .A(n3577), .B(n2153), .Z(n3628) );
  ANDN U3201 ( .B(n2154), .A(n2166), .Z(n2155) );
  XNOR U3202 ( .A(n2156), .B(n2155), .Z(n2169) );
  XNOR U3203 ( .A(n2158), .B(n2157), .Z(n2159) );
  NANDN U3204 ( .A(n2169), .B(n2159), .Z(n3563) );
  XOR U3205 ( .A(n3563), .B(n2160), .Z(n3633) );
  OR U3206 ( .A(n3633), .B(n2161), .Z(n2162) );
  XNOR U3207 ( .A(n3628), .B(n2162), .Z(n3585) );
  OR U3208 ( .A(n2164), .B(n2163), .Z(n3559) );
  NOR U3209 ( .A(n2166), .B(n2165), .Z(n2170) );
  XOR U3210 ( .A(n3559), .B(n2170), .Z(n3557) );
  ANDN U3211 ( .B(n2167), .A(n3557), .Z(n3640) );
  OR U3212 ( .A(n2169), .B(n2168), .Z(n3560) );
  XOR U3213 ( .A(n3560), .B(n2170), .Z(n3568) );
  OR U3214 ( .A(n3568), .B(n2171), .Z(n2172) );
  XOR U3215 ( .A(n3640), .B(n2172), .Z(n3650) );
  XNOR U3216 ( .A(n3585), .B(n3650), .Z(z[10]) );
  IV U3217 ( .A(x[20]), .Z(n2173) );
  IV U3218 ( .A(x[16]), .Z(n2258) );
  XOR U3219 ( .A(n2258), .B(x[22]), .Z(n2174) );
  XOR U3220 ( .A(n2174), .B(x[21]), .Z(n2198) );
  IV U3221 ( .A(n2198), .Z(n3682) );
  XOR U3222 ( .A(n2173), .B(n3682), .Z(n2247) );
  XOR U3223 ( .A(x[17]), .B(x[19]), .Z(n2175) );
  XOR U3224 ( .A(x[23]), .B(n2173), .Z(n2233) );
  XNOR U3225 ( .A(n2175), .B(n2233), .Z(n2212) );
  IV U3226 ( .A(n2212), .Z(n2190) );
  XOR U3227 ( .A(n2175), .B(n2174), .Z(n2176) );
  XOR U3228 ( .A(x[18]), .B(n2176), .Z(n3659) );
  XOR U3229 ( .A(n3659), .B(n2198), .Z(n2230) );
  XOR U3230 ( .A(n2190), .B(n2230), .Z(n2243) );
  IV U3231 ( .A(x[18]), .Z(n2186) );
  XOR U3232 ( .A(x[20]), .B(n2186), .Z(n2235) );
  NOR U3233 ( .A(n2243), .B(n2235), .Z(n2178) );
  XOR U3234 ( .A(x[23]), .B(n3682), .Z(n3667) );
  XOR U3235 ( .A(n3659), .B(n3667), .Z(n2177) );
  XNOR U3236 ( .A(n2178), .B(n2177), .Z(n2179) );
  XNOR U3237 ( .A(n2258), .B(n3659), .Z(n2242) );
  NOR U3238 ( .A(n2233), .B(n2242), .Z(n2188) );
  XNOR U3239 ( .A(n2179), .B(n2188), .Z(n2200) );
  IV U3240 ( .A(x[17]), .Z(n3681) );
  XNOR U3241 ( .A(n3681), .B(x[18]), .Z(n2180) );
  XNOR U3242 ( .A(n3667), .B(n2180), .Z(n2232) );
  ANDN U3243 ( .B(n2232), .A(x[16]), .Z(n2181) );
  XNOR U3244 ( .A(n2233), .B(n2180), .Z(n2237) );
  NANDN U3245 ( .A(n2190), .B(n2237), .Z(n2191) );
  XOR U3246 ( .A(n2181), .B(n2191), .Z(n2183) );
  OR U3247 ( .A(n2232), .B(n2212), .Z(n2182) );
  NAND U3248 ( .A(n2183), .B(n2182), .Z(n2184) );
  XOR U3249 ( .A(n2200), .B(n2184), .Z(n2185) );
  XOR U3250 ( .A(n2247), .B(n2185), .Z(n2226) );
  XNOR U3251 ( .A(n2190), .B(x[16]), .Z(n2213) );
  XNOR U3252 ( .A(n3682), .B(n2213), .Z(n2260) );
  IV U3253 ( .A(x[23]), .Z(n2189) );
  XOR U3254 ( .A(n2189), .B(n2186), .Z(n2252) );
  NANDN U3255 ( .A(n2260), .B(n2252), .Z(n2187) );
  XOR U3256 ( .A(n2188), .B(n2187), .Z(n2195) );
  XOR U3257 ( .A(n3681), .B(n2189), .Z(n3668) );
  NAND U3258 ( .A(n2230), .B(n3668), .Z(n2199) );
  ANDN U3259 ( .B(n2247), .A(n2258), .Z(n2193) );
  XNOR U3260 ( .A(n2191), .B(n2190), .Z(n2192) );
  XNOR U3261 ( .A(n2193), .B(n2192), .Z(n2194) );
  XNOR U3262 ( .A(n2195), .B(n2194), .Z(n2197) );
  XNOR U3263 ( .A(x[18]), .B(n3667), .Z(n2196) );
  XNOR U3264 ( .A(n2197), .B(n2196), .Z(n2227) );
  IV U3265 ( .A(n2227), .Z(n2219) );
  AND U3266 ( .A(n2222), .B(n2219), .Z(n2215) );
  XOR U3267 ( .A(n2226), .B(n2215), .Z(n2203) );
  ANDN U3268 ( .B(n2198), .A(x[17]), .Z(n2202) );
  XNOR U3269 ( .A(n2200), .B(n2199), .Z(n2201) );
  XNOR U3270 ( .A(n2202), .B(n2201), .Z(n2221) );
  ANDN U3271 ( .B(n2203), .A(n2221), .Z(n2210) );
  IV U3272 ( .A(n2222), .Z(n2207) );
  NANDN U3273 ( .A(n2207), .B(n2221), .Z(n2204) );
  NANDN U3274 ( .A(n2210), .B(n2204), .Z(n2234) );
  NANDN U3275 ( .A(n2222), .B(n2219), .Z(n2205) );
  NAND U3276 ( .A(n2205), .B(n2221), .Z(n2209) );
  XNOR U3277 ( .A(n2219), .B(n2226), .Z(n2206) );
  NANDN U3278 ( .A(n2207), .B(n2206), .Z(n2208) );
  AND U3279 ( .A(n2209), .B(n2208), .Z(n2259) );
  OR U3280 ( .A(n2234), .B(n2259), .Z(n2211) );
  ANDN U3281 ( .B(n2211), .A(n2210), .Z(n2238) );
  NANDN U3282 ( .A(n2238), .B(n2212), .Z(n3678) );
  NANDN U3283 ( .A(n2234), .B(n2213), .Z(n2214) );
  XOR U3284 ( .A(n3678), .B(n2214), .Z(n2246) );
  NANDN U3285 ( .A(n2219), .B(n2226), .Z(n2218) );
  XNOR U3286 ( .A(n2215), .B(n2221), .Z(n2216) );
  NANDN U3287 ( .A(n2226), .B(n2216), .Z(n2217) );
  AND U3288 ( .A(n2218), .B(n2217), .Z(n3684) );
  NANDN U3289 ( .A(n2219), .B(n2222), .Z(n2220) );
  NAND U3290 ( .A(n2226), .B(n2220), .Z(n2225) );
  XNOR U3291 ( .A(n2222), .B(n2221), .Z(n2223) );
  NANDN U3292 ( .A(n2227), .B(n2223), .Z(n2224) );
  NAND U3293 ( .A(n2225), .B(n2224), .Z(n3666) );
  IV U3294 ( .A(n3666), .Z(n3658) );
  NANDN U3295 ( .A(n3684), .B(n3658), .Z(n2229) );
  NANDN U3296 ( .A(n2227), .B(n2226), .Z(n2228) );
  NAND U3297 ( .A(n2229), .B(n2228), .Z(n3669) );
  NANDN U3298 ( .A(n3669), .B(n2230), .Z(n3661) );
  NANDN U3299 ( .A(n3684), .B(n3682), .Z(n2231) );
  XNOR U3300 ( .A(n3661), .B(n2231), .Z(n2248) );
  XOR U3301 ( .A(n2246), .B(n2248), .Z(z[18]) );
  NOR U3302 ( .A(n2234), .B(n2232), .Z(n2240) );
  XOR U3303 ( .A(n3658), .B(n2259), .Z(n2241) );
  NANDN U3304 ( .A(n2233), .B(n2241), .Z(n2254) );
  XOR U3305 ( .A(n2234), .B(n3684), .Z(n2261) );
  XNOR U3306 ( .A(n2241), .B(n2261), .Z(n2244) );
  OR U3307 ( .A(n2235), .B(n2244), .Z(n2236) );
  XNOR U3308 ( .A(n2254), .B(n2236), .Z(n3677) );
  NANDN U3309 ( .A(n2238), .B(n2237), .Z(n2249) );
  XNOR U3310 ( .A(n3677), .B(n2249), .Z(n2239) );
  XOR U3311 ( .A(n2240), .B(n2239), .Z(n3674) );
  NANDN U3312 ( .A(n2242), .B(n2241), .Z(n3662) );
  OR U3313 ( .A(n2244), .B(n2243), .Z(n2245) );
  XOR U3314 ( .A(n3662), .B(n2245), .Z(n2255) );
  XOR U3315 ( .A(n2255), .B(n2246), .Z(n3665) );
  XOR U3316 ( .A(n3674), .B(n3665), .Z(n3692) );
  ANDN U3317 ( .B(n2259), .A(n2247), .Z(n2251) );
  XNOR U3318 ( .A(n2249), .B(n2248), .Z(n2250) );
  XNOR U3319 ( .A(n2251), .B(n2250), .Z(n2257) );
  NAND U3320 ( .A(n2252), .B(n2261), .Z(n2253) );
  XNOR U3321 ( .A(n2254), .B(n2253), .Z(n3670) );
  XOR U3322 ( .A(n2255), .B(n3670), .Z(n2256) );
  XOR U3323 ( .A(n2257), .B(n2256), .Z(n3673) );
  XNOR U3324 ( .A(n3692), .B(n3673), .Z(z[17]) );
  ANDN U3325 ( .B(n2259), .A(n2258), .Z(n3680) );
  ANDN U3326 ( .B(n2261), .A(n2260), .Z(n3664) );
  XNOR U3327 ( .A(n3662), .B(z[17]), .Z(n2262) );
  XNOR U3328 ( .A(n3664), .B(n2262), .Z(n2263) );
  XOR U3329 ( .A(n3678), .B(n2263), .Z(n2264) );
  XOR U3330 ( .A(n3680), .B(n2264), .Z(z[23]) );
  IV U3331 ( .A(x[28]), .Z(n2265) );
  IV U3332 ( .A(x[24]), .Z(n2350) );
  XOR U3333 ( .A(n2350), .B(x[30]), .Z(n2266) );
  XOR U3334 ( .A(n2266), .B(x[29]), .Z(n2290) );
  IV U3335 ( .A(n2290), .Z(n3717) );
  XOR U3336 ( .A(n2265), .B(n3717), .Z(n2339) );
  XOR U3337 ( .A(x[25]), .B(x[27]), .Z(n2267) );
  XOR U3338 ( .A(x[31]), .B(n2265), .Z(n2325) );
  XNOR U3339 ( .A(n2267), .B(n2325), .Z(n2304) );
  IV U3340 ( .A(n2304), .Z(n2282) );
  XOR U3341 ( .A(n2267), .B(n2266), .Z(n2268) );
  XOR U3342 ( .A(x[26]), .B(n2268), .Z(n3694) );
  XOR U3343 ( .A(n3694), .B(n2290), .Z(n2322) );
  XOR U3344 ( .A(n2282), .B(n2322), .Z(n2335) );
  IV U3345 ( .A(x[26]), .Z(n2278) );
  XOR U3346 ( .A(x[28]), .B(n2278), .Z(n2327) );
  NOR U3347 ( .A(n2335), .B(n2327), .Z(n2270) );
  XOR U3348 ( .A(x[31]), .B(n3717), .Z(n3702) );
  XOR U3349 ( .A(n3694), .B(n3702), .Z(n2269) );
  XNOR U3350 ( .A(n2270), .B(n2269), .Z(n2271) );
  XNOR U3351 ( .A(n2350), .B(n3694), .Z(n2334) );
  NOR U3352 ( .A(n2325), .B(n2334), .Z(n2280) );
  XNOR U3353 ( .A(n2271), .B(n2280), .Z(n2292) );
  IV U3354 ( .A(x[25]), .Z(n3716) );
  XNOR U3355 ( .A(n3716), .B(x[26]), .Z(n2272) );
  XNOR U3356 ( .A(n3702), .B(n2272), .Z(n2324) );
  ANDN U3357 ( .B(n2324), .A(x[24]), .Z(n2273) );
  XNOR U3358 ( .A(n2325), .B(n2272), .Z(n2329) );
  NANDN U3359 ( .A(n2282), .B(n2329), .Z(n2283) );
  XOR U3360 ( .A(n2273), .B(n2283), .Z(n2275) );
  OR U3361 ( .A(n2324), .B(n2304), .Z(n2274) );
  NAND U3362 ( .A(n2275), .B(n2274), .Z(n2276) );
  XOR U3363 ( .A(n2292), .B(n2276), .Z(n2277) );
  XOR U3364 ( .A(n2339), .B(n2277), .Z(n2318) );
  XNOR U3365 ( .A(n2282), .B(x[24]), .Z(n2305) );
  XNOR U3366 ( .A(n3717), .B(n2305), .Z(n2352) );
  IV U3367 ( .A(x[31]), .Z(n2281) );
  XOR U3368 ( .A(n2281), .B(n2278), .Z(n2344) );
  NANDN U3369 ( .A(n2352), .B(n2344), .Z(n2279) );
  XOR U3370 ( .A(n2280), .B(n2279), .Z(n2287) );
  XOR U3371 ( .A(n3716), .B(n2281), .Z(n3703) );
  NAND U3372 ( .A(n2322), .B(n3703), .Z(n2291) );
  ANDN U3373 ( .B(n2339), .A(n2350), .Z(n2285) );
  XNOR U3374 ( .A(n2283), .B(n2282), .Z(n2284) );
  XNOR U3375 ( .A(n2285), .B(n2284), .Z(n2286) );
  XNOR U3376 ( .A(n2287), .B(n2286), .Z(n2289) );
  XNOR U3377 ( .A(x[26]), .B(n3702), .Z(n2288) );
  XNOR U3378 ( .A(n2289), .B(n2288), .Z(n2319) );
  IV U3379 ( .A(n2319), .Z(n2311) );
  AND U3380 ( .A(n2314), .B(n2311), .Z(n2307) );
  XOR U3381 ( .A(n2318), .B(n2307), .Z(n2295) );
  ANDN U3382 ( .B(n2290), .A(x[25]), .Z(n2294) );
  XNOR U3383 ( .A(n2292), .B(n2291), .Z(n2293) );
  XNOR U3384 ( .A(n2294), .B(n2293), .Z(n2313) );
  ANDN U3385 ( .B(n2295), .A(n2313), .Z(n2302) );
  IV U3386 ( .A(n2314), .Z(n2299) );
  NANDN U3387 ( .A(n2299), .B(n2313), .Z(n2296) );
  NANDN U3388 ( .A(n2302), .B(n2296), .Z(n2326) );
  NANDN U3389 ( .A(n2314), .B(n2311), .Z(n2297) );
  NAND U3390 ( .A(n2297), .B(n2313), .Z(n2301) );
  XNOR U3391 ( .A(n2311), .B(n2318), .Z(n2298) );
  NANDN U3392 ( .A(n2299), .B(n2298), .Z(n2300) );
  AND U3393 ( .A(n2301), .B(n2300), .Z(n2351) );
  OR U3394 ( .A(n2326), .B(n2351), .Z(n2303) );
  ANDN U3395 ( .B(n2303), .A(n2302), .Z(n2330) );
  NANDN U3396 ( .A(n2330), .B(n2304), .Z(n3713) );
  NANDN U3397 ( .A(n2326), .B(n2305), .Z(n2306) );
  XOR U3398 ( .A(n3713), .B(n2306), .Z(n2338) );
  NANDN U3399 ( .A(n2311), .B(n2318), .Z(n2310) );
  XNOR U3400 ( .A(n2307), .B(n2313), .Z(n2308) );
  NANDN U3401 ( .A(n2318), .B(n2308), .Z(n2309) );
  AND U3402 ( .A(n2310), .B(n2309), .Z(n3719) );
  NANDN U3403 ( .A(n2311), .B(n2314), .Z(n2312) );
  NAND U3404 ( .A(n2318), .B(n2312), .Z(n2317) );
  XNOR U3405 ( .A(n2314), .B(n2313), .Z(n2315) );
  NANDN U3406 ( .A(n2319), .B(n2315), .Z(n2316) );
  NAND U3407 ( .A(n2317), .B(n2316), .Z(n3701) );
  IV U3408 ( .A(n3701), .Z(n3693) );
  NANDN U3409 ( .A(n3719), .B(n3693), .Z(n2321) );
  NANDN U3410 ( .A(n2319), .B(n2318), .Z(n2320) );
  NAND U3411 ( .A(n2321), .B(n2320), .Z(n3704) );
  NANDN U3412 ( .A(n3704), .B(n2322), .Z(n3696) );
  NANDN U3413 ( .A(n3719), .B(n3717), .Z(n2323) );
  XNOR U3414 ( .A(n3696), .B(n2323), .Z(n2340) );
  XOR U3415 ( .A(n2338), .B(n2340), .Z(z[26]) );
  NOR U3416 ( .A(n2326), .B(n2324), .Z(n2332) );
  XOR U3417 ( .A(n3693), .B(n2351), .Z(n2333) );
  NANDN U3418 ( .A(n2325), .B(n2333), .Z(n2346) );
  XOR U3419 ( .A(n2326), .B(n3719), .Z(n2353) );
  XNOR U3420 ( .A(n2333), .B(n2353), .Z(n2336) );
  OR U3421 ( .A(n2327), .B(n2336), .Z(n2328) );
  XNOR U3422 ( .A(n2346), .B(n2328), .Z(n3712) );
  NANDN U3423 ( .A(n2330), .B(n2329), .Z(n2341) );
  XNOR U3424 ( .A(n3712), .B(n2341), .Z(n2331) );
  XOR U3425 ( .A(n2332), .B(n2331), .Z(n3709) );
  NANDN U3426 ( .A(n2334), .B(n2333), .Z(n3697) );
  OR U3427 ( .A(n2336), .B(n2335), .Z(n2337) );
  XOR U3428 ( .A(n3697), .B(n2337), .Z(n2347) );
  XOR U3429 ( .A(n2347), .B(n2338), .Z(n3700) );
  XOR U3430 ( .A(n3709), .B(n3700), .Z(n3727) );
  ANDN U3431 ( .B(n2351), .A(n2339), .Z(n2343) );
  XNOR U3432 ( .A(n2341), .B(n2340), .Z(n2342) );
  XNOR U3433 ( .A(n2343), .B(n2342), .Z(n2349) );
  NAND U3434 ( .A(n2344), .B(n2353), .Z(n2345) );
  XNOR U3435 ( .A(n2346), .B(n2345), .Z(n3705) );
  XOR U3436 ( .A(n2347), .B(n3705), .Z(n2348) );
  XOR U3437 ( .A(n2349), .B(n2348), .Z(n3708) );
  XNOR U3438 ( .A(n3727), .B(n3708), .Z(z[25]) );
  ANDN U3439 ( .B(n2351), .A(n2350), .Z(n3715) );
  ANDN U3440 ( .B(n2353), .A(n2352), .Z(n3699) );
  XNOR U3441 ( .A(n3697), .B(z[25]), .Z(n2354) );
  XNOR U3442 ( .A(n3699), .B(n2354), .Z(n2355) );
  XOR U3443 ( .A(n3713), .B(n2355), .Z(n2356) );
  XOR U3444 ( .A(n3715), .B(n2356), .Z(z[31]) );
  IV U3445 ( .A(x[36]), .Z(n2357) );
  IV U3446 ( .A(x[32]), .Z(n2442) );
  XOR U3447 ( .A(n2442), .B(x[38]), .Z(n2358) );
  XOR U3448 ( .A(n2358), .B(x[37]), .Z(n2382) );
  IV U3449 ( .A(n2382), .Z(n3752) );
  XOR U3450 ( .A(n2357), .B(n3752), .Z(n2431) );
  XOR U3451 ( .A(x[33]), .B(x[35]), .Z(n2359) );
  XOR U3452 ( .A(x[39]), .B(n2357), .Z(n2417) );
  XNOR U3453 ( .A(n2359), .B(n2417), .Z(n2396) );
  IV U3454 ( .A(n2396), .Z(n2374) );
  XOR U3455 ( .A(n2359), .B(n2358), .Z(n2360) );
  XOR U3456 ( .A(x[34]), .B(n2360), .Z(n3729) );
  XOR U3457 ( .A(n3729), .B(n2382), .Z(n2414) );
  XOR U3458 ( .A(n2374), .B(n2414), .Z(n2427) );
  IV U3459 ( .A(x[34]), .Z(n2370) );
  XOR U3460 ( .A(x[36]), .B(n2370), .Z(n2419) );
  NOR U3461 ( .A(n2427), .B(n2419), .Z(n2362) );
  XOR U3462 ( .A(x[39]), .B(n3752), .Z(n3737) );
  XOR U3463 ( .A(n3729), .B(n3737), .Z(n2361) );
  XNOR U3464 ( .A(n2362), .B(n2361), .Z(n2363) );
  XNOR U3465 ( .A(n2442), .B(n3729), .Z(n2426) );
  NOR U3466 ( .A(n2417), .B(n2426), .Z(n2372) );
  XNOR U3467 ( .A(n2363), .B(n2372), .Z(n2384) );
  IV U3468 ( .A(x[33]), .Z(n3751) );
  XNOR U3469 ( .A(n3751), .B(x[34]), .Z(n2364) );
  XNOR U3470 ( .A(n3737), .B(n2364), .Z(n2416) );
  ANDN U3471 ( .B(n2416), .A(x[32]), .Z(n2365) );
  XNOR U3472 ( .A(n2417), .B(n2364), .Z(n2421) );
  NANDN U3473 ( .A(n2374), .B(n2421), .Z(n2375) );
  XOR U3474 ( .A(n2365), .B(n2375), .Z(n2367) );
  OR U3475 ( .A(n2416), .B(n2396), .Z(n2366) );
  NAND U3476 ( .A(n2367), .B(n2366), .Z(n2368) );
  XOR U3477 ( .A(n2384), .B(n2368), .Z(n2369) );
  XOR U3478 ( .A(n2431), .B(n2369), .Z(n2410) );
  XNOR U3479 ( .A(n2374), .B(x[32]), .Z(n2397) );
  XNOR U3480 ( .A(n3752), .B(n2397), .Z(n2444) );
  IV U3481 ( .A(x[39]), .Z(n2373) );
  XOR U3482 ( .A(n2373), .B(n2370), .Z(n2436) );
  NANDN U3483 ( .A(n2444), .B(n2436), .Z(n2371) );
  XOR U3484 ( .A(n2372), .B(n2371), .Z(n2379) );
  XOR U3485 ( .A(n3751), .B(n2373), .Z(n3738) );
  NAND U3486 ( .A(n2414), .B(n3738), .Z(n2383) );
  ANDN U3487 ( .B(n2431), .A(n2442), .Z(n2377) );
  XNOR U3488 ( .A(n2375), .B(n2374), .Z(n2376) );
  XNOR U3489 ( .A(n2377), .B(n2376), .Z(n2378) );
  XNOR U3490 ( .A(n2379), .B(n2378), .Z(n2381) );
  XNOR U3491 ( .A(x[34]), .B(n3737), .Z(n2380) );
  XNOR U3492 ( .A(n2381), .B(n2380), .Z(n2411) );
  IV U3493 ( .A(n2411), .Z(n2403) );
  AND U3494 ( .A(n2406), .B(n2403), .Z(n2399) );
  XOR U3495 ( .A(n2410), .B(n2399), .Z(n2387) );
  ANDN U3496 ( .B(n2382), .A(x[33]), .Z(n2386) );
  XNOR U3497 ( .A(n2384), .B(n2383), .Z(n2385) );
  XNOR U3498 ( .A(n2386), .B(n2385), .Z(n2405) );
  ANDN U3499 ( .B(n2387), .A(n2405), .Z(n2394) );
  IV U3500 ( .A(n2406), .Z(n2391) );
  NANDN U3501 ( .A(n2391), .B(n2405), .Z(n2388) );
  NANDN U3502 ( .A(n2394), .B(n2388), .Z(n2418) );
  NANDN U3503 ( .A(n2406), .B(n2403), .Z(n2389) );
  NAND U3504 ( .A(n2389), .B(n2405), .Z(n2393) );
  XNOR U3505 ( .A(n2403), .B(n2410), .Z(n2390) );
  NANDN U3506 ( .A(n2391), .B(n2390), .Z(n2392) );
  AND U3507 ( .A(n2393), .B(n2392), .Z(n2443) );
  OR U3508 ( .A(n2418), .B(n2443), .Z(n2395) );
  ANDN U3509 ( .B(n2395), .A(n2394), .Z(n2422) );
  NANDN U3510 ( .A(n2422), .B(n2396), .Z(n3748) );
  NANDN U3511 ( .A(n2418), .B(n2397), .Z(n2398) );
  XOR U3512 ( .A(n3748), .B(n2398), .Z(n2430) );
  NANDN U3513 ( .A(n2403), .B(n2410), .Z(n2402) );
  XNOR U3514 ( .A(n2399), .B(n2405), .Z(n2400) );
  NANDN U3515 ( .A(n2410), .B(n2400), .Z(n2401) );
  AND U3516 ( .A(n2402), .B(n2401), .Z(n3754) );
  NANDN U3517 ( .A(n2403), .B(n2406), .Z(n2404) );
  NAND U3518 ( .A(n2410), .B(n2404), .Z(n2409) );
  XNOR U3519 ( .A(n2406), .B(n2405), .Z(n2407) );
  NANDN U3520 ( .A(n2411), .B(n2407), .Z(n2408) );
  NAND U3521 ( .A(n2409), .B(n2408), .Z(n3736) );
  IV U3522 ( .A(n3736), .Z(n3728) );
  NANDN U3523 ( .A(n3754), .B(n3728), .Z(n2413) );
  NANDN U3524 ( .A(n2411), .B(n2410), .Z(n2412) );
  NAND U3525 ( .A(n2413), .B(n2412), .Z(n3739) );
  NANDN U3526 ( .A(n3739), .B(n2414), .Z(n3731) );
  NANDN U3527 ( .A(n3754), .B(n3752), .Z(n2415) );
  XNOR U3528 ( .A(n3731), .B(n2415), .Z(n2432) );
  XOR U3529 ( .A(n2430), .B(n2432), .Z(z[34]) );
  NOR U3530 ( .A(n2418), .B(n2416), .Z(n2424) );
  XOR U3531 ( .A(n3728), .B(n2443), .Z(n2425) );
  NANDN U3532 ( .A(n2417), .B(n2425), .Z(n2438) );
  XOR U3533 ( .A(n2418), .B(n3754), .Z(n2445) );
  XNOR U3534 ( .A(n2425), .B(n2445), .Z(n2428) );
  OR U3535 ( .A(n2419), .B(n2428), .Z(n2420) );
  XNOR U3536 ( .A(n2438), .B(n2420), .Z(n3747) );
  NANDN U3537 ( .A(n2422), .B(n2421), .Z(n2433) );
  XNOR U3538 ( .A(n3747), .B(n2433), .Z(n2423) );
  XOR U3539 ( .A(n2424), .B(n2423), .Z(n3744) );
  NANDN U3540 ( .A(n2426), .B(n2425), .Z(n3732) );
  OR U3541 ( .A(n2428), .B(n2427), .Z(n2429) );
  XOR U3542 ( .A(n3732), .B(n2429), .Z(n2439) );
  XOR U3543 ( .A(n2439), .B(n2430), .Z(n3735) );
  XOR U3544 ( .A(n3744), .B(n3735), .Z(n3762) );
  ANDN U3545 ( .B(n2443), .A(n2431), .Z(n2435) );
  XNOR U3546 ( .A(n2433), .B(n2432), .Z(n2434) );
  XNOR U3547 ( .A(n2435), .B(n2434), .Z(n2441) );
  NAND U3548 ( .A(n2436), .B(n2445), .Z(n2437) );
  XNOR U3549 ( .A(n2438), .B(n2437), .Z(n3740) );
  XOR U3550 ( .A(n2439), .B(n3740), .Z(n2440) );
  XOR U3551 ( .A(n2441), .B(n2440), .Z(n3743) );
  XNOR U3552 ( .A(n3762), .B(n3743), .Z(z[33]) );
  ANDN U3553 ( .B(n2443), .A(n2442), .Z(n3750) );
  ANDN U3554 ( .B(n2445), .A(n2444), .Z(n3734) );
  XNOR U3555 ( .A(n3732), .B(z[33]), .Z(n2446) );
  XNOR U3556 ( .A(n3734), .B(n2446), .Z(n2447) );
  XOR U3557 ( .A(n3748), .B(n2447), .Z(n2448) );
  XOR U3558 ( .A(n3750), .B(n2448), .Z(z[39]) );
  IV U3559 ( .A(x[44]), .Z(n2449) );
  IV U3560 ( .A(x[40]), .Z(n2534) );
  XOR U3561 ( .A(n2534), .B(x[46]), .Z(n2450) );
  XOR U3562 ( .A(n2450), .B(x[45]), .Z(n2474) );
  IV U3563 ( .A(n2474), .Z(n3797) );
  XOR U3564 ( .A(n2449), .B(n3797), .Z(n2523) );
  XOR U3565 ( .A(x[41]), .B(x[43]), .Z(n2451) );
  XOR U3566 ( .A(x[47]), .B(n2449), .Z(n2509) );
  XNOR U3567 ( .A(n2451), .B(n2509), .Z(n2488) );
  IV U3568 ( .A(n2488), .Z(n2466) );
  XOR U3569 ( .A(n2451), .B(n2450), .Z(n2452) );
  XOR U3570 ( .A(x[42]), .B(n2452), .Z(n3774) );
  XOR U3571 ( .A(n3774), .B(n2474), .Z(n2506) );
  XOR U3572 ( .A(n2466), .B(n2506), .Z(n2519) );
  IV U3573 ( .A(x[42]), .Z(n2462) );
  XOR U3574 ( .A(x[44]), .B(n2462), .Z(n2511) );
  NOR U3575 ( .A(n2519), .B(n2511), .Z(n2454) );
  XOR U3576 ( .A(x[47]), .B(n3797), .Z(n3782) );
  XOR U3577 ( .A(n3774), .B(n3782), .Z(n2453) );
  XNOR U3578 ( .A(n2454), .B(n2453), .Z(n2455) );
  XNOR U3579 ( .A(n2534), .B(n3774), .Z(n2518) );
  NOR U3580 ( .A(n2509), .B(n2518), .Z(n2464) );
  XNOR U3581 ( .A(n2455), .B(n2464), .Z(n2476) );
  IV U3582 ( .A(x[41]), .Z(n3796) );
  XNOR U3583 ( .A(n3796), .B(x[42]), .Z(n2456) );
  XNOR U3584 ( .A(n3782), .B(n2456), .Z(n2508) );
  ANDN U3585 ( .B(n2508), .A(x[40]), .Z(n2457) );
  XNOR U3586 ( .A(n2509), .B(n2456), .Z(n2513) );
  NANDN U3587 ( .A(n2466), .B(n2513), .Z(n2467) );
  XOR U3588 ( .A(n2457), .B(n2467), .Z(n2459) );
  OR U3589 ( .A(n2508), .B(n2488), .Z(n2458) );
  NAND U3590 ( .A(n2459), .B(n2458), .Z(n2460) );
  XOR U3591 ( .A(n2476), .B(n2460), .Z(n2461) );
  XOR U3592 ( .A(n2523), .B(n2461), .Z(n2502) );
  XNOR U3593 ( .A(n2466), .B(x[40]), .Z(n2489) );
  XNOR U3594 ( .A(n3797), .B(n2489), .Z(n2536) );
  IV U3595 ( .A(x[47]), .Z(n2465) );
  XOR U3596 ( .A(n2465), .B(n2462), .Z(n2528) );
  NANDN U3597 ( .A(n2536), .B(n2528), .Z(n2463) );
  XOR U3598 ( .A(n2464), .B(n2463), .Z(n2471) );
  XOR U3599 ( .A(n3796), .B(n2465), .Z(n3783) );
  NAND U3600 ( .A(n2506), .B(n3783), .Z(n2475) );
  ANDN U3601 ( .B(n2523), .A(n2534), .Z(n2469) );
  XNOR U3602 ( .A(n2467), .B(n2466), .Z(n2468) );
  XNOR U3603 ( .A(n2469), .B(n2468), .Z(n2470) );
  XNOR U3604 ( .A(n2471), .B(n2470), .Z(n2473) );
  XNOR U3605 ( .A(x[42]), .B(n3782), .Z(n2472) );
  XNOR U3606 ( .A(n2473), .B(n2472), .Z(n2503) );
  IV U3607 ( .A(n2503), .Z(n2495) );
  AND U3608 ( .A(n2498), .B(n2495), .Z(n2491) );
  XOR U3609 ( .A(n2502), .B(n2491), .Z(n2479) );
  ANDN U3610 ( .B(n2474), .A(x[41]), .Z(n2478) );
  XNOR U3611 ( .A(n2476), .B(n2475), .Z(n2477) );
  XNOR U3612 ( .A(n2478), .B(n2477), .Z(n2497) );
  ANDN U3613 ( .B(n2479), .A(n2497), .Z(n2486) );
  IV U3614 ( .A(n2498), .Z(n2483) );
  NANDN U3615 ( .A(n2483), .B(n2497), .Z(n2480) );
  NANDN U3616 ( .A(n2486), .B(n2480), .Z(n2510) );
  NANDN U3617 ( .A(n2498), .B(n2495), .Z(n2481) );
  NAND U3618 ( .A(n2481), .B(n2497), .Z(n2485) );
  XNOR U3619 ( .A(n2495), .B(n2502), .Z(n2482) );
  NANDN U3620 ( .A(n2483), .B(n2482), .Z(n2484) );
  AND U3621 ( .A(n2485), .B(n2484), .Z(n2535) );
  OR U3622 ( .A(n2510), .B(n2535), .Z(n2487) );
  ANDN U3623 ( .B(n2487), .A(n2486), .Z(n2514) );
  NANDN U3624 ( .A(n2514), .B(n2488), .Z(n3793) );
  NANDN U3625 ( .A(n2510), .B(n2489), .Z(n2490) );
  XOR U3626 ( .A(n3793), .B(n2490), .Z(n2522) );
  NANDN U3627 ( .A(n2495), .B(n2502), .Z(n2494) );
  XNOR U3628 ( .A(n2491), .B(n2497), .Z(n2492) );
  NANDN U3629 ( .A(n2502), .B(n2492), .Z(n2493) );
  AND U3630 ( .A(n2494), .B(n2493), .Z(n3799) );
  NANDN U3631 ( .A(n2495), .B(n2498), .Z(n2496) );
  NAND U3632 ( .A(n2502), .B(n2496), .Z(n2501) );
  XNOR U3633 ( .A(n2498), .B(n2497), .Z(n2499) );
  NANDN U3634 ( .A(n2503), .B(n2499), .Z(n2500) );
  NAND U3635 ( .A(n2501), .B(n2500), .Z(n3781) );
  IV U3636 ( .A(n3781), .Z(n3773) );
  NANDN U3637 ( .A(n3799), .B(n3773), .Z(n2505) );
  NANDN U3638 ( .A(n2503), .B(n2502), .Z(n2504) );
  NAND U3639 ( .A(n2505), .B(n2504), .Z(n3784) );
  NANDN U3640 ( .A(n3784), .B(n2506), .Z(n3776) );
  NANDN U3641 ( .A(n3799), .B(n3797), .Z(n2507) );
  XNOR U3642 ( .A(n3776), .B(n2507), .Z(n2524) );
  XOR U3643 ( .A(n2522), .B(n2524), .Z(z[42]) );
  NOR U3644 ( .A(n2510), .B(n2508), .Z(n2516) );
  XOR U3645 ( .A(n3773), .B(n2535), .Z(n2517) );
  NANDN U3646 ( .A(n2509), .B(n2517), .Z(n2530) );
  XOR U3647 ( .A(n2510), .B(n3799), .Z(n2537) );
  XNOR U3648 ( .A(n2517), .B(n2537), .Z(n2520) );
  OR U3649 ( .A(n2511), .B(n2520), .Z(n2512) );
  XNOR U3650 ( .A(n2530), .B(n2512), .Z(n3792) );
  NANDN U3651 ( .A(n2514), .B(n2513), .Z(n2525) );
  XNOR U3652 ( .A(n3792), .B(n2525), .Z(n2515) );
  XOR U3653 ( .A(n2516), .B(n2515), .Z(n3789) );
  NANDN U3654 ( .A(n2518), .B(n2517), .Z(n3777) );
  OR U3655 ( .A(n2520), .B(n2519), .Z(n2521) );
  XOR U3656 ( .A(n3777), .B(n2521), .Z(n2531) );
  XOR U3657 ( .A(n2531), .B(n2522), .Z(n3780) );
  XOR U3658 ( .A(n3789), .B(n3780), .Z(n3807) );
  ANDN U3659 ( .B(n2535), .A(n2523), .Z(n2527) );
  XNOR U3660 ( .A(n2525), .B(n2524), .Z(n2526) );
  XNOR U3661 ( .A(n2527), .B(n2526), .Z(n2533) );
  NAND U3662 ( .A(n2528), .B(n2537), .Z(n2529) );
  XNOR U3663 ( .A(n2530), .B(n2529), .Z(n3785) );
  XOR U3664 ( .A(n2531), .B(n3785), .Z(n2532) );
  XOR U3665 ( .A(n2533), .B(n2532), .Z(n3788) );
  XNOR U3666 ( .A(n3807), .B(n3788), .Z(z[41]) );
  ANDN U3667 ( .B(n2535), .A(n2534), .Z(n3795) );
  ANDN U3668 ( .B(n2537), .A(n2536), .Z(n3779) );
  XNOR U3669 ( .A(n3777), .B(z[41]), .Z(n2538) );
  XNOR U3670 ( .A(n3779), .B(n2538), .Z(n2539) );
  XOR U3671 ( .A(n3793), .B(n2539), .Z(n2540) );
  XOR U3672 ( .A(n3795), .B(n2540), .Z(z[47]) );
  IV U3673 ( .A(x[52]), .Z(n2541) );
  IV U3674 ( .A(x[48]), .Z(n2626) );
  XOR U3675 ( .A(n2626), .B(x[54]), .Z(n2542) );
  XOR U3676 ( .A(n2542), .B(x[53]), .Z(n2566) );
  IV U3677 ( .A(n2566), .Z(n3833) );
  XOR U3678 ( .A(n2541), .B(n3833), .Z(n2615) );
  XOR U3679 ( .A(x[49]), .B(x[51]), .Z(n2543) );
  XOR U3680 ( .A(x[55]), .B(n2541), .Z(n2601) );
  XNOR U3681 ( .A(n2543), .B(n2601), .Z(n2580) );
  IV U3682 ( .A(n2580), .Z(n2558) );
  XOR U3683 ( .A(n2543), .B(n2542), .Z(n2544) );
  XOR U3684 ( .A(x[50]), .B(n2544), .Z(n3809) );
  XOR U3685 ( .A(n3809), .B(n2566), .Z(n2598) );
  XOR U3686 ( .A(n2558), .B(n2598), .Z(n2611) );
  IV U3687 ( .A(x[50]), .Z(n2554) );
  XOR U3688 ( .A(x[52]), .B(n2554), .Z(n2603) );
  NOR U3689 ( .A(n2611), .B(n2603), .Z(n2546) );
  XOR U3690 ( .A(x[55]), .B(n3833), .Z(n3818) );
  XOR U3691 ( .A(n3809), .B(n3818), .Z(n2545) );
  XNOR U3692 ( .A(n2546), .B(n2545), .Z(n2547) );
  XNOR U3693 ( .A(n2626), .B(n3809), .Z(n2610) );
  NOR U3694 ( .A(n2601), .B(n2610), .Z(n2556) );
  XNOR U3695 ( .A(n2547), .B(n2556), .Z(n2568) );
  IV U3696 ( .A(x[49]), .Z(n3832) );
  XNOR U3697 ( .A(n3832), .B(x[50]), .Z(n2548) );
  XNOR U3698 ( .A(n3818), .B(n2548), .Z(n2600) );
  ANDN U3699 ( .B(n2600), .A(x[48]), .Z(n2549) );
  XNOR U3700 ( .A(n2601), .B(n2548), .Z(n2605) );
  NANDN U3701 ( .A(n2558), .B(n2605), .Z(n2559) );
  XOR U3702 ( .A(n2549), .B(n2559), .Z(n2551) );
  OR U3703 ( .A(n2600), .B(n2580), .Z(n2550) );
  NAND U3704 ( .A(n2551), .B(n2550), .Z(n2552) );
  XOR U3705 ( .A(n2568), .B(n2552), .Z(n2553) );
  XOR U3706 ( .A(n2615), .B(n2553), .Z(n2594) );
  XNOR U3707 ( .A(n2558), .B(x[48]), .Z(n2581) );
  XNOR U3708 ( .A(n3833), .B(n2581), .Z(n2628) );
  IV U3709 ( .A(x[55]), .Z(n2557) );
  XOR U3710 ( .A(n2557), .B(n2554), .Z(n2620) );
  NANDN U3711 ( .A(n2628), .B(n2620), .Z(n2555) );
  XOR U3712 ( .A(n2556), .B(n2555), .Z(n2563) );
  XOR U3713 ( .A(n3832), .B(n2557), .Z(n3819) );
  NAND U3714 ( .A(n2598), .B(n3819), .Z(n2567) );
  ANDN U3715 ( .B(n2615), .A(n2626), .Z(n2561) );
  XNOR U3716 ( .A(n2559), .B(n2558), .Z(n2560) );
  XNOR U3717 ( .A(n2561), .B(n2560), .Z(n2562) );
  XNOR U3718 ( .A(n2563), .B(n2562), .Z(n2565) );
  XNOR U3719 ( .A(x[50]), .B(n3818), .Z(n2564) );
  XNOR U3720 ( .A(n2565), .B(n2564), .Z(n2595) );
  IV U3721 ( .A(n2595), .Z(n2587) );
  AND U3722 ( .A(n2590), .B(n2587), .Z(n2583) );
  XOR U3723 ( .A(n2594), .B(n2583), .Z(n2571) );
  ANDN U3724 ( .B(n2566), .A(x[49]), .Z(n2570) );
  XNOR U3725 ( .A(n2568), .B(n2567), .Z(n2569) );
  XNOR U3726 ( .A(n2570), .B(n2569), .Z(n2589) );
  ANDN U3727 ( .B(n2571), .A(n2589), .Z(n2578) );
  IV U3728 ( .A(n2590), .Z(n2575) );
  NANDN U3729 ( .A(n2575), .B(n2589), .Z(n2572) );
  NANDN U3730 ( .A(n2578), .B(n2572), .Z(n2602) );
  NANDN U3731 ( .A(n2590), .B(n2587), .Z(n2573) );
  NAND U3732 ( .A(n2573), .B(n2589), .Z(n2577) );
  XNOR U3733 ( .A(n2587), .B(n2594), .Z(n2574) );
  NANDN U3734 ( .A(n2575), .B(n2574), .Z(n2576) );
  AND U3735 ( .A(n2577), .B(n2576), .Z(n2627) );
  OR U3736 ( .A(n2602), .B(n2627), .Z(n2579) );
  ANDN U3737 ( .B(n2579), .A(n2578), .Z(n2606) );
  NANDN U3738 ( .A(n2606), .B(n2580), .Z(n3829) );
  NANDN U3739 ( .A(n2602), .B(n2581), .Z(n2582) );
  XOR U3740 ( .A(n3829), .B(n2582), .Z(n2614) );
  NANDN U3741 ( .A(n2587), .B(n2594), .Z(n2586) );
  XNOR U3742 ( .A(n2583), .B(n2589), .Z(n2584) );
  NANDN U3743 ( .A(n2594), .B(n2584), .Z(n2585) );
  AND U3744 ( .A(n2586), .B(n2585), .Z(n3835) );
  NANDN U3745 ( .A(n2587), .B(n2590), .Z(n2588) );
  NAND U3746 ( .A(n2594), .B(n2588), .Z(n2593) );
  XNOR U3747 ( .A(n2590), .B(n2589), .Z(n2591) );
  NANDN U3748 ( .A(n2595), .B(n2591), .Z(n2592) );
  NAND U3749 ( .A(n2593), .B(n2592), .Z(n3817) );
  IV U3750 ( .A(n3817), .Z(n3808) );
  NANDN U3751 ( .A(n3835), .B(n3808), .Z(n2597) );
  NANDN U3752 ( .A(n2595), .B(n2594), .Z(n2596) );
  NAND U3753 ( .A(n2597), .B(n2596), .Z(n3820) );
  NANDN U3754 ( .A(n3820), .B(n2598), .Z(n3811) );
  NANDN U3755 ( .A(n3835), .B(n3833), .Z(n2599) );
  XNOR U3756 ( .A(n3811), .B(n2599), .Z(n2616) );
  XOR U3757 ( .A(n2614), .B(n2616), .Z(z[50]) );
  NOR U3758 ( .A(n2602), .B(n2600), .Z(n2608) );
  XOR U3759 ( .A(n3808), .B(n2627), .Z(n2609) );
  NANDN U3760 ( .A(n2601), .B(n2609), .Z(n2622) );
  XOR U3761 ( .A(n2602), .B(n3835), .Z(n2629) );
  XNOR U3762 ( .A(n2609), .B(n2629), .Z(n2612) );
  OR U3763 ( .A(n2603), .B(n2612), .Z(n2604) );
  XNOR U3764 ( .A(n2622), .B(n2604), .Z(n3828) );
  NANDN U3765 ( .A(n2606), .B(n2605), .Z(n2617) );
  XNOR U3766 ( .A(n3828), .B(n2617), .Z(n2607) );
  XOR U3767 ( .A(n2608), .B(n2607), .Z(n3825) );
  NANDN U3768 ( .A(n2610), .B(n2609), .Z(n3812) );
  OR U3769 ( .A(n2612), .B(n2611), .Z(n2613) );
  XOR U3770 ( .A(n3812), .B(n2613), .Z(n2623) );
  XOR U3771 ( .A(n2623), .B(n2614), .Z(n3815) );
  XOR U3772 ( .A(n3825), .B(n3815), .Z(n3843) );
  ANDN U3773 ( .B(n2627), .A(n2615), .Z(n2619) );
  XNOR U3774 ( .A(n2617), .B(n2616), .Z(n2618) );
  XNOR U3775 ( .A(n2619), .B(n2618), .Z(n2625) );
  NAND U3776 ( .A(n2620), .B(n2629), .Z(n2621) );
  XNOR U3777 ( .A(n2622), .B(n2621), .Z(n3821) );
  XOR U3778 ( .A(n2623), .B(n3821), .Z(n2624) );
  XOR U3779 ( .A(n2625), .B(n2624), .Z(n3824) );
  XNOR U3780 ( .A(n3843), .B(n3824), .Z(z[49]) );
  ANDN U3781 ( .B(n2627), .A(n2626), .Z(n3831) );
  ANDN U3782 ( .B(n2629), .A(n2628), .Z(n3814) );
  XNOR U3783 ( .A(n3812), .B(z[49]), .Z(n2630) );
  XNOR U3784 ( .A(n3814), .B(n2630), .Z(n2631) );
  XOR U3785 ( .A(n3829), .B(n2631), .Z(n2632) );
  XOR U3786 ( .A(n3831), .B(n2632), .Z(z[55]) );
  IV U3787 ( .A(x[60]), .Z(n2633) );
  IV U3788 ( .A(x[56]), .Z(n2718) );
  XOR U3789 ( .A(n2718), .B(x[62]), .Z(n2634) );
  XOR U3790 ( .A(n2634), .B(x[61]), .Z(n2658) );
  IV U3791 ( .A(n2658), .Z(n3882) );
  XOR U3792 ( .A(n2633), .B(n3882), .Z(n2707) );
  XOR U3793 ( .A(x[57]), .B(x[59]), .Z(n2635) );
  XOR U3794 ( .A(x[63]), .B(n2633), .Z(n2693) );
  XNOR U3795 ( .A(n2635), .B(n2693), .Z(n2672) );
  IV U3796 ( .A(n2672), .Z(n2650) );
  XOR U3797 ( .A(n2635), .B(n2634), .Z(n2636) );
  XOR U3798 ( .A(x[58]), .B(n2636), .Z(n3845) );
  XOR U3799 ( .A(n3845), .B(n2658), .Z(n2690) );
  XOR U3800 ( .A(n2650), .B(n2690), .Z(n2703) );
  IV U3801 ( .A(x[58]), .Z(n2646) );
  XOR U3802 ( .A(x[60]), .B(n2646), .Z(n2695) );
  NOR U3803 ( .A(n2703), .B(n2695), .Z(n2638) );
  XOR U3804 ( .A(x[63]), .B(n3882), .Z(n3853) );
  XOR U3805 ( .A(n3845), .B(n3853), .Z(n2637) );
  XNOR U3806 ( .A(n2638), .B(n2637), .Z(n2639) );
  XNOR U3807 ( .A(n2718), .B(n3845), .Z(n2702) );
  NOR U3808 ( .A(n2693), .B(n2702), .Z(n2648) );
  XNOR U3809 ( .A(n2639), .B(n2648), .Z(n2660) );
  IV U3810 ( .A(x[57]), .Z(n3881) );
  XNOR U3811 ( .A(n3881), .B(x[58]), .Z(n2640) );
  XNOR U3812 ( .A(n3853), .B(n2640), .Z(n2692) );
  ANDN U3813 ( .B(n2692), .A(x[56]), .Z(n2641) );
  XNOR U3814 ( .A(n2693), .B(n2640), .Z(n2697) );
  NANDN U3815 ( .A(n2650), .B(n2697), .Z(n2651) );
  XOR U3816 ( .A(n2641), .B(n2651), .Z(n2643) );
  OR U3817 ( .A(n2692), .B(n2672), .Z(n2642) );
  NAND U3818 ( .A(n2643), .B(n2642), .Z(n2644) );
  XOR U3819 ( .A(n2660), .B(n2644), .Z(n2645) );
  XOR U3820 ( .A(n2707), .B(n2645), .Z(n2686) );
  XNOR U3821 ( .A(n2650), .B(x[56]), .Z(n2673) );
  XNOR U3822 ( .A(n3882), .B(n2673), .Z(n2720) );
  IV U3823 ( .A(x[63]), .Z(n2649) );
  XOR U3824 ( .A(n2649), .B(n2646), .Z(n2712) );
  NANDN U3825 ( .A(n2720), .B(n2712), .Z(n2647) );
  XOR U3826 ( .A(n2648), .B(n2647), .Z(n2655) );
  XOR U3827 ( .A(n3881), .B(n2649), .Z(n3854) );
  NAND U3828 ( .A(n2690), .B(n3854), .Z(n2659) );
  ANDN U3829 ( .B(n2707), .A(n2718), .Z(n2653) );
  XNOR U3830 ( .A(n2651), .B(n2650), .Z(n2652) );
  XNOR U3831 ( .A(n2653), .B(n2652), .Z(n2654) );
  XNOR U3832 ( .A(n2655), .B(n2654), .Z(n2657) );
  XNOR U3833 ( .A(x[58]), .B(n3853), .Z(n2656) );
  XNOR U3834 ( .A(n2657), .B(n2656), .Z(n2687) );
  IV U3835 ( .A(n2687), .Z(n2679) );
  AND U3836 ( .A(n2682), .B(n2679), .Z(n2675) );
  XOR U3837 ( .A(n2686), .B(n2675), .Z(n2663) );
  ANDN U3838 ( .B(n2658), .A(x[57]), .Z(n2662) );
  XNOR U3839 ( .A(n2660), .B(n2659), .Z(n2661) );
  XNOR U3840 ( .A(n2662), .B(n2661), .Z(n2681) );
  ANDN U3841 ( .B(n2663), .A(n2681), .Z(n2670) );
  IV U3842 ( .A(n2682), .Z(n2667) );
  NANDN U3843 ( .A(n2667), .B(n2681), .Z(n2664) );
  NANDN U3844 ( .A(n2670), .B(n2664), .Z(n2694) );
  NANDN U3845 ( .A(n2682), .B(n2679), .Z(n2665) );
  NAND U3846 ( .A(n2665), .B(n2681), .Z(n2669) );
  XNOR U3847 ( .A(n2679), .B(n2686), .Z(n2666) );
  NANDN U3848 ( .A(n2667), .B(n2666), .Z(n2668) );
  AND U3849 ( .A(n2669), .B(n2668), .Z(n2719) );
  OR U3850 ( .A(n2694), .B(n2719), .Z(n2671) );
  ANDN U3851 ( .B(n2671), .A(n2670), .Z(n2698) );
  NANDN U3852 ( .A(n2698), .B(n2672), .Z(n3878) );
  NANDN U3853 ( .A(n2694), .B(n2673), .Z(n2674) );
  XOR U3854 ( .A(n3878), .B(n2674), .Z(n2706) );
  NANDN U3855 ( .A(n2679), .B(n2686), .Z(n2678) );
  XNOR U3856 ( .A(n2675), .B(n2681), .Z(n2676) );
  NANDN U3857 ( .A(n2686), .B(n2676), .Z(n2677) );
  AND U3858 ( .A(n2678), .B(n2677), .Z(n3884) );
  NANDN U3859 ( .A(n2679), .B(n2682), .Z(n2680) );
  NAND U3860 ( .A(n2686), .B(n2680), .Z(n2685) );
  XNOR U3861 ( .A(n2682), .B(n2681), .Z(n2683) );
  NANDN U3862 ( .A(n2687), .B(n2683), .Z(n2684) );
  NAND U3863 ( .A(n2685), .B(n2684), .Z(n3852) );
  IV U3864 ( .A(n3852), .Z(n3844) );
  NANDN U3865 ( .A(n3884), .B(n3844), .Z(n2689) );
  NANDN U3866 ( .A(n2687), .B(n2686), .Z(n2688) );
  NAND U3867 ( .A(n2689), .B(n2688), .Z(n3855) );
  NANDN U3868 ( .A(n3855), .B(n2690), .Z(n3847) );
  NANDN U3869 ( .A(n3884), .B(n3882), .Z(n2691) );
  XNOR U3870 ( .A(n3847), .B(n2691), .Z(n2708) );
  XOR U3871 ( .A(n2706), .B(n2708), .Z(z[58]) );
  NOR U3872 ( .A(n2694), .B(n2692), .Z(n2700) );
  XOR U3873 ( .A(n3844), .B(n2719), .Z(n2701) );
  NANDN U3874 ( .A(n2693), .B(n2701), .Z(n2714) );
  XOR U3875 ( .A(n2694), .B(n3884), .Z(n2721) );
  XNOR U3876 ( .A(n2701), .B(n2721), .Z(n2704) );
  OR U3877 ( .A(n2695), .B(n2704), .Z(n2696) );
  XNOR U3878 ( .A(n2714), .B(n2696), .Z(n3877) );
  NANDN U3879 ( .A(n2698), .B(n2697), .Z(n2709) );
  XNOR U3880 ( .A(n3877), .B(n2709), .Z(n2699) );
  XOR U3881 ( .A(n2700), .B(n2699), .Z(n3860) );
  NANDN U3882 ( .A(n2702), .B(n2701), .Z(n3848) );
  OR U3883 ( .A(n2704), .B(n2703), .Z(n2705) );
  XOR U3884 ( .A(n3848), .B(n2705), .Z(n2715) );
  XOR U3885 ( .A(n2715), .B(n2706), .Z(n3851) );
  XOR U3886 ( .A(n3860), .B(n3851), .Z(n3892) );
  ANDN U3887 ( .B(n2719), .A(n2707), .Z(n2711) );
  XNOR U3888 ( .A(n2709), .B(n2708), .Z(n2710) );
  XNOR U3889 ( .A(n2711), .B(n2710), .Z(n2717) );
  NAND U3890 ( .A(n2712), .B(n2721), .Z(n2713) );
  XNOR U3891 ( .A(n2714), .B(n2713), .Z(n3856) );
  XOR U3892 ( .A(n2715), .B(n3856), .Z(n2716) );
  XOR U3893 ( .A(n2717), .B(n2716), .Z(n3859) );
  XNOR U3894 ( .A(n3892), .B(n3859), .Z(z[57]) );
  ANDN U3895 ( .B(n2719), .A(n2718), .Z(n3880) );
  ANDN U3896 ( .B(n2721), .A(n2720), .Z(n3850) );
  XNOR U3897 ( .A(n3848), .B(z[57]), .Z(n2722) );
  XNOR U3898 ( .A(n3850), .B(n2722), .Z(n2723) );
  XOR U3899 ( .A(n3878), .B(n2723), .Z(n2724) );
  XOR U3900 ( .A(n3880), .B(n2724), .Z(z[63]) );
  IV U3901 ( .A(x[68]), .Z(n2725) );
  IV U3902 ( .A(x[64]), .Z(n2810) );
  XOR U3903 ( .A(n2810), .B(x[70]), .Z(n2726) );
  XOR U3904 ( .A(n2726), .B(x[69]), .Z(n2750) );
  IV U3905 ( .A(n2750), .Z(n3917) );
  XOR U3906 ( .A(n2725), .B(n3917), .Z(n2799) );
  XOR U3907 ( .A(x[65]), .B(x[67]), .Z(n2727) );
  XOR U3908 ( .A(x[71]), .B(n2725), .Z(n2785) );
  XNOR U3909 ( .A(n2727), .B(n2785), .Z(n2764) );
  IV U3910 ( .A(n2764), .Z(n2742) );
  XOR U3911 ( .A(n2727), .B(n2726), .Z(n2728) );
  XOR U3912 ( .A(x[66]), .B(n2728), .Z(n3894) );
  XOR U3913 ( .A(n3894), .B(n2750), .Z(n2782) );
  XOR U3914 ( .A(n2742), .B(n2782), .Z(n2795) );
  IV U3915 ( .A(x[66]), .Z(n2738) );
  XOR U3916 ( .A(x[68]), .B(n2738), .Z(n2787) );
  NOR U3917 ( .A(n2795), .B(n2787), .Z(n2730) );
  XOR U3918 ( .A(x[71]), .B(n3917), .Z(n3902) );
  XOR U3919 ( .A(n3894), .B(n3902), .Z(n2729) );
  XNOR U3920 ( .A(n2730), .B(n2729), .Z(n2731) );
  XNOR U3921 ( .A(n2810), .B(n3894), .Z(n2794) );
  NOR U3922 ( .A(n2785), .B(n2794), .Z(n2740) );
  XNOR U3923 ( .A(n2731), .B(n2740), .Z(n2752) );
  IV U3924 ( .A(x[65]), .Z(n3916) );
  XNOR U3925 ( .A(n3916), .B(x[66]), .Z(n2732) );
  XNOR U3926 ( .A(n3902), .B(n2732), .Z(n2784) );
  ANDN U3927 ( .B(n2784), .A(x[64]), .Z(n2733) );
  XNOR U3928 ( .A(n2785), .B(n2732), .Z(n2789) );
  NANDN U3929 ( .A(n2742), .B(n2789), .Z(n2743) );
  XOR U3930 ( .A(n2733), .B(n2743), .Z(n2735) );
  OR U3931 ( .A(n2784), .B(n2764), .Z(n2734) );
  NAND U3932 ( .A(n2735), .B(n2734), .Z(n2736) );
  XOR U3933 ( .A(n2752), .B(n2736), .Z(n2737) );
  XOR U3934 ( .A(n2799), .B(n2737), .Z(n2778) );
  XNOR U3935 ( .A(n2742), .B(x[64]), .Z(n2765) );
  XNOR U3936 ( .A(n3917), .B(n2765), .Z(n2812) );
  IV U3937 ( .A(x[71]), .Z(n2741) );
  XOR U3938 ( .A(n2741), .B(n2738), .Z(n2804) );
  NANDN U3939 ( .A(n2812), .B(n2804), .Z(n2739) );
  XOR U3940 ( .A(n2740), .B(n2739), .Z(n2747) );
  XOR U3941 ( .A(n3916), .B(n2741), .Z(n3903) );
  NAND U3942 ( .A(n2782), .B(n3903), .Z(n2751) );
  ANDN U3943 ( .B(n2799), .A(n2810), .Z(n2745) );
  XNOR U3944 ( .A(n2743), .B(n2742), .Z(n2744) );
  XNOR U3945 ( .A(n2745), .B(n2744), .Z(n2746) );
  XNOR U3946 ( .A(n2747), .B(n2746), .Z(n2749) );
  XNOR U3947 ( .A(x[66]), .B(n3902), .Z(n2748) );
  XNOR U3948 ( .A(n2749), .B(n2748), .Z(n2779) );
  IV U3949 ( .A(n2779), .Z(n2771) );
  AND U3950 ( .A(n2774), .B(n2771), .Z(n2767) );
  XOR U3951 ( .A(n2778), .B(n2767), .Z(n2755) );
  ANDN U3952 ( .B(n2750), .A(x[65]), .Z(n2754) );
  XNOR U3953 ( .A(n2752), .B(n2751), .Z(n2753) );
  XNOR U3954 ( .A(n2754), .B(n2753), .Z(n2773) );
  ANDN U3955 ( .B(n2755), .A(n2773), .Z(n2762) );
  IV U3956 ( .A(n2774), .Z(n2759) );
  NANDN U3957 ( .A(n2759), .B(n2773), .Z(n2756) );
  NANDN U3958 ( .A(n2762), .B(n2756), .Z(n2786) );
  NANDN U3959 ( .A(n2774), .B(n2771), .Z(n2757) );
  NAND U3960 ( .A(n2757), .B(n2773), .Z(n2761) );
  XNOR U3961 ( .A(n2771), .B(n2778), .Z(n2758) );
  NANDN U3962 ( .A(n2759), .B(n2758), .Z(n2760) );
  AND U3963 ( .A(n2761), .B(n2760), .Z(n2811) );
  OR U3964 ( .A(n2786), .B(n2811), .Z(n2763) );
  ANDN U3965 ( .B(n2763), .A(n2762), .Z(n2790) );
  NANDN U3966 ( .A(n2790), .B(n2764), .Z(n3913) );
  NANDN U3967 ( .A(n2786), .B(n2765), .Z(n2766) );
  XOR U3968 ( .A(n3913), .B(n2766), .Z(n2798) );
  NANDN U3969 ( .A(n2771), .B(n2778), .Z(n2770) );
  XNOR U3970 ( .A(n2767), .B(n2773), .Z(n2768) );
  NANDN U3971 ( .A(n2778), .B(n2768), .Z(n2769) );
  AND U3972 ( .A(n2770), .B(n2769), .Z(n3919) );
  NANDN U3973 ( .A(n2771), .B(n2774), .Z(n2772) );
  NAND U3974 ( .A(n2778), .B(n2772), .Z(n2777) );
  XNOR U3975 ( .A(n2774), .B(n2773), .Z(n2775) );
  NANDN U3976 ( .A(n2779), .B(n2775), .Z(n2776) );
  NAND U3977 ( .A(n2777), .B(n2776), .Z(n3901) );
  IV U3978 ( .A(n3901), .Z(n3893) );
  NANDN U3979 ( .A(n3919), .B(n3893), .Z(n2781) );
  NANDN U3980 ( .A(n2779), .B(n2778), .Z(n2780) );
  NAND U3981 ( .A(n2781), .B(n2780), .Z(n3904) );
  NANDN U3982 ( .A(n3904), .B(n2782), .Z(n3896) );
  NANDN U3983 ( .A(n3919), .B(n3917), .Z(n2783) );
  XNOR U3984 ( .A(n3896), .B(n2783), .Z(n2800) );
  XOR U3985 ( .A(n2798), .B(n2800), .Z(z[66]) );
  NOR U3986 ( .A(n2786), .B(n2784), .Z(n2792) );
  XOR U3987 ( .A(n3893), .B(n2811), .Z(n2793) );
  NANDN U3988 ( .A(n2785), .B(n2793), .Z(n2806) );
  XOR U3989 ( .A(n2786), .B(n3919), .Z(n2813) );
  XNOR U3990 ( .A(n2793), .B(n2813), .Z(n2796) );
  OR U3991 ( .A(n2787), .B(n2796), .Z(n2788) );
  XNOR U3992 ( .A(n2806), .B(n2788), .Z(n3912) );
  NANDN U3993 ( .A(n2790), .B(n2789), .Z(n2801) );
  XNOR U3994 ( .A(n3912), .B(n2801), .Z(n2791) );
  XOR U3995 ( .A(n2792), .B(n2791), .Z(n3909) );
  NANDN U3996 ( .A(n2794), .B(n2793), .Z(n3897) );
  OR U3997 ( .A(n2796), .B(n2795), .Z(n2797) );
  XOR U3998 ( .A(n3897), .B(n2797), .Z(n2807) );
  XOR U3999 ( .A(n2807), .B(n2798), .Z(n3900) );
  XOR U4000 ( .A(n3909), .B(n3900), .Z(n3929) );
  ANDN U4001 ( .B(n2811), .A(n2799), .Z(n2803) );
  XNOR U4002 ( .A(n2801), .B(n2800), .Z(n2802) );
  XNOR U4003 ( .A(n2803), .B(n2802), .Z(n2809) );
  NAND U4004 ( .A(n2804), .B(n2813), .Z(n2805) );
  XNOR U4005 ( .A(n2806), .B(n2805), .Z(n3905) );
  XOR U4006 ( .A(n2807), .B(n3905), .Z(n2808) );
  XOR U4007 ( .A(n2809), .B(n2808), .Z(n3908) );
  XNOR U4008 ( .A(n3929), .B(n3908), .Z(z[65]) );
  ANDN U4009 ( .B(n2811), .A(n2810), .Z(n3915) );
  ANDN U4010 ( .B(n2813), .A(n2812), .Z(n3899) );
  XNOR U4011 ( .A(n3897), .B(z[65]), .Z(n2814) );
  XNOR U4012 ( .A(n3899), .B(n2814), .Z(n2815) );
  XOR U4013 ( .A(n3913), .B(n2815), .Z(n2816) );
  XOR U4014 ( .A(n3915), .B(n2816), .Z(z[71]) );
  IV U4015 ( .A(x[76]), .Z(n2817) );
  IV U4016 ( .A(x[72]), .Z(n2902) );
  XOR U4017 ( .A(n2902), .B(x[78]), .Z(n2818) );
  XOR U4018 ( .A(n2818), .B(x[77]), .Z(n2842) );
  IV U4019 ( .A(n2842), .Z(n3954) );
  XOR U4020 ( .A(n2817), .B(n3954), .Z(n2891) );
  XOR U4021 ( .A(x[73]), .B(x[75]), .Z(n2819) );
  XOR U4022 ( .A(x[79]), .B(n2817), .Z(n2877) );
  XNOR U4023 ( .A(n2819), .B(n2877), .Z(n2856) );
  IV U4024 ( .A(n2856), .Z(n2834) );
  XOR U4025 ( .A(n2819), .B(n2818), .Z(n2820) );
  XOR U4026 ( .A(x[74]), .B(n2820), .Z(n3931) );
  XOR U4027 ( .A(n3931), .B(n2842), .Z(n2874) );
  XOR U4028 ( .A(n2834), .B(n2874), .Z(n2887) );
  IV U4029 ( .A(x[74]), .Z(n2830) );
  XOR U4030 ( .A(x[76]), .B(n2830), .Z(n2879) );
  NOR U4031 ( .A(n2887), .B(n2879), .Z(n2822) );
  XOR U4032 ( .A(x[79]), .B(n3954), .Z(n3939) );
  XOR U4033 ( .A(n3931), .B(n3939), .Z(n2821) );
  XNOR U4034 ( .A(n2822), .B(n2821), .Z(n2823) );
  XNOR U4035 ( .A(n2902), .B(n3931), .Z(n2886) );
  NOR U4036 ( .A(n2877), .B(n2886), .Z(n2832) );
  XNOR U4037 ( .A(n2823), .B(n2832), .Z(n2844) );
  IV U4038 ( .A(x[73]), .Z(n3953) );
  XNOR U4039 ( .A(n3953), .B(x[74]), .Z(n2824) );
  XNOR U4040 ( .A(n3939), .B(n2824), .Z(n2876) );
  ANDN U4041 ( .B(n2876), .A(x[72]), .Z(n2825) );
  XNOR U4042 ( .A(n2877), .B(n2824), .Z(n2881) );
  NANDN U4043 ( .A(n2834), .B(n2881), .Z(n2835) );
  XOR U4044 ( .A(n2825), .B(n2835), .Z(n2827) );
  OR U4045 ( .A(n2876), .B(n2856), .Z(n2826) );
  NAND U4046 ( .A(n2827), .B(n2826), .Z(n2828) );
  XOR U4047 ( .A(n2844), .B(n2828), .Z(n2829) );
  XOR U4048 ( .A(n2891), .B(n2829), .Z(n2870) );
  XNOR U4049 ( .A(n2834), .B(x[72]), .Z(n2857) );
  XNOR U4050 ( .A(n3954), .B(n2857), .Z(n2904) );
  IV U4051 ( .A(x[79]), .Z(n2833) );
  XOR U4052 ( .A(n2833), .B(n2830), .Z(n2896) );
  NANDN U4053 ( .A(n2904), .B(n2896), .Z(n2831) );
  XOR U4054 ( .A(n2832), .B(n2831), .Z(n2839) );
  XOR U4055 ( .A(n3953), .B(n2833), .Z(n3940) );
  NAND U4056 ( .A(n2874), .B(n3940), .Z(n2843) );
  ANDN U4057 ( .B(n2891), .A(n2902), .Z(n2837) );
  XNOR U4058 ( .A(n2835), .B(n2834), .Z(n2836) );
  XNOR U4059 ( .A(n2837), .B(n2836), .Z(n2838) );
  XNOR U4060 ( .A(n2839), .B(n2838), .Z(n2841) );
  XNOR U4061 ( .A(x[74]), .B(n3939), .Z(n2840) );
  XNOR U4062 ( .A(n2841), .B(n2840), .Z(n2871) );
  IV U4063 ( .A(n2871), .Z(n2863) );
  AND U4064 ( .A(n2866), .B(n2863), .Z(n2859) );
  XOR U4065 ( .A(n2870), .B(n2859), .Z(n2847) );
  ANDN U4066 ( .B(n2842), .A(x[73]), .Z(n2846) );
  XNOR U4067 ( .A(n2844), .B(n2843), .Z(n2845) );
  XNOR U4068 ( .A(n2846), .B(n2845), .Z(n2865) );
  ANDN U4069 ( .B(n2847), .A(n2865), .Z(n2854) );
  IV U4070 ( .A(n2866), .Z(n2851) );
  NANDN U4071 ( .A(n2851), .B(n2865), .Z(n2848) );
  NANDN U4072 ( .A(n2854), .B(n2848), .Z(n2878) );
  NANDN U4073 ( .A(n2866), .B(n2863), .Z(n2849) );
  NAND U4074 ( .A(n2849), .B(n2865), .Z(n2853) );
  XNOR U4075 ( .A(n2863), .B(n2870), .Z(n2850) );
  NANDN U4076 ( .A(n2851), .B(n2850), .Z(n2852) );
  AND U4077 ( .A(n2853), .B(n2852), .Z(n2903) );
  OR U4078 ( .A(n2878), .B(n2903), .Z(n2855) );
  ANDN U4079 ( .B(n2855), .A(n2854), .Z(n2882) );
  NANDN U4080 ( .A(n2882), .B(n2856), .Z(n3950) );
  NANDN U4081 ( .A(n2878), .B(n2857), .Z(n2858) );
  XOR U4082 ( .A(n3950), .B(n2858), .Z(n2890) );
  NANDN U4083 ( .A(n2863), .B(n2870), .Z(n2862) );
  XNOR U4084 ( .A(n2859), .B(n2865), .Z(n2860) );
  NANDN U4085 ( .A(n2870), .B(n2860), .Z(n2861) );
  AND U4086 ( .A(n2862), .B(n2861), .Z(n3956) );
  NANDN U4087 ( .A(n2863), .B(n2866), .Z(n2864) );
  NAND U4088 ( .A(n2870), .B(n2864), .Z(n2869) );
  XNOR U4089 ( .A(n2866), .B(n2865), .Z(n2867) );
  NANDN U4090 ( .A(n2871), .B(n2867), .Z(n2868) );
  NAND U4091 ( .A(n2869), .B(n2868), .Z(n3938) );
  IV U4092 ( .A(n3938), .Z(n3930) );
  NANDN U4093 ( .A(n3956), .B(n3930), .Z(n2873) );
  NANDN U4094 ( .A(n2871), .B(n2870), .Z(n2872) );
  NAND U4095 ( .A(n2873), .B(n2872), .Z(n3941) );
  NANDN U4096 ( .A(n3941), .B(n2874), .Z(n3933) );
  NANDN U4097 ( .A(n3956), .B(n3954), .Z(n2875) );
  XNOR U4098 ( .A(n3933), .B(n2875), .Z(n2892) );
  XOR U4099 ( .A(n2890), .B(n2892), .Z(z[74]) );
  NOR U4100 ( .A(n2878), .B(n2876), .Z(n2884) );
  XOR U4101 ( .A(n3930), .B(n2903), .Z(n2885) );
  NANDN U4102 ( .A(n2877), .B(n2885), .Z(n2898) );
  XOR U4103 ( .A(n2878), .B(n3956), .Z(n2905) );
  XNOR U4104 ( .A(n2885), .B(n2905), .Z(n2888) );
  OR U4105 ( .A(n2879), .B(n2888), .Z(n2880) );
  XNOR U4106 ( .A(n2898), .B(n2880), .Z(n3949) );
  NANDN U4107 ( .A(n2882), .B(n2881), .Z(n2893) );
  XNOR U4108 ( .A(n3949), .B(n2893), .Z(n2883) );
  XOR U4109 ( .A(n2884), .B(n2883), .Z(n3946) );
  NANDN U4110 ( .A(n2886), .B(n2885), .Z(n3934) );
  OR U4111 ( .A(n2888), .B(n2887), .Z(n2889) );
  XOR U4112 ( .A(n3934), .B(n2889), .Z(n2899) );
  XOR U4113 ( .A(n2899), .B(n2890), .Z(n3937) );
  XOR U4114 ( .A(n3946), .B(n3937), .Z(n3964) );
  ANDN U4115 ( .B(n2903), .A(n2891), .Z(n2895) );
  XNOR U4116 ( .A(n2893), .B(n2892), .Z(n2894) );
  XNOR U4117 ( .A(n2895), .B(n2894), .Z(n2901) );
  NAND U4118 ( .A(n2896), .B(n2905), .Z(n2897) );
  XNOR U4119 ( .A(n2898), .B(n2897), .Z(n3942) );
  XOR U4120 ( .A(n2899), .B(n3942), .Z(n2900) );
  XOR U4121 ( .A(n2901), .B(n2900), .Z(n3945) );
  XNOR U4122 ( .A(n3964), .B(n3945), .Z(z[73]) );
  ANDN U4123 ( .B(n2903), .A(n2902), .Z(n3952) );
  ANDN U4124 ( .B(n2905), .A(n2904), .Z(n3936) );
  XNOR U4125 ( .A(n3934), .B(z[73]), .Z(n2906) );
  XNOR U4126 ( .A(n3936), .B(n2906), .Z(n2907) );
  XOR U4127 ( .A(n3950), .B(n2907), .Z(n2908) );
  XOR U4128 ( .A(n3952), .B(n2908), .Z(z[79]) );
  XOR U4129 ( .A(x[80]), .B(x[86]), .Z(n2909) );
  XOR U4130 ( .A(n2909), .B(x[85]), .Z(n3989) );
  IV U4131 ( .A(n3989), .Z(n2912) );
  XOR U4132 ( .A(x[84]), .B(n2912), .Z(n2978) );
  XNOR U4133 ( .A(x[87]), .B(n2912), .Z(n3974) );
  IV U4134 ( .A(x[81]), .Z(n3988) );
  IV U4135 ( .A(x[82]), .Z(n2916) );
  XOR U4136 ( .A(n3988), .B(n2916), .Z(n2920) );
  XOR U4137 ( .A(n3974), .B(n2920), .Z(n2963) );
  XOR U4138 ( .A(n3988), .B(x[83]), .Z(n2910) );
  IV U4139 ( .A(x[87]), .Z(n2925) );
  XOR U4140 ( .A(x[84]), .B(n2925), .Z(n2964) );
  XOR U4141 ( .A(n2910), .B(n2964), .Z(n2942) );
  IV U4142 ( .A(x[80]), .Z(n2989) );
  XOR U4143 ( .A(n2910), .B(n2909), .Z(n2911) );
  XOR U4144 ( .A(x[82]), .B(n2911), .Z(n3966) );
  XOR U4145 ( .A(n3966), .B(n2912), .Z(n2961) );
  XNOR U4146 ( .A(n2942), .B(n2961), .Z(n2974) );
  XOR U4147 ( .A(x[84]), .B(n2916), .Z(n2966) );
  NOR U4148 ( .A(n2974), .B(n2966), .Z(n2914) );
  XOR U4149 ( .A(n3966), .B(n3974), .Z(n2913) );
  XNOR U4150 ( .A(n2914), .B(n2913), .Z(n2915) );
  XNOR U4151 ( .A(n2989), .B(n3966), .Z(n2973) );
  NOR U4152 ( .A(n2964), .B(n2973), .Z(n2918) );
  XNOR U4153 ( .A(n2915), .B(n2918), .Z(n2932) );
  XOR U4154 ( .A(n2964), .B(n2920), .Z(n2968) );
  NANDN U4155 ( .A(n2968), .B(n2942), .Z(n2919) );
  IV U4156 ( .A(n2957), .Z(n2950) );
  XNOR U4157 ( .A(n2942), .B(n2989), .Z(n2943) );
  XNOR U4158 ( .A(n3989), .B(n2943), .Z(n2991) );
  XOR U4159 ( .A(x[87]), .B(n2916), .Z(n2983) );
  OR U4160 ( .A(n2991), .B(n2983), .Z(n2917) );
  XOR U4161 ( .A(n2918), .B(n2917), .Z(n2928) );
  XOR U4162 ( .A(n2919), .B(n2928), .Z(n2922) );
  XNOR U4163 ( .A(x[83]), .B(n2920), .Z(n2921) );
  XNOR U4164 ( .A(n2922), .B(n2921), .Z(n2924) );
  NANDN U4165 ( .A(x[80]), .B(n2978), .Z(n2923) );
  XNOR U4166 ( .A(n2924), .B(n2923), .Z(n2951) );
  ANDN U4167 ( .B(n3966), .A(n3974), .Z(n2926) );
  XOR U4168 ( .A(n3988), .B(n2925), .Z(n3975) );
  NAND U4169 ( .A(n2961), .B(n3975), .Z(n2930) );
  XOR U4170 ( .A(n2926), .B(n2930), .Z(n2927) );
  XNOR U4171 ( .A(n2928), .B(n2927), .Z(n2937) );
  IV U4172 ( .A(n2937), .Z(n2953) );
  AND U4173 ( .A(n2951), .B(n2953), .Z(n2945) );
  XNOR U4174 ( .A(n2950), .B(n2945), .Z(n2933) );
  ANDN U4175 ( .B(n3988), .A(n3989), .Z(n2929) );
  XOR U4176 ( .A(n2930), .B(n2929), .Z(n2931) );
  XOR U4177 ( .A(n2932), .B(n2931), .Z(n2952) );
  ANDN U4178 ( .B(n2933), .A(n2952), .Z(n2940) );
  NANDN U4179 ( .A(n2937), .B(n2952), .Z(n2934) );
  NANDN U4180 ( .A(n2940), .B(n2934), .Z(n2965) );
  NANDN U4181 ( .A(n2953), .B(n2951), .Z(n2935) );
  NAND U4182 ( .A(n2935), .B(n2952), .Z(n2939) );
  XNOR U4183 ( .A(n2951), .B(n2957), .Z(n2936) );
  NANDN U4184 ( .A(n2937), .B(n2936), .Z(n2938) );
  AND U4185 ( .A(n2939), .B(n2938), .Z(n2990) );
  OR U4186 ( .A(n2965), .B(n2990), .Z(n2941) );
  ANDN U4187 ( .B(n2941), .A(n2940), .Z(n2969) );
  NANDN U4188 ( .A(n2969), .B(n2942), .Z(n3985) );
  NANDN U4189 ( .A(n2965), .B(n2943), .Z(n2944) );
  XOR U4190 ( .A(n3985), .B(n2944), .Z(n2977) );
  NANDN U4191 ( .A(n2951), .B(n2957), .Z(n2948) );
  XNOR U4192 ( .A(n2945), .B(n2952), .Z(n2946) );
  NANDN U4193 ( .A(n2957), .B(n2946), .Z(n2947) );
  AND U4194 ( .A(n2948), .B(n2947), .Z(n3991) );
  NANDN U4195 ( .A(n2951), .B(n2953), .Z(n2949) );
  NANDN U4196 ( .A(n2950), .B(n2949), .Z(n2956) );
  IV U4197 ( .A(n2951), .Z(n2958) );
  XNOR U4198 ( .A(n2953), .B(n2952), .Z(n2954) );
  NANDN U4199 ( .A(n2958), .B(n2954), .Z(n2955) );
  NAND U4200 ( .A(n2956), .B(n2955), .Z(n3973) );
  IV U4201 ( .A(n3973), .Z(n3965) );
  NANDN U4202 ( .A(n3991), .B(n3965), .Z(n2960) );
  NANDN U4203 ( .A(n2958), .B(n2957), .Z(n2959) );
  NAND U4204 ( .A(n2960), .B(n2959), .Z(n3976) );
  NANDN U4205 ( .A(n3976), .B(n2961), .Z(n3968) );
  NANDN U4206 ( .A(n3991), .B(n3989), .Z(n2962) );
  XNOR U4207 ( .A(n3968), .B(n2962), .Z(n2979) );
  XOR U4208 ( .A(n2977), .B(n2979), .Z(z[82]) );
  ANDN U4209 ( .B(n2963), .A(n2965), .Z(n2971) );
  XOR U4210 ( .A(n3965), .B(n2990), .Z(n2972) );
  NANDN U4211 ( .A(n2964), .B(n2972), .Z(n2985) );
  XOR U4212 ( .A(n2965), .B(n3991), .Z(n2992) );
  XNOR U4213 ( .A(n2972), .B(n2992), .Z(n2975) );
  OR U4214 ( .A(n2966), .B(n2975), .Z(n2967) );
  XNOR U4215 ( .A(n2985), .B(n2967), .Z(n3984) );
  OR U4216 ( .A(n2969), .B(n2968), .Z(n2980) );
  XNOR U4217 ( .A(n3984), .B(n2980), .Z(n2970) );
  XOR U4218 ( .A(n2971), .B(n2970), .Z(n3981) );
  NANDN U4219 ( .A(n2973), .B(n2972), .Z(n3969) );
  OR U4220 ( .A(n2975), .B(n2974), .Z(n2976) );
  XOR U4221 ( .A(n3969), .B(n2976), .Z(n2986) );
  XOR U4222 ( .A(n2986), .B(n2977), .Z(n3972) );
  XOR U4223 ( .A(n3981), .B(n3972), .Z(n3999) );
  ANDN U4224 ( .B(n2990), .A(n2978), .Z(n2982) );
  XNOR U4225 ( .A(n2980), .B(n2979), .Z(n2981) );
  XNOR U4226 ( .A(n2982), .B(n2981), .Z(n2988) );
  NANDN U4227 ( .A(n2983), .B(n2992), .Z(n2984) );
  XNOR U4228 ( .A(n2985), .B(n2984), .Z(n3977) );
  XOR U4229 ( .A(n2986), .B(n3977), .Z(n2987) );
  XOR U4230 ( .A(n2988), .B(n2987), .Z(n3980) );
  XNOR U4231 ( .A(n3999), .B(n3980), .Z(z[81]) );
  ANDN U4232 ( .B(n2990), .A(n2989), .Z(n3987) );
  ANDN U4233 ( .B(n2992), .A(n2991), .Z(n3971) );
  XNOR U4234 ( .A(n3969), .B(z[81]), .Z(n2993) );
  XNOR U4235 ( .A(n3971), .B(n2993), .Z(n2994) );
  XOR U4236 ( .A(n3985), .B(n2994), .Z(n2995) );
  XOR U4237 ( .A(n3987), .B(n2995), .Z(z[87]) );
  XOR U4238 ( .A(x[88]), .B(x[94]), .Z(n2996) );
  XOR U4239 ( .A(n2996), .B(x[93]), .Z(n4026) );
  IV U4240 ( .A(n4026), .Z(n2999) );
  XOR U4241 ( .A(x[92]), .B(n2999), .Z(n3065) );
  XNOR U4242 ( .A(x[95]), .B(n2999), .Z(n4011) );
  IV U4243 ( .A(x[89]), .Z(n4025) );
  IV U4244 ( .A(x[90]), .Z(n3003) );
  XOR U4245 ( .A(n4025), .B(n3003), .Z(n3007) );
  XOR U4246 ( .A(n4011), .B(n3007), .Z(n3050) );
  XOR U4247 ( .A(n4025), .B(x[91]), .Z(n2997) );
  IV U4248 ( .A(x[95]), .Z(n3012) );
  XOR U4249 ( .A(x[92]), .B(n3012), .Z(n3051) );
  XOR U4250 ( .A(n2997), .B(n3051), .Z(n3029) );
  IV U4251 ( .A(x[88]), .Z(n3076) );
  XOR U4252 ( .A(n2997), .B(n2996), .Z(n2998) );
  XOR U4253 ( .A(x[90]), .B(n2998), .Z(n4001) );
  XOR U4254 ( .A(n4001), .B(n2999), .Z(n3048) );
  XNOR U4255 ( .A(n3029), .B(n3048), .Z(n3061) );
  XOR U4256 ( .A(x[92]), .B(n3003), .Z(n3053) );
  NOR U4257 ( .A(n3061), .B(n3053), .Z(n3001) );
  XOR U4258 ( .A(n4001), .B(n4011), .Z(n3000) );
  XNOR U4259 ( .A(n3001), .B(n3000), .Z(n3002) );
  XNOR U4260 ( .A(n3076), .B(n4001), .Z(n3060) );
  NOR U4261 ( .A(n3051), .B(n3060), .Z(n3005) );
  XNOR U4262 ( .A(n3002), .B(n3005), .Z(n3019) );
  XOR U4263 ( .A(n3051), .B(n3007), .Z(n3055) );
  NANDN U4264 ( .A(n3055), .B(n3029), .Z(n3006) );
  IV U4265 ( .A(n3044), .Z(n3037) );
  XNOR U4266 ( .A(n3029), .B(n3076), .Z(n3030) );
  XNOR U4267 ( .A(n4026), .B(n3030), .Z(n3078) );
  XOR U4268 ( .A(x[95]), .B(n3003), .Z(n3070) );
  OR U4269 ( .A(n3078), .B(n3070), .Z(n3004) );
  XOR U4270 ( .A(n3005), .B(n3004), .Z(n3015) );
  XOR U4271 ( .A(n3006), .B(n3015), .Z(n3009) );
  XNOR U4272 ( .A(x[91]), .B(n3007), .Z(n3008) );
  XNOR U4273 ( .A(n3009), .B(n3008), .Z(n3011) );
  NANDN U4274 ( .A(x[88]), .B(n3065), .Z(n3010) );
  XNOR U4275 ( .A(n3011), .B(n3010), .Z(n3038) );
  ANDN U4276 ( .B(n4001), .A(n4011), .Z(n3013) );
  XOR U4277 ( .A(n4025), .B(n3012), .Z(n4012) );
  NAND U4278 ( .A(n3048), .B(n4012), .Z(n3017) );
  XOR U4279 ( .A(n3013), .B(n3017), .Z(n3014) );
  XNOR U4280 ( .A(n3015), .B(n3014), .Z(n3024) );
  IV U4281 ( .A(n3024), .Z(n3040) );
  AND U4282 ( .A(n3038), .B(n3040), .Z(n3032) );
  XNOR U4283 ( .A(n3037), .B(n3032), .Z(n3020) );
  ANDN U4284 ( .B(n4025), .A(n4026), .Z(n3016) );
  XOR U4285 ( .A(n3017), .B(n3016), .Z(n3018) );
  XOR U4286 ( .A(n3019), .B(n3018), .Z(n3039) );
  ANDN U4287 ( .B(n3020), .A(n3039), .Z(n3027) );
  NANDN U4288 ( .A(n3024), .B(n3039), .Z(n3021) );
  NANDN U4289 ( .A(n3027), .B(n3021), .Z(n3052) );
  NANDN U4290 ( .A(n3040), .B(n3038), .Z(n3022) );
  NAND U4291 ( .A(n3022), .B(n3039), .Z(n3026) );
  XNOR U4292 ( .A(n3038), .B(n3044), .Z(n3023) );
  NANDN U4293 ( .A(n3024), .B(n3023), .Z(n3025) );
  AND U4294 ( .A(n3026), .B(n3025), .Z(n3077) );
  OR U4295 ( .A(n3052), .B(n3077), .Z(n3028) );
  ANDN U4296 ( .B(n3028), .A(n3027), .Z(n3056) );
  NANDN U4297 ( .A(n3056), .B(n3029), .Z(n4022) );
  NANDN U4298 ( .A(n3052), .B(n3030), .Z(n3031) );
  XOR U4299 ( .A(n4022), .B(n3031), .Z(n3064) );
  NANDN U4300 ( .A(n3038), .B(n3044), .Z(n3035) );
  XNOR U4301 ( .A(n3032), .B(n3039), .Z(n3033) );
  NANDN U4302 ( .A(n3044), .B(n3033), .Z(n3034) );
  AND U4303 ( .A(n3035), .B(n3034), .Z(n4028) );
  NANDN U4304 ( .A(n3038), .B(n3040), .Z(n3036) );
  NANDN U4305 ( .A(n3037), .B(n3036), .Z(n3043) );
  IV U4306 ( .A(n3038), .Z(n3045) );
  XNOR U4307 ( .A(n3040), .B(n3039), .Z(n3041) );
  NANDN U4308 ( .A(n3045), .B(n3041), .Z(n3042) );
  NAND U4309 ( .A(n3043), .B(n3042), .Z(n4010) );
  IV U4310 ( .A(n4010), .Z(n4000) );
  NANDN U4311 ( .A(n4028), .B(n4000), .Z(n3047) );
  NANDN U4312 ( .A(n3045), .B(n3044), .Z(n3046) );
  NAND U4313 ( .A(n3047), .B(n3046), .Z(n4013) );
  NANDN U4314 ( .A(n4013), .B(n3048), .Z(n4003) );
  NANDN U4315 ( .A(n4028), .B(n4026), .Z(n3049) );
  XNOR U4316 ( .A(n4003), .B(n3049), .Z(n3066) );
  XOR U4317 ( .A(n3064), .B(n3066), .Z(z[90]) );
  ANDN U4318 ( .B(n3050), .A(n3052), .Z(n3058) );
  XOR U4319 ( .A(n4000), .B(n3077), .Z(n3059) );
  NANDN U4320 ( .A(n3051), .B(n3059), .Z(n3072) );
  XOR U4321 ( .A(n3052), .B(n4028), .Z(n3079) );
  XNOR U4322 ( .A(n3059), .B(n3079), .Z(n3062) );
  OR U4323 ( .A(n3053), .B(n3062), .Z(n3054) );
  XNOR U4324 ( .A(n3072), .B(n3054), .Z(n4021) );
  OR U4325 ( .A(n3056), .B(n3055), .Z(n3067) );
  XNOR U4326 ( .A(n4021), .B(n3067), .Z(n3057) );
  XOR U4327 ( .A(n3058), .B(n3057), .Z(n4018) );
  NANDN U4328 ( .A(n3060), .B(n3059), .Z(n4004) );
  OR U4329 ( .A(n3062), .B(n3061), .Z(n3063) );
  XOR U4330 ( .A(n4004), .B(n3063), .Z(n3073) );
  XOR U4331 ( .A(n3073), .B(n3064), .Z(n4007) );
  XOR U4332 ( .A(n4018), .B(n4007), .Z(n4036) );
  ANDN U4333 ( .B(n3077), .A(n3065), .Z(n3069) );
  XNOR U4334 ( .A(n3067), .B(n3066), .Z(n3068) );
  XNOR U4335 ( .A(n3069), .B(n3068), .Z(n3075) );
  NANDN U4336 ( .A(n3070), .B(n3079), .Z(n3071) );
  XNOR U4337 ( .A(n3072), .B(n3071), .Z(n4014) );
  XOR U4338 ( .A(n3073), .B(n4014), .Z(n3074) );
  XOR U4339 ( .A(n3075), .B(n3074), .Z(n4017) );
  XNOR U4340 ( .A(n4036), .B(n4017), .Z(z[89]) );
  ANDN U4341 ( .B(n3077), .A(n3076), .Z(n4024) );
  ANDN U4342 ( .B(n3079), .A(n3078), .Z(n4006) );
  XNOR U4343 ( .A(n4004), .B(z[89]), .Z(n3080) );
  XNOR U4344 ( .A(n4006), .B(n3080), .Z(n3081) );
  XOR U4345 ( .A(n4022), .B(n3081), .Z(n3082) );
  XOR U4346 ( .A(n4024), .B(n3082), .Z(z[95]) );
  IV U4347 ( .A(x[97]), .Z(n3436) );
  IV U4348 ( .A(x[96]), .Z(n3105) );
  XNOR U4349 ( .A(n3105), .B(x[102]), .Z(n3083) );
  XNOR U4350 ( .A(x[101]), .B(n3083), .Z(n3437) );
  IV U4351 ( .A(n3437), .Z(n3085) );
  ANDN U4352 ( .B(n3436), .A(n3085), .Z(n3091) );
  XOR U4353 ( .A(x[97]), .B(x[103]), .Z(n3434) );
  XOR U4354 ( .A(x[97]), .B(x[99]), .Z(n3084) );
  XOR U4355 ( .A(n3430), .B(n3437), .Z(n3142) );
  NAND U4356 ( .A(n3434), .B(n3142), .Z(n3094) );
  XNOR U4357 ( .A(x[103]), .B(x[100]), .Z(n3443) );
  IV U4358 ( .A(n3443), .Z(n3088) );
  XOR U4359 ( .A(n3084), .B(n3088), .Z(n3108) );
  IV U4360 ( .A(n3108), .Z(n3124) );
  XOR U4361 ( .A(n3124), .B(n3142), .Z(n3459) );
  IV U4362 ( .A(x[100]), .Z(n3097) );
  XOR U4363 ( .A(x[98]), .B(n3097), .Z(n3445) );
  NOR U4364 ( .A(n3459), .B(n3445), .Z(n3087) );
  XOR U4365 ( .A(x[103]), .B(n3085), .Z(n3462) );
  XOR U4366 ( .A(n3430), .B(n3462), .Z(n3086) );
  XNOR U4367 ( .A(n3087), .B(n3086), .Z(n3089) );
  XNOR U4368 ( .A(n3105), .B(n3430), .Z(n3429) );
  ANDN U4369 ( .B(n3088), .A(n3429), .Z(n3093) );
  XNOR U4370 ( .A(n3089), .B(n3093), .Z(n3113) );
  XNOR U4371 ( .A(n3094), .B(n3113), .Z(n3090) );
  XNOR U4372 ( .A(n3091), .B(n3090), .Z(n3128) );
  NANDN U4373 ( .A(n3462), .B(n3430), .Z(n3096) );
  XOR U4374 ( .A(x[96]), .B(n3124), .Z(n3125) );
  XNOR U4375 ( .A(n3437), .B(n3125), .Z(n3428) );
  OR U4376 ( .A(n3465), .B(n3428), .Z(n3092) );
  XOR U4377 ( .A(n3093), .B(n3092), .Z(n3101) );
  XNOR U4378 ( .A(n3101), .B(n3094), .Z(n3095) );
  XNOR U4379 ( .A(n3096), .B(n3095), .Z(n3119) );
  XOR U4380 ( .A(x[98]), .B(n3436), .Z(n3104) );
  XNOR U4381 ( .A(n3443), .B(n3104), .Z(n3454) );
  OR U4382 ( .A(n3454), .B(n3124), .Z(n3106) );
  XOR U4383 ( .A(n3097), .B(n3437), .Z(n3472) );
  NOR U4384 ( .A(n3105), .B(n3472), .Z(n3099) );
  XNOR U4385 ( .A(x[98]), .B(n3108), .Z(n3098) );
  XNOR U4386 ( .A(n3099), .B(n3098), .Z(n3100) );
  XNOR U4387 ( .A(n3106), .B(n3100), .Z(n3103) );
  XOR U4388 ( .A(n3101), .B(n3462), .Z(n3102) );
  XNOR U4389 ( .A(n3103), .B(n3102), .Z(n3131) );
  IV U4390 ( .A(n3131), .Z(n3134) );
  NANDN U4391 ( .A(n3119), .B(n3134), .Z(n3136) );
  XNOR U4392 ( .A(n3462), .B(n3104), .Z(n3452) );
  ANDN U4393 ( .B(n3105), .A(n3452), .Z(n3107) );
  XOR U4394 ( .A(n3107), .B(n3106), .Z(n3110) );
  NANDN U4395 ( .A(n3108), .B(n3452), .Z(n3109) );
  NAND U4396 ( .A(n3110), .B(n3109), .Z(n3111) );
  XNOR U4397 ( .A(n3111), .B(n3472), .Z(n3112) );
  XOR U4398 ( .A(n3113), .B(n3112), .Z(n3139) );
  IV U4399 ( .A(n3139), .Z(n3135) );
  XNOR U4400 ( .A(n3136), .B(n3135), .Z(n3114) );
  NANDN U4401 ( .A(n3128), .B(n3114), .Z(n3116) );
  IV U4402 ( .A(n3128), .Z(n3137) );
  ANDN U4403 ( .B(n3119), .A(n3137), .Z(n3115) );
  ANDN U4404 ( .B(n3116), .A(n3115), .Z(n3451) );
  IV U4405 ( .A(n3119), .Z(n3129) );
  NANDN U4406 ( .A(n3129), .B(n3134), .Z(n3117) );
  NANDN U4407 ( .A(n3137), .B(n3117), .Z(n3121) );
  XNOR U4408 ( .A(n3134), .B(n3139), .Z(n3118) );
  NANDN U4409 ( .A(n3119), .B(n3118), .Z(n3120) );
  NAND U4410 ( .A(n3121), .B(n3120), .Z(n3471) );
  OR U4411 ( .A(n3451), .B(n3471), .Z(n3123) );
  NANDN U4412 ( .A(n3137), .B(n3129), .Z(n3122) );
  NAND U4413 ( .A(n3123), .B(n3122), .Z(n3453) );
  OR U4414 ( .A(n3453), .B(n3124), .Z(n3448) );
  OR U4415 ( .A(n3451), .B(n3125), .Z(n3126) );
  XNOR U4416 ( .A(n3448), .B(n3126), .Z(n3461) );
  NANDN U4417 ( .A(n3134), .B(n3129), .Z(n3127) );
  NANDN U4418 ( .A(n3135), .B(n3127), .Z(n3133) );
  XNOR U4419 ( .A(n3129), .B(n3128), .Z(n3130) );
  NANDN U4420 ( .A(n3131), .B(n3130), .Z(n3132) );
  AND U4421 ( .A(n3133), .B(n3132), .Z(n3463) );
  NANDN U4422 ( .A(n3135), .B(n3134), .Z(n3141) );
  XOR U4423 ( .A(n3137), .B(n3136), .Z(n3138) );
  NANDN U4424 ( .A(n3139), .B(n3138), .Z(n3140) );
  AND U4425 ( .A(n3141), .B(n3140), .Z(n3438) );
  XNOR U4426 ( .A(n3463), .B(n3438), .Z(n3435) );
  NANDN U4427 ( .A(n3435), .B(n3142), .Z(n3432) );
  ANDN U4428 ( .B(n3438), .A(n3437), .Z(n3143) );
  XNOR U4429 ( .A(n3432), .B(n3143), .Z(n3480) );
  XOR U4430 ( .A(n3461), .B(n3480), .Z(z[98]) );
  IV U4431 ( .A(x[108]), .Z(n3144) );
  IV U4432 ( .A(x[104]), .Z(n3229) );
  XOR U4433 ( .A(n3229), .B(x[110]), .Z(n3145) );
  XOR U4434 ( .A(n3145), .B(x[109]), .Z(n3169) );
  IV U4435 ( .A(n3169), .Z(n3511) );
  XOR U4436 ( .A(n3144), .B(n3511), .Z(n3218) );
  XOR U4437 ( .A(x[105]), .B(x[107]), .Z(n3146) );
  XOR U4438 ( .A(x[111]), .B(n3144), .Z(n3204) );
  XNOR U4439 ( .A(n3146), .B(n3204), .Z(n3183) );
  IV U4440 ( .A(n3183), .Z(n3161) );
  XOR U4441 ( .A(n3146), .B(n3145), .Z(n3147) );
  XOR U4442 ( .A(x[106]), .B(n3147), .Z(n3488) );
  XOR U4443 ( .A(n3488), .B(n3169), .Z(n3201) );
  XOR U4444 ( .A(n3161), .B(n3201), .Z(n3214) );
  IV U4445 ( .A(x[106]), .Z(n3157) );
  XOR U4446 ( .A(x[108]), .B(n3157), .Z(n3206) );
  NOR U4447 ( .A(n3214), .B(n3206), .Z(n3149) );
  XOR U4448 ( .A(x[111]), .B(n3511), .Z(n3496) );
  XOR U4449 ( .A(n3488), .B(n3496), .Z(n3148) );
  XNOR U4450 ( .A(n3149), .B(n3148), .Z(n3150) );
  XNOR U4451 ( .A(n3229), .B(n3488), .Z(n3213) );
  NOR U4452 ( .A(n3204), .B(n3213), .Z(n3159) );
  XNOR U4453 ( .A(n3150), .B(n3159), .Z(n3171) );
  IV U4454 ( .A(x[105]), .Z(n3510) );
  XNOR U4455 ( .A(n3510), .B(x[106]), .Z(n3151) );
  XNOR U4456 ( .A(n3496), .B(n3151), .Z(n3203) );
  ANDN U4457 ( .B(n3203), .A(x[104]), .Z(n3152) );
  XNOR U4458 ( .A(n3204), .B(n3151), .Z(n3208) );
  NANDN U4459 ( .A(n3161), .B(n3208), .Z(n3162) );
  XOR U4460 ( .A(n3152), .B(n3162), .Z(n3154) );
  OR U4461 ( .A(n3203), .B(n3183), .Z(n3153) );
  NAND U4462 ( .A(n3154), .B(n3153), .Z(n3155) );
  XOR U4463 ( .A(n3171), .B(n3155), .Z(n3156) );
  XOR U4464 ( .A(n3218), .B(n3156), .Z(n3197) );
  XNOR U4465 ( .A(n3161), .B(x[104]), .Z(n3184) );
  XNOR U4466 ( .A(n3511), .B(n3184), .Z(n3231) );
  IV U4467 ( .A(x[111]), .Z(n3160) );
  XOR U4468 ( .A(n3160), .B(n3157), .Z(n3223) );
  NANDN U4469 ( .A(n3231), .B(n3223), .Z(n3158) );
  XOR U4470 ( .A(n3159), .B(n3158), .Z(n3166) );
  XOR U4471 ( .A(n3510), .B(n3160), .Z(n3497) );
  NAND U4472 ( .A(n3201), .B(n3497), .Z(n3170) );
  ANDN U4473 ( .B(n3218), .A(n3229), .Z(n3164) );
  XNOR U4474 ( .A(n3162), .B(n3161), .Z(n3163) );
  XNOR U4475 ( .A(n3164), .B(n3163), .Z(n3165) );
  XNOR U4476 ( .A(n3166), .B(n3165), .Z(n3168) );
  XNOR U4477 ( .A(x[106]), .B(n3496), .Z(n3167) );
  XNOR U4478 ( .A(n3168), .B(n3167), .Z(n3198) );
  IV U4479 ( .A(n3198), .Z(n3190) );
  AND U4480 ( .A(n3193), .B(n3190), .Z(n3186) );
  XOR U4481 ( .A(n3197), .B(n3186), .Z(n3174) );
  ANDN U4482 ( .B(n3169), .A(x[105]), .Z(n3173) );
  XNOR U4483 ( .A(n3171), .B(n3170), .Z(n3172) );
  XNOR U4484 ( .A(n3173), .B(n3172), .Z(n3192) );
  ANDN U4485 ( .B(n3174), .A(n3192), .Z(n3181) );
  IV U4486 ( .A(n3193), .Z(n3178) );
  NANDN U4487 ( .A(n3178), .B(n3192), .Z(n3175) );
  NANDN U4488 ( .A(n3181), .B(n3175), .Z(n3205) );
  NANDN U4489 ( .A(n3193), .B(n3190), .Z(n3176) );
  NAND U4490 ( .A(n3176), .B(n3192), .Z(n3180) );
  XNOR U4491 ( .A(n3190), .B(n3197), .Z(n3177) );
  NANDN U4492 ( .A(n3178), .B(n3177), .Z(n3179) );
  AND U4493 ( .A(n3180), .B(n3179), .Z(n3230) );
  OR U4494 ( .A(n3205), .B(n3230), .Z(n3182) );
  ANDN U4495 ( .B(n3182), .A(n3181), .Z(n3209) );
  NANDN U4496 ( .A(n3209), .B(n3183), .Z(n3507) );
  NANDN U4497 ( .A(n3205), .B(n3184), .Z(n3185) );
  XOR U4498 ( .A(n3507), .B(n3185), .Z(n3217) );
  NANDN U4499 ( .A(n3190), .B(n3197), .Z(n3189) );
  XNOR U4500 ( .A(n3186), .B(n3192), .Z(n3187) );
  NANDN U4501 ( .A(n3197), .B(n3187), .Z(n3188) );
  AND U4502 ( .A(n3189), .B(n3188), .Z(n3513) );
  NANDN U4503 ( .A(n3190), .B(n3193), .Z(n3191) );
  NAND U4504 ( .A(n3197), .B(n3191), .Z(n3196) );
  XNOR U4505 ( .A(n3193), .B(n3192), .Z(n3194) );
  NANDN U4506 ( .A(n3198), .B(n3194), .Z(n3195) );
  NAND U4507 ( .A(n3196), .B(n3195), .Z(n3495) );
  IV U4508 ( .A(n3495), .Z(n3487) );
  NANDN U4509 ( .A(n3513), .B(n3487), .Z(n3200) );
  NANDN U4510 ( .A(n3198), .B(n3197), .Z(n3199) );
  NAND U4511 ( .A(n3200), .B(n3199), .Z(n3498) );
  NANDN U4512 ( .A(n3498), .B(n3201), .Z(n3490) );
  NANDN U4513 ( .A(n3513), .B(n3511), .Z(n3202) );
  XNOR U4514 ( .A(n3490), .B(n3202), .Z(n3219) );
  XOR U4515 ( .A(n3217), .B(n3219), .Z(z[106]) );
  NOR U4516 ( .A(n3205), .B(n3203), .Z(n3211) );
  XOR U4517 ( .A(n3487), .B(n3230), .Z(n3212) );
  NANDN U4518 ( .A(n3204), .B(n3212), .Z(n3225) );
  XOR U4519 ( .A(n3205), .B(n3513), .Z(n3232) );
  XNOR U4520 ( .A(n3212), .B(n3232), .Z(n3215) );
  OR U4521 ( .A(n3206), .B(n3215), .Z(n3207) );
  XNOR U4522 ( .A(n3225), .B(n3207), .Z(n3506) );
  NANDN U4523 ( .A(n3209), .B(n3208), .Z(n3220) );
  XNOR U4524 ( .A(n3506), .B(n3220), .Z(n3210) );
  XOR U4525 ( .A(n3211), .B(n3210), .Z(n3503) );
  NANDN U4526 ( .A(n3213), .B(n3212), .Z(n3491) );
  OR U4527 ( .A(n3215), .B(n3214), .Z(n3216) );
  XOR U4528 ( .A(n3491), .B(n3216), .Z(n3226) );
  XOR U4529 ( .A(n3226), .B(n3217), .Z(n3494) );
  XOR U4530 ( .A(n3503), .B(n3494), .Z(n3521) );
  ANDN U4531 ( .B(n3230), .A(n3218), .Z(n3222) );
  XNOR U4532 ( .A(n3220), .B(n3219), .Z(n3221) );
  XNOR U4533 ( .A(n3222), .B(n3221), .Z(n3228) );
  NAND U4534 ( .A(n3223), .B(n3232), .Z(n3224) );
  XNOR U4535 ( .A(n3225), .B(n3224), .Z(n3499) );
  XOR U4536 ( .A(n3226), .B(n3499), .Z(n3227) );
  XOR U4537 ( .A(n3228), .B(n3227), .Z(n3502) );
  XNOR U4538 ( .A(n3521), .B(n3502), .Z(z[105]) );
  ANDN U4539 ( .B(n3230), .A(n3229), .Z(n3509) );
  ANDN U4540 ( .B(n3232), .A(n3231), .Z(n3493) );
  XNOR U4541 ( .A(n3491), .B(z[105]), .Z(n3233) );
  XNOR U4542 ( .A(n3493), .B(n3233), .Z(n3234) );
  XOR U4543 ( .A(n3507), .B(n3234), .Z(n3235) );
  XOR U4544 ( .A(n3509), .B(n3235), .Z(z[111]) );
  IV U4545 ( .A(x[116]), .Z(n3236) );
  IV U4546 ( .A(x[112]), .Z(n3321) );
  XOR U4547 ( .A(n3321), .B(x[118]), .Z(n3237) );
  XOR U4548 ( .A(n3237), .B(x[117]), .Z(n3261) );
  IV U4549 ( .A(n3261), .Z(n3546) );
  XOR U4550 ( .A(n3236), .B(n3546), .Z(n3310) );
  XOR U4551 ( .A(x[113]), .B(x[115]), .Z(n3238) );
  XOR U4552 ( .A(x[119]), .B(n3236), .Z(n3296) );
  XNOR U4553 ( .A(n3238), .B(n3296), .Z(n3275) );
  IV U4554 ( .A(n3275), .Z(n3253) );
  XOR U4555 ( .A(n3238), .B(n3237), .Z(n3239) );
  XOR U4556 ( .A(x[114]), .B(n3239), .Z(n3523) );
  XOR U4557 ( .A(n3523), .B(n3261), .Z(n3293) );
  XOR U4558 ( .A(n3253), .B(n3293), .Z(n3306) );
  IV U4559 ( .A(x[114]), .Z(n3249) );
  XOR U4560 ( .A(x[116]), .B(n3249), .Z(n3298) );
  NOR U4561 ( .A(n3306), .B(n3298), .Z(n3241) );
  XOR U4562 ( .A(x[119]), .B(n3546), .Z(n3531) );
  XOR U4563 ( .A(n3523), .B(n3531), .Z(n3240) );
  XNOR U4564 ( .A(n3241), .B(n3240), .Z(n3242) );
  XNOR U4565 ( .A(n3321), .B(n3523), .Z(n3305) );
  NOR U4566 ( .A(n3296), .B(n3305), .Z(n3251) );
  XNOR U4567 ( .A(n3242), .B(n3251), .Z(n3263) );
  IV U4568 ( .A(x[113]), .Z(n3545) );
  XNOR U4569 ( .A(n3545), .B(x[114]), .Z(n3243) );
  XNOR U4570 ( .A(n3531), .B(n3243), .Z(n3295) );
  ANDN U4571 ( .B(n3295), .A(x[112]), .Z(n3244) );
  XNOR U4572 ( .A(n3296), .B(n3243), .Z(n3300) );
  NANDN U4573 ( .A(n3253), .B(n3300), .Z(n3254) );
  XOR U4574 ( .A(n3244), .B(n3254), .Z(n3246) );
  OR U4575 ( .A(n3295), .B(n3275), .Z(n3245) );
  NAND U4576 ( .A(n3246), .B(n3245), .Z(n3247) );
  XOR U4577 ( .A(n3263), .B(n3247), .Z(n3248) );
  XOR U4578 ( .A(n3310), .B(n3248), .Z(n3289) );
  XNOR U4579 ( .A(n3253), .B(x[112]), .Z(n3276) );
  XNOR U4580 ( .A(n3546), .B(n3276), .Z(n3323) );
  IV U4581 ( .A(x[119]), .Z(n3252) );
  XOR U4582 ( .A(n3252), .B(n3249), .Z(n3315) );
  NANDN U4583 ( .A(n3323), .B(n3315), .Z(n3250) );
  XOR U4584 ( .A(n3251), .B(n3250), .Z(n3258) );
  XOR U4585 ( .A(n3545), .B(n3252), .Z(n3532) );
  NAND U4586 ( .A(n3293), .B(n3532), .Z(n3262) );
  ANDN U4587 ( .B(n3310), .A(n3321), .Z(n3256) );
  XNOR U4588 ( .A(n3254), .B(n3253), .Z(n3255) );
  XNOR U4589 ( .A(n3256), .B(n3255), .Z(n3257) );
  XNOR U4590 ( .A(n3258), .B(n3257), .Z(n3260) );
  XNOR U4591 ( .A(x[114]), .B(n3531), .Z(n3259) );
  XNOR U4592 ( .A(n3260), .B(n3259), .Z(n3290) );
  IV U4593 ( .A(n3290), .Z(n3282) );
  AND U4594 ( .A(n3285), .B(n3282), .Z(n3278) );
  XOR U4595 ( .A(n3289), .B(n3278), .Z(n3266) );
  ANDN U4596 ( .B(n3261), .A(x[113]), .Z(n3265) );
  XNOR U4597 ( .A(n3263), .B(n3262), .Z(n3264) );
  XNOR U4598 ( .A(n3265), .B(n3264), .Z(n3284) );
  ANDN U4599 ( .B(n3266), .A(n3284), .Z(n3273) );
  IV U4600 ( .A(n3285), .Z(n3270) );
  NANDN U4601 ( .A(n3270), .B(n3284), .Z(n3267) );
  NANDN U4602 ( .A(n3273), .B(n3267), .Z(n3297) );
  NANDN U4603 ( .A(n3285), .B(n3282), .Z(n3268) );
  NAND U4604 ( .A(n3268), .B(n3284), .Z(n3272) );
  XNOR U4605 ( .A(n3282), .B(n3289), .Z(n3269) );
  NANDN U4606 ( .A(n3270), .B(n3269), .Z(n3271) );
  AND U4607 ( .A(n3272), .B(n3271), .Z(n3322) );
  OR U4608 ( .A(n3297), .B(n3322), .Z(n3274) );
  ANDN U4609 ( .B(n3274), .A(n3273), .Z(n3301) );
  NANDN U4610 ( .A(n3301), .B(n3275), .Z(n3542) );
  NANDN U4611 ( .A(n3297), .B(n3276), .Z(n3277) );
  XOR U4612 ( .A(n3542), .B(n3277), .Z(n3309) );
  NANDN U4613 ( .A(n3282), .B(n3289), .Z(n3281) );
  XNOR U4614 ( .A(n3278), .B(n3284), .Z(n3279) );
  NANDN U4615 ( .A(n3289), .B(n3279), .Z(n3280) );
  AND U4616 ( .A(n3281), .B(n3280), .Z(n3548) );
  NANDN U4617 ( .A(n3282), .B(n3285), .Z(n3283) );
  NAND U4618 ( .A(n3289), .B(n3283), .Z(n3288) );
  XNOR U4619 ( .A(n3285), .B(n3284), .Z(n3286) );
  NANDN U4620 ( .A(n3290), .B(n3286), .Z(n3287) );
  NAND U4621 ( .A(n3288), .B(n3287), .Z(n3530) );
  IV U4622 ( .A(n3530), .Z(n3522) );
  NANDN U4623 ( .A(n3548), .B(n3522), .Z(n3292) );
  NANDN U4624 ( .A(n3290), .B(n3289), .Z(n3291) );
  NAND U4625 ( .A(n3292), .B(n3291), .Z(n3533) );
  NANDN U4626 ( .A(n3533), .B(n3293), .Z(n3525) );
  NANDN U4627 ( .A(n3548), .B(n3546), .Z(n3294) );
  XNOR U4628 ( .A(n3525), .B(n3294), .Z(n3311) );
  XOR U4629 ( .A(n3309), .B(n3311), .Z(z[114]) );
  NOR U4630 ( .A(n3297), .B(n3295), .Z(n3303) );
  XOR U4631 ( .A(n3522), .B(n3322), .Z(n3304) );
  NANDN U4632 ( .A(n3296), .B(n3304), .Z(n3317) );
  XOR U4633 ( .A(n3297), .B(n3548), .Z(n3324) );
  XNOR U4634 ( .A(n3304), .B(n3324), .Z(n3307) );
  OR U4635 ( .A(n3298), .B(n3307), .Z(n3299) );
  XNOR U4636 ( .A(n3317), .B(n3299), .Z(n3541) );
  NANDN U4637 ( .A(n3301), .B(n3300), .Z(n3312) );
  XNOR U4638 ( .A(n3541), .B(n3312), .Z(n3302) );
  XOR U4639 ( .A(n3303), .B(n3302), .Z(n3538) );
  NANDN U4640 ( .A(n3305), .B(n3304), .Z(n3526) );
  OR U4641 ( .A(n3307), .B(n3306), .Z(n3308) );
  XOR U4642 ( .A(n3526), .B(n3308), .Z(n3318) );
  XOR U4643 ( .A(n3318), .B(n3309), .Z(n3529) );
  XOR U4644 ( .A(n3538), .B(n3529), .Z(n3556) );
  ANDN U4645 ( .B(n3322), .A(n3310), .Z(n3314) );
  XNOR U4646 ( .A(n3312), .B(n3311), .Z(n3313) );
  XNOR U4647 ( .A(n3314), .B(n3313), .Z(n3320) );
  NAND U4648 ( .A(n3315), .B(n3324), .Z(n3316) );
  XNOR U4649 ( .A(n3317), .B(n3316), .Z(n3534) );
  XOR U4650 ( .A(n3318), .B(n3534), .Z(n3319) );
  XOR U4651 ( .A(n3320), .B(n3319), .Z(n3537) );
  XNOR U4652 ( .A(n3556), .B(n3537), .Z(z[113]) );
  ANDN U4653 ( .B(n3322), .A(n3321), .Z(n3544) );
  ANDN U4654 ( .B(n3324), .A(n3323), .Z(n3528) );
  XNOR U4655 ( .A(n3526), .B(z[113]), .Z(n3325) );
  XNOR U4656 ( .A(n3528), .B(n3325), .Z(n3326) );
  XOR U4657 ( .A(n3542), .B(n3326), .Z(n3327) );
  XOR U4658 ( .A(n3544), .B(n3327), .Z(z[119]) );
  IV U4659 ( .A(x[124]), .Z(n3328) );
  IV U4660 ( .A(x[120]), .Z(n3413) );
  XOR U4661 ( .A(n3413), .B(x[126]), .Z(n3329) );
  XOR U4662 ( .A(n3329), .B(x[125]), .Z(n3353) );
  IV U4663 ( .A(n3353), .Z(n3612) );
  XOR U4664 ( .A(n3328), .B(n3612), .Z(n3402) );
  XOR U4665 ( .A(x[121]), .B(x[123]), .Z(n3330) );
  XOR U4666 ( .A(x[127]), .B(n3328), .Z(n3388) );
  XNOR U4667 ( .A(n3330), .B(n3388), .Z(n3367) );
  IV U4668 ( .A(n3367), .Z(n3345) );
  XOR U4669 ( .A(n3330), .B(n3329), .Z(n3331) );
  XOR U4670 ( .A(x[122]), .B(n3331), .Z(n3589) );
  XOR U4671 ( .A(n3589), .B(n3353), .Z(n3385) );
  XOR U4672 ( .A(n3345), .B(n3385), .Z(n3398) );
  IV U4673 ( .A(x[122]), .Z(n3341) );
  XOR U4674 ( .A(x[124]), .B(n3341), .Z(n3390) );
  NOR U4675 ( .A(n3398), .B(n3390), .Z(n3333) );
  XOR U4676 ( .A(x[127]), .B(n3612), .Z(n3597) );
  XOR U4677 ( .A(n3589), .B(n3597), .Z(n3332) );
  XNOR U4678 ( .A(n3333), .B(n3332), .Z(n3334) );
  XNOR U4679 ( .A(n3413), .B(n3589), .Z(n3397) );
  NOR U4680 ( .A(n3388), .B(n3397), .Z(n3343) );
  XNOR U4681 ( .A(n3334), .B(n3343), .Z(n3355) );
  IV U4682 ( .A(x[121]), .Z(n3611) );
  XNOR U4683 ( .A(n3611), .B(x[122]), .Z(n3335) );
  XNOR U4684 ( .A(n3597), .B(n3335), .Z(n3387) );
  ANDN U4685 ( .B(n3387), .A(x[120]), .Z(n3336) );
  XNOR U4686 ( .A(n3388), .B(n3335), .Z(n3392) );
  NANDN U4687 ( .A(n3345), .B(n3392), .Z(n3346) );
  XOR U4688 ( .A(n3336), .B(n3346), .Z(n3338) );
  OR U4689 ( .A(n3387), .B(n3367), .Z(n3337) );
  NAND U4690 ( .A(n3338), .B(n3337), .Z(n3339) );
  XOR U4691 ( .A(n3355), .B(n3339), .Z(n3340) );
  XOR U4692 ( .A(n3402), .B(n3340), .Z(n3381) );
  XNOR U4693 ( .A(n3345), .B(x[120]), .Z(n3368) );
  XNOR U4694 ( .A(n3612), .B(n3368), .Z(n3415) );
  IV U4695 ( .A(x[127]), .Z(n3344) );
  XOR U4696 ( .A(n3344), .B(n3341), .Z(n3407) );
  NANDN U4697 ( .A(n3415), .B(n3407), .Z(n3342) );
  XOR U4698 ( .A(n3343), .B(n3342), .Z(n3350) );
  XOR U4699 ( .A(n3611), .B(n3344), .Z(n3598) );
  NAND U4700 ( .A(n3385), .B(n3598), .Z(n3354) );
  ANDN U4701 ( .B(n3402), .A(n3413), .Z(n3348) );
  XNOR U4702 ( .A(n3346), .B(n3345), .Z(n3347) );
  XNOR U4703 ( .A(n3348), .B(n3347), .Z(n3349) );
  XNOR U4704 ( .A(n3350), .B(n3349), .Z(n3352) );
  XNOR U4705 ( .A(x[122]), .B(n3597), .Z(n3351) );
  XNOR U4706 ( .A(n3352), .B(n3351), .Z(n3382) );
  IV U4707 ( .A(n3382), .Z(n3374) );
  AND U4708 ( .A(n3377), .B(n3374), .Z(n3370) );
  XOR U4709 ( .A(n3381), .B(n3370), .Z(n3358) );
  ANDN U4710 ( .B(n3353), .A(x[121]), .Z(n3357) );
  XNOR U4711 ( .A(n3355), .B(n3354), .Z(n3356) );
  XNOR U4712 ( .A(n3357), .B(n3356), .Z(n3376) );
  ANDN U4713 ( .B(n3358), .A(n3376), .Z(n3365) );
  IV U4714 ( .A(n3377), .Z(n3362) );
  NANDN U4715 ( .A(n3362), .B(n3376), .Z(n3359) );
  NANDN U4716 ( .A(n3365), .B(n3359), .Z(n3389) );
  NANDN U4717 ( .A(n3377), .B(n3374), .Z(n3360) );
  NAND U4718 ( .A(n3360), .B(n3376), .Z(n3364) );
  XNOR U4719 ( .A(n3374), .B(n3381), .Z(n3361) );
  NANDN U4720 ( .A(n3362), .B(n3361), .Z(n3363) );
  AND U4721 ( .A(n3364), .B(n3363), .Z(n3414) );
  OR U4722 ( .A(n3389), .B(n3414), .Z(n3366) );
  ANDN U4723 ( .B(n3366), .A(n3365), .Z(n3393) );
  NANDN U4724 ( .A(n3393), .B(n3367), .Z(n3608) );
  NANDN U4725 ( .A(n3389), .B(n3368), .Z(n3369) );
  XOR U4726 ( .A(n3608), .B(n3369), .Z(n3401) );
  NANDN U4727 ( .A(n3374), .B(n3381), .Z(n3373) );
  XNOR U4728 ( .A(n3370), .B(n3376), .Z(n3371) );
  NANDN U4729 ( .A(n3381), .B(n3371), .Z(n3372) );
  AND U4730 ( .A(n3373), .B(n3372), .Z(n3614) );
  NANDN U4731 ( .A(n3374), .B(n3377), .Z(n3375) );
  NAND U4732 ( .A(n3381), .B(n3375), .Z(n3380) );
  XNOR U4733 ( .A(n3377), .B(n3376), .Z(n3378) );
  NANDN U4734 ( .A(n3382), .B(n3378), .Z(n3379) );
  NAND U4735 ( .A(n3380), .B(n3379), .Z(n3596) );
  IV U4736 ( .A(n3596), .Z(n3588) );
  NANDN U4737 ( .A(n3614), .B(n3588), .Z(n3384) );
  NANDN U4738 ( .A(n3382), .B(n3381), .Z(n3383) );
  NAND U4739 ( .A(n3384), .B(n3383), .Z(n3599) );
  NANDN U4740 ( .A(n3599), .B(n3385), .Z(n3591) );
  NANDN U4741 ( .A(n3614), .B(n3612), .Z(n3386) );
  XNOR U4742 ( .A(n3591), .B(n3386), .Z(n3403) );
  XOR U4743 ( .A(n3401), .B(n3403), .Z(z[122]) );
  NOR U4744 ( .A(n3389), .B(n3387), .Z(n3395) );
  XOR U4745 ( .A(n3588), .B(n3414), .Z(n3396) );
  NANDN U4746 ( .A(n3388), .B(n3396), .Z(n3409) );
  XOR U4747 ( .A(n3389), .B(n3614), .Z(n3416) );
  XNOR U4748 ( .A(n3396), .B(n3416), .Z(n3399) );
  OR U4749 ( .A(n3390), .B(n3399), .Z(n3391) );
  XNOR U4750 ( .A(n3409), .B(n3391), .Z(n3607) );
  NANDN U4751 ( .A(n3393), .B(n3392), .Z(n3404) );
  XNOR U4752 ( .A(n3607), .B(n3404), .Z(n3394) );
  XOR U4753 ( .A(n3395), .B(n3394), .Z(n3604) );
  NANDN U4754 ( .A(n3397), .B(n3396), .Z(n3592) );
  OR U4755 ( .A(n3399), .B(n3398), .Z(n3400) );
  XOR U4756 ( .A(n3592), .B(n3400), .Z(n3410) );
  XOR U4757 ( .A(n3410), .B(n3401), .Z(n3595) );
  XOR U4758 ( .A(n3604), .B(n3595), .Z(n3622) );
  ANDN U4759 ( .B(n3414), .A(n3402), .Z(n3406) );
  XNOR U4760 ( .A(n3404), .B(n3403), .Z(n3405) );
  XNOR U4761 ( .A(n3406), .B(n3405), .Z(n3412) );
  NAND U4762 ( .A(n3407), .B(n3416), .Z(n3408) );
  XNOR U4763 ( .A(n3409), .B(n3408), .Z(n3600) );
  XOR U4764 ( .A(n3410), .B(n3600), .Z(n3411) );
  XOR U4765 ( .A(n3412), .B(n3411), .Z(n3603) );
  XNOR U4766 ( .A(n3622), .B(n3603), .Z(z[121]) );
  ANDN U4767 ( .B(n3414), .A(n3413), .Z(n3610) );
  ANDN U4768 ( .B(n3416), .A(n3415), .Z(n3594) );
  XNOR U4769 ( .A(n3592), .B(z[121]), .Z(n3417) );
  XNOR U4770 ( .A(n3594), .B(n3417), .Z(n3418) );
  XOR U4771 ( .A(n3608), .B(n3418), .Z(n3419) );
  XOR U4772 ( .A(n3610), .B(n3419), .Z(z[127]) );
  NANDN U4773 ( .A(n3421), .B(n3420), .Z(n3422) );
  XNOR U4774 ( .A(n3423), .B(n3422), .Z(n3873) );
  XNOR U4775 ( .A(n3424), .B(n3873), .Z(n3425) );
  XOR U4776 ( .A(n3426), .B(n3425), .Z(n3816) );
  XOR U4777 ( .A(n3816), .B(n3427), .Z(z[0]) );
  XNOR U4778 ( .A(n3438), .B(n3451), .Z(n3464) );
  ANDN U4779 ( .B(n3464), .A(n3428), .Z(n3485) );
  NANDN U4780 ( .A(n3429), .B(n3444), .Z(n3483) );
  NANDN U4781 ( .A(n3430), .B(n3463), .Z(n3431) );
  XNOR U4782 ( .A(n3432), .B(n3431), .Z(n3442) );
  XNOR U4783 ( .A(n3483), .B(n3442), .Z(n3433) );
  XOR U4784 ( .A(n3485), .B(n3433), .Z(n4038) );
  XNOR U4785 ( .A(n4038), .B(z[98]), .Z(z[100]) );
  NANDN U4786 ( .A(n3435), .B(n3434), .Z(n3468) );
  XOR U4787 ( .A(n3437), .B(n3436), .Z(n3439) );
  NAND U4788 ( .A(n3439), .B(n3438), .Z(n3440) );
  XOR U4789 ( .A(n3468), .B(n3440), .Z(n3441) );
  XNOR U4790 ( .A(n3442), .B(n3441), .Z(n3450) );
  NANDN U4791 ( .A(n3443), .B(n3444), .Z(n3467) );
  XNOR U4792 ( .A(n3444), .B(n3464), .Z(n3458) );
  OR U4793 ( .A(n3458), .B(n3445), .Z(n3446) );
  XNOR U4794 ( .A(n3467), .B(n3446), .Z(n3455) );
  NANDN U4795 ( .A(n3471), .B(x[96]), .Z(n3447) );
  XNOR U4796 ( .A(n3448), .B(n3447), .Z(n3482) );
  XNOR U4797 ( .A(n3455), .B(n3482), .Z(n3449) );
  XOR U4798 ( .A(n3450), .B(n3449), .Z(z[101]) );
  ANDN U4799 ( .B(n3452), .A(n3451), .Z(n3457) );
  OR U4800 ( .A(n3454), .B(n3453), .Z(n3477) );
  XNOR U4801 ( .A(n3477), .B(n3455), .Z(n3456) );
  XOR U4802 ( .A(n3457), .B(n3456), .Z(n4039) );
  OR U4803 ( .A(n3459), .B(n3458), .Z(n3460) );
  XOR U4804 ( .A(n3483), .B(n3460), .Z(n3474) );
  XOR U4805 ( .A(n3474), .B(n3461), .Z(n4037) );
  XNOR U4806 ( .A(n4039), .B(n4037), .Z(n3481) );
  AND U4807 ( .A(n3463), .B(n3462), .Z(n3470) );
  NANDN U4808 ( .A(n3465), .B(n3464), .Z(n3466) );
  XNOR U4809 ( .A(n3467), .B(n3466), .Z(n3473) );
  XNOR U4810 ( .A(n3473), .B(n3468), .Z(n3469) );
  XOR U4811 ( .A(n3470), .B(n3469), .Z(n4042) );
  XNOR U4812 ( .A(n3481), .B(n4042), .Z(z[102]) );
  ANDN U4813 ( .B(n3472), .A(n3471), .Z(n3476) );
  XOR U4814 ( .A(n3474), .B(n3473), .Z(n3475) );
  XNOR U4815 ( .A(n3476), .B(n3475), .Z(n3478) );
  XNOR U4816 ( .A(n3478), .B(n3477), .Z(n3479) );
  XNOR U4817 ( .A(n3480), .B(n3479), .Z(n4040) );
  XNOR U4818 ( .A(n4040), .B(n3481), .Z(z[97]) );
  XNOR U4819 ( .A(n3483), .B(n3482), .Z(n3484) );
  XNOR U4820 ( .A(n3485), .B(n3484), .Z(n3486) );
  XOR U4821 ( .A(n3486), .B(z[97]), .Z(z[103]) );
  NANDN U4822 ( .A(n3488), .B(n3487), .Z(n3489) );
  XNOR U4823 ( .A(n3490), .B(n3489), .Z(n3517) );
  XNOR U4824 ( .A(n3491), .B(n3517), .Z(n3492) );
  XOR U4825 ( .A(n3493), .B(n3492), .Z(n3505) );
  XOR U4826 ( .A(n3505), .B(n3494), .Z(z[104]) );
  ANDN U4827 ( .B(n3496), .A(n3495), .Z(n3501) );
  NANDN U4828 ( .A(n3498), .B(n3497), .Z(n3515) );
  XNOR U4829 ( .A(n3499), .B(n3515), .Z(n3500) );
  XOR U4830 ( .A(n3501), .B(n3500), .Z(n3520) );
  XOR U4831 ( .A(n3503), .B(n3502), .Z(n3504) );
  XOR U4832 ( .A(n3520), .B(n3504), .Z(z[107]) );
  XNOR U4833 ( .A(n3505), .B(z[106]), .Z(z[108]) );
  XNOR U4834 ( .A(n3507), .B(n3506), .Z(n3508) );
  XNOR U4835 ( .A(n3509), .B(n3508), .Z(n3519) );
  XNOR U4836 ( .A(n3511), .B(n3510), .Z(n3512) );
  NANDN U4837 ( .A(n3513), .B(n3512), .Z(n3514) );
  XOR U4838 ( .A(n3515), .B(n3514), .Z(n3516) );
  XNOR U4839 ( .A(n3517), .B(n3516), .Z(n3518) );
  XNOR U4840 ( .A(n3519), .B(n3518), .Z(z[109]) );
  XNOR U4841 ( .A(n3521), .B(n3520), .Z(z[110]) );
  NANDN U4842 ( .A(n3523), .B(n3522), .Z(n3524) );
  XNOR U4843 ( .A(n3525), .B(n3524), .Z(n3552) );
  XNOR U4844 ( .A(n3526), .B(n3552), .Z(n3527) );
  XOR U4845 ( .A(n3528), .B(n3527), .Z(n3540) );
  XOR U4846 ( .A(n3540), .B(n3529), .Z(z[112]) );
  ANDN U4847 ( .B(n3531), .A(n3530), .Z(n3536) );
  NANDN U4848 ( .A(n3533), .B(n3532), .Z(n3550) );
  XNOR U4849 ( .A(n3534), .B(n3550), .Z(n3535) );
  XOR U4850 ( .A(n3536), .B(n3535), .Z(n3555) );
  XOR U4851 ( .A(n3538), .B(n3537), .Z(n3539) );
  XOR U4852 ( .A(n3555), .B(n3539), .Z(z[115]) );
  XNOR U4853 ( .A(n3540), .B(z[114]), .Z(z[116]) );
  XNOR U4854 ( .A(n3542), .B(n3541), .Z(n3543) );
  XNOR U4855 ( .A(n3544), .B(n3543), .Z(n3554) );
  XNOR U4856 ( .A(n3546), .B(n3545), .Z(n3547) );
  NANDN U4857 ( .A(n3548), .B(n3547), .Z(n3549) );
  XOR U4858 ( .A(n3550), .B(n3549), .Z(n3551) );
  XNOR U4859 ( .A(n3552), .B(n3551), .Z(n3553) );
  XNOR U4860 ( .A(n3554), .B(n3553), .Z(z[117]) );
  XNOR U4861 ( .A(n3556), .B(n3555), .Z(z[118]) );
  NOR U4862 ( .A(n3558), .B(n3557), .Z(n3571) );
  XNOR U4863 ( .A(n3560), .B(n3559), .Z(n3637) );
  OR U4864 ( .A(n3561), .B(n3637), .Z(n3562) );
  XOR U4865 ( .A(n3571), .B(n3562), .Z(n3656) );
  XNOR U4866 ( .A(n3564), .B(n3563), .Z(n3623) );
  ANDN U4867 ( .B(n3565), .A(n3623), .Z(n3579) );
  NOR U4868 ( .A(n3566), .B(n3568), .Z(n3573) );
  NANDN U4869 ( .A(n3567), .B(n3581), .Z(n3649) );
  XOR U4870 ( .A(n3633), .B(n3568), .Z(n3647) );
  XNOR U4871 ( .A(n3581), .B(n3647), .Z(n3582) );
  OR U4872 ( .A(n3582), .B(n3569), .Z(n3570) );
  XNOR U4873 ( .A(n3649), .B(n3570), .Z(n3643) );
  XOR U4874 ( .A(n3571), .B(n3643), .Z(n3572) );
  XOR U4875 ( .A(n3573), .B(n3572), .Z(n3655) );
  XOR U4876 ( .A(n3575), .B(n3574), .Z(n3576) );
  NANDN U4877 ( .A(n3577), .B(n3576), .Z(n3635) );
  XNOR U4878 ( .A(n3655), .B(n3635), .Z(n3578) );
  XOR U4879 ( .A(n3579), .B(n3578), .Z(n3652) );
  XOR U4880 ( .A(n3656), .B(n3652), .Z(n3587) );
  NAND U4881 ( .A(n3581), .B(n3580), .Z(n3627) );
  OR U4882 ( .A(n3583), .B(n3582), .Z(n3584) );
  XNOR U4883 ( .A(n3627), .B(n3584), .Z(n3651) );
  XNOR U4884 ( .A(n3651), .B(n3585), .Z(n3586) );
  XOR U4885 ( .A(n3587), .B(n3586), .Z(z[11]) );
  NANDN U4886 ( .A(n3589), .B(n3588), .Z(n3590) );
  XNOR U4887 ( .A(n3591), .B(n3590), .Z(n3618) );
  XNOR U4888 ( .A(n3592), .B(n3618), .Z(n3593) );
  XOR U4889 ( .A(n3594), .B(n3593), .Z(n3606) );
  XOR U4890 ( .A(n3606), .B(n3595), .Z(z[120]) );
  ANDN U4891 ( .B(n3597), .A(n3596), .Z(n3602) );
  NANDN U4892 ( .A(n3599), .B(n3598), .Z(n3616) );
  XNOR U4893 ( .A(n3600), .B(n3616), .Z(n3601) );
  XOR U4894 ( .A(n3602), .B(n3601), .Z(n3621) );
  XOR U4895 ( .A(n3604), .B(n3603), .Z(n3605) );
  XOR U4896 ( .A(n3621), .B(n3605), .Z(z[123]) );
  XNOR U4897 ( .A(n3606), .B(z[122]), .Z(z[124]) );
  XNOR U4898 ( .A(n3608), .B(n3607), .Z(n3609) );
  XNOR U4899 ( .A(n3610), .B(n3609), .Z(n3620) );
  XNOR U4900 ( .A(n3612), .B(n3611), .Z(n3613) );
  NANDN U4901 ( .A(n3614), .B(n3613), .Z(n3615) );
  XOR U4902 ( .A(n3616), .B(n3615), .Z(n3617) );
  XNOR U4903 ( .A(n3618), .B(n3617), .Z(n3619) );
  XNOR U4904 ( .A(n3620), .B(n3619), .Z(z[125]) );
  XNOR U4905 ( .A(n3622), .B(n3621), .Z(z[126]) );
  ANDN U4906 ( .B(n3624), .A(n3623), .Z(n3630) );
  NAND U4907 ( .A(n3647), .B(n3625), .Z(n3626) );
  XNOR U4908 ( .A(n3627), .B(n3626), .Z(n3639) );
  XNOR U4909 ( .A(n3628), .B(n3639), .Z(n3629) );
  XOR U4910 ( .A(n3630), .B(n3629), .Z(n4008) );
  XNOR U4911 ( .A(n4008), .B(z[10]), .Z(z[12]) );
  XOR U4912 ( .A(x[9]), .B(n3631), .Z(n3632) );
  NANDN U4913 ( .A(n3633), .B(n3632), .Z(n3634) );
  XOR U4914 ( .A(n3635), .B(n3634), .Z(n3636) );
  XNOR U4915 ( .A(n4008), .B(n3636), .Z(n3645) );
  NOR U4916 ( .A(n3638), .B(n3637), .Z(n3642) );
  XOR U4917 ( .A(n3640), .B(n3639), .Z(n3641) );
  XOR U4918 ( .A(n3642), .B(n3641), .Z(n3657) );
  XNOR U4919 ( .A(n3643), .B(n3657), .Z(n3644) );
  XOR U4920 ( .A(n3645), .B(n3644), .Z(z[13]) );
  AND U4921 ( .A(n3647), .B(n3646), .Z(n3648) );
  XNOR U4922 ( .A(n3649), .B(n3648), .Z(n3654) );
  XNOR U4923 ( .A(n3651), .B(n3650), .Z(n4009) );
  XNOR U4924 ( .A(n3652), .B(n4009), .Z(n3653) );
  XOR U4925 ( .A(n3654), .B(n3653), .Z(z[14]) );
  XNOR U4926 ( .A(n3657), .B(z[9]), .Z(z[15]) );
  NANDN U4927 ( .A(n3659), .B(n3658), .Z(n3660) );
  XNOR U4928 ( .A(n3661), .B(n3660), .Z(n3688) );
  XNOR U4929 ( .A(n3662), .B(n3688), .Z(n3663) );
  XOR U4930 ( .A(n3664), .B(n3663), .Z(n3676) );
  XOR U4931 ( .A(n3676), .B(n3665), .Z(z[16]) );
  ANDN U4932 ( .B(n3667), .A(n3666), .Z(n3672) );
  NANDN U4933 ( .A(n3669), .B(n3668), .Z(n3686) );
  XNOR U4934 ( .A(n3670), .B(n3686), .Z(n3671) );
  XOR U4935 ( .A(n3672), .B(n3671), .Z(n3691) );
  XOR U4936 ( .A(n3674), .B(n3673), .Z(n3675) );
  XOR U4937 ( .A(n3691), .B(n3675), .Z(z[19]) );
  XNOR U4938 ( .A(n3676), .B(z[18]), .Z(z[20]) );
  XNOR U4939 ( .A(n3678), .B(n3677), .Z(n3679) );
  XNOR U4940 ( .A(n3680), .B(n3679), .Z(n3690) );
  XNOR U4941 ( .A(n3682), .B(n3681), .Z(n3683) );
  NANDN U4942 ( .A(n3684), .B(n3683), .Z(n3685) );
  XOR U4943 ( .A(n3686), .B(n3685), .Z(n3687) );
  XNOR U4944 ( .A(n3688), .B(n3687), .Z(n3689) );
  XNOR U4945 ( .A(n3690), .B(n3689), .Z(z[21]) );
  XNOR U4946 ( .A(n3692), .B(n3691), .Z(z[22]) );
  NANDN U4947 ( .A(n3694), .B(n3693), .Z(n3695) );
  XNOR U4948 ( .A(n3696), .B(n3695), .Z(n3723) );
  XNOR U4949 ( .A(n3697), .B(n3723), .Z(n3698) );
  XOR U4950 ( .A(n3699), .B(n3698), .Z(n3711) );
  XOR U4951 ( .A(n3711), .B(n3700), .Z(z[24]) );
  ANDN U4952 ( .B(n3702), .A(n3701), .Z(n3707) );
  NANDN U4953 ( .A(n3704), .B(n3703), .Z(n3721) );
  XNOR U4954 ( .A(n3705), .B(n3721), .Z(n3706) );
  XOR U4955 ( .A(n3707), .B(n3706), .Z(n3726) );
  XOR U4956 ( .A(n3709), .B(n3708), .Z(n3710) );
  XOR U4957 ( .A(n3726), .B(n3710), .Z(z[27]) );
  XNOR U4958 ( .A(n3711), .B(z[26]), .Z(z[28]) );
  XNOR U4959 ( .A(n3713), .B(n3712), .Z(n3714) );
  XNOR U4960 ( .A(n3715), .B(n3714), .Z(n3725) );
  XNOR U4961 ( .A(n3717), .B(n3716), .Z(n3718) );
  NANDN U4962 ( .A(n3719), .B(n3718), .Z(n3720) );
  XOR U4963 ( .A(n3721), .B(n3720), .Z(n3722) );
  XNOR U4964 ( .A(n3723), .B(n3722), .Z(n3724) );
  XNOR U4965 ( .A(n3725), .B(n3724), .Z(z[29]) );
  XNOR U4966 ( .A(n3727), .B(n3726), .Z(z[30]) );
  NANDN U4967 ( .A(n3729), .B(n3728), .Z(n3730) );
  XNOR U4968 ( .A(n3731), .B(n3730), .Z(n3758) );
  XNOR U4969 ( .A(n3732), .B(n3758), .Z(n3733) );
  XOR U4970 ( .A(n3734), .B(n3733), .Z(n3746) );
  XOR U4971 ( .A(n3746), .B(n3735), .Z(z[32]) );
  ANDN U4972 ( .B(n3737), .A(n3736), .Z(n3742) );
  NANDN U4973 ( .A(n3739), .B(n3738), .Z(n3756) );
  XNOR U4974 ( .A(n3740), .B(n3756), .Z(n3741) );
  XOR U4975 ( .A(n3742), .B(n3741), .Z(n3761) );
  XOR U4976 ( .A(n3744), .B(n3743), .Z(n3745) );
  XOR U4977 ( .A(n3761), .B(n3745), .Z(z[35]) );
  XNOR U4978 ( .A(n3746), .B(z[34]), .Z(z[36]) );
  XNOR U4979 ( .A(n3748), .B(n3747), .Z(n3749) );
  XNOR U4980 ( .A(n3750), .B(n3749), .Z(n3760) );
  XNOR U4981 ( .A(n3752), .B(n3751), .Z(n3753) );
  NANDN U4982 ( .A(n3754), .B(n3753), .Z(n3755) );
  XOR U4983 ( .A(n3756), .B(n3755), .Z(n3757) );
  XNOR U4984 ( .A(n3758), .B(n3757), .Z(n3759) );
  XNOR U4985 ( .A(n3760), .B(n3759), .Z(z[37]) );
  XNOR U4986 ( .A(n3762), .B(n3761), .Z(z[38]) );
  ANDN U4987 ( .B(n3764), .A(n3763), .Z(n3769) );
  NANDN U4988 ( .A(n3766), .B(n3765), .Z(n3871) );
  XNOR U4989 ( .A(n3767), .B(n3871), .Z(n3768) );
  XOR U4990 ( .A(n3769), .B(n3768), .Z(n3926) );
  XOR U4991 ( .A(n3771), .B(n3770), .Z(n3772) );
  XOR U4992 ( .A(n3926), .B(n3772), .Z(z[3]) );
  NANDN U4993 ( .A(n3774), .B(n3773), .Z(n3775) );
  XNOR U4994 ( .A(n3776), .B(n3775), .Z(n3803) );
  XNOR U4995 ( .A(n3777), .B(n3803), .Z(n3778) );
  XOR U4996 ( .A(n3779), .B(n3778), .Z(n3791) );
  XOR U4997 ( .A(n3791), .B(n3780), .Z(z[40]) );
  ANDN U4998 ( .B(n3782), .A(n3781), .Z(n3787) );
  NANDN U4999 ( .A(n3784), .B(n3783), .Z(n3801) );
  XNOR U5000 ( .A(n3785), .B(n3801), .Z(n3786) );
  XOR U5001 ( .A(n3787), .B(n3786), .Z(n3806) );
  XOR U5002 ( .A(n3789), .B(n3788), .Z(n3790) );
  XOR U5003 ( .A(n3806), .B(n3790), .Z(z[43]) );
  XNOR U5004 ( .A(n3791), .B(z[42]), .Z(z[44]) );
  XNOR U5005 ( .A(n3793), .B(n3792), .Z(n3794) );
  XNOR U5006 ( .A(n3795), .B(n3794), .Z(n3805) );
  XNOR U5007 ( .A(n3797), .B(n3796), .Z(n3798) );
  NANDN U5008 ( .A(n3799), .B(n3798), .Z(n3800) );
  XOR U5009 ( .A(n3801), .B(n3800), .Z(n3802) );
  XNOR U5010 ( .A(n3803), .B(n3802), .Z(n3804) );
  XNOR U5011 ( .A(n3805), .B(n3804), .Z(z[45]) );
  XNOR U5012 ( .A(n3807), .B(n3806), .Z(z[46]) );
  NANDN U5013 ( .A(n3809), .B(n3808), .Z(n3810) );
  XNOR U5014 ( .A(n3811), .B(n3810), .Z(n3839) );
  XNOR U5015 ( .A(n3812), .B(n3839), .Z(n3813) );
  XOR U5016 ( .A(n3814), .B(n3813), .Z(n3827) );
  XOR U5017 ( .A(n3827), .B(n3815), .Z(z[48]) );
  XNOR U5018 ( .A(n3816), .B(z[2]), .Z(z[4]) );
  ANDN U5019 ( .B(n3818), .A(n3817), .Z(n3823) );
  NANDN U5020 ( .A(n3820), .B(n3819), .Z(n3837) );
  XNOR U5021 ( .A(n3821), .B(n3837), .Z(n3822) );
  XOR U5022 ( .A(n3823), .B(n3822), .Z(n3842) );
  XOR U5023 ( .A(n3825), .B(n3824), .Z(n3826) );
  XOR U5024 ( .A(n3842), .B(n3826), .Z(z[51]) );
  XNOR U5025 ( .A(n3827), .B(z[50]), .Z(z[52]) );
  XNOR U5026 ( .A(n3829), .B(n3828), .Z(n3830) );
  XNOR U5027 ( .A(n3831), .B(n3830), .Z(n3841) );
  XNOR U5028 ( .A(n3833), .B(n3832), .Z(n3834) );
  NANDN U5029 ( .A(n3835), .B(n3834), .Z(n3836) );
  XOR U5030 ( .A(n3837), .B(n3836), .Z(n3838) );
  XNOR U5031 ( .A(n3839), .B(n3838), .Z(n3840) );
  XNOR U5032 ( .A(n3841), .B(n3840), .Z(z[53]) );
  XNOR U5033 ( .A(n3843), .B(n3842), .Z(z[54]) );
  NANDN U5034 ( .A(n3845), .B(n3844), .Z(n3846) );
  XNOR U5035 ( .A(n3847), .B(n3846), .Z(n3888) );
  XNOR U5036 ( .A(n3848), .B(n3888), .Z(n3849) );
  XOR U5037 ( .A(n3850), .B(n3849), .Z(n3876) );
  XOR U5038 ( .A(n3876), .B(n3851), .Z(z[56]) );
  ANDN U5039 ( .B(n3853), .A(n3852), .Z(n3858) );
  NANDN U5040 ( .A(n3855), .B(n3854), .Z(n3886) );
  XNOR U5041 ( .A(n3856), .B(n3886), .Z(n3857) );
  XOR U5042 ( .A(n3858), .B(n3857), .Z(n3891) );
  XOR U5043 ( .A(n3860), .B(n3859), .Z(n3861) );
  XOR U5044 ( .A(n3891), .B(n3861), .Z(z[59]) );
  XNOR U5045 ( .A(n3863), .B(n3862), .Z(n3864) );
  XNOR U5046 ( .A(n3865), .B(n3864), .Z(n3875) );
  XNOR U5047 ( .A(n3867), .B(n3866), .Z(n3868) );
  NANDN U5048 ( .A(n3869), .B(n3868), .Z(n3870) );
  XOR U5049 ( .A(n3871), .B(n3870), .Z(n3872) );
  XNOR U5050 ( .A(n3873), .B(n3872), .Z(n3874) );
  XNOR U5051 ( .A(n3875), .B(n3874), .Z(z[5]) );
  XNOR U5052 ( .A(n3876), .B(z[58]), .Z(z[60]) );
  XNOR U5053 ( .A(n3878), .B(n3877), .Z(n3879) );
  XNOR U5054 ( .A(n3880), .B(n3879), .Z(n3890) );
  XNOR U5055 ( .A(n3882), .B(n3881), .Z(n3883) );
  NANDN U5056 ( .A(n3884), .B(n3883), .Z(n3885) );
  XOR U5057 ( .A(n3886), .B(n3885), .Z(n3887) );
  XNOR U5058 ( .A(n3888), .B(n3887), .Z(n3889) );
  XNOR U5059 ( .A(n3890), .B(n3889), .Z(z[61]) );
  XNOR U5060 ( .A(n3892), .B(n3891), .Z(z[62]) );
  NANDN U5061 ( .A(n3894), .B(n3893), .Z(n3895) );
  XNOR U5062 ( .A(n3896), .B(n3895), .Z(n3923) );
  XNOR U5063 ( .A(n3897), .B(n3923), .Z(n3898) );
  XOR U5064 ( .A(n3899), .B(n3898), .Z(n3911) );
  XOR U5065 ( .A(n3911), .B(n3900), .Z(z[64]) );
  ANDN U5066 ( .B(n3902), .A(n3901), .Z(n3907) );
  NANDN U5067 ( .A(n3904), .B(n3903), .Z(n3921) );
  XNOR U5068 ( .A(n3905), .B(n3921), .Z(n3906) );
  XOR U5069 ( .A(n3907), .B(n3906), .Z(n3928) );
  XOR U5070 ( .A(n3909), .B(n3908), .Z(n3910) );
  XOR U5071 ( .A(n3928), .B(n3910), .Z(z[67]) );
  XNOR U5072 ( .A(n3911), .B(z[66]), .Z(z[68]) );
  XNOR U5073 ( .A(n3913), .B(n3912), .Z(n3914) );
  XNOR U5074 ( .A(n3915), .B(n3914), .Z(n3925) );
  XNOR U5075 ( .A(n3917), .B(n3916), .Z(n3918) );
  NANDN U5076 ( .A(n3919), .B(n3918), .Z(n3920) );
  XOR U5077 ( .A(n3921), .B(n3920), .Z(n3922) );
  XNOR U5078 ( .A(n3923), .B(n3922), .Z(n3924) );
  XNOR U5079 ( .A(n3925), .B(n3924), .Z(z[69]) );
  XNOR U5080 ( .A(n3927), .B(n3926), .Z(z[6]) );
  XNOR U5081 ( .A(n3929), .B(n3928), .Z(z[70]) );
  NANDN U5082 ( .A(n3931), .B(n3930), .Z(n3932) );
  XNOR U5083 ( .A(n3933), .B(n3932), .Z(n3960) );
  XNOR U5084 ( .A(n3934), .B(n3960), .Z(n3935) );
  XOR U5085 ( .A(n3936), .B(n3935), .Z(n3948) );
  XOR U5086 ( .A(n3948), .B(n3937), .Z(z[72]) );
  ANDN U5087 ( .B(n3939), .A(n3938), .Z(n3944) );
  NANDN U5088 ( .A(n3941), .B(n3940), .Z(n3958) );
  XNOR U5089 ( .A(n3942), .B(n3958), .Z(n3943) );
  XOR U5090 ( .A(n3944), .B(n3943), .Z(n3963) );
  XOR U5091 ( .A(n3946), .B(n3945), .Z(n3947) );
  XOR U5092 ( .A(n3963), .B(n3947), .Z(z[75]) );
  XNOR U5093 ( .A(n3948), .B(z[74]), .Z(z[76]) );
  XNOR U5094 ( .A(n3950), .B(n3949), .Z(n3951) );
  XNOR U5095 ( .A(n3952), .B(n3951), .Z(n3962) );
  XNOR U5096 ( .A(n3954), .B(n3953), .Z(n3955) );
  NANDN U5097 ( .A(n3956), .B(n3955), .Z(n3957) );
  XOR U5098 ( .A(n3958), .B(n3957), .Z(n3959) );
  XNOR U5099 ( .A(n3960), .B(n3959), .Z(n3961) );
  XNOR U5100 ( .A(n3962), .B(n3961), .Z(z[77]) );
  XNOR U5101 ( .A(n3964), .B(n3963), .Z(z[78]) );
  NANDN U5102 ( .A(n3966), .B(n3965), .Z(n3967) );
  XNOR U5103 ( .A(n3968), .B(n3967), .Z(n3995) );
  XNOR U5104 ( .A(n3969), .B(n3995), .Z(n3970) );
  XOR U5105 ( .A(n3971), .B(n3970), .Z(n3983) );
  XOR U5106 ( .A(n3983), .B(n3972), .Z(z[80]) );
  ANDN U5107 ( .B(n3974), .A(n3973), .Z(n3979) );
  NANDN U5108 ( .A(n3976), .B(n3975), .Z(n3993) );
  XNOR U5109 ( .A(n3977), .B(n3993), .Z(n3978) );
  XOR U5110 ( .A(n3979), .B(n3978), .Z(n3998) );
  XOR U5111 ( .A(n3981), .B(n3980), .Z(n3982) );
  XOR U5112 ( .A(n3998), .B(n3982), .Z(z[83]) );
  XNOR U5113 ( .A(n3983), .B(z[82]), .Z(z[84]) );
  XNOR U5114 ( .A(n3985), .B(n3984), .Z(n3986) );
  XNOR U5115 ( .A(n3987), .B(n3986), .Z(n3997) );
  XNOR U5116 ( .A(n3989), .B(n3988), .Z(n3990) );
  NANDN U5117 ( .A(n3991), .B(n3990), .Z(n3992) );
  XOR U5118 ( .A(n3993), .B(n3992), .Z(n3994) );
  XNOR U5119 ( .A(n3995), .B(n3994), .Z(n3996) );
  XNOR U5120 ( .A(n3997), .B(n3996), .Z(z[85]) );
  XNOR U5121 ( .A(n3999), .B(n3998), .Z(z[86]) );
  NANDN U5122 ( .A(n4001), .B(n4000), .Z(n4002) );
  XNOR U5123 ( .A(n4003), .B(n4002), .Z(n4032) );
  XNOR U5124 ( .A(n4004), .B(n4032), .Z(n4005) );
  XOR U5125 ( .A(n4006), .B(n4005), .Z(n4020) );
  XOR U5126 ( .A(n4020), .B(n4007), .Z(z[88]) );
  XNOR U5127 ( .A(n4009), .B(n4008), .Z(z[8]) );
  ANDN U5128 ( .B(n4011), .A(n4010), .Z(n4016) );
  NANDN U5129 ( .A(n4013), .B(n4012), .Z(n4030) );
  XNOR U5130 ( .A(n4014), .B(n4030), .Z(n4015) );
  XOR U5131 ( .A(n4016), .B(n4015), .Z(n4035) );
  XOR U5132 ( .A(n4018), .B(n4017), .Z(n4019) );
  XOR U5133 ( .A(n4035), .B(n4019), .Z(z[91]) );
  XNOR U5134 ( .A(n4020), .B(z[90]), .Z(z[92]) );
  XNOR U5135 ( .A(n4022), .B(n4021), .Z(n4023) );
  XNOR U5136 ( .A(n4024), .B(n4023), .Z(n4034) );
  XNOR U5137 ( .A(n4026), .B(n4025), .Z(n4027) );
  NANDN U5138 ( .A(n4028), .B(n4027), .Z(n4029) );
  XOR U5139 ( .A(n4030), .B(n4029), .Z(n4031) );
  XNOR U5140 ( .A(n4032), .B(n4031), .Z(n4033) );
  XNOR U5141 ( .A(n4034), .B(n4033), .Z(z[93]) );
  XNOR U5142 ( .A(n4036), .B(n4035), .Z(z[94]) );
  XNOR U5143 ( .A(n4038), .B(n4037), .Z(z[96]) );
  XOR U5144 ( .A(n4040), .B(n4039), .Z(n4041) );
  XOR U5145 ( .A(n4042), .B(n4041), .Z(z[99]) );
endmodule


module aes_seq_CC5 ( clk, rst, msg, key, out );
  input [127:0] msg;
  input [255:0] key;
  output [127:0] out;
  input clk, rst;
  wire   init, \w0[1][127] , \w0[1][126] , \w0[1][125] , \w0[1][124] ,
         \w0[1][123] , \w0[1][122] , \w0[1][121] , \w0[1][120] , \w0[1][119] ,
         \w0[1][118] , \w0[1][117] , \w0[1][116] , \w0[1][115] , \w0[1][114] ,
         \w0[1][113] , \w0[1][112] , \w0[1][111] , \w0[1][110] , \w0[1][109] ,
         \w0[1][108] , \w0[1][107] , \w0[1][106] , \w0[1][105] , \w0[1][104] ,
         \w0[1][103] , \w0[1][102] , \w0[1][101] , \w0[1][100] , \w0[1][99] ,
         \w0[1][98] , \w0[1][97] , \w0[1][96] , \w0[1][95] , \w0[1][94] ,
         \w0[1][93] , \w0[1][92] , \w0[1][91] , \w0[1][90] , \w0[1][89] ,
         \w0[1][88] , \w0[1][87] , \w0[1][86] , \w0[1][85] , \w0[1][84] ,
         \w0[1][83] , \w0[1][82] , \w0[1][81] , \w0[1][80] , \w0[1][79] ,
         \w0[1][78] , \w0[1][77] , \w0[1][76] , \w0[1][75] , \w0[1][74] ,
         \w0[1][73] , \w0[1][72] , \w0[1][71] , \w0[1][70] , \w0[1][69] ,
         \w0[1][68] , \w0[1][67] , \w0[1][66] , \w0[1][65] , \w0[1][64] ,
         \w0[1][63] , \w0[1][62] , \w0[1][61] , \w0[1][60] , \w0[1][59] ,
         \w0[1][58] , \w0[1][57] , \w0[1][56] , \w0[1][55] , \w0[1][54] ,
         \w0[1][53] , \w0[1][52] , \w0[1][51] , \w0[1][50] , \w0[1][49] ,
         \w0[1][48] , \w0[1][47] , \w0[1][46] , \w0[1][45] , \w0[1][44] ,
         \w0[1][43] , \w0[1][42] , \w0[1][41] , \w0[1][40] , \w0[1][39] ,
         \w0[1][38] , \w0[1][37] , \w0[1][36] , \w0[1][35] , \w0[1][34] ,
         \w0[1][33] , \w0[1][32] , \w0[1][31] , \w0[1][30] , \w0[1][29] ,
         \w0[1][28] , \w0[1][27] , \w0[1][26] , \w0[1][25] , \w0[1][24] ,
         \w0[1][23] , \w0[1][22] , \w0[1][21] , \w0[1][20] , \w0[1][19] ,
         \w0[1][18] , \w0[1][17] , \w0[1][16] , \w0[1][15] , \w0[1][14] ,
         \w0[1][13] , \w0[1][12] , \w0[1][11] , \w0[1][10] , \w0[1][9] ,
         \w0[1][8] , \w0[1][7] , \w0[1][6] , \w0[1][5] , \w0[1][4] ,
         \w0[1][3] , \w0[1][2] , \w0[1][1] , \w0[1][0] , \w1[1][127] ,
         \w1[1][126] , \w1[1][125] , \w1[1][124] , \w1[1][123] , \w1[1][122] ,
         \w1[1][121] , \w1[1][120] , \w1[1][119] , \w1[1][118] , \w1[1][117] ,
         \w1[1][116] , \w1[1][115] , \w1[1][114] , \w1[1][113] , \w1[1][112] ,
         \w1[1][111] , \w1[1][110] , \w1[1][109] , \w1[1][108] , \w1[1][107] ,
         \w1[1][106] , \w1[1][105] , \w1[1][104] , \w1[1][103] , \w1[1][102] ,
         \w1[1][101] , \w1[1][100] , \w1[1][99] , \w1[1][98] , \w1[1][97] ,
         \w1[1][96] , \w1[1][95] , \w1[1][94] , \w1[1][93] , \w1[1][92] ,
         \w1[1][91] , \w1[1][90] , \w1[1][89] , \w1[1][88] , \w1[1][87] ,
         \w1[1][86] , \w1[1][85] , \w1[1][84] , \w1[1][83] , \w1[1][82] ,
         \w1[1][81] , \w1[1][80] , \w1[1][79] , \w1[1][78] , \w1[1][77] ,
         \w1[1][76] , \w1[1][75] , \w1[1][74] , \w1[1][73] , \w1[1][72] ,
         \w1[1][71] , \w1[1][70] , \w1[1][69] , \w1[1][68] , \w1[1][67] ,
         \w1[1][66] , \w1[1][65] , \w1[1][64] , \w1[1][63] , \w1[1][62] ,
         \w1[1][61] , \w1[1][60] , \w1[1][59] , \w1[1][58] , \w1[1][57] ,
         \w1[1][56] , \w1[1][55] , \w1[1][54] , \w1[1][53] , \w1[1][52] ,
         \w1[1][51] , \w1[1][50] , \w1[1][49] , \w1[1][48] , \w1[1][47] ,
         \w1[1][46] , \w1[1][45] , \w1[1][44] , \w1[1][43] , \w1[1][42] ,
         \w1[1][41] , \w1[1][40] , \w1[1][39] , \w1[1][38] , \w1[1][37] ,
         \w1[1][36] , \w1[1][35] , \w1[1][34] , \w1[1][33] , \w1[1][32] ,
         \w1[1][31] , \w1[1][30] , \w1[1][29] , \w1[1][28] , \w1[1][27] ,
         \w1[1][26] , \w1[1][25] , \w1[1][24] , \w1[1][23] , \w1[1][22] ,
         \w1[1][21] , \w1[1][20] , \w1[1][19] , \w1[1][18] , \w1[1][17] ,
         \w1[1][16] , \w1[1][15] , \w1[1][14] , \w1[1][13] , \w1[1][12] ,
         \w1[1][11] , \w1[1][10] , \w1[1][9] , \w1[1][8] , \w1[1][7] ,
         \w1[1][6] , \w1[1][5] , \w1[1][4] , \w1[1][3] , \w1[1][2] ,
         \w1[1][1] , \w1[1][0] , \w1[0][127] , \w1[0][126] , \w1[0][125] ,
         \w1[0][124] , \w1[0][123] , \w1[0][122] , \w1[0][121] , \w1[0][120] ,
         \w1[0][119] , \w1[0][118] , \w1[0][117] , \w1[0][116] , \w1[0][115] ,
         \w1[0][114] , \w1[0][113] , \w1[0][112] , \w1[0][111] , \w1[0][110] ,
         \w1[0][109] , \w1[0][108] , \w1[0][107] , \w1[0][106] , \w1[0][105] ,
         \w1[0][104] , \w1[0][103] , \w1[0][102] , \w1[0][101] , \w1[0][100] ,
         \w1[0][99] , \w1[0][98] , \w1[0][97] , \w1[0][96] , \w1[0][95] ,
         \w1[0][94] , \w1[0][93] , \w1[0][92] , \w1[0][91] , \w1[0][90] ,
         \w1[0][89] , \w1[0][88] , \w1[0][87] , \w1[0][86] , \w1[0][85] ,
         \w1[0][84] , \w1[0][83] , \w1[0][82] , \w1[0][81] , \w1[0][80] ,
         \w1[0][79] , \w1[0][78] , \w1[0][77] , \w1[0][76] , \w1[0][75] ,
         \w1[0][74] , \w1[0][73] , \w1[0][72] , \w1[0][71] , \w1[0][70] ,
         \w1[0][69] , \w1[0][68] , \w1[0][67] , \w1[0][66] , \w1[0][65] ,
         \w1[0][64] , \w1[0][63] , \w1[0][62] , \w1[0][61] , \w1[0][60] ,
         \w1[0][59] , \w1[0][58] , \w1[0][57] , \w1[0][56] , \w1[0][55] ,
         \w1[0][54] , \w1[0][53] , \w1[0][52] , \w1[0][51] , \w1[0][50] ,
         \w1[0][49] , \w1[0][48] , \w1[0][47] , \w1[0][46] , \w1[0][45] ,
         \w1[0][44] , \w1[0][43] , \w1[0][42] , \w1[0][41] , \w1[0][40] ,
         \w1[0][39] , \w1[0][38] , \w1[0][37] , \w1[0][36] , \w1[0][35] ,
         \w1[0][34] , \w1[0][33] , \w1[0][32] , \w1[0][31] , \w1[0][30] ,
         \w1[0][29] , \w1[0][28] , \w1[0][27] , \w1[0][26] , \w1[0][25] ,
         \w1[0][24] , \w1[0][23] , \w1[0][22] , \w1[0][21] , \w1[0][20] ,
         \w1[0][19] , \w1[0][18] , \w1[0][17] , \w1[0][16] , \w1[0][15] ,
         \w1[0][14] , \w1[0][13] , \w1[0][12] , \w1[0][11] , \w1[0][10] ,
         \w1[0][9] , \w1[0][8] , \w1[0][7] , \w1[0][6] , \w1[0][5] ,
         \w1[0][4] , \w1[0][3] , \w1[0][2] , \w1[0][1] , \w1[0][0] ,
         \w3[1][127] , \w3[1][126] , \w3[1][125] , \w3[1][124] , \w3[1][123] ,
         \w3[1][122] , \w3[1][121] , \w3[1][120] , \w3[1][119] , \w3[1][118] ,
         \w3[1][117] , \w3[1][116] , \w3[1][115] , \w3[1][114] , \w3[1][113] ,
         \w3[1][112] , \w3[1][111] , \w3[1][110] , \w3[1][109] , \w3[1][108] ,
         \w3[1][107] , \w3[1][106] , \w3[1][105] , \w3[1][104] , \w3[1][103] ,
         \w3[1][102] , \w3[1][101] , \w3[1][100] , \w3[1][99] , \w3[1][98] ,
         \w3[1][97] , \w3[1][96] , \w3[1][95] , \w3[1][94] , \w3[1][93] ,
         \w3[1][92] , \w3[1][91] , \w3[1][90] , \w3[1][89] , \w3[1][88] ,
         \w3[1][87] , \w3[1][86] , \w3[1][85] , \w3[1][84] , \w3[1][83] ,
         \w3[1][82] , \w3[1][81] , \w3[1][80] , \w3[1][79] , \w3[1][78] ,
         \w3[1][77] , \w3[1][76] , \w3[1][75] , \w3[1][74] , \w3[1][73] ,
         \w3[1][72] , \w3[1][71] , \w3[1][70] , \w3[1][69] , \w3[1][68] ,
         \w3[1][67] , \w3[1][66] , \w3[1][65] , \w3[1][64] , \w3[1][63] ,
         \w3[1][62] , \w3[1][61] , \w3[1][60] , \w3[1][59] , \w3[1][58] ,
         \w3[1][57] , \w3[1][56] , \w3[1][55] , \w3[1][54] , \w3[1][53] ,
         \w3[1][52] , \w3[1][51] , \w3[1][50] , \w3[1][49] , \w3[1][48] ,
         \w3[1][47] , \w3[1][46] , \w3[1][45] , \w3[1][44] , \w3[1][43] ,
         \w3[1][42] , \w3[1][41] , \w3[1][40] , \w3[1][39] , \w3[1][38] ,
         \w3[1][37] , \w3[1][36] , \w3[1][35] , \w3[1][34] , \w3[1][33] ,
         \w3[1][32] , \w3[1][31] , \w3[1][30] , \w3[1][29] , \w3[1][28] ,
         \w3[1][27] , \w3[1][26] , \w3[1][25] , \w3[1][24] , \w3[1][23] ,
         \w3[1][22] , \w3[1][21] , \w3[1][20] , \w3[1][19] , \w3[1][18] ,
         \w3[1][17] , \w3[1][16] , \w3[1][15] , \w3[1][14] , \w3[1][13] ,
         \w3[1][12] , \w3[1][11] , \w3[1][10] , \w3[1][9] , \w3[1][8] ,
         \w3[1][7] , \w3[1][6] , \w3[1][5] , \w3[1][4] , \w3[1][3] ,
         \w3[1][2] , \w3[1][1] , \w3[1][0] , \w3[0][127] , \w3[0][126] ,
         \w3[0][125] , \w3[0][124] , \w3[0][123] , \w3[0][122] , \w3[0][121] ,
         \w3[0][120] , \w3[0][119] , \w3[0][118] , \w3[0][117] , \w3[0][116] ,
         \w3[0][115] , \w3[0][114] , \w3[0][113] , \w3[0][112] , \w3[0][111] ,
         \w3[0][110] , \w3[0][109] , \w3[0][108] , \w3[0][107] , \w3[0][106] ,
         \w3[0][105] , \w3[0][104] , \w3[0][103] , \w3[0][102] , \w3[0][101] ,
         \w3[0][100] , \w3[0][99] , \w3[0][98] , \w3[0][97] , \w3[0][96] ,
         \w3[0][95] , \w3[0][94] , \w3[0][93] , \w3[0][92] , \w3[0][91] ,
         \w3[0][90] , \w3[0][89] , \w3[0][88] , \w3[0][87] , \w3[0][86] ,
         \w3[0][85] , \w3[0][84] , \w3[0][83] , \w3[0][82] , \w3[0][81] ,
         \w3[0][80] , \w3[0][79] , \w3[0][78] , \w3[0][77] , \w3[0][76] ,
         \w3[0][75] , \w3[0][74] , \w3[0][73] , \w3[0][72] , \w3[0][71] ,
         \w3[0][70] , \w3[0][69] , \w3[0][68] , \w3[0][67] , \w3[0][66] ,
         \w3[0][65] , \w3[0][64] , \w3[0][63] , \w3[0][62] , \w3[0][61] ,
         \w3[0][60] , \w3[0][59] , \w3[0][58] , \w3[0][57] , \w3[0][56] ,
         \w3[0][55] , \w3[0][54] , \w3[0][53] , \w3[0][52] , \w3[0][51] ,
         \w3[0][50] , \w3[0][49] , \w3[0][48] , \w3[0][47] , \w3[0][46] ,
         \w3[0][45] , \w3[0][44] , \w3[0][43] , \w3[0][42] , \w3[0][41] ,
         \w3[0][40] , \w3[0][39] , \w3[0][38] , \w3[0][37] , \w3[0][36] ,
         \w3[0][35] , \w3[0][34] , \w3[0][33] , \w3[0][32] , \w3[0][31] ,
         \w3[0][30] , \w3[0][29] , \w3[0][28] , \w3[0][27] , \w3[0][26] ,
         \w3[0][25] , \w3[0][24] , \w3[0][23] , \w3[0][22] , \w3[0][21] ,
         \w3[0][20] , \w3[0][19] , \w3[0][18] , \w3[0][17] , \w3[0][16] ,
         \w3[0][15] , \w3[0][14] , \w3[0][13] , \w3[0][12] , \w3[0][11] ,
         \w3[0][10] , \w3[0][9] , \w3[0][8] , \w3[0][7] , \w3[0][6] ,
         \w3[0][5] , \w3[0][4] , \w3[0][3] , \w3[0][2] , \w3[0][1] ,
         \w3[0][0] , n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396;
  wire   [127:0] state;

  SubBytes_0 \SUBBYTES[0].a  ( .x({\w1[0][127] , \w1[0][126] , \w1[0][125] , 
        \w1[0][124] , \w1[0][123] , \w1[0][122] , \w1[0][121] , \w1[0][120] , 
        \w1[0][119] , \w1[0][118] , \w1[0][117] , \w1[0][116] , \w1[0][115] , 
        \w1[0][114] , \w1[0][113] , \w1[0][112] , \w1[0][111] , \w1[0][110] , 
        \w1[0][109] , \w1[0][108] , \w1[0][107] , \w1[0][106] , \w1[0][105] , 
        \w1[0][104] , \w1[0][103] , \w1[0][102] , \w1[0][101] , \w1[0][100] , 
        \w1[0][99] , \w1[0][98] , \w1[0][97] , \w1[0][96] , \w1[0][95] , 
        \w1[0][94] , \w1[0][93] , \w1[0][92] , \w1[0][91] , \w1[0][90] , 
        \w1[0][89] , \w1[0][88] , \w1[0][87] , \w1[0][86] , \w1[0][85] , 
        \w1[0][84] , \w1[0][83] , \w1[0][82] , \w1[0][81] , \w1[0][80] , 
        \w1[0][79] , \w1[0][78] , \w1[0][77] , \w1[0][76] , \w1[0][75] , 
        \w1[0][74] , \w1[0][73] , \w1[0][72] , \w1[0][71] , \w1[0][70] , 
        \w1[0][69] , \w1[0][68] , \w1[0][67] , \w1[0][66] , \w1[0][65] , 
        \w1[0][64] , \w1[0][63] , \w1[0][62] , \w1[0][61] , \w1[0][60] , 
        \w1[0][59] , \w1[0][58] , \w1[0][57] , \w1[0][56] , \w1[0][55] , 
        \w1[0][54] , \w1[0][53] , \w1[0][52] , \w1[0][51] , \w1[0][50] , 
        \w1[0][49] , \w1[0][48] , \w1[0][47] , \w1[0][46] , \w1[0][45] , 
        \w1[0][44] , \w1[0][43] , \w1[0][42] , \w1[0][41] , \w1[0][40] , 
        \w1[0][39] , \w1[0][38] , \w1[0][37] , \w1[0][36] , \w1[0][35] , 
        \w1[0][34] , \w1[0][33] , \w1[0][32] , \w1[0][31] , \w1[0][30] , 
        \w1[0][29] , \w1[0][28] , \w1[0][27] , \w1[0][26] , \w1[0][25] , 
        \w1[0][24] , \w1[0][23] , \w1[0][22] , \w1[0][21] , \w1[0][20] , 
        \w1[0][19] , \w1[0][18] , \w1[0][17] , \w1[0][16] , \w1[0][15] , 
        \w1[0][14] , \w1[0][13] , \w1[0][12] , \w1[0][11] , \w1[0][10] , 
        \w1[0][9] , \w1[0][8] , \w1[0][7] , \w1[0][6] , \w1[0][5] , \w1[0][4] , 
        \w1[0][3] , \w1[0][2] , \w1[0][1] , \w1[0][0] }), .z({\w3[0][127] , 
        \w3[0][126] , \w3[0][125] , \w3[0][124] , \w3[0][123] , \w3[0][122] , 
        \w3[0][121] , \w3[0][120] , \w3[0][23] , \w3[0][22] , \w3[0][21] , 
        \w3[0][20] , \w3[0][19] , \w3[0][18] , \w3[0][17] , \w3[0][16] , 
        \w3[0][47] , \w3[0][46] , \w3[0][45] , \w3[0][44] , \w3[0][43] , 
        \w3[0][42] , \w3[0][41] , \w3[0][40] , \w3[0][71] , \w3[0][70] , 
        \w3[0][69] , \w3[0][68] , \w3[0][67] , \w3[0][66] , \w3[0][65] , 
        \w3[0][64] , \w3[0][95] , \w3[0][94] , \w3[0][93] , \w3[0][92] , 
        \w3[0][91] , \w3[0][90] , \w3[0][89] , \w3[0][88] , \w3[0][119] , 
        \w3[0][118] , \w3[0][117] , \w3[0][116] , \w3[0][115] , \w3[0][114] , 
        \w3[0][113] , \w3[0][112] , \w3[0][15] , \w3[0][14] , \w3[0][13] , 
        \w3[0][12] , \w3[0][11] , \w3[0][10] , \w3[0][9] , \w3[0][8] , 
        \w3[0][39] , \w3[0][38] , \w3[0][37] , \w3[0][36] , \w3[0][35] , 
        \w3[0][34] , \w3[0][33] , \w3[0][32] , \w3[0][63] , \w3[0][62] , 
        \w3[0][61] , \w3[0][60] , \w3[0][59] , \w3[0][58] , \w3[0][57] , 
        \w3[0][56] , \w3[0][87] , \w3[0][86] , \w3[0][85] , \w3[0][84] , 
        \w3[0][83] , \w3[0][82] , \w3[0][81] , \w3[0][80] , \w3[0][111] , 
        \w3[0][110] , \w3[0][109] , \w3[0][108] , \w3[0][107] , \w3[0][106] , 
        \w3[0][105] , \w3[0][104] , \w3[0][7] , \w3[0][6] , \w3[0][5] , 
        \w3[0][4] , \w3[0][3] , \w3[0][2] , \w3[0][1] , \w3[0][0] , 
        \w3[0][31] , \w3[0][30] , \w3[0][29] , \w3[0][28] , \w3[0][27] , 
        \w3[0][26] , \w3[0][25] , \w3[0][24] , \w3[0][55] , \w3[0][54] , 
        \w3[0][53] , \w3[0][52] , \w3[0][51] , \w3[0][50] , \w3[0][49] , 
        \w3[0][48] , \w3[0][79] , \w3[0][78] , \w3[0][77] , \w3[0][76] , 
        \w3[0][75] , \w3[0][74] , \w3[0][73] , \w3[0][72] , \w3[0][103] , 
        \w3[0][102] , \w3[0][101] , \w3[0][100] , \w3[0][99] , \w3[0][98] , 
        \w3[0][97] , \w3[0][96] }) );
  SubBytes_1 \SUBBYTES[1].a  ( .x({\w1[1][127] , \w1[1][126] , \w1[1][125] , 
        \w1[1][124] , \w1[1][123] , \w1[1][122] , \w1[1][121] , \w1[1][120] , 
        \w1[1][119] , \w1[1][118] , \w1[1][117] , \w1[1][116] , \w1[1][115] , 
        \w1[1][114] , \w1[1][113] , \w1[1][112] , \w1[1][111] , \w1[1][110] , 
        \w1[1][109] , \w1[1][108] , \w1[1][107] , \w1[1][106] , \w1[1][105] , 
        \w1[1][104] , \w1[1][103] , \w1[1][102] , \w1[1][101] , \w1[1][100] , 
        \w1[1][99] , \w1[1][98] , \w1[1][97] , \w1[1][96] , \w1[1][95] , 
        \w1[1][94] , \w1[1][93] , \w1[1][92] , \w1[1][91] , \w1[1][90] , 
        \w1[1][89] , \w1[1][88] , \w1[1][87] , \w1[1][86] , \w1[1][85] , 
        \w1[1][84] , \w1[1][83] , \w1[1][82] , \w1[1][81] , \w1[1][80] , 
        \w1[1][79] , \w1[1][78] , \w1[1][77] , \w1[1][76] , \w1[1][75] , 
        \w1[1][74] , \w1[1][73] , \w1[1][72] , \w1[1][71] , \w1[1][70] , 
        \w1[1][69] , \w1[1][68] , \w1[1][67] , \w1[1][66] , \w1[1][65] , 
        \w1[1][64] , \w1[1][63] , \w1[1][62] , \w1[1][61] , \w1[1][60] , 
        \w1[1][59] , \w1[1][58] , \w1[1][57] , \w1[1][56] , \w1[1][55] , 
        \w1[1][54] , \w1[1][53] , \w1[1][52] , \w1[1][51] , \w1[1][50] , 
        \w1[1][49] , \w1[1][48] , \w1[1][47] , \w1[1][46] , \w1[1][45] , 
        \w1[1][44] , \w1[1][43] , \w1[1][42] , \w1[1][41] , \w1[1][40] , 
        \w1[1][39] , \w1[1][38] , \w1[1][37] , \w1[1][36] , \w1[1][35] , 
        \w1[1][34] , \w1[1][33] , \w1[1][32] , \w1[1][31] , \w1[1][30] , 
        \w1[1][29] , \w1[1][28] , \w1[1][27] , \w1[1][26] , \w1[1][25] , 
        \w1[1][24] , \w1[1][23] , \w1[1][22] , \w1[1][21] , \w1[1][20] , 
        \w1[1][19] , \w1[1][18] , \w1[1][17] , \w1[1][16] , \w1[1][15] , 
        \w1[1][14] , \w1[1][13] , \w1[1][12] , \w1[1][11] , \w1[1][10] , 
        \w1[1][9] , \w1[1][8] , \w1[1][7] , \w1[1][6] , \w1[1][5] , \w1[1][4] , 
        \w1[1][3] , \w1[1][2] , \w1[1][1] , \w1[1][0] }), .z({\w3[1][127] , 
        \w3[1][126] , \w3[1][125] , \w3[1][124] , \w3[1][123] , \w3[1][122] , 
        \w3[1][121] , \w3[1][120] , \w3[1][23] , \w3[1][22] , \w3[1][21] , 
        \w3[1][20] , \w3[1][19] , \w3[1][18] , \w3[1][17] , \w3[1][16] , 
        \w3[1][47] , \w3[1][46] , \w3[1][45] , \w3[1][44] , \w3[1][43] , 
        \w3[1][42] , \w3[1][41] , \w3[1][40] , \w3[1][71] , \w3[1][70] , 
        \w3[1][69] , \w3[1][68] , \w3[1][67] , \w3[1][66] , \w3[1][65] , 
        \w3[1][64] , \w3[1][95] , \w3[1][94] , \w3[1][93] , \w3[1][92] , 
        \w3[1][91] , \w3[1][90] , \w3[1][89] , \w3[1][88] , \w3[1][119] , 
        \w3[1][118] , \w3[1][117] , \w3[1][116] , \w3[1][115] , \w3[1][114] , 
        \w3[1][113] , \w3[1][112] , \w3[1][15] , \w3[1][14] , \w3[1][13] , 
        \w3[1][12] , \w3[1][11] , \w3[1][10] , \w3[1][9] , \w3[1][8] , 
        \w3[1][39] , \w3[1][38] , \w3[1][37] , \w3[1][36] , \w3[1][35] , 
        \w3[1][34] , \w3[1][33] , \w3[1][32] , \w3[1][63] , \w3[1][62] , 
        \w3[1][61] , \w3[1][60] , \w3[1][59] , \w3[1][58] , \w3[1][57] , 
        \w3[1][56] , \w3[1][87] , \w3[1][86] , \w3[1][85] , \w3[1][84] , 
        \w3[1][83] , \w3[1][82] , \w3[1][81] , \w3[1][80] , \w3[1][111] , 
        \w3[1][110] , \w3[1][109] , \w3[1][108] , \w3[1][107] , \w3[1][106] , 
        \w3[1][105] , \w3[1][104] , \w3[1][7] , \w3[1][6] , \w3[1][5] , 
        \w3[1][4] , \w3[1][3] , \w3[1][2] , \w3[1][1] , \w3[1][0] , 
        \w3[1][31] , \w3[1][30] , \w3[1][29] , \w3[1][28] , \w3[1][27] , 
        \w3[1][26] , \w3[1][25] , \w3[1][24] , \w3[1][55] , \w3[1][54] , 
        \w3[1][53] , \w3[1][52] , \w3[1][51] , \w3[1][50] , \w3[1][49] , 
        \w3[1][48] , \w3[1][79] , \w3[1][78] , \w3[1][77] , \w3[1][76] , 
        \w3[1][75] , \w3[1][74] , \w3[1][73] , \w3[1][72] , \w3[1][103] , 
        \w3[1][102] , \w3[1][101] , \w3[1][100] , \w3[1][99] , \w3[1][98] , 
        \w3[1][97] , \w3[1][96] }) );
  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \state_reg[0]  ( .D(\w0[1][0] ), .CLK(clk), .RST(rst), .Q(state[0]) );
  DFF \state_reg[71]  ( .D(\w0[1][71] ), .CLK(clk), .RST(rst), .Q(state[71])
         );
  DFF \state_reg[88]  ( .D(\w0[1][88] ), .CLK(clk), .RST(rst), .Q(state[88])
         );
  DFF \state_reg[80]  ( .D(\w0[1][80] ), .CLK(clk), .RST(rst), .Q(state[80])
         );
  DFF \state_reg[81]  ( .D(\w0[1][81] ), .CLK(clk), .RST(rst), .Q(state[81])
         );
  DFF \state_reg[64]  ( .D(\w0[1][64] ), .CLK(clk), .RST(rst), .Q(state[64])
         );
  DFF \state_reg[72]  ( .D(\w0[1][72] ), .CLK(clk), .RST(rst), .Q(state[72])
         );
  DFF \state_reg[89]  ( .D(\w0[1][89] ), .CLK(clk), .RST(rst), .Q(state[89])
         );
  DFF \state_reg[82]  ( .D(\w0[1][82] ), .CLK(clk), .RST(rst), .Q(state[82])
         );
  DFF \state_reg[65]  ( .D(\w0[1][65] ), .CLK(clk), .RST(rst), .Q(state[65])
         );
  DFF \state_reg[73]  ( .D(\w0[1][73] ), .CLK(clk), .RST(rst), .Q(state[73])
         );
  DFF \state_reg[90]  ( .D(\w0[1][90] ), .CLK(clk), .RST(rst), .Q(state[90])
         );
  DFF \state_reg[83]  ( .D(\w0[1][83] ), .CLK(clk), .RST(rst), .Q(state[83])
         );
  DFF \state_reg[66]  ( .D(\w0[1][66] ), .CLK(clk), .RST(rst), .Q(state[66])
         );
  DFF \state_reg[74]  ( .D(\w0[1][74] ), .CLK(clk), .RST(rst), .Q(state[74])
         );
  DFF \state_reg[91]  ( .D(\w0[1][91] ), .CLK(clk), .RST(rst), .Q(state[91])
         );
  DFF \state_reg[75]  ( .D(\w0[1][75] ), .CLK(clk), .RST(rst), .Q(state[75])
         );
  DFF \state_reg[67]  ( .D(\w0[1][67] ), .CLK(clk), .RST(rst), .Q(state[67])
         );
  DFF \state_reg[84]  ( .D(\w0[1][84] ), .CLK(clk), .RST(rst), .Q(state[84])
         );
  DFF \state_reg[92]  ( .D(\w0[1][92] ), .CLK(clk), .RST(rst), .Q(state[92])
         );
  DFF \state_reg[76]  ( .D(\w0[1][76] ), .CLK(clk), .RST(rst), .Q(state[76])
         );
  DFF \state_reg[68]  ( .D(\w0[1][68] ), .CLK(clk), .RST(rst), .Q(state[68])
         );
  DFF \state_reg[85]  ( .D(\w0[1][85] ), .CLK(clk), .RST(rst), .Q(state[85])
         );
  DFF \state_reg[93]  ( .D(\w0[1][93] ), .CLK(clk), .RST(rst), .Q(state[93])
         );
  DFF \state_reg[86]  ( .D(\w0[1][86] ), .CLK(clk), .RST(rst), .Q(state[86])
         );
  DFF \state_reg[69]  ( .D(\w0[1][69] ), .CLK(clk), .RST(rst), .Q(state[69])
         );
  DFF \state_reg[77]  ( .D(\w0[1][77] ), .CLK(clk), .RST(rst), .Q(state[77])
         );
  DFF \state_reg[94]  ( .D(\w0[1][94] ), .CLK(clk), .RST(rst), .Q(state[94])
         );
  DFF \state_reg[78]  ( .D(\w0[1][78] ), .CLK(clk), .RST(rst), .Q(state[78])
         );
  DFF \state_reg[70]  ( .D(\w0[1][70] ), .CLK(clk), .RST(rst), .Q(state[70])
         );
  DFF \state_reg[87]  ( .D(\w0[1][87] ), .CLK(clk), .RST(rst), .Q(state[87])
         );
  DFF \state_reg[79]  ( .D(\w0[1][79] ), .CLK(clk), .RST(rst), .Q(state[79])
         );
  DFF \state_reg[95]  ( .D(\w0[1][95] ), .CLK(clk), .RST(rst), .Q(state[95])
         );
  DFF \state_reg[32]  ( .D(\w0[1][32] ), .CLK(clk), .RST(rst), .Q(state[32])
         );
  DFF \state_reg[56]  ( .D(\w0[1][56] ), .CLK(clk), .RST(rst), .Q(state[56])
         );
  DFF \state_reg[47]  ( .D(\w0[1][47] ), .CLK(clk), .RST(rst), .Q(state[47])
         );
  DFF \state_reg[57]  ( .D(\w0[1][57] ), .CLK(clk), .RST(rst), .Q(state[57])
         );
  DFF \state_reg[48]  ( .D(\w0[1][48] ), .CLK(clk), .RST(rst), .Q(state[48])
         );
  DFF \state_reg[33]  ( .D(\w0[1][33] ), .CLK(clk), .RST(rst), .Q(state[33])
         );
  DFF \state_reg[40]  ( .D(\w0[1][40] ), .CLK(clk), .RST(rst), .Q(state[40])
         );
  DFF \state_reg[58]  ( .D(\w0[1][58] ), .CLK(clk), .RST(rst), .Q(state[58])
         );
  DFF \state_reg[49]  ( .D(\w0[1][49] ), .CLK(clk), .RST(rst), .Q(state[49])
         );
  DFF \state_reg[34]  ( .D(\w0[1][34] ), .CLK(clk), .RST(rst), .Q(state[34])
         );
  DFF \state_reg[41]  ( .D(\w0[1][41] ), .CLK(clk), .RST(rst), .Q(state[41])
         );
  DFF \state_reg[50]  ( .D(\w0[1][50] ), .CLK(clk), .RST(rst), .Q(state[50])
         );
  DFF \state_reg[59]  ( .D(\w0[1][59] ), .CLK(clk), .RST(rst), .Q(state[59])
         );
  DFF \state_reg[35]  ( .D(\w0[1][35] ), .CLK(clk), .RST(rst), .Q(state[35])
         );
  DFF \state_reg[42]  ( .D(\w0[1][42] ), .CLK(clk), .RST(rst), .Q(state[42])
         );
  DFF \state_reg[60]  ( .D(\w0[1][60] ), .CLK(clk), .RST(rst), .Q(state[60])
         );
  DFF \state_reg[36]  ( .D(\w0[1][36] ), .CLK(clk), .RST(rst), .Q(state[36])
         );
  DFF \state_reg[51]  ( .D(\w0[1][51] ), .CLK(clk), .RST(rst), .Q(state[51])
         );
  DFF \state_reg[43]  ( .D(\w0[1][43] ), .CLK(clk), .RST(rst), .Q(state[43])
         );
  DFF \state_reg[61]  ( .D(\w0[1][61] ), .CLK(clk), .RST(rst), .Q(state[61])
         );
  DFF \state_reg[37]  ( .D(\w0[1][37] ), .CLK(clk), .RST(rst), .Q(state[37])
         );
  DFF \state_reg[52]  ( .D(\w0[1][52] ), .CLK(clk), .RST(rst), .Q(state[52])
         );
  DFF \state_reg[44]  ( .D(\w0[1][44] ), .CLK(clk), .RST(rst), .Q(state[44])
         );
  DFF \state_reg[53]  ( .D(\w0[1][53] ), .CLK(clk), .RST(rst), .Q(state[53])
         );
  DFF \state_reg[62]  ( .D(\w0[1][62] ), .CLK(clk), .RST(rst), .Q(state[62])
         );
  DFF \state_reg[38]  ( .D(\w0[1][38] ), .CLK(clk), .RST(rst), .Q(state[38])
         );
  DFF \state_reg[45]  ( .D(\w0[1][45] ), .CLK(clk), .RST(rst), .Q(state[45])
         );
  DFF \state_reg[63]  ( .D(\w0[1][63] ), .CLK(clk), .RST(rst), .Q(state[63])
         );
  DFF \state_reg[39]  ( .D(\w0[1][39] ), .CLK(clk), .RST(rst), .Q(state[39])
         );
  DFF \state_reg[55]  ( .D(\w0[1][55] ), .CLK(clk), .RST(rst), .Q(state[55])
         );
  DFF \state_reg[54]  ( .D(\w0[1][54] ), .CLK(clk), .RST(rst), .Q(state[54])
         );
  DFF \state_reg[46]  ( .D(\w0[1][46] ), .CLK(clk), .RST(rst), .Q(state[46])
         );
  DFF \state_reg[8]  ( .D(\w0[1][8] ), .CLK(clk), .RST(rst), .Q(state[8]) );
  DFF \state_reg[23]  ( .D(\w0[1][23] ), .CLK(clk), .RST(rst), .Q(state[23])
         );
  DFF \state_reg[1]  ( .D(\w0[1][1] ), .CLK(clk), .RST(rst), .Q(state[1]) );
  DFF \state_reg[16]  ( .D(\w0[1][16] ), .CLK(clk), .RST(rst), .Q(state[16])
         );
  DFF \state_reg[24]  ( .D(\w0[1][24] ), .CLK(clk), .RST(rst), .Q(state[24])
         );
  DFF \state_reg[9]  ( .D(\w0[1][9] ), .CLK(clk), .RST(rst), .Q(state[9]) );
  DFF \state_reg[10]  ( .D(\w0[1][10] ), .CLK(clk), .RST(rst), .Q(state[10])
         );
  DFF \state_reg[2]  ( .D(\w0[1][2] ), .CLK(clk), .RST(rst), .Q(state[2]) );
  DFF \state_reg[17]  ( .D(\w0[1][17] ), .CLK(clk), .RST(rst), .Q(state[17])
         );
  DFF \state_reg[25]  ( .D(\w0[1][25] ), .CLK(clk), .RST(rst), .Q(state[25])
         );
  DFF \state_reg[11]  ( .D(\w0[1][11] ), .CLK(clk), .RST(rst), .Q(state[11])
         );
  DFF \state_reg[3]  ( .D(\w0[1][3] ), .CLK(clk), .RST(rst), .Q(state[3]) );
  DFF \state_reg[18]  ( .D(\w0[1][18] ), .CLK(clk), .RST(rst), .Q(state[18])
         );
  DFF \state_reg[26]  ( .D(\w0[1][26] ), .CLK(clk), .RST(rst), .Q(state[26])
         );
  DFF \state_reg[12]  ( .D(\w0[1][12] ), .CLK(clk), .RST(rst), .Q(state[12])
         );
  DFF \state_reg[27]  ( .D(\w0[1][27] ), .CLK(clk), .RST(rst), .Q(state[27])
         );
  DFF \state_reg[19]  ( .D(\w0[1][19] ), .CLK(clk), .RST(rst), .Q(state[19])
         );
  DFF \state_reg[4]  ( .D(\w0[1][4] ), .CLK(clk), .RST(rst), .Q(state[4]) );
  DFF \state_reg[13]  ( .D(\w0[1][13] ), .CLK(clk), .RST(rst), .Q(state[13])
         );
  DFF \state_reg[28]  ( .D(\w0[1][28] ), .CLK(clk), .RST(rst), .Q(state[28])
         );
  DFF \state_reg[20]  ( .D(\w0[1][20] ), .CLK(clk), .RST(rst), .Q(state[20])
         );
  DFF \state_reg[5]  ( .D(\w0[1][5] ), .CLK(clk), .RST(rst), .Q(state[5]) );
  DFF \state_reg[14]  ( .D(\w0[1][14] ), .CLK(clk), .RST(rst), .Q(state[14])
         );
  DFF \state_reg[6]  ( .D(\w0[1][6] ), .CLK(clk), .RST(rst), .Q(state[6]) );
  DFF \state_reg[21]  ( .D(\w0[1][21] ), .CLK(clk), .RST(rst), .Q(state[21])
         );
  DFF \state_reg[29]  ( .D(\w0[1][29] ), .CLK(clk), .RST(rst), .Q(state[29])
         );
  DFF \state_reg[15]  ( .D(\w0[1][15] ), .CLK(clk), .RST(rst), .Q(state[15])
         );
  DFF \state_reg[30]  ( .D(\w0[1][30] ), .CLK(clk), .RST(rst), .Q(state[30])
         );
  DFF \state_reg[22]  ( .D(\w0[1][22] ), .CLK(clk), .RST(rst), .Q(state[22])
         );
  DFF \state_reg[7]  ( .D(\w0[1][7] ), .CLK(clk), .RST(rst), .Q(state[7]) );
  DFF \state_reg[31]  ( .D(\w0[1][31] ), .CLK(clk), .RST(rst), .Q(state[31])
         );
  DFF \state_reg[127]  ( .D(\w0[1][127] ), .CLK(clk), .RST(rst), .Q(state[127]) );
  DFF \state_reg[104]  ( .D(\w0[1][104] ), .CLK(clk), .RST(rst), .Q(state[104]) );
  DFF \state_reg[112]  ( .D(\w0[1][112] ), .CLK(clk), .RST(rst), .Q(state[112]) );
  DFF \state_reg[96]  ( .D(\w0[1][96] ), .CLK(clk), .RST(rst), .Q(state[96])
         );
  DFF \state_reg[113]  ( .D(\w0[1][113] ), .CLK(clk), .RST(rst), .Q(state[113]) );
  DFF \state_reg[105]  ( .D(\w0[1][105] ), .CLK(clk), .RST(rst), .Q(state[105]) );
  DFF \state_reg[120]  ( .D(\w0[1][120] ), .CLK(clk), .RST(rst), .Q(state[120]) );
  DFF \state_reg[97]  ( .D(\w0[1][97] ), .CLK(clk), .RST(rst), .Q(state[97])
         );
  DFF \state_reg[114]  ( .D(\w0[1][114] ), .CLK(clk), .RST(rst), .Q(state[114]) );
  DFF \state_reg[106]  ( .D(\w0[1][106] ), .CLK(clk), .RST(rst), .Q(state[106]) );
  DFF \state_reg[121]  ( .D(\w0[1][121] ), .CLK(clk), .RST(rst), .Q(state[121]) );
  DFF \state_reg[98]  ( .D(\w0[1][98] ), .CLK(clk), .RST(rst), .Q(state[98])
         );
  DFF \state_reg[115]  ( .D(\w0[1][115] ), .CLK(clk), .RST(rst), .Q(state[115]) );
  DFF \state_reg[107]  ( .D(\w0[1][107] ), .CLK(clk), .RST(rst), .Q(state[107]) );
  DFF \state_reg[122]  ( .D(\w0[1][122] ), .CLK(clk), .RST(rst), .Q(state[122]) );
  DFF \state_reg[116]  ( .D(\w0[1][116] ), .CLK(clk), .RST(rst), .Q(state[116]) );
  DFF \state_reg[108]  ( .D(\w0[1][108] ), .CLK(clk), .RST(rst), .Q(state[108]) );
  DFF \state_reg[99]  ( .D(\w0[1][99] ), .CLK(clk), .RST(rst), .Q(state[99])
         );
  DFF \state_reg[123]  ( .D(\w0[1][123] ), .CLK(clk), .RST(rst), .Q(state[123]) );
  DFF \state_reg[124]  ( .D(\w0[1][124] ), .CLK(clk), .RST(rst), .Q(state[124]) );
  DFF \state_reg[100]  ( .D(\w0[1][100] ), .CLK(clk), .RST(rst), .Q(state[100]) );
  DFF \state_reg[117]  ( .D(\w0[1][117] ), .CLK(clk), .RST(rst), .Q(state[117]) );
  DFF \state_reg[109]  ( .D(\w0[1][109] ), .CLK(clk), .RST(rst), .Q(state[109]) );
  DFF \state_reg[118]  ( .D(\w0[1][118] ), .CLK(clk), .RST(rst), .Q(state[118]) );
  DFF \state_reg[110]  ( .D(\w0[1][110] ), .CLK(clk), .RST(rst), .Q(state[110]) );
  DFF \state_reg[101]  ( .D(\w0[1][101] ), .CLK(clk), .RST(rst), .Q(state[101]) );
  DFF \state_reg[125]  ( .D(\w0[1][125] ), .CLK(clk), .RST(rst), .Q(state[125]) );
  DFF \state_reg[103]  ( .D(\w0[1][103] ), .CLK(clk), .RST(rst), .Q(state[103]) );
  DFF \state_reg[126]  ( .D(\w0[1][126] ), .CLK(clk), .RST(rst), .Q(state[126]) );
  DFF \state_reg[102]  ( .D(\w0[1][102] ), .CLK(clk), .RST(rst), .Q(state[102]) );
  DFF \state_reg[119]  ( .D(\w0[1][119] ), .CLK(clk), .RST(rst), .Q(state[119]) );
  DFF \state_reg[111]  ( .D(\w0[1][111] ), .CLK(clk), .RST(rst), .Q(state[111]) );
  XOR U1218 ( .A(n979), .B(\w3[0][7] ), .Z(n704) );
  XNOR U1219 ( .A(n950), .B(n704), .Z(\w0[1][31] ) );
  XOR U1220 ( .A(\w3[0][114] ), .B(\w3[0][122] ), .Z(n705) );
  XNOR U1221 ( .A(\w3[0][97] ), .B(n1003), .Z(n706) );
  XNOR U1222 ( .A(n705), .B(n706), .Z(\w0[1][121] ) );
  XNOR U1223 ( .A(\w3[0][13] ), .B(n826), .Z(n707) );
  XNOR U1224 ( .A(n797), .B(n707), .Z(\w0[1][21] ) );
  XOR U1225 ( .A(n979), .B(n978), .Z(n708) );
  XNOR U1226 ( .A(\w3[0][0] ), .B(\w3[0][1] ), .Z(n709) );
  XOR U1227 ( .A(n708), .B(n709), .Z(\w0[1][8] ) );
  XNOR U1228 ( .A(\w3[0][45] ), .B(n879), .Z(n710) );
  XNOR U1229 ( .A(n878), .B(n710), .Z(\w0[1][53] ) );
  XOR U1230 ( .A(\w3[0][41] ), .B(n893), .Z(n711) );
  XNOR U1231 ( .A(n866), .B(n711), .Z(\w0[1][49] ) );
  XNOR U1232 ( .A(\w3[0][77] ), .B(n964), .Z(n712) );
  XNOR U1233 ( .A(n963), .B(n712), .Z(\w0[1][85] ) );
  XOR U1234 ( .A(\w3[0][73] ), .B(n980), .Z(n713) );
  XNOR U1235 ( .A(n954), .B(n713), .Z(\w0[1][81] ) );
  IV U1236 ( .A(init), .Z(n714) );
  XOR U1237 ( .A(key[128]), .B(\w3[1][0] ), .Z(out[0]) );
  XOR U1238 ( .A(key[228]), .B(\w3[1][100] ), .Z(out[100]) );
  XOR U1239 ( .A(key[229]), .B(\w3[1][101] ), .Z(out[101]) );
  XOR U1240 ( .A(key[230]), .B(\w3[1][102] ), .Z(out[102]) );
  XOR U1241 ( .A(key[231]), .B(\w3[1][103] ), .Z(out[103]) );
  XOR U1242 ( .A(key[232]), .B(\w3[1][104] ), .Z(out[104]) );
  XOR U1243 ( .A(key[233]), .B(\w3[1][105] ), .Z(out[105]) );
  XOR U1244 ( .A(key[234]), .B(\w3[1][106] ), .Z(out[106]) );
  XOR U1245 ( .A(key[235]), .B(\w3[1][107] ), .Z(out[107]) );
  XOR U1246 ( .A(key[236]), .B(\w3[1][108] ), .Z(out[108]) );
  XOR U1247 ( .A(key[237]), .B(\w3[1][109] ), .Z(out[109]) );
  XOR U1248 ( .A(key[138]), .B(\w3[1][10] ), .Z(out[10]) );
  XOR U1249 ( .A(key[238]), .B(\w3[1][110] ), .Z(out[110]) );
  XOR U1250 ( .A(key[239]), .B(\w3[1][111] ), .Z(out[111]) );
  XOR U1251 ( .A(key[240]), .B(\w3[1][112] ), .Z(out[112]) );
  XOR U1252 ( .A(key[241]), .B(\w3[1][113] ), .Z(out[113]) );
  XOR U1253 ( .A(key[242]), .B(\w3[1][114] ), .Z(out[114]) );
  XOR U1254 ( .A(key[243]), .B(\w3[1][115] ), .Z(out[115]) );
  XOR U1255 ( .A(key[244]), .B(\w3[1][116] ), .Z(out[116]) );
  XOR U1256 ( .A(key[245]), .B(\w3[1][117] ), .Z(out[117]) );
  XOR U1257 ( .A(key[246]), .B(\w3[1][118] ), .Z(out[118]) );
  XOR U1258 ( .A(key[247]), .B(\w3[1][119] ), .Z(out[119]) );
  XOR U1259 ( .A(key[139]), .B(\w3[1][11] ), .Z(out[11]) );
  XOR U1260 ( .A(key[248]), .B(\w3[1][120] ), .Z(out[120]) );
  XOR U1261 ( .A(key[249]), .B(\w3[1][121] ), .Z(out[121]) );
  XOR U1262 ( .A(key[250]), .B(\w3[1][122] ), .Z(out[122]) );
  XOR U1263 ( .A(key[251]), .B(\w3[1][123] ), .Z(out[123]) );
  XOR U1264 ( .A(key[252]), .B(\w3[1][124] ), .Z(out[124]) );
  XOR U1265 ( .A(key[253]), .B(\w3[1][125] ), .Z(out[125]) );
  XOR U1266 ( .A(key[254]), .B(\w3[1][126] ), .Z(out[126]) );
  XOR U1267 ( .A(key[255]), .B(\w3[1][127] ), .Z(out[127]) );
  XOR U1268 ( .A(key[140]), .B(\w3[1][12] ), .Z(out[12]) );
  XOR U1269 ( .A(key[141]), .B(\w3[1][13] ), .Z(out[13]) );
  XOR U1270 ( .A(key[142]), .B(\w3[1][14] ), .Z(out[14]) );
  XOR U1271 ( .A(key[143]), .B(\w3[1][15] ), .Z(out[15]) );
  XOR U1272 ( .A(key[144]), .B(\w3[1][16] ), .Z(out[16]) );
  XOR U1273 ( .A(key[145]), .B(\w3[1][17] ), .Z(out[17]) );
  XOR U1274 ( .A(key[146]), .B(\w3[1][18] ), .Z(out[18]) );
  XOR U1275 ( .A(key[147]), .B(\w3[1][19] ), .Z(out[19]) );
  XOR U1276 ( .A(key[129]), .B(\w3[1][1] ), .Z(out[1]) );
  XOR U1277 ( .A(key[148]), .B(\w3[1][20] ), .Z(out[20]) );
  XOR U1278 ( .A(key[149]), .B(\w3[1][21] ), .Z(out[21]) );
  XOR U1279 ( .A(key[150]), .B(\w3[1][22] ), .Z(out[22]) );
  XOR U1280 ( .A(key[151]), .B(\w3[1][23] ), .Z(out[23]) );
  XOR U1281 ( .A(key[152]), .B(\w3[1][24] ), .Z(out[24]) );
  XOR U1282 ( .A(key[153]), .B(\w3[1][25] ), .Z(out[25]) );
  XOR U1283 ( .A(key[154]), .B(\w3[1][26] ), .Z(out[26]) );
  XOR U1284 ( .A(key[155]), .B(\w3[1][27] ), .Z(out[27]) );
  XOR U1285 ( .A(key[156]), .B(\w3[1][28] ), .Z(out[28]) );
  XOR U1286 ( .A(key[157]), .B(\w3[1][29] ), .Z(out[29]) );
  XOR U1287 ( .A(key[130]), .B(\w3[1][2] ), .Z(out[2]) );
  XOR U1288 ( .A(key[158]), .B(\w3[1][30] ), .Z(out[30]) );
  XOR U1289 ( .A(key[159]), .B(\w3[1][31] ), .Z(out[31]) );
  XOR U1290 ( .A(key[160]), .B(\w3[1][32] ), .Z(out[32]) );
  XOR U1291 ( .A(key[161]), .B(\w3[1][33] ), .Z(out[33]) );
  XOR U1292 ( .A(key[162]), .B(\w3[1][34] ), .Z(out[34]) );
  XOR U1293 ( .A(key[163]), .B(\w3[1][35] ), .Z(out[35]) );
  XOR U1294 ( .A(key[164]), .B(\w3[1][36] ), .Z(out[36]) );
  XOR U1295 ( .A(key[165]), .B(\w3[1][37] ), .Z(out[37]) );
  XOR U1296 ( .A(key[166]), .B(\w3[1][38] ), .Z(out[38]) );
  XOR U1297 ( .A(key[167]), .B(\w3[1][39] ), .Z(out[39]) );
  XOR U1298 ( .A(key[131]), .B(\w3[1][3] ), .Z(out[3]) );
  XOR U1299 ( .A(key[168]), .B(\w3[1][40] ), .Z(out[40]) );
  XOR U1300 ( .A(key[169]), .B(\w3[1][41] ), .Z(out[41]) );
  XOR U1301 ( .A(key[170]), .B(\w3[1][42] ), .Z(out[42]) );
  XOR U1302 ( .A(key[171]), .B(\w3[1][43] ), .Z(out[43]) );
  XOR U1303 ( .A(key[172]), .B(\w3[1][44] ), .Z(out[44]) );
  XOR U1304 ( .A(key[173]), .B(\w3[1][45] ), .Z(out[45]) );
  XOR U1305 ( .A(key[174]), .B(\w3[1][46] ), .Z(out[46]) );
  XOR U1306 ( .A(key[175]), .B(\w3[1][47] ), .Z(out[47]) );
  XOR U1307 ( .A(key[176]), .B(\w3[1][48] ), .Z(out[48]) );
  XOR U1308 ( .A(key[177]), .B(\w3[1][49] ), .Z(out[49]) );
  XOR U1309 ( .A(key[132]), .B(\w3[1][4] ), .Z(out[4]) );
  XOR U1310 ( .A(key[178]), .B(\w3[1][50] ), .Z(out[50]) );
  XOR U1311 ( .A(key[179]), .B(\w3[1][51] ), .Z(out[51]) );
  XOR U1312 ( .A(key[180]), .B(\w3[1][52] ), .Z(out[52]) );
  XOR U1313 ( .A(key[181]), .B(\w3[1][53] ), .Z(out[53]) );
  XOR U1314 ( .A(key[182]), .B(\w3[1][54] ), .Z(out[54]) );
  XOR U1315 ( .A(key[183]), .B(\w3[1][55] ), .Z(out[55]) );
  XOR U1316 ( .A(key[184]), .B(\w3[1][56] ), .Z(out[56]) );
  XOR U1317 ( .A(key[185]), .B(\w3[1][57] ), .Z(out[57]) );
  XOR U1318 ( .A(key[186]), .B(\w3[1][58] ), .Z(out[58]) );
  XOR U1319 ( .A(key[187]), .B(\w3[1][59] ), .Z(out[59]) );
  XOR U1320 ( .A(key[133]), .B(\w3[1][5] ), .Z(out[5]) );
  XOR U1321 ( .A(key[188]), .B(\w3[1][60] ), .Z(out[60]) );
  XOR U1322 ( .A(key[189]), .B(\w3[1][61] ), .Z(out[61]) );
  XOR U1323 ( .A(key[190]), .B(\w3[1][62] ), .Z(out[62]) );
  XOR U1324 ( .A(key[191]), .B(\w3[1][63] ), .Z(out[63]) );
  XOR U1325 ( .A(key[192]), .B(\w3[1][64] ), .Z(out[64]) );
  XOR U1326 ( .A(key[193]), .B(\w3[1][65] ), .Z(out[65]) );
  XOR U1327 ( .A(key[194]), .B(\w3[1][66] ), .Z(out[66]) );
  XOR U1328 ( .A(key[195]), .B(\w3[1][67] ), .Z(out[67]) );
  XOR U1329 ( .A(key[196]), .B(\w3[1][68] ), .Z(out[68]) );
  XOR U1330 ( .A(key[197]), .B(\w3[1][69] ), .Z(out[69]) );
  XOR U1331 ( .A(key[134]), .B(\w3[1][6] ), .Z(out[6]) );
  XOR U1332 ( .A(key[198]), .B(\w3[1][70] ), .Z(out[70]) );
  XOR U1333 ( .A(key[199]), .B(\w3[1][71] ), .Z(out[71]) );
  XOR U1334 ( .A(key[200]), .B(\w3[1][72] ), .Z(out[72]) );
  XOR U1335 ( .A(key[201]), .B(\w3[1][73] ), .Z(out[73]) );
  XOR U1336 ( .A(key[202]), .B(\w3[1][74] ), .Z(out[74]) );
  XOR U1337 ( .A(key[203]), .B(\w3[1][75] ), .Z(out[75]) );
  XOR U1338 ( .A(key[204]), .B(\w3[1][76] ), .Z(out[76]) );
  XOR U1339 ( .A(key[205]), .B(\w3[1][77] ), .Z(out[77]) );
  XOR U1340 ( .A(key[206]), .B(\w3[1][78] ), .Z(out[78]) );
  XOR U1341 ( .A(key[207]), .B(\w3[1][79] ), .Z(out[79]) );
  XOR U1342 ( .A(key[135]), .B(\w3[1][7] ), .Z(out[7]) );
  XOR U1343 ( .A(key[208]), .B(\w3[1][80] ), .Z(out[80]) );
  XOR U1344 ( .A(key[209]), .B(\w3[1][81] ), .Z(out[81]) );
  XOR U1345 ( .A(key[210]), .B(\w3[1][82] ), .Z(out[82]) );
  XOR U1346 ( .A(key[211]), .B(\w3[1][83] ), .Z(out[83]) );
  XOR U1347 ( .A(key[212]), .B(\w3[1][84] ), .Z(out[84]) );
  XOR U1348 ( .A(key[213]), .B(\w3[1][85] ), .Z(out[85]) );
  XOR U1349 ( .A(key[214]), .B(\w3[1][86] ), .Z(out[86]) );
  XOR U1350 ( .A(key[215]), .B(\w3[1][87] ), .Z(out[87]) );
  XOR U1351 ( .A(key[216]), .B(\w3[1][88] ), .Z(out[88]) );
  XOR U1352 ( .A(key[217]), .B(\w3[1][89] ), .Z(out[89]) );
  XOR U1353 ( .A(key[136]), .B(\w3[1][8] ), .Z(out[8]) );
  XOR U1354 ( .A(key[218]), .B(\w3[1][90] ), .Z(out[90]) );
  XOR U1355 ( .A(key[219]), .B(\w3[1][91] ), .Z(out[91]) );
  XOR U1356 ( .A(key[220]), .B(\w3[1][92] ), .Z(out[92]) );
  XOR U1357 ( .A(key[221]), .B(\w3[1][93] ), .Z(out[93]) );
  XOR U1358 ( .A(key[222]), .B(\w3[1][94] ), .Z(out[94]) );
  XOR U1359 ( .A(key[223]), .B(\w3[1][95] ), .Z(out[95]) );
  XOR U1360 ( .A(key[224]), .B(\w3[1][96] ), .Z(out[96]) );
  XOR U1361 ( .A(key[225]), .B(\w3[1][97] ), .Z(out[97]) );
  XOR U1362 ( .A(key[226]), .B(\w3[1][98] ), .Z(out[98]) );
  XOR U1363 ( .A(key[227]), .B(\w3[1][99] ), .Z(out[99]) );
  XOR U1364 ( .A(key[137]), .B(\w3[1][9] ), .Z(out[9]) );
  XNOR U1365 ( .A(\w3[0][1] ), .B(\w3[0][25] ), .Z(n1010) );
  XOR U1366 ( .A(\w3[0][16] ), .B(\w3[0][24] ), .Z(n979) );
  XOR U1367 ( .A(n1010), .B(n979), .Z(n715) );
  XNOR U1368 ( .A(\w3[0][8] ), .B(n715), .Z(\w0[1][0] ) );
  XOR U1369 ( .A(\w3[0][96] ), .B(\w3[0][101] ), .Z(n733) );
  XOR U1370 ( .A(\w3[0][108] ), .B(\w3[0][116] ), .Z(n717) );
  IV U1371 ( .A(\w3[0][120] ), .Z(n765) );
  XOR U1372 ( .A(n765), .B(\w3[0][125] ), .Z(n716) );
  XOR U1373 ( .A(n717), .B(n716), .Z(n770) );
  XOR U1374 ( .A(\w3[0][124] ), .B(n770), .Z(n718) );
  XNOR U1375 ( .A(n733), .B(n718), .Z(\w0[1][100] ) );
  XNOR U1376 ( .A(\w3[0][102] ), .B(\w3[0][126] ), .Z(n739) );
  XNOR U1377 ( .A(\w3[0][109] ), .B(\w3[0][117] ), .Z(n773) );
  XOR U1378 ( .A(\w3[0][125] ), .B(n773), .Z(n719) );
  XOR U1379 ( .A(n739), .B(n719), .Z(\w0[1][101] ) );
  XOR U1380 ( .A(\w3[0][96] ), .B(\w3[0][103] ), .Z(n740) );
  XNOR U1381 ( .A(\w3[0][110] ), .B(\w3[0][118] ), .Z(n750) );
  XNOR U1382 ( .A(n765), .B(\w3[0][127] ), .Z(n721) );
  XOR U1383 ( .A(n750), .B(n721), .Z(n776) );
  XOR U1384 ( .A(\w3[0][126] ), .B(n776), .Z(n720) );
  XNOR U1385 ( .A(n740), .B(n720), .Z(\w0[1][102] ) );
  XOR U1386 ( .A(\w3[0][111] ), .B(\w3[0][119] ), .Z(n780) );
  XOR U1387 ( .A(\w3[0][96] ), .B(n721), .Z(n722) );
  XOR U1388 ( .A(n780), .B(n722), .Z(\w0[1][103] ) );
  XNOR U1389 ( .A(\w3[0][120] ), .B(\w3[0][112] ), .Z(n999) );
  XNOR U1390 ( .A(n999), .B(\w3[0][97] ), .Z(n724) );
  XNOR U1391 ( .A(\w3[0][96] ), .B(\w3[0][105] ), .Z(n723) );
  XNOR U1392 ( .A(n724), .B(n723), .Z(\w0[1][104] ) );
  XNOR U1393 ( .A(\w3[0][97] ), .B(\w3[0][121] ), .Z(n998) );
  XNOR U1394 ( .A(\w3[0][113] ), .B(n998), .Z(n726) );
  XNOR U1395 ( .A(\w3[0][106] ), .B(\w3[0][98] ), .Z(n725) );
  XNOR U1396 ( .A(n726), .B(n725), .Z(\w0[1][105] ) );
  XOR U1397 ( .A(\w3[0][98] ), .B(\w3[0][122] ), .Z(n1001) );
  XOR U1398 ( .A(\w3[0][99] ), .B(n1001), .Z(n728) );
  XNOR U1399 ( .A(\w3[0][107] ), .B(\w3[0][114] ), .Z(n727) );
  XNOR U1400 ( .A(n728), .B(n727), .Z(\w0[1][106] ) );
  XNOR U1401 ( .A(\w3[0][99] ), .B(\w3[0][123] ), .Z(n1004) );
  XOR U1402 ( .A(\w3[0][108] ), .B(n1004), .Z(n729) );
  XOR U1403 ( .A(\w3[0][104] ), .B(n729), .Z(n746) );
  XNOR U1404 ( .A(\w3[0][96] ), .B(\w3[0][100] ), .Z(n1007) );
  XOR U1405 ( .A(\w3[0][115] ), .B(n1007), .Z(n730) );
  XOR U1406 ( .A(n746), .B(n730), .Z(\w0[1][107] ) );
  XOR U1407 ( .A(\w3[0][100] ), .B(\w3[0][104] ), .Z(n732) );
  XNOR U1408 ( .A(\w3[0][124] ), .B(\w3[0][109] ), .Z(n731) );
  XOR U1409 ( .A(n732), .B(n731), .Z(n748) );
  XNOR U1410 ( .A(\w3[0][116] ), .B(n733), .Z(n734) );
  XOR U1411 ( .A(n748), .B(n734), .Z(\w0[1][108] ) );
  XNOR U1412 ( .A(\w3[0][125] ), .B(\w3[0][101] ), .Z(n752) );
  XNOR U1413 ( .A(\w3[0][110] ), .B(n752), .Z(n736) );
  XNOR U1414 ( .A(\w3[0][117] ), .B(\w3[0][102] ), .Z(n735) );
  XNOR U1415 ( .A(n736), .B(n735), .Z(\w0[1][109] ) );
  XNOR U1416 ( .A(\w3[0][2] ), .B(\w3[0][26] ), .Z(n793) );
  XNOR U1417 ( .A(\w3[0][3] ), .B(n793), .Z(n738) );
  XNOR U1418 ( .A(\w3[0][11] ), .B(\w3[0][18] ), .Z(n737) );
  XNOR U1419 ( .A(n738), .B(n737), .Z(\w0[1][10] ) );
  XOR U1420 ( .A(\w3[0][111] ), .B(\w3[0][104] ), .Z(n757) );
  XOR U1421 ( .A(n739), .B(n757), .Z(n753) );
  XNOR U1422 ( .A(\w3[0][118] ), .B(n740), .Z(n741) );
  XOR U1423 ( .A(n753), .B(n741), .Z(\w0[1][110] ) );
  XOR U1424 ( .A(\w3[0][127] ), .B(\w3[0][103] ), .Z(n755) );
  XNOR U1425 ( .A(\w3[0][96] ), .B(\w3[0][104] ), .Z(n760) );
  XOR U1426 ( .A(\w3[0][119] ), .B(n760), .Z(n742) );
  XNOR U1427 ( .A(n755), .B(n742), .Z(\w0[1][111] ) );
  XOR U1428 ( .A(\w3[0][105] ), .B(\w3[0][113] ), .Z(n1003) );
  XNOR U1429 ( .A(n765), .B(n760), .Z(n743) );
  XNOR U1430 ( .A(n1003), .B(n743), .Z(\w0[1][112] ) );
  XOR U1431 ( .A(\w3[0][106] ), .B(\w3[0][114] ), .Z(n1006) );
  XOR U1432 ( .A(\w3[0][105] ), .B(n998), .Z(n744) );
  XNOR U1433 ( .A(n1006), .B(n744), .Z(\w0[1][113] ) );
  XNOR U1434 ( .A(\w3[0][107] ), .B(\w3[0][115] ), .Z(n767) );
  XNOR U1435 ( .A(\w3[0][106] ), .B(n1001), .Z(n745) );
  XOR U1436 ( .A(n767), .B(n745), .Z(\w0[1][114] ) );
  XNOR U1437 ( .A(\w3[0][116] ), .B(\w3[0][112] ), .Z(n768) );
  XOR U1438 ( .A(\w3[0][107] ), .B(n746), .Z(n747) );
  XOR U1439 ( .A(n768), .B(n747), .Z(\w0[1][115] ) );
  XNOR U1440 ( .A(\w3[0][117] ), .B(\w3[0][112] ), .Z(n772) );
  XOR U1441 ( .A(\w3[0][108] ), .B(n748), .Z(n749) );
  XOR U1442 ( .A(n772), .B(n749), .Z(\w0[1][116] ) );
  XOR U1443 ( .A(\w3[0][109] ), .B(n750), .Z(n751) );
  XOR U1444 ( .A(n752), .B(n751), .Z(\w0[1][117] ) );
  XNOR U1445 ( .A(\w3[0][119] ), .B(\w3[0][112] ), .Z(n778) );
  XOR U1446 ( .A(\w3[0][110] ), .B(n753), .Z(n754) );
  XOR U1447 ( .A(n778), .B(n754), .Z(\w0[1][118] ) );
  XOR U1448 ( .A(\w3[0][112] ), .B(n755), .Z(n756) );
  XOR U1449 ( .A(n757), .B(n756), .Z(\w0[1][119] ) );
  XNOR U1450 ( .A(\w3[0][3] ), .B(\w3[0][27] ), .Z(n822) );
  XNOR U1451 ( .A(\w3[0][8] ), .B(\w3[0][12] ), .Z(n758) );
  XNOR U1452 ( .A(n822), .B(n758), .Z(n791) );
  XNOR U1453 ( .A(\w3[0][0] ), .B(\w3[0][4] ), .Z(n841) );
  XOR U1454 ( .A(\w3[0][19] ), .B(n841), .Z(n759) );
  XOR U1455 ( .A(n791), .B(n759), .Z(\w0[1][11] ) );
  XNOR U1456 ( .A(\w3[0][121] ), .B(n760), .Z(n762) );
  XNOR U1457 ( .A(\w3[0][112] ), .B(\w3[0][113] ), .Z(n761) );
  XNOR U1458 ( .A(n762), .B(n761), .Z(\w0[1][120] ) );
  XOR U1459 ( .A(\w3[0][123] ), .B(n1006), .Z(n764) );
  XNOR U1460 ( .A(\w3[0][98] ), .B(\w3[0][115] ), .Z(n763) );
  XNOR U1461 ( .A(n764), .B(n763), .Z(\w0[1][122] ) );
  XOR U1462 ( .A(\w3[0][124] ), .B(n765), .Z(n766) );
  XOR U1463 ( .A(n767), .B(n766), .Z(n1009) );
  XOR U1464 ( .A(\w3[0][99] ), .B(n768), .Z(n769) );
  XNOR U1465 ( .A(n1009), .B(n769), .Z(\w0[1][123] ) );
  XOR U1466 ( .A(n770), .B(\w3[0][100] ), .Z(n771) );
  XOR U1467 ( .A(n772), .B(n771), .Z(\w0[1][124] ) );
  XOR U1468 ( .A(\w3[0][126] ), .B(\w3[0][118] ), .Z(n775) );
  XOR U1469 ( .A(\w3[0][101] ), .B(n773), .Z(n774) );
  XNOR U1470 ( .A(n775), .B(n774), .Z(\w0[1][125] ) );
  XOR U1471 ( .A(\w3[0][102] ), .B(n776), .Z(n777) );
  XOR U1472 ( .A(n778), .B(n777), .Z(\w0[1][126] ) );
  XNOR U1473 ( .A(\w3[0][103] ), .B(n999), .Z(n779) );
  XOR U1474 ( .A(n780), .B(n779), .Z(\w0[1][127] ) );
  XOR U1475 ( .A(\w3[0][13] ), .B(\w3[0][28] ), .Z(n782) );
  XNOR U1476 ( .A(\w3[0][8] ), .B(\w3[0][4] ), .Z(n781) );
  XOR U1477 ( .A(n782), .B(n781), .Z(n795) );
  XNOR U1478 ( .A(\w3[0][0] ), .B(\w3[0][5] ), .Z(n867) );
  XOR U1479 ( .A(\w3[0][20] ), .B(n867), .Z(n783) );
  XOR U1480 ( .A(n795), .B(n783), .Z(\w0[1][12] ) );
  XNOR U1481 ( .A(\w3[0][5] ), .B(\w3[0][29] ), .Z(n797) );
  XNOR U1482 ( .A(\w3[0][21] ), .B(n797), .Z(n785) );
  XNOR U1483 ( .A(\w3[0][14] ), .B(\w3[0][6] ), .Z(n784) );
  XNOR U1484 ( .A(n785), .B(n784), .Z(\w0[1][13] ) );
  XNOR U1485 ( .A(\w3[0][6] ), .B(\w3[0][30] ), .Z(n899) );
  XOR U1486 ( .A(\w3[0][8] ), .B(\w3[0][15] ), .Z(n802) );
  XOR U1487 ( .A(n899), .B(n802), .Z(n798) );
  XNOR U1488 ( .A(\w3[0][0] ), .B(\w3[0][7] ), .Z(n923) );
  XOR U1489 ( .A(\w3[0][22] ), .B(n923), .Z(n786) );
  XOR U1490 ( .A(n798), .B(n786), .Z(\w0[1][14] ) );
  XNOR U1491 ( .A(\w3[0][7] ), .B(\w3[0][31] ), .Z(n800) );
  XOR U1492 ( .A(\w3[0][8] ), .B(\w3[0][0] ), .Z(n803) );
  XNOR U1493 ( .A(\w3[0][23] ), .B(n803), .Z(n787) );
  XOR U1494 ( .A(n800), .B(n787), .Z(\w0[1][15] ) );
  XOR U1495 ( .A(\w3[0][17] ), .B(\w3[0][9] ), .Z(n806) );
  XNOR U1496 ( .A(\w3[0][24] ), .B(n803), .Z(n788) );
  XNOR U1497 ( .A(n806), .B(n788), .Z(\w0[1][16] ) );
  XOR U1498 ( .A(\w3[0][18] ), .B(\w3[0][10] ), .Z(n824) );
  IV U1499 ( .A(\w3[0][9] ), .Z(n978) );
  XNOR U1500 ( .A(n1010), .B(n978), .Z(n789) );
  XNOR U1501 ( .A(n824), .B(n789), .Z(\w0[1][17] ) );
  XNOR U1502 ( .A(\w3[0][11] ), .B(\w3[0][19] ), .Z(n812) );
  XOR U1503 ( .A(n793), .B(\w3[0][10] ), .Z(n790) );
  XOR U1504 ( .A(n812), .B(n790), .Z(\w0[1][18] ) );
  XNOR U1505 ( .A(\w3[0][16] ), .B(\w3[0][20] ), .Z(n813) );
  XOR U1506 ( .A(\w3[0][11] ), .B(n791), .Z(n792) );
  XOR U1507 ( .A(n813), .B(n792), .Z(\w0[1][19] ) );
  XOR U1508 ( .A(\w3[0][25] ), .B(n793), .Z(n794) );
  XNOR U1509 ( .A(n806), .B(n794), .Z(\w0[1][1] ) );
  IV U1510 ( .A(\w3[0][21] ), .Z(n819) );
  XOR U1511 ( .A(\w3[0][16] ), .B(n819), .Z(n817) );
  XOR U1512 ( .A(\w3[0][12] ), .B(n795), .Z(n796) );
  XOR U1513 ( .A(n817), .B(n796), .Z(\w0[1][20] ) );
  XNOR U1514 ( .A(\w3[0][14] ), .B(\w3[0][22] ), .Z(n826) );
  XNOR U1515 ( .A(\w3[0][16] ), .B(\w3[0][23] ), .Z(n827) );
  XOR U1516 ( .A(\w3[0][14] ), .B(n798), .Z(n799) );
  XOR U1517 ( .A(n827), .B(n799), .Z(\w0[1][22] ) );
  XNOR U1518 ( .A(\w3[0][16] ), .B(n800), .Z(n801) );
  XOR U1519 ( .A(n802), .B(n801), .Z(\w0[1][23] ) );
  XOR U1520 ( .A(n803), .B(\w3[0][17] ), .Z(n805) );
  XNOR U1521 ( .A(\w3[0][25] ), .B(\w3[0][16] ), .Z(n804) );
  XNOR U1522 ( .A(n805), .B(n804), .Z(\w0[1][24] ) );
  XOR U1523 ( .A(\w3[0][26] ), .B(n806), .Z(n808) );
  XNOR U1524 ( .A(\w3[0][1] ), .B(\w3[0][18] ), .Z(n807) );
  XNOR U1525 ( .A(n808), .B(n807), .Z(\w0[1][25] ) );
  XOR U1526 ( .A(\w3[0][27] ), .B(n824), .Z(n810) );
  XNOR U1527 ( .A(\w3[0][2] ), .B(\w3[0][19] ), .Z(n809) );
  XNOR U1528 ( .A(n810), .B(n809), .Z(\w0[1][26] ) );
  IV U1529 ( .A(\w3[0][24] ), .Z(n825) );
  XOR U1530 ( .A(n825), .B(\w3[0][28] ), .Z(n811) );
  XOR U1531 ( .A(n812), .B(n811), .Z(n843) );
  XOR U1532 ( .A(\w3[0][3] ), .B(n813), .Z(n814) );
  XNOR U1533 ( .A(n843), .B(n814), .Z(\w0[1][27] ) );
  XOR U1534 ( .A(\w3[0][20] ), .B(\w3[0][29] ), .Z(n816) );
  XOR U1535 ( .A(n825), .B(\w3[0][12] ), .Z(n815) );
  XOR U1536 ( .A(n816), .B(n815), .Z(n869) );
  XOR U1537 ( .A(\w3[0][4] ), .B(n817), .Z(n818) );
  XOR U1538 ( .A(n869), .B(n818), .Z(\w0[1][28] ) );
  XOR U1539 ( .A(\w3[0][13] ), .B(n819), .Z(n901) );
  XNOR U1540 ( .A(\w3[0][30] ), .B(n901), .Z(n821) );
  XNOR U1541 ( .A(\w3[0][5] ), .B(\w3[0][22] ), .Z(n820) );
  XNOR U1542 ( .A(n821), .B(n820), .Z(\w0[1][29] ) );
  XOR U1543 ( .A(\w3[0][26] ), .B(n822), .Z(n823) );
  XNOR U1544 ( .A(n824), .B(n823), .Z(\w0[1][2] ) );
  XNOR U1545 ( .A(n825), .B(\w3[0][31] ), .Z(n952) );
  XOR U1546 ( .A(n826), .B(n952), .Z(n925) );
  XOR U1547 ( .A(\w3[0][6] ), .B(n827), .Z(n828) );
  XOR U1548 ( .A(n925), .B(n828), .Z(\w0[1][30] ) );
  XNOR U1549 ( .A(\w3[0][15] ), .B(\w3[0][23] ), .Z(n950) );
  XOR U1550 ( .A(\w3[0][33] ), .B(\w3[0][57] ), .Z(n866) );
  XNOR U1551 ( .A(\w3[0][48] ), .B(\w3[0][56] ), .Z(n911) );
  XOR U1552 ( .A(n911), .B(\w3[0][40] ), .Z(n829) );
  XNOR U1553 ( .A(n866), .B(n829), .Z(\w0[1][32] ) );
  XOR U1554 ( .A(\w3[0][34] ), .B(\w3[0][58] ), .Z(n870) );
  XOR U1555 ( .A(\w3[0][41] ), .B(\w3[0][49] ), .Z(n889) );
  XNOR U1556 ( .A(\w3[0][57] ), .B(n889), .Z(n830) );
  XNOR U1557 ( .A(n870), .B(n830), .Z(\w0[1][33] ) );
  XNOR U1558 ( .A(\w3[0][35] ), .B(\w3[0][59] ), .Z(n850) );
  XNOR U1559 ( .A(\w3[0][42] ), .B(\w3[0][50] ), .Z(n893) );
  XOR U1560 ( .A(\w3[0][58] ), .B(n893), .Z(n831) );
  XOR U1561 ( .A(n850), .B(n831), .Z(\w0[1][34] ) );
  XOR U1562 ( .A(\w3[0][36] ), .B(\w3[0][32] ), .Z(n852) );
  XNOR U1563 ( .A(\w3[0][43] ), .B(\w3[0][51] ), .Z(n872) );
  XOR U1564 ( .A(\w3[0][56] ), .B(n872), .Z(n832) );
  XNOR U1565 ( .A(\w3[0][60] ), .B(n832), .Z(n896) );
  XNOR U1566 ( .A(\w3[0][59] ), .B(n896), .Z(n833) );
  XNOR U1567 ( .A(n852), .B(n833), .Z(\w0[1][35] ) );
  XOR U1568 ( .A(\w3[0][32] ), .B(\w3[0][37] ), .Z(n856) );
  XOR U1569 ( .A(\w3[0][44] ), .B(\w3[0][52] ), .Z(n835) );
  XNOR U1570 ( .A(\w3[0][56] ), .B(\w3[0][61] ), .Z(n834) );
  XOR U1571 ( .A(n835), .B(n834), .Z(n902) );
  XOR U1572 ( .A(\w3[0][60] ), .B(n902), .Z(n836) );
  XNOR U1573 ( .A(n856), .B(n836), .Z(\w0[1][36] ) );
  XNOR U1574 ( .A(\w3[0][38] ), .B(\w3[0][62] ), .Z(n861) );
  IV U1575 ( .A(\w3[0][53] ), .Z(n875) );
  XOR U1576 ( .A(\w3[0][45] ), .B(n875), .Z(n905) );
  XOR U1577 ( .A(\w3[0][61] ), .B(n905), .Z(n837) );
  XOR U1578 ( .A(n861), .B(n837), .Z(\w0[1][37] ) );
  XOR U1579 ( .A(\w3[0][32] ), .B(\w3[0][39] ), .Z(n862) );
  XNOR U1580 ( .A(\w3[0][46] ), .B(\w3[0][54] ), .Z(n878) );
  XOR U1581 ( .A(\w3[0][56] ), .B(\w3[0][63] ), .Z(n839) );
  XOR U1582 ( .A(n878), .B(n839), .Z(n908) );
  XOR U1583 ( .A(\w3[0][62] ), .B(n908), .Z(n838) );
  XNOR U1584 ( .A(n862), .B(n838), .Z(\w0[1][38] ) );
  XOR U1585 ( .A(\w3[0][47] ), .B(\w3[0][55] ), .Z(n913) );
  XOR U1586 ( .A(\w3[0][32] ), .B(n839), .Z(n840) );
  XOR U1587 ( .A(n913), .B(n840), .Z(\w0[1][39] ) );
  XOR U1588 ( .A(n841), .B(\w3[0][27] ), .Z(n842) );
  XNOR U1589 ( .A(n843), .B(n842), .Z(\w0[1][3] ) );
  XOR U1590 ( .A(\w3[0][41] ), .B(\w3[0][32] ), .Z(n845) );
  IV U1591 ( .A(\w3[0][33] ), .Z(n890) );
  XNOR U1592 ( .A(n911), .B(n890), .Z(n844) );
  XNOR U1593 ( .A(n845), .B(n844), .Z(\w0[1][40] ) );
  XOR U1594 ( .A(\w3[0][34] ), .B(\w3[0][42] ), .Z(n847) );
  XNOR U1595 ( .A(n866), .B(\w3[0][49] ), .Z(n846) );
  XNOR U1596 ( .A(n847), .B(n846), .Z(\w0[1][41] ) );
  XOR U1597 ( .A(\w3[0][35] ), .B(\w3[0][43] ), .Z(n849) );
  XNOR U1598 ( .A(n870), .B(\w3[0][50] ), .Z(n848) );
  XNOR U1599 ( .A(n849), .B(n848), .Z(\w0[1][42] ) );
  IV U1600 ( .A(\w3[0][40] ), .Z(n860) );
  XNOR U1601 ( .A(n860), .B(n850), .Z(n851) );
  XOR U1602 ( .A(\w3[0][44] ), .B(n851), .Z(n873) );
  XNOR U1603 ( .A(\w3[0][51] ), .B(n852), .Z(n853) );
  XOR U1604 ( .A(n873), .B(n853), .Z(\w0[1][43] ) );
  XOR U1605 ( .A(\w3[0][36] ), .B(\w3[0][45] ), .Z(n855) );
  XOR U1606 ( .A(n860), .B(\w3[0][60] ), .Z(n854) );
  XOR U1607 ( .A(n855), .B(n854), .Z(n876) );
  XNOR U1608 ( .A(\w3[0][52] ), .B(n856), .Z(n857) );
  XOR U1609 ( .A(n876), .B(n857), .Z(\w0[1][44] ) );
  XNOR U1610 ( .A(\w3[0][61] ), .B(\w3[0][37] ), .Z(n879) );
  XNOR U1611 ( .A(\w3[0][46] ), .B(n879), .Z(n859) );
  XOR U1612 ( .A(n875), .B(\w3[0][38] ), .Z(n858) );
  XNOR U1613 ( .A(n859), .B(n858), .Z(\w0[1][45] ) );
  XNOR U1614 ( .A(n860), .B(\w3[0][47] ), .Z(n884) );
  XOR U1615 ( .A(n861), .B(n884), .Z(n880) );
  XNOR U1616 ( .A(\w3[0][54] ), .B(n862), .Z(n863) );
  XOR U1617 ( .A(n880), .B(n863), .Z(\w0[1][46] ) );
  XOR U1618 ( .A(\w3[0][63] ), .B(\w3[0][39] ), .Z(n882) );
  XNOR U1619 ( .A(\w3[0][40] ), .B(\w3[0][32] ), .Z(n885) );
  XOR U1620 ( .A(\w3[0][55] ), .B(n885), .Z(n864) );
  XNOR U1621 ( .A(n882), .B(n864), .Z(\w0[1][47] ) );
  XNOR U1622 ( .A(\w3[0][56] ), .B(n889), .Z(n865) );
  XOR U1623 ( .A(n885), .B(n865), .Z(\w0[1][48] ) );
  XOR U1624 ( .A(n867), .B(\w3[0][28] ), .Z(n868) );
  XOR U1625 ( .A(n869), .B(n868), .Z(\w0[1][4] ) );
  XNOR U1626 ( .A(n870), .B(\w3[0][42] ), .Z(n871) );
  XOR U1627 ( .A(n872), .B(n871), .Z(\w0[1][50] ) );
  IV U1628 ( .A(\w3[0][48] ), .Z(n886) );
  XOR U1629 ( .A(n886), .B(\w3[0][52] ), .Z(n898) );
  XOR U1630 ( .A(\w3[0][43] ), .B(n873), .Z(n874) );
  XOR U1631 ( .A(n898), .B(n874), .Z(\w0[1][51] ) );
  XOR U1632 ( .A(\w3[0][48] ), .B(n875), .Z(n904) );
  XOR U1633 ( .A(\w3[0][44] ), .B(n876), .Z(n877) );
  XOR U1634 ( .A(n904), .B(n877), .Z(\w0[1][52] ) );
  XOR U1635 ( .A(n886), .B(\w3[0][55] ), .Z(n910) );
  XOR U1636 ( .A(\w3[0][46] ), .B(n880), .Z(n881) );
  XOR U1637 ( .A(n910), .B(n881), .Z(\w0[1][54] ) );
  XOR U1638 ( .A(\w3[0][48] ), .B(n882), .Z(n883) );
  XOR U1639 ( .A(n884), .B(n883), .Z(\w0[1][55] ) );
  XNOR U1640 ( .A(\w3[0][49] ), .B(n885), .Z(n888) );
  XOR U1641 ( .A(n886), .B(\w3[0][57] ), .Z(n887) );
  XNOR U1642 ( .A(n888), .B(n887), .Z(\w0[1][56] ) );
  XOR U1643 ( .A(\w3[0][58] ), .B(\w3[0][50] ), .Z(n892) );
  XOR U1644 ( .A(n890), .B(n889), .Z(n891) );
  XNOR U1645 ( .A(n892), .B(n891), .Z(\w0[1][57] ) );
  XOR U1646 ( .A(\w3[0][59] ), .B(\w3[0][51] ), .Z(n895) );
  XOR U1647 ( .A(\w3[0][34] ), .B(n893), .Z(n894) );
  XNOR U1648 ( .A(n895), .B(n894), .Z(\w0[1][58] ) );
  XNOR U1649 ( .A(\w3[0][35] ), .B(n896), .Z(n897) );
  XOR U1650 ( .A(n898), .B(n897), .Z(\w0[1][59] ) );
  XOR U1651 ( .A(\w3[0][29] ), .B(n899), .Z(n900) );
  XOR U1652 ( .A(n901), .B(n900), .Z(\w0[1][5] ) );
  XOR U1653 ( .A(\w3[0][36] ), .B(n902), .Z(n903) );
  XOR U1654 ( .A(n904), .B(n903), .Z(\w0[1][60] ) );
  XOR U1655 ( .A(\w3[0][62] ), .B(\w3[0][54] ), .Z(n907) );
  XOR U1656 ( .A(\w3[0][37] ), .B(n905), .Z(n906) );
  XNOR U1657 ( .A(n907), .B(n906), .Z(\w0[1][61] ) );
  XOR U1658 ( .A(\w3[0][38] ), .B(n908), .Z(n909) );
  XOR U1659 ( .A(n910), .B(n909), .Z(\w0[1][62] ) );
  XNOR U1660 ( .A(n911), .B(\w3[0][39] ), .Z(n912) );
  XOR U1661 ( .A(n913), .B(n912), .Z(\w0[1][63] ) );
  XOR U1662 ( .A(\w3[0][65] ), .B(\w3[0][89] ), .Z(n954) );
  XNOR U1663 ( .A(\w3[0][80] ), .B(\w3[0][88] ), .Z(n995) );
  XOR U1664 ( .A(n995), .B(\w3[0][72] ), .Z(n914) );
  XNOR U1665 ( .A(n954), .B(n914), .Z(\w0[1][64] ) );
  XOR U1666 ( .A(\w3[0][66] ), .B(\w3[0][90] ), .Z(n955) );
  XOR U1667 ( .A(\w3[0][73] ), .B(\w3[0][81] ), .Z(n974) );
  XNOR U1668 ( .A(\w3[0][89] ), .B(n974), .Z(n915) );
  XNOR U1669 ( .A(n955), .B(n915), .Z(\w0[1][65] ) );
  XNOR U1670 ( .A(\w3[0][67] ), .B(\w3[0][91] ), .Z(n935) );
  XNOR U1671 ( .A(\w3[0][74] ), .B(\w3[0][82] ), .Z(n980) );
  XOR U1672 ( .A(\w3[0][90] ), .B(n980), .Z(n916) );
  XOR U1673 ( .A(n935), .B(n916), .Z(\w0[1][66] ) );
  XOR U1674 ( .A(\w3[0][68] ), .B(\w3[0][64] ), .Z(n937) );
  XNOR U1675 ( .A(\w3[0][75] ), .B(\w3[0][83] ), .Z(n957) );
  XOR U1676 ( .A(\w3[0][88] ), .B(n957), .Z(n917) );
  XNOR U1677 ( .A(\w3[0][92] ), .B(n917), .Z(n983) );
  XNOR U1678 ( .A(\w3[0][91] ), .B(n983), .Z(n918) );
  XNOR U1679 ( .A(n937), .B(n918), .Z(\w0[1][67] ) );
  XOR U1680 ( .A(\w3[0][64] ), .B(\w3[0][69] ), .Z(n941) );
  XOR U1681 ( .A(\w3[0][76] ), .B(\w3[0][84] ), .Z(n920) );
  XNOR U1682 ( .A(\w3[0][88] ), .B(\w3[0][93] ), .Z(n919) );
  XOR U1683 ( .A(n920), .B(n919), .Z(n986) );
  XOR U1684 ( .A(\w3[0][92] ), .B(n986), .Z(n921) );
  XNOR U1685 ( .A(n941), .B(n921), .Z(\w0[1][68] ) );
  XNOR U1686 ( .A(\w3[0][70] ), .B(\w3[0][94] ), .Z(n946) );
  IV U1687 ( .A(\w3[0][85] ), .Z(n960) );
  XOR U1688 ( .A(\w3[0][77] ), .B(n960), .Z(n989) );
  XOR U1689 ( .A(\w3[0][93] ), .B(n989), .Z(n922) );
  XOR U1690 ( .A(n946), .B(n922), .Z(\w0[1][69] ) );
  XOR U1691 ( .A(n923), .B(\w3[0][30] ), .Z(n924) );
  XOR U1692 ( .A(n925), .B(n924), .Z(\w0[1][6] ) );
  XOR U1693 ( .A(\w3[0][64] ), .B(\w3[0][71] ), .Z(n947) );
  XNOR U1694 ( .A(\w3[0][78] ), .B(\w3[0][86] ), .Z(n963) );
  XOR U1695 ( .A(\w3[0][88] ), .B(\w3[0][95] ), .Z(n927) );
  XOR U1696 ( .A(n963), .B(n927), .Z(n992) );
  XOR U1697 ( .A(\w3[0][94] ), .B(n992), .Z(n926) );
  XNOR U1698 ( .A(n947), .B(n926), .Z(\w0[1][70] ) );
  XOR U1699 ( .A(\w3[0][79] ), .B(\w3[0][87] ), .Z(n997) );
  XOR U1700 ( .A(\w3[0][64] ), .B(n927), .Z(n928) );
  XOR U1701 ( .A(n997), .B(n928), .Z(\w0[1][71] ) );
  XOR U1702 ( .A(\w3[0][73] ), .B(\w3[0][64] ), .Z(n930) );
  IV U1703 ( .A(\w3[0][65] ), .Z(n975) );
  XNOR U1704 ( .A(n995), .B(n975), .Z(n929) );
  XNOR U1705 ( .A(n930), .B(n929), .Z(\w0[1][72] ) );
  XOR U1706 ( .A(\w3[0][66] ), .B(\w3[0][74] ), .Z(n932) );
  XNOR U1707 ( .A(n954), .B(\w3[0][81] ), .Z(n931) );
  XNOR U1708 ( .A(n932), .B(n931), .Z(\w0[1][73] ) );
  XOR U1709 ( .A(\w3[0][67] ), .B(\w3[0][75] ), .Z(n934) );
  XNOR U1710 ( .A(n955), .B(\w3[0][82] ), .Z(n933) );
  XNOR U1711 ( .A(n934), .B(n933), .Z(\w0[1][74] ) );
  IV U1712 ( .A(\w3[0][72] ), .Z(n945) );
  XNOR U1713 ( .A(n945), .B(n935), .Z(n936) );
  XOR U1714 ( .A(\w3[0][76] ), .B(n936), .Z(n958) );
  XNOR U1715 ( .A(\w3[0][83] ), .B(n937), .Z(n938) );
  XOR U1716 ( .A(n958), .B(n938), .Z(\w0[1][75] ) );
  XOR U1717 ( .A(\w3[0][68] ), .B(\w3[0][77] ), .Z(n940) );
  XOR U1718 ( .A(n945), .B(\w3[0][92] ), .Z(n939) );
  XOR U1719 ( .A(n940), .B(n939), .Z(n961) );
  XNOR U1720 ( .A(\w3[0][84] ), .B(n941), .Z(n942) );
  XOR U1721 ( .A(n961), .B(n942), .Z(\w0[1][76] ) );
  XNOR U1722 ( .A(\w3[0][93] ), .B(\w3[0][69] ), .Z(n964) );
  XNOR U1723 ( .A(\w3[0][78] ), .B(n964), .Z(n944) );
  XOR U1724 ( .A(n960), .B(\w3[0][70] ), .Z(n943) );
  XNOR U1725 ( .A(n944), .B(n943), .Z(\w0[1][77] ) );
  XNOR U1726 ( .A(n945), .B(\w3[0][79] ), .Z(n969) );
  XOR U1727 ( .A(n946), .B(n969), .Z(n965) );
  XNOR U1728 ( .A(\w3[0][86] ), .B(n947), .Z(n948) );
  XOR U1729 ( .A(n965), .B(n948), .Z(\w0[1][78] ) );
  XOR U1730 ( .A(\w3[0][95] ), .B(\w3[0][71] ), .Z(n967) );
  XNOR U1731 ( .A(\w3[0][72] ), .B(\w3[0][64] ), .Z(n970) );
  XOR U1732 ( .A(\w3[0][87] ), .B(n970), .Z(n949) );
  XNOR U1733 ( .A(n967), .B(n949), .Z(\w0[1][79] ) );
  XNOR U1734 ( .A(\w3[0][0] ), .B(n950), .Z(n951) );
  XOR U1735 ( .A(n952), .B(n951), .Z(\w0[1][7] ) );
  XNOR U1736 ( .A(\w3[0][88] ), .B(n974), .Z(n953) );
  XOR U1737 ( .A(n970), .B(n953), .Z(\w0[1][80] ) );
  XNOR U1738 ( .A(n955), .B(\w3[0][74] ), .Z(n956) );
  XOR U1739 ( .A(n957), .B(n956), .Z(\w0[1][82] ) );
  IV U1740 ( .A(\w3[0][80] ), .Z(n971) );
  XOR U1741 ( .A(n971), .B(\w3[0][84] ), .Z(n985) );
  XOR U1742 ( .A(\w3[0][75] ), .B(n958), .Z(n959) );
  XOR U1743 ( .A(n985), .B(n959), .Z(\w0[1][83] ) );
  XOR U1744 ( .A(\w3[0][80] ), .B(n960), .Z(n988) );
  XOR U1745 ( .A(\w3[0][76] ), .B(n961), .Z(n962) );
  XOR U1746 ( .A(n988), .B(n962), .Z(\w0[1][84] ) );
  XOR U1747 ( .A(n971), .B(\w3[0][87] ), .Z(n994) );
  XOR U1748 ( .A(\w3[0][78] ), .B(n965), .Z(n966) );
  XOR U1749 ( .A(n994), .B(n966), .Z(\w0[1][86] ) );
  XOR U1750 ( .A(\w3[0][80] ), .B(n967), .Z(n968) );
  XOR U1751 ( .A(n969), .B(n968), .Z(\w0[1][87] ) );
  XNOR U1752 ( .A(\w3[0][81] ), .B(n970), .Z(n973) );
  XOR U1753 ( .A(n971), .B(\w3[0][89] ), .Z(n972) );
  XNOR U1754 ( .A(n973), .B(n972), .Z(\w0[1][88] ) );
  XOR U1755 ( .A(\w3[0][90] ), .B(\w3[0][82] ), .Z(n977) );
  XOR U1756 ( .A(n975), .B(n974), .Z(n976) );
  XNOR U1757 ( .A(n977), .B(n976), .Z(\w0[1][89] ) );
  XOR U1758 ( .A(\w3[0][91] ), .B(\w3[0][83] ), .Z(n982) );
  XOR U1759 ( .A(\w3[0][66] ), .B(n980), .Z(n981) );
  XNOR U1760 ( .A(n982), .B(n981), .Z(\w0[1][90] ) );
  XNOR U1761 ( .A(\w3[0][67] ), .B(n983), .Z(n984) );
  XOR U1762 ( .A(n985), .B(n984), .Z(\w0[1][91] ) );
  XOR U1763 ( .A(\w3[0][68] ), .B(n986), .Z(n987) );
  XOR U1764 ( .A(n988), .B(n987), .Z(\w0[1][92] ) );
  XOR U1765 ( .A(\w3[0][94] ), .B(\w3[0][86] ), .Z(n991) );
  XOR U1766 ( .A(\w3[0][69] ), .B(n989), .Z(n990) );
  XNOR U1767 ( .A(n991), .B(n990), .Z(\w0[1][93] ) );
  XOR U1768 ( .A(\w3[0][70] ), .B(n992), .Z(n993) );
  XOR U1769 ( .A(n994), .B(n993), .Z(\w0[1][94] ) );
  XNOR U1770 ( .A(n995), .B(\w3[0][71] ), .Z(n996) );
  XOR U1771 ( .A(n997), .B(n996), .Z(\w0[1][95] ) );
  XNOR U1772 ( .A(n999), .B(n998), .Z(n1000) );
  XNOR U1773 ( .A(\w3[0][104] ), .B(n1000), .Z(\w0[1][96] ) );
  XNOR U1774 ( .A(\w3[0][121] ), .B(n1001), .Z(n1002) );
  XNOR U1775 ( .A(n1003), .B(n1002), .Z(\w0[1][97] ) );
  XOR U1776 ( .A(\w3[0][122] ), .B(n1004), .Z(n1005) );
  XNOR U1777 ( .A(n1006), .B(n1005), .Z(\w0[1][98] ) );
  XOR U1778 ( .A(n1007), .B(\w3[0][123] ), .Z(n1008) );
  XNOR U1779 ( .A(n1009), .B(n1008), .Z(\w0[1][99] ) );
  XOR U1780 ( .A(\w3[0][17] ), .B(\w3[0][10] ), .Z(n1012) );
  XOR U1781 ( .A(n1010), .B(\w3[0][2] ), .Z(n1011) );
  XNOR U1782 ( .A(n1012), .B(n1011), .Z(\w0[1][9] ) );
  NANDN U1783 ( .A(n714), .B(state[0]), .Z(n1014) );
  NANDN U1784 ( .A(init), .B(msg[0]), .Z(n1013) );
  NAND U1785 ( .A(n1014), .B(n1013), .Z(n1015) );
  XOR U1786 ( .A(key[0]), .B(n1015), .Z(\w1[0][0] ) );
  NANDN U1787 ( .A(n714), .B(state[100]), .Z(n1017) );
  NANDN U1788 ( .A(init), .B(msg[100]), .Z(n1016) );
  NAND U1789 ( .A(n1017), .B(n1016), .Z(n1018) );
  XOR U1790 ( .A(key[100]), .B(n1018), .Z(\w1[0][100] ) );
  NANDN U1791 ( .A(n714), .B(state[101]), .Z(n1020) );
  NANDN U1792 ( .A(init), .B(msg[101]), .Z(n1019) );
  NAND U1793 ( .A(n1020), .B(n1019), .Z(n1021) );
  XOR U1794 ( .A(key[101]), .B(n1021), .Z(\w1[0][101] ) );
  NANDN U1795 ( .A(n714), .B(state[102]), .Z(n1023) );
  NANDN U1796 ( .A(init), .B(msg[102]), .Z(n1022) );
  NAND U1797 ( .A(n1023), .B(n1022), .Z(n1024) );
  XOR U1798 ( .A(key[102]), .B(n1024), .Z(\w1[0][102] ) );
  NANDN U1799 ( .A(n714), .B(state[103]), .Z(n1026) );
  NANDN U1800 ( .A(init), .B(msg[103]), .Z(n1025) );
  NAND U1801 ( .A(n1026), .B(n1025), .Z(n1027) );
  XOR U1802 ( .A(key[103]), .B(n1027), .Z(\w1[0][103] ) );
  NANDN U1803 ( .A(n714), .B(state[104]), .Z(n1029) );
  NANDN U1804 ( .A(init), .B(msg[104]), .Z(n1028) );
  NAND U1805 ( .A(n1029), .B(n1028), .Z(n1030) );
  XOR U1806 ( .A(key[104]), .B(n1030), .Z(\w1[0][104] ) );
  NANDN U1807 ( .A(n714), .B(state[105]), .Z(n1032) );
  NANDN U1808 ( .A(init), .B(msg[105]), .Z(n1031) );
  NAND U1809 ( .A(n1032), .B(n1031), .Z(n1033) );
  XOR U1810 ( .A(key[105]), .B(n1033), .Z(\w1[0][105] ) );
  NANDN U1811 ( .A(n714), .B(state[106]), .Z(n1035) );
  NANDN U1812 ( .A(init), .B(msg[106]), .Z(n1034) );
  NAND U1813 ( .A(n1035), .B(n1034), .Z(n1036) );
  XOR U1814 ( .A(key[106]), .B(n1036), .Z(\w1[0][106] ) );
  NANDN U1815 ( .A(n714), .B(state[107]), .Z(n1038) );
  NANDN U1816 ( .A(init), .B(msg[107]), .Z(n1037) );
  NAND U1817 ( .A(n1038), .B(n1037), .Z(n1039) );
  XOR U1818 ( .A(key[107]), .B(n1039), .Z(\w1[0][107] ) );
  NANDN U1819 ( .A(n714), .B(state[108]), .Z(n1041) );
  NANDN U1820 ( .A(init), .B(msg[108]), .Z(n1040) );
  NAND U1821 ( .A(n1041), .B(n1040), .Z(n1042) );
  XOR U1822 ( .A(key[108]), .B(n1042), .Z(\w1[0][108] ) );
  NANDN U1823 ( .A(n714), .B(state[109]), .Z(n1044) );
  NANDN U1824 ( .A(init), .B(msg[109]), .Z(n1043) );
  NAND U1825 ( .A(n1044), .B(n1043), .Z(n1045) );
  XOR U1826 ( .A(key[109]), .B(n1045), .Z(\w1[0][109] ) );
  NANDN U1827 ( .A(n714), .B(state[10]), .Z(n1047) );
  NANDN U1828 ( .A(init), .B(msg[10]), .Z(n1046) );
  NAND U1829 ( .A(n1047), .B(n1046), .Z(n1048) );
  XOR U1830 ( .A(key[10]), .B(n1048), .Z(\w1[0][10] ) );
  NANDN U1831 ( .A(n714), .B(state[110]), .Z(n1050) );
  NANDN U1832 ( .A(init), .B(msg[110]), .Z(n1049) );
  NAND U1833 ( .A(n1050), .B(n1049), .Z(n1051) );
  XOR U1834 ( .A(key[110]), .B(n1051), .Z(\w1[0][110] ) );
  NANDN U1835 ( .A(n714), .B(state[111]), .Z(n1053) );
  NANDN U1836 ( .A(init), .B(msg[111]), .Z(n1052) );
  NAND U1837 ( .A(n1053), .B(n1052), .Z(n1054) );
  XOR U1838 ( .A(key[111]), .B(n1054), .Z(\w1[0][111] ) );
  NANDN U1839 ( .A(n714), .B(state[112]), .Z(n1056) );
  NANDN U1840 ( .A(init), .B(msg[112]), .Z(n1055) );
  NAND U1841 ( .A(n1056), .B(n1055), .Z(n1057) );
  XOR U1842 ( .A(key[112]), .B(n1057), .Z(\w1[0][112] ) );
  NANDN U1843 ( .A(n714), .B(state[113]), .Z(n1059) );
  NANDN U1844 ( .A(init), .B(msg[113]), .Z(n1058) );
  NAND U1845 ( .A(n1059), .B(n1058), .Z(n1060) );
  XOR U1846 ( .A(key[113]), .B(n1060), .Z(\w1[0][113] ) );
  NANDN U1847 ( .A(n714), .B(state[114]), .Z(n1062) );
  NANDN U1848 ( .A(init), .B(msg[114]), .Z(n1061) );
  NAND U1849 ( .A(n1062), .B(n1061), .Z(n1063) );
  XOR U1850 ( .A(key[114]), .B(n1063), .Z(\w1[0][114] ) );
  NANDN U1851 ( .A(n714), .B(state[115]), .Z(n1065) );
  NANDN U1852 ( .A(init), .B(msg[115]), .Z(n1064) );
  NAND U1853 ( .A(n1065), .B(n1064), .Z(n1066) );
  XOR U1854 ( .A(key[115]), .B(n1066), .Z(\w1[0][115] ) );
  NANDN U1855 ( .A(n714), .B(state[116]), .Z(n1068) );
  NANDN U1856 ( .A(init), .B(msg[116]), .Z(n1067) );
  NAND U1857 ( .A(n1068), .B(n1067), .Z(n1069) );
  XOR U1858 ( .A(key[116]), .B(n1069), .Z(\w1[0][116] ) );
  NANDN U1859 ( .A(n714), .B(state[117]), .Z(n1071) );
  NANDN U1860 ( .A(init), .B(msg[117]), .Z(n1070) );
  NAND U1861 ( .A(n1071), .B(n1070), .Z(n1072) );
  XOR U1862 ( .A(key[117]), .B(n1072), .Z(\w1[0][117] ) );
  NANDN U1863 ( .A(n714), .B(state[118]), .Z(n1074) );
  NANDN U1864 ( .A(init), .B(msg[118]), .Z(n1073) );
  NAND U1865 ( .A(n1074), .B(n1073), .Z(n1075) );
  XOR U1866 ( .A(key[118]), .B(n1075), .Z(\w1[0][118] ) );
  NANDN U1867 ( .A(n714), .B(state[119]), .Z(n1077) );
  NANDN U1868 ( .A(init), .B(msg[119]), .Z(n1076) );
  NAND U1869 ( .A(n1077), .B(n1076), .Z(n1078) );
  XOR U1870 ( .A(key[119]), .B(n1078), .Z(\w1[0][119] ) );
  NANDN U1871 ( .A(n714), .B(state[11]), .Z(n1080) );
  NANDN U1872 ( .A(init), .B(msg[11]), .Z(n1079) );
  NAND U1873 ( .A(n1080), .B(n1079), .Z(n1081) );
  XOR U1874 ( .A(key[11]), .B(n1081), .Z(\w1[0][11] ) );
  NANDN U1875 ( .A(n714), .B(state[120]), .Z(n1083) );
  NANDN U1876 ( .A(init), .B(msg[120]), .Z(n1082) );
  NAND U1877 ( .A(n1083), .B(n1082), .Z(n1084) );
  XOR U1878 ( .A(key[120]), .B(n1084), .Z(\w1[0][120] ) );
  NANDN U1879 ( .A(n714), .B(state[121]), .Z(n1086) );
  NANDN U1880 ( .A(init), .B(msg[121]), .Z(n1085) );
  NAND U1881 ( .A(n1086), .B(n1085), .Z(n1087) );
  XOR U1882 ( .A(key[121]), .B(n1087), .Z(\w1[0][121] ) );
  NANDN U1883 ( .A(n714), .B(state[122]), .Z(n1089) );
  NANDN U1884 ( .A(init), .B(msg[122]), .Z(n1088) );
  NAND U1885 ( .A(n1089), .B(n1088), .Z(n1090) );
  XOR U1886 ( .A(key[122]), .B(n1090), .Z(\w1[0][122] ) );
  NANDN U1887 ( .A(n714), .B(state[123]), .Z(n1092) );
  NANDN U1888 ( .A(init), .B(msg[123]), .Z(n1091) );
  NAND U1889 ( .A(n1092), .B(n1091), .Z(n1093) );
  XOR U1890 ( .A(key[123]), .B(n1093), .Z(\w1[0][123] ) );
  NANDN U1891 ( .A(n714), .B(state[124]), .Z(n1095) );
  NANDN U1892 ( .A(init), .B(msg[124]), .Z(n1094) );
  NAND U1893 ( .A(n1095), .B(n1094), .Z(n1096) );
  XOR U1894 ( .A(key[124]), .B(n1096), .Z(\w1[0][124] ) );
  NANDN U1895 ( .A(n714), .B(state[125]), .Z(n1098) );
  NANDN U1896 ( .A(init), .B(msg[125]), .Z(n1097) );
  NAND U1897 ( .A(n1098), .B(n1097), .Z(n1099) );
  XOR U1898 ( .A(key[125]), .B(n1099), .Z(\w1[0][125] ) );
  NANDN U1899 ( .A(n714), .B(state[126]), .Z(n1101) );
  NANDN U1900 ( .A(init), .B(msg[126]), .Z(n1100) );
  NAND U1901 ( .A(n1101), .B(n1100), .Z(n1102) );
  XOR U1902 ( .A(key[126]), .B(n1102), .Z(\w1[0][126] ) );
  NANDN U1903 ( .A(n714), .B(state[127]), .Z(n1104) );
  NANDN U1904 ( .A(init), .B(msg[127]), .Z(n1103) );
  NAND U1905 ( .A(n1104), .B(n1103), .Z(n1105) );
  XOR U1906 ( .A(key[127]), .B(n1105), .Z(\w1[0][127] ) );
  NANDN U1907 ( .A(n714), .B(state[12]), .Z(n1107) );
  NANDN U1908 ( .A(init), .B(msg[12]), .Z(n1106) );
  NAND U1909 ( .A(n1107), .B(n1106), .Z(n1108) );
  XOR U1910 ( .A(key[12]), .B(n1108), .Z(\w1[0][12] ) );
  NANDN U1911 ( .A(n714), .B(state[13]), .Z(n1110) );
  NANDN U1912 ( .A(init), .B(msg[13]), .Z(n1109) );
  NAND U1913 ( .A(n1110), .B(n1109), .Z(n1111) );
  XOR U1914 ( .A(key[13]), .B(n1111), .Z(\w1[0][13] ) );
  NANDN U1915 ( .A(n714), .B(state[14]), .Z(n1113) );
  NANDN U1916 ( .A(init), .B(msg[14]), .Z(n1112) );
  NAND U1917 ( .A(n1113), .B(n1112), .Z(n1114) );
  XOR U1918 ( .A(key[14]), .B(n1114), .Z(\w1[0][14] ) );
  NANDN U1919 ( .A(n714), .B(state[15]), .Z(n1116) );
  NANDN U1920 ( .A(init), .B(msg[15]), .Z(n1115) );
  NAND U1921 ( .A(n1116), .B(n1115), .Z(n1117) );
  XOR U1922 ( .A(key[15]), .B(n1117), .Z(\w1[0][15] ) );
  NANDN U1923 ( .A(n714), .B(state[16]), .Z(n1119) );
  NANDN U1924 ( .A(init), .B(msg[16]), .Z(n1118) );
  NAND U1925 ( .A(n1119), .B(n1118), .Z(n1120) );
  XOR U1926 ( .A(key[16]), .B(n1120), .Z(\w1[0][16] ) );
  NANDN U1927 ( .A(n714), .B(state[17]), .Z(n1122) );
  NANDN U1928 ( .A(init), .B(msg[17]), .Z(n1121) );
  NAND U1929 ( .A(n1122), .B(n1121), .Z(n1123) );
  XOR U1930 ( .A(key[17]), .B(n1123), .Z(\w1[0][17] ) );
  NANDN U1931 ( .A(n714), .B(state[18]), .Z(n1125) );
  NANDN U1932 ( .A(init), .B(msg[18]), .Z(n1124) );
  NAND U1933 ( .A(n1125), .B(n1124), .Z(n1126) );
  XOR U1934 ( .A(key[18]), .B(n1126), .Z(\w1[0][18] ) );
  NANDN U1935 ( .A(n714), .B(state[19]), .Z(n1128) );
  NANDN U1936 ( .A(init), .B(msg[19]), .Z(n1127) );
  NAND U1937 ( .A(n1128), .B(n1127), .Z(n1129) );
  XOR U1938 ( .A(key[19]), .B(n1129), .Z(\w1[0][19] ) );
  NANDN U1939 ( .A(n714), .B(state[1]), .Z(n1131) );
  NANDN U1940 ( .A(init), .B(msg[1]), .Z(n1130) );
  NAND U1941 ( .A(n1131), .B(n1130), .Z(n1132) );
  XOR U1942 ( .A(key[1]), .B(n1132), .Z(\w1[0][1] ) );
  NANDN U1943 ( .A(n714), .B(state[20]), .Z(n1134) );
  NANDN U1944 ( .A(init), .B(msg[20]), .Z(n1133) );
  NAND U1945 ( .A(n1134), .B(n1133), .Z(n1135) );
  XOR U1946 ( .A(key[20]), .B(n1135), .Z(\w1[0][20] ) );
  NANDN U1947 ( .A(n714), .B(state[21]), .Z(n1137) );
  NANDN U1948 ( .A(init), .B(msg[21]), .Z(n1136) );
  NAND U1949 ( .A(n1137), .B(n1136), .Z(n1138) );
  XOR U1950 ( .A(key[21]), .B(n1138), .Z(\w1[0][21] ) );
  NANDN U1951 ( .A(n714), .B(state[22]), .Z(n1140) );
  NANDN U1952 ( .A(init), .B(msg[22]), .Z(n1139) );
  NAND U1953 ( .A(n1140), .B(n1139), .Z(n1141) );
  XOR U1954 ( .A(key[22]), .B(n1141), .Z(\w1[0][22] ) );
  NANDN U1955 ( .A(n714), .B(state[23]), .Z(n1143) );
  NANDN U1956 ( .A(init), .B(msg[23]), .Z(n1142) );
  NAND U1957 ( .A(n1143), .B(n1142), .Z(n1144) );
  XOR U1958 ( .A(key[23]), .B(n1144), .Z(\w1[0][23] ) );
  NANDN U1959 ( .A(n714), .B(state[24]), .Z(n1146) );
  NANDN U1960 ( .A(init), .B(msg[24]), .Z(n1145) );
  NAND U1961 ( .A(n1146), .B(n1145), .Z(n1147) );
  XOR U1962 ( .A(key[24]), .B(n1147), .Z(\w1[0][24] ) );
  NANDN U1963 ( .A(n714), .B(state[25]), .Z(n1149) );
  NANDN U1964 ( .A(init), .B(msg[25]), .Z(n1148) );
  NAND U1965 ( .A(n1149), .B(n1148), .Z(n1150) );
  XOR U1966 ( .A(key[25]), .B(n1150), .Z(\w1[0][25] ) );
  NANDN U1967 ( .A(n714), .B(state[26]), .Z(n1152) );
  NANDN U1968 ( .A(init), .B(msg[26]), .Z(n1151) );
  NAND U1969 ( .A(n1152), .B(n1151), .Z(n1153) );
  XOR U1970 ( .A(key[26]), .B(n1153), .Z(\w1[0][26] ) );
  NANDN U1971 ( .A(n714), .B(state[27]), .Z(n1155) );
  NANDN U1972 ( .A(init), .B(msg[27]), .Z(n1154) );
  NAND U1973 ( .A(n1155), .B(n1154), .Z(n1156) );
  XOR U1974 ( .A(key[27]), .B(n1156), .Z(\w1[0][27] ) );
  NANDN U1975 ( .A(n714), .B(state[28]), .Z(n1158) );
  NANDN U1976 ( .A(init), .B(msg[28]), .Z(n1157) );
  NAND U1977 ( .A(n1158), .B(n1157), .Z(n1159) );
  XOR U1978 ( .A(key[28]), .B(n1159), .Z(\w1[0][28] ) );
  NANDN U1979 ( .A(n714), .B(state[29]), .Z(n1161) );
  NANDN U1980 ( .A(init), .B(msg[29]), .Z(n1160) );
  NAND U1981 ( .A(n1161), .B(n1160), .Z(n1162) );
  XOR U1982 ( .A(key[29]), .B(n1162), .Z(\w1[0][29] ) );
  NANDN U1983 ( .A(n714), .B(state[2]), .Z(n1164) );
  NANDN U1984 ( .A(init), .B(msg[2]), .Z(n1163) );
  NAND U1985 ( .A(n1164), .B(n1163), .Z(n1165) );
  XOR U1986 ( .A(key[2]), .B(n1165), .Z(\w1[0][2] ) );
  NANDN U1987 ( .A(n714), .B(state[30]), .Z(n1167) );
  NANDN U1988 ( .A(init), .B(msg[30]), .Z(n1166) );
  NAND U1989 ( .A(n1167), .B(n1166), .Z(n1168) );
  XOR U1990 ( .A(key[30]), .B(n1168), .Z(\w1[0][30] ) );
  NANDN U1991 ( .A(n714), .B(state[31]), .Z(n1170) );
  NANDN U1992 ( .A(init), .B(msg[31]), .Z(n1169) );
  NAND U1993 ( .A(n1170), .B(n1169), .Z(n1171) );
  XOR U1994 ( .A(key[31]), .B(n1171), .Z(\w1[0][31] ) );
  NANDN U1995 ( .A(n714), .B(state[32]), .Z(n1173) );
  NANDN U1996 ( .A(init), .B(msg[32]), .Z(n1172) );
  NAND U1997 ( .A(n1173), .B(n1172), .Z(n1174) );
  XOR U1998 ( .A(key[32]), .B(n1174), .Z(\w1[0][32] ) );
  NANDN U1999 ( .A(n714), .B(state[33]), .Z(n1176) );
  NANDN U2000 ( .A(init), .B(msg[33]), .Z(n1175) );
  NAND U2001 ( .A(n1176), .B(n1175), .Z(n1177) );
  XOR U2002 ( .A(key[33]), .B(n1177), .Z(\w1[0][33] ) );
  NANDN U2003 ( .A(n714), .B(state[34]), .Z(n1179) );
  NANDN U2004 ( .A(init), .B(msg[34]), .Z(n1178) );
  NAND U2005 ( .A(n1179), .B(n1178), .Z(n1180) );
  XOR U2006 ( .A(key[34]), .B(n1180), .Z(\w1[0][34] ) );
  NANDN U2007 ( .A(n714), .B(state[35]), .Z(n1182) );
  NANDN U2008 ( .A(init), .B(msg[35]), .Z(n1181) );
  NAND U2009 ( .A(n1182), .B(n1181), .Z(n1183) );
  XOR U2010 ( .A(key[35]), .B(n1183), .Z(\w1[0][35] ) );
  NANDN U2011 ( .A(n714), .B(state[36]), .Z(n1185) );
  NANDN U2012 ( .A(init), .B(msg[36]), .Z(n1184) );
  NAND U2013 ( .A(n1185), .B(n1184), .Z(n1186) );
  XOR U2014 ( .A(key[36]), .B(n1186), .Z(\w1[0][36] ) );
  NANDN U2015 ( .A(n714), .B(state[37]), .Z(n1188) );
  NANDN U2016 ( .A(init), .B(msg[37]), .Z(n1187) );
  NAND U2017 ( .A(n1188), .B(n1187), .Z(n1189) );
  XOR U2018 ( .A(key[37]), .B(n1189), .Z(\w1[0][37] ) );
  NANDN U2019 ( .A(n714), .B(state[38]), .Z(n1191) );
  NANDN U2020 ( .A(init), .B(msg[38]), .Z(n1190) );
  NAND U2021 ( .A(n1191), .B(n1190), .Z(n1192) );
  XOR U2022 ( .A(key[38]), .B(n1192), .Z(\w1[0][38] ) );
  NANDN U2023 ( .A(n714), .B(state[39]), .Z(n1194) );
  NANDN U2024 ( .A(init), .B(msg[39]), .Z(n1193) );
  NAND U2025 ( .A(n1194), .B(n1193), .Z(n1195) );
  XOR U2026 ( .A(key[39]), .B(n1195), .Z(\w1[0][39] ) );
  NANDN U2027 ( .A(n714), .B(state[3]), .Z(n1197) );
  NANDN U2028 ( .A(init), .B(msg[3]), .Z(n1196) );
  NAND U2029 ( .A(n1197), .B(n1196), .Z(n1198) );
  XOR U2030 ( .A(key[3]), .B(n1198), .Z(\w1[0][3] ) );
  NANDN U2031 ( .A(n714), .B(state[40]), .Z(n1200) );
  NANDN U2032 ( .A(init), .B(msg[40]), .Z(n1199) );
  NAND U2033 ( .A(n1200), .B(n1199), .Z(n1201) );
  XOR U2034 ( .A(key[40]), .B(n1201), .Z(\w1[0][40] ) );
  NANDN U2035 ( .A(n714), .B(state[41]), .Z(n1203) );
  NANDN U2036 ( .A(init), .B(msg[41]), .Z(n1202) );
  NAND U2037 ( .A(n1203), .B(n1202), .Z(n1204) );
  XOR U2038 ( .A(key[41]), .B(n1204), .Z(\w1[0][41] ) );
  NANDN U2039 ( .A(n714), .B(state[42]), .Z(n1206) );
  NANDN U2040 ( .A(init), .B(msg[42]), .Z(n1205) );
  NAND U2041 ( .A(n1206), .B(n1205), .Z(n1207) );
  XOR U2042 ( .A(key[42]), .B(n1207), .Z(\w1[0][42] ) );
  NANDN U2043 ( .A(n714), .B(state[43]), .Z(n1209) );
  NANDN U2044 ( .A(init), .B(msg[43]), .Z(n1208) );
  NAND U2045 ( .A(n1209), .B(n1208), .Z(n1210) );
  XOR U2046 ( .A(key[43]), .B(n1210), .Z(\w1[0][43] ) );
  NANDN U2047 ( .A(n714), .B(state[44]), .Z(n1212) );
  NANDN U2048 ( .A(init), .B(msg[44]), .Z(n1211) );
  NAND U2049 ( .A(n1212), .B(n1211), .Z(n1213) );
  XOR U2050 ( .A(key[44]), .B(n1213), .Z(\w1[0][44] ) );
  NANDN U2051 ( .A(n714), .B(state[45]), .Z(n1215) );
  NANDN U2052 ( .A(init), .B(msg[45]), .Z(n1214) );
  NAND U2053 ( .A(n1215), .B(n1214), .Z(n1216) );
  XOR U2054 ( .A(key[45]), .B(n1216), .Z(\w1[0][45] ) );
  NANDN U2055 ( .A(n714), .B(state[46]), .Z(n1218) );
  NANDN U2056 ( .A(init), .B(msg[46]), .Z(n1217) );
  NAND U2057 ( .A(n1218), .B(n1217), .Z(n1219) );
  XOR U2058 ( .A(key[46]), .B(n1219), .Z(\w1[0][46] ) );
  NANDN U2059 ( .A(n714), .B(state[47]), .Z(n1221) );
  NANDN U2060 ( .A(init), .B(msg[47]), .Z(n1220) );
  NAND U2061 ( .A(n1221), .B(n1220), .Z(n1222) );
  XOR U2062 ( .A(key[47]), .B(n1222), .Z(\w1[0][47] ) );
  NANDN U2063 ( .A(n714), .B(state[48]), .Z(n1224) );
  NANDN U2064 ( .A(init), .B(msg[48]), .Z(n1223) );
  NAND U2065 ( .A(n1224), .B(n1223), .Z(n1225) );
  XOR U2066 ( .A(key[48]), .B(n1225), .Z(\w1[0][48] ) );
  NANDN U2067 ( .A(n714), .B(state[49]), .Z(n1227) );
  NANDN U2068 ( .A(init), .B(msg[49]), .Z(n1226) );
  NAND U2069 ( .A(n1227), .B(n1226), .Z(n1228) );
  XOR U2070 ( .A(key[49]), .B(n1228), .Z(\w1[0][49] ) );
  NANDN U2071 ( .A(n714), .B(state[4]), .Z(n1230) );
  NANDN U2072 ( .A(init), .B(msg[4]), .Z(n1229) );
  NAND U2073 ( .A(n1230), .B(n1229), .Z(n1231) );
  XOR U2074 ( .A(key[4]), .B(n1231), .Z(\w1[0][4] ) );
  NANDN U2075 ( .A(n714), .B(state[50]), .Z(n1233) );
  NANDN U2076 ( .A(init), .B(msg[50]), .Z(n1232) );
  NAND U2077 ( .A(n1233), .B(n1232), .Z(n1234) );
  XOR U2078 ( .A(key[50]), .B(n1234), .Z(\w1[0][50] ) );
  NANDN U2079 ( .A(n714), .B(state[51]), .Z(n1236) );
  NANDN U2080 ( .A(init), .B(msg[51]), .Z(n1235) );
  NAND U2081 ( .A(n1236), .B(n1235), .Z(n1237) );
  XOR U2082 ( .A(key[51]), .B(n1237), .Z(\w1[0][51] ) );
  NANDN U2083 ( .A(n714), .B(state[52]), .Z(n1239) );
  NANDN U2084 ( .A(init), .B(msg[52]), .Z(n1238) );
  NAND U2085 ( .A(n1239), .B(n1238), .Z(n1240) );
  XOR U2086 ( .A(key[52]), .B(n1240), .Z(\w1[0][52] ) );
  NANDN U2087 ( .A(n714), .B(state[53]), .Z(n1242) );
  NANDN U2088 ( .A(init), .B(msg[53]), .Z(n1241) );
  NAND U2089 ( .A(n1242), .B(n1241), .Z(n1243) );
  XOR U2090 ( .A(key[53]), .B(n1243), .Z(\w1[0][53] ) );
  NANDN U2091 ( .A(n714), .B(state[54]), .Z(n1245) );
  NANDN U2092 ( .A(init), .B(msg[54]), .Z(n1244) );
  NAND U2093 ( .A(n1245), .B(n1244), .Z(n1246) );
  XOR U2094 ( .A(key[54]), .B(n1246), .Z(\w1[0][54] ) );
  NANDN U2095 ( .A(n714), .B(state[55]), .Z(n1248) );
  NANDN U2096 ( .A(init), .B(msg[55]), .Z(n1247) );
  NAND U2097 ( .A(n1248), .B(n1247), .Z(n1249) );
  XOR U2098 ( .A(key[55]), .B(n1249), .Z(\w1[0][55] ) );
  NANDN U2099 ( .A(n714), .B(state[56]), .Z(n1251) );
  NANDN U2100 ( .A(init), .B(msg[56]), .Z(n1250) );
  NAND U2101 ( .A(n1251), .B(n1250), .Z(n1252) );
  XOR U2102 ( .A(key[56]), .B(n1252), .Z(\w1[0][56] ) );
  NANDN U2103 ( .A(n714), .B(state[57]), .Z(n1254) );
  NANDN U2104 ( .A(init), .B(msg[57]), .Z(n1253) );
  NAND U2105 ( .A(n1254), .B(n1253), .Z(n1255) );
  XOR U2106 ( .A(key[57]), .B(n1255), .Z(\w1[0][57] ) );
  NANDN U2107 ( .A(n714), .B(state[58]), .Z(n1257) );
  NANDN U2108 ( .A(init), .B(msg[58]), .Z(n1256) );
  NAND U2109 ( .A(n1257), .B(n1256), .Z(n1258) );
  XOR U2110 ( .A(key[58]), .B(n1258), .Z(\w1[0][58] ) );
  NANDN U2111 ( .A(n714), .B(state[59]), .Z(n1260) );
  NANDN U2112 ( .A(init), .B(msg[59]), .Z(n1259) );
  NAND U2113 ( .A(n1260), .B(n1259), .Z(n1261) );
  XOR U2114 ( .A(key[59]), .B(n1261), .Z(\w1[0][59] ) );
  NANDN U2115 ( .A(n714), .B(state[5]), .Z(n1263) );
  NANDN U2116 ( .A(init), .B(msg[5]), .Z(n1262) );
  NAND U2117 ( .A(n1263), .B(n1262), .Z(n1264) );
  XOR U2118 ( .A(key[5]), .B(n1264), .Z(\w1[0][5] ) );
  NANDN U2119 ( .A(n714), .B(state[60]), .Z(n1266) );
  NANDN U2120 ( .A(init), .B(msg[60]), .Z(n1265) );
  NAND U2121 ( .A(n1266), .B(n1265), .Z(n1267) );
  XOR U2122 ( .A(key[60]), .B(n1267), .Z(\w1[0][60] ) );
  NANDN U2123 ( .A(n714), .B(state[61]), .Z(n1269) );
  NANDN U2124 ( .A(init), .B(msg[61]), .Z(n1268) );
  NAND U2125 ( .A(n1269), .B(n1268), .Z(n1270) );
  XOR U2126 ( .A(key[61]), .B(n1270), .Z(\w1[0][61] ) );
  NANDN U2127 ( .A(n714), .B(state[62]), .Z(n1272) );
  NANDN U2128 ( .A(init), .B(msg[62]), .Z(n1271) );
  NAND U2129 ( .A(n1272), .B(n1271), .Z(n1273) );
  XOR U2130 ( .A(key[62]), .B(n1273), .Z(\w1[0][62] ) );
  NANDN U2131 ( .A(n714), .B(state[63]), .Z(n1275) );
  NANDN U2132 ( .A(init), .B(msg[63]), .Z(n1274) );
  NAND U2133 ( .A(n1275), .B(n1274), .Z(n1276) );
  XOR U2134 ( .A(key[63]), .B(n1276), .Z(\w1[0][63] ) );
  NANDN U2135 ( .A(n714), .B(state[64]), .Z(n1278) );
  NANDN U2136 ( .A(init), .B(msg[64]), .Z(n1277) );
  NAND U2137 ( .A(n1278), .B(n1277), .Z(n1279) );
  XOR U2138 ( .A(key[64]), .B(n1279), .Z(\w1[0][64] ) );
  NANDN U2139 ( .A(n714), .B(state[65]), .Z(n1281) );
  NANDN U2140 ( .A(init), .B(msg[65]), .Z(n1280) );
  NAND U2141 ( .A(n1281), .B(n1280), .Z(n1282) );
  XOR U2142 ( .A(key[65]), .B(n1282), .Z(\w1[0][65] ) );
  NANDN U2143 ( .A(n714), .B(state[66]), .Z(n1284) );
  NANDN U2144 ( .A(init), .B(msg[66]), .Z(n1283) );
  NAND U2145 ( .A(n1284), .B(n1283), .Z(n1285) );
  XOR U2146 ( .A(key[66]), .B(n1285), .Z(\w1[0][66] ) );
  NANDN U2147 ( .A(n714), .B(state[67]), .Z(n1287) );
  NANDN U2148 ( .A(init), .B(msg[67]), .Z(n1286) );
  NAND U2149 ( .A(n1287), .B(n1286), .Z(n1288) );
  XOR U2150 ( .A(key[67]), .B(n1288), .Z(\w1[0][67] ) );
  NANDN U2151 ( .A(n714), .B(state[68]), .Z(n1290) );
  NANDN U2152 ( .A(init), .B(msg[68]), .Z(n1289) );
  NAND U2153 ( .A(n1290), .B(n1289), .Z(n1291) );
  XOR U2154 ( .A(key[68]), .B(n1291), .Z(\w1[0][68] ) );
  NANDN U2155 ( .A(n714), .B(state[69]), .Z(n1293) );
  NANDN U2156 ( .A(init), .B(msg[69]), .Z(n1292) );
  NAND U2157 ( .A(n1293), .B(n1292), .Z(n1294) );
  XOR U2158 ( .A(key[69]), .B(n1294), .Z(\w1[0][69] ) );
  NANDN U2159 ( .A(n714), .B(state[6]), .Z(n1296) );
  NANDN U2160 ( .A(init), .B(msg[6]), .Z(n1295) );
  NAND U2161 ( .A(n1296), .B(n1295), .Z(n1297) );
  XOR U2162 ( .A(key[6]), .B(n1297), .Z(\w1[0][6] ) );
  NANDN U2163 ( .A(n714), .B(state[70]), .Z(n1299) );
  NANDN U2164 ( .A(init), .B(msg[70]), .Z(n1298) );
  NAND U2165 ( .A(n1299), .B(n1298), .Z(n1300) );
  XOR U2166 ( .A(key[70]), .B(n1300), .Z(\w1[0][70] ) );
  NANDN U2167 ( .A(n714), .B(state[71]), .Z(n1302) );
  NANDN U2168 ( .A(init), .B(msg[71]), .Z(n1301) );
  NAND U2169 ( .A(n1302), .B(n1301), .Z(n1303) );
  XOR U2170 ( .A(key[71]), .B(n1303), .Z(\w1[0][71] ) );
  NANDN U2171 ( .A(n714), .B(state[72]), .Z(n1305) );
  NANDN U2172 ( .A(init), .B(msg[72]), .Z(n1304) );
  NAND U2173 ( .A(n1305), .B(n1304), .Z(n1306) );
  XOR U2174 ( .A(key[72]), .B(n1306), .Z(\w1[0][72] ) );
  NANDN U2175 ( .A(n714), .B(state[73]), .Z(n1308) );
  NANDN U2176 ( .A(init), .B(msg[73]), .Z(n1307) );
  NAND U2177 ( .A(n1308), .B(n1307), .Z(n1309) );
  XOR U2178 ( .A(key[73]), .B(n1309), .Z(\w1[0][73] ) );
  NANDN U2179 ( .A(n714), .B(state[74]), .Z(n1311) );
  NANDN U2180 ( .A(init), .B(msg[74]), .Z(n1310) );
  NAND U2181 ( .A(n1311), .B(n1310), .Z(n1312) );
  XOR U2182 ( .A(key[74]), .B(n1312), .Z(\w1[0][74] ) );
  NANDN U2183 ( .A(n714), .B(state[75]), .Z(n1314) );
  NANDN U2184 ( .A(init), .B(msg[75]), .Z(n1313) );
  NAND U2185 ( .A(n1314), .B(n1313), .Z(n1315) );
  XOR U2186 ( .A(key[75]), .B(n1315), .Z(\w1[0][75] ) );
  NANDN U2187 ( .A(n714), .B(state[76]), .Z(n1317) );
  NANDN U2188 ( .A(init), .B(msg[76]), .Z(n1316) );
  NAND U2189 ( .A(n1317), .B(n1316), .Z(n1318) );
  XOR U2190 ( .A(key[76]), .B(n1318), .Z(\w1[0][76] ) );
  NANDN U2191 ( .A(n714), .B(state[77]), .Z(n1320) );
  NANDN U2192 ( .A(init), .B(msg[77]), .Z(n1319) );
  NAND U2193 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U2194 ( .A(key[77]), .B(n1321), .Z(\w1[0][77] ) );
  NANDN U2195 ( .A(n714), .B(state[78]), .Z(n1323) );
  NANDN U2196 ( .A(init), .B(msg[78]), .Z(n1322) );
  NAND U2197 ( .A(n1323), .B(n1322), .Z(n1324) );
  XOR U2198 ( .A(key[78]), .B(n1324), .Z(\w1[0][78] ) );
  NANDN U2199 ( .A(n714), .B(state[79]), .Z(n1326) );
  NANDN U2200 ( .A(init), .B(msg[79]), .Z(n1325) );
  NAND U2201 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U2202 ( .A(key[79]), .B(n1327), .Z(\w1[0][79] ) );
  NANDN U2203 ( .A(n714), .B(state[7]), .Z(n1329) );
  NANDN U2204 ( .A(init), .B(msg[7]), .Z(n1328) );
  NAND U2205 ( .A(n1329), .B(n1328), .Z(n1330) );
  XOR U2206 ( .A(key[7]), .B(n1330), .Z(\w1[0][7] ) );
  NANDN U2207 ( .A(n714), .B(state[80]), .Z(n1332) );
  NANDN U2208 ( .A(init), .B(msg[80]), .Z(n1331) );
  NAND U2209 ( .A(n1332), .B(n1331), .Z(n1333) );
  XOR U2210 ( .A(key[80]), .B(n1333), .Z(\w1[0][80] ) );
  NANDN U2211 ( .A(n714), .B(state[81]), .Z(n1335) );
  NANDN U2212 ( .A(init), .B(msg[81]), .Z(n1334) );
  NAND U2213 ( .A(n1335), .B(n1334), .Z(n1336) );
  XOR U2214 ( .A(key[81]), .B(n1336), .Z(\w1[0][81] ) );
  NANDN U2215 ( .A(n714), .B(state[82]), .Z(n1338) );
  NANDN U2216 ( .A(init), .B(msg[82]), .Z(n1337) );
  NAND U2217 ( .A(n1338), .B(n1337), .Z(n1339) );
  XOR U2218 ( .A(key[82]), .B(n1339), .Z(\w1[0][82] ) );
  NANDN U2219 ( .A(n714), .B(state[83]), .Z(n1341) );
  NANDN U2220 ( .A(init), .B(msg[83]), .Z(n1340) );
  NAND U2221 ( .A(n1341), .B(n1340), .Z(n1342) );
  XOR U2222 ( .A(key[83]), .B(n1342), .Z(\w1[0][83] ) );
  NANDN U2223 ( .A(n714), .B(state[84]), .Z(n1344) );
  NANDN U2224 ( .A(init), .B(msg[84]), .Z(n1343) );
  NAND U2225 ( .A(n1344), .B(n1343), .Z(n1345) );
  XOR U2226 ( .A(key[84]), .B(n1345), .Z(\w1[0][84] ) );
  NANDN U2227 ( .A(n714), .B(state[85]), .Z(n1347) );
  NANDN U2228 ( .A(init), .B(msg[85]), .Z(n1346) );
  NAND U2229 ( .A(n1347), .B(n1346), .Z(n1348) );
  XOR U2230 ( .A(key[85]), .B(n1348), .Z(\w1[0][85] ) );
  NANDN U2231 ( .A(n714), .B(state[86]), .Z(n1350) );
  NANDN U2232 ( .A(init), .B(msg[86]), .Z(n1349) );
  NAND U2233 ( .A(n1350), .B(n1349), .Z(n1351) );
  XOR U2234 ( .A(key[86]), .B(n1351), .Z(\w1[0][86] ) );
  NANDN U2235 ( .A(n714), .B(state[87]), .Z(n1353) );
  NANDN U2236 ( .A(init), .B(msg[87]), .Z(n1352) );
  NAND U2237 ( .A(n1353), .B(n1352), .Z(n1354) );
  XOR U2238 ( .A(key[87]), .B(n1354), .Z(\w1[0][87] ) );
  NANDN U2239 ( .A(n714), .B(state[88]), .Z(n1356) );
  NANDN U2240 ( .A(init), .B(msg[88]), .Z(n1355) );
  NAND U2241 ( .A(n1356), .B(n1355), .Z(n1357) );
  XOR U2242 ( .A(key[88]), .B(n1357), .Z(\w1[0][88] ) );
  NANDN U2243 ( .A(n714), .B(state[89]), .Z(n1359) );
  NANDN U2244 ( .A(init), .B(msg[89]), .Z(n1358) );
  NAND U2245 ( .A(n1359), .B(n1358), .Z(n1360) );
  XOR U2246 ( .A(key[89]), .B(n1360), .Z(\w1[0][89] ) );
  NANDN U2247 ( .A(n714), .B(state[8]), .Z(n1362) );
  NANDN U2248 ( .A(init), .B(msg[8]), .Z(n1361) );
  NAND U2249 ( .A(n1362), .B(n1361), .Z(n1363) );
  XOR U2250 ( .A(key[8]), .B(n1363), .Z(\w1[0][8] ) );
  NANDN U2251 ( .A(n714), .B(state[90]), .Z(n1365) );
  NANDN U2252 ( .A(init), .B(msg[90]), .Z(n1364) );
  NAND U2253 ( .A(n1365), .B(n1364), .Z(n1366) );
  XOR U2254 ( .A(key[90]), .B(n1366), .Z(\w1[0][90] ) );
  NANDN U2255 ( .A(n714), .B(state[91]), .Z(n1368) );
  NANDN U2256 ( .A(init), .B(msg[91]), .Z(n1367) );
  NAND U2257 ( .A(n1368), .B(n1367), .Z(n1369) );
  XOR U2258 ( .A(key[91]), .B(n1369), .Z(\w1[0][91] ) );
  NANDN U2259 ( .A(n714), .B(state[92]), .Z(n1371) );
  NANDN U2260 ( .A(init), .B(msg[92]), .Z(n1370) );
  NAND U2261 ( .A(n1371), .B(n1370), .Z(n1372) );
  XOR U2262 ( .A(key[92]), .B(n1372), .Z(\w1[0][92] ) );
  NANDN U2263 ( .A(n714), .B(state[93]), .Z(n1374) );
  NANDN U2264 ( .A(init), .B(msg[93]), .Z(n1373) );
  NAND U2265 ( .A(n1374), .B(n1373), .Z(n1375) );
  XOR U2266 ( .A(key[93]), .B(n1375), .Z(\w1[0][93] ) );
  NANDN U2267 ( .A(n714), .B(state[94]), .Z(n1377) );
  NANDN U2268 ( .A(init), .B(msg[94]), .Z(n1376) );
  NAND U2269 ( .A(n1377), .B(n1376), .Z(n1378) );
  XOR U2270 ( .A(key[94]), .B(n1378), .Z(\w1[0][94] ) );
  NANDN U2271 ( .A(n714), .B(state[95]), .Z(n1380) );
  NANDN U2272 ( .A(init), .B(msg[95]), .Z(n1379) );
  NAND U2273 ( .A(n1380), .B(n1379), .Z(n1381) );
  XOR U2274 ( .A(key[95]), .B(n1381), .Z(\w1[0][95] ) );
  NANDN U2275 ( .A(n714), .B(state[96]), .Z(n1383) );
  NANDN U2276 ( .A(init), .B(msg[96]), .Z(n1382) );
  NAND U2277 ( .A(n1383), .B(n1382), .Z(n1384) );
  XOR U2278 ( .A(key[96]), .B(n1384), .Z(\w1[0][96] ) );
  NANDN U2279 ( .A(n714), .B(state[97]), .Z(n1386) );
  NANDN U2280 ( .A(init), .B(msg[97]), .Z(n1385) );
  NAND U2281 ( .A(n1386), .B(n1385), .Z(n1387) );
  XOR U2282 ( .A(key[97]), .B(n1387), .Z(\w1[0][97] ) );
  NANDN U2283 ( .A(n714), .B(state[98]), .Z(n1389) );
  NANDN U2284 ( .A(init), .B(msg[98]), .Z(n1388) );
  NAND U2285 ( .A(n1389), .B(n1388), .Z(n1390) );
  XOR U2286 ( .A(key[98]), .B(n1390), .Z(\w1[0][98] ) );
  NANDN U2287 ( .A(n714), .B(state[99]), .Z(n1392) );
  NANDN U2288 ( .A(init), .B(msg[99]), .Z(n1391) );
  NAND U2289 ( .A(n1392), .B(n1391), .Z(n1393) );
  XOR U2290 ( .A(key[99]), .B(n1393), .Z(\w1[0][99] ) );
  NANDN U2291 ( .A(n714), .B(state[9]), .Z(n1395) );
  NANDN U2292 ( .A(init), .B(msg[9]), .Z(n1394) );
  NAND U2293 ( .A(n1395), .B(n1394), .Z(n1396) );
  XOR U2294 ( .A(key[9]), .B(n1396), .Z(\w1[0][9] ) );
  XOR U2295 ( .A(key[128]), .B(\w0[1][0] ), .Z(\w1[1][0] ) );
  XOR U2296 ( .A(key[228]), .B(\w0[1][100] ), .Z(\w1[1][100] ) );
  XOR U2297 ( .A(key[229]), .B(\w0[1][101] ), .Z(\w1[1][101] ) );
  XOR U2298 ( .A(key[230]), .B(\w0[1][102] ), .Z(\w1[1][102] ) );
  XOR U2299 ( .A(key[231]), .B(\w0[1][103] ), .Z(\w1[1][103] ) );
  XOR U2300 ( .A(key[232]), .B(\w0[1][104] ), .Z(\w1[1][104] ) );
  XOR U2301 ( .A(key[233]), .B(\w0[1][105] ), .Z(\w1[1][105] ) );
  XOR U2302 ( .A(key[234]), .B(\w0[1][106] ), .Z(\w1[1][106] ) );
  XOR U2303 ( .A(key[235]), .B(\w0[1][107] ), .Z(\w1[1][107] ) );
  XOR U2304 ( .A(key[236]), .B(\w0[1][108] ), .Z(\w1[1][108] ) );
  XOR U2305 ( .A(key[237]), .B(\w0[1][109] ), .Z(\w1[1][109] ) );
  XOR U2306 ( .A(key[138]), .B(\w0[1][10] ), .Z(\w1[1][10] ) );
  XOR U2307 ( .A(key[238]), .B(\w0[1][110] ), .Z(\w1[1][110] ) );
  XOR U2308 ( .A(key[239]), .B(\w0[1][111] ), .Z(\w1[1][111] ) );
  XOR U2309 ( .A(key[240]), .B(\w0[1][112] ), .Z(\w1[1][112] ) );
  XOR U2310 ( .A(key[241]), .B(\w0[1][113] ), .Z(\w1[1][113] ) );
  XOR U2311 ( .A(key[242]), .B(\w0[1][114] ), .Z(\w1[1][114] ) );
  XOR U2312 ( .A(key[243]), .B(\w0[1][115] ), .Z(\w1[1][115] ) );
  XOR U2313 ( .A(key[244]), .B(\w0[1][116] ), .Z(\w1[1][116] ) );
  XOR U2314 ( .A(key[245]), .B(\w0[1][117] ), .Z(\w1[1][117] ) );
  XOR U2315 ( .A(key[246]), .B(\w0[1][118] ), .Z(\w1[1][118] ) );
  XOR U2316 ( .A(key[247]), .B(\w0[1][119] ), .Z(\w1[1][119] ) );
  XOR U2317 ( .A(key[139]), .B(\w0[1][11] ), .Z(\w1[1][11] ) );
  XOR U2318 ( .A(key[248]), .B(\w0[1][120] ), .Z(\w1[1][120] ) );
  XOR U2319 ( .A(key[249]), .B(\w0[1][121] ), .Z(\w1[1][121] ) );
  XOR U2320 ( .A(key[250]), .B(\w0[1][122] ), .Z(\w1[1][122] ) );
  XOR U2321 ( .A(key[251]), .B(\w0[1][123] ), .Z(\w1[1][123] ) );
  XOR U2322 ( .A(key[252]), .B(\w0[1][124] ), .Z(\w1[1][124] ) );
  XOR U2323 ( .A(key[253]), .B(\w0[1][125] ), .Z(\w1[1][125] ) );
  XOR U2324 ( .A(key[254]), .B(\w0[1][126] ), .Z(\w1[1][126] ) );
  XOR U2325 ( .A(key[255]), .B(\w0[1][127] ), .Z(\w1[1][127] ) );
  XOR U2326 ( .A(key[140]), .B(\w0[1][12] ), .Z(\w1[1][12] ) );
  XOR U2327 ( .A(key[141]), .B(\w0[1][13] ), .Z(\w1[1][13] ) );
  XOR U2328 ( .A(key[142]), .B(\w0[1][14] ), .Z(\w1[1][14] ) );
  XOR U2329 ( .A(key[143]), .B(\w0[1][15] ), .Z(\w1[1][15] ) );
  XOR U2330 ( .A(key[144]), .B(\w0[1][16] ), .Z(\w1[1][16] ) );
  XOR U2331 ( .A(key[145]), .B(\w0[1][17] ), .Z(\w1[1][17] ) );
  XOR U2332 ( .A(key[146]), .B(\w0[1][18] ), .Z(\w1[1][18] ) );
  XOR U2333 ( .A(key[147]), .B(\w0[1][19] ), .Z(\w1[1][19] ) );
  XOR U2334 ( .A(key[129]), .B(\w0[1][1] ), .Z(\w1[1][1] ) );
  XOR U2335 ( .A(key[148]), .B(\w0[1][20] ), .Z(\w1[1][20] ) );
  XOR U2336 ( .A(key[149]), .B(\w0[1][21] ), .Z(\w1[1][21] ) );
  XOR U2337 ( .A(key[150]), .B(\w0[1][22] ), .Z(\w1[1][22] ) );
  XOR U2338 ( .A(key[151]), .B(\w0[1][23] ), .Z(\w1[1][23] ) );
  XOR U2339 ( .A(key[152]), .B(\w0[1][24] ), .Z(\w1[1][24] ) );
  XOR U2340 ( .A(key[153]), .B(\w0[1][25] ), .Z(\w1[1][25] ) );
  XOR U2341 ( .A(key[154]), .B(\w0[1][26] ), .Z(\w1[1][26] ) );
  XOR U2342 ( .A(key[155]), .B(\w0[1][27] ), .Z(\w1[1][27] ) );
  XOR U2343 ( .A(key[156]), .B(\w0[1][28] ), .Z(\w1[1][28] ) );
  XOR U2344 ( .A(key[157]), .B(\w0[1][29] ), .Z(\w1[1][29] ) );
  XOR U2345 ( .A(key[130]), .B(\w0[1][2] ), .Z(\w1[1][2] ) );
  XOR U2346 ( .A(key[158]), .B(\w0[1][30] ), .Z(\w1[1][30] ) );
  XOR U2347 ( .A(key[159]), .B(\w0[1][31] ), .Z(\w1[1][31] ) );
  XOR U2348 ( .A(key[160]), .B(\w0[1][32] ), .Z(\w1[1][32] ) );
  XOR U2349 ( .A(key[161]), .B(\w0[1][33] ), .Z(\w1[1][33] ) );
  XOR U2350 ( .A(key[162]), .B(\w0[1][34] ), .Z(\w1[1][34] ) );
  XOR U2351 ( .A(key[163]), .B(\w0[1][35] ), .Z(\w1[1][35] ) );
  XOR U2352 ( .A(key[164]), .B(\w0[1][36] ), .Z(\w1[1][36] ) );
  XOR U2353 ( .A(key[165]), .B(\w0[1][37] ), .Z(\w1[1][37] ) );
  XOR U2354 ( .A(key[166]), .B(\w0[1][38] ), .Z(\w1[1][38] ) );
  XOR U2355 ( .A(key[167]), .B(\w0[1][39] ), .Z(\w1[1][39] ) );
  XOR U2356 ( .A(key[131]), .B(\w0[1][3] ), .Z(\w1[1][3] ) );
  XOR U2357 ( .A(key[168]), .B(\w0[1][40] ), .Z(\w1[1][40] ) );
  XOR U2358 ( .A(key[169]), .B(\w0[1][41] ), .Z(\w1[1][41] ) );
  XOR U2359 ( .A(key[170]), .B(\w0[1][42] ), .Z(\w1[1][42] ) );
  XOR U2360 ( .A(key[171]), .B(\w0[1][43] ), .Z(\w1[1][43] ) );
  XOR U2361 ( .A(key[172]), .B(\w0[1][44] ), .Z(\w1[1][44] ) );
  XOR U2362 ( .A(key[173]), .B(\w0[1][45] ), .Z(\w1[1][45] ) );
  XOR U2363 ( .A(key[174]), .B(\w0[1][46] ), .Z(\w1[1][46] ) );
  XOR U2364 ( .A(key[175]), .B(\w0[1][47] ), .Z(\w1[1][47] ) );
  XOR U2365 ( .A(key[176]), .B(\w0[1][48] ), .Z(\w1[1][48] ) );
  XOR U2366 ( .A(key[177]), .B(\w0[1][49] ), .Z(\w1[1][49] ) );
  XOR U2367 ( .A(key[132]), .B(\w0[1][4] ), .Z(\w1[1][4] ) );
  XOR U2368 ( .A(key[178]), .B(\w0[1][50] ), .Z(\w1[1][50] ) );
  XOR U2369 ( .A(key[179]), .B(\w0[1][51] ), .Z(\w1[1][51] ) );
  XOR U2370 ( .A(key[180]), .B(\w0[1][52] ), .Z(\w1[1][52] ) );
  XOR U2371 ( .A(key[181]), .B(\w0[1][53] ), .Z(\w1[1][53] ) );
  XOR U2372 ( .A(key[182]), .B(\w0[1][54] ), .Z(\w1[1][54] ) );
  XOR U2373 ( .A(key[183]), .B(\w0[1][55] ), .Z(\w1[1][55] ) );
  XOR U2374 ( .A(key[184]), .B(\w0[1][56] ), .Z(\w1[1][56] ) );
  XOR U2375 ( .A(key[185]), .B(\w0[1][57] ), .Z(\w1[1][57] ) );
  XOR U2376 ( .A(key[186]), .B(\w0[1][58] ), .Z(\w1[1][58] ) );
  XOR U2377 ( .A(key[187]), .B(\w0[1][59] ), .Z(\w1[1][59] ) );
  XOR U2378 ( .A(key[133]), .B(\w0[1][5] ), .Z(\w1[1][5] ) );
  XOR U2379 ( .A(key[188]), .B(\w0[1][60] ), .Z(\w1[1][60] ) );
  XOR U2380 ( .A(key[189]), .B(\w0[1][61] ), .Z(\w1[1][61] ) );
  XOR U2381 ( .A(key[190]), .B(\w0[1][62] ), .Z(\w1[1][62] ) );
  XOR U2382 ( .A(key[191]), .B(\w0[1][63] ), .Z(\w1[1][63] ) );
  XOR U2383 ( .A(key[192]), .B(\w0[1][64] ), .Z(\w1[1][64] ) );
  XOR U2384 ( .A(key[193]), .B(\w0[1][65] ), .Z(\w1[1][65] ) );
  XOR U2385 ( .A(key[194]), .B(\w0[1][66] ), .Z(\w1[1][66] ) );
  XOR U2386 ( .A(key[195]), .B(\w0[1][67] ), .Z(\w1[1][67] ) );
  XOR U2387 ( .A(key[196]), .B(\w0[1][68] ), .Z(\w1[1][68] ) );
  XOR U2388 ( .A(key[197]), .B(\w0[1][69] ), .Z(\w1[1][69] ) );
  XOR U2389 ( .A(key[134]), .B(\w0[1][6] ), .Z(\w1[1][6] ) );
  XOR U2390 ( .A(key[198]), .B(\w0[1][70] ), .Z(\w1[1][70] ) );
  XOR U2391 ( .A(key[199]), .B(\w0[1][71] ), .Z(\w1[1][71] ) );
  XOR U2392 ( .A(key[200]), .B(\w0[1][72] ), .Z(\w1[1][72] ) );
  XOR U2393 ( .A(key[201]), .B(\w0[1][73] ), .Z(\w1[1][73] ) );
  XOR U2394 ( .A(key[202]), .B(\w0[1][74] ), .Z(\w1[1][74] ) );
  XOR U2395 ( .A(key[203]), .B(\w0[1][75] ), .Z(\w1[1][75] ) );
  XOR U2396 ( .A(key[204]), .B(\w0[1][76] ), .Z(\w1[1][76] ) );
  XOR U2397 ( .A(key[205]), .B(\w0[1][77] ), .Z(\w1[1][77] ) );
  XOR U2398 ( .A(key[206]), .B(\w0[1][78] ), .Z(\w1[1][78] ) );
  XOR U2399 ( .A(key[207]), .B(\w0[1][79] ), .Z(\w1[1][79] ) );
  XOR U2400 ( .A(key[135]), .B(\w0[1][7] ), .Z(\w1[1][7] ) );
  XOR U2401 ( .A(key[208]), .B(\w0[1][80] ), .Z(\w1[1][80] ) );
  XOR U2402 ( .A(key[209]), .B(\w0[1][81] ), .Z(\w1[1][81] ) );
  XOR U2403 ( .A(key[210]), .B(\w0[1][82] ), .Z(\w1[1][82] ) );
  XOR U2404 ( .A(key[211]), .B(\w0[1][83] ), .Z(\w1[1][83] ) );
  XOR U2405 ( .A(key[212]), .B(\w0[1][84] ), .Z(\w1[1][84] ) );
  XOR U2406 ( .A(key[213]), .B(\w0[1][85] ), .Z(\w1[1][85] ) );
  XOR U2407 ( .A(key[214]), .B(\w0[1][86] ), .Z(\w1[1][86] ) );
  XOR U2408 ( .A(key[215]), .B(\w0[1][87] ), .Z(\w1[1][87] ) );
  XOR U2409 ( .A(key[216]), .B(\w0[1][88] ), .Z(\w1[1][88] ) );
  XOR U2410 ( .A(key[217]), .B(\w0[1][89] ), .Z(\w1[1][89] ) );
  XOR U2411 ( .A(key[136]), .B(\w0[1][8] ), .Z(\w1[1][8] ) );
  XOR U2412 ( .A(key[218]), .B(\w0[1][90] ), .Z(\w1[1][90] ) );
  XOR U2413 ( .A(key[219]), .B(\w0[1][91] ), .Z(\w1[1][91] ) );
  XOR U2414 ( .A(key[220]), .B(\w0[1][92] ), .Z(\w1[1][92] ) );
  XOR U2415 ( .A(key[221]), .B(\w0[1][93] ), .Z(\w1[1][93] ) );
  XOR U2416 ( .A(key[222]), .B(\w0[1][94] ), .Z(\w1[1][94] ) );
  XOR U2417 ( .A(key[223]), .B(\w0[1][95] ), .Z(\w1[1][95] ) );
  XOR U2418 ( .A(key[224]), .B(\w0[1][96] ), .Z(\w1[1][96] ) );
  XOR U2419 ( .A(key[225]), .B(\w0[1][97] ), .Z(\w1[1][97] ) );
  XOR U2420 ( .A(key[226]), .B(\w0[1][98] ), .Z(\w1[1][98] ) );
  XOR U2421 ( .A(key[227]), .B(\w0[1][99] ), .Z(\w1[1][99] ) );
  XOR U2422 ( .A(key[137]), .B(\w0[1][9] ), .Z(\w1[1][9] ) );
endmodule

