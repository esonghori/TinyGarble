
module compare_N16384_CC128 ( clk, rst, x, y, g, e );
  input [127:0] x;
  input [127:0] y;
  input clk, rst;
  output g, e;
  wire   ebreg, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649;

  DFF ebreg_reg ( .D(n5), .CLK(clk), .RST(rst), .Q(ebreg) );
  DFF greg_reg ( .D(n4), .CLK(clk), .RST(rst), .Q(g) );
  IV U10 ( .A(ebreg), .Z(e) );
  XNOR U11 ( .A(y[95]), .B(x[95]), .Z(n9) );
  NANDN U12 ( .A(x[94]), .B(y[94]), .Z(n8) );
  NAND U13 ( .A(n9), .B(n8), .Z(n547) );
  XNOR U14 ( .A(y[89]), .B(x[89]), .Z(n11) );
  NANDN U15 ( .A(x[88]), .B(y[88]), .Z(n10) );
  NAND U16 ( .A(n11), .B(n10), .Z(n529) );
  NOR U17 ( .A(n547), .B(n529), .Z(n17) );
  XNOR U18 ( .A(y[93]), .B(x[93]), .Z(n13) );
  NANDN U19 ( .A(x[92]), .B(y[92]), .Z(n12) );
  NAND U20 ( .A(n13), .B(n12), .Z(n541) );
  XNOR U21 ( .A(y[91]), .B(x[91]), .Z(n15) );
  NANDN U22 ( .A(x[90]), .B(y[90]), .Z(n14) );
  NAND U23 ( .A(n15), .B(n14), .Z(n535) );
  NOR U24 ( .A(n541), .B(n535), .Z(n16) );
  AND U25 ( .A(n17), .B(n16), .Z(n29) );
  XNOR U26 ( .A(y[71]), .B(x[71]), .Z(n19) );
  NANDN U27 ( .A(x[70]), .B(y[70]), .Z(n18) );
  NAND U28 ( .A(n19), .B(n18), .Z(n475) );
  XNOR U29 ( .A(y[65]), .B(x[65]), .Z(n21) );
  NANDN U30 ( .A(x[64]), .B(y[64]), .Z(n20) );
  NAND U31 ( .A(n21), .B(n20), .Z(n457) );
  NOR U32 ( .A(n475), .B(n457), .Z(n27) );
  XNOR U33 ( .A(y[69]), .B(x[69]), .Z(n23) );
  NANDN U34 ( .A(x[68]), .B(y[68]), .Z(n22) );
  NAND U35 ( .A(n23), .B(n22), .Z(n469) );
  XNOR U36 ( .A(y[67]), .B(x[67]), .Z(n25) );
  NANDN U37 ( .A(x[66]), .B(y[66]), .Z(n24) );
  NAND U38 ( .A(n25), .B(n24), .Z(n463) );
  NOR U39 ( .A(n469), .B(n463), .Z(n26) );
  AND U40 ( .A(n27), .B(n26), .Z(n28) );
  AND U41 ( .A(n29), .B(n28), .Z(n53) );
  XNOR U42 ( .A(y[87]), .B(x[87]), .Z(n31) );
  NANDN U43 ( .A(x[86]), .B(y[86]), .Z(n30) );
  NAND U44 ( .A(n31), .B(n30), .Z(n523) );
  XNOR U45 ( .A(y[81]), .B(x[81]), .Z(n33) );
  NANDN U46 ( .A(x[80]), .B(y[80]), .Z(n32) );
  NAND U47 ( .A(n33), .B(n32), .Z(n505) );
  NOR U48 ( .A(n523), .B(n505), .Z(n39) );
  XNOR U49 ( .A(y[85]), .B(x[85]), .Z(n35) );
  NANDN U50 ( .A(x[84]), .B(y[84]), .Z(n34) );
  NAND U51 ( .A(n35), .B(n34), .Z(n517) );
  XNOR U52 ( .A(y[83]), .B(x[83]), .Z(n37) );
  NANDN U53 ( .A(x[82]), .B(y[82]), .Z(n36) );
  NAND U54 ( .A(n37), .B(n36), .Z(n511) );
  NOR U55 ( .A(n517), .B(n511), .Z(n38) );
  AND U56 ( .A(n39), .B(n38), .Z(n51) );
  XNOR U57 ( .A(y[79]), .B(x[79]), .Z(n41) );
  NANDN U58 ( .A(x[78]), .B(y[78]), .Z(n40) );
  NAND U59 ( .A(n41), .B(n40), .Z(n499) );
  XNOR U60 ( .A(y[73]), .B(x[73]), .Z(n43) );
  NANDN U61 ( .A(x[72]), .B(y[72]), .Z(n42) );
  NAND U62 ( .A(n43), .B(n42), .Z(n481) );
  NOR U63 ( .A(n499), .B(n481), .Z(n49) );
  XNOR U64 ( .A(y[77]), .B(x[77]), .Z(n45) );
  NANDN U65 ( .A(x[76]), .B(y[76]), .Z(n44) );
  NAND U66 ( .A(n45), .B(n44), .Z(n493) );
  XNOR U67 ( .A(y[75]), .B(x[75]), .Z(n47) );
  NANDN U68 ( .A(x[74]), .B(y[74]), .Z(n46) );
  NAND U69 ( .A(n47), .B(n46), .Z(n487) );
  NOR U70 ( .A(n493), .B(n487), .Z(n48) );
  AND U71 ( .A(n49), .B(n48), .Z(n50) );
  AND U72 ( .A(n51), .B(n50), .Z(n52) );
  AND U73 ( .A(n53), .B(n52), .Z(n262) );
  XNOR U74 ( .A(y[23]), .B(x[23]), .Z(n55) );
  NANDN U75 ( .A(x[22]), .B(y[22]), .Z(n54) );
  NAND U76 ( .A(n55), .B(n54), .Z(n331) );
  XNOR U77 ( .A(y[17]), .B(x[17]), .Z(n57) );
  NANDN U78 ( .A(x[16]), .B(y[16]), .Z(n56) );
  NAND U79 ( .A(n57), .B(n56), .Z(n313) );
  NOR U80 ( .A(n331), .B(n313), .Z(n63) );
  XNOR U81 ( .A(y[21]), .B(x[21]), .Z(n59) );
  NANDN U82 ( .A(x[20]), .B(y[20]), .Z(n58) );
  NAND U83 ( .A(n59), .B(n58), .Z(n325) );
  XNOR U84 ( .A(y[19]), .B(x[19]), .Z(n61) );
  NANDN U85 ( .A(x[18]), .B(y[18]), .Z(n60) );
  NAND U86 ( .A(n61), .B(n60), .Z(n319) );
  NOR U87 ( .A(n325), .B(n319), .Z(n62) );
  AND U88 ( .A(n63), .B(n62), .Z(n76) );
  XNOR U89 ( .A(y[1]), .B(x[1]), .Z(n65) );
  NANDN U90 ( .A(x[0]), .B(y[0]), .Z(n64) );
  AND U91 ( .A(n65), .B(n64), .Z(n68) );
  XNOR U92 ( .A(y[13]), .B(x[13]), .Z(n67) );
  NANDN U93 ( .A(x[12]), .B(y[12]), .Z(n66) );
  NAND U94 ( .A(n67), .B(n66), .Z(n300) );
  ANDN U95 ( .B(n68), .A(n300), .Z(n74) );
  XNOR U96 ( .A(x[3]), .B(y[3]), .Z(n70) );
  NANDN U97 ( .A(x[2]), .B(y[2]), .Z(n69) );
  NAND U98 ( .A(n70), .B(n69), .Z(n281) );
  XNOR U99 ( .A(y[15]), .B(x[15]), .Z(n72) );
  NANDN U100 ( .A(x[14]), .B(y[14]), .Z(n71) );
  NAND U101 ( .A(n72), .B(n71), .Z(n307) );
  NOR U102 ( .A(n281), .B(n307), .Z(n73) );
  AND U103 ( .A(n74), .B(n73), .Z(n75) );
  AND U104 ( .A(n76), .B(n75), .Z(n100) );
  XNOR U105 ( .A(y[31]), .B(x[31]), .Z(n78) );
  NANDN U106 ( .A(x[30]), .B(y[30]), .Z(n77) );
  NAND U107 ( .A(n78), .B(n77), .Z(n355) );
  XNOR U108 ( .A(y[25]), .B(x[25]), .Z(n80) );
  NANDN U109 ( .A(x[24]), .B(y[24]), .Z(n79) );
  NAND U110 ( .A(n80), .B(n79), .Z(n337) );
  NOR U111 ( .A(n355), .B(n337), .Z(n86) );
  XNOR U112 ( .A(y[29]), .B(x[29]), .Z(n82) );
  NANDN U113 ( .A(x[28]), .B(y[28]), .Z(n81) );
  NAND U114 ( .A(n82), .B(n81), .Z(n349) );
  XNOR U115 ( .A(y[27]), .B(x[27]), .Z(n84) );
  NANDN U116 ( .A(x[26]), .B(y[26]), .Z(n83) );
  NAND U117 ( .A(n84), .B(n83), .Z(n343) );
  NOR U118 ( .A(n349), .B(n343), .Z(n85) );
  AND U119 ( .A(n86), .B(n85), .Z(n98) );
  XNOR U120 ( .A(y[11]), .B(x[11]), .Z(n88) );
  NANDN U121 ( .A(x[10]), .B(y[10]), .Z(n87) );
  NAND U122 ( .A(n88), .B(n87), .Z(n297) );
  XNOR U123 ( .A(y[5]), .B(x[5]), .Z(n90) );
  NANDN U124 ( .A(x[4]), .B(y[4]), .Z(n89) );
  NAND U125 ( .A(n90), .B(n89), .Z(n285) );
  NOR U126 ( .A(n297), .B(n285), .Z(n96) );
  XNOR U127 ( .A(y[9]), .B(x[9]), .Z(n92) );
  NANDN U128 ( .A(x[8]), .B(y[8]), .Z(n91) );
  NAND U129 ( .A(n92), .B(n91), .Z(n293) );
  XNOR U130 ( .A(y[7]), .B(x[7]), .Z(n94) );
  NANDN U131 ( .A(x[6]), .B(y[6]), .Z(n93) );
  NAND U132 ( .A(n94), .B(n93), .Z(n289) );
  NOR U133 ( .A(n293), .B(n289), .Z(n95) );
  AND U134 ( .A(n96), .B(n95), .Z(n97) );
  AND U135 ( .A(n98), .B(n97), .Z(n99) );
  AND U136 ( .A(n100), .B(n99), .Z(n148) );
  XNOR U137 ( .A(y[127]), .B(x[127]), .Z(n102) );
  NANDN U138 ( .A(x[126]), .B(y[126]), .Z(n101) );
  NAND U139 ( .A(n102), .B(n101), .Z(n643) );
  XNOR U140 ( .A(y[121]), .B(x[121]), .Z(n104) );
  NANDN U141 ( .A(x[120]), .B(y[120]), .Z(n103) );
  NAND U142 ( .A(n104), .B(n103), .Z(n625) );
  NOR U143 ( .A(n643), .B(n625), .Z(n110) );
  XNOR U144 ( .A(y[125]), .B(x[125]), .Z(n106) );
  NANDN U145 ( .A(x[124]), .B(y[124]), .Z(n105) );
  NAND U146 ( .A(n106), .B(n105), .Z(n637) );
  XNOR U147 ( .A(y[123]), .B(x[123]), .Z(n108) );
  NANDN U148 ( .A(x[122]), .B(y[122]), .Z(n107) );
  NAND U149 ( .A(n108), .B(n107), .Z(n631) );
  NOR U150 ( .A(n637), .B(n631), .Z(n109) );
  AND U151 ( .A(n110), .B(n109), .Z(n122) );
  XNOR U152 ( .A(y[103]), .B(x[103]), .Z(n112) );
  NANDN U153 ( .A(x[102]), .B(y[102]), .Z(n111) );
  NAND U154 ( .A(n112), .B(n111), .Z(n571) );
  XNOR U155 ( .A(y[97]), .B(x[97]), .Z(n114) );
  NANDN U156 ( .A(x[96]), .B(y[96]), .Z(n113) );
  NAND U157 ( .A(n114), .B(n113), .Z(n553) );
  NOR U158 ( .A(n571), .B(n553), .Z(n120) );
  XNOR U159 ( .A(y[101]), .B(x[101]), .Z(n116) );
  NANDN U160 ( .A(x[100]), .B(y[100]), .Z(n115) );
  NAND U161 ( .A(n116), .B(n115), .Z(n565) );
  XNOR U162 ( .A(y[99]), .B(x[99]), .Z(n118) );
  NANDN U163 ( .A(x[98]), .B(y[98]), .Z(n117) );
  NAND U164 ( .A(n118), .B(n117), .Z(n559) );
  NOR U165 ( .A(n565), .B(n559), .Z(n119) );
  AND U166 ( .A(n120), .B(n119), .Z(n121) );
  AND U167 ( .A(n122), .B(n121), .Z(n146) );
  XNOR U168 ( .A(y[119]), .B(x[119]), .Z(n124) );
  NANDN U169 ( .A(x[118]), .B(y[118]), .Z(n123) );
  NAND U170 ( .A(n124), .B(n123), .Z(n619) );
  XNOR U171 ( .A(y[113]), .B(x[113]), .Z(n126) );
  NANDN U172 ( .A(x[112]), .B(y[112]), .Z(n125) );
  NAND U173 ( .A(n126), .B(n125), .Z(n601) );
  NOR U174 ( .A(n619), .B(n601), .Z(n132) );
  XNOR U175 ( .A(y[117]), .B(x[117]), .Z(n128) );
  NANDN U176 ( .A(x[116]), .B(y[116]), .Z(n127) );
  NAND U177 ( .A(n128), .B(n127), .Z(n613) );
  XNOR U178 ( .A(y[115]), .B(x[115]), .Z(n130) );
  NANDN U179 ( .A(x[114]), .B(y[114]), .Z(n129) );
  NAND U180 ( .A(n130), .B(n129), .Z(n607) );
  NOR U181 ( .A(n613), .B(n607), .Z(n131) );
  AND U182 ( .A(n132), .B(n131), .Z(n144) );
  XNOR U183 ( .A(y[111]), .B(x[111]), .Z(n134) );
  NANDN U184 ( .A(x[110]), .B(y[110]), .Z(n133) );
  NAND U185 ( .A(n134), .B(n133), .Z(n595) );
  XNOR U186 ( .A(y[105]), .B(x[105]), .Z(n136) );
  NANDN U187 ( .A(x[104]), .B(y[104]), .Z(n135) );
  NAND U188 ( .A(n136), .B(n135), .Z(n577) );
  NOR U189 ( .A(n595), .B(n577), .Z(n142) );
  XNOR U190 ( .A(y[109]), .B(x[109]), .Z(n138) );
  NANDN U191 ( .A(x[108]), .B(y[108]), .Z(n137) );
  NAND U192 ( .A(n138), .B(n137), .Z(n589) );
  XNOR U193 ( .A(y[107]), .B(x[107]), .Z(n140) );
  NANDN U194 ( .A(x[106]), .B(y[106]), .Z(n139) );
  NAND U195 ( .A(n140), .B(n139), .Z(n583) );
  NOR U196 ( .A(n589), .B(n583), .Z(n141) );
  AND U197 ( .A(n142), .B(n141), .Z(n143) );
  AND U198 ( .A(n144), .B(n143), .Z(n145) );
  AND U199 ( .A(n146), .B(n145), .Z(n147) );
  AND U200 ( .A(n148), .B(n147), .Z(n260) );
  XNOR U201 ( .A(y[55]), .B(x[55]), .Z(n150) );
  NANDN U202 ( .A(x[54]), .B(y[54]), .Z(n149) );
  NAND U203 ( .A(n150), .B(n149), .Z(n427) );
  XNOR U204 ( .A(y[49]), .B(x[49]), .Z(n152) );
  NANDN U205 ( .A(x[48]), .B(y[48]), .Z(n151) );
  NAND U206 ( .A(n152), .B(n151), .Z(n409) );
  NOR U207 ( .A(n427), .B(n409), .Z(n158) );
  XNOR U208 ( .A(y[53]), .B(x[53]), .Z(n154) );
  NANDN U209 ( .A(x[52]), .B(y[52]), .Z(n153) );
  NAND U210 ( .A(n154), .B(n153), .Z(n421) );
  XNOR U211 ( .A(y[51]), .B(x[51]), .Z(n156) );
  NANDN U212 ( .A(x[50]), .B(y[50]), .Z(n155) );
  NAND U213 ( .A(n156), .B(n155), .Z(n415) );
  NOR U214 ( .A(n421), .B(n415), .Z(n157) );
  AND U215 ( .A(n158), .B(n157), .Z(n170) );
  XNOR U216 ( .A(y[47]), .B(x[47]), .Z(n160) );
  NANDN U217 ( .A(x[46]), .B(y[46]), .Z(n159) );
  NAND U218 ( .A(n160), .B(n159), .Z(n403) );
  XNOR U219 ( .A(y[41]), .B(x[41]), .Z(n162) );
  NANDN U220 ( .A(x[40]), .B(y[40]), .Z(n161) );
  NAND U221 ( .A(n162), .B(n161), .Z(n385) );
  NOR U222 ( .A(n403), .B(n385), .Z(n168) );
  XNOR U223 ( .A(y[45]), .B(x[45]), .Z(n164) );
  NANDN U224 ( .A(x[44]), .B(y[44]), .Z(n163) );
  NAND U225 ( .A(n164), .B(n163), .Z(n397) );
  XNOR U226 ( .A(y[43]), .B(x[43]), .Z(n166) );
  NANDN U227 ( .A(x[42]), .B(y[42]), .Z(n165) );
  NAND U228 ( .A(n166), .B(n165), .Z(n391) );
  NOR U229 ( .A(n397), .B(n391), .Z(n167) );
  AND U230 ( .A(n168), .B(n167), .Z(n169) );
  AND U231 ( .A(n170), .B(n169), .Z(n194) );
  XNOR U232 ( .A(y[63]), .B(x[63]), .Z(n172) );
  NANDN U233 ( .A(x[62]), .B(y[62]), .Z(n171) );
  NAND U234 ( .A(n172), .B(n171), .Z(n451) );
  XNOR U235 ( .A(y[57]), .B(x[57]), .Z(n174) );
  NANDN U236 ( .A(x[56]), .B(y[56]), .Z(n173) );
  NAND U237 ( .A(n174), .B(n173), .Z(n433) );
  NOR U238 ( .A(n451), .B(n433), .Z(n180) );
  XNOR U239 ( .A(y[61]), .B(x[61]), .Z(n176) );
  NANDN U240 ( .A(x[60]), .B(y[60]), .Z(n175) );
  NAND U241 ( .A(n176), .B(n175), .Z(n445) );
  XNOR U242 ( .A(y[59]), .B(x[59]), .Z(n178) );
  NANDN U243 ( .A(x[58]), .B(y[58]), .Z(n177) );
  NAND U244 ( .A(n178), .B(n177), .Z(n439) );
  NOR U245 ( .A(n445), .B(n439), .Z(n179) );
  AND U246 ( .A(n180), .B(n179), .Z(n192) );
  XNOR U247 ( .A(y[39]), .B(x[39]), .Z(n182) );
  NANDN U248 ( .A(x[38]), .B(y[38]), .Z(n181) );
  NAND U249 ( .A(n182), .B(n181), .Z(n379) );
  XNOR U250 ( .A(y[33]), .B(x[33]), .Z(n184) );
  NANDN U251 ( .A(x[32]), .B(y[32]), .Z(n183) );
  NAND U252 ( .A(n184), .B(n183), .Z(n361) );
  NOR U253 ( .A(n379), .B(n361), .Z(n190) );
  XNOR U254 ( .A(y[37]), .B(x[37]), .Z(n186) );
  NANDN U255 ( .A(x[36]), .B(y[36]), .Z(n185) );
  NAND U256 ( .A(n186), .B(n185), .Z(n373) );
  XNOR U257 ( .A(y[35]), .B(x[35]), .Z(n188) );
  NANDN U258 ( .A(x[34]), .B(y[34]), .Z(n187) );
  NAND U259 ( .A(n188), .B(n187), .Z(n367) );
  NOR U260 ( .A(n373), .B(n367), .Z(n189) );
  AND U261 ( .A(n190), .B(n189), .Z(n191) );
  AND U262 ( .A(n192), .B(n191), .Z(n193) );
  AND U263 ( .A(n194), .B(n193), .Z(n258) );
  ANDN U264 ( .B(x[126]), .A(y[126]), .Z(n639) );
  ANDN U265 ( .B(x[120]), .A(y[120]), .Z(n621) );
  NOR U266 ( .A(n639), .B(n621), .Z(n196) );
  ANDN U267 ( .B(x[124]), .A(y[124]), .Z(n633) );
  ANDN U268 ( .B(x[122]), .A(y[122]), .Z(n627) );
  NOR U269 ( .A(n633), .B(n627), .Z(n195) );
  AND U270 ( .A(n196), .B(n195), .Z(n200) );
  ANDN U271 ( .B(x[102]), .A(y[102]), .Z(n567) );
  ANDN U272 ( .B(x[96]), .A(y[96]), .Z(n549) );
  NOR U273 ( .A(n567), .B(n549), .Z(n198) );
  ANDN U274 ( .B(x[100]), .A(y[100]), .Z(n561) );
  ANDN U275 ( .B(x[98]), .A(y[98]), .Z(n555) );
  NOR U276 ( .A(n561), .B(n555), .Z(n197) );
  AND U277 ( .A(n198), .B(n197), .Z(n199) );
  AND U278 ( .A(n200), .B(n199), .Z(n208) );
  ANDN U279 ( .B(x[118]), .A(y[118]), .Z(n615) );
  ANDN U280 ( .B(x[112]), .A(y[112]), .Z(n597) );
  NOR U281 ( .A(n615), .B(n597), .Z(n202) );
  ANDN U282 ( .B(x[116]), .A(y[116]), .Z(n609) );
  ANDN U283 ( .B(x[114]), .A(y[114]), .Z(n603) );
  NOR U284 ( .A(n609), .B(n603), .Z(n201) );
  AND U285 ( .A(n202), .B(n201), .Z(n206) );
  ANDN U286 ( .B(x[110]), .A(y[110]), .Z(n591) );
  ANDN U287 ( .B(x[104]), .A(y[104]), .Z(n573) );
  NOR U288 ( .A(n591), .B(n573), .Z(n204) );
  ANDN U289 ( .B(x[108]), .A(y[108]), .Z(n585) );
  ANDN U290 ( .B(x[106]), .A(y[106]), .Z(n579) );
  NOR U291 ( .A(n585), .B(n579), .Z(n203) );
  AND U292 ( .A(n204), .B(n203), .Z(n205) );
  AND U293 ( .A(n206), .B(n205), .Z(n207) );
  AND U294 ( .A(n208), .B(n207), .Z(n224) );
  ANDN U295 ( .B(x[30]), .A(y[30]), .Z(n353) );
  ANDN U296 ( .B(x[24]), .A(y[24]), .Z(n335) );
  NOR U297 ( .A(n353), .B(n335), .Z(n210) );
  ANDN U298 ( .B(x[28]), .A(y[28]), .Z(n347) );
  ANDN U299 ( .B(x[26]), .A(y[26]), .Z(n341) );
  NOR U300 ( .A(n347), .B(n341), .Z(n209) );
  AND U301 ( .A(n210), .B(n209), .Z(n214) );
  ANDN U302 ( .B(x[6]), .A(y[6]), .Z(n270) );
  ANDN U303 ( .B(x[4]), .A(y[4]), .Z(n272) );
  NOR U304 ( .A(n270), .B(n272), .Z(n212) );
  NANDN U305 ( .A(y[0]), .B(x[0]), .Z(n274) );
  ANDN U306 ( .B(x[2]), .A(y[2]), .Z(n278) );
  ANDN U307 ( .B(n274), .A(n278), .Z(n211) );
  AND U308 ( .A(n212), .B(n211), .Z(n213) );
  AND U309 ( .A(n214), .B(n213), .Z(n222) );
  ANDN U310 ( .B(x[22]), .A(y[22]), .Z(n329) );
  ANDN U311 ( .B(x[16]), .A(y[16]), .Z(n311) );
  NOR U312 ( .A(n329), .B(n311), .Z(n216) );
  ANDN U313 ( .B(x[20]), .A(y[20]), .Z(n323) );
  ANDN U314 ( .B(x[18]), .A(y[18]), .Z(n317) );
  NOR U315 ( .A(n323), .B(n317), .Z(n215) );
  AND U316 ( .A(n216), .B(n215), .Z(n220) );
  ANDN U317 ( .B(x[14]), .A(y[14]), .Z(n305) );
  ANDN U318 ( .B(x[8]), .A(y[8]), .Z(n268) );
  NOR U319 ( .A(n305), .B(n268), .Z(n218) );
  ANDN U320 ( .B(x[12]), .A(y[12]), .Z(n264) );
  ANDN U321 ( .B(x[10]), .A(y[10]), .Z(n266) );
  NOR U322 ( .A(n264), .B(n266), .Z(n217) );
  AND U323 ( .A(n218), .B(n217), .Z(n219) );
  AND U324 ( .A(n220), .B(n219), .Z(n221) );
  AND U325 ( .A(n222), .B(n221), .Z(n223) );
  AND U326 ( .A(n224), .B(n223), .Z(n256) );
  ANDN U327 ( .B(x[94]), .A(y[94]), .Z(n543) );
  ANDN U328 ( .B(x[88]), .A(y[88]), .Z(n525) );
  NOR U329 ( .A(n543), .B(n525), .Z(n226) );
  ANDN U330 ( .B(x[92]), .A(y[92]), .Z(n537) );
  ANDN U331 ( .B(x[90]), .A(y[90]), .Z(n531) );
  NOR U332 ( .A(n537), .B(n531), .Z(n225) );
  AND U333 ( .A(n226), .B(n225), .Z(n230) );
  ANDN U334 ( .B(x[70]), .A(y[70]), .Z(n471) );
  ANDN U335 ( .B(x[64]), .A(y[64]), .Z(n455) );
  NOR U336 ( .A(n471), .B(n455), .Z(n228) );
  ANDN U337 ( .B(x[68]), .A(y[68]), .Z(n465) );
  ANDN U338 ( .B(x[66]), .A(y[66]), .Z(n459) );
  NOR U339 ( .A(n465), .B(n459), .Z(n227) );
  AND U340 ( .A(n228), .B(n227), .Z(n229) );
  AND U341 ( .A(n230), .B(n229), .Z(n238) );
  ANDN U342 ( .B(x[86]), .A(y[86]), .Z(n519) );
  ANDN U343 ( .B(x[80]), .A(y[80]), .Z(n501) );
  NOR U344 ( .A(n519), .B(n501), .Z(n232) );
  ANDN U345 ( .B(x[84]), .A(y[84]), .Z(n513) );
  ANDN U346 ( .B(x[82]), .A(y[82]), .Z(n507) );
  NOR U347 ( .A(n513), .B(n507), .Z(n231) );
  AND U348 ( .A(n232), .B(n231), .Z(n236) );
  ANDN U349 ( .B(x[78]), .A(y[78]), .Z(n495) );
  ANDN U350 ( .B(x[72]), .A(y[72]), .Z(n477) );
  NOR U351 ( .A(n495), .B(n477), .Z(n234) );
  ANDN U352 ( .B(x[76]), .A(y[76]), .Z(n489) );
  ANDN U353 ( .B(x[74]), .A(y[74]), .Z(n483) );
  NOR U354 ( .A(n489), .B(n483), .Z(n233) );
  AND U355 ( .A(n234), .B(n233), .Z(n235) );
  AND U356 ( .A(n236), .B(n235), .Z(n237) );
  AND U357 ( .A(n238), .B(n237), .Z(n254) );
  ANDN U358 ( .B(x[62]), .A(y[62]), .Z(n449) );
  ANDN U359 ( .B(x[56]), .A(y[56]), .Z(n431) );
  NOR U360 ( .A(n449), .B(n431), .Z(n240) );
  ANDN U361 ( .B(x[60]), .A(y[60]), .Z(n443) );
  ANDN U362 ( .B(x[58]), .A(y[58]), .Z(n437) );
  NOR U363 ( .A(n443), .B(n437), .Z(n239) );
  AND U364 ( .A(n240), .B(n239), .Z(n244) );
  ANDN U365 ( .B(x[38]), .A(y[38]), .Z(n377) );
  ANDN U366 ( .B(x[32]), .A(y[32]), .Z(n359) );
  NOR U367 ( .A(n377), .B(n359), .Z(n242) );
  ANDN U368 ( .B(x[36]), .A(y[36]), .Z(n371) );
  ANDN U369 ( .B(x[34]), .A(y[34]), .Z(n365) );
  NOR U370 ( .A(n371), .B(n365), .Z(n241) );
  AND U371 ( .A(n242), .B(n241), .Z(n243) );
  AND U372 ( .A(n244), .B(n243), .Z(n252) );
  ANDN U373 ( .B(x[54]), .A(y[54]), .Z(n425) );
  ANDN U374 ( .B(x[48]), .A(y[48]), .Z(n407) );
  NOR U375 ( .A(n425), .B(n407), .Z(n246) );
  ANDN U376 ( .B(x[52]), .A(y[52]), .Z(n419) );
  ANDN U377 ( .B(x[50]), .A(y[50]), .Z(n413) );
  NOR U378 ( .A(n419), .B(n413), .Z(n245) );
  AND U379 ( .A(n246), .B(n245), .Z(n250) );
  ANDN U380 ( .B(x[46]), .A(y[46]), .Z(n401) );
  ANDN U381 ( .B(x[40]), .A(y[40]), .Z(n383) );
  NOR U382 ( .A(n401), .B(n383), .Z(n248) );
  ANDN U383 ( .B(x[44]), .A(y[44]), .Z(n395) );
  ANDN U384 ( .B(x[42]), .A(y[42]), .Z(n389) );
  NOR U385 ( .A(n395), .B(n389), .Z(n247) );
  AND U386 ( .A(n248), .B(n247), .Z(n249) );
  AND U387 ( .A(n250), .B(n249), .Z(n251) );
  AND U388 ( .A(n252), .B(n251), .Z(n253) );
  AND U389 ( .A(n254), .B(n253), .Z(n255) );
  AND U390 ( .A(n256), .B(n255), .Z(n257) );
  AND U391 ( .A(n258), .B(n257), .Z(n259) );
  AND U392 ( .A(n260), .B(n259), .Z(n261) );
  AND U393 ( .A(n262), .B(n261), .Z(n263) );
  NAND U394 ( .A(e), .B(n263), .Z(n5) );
  NANDN U395 ( .A(n263), .B(e), .Z(n647) );
  ANDN U396 ( .B(x[127]), .A(y[127]), .Z(n645) );
  ANDN U397 ( .B(x[63]), .A(y[63]), .Z(n453) );
  ANDN U398 ( .B(x[61]), .A(y[61]), .Z(n447) );
  ANDN U399 ( .B(x[59]), .A(y[59]), .Z(n441) );
  ANDN U400 ( .B(x[57]), .A(y[57]), .Z(n435) );
  ANDN U401 ( .B(x[55]), .A(y[55]), .Z(n429) );
  ANDN U402 ( .B(x[53]), .A(y[53]), .Z(n423) );
  ANDN U403 ( .B(x[51]), .A(y[51]), .Z(n417) );
  ANDN U404 ( .B(x[49]), .A(y[49]), .Z(n411) );
  ANDN U405 ( .B(x[47]), .A(y[47]), .Z(n405) );
  ANDN U406 ( .B(x[45]), .A(y[45]), .Z(n399) );
  ANDN U407 ( .B(x[43]), .A(y[43]), .Z(n393) );
  ANDN U408 ( .B(x[41]), .A(y[41]), .Z(n387) );
  ANDN U409 ( .B(x[39]), .A(y[39]), .Z(n381) );
  ANDN U410 ( .B(x[37]), .A(y[37]), .Z(n375) );
  ANDN U411 ( .B(x[35]), .A(y[35]), .Z(n369) );
  ANDN U412 ( .B(x[33]), .A(y[33]), .Z(n363) );
  ANDN U413 ( .B(x[31]), .A(y[31]), .Z(n357) );
  ANDN U414 ( .B(x[29]), .A(y[29]), .Z(n351) );
  ANDN U415 ( .B(x[27]), .A(y[27]), .Z(n345) );
  ANDN U416 ( .B(x[25]), .A(y[25]), .Z(n339) );
  ANDN U417 ( .B(x[23]), .A(y[23]), .Z(n333) );
  ANDN U418 ( .B(x[21]), .A(y[21]), .Z(n327) );
  ANDN U419 ( .B(x[19]), .A(y[19]), .Z(n321) );
  ANDN U420 ( .B(x[17]), .A(y[17]), .Z(n315) );
  ANDN U421 ( .B(x[15]), .A(y[15]), .Z(n309) );
  NANDN U422 ( .A(y[13]), .B(x[13]), .Z(n303) );
  NANDN U423 ( .A(y[11]), .B(x[11]), .Z(n265) );
  ANDN U424 ( .B(n265), .A(n264), .Z(n299) );
  NANDN U425 ( .A(y[9]), .B(x[9]), .Z(n267) );
  ANDN U426 ( .B(n267), .A(n266), .Z(n295) );
  NANDN U427 ( .A(y[7]), .B(x[7]), .Z(n269) );
  ANDN U428 ( .B(n269), .A(n268), .Z(n291) );
  NANDN U429 ( .A(y[5]), .B(x[5]), .Z(n271) );
  ANDN U430 ( .B(n271), .A(n270), .Z(n287) );
  NANDN U431 ( .A(y[3]), .B(x[3]), .Z(n273) );
  ANDN U432 ( .B(n273), .A(n272), .Z(n283) );
  NANDN U433 ( .A(x[1]), .B(n274), .Z(n277) );
  XNOR U434 ( .A(n274), .B(x[1]), .Z(n275) );
  NAND U435 ( .A(n275), .B(y[1]), .Z(n276) );
  NAND U436 ( .A(n277), .B(n276), .Z(n279) );
  ANDN U437 ( .B(n279), .A(n278), .Z(n280) );
  OR U438 ( .A(n281), .B(n280), .Z(n282) );
  AND U439 ( .A(n283), .B(n282), .Z(n284) );
  OR U440 ( .A(n285), .B(n284), .Z(n286) );
  AND U441 ( .A(n287), .B(n286), .Z(n288) );
  OR U442 ( .A(n289), .B(n288), .Z(n290) );
  AND U443 ( .A(n291), .B(n290), .Z(n292) );
  OR U444 ( .A(n293), .B(n292), .Z(n294) );
  AND U445 ( .A(n295), .B(n294), .Z(n296) );
  OR U446 ( .A(n297), .B(n296), .Z(n298) );
  AND U447 ( .A(n299), .B(n298), .Z(n301) );
  OR U448 ( .A(n301), .B(n300), .Z(n302) );
  AND U449 ( .A(n303), .B(n302), .Z(n304) );
  NANDN U450 ( .A(n305), .B(n304), .Z(n306) );
  NANDN U451 ( .A(n307), .B(n306), .Z(n308) );
  NANDN U452 ( .A(n309), .B(n308), .Z(n310) );
  OR U453 ( .A(n311), .B(n310), .Z(n312) );
  NANDN U454 ( .A(n313), .B(n312), .Z(n314) );
  NANDN U455 ( .A(n315), .B(n314), .Z(n316) );
  OR U456 ( .A(n317), .B(n316), .Z(n318) );
  NANDN U457 ( .A(n319), .B(n318), .Z(n320) );
  NANDN U458 ( .A(n321), .B(n320), .Z(n322) );
  OR U459 ( .A(n323), .B(n322), .Z(n324) );
  NANDN U460 ( .A(n325), .B(n324), .Z(n326) );
  NANDN U461 ( .A(n327), .B(n326), .Z(n328) );
  OR U462 ( .A(n329), .B(n328), .Z(n330) );
  NANDN U463 ( .A(n331), .B(n330), .Z(n332) );
  NANDN U464 ( .A(n333), .B(n332), .Z(n334) );
  OR U465 ( .A(n335), .B(n334), .Z(n336) );
  NANDN U466 ( .A(n337), .B(n336), .Z(n338) );
  NANDN U467 ( .A(n339), .B(n338), .Z(n340) );
  OR U468 ( .A(n341), .B(n340), .Z(n342) );
  NANDN U469 ( .A(n343), .B(n342), .Z(n344) );
  NANDN U470 ( .A(n345), .B(n344), .Z(n346) );
  OR U471 ( .A(n347), .B(n346), .Z(n348) );
  NANDN U472 ( .A(n349), .B(n348), .Z(n350) );
  NANDN U473 ( .A(n351), .B(n350), .Z(n352) );
  OR U474 ( .A(n353), .B(n352), .Z(n354) );
  NANDN U475 ( .A(n355), .B(n354), .Z(n356) );
  NANDN U476 ( .A(n357), .B(n356), .Z(n358) );
  OR U477 ( .A(n359), .B(n358), .Z(n360) );
  NANDN U478 ( .A(n361), .B(n360), .Z(n362) );
  NANDN U479 ( .A(n363), .B(n362), .Z(n364) );
  OR U480 ( .A(n365), .B(n364), .Z(n366) );
  NANDN U481 ( .A(n367), .B(n366), .Z(n368) );
  NANDN U482 ( .A(n369), .B(n368), .Z(n370) );
  OR U483 ( .A(n371), .B(n370), .Z(n372) );
  NANDN U484 ( .A(n373), .B(n372), .Z(n374) );
  NANDN U485 ( .A(n375), .B(n374), .Z(n376) );
  OR U486 ( .A(n377), .B(n376), .Z(n378) );
  NANDN U487 ( .A(n379), .B(n378), .Z(n380) );
  NANDN U488 ( .A(n381), .B(n380), .Z(n382) );
  OR U489 ( .A(n383), .B(n382), .Z(n384) );
  NANDN U490 ( .A(n385), .B(n384), .Z(n386) );
  NANDN U491 ( .A(n387), .B(n386), .Z(n388) );
  OR U492 ( .A(n389), .B(n388), .Z(n390) );
  NANDN U493 ( .A(n391), .B(n390), .Z(n392) );
  NANDN U494 ( .A(n393), .B(n392), .Z(n394) );
  OR U495 ( .A(n395), .B(n394), .Z(n396) );
  NANDN U496 ( .A(n397), .B(n396), .Z(n398) );
  NANDN U497 ( .A(n399), .B(n398), .Z(n400) );
  OR U498 ( .A(n401), .B(n400), .Z(n402) );
  NANDN U499 ( .A(n403), .B(n402), .Z(n404) );
  NANDN U500 ( .A(n405), .B(n404), .Z(n406) );
  OR U501 ( .A(n407), .B(n406), .Z(n408) );
  NANDN U502 ( .A(n409), .B(n408), .Z(n410) );
  NANDN U503 ( .A(n411), .B(n410), .Z(n412) );
  OR U504 ( .A(n413), .B(n412), .Z(n414) );
  NANDN U505 ( .A(n415), .B(n414), .Z(n416) );
  NANDN U506 ( .A(n417), .B(n416), .Z(n418) );
  OR U507 ( .A(n419), .B(n418), .Z(n420) );
  NANDN U508 ( .A(n421), .B(n420), .Z(n422) );
  NANDN U509 ( .A(n423), .B(n422), .Z(n424) );
  OR U510 ( .A(n425), .B(n424), .Z(n426) );
  NANDN U511 ( .A(n427), .B(n426), .Z(n428) );
  NANDN U512 ( .A(n429), .B(n428), .Z(n430) );
  OR U513 ( .A(n431), .B(n430), .Z(n432) );
  NANDN U514 ( .A(n433), .B(n432), .Z(n434) );
  NANDN U515 ( .A(n435), .B(n434), .Z(n436) );
  OR U516 ( .A(n437), .B(n436), .Z(n438) );
  NANDN U517 ( .A(n439), .B(n438), .Z(n440) );
  NANDN U518 ( .A(n441), .B(n440), .Z(n442) );
  OR U519 ( .A(n443), .B(n442), .Z(n444) );
  NANDN U520 ( .A(n445), .B(n444), .Z(n446) );
  NANDN U521 ( .A(n447), .B(n446), .Z(n448) );
  OR U522 ( .A(n449), .B(n448), .Z(n450) );
  NANDN U523 ( .A(n451), .B(n450), .Z(n452) );
  NANDN U524 ( .A(n453), .B(n452), .Z(n454) );
  OR U525 ( .A(n455), .B(n454), .Z(n456) );
  NANDN U526 ( .A(n457), .B(n456), .Z(n458) );
  NANDN U527 ( .A(n459), .B(n458), .Z(n461) );
  ANDN U528 ( .B(x[65]), .A(y[65]), .Z(n460) );
  OR U529 ( .A(n461), .B(n460), .Z(n462) );
  NANDN U530 ( .A(n463), .B(n462), .Z(n464) );
  NANDN U531 ( .A(n465), .B(n464), .Z(n467) );
  ANDN U532 ( .B(x[67]), .A(y[67]), .Z(n466) );
  OR U533 ( .A(n467), .B(n466), .Z(n468) );
  NANDN U534 ( .A(n469), .B(n468), .Z(n470) );
  NANDN U535 ( .A(n471), .B(n470), .Z(n473) );
  ANDN U536 ( .B(x[69]), .A(y[69]), .Z(n472) );
  OR U537 ( .A(n473), .B(n472), .Z(n474) );
  NANDN U538 ( .A(n475), .B(n474), .Z(n476) );
  NANDN U539 ( .A(n477), .B(n476), .Z(n479) );
  ANDN U540 ( .B(x[71]), .A(y[71]), .Z(n478) );
  OR U541 ( .A(n479), .B(n478), .Z(n480) );
  NANDN U542 ( .A(n481), .B(n480), .Z(n482) );
  NANDN U543 ( .A(n483), .B(n482), .Z(n485) );
  ANDN U544 ( .B(x[73]), .A(y[73]), .Z(n484) );
  OR U545 ( .A(n485), .B(n484), .Z(n486) );
  NANDN U546 ( .A(n487), .B(n486), .Z(n488) );
  NANDN U547 ( .A(n489), .B(n488), .Z(n491) );
  ANDN U548 ( .B(x[75]), .A(y[75]), .Z(n490) );
  OR U549 ( .A(n491), .B(n490), .Z(n492) );
  NANDN U550 ( .A(n493), .B(n492), .Z(n494) );
  NANDN U551 ( .A(n495), .B(n494), .Z(n497) );
  ANDN U552 ( .B(x[77]), .A(y[77]), .Z(n496) );
  OR U553 ( .A(n497), .B(n496), .Z(n498) );
  NANDN U554 ( .A(n499), .B(n498), .Z(n500) );
  NANDN U555 ( .A(n501), .B(n500), .Z(n503) );
  ANDN U556 ( .B(x[79]), .A(y[79]), .Z(n502) );
  OR U557 ( .A(n503), .B(n502), .Z(n504) );
  NANDN U558 ( .A(n505), .B(n504), .Z(n506) );
  NANDN U559 ( .A(n507), .B(n506), .Z(n509) );
  ANDN U560 ( .B(x[81]), .A(y[81]), .Z(n508) );
  OR U561 ( .A(n509), .B(n508), .Z(n510) );
  NANDN U562 ( .A(n511), .B(n510), .Z(n512) );
  NANDN U563 ( .A(n513), .B(n512), .Z(n515) );
  ANDN U564 ( .B(x[83]), .A(y[83]), .Z(n514) );
  OR U565 ( .A(n515), .B(n514), .Z(n516) );
  NANDN U566 ( .A(n517), .B(n516), .Z(n518) );
  NANDN U567 ( .A(n519), .B(n518), .Z(n521) );
  ANDN U568 ( .B(x[85]), .A(y[85]), .Z(n520) );
  OR U569 ( .A(n521), .B(n520), .Z(n522) );
  NANDN U570 ( .A(n523), .B(n522), .Z(n524) );
  NANDN U571 ( .A(n525), .B(n524), .Z(n527) );
  ANDN U572 ( .B(x[87]), .A(y[87]), .Z(n526) );
  OR U573 ( .A(n527), .B(n526), .Z(n528) );
  NANDN U574 ( .A(n529), .B(n528), .Z(n530) );
  NANDN U575 ( .A(n531), .B(n530), .Z(n533) );
  ANDN U576 ( .B(x[89]), .A(y[89]), .Z(n532) );
  OR U577 ( .A(n533), .B(n532), .Z(n534) );
  NANDN U578 ( .A(n535), .B(n534), .Z(n536) );
  NANDN U579 ( .A(n537), .B(n536), .Z(n539) );
  ANDN U580 ( .B(x[91]), .A(y[91]), .Z(n538) );
  OR U581 ( .A(n539), .B(n538), .Z(n540) );
  NANDN U582 ( .A(n541), .B(n540), .Z(n542) );
  NANDN U583 ( .A(n543), .B(n542), .Z(n545) );
  ANDN U584 ( .B(x[93]), .A(y[93]), .Z(n544) );
  OR U585 ( .A(n545), .B(n544), .Z(n546) );
  NANDN U586 ( .A(n547), .B(n546), .Z(n548) );
  NANDN U587 ( .A(n549), .B(n548), .Z(n551) );
  ANDN U588 ( .B(x[95]), .A(y[95]), .Z(n550) );
  OR U589 ( .A(n551), .B(n550), .Z(n552) );
  NANDN U590 ( .A(n553), .B(n552), .Z(n554) );
  NANDN U591 ( .A(n555), .B(n554), .Z(n557) );
  ANDN U592 ( .B(x[97]), .A(y[97]), .Z(n556) );
  OR U593 ( .A(n557), .B(n556), .Z(n558) );
  NANDN U594 ( .A(n559), .B(n558), .Z(n560) );
  NANDN U595 ( .A(n561), .B(n560), .Z(n563) );
  ANDN U596 ( .B(x[99]), .A(y[99]), .Z(n562) );
  OR U597 ( .A(n563), .B(n562), .Z(n564) );
  NANDN U598 ( .A(n565), .B(n564), .Z(n566) );
  NANDN U599 ( .A(n567), .B(n566), .Z(n569) );
  ANDN U600 ( .B(x[101]), .A(y[101]), .Z(n568) );
  OR U601 ( .A(n569), .B(n568), .Z(n570) );
  NANDN U602 ( .A(n571), .B(n570), .Z(n572) );
  NANDN U603 ( .A(n573), .B(n572), .Z(n575) );
  ANDN U604 ( .B(x[103]), .A(y[103]), .Z(n574) );
  OR U605 ( .A(n575), .B(n574), .Z(n576) );
  NANDN U606 ( .A(n577), .B(n576), .Z(n578) );
  NANDN U607 ( .A(n579), .B(n578), .Z(n581) );
  ANDN U608 ( .B(x[105]), .A(y[105]), .Z(n580) );
  OR U609 ( .A(n581), .B(n580), .Z(n582) );
  NANDN U610 ( .A(n583), .B(n582), .Z(n584) );
  NANDN U611 ( .A(n585), .B(n584), .Z(n587) );
  ANDN U612 ( .B(x[107]), .A(y[107]), .Z(n586) );
  OR U613 ( .A(n587), .B(n586), .Z(n588) );
  NANDN U614 ( .A(n589), .B(n588), .Z(n590) );
  NANDN U615 ( .A(n591), .B(n590), .Z(n593) );
  ANDN U616 ( .B(x[109]), .A(y[109]), .Z(n592) );
  OR U617 ( .A(n593), .B(n592), .Z(n594) );
  NANDN U618 ( .A(n595), .B(n594), .Z(n596) );
  NANDN U619 ( .A(n597), .B(n596), .Z(n599) );
  ANDN U620 ( .B(x[111]), .A(y[111]), .Z(n598) );
  OR U621 ( .A(n599), .B(n598), .Z(n600) );
  NANDN U622 ( .A(n601), .B(n600), .Z(n602) );
  NANDN U623 ( .A(n603), .B(n602), .Z(n605) );
  ANDN U624 ( .B(x[113]), .A(y[113]), .Z(n604) );
  OR U625 ( .A(n605), .B(n604), .Z(n606) );
  NANDN U626 ( .A(n607), .B(n606), .Z(n608) );
  NANDN U627 ( .A(n609), .B(n608), .Z(n611) );
  ANDN U628 ( .B(x[115]), .A(y[115]), .Z(n610) );
  OR U629 ( .A(n611), .B(n610), .Z(n612) );
  NANDN U630 ( .A(n613), .B(n612), .Z(n614) );
  NANDN U631 ( .A(n615), .B(n614), .Z(n617) );
  ANDN U632 ( .B(x[117]), .A(y[117]), .Z(n616) );
  OR U633 ( .A(n617), .B(n616), .Z(n618) );
  NANDN U634 ( .A(n619), .B(n618), .Z(n620) );
  NANDN U635 ( .A(n621), .B(n620), .Z(n623) );
  ANDN U636 ( .B(x[119]), .A(y[119]), .Z(n622) );
  OR U637 ( .A(n623), .B(n622), .Z(n624) );
  NANDN U638 ( .A(n625), .B(n624), .Z(n626) );
  NANDN U639 ( .A(n627), .B(n626), .Z(n629) );
  ANDN U640 ( .B(x[121]), .A(y[121]), .Z(n628) );
  OR U641 ( .A(n629), .B(n628), .Z(n630) );
  NANDN U642 ( .A(n631), .B(n630), .Z(n632) );
  NANDN U643 ( .A(n633), .B(n632), .Z(n635) );
  ANDN U644 ( .B(x[123]), .A(y[123]), .Z(n634) );
  OR U645 ( .A(n635), .B(n634), .Z(n636) );
  NANDN U646 ( .A(n637), .B(n636), .Z(n638) );
  NANDN U647 ( .A(n639), .B(n638), .Z(n641) );
  ANDN U648 ( .B(x[125]), .A(y[125]), .Z(n640) );
  OR U649 ( .A(n641), .B(n640), .Z(n642) );
  NANDN U650 ( .A(n643), .B(n642), .Z(n644) );
  NANDN U651 ( .A(n645), .B(n644), .Z(n646) );
  NANDN U652 ( .A(n647), .B(n646), .Z(n649) );
  NAND U653 ( .A(n647), .B(g), .Z(n648) );
  NAND U654 ( .A(n649), .B(n648), .Z(n4) );
endmodule

