
module hamming_N1600_CC4 ( clk, rst, x, y, o );
  input [399:0] x;
  input [399:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  XOR U403 ( .A(n1610), .B(n1608), .Z(n1) );
  NANDN U404 ( .A(n1609), .B(n1), .Z(n2) );
  NAND U405 ( .A(n1610), .B(n1608), .Z(n3) );
  AND U406 ( .A(n2), .B(n3), .Z(n2044) );
  XOR U407 ( .A(n1843), .B(n1841), .Z(n4) );
  NANDN U408 ( .A(n1842), .B(n4), .Z(n5) );
  NAND U409 ( .A(n1843), .B(n1841), .Z(n6) );
  AND U410 ( .A(n5), .B(n6), .Z(n2037) );
  NAND U411 ( .A(n1622), .B(n1623), .Z(n7) );
  XOR U412 ( .A(n1622), .B(n1623), .Z(n8) );
  NANDN U413 ( .A(n1621), .B(n8), .Z(n9) );
  NAND U414 ( .A(n7), .B(n9), .Z(n2060) );
  NAND U415 ( .A(n2033), .B(n2032), .Z(n10) );
  NANDN U416 ( .A(n2033), .B(n2031), .Z(n11) );
  NANDN U417 ( .A(n2034), .B(n11), .Z(n12) );
  NAND U418 ( .A(n10), .B(n12), .Z(n2211) );
  XOR U419 ( .A(n2065), .B(n2063), .Z(n13) );
  NANDN U420 ( .A(n2064), .B(n13), .Z(n14) );
  NAND U421 ( .A(n2065), .B(n2063), .Z(n15) );
  AND U422 ( .A(n14), .B(n15), .Z(n2206) );
  XOR U423 ( .A(n1607), .B(n1605), .Z(n16) );
  NANDN U424 ( .A(n1606), .B(n16), .Z(n17) );
  NAND U425 ( .A(n1607), .B(n1605), .Z(n18) );
  AND U426 ( .A(n17), .B(n18), .Z(n2045) );
  NAND U427 ( .A(n1547), .B(n1548), .Z(n19) );
  XOR U428 ( .A(n1547), .B(n1548), .Z(n20) );
  NANDN U429 ( .A(n1546), .B(n20), .Z(n21) );
  NAND U430 ( .A(n19), .B(n21), .Z(n2035) );
  XOR U431 ( .A(n1698), .B(n1696), .Z(n22) );
  NANDN U432 ( .A(n1697), .B(n22), .Z(n23) );
  NAND U433 ( .A(n1698), .B(n1696), .Z(n24) );
  AND U434 ( .A(n23), .B(n24), .Z(n2063) );
  XOR U435 ( .A(n2043), .B(n2041), .Z(n25) );
  NANDN U436 ( .A(n2042), .B(n25), .Z(n26) );
  NAND U437 ( .A(n2043), .B(n2041), .Z(n27) );
  AND U438 ( .A(n26), .B(n27), .Z(n2213) );
  XOR U439 ( .A(n2037), .B(n2038), .Z(n28) );
  NANDN U440 ( .A(n2039), .B(n28), .Z(n29) );
  NAND U441 ( .A(n2037), .B(n2038), .Z(n30) );
  AND U442 ( .A(n29), .B(n30), .Z(n2209) );
  NAND U443 ( .A(n2061), .B(n2062), .Z(n31) );
  XOR U444 ( .A(n2061), .B(n2062), .Z(n32) );
  NANDN U445 ( .A(n2060), .B(n32), .Z(n33) );
  NAND U446 ( .A(n31), .B(n33), .Z(n2207) );
  NAND U447 ( .A(n1975), .B(n1976), .Z(n34) );
  XOR U448 ( .A(n1975), .B(n1976), .Z(n35) );
  NANDN U449 ( .A(n1974), .B(n35), .Z(n36) );
  NAND U450 ( .A(n34), .B(n36), .Z(n2273) );
  NAND U451 ( .A(n1694), .B(n1695), .Z(n37) );
  XOR U452 ( .A(n1694), .B(n1695), .Z(n38) );
  NANDN U453 ( .A(n1693), .B(n38), .Z(n39) );
  NAND U454 ( .A(n37), .B(n39), .Z(n2064) );
  XOR U455 ( .A(n1620), .B(n1618), .Z(n40) );
  NANDN U456 ( .A(n1619), .B(n40), .Z(n41) );
  NAND U457 ( .A(n1620), .B(n1618), .Z(n42) );
  AND U458 ( .A(n41), .B(n42), .Z(n2061) );
  NAND U459 ( .A(n2045), .B(n2044), .Z(n43) );
  XOR U460 ( .A(n2045), .B(n2044), .Z(n44) );
  NANDN U461 ( .A(n2046), .B(n44), .Z(n45) );
  NAND U462 ( .A(n43), .B(n45), .Z(n2212) );
  XOR U463 ( .A(n2059), .B(n2058), .Z(n46) );
  NAND U464 ( .A(n46), .B(n2057), .Z(n47) );
  NAND U465 ( .A(n2059), .B(n2058), .Z(n48) );
  AND U466 ( .A(n47), .B(n48), .Z(n2208) );
  NAND U467 ( .A(n2210), .B(n2211), .Z(n49) );
  XOR U468 ( .A(n2210), .B(n2211), .Z(n50) );
  NANDN U469 ( .A(n2209), .B(n50), .Z(n51) );
  NAND U470 ( .A(n49), .B(n51), .Z(n2334) );
  XOR U471 ( .A(n2300), .B(n2299), .Z(n2321) );
  XNOR U472 ( .A(n2294), .B(n2293), .Z(n2283) );
  XOR U473 ( .A(n2273), .B(n2272), .Z(n52) );
  NANDN U474 ( .A(n2274), .B(n52), .Z(n53) );
  NAND U475 ( .A(n2273), .B(n2272), .Z(n54) );
  AND U476 ( .A(n53), .B(n54), .Z(n2288) );
  XOR U477 ( .A(n1840), .B(n1838), .Z(n55) );
  NANDN U478 ( .A(n1839), .B(n55), .Z(n56) );
  NAND U479 ( .A(n1840), .B(n1838), .Z(n57) );
  AND U480 ( .A(n56), .B(n57), .Z(n2038) );
  XOR U481 ( .A(oglobal[2]), .B(n2035), .Z(n58) );
  NANDN U482 ( .A(n2036), .B(n58), .Z(n59) );
  NAND U483 ( .A(oglobal[2]), .B(n2035), .Z(n60) );
  AND U484 ( .A(n59), .B(n60), .Z(n2210) );
  NAND U485 ( .A(n2212), .B(n2213), .Z(n61) );
  XOR U486 ( .A(n2212), .B(n2213), .Z(n62) );
  NANDN U487 ( .A(oglobal[3]), .B(n62), .Z(n63) );
  NAND U488 ( .A(n61), .B(n63), .Z(n2333) );
  XNOR U489 ( .A(n1757), .B(n1756), .Z(n1530) );
  NANDN U490 ( .A(n1448), .B(n1447), .Z(n64) );
  NANDN U491 ( .A(n1445), .B(n1446), .Z(n65) );
  AND U492 ( .A(n64), .B(n65), .Z(n1870) );
  NAND U493 ( .A(n2055), .B(n2056), .Z(n66) );
  XOR U494 ( .A(n2055), .B(n2056), .Z(n67) );
  NANDN U495 ( .A(n2054), .B(n67), .Z(n68) );
  NAND U496 ( .A(n66), .B(n68), .Z(n2171) );
  NAND U497 ( .A(n2207), .B(n2208), .Z(n69) );
  XOR U498 ( .A(n2207), .B(n2208), .Z(n70) );
  NANDN U499 ( .A(n2206), .B(n70), .Z(n71) );
  NAND U500 ( .A(n69), .B(n71), .Z(n2335) );
  XOR U501 ( .A(n1638), .B(n1637), .Z(n1639) );
  XOR U502 ( .A(n1990), .B(n1989), .Z(n1991) );
  XNOR U503 ( .A(n2261), .B(n2260), .Z(n2263) );
  NANDN U504 ( .A(n2220), .B(n2223), .Z(n72) );
  OR U505 ( .A(n2223), .B(n2221), .Z(n73) );
  NAND U506 ( .A(n2222), .B(n73), .Z(n74) );
  NAND U507 ( .A(n72), .B(n74), .Z(n2298) );
  XOR U508 ( .A(n1978), .B(n1977), .Z(n1980) );
  NAND U509 ( .A(n2289), .B(n2290), .Z(n75) );
  XOR U510 ( .A(n2289), .B(n2290), .Z(n76) );
  NANDN U511 ( .A(n2288), .B(n76), .Z(n77) );
  NAND U512 ( .A(n75), .B(n77), .Z(n2361) );
  NAND U513 ( .A(n2414), .B(n2415), .Z(n78) );
  XOR U514 ( .A(n2414), .B(n2415), .Z(n79) );
  NANDN U515 ( .A(n2413), .B(n79), .Z(n80) );
  NAND U516 ( .A(n78), .B(n80), .Z(n2423) );
  XOR U517 ( .A(x[338]), .B(y[338]), .Z(n615) );
  XOR U518 ( .A(x[29]), .B(y[29]), .Z(n612) );
  XNOR U519 ( .A(x[340]), .B(y[340]), .Z(n613) );
  XNOR U520 ( .A(n612), .B(n613), .Z(n614) );
  XOR U521 ( .A(n615), .B(n614), .Z(n452) );
  XOR U522 ( .A(x[334]), .B(y[334]), .Z(n567) );
  XOR U523 ( .A(x[336]), .B(y[336]), .Z(n564) );
  XNOR U524 ( .A(x[385]), .B(y[385]), .Z(n565) );
  XNOR U525 ( .A(n564), .B(n565), .Z(n566) );
  XOR U526 ( .A(n567), .B(n566), .Z(n451) );
  XOR U527 ( .A(x[370]), .B(y[370]), .Z(n1063) );
  XOR U528 ( .A(x[13]), .B(y[13]), .Z(n1060) );
  XNOR U529 ( .A(x[372]), .B(y[372]), .Z(n1061) );
  XNOR U530 ( .A(n1060), .B(n1061), .Z(n1062) );
  XNOR U531 ( .A(n1063), .B(n1062), .Z(n450) );
  XOR U532 ( .A(n451), .B(n450), .Z(n453) );
  XOR U533 ( .A(n452), .B(n453), .Z(n585) );
  XOR U534 ( .A(x[362]), .B(y[362]), .Z(n663) );
  XOR U535 ( .A(x[17]), .B(y[17]), .Z(n661) );
  XNOR U536 ( .A(x[364]), .B(y[364]), .Z(n662) );
  XOR U537 ( .A(n661), .B(n662), .Z(n664) );
  XNOR U538 ( .A(n663), .B(n664), .Z(n1266) );
  XOR U539 ( .A(x[366]), .B(y[366]), .Z(n1080) );
  XOR U540 ( .A(x[368]), .B(y[368]), .Z(n1078) );
  XNOR U541 ( .A(x[393]), .B(y[393]), .Z(n1079) );
  XOR U542 ( .A(n1078), .B(n1079), .Z(n1081) );
  XOR U543 ( .A(n1080), .B(n1081), .Z(n1267) );
  XNOR U544 ( .A(n1266), .B(n1267), .Z(n1268) );
  XOR U545 ( .A(x[342]), .B(y[342]), .Z(n494) );
  XOR U546 ( .A(x[344]), .B(y[344]), .Z(n492) );
  XNOR U547 ( .A(x[387]), .B(y[387]), .Z(n493) );
  XOR U548 ( .A(n492), .B(n493), .Z(n495) );
  XOR U549 ( .A(n494), .B(n495), .Z(n1269) );
  XNOR U550 ( .A(n1268), .B(n1269), .Z(n582) );
  XOR U551 ( .A(x[354]), .B(y[354]), .Z(n749) );
  XOR U552 ( .A(x[21]), .B(y[21]), .Z(n747) );
  XNOR U553 ( .A(x[356]), .B(y[356]), .Z(n748) );
  XOR U554 ( .A(n747), .B(n748), .Z(n750) );
  XOR U555 ( .A(n749), .B(n750), .Z(n583) );
  XNOR U556 ( .A(n582), .B(n583), .Z(n584) );
  XOR U557 ( .A(n585), .B(n584), .Z(n857) );
  XOR U558 ( .A(x[310]), .B(y[310]), .Z(n700) );
  XOR U559 ( .A(x[312]), .B(y[312]), .Z(n698) );
  XNOR U560 ( .A(x[379]), .B(y[379]), .Z(n699) );
  XOR U561 ( .A(n698), .B(n699), .Z(n701) );
  XNOR U562 ( .A(n700), .B(n701), .Z(n153) );
  XOR U563 ( .A(x[382]), .B(y[382]), .Z(n1116) );
  XOR U564 ( .A(x[384]), .B(y[384]), .Z(n1114) );
  XNOR U565 ( .A(x[397]), .B(y[397]), .Z(n1115) );
  XOR U566 ( .A(n1114), .B(n1115), .Z(n1117) );
  XOR U567 ( .A(n1116), .B(n1117), .Z(n154) );
  XNOR U568 ( .A(n153), .B(n154), .Z(n156) );
  XOR U569 ( .A(x[314]), .B(y[314]), .Z(n694) );
  XOR U570 ( .A(x[41]), .B(y[41]), .Z(n692) );
  XNOR U571 ( .A(x[316]), .B(y[316]), .Z(n693) );
  XOR U572 ( .A(n692), .B(n693), .Z(n695) );
  XNOR U573 ( .A(n694), .B(n695), .Z(n155) );
  XOR U574 ( .A(n156), .B(n155), .Z(n100) );
  XOR U575 ( .A(x[306]), .B(y[306]), .Z(n531) );
  XOR U576 ( .A(x[45]), .B(y[45]), .Z(n528) );
  XNOR U577 ( .A(x[308]), .B(y[308]), .Z(n529) );
  XNOR U578 ( .A(n528), .B(n529), .Z(n530) );
  XOR U579 ( .A(n531), .B(n530), .Z(n228) );
  XOR U580 ( .A(x[386]), .B(y[386]), .Z(n393) );
  XOR U581 ( .A(x[5]), .B(y[5]), .Z(n390) );
  XNOR U582 ( .A(x[388]), .B(y[388]), .Z(n391) );
  XNOR U583 ( .A(n390), .B(n391), .Z(n392) );
  XOR U584 ( .A(n393), .B(n392), .Z(n226) );
  XOR U585 ( .A(x[302]), .B(y[302]), .Z(n465) );
  XOR U586 ( .A(x[304]), .B(y[304]), .Z(n462) );
  XNOR U587 ( .A(x[377]), .B(y[377]), .Z(n463) );
  XNOR U588 ( .A(n462), .B(n463), .Z(n464) );
  XNOR U589 ( .A(n465), .B(n464), .Z(n225) );
  XNOR U590 ( .A(n226), .B(n225), .Z(n227) );
  XNOR U591 ( .A(n228), .B(n227), .Z(n99) );
  XNOR U592 ( .A(n100), .B(n99), .Z(n101) );
  XOR U593 ( .A(x[298]), .B(y[298]), .Z(n689) );
  XOR U594 ( .A(x[49]), .B(y[49]), .Z(n686) );
  XNOR U595 ( .A(x[300]), .B(y[300]), .Z(n687) );
  XNOR U596 ( .A(n686), .B(n687), .Z(n688) );
  XOR U597 ( .A(n689), .B(n688), .Z(n216) );
  XOR U598 ( .A(x[390]), .B(y[390]), .Z(n338) );
  XOR U599 ( .A(x[392]), .B(y[392]), .Z(n335) );
  XNOR U600 ( .A(x[399]), .B(y[399]), .Z(n336) );
  XNOR U601 ( .A(n335), .B(n336), .Z(n337) );
  XOR U602 ( .A(n338), .B(n337), .Z(n214) );
  XOR U603 ( .A(x[294]), .B(y[294]), .Z(n543) );
  XOR U604 ( .A(x[296]), .B(y[296]), .Z(n540) );
  XNOR U605 ( .A(x[375]), .B(y[375]), .Z(n541) );
  XNOR U606 ( .A(n540), .B(n541), .Z(n542) );
  XNOR U607 ( .A(n543), .B(n542), .Z(n213) );
  XNOR U608 ( .A(n214), .B(n213), .Z(n215) );
  XOR U609 ( .A(n216), .B(n215), .Z(n102) );
  XNOR U610 ( .A(n101), .B(n102), .Z(n856) );
  XOR U611 ( .A(n857), .B(n856), .Z(n859) );
  XOR U612 ( .A(x[318]), .B(y[318]), .Z(n476) );
  XOR U613 ( .A(x[320]), .B(y[320]), .Z(n474) );
  XNOR U614 ( .A(x[381]), .B(y[381]), .Z(n475) );
  XOR U615 ( .A(n474), .B(n475), .Z(n477) );
  XNOR U616 ( .A(n476), .B(n477), .Z(n159) );
  XOR U617 ( .A(x[378]), .B(y[378]), .Z(n1243) );
  XOR U618 ( .A(x[9]), .B(y[9]), .Z(n1241) );
  XNOR U619 ( .A(x[380]), .B(y[380]), .Z(n1242) );
  XOR U620 ( .A(n1241), .B(n1242), .Z(n1244) );
  XOR U621 ( .A(n1243), .B(n1244), .Z(n160) );
  XNOR U622 ( .A(n159), .B(n160), .Z(n162) );
  XOR U623 ( .A(x[322]), .B(y[322]), .Z(n470) );
  XOR U624 ( .A(x[37]), .B(y[37]), .Z(n468) );
  XNOR U625 ( .A(x[324]), .B(y[324]), .Z(n469) );
  XOR U626 ( .A(n468), .B(n469), .Z(n471) );
  XNOR U627 ( .A(n470), .B(n471), .Z(n161) );
  XOR U628 ( .A(n162), .B(n161), .Z(n204) );
  XOR U629 ( .A(x[326]), .B(y[326]), .Z(n639) );
  XOR U630 ( .A(x[328]), .B(y[328]), .Z(n637) );
  XNOR U631 ( .A(x[383]), .B(y[383]), .Z(n638) );
  XOR U632 ( .A(n637), .B(n638), .Z(n640) );
  XNOR U633 ( .A(n639), .B(n640), .Z(n171) );
  XOR U634 ( .A(x[374]), .B(y[374]), .Z(n1044) );
  XOR U635 ( .A(x[376]), .B(y[376]), .Z(n1042) );
  XNOR U636 ( .A(x[395]), .B(y[395]), .Z(n1043) );
  XOR U637 ( .A(n1042), .B(n1043), .Z(n1045) );
  XOR U638 ( .A(n1044), .B(n1045), .Z(n172) );
  XNOR U639 ( .A(n171), .B(n172), .Z(n174) );
  XOR U640 ( .A(x[330]), .B(y[330]), .Z(n633) );
  XOR U641 ( .A(x[33]), .B(y[33]), .Z(n631) );
  XNOR U642 ( .A(x[332]), .B(y[332]), .Z(n632) );
  XOR U643 ( .A(n631), .B(n632), .Z(n634) );
  XNOR U644 ( .A(n633), .B(n634), .Z(n173) );
  XOR U645 ( .A(n174), .B(n173), .Z(n202) );
  XOR U646 ( .A(x[346]), .B(y[346]), .Z(n834) );
  XOR U647 ( .A(x[25]), .B(y[25]), .Z(n832) );
  XNOR U648 ( .A(x[348]), .B(y[348]), .Z(n833) );
  XOR U649 ( .A(n832), .B(n833), .Z(n835) );
  XNOR U650 ( .A(n834), .B(n835), .Z(n1168) );
  XOR U651 ( .A(x[358]), .B(y[358]), .Z(n670) );
  XOR U652 ( .A(x[360]), .B(y[360]), .Z(n668) );
  XNOR U653 ( .A(x[391]), .B(y[391]), .Z(n669) );
  XOR U654 ( .A(n668), .B(n669), .Z(n671) );
  XOR U655 ( .A(n670), .B(n671), .Z(n1169) );
  XNOR U656 ( .A(n1168), .B(n1169), .Z(n1171) );
  XOR U657 ( .A(x[350]), .B(y[350]), .Z(n797) );
  XOR U658 ( .A(x[352]), .B(y[352]), .Z(n795) );
  XNOR U659 ( .A(x[389]), .B(y[389]), .Z(n796) );
  XOR U660 ( .A(n795), .B(n796), .Z(n798) );
  XNOR U661 ( .A(n797), .B(n798), .Z(n1170) );
  XNOR U662 ( .A(n1171), .B(n1170), .Z(n201) );
  XNOR U663 ( .A(n202), .B(n201), .Z(n203) );
  XNOR U664 ( .A(n204), .B(n203), .Z(n858) );
  XOR U665 ( .A(n859), .B(n858), .Z(n724) );
  XOR U666 ( .A(x[0]), .B(y[0]), .Z(n429) );
  XOR U667 ( .A(x[2]), .B(y[2]), .Z(n426) );
  XNOR U668 ( .A(x[4]), .B(y[4]), .Z(n427) );
  XNOR U669 ( .A(n426), .B(n427), .Z(n428) );
  XOR U670 ( .A(n429), .B(n428), .Z(n591) );
  XOR U671 ( .A(x[7]), .B(y[7]), .Z(n417) );
  XOR U672 ( .A(x[1]), .B(y[1]), .Z(n414) );
  XNOR U673 ( .A(x[3]), .B(y[3]), .Z(n415) );
  XNOR U674 ( .A(n414), .B(n415), .Z(n416) );
  XOR U675 ( .A(n417), .B(n416), .Z(n589) );
  XOR U676 ( .A(x[19]), .B(y[19]), .Z(n423) );
  XOR U677 ( .A(x[11]), .B(y[11]), .Z(n420) );
  XNOR U678 ( .A(x[15]), .B(y[15]), .Z(n421) );
  XNOR U679 ( .A(n420), .B(n421), .Z(n422) );
  XNOR U680 ( .A(n423), .B(n422), .Z(n588) );
  XNOR U681 ( .A(n589), .B(n588), .Z(n590) );
  XNOR U682 ( .A(n591), .B(n590), .Z(n1036) );
  XOR U683 ( .A(x[31]), .B(y[31]), .Z(n192) );
  XOR U684 ( .A(x[23]), .B(y[23]), .Z(n189) );
  XNOR U685 ( .A(x[27]), .B(y[27]), .Z(n190) );
  XNOR U686 ( .A(n189), .B(n190), .Z(n191) );
  XOR U687 ( .A(n192), .B(n191), .Z(n489) );
  XOR U688 ( .A(x[43]), .B(y[43]), .Z(n180) );
  XOR U689 ( .A(x[35]), .B(y[35]), .Z(n177) );
  XNOR U690 ( .A(x[39]), .B(y[39]), .Z(n178) );
  XNOR U691 ( .A(n177), .B(n178), .Z(n179) );
  XOR U692 ( .A(n180), .B(n179), .Z(n487) );
  XOR U693 ( .A(x[55]), .B(y[55]), .Z(n186) );
  XOR U694 ( .A(x[47]), .B(y[47]), .Z(n183) );
  XNOR U695 ( .A(x[51]), .B(y[51]), .Z(n184) );
  XNOR U696 ( .A(n183), .B(n184), .Z(n185) );
  XNOR U697 ( .A(n186), .B(n185), .Z(n486) );
  XNOR U698 ( .A(n487), .B(n486), .Z(n488) );
  XOR U699 ( .A(n489), .B(n488), .Z(n1037) );
  XNOR U700 ( .A(n1036), .B(n1037), .Z(n1038) );
  XOR U701 ( .A(x[67]), .B(y[67]), .Z(n1147) );
  XOR U702 ( .A(x[59]), .B(y[59]), .Z(n1144) );
  XNOR U703 ( .A(x[63]), .B(y[63]), .Z(n1145) );
  XNOR U704 ( .A(n1144), .B(n1145), .Z(n1146) );
  XOR U705 ( .A(n1147), .B(n1146), .Z(n829) );
  XOR U706 ( .A(x[79]), .B(y[79]), .Z(n1135) );
  XOR U707 ( .A(x[71]), .B(y[71]), .Z(n1132) );
  XNOR U708 ( .A(x[75]), .B(y[75]), .Z(n1133) );
  XNOR U709 ( .A(n1132), .B(n1133), .Z(n1134) );
  XOR U710 ( .A(n1135), .B(n1134), .Z(n827) );
  XOR U711 ( .A(x[91]), .B(y[91]), .Z(n1214) );
  XOR U712 ( .A(x[83]), .B(y[83]), .Z(n1211) );
  XNOR U713 ( .A(x[87]), .B(y[87]), .Z(n1212) );
  XNOR U714 ( .A(n1211), .B(n1212), .Z(n1213) );
  XNOR U715 ( .A(n1214), .B(n1213), .Z(n826) );
  XNOR U716 ( .A(n827), .B(n826), .Z(n828) );
  XOR U717 ( .A(n829), .B(n828), .Z(n1039) );
  XNOR U718 ( .A(n1038), .B(n1039), .Z(n237) );
  XOR U719 ( .A(x[245]), .B(y[245]), .Z(n888) );
  XOR U720 ( .A(x[243]), .B(y[243]), .Z(n886) );
  XNOR U721 ( .A(x[323]), .B(y[323]), .Z(n887) );
  XOR U722 ( .A(n886), .B(n887), .Z(n889) );
  XNOR U723 ( .A(n888), .B(n889), .Z(n552) );
  XOR U724 ( .A(x[241]), .B(y[241]), .Z(n936) );
  XOR U725 ( .A(x[239]), .B(y[239]), .Z(n934) );
  XNOR U726 ( .A(x[325]), .B(y[325]), .Z(n935) );
  XOR U727 ( .A(n934), .B(n935), .Z(n937) );
  XOR U728 ( .A(n936), .B(n937), .Z(n553) );
  XNOR U729 ( .A(n552), .B(n553), .Z(n555) );
  XOR U730 ( .A(x[237]), .B(y[237]), .Z(n930) );
  XOR U731 ( .A(x[235]), .B(y[235]), .Z(n928) );
  XNOR U732 ( .A(x[327]), .B(y[327]), .Z(n929) );
  XOR U733 ( .A(n928), .B(n929), .Z(n931) );
  XNOR U734 ( .A(n930), .B(n931), .Z(n554) );
  XOR U735 ( .A(n555), .B(n554), .Z(n823) );
  XOR U736 ( .A(x[269]), .B(y[269]), .Z(n978) );
  XOR U737 ( .A(x[267]), .B(y[267]), .Z(n976) );
  XNOR U738 ( .A(x[311]), .B(y[311]), .Z(n977) );
  XOR U739 ( .A(n976), .B(n977), .Z(n979) );
  XNOR U740 ( .A(n978), .B(n979), .Z(n741) );
  XOR U741 ( .A(x[265]), .B(y[265]), .Z(n990) );
  XOR U742 ( .A(x[263]), .B(y[263]), .Z(n988) );
  XNOR U743 ( .A(x[313]), .B(y[313]), .Z(n989) );
  XOR U744 ( .A(n988), .B(n989), .Z(n991) );
  XOR U745 ( .A(n990), .B(n991), .Z(n742) );
  XNOR U746 ( .A(n741), .B(n742), .Z(n744) );
  XOR U747 ( .A(x[261]), .B(y[261]), .Z(n984) );
  XOR U748 ( .A(x[259]), .B(y[259]), .Z(n982) );
  XNOR U749 ( .A(x[315]), .B(y[315]), .Z(n983) );
  XOR U750 ( .A(n982), .B(n983), .Z(n985) );
  XNOR U751 ( .A(n984), .B(n985), .Z(n743) );
  XOR U752 ( .A(n744), .B(n743), .Z(n821) );
  XOR U753 ( .A(x[257]), .B(y[257]), .Z(n996) );
  XOR U754 ( .A(x[255]), .B(y[255]), .Z(n994) );
  XNOR U755 ( .A(x[317]), .B(y[317]), .Z(n995) );
  XOR U756 ( .A(n994), .B(n995), .Z(n997) );
  XNOR U757 ( .A(n996), .B(n997), .Z(n594) );
  XOR U758 ( .A(x[253]), .B(y[253]), .Z(n882) );
  XOR U759 ( .A(x[251]), .B(y[251]), .Z(n880) );
  XNOR U760 ( .A(x[319]), .B(y[319]), .Z(n881) );
  XOR U761 ( .A(n880), .B(n881), .Z(n883) );
  XOR U762 ( .A(n882), .B(n883), .Z(n595) );
  XNOR U763 ( .A(n594), .B(n595), .Z(n597) );
  XOR U764 ( .A(x[249]), .B(y[249]), .Z(n876) );
  XOR U765 ( .A(x[247]), .B(y[247]), .Z(n874) );
  XNOR U766 ( .A(x[321]), .B(y[321]), .Z(n875) );
  XOR U767 ( .A(n874), .B(n875), .Z(n877) );
  XNOR U768 ( .A(n876), .B(n877), .Z(n596) );
  XNOR U769 ( .A(n597), .B(n596), .Z(n820) );
  XNOR U770 ( .A(n821), .B(n820), .Z(n822) );
  XOR U771 ( .A(n823), .B(n822), .Z(n238) );
  XNOR U772 ( .A(n237), .B(n238), .Z(n240) );
  XOR U773 ( .A(x[24]), .B(y[24]), .Z(n374) );
  XOR U774 ( .A(x[26]), .B(y[26]), .Z(n372) );
  XNOR U775 ( .A(x[28]), .B(y[28]), .Z(n373) );
  XOR U776 ( .A(n372), .B(n373), .Z(n375) );
  XNOR U777 ( .A(n374), .B(n375), .Z(n783) );
  XOR U778 ( .A(x[30]), .B(y[30]), .Z(n380) );
  XOR U779 ( .A(x[32]), .B(y[32]), .Z(n378) );
  XNOR U780 ( .A(x[34]), .B(y[34]), .Z(n379) );
  XOR U781 ( .A(n378), .B(n379), .Z(n381) );
  XOR U782 ( .A(n380), .B(n381), .Z(n784) );
  XNOR U783 ( .A(n783), .B(n784), .Z(n786) );
  XOR U784 ( .A(x[36]), .B(y[36]), .Z(n386) );
  XOR U785 ( .A(x[38]), .B(y[38]), .Z(n384) );
  XNOR U786 ( .A(x[40]), .B(y[40]), .Z(n385) );
  XOR U787 ( .A(n384), .B(n385), .Z(n387) );
  XNOR U788 ( .A(n386), .B(n387), .Z(n785) );
  XOR U789 ( .A(n786), .B(n785), .Z(n772) );
  XOR U790 ( .A(x[54]), .B(y[54]), .Z(n363) );
  XOR U791 ( .A(x[56]), .B(y[56]), .Z(n360) );
  XNOR U792 ( .A(x[58]), .B(y[58]), .Z(n361) );
  XNOR U793 ( .A(n360), .B(n361), .Z(n362) );
  XOR U794 ( .A(n363), .B(n362), .Z(n853) );
  XOR U795 ( .A(x[48]), .B(y[48]), .Z(n351) );
  XOR U796 ( .A(x[50]), .B(y[50]), .Z(n348) );
  XNOR U797 ( .A(x[52]), .B(y[52]), .Z(n349) );
  XNOR U798 ( .A(n348), .B(n349), .Z(n350) );
  XOR U799 ( .A(n351), .B(n350), .Z(n851) );
  XOR U800 ( .A(x[42]), .B(y[42]), .Z(n357) );
  XOR U801 ( .A(x[44]), .B(y[44]), .Z(n354) );
  XNOR U802 ( .A(x[46]), .B(y[46]), .Z(n355) );
  XNOR U803 ( .A(n354), .B(n355), .Z(n356) );
  XNOR U804 ( .A(n357), .B(n356), .Z(n850) );
  XNOR U805 ( .A(n851), .B(n850), .Z(n852) );
  XNOR U806 ( .A(n853), .B(n852), .Z(n771) );
  XNOR U807 ( .A(n772), .B(n771), .Z(n773) );
  XOR U808 ( .A(x[18]), .B(y[18]), .Z(n447) );
  XOR U809 ( .A(x[20]), .B(y[20]), .Z(n444) );
  XNOR U810 ( .A(x[22]), .B(y[22]), .Z(n445) );
  XNOR U811 ( .A(n444), .B(n445), .Z(n446) );
  XOR U812 ( .A(n447), .B(n446), .Z(n513) );
  XOR U813 ( .A(x[12]), .B(y[12]), .Z(n435) );
  XOR U814 ( .A(x[14]), .B(y[14]), .Z(n432) );
  XNOR U815 ( .A(x[16]), .B(y[16]), .Z(n433) );
  XNOR U816 ( .A(n432), .B(n433), .Z(n434) );
  XOR U817 ( .A(n435), .B(n434), .Z(n511) );
  XOR U818 ( .A(x[6]), .B(y[6]), .Z(n441) );
  XOR U819 ( .A(x[8]), .B(y[8]), .Z(n438) );
  XNOR U820 ( .A(x[10]), .B(y[10]), .Z(n439) );
  XNOR U821 ( .A(n438), .B(n439), .Z(n440) );
  XNOR U822 ( .A(n441), .B(n440), .Z(n510) );
  XNOR U823 ( .A(n511), .B(n510), .Z(n512) );
  XOR U824 ( .A(n513), .B(n512), .Z(n774) );
  XNOR U825 ( .A(n773), .B(n774), .Z(n239) );
  XNOR U826 ( .A(n240), .B(n239), .Z(n723) );
  XNOR U827 ( .A(n724), .B(n723), .Z(n726) );
  XOR U828 ( .A(x[154]), .B(y[154]), .Z(n1050) );
  XOR U829 ( .A(x[156]), .B(y[156]), .Z(n1048) );
  XNOR U830 ( .A(x[341]), .B(y[341]), .Z(n1049) );
  XOR U831 ( .A(n1048), .B(n1049), .Z(n1051) );
  XNOR U832 ( .A(n1050), .B(n1051), .Z(n219) );
  XOR U833 ( .A(x[158]), .B(y[158]), .Z(n1056) );
  XOR U834 ( .A(x[117]), .B(y[117]), .Z(n1054) );
  XNOR U835 ( .A(x[160]), .B(y[160]), .Z(n1055) );
  XOR U836 ( .A(n1054), .B(n1055), .Z(n1057) );
  XOR U837 ( .A(n1056), .B(n1057), .Z(n220) );
  XNOR U838 ( .A(n219), .B(n220), .Z(n222) );
  XOR U839 ( .A(x[162]), .B(y[162]), .Z(n1068) );
  XOR U840 ( .A(x[164]), .B(y[164]), .Z(n1066) );
  XNOR U841 ( .A(x[343]), .B(y[343]), .Z(n1067) );
  XOR U842 ( .A(n1066), .B(n1067), .Z(n1069) );
  XNOR U843 ( .A(n1068), .B(n1069), .Z(n221) );
  XOR U844 ( .A(n222), .B(n221), .Z(n817) );
  XOR U845 ( .A(x[166]), .B(y[166]), .Z(n1074) );
  XOR U846 ( .A(x[113]), .B(y[113]), .Z(n1072) );
  XNOR U847 ( .A(x[168]), .B(y[168]), .Z(n1073) );
  XOR U848 ( .A(n1072), .B(n1073), .Z(n1075) );
  XNOR U849 ( .A(n1074), .B(n1075), .Z(n87) );
  XOR U850 ( .A(x[170]), .B(y[170]), .Z(n1086) );
  XOR U851 ( .A(x[172]), .B(y[172]), .Z(n1084) );
  XNOR U852 ( .A(x[345]), .B(y[345]), .Z(n1085) );
  XOR U853 ( .A(n1084), .B(n1085), .Z(n1087) );
  XOR U854 ( .A(n1086), .B(n1087), .Z(n88) );
  XNOR U855 ( .A(n87), .B(n88), .Z(n90) );
  XOR U856 ( .A(x[174]), .B(y[174]), .Z(n1092) );
  XOR U857 ( .A(x[109]), .B(y[109]), .Z(n1090) );
  XNOR U858 ( .A(x[176]), .B(y[176]), .Z(n1091) );
  XOR U859 ( .A(n1090), .B(n1091), .Z(n1093) );
  XNOR U860 ( .A(n1092), .B(n1093), .Z(n89) );
  XOR U861 ( .A(n90), .B(n89), .Z(n815) );
  XOR U862 ( .A(x[186]), .B(y[186]), .Z(n961) );
  XOR U863 ( .A(x[188]), .B(y[188]), .Z(n958) );
  XNOR U864 ( .A(x[349]), .B(y[349]), .Z(n959) );
  XNOR U865 ( .A(n958), .B(n959), .Z(n960) );
  XOR U866 ( .A(n961), .B(n960), .Z(n108) );
  XOR U867 ( .A(x[182]), .B(y[182]), .Z(n652) );
  XOR U868 ( .A(x[105]), .B(y[105]), .Z(n649) );
  XNOR U869 ( .A(x[184]), .B(y[184]), .Z(n650) );
  XNOR U870 ( .A(n649), .B(n650), .Z(n651) );
  XOR U871 ( .A(n652), .B(n651), .Z(n106) );
  XOR U872 ( .A(x[178]), .B(y[178]), .Z(n658) );
  XOR U873 ( .A(x[180]), .B(y[180]), .Z(n655) );
  XNOR U874 ( .A(x[347]), .B(y[347]), .Z(n656) );
  XNOR U875 ( .A(n655), .B(n656), .Z(n657) );
  XNOR U876 ( .A(n658), .B(n657), .Z(n105) );
  XNOR U877 ( .A(n106), .B(n105), .Z(n107) );
  XNOR U878 ( .A(n108), .B(n107), .Z(n814) );
  XNOR U879 ( .A(n815), .B(n814), .Z(n816) );
  XNOR U880 ( .A(n817), .B(n816), .Z(n234) );
  XOR U881 ( .A(x[150]), .B(y[150]), .Z(n1232) );
  XOR U882 ( .A(x[121]), .B(y[121]), .Z(n1229) );
  XNOR U883 ( .A(x[152]), .B(y[152]), .Z(n1230) );
  XNOR U884 ( .A(n1229), .B(n1230), .Z(n1231) );
  XOR U885 ( .A(n1232), .B(n1231), .Z(n168) );
  XOR U886 ( .A(x[146]), .B(y[146]), .Z(n1238) );
  XOR U887 ( .A(x[148]), .B(y[148]), .Z(n1235) );
  XNOR U888 ( .A(x[339]), .B(y[339]), .Z(n1236) );
  XNOR U889 ( .A(n1235), .B(n1236), .Z(n1237) );
  XOR U890 ( .A(n1238), .B(n1237), .Z(n166) );
  XOR U891 ( .A(x[142]), .B(y[142]), .Z(n1129) );
  XOR U892 ( .A(x[125]), .B(y[125]), .Z(n1126) );
  XNOR U893 ( .A(x[144]), .B(y[144]), .Z(n1127) );
  XNOR U894 ( .A(n1126), .B(n1127), .Z(n1128) );
  XNOR U895 ( .A(n1129), .B(n1128), .Z(n165) );
  XNOR U896 ( .A(n166), .B(n165), .Z(n167) );
  XNOR U897 ( .A(n168), .B(n167), .Z(n705) );
  XOR U898 ( .A(x[138]), .B(y[138]), .Z(n1123) );
  XOR U899 ( .A(x[140]), .B(y[140]), .Z(n1120) );
  XNOR U900 ( .A(x[337]), .B(y[337]), .Z(n1121) );
  XNOR U901 ( .A(n1120), .B(n1121), .Z(n1122) );
  XOR U902 ( .A(n1123), .B(n1122), .Z(n198) );
  XOR U903 ( .A(x[134]), .B(y[134]), .Z(n405) );
  XOR U904 ( .A(x[129]), .B(y[129]), .Z(n402) );
  XNOR U905 ( .A(x[136]), .B(y[136]), .Z(n403) );
  XNOR U906 ( .A(n402), .B(n403), .Z(n404) );
  XOR U907 ( .A(n405), .B(n404), .Z(n196) );
  XOR U908 ( .A(x[130]), .B(y[130]), .Z(n399) );
  XOR U909 ( .A(x[132]), .B(y[132]), .Z(n396) );
  XNOR U910 ( .A(x[335]), .B(y[335]), .Z(n397) );
  XNOR U911 ( .A(n396), .B(n397), .Z(n398) );
  XNOR U912 ( .A(n399), .B(n398), .Z(n195) );
  XNOR U913 ( .A(n196), .B(n195), .Z(n197) );
  XOR U914 ( .A(n198), .B(n197), .Z(n706) );
  XNOR U915 ( .A(n705), .B(n706), .Z(n707) );
  XOR U916 ( .A(x[126]), .B(y[126]), .Z(n332) );
  XOR U917 ( .A(x[128]), .B(y[128]), .Z(n329) );
  XNOR U918 ( .A(x[133]), .B(y[133]), .Z(n330) );
  XNOR U919 ( .A(n329), .B(n330), .Z(n331) );
  XOR U920 ( .A(n332), .B(n331), .Z(n252) );
  XOR U921 ( .A(x[120]), .B(y[120]), .Z(n344) );
  XOR U922 ( .A(x[122]), .B(y[122]), .Z(n341) );
  XNOR U923 ( .A(x[124]), .B(y[124]), .Z(n342) );
  XNOR U924 ( .A(n341), .B(n342), .Z(n343) );
  XOR U925 ( .A(n344), .B(n343), .Z(n250) );
  XOR U926 ( .A(x[114]), .B(y[114]), .Z(n1281) );
  XOR U927 ( .A(x[116]), .B(y[116]), .Z(n1278) );
  XNOR U928 ( .A(x[118]), .B(y[118]), .Z(n1279) );
  XNOR U929 ( .A(n1278), .B(n1279), .Z(n1280) );
  XNOR U930 ( .A(n1281), .B(n1280), .Z(n249) );
  XNOR U931 ( .A(n250), .B(n249), .Z(n251) );
  XOR U932 ( .A(n252), .B(n251), .Z(n708) );
  XNOR U933 ( .A(n707), .B(n708), .Z(n231) );
  XOR U934 ( .A(x[78]), .B(y[78]), .Z(n1158) );
  XOR U935 ( .A(x[80]), .B(y[80]), .Z(n1156) );
  XNOR U936 ( .A(x[82]), .B(y[82]), .Z(n1157) );
  XOR U937 ( .A(n1156), .B(n1157), .Z(n1159) );
  XNOR U938 ( .A(n1158), .B(n1159), .Z(n366) );
  XOR U939 ( .A(x[84]), .B(y[84]), .Z(n1152) );
  XOR U940 ( .A(x[86]), .B(y[86]), .Z(n1150) );
  XNOR U941 ( .A(x[88]), .B(y[88]), .Z(n1151) );
  XOR U942 ( .A(n1150), .B(n1151), .Z(n1153) );
  XOR U943 ( .A(n1152), .B(n1153), .Z(n367) );
  XNOR U944 ( .A(n366), .B(n367), .Z(n369) );
  XOR U945 ( .A(x[90]), .B(y[90]), .Z(n1164) );
  XOR U946 ( .A(x[92]), .B(y[92]), .Z(n1162) );
  XNOR U947 ( .A(x[94]), .B(y[94]), .Z(n1163) );
  XOR U948 ( .A(n1162), .B(n1163), .Z(n1165) );
  XNOR U949 ( .A(n1164), .B(n1165), .Z(n368) );
  XOR U950 ( .A(n369), .B(n368), .Z(n712) );
  XOR U951 ( .A(x[108]), .B(y[108]), .Z(n1275) );
  XOR U952 ( .A(x[110]), .B(y[110]), .Z(n1272) );
  XNOR U953 ( .A(x[112]), .B(y[112]), .Z(n1273) );
  XNOR U954 ( .A(n1272), .B(n1273), .Z(n1274) );
  XOR U955 ( .A(n1275), .B(n1274), .Z(n326) );
  XOR U956 ( .A(x[102]), .B(y[102]), .Z(n1208) );
  XOR U957 ( .A(x[104]), .B(y[104]), .Z(n1205) );
  XNOR U958 ( .A(x[106]), .B(y[106]), .Z(n1206) );
  XNOR U959 ( .A(n1205), .B(n1206), .Z(n1207) );
  XOR U960 ( .A(n1208), .B(n1207), .Z(n324) );
  XOR U961 ( .A(x[96]), .B(y[96]), .Z(n1202) );
  XOR U962 ( .A(x[98]), .B(y[98]), .Z(n1199) );
  XNOR U963 ( .A(x[100]), .B(y[100]), .Z(n1200) );
  XNOR U964 ( .A(n1199), .B(n1200), .Z(n1201) );
  XNOR U965 ( .A(n1202), .B(n1201), .Z(n323) );
  XNOR U966 ( .A(n324), .B(n323), .Z(n325) );
  XNOR U967 ( .A(n326), .B(n325), .Z(n711) );
  XNOR U968 ( .A(n712), .B(n711), .Z(n713) );
  XOR U969 ( .A(x[72]), .B(y[72]), .Z(n1263) );
  XOR U970 ( .A(x[74]), .B(y[74]), .Z(n1260) );
  XNOR U971 ( .A(x[76]), .B(y[76]), .Z(n1261) );
  XNOR U972 ( .A(n1260), .B(n1261), .Z(n1262) );
  XOR U973 ( .A(n1263), .B(n1262), .Z(n780) );
  XOR U974 ( .A(x[66]), .B(y[66]), .Z(n1251) );
  XOR U975 ( .A(x[68]), .B(y[68]), .Z(n1248) );
  XNOR U976 ( .A(x[70]), .B(y[70]), .Z(n1249) );
  XNOR U977 ( .A(n1248), .B(n1249), .Z(n1250) );
  XOR U978 ( .A(n1251), .B(n1250), .Z(n778) );
  XOR U979 ( .A(x[60]), .B(y[60]), .Z(n1257) );
  XOR U980 ( .A(x[62]), .B(y[62]), .Z(n1254) );
  XNOR U981 ( .A(x[64]), .B(y[64]), .Z(n1255) );
  XNOR U982 ( .A(n1254), .B(n1255), .Z(n1256) );
  XNOR U983 ( .A(n1257), .B(n1256), .Z(n777) );
  XNOR U984 ( .A(n778), .B(n777), .Z(n779) );
  XOR U985 ( .A(n780), .B(n779), .Z(n714) );
  XOR U986 ( .A(n713), .B(n714), .Z(n232) );
  XNOR U987 ( .A(n231), .B(n232), .Z(n233) );
  XOR U988 ( .A(n234), .B(n233), .Z(n718) );
  XOR U989 ( .A(x[278]), .B(y[278]), .Z(n572) );
  XOR U990 ( .A(x[280]), .B(y[280]), .Z(n570) );
  XNOR U991 ( .A(x[371]), .B(y[371]), .Z(n571) );
  XOR U992 ( .A(n570), .B(n571), .Z(n573) );
  XNOR U993 ( .A(n572), .B(n573), .Z(n81) );
  XOR U994 ( .A(x[194]), .B(y[194]), .Z(n1195) );
  XOR U995 ( .A(x[196]), .B(y[196]), .Z(n1193) );
  XNOR U996 ( .A(x[398]), .B(y[398]), .Z(n1194) );
  XOR U997 ( .A(n1193), .B(n1194), .Z(n1196) );
  XOR U998 ( .A(n1195), .B(n1196), .Z(n82) );
  XNOR U999 ( .A(n81), .B(n82), .Z(n84) );
  XOR U1000 ( .A(x[282]), .B(y[282]), .Z(n536) );
  XOR U1001 ( .A(x[57]), .B(y[57]), .Z(n534) );
  XNOR U1002 ( .A(x[284]), .B(y[284]), .Z(n535) );
  XOR U1003 ( .A(n534), .B(n535), .Z(n537) );
  XNOR U1004 ( .A(n536), .B(n537), .Z(n83) );
  XOR U1005 ( .A(n84), .B(n83), .Z(n208) );
  XOR U1006 ( .A(x[286]), .B(y[286]), .Z(n627) );
  XOR U1007 ( .A(x[288]), .B(y[288]), .Z(n625) );
  XNOR U1008 ( .A(x[373]), .B(y[373]), .Z(n626) );
  XOR U1009 ( .A(n625), .B(n626), .Z(n628) );
  XNOR U1010 ( .A(n627), .B(n628), .Z(n93) );
  XOR U1011 ( .A(x[394]), .B(y[394]), .Z(n1285) );
  XNOR U1012 ( .A(x[396]), .B(y[396]), .Z(n1284) );
  XOR U1013 ( .A(oglobal[0]), .B(n1284), .Z(n1286) );
  XOR U1014 ( .A(n1285), .B(n1286), .Z(n94) );
  XNOR U1015 ( .A(n93), .B(n94), .Z(n96) );
  XOR U1016 ( .A(x[290]), .B(y[290]), .Z(n560) );
  XOR U1017 ( .A(x[53]), .B(y[53]), .Z(n558) );
  XNOR U1018 ( .A(x[292]), .B(y[292]), .Z(n559) );
  XOR U1019 ( .A(n558), .B(n559), .Z(n561) );
  XNOR U1020 ( .A(n560), .B(n561), .Z(n95) );
  XNOR U1021 ( .A(n96), .B(n95), .Z(n207) );
  XNOR U1022 ( .A(n208), .B(n207), .Z(n210) );
  XOR U1023 ( .A(x[274]), .B(y[274]), .Z(n603) );
  XOR U1024 ( .A(x[61]), .B(y[61]), .Z(n600) );
  XNOR U1025 ( .A(x[276]), .B(y[276]), .Z(n601) );
  XNOR U1026 ( .A(n600), .B(n601), .Z(n602) );
  XOR U1027 ( .A(n603), .B(n602), .Z(n114) );
  XOR U1028 ( .A(x[270]), .B(y[270]), .Z(n609) );
  XOR U1029 ( .A(x[272]), .B(y[272]), .Z(n606) );
  XNOR U1030 ( .A(x[369]), .B(y[369]), .Z(n607) );
  XNOR U1031 ( .A(n606), .B(n607), .Z(n608) );
  XOR U1032 ( .A(n609), .B(n608), .Z(n112) );
  XOR U1033 ( .A(x[266]), .B(y[266]), .Z(n507) );
  XOR U1034 ( .A(x[65]), .B(y[65]), .Z(n504) );
  XNOR U1035 ( .A(x[268]), .B(y[268]), .Z(n505) );
  XNOR U1036 ( .A(n504), .B(n505), .Z(n506) );
  XNOR U1037 ( .A(n507), .B(n506), .Z(n111) );
  XNOR U1038 ( .A(n112), .B(n111), .Z(n113) );
  XNOR U1039 ( .A(n114), .B(n113), .Z(n209) );
  XOR U1040 ( .A(n210), .B(n209), .Z(n871) );
  XOR U1041 ( .A(x[262]), .B(y[262]), .Z(n501) );
  XOR U1042 ( .A(x[264]), .B(y[264]), .Z(n498) );
  XNOR U1043 ( .A(x[367]), .B(y[367]), .Z(n499) );
  XNOR U1044 ( .A(n498), .B(n499), .Z(n500) );
  XOR U1045 ( .A(n501), .B(n500), .Z(n150) );
  XOR U1046 ( .A(x[258]), .B(y[258]), .Z(n847) );
  XOR U1047 ( .A(x[69]), .B(y[69]), .Z(n844) );
  XNOR U1048 ( .A(x[260]), .B(y[260]), .Z(n845) );
  XNOR U1049 ( .A(n844), .B(n845), .Z(n846) );
  XOR U1050 ( .A(n847), .B(n846), .Z(n148) );
  XOR U1051 ( .A(x[254]), .B(y[254]), .Z(n841) );
  XOR U1052 ( .A(x[256]), .B(y[256]), .Z(n838) );
  XNOR U1053 ( .A(x[365]), .B(y[365]), .Z(n839) );
  XNOR U1054 ( .A(n838), .B(n839), .Z(n840) );
  XNOR U1055 ( .A(n841), .B(n840), .Z(n147) );
  XNOR U1056 ( .A(n148), .B(n147), .Z(n149) );
  XNOR U1057 ( .A(n150), .B(n149), .Z(n243) );
  XOR U1058 ( .A(x[250]), .B(y[250]), .Z(n792) );
  XOR U1059 ( .A(x[73]), .B(y[73]), .Z(n789) );
  XNOR U1060 ( .A(x[252]), .B(y[252]), .Z(n790) );
  XNOR U1061 ( .A(n789), .B(n790), .Z(n791) );
  XOR U1062 ( .A(n792), .B(n791), .Z(n138) );
  XOR U1063 ( .A(x[246]), .B(y[246]), .Z(n804) );
  XOR U1064 ( .A(x[248]), .B(y[248]), .Z(n801) );
  XNOR U1065 ( .A(x[363]), .B(y[363]), .Z(n802) );
  XNOR U1066 ( .A(n801), .B(n802), .Z(n803) );
  XOR U1067 ( .A(n804), .B(n803), .Z(n136) );
  XOR U1068 ( .A(x[242]), .B(y[242]), .Z(n762) );
  XOR U1069 ( .A(x[77]), .B(y[77]), .Z(n759) );
  XNOR U1070 ( .A(x[244]), .B(y[244]), .Z(n760) );
  XNOR U1071 ( .A(n759), .B(n760), .Z(n761) );
  XNOR U1072 ( .A(n762), .B(n761), .Z(n135) );
  XNOR U1073 ( .A(n136), .B(n135), .Z(n137) );
  XOR U1074 ( .A(n138), .B(n137), .Z(n244) );
  XNOR U1075 ( .A(n243), .B(n244), .Z(n246) );
  XOR U1076 ( .A(x[238]), .B(y[238]), .Z(n756) );
  XOR U1077 ( .A(x[240]), .B(y[240]), .Z(n753) );
  XNOR U1078 ( .A(x[361]), .B(y[361]), .Z(n754) );
  XNOR U1079 ( .A(n753), .B(n754), .Z(n755) );
  XOR U1080 ( .A(n756), .B(n755), .Z(n144) );
  XOR U1081 ( .A(x[234]), .B(y[234]), .Z(n683) );
  XOR U1082 ( .A(x[81]), .B(y[81]), .Z(n681) );
  XOR U1083 ( .A(x[236]), .B(y[236]), .Z(n680) );
  XOR U1084 ( .A(n681), .B(n680), .Z(n682) );
  XOR U1085 ( .A(n683), .B(n682), .Z(n142) );
  XOR U1086 ( .A(x[230]), .B(y[230]), .Z(n677) );
  XOR U1087 ( .A(x[232]), .B(y[232]), .Z(n675) );
  XOR U1088 ( .A(x[359]), .B(y[359]), .Z(n674) );
  XOR U1089 ( .A(n675), .B(n674), .Z(n676) );
  XNOR U1090 ( .A(n677), .B(n676), .Z(n141) );
  XNOR U1091 ( .A(n142), .B(n141), .Z(n143) );
  XNOR U1092 ( .A(n144), .B(n143), .Z(n245) );
  XOR U1093 ( .A(n246), .B(n245), .Z(n869) );
  XOR U1094 ( .A(x[226]), .B(y[226]), .Z(n1220) );
  XOR U1095 ( .A(x[85]), .B(y[85]), .Z(n1217) );
  XNOR U1096 ( .A(x[228]), .B(y[228]), .Z(n1218) );
  XNOR U1097 ( .A(n1217), .B(n1218), .Z(n1219) );
  XOR U1098 ( .A(n1220), .B(n1219), .Z(n126) );
  XOR U1099 ( .A(x[222]), .B(y[222]), .Z(n1226) );
  XOR U1100 ( .A(x[224]), .B(y[224]), .Z(n1223) );
  XNOR U1101 ( .A(x[357]), .B(y[357]), .Z(n1224) );
  XNOR U1102 ( .A(n1223), .B(n1224), .Z(n1225) );
  XOR U1103 ( .A(n1226), .B(n1225), .Z(n124) );
  XOR U1104 ( .A(x[218]), .B(y[218]), .Z(n313) );
  XOR U1105 ( .A(x[89]), .B(y[89]), .Z(n310) );
  XNOR U1106 ( .A(x[220]), .B(y[220]), .Z(n311) );
  XNOR U1107 ( .A(n310), .B(n311), .Z(n312) );
  XNOR U1108 ( .A(n313), .B(n312), .Z(n123) );
  XNOR U1109 ( .A(n124), .B(n123), .Z(n125) );
  XNOR U1110 ( .A(n126), .B(n125), .Z(n516) );
  XOR U1111 ( .A(x[214]), .B(y[214]), .Z(n1183) );
  XOR U1112 ( .A(x[216]), .B(y[216]), .Z(n1180) );
  XNOR U1113 ( .A(x[355]), .B(y[355]), .Z(n1181) );
  XNOR U1114 ( .A(n1180), .B(n1181), .Z(n1182) );
  XOR U1115 ( .A(n1183), .B(n1182), .Z(n132) );
  XOR U1116 ( .A(x[210]), .B(y[210]), .Z(n907) );
  XOR U1117 ( .A(x[93]), .B(y[93]), .Z(n904) );
  XNOR U1118 ( .A(x[212]), .B(y[212]), .Z(n905) );
  XNOR U1119 ( .A(n904), .B(n905), .Z(n906) );
  XOR U1120 ( .A(n907), .B(n906), .Z(n130) );
  XOR U1121 ( .A(x[206]), .B(y[206]), .Z(n1177) );
  XOR U1122 ( .A(x[208]), .B(y[208]), .Z(n1174) );
  XNOR U1123 ( .A(x[353]), .B(y[353]), .Z(n1175) );
  XNOR U1124 ( .A(n1174), .B(n1175), .Z(n1176) );
  XNOR U1125 ( .A(n1177), .B(n1176), .Z(n129) );
  XNOR U1126 ( .A(n130), .B(n129), .Z(n131) );
  XOR U1127 ( .A(n132), .B(n131), .Z(n517) );
  XNOR U1128 ( .A(n516), .B(n517), .Z(n519) );
  XOR U1129 ( .A(x[202]), .B(y[202]), .Z(n955) );
  XOR U1130 ( .A(x[97]), .B(y[97]), .Z(n952) );
  XNOR U1131 ( .A(x[204]), .B(y[204]), .Z(n953) );
  XNOR U1132 ( .A(n952), .B(n953), .Z(n954) );
  XOR U1133 ( .A(n955), .B(n954), .Z(n120) );
  XOR U1134 ( .A(x[198]), .B(y[198]), .Z(n1015) );
  XOR U1135 ( .A(x[200]), .B(y[200]), .Z(n1012) );
  XNOR U1136 ( .A(x[351]), .B(y[351]), .Z(n1013) );
  XNOR U1137 ( .A(n1012), .B(n1013), .Z(n1014) );
  XOR U1138 ( .A(n1015), .B(n1014), .Z(n118) );
  XOR U1139 ( .A(x[190]), .B(y[190]), .Z(n1009) );
  XOR U1140 ( .A(x[101]), .B(y[101]), .Z(n1006) );
  XNOR U1141 ( .A(x[192]), .B(y[192]), .Z(n1007) );
  XNOR U1142 ( .A(n1006), .B(n1007), .Z(n1008) );
  XNOR U1143 ( .A(n1009), .B(n1008), .Z(n117) );
  XNOR U1144 ( .A(n118), .B(n117), .Z(n119) );
  XNOR U1145 ( .A(n120), .B(n119), .Z(n518) );
  XNOR U1146 ( .A(n519), .B(n518), .Z(n868) );
  XNOR U1147 ( .A(n869), .B(n868), .Z(n870) );
  XNOR U1148 ( .A(n871), .B(n870), .Z(n717) );
  XNOR U1149 ( .A(n718), .B(n717), .Z(n719) );
  XOR U1150 ( .A(x[103]), .B(y[103]), .Z(n1141) );
  XOR U1151 ( .A(x[95]), .B(y[95]), .Z(n1138) );
  XNOR U1152 ( .A(x[99]), .B(y[99]), .Z(n1139) );
  XNOR U1153 ( .A(n1138), .B(n1139), .Z(n1140) );
  XOR U1154 ( .A(n1141), .B(n1140), .Z(n622) );
  XOR U1155 ( .A(x[115]), .B(y[115]), .Z(n319) );
  XOR U1156 ( .A(x[107]), .B(y[107]), .Z(n316) );
  XNOR U1157 ( .A(x[111]), .B(y[111]), .Z(n317) );
  XNOR U1158 ( .A(n316), .B(n317), .Z(n318) );
  XOR U1159 ( .A(n319), .B(n318), .Z(n620) );
  XOR U1160 ( .A(x[127]), .B(y[127]), .Z(n1189) );
  XOR U1161 ( .A(x[119]), .B(y[119]), .Z(n1186) );
  XNOR U1162 ( .A(x[123]), .B(y[123]), .Z(n1187) );
  XNOR U1163 ( .A(n1186), .B(n1187), .Z(n1188) );
  XNOR U1164 ( .A(n1189), .B(n1188), .Z(n619) );
  XNOR U1165 ( .A(n620), .B(n619), .Z(n621) );
  XNOR U1166 ( .A(n622), .B(n621), .Z(n765) );
  XOR U1167 ( .A(x[137]), .B(y[137]), .Z(n307) );
  XOR U1168 ( .A(x[131]), .B(y[131]), .Z(n304) );
  XNOR U1169 ( .A(x[135]), .B(y[135]), .Z(n305) );
  XNOR U1170 ( .A(n304), .B(n305), .Z(n306) );
  XOR U1171 ( .A(n307), .B(n306), .Z(n459) );
  XOR U1172 ( .A(x[143]), .B(y[143]), .Z(n895) );
  XOR U1173 ( .A(x[139]), .B(y[139]), .Z(n892) );
  XNOR U1174 ( .A(x[141]), .B(y[141]), .Z(n893) );
  XNOR U1175 ( .A(n892), .B(n893), .Z(n894) );
  XOR U1176 ( .A(n895), .B(n894), .Z(n457) );
  XOR U1177 ( .A(x[149]), .B(y[149]), .Z(n949) );
  XOR U1178 ( .A(x[145]), .B(y[145]), .Z(n946) );
  XNOR U1179 ( .A(x[147]), .B(y[147]), .Z(n947) );
  XNOR U1180 ( .A(n946), .B(n947), .Z(n948) );
  XNOR U1181 ( .A(n949), .B(n948), .Z(n456) );
  XNOR U1182 ( .A(n457), .B(n456), .Z(n458) );
  XOR U1183 ( .A(n459), .B(n458), .Z(n766) );
  XNOR U1184 ( .A(n765), .B(n766), .Z(n768) );
  XOR U1185 ( .A(x[155]), .B(y[155]), .Z(n1003) );
  XOR U1186 ( .A(x[151]), .B(y[151]), .Z(n1000) );
  XNOR U1187 ( .A(x[153]), .B(y[153]), .Z(n1001) );
  XNOR U1188 ( .A(n1000), .B(n1001), .Z(n1002) );
  XOR U1189 ( .A(n1003), .B(n1002), .Z(n525) );
  XOR U1190 ( .A(x[161]), .B(y[161]), .Z(n901) );
  XOR U1191 ( .A(x[157]), .B(y[157]), .Z(n898) );
  XNOR U1192 ( .A(x[159]), .B(y[159]), .Z(n899) );
  XNOR U1193 ( .A(n898), .B(n899), .Z(n900) );
  XOR U1194 ( .A(n901), .B(n900), .Z(n523) );
  XOR U1195 ( .A(x[167]), .B(y[167]), .Z(n288) );
  XOR U1196 ( .A(x[163]), .B(y[163]), .Z(n285) );
  XNOR U1197 ( .A(x[165]), .B(y[165]), .Z(n286) );
  XNOR U1198 ( .A(n285), .B(n286), .Z(n287) );
  XNOR U1199 ( .A(n288), .B(n287), .Z(n522) );
  XNOR U1200 ( .A(n523), .B(n522), .Z(n524) );
  XNOR U1201 ( .A(n525), .B(n524), .Z(n767) );
  XOR U1202 ( .A(n768), .B(n767), .Z(n865) );
  XOR U1203 ( .A(x[275]), .B(y[275]), .Z(n281) );
  XOR U1204 ( .A(x[289]), .B(y[289]), .Z(n279) );
  XNOR U1205 ( .A(x[301]), .B(y[301]), .Z(n280) );
  XOR U1206 ( .A(n279), .B(n280), .Z(n282) );
  XNOR U1207 ( .A(n281), .B(n282), .Z(n735) );
  XOR U1208 ( .A(x[273]), .B(y[273]), .Z(n966) );
  XOR U1209 ( .A(x[271]), .B(y[271]), .Z(n964) );
  XNOR U1210 ( .A(x[309]), .B(y[309]), .Z(n965) );
  XOR U1211 ( .A(n964), .B(n965), .Z(n967) );
  XOR U1212 ( .A(n966), .B(n967), .Z(n736) );
  XNOR U1213 ( .A(n735), .B(n736), .Z(n738) );
  XOR U1214 ( .A(x[283]), .B(y[283]), .Z(n267) );
  XNOR U1215 ( .A(x[285]), .B(y[285]), .Z(n268) );
  XNOR U1216 ( .A(n267), .B(n268), .Z(n269) );
  XOR U1217 ( .A(x[277]), .B(y[277]), .Z(n263) );
  XOR U1218 ( .A(x[279]), .B(y[279]), .Z(n261) );
  XNOR U1219 ( .A(x[293]), .B(y[293]), .Z(n262) );
  XOR U1220 ( .A(n261), .B(n262), .Z(n264) );
  XOR U1221 ( .A(n263), .B(n264), .Z(n270) );
  XNOR U1222 ( .A(n269), .B(n270), .Z(n737) );
  XOR U1223 ( .A(n738), .B(n737), .Z(n809) );
  XOR U1224 ( .A(x[209]), .B(y[209]), .Z(n1021) );
  XOR U1225 ( .A(x[205]), .B(y[205]), .Z(n1019) );
  XOR U1226 ( .A(x[207]), .B(y[207]), .Z(n1018) );
  XOR U1227 ( .A(n1019), .B(n1018), .Z(n1020) );
  XOR U1228 ( .A(n1021), .B(n1020), .Z(n646) );
  XOR U1229 ( .A(x[215]), .B(y[215]), .Z(n1027) );
  XOR U1230 ( .A(x[211]), .B(y[211]), .Z(n1025) );
  XOR U1231 ( .A(x[213]), .B(y[213]), .Z(n1024) );
  XOR U1232 ( .A(n1025), .B(n1024), .Z(n1026) );
  XOR U1233 ( .A(n1027), .B(n1026), .Z(n644) );
  XOR U1234 ( .A(x[221]), .B(y[221]), .Z(n1111) );
  XOR U1235 ( .A(x[217]), .B(y[217]), .Z(n1108) );
  XNOR U1236 ( .A(x[219]), .B(y[219]), .Z(n1109) );
  XNOR U1237 ( .A(n1108), .B(n1109), .Z(n1110) );
  XNOR U1238 ( .A(n1111), .B(n1110), .Z(n643) );
  XNOR U1239 ( .A(n644), .B(n643), .Z(n645) );
  XNOR U1240 ( .A(n646), .B(n645), .Z(n808) );
  XNOR U1241 ( .A(n809), .B(n808), .Z(n811) );
  XOR U1242 ( .A(x[225]), .B(y[225]), .Z(n1099) );
  XOR U1243 ( .A(x[223]), .B(y[223]), .Z(n1096) );
  XNOR U1244 ( .A(x[333]), .B(y[333]), .Z(n1097) );
  XNOR U1245 ( .A(n1096), .B(n1097), .Z(n1098) );
  XOR U1246 ( .A(n1099), .B(n1098), .Z(n579) );
  XOR U1247 ( .A(x[229]), .B(y[229]), .Z(n1105) );
  XOR U1248 ( .A(x[227]), .B(y[227]), .Z(n1102) );
  XNOR U1249 ( .A(x[331]), .B(y[331]), .Z(n1103) );
  XNOR U1250 ( .A(n1102), .B(n1103), .Z(n1104) );
  XOR U1251 ( .A(n1105), .B(n1104), .Z(n577) );
  XOR U1252 ( .A(x[233]), .B(y[233]), .Z(n943) );
  XOR U1253 ( .A(x[231]), .B(y[231]), .Z(n940) );
  XNOR U1254 ( .A(x[329]), .B(y[329]), .Z(n941) );
  XNOR U1255 ( .A(n940), .B(n941), .Z(n942) );
  XNOR U1256 ( .A(n943), .B(n942), .Z(n576) );
  XNOR U1257 ( .A(n577), .B(n576), .Z(n578) );
  XNOR U1258 ( .A(n579), .B(n578), .Z(n810) );
  XOR U1259 ( .A(n811), .B(n810), .Z(n863) );
  XOR U1260 ( .A(x[287]), .B(y[287]), .Z(n275) );
  XOR U1261 ( .A(x[281]), .B(y[281]), .Z(n273) );
  XNOR U1262 ( .A(x[291]), .B(y[291]), .Z(n274) );
  XOR U1263 ( .A(n273), .B(n274), .Z(n276) );
  XNOR U1264 ( .A(n275), .B(n276), .Z(n408) );
  XOR U1265 ( .A(x[295]), .B(y[295]), .Z(n257) );
  XOR U1266 ( .A(x[297]), .B(y[297]), .Z(n255) );
  XNOR U1267 ( .A(x[299]), .B(y[299]), .Z(n256) );
  XOR U1268 ( .A(n255), .B(n256), .Z(n258) );
  XOR U1269 ( .A(n257), .B(n258), .Z(n409) );
  XNOR U1270 ( .A(n408), .B(n409), .Z(n411) );
  XOR U1271 ( .A(x[303]), .B(y[303]), .Z(n972) );
  XOR U1272 ( .A(x[305]), .B(y[305]), .Z(n970) );
  XNOR U1273 ( .A(x[307]), .B(y[307]), .Z(n971) );
  XOR U1274 ( .A(n970), .B(n971), .Z(n973) );
  XNOR U1275 ( .A(n972), .B(n973), .Z(n410) );
  XOR U1276 ( .A(n411), .B(n410), .Z(n730) );
  XOR U1277 ( .A(x[173]), .B(y[173]), .Z(n300) );
  XOR U1278 ( .A(x[169]), .B(y[169]), .Z(n297) );
  XNOR U1279 ( .A(x[171]), .B(y[171]), .Z(n298) );
  XNOR U1280 ( .A(n297), .B(n298), .Z(n299) );
  XOR U1281 ( .A(n300), .B(n299), .Z(n549) );
  XOR U1282 ( .A(x[179]), .B(y[179]), .Z(n294) );
  XOR U1283 ( .A(x[175]), .B(y[175]), .Z(n291) );
  XNOR U1284 ( .A(x[177]), .B(y[177]), .Z(n292) );
  XNOR U1285 ( .A(n291), .B(n292), .Z(n293) );
  XOR U1286 ( .A(n294), .B(n293), .Z(n547) );
  XOR U1287 ( .A(x[185]), .B(y[185]), .Z(n925) );
  XOR U1288 ( .A(x[181]), .B(y[181]), .Z(n922) );
  XNOR U1289 ( .A(x[183]), .B(y[183]), .Z(n923) );
  XNOR U1290 ( .A(n922), .B(n923), .Z(n924) );
  XNOR U1291 ( .A(n925), .B(n924), .Z(n546) );
  XNOR U1292 ( .A(n547), .B(n546), .Z(n548) );
  XNOR U1293 ( .A(n549), .B(n548), .Z(n729) );
  XNOR U1294 ( .A(n730), .B(n729), .Z(n732) );
  XOR U1295 ( .A(x[191]), .B(y[191]), .Z(n913) );
  XOR U1296 ( .A(x[187]), .B(y[187]), .Z(n911) );
  XOR U1297 ( .A(x[189]), .B(y[189]), .Z(n910) );
  XOR U1298 ( .A(n911), .B(n910), .Z(n912) );
  XOR U1299 ( .A(n913), .B(n912), .Z(n483) );
  XOR U1300 ( .A(x[197]), .B(y[197]), .Z(n919) );
  XOR U1301 ( .A(x[193]), .B(y[193]), .Z(n917) );
  XOR U1302 ( .A(x[195]), .B(y[195]), .Z(n916) );
  XOR U1303 ( .A(n917), .B(n916), .Z(n918) );
  XOR U1304 ( .A(n919), .B(n918), .Z(n481) );
  XOR U1305 ( .A(x[203]), .B(y[203]), .Z(n1033) );
  XOR U1306 ( .A(x[199]), .B(y[199]), .Z(n1031) );
  XOR U1307 ( .A(x[201]), .B(y[201]), .Z(n1030) );
  XOR U1308 ( .A(n1031), .B(n1030), .Z(n1032) );
  XNOR U1309 ( .A(n1033), .B(n1032), .Z(n480) );
  XNOR U1310 ( .A(n481), .B(n480), .Z(n482) );
  XNOR U1311 ( .A(n483), .B(n482), .Z(n731) );
  XNOR U1312 ( .A(n732), .B(n731), .Z(n862) );
  XNOR U1313 ( .A(n863), .B(n862), .Z(n864) );
  XOR U1314 ( .A(n865), .B(n864), .Z(n720) );
  XNOR U1315 ( .A(n719), .B(n720), .Z(n725) );
  XOR U1316 ( .A(n726), .B(n725), .Z(o[0]) );
  NANDN U1317 ( .A(n82), .B(n81), .Z(n86) );
  NAND U1318 ( .A(n84), .B(n83), .Z(n85) );
  AND U1319 ( .A(n86), .B(n85), .Z(n1339) );
  NANDN U1320 ( .A(n88), .B(n87), .Z(n92) );
  NAND U1321 ( .A(n90), .B(n89), .Z(n91) );
  AND U1322 ( .A(n92), .B(n91), .Z(n1338) );
  NANDN U1323 ( .A(n94), .B(n93), .Z(n98) );
  NAND U1324 ( .A(n96), .B(n95), .Z(n97) );
  NAND U1325 ( .A(n98), .B(n97), .Z(n1337) );
  XOR U1326 ( .A(n1338), .B(n1337), .Z(n1340) );
  XOR U1327 ( .A(n1339), .B(n1340), .Z(n1749) );
  NANDN U1328 ( .A(n100), .B(n99), .Z(n104) );
  NANDN U1329 ( .A(n102), .B(n101), .Z(n103) );
  NAND U1330 ( .A(n104), .B(n103), .Z(n1748) );
  XNOR U1331 ( .A(n1749), .B(n1748), .Z(n1751) );
  NANDN U1332 ( .A(n106), .B(n105), .Z(n110) );
  NANDN U1333 ( .A(n108), .B(n107), .Z(n109) );
  AND U1334 ( .A(n110), .B(n109), .Z(n1725) );
  NANDN U1335 ( .A(n112), .B(n111), .Z(n116) );
  NANDN U1336 ( .A(n114), .B(n113), .Z(n115) );
  AND U1337 ( .A(n116), .B(n115), .Z(n1724) );
  XOR U1338 ( .A(n1725), .B(n1724), .Z(n1727) );
  NANDN U1339 ( .A(n118), .B(n117), .Z(n122) );
  NANDN U1340 ( .A(n120), .B(n119), .Z(n121) );
  AND U1341 ( .A(n122), .B(n121), .Z(n1726) );
  XOR U1342 ( .A(n1727), .B(n1726), .Z(n1537) );
  NANDN U1343 ( .A(n124), .B(n123), .Z(n128) );
  NANDN U1344 ( .A(n126), .B(n125), .Z(n127) );
  AND U1345 ( .A(n128), .B(n127), .Z(n1535) );
  NANDN U1346 ( .A(n130), .B(n129), .Z(n134) );
  NANDN U1347 ( .A(n132), .B(n131), .Z(n133) );
  NAND U1348 ( .A(n134), .B(n133), .Z(n1534) );
  XNOR U1349 ( .A(n1535), .B(n1534), .Z(n1536) );
  XNOR U1350 ( .A(n1537), .B(n1536), .Z(n1750) );
  XOR U1351 ( .A(n1751), .B(n1750), .Z(n1448) );
  NANDN U1352 ( .A(n136), .B(n135), .Z(n140) );
  NANDN U1353 ( .A(n138), .B(n137), .Z(n139) );
  AND U1354 ( .A(n140), .B(n139), .Z(n1732) );
  NANDN U1355 ( .A(n142), .B(n141), .Z(n146) );
  NANDN U1356 ( .A(n144), .B(n143), .Z(n145) );
  AND U1357 ( .A(n146), .B(n145), .Z(n1730) );
  NANDN U1358 ( .A(n148), .B(n147), .Z(n152) );
  NANDN U1359 ( .A(n150), .B(n149), .Z(n151) );
  NAND U1360 ( .A(n152), .B(n151), .Z(n1731) );
  XOR U1361 ( .A(n1730), .B(n1731), .Z(n1733) );
  XNOR U1362 ( .A(n1732), .B(n1733), .Z(n1857) );
  NANDN U1363 ( .A(n154), .B(n153), .Z(n158) );
  NAND U1364 ( .A(n156), .B(n155), .Z(n157) );
  AND U1365 ( .A(n158), .B(n157), .Z(n1316) );
  NANDN U1366 ( .A(n160), .B(n159), .Z(n164) );
  NAND U1367 ( .A(n162), .B(n161), .Z(n163) );
  AND U1368 ( .A(n164), .B(n163), .Z(n1314) );
  NANDN U1369 ( .A(n166), .B(n165), .Z(n170) );
  NANDN U1370 ( .A(n168), .B(n167), .Z(n169) );
  AND U1371 ( .A(n170), .B(n169), .Z(n1313) );
  XNOR U1372 ( .A(n1314), .B(n1313), .Z(n1315) );
  XOR U1373 ( .A(n1316), .B(n1315), .Z(n1858) );
  XNOR U1374 ( .A(n1857), .B(n1858), .Z(n1859) );
  NANDN U1375 ( .A(n172), .B(n171), .Z(n176) );
  NAND U1376 ( .A(n174), .B(n173), .Z(n175) );
  AND U1377 ( .A(n176), .B(n175), .Z(n1322) );
  NANDN U1378 ( .A(n178), .B(n177), .Z(n182) );
  NAND U1379 ( .A(n180), .B(n179), .Z(n181) );
  AND U1380 ( .A(n182), .B(n181), .Z(n1587) );
  NANDN U1381 ( .A(n184), .B(n183), .Z(n188) );
  NAND U1382 ( .A(n186), .B(n185), .Z(n187) );
  NAND U1383 ( .A(n188), .B(n187), .Z(n1588) );
  XNOR U1384 ( .A(n1587), .B(n1588), .Z(n1590) );
  NANDN U1385 ( .A(n190), .B(n189), .Z(n194) );
  NAND U1386 ( .A(n192), .B(n191), .Z(n193) );
  AND U1387 ( .A(n194), .B(n193), .Z(n1589) );
  XOR U1388 ( .A(n1590), .B(n1589), .Z(n1320) );
  NANDN U1389 ( .A(n196), .B(n195), .Z(n200) );
  NANDN U1390 ( .A(n198), .B(n197), .Z(n199) );
  AND U1391 ( .A(n200), .B(n199), .Z(n1319) );
  XNOR U1392 ( .A(n1320), .B(n1319), .Z(n1321) );
  XOR U1393 ( .A(n1322), .B(n1321), .Z(n1860) );
  XNOR U1394 ( .A(n1859), .B(n1860), .Z(n1446) );
  NANDN U1395 ( .A(n202), .B(n201), .Z(n206) );
  NANDN U1396 ( .A(n204), .B(n203), .Z(n205) );
  AND U1397 ( .A(n206), .B(n205), .Z(n1775) );
  NANDN U1398 ( .A(n208), .B(n207), .Z(n212) );
  NAND U1399 ( .A(n210), .B(n209), .Z(n211) );
  AND U1400 ( .A(n212), .B(n211), .Z(n1772) );
  NANDN U1401 ( .A(n214), .B(n213), .Z(n218) );
  NANDN U1402 ( .A(n216), .B(n215), .Z(n217) );
  AND U1403 ( .A(n218), .B(n217), .Z(n1333) );
  NANDN U1404 ( .A(n220), .B(n219), .Z(n224) );
  NAND U1405 ( .A(n222), .B(n221), .Z(n223) );
  AND U1406 ( .A(n224), .B(n223), .Z(n1332) );
  NANDN U1407 ( .A(n226), .B(n225), .Z(n230) );
  NANDN U1408 ( .A(n228), .B(n227), .Z(n229) );
  AND U1409 ( .A(n230), .B(n229), .Z(n1331) );
  XOR U1410 ( .A(n1332), .B(n1331), .Z(n1334) );
  XOR U1411 ( .A(n1333), .B(n1334), .Z(n1773) );
  XNOR U1412 ( .A(n1772), .B(n1773), .Z(n1774) );
  XNOR U1413 ( .A(n1775), .B(n1774), .Z(n1445) );
  XNOR U1414 ( .A(n1446), .B(n1445), .Z(n1447) );
  XOR U1415 ( .A(n1448), .B(n1447), .Z(n1791) );
  NANDN U1416 ( .A(n232), .B(n231), .Z(n236) );
  NAND U1417 ( .A(n234), .B(n233), .Z(n235) );
  NAND U1418 ( .A(n236), .B(n235), .Z(n1790) );
  XOR U1419 ( .A(n1791), .B(n1790), .Z(n1792) );
  NANDN U1420 ( .A(n238), .B(n237), .Z(n242) );
  NAND U1421 ( .A(n240), .B(n239), .Z(n241) );
  AND U1422 ( .A(n242), .B(n241), .Z(n1442) );
  NANDN U1423 ( .A(n244), .B(n243), .Z(n248) );
  NAND U1424 ( .A(n246), .B(n245), .Z(n247) );
  AND U1425 ( .A(n248), .B(n247), .Z(n1781) );
  NANDN U1426 ( .A(n250), .B(n249), .Z(n254) );
  NANDN U1427 ( .A(n252), .B(n251), .Z(n253) );
  AND U1428 ( .A(n254), .B(n253), .Z(n1504) );
  NANDN U1429 ( .A(n256), .B(n255), .Z(n260) );
  NANDN U1430 ( .A(n258), .B(n257), .Z(n259) );
  AND U1431 ( .A(n260), .B(n259), .Z(n1357) );
  NANDN U1432 ( .A(n262), .B(n261), .Z(n266) );
  NANDN U1433 ( .A(n264), .B(n263), .Z(n265) );
  AND U1434 ( .A(n266), .B(n265), .Z(n1355) );
  XNOR U1435 ( .A(n1355), .B(oglobal[1]), .Z(n1356) );
  XOR U1436 ( .A(n1357), .B(n1356), .Z(n1505) );
  XNOR U1437 ( .A(n1504), .B(n1505), .Z(n1506) );
  NANDN U1438 ( .A(n268), .B(n267), .Z(n272) );
  NANDN U1439 ( .A(n270), .B(n269), .Z(n271) );
  AND U1440 ( .A(n272), .B(n271), .Z(n1352) );
  NANDN U1441 ( .A(n274), .B(n273), .Z(n278) );
  NANDN U1442 ( .A(n276), .B(n275), .Z(n277) );
  AND U1443 ( .A(n278), .B(n277), .Z(n1350) );
  NANDN U1444 ( .A(n280), .B(n279), .Z(n284) );
  NANDN U1445 ( .A(n282), .B(n281), .Z(n283) );
  NAND U1446 ( .A(n284), .B(n283), .Z(n1349) );
  XNOR U1447 ( .A(n1350), .B(n1349), .Z(n1351) );
  XOR U1448 ( .A(n1352), .B(n1351), .Z(n1507) );
  XNOR U1449 ( .A(n1506), .B(n1507), .Z(n1779) );
  NANDN U1450 ( .A(n286), .B(n285), .Z(n290) );
  NAND U1451 ( .A(n288), .B(n287), .Z(n289) );
  NAND U1452 ( .A(n290), .B(n289), .Z(n1698) );
  NANDN U1453 ( .A(n292), .B(n291), .Z(n296) );
  NAND U1454 ( .A(n294), .B(n293), .Z(n295) );
  AND U1455 ( .A(n296), .B(n295), .Z(n1697) );
  NANDN U1456 ( .A(n298), .B(n297), .Z(n302) );
  NAND U1457 ( .A(n300), .B(n299), .Z(n301) );
  NAND U1458 ( .A(n302), .B(n301), .Z(n1696) );
  XOR U1459 ( .A(n1697), .B(n1696), .Z(n303) );
  XOR U1460 ( .A(n1698), .B(n303), .Z(n1494) );
  NANDN U1461 ( .A(n305), .B(n304), .Z(n309) );
  NAND U1462 ( .A(n307), .B(n306), .Z(n308) );
  NAND U1463 ( .A(n309), .B(n308), .Z(n1843) );
  NANDN U1464 ( .A(n311), .B(n310), .Z(n315) );
  NAND U1465 ( .A(n313), .B(n312), .Z(n314) );
  AND U1466 ( .A(n315), .B(n314), .Z(n1842) );
  NANDN U1467 ( .A(n317), .B(n316), .Z(n321) );
  NAND U1468 ( .A(n319), .B(n318), .Z(n320) );
  NAND U1469 ( .A(n321), .B(n320), .Z(n1841) );
  XOR U1470 ( .A(n1842), .B(n1841), .Z(n322) );
  XOR U1471 ( .A(n1843), .B(n322), .Z(n1493) );
  NANDN U1472 ( .A(n324), .B(n323), .Z(n328) );
  NANDN U1473 ( .A(n326), .B(n325), .Z(n327) );
  AND U1474 ( .A(n328), .B(n327), .Z(n1492) );
  XOR U1475 ( .A(n1493), .B(n1492), .Z(n1495) );
  XOR U1476 ( .A(n1494), .B(n1495), .Z(n1778) );
  XOR U1477 ( .A(n1779), .B(n1778), .Z(n1780) );
  XOR U1478 ( .A(n1781), .B(n1780), .Z(n1440) );
  NANDN U1479 ( .A(n330), .B(n329), .Z(n334) );
  NAND U1480 ( .A(n332), .B(n331), .Z(n333) );
  NAND U1481 ( .A(n334), .B(n333), .Z(n1548) );
  NANDN U1482 ( .A(n336), .B(n335), .Z(n340) );
  NAND U1483 ( .A(n338), .B(n337), .Z(n339) );
  NAND U1484 ( .A(n340), .B(n339), .Z(n1547) );
  NANDN U1485 ( .A(n342), .B(n341), .Z(n346) );
  NAND U1486 ( .A(n344), .B(n343), .Z(n345) );
  AND U1487 ( .A(n346), .B(n345), .Z(n1546) );
  XOR U1488 ( .A(n1547), .B(n1546), .Z(n347) );
  XOR U1489 ( .A(n1548), .B(n347), .Z(n1476) );
  NANDN U1490 ( .A(n349), .B(n348), .Z(n353) );
  NAND U1491 ( .A(n351), .B(n350), .Z(n352) );
  AND U1492 ( .A(n353), .B(n352), .Z(n1826) );
  NANDN U1493 ( .A(n355), .B(n354), .Z(n359) );
  NAND U1494 ( .A(n357), .B(n356), .Z(n358) );
  NAND U1495 ( .A(n359), .B(n358), .Z(n1827) );
  XNOR U1496 ( .A(n1826), .B(n1827), .Z(n1829) );
  NANDN U1497 ( .A(n361), .B(n360), .Z(n365) );
  NAND U1498 ( .A(n363), .B(n362), .Z(n364) );
  AND U1499 ( .A(n365), .B(n364), .Z(n1828) );
  XOR U1500 ( .A(n1829), .B(n1828), .Z(n1474) );
  NANDN U1501 ( .A(n367), .B(n366), .Z(n371) );
  NAND U1502 ( .A(n369), .B(n368), .Z(n370) );
  NAND U1503 ( .A(n371), .B(n370), .Z(n1473) );
  XNOR U1504 ( .A(n1474), .B(n1473), .Z(n1475) );
  XNOR U1505 ( .A(n1476), .B(n1475), .Z(n1851) );
  NANDN U1506 ( .A(n373), .B(n372), .Z(n377) );
  NANDN U1507 ( .A(n375), .B(n374), .Z(n376) );
  AND U1508 ( .A(n377), .B(n376), .Z(n1814) );
  NANDN U1509 ( .A(n379), .B(n378), .Z(n383) );
  NANDN U1510 ( .A(n381), .B(n380), .Z(n382) );
  NAND U1511 ( .A(n383), .B(n382), .Z(n1815) );
  XNOR U1512 ( .A(n1814), .B(n1815), .Z(n1817) );
  NANDN U1513 ( .A(n385), .B(n384), .Z(n389) );
  NANDN U1514 ( .A(n387), .B(n386), .Z(n388) );
  AND U1515 ( .A(n389), .B(n388), .Z(n1816) );
  XOR U1516 ( .A(n1817), .B(n1816), .Z(n1482) );
  NANDN U1517 ( .A(n391), .B(n390), .Z(n395) );
  NAND U1518 ( .A(n393), .B(n392), .Z(n394) );
  AND U1519 ( .A(n395), .B(n394), .Z(n1360) );
  NANDN U1520 ( .A(n397), .B(n396), .Z(n401) );
  NAND U1521 ( .A(n399), .B(n398), .Z(n400) );
  NAND U1522 ( .A(n401), .B(n400), .Z(n1361) );
  XNOR U1523 ( .A(n1360), .B(n1361), .Z(n1363) );
  NANDN U1524 ( .A(n403), .B(n402), .Z(n407) );
  NAND U1525 ( .A(n405), .B(n404), .Z(n406) );
  AND U1526 ( .A(n407), .B(n406), .Z(n1362) );
  XOR U1527 ( .A(n1363), .B(n1362), .Z(n1480) );
  NANDN U1528 ( .A(n409), .B(n408), .Z(n413) );
  NAND U1529 ( .A(n411), .B(n410), .Z(n412) );
  NAND U1530 ( .A(n413), .B(n412), .Z(n1479) );
  XNOR U1531 ( .A(n1480), .B(n1479), .Z(n1481) );
  XOR U1532 ( .A(n1482), .B(n1481), .Z(n1852) );
  XNOR U1533 ( .A(n1851), .B(n1852), .Z(n1854) );
  NANDN U1534 ( .A(n415), .B(n414), .Z(n419) );
  NAND U1535 ( .A(n417), .B(n416), .Z(n418) );
  AND U1536 ( .A(n419), .B(n418), .Z(n1575) );
  NANDN U1537 ( .A(n421), .B(n420), .Z(n425) );
  NAND U1538 ( .A(n423), .B(n422), .Z(n424) );
  NAND U1539 ( .A(n425), .B(n424), .Z(n1576) );
  XNOR U1540 ( .A(n1575), .B(n1576), .Z(n1578) );
  NANDN U1541 ( .A(n427), .B(n426), .Z(n431) );
  NAND U1542 ( .A(n429), .B(n428), .Z(n430) );
  AND U1543 ( .A(n431), .B(n430), .Z(n1577) );
  XOR U1544 ( .A(n1578), .B(n1577), .Z(n1458) );
  NANDN U1545 ( .A(n433), .B(n432), .Z(n437) );
  NAND U1546 ( .A(n435), .B(n434), .Z(n436) );
  AND U1547 ( .A(n437), .B(n436), .Z(n1820) );
  NANDN U1548 ( .A(n439), .B(n438), .Z(n443) );
  NAND U1549 ( .A(n441), .B(n440), .Z(n442) );
  NAND U1550 ( .A(n443), .B(n442), .Z(n1821) );
  XNOR U1551 ( .A(n1820), .B(n1821), .Z(n1823) );
  NANDN U1552 ( .A(n445), .B(n444), .Z(n449) );
  NAND U1553 ( .A(n447), .B(n446), .Z(n448) );
  AND U1554 ( .A(n449), .B(n448), .Z(n1822) );
  XOR U1555 ( .A(n1823), .B(n1822), .Z(n1456) );
  NANDN U1556 ( .A(n451), .B(n450), .Z(n455) );
  OR U1557 ( .A(n453), .B(n452), .Z(n454) );
  AND U1558 ( .A(n455), .B(n454), .Z(n1455) );
  XNOR U1559 ( .A(n1456), .B(n1455), .Z(n1457) );
  XNOR U1560 ( .A(n1458), .B(n1457), .Z(n1853) );
  XNOR U1561 ( .A(n1854), .B(n1853), .Z(n1439) );
  XNOR U1562 ( .A(n1440), .B(n1439), .Z(n1441) );
  XOR U1563 ( .A(n1442), .B(n1441), .Z(n1793) );
  XNOR U1564 ( .A(n1792), .B(n1793), .Z(n1787) );
  NANDN U1565 ( .A(n457), .B(n456), .Z(n461) );
  NANDN U1566 ( .A(n459), .B(n458), .Z(n460) );
  AND U1567 ( .A(n461), .B(n460), .Z(n1553) );
  NANDN U1568 ( .A(n463), .B(n462), .Z(n467) );
  NAND U1569 ( .A(n465), .B(n464), .Z(n466) );
  AND U1570 ( .A(n467), .B(n466), .Z(n1612) );
  NANDN U1571 ( .A(n469), .B(n468), .Z(n473) );
  NANDN U1572 ( .A(n471), .B(n470), .Z(n472) );
  NAND U1573 ( .A(n473), .B(n472), .Z(n1613) );
  XNOR U1574 ( .A(n1612), .B(n1613), .Z(n1615) );
  NANDN U1575 ( .A(n475), .B(n474), .Z(n479) );
  NANDN U1576 ( .A(n477), .B(n476), .Z(n478) );
  AND U1577 ( .A(n479), .B(n478), .Z(n1614) );
  XOR U1578 ( .A(n1615), .B(n1614), .Z(n1551) );
  NANDN U1579 ( .A(n481), .B(n480), .Z(n485) );
  NANDN U1580 ( .A(n483), .B(n482), .Z(n484) );
  AND U1581 ( .A(n485), .B(n484), .Z(n1550) );
  XNOR U1582 ( .A(n1551), .B(n1550), .Z(n1552) );
  XOR U1583 ( .A(n1553), .B(n1552), .Z(n1745) );
  NANDN U1584 ( .A(n487), .B(n486), .Z(n491) );
  NANDN U1585 ( .A(n489), .B(n488), .Z(n490) );
  AND U1586 ( .A(n491), .B(n490), .Z(n1684) );
  NANDN U1587 ( .A(n493), .B(n492), .Z(n497) );
  NANDN U1588 ( .A(n495), .B(n494), .Z(n496) );
  AND U1589 ( .A(n497), .B(n496), .Z(n1674) );
  NANDN U1590 ( .A(n499), .B(n498), .Z(n503) );
  NAND U1591 ( .A(n501), .B(n500), .Z(n502) );
  NAND U1592 ( .A(n503), .B(n502), .Z(n1675) );
  XNOR U1593 ( .A(n1674), .B(n1675), .Z(n1677) );
  NANDN U1594 ( .A(n505), .B(n504), .Z(n509) );
  NAND U1595 ( .A(n507), .B(n506), .Z(n508) );
  AND U1596 ( .A(n509), .B(n508), .Z(n1676) );
  XOR U1597 ( .A(n1677), .B(n1676), .Z(n1682) );
  NANDN U1598 ( .A(n511), .B(n510), .Z(n515) );
  NANDN U1599 ( .A(n513), .B(n512), .Z(n514) );
  AND U1600 ( .A(n515), .B(n514), .Z(n1681) );
  XNOR U1601 ( .A(n1682), .B(n1681), .Z(n1683) );
  XOR U1602 ( .A(n1684), .B(n1683), .Z(n1743) );
  NANDN U1603 ( .A(n517), .B(n516), .Z(n521) );
  NAND U1604 ( .A(n519), .B(n518), .Z(n520) );
  NAND U1605 ( .A(n521), .B(n520), .Z(n1742) );
  XNOR U1606 ( .A(n1743), .B(n1742), .Z(n1744) );
  XOR U1607 ( .A(n1745), .B(n1744), .Z(n1302) );
  NANDN U1608 ( .A(n523), .B(n522), .Z(n527) );
  NANDN U1609 ( .A(n525), .B(n524), .Z(n526) );
  AND U1610 ( .A(n527), .B(n526), .Z(n1370) );
  NANDN U1611 ( .A(n529), .B(n528), .Z(n533) );
  NAND U1612 ( .A(n531), .B(n530), .Z(n532) );
  AND U1613 ( .A(n533), .B(n532), .Z(n1373) );
  NANDN U1614 ( .A(n535), .B(n534), .Z(n539) );
  NANDN U1615 ( .A(n537), .B(n536), .Z(n538) );
  NAND U1616 ( .A(n539), .B(n538), .Z(n1374) );
  XNOR U1617 ( .A(n1373), .B(n1374), .Z(n1376) );
  NANDN U1618 ( .A(n541), .B(n540), .Z(n545) );
  NAND U1619 ( .A(n543), .B(n542), .Z(n544) );
  AND U1620 ( .A(n545), .B(n544), .Z(n1375) );
  XOR U1621 ( .A(n1376), .B(n1375), .Z(n1368) );
  NANDN U1622 ( .A(n547), .B(n546), .Z(n551) );
  NANDN U1623 ( .A(n549), .B(n548), .Z(n550) );
  AND U1624 ( .A(n551), .B(n550), .Z(n1367) );
  XNOR U1625 ( .A(n1368), .B(n1367), .Z(n1369) );
  XOR U1626 ( .A(n1370), .B(n1369), .Z(n1805) );
  NANDN U1627 ( .A(n553), .B(n552), .Z(n557) );
  NAND U1628 ( .A(n555), .B(n554), .Z(n556) );
  AND U1629 ( .A(n557), .B(n556), .Z(n1627) );
  NANDN U1630 ( .A(n559), .B(n558), .Z(n563) );
  NANDN U1631 ( .A(n561), .B(n560), .Z(n562) );
  AND U1632 ( .A(n563), .B(n562), .Z(n1668) );
  NANDN U1633 ( .A(n565), .B(n564), .Z(n569) );
  NAND U1634 ( .A(n567), .B(n566), .Z(n568) );
  NAND U1635 ( .A(n569), .B(n568), .Z(n1669) );
  XNOR U1636 ( .A(n1668), .B(n1669), .Z(n1671) );
  NANDN U1637 ( .A(n571), .B(n570), .Z(n575) );
  NANDN U1638 ( .A(n573), .B(n572), .Z(n574) );
  AND U1639 ( .A(n575), .B(n574), .Z(n1670) );
  XOR U1640 ( .A(n1671), .B(n1670), .Z(n1626) );
  NANDN U1641 ( .A(n577), .B(n576), .Z(n581) );
  NANDN U1642 ( .A(n579), .B(n578), .Z(n580) );
  AND U1643 ( .A(n581), .B(n580), .Z(n1625) );
  XOR U1644 ( .A(n1626), .B(n1625), .Z(n1628) );
  XOR U1645 ( .A(n1627), .B(n1628), .Z(n1803) );
  NANDN U1646 ( .A(n583), .B(n582), .Z(n587) );
  NANDN U1647 ( .A(n585), .B(n584), .Z(n586) );
  AND U1648 ( .A(n587), .B(n586), .Z(n1802) );
  XNOR U1649 ( .A(n1803), .B(n1802), .Z(n1804) );
  XOR U1650 ( .A(n1805), .B(n1804), .Z(n1301) );
  XOR U1651 ( .A(n1302), .B(n1301), .Z(n1304) );
  NANDN U1652 ( .A(n589), .B(n588), .Z(n593) );
  NANDN U1653 ( .A(n591), .B(n590), .Z(n592) );
  AND U1654 ( .A(n593), .B(n592), .Z(n1847) );
  NANDN U1655 ( .A(n595), .B(n594), .Z(n599) );
  NAND U1656 ( .A(n597), .B(n596), .Z(n598) );
  AND U1657 ( .A(n599), .B(n598), .Z(n1846) );
  NANDN U1658 ( .A(n601), .B(n600), .Z(n605) );
  NAND U1659 ( .A(n603), .B(n602), .Z(n604) );
  NAND U1660 ( .A(n605), .B(n604), .Z(n1610) );
  NANDN U1661 ( .A(n607), .B(n606), .Z(n611) );
  NAND U1662 ( .A(n609), .B(n608), .Z(n610) );
  AND U1663 ( .A(n611), .B(n610), .Z(n1609) );
  NANDN U1664 ( .A(n613), .B(n612), .Z(n617) );
  NAND U1665 ( .A(n615), .B(n614), .Z(n616) );
  NAND U1666 ( .A(n617), .B(n616), .Z(n1608) );
  XOR U1667 ( .A(n1609), .B(n1608), .Z(n618) );
  XNOR U1668 ( .A(n1610), .B(n618), .Z(n1845) );
  XOR U1669 ( .A(n1846), .B(n1845), .Z(n1848) );
  XOR U1670 ( .A(n1847), .B(n1848), .Z(n1756) );
  NANDN U1671 ( .A(n620), .B(n619), .Z(n624) );
  NANDN U1672 ( .A(n622), .B(n621), .Z(n623) );
  AND U1673 ( .A(n624), .B(n623), .Z(n1417) );
  NANDN U1674 ( .A(n626), .B(n625), .Z(n630) );
  NANDN U1675 ( .A(n628), .B(n627), .Z(n629) );
  AND U1676 ( .A(n630), .B(n629), .Z(n1599) );
  NANDN U1677 ( .A(n632), .B(n631), .Z(n636) );
  NANDN U1678 ( .A(n634), .B(n633), .Z(n635) );
  NAND U1679 ( .A(n636), .B(n635), .Z(n1600) );
  XNOR U1680 ( .A(n1599), .B(n1600), .Z(n1602) );
  NANDN U1681 ( .A(n638), .B(n637), .Z(n642) );
  NANDN U1682 ( .A(n640), .B(n639), .Z(n641) );
  AND U1683 ( .A(n642), .B(n641), .Z(n1601) );
  XOR U1684 ( .A(n1602), .B(n1601), .Z(n1416) );
  NANDN U1685 ( .A(n644), .B(n643), .Z(n648) );
  NANDN U1686 ( .A(n646), .B(n645), .Z(n647) );
  AND U1687 ( .A(n648), .B(n647), .Z(n1415) );
  XOR U1688 ( .A(n1416), .B(n1415), .Z(n1418) );
  XOR U1689 ( .A(n1417), .B(n1418), .Z(n1755) );
  NANDN U1690 ( .A(n650), .B(n649), .Z(n654) );
  NAND U1691 ( .A(n652), .B(n651), .Z(n653) );
  NAND U1692 ( .A(n654), .B(n653), .Z(n1840) );
  NANDN U1693 ( .A(n656), .B(n655), .Z(n660) );
  NAND U1694 ( .A(n658), .B(n657), .Z(n659) );
  AND U1695 ( .A(n660), .B(n659), .Z(n1839) );
  NANDN U1696 ( .A(n662), .B(n661), .Z(n666) );
  NANDN U1697 ( .A(n664), .B(n663), .Z(n665) );
  NAND U1698 ( .A(n666), .B(n665), .Z(n1838) );
  XOR U1699 ( .A(n1839), .B(n1838), .Z(n667) );
  XOR U1700 ( .A(n1840), .B(n667), .Z(n1310) );
  NANDN U1701 ( .A(n669), .B(n668), .Z(n673) );
  NANDN U1702 ( .A(n671), .B(n670), .Z(n672) );
  AND U1703 ( .A(n673), .B(n672), .Z(n1706) );
  NAND U1704 ( .A(n675), .B(n674), .Z(n679) );
  NAND U1705 ( .A(n677), .B(n676), .Z(n678) );
  NAND U1706 ( .A(n679), .B(n678), .Z(n1707) );
  XNOR U1707 ( .A(n1706), .B(n1707), .Z(n1709) );
  NAND U1708 ( .A(n681), .B(n680), .Z(n685) );
  NAND U1709 ( .A(n683), .B(n682), .Z(n684) );
  AND U1710 ( .A(n685), .B(n684), .Z(n1708) );
  XOR U1711 ( .A(n1709), .B(n1708), .Z(n1308) );
  NANDN U1712 ( .A(n687), .B(n686), .Z(n691) );
  NAND U1713 ( .A(n689), .B(n688), .Z(n690) );
  NAND U1714 ( .A(n691), .B(n690), .Z(n1623) );
  NANDN U1715 ( .A(n693), .B(n692), .Z(n697) );
  NANDN U1716 ( .A(n695), .B(n694), .Z(n696) );
  NAND U1717 ( .A(n697), .B(n696), .Z(n1622) );
  NANDN U1718 ( .A(n699), .B(n698), .Z(n703) );
  NANDN U1719 ( .A(n701), .B(n700), .Z(n702) );
  AND U1720 ( .A(n703), .B(n702), .Z(n1621) );
  XOR U1721 ( .A(n1622), .B(n1621), .Z(n704) );
  XNOR U1722 ( .A(n1623), .B(n704), .Z(n1307) );
  XNOR U1723 ( .A(n1308), .B(n1307), .Z(n1309) );
  XOR U1724 ( .A(n1310), .B(n1309), .Z(n1754) );
  XOR U1725 ( .A(n1755), .B(n1754), .Z(n1757) );
  NANDN U1726 ( .A(n706), .B(n705), .Z(n710) );
  NANDN U1727 ( .A(n708), .B(n707), .Z(n709) );
  AND U1728 ( .A(n710), .B(n709), .Z(n1528) );
  NANDN U1729 ( .A(n712), .B(n711), .Z(n716) );
  NANDN U1730 ( .A(n714), .B(n713), .Z(n715) );
  NAND U1731 ( .A(n716), .B(n715), .Z(n1529) );
  XNOR U1732 ( .A(n1528), .B(n1529), .Z(n1531) );
  XOR U1733 ( .A(n1530), .B(n1531), .Z(n1303) );
  XOR U1734 ( .A(n1304), .B(n1303), .Z(n1785) );
  NANDN U1735 ( .A(n718), .B(n717), .Z(n722) );
  NANDN U1736 ( .A(n720), .B(n719), .Z(n721) );
  AND U1737 ( .A(n722), .B(n721), .Z(n1784) );
  XNOR U1738 ( .A(n1785), .B(n1784), .Z(n1786) );
  XOR U1739 ( .A(n1787), .B(n1786), .Z(n1290) );
  NANDN U1740 ( .A(n724), .B(n723), .Z(n728) );
  NAND U1741 ( .A(n726), .B(n725), .Z(n727) );
  NAND U1742 ( .A(n728), .B(n727), .Z(n1289) );
  XNOR U1743 ( .A(n1290), .B(n1289), .Z(n1292) );
  NANDN U1744 ( .A(n730), .B(n729), .Z(n734) );
  NAND U1745 ( .A(n732), .B(n731), .Z(n733) );
  AND U1746 ( .A(n734), .B(n733), .Z(n1394) );
  NANDN U1747 ( .A(n736), .B(n735), .Z(n740) );
  NAND U1748 ( .A(n738), .B(n737), .Z(n739) );
  AND U1749 ( .A(n740), .B(n739), .Z(n1345) );
  NANDN U1750 ( .A(n742), .B(n741), .Z(n746) );
  NAND U1751 ( .A(n744), .B(n743), .Z(n745) );
  AND U1752 ( .A(n746), .B(n745), .Z(n1344) );
  NANDN U1753 ( .A(n748), .B(n747), .Z(n752) );
  NANDN U1754 ( .A(n750), .B(n749), .Z(n751) );
  AND U1755 ( .A(n752), .B(n751), .Z(n1662) );
  NANDN U1756 ( .A(n754), .B(n753), .Z(n758) );
  NAND U1757 ( .A(n756), .B(n755), .Z(n757) );
  NAND U1758 ( .A(n758), .B(n757), .Z(n1663) );
  XNOR U1759 ( .A(n1662), .B(n1663), .Z(n1665) );
  NANDN U1760 ( .A(n760), .B(n759), .Z(n764) );
  NAND U1761 ( .A(n762), .B(n761), .Z(n763) );
  AND U1762 ( .A(n764), .B(n763), .Z(n1664) );
  XNOR U1763 ( .A(n1665), .B(n1664), .Z(n1343) );
  XOR U1764 ( .A(n1344), .B(n1343), .Z(n1346) );
  XOR U1765 ( .A(n1345), .B(n1346), .Z(n1392) );
  NANDN U1766 ( .A(n766), .B(n765), .Z(n770) );
  NAND U1767 ( .A(n768), .B(n767), .Z(n769) );
  NAND U1768 ( .A(n770), .B(n769), .Z(n1391) );
  XNOR U1769 ( .A(n1392), .B(n1391), .Z(n1393) );
  XOR U1770 ( .A(n1394), .B(n1393), .Z(n1798) );
  NANDN U1771 ( .A(n772), .B(n771), .Z(n776) );
  NANDN U1772 ( .A(n774), .B(n773), .Z(n775) );
  AND U1773 ( .A(n776), .B(n775), .Z(n1328) );
  NANDN U1774 ( .A(n778), .B(n777), .Z(n782) );
  NANDN U1775 ( .A(n780), .B(n779), .Z(n781) );
  AND U1776 ( .A(n782), .B(n781), .Z(n1739) );
  NANDN U1777 ( .A(n784), .B(n783), .Z(n788) );
  NAND U1778 ( .A(n786), .B(n785), .Z(n787) );
  AND U1779 ( .A(n788), .B(n787), .Z(n1737) );
  NANDN U1780 ( .A(n790), .B(n789), .Z(n794) );
  NAND U1781 ( .A(n792), .B(n791), .Z(n793) );
  NAND U1782 ( .A(n794), .B(n793), .Z(n1695) );
  NANDN U1783 ( .A(n796), .B(n795), .Z(n800) );
  NANDN U1784 ( .A(n798), .B(n797), .Z(n799) );
  NAND U1785 ( .A(n800), .B(n799), .Z(n1694) );
  NANDN U1786 ( .A(n802), .B(n801), .Z(n806) );
  NAND U1787 ( .A(n804), .B(n803), .Z(n805) );
  AND U1788 ( .A(n806), .B(n805), .Z(n1693) );
  XOR U1789 ( .A(n1694), .B(n1693), .Z(n807) );
  XNOR U1790 ( .A(n1695), .B(n807), .Z(n1736) );
  XNOR U1791 ( .A(n1737), .B(n1736), .Z(n1738) );
  XOR U1792 ( .A(n1739), .B(n1738), .Z(n1326) );
  NANDN U1793 ( .A(n809), .B(n808), .Z(n813) );
  NAND U1794 ( .A(n811), .B(n810), .Z(n812) );
  NAND U1795 ( .A(n813), .B(n812), .Z(n1325) );
  XNOR U1796 ( .A(n1326), .B(n1325), .Z(n1327) );
  XOR U1797 ( .A(n1328), .B(n1327), .Z(n1796) );
  NANDN U1798 ( .A(n815), .B(n814), .Z(n819) );
  NANDN U1799 ( .A(n817), .B(n816), .Z(n818) );
  AND U1800 ( .A(n819), .B(n818), .Z(n1769) );
  NANDN U1801 ( .A(n821), .B(n820), .Z(n825) );
  NANDN U1802 ( .A(n823), .B(n822), .Z(n824) );
  AND U1803 ( .A(n825), .B(n824), .Z(n1766) );
  NANDN U1804 ( .A(n827), .B(n826), .Z(n831) );
  NANDN U1805 ( .A(n829), .B(n828), .Z(n830) );
  AND U1806 ( .A(n831), .B(n830), .Z(n1702) );
  NANDN U1807 ( .A(n833), .B(n832), .Z(n837) );
  NANDN U1808 ( .A(n835), .B(n834), .Z(n836) );
  AND U1809 ( .A(n837), .B(n836), .Z(n1649) );
  NANDN U1810 ( .A(n839), .B(n838), .Z(n843) );
  NAND U1811 ( .A(n841), .B(n840), .Z(n842) );
  NAND U1812 ( .A(n843), .B(n842), .Z(n1650) );
  XNOR U1813 ( .A(n1649), .B(n1650), .Z(n1652) );
  NANDN U1814 ( .A(n845), .B(n844), .Z(n849) );
  NAND U1815 ( .A(n847), .B(n846), .Z(n848) );
  AND U1816 ( .A(n849), .B(n848), .Z(n1651) );
  XOR U1817 ( .A(n1652), .B(n1651), .Z(n1701) );
  NANDN U1818 ( .A(n851), .B(n850), .Z(n855) );
  NANDN U1819 ( .A(n853), .B(n852), .Z(n854) );
  AND U1820 ( .A(n855), .B(n854), .Z(n1700) );
  XOR U1821 ( .A(n1701), .B(n1700), .Z(n1703) );
  XOR U1822 ( .A(n1702), .B(n1703), .Z(n1767) );
  XNOR U1823 ( .A(n1766), .B(n1767), .Z(n1768) );
  XOR U1824 ( .A(n1769), .B(n1768), .Z(n1797) );
  XOR U1825 ( .A(n1796), .B(n1797), .Z(n1799) );
  XNOR U1826 ( .A(n1798), .B(n1799), .Z(n1297) );
  NAND U1827 ( .A(n857), .B(n856), .Z(n861) );
  NAND U1828 ( .A(n859), .B(n858), .Z(n860) );
  NAND U1829 ( .A(n861), .B(n860), .Z(n1631) );
  NANDN U1830 ( .A(n863), .B(n862), .Z(n867) );
  NANDN U1831 ( .A(n865), .B(n864), .Z(n866) );
  AND U1832 ( .A(n867), .B(n866), .Z(n1632) );
  XOR U1833 ( .A(n1631), .B(n1632), .Z(n1634) );
  NANDN U1834 ( .A(n869), .B(n868), .Z(n873) );
  NANDN U1835 ( .A(n871), .B(n870), .Z(n872) );
  AND U1836 ( .A(n873), .B(n872), .Z(n1633) );
  XOR U1837 ( .A(n1634), .B(n1633), .Z(n1295) );
  NANDN U1838 ( .A(n875), .B(n874), .Z(n879) );
  NANDN U1839 ( .A(n877), .B(n876), .Z(n878) );
  AND U1840 ( .A(n879), .B(n878), .Z(n1397) );
  NANDN U1841 ( .A(n881), .B(n880), .Z(n885) );
  NANDN U1842 ( .A(n883), .B(n882), .Z(n884) );
  NAND U1843 ( .A(n885), .B(n884), .Z(n1398) );
  XNOR U1844 ( .A(n1397), .B(n1398), .Z(n1400) );
  NANDN U1845 ( .A(n887), .B(n886), .Z(n891) );
  NANDN U1846 ( .A(n889), .B(n888), .Z(n890) );
  AND U1847 ( .A(n891), .B(n890), .Z(n1399) );
  XOR U1848 ( .A(n1400), .B(n1399), .Z(n1488) );
  NANDN U1849 ( .A(n893), .B(n892), .Z(n897) );
  NAND U1850 ( .A(n895), .B(n894), .Z(n896) );
  AND U1851 ( .A(n897), .B(n896), .Z(n1643) );
  NANDN U1852 ( .A(n899), .B(n898), .Z(n903) );
  NAND U1853 ( .A(n901), .B(n900), .Z(n902) );
  NAND U1854 ( .A(n903), .B(n902), .Z(n1644) );
  XNOR U1855 ( .A(n1643), .B(n1644), .Z(n1646) );
  NANDN U1856 ( .A(n905), .B(n904), .Z(n909) );
  NAND U1857 ( .A(n907), .B(n906), .Z(n908) );
  AND U1858 ( .A(n909), .B(n908), .Z(n1645) );
  XOR U1859 ( .A(n1646), .B(n1645), .Z(n1486) );
  NAND U1860 ( .A(n911), .B(n910), .Z(n915) );
  NAND U1861 ( .A(n913), .B(n912), .Z(n914) );
  AND U1862 ( .A(n915), .B(n914), .Z(n1718) );
  NAND U1863 ( .A(n917), .B(n916), .Z(n921) );
  NAND U1864 ( .A(n919), .B(n918), .Z(n920) );
  NAND U1865 ( .A(n921), .B(n920), .Z(n1719) );
  XNOR U1866 ( .A(n1718), .B(n1719), .Z(n1721) );
  NANDN U1867 ( .A(n923), .B(n922), .Z(n927) );
  NAND U1868 ( .A(n925), .B(n924), .Z(n926) );
  AND U1869 ( .A(n927), .B(n926), .Z(n1720) );
  XNOR U1870 ( .A(n1721), .B(n1720), .Z(n1485) );
  XNOR U1871 ( .A(n1486), .B(n1485), .Z(n1487) );
  XNOR U1872 ( .A(n1488), .B(n1487), .Z(n1760) );
  NANDN U1873 ( .A(n929), .B(n928), .Z(n933) );
  NANDN U1874 ( .A(n931), .B(n930), .Z(n932) );
  AND U1875 ( .A(n933), .B(n932), .Z(n1427) );
  NANDN U1876 ( .A(n935), .B(n934), .Z(n939) );
  NANDN U1877 ( .A(n937), .B(n936), .Z(n938) );
  NAND U1878 ( .A(n939), .B(n938), .Z(n1428) );
  XNOR U1879 ( .A(n1427), .B(n1428), .Z(n1430) );
  NANDN U1880 ( .A(n941), .B(n940), .Z(n945) );
  NAND U1881 ( .A(n943), .B(n942), .Z(n944) );
  AND U1882 ( .A(n945), .B(n944), .Z(n1429) );
  XOR U1883 ( .A(n1430), .B(n1429), .Z(n1464) );
  NANDN U1884 ( .A(n947), .B(n946), .Z(n951) );
  NAND U1885 ( .A(n949), .B(n948), .Z(n950) );
  AND U1886 ( .A(n951), .B(n950), .Z(n1655) );
  NANDN U1887 ( .A(n953), .B(n952), .Z(n957) );
  NAND U1888 ( .A(n955), .B(n954), .Z(n956) );
  NAND U1889 ( .A(n957), .B(n956), .Z(n1656) );
  XNOR U1890 ( .A(n1655), .B(n1656), .Z(n1658) );
  NANDN U1891 ( .A(n959), .B(n958), .Z(n963) );
  NAND U1892 ( .A(n961), .B(n960), .Z(n962) );
  AND U1893 ( .A(n963), .B(n962), .Z(n1657) );
  XOR U1894 ( .A(n1658), .B(n1657), .Z(n1462) );
  NANDN U1895 ( .A(n965), .B(n964), .Z(n969) );
  NANDN U1896 ( .A(n967), .B(n966), .Z(n968) );
  AND U1897 ( .A(n969), .B(n968), .Z(n1385) );
  NANDN U1898 ( .A(n971), .B(n970), .Z(n975) );
  NANDN U1899 ( .A(n973), .B(n972), .Z(n974) );
  NAND U1900 ( .A(n975), .B(n974), .Z(n1386) );
  XNOR U1901 ( .A(n1385), .B(n1386), .Z(n1388) );
  NANDN U1902 ( .A(n977), .B(n976), .Z(n981) );
  NANDN U1903 ( .A(n979), .B(n978), .Z(n980) );
  AND U1904 ( .A(n981), .B(n980), .Z(n1387) );
  XNOR U1905 ( .A(n1388), .B(n1387), .Z(n1461) );
  XNOR U1906 ( .A(n1462), .B(n1461), .Z(n1463) );
  XOR U1907 ( .A(n1464), .B(n1463), .Z(n1761) );
  XNOR U1908 ( .A(n1760), .B(n1761), .Z(n1762) );
  NANDN U1909 ( .A(n983), .B(n982), .Z(n987) );
  NANDN U1910 ( .A(n985), .B(n984), .Z(n986) );
  AND U1911 ( .A(n987), .B(n986), .Z(n1403) );
  NANDN U1912 ( .A(n989), .B(n988), .Z(n993) );
  NANDN U1913 ( .A(n991), .B(n990), .Z(n992) );
  NAND U1914 ( .A(n993), .B(n992), .Z(n1404) );
  XNOR U1915 ( .A(n1403), .B(n1404), .Z(n1406) );
  NANDN U1916 ( .A(n995), .B(n994), .Z(n999) );
  NANDN U1917 ( .A(n997), .B(n996), .Z(n998) );
  AND U1918 ( .A(n999), .B(n998), .Z(n1405) );
  XOR U1919 ( .A(n1406), .B(n1405), .Z(n1452) );
  NANDN U1920 ( .A(n1001), .B(n1000), .Z(n1005) );
  NAND U1921 ( .A(n1003), .B(n1002), .Z(n1004) );
  AND U1922 ( .A(n1005), .B(n1004), .Z(n1687) );
  NANDN U1923 ( .A(n1007), .B(n1006), .Z(n1011) );
  NAND U1924 ( .A(n1009), .B(n1008), .Z(n1010) );
  NAND U1925 ( .A(n1011), .B(n1010), .Z(n1688) );
  XNOR U1926 ( .A(n1687), .B(n1688), .Z(n1690) );
  NANDN U1927 ( .A(n1013), .B(n1012), .Z(n1017) );
  NAND U1928 ( .A(n1015), .B(n1014), .Z(n1016) );
  AND U1929 ( .A(n1017), .B(n1016), .Z(n1689) );
  XOR U1930 ( .A(n1690), .B(n1689), .Z(n1450) );
  NAND U1931 ( .A(n1019), .B(n1018), .Z(n1023) );
  NAND U1932 ( .A(n1021), .B(n1020), .Z(n1022) );
  AND U1933 ( .A(n1023), .B(n1022), .Z(n1712) );
  NAND U1934 ( .A(n1025), .B(n1024), .Z(n1029) );
  NAND U1935 ( .A(n1027), .B(n1026), .Z(n1028) );
  NAND U1936 ( .A(n1029), .B(n1028), .Z(n1713) );
  XNOR U1937 ( .A(n1712), .B(n1713), .Z(n1715) );
  NAND U1938 ( .A(n1031), .B(n1030), .Z(n1035) );
  NAND U1939 ( .A(n1033), .B(n1032), .Z(n1034) );
  AND U1940 ( .A(n1035), .B(n1034), .Z(n1714) );
  XNOR U1941 ( .A(n1715), .B(n1714), .Z(n1449) );
  XNOR U1942 ( .A(n1450), .B(n1449), .Z(n1451) );
  XOR U1943 ( .A(n1452), .B(n1451), .Z(n1763) );
  XOR U1944 ( .A(n1762), .B(n1763), .Z(n1638) );
  NANDN U1945 ( .A(n1037), .B(n1036), .Z(n1041) );
  NANDN U1946 ( .A(n1039), .B(n1038), .Z(n1040) );
  AND U1947 ( .A(n1041), .B(n1040), .Z(n1811) );
  NANDN U1948 ( .A(n1043), .B(n1042), .Z(n1047) );
  NANDN U1949 ( .A(n1045), .B(n1044), .Z(n1046) );
  AND U1950 ( .A(n1047), .B(n1046), .Z(n1409) );
  NANDN U1951 ( .A(n1049), .B(n1048), .Z(n1053) );
  NANDN U1952 ( .A(n1051), .B(n1050), .Z(n1052) );
  NAND U1953 ( .A(n1053), .B(n1052), .Z(n1410) );
  XNOR U1954 ( .A(n1409), .B(n1410), .Z(n1412) );
  NANDN U1955 ( .A(n1055), .B(n1054), .Z(n1059) );
  NANDN U1956 ( .A(n1057), .B(n1056), .Z(n1058) );
  AND U1957 ( .A(n1059), .B(n1058), .Z(n1411) );
  XOR U1958 ( .A(n1412), .B(n1411), .Z(n1500) );
  NANDN U1959 ( .A(n1061), .B(n1060), .Z(n1065) );
  NAND U1960 ( .A(n1063), .B(n1062), .Z(n1064) );
  AND U1961 ( .A(n1065), .B(n1064), .Z(n1832) );
  NANDN U1962 ( .A(n1067), .B(n1066), .Z(n1071) );
  NANDN U1963 ( .A(n1069), .B(n1068), .Z(n1070) );
  NAND U1964 ( .A(n1071), .B(n1070), .Z(n1833) );
  XNOR U1965 ( .A(n1832), .B(n1833), .Z(n1835) );
  NANDN U1966 ( .A(n1073), .B(n1072), .Z(n1077) );
  NANDN U1967 ( .A(n1075), .B(n1074), .Z(n1076) );
  AND U1968 ( .A(n1077), .B(n1076), .Z(n1834) );
  XOR U1969 ( .A(n1835), .B(n1834), .Z(n1499) );
  NANDN U1970 ( .A(n1079), .B(n1078), .Z(n1083) );
  NANDN U1971 ( .A(n1081), .B(n1080), .Z(n1082) );
  AND U1972 ( .A(n1083), .B(n1082), .Z(n1433) );
  NANDN U1973 ( .A(n1085), .B(n1084), .Z(n1089) );
  NANDN U1974 ( .A(n1087), .B(n1086), .Z(n1088) );
  NAND U1975 ( .A(n1089), .B(n1088), .Z(n1434) );
  XNOR U1976 ( .A(n1433), .B(n1434), .Z(n1436) );
  NANDN U1977 ( .A(n1091), .B(n1090), .Z(n1095) );
  NANDN U1978 ( .A(n1093), .B(n1092), .Z(n1094) );
  AND U1979 ( .A(n1095), .B(n1094), .Z(n1435) );
  XNOR U1980 ( .A(n1436), .B(n1435), .Z(n1498) );
  XOR U1981 ( .A(n1499), .B(n1498), .Z(n1501) );
  XOR U1982 ( .A(n1500), .B(n1501), .Z(n1809) );
  NANDN U1983 ( .A(n1097), .B(n1096), .Z(n1101) );
  NAND U1984 ( .A(n1099), .B(n1098), .Z(n1100) );
  AND U1985 ( .A(n1101), .B(n1100), .Z(n1421) );
  NANDN U1986 ( .A(n1103), .B(n1102), .Z(n1107) );
  NAND U1987 ( .A(n1105), .B(n1104), .Z(n1106) );
  NAND U1988 ( .A(n1107), .B(n1106), .Z(n1422) );
  XNOR U1989 ( .A(n1421), .B(n1422), .Z(n1424) );
  NANDN U1990 ( .A(n1109), .B(n1108), .Z(n1113) );
  NAND U1991 ( .A(n1111), .B(n1110), .Z(n1112) );
  AND U1992 ( .A(n1113), .B(n1112), .Z(n1423) );
  XOR U1993 ( .A(n1424), .B(n1423), .Z(n1469) );
  NANDN U1994 ( .A(n1115), .B(n1114), .Z(n1119) );
  NANDN U1995 ( .A(n1117), .B(n1116), .Z(n1118) );
  AND U1996 ( .A(n1119), .B(n1118), .Z(n1379) );
  NANDN U1997 ( .A(n1121), .B(n1120), .Z(n1125) );
  NAND U1998 ( .A(n1123), .B(n1122), .Z(n1124) );
  NAND U1999 ( .A(n1125), .B(n1124), .Z(n1380) );
  XNOR U2000 ( .A(n1379), .B(n1380), .Z(n1382) );
  NANDN U2001 ( .A(n1127), .B(n1126), .Z(n1131) );
  NAND U2002 ( .A(n1129), .B(n1128), .Z(n1130) );
  AND U2003 ( .A(n1131), .B(n1130), .Z(n1381) );
  XOR U2004 ( .A(n1382), .B(n1381), .Z(n1468) );
  NANDN U2005 ( .A(n1133), .B(n1132), .Z(n1137) );
  NAND U2006 ( .A(n1135), .B(n1134), .Z(n1136) );
  AND U2007 ( .A(n1137), .B(n1136), .Z(n1557) );
  NANDN U2008 ( .A(n1139), .B(n1138), .Z(n1143) );
  NAND U2009 ( .A(n1141), .B(n1140), .Z(n1142) );
  NAND U2010 ( .A(n1143), .B(n1142), .Z(n1558) );
  XNOR U2011 ( .A(n1557), .B(n1558), .Z(n1560) );
  NANDN U2012 ( .A(n1145), .B(n1144), .Z(n1149) );
  NAND U2013 ( .A(n1147), .B(n1146), .Z(n1148) );
  AND U2014 ( .A(n1149), .B(n1148), .Z(n1559) );
  XNOR U2015 ( .A(n1560), .B(n1559), .Z(n1467) );
  XOR U2016 ( .A(n1468), .B(n1467), .Z(n1470) );
  XNOR U2017 ( .A(n1469), .B(n1470), .Z(n1808) );
  XNOR U2018 ( .A(n1809), .B(n1808), .Z(n1810) );
  XNOR U2019 ( .A(n1811), .B(n1810), .Z(n1637) );
  NANDN U2020 ( .A(n1151), .B(n1150), .Z(n1155) );
  NANDN U2021 ( .A(n1153), .B(n1152), .Z(n1154) );
  AND U2022 ( .A(n1155), .B(n1154), .Z(n1593) );
  NANDN U2023 ( .A(n1157), .B(n1156), .Z(n1161) );
  NANDN U2024 ( .A(n1159), .B(n1158), .Z(n1160) );
  NAND U2025 ( .A(n1161), .B(n1160), .Z(n1594) );
  XNOR U2026 ( .A(n1593), .B(n1594), .Z(n1596) );
  NANDN U2027 ( .A(n1163), .B(n1162), .Z(n1167) );
  NANDN U2028 ( .A(n1165), .B(n1164), .Z(n1166) );
  AND U2029 ( .A(n1167), .B(n1166), .Z(n1595) );
  XOR U2030 ( .A(n1596), .B(n1595), .Z(n1512) );
  NANDN U2031 ( .A(n1169), .B(n1168), .Z(n1173) );
  NAND U2032 ( .A(n1171), .B(n1170), .Z(n1172) );
  AND U2033 ( .A(n1173), .B(n1172), .Z(n1511) );
  NANDN U2034 ( .A(n1175), .B(n1174), .Z(n1179) );
  NAND U2035 ( .A(n1177), .B(n1176), .Z(n1178) );
  NAND U2036 ( .A(n1179), .B(n1178), .Z(n1607) );
  NANDN U2037 ( .A(n1181), .B(n1180), .Z(n1185) );
  NAND U2038 ( .A(n1183), .B(n1182), .Z(n1184) );
  AND U2039 ( .A(n1185), .B(n1184), .Z(n1606) );
  NANDN U2040 ( .A(n1187), .B(n1186), .Z(n1191) );
  NAND U2041 ( .A(n1189), .B(n1188), .Z(n1190) );
  NAND U2042 ( .A(n1191), .B(n1190), .Z(n1605) );
  XOR U2043 ( .A(n1606), .B(n1605), .Z(n1192) );
  XNOR U2044 ( .A(n1607), .B(n1192), .Z(n1510) );
  XOR U2045 ( .A(n1511), .B(n1510), .Z(n1513) );
  XOR U2046 ( .A(n1512), .B(n1513), .Z(n1866) );
  NANDN U2047 ( .A(n1194), .B(n1193), .Z(n1198) );
  NANDN U2048 ( .A(n1196), .B(n1195), .Z(n1197) );
  AND U2049 ( .A(n1198), .B(n1197), .Z(n1563) );
  NANDN U2050 ( .A(n1200), .B(n1199), .Z(n1204) );
  NAND U2051 ( .A(n1202), .B(n1201), .Z(n1203) );
  NAND U2052 ( .A(n1204), .B(n1203), .Z(n1564) );
  XNOR U2053 ( .A(n1563), .B(n1564), .Z(n1566) );
  NANDN U2054 ( .A(n1206), .B(n1205), .Z(n1210) );
  NAND U2055 ( .A(n1208), .B(n1207), .Z(n1209) );
  AND U2056 ( .A(n1210), .B(n1209), .Z(n1565) );
  XOR U2057 ( .A(n1566), .B(n1565), .Z(n1518) );
  NANDN U2058 ( .A(n1212), .B(n1211), .Z(n1216) );
  NAND U2059 ( .A(n1214), .B(n1213), .Z(n1215) );
  AND U2060 ( .A(n1216), .B(n1215), .Z(n1569) );
  NANDN U2061 ( .A(n1218), .B(n1217), .Z(n1222) );
  NAND U2062 ( .A(n1220), .B(n1219), .Z(n1221) );
  NAND U2063 ( .A(n1222), .B(n1221), .Z(n1570) );
  XNOR U2064 ( .A(n1569), .B(n1570), .Z(n1572) );
  NANDN U2065 ( .A(n1224), .B(n1223), .Z(n1228) );
  NAND U2066 ( .A(n1226), .B(n1225), .Z(n1227) );
  AND U2067 ( .A(n1228), .B(n1227), .Z(n1571) );
  XOR U2068 ( .A(n1572), .B(n1571), .Z(n1517) );
  NANDN U2069 ( .A(n1230), .B(n1229), .Z(n1234) );
  NAND U2070 ( .A(n1232), .B(n1231), .Z(n1233) );
  NAND U2071 ( .A(n1234), .B(n1233), .Z(n1620) );
  NANDN U2072 ( .A(n1236), .B(n1235), .Z(n1240) );
  NAND U2073 ( .A(n1238), .B(n1237), .Z(n1239) );
  AND U2074 ( .A(n1240), .B(n1239), .Z(n1619) );
  NANDN U2075 ( .A(n1242), .B(n1241), .Z(n1246) );
  NANDN U2076 ( .A(n1244), .B(n1243), .Z(n1245) );
  NAND U2077 ( .A(n1246), .B(n1245), .Z(n1618) );
  XOR U2078 ( .A(n1619), .B(n1618), .Z(n1247) );
  XNOR U2079 ( .A(n1620), .B(n1247), .Z(n1516) );
  XOR U2080 ( .A(n1517), .B(n1516), .Z(n1519) );
  XOR U2081 ( .A(n1518), .B(n1519), .Z(n1864) );
  NANDN U2082 ( .A(n1249), .B(n1248), .Z(n1253) );
  NAND U2083 ( .A(n1251), .B(n1250), .Z(n1252) );
  AND U2084 ( .A(n1253), .B(n1252), .Z(n1581) );
  NANDN U2085 ( .A(n1255), .B(n1254), .Z(n1259) );
  NAND U2086 ( .A(n1257), .B(n1256), .Z(n1258) );
  NAND U2087 ( .A(n1259), .B(n1258), .Z(n1582) );
  XNOR U2088 ( .A(n1581), .B(n1582), .Z(n1584) );
  NANDN U2089 ( .A(n1261), .B(n1260), .Z(n1265) );
  NAND U2090 ( .A(n1263), .B(n1262), .Z(n1264) );
  AND U2091 ( .A(n1265), .B(n1264), .Z(n1583) );
  XOR U2092 ( .A(n1584), .B(n1583), .Z(n1524) );
  NANDN U2093 ( .A(n1267), .B(n1266), .Z(n1271) );
  NANDN U2094 ( .A(n1269), .B(n1268), .Z(n1270) );
  AND U2095 ( .A(n1271), .B(n1270), .Z(n1523) );
  NANDN U2096 ( .A(n1273), .B(n1272), .Z(n1277) );
  NAND U2097 ( .A(n1275), .B(n1274), .Z(n1276) );
  AND U2098 ( .A(n1277), .B(n1276), .Z(n1540) );
  NANDN U2099 ( .A(n1279), .B(n1278), .Z(n1283) );
  NAND U2100 ( .A(n1281), .B(n1280), .Z(n1282) );
  NAND U2101 ( .A(n1283), .B(n1282), .Z(n1541) );
  XNOR U2102 ( .A(n1540), .B(n1541), .Z(n1543) );
  NANDN U2103 ( .A(n1284), .B(oglobal[0]), .Z(n1288) );
  NANDN U2104 ( .A(n1286), .B(n1285), .Z(n1287) );
  AND U2105 ( .A(n1288), .B(n1287), .Z(n1542) );
  XNOR U2106 ( .A(n1543), .B(n1542), .Z(n1522) );
  XOR U2107 ( .A(n1523), .B(n1522), .Z(n1525) );
  XNOR U2108 ( .A(n1524), .B(n1525), .Z(n1863) );
  XNOR U2109 ( .A(n1864), .B(n1863), .Z(n1865) );
  XOR U2110 ( .A(n1866), .B(n1865), .Z(n1640) );
  XNOR U2111 ( .A(n1639), .B(n1640), .Z(n1296) );
  XNOR U2112 ( .A(n1295), .B(n1296), .Z(n1298) );
  XOR U2113 ( .A(n1297), .B(n1298), .Z(n1291) );
  XOR U2114 ( .A(n1292), .B(n1291), .Z(o[1]) );
  NANDN U2115 ( .A(n1290), .B(n1289), .Z(n1294) );
  NAND U2116 ( .A(n1292), .B(n1291), .Z(n1293) );
  NAND U2117 ( .A(n1294), .B(n1293), .Z(n1974) );
  NAND U2118 ( .A(n1296), .B(n1295), .Z(n1300) );
  NANDN U2119 ( .A(n1298), .B(n1297), .Z(n1299) );
  AND U2120 ( .A(n1300), .B(n1299), .Z(n1963) );
  NAND U2121 ( .A(n1302), .B(n1301), .Z(n1306) );
  NAND U2122 ( .A(n1304), .B(n1303), .Z(n1305) );
  AND U2123 ( .A(n1306), .B(n1305), .Z(n1951) );
  NANDN U2124 ( .A(n1308), .B(n1307), .Z(n1312) );
  NANDN U2125 ( .A(n1310), .B(n1309), .Z(n1311) );
  AND U2126 ( .A(n1312), .B(n1311), .Z(n2048) );
  NANDN U2127 ( .A(n1314), .B(n1313), .Z(n1318) );
  NANDN U2128 ( .A(n1316), .B(n1315), .Z(n1317) );
  NAND U2129 ( .A(n1318), .B(n1317), .Z(n2049) );
  XNOR U2130 ( .A(n2048), .B(n2049), .Z(n2051) );
  NANDN U2131 ( .A(n1320), .B(n1319), .Z(n1324) );
  NANDN U2132 ( .A(n1322), .B(n1321), .Z(n1323) );
  AND U2133 ( .A(n1324), .B(n1323), .Z(n2050) );
  XOR U2134 ( .A(n2051), .B(n2050), .Z(n2118) );
  NANDN U2135 ( .A(n1326), .B(n1325), .Z(n1330) );
  NANDN U2136 ( .A(n1328), .B(n1327), .Z(n1329) );
  AND U2137 ( .A(n1330), .B(n1329), .Z(n2115) );
  NANDN U2138 ( .A(n1332), .B(n1331), .Z(n1336) );
  NANDN U2139 ( .A(n1334), .B(n1333), .Z(n1335) );
  AND U2140 ( .A(n1336), .B(n1335), .Z(n1934) );
  NANDN U2141 ( .A(n1338), .B(n1337), .Z(n1342) );
  OR U2142 ( .A(n1340), .B(n1339), .Z(n1341) );
  AND U2143 ( .A(n1342), .B(n1341), .Z(n1932) );
  NANDN U2144 ( .A(n1344), .B(n1343), .Z(n1348) );
  OR U2145 ( .A(n1346), .B(n1345), .Z(n1347) );
  NAND U2146 ( .A(n1348), .B(n1347), .Z(n1931) );
  XNOR U2147 ( .A(n1932), .B(n1931), .Z(n1933) );
  XOR U2148 ( .A(n1934), .B(n1933), .Z(n2116) );
  XNOR U2149 ( .A(n2115), .B(n2116), .Z(n2117) );
  XNOR U2150 ( .A(n2118), .B(n2117), .Z(n1950) );
  XNOR U2151 ( .A(n1951), .B(n1950), .Z(n1953) );
  NANDN U2152 ( .A(n1350), .B(n1349), .Z(n1354) );
  NANDN U2153 ( .A(n1352), .B(n1351), .Z(n1353) );
  NAND U2154 ( .A(n1354), .B(n1353), .Z(n2034) );
  NANDN U2155 ( .A(n1355), .B(oglobal[1]), .Z(n1359) );
  NANDN U2156 ( .A(n1357), .B(n1356), .Z(n1358) );
  AND U2157 ( .A(n1359), .B(n1358), .Z(n2033) );
  NANDN U2158 ( .A(n1361), .B(n1360), .Z(n1365) );
  NAND U2159 ( .A(n1363), .B(n1362), .Z(n1364) );
  NAND U2160 ( .A(n1365), .B(n1364), .Z(n2032) );
  IV U2161 ( .A(n2032), .Z(n2031) );
  XNOR U2162 ( .A(n2033), .B(n2031), .Z(n1366) );
  XNOR U2163 ( .A(n2034), .B(n1366), .Z(n2133) );
  NANDN U2164 ( .A(n1368), .B(n1367), .Z(n1372) );
  NAND U2165 ( .A(n1370), .B(n1369), .Z(n1371) );
  NAND U2166 ( .A(n1372), .B(n1371), .Z(n2134) );
  XNOR U2167 ( .A(n2133), .B(n2134), .Z(n2136) );
  NANDN U2168 ( .A(n1374), .B(n1373), .Z(n1378) );
  NAND U2169 ( .A(n1376), .B(n1375), .Z(n1377) );
  AND U2170 ( .A(n1378), .B(n1377), .Z(n2088) );
  NANDN U2171 ( .A(n1380), .B(n1379), .Z(n1384) );
  NAND U2172 ( .A(n1382), .B(n1381), .Z(n1383) );
  AND U2173 ( .A(n1384), .B(n1383), .Z(n2086) );
  NANDN U2174 ( .A(n1386), .B(n1385), .Z(n1390) );
  NAND U2175 ( .A(n1388), .B(n1387), .Z(n1389) );
  NAND U2176 ( .A(n1390), .B(n1389), .Z(n2085) );
  XNOR U2177 ( .A(n2086), .B(n2085), .Z(n2087) );
  XNOR U2178 ( .A(n2088), .B(n2087), .Z(n2135) );
  XOR U2179 ( .A(n2136), .B(n2135), .Z(n1920) );
  NANDN U2180 ( .A(n1392), .B(n1391), .Z(n1396) );
  NANDN U2181 ( .A(n1394), .B(n1393), .Z(n1395) );
  AND U2182 ( .A(n1396), .B(n1395), .Z(n1919) );
  XNOR U2183 ( .A(n1920), .B(n1919), .Z(n1921) );
  NANDN U2184 ( .A(n1398), .B(n1397), .Z(n1402) );
  NAND U2185 ( .A(n1400), .B(n1399), .Z(n1401) );
  AND U2186 ( .A(n1402), .B(n1401), .Z(n2075) );
  NANDN U2187 ( .A(n1404), .B(n1403), .Z(n1408) );
  NAND U2188 ( .A(n1406), .B(n1405), .Z(n1407) );
  AND U2189 ( .A(n1408), .B(n1407), .Z(n2074) );
  NANDN U2190 ( .A(n1410), .B(n1409), .Z(n1414) );
  NAND U2191 ( .A(n1412), .B(n1411), .Z(n1413) );
  NAND U2192 ( .A(n1414), .B(n1413), .Z(n2073) );
  XOR U2193 ( .A(n2074), .B(n2073), .Z(n2076) );
  XOR U2194 ( .A(n2075), .B(n2076), .Z(n2016) );
  NANDN U2195 ( .A(n1416), .B(n1415), .Z(n1420) );
  NANDN U2196 ( .A(n1418), .B(n1417), .Z(n1419) );
  AND U2197 ( .A(n1420), .B(n1419), .Z(n2014) );
  NANDN U2198 ( .A(n1422), .B(n1421), .Z(n1426) );
  NAND U2199 ( .A(n1424), .B(n1423), .Z(n1425) );
  AND U2200 ( .A(n1426), .B(n1425), .Z(n2081) );
  NANDN U2201 ( .A(n1428), .B(n1427), .Z(n1432) );
  NAND U2202 ( .A(n1430), .B(n1429), .Z(n1431) );
  AND U2203 ( .A(n1432), .B(n1431), .Z(n2080) );
  NANDN U2204 ( .A(n1434), .B(n1433), .Z(n1438) );
  NAND U2205 ( .A(n1436), .B(n1435), .Z(n1437) );
  NAND U2206 ( .A(n1438), .B(n1437), .Z(n2079) );
  XOR U2207 ( .A(n2080), .B(n2079), .Z(n2082) );
  XNOR U2208 ( .A(n2081), .B(n2082), .Z(n2013) );
  XNOR U2209 ( .A(n2014), .B(n2013), .Z(n2015) );
  XOR U2210 ( .A(n2016), .B(n2015), .Z(n1922) );
  XNOR U2211 ( .A(n1921), .B(n1922), .Z(n1952) );
  XOR U2212 ( .A(n1953), .B(n1952), .Z(n1873) );
  NANDN U2213 ( .A(n1440), .B(n1439), .Z(n1444) );
  NANDN U2214 ( .A(n1442), .B(n1441), .Z(n1443) );
  AND U2215 ( .A(n1444), .B(n1443), .Z(n1871) );
  XNOR U2216 ( .A(n1871), .B(n1870), .Z(n1872) );
  XNOR U2217 ( .A(n1873), .B(n1872), .Z(n1962) );
  XNOR U2218 ( .A(n1963), .B(n1962), .Z(n1965) );
  NANDN U2219 ( .A(n1450), .B(n1449), .Z(n1454) );
  NANDN U2220 ( .A(n1452), .B(n1451), .Z(n1453) );
  AND U2221 ( .A(n1454), .B(n1453), .Z(n1937) );
  NANDN U2222 ( .A(n1456), .B(n1455), .Z(n1460) );
  NANDN U2223 ( .A(n1458), .B(n1457), .Z(n1459) );
  NAND U2224 ( .A(n1460), .B(n1459), .Z(n1938) );
  XNOR U2225 ( .A(n1937), .B(n1938), .Z(n1939) );
  NANDN U2226 ( .A(n1462), .B(n1461), .Z(n1466) );
  NANDN U2227 ( .A(n1464), .B(n1463), .Z(n1465) );
  NAND U2228 ( .A(n1466), .B(n1465), .Z(n1940) );
  XOR U2229 ( .A(n1939), .B(n1940), .Z(n2054) );
  NANDN U2230 ( .A(n1468), .B(n1467), .Z(n1472) );
  OR U2231 ( .A(n1470), .B(n1469), .Z(n1471) );
  AND U2232 ( .A(n1472), .B(n1471), .Z(n1925) );
  NANDN U2233 ( .A(n1474), .B(n1473), .Z(n1478) );
  NANDN U2234 ( .A(n1476), .B(n1475), .Z(n1477) );
  NAND U2235 ( .A(n1478), .B(n1477), .Z(n1926) );
  XNOR U2236 ( .A(n1925), .B(n1926), .Z(n1927) );
  NANDN U2237 ( .A(n1480), .B(n1479), .Z(n1484) );
  NANDN U2238 ( .A(n1482), .B(n1481), .Z(n1483) );
  NAND U2239 ( .A(n1484), .B(n1483), .Z(n1928) );
  XNOR U2240 ( .A(n1927), .B(n1928), .Z(n2056) );
  NANDN U2241 ( .A(n1486), .B(n1485), .Z(n1490) );
  NANDN U2242 ( .A(n1488), .B(n1487), .Z(n1489) );
  AND U2243 ( .A(n1490), .B(n1489), .Z(n2055) );
  XNOR U2244 ( .A(n2056), .B(n2055), .Z(n1491) );
  XNOR U2245 ( .A(n2054), .B(n1491), .Z(n1958) );
  NANDN U2246 ( .A(n1493), .B(n1492), .Z(n1497) );
  OR U2247 ( .A(n1495), .B(n1494), .Z(n1496) );
  AND U2248 ( .A(n1497), .B(n1496), .Z(n2129) );
  NANDN U2249 ( .A(n1499), .B(n1498), .Z(n1503) );
  OR U2250 ( .A(n1501), .B(n1500), .Z(n1502) );
  AND U2251 ( .A(n1503), .B(n1502), .Z(n2128) );
  NANDN U2252 ( .A(n1505), .B(n1504), .Z(n1509) );
  NANDN U2253 ( .A(n1507), .B(n1506), .Z(n1508) );
  NAND U2254 ( .A(n1509), .B(n1508), .Z(n2127) );
  XOR U2255 ( .A(n2128), .B(n2127), .Z(n2130) );
  XOR U2256 ( .A(n2129), .B(n2130), .Z(n2020) );
  NANDN U2257 ( .A(n1511), .B(n1510), .Z(n1515) );
  OR U2258 ( .A(n1513), .B(n1512), .Z(n1514) );
  AND U2259 ( .A(n1515), .B(n1514), .Z(n2123) );
  NANDN U2260 ( .A(n1517), .B(n1516), .Z(n1521) );
  OR U2261 ( .A(n1519), .B(n1518), .Z(n1520) );
  AND U2262 ( .A(n1521), .B(n1520), .Z(n2122) );
  NANDN U2263 ( .A(n1523), .B(n1522), .Z(n1527) );
  OR U2264 ( .A(n1525), .B(n1524), .Z(n1526) );
  NAND U2265 ( .A(n1527), .B(n1526), .Z(n2121) );
  XOR U2266 ( .A(n2122), .B(n2121), .Z(n2124) );
  XNOR U2267 ( .A(n2123), .B(n2124), .Z(n2019) );
  XNOR U2268 ( .A(n2020), .B(n2019), .Z(n2022) );
  NANDN U2269 ( .A(n1529), .B(n1528), .Z(n1533) );
  NAND U2270 ( .A(n1531), .B(n1530), .Z(n1532) );
  AND U2271 ( .A(n1533), .B(n1532), .Z(n2021) );
  XOR U2272 ( .A(n2022), .B(n2021), .Z(n1957) );
  NANDN U2273 ( .A(n1535), .B(n1534), .Z(n1539) );
  NANDN U2274 ( .A(n1537), .B(n1536), .Z(n1538) );
  NAND U2275 ( .A(n1539), .B(n1538), .Z(n1891) );
  NANDN U2276 ( .A(n1541), .B(n1540), .Z(n1545) );
  NAND U2277 ( .A(n1543), .B(n1542), .Z(n1544) );
  NAND U2278 ( .A(n1545), .B(n1544), .Z(n2036) );
  XNOR U2279 ( .A(n2035), .B(oglobal[2]), .Z(n1549) );
  XNOR U2280 ( .A(n2036), .B(n1549), .Z(n1889) );
  IV U2281 ( .A(n1889), .Z(n1888) );
  NANDN U2282 ( .A(n1551), .B(n1550), .Z(n1555) );
  NAND U2283 ( .A(n1553), .B(n1552), .Z(n1554) );
  AND U2284 ( .A(n1555), .B(n1554), .Z(n1890) );
  XNOR U2285 ( .A(n1888), .B(n1890), .Z(n1556) );
  XNOR U2286 ( .A(n1891), .B(n1556), .Z(n1998) );
  NANDN U2287 ( .A(n1558), .B(n1557), .Z(n1562) );
  NAND U2288 ( .A(n1560), .B(n1559), .Z(n1561) );
  AND U2289 ( .A(n1562), .B(n1561), .Z(n1909) );
  NANDN U2290 ( .A(n1564), .B(n1563), .Z(n1568) );
  NAND U2291 ( .A(n1566), .B(n1565), .Z(n1567) );
  AND U2292 ( .A(n1568), .B(n1567), .Z(n1908) );
  NANDN U2293 ( .A(n1570), .B(n1569), .Z(n1574) );
  NAND U2294 ( .A(n1572), .B(n1571), .Z(n1573) );
  NAND U2295 ( .A(n1574), .B(n1573), .Z(n1907) );
  XOR U2296 ( .A(n1908), .B(n1907), .Z(n1910) );
  XOR U2297 ( .A(n1909), .B(n1910), .Z(n1898) );
  NANDN U2298 ( .A(n1576), .B(n1575), .Z(n1580) );
  NAND U2299 ( .A(n1578), .B(n1577), .Z(n1579) );
  AND U2300 ( .A(n1580), .B(n1579), .Z(n1903) );
  NANDN U2301 ( .A(n1582), .B(n1581), .Z(n1586) );
  NAND U2302 ( .A(n1584), .B(n1583), .Z(n1585) );
  AND U2303 ( .A(n1586), .B(n1585), .Z(n1902) );
  NANDN U2304 ( .A(n1588), .B(n1587), .Z(n1592) );
  NAND U2305 ( .A(n1590), .B(n1589), .Z(n1591) );
  NAND U2306 ( .A(n1592), .B(n1591), .Z(n1901) );
  XOR U2307 ( .A(n1902), .B(n1901), .Z(n1904) );
  XOR U2308 ( .A(n1903), .B(n1904), .Z(n1896) );
  NANDN U2309 ( .A(n1594), .B(n1593), .Z(n1598) );
  NAND U2310 ( .A(n1596), .B(n1595), .Z(n1597) );
  AND U2311 ( .A(n1598), .B(n1597), .Z(n1895) );
  XNOR U2312 ( .A(n1896), .B(n1895), .Z(n1897) );
  XNOR U2313 ( .A(n1898), .B(n1897), .Z(n1995) );
  NANDN U2314 ( .A(n1600), .B(n1599), .Z(n1604) );
  NAND U2315 ( .A(n1602), .B(n1601), .Z(n1603) );
  AND U2316 ( .A(n1604), .B(n1603), .Z(n2046) );
  XNOR U2317 ( .A(n2045), .B(n2044), .Z(n1611) );
  XNOR U2318 ( .A(n2046), .B(n1611), .Z(n2099) );
  NANDN U2319 ( .A(n1613), .B(n1612), .Z(n1617) );
  NAND U2320 ( .A(n1615), .B(n1614), .Z(n1616) );
  NAND U2321 ( .A(n1617), .B(n1616), .Z(n2062) );
  XNOR U2322 ( .A(n2061), .B(n2060), .Z(n1624) );
  XNOR U2323 ( .A(n2062), .B(n1624), .Z(n2097) );
  NANDN U2324 ( .A(n1626), .B(n1625), .Z(n1630) );
  OR U2325 ( .A(n1628), .B(n1627), .Z(n1629) );
  AND U2326 ( .A(n1630), .B(n1629), .Z(n2098) );
  XOR U2327 ( .A(n2097), .B(n2098), .Z(n2100) );
  XOR U2328 ( .A(n2099), .B(n2100), .Z(n1996) );
  XNOR U2329 ( .A(n1995), .B(n1996), .Z(n1997) );
  XOR U2330 ( .A(n1998), .B(n1997), .Z(n1956) );
  XNOR U2331 ( .A(n1957), .B(n1956), .Z(n1959) );
  XNOR U2332 ( .A(n1958), .B(n1959), .Z(n1978) );
  NAND U2333 ( .A(n1632), .B(n1631), .Z(n1636) );
  NAND U2334 ( .A(n1634), .B(n1633), .Z(n1635) );
  NAND U2335 ( .A(n1636), .B(n1635), .Z(n1985) );
  NAND U2336 ( .A(n1638), .B(n1637), .Z(n1642) );
  NANDN U2337 ( .A(n1640), .B(n1639), .Z(n1641) );
  NAND U2338 ( .A(n1642), .B(n1641), .Z(n1983) );
  NANDN U2339 ( .A(n1644), .B(n1643), .Z(n1648) );
  NAND U2340 ( .A(n1646), .B(n1645), .Z(n1647) );
  AND U2341 ( .A(n1648), .B(n1647), .Z(n2059) );
  NANDN U2342 ( .A(n1650), .B(n1649), .Z(n1654) );
  NAND U2343 ( .A(n1652), .B(n1651), .Z(n1653) );
  AND U2344 ( .A(n1654), .B(n1653), .Z(n2057) );
  NANDN U2345 ( .A(n1656), .B(n1655), .Z(n1660) );
  NAND U2346 ( .A(n1658), .B(n1657), .Z(n1659) );
  AND U2347 ( .A(n1660), .B(n1659), .Z(n2058) );
  XNOR U2348 ( .A(n2057), .B(n2058), .Z(n1661) );
  XNOR U2349 ( .A(n2059), .B(n1661), .Z(n2094) );
  NANDN U2350 ( .A(n1663), .B(n1662), .Z(n1667) );
  NAND U2351 ( .A(n1665), .B(n1664), .Z(n1666) );
  AND U2352 ( .A(n1667), .B(n1666), .Z(n2043) );
  NANDN U2353 ( .A(n1669), .B(n1668), .Z(n1673) );
  NAND U2354 ( .A(n1671), .B(n1670), .Z(n1672) );
  NAND U2355 ( .A(n1673), .B(n1672), .Z(n2042) );
  NANDN U2356 ( .A(n1675), .B(n1674), .Z(n1679) );
  NAND U2357 ( .A(n1677), .B(n1676), .Z(n1678) );
  AND U2358 ( .A(n1679), .B(n1678), .Z(n2041) );
  XOR U2359 ( .A(n2042), .B(n2041), .Z(n1680) );
  XNOR U2360 ( .A(n2043), .B(n1680), .Z(n2091) );
  NANDN U2361 ( .A(n1682), .B(n1681), .Z(n1686) );
  NAND U2362 ( .A(n1684), .B(n1683), .Z(n1685) );
  AND U2363 ( .A(n1686), .B(n1685), .Z(n2092) );
  XNOR U2364 ( .A(n2091), .B(n2092), .Z(n2093) );
  XOR U2365 ( .A(n2094), .B(n2093), .Z(n1947) );
  NANDN U2366 ( .A(n1688), .B(n1687), .Z(n1692) );
  NAND U2367 ( .A(n1690), .B(n1689), .Z(n1691) );
  NAND U2368 ( .A(n1692), .B(n1691), .Z(n2065) );
  XNOR U2369 ( .A(n2064), .B(n2063), .Z(n1699) );
  XNOR U2370 ( .A(n2065), .B(n1699), .Z(n2004) );
  NANDN U2371 ( .A(n1701), .B(n1700), .Z(n1705) );
  NANDN U2372 ( .A(n1703), .B(n1702), .Z(n1704) );
  AND U2373 ( .A(n1705), .B(n1704), .Z(n2002) );
  NANDN U2374 ( .A(n1707), .B(n1706), .Z(n1711) );
  NAND U2375 ( .A(n1709), .B(n1708), .Z(n1710) );
  NAND U2376 ( .A(n1711), .B(n1710), .Z(n2068) );
  NANDN U2377 ( .A(n1713), .B(n1712), .Z(n1717) );
  NAND U2378 ( .A(n1715), .B(n1714), .Z(n1716) );
  NAND U2379 ( .A(n1717), .B(n1716), .Z(n2067) );
  XOR U2380 ( .A(n2068), .B(n2067), .Z(n2070) );
  NANDN U2381 ( .A(n1719), .B(n1718), .Z(n1723) );
  NAND U2382 ( .A(n1721), .B(n1720), .Z(n1722) );
  NAND U2383 ( .A(n1723), .B(n1722), .Z(n2069) );
  XNOR U2384 ( .A(n2070), .B(n2069), .Z(n2001) );
  XNOR U2385 ( .A(n2002), .B(n2001), .Z(n2003) );
  XOR U2386 ( .A(n2004), .B(n2003), .Z(n1945) );
  NAND U2387 ( .A(n1725), .B(n1724), .Z(n1729) );
  NAND U2388 ( .A(n1727), .B(n1726), .Z(n1728) );
  AND U2389 ( .A(n1729), .B(n1728), .Z(n2009) );
  NANDN U2390 ( .A(n1731), .B(n1730), .Z(n1735) );
  NANDN U2391 ( .A(n1733), .B(n1732), .Z(n1734) );
  AND U2392 ( .A(n1735), .B(n1734), .Z(n2008) );
  NANDN U2393 ( .A(n1737), .B(n1736), .Z(n1741) );
  NAND U2394 ( .A(n1739), .B(n1738), .Z(n1740) );
  NAND U2395 ( .A(n1741), .B(n1740), .Z(n2007) );
  XOR U2396 ( .A(n2008), .B(n2007), .Z(n2010) );
  XNOR U2397 ( .A(n2009), .B(n2010), .Z(n1944) );
  XNOR U2398 ( .A(n1945), .B(n1944), .Z(n1946) );
  XNOR U2399 ( .A(n1947), .B(n1946), .Z(n1984) );
  XOR U2400 ( .A(n1983), .B(n1984), .Z(n1986) );
  XOR U2401 ( .A(n1985), .B(n1986), .Z(n1977) );
  NANDN U2402 ( .A(n1743), .B(n1742), .Z(n1747) );
  NANDN U2403 ( .A(n1745), .B(n1744), .Z(n1746) );
  AND U2404 ( .A(n1747), .B(n1746), .Z(n1885) );
  NANDN U2405 ( .A(n1749), .B(n1748), .Z(n1753) );
  NAND U2406 ( .A(n1751), .B(n1750), .Z(n1752) );
  AND U2407 ( .A(n1753), .B(n1752), .Z(n1883) );
  NAND U2408 ( .A(n1755), .B(n1754), .Z(n1759) );
  NAND U2409 ( .A(n1757), .B(n1756), .Z(n1758) );
  NAND U2410 ( .A(n1759), .B(n1758), .Z(n1882) );
  XNOR U2411 ( .A(n1883), .B(n1882), .Z(n1884) );
  XNOR U2412 ( .A(n1885), .B(n1884), .Z(n1992) );
  NANDN U2413 ( .A(n1761), .B(n1760), .Z(n1765) );
  NANDN U2414 ( .A(n1763), .B(n1762), .Z(n1764) );
  AND U2415 ( .A(n1765), .B(n1764), .Z(n1879) );
  NANDN U2416 ( .A(n1767), .B(n1766), .Z(n1771) );
  NAND U2417 ( .A(n1769), .B(n1768), .Z(n1770) );
  AND U2418 ( .A(n1771), .B(n1770), .Z(n1877) );
  NANDN U2419 ( .A(n1773), .B(n1772), .Z(n1777) );
  NAND U2420 ( .A(n1775), .B(n1774), .Z(n1776) );
  NAND U2421 ( .A(n1777), .B(n1776), .Z(n1876) );
  XNOR U2422 ( .A(n1877), .B(n1876), .Z(n1878) );
  XOR U2423 ( .A(n1879), .B(n1878), .Z(n1990) );
  NAND U2424 ( .A(n1779), .B(n1778), .Z(n1783) );
  NAND U2425 ( .A(n1781), .B(n1780), .Z(n1782) );
  AND U2426 ( .A(n1783), .B(n1782), .Z(n1989) );
  XOR U2427 ( .A(n1992), .B(n1991), .Z(n1979) );
  XOR U2428 ( .A(n1980), .B(n1979), .Z(n1964) );
  XOR U2429 ( .A(n1965), .B(n1964), .Z(n1975) );
  NANDN U2430 ( .A(n1785), .B(n1784), .Z(n1789) );
  NAND U2431 ( .A(n1787), .B(n1786), .Z(n1788) );
  AND U2432 ( .A(n1789), .B(n1788), .Z(n1971) );
  NAND U2433 ( .A(n1791), .B(n1790), .Z(n1795) );
  NANDN U2434 ( .A(n1793), .B(n1792), .Z(n1794) );
  AND U2435 ( .A(n1795), .B(n1794), .Z(n1969) );
  NAND U2436 ( .A(n1797), .B(n1796), .Z(n1801) );
  NAND U2437 ( .A(n1799), .B(n1798), .Z(n1800) );
  AND U2438 ( .A(n1801), .B(n1800), .Z(n2140) );
  NANDN U2439 ( .A(n1803), .B(n1802), .Z(n1807) );
  NANDN U2440 ( .A(n1805), .B(n1804), .Z(n1806) );
  AND U2441 ( .A(n1807), .B(n1806), .Z(n2112) );
  NANDN U2442 ( .A(n1809), .B(n1808), .Z(n1813) );
  NANDN U2443 ( .A(n1811), .B(n1810), .Z(n1812) );
  AND U2444 ( .A(n1813), .B(n1812), .Z(n2109) );
  NANDN U2445 ( .A(n1815), .B(n1814), .Z(n1819) );
  NAND U2446 ( .A(n1817), .B(n1816), .Z(n1818) );
  AND U2447 ( .A(n1819), .B(n1818), .Z(n1915) );
  NANDN U2448 ( .A(n1821), .B(n1820), .Z(n1825) );
  NAND U2449 ( .A(n1823), .B(n1822), .Z(n1824) );
  AND U2450 ( .A(n1825), .B(n1824), .Z(n1914) );
  NANDN U2451 ( .A(n1827), .B(n1826), .Z(n1831) );
  NAND U2452 ( .A(n1829), .B(n1828), .Z(n1830) );
  NAND U2453 ( .A(n1831), .B(n1830), .Z(n1913) );
  XOR U2454 ( .A(n1914), .B(n1913), .Z(n1916) );
  XOR U2455 ( .A(n1915), .B(n1916), .Z(n2106) );
  NANDN U2456 ( .A(n1833), .B(n1832), .Z(n1837) );
  NAND U2457 ( .A(n1835), .B(n1834), .Z(n1836) );
  AND U2458 ( .A(n1837), .B(n1836), .Z(n2039) );
  XNOR U2459 ( .A(n2038), .B(n2037), .Z(n1844) );
  XNOR U2460 ( .A(n2039), .B(n1844), .Z(n2103) );
  NANDN U2461 ( .A(n1846), .B(n1845), .Z(n1850) );
  NANDN U2462 ( .A(n1848), .B(n1847), .Z(n1849) );
  AND U2463 ( .A(n1850), .B(n1849), .Z(n2104) );
  XNOR U2464 ( .A(n2103), .B(n2104), .Z(n2105) );
  XOR U2465 ( .A(n2106), .B(n2105), .Z(n2110) );
  XNOR U2466 ( .A(n2109), .B(n2110), .Z(n2111) );
  XOR U2467 ( .A(n2112), .B(n2111), .Z(n2139) );
  XNOR U2468 ( .A(n2140), .B(n2139), .Z(n2142) );
  NANDN U2469 ( .A(n1852), .B(n1851), .Z(n1856) );
  NAND U2470 ( .A(n1854), .B(n1853), .Z(n1855) );
  AND U2471 ( .A(n1856), .B(n1855), .Z(n2028) );
  NANDN U2472 ( .A(n1858), .B(n1857), .Z(n1862) );
  NANDN U2473 ( .A(n1860), .B(n1859), .Z(n1861) );
  AND U2474 ( .A(n1862), .B(n1861), .Z(n2026) );
  NANDN U2475 ( .A(n1864), .B(n1863), .Z(n1868) );
  NANDN U2476 ( .A(n1866), .B(n1865), .Z(n1867) );
  AND U2477 ( .A(n1868), .B(n1867), .Z(n2025) );
  XNOR U2478 ( .A(n2026), .B(n2025), .Z(n2027) );
  XNOR U2479 ( .A(n2028), .B(n2027), .Z(n2141) );
  XNOR U2480 ( .A(n2142), .B(n2141), .Z(n1968) );
  XNOR U2481 ( .A(n1969), .B(n1968), .Z(n1970) );
  XNOR U2482 ( .A(n1971), .B(n1970), .Z(n1976) );
  XNOR U2483 ( .A(n1975), .B(n1976), .Z(n1869) );
  XNOR U2484 ( .A(n1974), .B(n1869), .Z(o[2]) );
  NANDN U2485 ( .A(n1871), .B(n1870), .Z(n1875) );
  NANDN U2486 ( .A(n1873), .B(n1872), .Z(n1874) );
  NAND U2487 ( .A(n1875), .B(n1874), .Z(n2262) );
  NANDN U2488 ( .A(n1877), .B(n1876), .Z(n1881) );
  NANDN U2489 ( .A(n1879), .B(n1878), .Z(n1880) );
  AND U2490 ( .A(n1881), .B(n1880), .Z(n2255) );
  NANDN U2491 ( .A(n1883), .B(n1882), .Z(n1887) );
  NANDN U2492 ( .A(n1885), .B(n1884), .Z(n1886) );
  AND U2493 ( .A(n1887), .B(n1886), .Z(n2254) );
  XNOR U2494 ( .A(n2255), .B(n2254), .Z(n2256) );
  NANDN U2495 ( .A(n1890), .B(n1888), .Z(n1894) );
  AND U2496 ( .A(n1890), .B(n1889), .Z(n1892) );
  OR U2497 ( .A(n1892), .B(n1891), .Z(n1893) );
  AND U2498 ( .A(n1894), .B(n1893), .Z(n2227) );
  NANDN U2499 ( .A(n1896), .B(n1895), .Z(n1900) );
  NANDN U2500 ( .A(n1898), .B(n1897), .Z(n1899) );
  AND U2501 ( .A(n1900), .B(n1899), .Z(n2225) );
  NANDN U2502 ( .A(n1902), .B(n1901), .Z(n1906) );
  OR U2503 ( .A(n1904), .B(n1903), .Z(n1905) );
  AND U2504 ( .A(n1906), .B(n1905), .Z(n2196) );
  NANDN U2505 ( .A(n1908), .B(n1907), .Z(n1912) );
  OR U2506 ( .A(n1910), .B(n1909), .Z(n1911) );
  AND U2507 ( .A(n1912), .B(n1911), .Z(n2194) );
  NANDN U2508 ( .A(n1914), .B(n1913), .Z(n1918) );
  OR U2509 ( .A(n1916), .B(n1915), .Z(n1917) );
  NAND U2510 ( .A(n1918), .B(n1917), .Z(n2195) );
  XOR U2511 ( .A(n2194), .B(n2195), .Z(n2197) );
  XNOR U2512 ( .A(n2196), .B(n2197), .Z(n2224) );
  XNOR U2513 ( .A(n2225), .B(n2224), .Z(n2226) );
  XOR U2514 ( .A(n2227), .B(n2226), .Z(n2257) );
  XOR U2515 ( .A(n2256), .B(n2257), .Z(n2261) );
  NANDN U2516 ( .A(n1920), .B(n1919), .Z(n1924) );
  NANDN U2517 ( .A(n1922), .B(n1921), .Z(n1923) );
  NAND U2518 ( .A(n1924), .B(n1923), .Z(n2167) );
  NANDN U2519 ( .A(n1926), .B(n1925), .Z(n1930) );
  NANDN U2520 ( .A(n1928), .B(n1927), .Z(n1929) );
  NAND U2521 ( .A(n1930), .B(n1929), .Z(n2223) );
  NANDN U2522 ( .A(n1932), .B(n1931), .Z(n1936) );
  NANDN U2523 ( .A(n1934), .B(n1933), .Z(n1935) );
  AND U2524 ( .A(n1936), .B(n1935), .Z(n2222) );
  NANDN U2525 ( .A(n1938), .B(n1937), .Z(n1942) );
  NANDN U2526 ( .A(n1940), .B(n1939), .Z(n1941) );
  NAND U2527 ( .A(n1942), .B(n1941), .Z(n2221) );
  IV U2528 ( .A(n2221), .Z(n2220) );
  XNOR U2529 ( .A(n2222), .B(n2220), .Z(n1943) );
  XNOR U2530 ( .A(n2223), .B(n1943), .Z(n2164) );
  NANDN U2531 ( .A(n1945), .B(n1944), .Z(n1949) );
  NANDN U2532 ( .A(n1947), .B(n1946), .Z(n1948) );
  NAND U2533 ( .A(n1949), .B(n1948), .Z(n2165) );
  XNOR U2534 ( .A(n2164), .B(n2165), .Z(n2166) );
  XNOR U2535 ( .A(n2167), .B(n2166), .Z(n2260) );
  XOR U2536 ( .A(n2262), .B(n2263), .Z(n2154) );
  NANDN U2537 ( .A(n1951), .B(n1950), .Z(n1955) );
  NAND U2538 ( .A(n1953), .B(n1952), .Z(n1954) );
  AND U2539 ( .A(n1955), .B(n1954), .Z(n2153) );
  NANDN U2540 ( .A(n1957), .B(n1956), .Z(n1961) );
  NAND U2541 ( .A(n1959), .B(n1958), .Z(n1960) );
  NAND U2542 ( .A(n1961), .B(n1960), .Z(n2152) );
  XNOR U2543 ( .A(n2153), .B(n2152), .Z(n2155) );
  XNOR U2544 ( .A(n2154), .B(n2155), .Z(n2277) );
  NANDN U2545 ( .A(n1963), .B(n1962), .Z(n1967) );
  NAND U2546 ( .A(n1965), .B(n1964), .Z(n1966) );
  AND U2547 ( .A(n1967), .B(n1966), .Z(n2276) );
  NANDN U2548 ( .A(n1969), .B(n1968), .Z(n1973) );
  NANDN U2549 ( .A(n1971), .B(n1970), .Z(n1972) );
  NAND U2550 ( .A(n1973), .B(n1972), .Z(n2275) );
  XNOR U2551 ( .A(n2276), .B(n2275), .Z(n2278) );
  XNOR U2552 ( .A(n2277), .B(n2278), .Z(n2274) );
  NAND U2553 ( .A(n1978), .B(n1977), .Z(n1982) );
  NAND U2554 ( .A(n1980), .B(n1979), .Z(n1981) );
  NAND U2555 ( .A(n1982), .B(n1981), .Z(n2148) );
  NAND U2556 ( .A(n1984), .B(n1983), .Z(n1988) );
  NAND U2557 ( .A(n1986), .B(n1985), .Z(n1987) );
  NAND U2558 ( .A(n1988), .B(n1987), .Z(n2268) );
  NAND U2559 ( .A(n1990), .B(n1989), .Z(n1994) );
  NAND U2560 ( .A(n1992), .B(n1991), .Z(n1993) );
  NAND U2561 ( .A(n1994), .B(n1993), .Z(n2266) );
  NANDN U2562 ( .A(n1996), .B(n1995), .Z(n2000) );
  NAND U2563 ( .A(n1998), .B(n1997), .Z(n1999) );
  AND U2564 ( .A(n2000), .B(n1999), .Z(n2245) );
  NANDN U2565 ( .A(n2002), .B(n2001), .Z(n2006) );
  NAND U2566 ( .A(n2004), .B(n2003), .Z(n2005) );
  AND U2567 ( .A(n2006), .B(n2005), .Z(n2238) );
  NANDN U2568 ( .A(n2008), .B(n2007), .Z(n2012) );
  OR U2569 ( .A(n2010), .B(n2009), .Z(n2011) );
  AND U2570 ( .A(n2012), .B(n2011), .Z(n2237) );
  NANDN U2571 ( .A(n2014), .B(n2013), .Z(n2018) );
  NANDN U2572 ( .A(n2016), .B(n2015), .Z(n2017) );
  NAND U2573 ( .A(n2018), .B(n2017), .Z(n2236) );
  XOR U2574 ( .A(n2237), .B(n2236), .Z(n2239) );
  XOR U2575 ( .A(n2238), .B(n2239), .Z(n2243) );
  NANDN U2576 ( .A(n2020), .B(n2019), .Z(n2024) );
  NAND U2577 ( .A(n2022), .B(n2021), .Z(n2023) );
  NAND U2578 ( .A(n2024), .B(n2023), .Z(n2242) );
  XNOR U2579 ( .A(n2243), .B(n2242), .Z(n2244) );
  XOR U2580 ( .A(n2245), .B(n2244), .Z(n2267) );
  XOR U2581 ( .A(n2266), .B(n2267), .Z(n2269) );
  XOR U2582 ( .A(n2268), .B(n2269), .Z(n2147) );
  NANDN U2583 ( .A(n2026), .B(n2025), .Z(n2030) );
  NANDN U2584 ( .A(n2028), .B(n2027), .Z(n2029) );
  AND U2585 ( .A(n2030), .B(n2029), .Z(n2161) );
  XNOR U2586 ( .A(n2210), .B(n2209), .Z(n2040) );
  XOR U2587 ( .A(n2211), .B(n2040), .Z(n2191) );
  XNOR U2588 ( .A(n2212), .B(oglobal[3]), .Z(n2047) );
  XOR U2589 ( .A(n2213), .B(n2047), .Z(n2189) );
  NANDN U2590 ( .A(n2049), .B(n2048), .Z(n2053) );
  NAND U2591 ( .A(n2051), .B(n2050), .Z(n2052) );
  AND U2592 ( .A(n2053), .B(n2052), .Z(n2188) );
  XNOR U2593 ( .A(n2189), .B(n2188), .Z(n2190) );
  XNOR U2594 ( .A(n2191), .B(n2190), .Z(n2172) );
  XNOR U2595 ( .A(n2207), .B(n2206), .Z(n2066) );
  XOR U2596 ( .A(n2208), .B(n2066), .Z(n2215) );
  NAND U2597 ( .A(n2068), .B(n2067), .Z(n2072) );
  NAND U2598 ( .A(n2070), .B(n2069), .Z(n2071) );
  AND U2599 ( .A(n2072), .B(n2071), .Z(n2214) );
  XNOR U2600 ( .A(n2215), .B(n2214), .Z(n2216) );
  NANDN U2601 ( .A(n2074), .B(n2073), .Z(n2078) );
  OR U2602 ( .A(n2076), .B(n2075), .Z(n2077) );
  AND U2603 ( .A(n2078), .B(n2077), .Z(n2202) );
  NANDN U2604 ( .A(n2080), .B(n2079), .Z(n2084) );
  OR U2605 ( .A(n2082), .B(n2081), .Z(n2083) );
  AND U2606 ( .A(n2084), .B(n2083), .Z(n2200) );
  NANDN U2607 ( .A(n2086), .B(n2085), .Z(n2090) );
  NANDN U2608 ( .A(n2088), .B(n2087), .Z(n2089) );
  NAND U2609 ( .A(n2090), .B(n2089), .Z(n2201) );
  XOR U2610 ( .A(n2200), .B(n2201), .Z(n2203) );
  XOR U2611 ( .A(n2202), .B(n2203), .Z(n2217) );
  XNOR U2612 ( .A(n2216), .B(n2217), .Z(n2170) );
  XOR U2613 ( .A(n2171), .B(n2170), .Z(n2173) );
  XNOR U2614 ( .A(n2172), .B(n2173), .Z(n2158) );
  NANDN U2615 ( .A(n2092), .B(n2091), .Z(n2096) );
  NAND U2616 ( .A(n2094), .B(n2093), .Z(n2095) );
  AND U2617 ( .A(n2096), .B(n2095), .Z(n2233) );
  NANDN U2618 ( .A(n2098), .B(n2097), .Z(n2102) );
  NANDN U2619 ( .A(n2100), .B(n2099), .Z(n2101) );
  AND U2620 ( .A(n2102), .B(n2101), .Z(n2231) );
  NANDN U2621 ( .A(n2104), .B(n2103), .Z(n2108) );
  NANDN U2622 ( .A(n2106), .B(n2105), .Z(n2107) );
  NAND U2623 ( .A(n2108), .B(n2107), .Z(n2230) );
  XNOR U2624 ( .A(n2231), .B(n2230), .Z(n2232) );
  XOR U2625 ( .A(n2233), .B(n2232), .Z(n2159) );
  XNOR U2626 ( .A(n2158), .B(n2159), .Z(n2160) );
  XOR U2627 ( .A(n2161), .B(n2160), .Z(n2178) );
  NANDN U2628 ( .A(n2110), .B(n2109), .Z(n2114) );
  NAND U2629 ( .A(n2112), .B(n2111), .Z(n2113) );
  AND U2630 ( .A(n2114), .B(n2113), .Z(n2251) );
  NANDN U2631 ( .A(n2116), .B(n2115), .Z(n2120) );
  NANDN U2632 ( .A(n2118), .B(n2117), .Z(n2119) );
  AND U2633 ( .A(n2120), .B(n2119), .Z(n2249) );
  NANDN U2634 ( .A(n2122), .B(n2121), .Z(n2126) );
  OR U2635 ( .A(n2124), .B(n2123), .Z(n2125) );
  AND U2636 ( .A(n2126), .B(n2125), .Z(n2185) );
  NANDN U2637 ( .A(n2128), .B(n2127), .Z(n2132) );
  OR U2638 ( .A(n2130), .B(n2129), .Z(n2131) );
  AND U2639 ( .A(n2132), .B(n2131), .Z(n2183) );
  NANDN U2640 ( .A(n2134), .B(n2133), .Z(n2138) );
  NAND U2641 ( .A(n2136), .B(n2135), .Z(n2137) );
  AND U2642 ( .A(n2138), .B(n2137), .Z(n2182) );
  XNOR U2643 ( .A(n2183), .B(n2182), .Z(n2184) );
  XNOR U2644 ( .A(n2185), .B(n2184), .Z(n2248) );
  XNOR U2645 ( .A(n2249), .B(n2248), .Z(n2250) );
  XOR U2646 ( .A(n2251), .B(n2250), .Z(n2176) );
  NANDN U2647 ( .A(n2140), .B(n2139), .Z(n2144) );
  NAND U2648 ( .A(n2142), .B(n2141), .Z(n2143) );
  AND U2649 ( .A(n2144), .B(n2143), .Z(n2177) );
  XOR U2650 ( .A(n2176), .B(n2177), .Z(n2179) );
  XOR U2651 ( .A(n2178), .B(n2179), .Z(n2146) );
  XOR U2652 ( .A(n2147), .B(n2146), .Z(n2149) );
  XOR U2653 ( .A(n2148), .B(n2149), .Z(n2272) );
  XNOR U2654 ( .A(n2273), .B(n2272), .Z(n2145) );
  XNOR U2655 ( .A(n2274), .B(n2145), .Z(o[3]) );
  NAND U2656 ( .A(n2147), .B(n2146), .Z(n2151) );
  NAND U2657 ( .A(n2149), .B(n2148), .Z(n2150) );
  AND U2658 ( .A(n2151), .B(n2150), .Z(n2285) );
  NANDN U2659 ( .A(n2153), .B(n2152), .Z(n2157) );
  NAND U2660 ( .A(n2155), .B(n2154), .Z(n2156) );
  AND U2661 ( .A(n2157), .B(n2156), .Z(n2318) );
  NANDN U2662 ( .A(n2159), .B(n2158), .Z(n2163) );
  NANDN U2663 ( .A(n2161), .B(n2160), .Z(n2162) );
  AND U2664 ( .A(n2163), .B(n2162), .Z(n2306) );
  NANDN U2665 ( .A(n2165), .B(n2164), .Z(n2169) );
  NAND U2666 ( .A(n2167), .B(n2166), .Z(n2168) );
  AND U2667 ( .A(n2169), .B(n2168), .Z(n2303) );
  NANDN U2668 ( .A(n2171), .B(n2170), .Z(n2175) );
  NANDN U2669 ( .A(n2173), .B(n2172), .Z(n2174) );
  NAND U2670 ( .A(n2175), .B(n2174), .Z(n2304) );
  XNOR U2671 ( .A(n2303), .B(n2304), .Z(n2305) );
  XOR U2672 ( .A(n2306), .B(n2305), .Z(n2316) );
  NAND U2673 ( .A(n2177), .B(n2176), .Z(n2181) );
  NAND U2674 ( .A(n2179), .B(n2178), .Z(n2180) );
  AND U2675 ( .A(n2181), .B(n2180), .Z(n2315) );
  XNOR U2676 ( .A(n2316), .B(n2315), .Z(n2317) );
  XNOR U2677 ( .A(n2318), .B(n2317), .Z(n2282) );
  NANDN U2678 ( .A(n2183), .B(n2182), .Z(n2187) );
  NANDN U2679 ( .A(n2185), .B(n2184), .Z(n2186) );
  AND U2680 ( .A(n2187), .B(n2186), .Z(n2324) );
  NANDN U2681 ( .A(n2189), .B(n2188), .Z(n2193) );
  NANDN U2682 ( .A(n2191), .B(n2190), .Z(n2192) );
  AND U2683 ( .A(n2193), .B(n2192), .Z(n2322) );
  NANDN U2684 ( .A(n2195), .B(n2194), .Z(n2199) );
  NANDN U2685 ( .A(n2197), .B(n2196), .Z(n2198) );
  AND U2686 ( .A(n2199), .B(n2198), .Z(n2343) );
  NANDN U2687 ( .A(n2201), .B(n2200), .Z(n2205) );
  NANDN U2688 ( .A(n2203), .B(n2202), .Z(n2204) );
  AND U2689 ( .A(n2205), .B(n2204), .Z(n2341) );
  XOR U2690 ( .A(n2335), .B(n2334), .Z(n2336) );
  XOR U2691 ( .A(n2333), .B(oglobal[4]), .Z(n2337) );
  XNOR U2692 ( .A(n2336), .B(n2337), .Z(n2340) );
  XNOR U2693 ( .A(n2341), .B(n2340), .Z(n2342) );
  XNOR U2694 ( .A(n2343), .B(n2342), .Z(n2299) );
  NANDN U2695 ( .A(n2215), .B(n2214), .Z(n2219) );
  NANDN U2696 ( .A(n2217), .B(n2216), .Z(n2218) );
  NAND U2697 ( .A(n2219), .B(n2218), .Z(n2297) );
  XNOR U2698 ( .A(n2297), .B(n2298), .Z(n2300) );
  XNOR U2699 ( .A(n2322), .B(n2321), .Z(n2323) );
  XNOR U2700 ( .A(n2324), .B(n2323), .Z(n2312) );
  NANDN U2701 ( .A(n2225), .B(n2224), .Z(n2229) );
  NANDN U2702 ( .A(n2227), .B(n2226), .Z(n2228) );
  AND U2703 ( .A(n2229), .B(n2228), .Z(n2327) );
  NANDN U2704 ( .A(n2231), .B(n2230), .Z(n2235) );
  NANDN U2705 ( .A(n2233), .B(n2232), .Z(n2234) );
  NAND U2706 ( .A(n2235), .B(n2234), .Z(n2328) );
  XNOR U2707 ( .A(n2327), .B(n2328), .Z(n2330) );
  NANDN U2708 ( .A(n2237), .B(n2236), .Z(n2241) );
  OR U2709 ( .A(n2239), .B(n2238), .Z(n2240) );
  AND U2710 ( .A(n2241), .B(n2240), .Z(n2329) );
  XOR U2711 ( .A(n2330), .B(n2329), .Z(n2310) );
  NANDN U2712 ( .A(n2243), .B(n2242), .Z(n2247) );
  NAND U2713 ( .A(n2245), .B(n2244), .Z(n2246) );
  AND U2714 ( .A(n2247), .B(n2246), .Z(n2309) );
  XNOR U2715 ( .A(n2310), .B(n2309), .Z(n2311) );
  XOR U2716 ( .A(n2312), .B(n2311), .Z(n2349) );
  NANDN U2717 ( .A(n2249), .B(n2248), .Z(n2253) );
  NANDN U2718 ( .A(n2251), .B(n2250), .Z(n2252) );
  AND U2719 ( .A(n2253), .B(n2252), .Z(n2346) );
  NANDN U2720 ( .A(n2255), .B(n2254), .Z(n2259) );
  NANDN U2721 ( .A(n2257), .B(n2256), .Z(n2258) );
  NAND U2722 ( .A(n2259), .B(n2258), .Z(n2347) );
  XNOR U2723 ( .A(n2346), .B(n2347), .Z(n2348) );
  XOR U2724 ( .A(n2349), .B(n2348), .Z(n2294) );
  NAND U2725 ( .A(n2261), .B(n2260), .Z(n2265) );
  NANDN U2726 ( .A(n2263), .B(n2262), .Z(n2264) );
  AND U2727 ( .A(n2265), .B(n2264), .Z(n2292) );
  NAND U2728 ( .A(n2267), .B(n2266), .Z(n2271) );
  NAND U2729 ( .A(n2269), .B(n2268), .Z(n2270) );
  AND U2730 ( .A(n2271), .B(n2270), .Z(n2291) );
  XOR U2731 ( .A(n2292), .B(n2291), .Z(n2293) );
  XNOR U2732 ( .A(n2282), .B(n2283), .Z(n2284) );
  XNOR U2733 ( .A(n2285), .B(n2284), .Z(n2290) );
  NANDN U2734 ( .A(n2276), .B(n2275), .Z(n2280) );
  NAND U2735 ( .A(n2278), .B(n2277), .Z(n2279) );
  NAND U2736 ( .A(n2280), .B(n2279), .Z(n2289) );
  XNOR U2737 ( .A(n2288), .B(n2289), .Z(n2281) );
  XNOR U2738 ( .A(n2290), .B(n2281), .Z(o[4]) );
  NANDN U2739 ( .A(n2283), .B(n2282), .Z(n2287) );
  NAND U2740 ( .A(n2285), .B(n2284), .Z(n2286) );
  AND U2741 ( .A(n2287), .B(n2286), .Z(n2362) );
  NAND U2742 ( .A(n2292), .B(n2291), .Z(n2296) );
  NAND U2743 ( .A(n2294), .B(n2293), .Z(n2295) );
  NAND U2744 ( .A(n2296), .B(n2295), .Z(n2354) );
  NANDN U2745 ( .A(n2298), .B(n2297), .Z(n2302) );
  NAND U2746 ( .A(n2300), .B(n2299), .Z(n2301) );
  AND U2747 ( .A(n2302), .B(n2301), .Z(n2375) );
  NANDN U2748 ( .A(n2304), .B(n2303), .Z(n2308) );
  NAND U2749 ( .A(n2306), .B(n2305), .Z(n2307) );
  AND U2750 ( .A(n2308), .B(n2307), .Z(n2373) );
  NANDN U2751 ( .A(n2310), .B(n2309), .Z(n2314) );
  NAND U2752 ( .A(n2312), .B(n2311), .Z(n2313) );
  AND U2753 ( .A(n2314), .B(n2313), .Z(n2372) );
  XNOR U2754 ( .A(n2373), .B(n2372), .Z(n2374) );
  XNOR U2755 ( .A(n2375), .B(n2374), .Z(n2353) );
  XOR U2756 ( .A(n2354), .B(n2353), .Z(n2356) );
  NANDN U2757 ( .A(n2316), .B(n2315), .Z(n2320) );
  NANDN U2758 ( .A(n2318), .B(n2317), .Z(n2319) );
  AND U2759 ( .A(n2320), .B(n2319), .Z(n2369) );
  NANDN U2760 ( .A(n2322), .B(n2321), .Z(n2326) );
  NANDN U2761 ( .A(n2324), .B(n2323), .Z(n2325) );
  AND U2762 ( .A(n2326), .B(n2325), .Z(n2381) );
  NANDN U2763 ( .A(n2328), .B(n2327), .Z(n2332) );
  NAND U2764 ( .A(n2330), .B(n2329), .Z(n2331) );
  AND U2765 ( .A(n2332), .B(n2331), .Z(n2379) );
  ANDN U2766 ( .B(oglobal[4]), .A(n2333), .Z(n2384) );
  XOR U2767 ( .A(n2384), .B(oglobal[5]), .Z(n2386) );
  OR U2768 ( .A(n2335), .B(n2334), .Z(n2339) );
  NANDN U2769 ( .A(n2337), .B(n2336), .Z(n2338) );
  AND U2770 ( .A(n2339), .B(n2338), .Z(n2385) );
  XNOR U2771 ( .A(n2386), .B(n2385), .Z(n2387) );
  NANDN U2772 ( .A(n2341), .B(n2340), .Z(n2345) );
  NANDN U2773 ( .A(n2343), .B(n2342), .Z(n2344) );
  NAND U2774 ( .A(n2345), .B(n2344), .Z(n2388) );
  XNOR U2775 ( .A(n2387), .B(n2388), .Z(n2378) );
  XNOR U2776 ( .A(n2379), .B(n2378), .Z(n2380) );
  XOR U2777 ( .A(n2381), .B(n2380), .Z(n2367) );
  NANDN U2778 ( .A(n2347), .B(n2346), .Z(n2351) );
  NANDN U2779 ( .A(n2349), .B(n2348), .Z(n2350) );
  AND U2780 ( .A(n2351), .B(n2350), .Z(n2366) );
  XNOR U2781 ( .A(n2367), .B(n2366), .Z(n2368) );
  XNOR U2782 ( .A(n2369), .B(n2368), .Z(n2355) );
  XNOR U2783 ( .A(n2356), .B(n2355), .Z(n2360) );
  IV U2784 ( .A(n2360), .Z(n2359) );
  XNOR U2785 ( .A(n2361), .B(n2359), .Z(n2352) );
  XNOR U2786 ( .A(n2362), .B(n2352), .Z(o[5]) );
  NAND U2787 ( .A(n2354), .B(n2353), .Z(n2358) );
  NAND U2788 ( .A(n2356), .B(n2355), .Z(n2357) );
  NAND U2789 ( .A(n2358), .B(n2357), .Z(n2402) );
  NANDN U2790 ( .A(n2361), .B(n2359), .Z(n2365) );
  AND U2791 ( .A(n2361), .B(n2360), .Z(n2363) );
  OR U2792 ( .A(n2363), .B(n2362), .Z(n2364) );
  AND U2793 ( .A(n2365), .B(n2364), .Z(n2400) );
  NANDN U2794 ( .A(n2367), .B(n2366), .Z(n2371) );
  NANDN U2795 ( .A(n2369), .B(n2368), .Z(n2370) );
  AND U2796 ( .A(n2371), .B(n2370), .Z(n2409) );
  NANDN U2797 ( .A(n2373), .B(n2372), .Z(n2377) );
  NAND U2798 ( .A(n2375), .B(n2374), .Z(n2376) );
  AND U2799 ( .A(n2377), .B(n2376), .Z(n2407) );
  NANDN U2800 ( .A(n2379), .B(n2378), .Z(n2383) );
  NAND U2801 ( .A(n2381), .B(n2380), .Z(n2382) );
  AND U2802 ( .A(n2383), .B(n2382), .Z(n2396) );
  AND U2803 ( .A(n2384), .B(oglobal[5]), .Z(n2392) );
  XOR U2804 ( .A(n2392), .B(oglobal[6]), .Z(n2394) );
  NANDN U2805 ( .A(n2386), .B(n2385), .Z(n2390) );
  NANDN U2806 ( .A(n2388), .B(n2387), .Z(n2389) );
  NAND U2807 ( .A(n2390), .B(n2389), .Z(n2393) );
  XNOR U2808 ( .A(n2394), .B(n2393), .Z(n2395) );
  XNOR U2809 ( .A(n2396), .B(n2395), .Z(n2406) );
  XNOR U2810 ( .A(n2407), .B(n2406), .Z(n2408) );
  XNOR U2811 ( .A(n2409), .B(n2408), .Z(n2401) );
  IV U2812 ( .A(n2401), .Z(n2399) );
  XNOR U2813 ( .A(n2400), .B(n2399), .Z(n2391) );
  XNOR U2814 ( .A(n2402), .B(n2391), .Z(o[6]) );
  NAND U2815 ( .A(n2392), .B(oglobal[6]), .Z(n2416) );
  XNOR U2816 ( .A(oglobal[7]), .B(n2416), .Z(n2418) );
  NANDN U2817 ( .A(n2394), .B(n2393), .Z(n2398) );
  NANDN U2818 ( .A(n2396), .B(n2395), .Z(n2397) );
  AND U2819 ( .A(n2398), .B(n2397), .Z(n2417) );
  XNOR U2820 ( .A(n2418), .B(n2417), .Z(n2415) );
  NAND U2821 ( .A(n2399), .B(n2400), .Z(n2405) );
  ANDN U2822 ( .B(n2401), .A(n2400), .Z(n2403) );
  OR U2823 ( .A(n2403), .B(n2402), .Z(n2404) );
  AND U2824 ( .A(n2405), .B(n2404), .Z(n2413) );
  NANDN U2825 ( .A(n2407), .B(n2406), .Z(n2411) );
  NAND U2826 ( .A(n2409), .B(n2408), .Z(n2410) );
  NAND U2827 ( .A(n2411), .B(n2410), .Z(n2414) );
  XNOR U2828 ( .A(n2413), .B(n2414), .Z(n2412) );
  XNOR U2829 ( .A(n2415), .B(n2412), .Z(o[7]) );
  NANDN U2830 ( .A(n2416), .B(oglobal[7]), .Z(n2420) );
  NAND U2831 ( .A(n2418), .B(n2417), .Z(n2419) );
  AND U2832 ( .A(n2420), .B(n2419), .Z(n2421) );
  XNOR U2833 ( .A(n2421), .B(oglobal[8]), .Z(n2422) );
  XNOR U2834 ( .A(n2423), .B(n2422), .Z(o[8]) );
  NANDN U2835 ( .A(n2421), .B(oglobal[8]), .Z(n2425) );
  NANDN U2836 ( .A(n2423), .B(n2422), .Z(n2424) );
  AND U2837 ( .A(n2425), .B(n2424), .Z(n2426) );
  XNOR U2838 ( .A(n2426), .B(oglobal[9]), .Z(o[9]) );
  NANDN U2839 ( .A(n2426), .B(oglobal[9]), .Z(n2427) );
  XNOR U2840 ( .A(oglobal[10]), .B(n2427), .Z(o[10]) );
endmodule

