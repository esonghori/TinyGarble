
module matrixMult_N_M_3_N8_M32 ( clk, rst, x, y, o );
  input [31:0] x;
  input [31:0] y;
  output [31:0] o;
  input clk, rst;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350,
         n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361,
         n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006;

  DFF \o_reg[31]  ( .D(N64), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \o_reg[30]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \o_reg[29]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \o_reg[28]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \o_reg[27]  ( .D(N60), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \o_reg[26]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \o_reg[25]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \o_reg[24]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \o_reg[23]  ( .D(N56), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \o_reg[22]  ( .D(N55), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \o_reg[21]  ( .D(N54), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \o_reg[20]  ( .D(N53), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \o_reg[19]  ( .D(N52), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \o_reg[18]  ( .D(N51), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \o_reg[17]  ( .D(N50), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \o_reg[16]  ( .D(N49), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \o_reg[15]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \o_reg[14]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \o_reg[13]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \o_reg[12]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \o_reg[11]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \o_reg[10]  ( .D(N43), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \o_reg[9]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \o_reg[8]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \o_reg[7]  ( .D(N40), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \o_reg[6]  ( .D(N39), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \o_reg[5]  ( .D(N38), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \o_reg[4]  ( .D(N37), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \o_reg[3]  ( .D(N36), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \o_reg[2]  ( .D(N35), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \o_reg[1]  ( .D(N34), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \o_reg[0]  ( .D(N33), .CLK(clk), .RST(rst), .Q(o[0]) );
  XNOR U3 ( .A(n642), .B(n643), .Z(n645) );
  XOR U4 ( .A(n914), .B(n915), .Z(n946) );
  XOR U5 ( .A(n1473), .B(n1474), .Z(n1475) );
  AND U6 ( .A(y[11]), .B(x[14]), .Z(n1964) );
  XNOR U7 ( .A(n542), .B(n543), .Z(n532) );
  XNOR U8 ( .A(n653), .B(n654), .Z(n610) );
  XOR U9 ( .A(n645), .B(n644), .Z(n604) );
  XOR U10 ( .A(n1274), .B(n1275), .Z(n1300) );
  OR U11 ( .A(n1171), .B(n214), .Z(n1) );
  OR U12 ( .A(n212), .B(n213), .Z(n2) );
  NAND U13 ( .A(n1), .B(n2), .Z(n277) );
  XNOR U14 ( .A(n392), .B(n393), .Z(n375) );
  XOR U15 ( .A(n1263), .B(n1262), .Z(n1306) );
  XOR U16 ( .A(n1695), .B(n1696), .Z(n1595) );
  XNOR U17 ( .A(n1886), .B(n1887), .Z(n1888) );
  NAND U18 ( .A(n1163), .B(n372), .Z(n3) );
  XOR U19 ( .A(n372), .B(n1163), .Z(n4) );
  NANDN U20 ( .A(n373), .B(n4), .Z(n5) );
  NAND U21 ( .A(n3), .B(n5), .Z(n444) );
  XOR U22 ( .A(n2364), .B(n2363), .Z(n2365) );
  XNOR U23 ( .A(n2595), .B(n2596), .Z(n2550) );
  XOR U24 ( .A(n2395), .B(n2396), .Z(n2514) );
  XNOR U25 ( .A(n1747), .B(n1748), .Z(n1749) );
  XNOR U26 ( .A(n755), .B(n756), .Z(n757) );
  XOR U27 ( .A(n788), .B(n789), .Z(n791) );
  XNOR U28 ( .A(n952), .B(n953), .Z(n955) );
  XNOR U29 ( .A(n929), .B(n930), .Z(n896) );
  XNOR U30 ( .A(n1001), .B(n1002), .Z(n988) );
  XNOR U31 ( .A(n1185), .B(n1186), .Z(n1187) );
  XNOR U32 ( .A(n1354), .B(n1355), .Z(n1356) );
  XNOR U33 ( .A(n1772), .B(n1773), .Z(n1774) );
  XOR U34 ( .A(n1766), .B(n1767), .Z(n1769) );
  XOR U35 ( .A(n354), .B(n355), .Z(n356) );
  XOR U36 ( .A(n482), .B(n483), .Z(n477) );
  XOR U37 ( .A(n1228), .B(n1227), .Z(n1229) );
  XNOR U38 ( .A(n1221), .B(n1222), .Z(n1223) );
  ANDN U39 ( .B(x[15]), .A(n2499), .Z(n2086) );
  XOR U40 ( .A(n2303), .B(n2304), .Z(n2291) );
  XOR U41 ( .A(n375), .B(n374), .Z(n376) );
  XOR U42 ( .A(n494), .B(n1180), .Z(n458) );
  XOR U43 ( .A(n686), .B(n687), .Z(n762) );
  XOR U44 ( .A(n1314), .B(n1315), .Z(n1307) );
  XOR U45 ( .A(n1336), .B(n1337), .Z(n1339) );
  XNOR U46 ( .A(n1603), .B(n1604), .Z(n1613) );
  XOR U47 ( .A(n1665), .B(n1666), .Z(n1598) );
  XNOR U48 ( .A(n1778), .B(n1779), .Z(n1780) );
  XNOR U49 ( .A(n2012), .B(n2013), .Z(n2014) );
  XOR U50 ( .A(n2168), .B(n2169), .Z(n2117) );
  AND U51 ( .A(y[4]), .B(x[24]), .Z(n2471) );
  XNOR U52 ( .A(n90), .B(n91), .Z(n76) );
  XOR U53 ( .A(n606), .B(n607), .Z(n598) );
  XNOR U54 ( .A(n2436), .B(n2437), .Z(n2364) );
  XOR U55 ( .A(n2383), .B(n2384), .Z(n2359) );
  XOR U56 ( .A(n2550), .B(n2549), .Z(n2551) );
  OR U57 ( .A(n2621), .B(n2622), .Z(n6) );
  OR U58 ( .A(n2890), .B(n2620), .Z(n7) );
  AND U59 ( .A(n6), .B(n7), .Z(n2733) );
  XOR U60 ( .A(n2880), .B(n2881), .Z(n2878) );
  XNOR U61 ( .A(n2503), .B(n2504), .Z(n2515) );
  OR U62 ( .A(n2584), .B(n2585), .Z(n8) );
  OR U63 ( .A(n2848), .B(n2583), .Z(n9) );
  AND U64 ( .A(n8), .B(n9), .Z(n2724) );
  XNOR U65 ( .A(n663), .B(n662), .Z(n644) );
  XNOR U66 ( .A(n884), .B(n885), .Z(n886) );
  XNOR U67 ( .A(n1125), .B(n1239), .Z(n1156) );
  XNOR U68 ( .A(n1342), .B(n1343), .Z(n1344) );
  XOR U69 ( .A(n1467), .B(n1468), .Z(n1469) );
  AND U70 ( .A(x[12]), .B(y[13]), .Z(n1946) );
  XNOR U71 ( .A(n1910), .B(n1911), .Z(n1912) );
  XOR U72 ( .A(n337), .B(n338), .Z(n340) );
  XNOR U73 ( .A(n386), .B(n387), .Z(n388) );
  XOR U74 ( .A(n569), .B(n568), .Z(n570) );
  XOR U75 ( .A(n611), .B(n610), .Z(n612) );
  XNOR U76 ( .A(n735), .B(n736), .Z(n737) );
  XOR U77 ( .A(n955), .B(n954), .Z(n872) );
  XOR U78 ( .A(n989), .B(n988), .Z(n990) );
  XOR U79 ( .A(n1046), .B(n1047), .Z(n1049) );
  XOR U80 ( .A(n1188), .B(n1187), .Z(n1100) );
  XOR U81 ( .A(n1366), .B(n1367), .Z(n1368) );
  XNOR U82 ( .A(n1360), .B(n1361), .Z(n1362) );
  XNOR U83 ( .A(n1565), .B(n1566), .Z(n1567) );
  XNOR U84 ( .A(n1693), .B(n1694), .Z(n1695) );
  XOR U85 ( .A(n1485), .B(n1486), .Z(n1487) );
  XOR U86 ( .A(n1768), .B(n1769), .Z(n1796) );
  XNOR U87 ( .A(n1790), .B(n1791), .Z(n1792) );
  XOR U88 ( .A(n2086), .B(n2087), .Z(n2089) );
  XNOR U89 ( .A(n2136), .B(n2137), .Z(n2100) );
  XNOR U90 ( .A(n2112), .B(n2113), .Z(n2068) );
  XOR U91 ( .A(n346), .B(n345), .Z(n312) );
  XNOR U92 ( .A(n366), .B(n367), .Z(n368) );
  XOR U93 ( .A(n478), .B(n479), .Z(n501) );
  XOR U94 ( .A(n532), .B(n531), .Z(n533) );
  XOR U95 ( .A(n470), .B(n471), .Z(n473) );
  XOR U96 ( .A(n527), .B(n528), .Z(n519) );
  XOR U97 ( .A(n802), .B(n803), .Z(n809) );
  XOR U98 ( .A(n984), .B(n985), .Z(n970) );
  XNOR U99 ( .A(n1042), .B(n1043), .Z(n1052) );
  XNOR U100 ( .A(n1260), .B(n1261), .Z(n1263) );
  XOR U101 ( .A(n1445), .B(n1446), .Z(n1438) );
  XNOR U102 ( .A(n1928), .B(n1929), .Z(n1930) );
  XNOR U103 ( .A(n1784), .B(n1785), .Z(n1786) );
  XNOR U104 ( .A(n2006), .B(n2007), .Z(n2008) );
  XOR U105 ( .A(n2267), .B(n2268), .Z(n2274) );
  XNOR U106 ( .A(n2407), .B(n2408), .Z(n2384) );
  XOR U107 ( .A(n2448), .B(n2449), .Z(n2460) );
  AND U108 ( .A(y[16]), .B(x[12]), .Z(n2477) );
  XNOR U109 ( .A(n443), .B(n444), .Z(n445) );
  XOR U110 ( .A(n599), .B(n598), .Z(n600) );
  XNOR U111 ( .A(n1615), .B(n1616), .Z(n1589) );
  XOR U112 ( .A(n2339), .B(n2340), .Z(n2342) );
  XOR U113 ( .A(n2401), .B(n2402), .Z(n2366) );
  XOR U114 ( .A(n2641), .B(n2642), .Z(n2552) );
  XOR U115 ( .A(n2672), .B(n2673), .Z(n2677) );
  AND U116 ( .A(y[13]), .B(x[16]), .Z(n2586) );
  OR U117 ( .A(n2896), .B(n2601), .Z(n10) );
  OR U118 ( .A(n2599), .B(n2600), .Z(n11) );
  NAND U119 ( .A(n10), .B(n11), .Z(n2879) );
  XOR U120 ( .A(n2754), .B(n2755), .Z(n2753) );
  XNOR U121 ( .A(n2763), .B(n2764), .Z(n2744) );
  XNOR U122 ( .A(n2509), .B(n2510), .Z(n2525) );
  NAND U123 ( .A(n89), .B(n59), .Z(n12) );
  XOR U124 ( .A(n59), .B(n89), .Z(n13) );
  NANDN U125 ( .A(n60), .B(n13), .Z(n14) );
  NAND U126 ( .A(n12), .B(n14), .Z(n71) );
  XOR U127 ( .A(n77), .B(n76), .Z(n78) );
  XOR U128 ( .A(n278), .B(n279), .Z(n256) );
  XNOR U129 ( .A(n678), .B(n679), .Z(n680) );
  XNOR U130 ( .A(n1209), .B(n1210), .Z(n1211) );
  XNOR U131 ( .A(n1455), .B(n1456), .Z(n1457) );
  XOR U132 ( .A(n1864), .B(n1865), .Z(n1732) );
  XNOR U133 ( .A(n2024), .B(n2025), .Z(n2026) );
  OR U134 ( .A(n2658), .B(n2659), .Z(n15) );
  OR U135 ( .A(n2760), .B(n2657), .Z(n16) );
  NAND U136 ( .A(n15), .B(n16), .Z(n2931) );
  XNOR U137 ( .A(n2696), .B(n2697), .Z(n2703) );
  XOR U138 ( .A(n134), .B(n135), .Z(n129) );
  XOR U139 ( .A(n2186), .B(n2187), .Z(n2181) );
  XNOR U140 ( .A(n2997), .B(n2998), .Z(n2993) );
  IV U141 ( .A(y[0]), .Z(n17) );
  IV U142 ( .A(y[1]), .Z(n18) );
  IV U143 ( .A(y[2]), .Z(n19) );
  IV U144 ( .A(y[3]), .Z(n20) );
  IV U145 ( .A(y[4]), .Z(n21) );
  IV U146 ( .A(y[5]), .Z(n22) );
  IV U147 ( .A(y[6]), .Z(n23) );
  IV U148 ( .A(x[0]), .Z(n24) );
  IV U149 ( .A(x[1]), .Z(n25) );
  IV U150 ( .A(x[2]), .Z(n26) );
  IV U151 ( .A(x[3]), .Z(n27) );
  IV U152 ( .A(x[7]), .Z(n28) );
  IV U153 ( .A(x[8]), .Z(n29) );
  AND U154 ( .A(y[0]), .B(x[0]), .Z(n707) );
  XOR U155 ( .A(n707), .B(o[0]), .Z(N33) );
  AND U156 ( .A(y[0]), .B(x[1]), .Z(n30) );
  NAND U157 ( .A(y[1]), .B(x[0]), .Z(n36) );
  XNOR U158 ( .A(n36), .B(o[1]), .Z(n31) );
  XOR U159 ( .A(n30), .B(n31), .Z(n32) );
  AND U160 ( .A(o[0]), .B(n707), .Z(n33) );
  XOR U161 ( .A(n32), .B(n33), .Z(N34) );
  OR U162 ( .A(n31), .B(n30), .Z(n35) );
  NANDN U163 ( .A(n33), .B(n32), .Z(n34) );
  NAND U164 ( .A(n35), .B(n34), .Z(n38) );
  NAND U165 ( .A(y[2]), .B(x[0]), .Z(n49) );
  XOR U166 ( .A(n49), .B(o[2]), .Z(n37) );
  XNOR U167 ( .A(n38), .B(n37), .Z(n40) );
  ANDN U168 ( .B(o[1]), .A(n36), .Z(n43) );
  ANDN U169 ( .B(x[2]), .A(n17), .Z(n44) );
  XNOR U170 ( .A(n43), .B(n44), .Z(n46) );
  ANDN U171 ( .B(x[1]), .A(n18), .Z(n45) );
  XNOR U172 ( .A(n46), .B(n45), .Z(n39) );
  XNOR U173 ( .A(n40), .B(n39), .Z(N35) );
  NAND U174 ( .A(n38), .B(n37), .Z(n42) );
  OR U175 ( .A(n40), .B(n39), .Z(n41) );
  NAND U176 ( .A(n42), .B(n41), .Z(n53) );
  OR U177 ( .A(n44), .B(n43), .Z(n48) );
  OR U178 ( .A(n46), .B(n45), .Z(n47) );
  AND U179 ( .A(n48), .B(n47), .Z(n54) );
  XNOR U180 ( .A(n53), .B(n54), .Z(n55) );
  NAND U181 ( .A(y[1]), .B(x[2]), .Z(n65) );
  XNOR U182 ( .A(n65), .B(o[3]), .Z(n59) );
  NANDN U183 ( .A(n49), .B(o[2]), .Z(n62) );
  AND U184 ( .A(x[0]), .B(y[3]), .Z(n51) );
  NAND U185 ( .A(x[3]), .B(y[0]), .Z(n50) );
  XOR U186 ( .A(n51), .B(n50), .Z(n61) );
  XNOR U187 ( .A(n62), .B(n61), .Z(n60) );
  ANDN U188 ( .B(x[1]), .A(n19), .Z(n89) );
  XOR U189 ( .A(n60), .B(n89), .Z(n52) );
  XOR U190 ( .A(n59), .B(n52), .Z(n56) );
  XNOR U191 ( .A(n55), .B(n56), .Z(N36) );
  NANDN U192 ( .A(n54), .B(n53), .Z(n58) );
  NAND U193 ( .A(n56), .B(n55), .Z(n57) );
  NAND U194 ( .A(n58), .B(n57), .Z(n70) );
  XNOR U195 ( .A(n70), .B(n71), .Z(n72) );
  ANDN U196 ( .B(y[3]), .A(n27), .Z(n138) );
  NAND U197 ( .A(n707), .B(n138), .Z(n64) );
  OR U198 ( .A(n62), .B(n61), .Z(n63) );
  NAND U199 ( .A(n64), .B(n63), .Z(n79) );
  NANDN U200 ( .A(n65), .B(o[3]), .Z(n86) );
  AND U201 ( .A(x[0]), .B(y[4]), .Z(n67) );
  AND U202 ( .A(y[0]), .B(x[4]), .Z(n66) );
  XNOR U203 ( .A(n67), .B(n66), .Z(n85) );
  XOR U204 ( .A(n86), .B(n85), .Z(n77) );
  AND U205 ( .A(y[3]), .B(x[1]), .Z(n69) );
  NAND U206 ( .A(y[2]), .B(x[2]), .Z(n68) );
  XOR U207 ( .A(n69), .B(n68), .Z(n91) );
  NAND U208 ( .A(x[3]), .B(y[1]), .Z(n82) );
  XNOR U209 ( .A(n82), .B(o[4]), .Z(n90) );
  XOR U210 ( .A(n79), .B(n78), .Z(n73) );
  XOR U211 ( .A(n72), .B(n73), .Z(N37) );
  NANDN U212 ( .A(n71), .B(n70), .Z(n75) );
  NANDN U213 ( .A(n73), .B(n72), .Z(n74) );
  NAND U214 ( .A(n75), .B(n74), .Z(n94) );
  NAND U215 ( .A(n77), .B(n76), .Z(n81) );
  NAND U216 ( .A(n79), .B(n78), .Z(n80) );
  NAND U217 ( .A(n81), .B(n80), .Z(n95) );
  XNOR U218 ( .A(n94), .B(n95), .Z(n96) );
  NANDN U219 ( .A(n82), .B(o[4]), .Z(n114) );
  AND U220 ( .A(y[5]), .B(x[0]), .Z(n84) );
  AND U221 ( .A(x[5]), .B(y[0]), .Z(n83) );
  XNOR U222 ( .A(n84), .B(n83), .Z(n113) );
  XOR U223 ( .A(n114), .B(n113), .Z(n108) );
  ANDN U224 ( .B(y[3]), .A(n26), .Z(n106) );
  ANDN U225 ( .B(x[1]), .A(n21), .Z(n122) );
  ANDN U226 ( .B(x[4]), .A(n18), .Z(n117) );
  XOR U227 ( .A(o[5]), .B(n117), .Z(n120) );
  ANDN U228 ( .B(x[3]), .A(n19), .Z(n121) );
  XNOR U229 ( .A(n120), .B(n121), .Z(n123) );
  XNOR U230 ( .A(n122), .B(n123), .Z(n107) );
  XNOR U231 ( .A(n106), .B(n107), .Z(n109) );
  XNOR U232 ( .A(n108), .B(n109), .Z(n103) );
  IV U233 ( .A(x[4]), .Z(n2454) );
  ANDN U234 ( .B(y[4]), .A(n2454), .Z(n212) );
  NAND U235 ( .A(n707), .B(n212), .Z(n88) );
  OR U236 ( .A(n86), .B(n85), .Z(n87) );
  NAND U237 ( .A(n88), .B(n87), .Z(n101) );
  NAND U238 ( .A(n89), .B(n106), .Z(n93) );
  NANDN U239 ( .A(n91), .B(n90), .Z(n92) );
  NAND U240 ( .A(n93), .B(n92), .Z(n100) );
  XNOR U241 ( .A(n101), .B(n100), .Z(n102) );
  XNOR U242 ( .A(n103), .B(n102), .Z(n97) );
  XOR U243 ( .A(n96), .B(n97), .Z(N38) );
  NANDN U244 ( .A(n95), .B(n94), .Z(n99) );
  NANDN U245 ( .A(n97), .B(n96), .Z(n98) );
  NAND U246 ( .A(n99), .B(n98), .Z(n126) );
  OR U247 ( .A(n101), .B(n100), .Z(n105) );
  OR U248 ( .A(n103), .B(n102), .Z(n104) );
  AND U249 ( .A(n105), .B(n104), .Z(n127) );
  XNOR U250 ( .A(n126), .B(n127), .Z(n128) );
  OR U251 ( .A(n107), .B(n106), .Z(n111) );
  OR U252 ( .A(n109), .B(n108), .Z(n110) );
  AND U253 ( .A(n111), .B(n110), .Z(n132) );
  AND U254 ( .A(y[5]), .B(x[5]), .Z(n112) );
  NAND U255 ( .A(n707), .B(n112), .Z(n116) );
  OR U256 ( .A(n114), .B(n113), .Z(n115) );
  NAND U257 ( .A(n116), .B(n115), .Z(n154) );
  NAND U258 ( .A(n117), .B(o[5]), .Z(n145) );
  AND U259 ( .A(x[0]), .B(y[6]), .Z(n119) );
  AND U260 ( .A(x[6]), .B(y[0]), .Z(n118) );
  XNOR U261 ( .A(n119), .B(n118), .Z(n144) );
  XOR U262 ( .A(n145), .B(n144), .Z(n153) );
  XNOR U263 ( .A(n154), .B(n153), .Z(n156) );
  ANDN U264 ( .B(x[4]), .A(n19), .Z(n492) );
  ANDN U265 ( .B(x[1]), .A(n22), .Z(n413) );
  AND U266 ( .A(x[5]), .B(y[1]), .Z(n148) );
  XNOR U267 ( .A(o[6]), .B(n148), .Z(n149) );
  XOR U268 ( .A(n413), .B(n149), .Z(n150) );
  XOR U269 ( .A(n492), .B(n150), .Z(n139) );
  AND U270 ( .A(x[2]), .B(y[4]), .Z(n559) );
  XNOR U271 ( .A(n138), .B(n559), .Z(n140) );
  XOR U272 ( .A(n139), .B(n140), .Z(n155) );
  XNOR U273 ( .A(n156), .B(n155), .Z(n133) );
  XOR U274 ( .A(n132), .B(n133), .Z(n134) );
  OR U275 ( .A(n121), .B(n120), .Z(n125) );
  OR U276 ( .A(n123), .B(n122), .Z(n124) );
  AND U277 ( .A(n125), .B(n124), .Z(n135) );
  XOR U278 ( .A(n128), .B(n129), .Z(N39) );
  NANDN U279 ( .A(n127), .B(n126), .Z(n131) );
  NANDN U280 ( .A(n129), .B(n128), .Z(n130) );
  NAND U281 ( .A(n131), .B(n130), .Z(n188) );
  OR U282 ( .A(n133), .B(n132), .Z(n137) );
  NANDN U283 ( .A(n135), .B(n134), .Z(n136) );
  AND U284 ( .A(n137), .B(n136), .Z(n189) );
  XNOR U285 ( .A(n188), .B(n189), .Z(n190) );
  OR U286 ( .A(n138), .B(n559), .Z(n142) );
  NANDN U287 ( .A(n140), .B(n139), .Z(n141) );
  NAND U288 ( .A(n142), .B(n141), .Z(n185) );
  AND U289 ( .A(y[6]), .B(x[6]), .Z(n143) );
  NAND U290 ( .A(n707), .B(n143), .Z(n147) );
  OR U291 ( .A(n145), .B(n144), .Z(n146) );
  AND U292 ( .A(n147), .B(n146), .Z(n183) );
  IV U293 ( .A(x[5]), .Z(n2252) );
  ANDN U294 ( .B(y[2]), .A(n2252), .Z(n332) );
  ANDN U295 ( .B(x[1]), .A(n23), .Z(n541) );
  NAND U296 ( .A(x[6]), .B(y[1]), .Z(n171) );
  XNOR U297 ( .A(o[7]), .B(n171), .Z(n172) );
  XNOR U298 ( .A(n541), .B(n172), .Z(n173) );
  XNOR U299 ( .A(n332), .B(n173), .Z(n182) );
  XOR U300 ( .A(n183), .B(n182), .Z(n184) );
  XNOR U301 ( .A(n185), .B(n184), .Z(n194) );
  ANDN U302 ( .B(x[2]), .A(n22), .Z(n616) );
  ANDN U303 ( .B(y[3]), .A(n2454), .Z(n360) );
  ANDN U304 ( .B(y[4]), .A(n27), .Z(n167) );
  XNOR U305 ( .A(n360), .B(n167), .Z(n168) );
  XOR U306 ( .A(n616), .B(n168), .Z(n176) );
  NAND U307 ( .A(x[0]), .B(y[7]), .Z(n164) );
  AND U308 ( .A(n148), .B(o[6]), .Z(n162) );
  NAND U309 ( .A(x[7]), .B(y[0]), .Z(n161) );
  XNOR U310 ( .A(n162), .B(n161), .Z(n163) );
  XOR U311 ( .A(n164), .B(n163), .Z(n177) );
  XNOR U312 ( .A(n176), .B(n177), .Z(n179) );
  NANDN U313 ( .A(n149), .B(n413), .Z(n152) );
  NANDN U314 ( .A(n150), .B(n492), .Z(n151) );
  AND U315 ( .A(n152), .B(n151), .Z(n178) );
  XOR U316 ( .A(n179), .B(n178), .Z(n195) );
  XOR U317 ( .A(n194), .B(n195), .Z(n197) );
  OR U318 ( .A(n154), .B(n153), .Z(n158) );
  OR U319 ( .A(n156), .B(n155), .Z(n157) );
  AND U320 ( .A(n158), .B(n157), .Z(n196) );
  XOR U321 ( .A(n197), .B(n196), .Z(n191) );
  XNOR U322 ( .A(n190), .B(n191), .Z(N40) );
  AND U323 ( .A(y[0]), .B(x[8]), .Z(n160) );
  NAND U324 ( .A(y[8]), .B(x[0]), .Z(n159) );
  XOR U325 ( .A(n160), .B(n159), .Z(n222) );
  NAND U326 ( .A(y[1]), .B(x[7]), .Z(n225) );
  XNOR U327 ( .A(n225), .B(o[8]), .Z(n221) );
  XOR U328 ( .A(n222), .B(n221), .Z(n243) );
  NANDN U329 ( .A(n162), .B(n161), .Z(n166) );
  NAND U330 ( .A(n164), .B(n163), .Z(n165) );
  NAND U331 ( .A(n166), .B(n165), .Z(n242) );
  XOR U332 ( .A(n243), .B(n242), .Z(n244) );
  OR U333 ( .A(n167), .B(n360), .Z(n170) );
  OR U334 ( .A(n168), .B(n616), .Z(n169) );
  NAND U335 ( .A(n170), .B(n169), .Z(n245) );
  XNOR U336 ( .A(n244), .B(n245), .Z(n208) );
  ANDN U337 ( .B(x[6]), .A(n19), .Z(n213) );
  XNOR U338 ( .A(n212), .B(n213), .Z(n214) );
  NOR U339 ( .A(n26), .B(n23), .Z(n1171) );
  XNOR U340 ( .A(n214), .B(n1171), .Z(n215) );
  ANDN U341 ( .B(x[3]), .A(n22), .Z(n1020) );
  XNOR U342 ( .A(n215), .B(n1020), .Z(n217) );
  NANDN U343 ( .A(n171), .B(o[7]), .Z(n233) );
  AND U344 ( .A(y[7]), .B(x[1]), .Z(n712) );
  AND U345 ( .A(x[5]), .B(y[3]), .Z(n847) );
  XNOR U346 ( .A(n712), .B(n847), .Z(n232) );
  XOR U347 ( .A(n233), .B(n232), .Z(n216) );
  XNOR U348 ( .A(n217), .B(n216), .Z(n236) );
  NAND U349 ( .A(n541), .B(n172), .Z(n175) );
  NANDN U350 ( .A(n173), .B(n332), .Z(n174) );
  AND U351 ( .A(n175), .B(n174), .Z(n237) );
  XOR U352 ( .A(n236), .B(n237), .Z(n239) );
  OR U353 ( .A(n177), .B(n176), .Z(n181) );
  OR U354 ( .A(n179), .B(n178), .Z(n180) );
  AND U355 ( .A(n181), .B(n180), .Z(n238) );
  XOR U356 ( .A(n239), .B(n238), .Z(n206) );
  NANDN U357 ( .A(n183), .B(n182), .Z(n187) );
  OR U358 ( .A(n185), .B(n184), .Z(n186) );
  NAND U359 ( .A(n187), .B(n186), .Z(n207) );
  XNOR U360 ( .A(n206), .B(n207), .Z(n209) );
  XNOR U361 ( .A(n208), .B(n209), .Z(n203) );
  NANDN U362 ( .A(n189), .B(n188), .Z(n193) );
  NAND U363 ( .A(n191), .B(n190), .Z(n192) );
  NAND U364 ( .A(n193), .B(n192), .Z(n200) );
  NANDN U365 ( .A(n195), .B(n194), .Z(n199) );
  OR U366 ( .A(n197), .B(n196), .Z(n198) );
  AND U367 ( .A(n199), .B(n198), .Z(n201) );
  XNOR U368 ( .A(n200), .B(n201), .Z(n202) );
  XOR U369 ( .A(n203), .B(n202), .Z(N41) );
  NANDN U370 ( .A(n201), .B(n200), .Z(n205) );
  NANDN U371 ( .A(n203), .B(n202), .Z(n204) );
  NAND U372 ( .A(n205), .B(n204), .Z(n248) );
  OR U373 ( .A(n207), .B(n206), .Z(n211) );
  OR U374 ( .A(n209), .B(n208), .Z(n210) );
  AND U375 ( .A(n211), .B(n210), .Z(n249) );
  XNOR U376 ( .A(n248), .B(n249), .Z(n250) );
  OR U377 ( .A(n215), .B(n1020), .Z(n219) );
  OR U378 ( .A(n217), .B(n216), .Z(n218) );
  NAND U379 ( .A(n219), .B(n218), .Z(n276) );
  XOR U380 ( .A(n277), .B(n276), .Z(n278) );
  AND U381 ( .A(x[8]), .B(y[8]), .Z(n220) );
  NAND U382 ( .A(n707), .B(n220), .Z(n224) );
  NANDN U383 ( .A(n222), .B(n221), .Z(n223) );
  NAND U384 ( .A(n224), .B(n223), .Z(n263) );
  NANDN U385 ( .A(n225), .B(o[8]), .Z(n283) );
  AND U386 ( .A(y[2]), .B(x[7]), .Z(n227) );
  AND U387 ( .A(x[5]), .B(y[4]), .Z(n226) );
  XNOR U388 ( .A(n227), .B(n226), .Z(n282) );
  XOR U389 ( .A(n283), .B(n282), .Z(n261) );
  AND U390 ( .A(x[0]), .B(y[9]), .Z(n229) );
  NAND U391 ( .A(y[0]), .B(x[9]), .Z(n228) );
  XOR U392 ( .A(n229), .B(n228), .Z(n296) );
  NAND U393 ( .A(y[1]), .B(x[8]), .Z(n289) );
  XOR U394 ( .A(n289), .B(o[9]), .Z(n295) );
  XNOR U395 ( .A(n296), .B(n295), .Z(n260) );
  XOR U396 ( .A(n261), .B(n260), .Z(n262) );
  XNOR U397 ( .A(n263), .B(n262), .Z(n272) );
  NAND U398 ( .A(y[5]), .B(x[4]), .Z(n719) );
  AND U399 ( .A(x[6]), .B(y[3]), .Z(n231) );
  NAND U400 ( .A(y[8]), .B(x[1]), .Z(n230) );
  XNOR U401 ( .A(n231), .B(n230), .Z(n291) );
  XNOR U402 ( .A(n719), .B(n291), .Z(n266) );
  IV U403 ( .A(y[7]), .Z(n2433) );
  ANDN U404 ( .B(x[2]), .A(n2433), .Z(n933) );
  NAND U405 ( .A(y[6]), .B(x[3]), .Z(n648) );
  XOR U406 ( .A(n933), .B(n648), .Z(n267) );
  XNOR U407 ( .A(n266), .B(n267), .Z(n270) );
  NAND U408 ( .A(y[3]), .B(x[1]), .Z(n290) );
  ANDN U409 ( .B(y[7]), .A(n2252), .Z(n456) );
  NANDN U410 ( .A(n290), .B(n456), .Z(n235) );
  OR U411 ( .A(n233), .B(n232), .Z(n234) );
  AND U412 ( .A(n235), .B(n234), .Z(n271) );
  XOR U413 ( .A(n270), .B(n271), .Z(n273) );
  XOR U414 ( .A(n272), .B(n273), .Z(n279) );
  NANDN U415 ( .A(n237), .B(n236), .Z(n241) );
  OR U416 ( .A(n239), .B(n238), .Z(n240) );
  NAND U417 ( .A(n241), .B(n240), .Z(n255) );
  OR U418 ( .A(n243), .B(n242), .Z(n247) );
  NANDN U419 ( .A(n245), .B(n244), .Z(n246) );
  NAND U420 ( .A(n247), .B(n246), .Z(n254) );
  XOR U421 ( .A(n255), .B(n254), .Z(n257) );
  XNOR U422 ( .A(n256), .B(n257), .Z(n251) );
  XOR U423 ( .A(n250), .B(n251), .Z(N42) );
  NANDN U424 ( .A(n249), .B(n248), .Z(n253) );
  NANDN U425 ( .A(n251), .B(n250), .Z(n252) );
  NAND U426 ( .A(n253), .B(n252), .Z(n299) );
  OR U427 ( .A(n255), .B(n254), .Z(n259) );
  NAND U428 ( .A(n257), .B(n256), .Z(n258) );
  AND U429 ( .A(n259), .B(n258), .Z(n300) );
  XNOR U430 ( .A(n299), .B(n300), .Z(n301) );
  NANDN U431 ( .A(n261), .B(n260), .Z(n265) );
  OR U432 ( .A(n263), .B(n262), .Z(n264) );
  NAND U433 ( .A(n265), .B(n264), .Z(n318) );
  NANDN U434 ( .A(n933), .B(n648), .Z(n269) );
  OR U435 ( .A(n267), .B(n266), .Z(n268) );
  NAND U436 ( .A(n269), .B(n268), .Z(n317) );
  XOR U437 ( .A(n318), .B(n317), .Z(n319) );
  NANDN U438 ( .A(n271), .B(n270), .Z(n275) );
  NANDN U439 ( .A(n273), .B(n272), .Z(n274) );
  AND U440 ( .A(n275), .B(n274), .Z(n320) );
  XNOR U441 ( .A(n319), .B(n320), .Z(n307) );
  OR U442 ( .A(n277), .B(n276), .Z(n281) );
  NANDN U443 ( .A(n279), .B(n278), .Z(n280) );
  NAND U444 ( .A(n281), .B(n280), .Z(n306) );
  AND U445 ( .A(x[7]), .B(y[4]), .Z(n324) );
  NAND U446 ( .A(n324), .B(n332), .Z(n285) );
  OR U447 ( .A(n283), .B(n282), .Z(n284) );
  AND U448 ( .A(n285), .B(n284), .Z(n339) );
  AND U449 ( .A(y[2]), .B(x[8]), .Z(n546) );
  NAND U450 ( .A(x[5]), .B(y[5]), .Z(n286) );
  XOR U451 ( .A(n546), .B(n286), .Z(n334) );
  NAND U452 ( .A(x[9]), .B(y[1]), .Z(n349) );
  XOR U453 ( .A(o[10]), .B(n349), .Z(n333) );
  XOR U454 ( .A(n334), .B(n333), .Z(n337) );
  AND U455 ( .A(y[3]), .B(x[7]), .Z(n288) );
  NAND U456 ( .A(x[4]), .B(y[6]), .Z(n287) );
  XOR U457 ( .A(n288), .B(n287), .Z(n363) );
  NAND U458 ( .A(x[6]), .B(y[4]), .Z(n362) );
  XNOR U459 ( .A(n363), .B(n362), .Z(n338) );
  XNOR U460 ( .A(n339), .B(n340), .Z(n313) );
  ANDN U461 ( .B(y[10]), .A(n24), .Z(n357) );
  NANDN U462 ( .A(n289), .B(o[9]), .Z(n354) );
  ANDN U463 ( .B(x[10]), .A(n17), .Z(n355) );
  XNOR U464 ( .A(n357), .B(n356), .Z(n345) );
  IV U465 ( .A(y[9]), .Z(n2314) );
  ANDN U466 ( .B(x[1]), .A(n2314), .Z(n1289) );
  ANDN U467 ( .B(x[3]), .A(n2433), .Z(n1250) );
  NANDN U468 ( .A(n26), .B(y[8]), .Z(n328) );
  XNOR U469 ( .A(n1250), .B(n328), .Z(n329) );
  XNOR U470 ( .A(n1289), .B(n329), .Z(n344) );
  IV U471 ( .A(y[8]), .Z(n2430) );
  ANDN U472 ( .B(x[6]), .A(n2430), .Z(n633) );
  NANDN U473 ( .A(n290), .B(n633), .Z(n293) );
  NANDN U474 ( .A(n719), .B(n291), .Z(n292) );
  AND U475 ( .A(n293), .B(n292), .Z(n343) );
  XOR U476 ( .A(n344), .B(n343), .Z(n346) );
  AND U477 ( .A(x[9]), .B(y[9]), .Z(n294) );
  NAND U478 ( .A(n707), .B(n294), .Z(n298) );
  OR U479 ( .A(n296), .B(n295), .Z(n297) );
  NAND U480 ( .A(n298), .B(n297), .Z(n311) );
  XNOR U481 ( .A(n312), .B(n311), .Z(n314) );
  XOR U482 ( .A(n313), .B(n314), .Z(n305) );
  XNOR U483 ( .A(n306), .B(n305), .Z(n308) );
  XNOR U484 ( .A(n307), .B(n308), .Z(n302) );
  XOR U485 ( .A(n301), .B(n302), .Z(N43) );
  NANDN U486 ( .A(n300), .B(n299), .Z(n304) );
  NANDN U487 ( .A(n302), .B(n301), .Z(n303) );
  NAND U488 ( .A(n304), .B(n303), .Z(n419) );
  OR U489 ( .A(n306), .B(n305), .Z(n310) );
  OR U490 ( .A(n308), .B(n307), .Z(n309) );
  AND U491 ( .A(n310), .B(n309), .Z(n420) );
  XNOR U492 ( .A(n419), .B(n420), .Z(n421) );
  OR U493 ( .A(n312), .B(n311), .Z(n316) );
  NANDN U494 ( .A(n314), .B(n313), .Z(n315) );
  AND U495 ( .A(n316), .B(n315), .Z(n425) );
  OR U496 ( .A(n318), .B(n317), .Z(n322) );
  NANDN U497 ( .A(n320), .B(n319), .Z(n321) );
  NAND U498 ( .A(n322), .B(n321), .Z(n426) );
  XOR U499 ( .A(n425), .B(n426), .Z(n428) );
  NAND U500 ( .A(y[2]), .B(x[9]), .Z(n323) );
  XOR U501 ( .A(n324), .B(n323), .Z(n398) );
  NAND U502 ( .A(y[3]), .B(x[8]), .Z(n397) );
  XNOR U503 ( .A(n398), .B(n397), .Z(n373) );
  ANDN U504 ( .B(x[3]), .A(n2430), .Z(n1163) );
  AND U505 ( .A(y[9]), .B(x[2]), .Z(n326) );
  NAND U506 ( .A(x[5]), .B(y[6]), .Z(n325) );
  XOR U507 ( .A(n326), .B(n325), .Z(n410) );
  NAND U508 ( .A(y[7]), .B(x[4]), .Z(n409) );
  XOR U509 ( .A(n410), .B(n409), .Z(n372) );
  XOR U510 ( .A(n1163), .B(n372), .Z(n327) );
  XOR U511 ( .A(n373), .B(n327), .Z(n389) );
  NANDN U512 ( .A(n1250), .B(n328), .Z(n331) );
  NANDN U513 ( .A(n1289), .B(n329), .Z(n330) );
  NAND U514 ( .A(n331), .B(n330), .Z(n386) );
  NAND U515 ( .A(y[5]), .B(x[8]), .Z(n1140) );
  NANDN U516 ( .A(n1140), .B(n332), .Z(n336) );
  OR U517 ( .A(n334), .B(n333), .Z(n335) );
  NAND U518 ( .A(n336), .B(n335), .Z(n387) );
  XOR U519 ( .A(n389), .B(n388), .Z(n380) );
  NANDN U520 ( .A(n338), .B(n337), .Z(n342) );
  OR U521 ( .A(n340), .B(n339), .Z(n341) );
  AND U522 ( .A(n342), .B(n341), .Z(n381) );
  XNOR U523 ( .A(n380), .B(n381), .Z(n383) );
  OR U524 ( .A(n344), .B(n343), .Z(n348) );
  NAND U525 ( .A(n346), .B(n345), .Z(n347) );
  NAND U526 ( .A(n348), .B(n347), .Z(n369) );
  NANDN U527 ( .A(n349), .B(o[10]), .Z(n393) );
  AND U528 ( .A(x[0]), .B(y[11]), .Z(n351) );
  NAND U529 ( .A(y[0]), .B(x[11]), .Z(n350) );
  XNOR U530 ( .A(n351), .B(n350), .Z(n392) );
  AND U531 ( .A(y[10]), .B(x[1]), .Z(n353) );
  NAND U532 ( .A(x[6]), .B(y[5]), .Z(n352) );
  XOR U533 ( .A(n353), .B(n352), .Z(n416) );
  NAND U534 ( .A(x[10]), .B(y[1]), .Z(n401) );
  XOR U535 ( .A(o[11]), .B(n401), .Z(n415) );
  XOR U536 ( .A(n416), .B(n415), .Z(n374) );
  NANDN U537 ( .A(n355), .B(n354), .Z(n359) );
  OR U538 ( .A(n357), .B(n356), .Z(n358) );
  NAND U539 ( .A(n359), .B(n358), .Z(n377) );
  XOR U540 ( .A(n376), .B(n377), .Z(n366) );
  AND U541 ( .A(x[7]), .B(y[6]), .Z(n361) );
  NAND U542 ( .A(n361), .B(n360), .Z(n365) );
  OR U543 ( .A(n363), .B(n362), .Z(n364) );
  NAND U544 ( .A(n365), .B(n364), .Z(n367) );
  XNOR U545 ( .A(n369), .B(n368), .Z(n382) );
  XNOR U546 ( .A(n383), .B(n382), .Z(n427) );
  XNOR U547 ( .A(n428), .B(n427), .Z(n422) );
  XOR U548 ( .A(n421), .B(n422), .Z(N44) );
  NANDN U549 ( .A(n367), .B(n366), .Z(n371) );
  NANDN U550 ( .A(n369), .B(n368), .Z(n370) );
  NAND U551 ( .A(n371), .B(n370), .Z(n446) );
  NAND U552 ( .A(n375), .B(n374), .Z(n379) );
  NANDN U553 ( .A(n377), .B(n376), .Z(n378) );
  AND U554 ( .A(n379), .B(n378), .Z(n443) );
  XNOR U555 ( .A(n446), .B(n445), .Z(n440) );
  OR U556 ( .A(n381), .B(n380), .Z(n385) );
  OR U557 ( .A(n383), .B(n382), .Z(n384) );
  NAND U558 ( .A(n385), .B(n384), .Z(n438) );
  NANDN U559 ( .A(n387), .B(n386), .Z(n391) );
  NAND U560 ( .A(n389), .B(n388), .Z(n390) );
  NAND U561 ( .A(n391), .B(n390), .Z(n503) );
  IV U562 ( .A(y[11]), .Z(n2499) );
  ANDN U563 ( .B(x[11]), .A(n2499), .Z(n1492) );
  NAND U564 ( .A(n707), .B(n1492), .Z(n395) );
  NANDN U565 ( .A(n393), .B(n392), .Z(n394) );
  NAND U566 ( .A(n395), .B(n394), .Z(n478) );
  NAND U567 ( .A(y[2]), .B(x[7]), .Z(n620) );
  AND U568 ( .A(y[4]), .B(x[9]), .Z(n396) );
  NANDN U569 ( .A(n620), .B(n396), .Z(n400) );
  OR U570 ( .A(n398), .B(n397), .Z(n399) );
  NAND U571 ( .A(n400), .B(n399), .Z(n476) );
  NANDN U572 ( .A(n401), .B(o[11]), .Z(n483) );
  AND U573 ( .A(x[1]), .B(y[11]), .Z(n403) );
  NAND U574 ( .A(x[6]), .B(y[6]), .Z(n402) );
  XNOR U575 ( .A(n403), .B(n402), .Z(n482) );
  XOR U576 ( .A(n476), .B(n477), .Z(n479) );
  AND U577 ( .A(x[0]), .B(y[12]), .Z(n405) );
  NAND U578 ( .A(y[0]), .B(x[12]), .Z(n404) );
  XOR U579 ( .A(n405), .B(n404), .Z(n487) );
  NAND U580 ( .A(x[11]), .B(y[1]), .Z(n465) );
  XOR U581 ( .A(o[12]), .B(n465), .Z(n486) );
  XOR U582 ( .A(n487), .B(n486), .Z(n472) );
  AND U583 ( .A(x[8]), .B(y[4]), .Z(n407) );
  NAND U584 ( .A(y[10]), .B(x[2]), .Z(n406) );
  XOR U585 ( .A(n407), .B(n406), .Z(n462) );
  NAND U586 ( .A(y[9]), .B(x[3]), .Z(n461) );
  XOR U587 ( .A(n462), .B(n461), .Z(n470) );
  IV U588 ( .A(x[9]), .Z(n2452) );
  ANDN U589 ( .B(y[3]), .A(n2452), .Z(n1180) );
  AND U590 ( .A(y[2]), .B(x[10]), .Z(n1145) );
  NAND U591 ( .A(y[8]), .B(x[4]), .Z(n408) );
  XNOR U592 ( .A(n1145), .B(n408), .Z(n494) );
  NAND U593 ( .A(x[7]), .B(y[5]), .Z(n455) );
  XNOR U594 ( .A(n456), .B(n455), .Z(n457) );
  XNOR U595 ( .A(n458), .B(n457), .Z(n471) );
  XOR U596 ( .A(n472), .B(n473), .Z(n451) );
  ANDN U597 ( .B(y[9]), .A(n2252), .Z(n649) );
  NAND U598 ( .A(n1171), .B(n649), .Z(n412) );
  OR U599 ( .A(n410), .B(n409), .Z(n411) );
  NAND U600 ( .A(n412), .B(n411), .Z(n450) );
  AND U601 ( .A(y[10]), .B(x[6]), .Z(n414) );
  NAND U602 ( .A(n414), .B(n413), .Z(n418) );
  OR U603 ( .A(n416), .B(n415), .Z(n417) );
  NAND U604 ( .A(n418), .B(n417), .Z(n449) );
  XOR U605 ( .A(n450), .B(n449), .Z(n452) );
  XNOR U606 ( .A(n451), .B(n452), .Z(n502) );
  XOR U607 ( .A(n501), .B(n502), .Z(n504) );
  XOR U608 ( .A(n503), .B(n504), .Z(n437) );
  XNOR U609 ( .A(n438), .B(n437), .Z(n439) );
  XNOR U610 ( .A(n440), .B(n439), .Z(n434) );
  NANDN U611 ( .A(n420), .B(n419), .Z(n424) );
  NANDN U612 ( .A(n422), .B(n421), .Z(n423) );
  NAND U613 ( .A(n424), .B(n423), .Z(n431) );
  OR U614 ( .A(n426), .B(n425), .Z(n430) );
  NAND U615 ( .A(n428), .B(n427), .Z(n429) );
  AND U616 ( .A(n430), .B(n429), .Z(n432) );
  XNOR U617 ( .A(n431), .B(n432), .Z(n433) );
  XOR U618 ( .A(n434), .B(n433), .Z(N45) );
  NANDN U619 ( .A(n432), .B(n431), .Z(n436) );
  NANDN U620 ( .A(n434), .B(n433), .Z(n435) );
  NAND U621 ( .A(n436), .B(n435), .Z(n574) );
  OR U622 ( .A(n438), .B(n437), .Z(n442) );
  OR U623 ( .A(n440), .B(n439), .Z(n441) );
  AND U624 ( .A(n442), .B(n441), .Z(n575) );
  XNOR U625 ( .A(n574), .B(n575), .Z(n576) );
  NANDN U626 ( .A(n444), .B(n443), .Z(n448) );
  NAND U627 ( .A(n446), .B(n445), .Z(n447) );
  NAND U628 ( .A(n448), .B(n447), .Z(n583) );
  OR U629 ( .A(n450), .B(n449), .Z(n454) );
  NAND U630 ( .A(n452), .B(n451), .Z(n453) );
  AND U631 ( .A(n454), .B(n453), .Z(n513) );
  NANDN U632 ( .A(n456), .B(n455), .Z(n460) );
  NANDN U633 ( .A(n458), .B(n457), .Z(n459) );
  NAND U634 ( .A(n460), .B(n459), .Z(n508) );
  AND U635 ( .A(x[8]), .B(y[10]), .Z(n909) );
  NAND U636 ( .A(n909), .B(n559), .Z(n464) );
  OR U637 ( .A(n462), .B(n461), .Z(n463) );
  NAND U638 ( .A(n464), .B(n463), .Z(n534) );
  NANDN U639 ( .A(n465), .B(o[12]), .Z(n543) );
  AND U640 ( .A(y[12]), .B(x[1]), .Z(n467) );
  NAND U641 ( .A(y[6]), .B(x[7]), .Z(n466) );
  XNOR U642 ( .A(n467), .B(n466), .Z(n542) );
  AND U643 ( .A(x[2]), .B(y[11]), .Z(n469) );
  NAND U644 ( .A(x[9]), .B(y[4]), .Z(n468) );
  XOR U645 ( .A(n469), .B(n468), .Z(n561) );
  NAND U646 ( .A(x[6]), .B(y[7]), .Z(n560) );
  XOR U647 ( .A(n561), .B(n560), .Z(n531) );
  XNOR U648 ( .A(n534), .B(n533), .Z(n507) );
  XNOR U649 ( .A(n508), .B(n507), .Z(n510) );
  NANDN U650 ( .A(n471), .B(n470), .Z(n475) );
  NANDN U651 ( .A(n473), .B(n472), .Z(n474) );
  AND U652 ( .A(n475), .B(n474), .Z(n509) );
  XOR U653 ( .A(n510), .B(n509), .Z(n514) );
  XOR U654 ( .A(n513), .B(n514), .Z(n515) );
  NANDN U655 ( .A(n477), .B(n476), .Z(n481) );
  NANDN U656 ( .A(n479), .B(n478), .Z(n480) );
  NAND U657 ( .A(n481), .B(n480), .Z(n522) );
  IV U658 ( .A(x[6]), .Z(n2313) );
  ANDN U659 ( .B(y[11]), .A(n2313), .Z(n941) );
  NAND U660 ( .A(n541), .B(n941), .Z(n485) );
  NANDN U661 ( .A(n483), .B(n482), .Z(n484) );
  NAND U662 ( .A(n485), .B(n484), .Z(n527) );
  IV U663 ( .A(y[12]), .Z(n2245) );
  ANDN U664 ( .B(x[12]), .A(n2245), .Z(n1819) );
  NAND U665 ( .A(n707), .B(n1819), .Z(n489) );
  OR U666 ( .A(n487), .B(n486), .Z(n488) );
  NAND U667 ( .A(n489), .B(n488), .Z(n525) );
  AND U668 ( .A(y[5]), .B(x[8]), .Z(n491) );
  NAND U669 ( .A(y[2]), .B(x[11]), .Z(n490) );
  XOR U670 ( .A(n491), .B(n490), .Z(n548) );
  NAND U671 ( .A(y[3]), .B(x[10]), .Z(n547) );
  XNOR U672 ( .A(n548), .B(n547), .Z(n526) );
  XOR U673 ( .A(n525), .B(n526), .Z(n528) );
  AND U674 ( .A(x[10]), .B(y[8]), .Z(n493) );
  NAND U675 ( .A(n493), .B(n492), .Z(n496) );
  NAND U676 ( .A(n494), .B(n1180), .Z(n495) );
  NAND U677 ( .A(n496), .B(n495), .Z(n571) );
  AND U678 ( .A(x[0]), .B(y[13]), .Z(n498) );
  NAND U679 ( .A(x[13]), .B(y[0]), .Z(n497) );
  XOR U680 ( .A(n498), .B(n497), .Z(n556) );
  NAND U681 ( .A(x[12]), .B(y[1]), .Z(n565) );
  XOR U682 ( .A(o[13]), .B(n565), .Z(n555) );
  XOR U683 ( .A(n556), .B(n555), .Z(n569) );
  AND U684 ( .A(x[3]), .B(y[10]), .Z(n500) );
  NAND U685 ( .A(x[5]), .B(y[8]), .Z(n499) );
  XOR U686 ( .A(n500), .B(n499), .Z(n552) );
  NAND U687 ( .A(y[9]), .B(x[4]), .Z(n551) );
  XOR U688 ( .A(n552), .B(n551), .Z(n568) );
  XOR U689 ( .A(n571), .B(n570), .Z(n520) );
  XNOR U690 ( .A(n519), .B(n520), .Z(n521) );
  XOR U691 ( .A(n522), .B(n521), .Z(n516) );
  XNOR U692 ( .A(n515), .B(n516), .Z(n580) );
  NANDN U693 ( .A(n502), .B(n501), .Z(n506) );
  NANDN U694 ( .A(n504), .B(n503), .Z(n505) );
  NAND U695 ( .A(n506), .B(n505), .Z(n581) );
  XOR U696 ( .A(n580), .B(n581), .Z(n582) );
  XNOR U697 ( .A(n583), .B(n582), .Z(n577) );
  XOR U698 ( .A(n576), .B(n577), .Z(N46) );
  OR U699 ( .A(n508), .B(n507), .Z(n512) );
  OR U700 ( .A(n510), .B(n509), .Z(n511) );
  NAND U701 ( .A(n512), .B(n511), .Z(n595) );
  OR U702 ( .A(n514), .B(n513), .Z(n518) );
  NANDN U703 ( .A(n516), .B(n515), .Z(n517) );
  AND U704 ( .A(n518), .B(n517), .Z(n592) );
  NANDN U705 ( .A(n520), .B(n519), .Z(n524) );
  NANDN U706 ( .A(n522), .B(n521), .Z(n523) );
  AND U707 ( .A(n524), .B(n523), .Z(n601) );
  NANDN U708 ( .A(n526), .B(n525), .Z(n530) );
  NANDN U709 ( .A(n528), .B(n527), .Z(n529) );
  NAND U710 ( .A(n530), .B(n529), .Z(n606) );
  NAND U711 ( .A(n532), .B(n531), .Z(n536) );
  NAND U712 ( .A(n534), .B(n533), .Z(n535) );
  AND U713 ( .A(n536), .B(n535), .Z(n605) );
  AND U714 ( .A(y[6]), .B(x[8]), .Z(n538) );
  NAND U715 ( .A(x[3]), .B(y[11]), .Z(n537) );
  XNOR U716 ( .A(n538), .B(n537), .Z(n650) );
  XNOR U717 ( .A(n649), .B(n650), .Z(n662) );
  ANDN U718 ( .B(y[10]), .A(n2454), .Z(n1012) );
  IV U719 ( .A(x[10]), .Z(n2455) );
  ANDN U720 ( .B(y[4]), .A(n2455), .Z(n1255) );
  AND U721 ( .A(y[12]), .B(x[2]), .Z(n540) );
  NAND U722 ( .A(y[5]), .B(x[9]), .Z(n539) );
  XOR U723 ( .A(n540), .B(n539), .Z(n617) );
  XOR U724 ( .A(n1255), .B(n617), .Z(n661) );
  XNOR U725 ( .A(n1012), .B(n661), .Z(n663) );
  ANDN U726 ( .B(x[7]), .A(n2245), .Z(n1164) );
  NAND U727 ( .A(n1164), .B(n541), .Z(n545) );
  NANDN U728 ( .A(n543), .B(n542), .Z(n544) );
  NAND U729 ( .A(n545), .B(n544), .Z(n642) );
  AND U730 ( .A(x[11]), .B(y[5]), .Z(n734) );
  NAND U731 ( .A(n546), .B(n734), .Z(n550) );
  OR U732 ( .A(n548), .B(n547), .Z(n549) );
  AND U733 ( .A(n550), .B(n549), .Z(n643) );
  XOR U734 ( .A(n605), .B(n604), .Z(n607) );
  ANDN U735 ( .B(y[10]), .A(n2252), .Z(n702) );
  NAND U736 ( .A(n1163), .B(n702), .Z(n554) );
  OR U737 ( .A(n552), .B(n551), .Z(n553) );
  NAND U738 ( .A(n554), .B(n553), .Z(n638) );
  ANDN U739 ( .B(y[13]), .A(n25), .Z(n631) );
  ANDN U740 ( .B(x[11]), .A(n20), .Z(n630) );
  XNOR U741 ( .A(n631), .B(n630), .Z(n632) );
  XOR U742 ( .A(n633), .B(n632), .Z(n637) );
  AND U743 ( .A(x[13]), .B(y[13]), .Z(n2147) );
  NAND U744 ( .A(n707), .B(n2147), .Z(n558) );
  OR U745 ( .A(n556), .B(n555), .Z(n557) );
  AND U746 ( .A(n558), .B(n557), .Z(n636) );
  XNOR U747 ( .A(n637), .B(n636), .Z(n639) );
  XOR U748 ( .A(n638), .B(n639), .Z(n668) );
  AND U749 ( .A(y[11]), .B(x[9]), .Z(n1179) );
  NAND U750 ( .A(n1179), .B(n559), .Z(n563) );
  OR U751 ( .A(n561), .B(n560), .Z(n562) );
  AND U752 ( .A(n563), .B(n562), .Z(n613) );
  AND U753 ( .A(y[2]), .B(x[12]), .Z(n1284) );
  NAND U754 ( .A(y[7]), .B(x[7]), .Z(n564) );
  XOR U755 ( .A(n1284), .B(n564), .Z(n622) );
  NAND U756 ( .A(y[1]), .B(x[13]), .Z(n627) );
  XOR U757 ( .A(o[14]), .B(n627), .Z(n621) );
  XOR U758 ( .A(n622), .B(n621), .Z(n611) );
  NANDN U759 ( .A(n565), .B(o[13]), .Z(n654) );
  AND U760 ( .A(x[0]), .B(y[14]), .Z(n567) );
  NAND U761 ( .A(y[0]), .B(x[14]), .Z(n566) );
  XNOR U762 ( .A(n567), .B(n566), .Z(n653) );
  XOR U763 ( .A(n613), .B(n612), .Z(n666) );
  NAND U764 ( .A(n569), .B(n568), .Z(n573) );
  NAND U765 ( .A(n571), .B(n570), .Z(n572) );
  NAND U766 ( .A(n573), .B(n572), .Z(n667) );
  XOR U767 ( .A(n666), .B(n667), .Z(n669) );
  XNOR U768 ( .A(n668), .B(n669), .Z(n599) );
  XOR U769 ( .A(n601), .B(n600), .Z(n593) );
  XNOR U770 ( .A(n592), .B(n593), .Z(n594) );
  XNOR U771 ( .A(n595), .B(n594), .Z(n589) );
  NANDN U772 ( .A(n575), .B(n574), .Z(n579) );
  NANDN U773 ( .A(n577), .B(n576), .Z(n578) );
  NAND U774 ( .A(n579), .B(n578), .Z(n586) );
  OR U775 ( .A(n581), .B(n580), .Z(n585) );
  NANDN U776 ( .A(n583), .B(n582), .Z(n584) );
  NAND U777 ( .A(n585), .B(n584), .Z(n587) );
  XNOR U778 ( .A(n586), .B(n587), .Z(n588) );
  XOR U779 ( .A(n589), .B(n588), .Z(N47) );
  NANDN U780 ( .A(n587), .B(n586), .Z(n591) );
  NANDN U781 ( .A(n589), .B(n588), .Z(n590) );
  NAND U782 ( .A(n591), .B(n590), .Z(n672) );
  OR U783 ( .A(n593), .B(n592), .Z(n597) );
  OR U784 ( .A(n595), .B(n594), .Z(n596) );
  AND U785 ( .A(n597), .B(n596), .Z(n673) );
  XNOR U786 ( .A(n672), .B(n673), .Z(n674) );
  NAND U787 ( .A(n599), .B(n598), .Z(n603) );
  NANDN U788 ( .A(n601), .B(n600), .Z(n602) );
  NAND U789 ( .A(n603), .B(n602), .Z(n681) );
  NANDN U790 ( .A(n605), .B(n604), .Z(n609) );
  NANDN U791 ( .A(n607), .B(n606), .Z(n608) );
  NAND U792 ( .A(n609), .B(n608), .Z(n764) );
  NAND U793 ( .A(n611), .B(n610), .Z(n615) );
  NANDN U794 ( .A(n613), .B(n612), .Z(n614) );
  AND U795 ( .A(n615), .B(n614), .Z(n684) );
  ANDN U796 ( .B(y[12]), .A(n2452), .Z(n1372) );
  NAND U797 ( .A(n616), .B(n1372), .Z(n619) );
  NANDN U798 ( .A(n617), .B(n1255), .Z(n618) );
  NAND U799 ( .A(n619), .B(n618), .Z(n697) );
  ANDN U800 ( .B(x[12]), .A(n2433), .Z(n1172) );
  NANDN U801 ( .A(n620), .B(n1172), .Z(n624) );
  OR U802 ( .A(n622), .B(n621), .Z(n623) );
  NAND U803 ( .A(n624), .B(n623), .Z(n758) );
  NAND U804 ( .A(y[3]), .B(x[12]), .Z(n752) );
  AND U805 ( .A(y[4]), .B(x[11]), .Z(n626) );
  NAND U806 ( .A(y[2]), .B(x[13]), .Z(n625) );
  XOR U807 ( .A(n626), .B(n625), .Z(n751) );
  XNOR U808 ( .A(n752), .B(n751), .Z(n755) );
  NANDN U809 ( .A(n627), .B(o[14]), .Z(n709) );
  AND U810 ( .A(y[0]), .B(x[15]), .Z(n629) );
  NAND U811 ( .A(y[15]), .B(x[0]), .Z(n628) );
  XOR U812 ( .A(n629), .B(n628), .Z(n708) );
  XOR U813 ( .A(n709), .B(n708), .Z(n756) );
  XOR U814 ( .A(n758), .B(n757), .Z(n696) );
  XOR U815 ( .A(n697), .B(n696), .Z(n698) );
  OR U816 ( .A(n631), .B(n630), .Z(n635) );
  OR U817 ( .A(n633), .B(n632), .Z(n634) );
  AND U818 ( .A(n635), .B(n634), .Z(n699) );
  XNOR U819 ( .A(n698), .B(n699), .Z(n685) );
  XOR U820 ( .A(n684), .B(n685), .Z(n686) );
  OR U821 ( .A(n637), .B(n636), .Z(n641) );
  NANDN U822 ( .A(n639), .B(n638), .Z(n640) );
  AND U823 ( .A(n641), .B(n640), .Z(n687) );
  NANDN U824 ( .A(n643), .B(n642), .Z(n647) );
  NAND U825 ( .A(n645), .B(n644), .Z(n646) );
  AND U826 ( .A(n647), .B(n646), .Z(n692) );
  AND U827 ( .A(y[11]), .B(x[8]), .Z(n1030) );
  NANDN U828 ( .A(n648), .B(n1030), .Z(n652) );
  NAND U829 ( .A(n650), .B(n649), .Z(n651) );
  NAND U830 ( .A(n652), .B(n651), .Z(n736) );
  IV U831 ( .A(y[14]), .Z(n2429) );
  ANDN U832 ( .B(x[14]), .A(n2429), .Z(n2466) );
  NAND U833 ( .A(n707), .B(n2466), .Z(n656) );
  NANDN U834 ( .A(n654), .B(n653), .Z(n655) );
  AND U835 ( .A(n656), .B(n655), .Z(n735) );
  NAND U836 ( .A(y[8]), .B(x[7]), .Z(n721) );
  AND U837 ( .A(x[4]), .B(y[11]), .Z(n658) );
  NAND U838 ( .A(y[5]), .B(x[10]), .Z(n657) );
  XOR U839 ( .A(n658), .B(n657), .Z(n720) );
  XNOR U840 ( .A(n721), .B(n720), .Z(n703) );
  AND U841 ( .A(x[6]), .B(y[9]), .Z(n830) );
  XNOR U842 ( .A(n702), .B(n830), .Z(n704) );
  XOR U843 ( .A(n703), .B(n704), .Z(n744) );
  NAND U844 ( .A(x[14]), .B(y[1]), .Z(n724) );
  XOR U845 ( .A(o[15]), .B(n724), .Z(n714) );
  AND U846 ( .A(y[14]), .B(x[1]), .Z(n660) );
  NAND U847 ( .A(y[7]), .B(x[8]), .Z(n659) );
  XOR U848 ( .A(n660), .B(n659), .Z(n713) );
  XNOR U849 ( .A(n714), .B(n713), .Z(n741) );
  ANDN U850 ( .B(x[9]), .A(n23), .Z(n730) );
  ANDN U851 ( .B(y[12]), .A(n27), .Z(n728) );
  ANDN U852 ( .B(y[13]), .A(n26), .Z(n727) );
  XNOR U853 ( .A(n728), .B(n727), .Z(n729) );
  XNOR U854 ( .A(n730), .B(n729), .Z(n742) );
  XOR U855 ( .A(n741), .B(n742), .Z(n743) );
  XNOR U856 ( .A(n744), .B(n743), .Z(n738) );
  XNOR U857 ( .A(n737), .B(n738), .Z(n690) );
  NANDN U858 ( .A(n1012), .B(n661), .Z(n665) );
  NAND U859 ( .A(n663), .B(n662), .Z(n664) );
  NAND U860 ( .A(n665), .B(n664), .Z(n691) );
  XNOR U861 ( .A(n690), .B(n691), .Z(n693) );
  XOR U862 ( .A(n692), .B(n693), .Z(n761) );
  XNOR U863 ( .A(n762), .B(n761), .Z(n763) );
  XNOR U864 ( .A(n764), .B(n763), .Z(n679) );
  NANDN U865 ( .A(n667), .B(n666), .Z(n671) );
  NANDN U866 ( .A(n669), .B(n668), .Z(n670) );
  AND U867 ( .A(n671), .B(n670), .Z(n678) );
  XNOR U868 ( .A(n681), .B(n680), .Z(n675) );
  XOR U869 ( .A(n674), .B(n675), .Z(N48) );
  NANDN U870 ( .A(n673), .B(n672), .Z(n677) );
  NANDN U871 ( .A(n675), .B(n674), .Z(n676) );
  NAND U872 ( .A(n677), .B(n676), .Z(n767) );
  NANDN U873 ( .A(n679), .B(n678), .Z(n683) );
  NANDN U874 ( .A(n681), .B(n680), .Z(n682) );
  NAND U875 ( .A(n683), .B(n682), .Z(n768) );
  XNOR U876 ( .A(n767), .B(n768), .Z(n769) );
  OR U877 ( .A(n685), .B(n684), .Z(n689) );
  NANDN U878 ( .A(n687), .B(n686), .Z(n688) );
  NAND U879 ( .A(n689), .B(n688), .Z(n857) );
  OR U880 ( .A(n691), .B(n690), .Z(n695) );
  OR U881 ( .A(n693), .B(n692), .Z(n694) );
  NAND U882 ( .A(n695), .B(n694), .Z(n855) );
  OR U883 ( .A(n697), .B(n696), .Z(n701) );
  NANDN U884 ( .A(n699), .B(n698), .Z(n700) );
  AND U885 ( .A(n701), .B(n700), .Z(n854) );
  XOR U886 ( .A(n855), .B(n854), .Z(n856) );
  XNOR U887 ( .A(n857), .B(n856), .Z(n776) );
  OR U888 ( .A(n702), .B(n830), .Z(n706) );
  NANDN U889 ( .A(n704), .B(n703), .Z(n705) );
  AND U890 ( .A(n706), .B(n705), .Z(n812) );
  NAND U891 ( .A(x[15]), .B(y[15]), .Z(n2764) );
  NANDN U892 ( .A(n2764), .B(n707), .Z(n711) );
  OR U893 ( .A(n709), .B(n708), .Z(n710) );
  AND U894 ( .A(n711), .B(n710), .Z(n794) );
  ANDN U895 ( .B(y[14]), .A(n29), .Z(n1645) );
  NAND U896 ( .A(n712), .B(n1645), .Z(n716) );
  OR U897 ( .A(n714), .B(n713), .Z(n715) );
  AND U898 ( .A(n716), .B(n715), .Z(n795) );
  XOR U899 ( .A(n794), .B(n795), .Z(n796) );
  NAND U900 ( .A(x[0]), .B(y[16]), .Z(n840) );
  NAND U901 ( .A(x[16]), .B(y[0]), .Z(n839) );
  XOR U902 ( .A(n840), .B(n839), .Z(n841) );
  NAND U903 ( .A(x[15]), .B(y[1]), .Z(n851) );
  XOR U904 ( .A(o[16]), .B(n851), .Z(n842) );
  XOR U905 ( .A(n841), .B(n842), .Z(n825) );
  AND U906 ( .A(y[9]), .B(x[7]), .Z(n718) );
  NAND U907 ( .A(x[6]), .B(y[10]), .Z(n717) );
  XOR U908 ( .A(n718), .B(n717), .Z(n832) );
  NAND U909 ( .A(y[6]), .B(x[10]), .Z(n831) );
  XNOR U910 ( .A(n832), .B(n831), .Z(n824) );
  XNOR U911 ( .A(n825), .B(n824), .Z(n827) );
  ANDN U912 ( .B(y[11]), .A(n2455), .Z(n1413) );
  NANDN U913 ( .A(n719), .B(n1413), .Z(n723) );
  OR U914 ( .A(n721), .B(n720), .Z(n722) );
  AND U915 ( .A(n723), .B(n722), .Z(n826) );
  XNOR U916 ( .A(n827), .B(n826), .Z(n797) );
  XNOR U917 ( .A(n796), .B(n797), .Z(n813) );
  XOR U918 ( .A(n812), .B(n813), .Z(n814) );
  NANDN U919 ( .A(n724), .B(o[15]), .Z(n836) );
  AND U920 ( .A(y[15]), .B(x[1]), .Z(n726) );
  NAND U921 ( .A(y[8]), .B(x[8]), .Z(n725) );
  XOR U922 ( .A(n726), .B(n725), .Z(n835) );
  XNOR U923 ( .A(n836), .B(n835), .Z(n820) );
  OR U924 ( .A(n728), .B(n727), .Z(n732) );
  OR U925 ( .A(n730), .B(n729), .Z(n731) );
  AND U926 ( .A(n732), .B(n731), .Z(n818) );
  NAND U927 ( .A(y[2]), .B(x[14]), .Z(n733) );
  XOR U928 ( .A(n734), .B(n733), .Z(n785) );
  NAND U929 ( .A(y[12]), .B(x[4]), .Z(n784) );
  XOR U930 ( .A(n785), .B(n784), .Z(n819) );
  XNOR U931 ( .A(n818), .B(n819), .Z(n821) );
  XOR U932 ( .A(n820), .B(n821), .Z(n815) );
  XOR U933 ( .A(n814), .B(n815), .Z(n807) );
  NANDN U934 ( .A(n736), .B(n735), .Z(n740) );
  NANDN U935 ( .A(n738), .B(n737), .Z(n739) );
  AND U936 ( .A(n740), .B(n739), .Z(n806) );
  XOR U937 ( .A(n807), .B(n806), .Z(n808) );
  NANDN U938 ( .A(n742), .B(n741), .Z(n746) );
  OR U939 ( .A(n744), .B(n743), .Z(n745) );
  AND U940 ( .A(n746), .B(n745), .Z(n800) );
  AND U941 ( .A(x[2]), .B(y[14]), .Z(n748) );
  NAND U942 ( .A(y[7]), .B(x[9]), .Z(n747) );
  XOR U943 ( .A(n748), .B(n747), .Z(n780) );
  NAND U944 ( .A(y[13]), .B(x[3]), .Z(n779) );
  XOR U945 ( .A(n780), .B(n779), .Z(n788) );
  ANDN U946 ( .B(x[12]), .A(n21), .Z(n1512) );
  AND U947 ( .A(x[13]), .B(y[3]), .Z(n750) );
  NAND U948 ( .A(x[5]), .B(y[11]), .Z(n749) );
  XOR U949 ( .A(n750), .B(n749), .Z(n848) );
  XOR U950 ( .A(n1512), .B(n848), .Z(n789) );
  ANDN U951 ( .B(x[11]), .A(n19), .Z(n1037) );
  IV U952 ( .A(x[13]), .Z(n2049) );
  ANDN U953 ( .B(y[4]), .A(n2049), .Z(n913) );
  NAND U954 ( .A(n1037), .B(n913), .Z(n754) );
  OR U955 ( .A(n752), .B(n751), .Z(n753) );
  AND U956 ( .A(n754), .B(n753), .Z(n790) );
  XOR U957 ( .A(n791), .B(n790), .Z(n801) );
  XOR U958 ( .A(n800), .B(n801), .Z(n802) );
  NANDN U959 ( .A(n756), .B(n755), .Z(n760) );
  NANDN U960 ( .A(n758), .B(n757), .Z(n759) );
  AND U961 ( .A(n760), .B(n759), .Z(n803) );
  XNOR U962 ( .A(n808), .B(n809), .Z(n774) );
  NANDN U963 ( .A(n762), .B(n761), .Z(n766) );
  NAND U964 ( .A(n764), .B(n763), .Z(n765) );
  AND U965 ( .A(n766), .B(n765), .Z(n773) );
  XOR U966 ( .A(n774), .B(n773), .Z(n775) );
  XNOR U967 ( .A(n776), .B(n775), .Z(n770) );
  XOR U968 ( .A(n769), .B(n770), .Z(N49) );
  NANDN U969 ( .A(n768), .B(n767), .Z(n772) );
  NANDN U970 ( .A(n770), .B(n769), .Z(n771) );
  NAND U971 ( .A(n772), .B(n771), .Z(n860) );
  OR U972 ( .A(n774), .B(n773), .Z(n778) );
  NANDN U973 ( .A(n776), .B(n775), .Z(n777) );
  NAND U974 ( .A(n778), .B(n777), .Z(n861) );
  XNOR U975 ( .A(n860), .B(n861), .Z(n862) );
  AND U976 ( .A(x[7]), .B(y[10]), .Z(n948) );
  ANDN U977 ( .B(y[13]), .A(n2454), .Z(n915) );
  ANDN U978 ( .B(x[11]), .A(n23), .Z(n912) );
  XOR U979 ( .A(n913), .B(n912), .Z(n914) );
  ANDN U980 ( .B(y[12]), .A(n2252), .Z(n943) );
  ANDN U981 ( .B(x[8]), .A(n2314), .Z(n940) );
  XOR U982 ( .A(n941), .B(n940), .Z(n942) );
  XNOR U983 ( .A(n943), .B(n942), .Z(n947) );
  XNOR U984 ( .A(n946), .B(n947), .Z(n949) );
  XNOR U985 ( .A(n948), .B(n949), .Z(n954) );
  AND U986 ( .A(y[14]), .B(x[9]), .Z(n1491) );
  NAND U987 ( .A(n1491), .B(n933), .Z(n782) );
  OR U988 ( .A(n780), .B(n779), .Z(n781) );
  NAND U989 ( .A(n782), .B(n781), .Z(n953) );
  AND U990 ( .A(x[14]), .B(y[5]), .Z(n783) );
  NAND U991 ( .A(n783), .B(n1037), .Z(n787) );
  OR U992 ( .A(n785), .B(n784), .Z(n786) );
  AND U993 ( .A(n787), .B(n786), .Z(n952) );
  NANDN U994 ( .A(n789), .B(n788), .Z(n793) );
  OR U995 ( .A(n791), .B(n790), .Z(n792) );
  NAND U996 ( .A(n793), .B(n792), .Z(n873) );
  XOR U997 ( .A(n872), .B(n873), .Z(n875) );
  OR U998 ( .A(n795), .B(n794), .Z(n799) );
  NANDN U999 ( .A(n797), .B(n796), .Z(n798) );
  NAND U1000 ( .A(n799), .B(n798), .Z(n874) );
  XOR U1001 ( .A(n875), .B(n874), .Z(n958) );
  OR U1002 ( .A(n801), .B(n800), .Z(n805) );
  NANDN U1003 ( .A(n803), .B(n802), .Z(n804) );
  NAND U1004 ( .A(n805), .B(n804), .Z(n959) );
  XNOR U1005 ( .A(n958), .B(n959), .Z(n961) );
  OR U1006 ( .A(n807), .B(n806), .Z(n811) );
  NANDN U1007 ( .A(n809), .B(n808), .Z(n810) );
  NAND U1008 ( .A(n811), .B(n810), .Z(n960) );
  XOR U1009 ( .A(n961), .B(n960), .Z(n868) );
  OR U1010 ( .A(n813), .B(n812), .Z(n817) );
  NANDN U1011 ( .A(n815), .B(n814), .Z(n816) );
  NAND U1012 ( .A(n817), .B(n816), .Z(n967) );
  OR U1013 ( .A(n819), .B(n818), .Z(n823) );
  NANDN U1014 ( .A(n821), .B(n820), .Z(n822) );
  NAND U1015 ( .A(n823), .B(n822), .Z(n965) );
  OR U1016 ( .A(n825), .B(n824), .Z(n829) );
  OR U1017 ( .A(n827), .B(n826), .Z(n828) );
  NAND U1018 ( .A(n829), .B(n828), .Z(n881) );
  NAND U1019 ( .A(n948), .B(n830), .Z(n834) );
  OR U1020 ( .A(n832), .B(n831), .Z(n833) );
  NAND U1021 ( .A(n834), .B(n833), .Z(n884) );
  NAND U1022 ( .A(y[15]), .B(x[8]), .Z(n1507) );
  ANDN U1023 ( .B(x[1]), .A(n2430), .Z(n1000) );
  NANDN U1024 ( .A(n1507), .B(n1000), .Z(n838) );
  OR U1025 ( .A(n836), .B(n835), .Z(n837) );
  AND U1026 ( .A(n838), .B(n837), .Z(n885) );
  OR U1027 ( .A(n840), .B(n839), .Z(n844) );
  NANDN U1028 ( .A(n842), .B(n841), .Z(n843) );
  NAND U1029 ( .A(n844), .B(n843), .Z(n891) );
  AND U1030 ( .A(y[15]), .B(x[2]), .Z(n846) );
  NAND U1031 ( .A(y[7]), .B(x[10]), .Z(n845) );
  XOR U1032 ( .A(n846), .B(n845), .Z(n935) );
  NAND U1033 ( .A(y[14]), .B(x[3]), .Z(n934) );
  XOR U1034 ( .A(n935), .B(n934), .Z(n890) );
  XNOR U1035 ( .A(n891), .B(n890), .Z(n893) );
  NAND U1036 ( .A(x[16]), .B(y[1]), .Z(n920) );
  XOR U1037 ( .A(o[17]), .B(n920), .Z(n903) );
  AND U1038 ( .A(y[0]), .B(x[17]), .Z(n902) );
  XOR U1039 ( .A(n903), .B(n902), .Z(n905) );
  AND U1040 ( .A(y[17]), .B(x[0]), .Z(n904) );
  XNOR U1041 ( .A(n905), .B(n904), .Z(n892) );
  XOR U1042 ( .A(n893), .B(n892), .Z(n887) );
  XNOR U1043 ( .A(n886), .B(n887), .Z(n878) );
  ANDN U1044 ( .B(y[11]), .A(n2049), .Z(n1813) );
  NAND U1045 ( .A(n847), .B(n1813), .Z(n850) );
  NANDN U1046 ( .A(n848), .B(n1512), .Z(n849) );
  NAND U1047 ( .A(n850), .B(n849), .Z(n898) );
  NAND U1048 ( .A(x[12]), .B(y[5]), .Z(n925) );
  ANDN U1049 ( .B(x[14]), .A(n20), .Z(n924) );
  NAND U1050 ( .A(x[15]), .B(y[2]), .Z(n923) );
  XOR U1051 ( .A(n924), .B(n923), .Z(n926) );
  XNOR U1052 ( .A(n925), .B(n926), .Z(n897) );
  NANDN U1053 ( .A(n851), .B(o[16]), .Z(n930) );
  AND U1054 ( .A(x[1]), .B(y[16]), .Z(n853) );
  NAND U1055 ( .A(y[8]), .B(x[9]), .Z(n852) );
  XNOR U1056 ( .A(n853), .B(n852), .Z(n929) );
  XOR U1057 ( .A(n897), .B(n896), .Z(n899) );
  XNOR U1058 ( .A(n898), .B(n899), .Z(n879) );
  XNOR U1059 ( .A(n878), .B(n879), .Z(n880) );
  XOR U1060 ( .A(n881), .B(n880), .Z(n964) );
  XNOR U1061 ( .A(n965), .B(n964), .Z(n966) );
  XNOR U1062 ( .A(n967), .B(n966), .Z(n866) );
  OR U1063 ( .A(n855), .B(n854), .Z(n859) );
  NANDN U1064 ( .A(n857), .B(n856), .Z(n858) );
  AND U1065 ( .A(n859), .B(n858), .Z(n867) );
  XOR U1066 ( .A(n866), .B(n867), .Z(n869) );
  XNOR U1067 ( .A(n868), .B(n869), .Z(n863) );
  XOR U1068 ( .A(n862), .B(n863), .Z(N50) );
  NANDN U1069 ( .A(n861), .B(n860), .Z(n865) );
  NANDN U1070 ( .A(n863), .B(n862), .Z(n864) );
  NAND U1071 ( .A(n865), .B(n864), .Z(n1070) );
  NANDN U1072 ( .A(n867), .B(n866), .Z(n871) );
  OR U1073 ( .A(n869), .B(n868), .Z(n870) );
  AND U1074 ( .A(n871), .B(n870), .Z(n1071) );
  XNOR U1075 ( .A(n1070), .B(n1071), .Z(n1072) );
  NANDN U1076 ( .A(n873), .B(n872), .Z(n877) );
  OR U1077 ( .A(n875), .B(n874), .Z(n876) );
  AND U1078 ( .A(n877), .B(n876), .Z(n976) );
  OR U1079 ( .A(n879), .B(n878), .Z(n883) );
  OR U1080 ( .A(n881), .B(n880), .Z(n882) );
  AND U1081 ( .A(n883), .B(n882), .Z(n977) );
  XOR U1082 ( .A(n976), .B(n977), .Z(n979) );
  NANDN U1083 ( .A(n885), .B(n884), .Z(n889) );
  NANDN U1084 ( .A(n887), .B(n886), .Z(n888) );
  NAND U1085 ( .A(n889), .B(n888), .Z(n1048) );
  NAND U1086 ( .A(n891), .B(n890), .Z(n895) );
  NANDN U1087 ( .A(n893), .B(n892), .Z(n894) );
  NAND U1088 ( .A(n895), .B(n894), .Z(n1046) );
  NANDN U1089 ( .A(n897), .B(n896), .Z(n901) );
  NANDN U1090 ( .A(n899), .B(n898), .Z(n900) );
  AND U1091 ( .A(n901), .B(n900), .Z(n1047) );
  XOR U1092 ( .A(n1048), .B(n1049), .Z(n972) );
  NANDN U1093 ( .A(n903), .B(n902), .Z(n907) );
  NANDN U1094 ( .A(n905), .B(n904), .Z(n906) );
  NAND U1095 ( .A(n907), .B(n906), .Z(n1053) );
  NAND U1096 ( .A(x[4]), .B(y[14]), .Z(n908) );
  XOR U1097 ( .A(n909), .B(n908), .Z(n1014) );
  NAND U1098 ( .A(x[7]), .B(y[11]), .Z(n1013) );
  XNOR U1099 ( .A(n1014), .B(n1013), .Z(n1042) );
  ANDN U1100 ( .B(y[12]), .A(n2313), .Z(n1536) );
  NAND U1101 ( .A(y[13]), .B(x[5]), .Z(n1124) );
  XOR U1102 ( .A(n1536), .B(n1124), .Z(n1043) );
  XNOR U1103 ( .A(n1053), .B(n1052), .Z(n1054) );
  NAND U1104 ( .A(x[2]), .B(y[16]), .Z(n1039) );
  AND U1105 ( .A(y[2]), .B(x[16]), .Z(n911) );
  NAND U1106 ( .A(y[7]), .B(x[11]), .Z(n910) );
  XOR U1107 ( .A(n911), .B(n910), .Z(n1038) );
  XOR U1108 ( .A(n1039), .B(n1038), .Z(n1055) );
  XOR U1109 ( .A(n1054), .B(n1055), .Z(n1066) );
  OR U1110 ( .A(n913), .B(n912), .Z(n917) );
  NANDN U1111 ( .A(n915), .B(n914), .Z(n916) );
  NAND U1112 ( .A(n917), .B(n916), .Z(n991) );
  AND U1113 ( .A(y[3]), .B(x[15]), .Z(n919) );
  NAND U1114 ( .A(y[9]), .B(x[9]), .Z(n918) );
  XOR U1115 ( .A(n919), .B(n918), .Z(n1032) );
  NAND U1116 ( .A(x[14]), .B(y[4]), .Z(n1031) );
  XOR U1117 ( .A(n1032), .B(n1031), .Z(n989) );
  NANDN U1118 ( .A(n920), .B(o[17]), .Z(n1002) );
  AND U1119 ( .A(y[17]), .B(x[1]), .Z(n922) );
  NAND U1120 ( .A(y[8]), .B(x[10]), .Z(n921) );
  XNOR U1121 ( .A(n922), .B(n921), .Z(n1001) );
  XOR U1122 ( .A(n991), .B(n990), .Z(n1065) );
  NANDN U1123 ( .A(n924), .B(n923), .Z(n928) );
  NANDN U1124 ( .A(n926), .B(n925), .Z(n927) );
  AND U1125 ( .A(n928), .B(n927), .Z(n1064) );
  XOR U1126 ( .A(n1065), .B(n1064), .Z(n1067) );
  XNOR U1127 ( .A(n1066), .B(n1067), .Z(n971) );
  IV U1128 ( .A(y[16]), .Z(n1162) );
  ANDN U1129 ( .B(x[9]), .A(n1162), .Z(n1904) );
  NAND U1130 ( .A(n1904), .B(n1000), .Z(n932) );
  NANDN U1131 ( .A(n930), .B(n929), .Z(n931) );
  NAND U1132 ( .A(n932), .B(n931), .Z(n1061) );
  IV U1133 ( .A(y[15]), .Z(n2048) );
  ANDN U1134 ( .B(x[10]), .A(n2048), .Z(n1905) );
  NAND U1135 ( .A(n933), .B(n1905), .Z(n937) );
  OR U1136 ( .A(n935), .B(n934), .Z(n936) );
  NAND U1137 ( .A(n937), .B(n936), .Z(n997) );
  NAND U1138 ( .A(x[0]), .B(y[18]), .Z(n1006) );
  NAND U1139 ( .A(y[0]), .B(x[18]), .Z(n1005) );
  XOR U1140 ( .A(n1006), .B(n1005), .Z(n1007) );
  NAND U1141 ( .A(x[17]), .B(y[1]), .Z(n1019) );
  XOR U1142 ( .A(o[18]), .B(n1019), .Z(n1008) );
  XOR U1143 ( .A(n1007), .B(n1008), .Z(n995) );
  AND U1144 ( .A(y[15]), .B(x[3]), .Z(n939) );
  NAND U1145 ( .A(x[13]), .B(y[5]), .Z(n938) );
  XOR U1146 ( .A(n939), .B(n938), .Z(n1022) );
  NAND U1147 ( .A(x[12]), .B(y[6]), .Z(n1021) );
  XOR U1148 ( .A(n1022), .B(n1021), .Z(n994) );
  XNOR U1149 ( .A(n995), .B(n994), .Z(n996) );
  XOR U1150 ( .A(n997), .B(n996), .Z(n1058) );
  OR U1151 ( .A(n941), .B(n940), .Z(n945) );
  NANDN U1152 ( .A(n943), .B(n942), .Z(n944) );
  AND U1153 ( .A(n945), .B(n944), .Z(n1059) );
  XNOR U1154 ( .A(n1058), .B(n1059), .Z(n1060) );
  XNOR U1155 ( .A(n1061), .B(n1060), .Z(n982) );
  NANDN U1156 ( .A(n947), .B(n946), .Z(n951) );
  NAND U1157 ( .A(n949), .B(n948), .Z(n950) );
  AND U1158 ( .A(n951), .B(n950), .Z(n983) );
  XOR U1159 ( .A(n982), .B(n983), .Z(n985) );
  NANDN U1160 ( .A(n953), .B(n952), .Z(n957) );
  NAND U1161 ( .A(n955), .B(n954), .Z(n956) );
  AND U1162 ( .A(n957), .B(n956), .Z(n984) );
  XOR U1163 ( .A(n971), .B(n970), .Z(n973) );
  XNOR U1164 ( .A(n972), .B(n973), .Z(n978) );
  XNOR U1165 ( .A(n979), .B(n978), .Z(n1079) );
  OR U1166 ( .A(n959), .B(n958), .Z(n963) );
  OR U1167 ( .A(n961), .B(n960), .Z(n962) );
  NAND U1168 ( .A(n963), .B(n962), .Z(n1077) );
  OR U1169 ( .A(n965), .B(n964), .Z(n969) );
  OR U1170 ( .A(n967), .B(n966), .Z(n968) );
  NAND U1171 ( .A(n969), .B(n968), .Z(n1076) );
  XNOR U1172 ( .A(n1077), .B(n1076), .Z(n1078) );
  XNOR U1173 ( .A(n1079), .B(n1078), .Z(n1073) );
  XOR U1174 ( .A(n1072), .B(n1073), .Z(N51) );
  NANDN U1175 ( .A(n971), .B(n970), .Z(n975) );
  NANDN U1176 ( .A(n973), .B(n972), .Z(n974) );
  AND U1177 ( .A(n975), .B(n974), .Z(n1088) );
  OR U1178 ( .A(n977), .B(n976), .Z(n981) );
  NAND U1179 ( .A(n979), .B(n978), .Z(n980) );
  AND U1180 ( .A(n981), .B(n980), .Z(n1089) );
  XNOR U1181 ( .A(n1088), .B(n1089), .Z(n1091) );
  NANDN U1182 ( .A(n983), .B(n982), .Z(n987) );
  NANDN U1183 ( .A(n985), .B(n984), .Z(n986) );
  NAND U1184 ( .A(n987), .B(n986), .Z(n1097) );
  NAND U1185 ( .A(n989), .B(n988), .Z(n993) );
  NANDN U1186 ( .A(n991), .B(n990), .Z(n992) );
  NAND U1187 ( .A(n993), .B(n992), .Z(n1113) );
  NANDN U1188 ( .A(n995), .B(n994), .Z(n999) );
  NAND U1189 ( .A(n997), .B(n996), .Z(n998) );
  NAND U1190 ( .A(n999), .B(n998), .Z(n1112) );
  XOR U1191 ( .A(n1113), .B(n1112), .Z(n1114) );
  ANDN U1192 ( .B(y[17]), .A(n2455), .Z(n2302) );
  NAND U1193 ( .A(n1000), .B(n2302), .Z(n1004) );
  NANDN U1194 ( .A(n1002), .B(n1001), .Z(n1003) );
  AND U1195 ( .A(n1004), .B(n1003), .Z(n1120) );
  OR U1196 ( .A(n1006), .B(n1005), .Z(n1010) );
  NANDN U1197 ( .A(n1008), .B(n1007), .Z(n1009) );
  NAND U1198 ( .A(n1010), .B(n1009), .Z(n1119) );
  AND U1199 ( .A(x[16]), .B(y[3]), .Z(n1651) );
  NAND U1200 ( .A(y[10]), .B(x[9]), .Z(n1011) );
  XOR U1201 ( .A(n1651), .B(n1011), .Z(n1182) );
  NAND U1202 ( .A(x[15]), .B(y[4]), .Z(n1181) );
  XOR U1203 ( .A(n1182), .B(n1181), .Z(n1118) );
  XNOR U1204 ( .A(n1119), .B(n1118), .Z(n1121) );
  XNOR U1205 ( .A(n1120), .B(n1121), .Z(n1108) );
  NAND U1206 ( .A(n1012), .B(n1645), .Z(n1016) );
  OR U1207 ( .A(n1014), .B(n1013), .Z(n1015) );
  NAND U1208 ( .A(n1016), .B(n1015), .Z(n1157) );
  NAND U1209 ( .A(y[15]), .B(x[4]), .Z(n1239) );
  AND U1210 ( .A(x[6]), .B(y[13]), .Z(n1018) );
  NAND U1211 ( .A(x[5]), .B(y[14]), .Z(n1017) );
  XNOR U1212 ( .A(n1018), .B(n1017), .Z(n1125) );
  XNOR U1213 ( .A(n1157), .B(n1156), .Z(n1159) );
  NANDN U1214 ( .A(n1019), .B(o[18]), .Z(n1131) );
  NAND U1215 ( .A(x[0]), .B(y[19]), .Z(n1129) );
  NAND U1216 ( .A(y[0]), .B(x[19]), .Z(n1128) );
  XOR U1217 ( .A(n1129), .B(n1128), .Z(n1130) );
  XNOR U1218 ( .A(n1131), .B(n1130), .Z(n1158) );
  XOR U1219 ( .A(n1159), .B(n1158), .Z(n1106) );
  ANDN U1220 ( .B(y[15]), .A(n2049), .Z(n2442) );
  NAND U1221 ( .A(n1020), .B(n2442), .Z(n1024) );
  OR U1222 ( .A(n1022), .B(n1021), .Z(n1023) );
  NAND U1223 ( .A(n1024), .B(n1023), .Z(n1153) );
  AND U1224 ( .A(x[3]), .B(y[16]), .Z(n1026) );
  NAND U1225 ( .A(y[8]), .B(x[11]), .Z(n1025) );
  XOR U1226 ( .A(n1026), .B(n1025), .Z(n1165) );
  XOR U1227 ( .A(n1164), .B(n1165), .Z(n1150) );
  NAND U1228 ( .A(y[1]), .B(x[18]), .Z(n1170) );
  XOR U1229 ( .A(o[19]), .B(n1170), .Z(n1147) );
  AND U1230 ( .A(y[9]), .B(x[10]), .Z(n1028) );
  NAND U1231 ( .A(y[2]), .B(x[17]), .Z(n1027) );
  XOR U1232 ( .A(n1028), .B(n1027), .Z(n1146) );
  XOR U1233 ( .A(n1147), .B(n1146), .Z(n1151) );
  XNOR U1234 ( .A(n1150), .B(n1151), .Z(n1152) );
  XOR U1235 ( .A(n1153), .B(n1152), .Z(n1107) );
  XOR U1236 ( .A(n1106), .B(n1107), .Z(n1109) );
  XOR U1237 ( .A(n1108), .B(n1109), .Z(n1115) );
  XOR U1238 ( .A(n1114), .B(n1115), .Z(n1095) );
  NAND U1239 ( .A(y[5]), .B(x[14]), .Z(n1029) );
  XOR U1240 ( .A(n1030), .B(n1029), .Z(n1142) );
  NAND U1241 ( .A(x[1]), .B(y[18]), .Z(n1141) );
  XOR U1242 ( .A(n1142), .B(n1141), .Z(n1188) );
  ANDN U1243 ( .B(x[15]), .A(n2314), .Z(n1838) );
  NAND U1244 ( .A(n1838), .B(n1180), .Z(n1034) );
  OR U1245 ( .A(n1032), .B(n1031), .Z(n1033) );
  NAND U1246 ( .A(n1034), .B(n1033), .Z(n1185) );
  AND U1247 ( .A(y[17]), .B(x[2]), .Z(n1036) );
  NAND U1248 ( .A(x[13]), .B(y[6]), .Z(n1035) );
  XNOR U1249 ( .A(n1036), .B(n1035), .Z(n1173) );
  XNOR U1250 ( .A(n1172), .B(n1173), .Z(n1186) );
  AND U1251 ( .A(x[16]), .B(y[7]), .Z(n1505) );
  NAND U1252 ( .A(n1505), .B(n1037), .Z(n1041) );
  OR U1253 ( .A(n1039), .B(n1038), .Z(n1040) );
  AND U1254 ( .A(n1041), .B(n1040), .Z(n1101) );
  XOR U1255 ( .A(n1100), .B(n1101), .Z(n1103) );
  NANDN U1256 ( .A(n1536), .B(n1124), .Z(n1045) );
  NANDN U1257 ( .A(n1043), .B(n1042), .Z(n1044) );
  NAND U1258 ( .A(n1045), .B(n1044), .Z(n1102) );
  XOR U1259 ( .A(n1103), .B(n1102), .Z(n1094) );
  XOR U1260 ( .A(n1095), .B(n1094), .Z(n1096) );
  XOR U1261 ( .A(n1097), .B(n1096), .Z(n1194) );
  NANDN U1262 ( .A(n1047), .B(n1046), .Z(n1051) );
  NANDN U1263 ( .A(n1049), .B(n1048), .Z(n1050) );
  NAND U1264 ( .A(n1051), .B(n1050), .Z(n1192) );
  NANDN U1265 ( .A(n1053), .B(n1052), .Z(n1057) );
  NANDN U1266 ( .A(n1055), .B(n1054), .Z(n1056) );
  AND U1267 ( .A(n1057), .B(n1056), .Z(n1200) );
  OR U1268 ( .A(n1059), .B(n1058), .Z(n1063) );
  OR U1269 ( .A(n1061), .B(n1060), .Z(n1062) );
  AND U1270 ( .A(n1063), .B(n1062), .Z(n1197) );
  NANDN U1271 ( .A(n1065), .B(n1064), .Z(n1069) );
  NANDN U1272 ( .A(n1067), .B(n1066), .Z(n1068) );
  NAND U1273 ( .A(n1069), .B(n1068), .Z(n1198) );
  XNOR U1274 ( .A(n1197), .B(n1198), .Z(n1199) );
  XOR U1275 ( .A(n1200), .B(n1199), .Z(n1191) );
  XNOR U1276 ( .A(n1192), .B(n1191), .Z(n1193) );
  XOR U1277 ( .A(n1194), .B(n1193), .Z(n1090) );
  XOR U1278 ( .A(n1091), .B(n1090), .Z(n1084) );
  NANDN U1279 ( .A(n1071), .B(n1070), .Z(n1075) );
  NANDN U1280 ( .A(n1073), .B(n1072), .Z(n1074) );
  NAND U1281 ( .A(n1075), .B(n1074), .Z(n1082) );
  OR U1282 ( .A(n1077), .B(n1076), .Z(n1081) );
  OR U1283 ( .A(n1079), .B(n1078), .Z(n1080) );
  AND U1284 ( .A(n1081), .B(n1080), .Z(n1083) );
  XNOR U1285 ( .A(n1082), .B(n1083), .Z(n1085) );
  XNOR U1286 ( .A(n1084), .B(n1085), .Z(N52) );
  NANDN U1287 ( .A(n1083), .B(n1082), .Z(n1087) );
  NAND U1288 ( .A(n1085), .B(n1084), .Z(n1086) );
  NAND U1289 ( .A(n1087), .B(n1086), .Z(n1203) );
  OR U1290 ( .A(n1089), .B(n1088), .Z(n1093) );
  OR U1291 ( .A(n1091), .B(n1090), .Z(n1092) );
  AND U1292 ( .A(n1093), .B(n1092), .Z(n1204) );
  XNOR U1293 ( .A(n1203), .B(n1204), .Z(n1205) );
  OR U1294 ( .A(n1095), .B(n1094), .Z(n1099) );
  NANDN U1295 ( .A(n1097), .B(n1096), .Z(n1098) );
  NAND U1296 ( .A(n1099), .B(n1098), .Z(n1309) );
  NANDN U1297 ( .A(n1101), .B(n1100), .Z(n1105) );
  OR U1298 ( .A(n1103), .B(n1102), .Z(n1104) );
  AND U1299 ( .A(n1105), .B(n1104), .Z(n1315) );
  NANDN U1300 ( .A(n1107), .B(n1106), .Z(n1111) );
  NANDN U1301 ( .A(n1109), .B(n1108), .Z(n1110) );
  NAND U1302 ( .A(n1111), .B(n1110), .Z(n1313) );
  OR U1303 ( .A(n1113), .B(n1112), .Z(n1117) );
  NANDN U1304 ( .A(n1115), .B(n1114), .Z(n1116) );
  NAND U1305 ( .A(n1117), .B(n1116), .Z(n1312) );
  XOR U1306 ( .A(n1313), .B(n1312), .Z(n1314) );
  NAND U1307 ( .A(n1119), .B(n1118), .Z(n1123) );
  OR U1308 ( .A(n1121), .B(n1120), .Z(n1122) );
  NAND U1309 ( .A(n1123), .B(n1122), .Z(n1303) );
  ANDN U1310 ( .B(y[14]), .A(n2313), .Z(n1278) );
  NANDN U1311 ( .A(n1124), .B(n1278), .Z(n1127) );
  NANDN U1312 ( .A(n1239), .B(n1125), .Z(n1126) );
  NAND U1313 ( .A(n1127), .B(n1126), .Z(n1274) );
  OR U1314 ( .A(n1129), .B(n1128), .Z(n1133) );
  NANDN U1315 ( .A(n1131), .B(n1130), .Z(n1132) );
  NAND U1316 ( .A(n1133), .B(n1132), .Z(n1272) );
  AND U1317 ( .A(x[18]), .B(y[2]), .Z(n1135) );
  NAND U1318 ( .A(y[8]), .B(x[12]), .Z(n1134) );
  XOR U1319 ( .A(n1135), .B(n1134), .Z(n1286) );
  NAND U1320 ( .A(y[3]), .B(x[17]), .Z(n1285) );
  XNOR U1321 ( .A(n1286), .B(n1285), .Z(n1273) );
  XOR U1322 ( .A(n1272), .B(n1273), .Z(n1275) );
  AND U1323 ( .A(y[17]), .B(x[3]), .Z(n1137) );
  NAND U1324 ( .A(y[7]), .B(x[13]), .Z(n1136) );
  XOR U1325 ( .A(n1137), .B(n1136), .Z(n1252) );
  NAND U1326 ( .A(y[12]), .B(x[8]), .Z(n1251) );
  XOR U1327 ( .A(n1252), .B(n1251), .Z(n1280) );
  AND U1328 ( .A(x[4]), .B(y[16]), .Z(n1139) );
  NAND U1329 ( .A(x[5]), .B(y[15]), .Z(n1138) );
  XOR U1330 ( .A(n1139), .B(n1138), .Z(n1241) );
  NAND U1331 ( .A(y[13]), .B(x[7]), .Z(n1240) );
  XOR U1332 ( .A(n1241), .B(n1240), .Z(n1279) );
  XNOR U1333 ( .A(n1278), .B(n1279), .Z(n1281) );
  XOR U1334 ( .A(n1280), .B(n1281), .Z(n1224) );
  NANDN U1335 ( .A(n1140), .B(n1964), .Z(n1144) );
  OR U1336 ( .A(n1142), .B(n1141), .Z(n1143) );
  NAND U1337 ( .A(n1144), .B(n1143), .Z(n1222) );
  IV U1338 ( .A(x[17]), .Z(n2483) );
  ANDN U1339 ( .B(y[9]), .A(n2483), .Z(n2094) );
  NAND U1340 ( .A(n1145), .B(n2094), .Z(n1149) );
  OR U1341 ( .A(n1147), .B(n1146), .Z(n1148) );
  AND U1342 ( .A(n1149), .B(n1148), .Z(n1221) );
  XNOR U1343 ( .A(n1224), .B(n1223), .Z(n1301) );
  XNOR U1344 ( .A(n1300), .B(n1301), .Z(n1302) );
  XOR U1345 ( .A(n1303), .B(n1302), .Z(n1260) );
  NANDN U1346 ( .A(n1151), .B(n1150), .Z(n1155) );
  NANDN U1347 ( .A(n1153), .B(n1152), .Z(n1154) );
  NAND U1348 ( .A(n1155), .B(n1154), .Z(n1261) );
  NAND U1349 ( .A(n1157), .B(n1156), .Z(n1161) );
  NANDN U1350 ( .A(n1159), .B(n1158), .Z(n1160) );
  AND U1351 ( .A(n1161), .B(n1160), .Z(n1269) );
  IV U1352 ( .A(x[11]), .Z(n2482) );
  NOR U1353 ( .A(n1162), .B(n2482), .Z(n2303) );
  NAND U1354 ( .A(n2303), .B(n1163), .Z(n1167) );
  NANDN U1355 ( .A(n1165), .B(n1164), .Z(n1166) );
  NAND U1356 ( .A(n1167), .B(n1166), .Z(n1235) );
  AND U1357 ( .A(y[19]), .B(x[1]), .Z(n1169) );
  NAND U1358 ( .A(y[9]), .B(x[11]), .Z(n1168) );
  XOR U1359 ( .A(n1169), .B(n1168), .Z(n1291) );
  AND U1360 ( .A(x[19]), .B(y[1]), .Z(n1299) );
  XOR U1361 ( .A(o[20]), .B(n1299), .Z(n1290) );
  XOR U1362 ( .A(n1291), .B(n1290), .Z(n1234) );
  NANDN U1363 ( .A(n1170), .B(o[19]), .Z(n1247) );
  NAND U1364 ( .A(x[0]), .B(y[20]), .Z(n1245) );
  NAND U1365 ( .A(y[0]), .B(x[20]), .Z(n1244) );
  XOR U1366 ( .A(n1245), .B(n1244), .Z(n1246) );
  XNOR U1367 ( .A(n1247), .B(n1246), .Z(n1233) );
  XOR U1368 ( .A(n1234), .B(n1233), .Z(n1236) );
  XOR U1369 ( .A(n1235), .B(n1236), .Z(n1217) );
  NAND U1370 ( .A(x[13]), .B(y[17]), .Z(n2660) );
  NANDN U1371 ( .A(n2660), .B(n1171), .Z(n1175) );
  NAND U1372 ( .A(n1173), .B(n1172), .Z(n1174) );
  AND U1373 ( .A(n1175), .B(n1174), .Z(n1230) );
  AND U1374 ( .A(x[16]), .B(y[4]), .Z(n1177) );
  NAND U1375 ( .A(y[10]), .B(x[10]), .Z(n1176) );
  XOR U1376 ( .A(n1177), .B(n1176), .Z(n1257) );
  NAND U1377 ( .A(x[2]), .B(y[18]), .Z(n1256) );
  XOR U1378 ( .A(n1257), .B(n1256), .Z(n1228) );
  NAND U1379 ( .A(y[5]), .B(x[15]), .Z(n1178) );
  XOR U1380 ( .A(n1179), .B(n1178), .Z(n1296) );
  NAND U1381 ( .A(x[14]), .B(y[6]), .Z(n1295) );
  XOR U1382 ( .A(n1296), .B(n1295), .Z(n1227) );
  XOR U1383 ( .A(n1230), .B(n1229), .Z(n1215) );
  IV U1384 ( .A(y[10]), .Z(n2500) );
  ANDN U1385 ( .B(x[16]), .A(n2500), .Z(n2081) );
  NAND U1386 ( .A(n1180), .B(n2081), .Z(n1184) );
  OR U1387 ( .A(n1182), .B(n1181), .Z(n1183) );
  NAND U1388 ( .A(n1184), .B(n1183), .Z(n1216) );
  XOR U1389 ( .A(n1215), .B(n1216), .Z(n1218) );
  XNOR U1390 ( .A(n1217), .B(n1218), .Z(n1267) );
  NANDN U1391 ( .A(n1186), .B(n1185), .Z(n1190) );
  NAND U1392 ( .A(n1188), .B(n1187), .Z(n1189) );
  AND U1393 ( .A(n1190), .B(n1189), .Z(n1266) );
  XNOR U1394 ( .A(n1267), .B(n1266), .Z(n1268) );
  XOR U1395 ( .A(n1269), .B(n1268), .Z(n1262) );
  XOR U1396 ( .A(n1307), .B(n1306), .Z(n1308) );
  XNOR U1397 ( .A(n1309), .B(n1308), .Z(n1210) );
  NANDN U1398 ( .A(n1192), .B(n1191), .Z(n1196) );
  NANDN U1399 ( .A(n1194), .B(n1193), .Z(n1195) );
  AND U1400 ( .A(n1196), .B(n1195), .Z(n1209) );
  OR U1401 ( .A(n1198), .B(n1197), .Z(n1202) );
  OR U1402 ( .A(n1200), .B(n1199), .Z(n1201) );
  NAND U1403 ( .A(n1202), .B(n1201), .Z(n1212) );
  XNOR U1404 ( .A(n1211), .B(n1212), .Z(n1206) );
  XOR U1405 ( .A(n1205), .B(n1206), .Z(N53) );
  NANDN U1406 ( .A(n1204), .B(n1203), .Z(n1208) );
  NANDN U1407 ( .A(n1206), .B(n1205), .Z(n1207) );
  NAND U1408 ( .A(n1208), .B(n1207), .Z(n1318) );
  NANDN U1409 ( .A(n1210), .B(n1209), .Z(n1214) );
  NANDN U1410 ( .A(n1212), .B(n1211), .Z(n1213) );
  NAND U1411 ( .A(n1214), .B(n1213), .Z(n1319) );
  XNOR U1412 ( .A(n1318), .B(n1319), .Z(n1320) );
  NANDN U1413 ( .A(n1216), .B(n1215), .Z(n1220) );
  NANDN U1414 ( .A(n1218), .B(n1217), .Z(n1219) );
  NAND U1415 ( .A(n1220), .B(n1219), .Z(n1439) );
  NANDN U1416 ( .A(n1222), .B(n1221), .Z(n1226) );
  NAND U1417 ( .A(n1224), .B(n1223), .Z(n1225) );
  AND U1418 ( .A(n1226), .B(n1225), .Z(n1443) );
  NAND U1419 ( .A(n1228), .B(n1227), .Z(n1232) );
  NANDN U1420 ( .A(n1230), .B(n1229), .Z(n1231) );
  NAND U1421 ( .A(n1232), .B(n1231), .Z(n1444) );
  XOR U1422 ( .A(n1443), .B(n1444), .Z(n1445) );
  NANDN U1423 ( .A(n1234), .B(n1233), .Z(n1238) );
  NANDN U1424 ( .A(n1236), .B(n1235), .Z(n1237) );
  NAND U1425 ( .A(n1238), .B(n1237), .Z(n1446) );
  ANDN U1426 ( .B(y[16]), .A(n2252), .Z(n1416) );
  NANDN U1427 ( .A(n1239), .B(n1416), .Z(n1243) );
  OR U1428 ( .A(n1241), .B(n1240), .Z(n1242) );
  NAND U1429 ( .A(n1243), .B(n1242), .Z(n1342) );
  OR U1430 ( .A(n1245), .B(n1244), .Z(n1249) );
  NANDN U1431 ( .A(n1247), .B(n1246), .Z(n1248) );
  AND U1432 ( .A(n1249), .B(n1248), .Z(n1343) );
  ANDN U1433 ( .B(x[13]), .A(n2430), .Z(n1426) );
  ANDN U1434 ( .B(y[17]), .A(n2454), .Z(n1424) );
  ANDN U1435 ( .B(y[18]), .A(n27), .Z(n1425) );
  XNOR U1436 ( .A(n1424), .B(n1425), .Z(n1427) );
  XNOR U1437 ( .A(n1426), .B(n1427), .Z(n1432) );
  ANDN U1438 ( .B(y[15]), .A(n2313), .Z(n1398) );
  ANDN U1439 ( .B(y[14]), .A(n28), .Z(n1506) );
  ANDN U1440 ( .B(x[14]), .A(n2433), .Z(n1397) );
  XNOR U1441 ( .A(n1506), .B(n1397), .Z(n1399) );
  XNOR U1442 ( .A(n1398), .B(n1399), .Z(n1374) );
  NAND U1443 ( .A(y[13]), .B(x[8]), .Z(n1808) );
  XOR U1444 ( .A(n1372), .B(n1808), .Z(n1373) );
  XNOR U1445 ( .A(n1374), .B(n1373), .Z(n1431) );
  XNOR U1446 ( .A(n1432), .B(n1431), .Z(n1434) );
  ANDN U1447 ( .B(x[12]), .A(n2314), .Z(n1379) );
  IV U1448 ( .A(y[19]), .Z(n2140) );
  ANDN U1449 ( .B(x[2]), .A(n2140), .Z(n1377) );
  ANDN U1450 ( .B(y[4]), .A(n2483), .Z(n1378) );
  XNOR U1451 ( .A(n1377), .B(n1378), .Z(n1380) );
  XNOR U1452 ( .A(n1379), .B(n1380), .Z(n1433) );
  XOR U1453 ( .A(n1434), .B(n1433), .Z(n1345) );
  XNOR U1454 ( .A(n1344), .B(n1345), .Z(n1369) );
  NAND U1455 ( .A(y[10]), .B(x[11]), .Z(n1388) );
  NAND U1456 ( .A(y[1]), .B(x[20]), .Z(n1430) );
  XOR U1457 ( .A(o[21]), .B(n1430), .Z(n1386) );
  NAND U1458 ( .A(y[2]), .B(x[19]), .Z(n1385) );
  XNOR U1459 ( .A(n1386), .B(n1385), .Z(n1387) );
  XNOR U1460 ( .A(n1388), .B(n1387), .Z(n1349) );
  IV U1461 ( .A(y[20]), .Z(n2453) );
  ANDN U1462 ( .B(x[1]), .A(n2453), .Z(n1411) );
  NAND U1463 ( .A(y[3]), .B(x[18]), .Z(n1410) );
  XOR U1464 ( .A(n1411), .B(n1410), .Z(n1412) );
  XOR U1465 ( .A(n1413), .B(n1412), .Z(n1348) );
  XOR U1466 ( .A(n1349), .B(n1348), .Z(n1350) );
  NANDN U1467 ( .A(n2660), .B(n1250), .Z(n1254) );
  OR U1468 ( .A(n1252), .B(n1251), .Z(n1253) );
  AND U1469 ( .A(n1254), .B(n1253), .Z(n1351) );
  XOR U1470 ( .A(n1350), .B(n1351), .Z(n1366) );
  NAND U1471 ( .A(n1255), .B(n2081), .Z(n1259) );
  OR U1472 ( .A(n1257), .B(n1256), .Z(n1258) );
  NAND U1473 ( .A(n1259), .B(n1258), .Z(n1367) );
  XOR U1474 ( .A(n1369), .B(n1368), .Z(n1437) );
  XOR U1475 ( .A(n1438), .B(n1437), .Z(n1440) );
  XOR U1476 ( .A(n1439), .B(n1440), .Z(n1330) );
  NANDN U1477 ( .A(n1261), .B(n1260), .Z(n1265) );
  NAND U1478 ( .A(n1263), .B(n1262), .Z(n1264) );
  AND U1479 ( .A(n1265), .B(n1264), .Z(n1331) );
  XOR U1480 ( .A(n1330), .B(n1331), .Z(n1332) );
  OR U1481 ( .A(n1267), .B(n1266), .Z(n1271) );
  OR U1482 ( .A(n1269), .B(n1268), .Z(n1270) );
  NAND U1483 ( .A(n1271), .B(n1270), .Z(n1338) );
  NANDN U1484 ( .A(n1273), .B(n1272), .Z(n1277) );
  NANDN U1485 ( .A(n1275), .B(n1274), .Z(n1276) );
  NAND U1486 ( .A(n1277), .B(n1276), .Z(n1363) );
  NAND U1487 ( .A(n1279), .B(n1278), .Z(n1283) );
  NANDN U1488 ( .A(n1281), .B(n1280), .Z(n1282) );
  NAND U1489 ( .A(n1283), .B(n1282), .Z(n1360) );
  ANDN U1490 ( .B(x[18]), .A(n2430), .Z(n2092) );
  NAND U1491 ( .A(n1284), .B(n2092), .Z(n1288) );
  OR U1492 ( .A(n1286), .B(n1285), .Z(n1287) );
  NAND U1493 ( .A(n1288), .B(n1287), .Z(n1357) );
  NAND U1494 ( .A(x[11]), .B(y[19]), .Z(n2834) );
  NANDN U1495 ( .A(n2834), .B(n1289), .Z(n1293) );
  NANDN U1496 ( .A(n1291), .B(n1290), .Z(n1292) );
  NAND U1497 ( .A(n1293), .B(n1292), .Z(n1354) );
  NAND U1498 ( .A(x[16]), .B(y[5]), .Z(n1417) );
  XOR U1499 ( .A(n1416), .B(n1417), .Z(n1419) );
  NAND U1500 ( .A(x[15]), .B(y[6]), .Z(n1418) );
  XOR U1501 ( .A(n1419), .B(n1418), .Z(n1391) );
  AND U1502 ( .A(x[9]), .B(y[5]), .Z(n1294) );
  NAND U1503 ( .A(n2086), .B(n1294), .Z(n1298) );
  OR U1504 ( .A(n1296), .B(n1295), .Z(n1297) );
  NAND U1505 ( .A(n1298), .B(n1297), .Z(n1392) );
  XNOR U1506 ( .A(n1391), .B(n1392), .Z(n1394) );
  IV U1507 ( .A(y[21]), .Z(n2457) );
  ANDN U1508 ( .B(x[0]), .A(n2457), .Z(n1406) );
  AND U1509 ( .A(n1299), .B(o[20]), .Z(n1404) );
  IV U1510 ( .A(x[21]), .Z(n2431) );
  ANDN U1511 ( .B(y[0]), .A(n2431), .Z(n1405) );
  XNOR U1512 ( .A(n1404), .B(n1405), .Z(n1407) );
  XNOR U1513 ( .A(n1406), .B(n1407), .Z(n1393) );
  XOR U1514 ( .A(n1394), .B(n1393), .Z(n1355) );
  XNOR U1515 ( .A(n1357), .B(n1356), .Z(n1361) );
  XNOR U1516 ( .A(n1363), .B(n1362), .Z(n1337) );
  NANDN U1517 ( .A(n1301), .B(n1300), .Z(n1305) );
  NANDN U1518 ( .A(n1303), .B(n1302), .Z(n1304) );
  AND U1519 ( .A(n1305), .B(n1304), .Z(n1336) );
  XOR U1520 ( .A(n1338), .B(n1339), .Z(n1333) );
  XOR U1521 ( .A(n1332), .B(n1333), .Z(n1327) );
  NANDN U1522 ( .A(n1307), .B(n1306), .Z(n1311) );
  OR U1523 ( .A(n1309), .B(n1308), .Z(n1310) );
  NAND U1524 ( .A(n1311), .B(n1310), .Z(n1325) );
  OR U1525 ( .A(n1313), .B(n1312), .Z(n1317) );
  NANDN U1526 ( .A(n1315), .B(n1314), .Z(n1316) );
  NAND U1527 ( .A(n1317), .B(n1316), .Z(n1324) );
  XOR U1528 ( .A(n1325), .B(n1324), .Z(n1326) );
  XOR U1529 ( .A(n1327), .B(n1326), .Z(n1321) );
  XOR U1530 ( .A(n1320), .B(n1321), .Z(N54) );
  NANDN U1531 ( .A(n1319), .B(n1318), .Z(n1323) );
  NANDN U1532 ( .A(n1321), .B(n1320), .Z(n1322) );
  NAND U1533 ( .A(n1323), .B(n1322), .Z(n1449) );
  OR U1534 ( .A(n1325), .B(n1324), .Z(n1329) );
  NANDN U1535 ( .A(n1327), .B(n1326), .Z(n1328) );
  AND U1536 ( .A(n1329), .B(n1328), .Z(n1450) );
  XNOR U1537 ( .A(n1449), .B(n1450), .Z(n1451) );
  NANDN U1538 ( .A(n1331), .B(n1330), .Z(n1335) );
  OR U1539 ( .A(n1333), .B(n1332), .Z(n1334) );
  NAND U1540 ( .A(n1335), .B(n1334), .Z(n1458) );
  NANDN U1541 ( .A(n1337), .B(n1336), .Z(n1341) );
  NANDN U1542 ( .A(n1339), .B(n1338), .Z(n1340) );
  NAND U1543 ( .A(n1341), .B(n1340), .Z(n1455) );
  NANDN U1544 ( .A(n1343), .B(n1342), .Z(n1347) );
  NANDN U1545 ( .A(n1345), .B(n1344), .Z(n1346) );
  NAND U1546 ( .A(n1347), .B(n1346), .Z(n1548) );
  OR U1547 ( .A(n1349), .B(n1348), .Z(n1353) );
  NANDN U1548 ( .A(n1351), .B(n1350), .Z(n1352) );
  NAND U1549 ( .A(n1353), .B(n1352), .Z(n1547) );
  XOR U1550 ( .A(n1548), .B(n1547), .Z(n1549) );
  NANDN U1551 ( .A(n1355), .B(n1354), .Z(n1359) );
  NAND U1552 ( .A(n1357), .B(n1356), .Z(n1358) );
  NAND U1553 ( .A(n1359), .B(n1358), .Z(n1550) );
  XNOR U1554 ( .A(n1549), .B(n1550), .Z(n1461) );
  NANDN U1555 ( .A(n1361), .B(n1360), .Z(n1365) );
  NAND U1556 ( .A(n1363), .B(n1362), .Z(n1364) );
  AND U1557 ( .A(n1365), .B(n1364), .Z(n1462) );
  XNOR U1558 ( .A(n1461), .B(n1462), .Z(n1464) );
  NANDN U1559 ( .A(n1367), .B(n1366), .Z(n1371) );
  OR U1560 ( .A(n1369), .B(n1368), .Z(n1370) );
  NAND U1561 ( .A(n1371), .B(n1370), .Z(n1556) );
  NANDN U1562 ( .A(n1372), .B(n1808), .Z(n1376) );
  OR U1563 ( .A(n1374), .B(n1373), .Z(n1375) );
  AND U1564 ( .A(n1376), .B(n1375), .Z(n1573) );
  OR U1565 ( .A(n1378), .B(n1377), .Z(n1382) );
  OR U1566 ( .A(n1380), .B(n1379), .Z(n1381) );
  NAND U1567 ( .A(n1382), .B(n1381), .Z(n1488) );
  AND U1568 ( .A(x[18]), .B(y[4]), .Z(n1384) );
  NAND U1569 ( .A(y[10]), .B(x[12]), .Z(n1383) );
  XOR U1570 ( .A(n1384), .B(n1383), .Z(n1514) );
  NAND U1571 ( .A(x[4]), .B(y[18]), .Z(n1513) );
  XOR U1572 ( .A(n1514), .B(n1513), .Z(n1485) );
  NAND U1573 ( .A(x[5]), .B(y[17]), .Z(n1530) );
  NAND U1574 ( .A(x[17]), .B(y[5]), .Z(n1529) );
  XOR U1575 ( .A(n1530), .B(n1529), .Z(n1531) );
  NAND U1576 ( .A(x[16]), .B(y[6]), .Z(n1532) );
  XOR U1577 ( .A(n1531), .B(n1532), .Z(n1486) );
  XOR U1578 ( .A(n1488), .B(n1487), .Z(n1571) );
  OR U1579 ( .A(n1386), .B(n1385), .Z(n1390) );
  OR U1580 ( .A(n1388), .B(n1387), .Z(n1389) );
  NAND U1581 ( .A(n1390), .B(n1389), .Z(n1572) );
  XNOR U1582 ( .A(n1571), .B(n1572), .Z(n1574) );
  XOR U1583 ( .A(n1573), .B(n1574), .Z(n1554) );
  OR U1584 ( .A(n1392), .B(n1391), .Z(n1396) );
  OR U1585 ( .A(n1394), .B(n1393), .Z(n1395) );
  NAND U1586 ( .A(n1396), .B(n1395), .Z(n1560) );
  OR U1587 ( .A(n1397), .B(n1506), .Z(n1401) );
  OR U1588 ( .A(n1399), .B(n1398), .Z(n1400) );
  NAND U1589 ( .A(n1401), .B(n1400), .Z(n1470) );
  AND U1590 ( .A(x[8]), .B(y[14]), .Z(n1403) );
  NAND U1591 ( .A(y[15]), .B(x[7]), .Z(n1402) );
  XOR U1592 ( .A(n1403), .B(n1402), .Z(n1509) );
  NAND U1593 ( .A(y[13]), .B(x[9]), .Z(n1508) );
  XOR U1594 ( .A(n1509), .B(n1508), .Z(n1467) );
  NAND U1595 ( .A(x[0]), .B(y[22]), .Z(n1518) );
  NAND U1596 ( .A(y[0]), .B(x[22]), .Z(n1517) );
  XOR U1597 ( .A(n1518), .B(n1517), .Z(n1519) );
  NAND U1598 ( .A(y[1]), .B(x[21]), .Z(n1535) );
  XOR U1599 ( .A(o[22]), .B(n1535), .Z(n1520) );
  XOR U1600 ( .A(n1519), .B(n1520), .Z(n1468) );
  XOR U1601 ( .A(n1470), .B(n1469), .Z(n1482) );
  OR U1602 ( .A(n1405), .B(n1404), .Z(n1409) );
  OR U1603 ( .A(n1407), .B(n1406), .Z(n1408) );
  AND U1604 ( .A(n1409), .B(n1408), .Z(n1479) );
  NANDN U1605 ( .A(n1411), .B(n1410), .Z(n1415) );
  OR U1606 ( .A(n1413), .B(n1412), .Z(n1414) );
  AND U1607 ( .A(n1415), .B(n1414), .Z(n1480) );
  XOR U1608 ( .A(n1479), .B(n1480), .Z(n1481) );
  XOR U1609 ( .A(n1482), .B(n1481), .Z(n1568) );
  NAND U1610 ( .A(x[13]), .B(y[9]), .Z(n1542) );
  NAND U1611 ( .A(x[2]), .B(y[20]), .Z(n1541) );
  XOR U1612 ( .A(n1542), .B(n1541), .Z(n1543) );
  NAND U1613 ( .A(y[2]), .B(x[20]), .Z(n1544) );
  XOR U1614 ( .A(n1543), .B(n1544), .Z(n1526) );
  NANDN U1615 ( .A(n1417), .B(n1416), .Z(n1421) );
  OR U1616 ( .A(n1419), .B(n1418), .Z(n1420) );
  AND U1617 ( .A(n1421), .B(n1420), .Z(n1524) );
  AND U1618 ( .A(x[10]), .B(y[12]), .Z(n1423) );
  NAND U1619 ( .A(x[6]), .B(y[16]), .Z(n1422) );
  XOR U1620 ( .A(n1423), .B(n1422), .Z(n1538) );
  NAND U1621 ( .A(x[15]), .B(y[7]), .Z(n1537) );
  XNOR U1622 ( .A(n1538), .B(n1537), .Z(n1523) );
  XOR U1623 ( .A(n1524), .B(n1523), .Z(n1525) );
  XNOR U1624 ( .A(n1526), .B(n1525), .Z(n1565) );
  OR U1625 ( .A(n1425), .B(n1424), .Z(n1429) );
  OR U1626 ( .A(n1427), .B(n1426), .Z(n1428) );
  NAND U1627 ( .A(n1429), .B(n1428), .Z(n1476) );
  NAND U1628 ( .A(y[8]), .B(x[14]), .Z(n1499) );
  NAND U1629 ( .A(y[19]), .B(x[3]), .Z(n1498) );
  XOR U1630 ( .A(n1499), .B(n1498), .Z(n1500) );
  NAND U1631 ( .A(y[3]), .B(x[19]), .Z(n1501) );
  XOR U1632 ( .A(n1500), .B(n1501), .Z(n1474) );
  NANDN U1633 ( .A(n1430), .B(o[21]), .Z(n1495) );
  NAND U1634 ( .A(x[1]), .B(y[21]), .Z(n1493) );
  XOR U1635 ( .A(n1492), .B(n1493), .Z(n1494) );
  XOR U1636 ( .A(n1495), .B(n1494), .Z(n1473) );
  XNOR U1637 ( .A(n1476), .B(n1475), .Z(n1566) );
  XNOR U1638 ( .A(n1568), .B(n1567), .Z(n1559) );
  XNOR U1639 ( .A(n1560), .B(n1559), .Z(n1562) );
  OR U1640 ( .A(n1432), .B(n1431), .Z(n1436) );
  OR U1641 ( .A(n1434), .B(n1433), .Z(n1435) );
  NAND U1642 ( .A(n1436), .B(n1435), .Z(n1561) );
  XOR U1643 ( .A(n1562), .B(n1561), .Z(n1553) );
  XOR U1644 ( .A(n1554), .B(n1553), .Z(n1555) );
  XNOR U1645 ( .A(n1556), .B(n1555), .Z(n1463) );
  XNOR U1646 ( .A(n1464), .B(n1463), .Z(n1580) );
  NANDN U1647 ( .A(n1438), .B(n1437), .Z(n1442) );
  NANDN U1648 ( .A(n1440), .B(n1439), .Z(n1441) );
  NAND U1649 ( .A(n1442), .B(n1441), .Z(n1578) );
  OR U1650 ( .A(n1444), .B(n1443), .Z(n1448) );
  NANDN U1651 ( .A(n1446), .B(n1445), .Z(n1447) );
  NAND U1652 ( .A(n1448), .B(n1447), .Z(n1577) );
  XNOR U1653 ( .A(n1578), .B(n1577), .Z(n1579) );
  XNOR U1654 ( .A(n1580), .B(n1579), .Z(n1456) );
  XOR U1655 ( .A(n1458), .B(n1457), .Z(n1452) );
  XOR U1656 ( .A(n1451), .B(n1452), .Z(N55) );
  NANDN U1657 ( .A(n1450), .B(n1449), .Z(n1454) );
  NANDN U1658 ( .A(n1452), .B(n1451), .Z(n1453) );
  NAND U1659 ( .A(n1454), .B(n1453), .Z(n1583) );
  NANDN U1660 ( .A(n1456), .B(n1455), .Z(n1460) );
  NAND U1661 ( .A(n1458), .B(n1457), .Z(n1459) );
  NAND U1662 ( .A(n1460), .B(n1459), .Z(n1584) );
  XNOR U1663 ( .A(n1583), .B(n1584), .Z(n1585) );
  OR U1664 ( .A(n1462), .B(n1461), .Z(n1466) );
  OR U1665 ( .A(n1464), .B(n1463), .Z(n1465) );
  NAND U1666 ( .A(n1466), .B(n1465), .Z(n1590) );
  NANDN U1667 ( .A(n1468), .B(n1467), .Z(n1472) );
  OR U1668 ( .A(n1470), .B(n1469), .Z(n1471) );
  AND U1669 ( .A(n1472), .B(n1471), .Z(n1663) );
  NANDN U1670 ( .A(n1474), .B(n1473), .Z(n1478) );
  OR U1671 ( .A(n1476), .B(n1475), .Z(n1477) );
  AND U1672 ( .A(n1478), .B(n1477), .Z(n1664) );
  XOR U1673 ( .A(n1663), .B(n1664), .Z(n1665) );
  OR U1674 ( .A(n1480), .B(n1479), .Z(n1484) );
  NANDN U1675 ( .A(n1482), .B(n1481), .Z(n1483) );
  NAND U1676 ( .A(n1484), .B(n1483), .Z(n1666) );
  NANDN U1677 ( .A(n1486), .B(n1485), .Z(n1490) );
  OR U1678 ( .A(n1488), .B(n1487), .Z(n1489) );
  AND U1679 ( .A(n1490), .B(n1489), .Z(n1596) );
  XOR U1680 ( .A(n1491), .B(n1507), .Z(n1648) );
  NAND U1681 ( .A(y[16]), .B(x[7]), .Z(n1647) );
  XOR U1682 ( .A(n1648), .B(n1647), .Z(n1669) );
  NAND U1683 ( .A(y[13]), .B(x[10]), .Z(n1670) );
  XOR U1684 ( .A(n1669), .B(n1670), .Z(n1672) );
  NAND U1685 ( .A(x[6]), .B(y[17]), .Z(n1640) );
  NAND U1686 ( .A(x[15]), .B(y[8]), .Z(n1639) );
  XOR U1687 ( .A(n1640), .B(n1639), .Z(n1641) );
  NAND U1688 ( .A(x[11]), .B(y[12]), .Z(n1642) );
  XNOR U1689 ( .A(n1641), .B(n1642), .Z(n1671) );
  XNOR U1690 ( .A(n1672), .B(n1671), .Z(n1696) );
  NANDN U1691 ( .A(n1493), .B(n1492), .Z(n1497) );
  OR U1692 ( .A(n1495), .B(n1494), .Z(n1496) );
  NAND U1693 ( .A(n1497), .B(n1496), .Z(n1694) );
  OR U1694 ( .A(n1499), .B(n1498), .Z(n1503) );
  NANDN U1695 ( .A(n1501), .B(n1500), .Z(n1502) );
  AND U1696 ( .A(n1503), .B(n1502), .Z(n1693) );
  XOR U1697 ( .A(n1596), .B(n1595), .Z(n1597) );
  XOR U1698 ( .A(n1598), .B(n1597), .Z(n1608) );
  NAND U1699 ( .A(y[23]), .B(x[0]), .Z(n1628) );
  NAND U1700 ( .A(y[0]), .B(x[23]), .Z(n1627) );
  XOR U1701 ( .A(n1628), .B(n1627), .Z(n1629) );
  NAND U1702 ( .A(y[1]), .B(x[22]), .Z(n1656) );
  XOR U1703 ( .A(o[23]), .B(n1656), .Z(n1630) );
  XNOR U1704 ( .A(n1629), .B(n1630), .Z(n1707) );
  NAND U1705 ( .A(x[20]), .B(y[3]), .Z(n1504) );
  XOR U1706 ( .A(n1505), .B(n1504), .Z(n1653) );
  NAND U1707 ( .A(y[4]), .B(x[19]), .Z(n1652) );
  XOR U1708 ( .A(n1653), .B(n1652), .Z(n1705) );
  NANDN U1709 ( .A(n1507), .B(n1506), .Z(n1511) );
  OR U1710 ( .A(n1509), .B(n1508), .Z(n1510) );
  NAND U1711 ( .A(n1511), .B(n1510), .Z(n1706) );
  XNOR U1712 ( .A(n1705), .B(n1706), .Z(n1708) );
  XNOR U1713 ( .A(n1707), .B(n1708), .Z(n1713) );
  ANDN U1714 ( .B(x[18]), .A(n2500), .Z(n2485) );
  NAND U1715 ( .A(n1512), .B(n2485), .Z(n1516) );
  OR U1716 ( .A(n1514), .B(n1513), .Z(n1515) );
  AND U1717 ( .A(n1516), .B(n1515), .Z(n1712) );
  OR U1718 ( .A(n1518), .B(n1517), .Z(n1522) );
  NANDN U1719 ( .A(n1520), .B(n1519), .Z(n1521) );
  AND U1720 ( .A(n1522), .B(n1521), .Z(n1711) );
  XNOR U1721 ( .A(n1712), .B(n1711), .Z(n1714) );
  XOR U1722 ( .A(n1713), .B(n1714), .Z(n1619) );
  OR U1723 ( .A(n1524), .B(n1523), .Z(n1528) );
  NANDN U1724 ( .A(n1526), .B(n1525), .Z(n1527) );
  NAND U1725 ( .A(n1528), .B(n1527), .Z(n1620) );
  XOR U1726 ( .A(n1619), .B(n1620), .Z(n1622) );
  NAND U1727 ( .A(x[13]), .B(y[10]), .Z(n1682) );
  NAND U1728 ( .A(x[2]), .B(y[21]), .Z(n1681) );
  XOR U1729 ( .A(n1682), .B(n1681), .Z(n1683) );
  NAND U1730 ( .A(y[2]), .B(x[21]), .Z(n1684) );
  XOR U1731 ( .A(n1683), .B(n1684), .Z(n1720) );
  OR U1732 ( .A(n1530), .B(n1529), .Z(n1534) );
  NANDN U1733 ( .A(n1532), .B(n1531), .Z(n1533) );
  AND U1734 ( .A(n1534), .B(n1533), .Z(n1717) );
  NANDN U1735 ( .A(n1535), .B(o[22]), .Z(n1636) );
  NAND U1736 ( .A(y[11]), .B(x[12]), .Z(n1634) );
  NAND U1737 ( .A(x[1]), .B(y[22]), .Z(n1633) );
  XOR U1738 ( .A(n1634), .B(n1633), .Z(n1635) );
  XOR U1739 ( .A(n1636), .B(n1635), .Z(n1718) );
  XNOR U1740 ( .A(n1717), .B(n1718), .Z(n1719) );
  XOR U1741 ( .A(n1720), .B(n1719), .Z(n1660) );
  ANDN U1742 ( .B(y[16]), .A(n2455), .Z(n2052) );
  NAND U1743 ( .A(n1536), .B(n2052), .Z(n1540) );
  OR U1744 ( .A(n1538), .B(n1537), .Z(n1539) );
  AND U1745 ( .A(n1540), .B(n1539), .Z(n1699) );
  NAND U1746 ( .A(x[5]), .B(y[18]), .Z(n1688) );
  NAND U1747 ( .A(y[5]), .B(x[18]), .Z(n1687) );
  XOR U1748 ( .A(n1688), .B(n1687), .Z(n1689) );
  NAND U1749 ( .A(y[6]), .B(x[17]), .Z(n1690) );
  XOR U1750 ( .A(n1689), .B(n1690), .Z(n1700) );
  XNOR U1751 ( .A(n1699), .B(n1700), .Z(n1702) );
  NAND U1752 ( .A(y[9]), .B(x[14]), .Z(n1676) );
  NAND U1753 ( .A(y[20]), .B(x[3]), .Z(n1675) );
  XOR U1754 ( .A(n1676), .B(n1675), .Z(n1677) );
  NAND U1755 ( .A(y[19]), .B(x[4]), .Z(n1678) );
  XOR U1756 ( .A(n1677), .B(n1678), .Z(n1701) );
  XOR U1757 ( .A(n1702), .B(n1701), .Z(n1657) );
  OR U1758 ( .A(n1542), .B(n1541), .Z(n1546) );
  NANDN U1759 ( .A(n1544), .B(n1543), .Z(n1545) );
  NAND U1760 ( .A(n1546), .B(n1545), .Z(n1658) );
  XOR U1761 ( .A(n1657), .B(n1658), .Z(n1659) );
  XNOR U1762 ( .A(n1660), .B(n1659), .Z(n1621) );
  XNOR U1763 ( .A(n1622), .B(n1621), .Z(n1607) );
  XOR U1764 ( .A(n1608), .B(n1607), .Z(n1610) );
  OR U1765 ( .A(n1548), .B(n1547), .Z(n1552) );
  NANDN U1766 ( .A(n1550), .B(n1549), .Z(n1551) );
  AND U1767 ( .A(n1552), .B(n1551), .Z(n1609) );
  XOR U1768 ( .A(n1610), .B(n1609), .Z(n1615) );
  NANDN U1769 ( .A(n1554), .B(n1553), .Z(n1558) );
  OR U1770 ( .A(n1556), .B(n1555), .Z(n1557) );
  NAND U1771 ( .A(n1558), .B(n1557), .Z(n1614) );
  OR U1772 ( .A(n1560), .B(n1559), .Z(n1564) );
  OR U1773 ( .A(n1562), .B(n1561), .Z(n1563) );
  NAND U1774 ( .A(n1564), .B(n1563), .Z(n1604) );
  NANDN U1775 ( .A(n1566), .B(n1565), .Z(n1570) );
  NAND U1776 ( .A(n1568), .B(n1567), .Z(n1569) );
  NAND U1777 ( .A(n1570), .B(n1569), .Z(n1602) );
  OR U1778 ( .A(n1572), .B(n1571), .Z(n1576) );
  OR U1779 ( .A(n1574), .B(n1573), .Z(n1575) );
  AND U1780 ( .A(n1576), .B(n1575), .Z(n1601) );
  XOR U1781 ( .A(n1602), .B(n1601), .Z(n1603) );
  XOR U1782 ( .A(n1614), .B(n1613), .Z(n1616) );
  XOR U1783 ( .A(n1590), .B(n1589), .Z(n1592) );
  OR U1784 ( .A(n1578), .B(n1577), .Z(n1582) );
  OR U1785 ( .A(n1580), .B(n1579), .Z(n1581) );
  NAND U1786 ( .A(n1582), .B(n1581), .Z(n1591) );
  XOR U1787 ( .A(n1592), .B(n1591), .Z(n1586) );
  XNOR U1788 ( .A(n1585), .B(n1586), .Z(N56) );
  NANDN U1789 ( .A(n1584), .B(n1583), .Z(n1588) );
  NAND U1790 ( .A(n1586), .B(n1585), .Z(n1587) );
  NAND U1791 ( .A(n1588), .B(n1587), .Z(n1723) );
  NANDN U1792 ( .A(n1590), .B(n1589), .Z(n1594) );
  OR U1793 ( .A(n1592), .B(n1591), .Z(n1593) );
  AND U1794 ( .A(n1594), .B(n1593), .Z(n1724) );
  XNOR U1795 ( .A(n1723), .B(n1724), .Z(n1725) );
  NANDN U1796 ( .A(n1596), .B(n1595), .Z(n1600) );
  OR U1797 ( .A(n1598), .B(n1597), .Z(n1599) );
  NAND U1798 ( .A(n1600), .B(n1599), .Z(n1863) );
  OR U1799 ( .A(n1602), .B(n1601), .Z(n1606) );
  NANDN U1800 ( .A(n1604), .B(n1603), .Z(n1605) );
  AND U1801 ( .A(n1606), .B(n1605), .Z(n1862) );
  XOR U1802 ( .A(n1863), .B(n1862), .Z(n1864) );
  NANDN U1803 ( .A(n1608), .B(n1607), .Z(n1612) );
  OR U1804 ( .A(n1610), .B(n1609), .Z(n1611) );
  AND U1805 ( .A(n1612), .B(n1611), .Z(n1865) );
  NANDN U1806 ( .A(n1614), .B(n1613), .Z(n1618) );
  NANDN U1807 ( .A(n1616), .B(n1615), .Z(n1617) );
  AND U1808 ( .A(n1618), .B(n1617), .Z(n1730) );
  NANDN U1809 ( .A(n1620), .B(n1619), .Z(n1624) );
  NANDN U1810 ( .A(n1622), .B(n1621), .Z(n1623) );
  NAND U1811 ( .A(n1624), .B(n1623), .Z(n1853) );
  NAND U1812 ( .A(y[10]), .B(x[14]), .Z(n1810) );
  AND U1813 ( .A(y[13]), .B(x[11]), .Z(n1626) );
  NAND U1814 ( .A(x[8]), .B(y[16]), .Z(n1625) );
  XOR U1815 ( .A(n1626), .B(n1625), .Z(n1809) );
  XNOR U1816 ( .A(n1810), .B(n1809), .Z(n1805) );
  NOR U1817 ( .A(n2452), .B(n2048), .Z(n1646) );
  IV U1818 ( .A(n1646), .Z(n1802) );
  ANDN U1819 ( .B(y[14]), .A(n2455), .Z(n1803) );
  XNOR U1820 ( .A(n1802), .B(n1803), .Z(n1804) );
  XOR U1821 ( .A(n1805), .B(n1804), .Z(n1846) );
  OR U1822 ( .A(n1628), .B(n1627), .Z(n1632) );
  NANDN U1823 ( .A(n1630), .B(n1629), .Z(n1631) );
  NAND U1824 ( .A(n1632), .B(n1631), .Z(n1844) );
  NAND U1825 ( .A(x[4]), .B(y[20]), .Z(n1841) );
  NAND U1826 ( .A(x[3]), .B(y[21]), .Z(n1839) );
  XOR U1827 ( .A(n1838), .B(n1839), .Z(n1840) );
  XNOR U1828 ( .A(n1841), .B(n1840), .Z(n1845) );
  XOR U1829 ( .A(n1844), .B(n1845), .Z(n1847) );
  XOR U1830 ( .A(n1846), .B(n1847), .Z(n1798) );
  OR U1831 ( .A(n1634), .B(n1633), .Z(n1638) );
  NANDN U1832 ( .A(n1636), .B(n1635), .Z(n1637) );
  NAND U1833 ( .A(n1638), .B(n1637), .Z(n1768) );
  NAND U1834 ( .A(x[21]), .B(y[3]), .Z(n1761) );
  NAND U1835 ( .A(x[5]), .B(y[19]), .Z(n1759) );
  NAND U1836 ( .A(x[16]), .B(y[8]), .Z(n1758) );
  XOR U1837 ( .A(n1759), .B(n1758), .Z(n1760) );
  XOR U1838 ( .A(n1761), .B(n1760), .Z(n1744) );
  OR U1839 ( .A(n1640), .B(n1639), .Z(n1644) );
  NANDN U1840 ( .A(n1642), .B(n1641), .Z(n1643) );
  AND U1841 ( .A(n1644), .B(n1643), .Z(n1741) );
  NAND U1842 ( .A(y[5]), .B(x[19]), .Z(n1755) );
  AND U1843 ( .A(y[4]), .B(x[20]), .Z(n1940) );
  NAND U1844 ( .A(x[6]), .B(y[18]), .Z(n1753) );
  XOR U1845 ( .A(n1940), .B(n1753), .Z(n1754) );
  XNOR U1846 ( .A(n1755), .B(n1754), .Z(n1742) );
  XNOR U1847 ( .A(n1741), .B(n1742), .Z(n1743) );
  XNOR U1848 ( .A(n1744), .B(n1743), .Z(n1767) );
  NAND U1849 ( .A(n1646), .B(n1645), .Z(n1650) );
  OR U1850 ( .A(n1648), .B(n1647), .Z(n1649) );
  NAND U1851 ( .A(n1650), .B(n1649), .Z(n1766) );
  NAND U1852 ( .A(x[2]), .B(y[22]), .Z(n1820) );
  XOR U1853 ( .A(n1819), .B(n1820), .Z(n1822) );
  NAND U1854 ( .A(y[2]), .B(x[22]), .Z(n1821) );
  XOR U1855 ( .A(n1822), .B(n1821), .Z(n1737) );
  IV U1856 ( .A(x[20]), .Z(n2432) );
  ANDN U1857 ( .B(y[7]), .A(n2432), .Z(n2247) );
  NAND U1858 ( .A(n1651), .B(n2247), .Z(n1655) );
  OR U1859 ( .A(n1653), .B(n1652), .Z(n1654) );
  NAND U1860 ( .A(n1655), .B(n1654), .Z(n1736) );
  NANDN U1861 ( .A(n1656), .B(o[23]), .Z(n1816) );
  NAND U1862 ( .A(x[1]), .B(y[23]), .Z(n1814) );
  XOR U1863 ( .A(n1813), .B(n1814), .Z(n1815) );
  XOR U1864 ( .A(n1816), .B(n1815), .Z(n1735) );
  XNOR U1865 ( .A(n1736), .B(n1735), .Z(n1738) );
  XNOR U1866 ( .A(n1737), .B(n1738), .Z(n1797) );
  XOR U1867 ( .A(n1796), .B(n1797), .Z(n1799) );
  XOR U1868 ( .A(n1798), .B(n1799), .Z(n1850) );
  OR U1869 ( .A(n1658), .B(n1657), .Z(n1662) );
  NANDN U1870 ( .A(n1660), .B(n1659), .Z(n1661) );
  NAND U1871 ( .A(n1662), .B(n1661), .Z(n1851) );
  XOR U1872 ( .A(n1850), .B(n1851), .Z(n1852) );
  XOR U1873 ( .A(n1853), .B(n1852), .Z(n1858) );
  OR U1874 ( .A(n1664), .B(n1663), .Z(n1668) );
  NANDN U1875 ( .A(n1666), .B(n1665), .Z(n1667) );
  NAND U1876 ( .A(n1668), .B(n1667), .Z(n1857) );
  NANDN U1877 ( .A(n1670), .B(n1669), .Z(n1674) );
  NANDN U1878 ( .A(n1672), .B(n1671), .Z(n1673) );
  NAND U1879 ( .A(n1674), .B(n1673), .Z(n1790) );
  OR U1880 ( .A(n1676), .B(n1675), .Z(n1680) );
  NANDN U1881 ( .A(n1678), .B(n1677), .Z(n1679) );
  NAND U1882 ( .A(n1680), .B(n1679), .Z(n1772) );
  OR U1883 ( .A(n1682), .B(n1681), .Z(n1686) );
  NANDN U1884 ( .A(n1684), .B(n1683), .Z(n1685) );
  AND U1885 ( .A(n1686), .B(n1685), .Z(n1773) );
  NAND U1886 ( .A(x[7]), .B(y[17]), .Z(n1827) );
  NAND U1887 ( .A(x[17]), .B(y[7]), .Z(n1826) );
  XOR U1888 ( .A(n1827), .B(n1826), .Z(n1828) );
  NAND U1889 ( .A(y[6]), .B(x[18]), .Z(n1829) );
  XOR U1890 ( .A(n1828), .B(n1829), .Z(n1747) );
  NAND U1891 ( .A(x[0]), .B(y[24]), .Z(n1833) );
  AND U1892 ( .A(y[0]), .B(x[24]), .Z(n1832) );
  XNOR U1893 ( .A(n1833), .B(n1832), .Z(n1834) );
  NAND U1894 ( .A(y[1]), .B(x[23]), .Z(n1825) );
  XOR U1895 ( .A(o[24]), .B(n1825), .Z(n1835) );
  XNOR U1896 ( .A(n1834), .B(n1835), .Z(n1748) );
  OR U1897 ( .A(n1688), .B(n1687), .Z(n1692) );
  NANDN U1898 ( .A(n1690), .B(n1689), .Z(n1691) );
  NAND U1899 ( .A(n1692), .B(n1691), .Z(n1750) );
  XOR U1900 ( .A(n1749), .B(n1750), .Z(n1775) );
  XNOR U1901 ( .A(n1774), .B(n1775), .Z(n1791) );
  NANDN U1902 ( .A(n1694), .B(n1693), .Z(n1698) );
  NANDN U1903 ( .A(n1696), .B(n1695), .Z(n1697) );
  AND U1904 ( .A(n1698), .B(n1697), .Z(n1793) );
  XNOR U1905 ( .A(n1792), .B(n1793), .Z(n1787) );
  OR U1906 ( .A(n1700), .B(n1699), .Z(n1704) );
  OR U1907 ( .A(n1702), .B(n1701), .Z(n1703) );
  NAND U1908 ( .A(n1704), .B(n1703), .Z(n1781) );
  OR U1909 ( .A(n1706), .B(n1705), .Z(n1710) );
  OR U1910 ( .A(n1708), .B(n1707), .Z(n1709) );
  NAND U1911 ( .A(n1710), .B(n1709), .Z(n1778) );
  OR U1912 ( .A(n1712), .B(n1711), .Z(n1716) );
  NANDN U1913 ( .A(n1714), .B(n1713), .Z(n1715) );
  NAND U1914 ( .A(n1716), .B(n1715), .Z(n1779) );
  XOR U1915 ( .A(n1781), .B(n1780), .Z(n1784) );
  OR U1916 ( .A(n1718), .B(n1717), .Z(n1722) );
  OR U1917 ( .A(n1720), .B(n1719), .Z(n1721) );
  AND U1918 ( .A(n1722), .B(n1721), .Z(n1785) );
  XNOR U1919 ( .A(n1787), .B(n1786), .Z(n1856) );
  XNOR U1920 ( .A(n1857), .B(n1856), .Z(n1859) );
  XNOR U1921 ( .A(n1858), .B(n1859), .Z(n1729) );
  XOR U1922 ( .A(n1730), .B(n1729), .Z(n1731) );
  XNOR U1923 ( .A(n1732), .B(n1731), .Z(n1726) );
  XOR U1924 ( .A(n1725), .B(n1726), .Z(N57) );
  NANDN U1925 ( .A(n1724), .B(n1723), .Z(n1728) );
  NANDN U1926 ( .A(n1726), .B(n1725), .Z(n1727) );
  NAND U1927 ( .A(n1728), .B(n1727), .Z(n1868) );
  NANDN U1928 ( .A(n1730), .B(n1729), .Z(n1734) );
  OR U1929 ( .A(n1732), .B(n1731), .Z(n1733) );
  AND U1930 ( .A(n1734), .B(n1733), .Z(n1869) );
  XNOR U1931 ( .A(n1868), .B(n1869), .Z(n1870) );
  NAND U1932 ( .A(n1736), .B(n1735), .Z(n1740) );
  NANDN U1933 ( .A(n1738), .B(n1737), .Z(n1739) );
  AND U1934 ( .A(n1740), .B(n1739), .Z(n2002) );
  OR U1935 ( .A(n1742), .B(n1741), .Z(n1746) );
  OR U1936 ( .A(n1744), .B(n1743), .Z(n1745) );
  AND U1937 ( .A(n1746), .B(n1745), .Z(n2000) );
  NANDN U1938 ( .A(n1748), .B(n1747), .Z(n1752) );
  NANDN U1939 ( .A(n1750), .B(n1749), .Z(n1751) );
  NAND U1940 ( .A(n1752), .B(n1751), .Z(n1925) );
  ANDN U1941 ( .B(x[23]), .A(n19), .Z(n1960) );
  ANDN U1942 ( .B(x[4]), .A(n2457), .Z(n1958) );
  ANDN U1943 ( .B(x[16]), .A(n2314), .Z(n1959) );
  XNOR U1944 ( .A(n1958), .B(n1959), .Z(n1961) );
  XOR U1945 ( .A(n1960), .B(n1961), .Z(n1984) );
  ANDN U1946 ( .B(x[15]), .A(n2500), .Z(n1936) );
  ANDN U1947 ( .B(x[18]), .A(n2433), .Z(n1934) );
  ANDN U1948 ( .B(y[19]), .A(n2313), .Z(n1935) );
  XNOR U1949 ( .A(n1934), .B(n1935), .Z(n1937) );
  XOR U1950 ( .A(n1936), .B(n1937), .Z(n1982) );
  NANDN U1951 ( .A(n1753), .B(n1940), .Z(n1757) );
  OR U1952 ( .A(n1755), .B(n1754), .Z(n1756) );
  AND U1953 ( .A(n1757), .B(n1756), .Z(n1983) );
  XNOR U1954 ( .A(n1982), .B(n1983), .Z(n1985) );
  XNOR U1955 ( .A(n1984), .B(n1985), .Z(n1923) );
  OR U1956 ( .A(n1759), .B(n1758), .Z(n1763) );
  NANDN U1957 ( .A(n1761), .B(n1760), .Z(n1762) );
  AND U1958 ( .A(n1763), .B(n1762), .Z(n1990) );
  ANDN U1959 ( .B(x[22]), .A(n20), .Z(n1954) );
  ANDN U1960 ( .B(y[20]), .A(n2252), .Z(n1952) );
  ANDN U1961 ( .B(x[17]), .A(n2430), .Z(n1953) );
  XNOR U1962 ( .A(n1952), .B(n1953), .Z(n1955) );
  XOR U1963 ( .A(n1954), .B(n1955), .Z(n1989) );
  NAND U1964 ( .A(y[6]), .B(x[19]), .Z(n1942) );
  AND U1965 ( .A(x[21]), .B(y[4]), .Z(n1765) );
  AND U1966 ( .A(x[20]), .B(y[5]), .Z(n1764) );
  XNOR U1967 ( .A(n1765), .B(n1764), .Z(n1941) );
  XOR U1968 ( .A(n1942), .B(n1941), .Z(n1988) );
  XOR U1969 ( .A(n1989), .B(n1988), .Z(n1991) );
  XOR U1970 ( .A(n1990), .B(n1991), .Z(n1922) );
  XNOR U1971 ( .A(n1923), .B(n1922), .Z(n1924) );
  XOR U1972 ( .A(n1925), .B(n1924), .Z(n2001) );
  XNOR U1973 ( .A(n2000), .B(n2001), .Z(n2003) );
  XNOR U1974 ( .A(n2002), .B(n2003), .Z(n1931) );
  NANDN U1975 ( .A(n1767), .B(n1766), .Z(n1771) );
  NANDN U1976 ( .A(n1769), .B(n1768), .Z(n1770) );
  NAND U1977 ( .A(n1771), .B(n1770), .Z(n1929) );
  NANDN U1978 ( .A(n1773), .B(n1772), .Z(n1777) );
  NAND U1979 ( .A(n1775), .B(n1774), .Z(n1776) );
  AND U1980 ( .A(n1777), .B(n1776), .Z(n1928) );
  XNOR U1981 ( .A(n1931), .B(n1930), .Z(n1881) );
  NANDN U1982 ( .A(n1779), .B(n1778), .Z(n1783) );
  NANDN U1983 ( .A(n1781), .B(n1780), .Z(n1782) );
  AND U1984 ( .A(n1783), .B(n1782), .Z(n1880) );
  XOR U1985 ( .A(n1881), .B(n1880), .Z(n1882) );
  NANDN U1986 ( .A(n1785), .B(n1784), .Z(n1789) );
  NANDN U1987 ( .A(n1787), .B(n1786), .Z(n1788) );
  NAND U1988 ( .A(n1789), .B(n1788), .Z(n1883) );
  XNOR U1989 ( .A(n1882), .B(n1883), .Z(n1889) );
  NANDN U1990 ( .A(n1791), .B(n1790), .Z(n1795) );
  NAND U1991 ( .A(n1793), .B(n1792), .Z(n1794) );
  NAND U1992 ( .A(n1795), .B(n1794), .Z(n2015) );
  NANDN U1993 ( .A(n1797), .B(n1796), .Z(n1801) );
  OR U1994 ( .A(n1799), .B(n1798), .Z(n1800) );
  NAND U1995 ( .A(n1801), .B(n1800), .Z(n2012) );
  NANDN U1996 ( .A(n1803), .B(n1802), .Z(n1807) );
  NAND U1997 ( .A(n1805), .B(n1804), .Z(n1806) );
  NAND U1998 ( .A(n1807), .B(n1806), .Z(n1917) );
  NANDN U1999 ( .A(n1808), .B(n2303), .Z(n1812) );
  OR U2000 ( .A(n1810), .B(n1809), .Z(n1811) );
  AND U2001 ( .A(n1812), .B(n1811), .Z(n1978) );
  NAND U2002 ( .A(x[1]), .B(y[24]), .Z(n1971) );
  AND U2003 ( .A(x[13]), .B(y[12]), .Z(n1970) );
  XNOR U2004 ( .A(n1971), .B(n1970), .Z(n1973) );
  NAND U2005 ( .A(y[1]), .B(x[24]), .Z(n1945) );
  XNOR U2006 ( .A(n1945), .B(o[25]), .Z(n1972) );
  XNOR U2007 ( .A(n1973), .B(n1972), .Z(n1977) );
  ANDN U2008 ( .B(x[11]), .A(n2429), .Z(n1948) );
  ANDN U2009 ( .B(y[18]), .A(n28), .Z(n1947) );
  XNOR U2010 ( .A(n1946), .B(n1947), .Z(n1949) );
  XOR U2011 ( .A(n1948), .B(n1949), .Z(n1976) );
  XNOR U2012 ( .A(n1977), .B(n1976), .Z(n1979) );
  XOR U2013 ( .A(n1978), .B(n1979), .Z(n1916) );
  XNOR U2014 ( .A(n1917), .B(n1916), .Z(n1918) );
  NANDN U2015 ( .A(n1814), .B(n1813), .Z(n1818) );
  OR U2016 ( .A(n1816), .B(n1815), .Z(n1817) );
  NAND U2017 ( .A(n1818), .B(n1817), .Z(n1913) );
  NANDN U2018 ( .A(n1820), .B(n1819), .Z(n1824) );
  OR U2019 ( .A(n1822), .B(n1821), .Z(n1823) );
  NAND U2020 ( .A(n1824), .B(n1823), .Z(n1910) );
  NAND U2021 ( .A(x[8]), .B(y[17]), .Z(n1906) );
  XNOR U2022 ( .A(n1905), .B(n1904), .Z(n1907) );
  XOR U2023 ( .A(n1906), .B(n1907), .Z(n1892) );
  NANDN U2024 ( .A(n1825), .B(o[24]), .Z(n1900) );
  IV U2025 ( .A(x[25]), .Z(n2484) );
  ANDN U2026 ( .B(y[0]), .A(n2484), .Z(n1899) );
  NAND U2027 ( .A(x[0]), .B(y[25]), .Z(n1898) );
  XOR U2028 ( .A(n1899), .B(n1898), .Z(n1901) );
  XNOR U2029 ( .A(n1900), .B(n1901), .Z(n1893) );
  XOR U2030 ( .A(n1892), .B(n1893), .Z(n1895) );
  OR U2031 ( .A(n1827), .B(n1826), .Z(n1831) );
  NANDN U2032 ( .A(n1829), .B(n1828), .Z(n1830) );
  NAND U2033 ( .A(n1831), .B(n1830), .Z(n1894) );
  XOR U2034 ( .A(n1895), .B(n1894), .Z(n1911) );
  XNOR U2035 ( .A(n1913), .B(n1912), .Z(n1919) );
  XOR U2036 ( .A(n1918), .B(n1919), .Z(n2009) );
  NAND U2037 ( .A(y[23]), .B(x[2]), .Z(n1967) );
  NAND U2038 ( .A(x[3]), .B(y[22]), .Z(n1965) );
  XOR U2039 ( .A(n1964), .B(n1965), .Z(n1966) );
  XOR U2040 ( .A(n1967), .B(n1966), .Z(n1994) );
  NANDN U2041 ( .A(n1833), .B(n1832), .Z(n1837) );
  NANDN U2042 ( .A(n1835), .B(n1834), .Z(n1836) );
  NAND U2043 ( .A(n1837), .B(n1836), .Z(n1995) );
  XNOR U2044 ( .A(n1994), .B(n1995), .Z(n1997) );
  NANDN U2045 ( .A(n1839), .B(n1838), .Z(n1843) );
  OR U2046 ( .A(n1841), .B(n1840), .Z(n1842) );
  AND U2047 ( .A(n1843), .B(n1842), .Z(n1996) );
  XNOR U2048 ( .A(n1997), .B(n1996), .Z(n2006) );
  NANDN U2049 ( .A(n1845), .B(n1844), .Z(n1849) );
  OR U2050 ( .A(n1847), .B(n1846), .Z(n1848) );
  NAND U2051 ( .A(n1849), .B(n1848), .Z(n2007) );
  XNOR U2052 ( .A(n2009), .B(n2008), .Z(n2013) );
  XOR U2053 ( .A(n2015), .B(n2014), .Z(n1886) );
  OR U2054 ( .A(n1851), .B(n1850), .Z(n1855) );
  NANDN U2055 ( .A(n1853), .B(n1852), .Z(n1854) );
  AND U2056 ( .A(n1855), .B(n1854), .Z(n1887) );
  XNOR U2057 ( .A(n1889), .B(n1888), .Z(n1874) );
  OR U2058 ( .A(n1857), .B(n1856), .Z(n1861) );
  NANDN U2059 ( .A(n1859), .B(n1858), .Z(n1860) );
  AND U2060 ( .A(n1861), .B(n1860), .Z(n1875) );
  XNOR U2061 ( .A(n1874), .B(n1875), .Z(n1877) );
  OR U2062 ( .A(n1863), .B(n1862), .Z(n1867) );
  NANDN U2063 ( .A(n1865), .B(n1864), .Z(n1866) );
  AND U2064 ( .A(n1867), .B(n1866), .Z(n1876) );
  XOR U2065 ( .A(n1877), .B(n1876), .Z(n1871) );
  XNOR U2066 ( .A(n1870), .B(n1871), .Z(N58) );
  NANDN U2067 ( .A(n1869), .B(n1868), .Z(n1873) );
  NAND U2068 ( .A(n1871), .B(n1870), .Z(n1872) );
  NAND U2069 ( .A(n1873), .B(n1872), .Z(n2018) );
  OR U2070 ( .A(n1875), .B(n1874), .Z(n1879) );
  OR U2071 ( .A(n1877), .B(n1876), .Z(n1878) );
  AND U2072 ( .A(n1879), .B(n1878), .Z(n2019) );
  XNOR U2073 ( .A(n2018), .B(n2019), .Z(n2020) );
  OR U2074 ( .A(n1881), .B(n1880), .Z(n1885) );
  NANDN U2075 ( .A(n1883), .B(n1882), .Z(n1884) );
  NAND U2076 ( .A(n1885), .B(n1884), .Z(n2027) );
  NANDN U2077 ( .A(n1887), .B(n1886), .Z(n1891) );
  NANDN U2078 ( .A(n1889), .B(n1888), .Z(n1890) );
  NAND U2079 ( .A(n1891), .B(n1890), .Z(n2024) );
  NANDN U2080 ( .A(n1893), .B(n1892), .Z(n1897) );
  NANDN U2081 ( .A(n1895), .B(n1894), .Z(n1896) );
  AND U2082 ( .A(n1897), .B(n1896), .Z(n2160) );
  NAND U2083 ( .A(x[2]), .B(y[24]), .Z(n2087) );
  AND U2084 ( .A(y[2]), .B(x[24]), .Z(n2088) );
  XOR U2085 ( .A(n2089), .B(n2088), .Z(n2037) );
  NANDN U2086 ( .A(n1899), .B(n1898), .Z(n1903) );
  NANDN U2087 ( .A(n1901), .B(n1900), .Z(n1902) );
  NAND U2088 ( .A(n1903), .B(n1902), .Z(n2036) );
  XNOR U2089 ( .A(n2037), .B(n2036), .Z(n2039) );
  OR U2090 ( .A(n1905), .B(n1904), .Z(n1909) );
  NANDN U2091 ( .A(n1907), .B(n1906), .Z(n1908) );
  NAND U2092 ( .A(n1909), .B(n1908), .Z(n2038) );
  XNOR U2093 ( .A(n2039), .B(n2038), .Z(n2161) );
  XNOR U2094 ( .A(n2160), .B(n2161), .Z(n2163) );
  NANDN U2095 ( .A(n1911), .B(n1910), .Z(n1915) );
  NAND U2096 ( .A(n1913), .B(n1912), .Z(n1914) );
  AND U2097 ( .A(n1915), .B(n1914), .Z(n2162) );
  XOR U2098 ( .A(n2163), .B(n2162), .Z(n2125) );
  NANDN U2099 ( .A(n1917), .B(n1916), .Z(n1921) );
  NANDN U2100 ( .A(n1919), .B(n1918), .Z(n1920) );
  NAND U2101 ( .A(n1921), .B(n1920), .Z(n2123) );
  NANDN U2102 ( .A(n1923), .B(n1922), .Z(n1927) );
  NANDN U2103 ( .A(n1925), .B(n1924), .Z(n1926) );
  NAND U2104 ( .A(n1927), .B(n1926), .Z(n2122) );
  XOR U2105 ( .A(n2123), .B(n2122), .Z(n2124) );
  XOR U2106 ( .A(n2125), .B(n2124), .Z(n2033) );
  NANDN U2107 ( .A(n1929), .B(n1928), .Z(n1933) );
  NAND U2108 ( .A(n1931), .B(n1930), .Z(n1932) );
  AND U2109 ( .A(n1933), .B(n1932), .Z(n2030) );
  ANDN U2110 ( .B(y[22]), .A(n2454), .Z(n2093) );
  XNOR U2111 ( .A(n2092), .B(n2093), .Z(n2095) );
  XNOR U2112 ( .A(n2094), .B(n2095), .Z(n2098) );
  OR U2113 ( .A(n1935), .B(n1934), .Z(n1939) );
  OR U2114 ( .A(n1937), .B(n1936), .Z(n1938) );
  NAND U2115 ( .A(n1939), .B(n1938), .Z(n2099) );
  XOR U2116 ( .A(n2098), .B(n2099), .Z(n2101) );
  NAND U2117 ( .A(y[7]), .B(x[19]), .Z(n2135) );
  AND U2118 ( .A(y[15]), .B(x[11]), .Z(n2134) );
  XNOR U2119 ( .A(n2135), .B(n2134), .Z(n2136) );
  NAND U2120 ( .A(y[23]), .B(x[3]), .Z(n2137) );
  XNOR U2121 ( .A(n2101), .B(n2100), .Z(n2062) );
  ANDN U2122 ( .B(y[5]), .A(n2431), .Z(n2148) );
  NAND U2123 ( .A(n1940), .B(n2148), .Z(n1944) );
  OR U2124 ( .A(n1942), .B(n1941), .Z(n1943) );
  NAND U2125 ( .A(n1944), .B(n1943), .Z(n2075) );
  NAND U2126 ( .A(y[4]), .B(x[22]), .Z(n2083) );
  NAND U2127 ( .A(y[3]), .B(x[23]), .Z(n2080) );
  XNOR U2128 ( .A(n2081), .B(n2080), .Z(n2082) );
  XNOR U2129 ( .A(n2083), .B(n2082), .Z(n2074) );
  XNOR U2130 ( .A(n2075), .B(n2074), .Z(n2077) );
  NAND U2131 ( .A(y[6]), .B(x[20]), .Z(n2149) );
  XNOR U2132 ( .A(n2148), .B(n2147), .Z(n2150) );
  XOR U2133 ( .A(n2149), .B(n2150), .Z(n2076) );
  XNOR U2134 ( .A(n2077), .B(n2076), .Z(n2063) );
  XNOR U2135 ( .A(n2062), .B(n2063), .Z(n2065) );
  ANDN U2136 ( .B(o[25]), .A(n1945), .Z(n2143) );
  ANDN U2137 ( .B(x[14]), .A(n2245), .Z(n2141) );
  ANDN U2138 ( .B(y[25]), .A(n25), .Z(n2142) );
  XNOR U2139 ( .A(n2141), .B(n2142), .Z(n2144) );
  XOR U2140 ( .A(n2143), .B(n2144), .Z(n2042) );
  NAND U2141 ( .A(x[0]), .B(y[26]), .Z(n2057) );
  AND U2142 ( .A(x[26]), .B(y[0]), .Z(n2056) );
  XNOR U2143 ( .A(n2057), .B(n2056), .Z(n2059) );
  NAND U2144 ( .A(x[25]), .B(y[1]), .Z(n2153) );
  XNOR U2145 ( .A(n2153), .B(o[26]), .Z(n2058) );
  XNOR U2146 ( .A(n2059), .B(n2058), .Z(n2043) );
  XNOR U2147 ( .A(n2042), .B(n2043), .Z(n2045) );
  OR U2148 ( .A(n1947), .B(n1946), .Z(n1951) );
  OR U2149 ( .A(n1949), .B(n1948), .Z(n1950) );
  NAND U2150 ( .A(n1951), .B(n1950), .Z(n2044) );
  XOR U2151 ( .A(n2045), .B(n2044), .Z(n2107) );
  OR U2152 ( .A(n1953), .B(n1952), .Z(n1957) );
  OR U2153 ( .A(n1955), .B(n1954), .Z(n1956) );
  AND U2154 ( .A(n1957), .B(n1956), .Z(n2105) );
  OR U2155 ( .A(n1959), .B(n1958), .Z(n1963) );
  OR U2156 ( .A(n1961), .B(n1960), .Z(n1962) );
  AND U2157 ( .A(n1963), .B(n1962), .Z(n2104) );
  XNOR U2158 ( .A(n2105), .B(n2104), .Z(n2106) );
  XNOR U2159 ( .A(n2107), .B(n2106), .Z(n2064) );
  XNOR U2160 ( .A(n2065), .B(n2064), .Z(n2070) );
  NANDN U2161 ( .A(n1965), .B(n1964), .Z(n1969) );
  OR U2162 ( .A(n1967), .B(n1966), .Z(n1968) );
  NAND U2163 ( .A(n1969), .B(n1968), .Z(n2111) );
  NANDN U2164 ( .A(n1971), .B(n1970), .Z(n1975) );
  NAND U2165 ( .A(n1973), .B(n1972), .Z(n1974) );
  NAND U2166 ( .A(n1975), .B(n1974), .Z(n2110) );
  XOR U2167 ( .A(n2111), .B(n2110), .Z(n2112) );
  ANDN U2168 ( .B(y[17]), .A(n2452), .Z(n2156) );
  ANDN U2169 ( .B(y[20]), .A(n2313), .Z(n2154) );
  ANDN U2170 ( .B(y[18]), .A(n29), .Z(n2155) );
  XNOR U2171 ( .A(n2154), .B(n2155), .Z(n2157) );
  XNOR U2172 ( .A(n2156), .B(n2157), .Z(n2131) );
  ANDN U2173 ( .B(x[7]), .A(n2140), .Z(n2128) );
  ANDN U2174 ( .B(x[12]), .A(n2429), .Z(n2050) );
  ANDN U2175 ( .B(y[21]), .A(n2252), .Z(n2051) );
  XNOR U2176 ( .A(n2050), .B(n2051), .Z(n2053) );
  XNOR U2177 ( .A(n2052), .B(n2053), .Z(n2129) );
  XNOR U2178 ( .A(n2128), .B(n2129), .Z(n2130) );
  XNOR U2179 ( .A(n2131), .B(n2130), .Z(n2113) );
  OR U2180 ( .A(n1977), .B(n1976), .Z(n1981) );
  OR U2181 ( .A(n1979), .B(n1978), .Z(n1980) );
  AND U2182 ( .A(n1981), .B(n1980), .Z(n2069) );
  XNOR U2183 ( .A(n2068), .B(n2069), .Z(n2071) );
  XNOR U2184 ( .A(n2070), .B(n2071), .Z(n2116) );
  OR U2185 ( .A(n1983), .B(n1982), .Z(n1987) );
  OR U2186 ( .A(n1985), .B(n1984), .Z(n1986) );
  NAND U2187 ( .A(n1987), .B(n1986), .Z(n2167) );
  NANDN U2188 ( .A(n1989), .B(n1988), .Z(n1993) );
  OR U2189 ( .A(n1991), .B(n1990), .Z(n1992) );
  NAND U2190 ( .A(n1993), .B(n1992), .Z(n2166) );
  XOR U2191 ( .A(n2167), .B(n2166), .Z(n2168) );
  NAND U2192 ( .A(n1995), .B(n1994), .Z(n1999) );
  OR U2193 ( .A(n1997), .B(n1996), .Z(n1998) );
  NAND U2194 ( .A(n1999), .B(n1998), .Z(n2169) );
  XNOR U2195 ( .A(n2116), .B(n2117), .Z(n2119) );
  OR U2196 ( .A(n2001), .B(n2000), .Z(n2005) );
  OR U2197 ( .A(n2003), .B(n2002), .Z(n2004) );
  NAND U2198 ( .A(n2005), .B(n2004), .Z(n2118) );
  XNOR U2199 ( .A(n2119), .B(n2118), .Z(n2031) );
  XNOR U2200 ( .A(n2030), .B(n2031), .Z(n2032) );
  XNOR U2201 ( .A(n2033), .B(n2032), .Z(n2174) );
  NANDN U2202 ( .A(n2007), .B(n2006), .Z(n2011) );
  NAND U2203 ( .A(n2009), .B(n2008), .Z(n2010) );
  NAND U2204 ( .A(n2011), .B(n2010), .Z(n2173) );
  NANDN U2205 ( .A(n2013), .B(n2012), .Z(n2017) );
  NANDN U2206 ( .A(n2015), .B(n2014), .Z(n2016) );
  NAND U2207 ( .A(n2017), .B(n2016), .Z(n2172) );
  XOR U2208 ( .A(n2173), .B(n2172), .Z(n2175) );
  XNOR U2209 ( .A(n2174), .B(n2175), .Z(n2025) );
  XNOR U2210 ( .A(n2027), .B(n2026), .Z(n2021) );
  XOR U2211 ( .A(n2020), .B(n2021), .Z(N59) );
  NANDN U2212 ( .A(n2019), .B(n2018), .Z(n2023) );
  NANDN U2213 ( .A(n2021), .B(n2020), .Z(n2022) );
  NAND U2214 ( .A(n2023), .B(n2022), .Z(n2178) );
  NANDN U2215 ( .A(n2025), .B(n2024), .Z(n2029) );
  NANDN U2216 ( .A(n2027), .B(n2026), .Z(n2028) );
  NAND U2217 ( .A(n2029), .B(n2028), .Z(n2179) );
  XNOR U2218 ( .A(n2178), .B(n2179), .Z(n2180) );
  OR U2219 ( .A(n2031), .B(n2030), .Z(n2035) );
  OR U2220 ( .A(n2033), .B(n2032), .Z(n2034) );
  AND U2221 ( .A(n2035), .B(n2034), .Z(n2184) );
  OR U2222 ( .A(n2037), .B(n2036), .Z(n2041) );
  OR U2223 ( .A(n2039), .B(n2038), .Z(n2040) );
  NAND U2224 ( .A(n2041), .B(n2040), .Z(n2318) );
  OR U2225 ( .A(n2043), .B(n2042), .Z(n2047) );
  OR U2226 ( .A(n2045), .B(n2044), .Z(n2046) );
  NAND U2227 ( .A(n2047), .B(n2046), .Z(n2316) );
  ANDN U2228 ( .B(x[12]), .A(n2048), .Z(n2289) );
  ANDN U2229 ( .B(y[14]), .A(n2049), .Z(n2290) );
  XNOR U2230 ( .A(n2289), .B(n2290), .Z(n2292) );
  NAND U2231 ( .A(y[11]), .B(x[16]), .Z(n2301) );
  XOR U2232 ( .A(n2302), .B(n2301), .Z(n2304) );
  XNOR U2233 ( .A(n2292), .B(n2291), .Z(n2222) );
  AND U2234 ( .A(y[24]), .B(x[3]), .Z(n2297) );
  ANDN U2235 ( .B(y[25]), .A(n26), .Z(n2295) );
  ANDN U2236 ( .B(x[15]), .A(n2245), .Z(n2296) );
  XNOR U2237 ( .A(n2295), .B(n2296), .Z(n2298) );
  XOR U2238 ( .A(n2297), .B(n2298), .Z(n2220) );
  NAND U2239 ( .A(y[21]), .B(x[6]), .Z(n2255) );
  ANDN U2240 ( .B(y[2]), .A(n2484), .Z(n2254) );
  NAND U2241 ( .A(y[8]), .B(x[19]), .Z(n2253) );
  XOR U2242 ( .A(n2254), .B(n2253), .Z(n2256) );
  XNOR U2243 ( .A(n2255), .B(n2256), .Z(n2221) );
  XNOR U2244 ( .A(n2220), .B(n2221), .Z(n2223) );
  XNOR U2245 ( .A(n2222), .B(n2223), .Z(n2279) );
  OR U2246 ( .A(n2051), .B(n2050), .Z(n2055) );
  OR U2247 ( .A(n2053), .B(n2052), .Z(n2054) );
  AND U2248 ( .A(n2055), .B(n2054), .Z(n2277) );
  NANDN U2249 ( .A(n2057), .B(n2056), .Z(n2061) );
  NAND U2250 ( .A(n2059), .B(n2058), .Z(n2060) );
  NAND U2251 ( .A(n2061), .B(n2060), .Z(n2278) );
  XOR U2252 ( .A(n2277), .B(n2278), .Z(n2280) );
  XNOR U2253 ( .A(n2279), .B(n2280), .Z(n2315) );
  XNOR U2254 ( .A(n2316), .B(n2315), .Z(n2317) );
  XNOR U2255 ( .A(n2318), .B(n2317), .Z(n2196) );
  OR U2256 ( .A(n2063), .B(n2062), .Z(n2067) );
  OR U2257 ( .A(n2065), .B(n2064), .Z(n2066) );
  NAND U2258 ( .A(n2067), .B(n2066), .Z(n2197) );
  XOR U2259 ( .A(n2196), .B(n2197), .Z(n2199) );
  OR U2260 ( .A(n2069), .B(n2068), .Z(n2073) );
  NANDN U2261 ( .A(n2071), .B(n2070), .Z(n2072) );
  AND U2262 ( .A(n2073), .B(n2072), .Z(n2198) );
  XOR U2263 ( .A(n2199), .B(n2198), .Z(n2341) );
  OR U2264 ( .A(n2075), .B(n2074), .Z(n2079) );
  OR U2265 ( .A(n2077), .B(n2076), .Z(n2078) );
  NAND U2266 ( .A(n2079), .B(n2078), .Z(n2203) );
  NANDN U2267 ( .A(n2081), .B(n2080), .Z(n2085) );
  NAND U2268 ( .A(n2083), .B(n2082), .Z(n2084) );
  AND U2269 ( .A(n2085), .B(n2084), .Z(n2271) );
  NANDN U2270 ( .A(n2087), .B(n2086), .Z(n2091) );
  NANDN U2271 ( .A(n2089), .B(n2088), .Z(n2090) );
  NAND U2272 ( .A(n2091), .B(n2090), .Z(n2272) );
  XOR U2273 ( .A(n2271), .B(n2272), .Z(n2273) );
  OR U2274 ( .A(n2093), .B(n2092), .Z(n2097) );
  OR U2275 ( .A(n2095), .B(n2094), .Z(n2096) );
  AND U2276 ( .A(n2097), .B(n2096), .Z(n2265) );
  ANDN U2277 ( .B(y[18]), .A(n2452), .Z(n2228) );
  ANDN U2278 ( .B(x[18]), .A(n2314), .Z(n2226) );
  ANDN U2279 ( .B(y[6]), .A(n2431), .Z(n2227) );
  XNOR U2280 ( .A(n2226), .B(n2227), .Z(n2229) );
  XNOR U2281 ( .A(n2228), .B(n2229), .Z(n2266) );
  XOR U2282 ( .A(n2265), .B(n2266), .Z(n2267) );
  ANDN U2283 ( .B(y[27]), .A(n24), .Z(n2235) );
  ANDN U2284 ( .B(x[26]), .A(n18), .Z(n2232) );
  XOR U2285 ( .A(o[27]), .B(n2232), .Z(n2233) );
  ANDN U2286 ( .B(x[27]), .A(n17), .Z(n2234) );
  XNOR U2287 ( .A(n2233), .B(n2234), .Z(n2236) );
  XNOR U2288 ( .A(n2235), .B(n2236), .Z(n2268) );
  XOR U2289 ( .A(n2273), .B(n2274), .Z(n2321) );
  NANDN U2290 ( .A(n2099), .B(n2098), .Z(n2103) );
  NANDN U2291 ( .A(n2101), .B(n2100), .Z(n2102) );
  AND U2292 ( .A(n2103), .B(n2102), .Z(n2322) );
  XOR U2293 ( .A(n2321), .B(n2322), .Z(n2324) );
  OR U2294 ( .A(n2105), .B(n2104), .Z(n2109) );
  OR U2295 ( .A(n2107), .B(n2106), .Z(n2108) );
  NAND U2296 ( .A(n2109), .B(n2108), .Z(n2323) );
  XNOR U2297 ( .A(n2324), .B(n2323), .Z(n2202) );
  XNOR U2298 ( .A(n2203), .B(n2202), .Z(n2205) );
  OR U2299 ( .A(n2111), .B(n2110), .Z(n2115) );
  NANDN U2300 ( .A(n2113), .B(n2112), .Z(n2114) );
  NAND U2301 ( .A(n2115), .B(n2114), .Z(n2204) );
  XOR U2302 ( .A(n2205), .B(n2204), .Z(n2339) );
  OR U2303 ( .A(n2117), .B(n2116), .Z(n2121) );
  OR U2304 ( .A(n2119), .B(n2118), .Z(n2120) );
  NAND U2305 ( .A(n2121), .B(n2120), .Z(n2340) );
  XOR U2306 ( .A(n2341), .B(n2342), .Z(n2335) );
  OR U2307 ( .A(n2123), .B(n2122), .Z(n2127) );
  NANDN U2308 ( .A(n2125), .B(n2124), .Z(n2126) );
  AND U2309 ( .A(n2127), .B(n2126), .Z(n2333) );
  OR U2310 ( .A(n2129), .B(n2128), .Z(n2133) );
  OR U2311 ( .A(n2131), .B(n2130), .Z(n2132) );
  AND U2312 ( .A(n2133), .B(n2132), .Z(n2192) );
  NANDN U2313 ( .A(n2135), .B(n2134), .Z(n2139) );
  NANDN U2314 ( .A(n2137), .B(n2136), .Z(n2138) );
  AND U2315 ( .A(n2139), .B(n2138), .Z(n2216) );
  ANDN U2316 ( .B(x[22]), .A(n22), .Z(n2309) );
  ANDN U2317 ( .B(x[23]), .A(n21), .Z(n2307) );
  ANDN U2318 ( .B(x[8]), .A(n2140), .Z(n2308) );
  XNOR U2319 ( .A(n2307), .B(n2308), .Z(n2310) );
  XOR U2320 ( .A(n2309), .B(n2310), .Z(n2214) );
  NAND U2321 ( .A(x[7]), .B(y[20]), .Z(n2248) );
  NAND U2322 ( .A(y[3]), .B(x[24]), .Z(n2246) );
  XOR U2323 ( .A(n2247), .B(n2246), .Z(n2249) );
  XNOR U2324 ( .A(n2248), .B(n2249), .Z(n2215) );
  XNOR U2325 ( .A(n2214), .B(n2215), .Z(n2217) );
  XOR U2326 ( .A(n2216), .B(n2217), .Z(n2190) );
  OR U2327 ( .A(n2142), .B(n2141), .Z(n2146) );
  OR U2328 ( .A(n2144), .B(n2143), .Z(n2145) );
  NAND U2329 ( .A(n2146), .B(n2145), .Z(n2209) );
  OR U2330 ( .A(n2148), .B(n2147), .Z(n2152) );
  NANDN U2331 ( .A(n2150), .B(n2149), .Z(n2151) );
  NAND U2332 ( .A(n2152), .B(n2151), .Z(n2208) );
  XOR U2333 ( .A(n2209), .B(n2208), .Z(n2211) );
  ANDN U2334 ( .B(y[10]), .A(n2483), .Z(n2241) );
  ANDN U2335 ( .B(y[22]), .A(n2252), .Z(n2239) );
  IV U2336 ( .A(y[23]), .Z(n2456) );
  ANDN U2337 ( .B(x[4]), .A(n2456), .Z(n2240) );
  XNOR U2338 ( .A(n2239), .B(n2240), .Z(n2242) );
  XOR U2339 ( .A(n2241), .B(n2242), .Z(n2259) );
  NAND U2340 ( .A(y[13]), .B(x[14]), .Z(n2285) );
  ANDN U2341 ( .B(o[26]), .A(n2153), .Z(n2284) );
  NAND U2342 ( .A(x[1]), .B(y[26]), .Z(n2283) );
  XOR U2343 ( .A(n2284), .B(n2283), .Z(n2286) );
  XNOR U2344 ( .A(n2285), .B(n2286), .Z(n2260) );
  XNOR U2345 ( .A(n2259), .B(n2260), .Z(n2262) );
  OR U2346 ( .A(n2155), .B(n2154), .Z(n2159) );
  OR U2347 ( .A(n2157), .B(n2156), .Z(n2158) );
  NAND U2348 ( .A(n2159), .B(n2158), .Z(n2261) );
  XOR U2349 ( .A(n2262), .B(n2261), .Z(n2210) );
  XOR U2350 ( .A(n2211), .B(n2210), .Z(n2191) );
  XNOR U2351 ( .A(n2190), .B(n2191), .Z(n2193) );
  XOR U2352 ( .A(n2192), .B(n2193), .Z(n2327) );
  OR U2353 ( .A(n2161), .B(n2160), .Z(n2165) );
  OR U2354 ( .A(n2163), .B(n2162), .Z(n2164) );
  AND U2355 ( .A(n2165), .B(n2164), .Z(n2328) );
  XNOR U2356 ( .A(n2327), .B(n2328), .Z(n2330) );
  OR U2357 ( .A(n2167), .B(n2166), .Z(n2171) );
  NANDN U2358 ( .A(n2169), .B(n2168), .Z(n2170) );
  NAND U2359 ( .A(n2171), .B(n2170), .Z(n2329) );
  XOR U2360 ( .A(n2330), .B(n2329), .Z(n2334) );
  XOR U2361 ( .A(n2333), .B(n2334), .Z(n2336) );
  XNOR U2362 ( .A(n2335), .B(n2336), .Z(n2185) );
  XOR U2363 ( .A(n2184), .B(n2185), .Z(n2186) );
  OR U2364 ( .A(n2173), .B(n2172), .Z(n2177) );
  NAND U2365 ( .A(n2175), .B(n2174), .Z(n2176) );
  NAND U2366 ( .A(n2177), .B(n2176), .Z(n2187) );
  XOR U2367 ( .A(n2180), .B(n2181), .Z(N60) );
  NANDN U2368 ( .A(n2179), .B(n2178), .Z(n2183) );
  NANDN U2369 ( .A(n2181), .B(n2180), .Z(n2182) );
  NAND U2370 ( .A(n2183), .B(n2182), .Z(n2345) );
  OR U2371 ( .A(n2185), .B(n2184), .Z(n2189) );
  NANDN U2372 ( .A(n2187), .B(n2186), .Z(n2188) );
  AND U2373 ( .A(n2189), .B(n2188), .Z(n2346) );
  XNOR U2374 ( .A(n2345), .B(n2346), .Z(n2347) );
  OR U2375 ( .A(n2191), .B(n2190), .Z(n2195) );
  OR U2376 ( .A(n2193), .B(n2192), .Z(n2194) );
  AND U2377 ( .A(n2195), .B(n2194), .Z(n2522) );
  NANDN U2378 ( .A(n2197), .B(n2196), .Z(n2201) );
  OR U2379 ( .A(n2199), .B(n2198), .Z(n2200) );
  NAND U2380 ( .A(n2201), .B(n2200), .Z(n2520) );
  OR U2381 ( .A(n2203), .B(n2202), .Z(n2207) );
  OR U2382 ( .A(n2205), .B(n2204), .Z(n2206) );
  NAND U2383 ( .A(n2207), .B(n2206), .Z(n2519) );
  XOR U2384 ( .A(n2520), .B(n2519), .Z(n2521) );
  XNOR U2385 ( .A(n2522), .B(n2521), .Z(n2527) );
  OR U2386 ( .A(n2209), .B(n2208), .Z(n2213) );
  NAND U2387 ( .A(n2211), .B(n2210), .Z(n2212) );
  AND U2388 ( .A(n2213), .B(n2212), .Z(n2396) );
  OR U2389 ( .A(n2215), .B(n2214), .Z(n2219) );
  OR U2390 ( .A(n2217), .B(n2216), .Z(n2218) );
  AND U2391 ( .A(n2219), .B(n2218), .Z(n2393) );
  OR U2392 ( .A(n2221), .B(n2220), .Z(n2225) );
  OR U2393 ( .A(n2223), .B(n2222), .Z(n2224) );
  AND U2394 ( .A(n2225), .B(n2224), .Z(n2394) );
  XOR U2395 ( .A(n2393), .B(n2394), .Z(n2395) );
  OR U2396 ( .A(n2227), .B(n2226), .Z(n2231) );
  OR U2397 ( .A(n2229), .B(n2228), .Z(n2230) );
  AND U2398 ( .A(n2231), .B(n2230), .Z(n2405) );
  ANDN U2399 ( .B(y[18]), .A(n2455), .Z(n2425) );
  ANDN U2400 ( .B(y[19]), .A(n2452), .Z(n2423) );
  ANDN U2401 ( .B(x[8]), .A(n2453), .Z(n2424) );
  XNOR U2402 ( .A(n2423), .B(n2424), .Z(n2426) );
  XNOR U2403 ( .A(n2425), .B(n2426), .Z(n2406) );
  XOR U2404 ( .A(n2405), .B(n2406), .Z(n2407) );
  NAND U2405 ( .A(x[0]), .B(y[28]), .Z(n2414) );
  AND U2406 ( .A(n2232), .B(o[27]), .Z(n2412) );
  NAND U2407 ( .A(y[0]), .B(x[28]), .Z(n2411) );
  XNOR U2408 ( .A(n2412), .B(n2411), .Z(n2413) );
  XNOR U2409 ( .A(n2414), .B(n2413), .Z(n2408) );
  OR U2410 ( .A(n2234), .B(n2233), .Z(n2238) );
  OR U2411 ( .A(n2236), .B(n2235), .Z(n2237) );
  NAND U2412 ( .A(n2238), .B(n2237), .Z(n2382) );
  OR U2413 ( .A(n2240), .B(n2239), .Z(n2244) );
  OR U2414 ( .A(n2242), .B(n2241), .Z(n2243) );
  NAND U2415 ( .A(n2244), .B(n2243), .Z(n2381) );
  XOR U2416 ( .A(n2382), .B(n2381), .Z(n2383) );
  ANDN U2417 ( .B(y[27]), .A(n25), .Z(n2464) );
  ANDN U2418 ( .B(y[3]), .A(n2484), .Z(n2465) );
  XNOR U2419 ( .A(n2464), .B(n2465), .Z(n2467) );
  XNOR U2420 ( .A(n2466), .B(n2467), .Z(n2371) );
  ANDN U2421 ( .B(x[16]), .A(n2245), .Z(n2472) );
  ANDN U2422 ( .B(y[26]), .A(n26), .Z(n2470) );
  XNOR U2423 ( .A(n2470), .B(n2471), .Z(n2473) );
  XOR U2424 ( .A(n2472), .B(n2473), .Z(n2369) );
  NANDN U2425 ( .A(n2247), .B(n2246), .Z(n2251) );
  NANDN U2426 ( .A(n2249), .B(n2248), .Z(n2250) );
  NAND U2427 ( .A(n2251), .B(n2250), .Z(n2370) );
  XNOR U2428 ( .A(n2369), .B(n2370), .Z(n2372) );
  XNOR U2429 ( .A(n2371), .B(n2372), .Z(n2357) );
  ANDN U2430 ( .B(x[23]), .A(n22), .Z(n2440) );
  ANDN U2431 ( .B(y[25]), .A(n27), .Z(n2441) );
  XNOR U2432 ( .A(n2440), .B(n2441), .Z(n2443) );
  XNOR U2433 ( .A(n2442), .B(n2443), .Z(n2377) );
  ANDN U2434 ( .B(y[23]), .A(n2252), .Z(n2493) );
  ANDN U2435 ( .B(y[8]), .A(n2432), .Z(n2491) );
  ANDN U2436 ( .B(x[21]), .A(n2433), .Z(n2492) );
  XNOR U2437 ( .A(n2491), .B(n2492), .Z(n2494) );
  XOR U2438 ( .A(n2493), .B(n2494), .Z(n2376) );
  NANDN U2439 ( .A(n2254), .B(n2253), .Z(n2258) );
  NANDN U2440 ( .A(n2256), .B(n2255), .Z(n2257) );
  NAND U2441 ( .A(n2258), .B(n2257), .Z(n2375) );
  XNOR U2442 ( .A(n2376), .B(n2375), .Z(n2378) );
  XNOR U2443 ( .A(n2377), .B(n2378), .Z(n2358) );
  XNOR U2444 ( .A(n2357), .B(n2358), .Z(n2360) );
  XNOR U2445 ( .A(n2359), .B(n2360), .Z(n2513) );
  XNOR U2446 ( .A(n2514), .B(n2513), .Z(n2516) );
  OR U2447 ( .A(n2260), .B(n2259), .Z(n2264) );
  OR U2448 ( .A(n2262), .B(n2261), .Z(n2263) );
  AND U2449 ( .A(n2264), .B(n2263), .Z(n2387) );
  OR U2450 ( .A(n2266), .B(n2265), .Z(n2270) );
  NANDN U2451 ( .A(n2268), .B(n2267), .Z(n2269) );
  NAND U2452 ( .A(n2270), .B(n2269), .Z(n2388) );
  XOR U2453 ( .A(n2387), .B(n2388), .Z(n2389) );
  OR U2454 ( .A(n2272), .B(n2271), .Z(n2276) );
  NANDN U2455 ( .A(n2274), .B(n2273), .Z(n2275) );
  NAND U2456 ( .A(n2276), .B(n2275), .Z(n2390) );
  XNOR U2457 ( .A(n2389), .B(n2390), .Z(n2504) );
  OR U2458 ( .A(n2278), .B(n2277), .Z(n2282) );
  NAND U2459 ( .A(n2280), .B(n2279), .Z(n2281) );
  AND U2460 ( .A(n2282), .B(n2281), .Z(n2501) );
  NANDN U2461 ( .A(n2284), .B(n2283), .Z(n2288) );
  NANDN U2462 ( .A(n2286), .B(n2285), .Z(n2287) );
  AND U2463 ( .A(n2288), .B(n2287), .Z(n2402) );
  OR U2464 ( .A(n2290), .B(n2289), .Z(n2294) );
  NANDN U2465 ( .A(n2292), .B(n2291), .Z(n2293) );
  AND U2466 ( .A(n2294), .B(n2293), .Z(n2399) );
  OR U2467 ( .A(n2296), .B(n2295), .Z(n2300) );
  OR U2468 ( .A(n2298), .B(n2297), .Z(n2299) );
  AND U2469 ( .A(n2300), .B(n2299), .Z(n2400) );
  XOR U2470 ( .A(n2399), .B(n2400), .Z(n2401) );
  ANDN U2471 ( .B(x[7]), .A(n2457), .Z(n2478) );
  ANDN U2472 ( .B(y[17]), .A(n2482), .Z(n2476) );
  XNOR U2473 ( .A(n2476), .B(n2477), .Z(n2479) );
  XOR U2474 ( .A(n2478), .B(n2479), .Z(n2458) );
  NANDN U2475 ( .A(n2302), .B(n2301), .Z(n2306) );
  OR U2476 ( .A(n2304), .B(n2303), .Z(n2305) );
  NAND U2477 ( .A(n2306), .B(n2305), .Z(n2459) );
  XNOR U2478 ( .A(n2458), .B(n2459), .Z(n2461) );
  NAND U2479 ( .A(y[13]), .B(x[15]), .Z(n2447) );
  AND U2480 ( .A(x[26]), .B(y[2]), .Z(n2446) );
  XNOR U2481 ( .A(n2447), .B(n2446), .Z(n2448) );
  AND U2482 ( .A(x[27]), .B(y[1]), .Z(n2588) );
  XNOR U2483 ( .A(o[28]), .B(n2588), .Z(n2449) );
  XNOR U2484 ( .A(n2461), .B(n2460), .Z(n2363) );
  OR U2485 ( .A(n2308), .B(n2307), .Z(n2312) );
  OR U2486 ( .A(n2310), .B(n2309), .Z(n2311) );
  AND U2487 ( .A(n2312), .B(n2311), .Z(n2434) );
  ANDN U2488 ( .B(y[22]), .A(n2313), .Z(n2487) );
  ANDN U2489 ( .B(x[19]), .A(n2314), .Z(n2486) );
  XNOR U2490 ( .A(n2485), .B(n2486), .Z(n2488) );
  XNOR U2491 ( .A(n2487), .B(n2488), .Z(n2435) );
  XOR U2492 ( .A(n2434), .B(n2435), .Z(n2436) );
  ANDN U2493 ( .B(y[11]), .A(n2483), .Z(n2419) );
  AND U2494 ( .A(y[24]), .B(x[4]), .Z(n2417) );
  ANDN U2495 ( .B(x[22]), .A(n23), .Z(n2418) );
  XNOR U2496 ( .A(n2417), .B(n2418), .Z(n2420) );
  XNOR U2497 ( .A(n2419), .B(n2420), .Z(n2437) );
  XOR U2498 ( .A(n2366), .B(n2365), .Z(n2502) );
  XOR U2499 ( .A(n2501), .B(n2502), .Z(n2503) );
  XOR U2500 ( .A(n2516), .B(n2515), .Z(n2510) );
  OR U2501 ( .A(n2316), .B(n2315), .Z(n2320) );
  OR U2502 ( .A(n2318), .B(n2317), .Z(n2319) );
  AND U2503 ( .A(n2320), .B(n2319), .Z(n2507) );
  NANDN U2504 ( .A(n2322), .B(n2321), .Z(n2326) );
  OR U2505 ( .A(n2324), .B(n2323), .Z(n2325) );
  NAND U2506 ( .A(n2326), .B(n2325), .Z(n2508) );
  XOR U2507 ( .A(n2507), .B(n2508), .Z(n2509) );
  OR U2508 ( .A(n2328), .B(n2327), .Z(n2332) );
  OR U2509 ( .A(n2330), .B(n2329), .Z(n2331) );
  AND U2510 ( .A(n2332), .B(n2331), .Z(n2526) );
  XNOR U2511 ( .A(n2525), .B(n2526), .Z(n2528) );
  XNOR U2512 ( .A(n2527), .B(n2528), .Z(n2351) );
  OR U2513 ( .A(n2334), .B(n2333), .Z(n2338) );
  NAND U2514 ( .A(n2336), .B(n2335), .Z(n2337) );
  AND U2515 ( .A(n2338), .B(n2337), .Z(n2352) );
  XOR U2516 ( .A(n2351), .B(n2352), .Z(n2354) );
  NANDN U2517 ( .A(n2340), .B(n2339), .Z(n2344) );
  NANDN U2518 ( .A(n2342), .B(n2341), .Z(n2343) );
  NAND U2519 ( .A(n2344), .B(n2343), .Z(n2353) );
  XOR U2520 ( .A(n2354), .B(n2353), .Z(n2348) );
  XNOR U2521 ( .A(n2347), .B(n2348), .Z(N61) );
  NANDN U2522 ( .A(n2346), .B(n2345), .Z(n2350) );
  NAND U2523 ( .A(n2348), .B(n2347), .Z(n2349) );
  NAND U2524 ( .A(n2350), .B(n2349), .Z(n2531) );
  NANDN U2525 ( .A(n2352), .B(n2351), .Z(n2356) );
  OR U2526 ( .A(n2354), .B(n2353), .Z(n2355) );
  AND U2527 ( .A(n2356), .B(n2355), .Z(n2532) );
  XNOR U2528 ( .A(n2531), .B(n2532), .Z(n2533) );
  OR U2529 ( .A(n2358), .B(n2357), .Z(n2362) );
  NANDN U2530 ( .A(n2360), .B(n2359), .Z(n2361) );
  AND U2531 ( .A(n2362), .B(n2361), .Z(n2684) );
  NAND U2532 ( .A(n2364), .B(n2363), .Z(n2368) );
  NANDN U2533 ( .A(n2366), .B(n2365), .Z(n2367) );
  NAND U2534 ( .A(n2368), .B(n2367), .Z(n2689) );
  OR U2535 ( .A(n2370), .B(n2369), .Z(n2374) );
  NANDN U2536 ( .A(n2372), .B(n2371), .Z(n2373) );
  NAND U2537 ( .A(n2374), .B(n2373), .Z(n2546) );
  OR U2538 ( .A(n2376), .B(n2375), .Z(n2380) );
  NANDN U2539 ( .A(n2378), .B(n2377), .Z(n2379) );
  NAND U2540 ( .A(n2380), .B(n2379), .Z(n2544) );
  OR U2541 ( .A(n2382), .B(n2381), .Z(n2386) );
  NANDN U2542 ( .A(n2384), .B(n2383), .Z(n2385) );
  NAND U2543 ( .A(n2386), .B(n2385), .Z(n2543) );
  XNOR U2544 ( .A(n2544), .B(n2543), .Z(n2545) );
  XNOR U2545 ( .A(n2546), .B(n2545), .Z(n2688) );
  XOR U2546 ( .A(n2689), .B(n2688), .Z(n2691) );
  OR U2547 ( .A(n2388), .B(n2387), .Z(n2392) );
  NANDN U2548 ( .A(n2390), .B(n2389), .Z(n2391) );
  AND U2549 ( .A(n2392), .B(n2391), .Z(n2690) );
  XOR U2550 ( .A(n2691), .B(n2690), .Z(n2682) );
  OR U2551 ( .A(n2394), .B(n2393), .Z(n2398) );
  NANDN U2552 ( .A(n2396), .B(n2395), .Z(n2397) );
  NAND U2553 ( .A(n2398), .B(n2397), .Z(n2683) );
  XNOR U2554 ( .A(n2682), .B(n2683), .Z(n2685) );
  XOR U2555 ( .A(n2684), .B(n2685), .Z(n2697) );
  OR U2556 ( .A(n2400), .B(n2399), .Z(n2404) );
  NANDN U2557 ( .A(n2402), .B(n2401), .Z(n2403) );
  AND U2558 ( .A(n2404), .B(n2403), .Z(n2678) );
  OR U2559 ( .A(n2406), .B(n2405), .Z(n2410) );
  NANDN U2560 ( .A(n2408), .B(n2407), .Z(n2409) );
  AND U2561 ( .A(n2410), .B(n2409), .Z(n2676) );
  NANDN U2562 ( .A(n2412), .B(n2411), .Z(n2416) );
  NAND U2563 ( .A(n2414), .B(n2413), .Z(n2415) );
  AND U2564 ( .A(n2416), .B(n2415), .Z(n2673) );
  OR U2565 ( .A(n2418), .B(n2417), .Z(n2422) );
  OR U2566 ( .A(n2420), .B(n2419), .Z(n2421) );
  AND U2567 ( .A(n2422), .B(n2421), .Z(n2670) );
  OR U2568 ( .A(n2424), .B(n2423), .Z(n2428) );
  OR U2569 ( .A(n2426), .B(n2425), .Z(n2427) );
  AND U2570 ( .A(n2428), .B(n2427), .Z(n2645) );
  ANDN U2571 ( .B(x[15]), .A(n2429), .Z(n2621) );
  NOR U2572 ( .A(n2431), .B(n2430), .Z(n2890) );
  ANDN U2573 ( .B(y[9]), .A(n2432), .Z(n2620) );
  XNOR U2574 ( .A(n2890), .B(n2620), .Z(n2622) );
  XNOR U2575 ( .A(n2621), .B(n2622), .Z(n2646) );
  XOR U2576 ( .A(n2645), .B(n2646), .Z(n2647) );
  AND U2577 ( .A(y[17]), .B(x[12]), .Z(n2836) );
  ANDN U2578 ( .B(x[22]), .A(n2433), .Z(n2616) );
  NAND U2579 ( .A(x[1]), .B(y[28]), .Z(n2615) );
  XOR U2580 ( .A(n2616), .B(n2615), .Z(n2617) );
  XNOR U2581 ( .A(n2836), .B(n2617), .Z(n2648) );
  XOR U2582 ( .A(n2647), .B(n2648), .Z(n2671) );
  XOR U2583 ( .A(n2670), .B(n2671), .Z(n2672) );
  XNOR U2584 ( .A(n2676), .B(n2677), .Z(n2679) );
  XOR U2585 ( .A(n2678), .B(n2679), .Z(n2633) );
  OR U2586 ( .A(n2435), .B(n2434), .Z(n2439) );
  NANDN U2587 ( .A(n2437), .B(n2436), .Z(n2438) );
  NAND U2588 ( .A(n2439), .B(n2438), .Z(n2634) );
  XNOR U2589 ( .A(n2633), .B(n2634), .Z(n2636) );
  OR U2590 ( .A(n2441), .B(n2440), .Z(n2445) );
  OR U2591 ( .A(n2443), .B(n2442), .Z(n2444) );
  AND U2592 ( .A(n2445), .B(n2444), .Z(n2561) );
  NANDN U2593 ( .A(n2447), .B(n2446), .Z(n2451) );
  NANDN U2594 ( .A(n2449), .B(n2448), .Z(n2450) );
  NAND U2595 ( .A(n2451), .B(n2450), .Z(n2562) );
  XOR U2596 ( .A(n2561), .B(n2562), .Z(n2563) );
  NOR U2597 ( .A(n2453), .B(n2452), .Z(n2760) );
  ANDN U2598 ( .B(y[25]), .A(n2454), .Z(n2584) );
  AND U2599 ( .A(y[24]), .B(x[5]), .Z(n2848) );
  ANDN U2600 ( .B(y[19]), .A(n2455), .Z(n2583) );
  XNOR U2601 ( .A(n2848), .B(n2583), .Z(n2585) );
  XNOR U2602 ( .A(n2584), .B(n2585), .Z(n2657) );
  XNOR U2603 ( .A(n2760), .B(n2657), .Z(n2659) );
  ANDN U2604 ( .B(x[6]), .A(n2456), .Z(n2609) );
  ANDN U2605 ( .B(x[8]), .A(n2457), .Z(n2607) );
  ANDN U2606 ( .B(y[22]), .A(n28), .Z(n2608) );
  XNOR U2607 ( .A(n2607), .B(n2608), .Z(n2610) );
  XNOR U2608 ( .A(n2609), .B(n2610), .Z(n2658) );
  XNOR U2609 ( .A(n2659), .B(n2658), .Z(n2564) );
  XOR U2610 ( .A(n2563), .B(n2564), .Z(n2557) );
  OR U2611 ( .A(n2459), .B(n2458), .Z(n2463) );
  OR U2612 ( .A(n2461), .B(n2460), .Z(n2462) );
  AND U2613 ( .A(n2463), .B(n2462), .Z(n2556) );
  OR U2614 ( .A(n2465), .B(n2464), .Z(n2469) );
  OR U2615 ( .A(n2467), .B(n2466), .Z(n2468) );
  AND U2616 ( .A(n2469), .B(n2468), .Z(n2642) );
  OR U2617 ( .A(n2471), .B(n2470), .Z(n2475) );
  OR U2618 ( .A(n2473), .B(n2472), .Z(n2474) );
  AND U2619 ( .A(n2475), .B(n2474), .Z(n2639) );
  OR U2620 ( .A(n2477), .B(n2476), .Z(n2481) );
  OR U2621 ( .A(n2479), .B(n2478), .Z(n2480) );
  AND U2622 ( .A(n2481), .B(n2480), .Z(n2567) );
  AND U2623 ( .A(y[26]), .B(x[3]), .Z(n2896) );
  ANDN U2624 ( .B(y[18]), .A(n2482), .Z(n2599) );
  ANDN U2625 ( .B(y[12]), .A(n2483), .Z(n2600) );
  XNOR U2626 ( .A(n2599), .B(n2600), .Z(n2601) );
  XNOR U2627 ( .A(n2896), .B(n2601), .Z(n2568) );
  XOR U2628 ( .A(n2567), .B(n2568), .Z(n2569) );
  NAND U2629 ( .A(y[16]), .B(x[13]), .Z(n2604) );
  AND U2630 ( .A(x[23]), .B(y[6]), .Z(n2771) );
  NAND U2631 ( .A(x[24]), .B(y[5]), .Z(n2602) );
  XNOR U2632 ( .A(n2771), .B(n2602), .Z(n2603) );
  XNOR U2633 ( .A(n2604), .B(n2603), .Z(n2570) );
  XOR U2634 ( .A(n2569), .B(n2570), .Z(n2640) );
  XOR U2635 ( .A(n2639), .B(n2640), .Z(n2641) );
  ANDN U2636 ( .B(y[29]), .A(n24), .Z(n2666) );
  ANDN U2637 ( .B(x[28]), .A(n18), .Z(n2623) );
  XOR U2638 ( .A(o[29]), .B(n2623), .Z(n2664) );
  ANDN U2639 ( .B(x[29]), .A(n17), .Z(n2665) );
  XNOR U2640 ( .A(n2664), .B(n2665), .Z(n2667) );
  XOR U2641 ( .A(n2666), .B(n2667), .Z(n2651) );
  NAND U2642 ( .A(x[14]), .B(y[15]), .Z(n2628) );
  ANDN U2643 ( .B(y[4]), .A(n2484), .Z(n2627) );
  NAND U2644 ( .A(y[3]), .B(x[26]), .Z(n2626) );
  XOR U2645 ( .A(n2627), .B(n2626), .Z(n2629) );
  XNOR U2646 ( .A(n2628), .B(n2629), .Z(n2652) );
  XNOR U2647 ( .A(n2651), .B(n2652), .Z(n2654) );
  OR U2648 ( .A(n2486), .B(n2485), .Z(n2490) );
  OR U2649 ( .A(n2488), .B(n2487), .Z(n2489) );
  NAND U2650 ( .A(n2490), .B(n2489), .Z(n2653) );
  XNOR U2651 ( .A(n2654), .B(n2653), .Z(n2549) );
  OR U2652 ( .A(n2492), .B(n2491), .Z(n2496) );
  OR U2653 ( .A(n2494), .B(n2493), .Z(n2495) );
  AND U2654 ( .A(n2496), .B(n2495), .Z(n2593) );
  NAND U2655 ( .A(y[1]), .B(o[28]), .Z(n2497) );
  XNOR U2656 ( .A(y[2]), .B(n2497), .Z(n2498) );
  NAND U2657 ( .A(n2498), .B(x[27]), .Z(n2587) );
  XNOR U2658 ( .A(n2587), .B(n2586), .Z(n2594) );
  XOR U2659 ( .A(n2593), .B(n2594), .Z(n2595) );
  ANDN U2660 ( .B(x[18]), .A(n2499), .Z(n2573) );
  ANDN U2661 ( .B(x[19]), .A(n2500), .Z(n2574) );
  XNOR U2662 ( .A(n2573), .B(n2574), .Z(n2576) );
  ANDN U2663 ( .B(y[27]), .A(n26), .Z(n2575) );
  XNOR U2664 ( .A(n2576), .B(n2575), .Z(n2596) );
  XOR U2665 ( .A(n2552), .B(n2551), .Z(n2555) );
  XOR U2666 ( .A(n2556), .B(n2555), .Z(n2558) );
  XNOR U2667 ( .A(n2557), .B(n2558), .Z(n2635) );
  XOR U2668 ( .A(n2636), .B(n2635), .Z(n2695) );
  OR U2669 ( .A(n2502), .B(n2501), .Z(n2506) );
  NANDN U2670 ( .A(n2504), .B(n2503), .Z(n2505) );
  NAND U2671 ( .A(n2506), .B(n2505), .Z(n2694) );
  XOR U2672 ( .A(n2695), .B(n2694), .Z(n2696) );
  OR U2673 ( .A(n2508), .B(n2507), .Z(n2512) );
  NANDN U2674 ( .A(n2510), .B(n2509), .Z(n2511) );
  AND U2675 ( .A(n2512), .B(n2511), .Z(n2700) );
  OR U2676 ( .A(n2514), .B(n2513), .Z(n2518) );
  OR U2677 ( .A(n2516), .B(n2515), .Z(n2517) );
  NAND U2678 ( .A(n2518), .B(n2517), .Z(n2701) );
  XOR U2679 ( .A(n2700), .B(n2701), .Z(n2702) );
  XOR U2680 ( .A(n2703), .B(n2702), .Z(n2540) );
  OR U2681 ( .A(n2520), .B(n2519), .Z(n2524) );
  NANDN U2682 ( .A(n2522), .B(n2521), .Z(n2523) );
  AND U2683 ( .A(n2524), .B(n2523), .Z(n2537) );
  OR U2684 ( .A(n2526), .B(n2525), .Z(n2530) );
  OR U2685 ( .A(n2528), .B(n2527), .Z(n2529) );
  NAND U2686 ( .A(n2530), .B(n2529), .Z(n2538) );
  XNOR U2687 ( .A(n2537), .B(n2538), .Z(n2539) );
  XOR U2688 ( .A(n2540), .B(n2539), .Z(n2534) );
  XNOR U2689 ( .A(n2533), .B(n2534), .Z(N62) );
  NANDN U2690 ( .A(n2532), .B(n2531), .Z(n2536) );
  NAND U2691 ( .A(n2534), .B(n2533), .Z(n2535) );
  AND U2692 ( .A(n2536), .B(n2535), .Z(n2708) );
  OR U2693 ( .A(n2538), .B(n2537), .Z(n2542) );
  OR U2694 ( .A(n2540), .B(n2539), .Z(n2541) );
  AND U2695 ( .A(n2542), .B(n2541), .Z(n2709) );
  XNOR U2696 ( .A(n2708), .B(n2709), .Z(n2707) );
  OR U2697 ( .A(n2544), .B(n2543), .Z(n2548) );
  OR U2698 ( .A(n2546), .B(n2545), .Z(n2547) );
  NAND U2699 ( .A(n2548), .B(n2547), .Z(n2980) );
  NAND U2700 ( .A(n2550), .B(n2549), .Z(n2554) );
  NANDN U2701 ( .A(n2552), .B(n2551), .Z(n2553) );
  NAND U2702 ( .A(n2554), .B(n2553), .Z(n2979) );
  IV U2703 ( .A(n2979), .Z(n2978) );
  XNOR U2704 ( .A(n2980), .B(n2978), .Z(n2632) );
  NANDN U2705 ( .A(n2556), .B(n2555), .Z(n2560) );
  NANDN U2706 ( .A(n2558), .B(n2557), .Z(n2559) );
  AND U2707 ( .A(n2560), .B(n2559), .Z(n2973) );
  OR U2708 ( .A(n2562), .B(n2561), .Z(n2566) );
  NANDN U2709 ( .A(n2564), .B(n2563), .Z(n2565) );
  AND U2710 ( .A(n2566), .B(n2565), .Z(n2720) );
  OR U2711 ( .A(n2568), .B(n2567), .Z(n2572) );
  NANDN U2712 ( .A(n2570), .B(n2569), .Z(n2571) );
  AND U2713 ( .A(n2572), .B(n2571), .Z(n2721) );
  XOR U2714 ( .A(n2720), .B(n2721), .Z(n2718) );
  OR U2715 ( .A(n2574), .B(n2573), .Z(n2578) );
  OR U2716 ( .A(n2576), .B(n2575), .Z(n2577) );
  NAND U2717 ( .A(n2578), .B(n2577), .Z(n2739) );
  AND U2718 ( .A(y[26]), .B(x[4]), .Z(n2580) );
  NAND U2719 ( .A(x[3]), .B(y[27]), .Z(n2579) );
  XOR U2720 ( .A(n2580), .B(n2579), .Z(n2895) );
  AND U2721 ( .A(x[18]), .B(y[12]), .Z(n2894) );
  XNOR U2722 ( .A(n2895), .B(n2894), .Z(n2736) );
  AND U2723 ( .A(y[24]), .B(x[6]), .Z(n2582) );
  NAND U2724 ( .A(x[5]), .B(y[25]), .Z(n2581) );
  XOR U2725 ( .A(n2582), .B(n2581), .Z(n2847) );
  AND U2726 ( .A(x[19]), .B(y[11]), .Z(n2846) );
  XOR U2727 ( .A(n2847), .B(n2846), .Z(n2737) );
  XOR U2728 ( .A(n2736), .B(n2737), .Z(n2738) );
  XOR U2729 ( .A(n2739), .B(n2738), .Z(n2725) );
  XNOR U2730 ( .A(n2725), .B(n2724), .Z(n2727) );
  OR U2731 ( .A(n2587), .B(n2586), .Z(n2592) );
  NAND U2732 ( .A(o[28]), .B(n2588), .Z(n2590) );
  NAND U2733 ( .A(y[2]), .B(x[27]), .Z(n2589) );
  AND U2734 ( .A(n2590), .B(n2589), .Z(n2591) );
  ANDN U2735 ( .B(n2592), .A(n2591), .Z(n2726) );
  XNOR U2736 ( .A(n2727), .B(n2726), .Z(n2719) );
  XOR U2737 ( .A(n2718), .B(n2719), .Z(n2970) );
  OR U2738 ( .A(n2594), .B(n2593), .Z(n2598) );
  NANDN U2739 ( .A(n2596), .B(n2595), .Z(n2597) );
  NAND U2740 ( .A(n2598), .B(n2597), .Z(n2955) );
  NAND U2741 ( .A(x[20]), .B(y[10]), .Z(n2843) );
  AND U2742 ( .A(x[14]), .B(y[16]), .Z(n2842) );
  XOR U2743 ( .A(n2843), .B(n2842), .Z(n2841) );
  AND U2744 ( .A(y[22]), .B(x[8]), .Z(n2840) );
  XOR U2745 ( .A(n2841), .B(n2840), .Z(n2881) );
  NAND U2746 ( .A(y[0]), .B(x[30]), .Z(n2779) );
  NAND U2747 ( .A(y[1]), .B(x[29]), .Z(n2782) );
  XNOR U2748 ( .A(o[30]), .B(n2782), .Z(n2778) );
  XOR U2749 ( .A(n2779), .B(n2778), .Z(n2777) );
  AND U2750 ( .A(y[30]), .B(x[0]), .Z(n2776) );
  XNOR U2751 ( .A(n2777), .B(n2776), .Z(n2880) );
  XOR U2752 ( .A(n2879), .B(n2878), .Z(n2936) );
  NANDN U2753 ( .A(n2771), .B(n2602), .Z(n2606) );
  NAND U2754 ( .A(n2604), .B(n2603), .Z(n2605) );
  AND U2755 ( .A(n2606), .B(n2605), .Z(n2937) );
  XNOR U2756 ( .A(n2936), .B(n2937), .Z(n2935) );
  OR U2757 ( .A(n2608), .B(n2607), .Z(n2612) );
  OR U2758 ( .A(n2610), .B(n2609), .Z(n2611) );
  AND U2759 ( .A(n2612), .B(n2611), .Z(n2873) );
  NAND U2760 ( .A(x[17]), .B(y[13]), .Z(n2909) );
  NAND U2761 ( .A(x[2]), .B(y[28]), .Z(n2911) );
  NAND U2762 ( .A(y[4]), .B(x[26]), .Z(n2910) );
  XNOR U2763 ( .A(n2911), .B(n2910), .Z(n2908) );
  XNOR U2764 ( .A(n2909), .B(n2908), .Z(n2874) );
  NAND U2765 ( .A(y[23]), .B(x[7]), .Z(n2889) );
  AND U2766 ( .A(y[9]), .B(x[21]), .Z(n2614) );
  AND U2767 ( .A(x[22]), .B(y[8]), .Z(n2613) );
  XNOR U2768 ( .A(n2614), .B(n2613), .Z(n2888) );
  XOR U2769 ( .A(n2889), .B(n2888), .Z(n2875) );
  XNOR U2770 ( .A(n2874), .B(n2875), .Z(n2872) );
  XOR U2771 ( .A(n2873), .B(n2872), .Z(n2934) );
  XNOR U2772 ( .A(n2935), .B(n2934), .Z(n2954) );
  XOR U2773 ( .A(n2955), .B(n2954), .Z(n2953) );
  NANDN U2774 ( .A(n2616), .B(n2615), .Z(n2619) );
  OR U2775 ( .A(n2617), .B(n2836), .Z(n2618) );
  AND U2776 ( .A(n2619), .B(n2618), .Z(n2755) );
  NAND U2777 ( .A(n2623), .B(o[29]), .Z(n2903) );
  NAND U2778 ( .A(y[2]), .B(x[28]), .Z(n2905) );
  NAND U2779 ( .A(x[16]), .B(y[14]), .Z(n2904) );
  XNOR U2780 ( .A(n2905), .B(n2904), .Z(n2902) );
  XNOR U2781 ( .A(n2903), .B(n2902), .Z(n2731) );
  NAND U2782 ( .A(x[25]), .B(y[5]), .Z(n2770) );
  AND U2783 ( .A(y[6]), .B(x[24]), .Z(n2625) );
  NAND U2784 ( .A(y[7]), .B(x[23]), .Z(n2624) );
  XOR U2785 ( .A(n2625), .B(n2624), .Z(n2769) );
  XOR U2786 ( .A(n2770), .B(n2769), .Z(n2730) );
  XOR U2787 ( .A(n2731), .B(n2730), .Z(n2732) );
  XOR U2788 ( .A(n2733), .B(n2732), .Z(n2754) );
  NANDN U2789 ( .A(n2627), .B(n2626), .Z(n2631) );
  NANDN U2790 ( .A(n2629), .B(n2628), .Z(n2630) );
  AND U2791 ( .A(n2631), .B(n2630), .Z(n2752) );
  XOR U2792 ( .A(n2753), .B(n2752), .Z(n2952) );
  XNOR U2793 ( .A(n2953), .B(n2952), .Z(n2971) );
  XNOR U2794 ( .A(n2970), .B(n2971), .Z(n2972) );
  XNOR U2795 ( .A(n2973), .B(n2972), .Z(n2981) );
  XOR U2796 ( .A(n2632), .B(n2981), .Z(n2967) );
  OR U2797 ( .A(n2634), .B(n2633), .Z(n2638) );
  NANDN U2798 ( .A(n2636), .B(n2635), .Z(n2637) );
  AND U2799 ( .A(n2638), .B(n2637), .Z(n2965) );
  OR U2800 ( .A(n2640), .B(n2639), .Z(n2644) );
  NANDN U2801 ( .A(n2642), .B(n2641), .Z(n2643) );
  AND U2802 ( .A(n2644), .B(n2643), .Z(n2714) );
  OR U2803 ( .A(n2646), .B(n2645), .Z(n2650) );
  NANDN U2804 ( .A(n2648), .B(n2647), .Z(n2649) );
  AND U2805 ( .A(n2650), .B(n2649), .Z(n2715) );
  XOR U2806 ( .A(n2714), .B(n2715), .Z(n2712) );
  OR U2807 ( .A(n2652), .B(n2651), .Z(n2656) );
  OR U2808 ( .A(n2654), .B(n2653), .Z(n2655) );
  NAND U2809 ( .A(n2656), .B(n2655), .Z(n2713) );
  XNOR U2810 ( .A(n2712), .B(n2713), .Z(n2949) );
  NAND U2811 ( .A(y[3]), .B(x[27]), .Z(n2766) );
  AND U2812 ( .A(y[29]), .B(x[1]), .Z(n2765) );
  XNOR U2813 ( .A(n2766), .B(n2765), .Z(n2763) );
  AND U2814 ( .A(y[18]), .B(x[12]), .Z(n2661) );
  XOR U2815 ( .A(n2661), .B(n2660), .Z(n2835) );
  XNOR U2816 ( .A(n2835), .B(n2834), .Z(n2759) );
  AND U2817 ( .A(x[10]), .B(y[20]), .Z(n2663) );
  AND U2818 ( .A(y[21]), .B(x[9]), .Z(n2662) );
  XNOR U2819 ( .A(n2663), .B(n2662), .Z(n2758) );
  XOR U2820 ( .A(n2759), .B(n2758), .Z(n2746) );
  OR U2821 ( .A(n2665), .B(n2664), .Z(n2669) );
  OR U2822 ( .A(n2667), .B(n2666), .Z(n2668) );
  AND U2823 ( .A(n2669), .B(n2668), .Z(n2747) );
  XNOR U2824 ( .A(n2746), .B(n2747), .Z(n2745) );
  XOR U2825 ( .A(n2744), .B(n2745), .Z(n2930) );
  XNOR U2826 ( .A(n2931), .B(n2930), .Z(n2929) );
  OR U2827 ( .A(n2671), .B(n2670), .Z(n2675) );
  NANDN U2828 ( .A(n2673), .B(n2672), .Z(n2674) );
  NAND U2829 ( .A(n2675), .B(n2674), .Z(n2928) );
  XOR U2830 ( .A(n2929), .B(n2928), .Z(n2948) );
  XOR U2831 ( .A(n2949), .B(n2948), .Z(n2947) );
  OR U2832 ( .A(n2677), .B(n2676), .Z(n2681) );
  OR U2833 ( .A(n2679), .B(n2678), .Z(n2680) );
  NAND U2834 ( .A(n2681), .B(n2680), .Z(n2946) );
  XNOR U2835 ( .A(n2947), .B(n2946), .Z(n2964) );
  XNOR U2836 ( .A(n2965), .B(n2964), .Z(n2966) );
  XOR U2837 ( .A(n2967), .B(n2966), .Z(n2994) );
  OR U2838 ( .A(n2683), .B(n2682), .Z(n2687) );
  OR U2839 ( .A(n2685), .B(n2684), .Z(n2686) );
  NAND U2840 ( .A(n2687), .B(n2686), .Z(n3000) );
  NANDN U2841 ( .A(n2689), .B(n2688), .Z(n2693) );
  OR U2842 ( .A(n2691), .B(n2690), .Z(n2692) );
  AND U2843 ( .A(n2693), .B(n2692), .Z(n2999) );
  XOR U2844 ( .A(n3000), .B(n2999), .Z(n2997) );
  OR U2845 ( .A(n2695), .B(n2694), .Z(n2699) );
  NANDN U2846 ( .A(n2697), .B(n2696), .Z(n2698) );
  AND U2847 ( .A(n2699), .B(n2698), .Z(n2998) );
  XOR U2848 ( .A(n2994), .B(n2993), .Z(n2992) );
  OR U2849 ( .A(n2701), .B(n2700), .Z(n2705) );
  NANDN U2850 ( .A(n2703), .B(n2702), .Z(n2704) );
  NAND U2851 ( .A(n2705), .B(n2704), .Z(n2991) );
  XOR U2852 ( .A(n2992), .B(n2991), .Z(n2706) );
  XNOR U2853 ( .A(n2707), .B(n2706), .Z(N63) );
  OR U2854 ( .A(n2707), .B(n2706), .Z(n2711) );
  OR U2855 ( .A(n2709), .B(n2708), .Z(n2710) );
  AND U2856 ( .A(n2711), .B(n2710), .Z(n2990) );
  NANDN U2857 ( .A(n2713), .B(n2712), .Z(n2717) );
  OR U2858 ( .A(n2715), .B(n2714), .Z(n2716) );
  AND U2859 ( .A(n2717), .B(n2716), .Z(n2963) );
  NANDN U2860 ( .A(n2719), .B(n2718), .Z(n2723) );
  OR U2861 ( .A(n2721), .B(n2720), .Z(n2722) );
  AND U2862 ( .A(n2723), .B(n2722), .Z(n2945) );
  NOR U2863 ( .A(n2725), .B(n2724), .Z(n2729) );
  NOR U2864 ( .A(n2727), .B(n2726), .Z(n2728) );
  NOR U2865 ( .A(n2729), .B(n2728), .Z(n2927) );
  ANDN U2866 ( .B(n2731), .A(n2730), .Z(n2735) );
  NOR U2867 ( .A(n2733), .B(n2732), .Z(n2734) );
  NOR U2868 ( .A(n2735), .B(n2734), .Z(n2743) );
  NANDN U2869 ( .A(n2737), .B(n2736), .Z(n2741) );
  OR U2870 ( .A(n2739), .B(n2738), .Z(n2740) );
  AND U2871 ( .A(n2741), .B(n2740), .Z(n2742) );
  XNOR U2872 ( .A(n2743), .B(n2742), .Z(n2751) );
  OR U2873 ( .A(n2745), .B(n2744), .Z(n2749) );
  OR U2874 ( .A(n2747), .B(n2746), .Z(n2748) );
  NAND U2875 ( .A(n2749), .B(n2748), .Z(n2750) );
  XNOR U2876 ( .A(n2751), .B(n2750), .Z(n2925) );
  OR U2877 ( .A(n2753), .B(n2752), .Z(n2757) );
  NANDN U2878 ( .A(n2755), .B(n2754), .Z(n2756) );
  AND U2879 ( .A(n2757), .B(n2756), .Z(n2923) );
  OR U2880 ( .A(n2759), .B(n2758), .Z(n2762) );
  NAND U2881 ( .A(y[21]), .B(x[10]), .Z(n2794) );
  NANDN U2882 ( .A(n2794), .B(n2760), .Z(n2761) );
  AND U2883 ( .A(n2762), .B(n2761), .Z(n2833) );
  NANDN U2884 ( .A(n2764), .B(n2763), .Z(n2768) );
  NANDN U2885 ( .A(n2766), .B(n2765), .Z(n2767) );
  AND U2886 ( .A(n2768), .B(n2767), .Z(n2775) );
  OR U2887 ( .A(n2770), .B(n2769), .Z(n2773) );
  NAND U2888 ( .A(y[7]), .B(x[24]), .Z(n2799) );
  NANDN U2889 ( .A(n2799), .B(n2771), .Z(n2772) );
  NAND U2890 ( .A(n2773), .B(n2772), .Z(n2774) );
  XNOR U2891 ( .A(n2775), .B(n2774), .Z(n2831) );
  NANDN U2892 ( .A(n2777), .B(n2776), .Z(n2781) );
  NANDN U2893 ( .A(n2779), .B(n2778), .Z(n2780) );
  AND U2894 ( .A(n2781), .B(n2780), .Z(n2829) );
  AND U2895 ( .A(x[21]), .B(y[10]), .Z(n2788) );
  ANDN U2896 ( .B(o[30]), .A(n2782), .Z(n2786) );
  NAND U2897 ( .A(y[9]), .B(x[22]), .Z(n2891) );
  XNOR U2898 ( .A(n2891), .B(o[31]), .Z(n2784) );
  NAND U2899 ( .A(x[4]), .B(y[27]), .Z(n2897) );
  NAND U2900 ( .A(x[6]), .B(y[25]), .Z(n2849) );
  XNOR U2901 ( .A(n2897), .B(n2849), .Z(n2783) );
  XNOR U2902 ( .A(n2784), .B(n2783), .Z(n2785) );
  XNOR U2903 ( .A(n2786), .B(n2785), .Z(n2787) );
  XNOR U2904 ( .A(n2788), .B(n2787), .Z(n2827) );
  AND U2905 ( .A(y[29]), .B(x[2]), .Z(n2790) );
  NAND U2906 ( .A(y[1]), .B(x[30]), .Z(n2789) );
  XNOR U2907 ( .A(n2790), .B(n2789), .Z(n2798) );
  AND U2908 ( .A(x[27]), .B(y[4]), .Z(n2796) );
  AND U2909 ( .A(x[17]), .B(y[14]), .Z(n2792) );
  NAND U2910 ( .A(y[8]), .B(x[23]), .Z(n2791) );
  XNOR U2911 ( .A(n2792), .B(n2791), .Z(n2793) );
  XOR U2912 ( .A(n2794), .B(n2793), .Z(n2795) );
  XNOR U2913 ( .A(n2796), .B(n2795), .Z(n2797) );
  XOR U2914 ( .A(n2798), .B(n2797), .Z(n2801) );
  NAND U2915 ( .A(x[13]), .B(y[18]), .Z(n2837) );
  XNOR U2916 ( .A(n2799), .B(n2837), .Z(n2800) );
  XNOR U2917 ( .A(n2801), .B(n2800), .Z(n2817) );
  AND U2918 ( .A(y[22]), .B(x[9]), .Z(n2803) );
  NAND U2919 ( .A(x[25]), .B(y[6]), .Z(n2802) );
  XNOR U2920 ( .A(n2803), .B(n2802), .Z(n2807) );
  AND U2921 ( .A(y[16]), .B(x[15]), .Z(n2805) );
  NAND U2922 ( .A(x[0]), .B(y[31]), .Z(n2804) );
  XNOR U2923 ( .A(n2805), .B(n2804), .Z(n2806) );
  XOR U2924 ( .A(n2807), .B(n2806), .Z(n2815) );
  AND U2925 ( .A(y[15]), .B(x[16]), .Z(n2809) );
  NAND U2926 ( .A(y[2]), .B(x[29]), .Z(n2808) );
  XNOR U2927 ( .A(n2809), .B(n2808), .Z(n2813) );
  AND U2928 ( .A(y[17]), .B(x[14]), .Z(n2811) );
  NAND U2929 ( .A(x[20]), .B(y[11]), .Z(n2810) );
  XNOR U2930 ( .A(n2811), .B(n2810), .Z(n2812) );
  XNOR U2931 ( .A(n2813), .B(n2812), .Z(n2814) );
  XNOR U2932 ( .A(n2815), .B(n2814), .Z(n2816) );
  XOR U2933 ( .A(n2817), .B(n2816), .Z(n2825) );
  AND U2934 ( .A(x[19]), .B(y[12]), .Z(n2819) );
  NAND U2935 ( .A(y[23]), .B(x[8]), .Z(n2818) );
  XNOR U2936 ( .A(n2819), .B(n2818), .Z(n2823) );
  AND U2937 ( .A(y[24]), .B(x[7]), .Z(n2821) );
  NAND U2938 ( .A(x[5]), .B(y[26]), .Z(n2820) );
  XNOR U2939 ( .A(n2821), .B(n2820), .Z(n2822) );
  XNOR U2940 ( .A(n2823), .B(n2822), .Z(n2824) );
  XNOR U2941 ( .A(n2825), .B(n2824), .Z(n2826) );
  XNOR U2942 ( .A(n2827), .B(n2826), .Z(n2828) );
  XNOR U2943 ( .A(n2829), .B(n2828), .Z(n2830) );
  XNOR U2944 ( .A(n2831), .B(n2830), .Z(n2832) );
  XNOR U2945 ( .A(n2833), .B(n2832), .Z(n2921) );
  OR U2946 ( .A(n2835), .B(n2834), .Z(n2839) );
  NANDN U2947 ( .A(n2837), .B(n2836), .Z(n2838) );
  AND U2948 ( .A(n2839), .B(n2838), .Z(n2871) );
  NANDN U2949 ( .A(n2841), .B(n2840), .Z(n2845) );
  NANDN U2950 ( .A(n2843), .B(n2842), .Z(n2844) );
  AND U2951 ( .A(n2845), .B(n2844), .Z(n2853) );
  NANDN U2952 ( .A(n2847), .B(n2846), .Z(n2851) );
  NANDN U2953 ( .A(n2849), .B(n2848), .Z(n2850) );
  NAND U2954 ( .A(n2851), .B(n2850), .Z(n2852) );
  XNOR U2955 ( .A(n2853), .B(n2852), .Z(n2869) );
  AND U2956 ( .A(y[20]), .B(x[11]), .Z(n2855) );
  NAND U2957 ( .A(y[19]), .B(x[12]), .Z(n2854) );
  XNOR U2958 ( .A(n2855), .B(n2854), .Z(n2859) );
  AND U2959 ( .A(y[30]), .B(x[1]), .Z(n2857) );
  NAND U2960 ( .A(y[3]), .B(x[28]), .Z(n2856) );
  XNOR U2961 ( .A(n2857), .B(n2856), .Z(n2858) );
  XOR U2962 ( .A(n2859), .B(n2858), .Z(n2867) );
  AND U2963 ( .A(x[18]), .B(y[13]), .Z(n2861) );
  NAND U2964 ( .A(y[5]), .B(x[26]), .Z(n2860) );
  XNOR U2965 ( .A(n2861), .B(n2860), .Z(n2865) );
  AND U2966 ( .A(x[31]), .B(y[0]), .Z(n2863) );
  NAND U2967 ( .A(x[3]), .B(y[28]), .Z(n2862) );
  XNOR U2968 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U2969 ( .A(n2865), .B(n2864), .Z(n2866) );
  XNOR U2970 ( .A(n2867), .B(n2866), .Z(n2868) );
  XNOR U2971 ( .A(n2869), .B(n2868), .Z(n2870) );
  XNOR U2972 ( .A(n2871), .B(n2870), .Z(n2887) );
  NANDN U2973 ( .A(n2873), .B(n2872), .Z(n2877) );
  NANDN U2974 ( .A(n2875), .B(n2874), .Z(n2876) );
  AND U2975 ( .A(n2877), .B(n2876), .Z(n2885) );
  OR U2976 ( .A(n2879), .B(n2878), .Z(n2883) );
  NANDN U2977 ( .A(n2881), .B(n2880), .Z(n2882) );
  NAND U2978 ( .A(n2883), .B(n2882), .Z(n2884) );
  XNOR U2979 ( .A(n2885), .B(n2884), .Z(n2886) );
  XOR U2980 ( .A(n2887), .B(n2886), .Z(n2919) );
  OR U2981 ( .A(n2889), .B(n2888), .Z(n2893) );
  NANDN U2982 ( .A(n2891), .B(n2890), .Z(n2892) );
  AND U2983 ( .A(n2893), .B(n2892), .Z(n2901) );
  NANDN U2984 ( .A(n2895), .B(n2894), .Z(n2899) );
  NANDN U2985 ( .A(n2897), .B(n2896), .Z(n2898) );
  NAND U2986 ( .A(n2899), .B(n2898), .Z(n2900) );
  XNOR U2987 ( .A(n2901), .B(n2900), .Z(n2917) );
  OR U2988 ( .A(n2903), .B(n2902), .Z(n2907) );
  OR U2989 ( .A(n2905), .B(n2904), .Z(n2906) );
  AND U2990 ( .A(n2907), .B(n2906), .Z(n2915) );
  OR U2991 ( .A(n2909), .B(n2908), .Z(n2913) );
  OR U2992 ( .A(n2911), .B(n2910), .Z(n2912) );
  NAND U2993 ( .A(n2913), .B(n2912), .Z(n2914) );
  XNOR U2994 ( .A(n2915), .B(n2914), .Z(n2916) );
  XNOR U2995 ( .A(n2917), .B(n2916), .Z(n2918) );
  XNOR U2996 ( .A(n2919), .B(n2918), .Z(n2920) );
  XNOR U2997 ( .A(n2921), .B(n2920), .Z(n2922) );
  XNOR U2998 ( .A(n2923), .B(n2922), .Z(n2924) );
  XOR U2999 ( .A(n2925), .B(n2924), .Z(n2926) );
  XNOR U3000 ( .A(n2927), .B(n2926), .Z(n2943) );
  OR U3001 ( .A(n2929), .B(n2928), .Z(n2933) );
  OR U3002 ( .A(n2931), .B(n2930), .Z(n2932) );
  AND U3003 ( .A(n2933), .B(n2932), .Z(n2941) );
  OR U3004 ( .A(n2935), .B(n2934), .Z(n2939) );
  OR U3005 ( .A(n2937), .B(n2936), .Z(n2938) );
  NAND U3006 ( .A(n2939), .B(n2938), .Z(n2940) );
  XNOR U3007 ( .A(n2941), .B(n2940), .Z(n2942) );
  XNOR U3008 ( .A(n2943), .B(n2942), .Z(n2944) );
  XNOR U3009 ( .A(n2945), .B(n2944), .Z(n2961) );
  OR U3010 ( .A(n2947), .B(n2946), .Z(n2951) );
  NANDN U3011 ( .A(n2949), .B(n2948), .Z(n2950) );
  AND U3012 ( .A(n2951), .B(n2950), .Z(n2959) );
  OR U3013 ( .A(n2953), .B(n2952), .Z(n2957) );
  NANDN U3014 ( .A(n2955), .B(n2954), .Z(n2956) );
  NAND U3015 ( .A(n2957), .B(n2956), .Z(n2958) );
  XNOR U3016 ( .A(n2959), .B(n2958), .Z(n2960) );
  XNOR U3017 ( .A(n2961), .B(n2960), .Z(n2962) );
  XNOR U3018 ( .A(n2963), .B(n2962), .Z(n2988) );
  NOR U3019 ( .A(n2965), .B(n2964), .Z(n2969) );
  ANDN U3020 ( .B(n2967), .A(n2966), .Z(n2968) );
  NOR U3021 ( .A(n2969), .B(n2968), .Z(n2977) );
  NANDN U3022 ( .A(n2971), .B(n2970), .Z(n2975) );
  NANDN U3023 ( .A(n2973), .B(n2972), .Z(n2974) );
  AND U3024 ( .A(n2975), .B(n2974), .Z(n2976) );
  XNOR U3025 ( .A(n2977), .B(n2976), .Z(n2986) );
  NANDN U3026 ( .A(n2980), .B(n2978), .Z(n2984) );
  XOR U3027 ( .A(n2980), .B(n2979), .Z(n2982) );
  NAND U3028 ( .A(n2982), .B(n2981), .Z(n2983) );
  AND U3029 ( .A(n2984), .B(n2983), .Z(n2985) );
  XNOR U3030 ( .A(n2986), .B(n2985), .Z(n2987) );
  XNOR U3031 ( .A(n2988), .B(n2987), .Z(n2989) );
  XNOR U3032 ( .A(n2990), .B(n2989), .Z(n3006) );
  OR U3033 ( .A(n2992), .B(n2991), .Z(n2996) );
  NANDN U3034 ( .A(n2994), .B(n2993), .Z(n2995) );
  AND U3035 ( .A(n2996), .B(n2995), .Z(n3004) );
  NANDN U3036 ( .A(n2998), .B(n2997), .Z(n3002) );
  OR U3037 ( .A(n3000), .B(n2999), .Z(n3001) );
  NAND U3038 ( .A(n3002), .B(n3001), .Z(n3003) );
  XNOR U3039 ( .A(n3004), .B(n3003), .Z(n3005) );
  XNOR U3040 ( .A(n3006), .B(n3005), .Z(N64) );
endmodule

