
module first_nns_comb_W15_N256 ( q, DB, min_val_out );
  input [14:0] q;
  input [3839:0] DB;
  output [14:0] min_val_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297,
         n36298, n36299, n36300, n36301, n36302, n36303, n36304, n36305,
         n36306, n36307, n36308, n36309, n36310, n36311, n36312, n36313,
         n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321,
         n36322, n36323, n36324, n36325, n36326, n36327, n36328, n36329,
         n36330, n36331, n36332, n36333, n36334, n36335, n36336, n36337,
         n36338, n36339, n36340, n36341, n36342, n36343, n36344, n36345,
         n36346, n36347, n36348, n36349, n36350, n36351, n36352, n36353,
         n36354, n36355, n36356, n36357, n36358, n36359, n36360, n36361,
         n36362, n36363, n36364, n36365, n36366, n36367, n36368, n36369,
         n36370, n36371, n36372, n36373, n36374, n36375, n36376, n36377,
         n36378, n36379, n36380, n36381, n36382, n36383, n36384, n36385,
         n36386, n36387, n36388, n36389, n36390, n36391, n36392, n36393,
         n36394, n36395, n36396, n36397, n36398, n36399, n36400, n36401,
         n36402, n36403, n36404, n36405, n36406, n36407, n36408, n36409,
         n36410, n36411, n36412, n36413, n36414, n36415, n36416, n36417,
         n36418, n36419, n36420, n36421, n36422, n36423, n36424, n36425,
         n36426, n36427, n36428, n36429, n36430, n36431, n36432, n36433,
         n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
         n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449,
         n36450, n36451, n36452, n36453, n36454, n36455, n36456, n36457,
         n36458, n36459, n36460, n36461, n36462, n36463, n36464, n36465,
         n36466, n36467, n36468, n36469, n36470, n36471, n36472, n36473,
         n36474, n36475, n36476, n36477, n36478, n36479, n36480, n36481,
         n36482, n36483, n36484, n36485, n36486, n36487, n36488, n36489,
         n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497,
         n36498, n36499, n36500, n36501, n36502, n36503, n36504, n36505,
         n36506, n36507, n36508, n36509, n36510, n36511, n36512, n36513,
         n36514, n36515, n36516, n36517, n36518, n36519, n36520, n36521,
         n36522, n36523, n36524, n36525, n36526, n36527, n36528, n36529,
         n36530, n36531, n36532, n36533, n36534, n36535, n36536, n36537,
         n36538, n36539, n36540, n36541, n36542, n36543, n36544, n36545,
         n36546, n36547, n36548, n36549, n36550, n36551, n36552, n36553,
         n36554, n36555, n36556, n36557, n36558, n36559, n36560, n36561,
         n36562, n36563, n36564, n36565, n36566, n36567, n36568, n36569,
         n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
         n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585,
         n36586, n36587, n36588, n36589, n36590, n36591, n36592, n36593,
         n36594, n36595, n36596, n36597, n36598, n36599, n36600, n36601,
         n36602, n36603, n36604, n36605, n36606, n36607, n36608, n36609,
         n36610, n36611, n36612, n36613, n36614, n36615, n36616, n36617,
         n36618, n36619, n36620, n36621, n36622, n36623, n36624, n36625,
         n36626, n36627, n36628, n36629, n36630, n36631, n36632, n36633,
         n36634, n36635, n36636, n36637, n36638, n36639, n36640, n36641,
         n36642, n36643, n36644, n36645, n36646, n36647, n36648, n36649,
         n36650, n36651, n36652, n36653, n36654, n36655, n36656, n36657,
         n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36665,
         n36666, n36667, n36668, n36669, n36670, n36671, n36672, n36673,
         n36674, n36675, n36676, n36677, n36678, n36679, n36680, n36681,
         n36682, n36683, n36684, n36685, n36686, n36687, n36688, n36689,
         n36690, n36691, n36692, n36693, n36694, n36695, n36696, n36697,
         n36698, n36699, n36700, n36701, n36702, n36703, n36704, n36705,
         n36706, n36707, n36708, n36709, n36710, n36711, n36712, n36713,
         n36714, n36715, n36716, n36717, n36718, n36719, n36720, n36721,
         n36722, n36723, n36724, n36725, n36726, n36727, n36728, n36729,
         n36730, n36731, n36732, n36733, n36734, n36735, n36736, n36737,
         n36738, n36739, n36740, n36741, n36742, n36743, n36744, n36745,
         n36746, n36747, n36748, n36749, n36750, n36751, n36752, n36753,
         n36754, n36755, n36756, n36757, n36758, n36759, n36760, n36761,
         n36762, n36763, n36764, n36765, n36766, n36767, n36768, n36769,
         n36770, n36771, n36772, n36773, n36774, n36775, n36776, n36777,
         n36778, n36779, n36780, n36781, n36782, n36783, n36784, n36785,
         n36786, n36787, n36788, n36789, n36790, n36791, n36792, n36793,
         n36794, n36795, n36796, n36797, n36798, n36799, n36800, n36801,
         n36802, n36803, n36804, n36805, n36806, n36807, n36808, n36809,
         n36810, n36811, n36812, n36813, n36814, n36815, n36816, n36817,
         n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
         n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833,
         n36834, n36835, n36836, n36837, n36838, n36839, n36840, n36841,
         n36842, n36843, n36844, n36845, n36846, n36847, n36848, n36849,
         n36850, n36851, n36852, n36853, n36854, n36855, n36856, n36857,
         n36858, n36859, n36860, n36861, n36862, n36863, n36864, n36865,
         n36866, n36867, n36868, n36869, n36870, n36871, n36872, n36873,
         n36874, n36875, n36876, n36877, n36878, n36879, n36880, n36881,
         n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
         n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897,
         n36898, n36899, n36900, n36901, n36902, n36903, n36904, n36905,
         n36906, n36907, n36908, n36909, n36910, n36911, n36912, n36913,
         n36914, n36915, n36916, n36917, n36918, n36919, n36920, n36921,
         n36922, n36923, n36924, n36925, n36926, n36927, n36928, n36929,
         n36930, n36931, n36932, n36933, n36934, n36935, n36936, n36937,
         n36938, n36939, n36940, n36941, n36942, n36943, n36944, n36945,
         n36946, n36947, n36948, n36949, n36950, n36951, n36952, n36953,
         n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
         n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969,
         n36970, n36971, n36972, n36973, n36974, n36975, n36976, n36977,
         n36978, n36979, n36980, n36981, n36982, n36983, n36984, n36985,
         n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
         n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001,
         n37002, n37003, n37004, n37005, n37006, n37007, n37008, n37009,
         n37010, n37011, n37012, n37013, n37014, n37015, n37016, n37017,
         n37018, n37019, n37020, n37021, n37022, n37023, n37024, n37025,
         n37026, n37027, n37028, n37029, n37030, n37031, n37032, n37033,
         n37034, n37035, n37036, n37037, n37038, n37039, n37040, n37041,
         n37042, n37043, n37044, n37045, n37046, n37047, n37048, n37049,
         n37050, n37051, n37052, n37053, n37054, n37055, n37056, n37057,
         n37058, n37059, n37060, n37061, n37062, n37063, n37064, n37065,
         n37066, n37067, n37068, n37069, n37070, n37071, n37072, n37073,
         n37074, n37075, n37076, n37077, n37078, n37079, n37080, n37081,
         n37082, n37083, n37084, n37085, n37086, n37087, n37088, n37089,
         n37090, n37091, n37092, n37093, n37094, n37095, n37096, n37097,
         n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
         n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113,
         n37114, n37115, n37116, n37117, n37118, n37119, n37120, n37121,
         n37122, n37123, n37124, n37125, n37126, n37127, n37128, n37129,
         n37130, n37131, n37132, n37133, n37134, n37135, n37136, n37137,
         n37138, n37139, n37140, n37141, n37142, n37143, n37144, n37145,
         n37146, n37147, n37148, n37149, n37150, n37151, n37152, n37153,
         n37154, n37155, n37156, n37157, n37158, n37159, n37160, n37161,
         n37162, n37163, n37164, n37165, n37166, n37167, n37168, n37169,
         n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
         n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185,
         n37186, n37187, n37188, n37189, n37190, n37191, n37192, n37193,
         n37194, n37195, n37196, n37197, n37198, n37199, n37200, n37201,
         n37202, n37203, n37204, n37205, n37206, n37207, n37208, n37209,
         n37210, n37211, n37212, n37213, n37214, n37215, n37216, n37217,
         n37218, n37219, n37220, n37221, n37222, n37223, n37224, n37225,
         n37226, n37227, n37228, n37229, n37230, n37231, n37232, n37233,
         n37234, n37235, n37236, n37237, n37238, n37239, n37240, n37241,
         n37242, n37243, n37244, n37245, n37246, n37247, n37248, n37249,
         n37250, n37251, n37252, n37253, n37254, n37255, n37256, n37257,
         n37258, n37259, n37260, n37261, n37262, n37263, n37264, n37265,
         n37266, n37267, n37268, n37269, n37270, n37271, n37272, n37273,
         n37274, n37275, n37276, n37277, n37278, n37279, n37280, n37281,
         n37282, n37283, n37284, n37285, n37286, n37287, n37288, n37289,
         n37290, n37291, n37292, n37293, n37294, n37295, n37296, n37297,
         n37298, n37299, n37300, n37301, n37302, n37303, n37304, n37305,
         n37306, n37307, n37308, n37309, n37310, n37311, n37312, n37313,
         n37314, n37315, n37316, n37317, n37318, n37319, n37320, n37321,
         n37322, n37323, n37324, n37325, n37326, n37327, n37328, n37329,
         n37330, n37331, n37332, n37333, n37334, n37335, n37336, n37337,
         n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
         n37346, n37347, n37348, n37349, n37350, n37351, n37352, n37353,
         n37354, n37355, n37356, n37357, n37358, n37359, n37360, n37361,
         n37362, n37363, n37364, n37365, n37366, n37367, n37368, n37369,
         n37370, n37371, n37372, n37373, n37374, n37375, n37376, n37377,
         n37378, n37379, n37380, n37381, n37382, n37383, n37384, n37385,
         n37386, n37387, n37388, n37389, n37390, n37391, n37392, n37393,
         n37394, n37395, n37396, n37397, n37398, n37399, n37400, n37401,
         n37402, n37403, n37404, n37405, n37406, n37407, n37408, n37409,
         n37410, n37411, n37412, n37413, n37414, n37415, n37416, n37417,
         n37418, n37419, n37420, n37421, n37422, n37423, n37424, n37425,
         n37426, n37427, n37428, n37429, n37430, n37431, n37432, n37433,
         n37434, n37435, n37436, n37437, n37438, n37439, n37440, n37441,
         n37442, n37443, n37444, n37445, n37446, n37447, n37448, n37449,
         n37450, n37451, n37452, n37453, n37454, n37455, n37456, n37457,
         n37458, n37459, n37460, n37461, n37462, n37463, n37464, n37465,
         n37466, n37467, n37468, n37469, n37470, n37471, n37472, n37473,
         n37474, n37475, n37476, n37477, n37478, n37479, n37480, n37481,
         n37482, n37483, n37484, n37485, n37486, n37487, n37488, n37489,
         n37490, n37491, n37492, n37493, n37494, n37495, n37496, n37497,
         n37498, n37499, n37500, n37501, n37502, n37503, n37504, n37505,
         n37506, n37507, n37508, n37509, n37510, n37511, n37512, n37513,
         n37514, n37515, n37516, n37517, n37518, n37519, n37520, n37521,
         n37522, n37523, n37524, n37525, n37526, n37527, n37528, n37529,
         n37530, n37531, n37532, n37533, n37534, n37535, n37536, n37537,
         n37538, n37539, n37540, n37541, n37542, n37543, n37544, n37545,
         n37546, n37547, n37548, n37549, n37550, n37551, n37552, n37553,
         n37554, n37555, n37556, n37557, n37558, n37559, n37560, n37561,
         n37562, n37563, n37564, n37565, n37566, n37567, n37568, n37569,
         n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577,
         n37578, n37579, n37580, n37581, n37582, n37583, n37584, n37585,
         n37586, n37587, n37588, n37589, n37590, n37591, n37592, n37593,
         n37594, n37595, n37596, n37597, n37598, n37599, n37600, n37601,
         n37602, n37603, n37604, n37605, n37606, n37607, n37608, n37609,
         n37610, n37611, n37612, n37613, n37614, n37615, n37616, n37617,
         n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
         n37626, n37627, n37628, n37629, n37630, n37631, n37632, n37633,
         n37634, n37635, n37636, n37637, n37638, n37639, n37640, n37641,
         n37642, n37643, n37644, n37645, n37646, n37647, n37648, n37649,
         n37650, n37651, n37652, n37653, n37654, n37655, n37656, n37657,
         n37658, n37659, n37660, n37661, n37662, n37663, n37664, n37665,
         n37666, n37667, n37668, n37669, n37670, n37671, n37672, n37673,
         n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
         n37682, n37683, n37684, n37685, n37686, n37687, n37688, n37689,
         n37690, n37691, n37692, n37693, n37694, n37695, n37696, n37697,
         n37698, n37699, n37700, n37701, n37702, n37703, n37704, n37705,
         n37706, n37707, n37708, n37709, n37710, n37711, n37712, n37713,
         n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
         n37722, n37723, n37724, n37725, n37726, n37727, n37728, n37729,
         n37730, n37731, n37732, n37733, n37734, n37735, n37736, n37737,
         n37738, n37739, n37740, n37741, n37742, n37743, n37744, n37745,
         n37746, n37747, n37748, n37749, n37750, n37751, n37752, n37753,
         n37754, n37755, n37756, n37757, n37758, n37759, n37760, n37761,
         n37762, n37763, n37764, n37765, n37766, n37767, n37768, n37769,
         n37770, n37771, n37772, n37773, n37774, n37775, n37776, n37777,
         n37778, n37779, n37780, n37781, n37782, n37783, n37784, n37785,
         n37786, n37787, n37788, n37789, n37790, n37791, n37792, n37793,
         n37794, n37795, n37796, n37797, n37798, n37799, n37800, n37801,
         n37802, n37803, n37804, n37805, n37806, n37807, n37808, n37809,
         n37810, n37811, n37812, n37813, n37814, n37815, n37816, n37817,
         n37818, n37819, n37820, n37821, n37822, n37823, n37824, n37825,
         n37826, n37827, n37828, n37829, n37830, n37831, n37832, n37833,
         n37834, n37835, n37836, n37837, n37838, n37839, n37840, n37841,
         n37842, n37843, n37844, n37845, n37846, n37847, n37848, n37849,
         n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
         n37858, n37859, n37860, n37861, n37862, n37863, n37864, n37865,
         n37866, n37867, n37868, n37869, n37870, n37871, n37872, n37873,
         n37874, n37875, n37876, n37877, n37878, n37879, n37880, n37881,
         n37882, n37883, n37884, n37885, n37886, n37887, n37888, n37889,
         n37890, n37891, n37892, n37893, n37894, n37895, n37896, n37897,
         n37898, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
         n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913,
         n37914, n37915, n37916, n37917, n37918, n37919, n37920, n37921,
         n37922, n37923, n37924, n37925, n37926, n37927, n37928, n37929,
         n37930, n37931, n37932, n37933, n37934, n37935, n37936, n37937,
         n37938, n37939, n37940, n37941, n37942, n37943, n37944, n37945,
         n37946, n37947, n37948, n37949, n37950, n37951, n37952, n37953,
         n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961,
         n37962, n37963, n37964, n37965, n37966, n37967, n37968, n37969,
         n37970, n37971, n37972, n37973, n37974, n37975, n37976, n37977,
         n37978, n37979, n37980, n37981, n37982, n37983, n37984, n37985,
         n37986, n37987, n37988, n37989, n37990, n37991, n37992, n37993,
         n37994, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
         n38002, n38003, n38004, n38005, n38006, n38007, n38008, n38009,
         n38010, n38011, n38012, n38013, n38014, n38015, n38016, n38017,
         n38018, n38019, n38020, n38021, n38022, n38023, n38024, n38025,
         n38026, n38027, n38028, n38029, n38030, n38031, n38032, n38033,
         n38034, n38035, n38036, n38037, n38038, n38039, n38040, n38041,
         n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
         n38050, n38051, n38052, n38053, n38054, n38055, n38056, n38057,
         n38058, n38059, n38060, n38061, n38062, n38063, n38064, n38065,
         n38066, n38067, n38068, n38069, n38070, n38071, n38072, n38073,
         n38074, n38075, n38076, n38077, n38078, n38079, n38080, n38081,
         n38082, n38083, n38084, n38085, n38086, n38087, n38088, n38089,
         n38090, n38091, n38092, n38093, n38094, n38095, n38096, n38097,
         n38098, n38099, n38100, n38101, n38102, n38103, n38104, n38105,
         n38106, n38107, n38108, n38109, n38110, n38111, n38112, n38113,
         n38114, n38115, n38116, n38117, n38118, n38119, n38120, n38121,
         n38122, n38123, n38124, n38125, n38126, n38127, n38128, n38129,
         n38130, n38131, n38132, n38133, n38134, n38135, n38136, n38137,
         n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
         n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38153,
         n38154, n38155, n38156, n38157, n38158, n38159, n38160, n38161,
         n38162, n38163, n38164, n38165, n38166, n38167, n38168, n38169,
         n38170, n38171, n38172, n38173, n38174, n38175, n38176, n38177,
         n38178, n38179, n38180, n38181, n38182, n38183, n38184, n38185,
         n38186, n38187, n38188, n38189, n38190, n38191, n38192, n38193,
         n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201,
         n38202, n38203, n38204, n38205, n38206, n38207, n38208, n38209,
         n38210, n38211, n38212, n38213, n38214, n38215, n38216, n38217,
         n38218, n38219, n38220, n38221, n38222, n38223, n38224, n38225,
         n38226, n38227, n38228, n38229, n38230, n38231, n38232, n38233,
         n38234, n38235, n38236, n38237, n38238, n38239, n38240, n38241,
         n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
         n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257,
         n38258, n38259, n38260, n38261, n38262, n38263, n38264, n38265,
         n38266, n38267, n38268, n38269, n38270, n38271, n38272, n38273,
         n38274, n38275, n38276, n38277, n38278, n38279, n38280, n38281,
         n38282, n38283, n38284, n38285, n38286, n38287, n38288, n38289,
         n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
         n38298, n38299, n38300, n38301, n38302, n38303, n38304, n38305,
         n38306, n38307, n38308, n38309, n38310, n38311, n38312, n38313,
         n38314, n38315, n38316, n38317, n38318, n38319, n38320, n38321,
         n38322, n38323, n38324, n38325, n38326, n38327, n38328, n38329,
         n38330, n38331, n38332, n38333, n38334, n38335, n38336, n38337,
         n38338, n38339, n38340, n38341, n38342, n38343, n38344, n38345,
         n38346, n38347, n38348, n38349, n38350, n38351, n38352, n38353,
         n38354, n38355, n38356, n38357, n38358, n38359, n38360, n38361,
         n38362, n38363, n38364, n38365, n38366, n38367, n38368, n38369,
         n38370, n38371, n38372, n38373, n38374, n38375, n38376, n38377,
         n38378, n38379, n38380, n38381, n38382, n38383, n38384, n38385,
         n38386, n38387, n38388, n38389, n38390, n38391, n38392, n38393,
         n38394, n38395, n38396, n38397, n38398, n38399, n38400, n38401,
         n38402, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
         n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417,
         n38418, n38419, n38420, n38421, n38422, n38423, n38424, n38425,
         n38426, n38427, n38428, n38429, n38430, n38431, n38432, n38433,
         n38434, n38435, n38436, n38437, n38438, n38439, n38440, n38441,
         n38442, n38443, n38444, n38445, n38446, n38447, n38448, n38449,
         n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
         n38458, n38459, n38460, n38461, n38462, n38463, n38464, n38465,
         n38466, n38467, n38468, n38469, n38470, n38471, n38472, n38473,
         n38474, n38475, n38476, n38477, n38478, n38479, n38480, n38481,
         n38482, n38483, n38484, n38485, n38486, n38487, n38488, n38489,
         n38490, n38491, n38492, n38493, n38494, n38495, n38496, n38497,
         n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505,
         n38506, n38507, n38508, n38509, n38510, n38511, n38512, n38513,
         n38514, n38515, n38516, n38517, n38518, n38519, n38520, n38521,
         n38522, n38523, n38524, n38525, n38526, n38527, n38528, n38529,
         n38530, n38531, n38532, n38533, n38534, n38535, n38536, n38537,
         n38538, n38539, n38540, n38541, n38542, n38543, n38544, n38545,
         n38546, n38547, n38548, n38549, n38550, n38551, n38552, n38553,
         n38554, n38555, n38556, n38557, n38558, n38559, n38560, n38561,
         n38562, n38563, n38564, n38565, n38566, n38567, n38568, n38569,
         n38570, n38571, n38572, n38573, n38574, n38575, n38576, n38577,
         n38578, n38579, n38580, n38581, n38582, n38583, n38584, n38585,
         n38586, n38587, n38588, n38589, n38590, n38591, n38592, n38593,
         n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601,
         n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609,
         n38610, n38611, n38612, n38613, n38614, n38615, n38616, n38617,
         n38618, n38619, n38620, n38621, n38622, n38623, n38624, n38625,
         n38626, n38627, n38628, n38629, n38630, n38631, n38632, n38633,
         n38634, n38635, n38636, n38637, n38638, n38639, n38640, n38641,
         n38642, n38643, n38644, n38645, n38646, n38647, n38648, n38649,
         n38650, n38651, n38652, n38653, n38654, n38655, n38656, n38657,
         n38658, n38659, n38660, n38661, n38662, n38663, n38664, n38665,
         n38666, n38667, n38668, n38669, n38670, n38671, n38672, n38673,
         n38674, n38675, n38676, n38677, n38678, n38679, n38680, n38681,
         n38682, n38683, n38684, n38685, n38686, n38687, n38688, n38689,
         n38690, n38691, n38692, n38693, n38694, n38695, n38696, n38697,
         n38698, n38699, n38700, n38701, n38702, n38703, n38704, n38705,
         n38706, n38707, n38708, n38709, n38710, n38711, n38712, n38713,
         n38714, n38715, n38716, n38717, n38718, n38719, n38720, n38721,
         n38722, n38723, n38724, n38725, n38726, n38727, n38728, n38729,
         n38730, n38731, n38732, n38733, n38734, n38735, n38736, n38737,
         n38738, n38739, n38740, n38741, n38742, n38743, n38744, n38745,
         n38746, n38747, n38748, n38749, n38750, n38751, n38752, n38753,
         n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761,
         n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769,
         n38770, n38771, n38772, n38773, n38774, n38775, n38776, n38777,
         n38778, n38779, n38780, n38781, n38782, n38783, n38784, n38785,
         n38786, n38787, n38788, n38789, n38790, n38791, n38792, n38793,
         n38794, n38795, n38796, n38797, n38798, n38799, n38800, n38801,
         n38802, n38803, n38804, n38805, n38806, n38807, n38808, n38809,
         n38810, n38811, n38812, n38813, n38814, n38815, n38816, n38817,
         n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825,
         n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833,
         n38834, n38835, n38836, n38837, n38838, n38839, n38840, n38841,
         n38842, n38843, n38844, n38845, n38846, n38847, n38848, n38849,
         n38850, n38851, n38852, n38853, n38854, n38855, n38856, n38857,
         n38858, n38859, n38860, n38861, n38862, n38863, n38864, n38865,
         n38866, n38867, n38868, n38869, n38870, n38871, n38872, n38873,
         n38874, n38875, n38876, n38877, n38878, n38879, n38880, n38881,
         n38882, n38883, n38884, n38885, n38886, n38887, n38888, n38889,
         n38890, n38891, n38892, n38893, n38894, n38895, n38896, n38897,
         n38898, n38899, n38900, n38901, n38902, n38903, n38904, n38905,
         n38906, n38907, n38908, n38909, n38910, n38911, n38912, n38913,
         n38914, n38915, n38916, n38917, n38918, n38919, n38920, n38921,
         n38922, n38923, n38924, n38925, n38926, n38927, n38928, n38929,
         n38930, n38931, n38932, n38933, n38934, n38935, n38936, n38937,
         n38938, n38939, n38940, n38941, n38942, n38943, n38944, n38945,
         n38946, n38947, n38948, n38949, n38950, n38951, n38952, n38953,
         n38954, n38955, n38956, n38957, n38958, n38959, n38960, n38961,
         n38962, n38963, n38964, n38965, n38966, n38967, n38968, n38969,
         n38970, n38971, n38972, n38973, n38974, n38975, n38976, n38977,
         n38978, n38979, n38980, n38981, n38982, n38983, n38984, n38985,
         n38986, n38987, n38988, n38989, n38990, n38991, n38992, n38993,
         n38994, n38995, n38996, n38997, n38998, n38999, n39000, n39001,
         n39002, n39003, n39004, n39005, n39006, n39007, n39008, n39009,
         n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017,
         n39018, n39019, n39020, n39021, n39022, n39023, n39024, n39025,
         n39026, n39027, n39028, n39029, n39030, n39031, n39032, n39033,
         n39034, n39035, n39036, n39037, n39038, n39039, n39040, n39041,
         n39042, n39043, n39044, n39045, n39046, n39047, n39048, n39049,
         n39050, n39051, n39052, n39053, n39054, n39055, n39056, n39057,
         n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065,
         n39066, n39067, n39068, n39069, n39070, n39071, n39072, n39073,
         n39074, n39075, n39076, n39077, n39078, n39079, n39080, n39081,
         n39082, n39083, n39084, n39085, n39086, n39087, n39088, n39089,
         n39090, n39091, n39092, n39093, n39094, n39095, n39096, n39097,
         n39098, n39099, n39100, n39101, n39102, n39103, n39104, n39105,
         n39106, n39107, n39108, n39109, n39110, n39111, n39112, n39113,
         n39114, n39115, n39116, n39117, n39118, n39119, n39120, n39121,
         n39122, n39123, n39124, n39125, n39126, n39127, n39128, n39129,
         n39130, n39131, n39132, n39133, n39134, n39135, n39136, n39137,
         n39138, n39139, n39140, n39141, n39142, n39143, n39144, n39145,
         n39146, n39147, n39148, n39149, n39150, n39151, n39152, n39153,
         n39154, n39155, n39156, n39157, n39158, n39159, n39160, n39161,
         n39162, n39163, n39164, n39165, n39166, n39167, n39168, n39169,
         n39170, n39171, n39172, n39173, n39174, n39175, n39176, n39177,
         n39178, n39179, n39180, n39181, n39182, n39183, n39184, n39185,
         n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193,
         n39194, n39195, n39196, n39197, n39198, n39199, n39200, n39201,
         n39202, n39203, n39204, n39205, n39206, n39207, n39208, n39209,
         n39210, n39211, n39212, n39213, n39214, n39215, n39216, n39217,
         n39218, n39219, n39220, n39221, n39222, n39223, n39224, n39225,
         n39226, n39227, n39228, n39229, n39230, n39231, n39232, n39233,
         n39234, n39235, n39236, n39237, n39238, n39239, n39240, n39241,
         n39242, n39243, n39244, n39245, n39246, n39247, n39248, n39249,
         n39250, n39251, n39252, n39253, n39254, n39255, n39256, n39257,
         n39258, n39259, n39260, n39261, n39262, n39263, n39264, n39265,
         n39266, n39267, n39268, n39269, n39270, n39271, n39272, n39273,
         n39274, n39275, n39276, n39277, n39278, n39279, n39280, n39281,
         n39282, n39283, n39284, n39285, n39286, n39287, n39288, n39289,
         n39290, n39291, n39292, n39293, n39294, n39295, n39296, n39297,
         n39298, n39299, n39300, n39301, n39302, n39303, n39304, n39305,
         n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
         n39314, n39315, n39316, n39317, n39318, n39319, n39320, n39321,
         n39322, n39323, n39324, n39325, n39326, n39327, n39328, n39329,
         n39330, n39331, n39332, n39333, n39334;

  XOR U3841 ( .A(DB[3834]), .B(n1), .Z(min_val_out[9]) );
  AND U3842 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3843 ( .A(n4), .B(n5), .Z(n3) );
  XOR U3844 ( .A(DB[3834]), .B(DB[3819]), .Z(n5) );
  AND U3845 ( .A(n6), .B(n7), .Z(n4) );
  XOR U3846 ( .A(n8), .B(n9), .Z(n7) );
  XOR U3847 ( .A(DB[3819]), .B(DB[3804]), .Z(n9) );
  AND U3848 ( .A(n10), .B(n11), .Z(n8) );
  XOR U3849 ( .A(n12), .B(n13), .Z(n11) );
  XOR U3850 ( .A(DB[3804]), .B(DB[3789]), .Z(n13) );
  AND U3851 ( .A(n14), .B(n15), .Z(n12) );
  XOR U3852 ( .A(n16), .B(n17), .Z(n15) );
  XOR U3853 ( .A(DB[3789]), .B(DB[3774]), .Z(n17) );
  AND U3854 ( .A(n18), .B(n19), .Z(n16) );
  XOR U3855 ( .A(n20), .B(n21), .Z(n19) );
  XOR U3856 ( .A(DB[3774]), .B(DB[3759]), .Z(n21) );
  AND U3857 ( .A(n22), .B(n23), .Z(n20) );
  XOR U3858 ( .A(n24), .B(n25), .Z(n23) );
  XOR U3859 ( .A(DB[3759]), .B(DB[3744]), .Z(n25) );
  AND U3860 ( .A(n26), .B(n27), .Z(n24) );
  XOR U3861 ( .A(n28), .B(n29), .Z(n27) );
  XOR U3862 ( .A(DB[3744]), .B(DB[3729]), .Z(n29) );
  AND U3863 ( .A(n30), .B(n31), .Z(n28) );
  XOR U3864 ( .A(n32), .B(n33), .Z(n31) );
  XOR U3865 ( .A(DB[3729]), .B(DB[3714]), .Z(n33) );
  AND U3866 ( .A(n34), .B(n35), .Z(n32) );
  XOR U3867 ( .A(n36), .B(n37), .Z(n35) );
  XOR U3868 ( .A(DB[3714]), .B(DB[3699]), .Z(n37) );
  AND U3869 ( .A(n38), .B(n39), .Z(n36) );
  XOR U3870 ( .A(n40), .B(n41), .Z(n39) );
  XOR U3871 ( .A(DB[3699]), .B(DB[3684]), .Z(n41) );
  AND U3872 ( .A(n42), .B(n43), .Z(n40) );
  XOR U3873 ( .A(n44), .B(n45), .Z(n43) );
  XOR U3874 ( .A(DB[3684]), .B(DB[3669]), .Z(n45) );
  AND U3875 ( .A(n46), .B(n47), .Z(n44) );
  XOR U3876 ( .A(n48), .B(n49), .Z(n47) );
  XOR U3877 ( .A(DB[3669]), .B(DB[3654]), .Z(n49) );
  AND U3878 ( .A(n50), .B(n51), .Z(n48) );
  XOR U3879 ( .A(n52), .B(n53), .Z(n51) );
  XOR U3880 ( .A(DB[3654]), .B(DB[3639]), .Z(n53) );
  AND U3881 ( .A(n54), .B(n55), .Z(n52) );
  XOR U3882 ( .A(n56), .B(n57), .Z(n55) );
  XOR U3883 ( .A(DB[3639]), .B(DB[3624]), .Z(n57) );
  AND U3884 ( .A(n58), .B(n59), .Z(n56) );
  XOR U3885 ( .A(n60), .B(n61), .Z(n59) );
  XOR U3886 ( .A(DB[3624]), .B(DB[3609]), .Z(n61) );
  AND U3887 ( .A(n62), .B(n63), .Z(n60) );
  XOR U3888 ( .A(n64), .B(n65), .Z(n63) );
  XOR U3889 ( .A(DB[3609]), .B(DB[3594]), .Z(n65) );
  AND U3890 ( .A(n66), .B(n67), .Z(n64) );
  XOR U3891 ( .A(n68), .B(n69), .Z(n67) );
  XOR U3892 ( .A(DB[3594]), .B(DB[3579]), .Z(n69) );
  AND U3893 ( .A(n70), .B(n71), .Z(n68) );
  XOR U3894 ( .A(n72), .B(n73), .Z(n71) );
  XOR U3895 ( .A(DB[3579]), .B(DB[3564]), .Z(n73) );
  AND U3896 ( .A(n74), .B(n75), .Z(n72) );
  XOR U3897 ( .A(n76), .B(n77), .Z(n75) );
  XOR U3898 ( .A(DB[3564]), .B(DB[3549]), .Z(n77) );
  AND U3899 ( .A(n78), .B(n79), .Z(n76) );
  XOR U3900 ( .A(n80), .B(n81), .Z(n79) );
  XOR U3901 ( .A(DB[3549]), .B(DB[3534]), .Z(n81) );
  AND U3902 ( .A(n82), .B(n83), .Z(n80) );
  XOR U3903 ( .A(n84), .B(n85), .Z(n83) );
  XOR U3904 ( .A(DB[3534]), .B(DB[3519]), .Z(n85) );
  AND U3905 ( .A(n86), .B(n87), .Z(n84) );
  XOR U3906 ( .A(n88), .B(n89), .Z(n87) );
  XOR U3907 ( .A(DB[3519]), .B(DB[3504]), .Z(n89) );
  AND U3908 ( .A(n90), .B(n91), .Z(n88) );
  XOR U3909 ( .A(n92), .B(n93), .Z(n91) );
  XOR U3910 ( .A(DB[3504]), .B(DB[3489]), .Z(n93) );
  AND U3911 ( .A(n94), .B(n95), .Z(n92) );
  XOR U3912 ( .A(n96), .B(n97), .Z(n95) );
  XOR U3913 ( .A(DB[3489]), .B(DB[3474]), .Z(n97) );
  AND U3914 ( .A(n98), .B(n99), .Z(n96) );
  XOR U3915 ( .A(n100), .B(n101), .Z(n99) );
  XOR U3916 ( .A(DB[3474]), .B(DB[3459]), .Z(n101) );
  AND U3917 ( .A(n102), .B(n103), .Z(n100) );
  XOR U3918 ( .A(n104), .B(n105), .Z(n103) );
  XOR U3919 ( .A(DB[3459]), .B(DB[3444]), .Z(n105) );
  AND U3920 ( .A(n106), .B(n107), .Z(n104) );
  XOR U3921 ( .A(n108), .B(n109), .Z(n107) );
  XOR U3922 ( .A(DB[3444]), .B(DB[3429]), .Z(n109) );
  AND U3923 ( .A(n110), .B(n111), .Z(n108) );
  XOR U3924 ( .A(n112), .B(n113), .Z(n111) );
  XOR U3925 ( .A(DB[3429]), .B(DB[3414]), .Z(n113) );
  AND U3926 ( .A(n114), .B(n115), .Z(n112) );
  XOR U3927 ( .A(n116), .B(n117), .Z(n115) );
  XOR U3928 ( .A(DB[3414]), .B(DB[3399]), .Z(n117) );
  AND U3929 ( .A(n118), .B(n119), .Z(n116) );
  XOR U3930 ( .A(n120), .B(n121), .Z(n119) );
  XOR U3931 ( .A(DB[3399]), .B(DB[3384]), .Z(n121) );
  AND U3932 ( .A(n122), .B(n123), .Z(n120) );
  XOR U3933 ( .A(n124), .B(n125), .Z(n123) );
  XOR U3934 ( .A(DB[3384]), .B(DB[3369]), .Z(n125) );
  AND U3935 ( .A(n126), .B(n127), .Z(n124) );
  XOR U3936 ( .A(n128), .B(n129), .Z(n127) );
  XOR U3937 ( .A(DB[3369]), .B(DB[3354]), .Z(n129) );
  AND U3938 ( .A(n130), .B(n131), .Z(n128) );
  XOR U3939 ( .A(n132), .B(n133), .Z(n131) );
  XOR U3940 ( .A(DB[3354]), .B(DB[3339]), .Z(n133) );
  AND U3941 ( .A(n134), .B(n135), .Z(n132) );
  XOR U3942 ( .A(n136), .B(n137), .Z(n135) );
  XOR U3943 ( .A(DB[3339]), .B(DB[3324]), .Z(n137) );
  AND U3944 ( .A(n138), .B(n139), .Z(n136) );
  XOR U3945 ( .A(n140), .B(n141), .Z(n139) );
  XOR U3946 ( .A(DB[3324]), .B(DB[3309]), .Z(n141) );
  AND U3947 ( .A(n142), .B(n143), .Z(n140) );
  XOR U3948 ( .A(n144), .B(n145), .Z(n143) );
  XOR U3949 ( .A(DB[3309]), .B(DB[3294]), .Z(n145) );
  AND U3950 ( .A(n146), .B(n147), .Z(n144) );
  XOR U3951 ( .A(n148), .B(n149), .Z(n147) );
  XOR U3952 ( .A(DB[3294]), .B(DB[3279]), .Z(n149) );
  AND U3953 ( .A(n150), .B(n151), .Z(n148) );
  XOR U3954 ( .A(n152), .B(n153), .Z(n151) );
  XOR U3955 ( .A(DB[3279]), .B(DB[3264]), .Z(n153) );
  AND U3956 ( .A(n154), .B(n155), .Z(n152) );
  XOR U3957 ( .A(n156), .B(n157), .Z(n155) );
  XOR U3958 ( .A(DB[3264]), .B(DB[3249]), .Z(n157) );
  AND U3959 ( .A(n158), .B(n159), .Z(n156) );
  XOR U3960 ( .A(n160), .B(n161), .Z(n159) );
  XOR U3961 ( .A(DB[3249]), .B(DB[3234]), .Z(n161) );
  AND U3962 ( .A(n162), .B(n163), .Z(n160) );
  XOR U3963 ( .A(n164), .B(n165), .Z(n163) );
  XOR U3964 ( .A(DB[3234]), .B(DB[3219]), .Z(n165) );
  AND U3965 ( .A(n166), .B(n167), .Z(n164) );
  XOR U3966 ( .A(n168), .B(n169), .Z(n167) );
  XOR U3967 ( .A(DB[3219]), .B(DB[3204]), .Z(n169) );
  AND U3968 ( .A(n170), .B(n171), .Z(n168) );
  XOR U3969 ( .A(n172), .B(n173), .Z(n171) );
  XOR U3970 ( .A(DB[3204]), .B(DB[3189]), .Z(n173) );
  AND U3971 ( .A(n174), .B(n175), .Z(n172) );
  XOR U3972 ( .A(n176), .B(n177), .Z(n175) );
  XOR U3973 ( .A(DB[3189]), .B(DB[3174]), .Z(n177) );
  AND U3974 ( .A(n178), .B(n179), .Z(n176) );
  XOR U3975 ( .A(n180), .B(n181), .Z(n179) );
  XOR U3976 ( .A(DB[3174]), .B(DB[3159]), .Z(n181) );
  AND U3977 ( .A(n182), .B(n183), .Z(n180) );
  XOR U3978 ( .A(n184), .B(n185), .Z(n183) );
  XOR U3979 ( .A(DB[3159]), .B(DB[3144]), .Z(n185) );
  AND U3980 ( .A(n186), .B(n187), .Z(n184) );
  XOR U3981 ( .A(n188), .B(n189), .Z(n187) );
  XOR U3982 ( .A(DB[3144]), .B(DB[3129]), .Z(n189) );
  AND U3983 ( .A(n190), .B(n191), .Z(n188) );
  XOR U3984 ( .A(n192), .B(n193), .Z(n191) );
  XOR U3985 ( .A(DB[3129]), .B(DB[3114]), .Z(n193) );
  AND U3986 ( .A(n194), .B(n195), .Z(n192) );
  XOR U3987 ( .A(n196), .B(n197), .Z(n195) );
  XOR U3988 ( .A(DB[3114]), .B(DB[3099]), .Z(n197) );
  AND U3989 ( .A(n198), .B(n199), .Z(n196) );
  XOR U3990 ( .A(n200), .B(n201), .Z(n199) );
  XOR U3991 ( .A(DB[3099]), .B(DB[3084]), .Z(n201) );
  AND U3992 ( .A(n202), .B(n203), .Z(n200) );
  XOR U3993 ( .A(n204), .B(n205), .Z(n203) );
  XOR U3994 ( .A(DB[3084]), .B(DB[3069]), .Z(n205) );
  AND U3995 ( .A(n206), .B(n207), .Z(n204) );
  XOR U3996 ( .A(n208), .B(n209), .Z(n207) );
  XOR U3997 ( .A(DB[3069]), .B(DB[3054]), .Z(n209) );
  AND U3998 ( .A(n210), .B(n211), .Z(n208) );
  XOR U3999 ( .A(n212), .B(n213), .Z(n211) );
  XOR U4000 ( .A(DB[3054]), .B(DB[3039]), .Z(n213) );
  AND U4001 ( .A(n214), .B(n215), .Z(n212) );
  XOR U4002 ( .A(n216), .B(n217), .Z(n215) );
  XOR U4003 ( .A(DB[3039]), .B(DB[3024]), .Z(n217) );
  AND U4004 ( .A(n218), .B(n219), .Z(n216) );
  XOR U4005 ( .A(n220), .B(n221), .Z(n219) );
  XOR U4006 ( .A(DB[3024]), .B(DB[3009]), .Z(n221) );
  AND U4007 ( .A(n222), .B(n223), .Z(n220) );
  XOR U4008 ( .A(n224), .B(n225), .Z(n223) );
  XOR U4009 ( .A(DB[3009]), .B(DB[2994]), .Z(n225) );
  AND U4010 ( .A(n226), .B(n227), .Z(n224) );
  XOR U4011 ( .A(n228), .B(n229), .Z(n227) );
  XOR U4012 ( .A(DB[2994]), .B(DB[2979]), .Z(n229) );
  AND U4013 ( .A(n230), .B(n231), .Z(n228) );
  XOR U4014 ( .A(n232), .B(n233), .Z(n231) );
  XOR U4015 ( .A(DB[2979]), .B(DB[2964]), .Z(n233) );
  AND U4016 ( .A(n234), .B(n235), .Z(n232) );
  XOR U4017 ( .A(n236), .B(n237), .Z(n235) );
  XOR U4018 ( .A(DB[2964]), .B(DB[2949]), .Z(n237) );
  AND U4019 ( .A(n238), .B(n239), .Z(n236) );
  XOR U4020 ( .A(n240), .B(n241), .Z(n239) );
  XOR U4021 ( .A(DB[2949]), .B(DB[2934]), .Z(n241) );
  AND U4022 ( .A(n242), .B(n243), .Z(n240) );
  XOR U4023 ( .A(n244), .B(n245), .Z(n243) );
  XOR U4024 ( .A(DB[2934]), .B(DB[2919]), .Z(n245) );
  AND U4025 ( .A(n246), .B(n247), .Z(n244) );
  XOR U4026 ( .A(n248), .B(n249), .Z(n247) );
  XOR U4027 ( .A(DB[2919]), .B(DB[2904]), .Z(n249) );
  AND U4028 ( .A(n250), .B(n251), .Z(n248) );
  XOR U4029 ( .A(n252), .B(n253), .Z(n251) );
  XOR U4030 ( .A(DB[2904]), .B(DB[2889]), .Z(n253) );
  AND U4031 ( .A(n254), .B(n255), .Z(n252) );
  XOR U4032 ( .A(n256), .B(n257), .Z(n255) );
  XOR U4033 ( .A(DB[2889]), .B(DB[2874]), .Z(n257) );
  AND U4034 ( .A(n258), .B(n259), .Z(n256) );
  XOR U4035 ( .A(n260), .B(n261), .Z(n259) );
  XOR U4036 ( .A(DB[2874]), .B(DB[2859]), .Z(n261) );
  AND U4037 ( .A(n262), .B(n263), .Z(n260) );
  XOR U4038 ( .A(n264), .B(n265), .Z(n263) );
  XOR U4039 ( .A(DB[2859]), .B(DB[2844]), .Z(n265) );
  AND U4040 ( .A(n266), .B(n267), .Z(n264) );
  XOR U4041 ( .A(n268), .B(n269), .Z(n267) );
  XOR U4042 ( .A(DB[2844]), .B(DB[2829]), .Z(n269) );
  AND U4043 ( .A(n270), .B(n271), .Z(n268) );
  XOR U4044 ( .A(n272), .B(n273), .Z(n271) );
  XOR U4045 ( .A(DB[2829]), .B(DB[2814]), .Z(n273) );
  AND U4046 ( .A(n274), .B(n275), .Z(n272) );
  XOR U4047 ( .A(n276), .B(n277), .Z(n275) );
  XOR U4048 ( .A(DB[2814]), .B(DB[2799]), .Z(n277) );
  AND U4049 ( .A(n278), .B(n279), .Z(n276) );
  XOR U4050 ( .A(n280), .B(n281), .Z(n279) );
  XOR U4051 ( .A(DB[2799]), .B(DB[2784]), .Z(n281) );
  AND U4052 ( .A(n282), .B(n283), .Z(n280) );
  XOR U4053 ( .A(n284), .B(n285), .Z(n283) );
  XOR U4054 ( .A(DB[2784]), .B(DB[2769]), .Z(n285) );
  AND U4055 ( .A(n286), .B(n287), .Z(n284) );
  XOR U4056 ( .A(n288), .B(n289), .Z(n287) );
  XOR U4057 ( .A(DB[2769]), .B(DB[2754]), .Z(n289) );
  AND U4058 ( .A(n290), .B(n291), .Z(n288) );
  XOR U4059 ( .A(n292), .B(n293), .Z(n291) );
  XOR U4060 ( .A(DB[2754]), .B(DB[2739]), .Z(n293) );
  AND U4061 ( .A(n294), .B(n295), .Z(n292) );
  XOR U4062 ( .A(n296), .B(n297), .Z(n295) );
  XOR U4063 ( .A(DB[2739]), .B(DB[2724]), .Z(n297) );
  AND U4064 ( .A(n298), .B(n299), .Z(n296) );
  XOR U4065 ( .A(n300), .B(n301), .Z(n299) );
  XOR U4066 ( .A(DB[2724]), .B(DB[2709]), .Z(n301) );
  AND U4067 ( .A(n302), .B(n303), .Z(n300) );
  XOR U4068 ( .A(n304), .B(n305), .Z(n303) );
  XOR U4069 ( .A(DB[2709]), .B(DB[2694]), .Z(n305) );
  AND U4070 ( .A(n306), .B(n307), .Z(n304) );
  XOR U4071 ( .A(n308), .B(n309), .Z(n307) );
  XOR U4072 ( .A(DB[2694]), .B(DB[2679]), .Z(n309) );
  AND U4073 ( .A(n310), .B(n311), .Z(n308) );
  XOR U4074 ( .A(n312), .B(n313), .Z(n311) );
  XOR U4075 ( .A(DB[2679]), .B(DB[2664]), .Z(n313) );
  AND U4076 ( .A(n314), .B(n315), .Z(n312) );
  XOR U4077 ( .A(n316), .B(n317), .Z(n315) );
  XOR U4078 ( .A(DB[2664]), .B(DB[2649]), .Z(n317) );
  AND U4079 ( .A(n318), .B(n319), .Z(n316) );
  XOR U4080 ( .A(n320), .B(n321), .Z(n319) );
  XOR U4081 ( .A(DB[2649]), .B(DB[2634]), .Z(n321) );
  AND U4082 ( .A(n322), .B(n323), .Z(n320) );
  XOR U4083 ( .A(n324), .B(n325), .Z(n323) );
  XOR U4084 ( .A(DB[2634]), .B(DB[2619]), .Z(n325) );
  AND U4085 ( .A(n326), .B(n327), .Z(n324) );
  XOR U4086 ( .A(n328), .B(n329), .Z(n327) );
  XOR U4087 ( .A(DB[2619]), .B(DB[2604]), .Z(n329) );
  AND U4088 ( .A(n330), .B(n331), .Z(n328) );
  XOR U4089 ( .A(n332), .B(n333), .Z(n331) );
  XOR U4090 ( .A(DB[2604]), .B(DB[2589]), .Z(n333) );
  AND U4091 ( .A(n334), .B(n335), .Z(n332) );
  XOR U4092 ( .A(n336), .B(n337), .Z(n335) );
  XOR U4093 ( .A(DB[2589]), .B(DB[2574]), .Z(n337) );
  AND U4094 ( .A(n338), .B(n339), .Z(n336) );
  XOR U4095 ( .A(n340), .B(n341), .Z(n339) );
  XOR U4096 ( .A(DB[2574]), .B(DB[2559]), .Z(n341) );
  AND U4097 ( .A(n342), .B(n343), .Z(n340) );
  XOR U4098 ( .A(n344), .B(n345), .Z(n343) );
  XOR U4099 ( .A(DB[2559]), .B(DB[2544]), .Z(n345) );
  AND U4100 ( .A(n346), .B(n347), .Z(n344) );
  XOR U4101 ( .A(n348), .B(n349), .Z(n347) );
  XOR U4102 ( .A(DB[2544]), .B(DB[2529]), .Z(n349) );
  AND U4103 ( .A(n350), .B(n351), .Z(n348) );
  XOR U4104 ( .A(n352), .B(n353), .Z(n351) );
  XOR U4105 ( .A(DB[2529]), .B(DB[2514]), .Z(n353) );
  AND U4106 ( .A(n354), .B(n355), .Z(n352) );
  XOR U4107 ( .A(n356), .B(n357), .Z(n355) );
  XOR U4108 ( .A(DB[2514]), .B(DB[2499]), .Z(n357) );
  AND U4109 ( .A(n358), .B(n359), .Z(n356) );
  XOR U4110 ( .A(n360), .B(n361), .Z(n359) );
  XOR U4111 ( .A(DB[2499]), .B(DB[2484]), .Z(n361) );
  AND U4112 ( .A(n362), .B(n363), .Z(n360) );
  XOR U4113 ( .A(n364), .B(n365), .Z(n363) );
  XOR U4114 ( .A(DB[2484]), .B(DB[2469]), .Z(n365) );
  AND U4115 ( .A(n366), .B(n367), .Z(n364) );
  XOR U4116 ( .A(n368), .B(n369), .Z(n367) );
  XOR U4117 ( .A(DB[2469]), .B(DB[2454]), .Z(n369) );
  AND U4118 ( .A(n370), .B(n371), .Z(n368) );
  XOR U4119 ( .A(n372), .B(n373), .Z(n371) );
  XOR U4120 ( .A(DB[2454]), .B(DB[2439]), .Z(n373) );
  AND U4121 ( .A(n374), .B(n375), .Z(n372) );
  XOR U4122 ( .A(n376), .B(n377), .Z(n375) );
  XOR U4123 ( .A(DB[2439]), .B(DB[2424]), .Z(n377) );
  AND U4124 ( .A(n378), .B(n379), .Z(n376) );
  XOR U4125 ( .A(n380), .B(n381), .Z(n379) );
  XOR U4126 ( .A(DB[2424]), .B(DB[2409]), .Z(n381) );
  AND U4127 ( .A(n382), .B(n383), .Z(n380) );
  XOR U4128 ( .A(n384), .B(n385), .Z(n383) );
  XOR U4129 ( .A(DB[2409]), .B(DB[2394]), .Z(n385) );
  AND U4130 ( .A(n386), .B(n387), .Z(n384) );
  XOR U4131 ( .A(n388), .B(n389), .Z(n387) );
  XOR U4132 ( .A(DB[2394]), .B(DB[2379]), .Z(n389) );
  AND U4133 ( .A(n390), .B(n391), .Z(n388) );
  XOR U4134 ( .A(n392), .B(n393), .Z(n391) );
  XOR U4135 ( .A(DB[2379]), .B(DB[2364]), .Z(n393) );
  AND U4136 ( .A(n394), .B(n395), .Z(n392) );
  XOR U4137 ( .A(n396), .B(n397), .Z(n395) );
  XOR U4138 ( .A(DB[2364]), .B(DB[2349]), .Z(n397) );
  AND U4139 ( .A(n398), .B(n399), .Z(n396) );
  XOR U4140 ( .A(n400), .B(n401), .Z(n399) );
  XOR U4141 ( .A(DB[2349]), .B(DB[2334]), .Z(n401) );
  AND U4142 ( .A(n402), .B(n403), .Z(n400) );
  XOR U4143 ( .A(n404), .B(n405), .Z(n403) );
  XOR U4144 ( .A(DB[2334]), .B(DB[2319]), .Z(n405) );
  AND U4145 ( .A(n406), .B(n407), .Z(n404) );
  XOR U4146 ( .A(n408), .B(n409), .Z(n407) );
  XOR U4147 ( .A(DB[2319]), .B(DB[2304]), .Z(n409) );
  AND U4148 ( .A(n410), .B(n411), .Z(n408) );
  XOR U4149 ( .A(n412), .B(n413), .Z(n411) );
  XOR U4150 ( .A(DB[2304]), .B(DB[2289]), .Z(n413) );
  AND U4151 ( .A(n414), .B(n415), .Z(n412) );
  XOR U4152 ( .A(n416), .B(n417), .Z(n415) );
  XOR U4153 ( .A(DB[2289]), .B(DB[2274]), .Z(n417) );
  AND U4154 ( .A(n418), .B(n419), .Z(n416) );
  XOR U4155 ( .A(n420), .B(n421), .Z(n419) );
  XOR U4156 ( .A(DB[2274]), .B(DB[2259]), .Z(n421) );
  AND U4157 ( .A(n422), .B(n423), .Z(n420) );
  XOR U4158 ( .A(n424), .B(n425), .Z(n423) );
  XOR U4159 ( .A(DB[2259]), .B(DB[2244]), .Z(n425) );
  AND U4160 ( .A(n426), .B(n427), .Z(n424) );
  XOR U4161 ( .A(n428), .B(n429), .Z(n427) );
  XOR U4162 ( .A(DB[2244]), .B(DB[2229]), .Z(n429) );
  AND U4163 ( .A(n430), .B(n431), .Z(n428) );
  XOR U4164 ( .A(n432), .B(n433), .Z(n431) );
  XOR U4165 ( .A(DB[2229]), .B(DB[2214]), .Z(n433) );
  AND U4166 ( .A(n434), .B(n435), .Z(n432) );
  XOR U4167 ( .A(n436), .B(n437), .Z(n435) );
  XOR U4168 ( .A(DB[2214]), .B(DB[2199]), .Z(n437) );
  AND U4169 ( .A(n438), .B(n439), .Z(n436) );
  XOR U4170 ( .A(n440), .B(n441), .Z(n439) );
  XOR U4171 ( .A(DB[2199]), .B(DB[2184]), .Z(n441) );
  AND U4172 ( .A(n442), .B(n443), .Z(n440) );
  XOR U4173 ( .A(n444), .B(n445), .Z(n443) );
  XOR U4174 ( .A(DB[2184]), .B(DB[2169]), .Z(n445) );
  AND U4175 ( .A(n446), .B(n447), .Z(n444) );
  XOR U4176 ( .A(n448), .B(n449), .Z(n447) );
  XOR U4177 ( .A(DB[2169]), .B(DB[2154]), .Z(n449) );
  AND U4178 ( .A(n450), .B(n451), .Z(n448) );
  XOR U4179 ( .A(n452), .B(n453), .Z(n451) );
  XOR U4180 ( .A(DB[2154]), .B(DB[2139]), .Z(n453) );
  AND U4181 ( .A(n454), .B(n455), .Z(n452) );
  XOR U4182 ( .A(n456), .B(n457), .Z(n455) );
  XOR U4183 ( .A(DB[2139]), .B(DB[2124]), .Z(n457) );
  AND U4184 ( .A(n458), .B(n459), .Z(n456) );
  XOR U4185 ( .A(n460), .B(n461), .Z(n459) );
  XOR U4186 ( .A(DB[2124]), .B(DB[2109]), .Z(n461) );
  AND U4187 ( .A(n462), .B(n463), .Z(n460) );
  XOR U4188 ( .A(n464), .B(n465), .Z(n463) );
  XOR U4189 ( .A(DB[2109]), .B(DB[2094]), .Z(n465) );
  AND U4190 ( .A(n466), .B(n467), .Z(n464) );
  XOR U4191 ( .A(n468), .B(n469), .Z(n467) );
  XOR U4192 ( .A(DB[2094]), .B(DB[2079]), .Z(n469) );
  AND U4193 ( .A(n470), .B(n471), .Z(n468) );
  XOR U4194 ( .A(n472), .B(n473), .Z(n471) );
  XOR U4195 ( .A(DB[2079]), .B(DB[2064]), .Z(n473) );
  AND U4196 ( .A(n474), .B(n475), .Z(n472) );
  XOR U4197 ( .A(n476), .B(n477), .Z(n475) );
  XOR U4198 ( .A(DB[2064]), .B(DB[2049]), .Z(n477) );
  AND U4199 ( .A(n478), .B(n479), .Z(n476) );
  XOR U4200 ( .A(n480), .B(n481), .Z(n479) );
  XOR U4201 ( .A(DB[2049]), .B(DB[2034]), .Z(n481) );
  AND U4202 ( .A(n482), .B(n483), .Z(n480) );
  XOR U4203 ( .A(n484), .B(n485), .Z(n483) );
  XOR U4204 ( .A(DB[2034]), .B(DB[2019]), .Z(n485) );
  AND U4205 ( .A(n486), .B(n487), .Z(n484) );
  XOR U4206 ( .A(n488), .B(n489), .Z(n487) );
  XOR U4207 ( .A(DB[2019]), .B(DB[2004]), .Z(n489) );
  AND U4208 ( .A(n490), .B(n491), .Z(n488) );
  XOR U4209 ( .A(n492), .B(n493), .Z(n491) );
  XOR U4210 ( .A(DB[2004]), .B(DB[1989]), .Z(n493) );
  AND U4211 ( .A(n494), .B(n495), .Z(n492) );
  XOR U4212 ( .A(n496), .B(n497), .Z(n495) );
  XOR U4213 ( .A(DB[1989]), .B(DB[1974]), .Z(n497) );
  AND U4214 ( .A(n498), .B(n499), .Z(n496) );
  XOR U4215 ( .A(n500), .B(n501), .Z(n499) );
  XOR U4216 ( .A(DB[1974]), .B(DB[1959]), .Z(n501) );
  AND U4217 ( .A(n502), .B(n503), .Z(n500) );
  XOR U4218 ( .A(n504), .B(n505), .Z(n503) );
  XOR U4219 ( .A(DB[1959]), .B(DB[1944]), .Z(n505) );
  AND U4220 ( .A(n506), .B(n507), .Z(n504) );
  XOR U4221 ( .A(n508), .B(n509), .Z(n507) );
  XOR U4222 ( .A(DB[1944]), .B(DB[1929]), .Z(n509) );
  AND U4223 ( .A(n510), .B(n511), .Z(n508) );
  XOR U4224 ( .A(n512), .B(n513), .Z(n511) );
  XOR U4225 ( .A(DB[1929]), .B(DB[1914]), .Z(n513) );
  AND U4226 ( .A(n514), .B(n515), .Z(n512) );
  XOR U4227 ( .A(n516), .B(n517), .Z(n515) );
  XOR U4228 ( .A(DB[1914]), .B(DB[1899]), .Z(n517) );
  AND U4229 ( .A(n518), .B(n519), .Z(n516) );
  XOR U4230 ( .A(n520), .B(n521), .Z(n519) );
  XOR U4231 ( .A(DB[1899]), .B(DB[1884]), .Z(n521) );
  AND U4232 ( .A(n522), .B(n523), .Z(n520) );
  XOR U4233 ( .A(n524), .B(n525), .Z(n523) );
  XOR U4234 ( .A(DB[1884]), .B(DB[1869]), .Z(n525) );
  AND U4235 ( .A(n526), .B(n527), .Z(n524) );
  XOR U4236 ( .A(n528), .B(n529), .Z(n527) );
  XOR U4237 ( .A(DB[1869]), .B(DB[1854]), .Z(n529) );
  AND U4238 ( .A(n530), .B(n531), .Z(n528) );
  XOR U4239 ( .A(n532), .B(n533), .Z(n531) );
  XOR U4240 ( .A(DB[1854]), .B(DB[1839]), .Z(n533) );
  AND U4241 ( .A(n534), .B(n535), .Z(n532) );
  XOR U4242 ( .A(n536), .B(n537), .Z(n535) );
  XOR U4243 ( .A(DB[1839]), .B(DB[1824]), .Z(n537) );
  AND U4244 ( .A(n538), .B(n539), .Z(n536) );
  XOR U4245 ( .A(n540), .B(n541), .Z(n539) );
  XOR U4246 ( .A(DB[1824]), .B(DB[1809]), .Z(n541) );
  AND U4247 ( .A(n542), .B(n543), .Z(n540) );
  XOR U4248 ( .A(n544), .B(n545), .Z(n543) );
  XOR U4249 ( .A(DB[1809]), .B(DB[1794]), .Z(n545) );
  AND U4250 ( .A(n546), .B(n547), .Z(n544) );
  XOR U4251 ( .A(n548), .B(n549), .Z(n547) );
  XOR U4252 ( .A(DB[1794]), .B(DB[1779]), .Z(n549) );
  AND U4253 ( .A(n550), .B(n551), .Z(n548) );
  XOR U4254 ( .A(n552), .B(n553), .Z(n551) );
  XOR U4255 ( .A(DB[1779]), .B(DB[1764]), .Z(n553) );
  AND U4256 ( .A(n554), .B(n555), .Z(n552) );
  XOR U4257 ( .A(n556), .B(n557), .Z(n555) );
  XOR U4258 ( .A(DB[1764]), .B(DB[1749]), .Z(n557) );
  AND U4259 ( .A(n558), .B(n559), .Z(n556) );
  XOR U4260 ( .A(n560), .B(n561), .Z(n559) );
  XOR U4261 ( .A(DB[1749]), .B(DB[1734]), .Z(n561) );
  AND U4262 ( .A(n562), .B(n563), .Z(n560) );
  XOR U4263 ( .A(n564), .B(n565), .Z(n563) );
  XOR U4264 ( .A(DB[1734]), .B(DB[1719]), .Z(n565) );
  AND U4265 ( .A(n566), .B(n567), .Z(n564) );
  XOR U4266 ( .A(n568), .B(n569), .Z(n567) );
  XOR U4267 ( .A(DB[1719]), .B(DB[1704]), .Z(n569) );
  AND U4268 ( .A(n570), .B(n571), .Z(n568) );
  XOR U4269 ( .A(n572), .B(n573), .Z(n571) );
  XOR U4270 ( .A(DB[1704]), .B(DB[1689]), .Z(n573) );
  AND U4271 ( .A(n574), .B(n575), .Z(n572) );
  XOR U4272 ( .A(n576), .B(n577), .Z(n575) );
  XOR U4273 ( .A(DB[1689]), .B(DB[1674]), .Z(n577) );
  AND U4274 ( .A(n578), .B(n579), .Z(n576) );
  XOR U4275 ( .A(n580), .B(n581), .Z(n579) );
  XOR U4276 ( .A(DB[1674]), .B(DB[1659]), .Z(n581) );
  AND U4277 ( .A(n582), .B(n583), .Z(n580) );
  XOR U4278 ( .A(n584), .B(n585), .Z(n583) );
  XOR U4279 ( .A(DB[1659]), .B(DB[1644]), .Z(n585) );
  AND U4280 ( .A(n586), .B(n587), .Z(n584) );
  XOR U4281 ( .A(n588), .B(n589), .Z(n587) );
  XOR U4282 ( .A(DB[1644]), .B(DB[1629]), .Z(n589) );
  AND U4283 ( .A(n590), .B(n591), .Z(n588) );
  XOR U4284 ( .A(n592), .B(n593), .Z(n591) );
  XOR U4285 ( .A(DB[1629]), .B(DB[1614]), .Z(n593) );
  AND U4286 ( .A(n594), .B(n595), .Z(n592) );
  XOR U4287 ( .A(n596), .B(n597), .Z(n595) );
  XOR U4288 ( .A(DB[1614]), .B(DB[1599]), .Z(n597) );
  AND U4289 ( .A(n598), .B(n599), .Z(n596) );
  XOR U4290 ( .A(n600), .B(n601), .Z(n599) );
  XOR U4291 ( .A(DB[1599]), .B(DB[1584]), .Z(n601) );
  AND U4292 ( .A(n602), .B(n603), .Z(n600) );
  XOR U4293 ( .A(n604), .B(n605), .Z(n603) );
  XOR U4294 ( .A(DB[1584]), .B(DB[1569]), .Z(n605) );
  AND U4295 ( .A(n606), .B(n607), .Z(n604) );
  XOR U4296 ( .A(n608), .B(n609), .Z(n607) );
  XOR U4297 ( .A(DB[1569]), .B(DB[1554]), .Z(n609) );
  AND U4298 ( .A(n610), .B(n611), .Z(n608) );
  XOR U4299 ( .A(n612), .B(n613), .Z(n611) );
  XOR U4300 ( .A(DB[1554]), .B(DB[1539]), .Z(n613) );
  AND U4301 ( .A(n614), .B(n615), .Z(n612) );
  XOR U4302 ( .A(n616), .B(n617), .Z(n615) );
  XOR U4303 ( .A(DB[1539]), .B(DB[1524]), .Z(n617) );
  AND U4304 ( .A(n618), .B(n619), .Z(n616) );
  XOR U4305 ( .A(n620), .B(n621), .Z(n619) );
  XOR U4306 ( .A(DB[1524]), .B(DB[1509]), .Z(n621) );
  AND U4307 ( .A(n622), .B(n623), .Z(n620) );
  XOR U4308 ( .A(n624), .B(n625), .Z(n623) );
  XOR U4309 ( .A(DB[1509]), .B(DB[1494]), .Z(n625) );
  AND U4310 ( .A(n626), .B(n627), .Z(n624) );
  XOR U4311 ( .A(n628), .B(n629), .Z(n627) );
  XOR U4312 ( .A(DB[1494]), .B(DB[1479]), .Z(n629) );
  AND U4313 ( .A(n630), .B(n631), .Z(n628) );
  XOR U4314 ( .A(n632), .B(n633), .Z(n631) );
  XOR U4315 ( .A(DB[1479]), .B(DB[1464]), .Z(n633) );
  AND U4316 ( .A(n634), .B(n635), .Z(n632) );
  XOR U4317 ( .A(n636), .B(n637), .Z(n635) );
  XOR U4318 ( .A(DB[1464]), .B(DB[1449]), .Z(n637) );
  AND U4319 ( .A(n638), .B(n639), .Z(n636) );
  XOR U4320 ( .A(n640), .B(n641), .Z(n639) );
  XOR U4321 ( .A(DB[1449]), .B(DB[1434]), .Z(n641) );
  AND U4322 ( .A(n642), .B(n643), .Z(n640) );
  XOR U4323 ( .A(n644), .B(n645), .Z(n643) );
  XOR U4324 ( .A(DB[1434]), .B(DB[1419]), .Z(n645) );
  AND U4325 ( .A(n646), .B(n647), .Z(n644) );
  XOR U4326 ( .A(n648), .B(n649), .Z(n647) );
  XOR U4327 ( .A(DB[1419]), .B(DB[1404]), .Z(n649) );
  AND U4328 ( .A(n650), .B(n651), .Z(n648) );
  XOR U4329 ( .A(n652), .B(n653), .Z(n651) );
  XOR U4330 ( .A(DB[1404]), .B(DB[1389]), .Z(n653) );
  AND U4331 ( .A(n654), .B(n655), .Z(n652) );
  XOR U4332 ( .A(n656), .B(n657), .Z(n655) );
  XOR U4333 ( .A(DB[1389]), .B(DB[1374]), .Z(n657) );
  AND U4334 ( .A(n658), .B(n659), .Z(n656) );
  XOR U4335 ( .A(n660), .B(n661), .Z(n659) );
  XOR U4336 ( .A(DB[1374]), .B(DB[1359]), .Z(n661) );
  AND U4337 ( .A(n662), .B(n663), .Z(n660) );
  XOR U4338 ( .A(n664), .B(n665), .Z(n663) );
  XOR U4339 ( .A(DB[1359]), .B(DB[1344]), .Z(n665) );
  AND U4340 ( .A(n666), .B(n667), .Z(n664) );
  XOR U4341 ( .A(n668), .B(n669), .Z(n667) );
  XOR U4342 ( .A(DB[1344]), .B(DB[1329]), .Z(n669) );
  AND U4343 ( .A(n670), .B(n671), .Z(n668) );
  XOR U4344 ( .A(n672), .B(n673), .Z(n671) );
  XOR U4345 ( .A(DB[1329]), .B(DB[1314]), .Z(n673) );
  AND U4346 ( .A(n674), .B(n675), .Z(n672) );
  XOR U4347 ( .A(n676), .B(n677), .Z(n675) );
  XOR U4348 ( .A(DB[1314]), .B(DB[1299]), .Z(n677) );
  AND U4349 ( .A(n678), .B(n679), .Z(n676) );
  XOR U4350 ( .A(n680), .B(n681), .Z(n679) );
  XOR U4351 ( .A(DB[1299]), .B(DB[1284]), .Z(n681) );
  AND U4352 ( .A(n682), .B(n683), .Z(n680) );
  XOR U4353 ( .A(n684), .B(n685), .Z(n683) );
  XOR U4354 ( .A(DB[1284]), .B(DB[1269]), .Z(n685) );
  AND U4355 ( .A(n686), .B(n687), .Z(n684) );
  XOR U4356 ( .A(n688), .B(n689), .Z(n687) );
  XOR U4357 ( .A(DB[1269]), .B(DB[1254]), .Z(n689) );
  AND U4358 ( .A(n690), .B(n691), .Z(n688) );
  XOR U4359 ( .A(n692), .B(n693), .Z(n691) );
  XOR U4360 ( .A(DB[1254]), .B(DB[1239]), .Z(n693) );
  AND U4361 ( .A(n694), .B(n695), .Z(n692) );
  XOR U4362 ( .A(n696), .B(n697), .Z(n695) );
  XOR U4363 ( .A(DB[1239]), .B(DB[1224]), .Z(n697) );
  AND U4364 ( .A(n698), .B(n699), .Z(n696) );
  XOR U4365 ( .A(n700), .B(n701), .Z(n699) );
  XOR U4366 ( .A(DB[1224]), .B(DB[1209]), .Z(n701) );
  AND U4367 ( .A(n702), .B(n703), .Z(n700) );
  XOR U4368 ( .A(n704), .B(n705), .Z(n703) );
  XOR U4369 ( .A(DB[1209]), .B(DB[1194]), .Z(n705) );
  AND U4370 ( .A(n706), .B(n707), .Z(n704) );
  XOR U4371 ( .A(n708), .B(n709), .Z(n707) );
  XOR U4372 ( .A(DB[1194]), .B(DB[1179]), .Z(n709) );
  AND U4373 ( .A(n710), .B(n711), .Z(n708) );
  XOR U4374 ( .A(n712), .B(n713), .Z(n711) );
  XOR U4375 ( .A(DB[1179]), .B(DB[1164]), .Z(n713) );
  AND U4376 ( .A(n714), .B(n715), .Z(n712) );
  XOR U4377 ( .A(n716), .B(n717), .Z(n715) );
  XOR U4378 ( .A(DB[1164]), .B(DB[1149]), .Z(n717) );
  AND U4379 ( .A(n718), .B(n719), .Z(n716) );
  XOR U4380 ( .A(n720), .B(n721), .Z(n719) );
  XOR U4381 ( .A(DB[1149]), .B(DB[1134]), .Z(n721) );
  AND U4382 ( .A(n722), .B(n723), .Z(n720) );
  XOR U4383 ( .A(n724), .B(n725), .Z(n723) );
  XOR U4384 ( .A(DB[1134]), .B(DB[1119]), .Z(n725) );
  AND U4385 ( .A(n726), .B(n727), .Z(n724) );
  XOR U4386 ( .A(n728), .B(n729), .Z(n727) );
  XOR U4387 ( .A(DB[1119]), .B(DB[1104]), .Z(n729) );
  AND U4388 ( .A(n730), .B(n731), .Z(n728) );
  XOR U4389 ( .A(n732), .B(n733), .Z(n731) );
  XOR U4390 ( .A(DB[1104]), .B(DB[1089]), .Z(n733) );
  AND U4391 ( .A(n734), .B(n735), .Z(n732) );
  XOR U4392 ( .A(n736), .B(n737), .Z(n735) );
  XOR U4393 ( .A(DB[1089]), .B(DB[1074]), .Z(n737) );
  AND U4394 ( .A(n738), .B(n739), .Z(n736) );
  XOR U4395 ( .A(n740), .B(n741), .Z(n739) );
  XOR U4396 ( .A(DB[1074]), .B(DB[1059]), .Z(n741) );
  AND U4397 ( .A(n742), .B(n743), .Z(n740) );
  XOR U4398 ( .A(n744), .B(n745), .Z(n743) );
  XOR U4399 ( .A(DB[1059]), .B(DB[1044]), .Z(n745) );
  AND U4400 ( .A(n746), .B(n747), .Z(n744) );
  XOR U4401 ( .A(n748), .B(n749), .Z(n747) );
  XOR U4402 ( .A(DB[1044]), .B(DB[1029]), .Z(n749) );
  AND U4403 ( .A(n750), .B(n751), .Z(n748) );
  XOR U4404 ( .A(n752), .B(n753), .Z(n751) );
  XOR U4405 ( .A(DB[1029]), .B(DB[1014]), .Z(n753) );
  AND U4406 ( .A(n754), .B(n755), .Z(n752) );
  XOR U4407 ( .A(n756), .B(n757), .Z(n755) );
  XOR U4408 ( .A(DB[999]), .B(DB[1014]), .Z(n757) );
  AND U4409 ( .A(n758), .B(n759), .Z(n756) );
  XOR U4410 ( .A(n760), .B(n761), .Z(n759) );
  XOR U4411 ( .A(DB[999]), .B(DB[984]), .Z(n761) );
  AND U4412 ( .A(n762), .B(n763), .Z(n760) );
  XOR U4413 ( .A(n764), .B(n765), .Z(n763) );
  XOR U4414 ( .A(DB[984]), .B(DB[969]), .Z(n765) );
  AND U4415 ( .A(n766), .B(n767), .Z(n764) );
  XOR U4416 ( .A(n768), .B(n769), .Z(n767) );
  XOR U4417 ( .A(DB[969]), .B(DB[954]), .Z(n769) );
  AND U4418 ( .A(n770), .B(n771), .Z(n768) );
  XOR U4419 ( .A(n772), .B(n773), .Z(n771) );
  XOR U4420 ( .A(DB[954]), .B(DB[939]), .Z(n773) );
  AND U4421 ( .A(n774), .B(n775), .Z(n772) );
  XOR U4422 ( .A(n776), .B(n777), .Z(n775) );
  XOR U4423 ( .A(DB[939]), .B(DB[924]), .Z(n777) );
  AND U4424 ( .A(n778), .B(n779), .Z(n776) );
  XOR U4425 ( .A(n780), .B(n781), .Z(n779) );
  XOR U4426 ( .A(DB[924]), .B(DB[909]), .Z(n781) );
  AND U4427 ( .A(n782), .B(n783), .Z(n780) );
  XOR U4428 ( .A(n784), .B(n785), .Z(n783) );
  XOR U4429 ( .A(DB[909]), .B(DB[894]), .Z(n785) );
  AND U4430 ( .A(n786), .B(n787), .Z(n784) );
  XOR U4431 ( .A(n788), .B(n789), .Z(n787) );
  XOR U4432 ( .A(DB[894]), .B(DB[879]), .Z(n789) );
  AND U4433 ( .A(n790), .B(n791), .Z(n788) );
  XOR U4434 ( .A(n792), .B(n793), .Z(n791) );
  XOR U4435 ( .A(DB[879]), .B(DB[864]), .Z(n793) );
  AND U4436 ( .A(n794), .B(n795), .Z(n792) );
  XOR U4437 ( .A(n796), .B(n797), .Z(n795) );
  XOR U4438 ( .A(DB[864]), .B(DB[849]), .Z(n797) );
  AND U4439 ( .A(n798), .B(n799), .Z(n796) );
  XOR U4440 ( .A(n800), .B(n801), .Z(n799) );
  XOR U4441 ( .A(DB[849]), .B(DB[834]), .Z(n801) );
  AND U4442 ( .A(n802), .B(n803), .Z(n800) );
  XOR U4443 ( .A(n804), .B(n805), .Z(n803) );
  XOR U4444 ( .A(DB[834]), .B(DB[819]), .Z(n805) );
  AND U4445 ( .A(n806), .B(n807), .Z(n804) );
  XOR U4446 ( .A(n808), .B(n809), .Z(n807) );
  XOR U4447 ( .A(DB[819]), .B(DB[804]), .Z(n809) );
  AND U4448 ( .A(n810), .B(n811), .Z(n808) );
  XOR U4449 ( .A(n812), .B(n813), .Z(n811) );
  XOR U4450 ( .A(DB[804]), .B(DB[789]), .Z(n813) );
  AND U4451 ( .A(n814), .B(n815), .Z(n812) );
  XOR U4452 ( .A(n816), .B(n817), .Z(n815) );
  XOR U4453 ( .A(DB[789]), .B(DB[774]), .Z(n817) );
  AND U4454 ( .A(n818), .B(n819), .Z(n816) );
  XOR U4455 ( .A(n820), .B(n821), .Z(n819) );
  XOR U4456 ( .A(DB[774]), .B(DB[759]), .Z(n821) );
  AND U4457 ( .A(n822), .B(n823), .Z(n820) );
  XOR U4458 ( .A(n824), .B(n825), .Z(n823) );
  XOR U4459 ( .A(DB[759]), .B(DB[744]), .Z(n825) );
  AND U4460 ( .A(n826), .B(n827), .Z(n824) );
  XOR U4461 ( .A(n828), .B(n829), .Z(n827) );
  XOR U4462 ( .A(DB[744]), .B(DB[729]), .Z(n829) );
  AND U4463 ( .A(n830), .B(n831), .Z(n828) );
  XOR U4464 ( .A(n832), .B(n833), .Z(n831) );
  XOR U4465 ( .A(DB[729]), .B(DB[714]), .Z(n833) );
  AND U4466 ( .A(n834), .B(n835), .Z(n832) );
  XOR U4467 ( .A(n836), .B(n837), .Z(n835) );
  XOR U4468 ( .A(DB[714]), .B(DB[699]), .Z(n837) );
  AND U4469 ( .A(n838), .B(n839), .Z(n836) );
  XOR U4470 ( .A(n840), .B(n841), .Z(n839) );
  XOR U4471 ( .A(DB[699]), .B(DB[684]), .Z(n841) );
  AND U4472 ( .A(n842), .B(n843), .Z(n840) );
  XOR U4473 ( .A(n844), .B(n845), .Z(n843) );
  XOR U4474 ( .A(DB[684]), .B(DB[669]), .Z(n845) );
  AND U4475 ( .A(n846), .B(n847), .Z(n844) );
  XOR U4476 ( .A(n848), .B(n849), .Z(n847) );
  XOR U4477 ( .A(DB[669]), .B(DB[654]), .Z(n849) );
  AND U4478 ( .A(n850), .B(n851), .Z(n848) );
  XOR U4479 ( .A(n852), .B(n853), .Z(n851) );
  XOR U4480 ( .A(DB[654]), .B(DB[639]), .Z(n853) );
  AND U4481 ( .A(n854), .B(n855), .Z(n852) );
  XOR U4482 ( .A(n856), .B(n857), .Z(n855) );
  XOR U4483 ( .A(DB[639]), .B(DB[624]), .Z(n857) );
  AND U4484 ( .A(n858), .B(n859), .Z(n856) );
  XOR U4485 ( .A(n860), .B(n861), .Z(n859) );
  XOR U4486 ( .A(DB[624]), .B(DB[609]), .Z(n861) );
  AND U4487 ( .A(n862), .B(n863), .Z(n860) );
  XOR U4488 ( .A(n864), .B(n865), .Z(n863) );
  XOR U4489 ( .A(DB[609]), .B(DB[594]), .Z(n865) );
  AND U4490 ( .A(n866), .B(n867), .Z(n864) );
  XOR U4491 ( .A(n868), .B(n869), .Z(n867) );
  XOR U4492 ( .A(DB[594]), .B(DB[579]), .Z(n869) );
  AND U4493 ( .A(n870), .B(n871), .Z(n868) );
  XOR U4494 ( .A(n872), .B(n873), .Z(n871) );
  XOR U4495 ( .A(DB[579]), .B(DB[564]), .Z(n873) );
  AND U4496 ( .A(n874), .B(n875), .Z(n872) );
  XOR U4497 ( .A(n876), .B(n877), .Z(n875) );
  XOR U4498 ( .A(DB[564]), .B(DB[549]), .Z(n877) );
  AND U4499 ( .A(n878), .B(n879), .Z(n876) );
  XOR U4500 ( .A(n880), .B(n881), .Z(n879) );
  XOR U4501 ( .A(DB[549]), .B(DB[534]), .Z(n881) );
  AND U4502 ( .A(n882), .B(n883), .Z(n880) );
  XOR U4503 ( .A(n884), .B(n885), .Z(n883) );
  XOR U4504 ( .A(DB[534]), .B(DB[519]), .Z(n885) );
  AND U4505 ( .A(n886), .B(n887), .Z(n884) );
  XOR U4506 ( .A(n888), .B(n889), .Z(n887) );
  XOR U4507 ( .A(DB[519]), .B(DB[504]), .Z(n889) );
  AND U4508 ( .A(n890), .B(n891), .Z(n888) );
  XOR U4509 ( .A(n892), .B(n893), .Z(n891) );
  XOR U4510 ( .A(DB[504]), .B(DB[489]), .Z(n893) );
  AND U4511 ( .A(n894), .B(n895), .Z(n892) );
  XOR U4512 ( .A(n896), .B(n897), .Z(n895) );
  XOR U4513 ( .A(DB[489]), .B(DB[474]), .Z(n897) );
  AND U4514 ( .A(n898), .B(n899), .Z(n896) );
  XOR U4515 ( .A(n900), .B(n901), .Z(n899) );
  XOR U4516 ( .A(DB[474]), .B(DB[459]), .Z(n901) );
  AND U4517 ( .A(n902), .B(n903), .Z(n900) );
  XOR U4518 ( .A(n904), .B(n905), .Z(n903) );
  XOR U4519 ( .A(DB[459]), .B(DB[444]), .Z(n905) );
  AND U4520 ( .A(n906), .B(n907), .Z(n904) );
  XOR U4521 ( .A(n908), .B(n909), .Z(n907) );
  XOR U4522 ( .A(DB[444]), .B(DB[429]), .Z(n909) );
  AND U4523 ( .A(n910), .B(n911), .Z(n908) );
  XOR U4524 ( .A(n912), .B(n913), .Z(n911) );
  XOR U4525 ( .A(DB[429]), .B(DB[414]), .Z(n913) );
  AND U4526 ( .A(n914), .B(n915), .Z(n912) );
  XOR U4527 ( .A(n916), .B(n917), .Z(n915) );
  XOR U4528 ( .A(DB[414]), .B(DB[399]), .Z(n917) );
  AND U4529 ( .A(n918), .B(n919), .Z(n916) );
  XOR U4530 ( .A(n920), .B(n921), .Z(n919) );
  XOR U4531 ( .A(DB[399]), .B(DB[384]), .Z(n921) );
  AND U4532 ( .A(n922), .B(n923), .Z(n920) );
  XOR U4533 ( .A(n924), .B(n925), .Z(n923) );
  XOR U4534 ( .A(DB[384]), .B(DB[369]), .Z(n925) );
  AND U4535 ( .A(n926), .B(n927), .Z(n924) );
  XOR U4536 ( .A(n928), .B(n929), .Z(n927) );
  XOR U4537 ( .A(DB[369]), .B(DB[354]), .Z(n929) );
  AND U4538 ( .A(n930), .B(n931), .Z(n928) );
  XOR U4539 ( .A(n932), .B(n933), .Z(n931) );
  XOR U4540 ( .A(DB[354]), .B(DB[339]), .Z(n933) );
  AND U4541 ( .A(n934), .B(n935), .Z(n932) );
  XOR U4542 ( .A(n936), .B(n937), .Z(n935) );
  XOR U4543 ( .A(DB[339]), .B(DB[324]), .Z(n937) );
  AND U4544 ( .A(n938), .B(n939), .Z(n936) );
  XOR U4545 ( .A(n940), .B(n941), .Z(n939) );
  XOR U4546 ( .A(DB[324]), .B(DB[309]), .Z(n941) );
  AND U4547 ( .A(n942), .B(n943), .Z(n940) );
  XOR U4548 ( .A(n944), .B(n945), .Z(n943) );
  XOR U4549 ( .A(DB[309]), .B(DB[294]), .Z(n945) );
  AND U4550 ( .A(n946), .B(n947), .Z(n944) );
  XOR U4551 ( .A(n948), .B(n949), .Z(n947) );
  XOR U4552 ( .A(DB[294]), .B(DB[279]), .Z(n949) );
  AND U4553 ( .A(n950), .B(n951), .Z(n948) );
  XOR U4554 ( .A(n952), .B(n953), .Z(n951) );
  XOR U4555 ( .A(DB[279]), .B(DB[264]), .Z(n953) );
  AND U4556 ( .A(n954), .B(n955), .Z(n952) );
  XOR U4557 ( .A(n956), .B(n957), .Z(n955) );
  XOR U4558 ( .A(DB[264]), .B(DB[249]), .Z(n957) );
  AND U4559 ( .A(n958), .B(n959), .Z(n956) );
  XOR U4560 ( .A(n960), .B(n961), .Z(n959) );
  XOR U4561 ( .A(DB[249]), .B(DB[234]), .Z(n961) );
  AND U4562 ( .A(n962), .B(n963), .Z(n960) );
  XOR U4563 ( .A(n964), .B(n965), .Z(n963) );
  XOR U4564 ( .A(DB[234]), .B(DB[219]), .Z(n965) );
  AND U4565 ( .A(n966), .B(n967), .Z(n964) );
  XOR U4566 ( .A(n968), .B(n969), .Z(n967) );
  XOR U4567 ( .A(DB[219]), .B(DB[204]), .Z(n969) );
  AND U4568 ( .A(n970), .B(n971), .Z(n968) );
  XOR U4569 ( .A(n972), .B(n973), .Z(n971) );
  XOR U4570 ( .A(DB[204]), .B(DB[189]), .Z(n973) );
  AND U4571 ( .A(n974), .B(n975), .Z(n972) );
  XOR U4572 ( .A(n976), .B(n977), .Z(n975) );
  XOR U4573 ( .A(DB[189]), .B(DB[174]), .Z(n977) );
  AND U4574 ( .A(n978), .B(n979), .Z(n976) );
  XOR U4575 ( .A(n980), .B(n981), .Z(n979) );
  XOR U4576 ( .A(DB[174]), .B(DB[159]), .Z(n981) );
  AND U4577 ( .A(n982), .B(n983), .Z(n980) );
  XOR U4578 ( .A(n984), .B(n985), .Z(n983) );
  XOR U4579 ( .A(DB[159]), .B(DB[144]), .Z(n985) );
  AND U4580 ( .A(n986), .B(n987), .Z(n984) );
  XOR U4581 ( .A(n988), .B(n989), .Z(n987) );
  XOR U4582 ( .A(DB[144]), .B(DB[129]), .Z(n989) );
  AND U4583 ( .A(n990), .B(n991), .Z(n988) );
  XOR U4584 ( .A(n992), .B(n993), .Z(n991) );
  XOR U4585 ( .A(DB[129]), .B(DB[114]), .Z(n993) );
  AND U4586 ( .A(n994), .B(n995), .Z(n992) );
  XOR U4587 ( .A(n996), .B(n997), .Z(n995) );
  XOR U4588 ( .A(DB[99]), .B(DB[114]), .Z(n997) );
  AND U4589 ( .A(n998), .B(n999), .Z(n996) );
  XOR U4590 ( .A(n1000), .B(n1001), .Z(n999) );
  XOR U4591 ( .A(DB[99]), .B(DB[84]), .Z(n1001) );
  AND U4592 ( .A(n1002), .B(n1003), .Z(n1000) );
  XOR U4593 ( .A(n1004), .B(n1005), .Z(n1003) );
  XOR U4594 ( .A(DB[84]), .B(DB[69]), .Z(n1005) );
  AND U4595 ( .A(n1006), .B(n1007), .Z(n1004) );
  XOR U4596 ( .A(n1008), .B(n1009), .Z(n1007) );
  XOR U4597 ( .A(DB[69]), .B(DB[54]), .Z(n1009) );
  AND U4598 ( .A(n1010), .B(n1011), .Z(n1008) );
  XOR U4599 ( .A(n1012), .B(n1013), .Z(n1011) );
  XOR U4600 ( .A(DB[54]), .B(DB[39]), .Z(n1013) );
  AND U4601 ( .A(n1014), .B(n1015), .Z(n1012) );
  XOR U4602 ( .A(n1016), .B(n1017), .Z(n1015) );
  XOR U4603 ( .A(DB[39]), .B(DB[24]), .Z(n1017) );
  AND U4604 ( .A(n1018), .B(n1019), .Z(n1016) );
  XOR U4605 ( .A(DB[9]), .B(DB[24]), .Z(n1019) );
  XOR U4606 ( .A(DB[3833]), .B(n1020), .Z(min_val_out[8]) );
  AND U4607 ( .A(n2), .B(n1021), .Z(n1020) );
  XOR U4608 ( .A(n1022), .B(n1023), .Z(n1021) );
  XOR U4609 ( .A(DB[3833]), .B(DB[3818]), .Z(n1023) );
  AND U4610 ( .A(n6), .B(n1024), .Z(n1022) );
  XOR U4611 ( .A(n1025), .B(n1026), .Z(n1024) );
  XOR U4612 ( .A(DB[3818]), .B(DB[3803]), .Z(n1026) );
  AND U4613 ( .A(n10), .B(n1027), .Z(n1025) );
  XOR U4614 ( .A(n1028), .B(n1029), .Z(n1027) );
  XOR U4615 ( .A(DB[3803]), .B(DB[3788]), .Z(n1029) );
  AND U4616 ( .A(n14), .B(n1030), .Z(n1028) );
  XOR U4617 ( .A(n1031), .B(n1032), .Z(n1030) );
  XOR U4618 ( .A(DB[3788]), .B(DB[3773]), .Z(n1032) );
  AND U4619 ( .A(n18), .B(n1033), .Z(n1031) );
  XOR U4620 ( .A(n1034), .B(n1035), .Z(n1033) );
  XOR U4621 ( .A(DB[3773]), .B(DB[3758]), .Z(n1035) );
  AND U4622 ( .A(n22), .B(n1036), .Z(n1034) );
  XOR U4623 ( .A(n1037), .B(n1038), .Z(n1036) );
  XOR U4624 ( .A(DB[3758]), .B(DB[3743]), .Z(n1038) );
  AND U4625 ( .A(n26), .B(n1039), .Z(n1037) );
  XOR U4626 ( .A(n1040), .B(n1041), .Z(n1039) );
  XOR U4627 ( .A(DB[3743]), .B(DB[3728]), .Z(n1041) );
  AND U4628 ( .A(n30), .B(n1042), .Z(n1040) );
  XOR U4629 ( .A(n1043), .B(n1044), .Z(n1042) );
  XOR U4630 ( .A(DB[3728]), .B(DB[3713]), .Z(n1044) );
  AND U4631 ( .A(n34), .B(n1045), .Z(n1043) );
  XOR U4632 ( .A(n1046), .B(n1047), .Z(n1045) );
  XOR U4633 ( .A(DB[3713]), .B(DB[3698]), .Z(n1047) );
  AND U4634 ( .A(n38), .B(n1048), .Z(n1046) );
  XOR U4635 ( .A(n1049), .B(n1050), .Z(n1048) );
  XOR U4636 ( .A(DB[3698]), .B(DB[3683]), .Z(n1050) );
  AND U4637 ( .A(n42), .B(n1051), .Z(n1049) );
  XOR U4638 ( .A(n1052), .B(n1053), .Z(n1051) );
  XOR U4639 ( .A(DB[3683]), .B(DB[3668]), .Z(n1053) );
  AND U4640 ( .A(n46), .B(n1054), .Z(n1052) );
  XOR U4641 ( .A(n1055), .B(n1056), .Z(n1054) );
  XOR U4642 ( .A(DB[3668]), .B(DB[3653]), .Z(n1056) );
  AND U4643 ( .A(n50), .B(n1057), .Z(n1055) );
  XOR U4644 ( .A(n1058), .B(n1059), .Z(n1057) );
  XOR U4645 ( .A(DB[3653]), .B(DB[3638]), .Z(n1059) );
  AND U4646 ( .A(n54), .B(n1060), .Z(n1058) );
  XOR U4647 ( .A(n1061), .B(n1062), .Z(n1060) );
  XOR U4648 ( .A(DB[3638]), .B(DB[3623]), .Z(n1062) );
  AND U4649 ( .A(n58), .B(n1063), .Z(n1061) );
  XOR U4650 ( .A(n1064), .B(n1065), .Z(n1063) );
  XOR U4651 ( .A(DB[3623]), .B(DB[3608]), .Z(n1065) );
  AND U4652 ( .A(n62), .B(n1066), .Z(n1064) );
  XOR U4653 ( .A(n1067), .B(n1068), .Z(n1066) );
  XOR U4654 ( .A(DB[3608]), .B(DB[3593]), .Z(n1068) );
  AND U4655 ( .A(n66), .B(n1069), .Z(n1067) );
  XOR U4656 ( .A(n1070), .B(n1071), .Z(n1069) );
  XOR U4657 ( .A(DB[3593]), .B(DB[3578]), .Z(n1071) );
  AND U4658 ( .A(n70), .B(n1072), .Z(n1070) );
  XOR U4659 ( .A(n1073), .B(n1074), .Z(n1072) );
  XOR U4660 ( .A(DB[3578]), .B(DB[3563]), .Z(n1074) );
  AND U4661 ( .A(n74), .B(n1075), .Z(n1073) );
  XOR U4662 ( .A(n1076), .B(n1077), .Z(n1075) );
  XOR U4663 ( .A(DB[3563]), .B(DB[3548]), .Z(n1077) );
  AND U4664 ( .A(n78), .B(n1078), .Z(n1076) );
  XOR U4665 ( .A(n1079), .B(n1080), .Z(n1078) );
  XOR U4666 ( .A(DB[3548]), .B(DB[3533]), .Z(n1080) );
  AND U4667 ( .A(n82), .B(n1081), .Z(n1079) );
  XOR U4668 ( .A(n1082), .B(n1083), .Z(n1081) );
  XOR U4669 ( .A(DB[3533]), .B(DB[3518]), .Z(n1083) );
  AND U4670 ( .A(n86), .B(n1084), .Z(n1082) );
  XOR U4671 ( .A(n1085), .B(n1086), .Z(n1084) );
  XOR U4672 ( .A(DB[3518]), .B(DB[3503]), .Z(n1086) );
  AND U4673 ( .A(n90), .B(n1087), .Z(n1085) );
  XOR U4674 ( .A(n1088), .B(n1089), .Z(n1087) );
  XOR U4675 ( .A(DB[3503]), .B(DB[3488]), .Z(n1089) );
  AND U4676 ( .A(n94), .B(n1090), .Z(n1088) );
  XOR U4677 ( .A(n1091), .B(n1092), .Z(n1090) );
  XOR U4678 ( .A(DB[3488]), .B(DB[3473]), .Z(n1092) );
  AND U4679 ( .A(n98), .B(n1093), .Z(n1091) );
  XOR U4680 ( .A(n1094), .B(n1095), .Z(n1093) );
  XOR U4681 ( .A(DB[3473]), .B(DB[3458]), .Z(n1095) );
  AND U4682 ( .A(n102), .B(n1096), .Z(n1094) );
  XOR U4683 ( .A(n1097), .B(n1098), .Z(n1096) );
  XOR U4684 ( .A(DB[3458]), .B(DB[3443]), .Z(n1098) );
  AND U4685 ( .A(n106), .B(n1099), .Z(n1097) );
  XOR U4686 ( .A(n1100), .B(n1101), .Z(n1099) );
  XOR U4687 ( .A(DB[3443]), .B(DB[3428]), .Z(n1101) );
  AND U4688 ( .A(n110), .B(n1102), .Z(n1100) );
  XOR U4689 ( .A(n1103), .B(n1104), .Z(n1102) );
  XOR U4690 ( .A(DB[3428]), .B(DB[3413]), .Z(n1104) );
  AND U4691 ( .A(n114), .B(n1105), .Z(n1103) );
  XOR U4692 ( .A(n1106), .B(n1107), .Z(n1105) );
  XOR U4693 ( .A(DB[3413]), .B(DB[3398]), .Z(n1107) );
  AND U4694 ( .A(n118), .B(n1108), .Z(n1106) );
  XOR U4695 ( .A(n1109), .B(n1110), .Z(n1108) );
  XOR U4696 ( .A(DB[3398]), .B(DB[3383]), .Z(n1110) );
  AND U4697 ( .A(n122), .B(n1111), .Z(n1109) );
  XOR U4698 ( .A(n1112), .B(n1113), .Z(n1111) );
  XOR U4699 ( .A(DB[3383]), .B(DB[3368]), .Z(n1113) );
  AND U4700 ( .A(n126), .B(n1114), .Z(n1112) );
  XOR U4701 ( .A(n1115), .B(n1116), .Z(n1114) );
  XOR U4702 ( .A(DB[3368]), .B(DB[3353]), .Z(n1116) );
  AND U4703 ( .A(n130), .B(n1117), .Z(n1115) );
  XOR U4704 ( .A(n1118), .B(n1119), .Z(n1117) );
  XOR U4705 ( .A(DB[3353]), .B(DB[3338]), .Z(n1119) );
  AND U4706 ( .A(n134), .B(n1120), .Z(n1118) );
  XOR U4707 ( .A(n1121), .B(n1122), .Z(n1120) );
  XOR U4708 ( .A(DB[3338]), .B(DB[3323]), .Z(n1122) );
  AND U4709 ( .A(n138), .B(n1123), .Z(n1121) );
  XOR U4710 ( .A(n1124), .B(n1125), .Z(n1123) );
  XOR U4711 ( .A(DB[3323]), .B(DB[3308]), .Z(n1125) );
  AND U4712 ( .A(n142), .B(n1126), .Z(n1124) );
  XOR U4713 ( .A(n1127), .B(n1128), .Z(n1126) );
  XOR U4714 ( .A(DB[3308]), .B(DB[3293]), .Z(n1128) );
  AND U4715 ( .A(n146), .B(n1129), .Z(n1127) );
  XOR U4716 ( .A(n1130), .B(n1131), .Z(n1129) );
  XOR U4717 ( .A(DB[3293]), .B(DB[3278]), .Z(n1131) );
  AND U4718 ( .A(n150), .B(n1132), .Z(n1130) );
  XOR U4719 ( .A(n1133), .B(n1134), .Z(n1132) );
  XOR U4720 ( .A(DB[3278]), .B(DB[3263]), .Z(n1134) );
  AND U4721 ( .A(n154), .B(n1135), .Z(n1133) );
  XOR U4722 ( .A(n1136), .B(n1137), .Z(n1135) );
  XOR U4723 ( .A(DB[3263]), .B(DB[3248]), .Z(n1137) );
  AND U4724 ( .A(n158), .B(n1138), .Z(n1136) );
  XOR U4725 ( .A(n1139), .B(n1140), .Z(n1138) );
  XOR U4726 ( .A(DB[3248]), .B(DB[3233]), .Z(n1140) );
  AND U4727 ( .A(n162), .B(n1141), .Z(n1139) );
  XOR U4728 ( .A(n1142), .B(n1143), .Z(n1141) );
  XOR U4729 ( .A(DB[3233]), .B(DB[3218]), .Z(n1143) );
  AND U4730 ( .A(n166), .B(n1144), .Z(n1142) );
  XOR U4731 ( .A(n1145), .B(n1146), .Z(n1144) );
  XOR U4732 ( .A(DB[3218]), .B(DB[3203]), .Z(n1146) );
  AND U4733 ( .A(n170), .B(n1147), .Z(n1145) );
  XOR U4734 ( .A(n1148), .B(n1149), .Z(n1147) );
  XOR U4735 ( .A(DB[3203]), .B(DB[3188]), .Z(n1149) );
  AND U4736 ( .A(n174), .B(n1150), .Z(n1148) );
  XOR U4737 ( .A(n1151), .B(n1152), .Z(n1150) );
  XOR U4738 ( .A(DB[3188]), .B(DB[3173]), .Z(n1152) );
  AND U4739 ( .A(n178), .B(n1153), .Z(n1151) );
  XOR U4740 ( .A(n1154), .B(n1155), .Z(n1153) );
  XOR U4741 ( .A(DB[3173]), .B(DB[3158]), .Z(n1155) );
  AND U4742 ( .A(n182), .B(n1156), .Z(n1154) );
  XOR U4743 ( .A(n1157), .B(n1158), .Z(n1156) );
  XOR U4744 ( .A(DB[3158]), .B(DB[3143]), .Z(n1158) );
  AND U4745 ( .A(n186), .B(n1159), .Z(n1157) );
  XOR U4746 ( .A(n1160), .B(n1161), .Z(n1159) );
  XOR U4747 ( .A(DB[3143]), .B(DB[3128]), .Z(n1161) );
  AND U4748 ( .A(n190), .B(n1162), .Z(n1160) );
  XOR U4749 ( .A(n1163), .B(n1164), .Z(n1162) );
  XOR U4750 ( .A(DB[3128]), .B(DB[3113]), .Z(n1164) );
  AND U4751 ( .A(n194), .B(n1165), .Z(n1163) );
  XOR U4752 ( .A(n1166), .B(n1167), .Z(n1165) );
  XOR U4753 ( .A(DB[3113]), .B(DB[3098]), .Z(n1167) );
  AND U4754 ( .A(n198), .B(n1168), .Z(n1166) );
  XOR U4755 ( .A(n1169), .B(n1170), .Z(n1168) );
  XOR U4756 ( .A(DB[3098]), .B(DB[3083]), .Z(n1170) );
  AND U4757 ( .A(n202), .B(n1171), .Z(n1169) );
  XOR U4758 ( .A(n1172), .B(n1173), .Z(n1171) );
  XOR U4759 ( .A(DB[3083]), .B(DB[3068]), .Z(n1173) );
  AND U4760 ( .A(n206), .B(n1174), .Z(n1172) );
  XOR U4761 ( .A(n1175), .B(n1176), .Z(n1174) );
  XOR U4762 ( .A(DB[3068]), .B(DB[3053]), .Z(n1176) );
  AND U4763 ( .A(n210), .B(n1177), .Z(n1175) );
  XOR U4764 ( .A(n1178), .B(n1179), .Z(n1177) );
  XOR U4765 ( .A(DB[3053]), .B(DB[3038]), .Z(n1179) );
  AND U4766 ( .A(n214), .B(n1180), .Z(n1178) );
  XOR U4767 ( .A(n1181), .B(n1182), .Z(n1180) );
  XOR U4768 ( .A(DB[3038]), .B(DB[3023]), .Z(n1182) );
  AND U4769 ( .A(n218), .B(n1183), .Z(n1181) );
  XOR U4770 ( .A(n1184), .B(n1185), .Z(n1183) );
  XOR U4771 ( .A(DB[3023]), .B(DB[3008]), .Z(n1185) );
  AND U4772 ( .A(n222), .B(n1186), .Z(n1184) );
  XOR U4773 ( .A(n1187), .B(n1188), .Z(n1186) );
  XOR U4774 ( .A(DB[3008]), .B(DB[2993]), .Z(n1188) );
  AND U4775 ( .A(n226), .B(n1189), .Z(n1187) );
  XOR U4776 ( .A(n1190), .B(n1191), .Z(n1189) );
  XOR U4777 ( .A(DB[2993]), .B(DB[2978]), .Z(n1191) );
  AND U4778 ( .A(n230), .B(n1192), .Z(n1190) );
  XOR U4779 ( .A(n1193), .B(n1194), .Z(n1192) );
  XOR U4780 ( .A(DB[2978]), .B(DB[2963]), .Z(n1194) );
  AND U4781 ( .A(n234), .B(n1195), .Z(n1193) );
  XOR U4782 ( .A(n1196), .B(n1197), .Z(n1195) );
  XOR U4783 ( .A(DB[2963]), .B(DB[2948]), .Z(n1197) );
  AND U4784 ( .A(n238), .B(n1198), .Z(n1196) );
  XOR U4785 ( .A(n1199), .B(n1200), .Z(n1198) );
  XOR U4786 ( .A(DB[2948]), .B(DB[2933]), .Z(n1200) );
  AND U4787 ( .A(n242), .B(n1201), .Z(n1199) );
  XOR U4788 ( .A(n1202), .B(n1203), .Z(n1201) );
  XOR U4789 ( .A(DB[2933]), .B(DB[2918]), .Z(n1203) );
  AND U4790 ( .A(n246), .B(n1204), .Z(n1202) );
  XOR U4791 ( .A(n1205), .B(n1206), .Z(n1204) );
  XOR U4792 ( .A(DB[2918]), .B(DB[2903]), .Z(n1206) );
  AND U4793 ( .A(n250), .B(n1207), .Z(n1205) );
  XOR U4794 ( .A(n1208), .B(n1209), .Z(n1207) );
  XOR U4795 ( .A(DB[2903]), .B(DB[2888]), .Z(n1209) );
  AND U4796 ( .A(n254), .B(n1210), .Z(n1208) );
  XOR U4797 ( .A(n1211), .B(n1212), .Z(n1210) );
  XOR U4798 ( .A(DB[2888]), .B(DB[2873]), .Z(n1212) );
  AND U4799 ( .A(n258), .B(n1213), .Z(n1211) );
  XOR U4800 ( .A(n1214), .B(n1215), .Z(n1213) );
  XOR U4801 ( .A(DB[2873]), .B(DB[2858]), .Z(n1215) );
  AND U4802 ( .A(n262), .B(n1216), .Z(n1214) );
  XOR U4803 ( .A(n1217), .B(n1218), .Z(n1216) );
  XOR U4804 ( .A(DB[2858]), .B(DB[2843]), .Z(n1218) );
  AND U4805 ( .A(n266), .B(n1219), .Z(n1217) );
  XOR U4806 ( .A(n1220), .B(n1221), .Z(n1219) );
  XOR U4807 ( .A(DB[2843]), .B(DB[2828]), .Z(n1221) );
  AND U4808 ( .A(n270), .B(n1222), .Z(n1220) );
  XOR U4809 ( .A(n1223), .B(n1224), .Z(n1222) );
  XOR U4810 ( .A(DB[2828]), .B(DB[2813]), .Z(n1224) );
  AND U4811 ( .A(n274), .B(n1225), .Z(n1223) );
  XOR U4812 ( .A(n1226), .B(n1227), .Z(n1225) );
  XOR U4813 ( .A(DB[2813]), .B(DB[2798]), .Z(n1227) );
  AND U4814 ( .A(n278), .B(n1228), .Z(n1226) );
  XOR U4815 ( .A(n1229), .B(n1230), .Z(n1228) );
  XOR U4816 ( .A(DB[2798]), .B(DB[2783]), .Z(n1230) );
  AND U4817 ( .A(n282), .B(n1231), .Z(n1229) );
  XOR U4818 ( .A(n1232), .B(n1233), .Z(n1231) );
  XOR U4819 ( .A(DB[2783]), .B(DB[2768]), .Z(n1233) );
  AND U4820 ( .A(n286), .B(n1234), .Z(n1232) );
  XOR U4821 ( .A(n1235), .B(n1236), .Z(n1234) );
  XOR U4822 ( .A(DB[2768]), .B(DB[2753]), .Z(n1236) );
  AND U4823 ( .A(n290), .B(n1237), .Z(n1235) );
  XOR U4824 ( .A(n1238), .B(n1239), .Z(n1237) );
  XOR U4825 ( .A(DB[2753]), .B(DB[2738]), .Z(n1239) );
  AND U4826 ( .A(n294), .B(n1240), .Z(n1238) );
  XOR U4827 ( .A(n1241), .B(n1242), .Z(n1240) );
  XOR U4828 ( .A(DB[2738]), .B(DB[2723]), .Z(n1242) );
  AND U4829 ( .A(n298), .B(n1243), .Z(n1241) );
  XOR U4830 ( .A(n1244), .B(n1245), .Z(n1243) );
  XOR U4831 ( .A(DB[2723]), .B(DB[2708]), .Z(n1245) );
  AND U4832 ( .A(n302), .B(n1246), .Z(n1244) );
  XOR U4833 ( .A(n1247), .B(n1248), .Z(n1246) );
  XOR U4834 ( .A(DB[2708]), .B(DB[2693]), .Z(n1248) );
  AND U4835 ( .A(n306), .B(n1249), .Z(n1247) );
  XOR U4836 ( .A(n1250), .B(n1251), .Z(n1249) );
  XOR U4837 ( .A(DB[2693]), .B(DB[2678]), .Z(n1251) );
  AND U4838 ( .A(n310), .B(n1252), .Z(n1250) );
  XOR U4839 ( .A(n1253), .B(n1254), .Z(n1252) );
  XOR U4840 ( .A(DB[2678]), .B(DB[2663]), .Z(n1254) );
  AND U4841 ( .A(n314), .B(n1255), .Z(n1253) );
  XOR U4842 ( .A(n1256), .B(n1257), .Z(n1255) );
  XOR U4843 ( .A(DB[2663]), .B(DB[2648]), .Z(n1257) );
  AND U4844 ( .A(n318), .B(n1258), .Z(n1256) );
  XOR U4845 ( .A(n1259), .B(n1260), .Z(n1258) );
  XOR U4846 ( .A(DB[2648]), .B(DB[2633]), .Z(n1260) );
  AND U4847 ( .A(n322), .B(n1261), .Z(n1259) );
  XOR U4848 ( .A(n1262), .B(n1263), .Z(n1261) );
  XOR U4849 ( .A(DB[2633]), .B(DB[2618]), .Z(n1263) );
  AND U4850 ( .A(n326), .B(n1264), .Z(n1262) );
  XOR U4851 ( .A(n1265), .B(n1266), .Z(n1264) );
  XOR U4852 ( .A(DB[2618]), .B(DB[2603]), .Z(n1266) );
  AND U4853 ( .A(n330), .B(n1267), .Z(n1265) );
  XOR U4854 ( .A(n1268), .B(n1269), .Z(n1267) );
  XOR U4855 ( .A(DB[2603]), .B(DB[2588]), .Z(n1269) );
  AND U4856 ( .A(n334), .B(n1270), .Z(n1268) );
  XOR U4857 ( .A(n1271), .B(n1272), .Z(n1270) );
  XOR U4858 ( .A(DB[2588]), .B(DB[2573]), .Z(n1272) );
  AND U4859 ( .A(n338), .B(n1273), .Z(n1271) );
  XOR U4860 ( .A(n1274), .B(n1275), .Z(n1273) );
  XOR U4861 ( .A(DB[2573]), .B(DB[2558]), .Z(n1275) );
  AND U4862 ( .A(n342), .B(n1276), .Z(n1274) );
  XOR U4863 ( .A(n1277), .B(n1278), .Z(n1276) );
  XOR U4864 ( .A(DB[2558]), .B(DB[2543]), .Z(n1278) );
  AND U4865 ( .A(n346), .B(n1279), .Z(n1277) );
  XOR U4866 ( .A(n1280), .B(n1281), .Z(n1279) );
  XOR U4867 ( .A(DB[2543]), .B(DB[2528]), .Z(n1281) );
  AND U4868 ( .A(n350), .B(n1282), .Z(n1280) );
  XOR U4869 ( .A(n1283), .B(n1284), .Z(n1282) );
  XOR U4870 ( .A(DB[2528]), .B(DB[2513]), .Z(n1284) );
  AND U4871 ( .A(n354), .B(n1285), .Z(n1283) );
  XOR U4872 ( .A(n1286), .B(n1287), .Z(n1285) );
  XOR U4873 ( .A(DB[2513]), .B(DB[2498]), .Z(n1287) );
  AND U4874 ( .A(n358), .B(n1288), .Z(n1286) );
  XOR U4875 ( .A(n1289), .B(n1290), .Z(n1288) );
  XOR U4876 ( .A(DB[2498]), .B(DB[2483]), .Z(n1290) );
  AND U4877 ( .A(n362), .B(n1291), .Z(n1289) );
  XOR U4878 ( .A(n1292), .B(n1293), .Z(n1291) );
  XOR U4879 ( .A(DB[2483]), .B(DB[2468]), .Z(n1293) );
  AND U4880 ( .A(n366), .B(n1294), .Z(n1292) );
  XOR U4881 ( .A(n1295), .B(n1296), .Z(n1294) );
  XOR U4882 ( .A(DB[2468]), .B(DB[2453]), .Z(n1296) );
  AND U4883 ( .A(n370), .B(n1297), .Z(n1295) );
  XOR U4884 ( .A(n1298), .B(n1299), .Z(n1297) );
  XOR U4885 ( .A(DB[2453]), .B(DB[2438]), .Z(n1299) );
  AND U4886 ( .A(n374), .B(n1300), .Z(n1298) );
  XOR U4887 ( .A(n1301), .B(n1302), .Z(n1300) );
  XOR U4888 ( .A(DB[2438]), .B(DB[2423]), .Z(n1302) );
  AND U4889 ( .A(n378), .B(n1303), .Z(n1301) );
  XOR U4890 ( .A(n1304), .B(n1305), .Z(n1303) );
  XOR U4891 ( .A(DB[2423]), .B(DB[2408]), .Z(n1305) );
  AND U4892 ( .A(n382), .B(n1306), .Z(n1304) );
  XOR U4893 ( .A(n1307), .B(n1308), .Z(n1306) );
  XOR U4894 ( .A(DB[2408]), .B(DB[2393]), .Z(n1308) );
  AND U4895 ( .A(n386), .B(n1309), .Z(n1307) );
  XOR U4896 ( .A(n1310), .B(n1311), .Z(n1309) );
  XOR U4897 ( .A(DB[2393]), .B(DB[2378]), .Z(n1311) );
  AND U4898 ( .A(n390), .B(n1312), .Z(n1310) );
  XOR U4899 ( .A(n1313), .B(n1314), .Z(n1312) );
  XOR U4900 ( .A(DB[2378]), .B(DB[2363]), .Z(n1314) );
  AND U4901 ( .A(n394), .B(n1315), .Z(n1313) );
  XOR U4902 ( .A(n1316), .B(n1317), .Z(n1315) );
  XOR U4903 ( .A(DB[2363]), .B(DB[2348]), .Z(n1317) );
  AND U4904 ( .A(n398), .B(n1318), .Z(n1316) );
  XOR U4905 ( .A(n1319), .B(n1320), .Z(n1318) );
  XOR U4906 ( .A(DB[2348]), .B(DB[2333]), .Z(n1320) );
  AND U4907 ( .A(n402), .B(n1321), .Z(n1319) );
  XOR U4908 ( .A(n1322), .B(n1323), .Z(n1321) );
  XOR U4909 ( .A(DB[2333]), .B(DB[2318]), .Z(n1323) );
  AND U4910 ( .A(n406), .B(n1324), .Z(n1322) );
  XOR U4911 ( .A(n1325), .B(n1326), .Z(n1324) );
  XOR U4912 ( .A(DB[2318]), .B(DB[2303]), .Z(n1326) );
  AND U4913 ( .A(n410), .B(n1327), .Z(n1325) );
  XOR U4914 ( .A(n1328), .B(n1329), .Z(n1327) );
  XOR U4915 ( .A(DB[2303]), .B(DB[2288]), .Z(n1329) );
  AND U4916 ( .A(n414), .B(n1330), .Z(n1328) );
  XOR U4917 ( .A(n1331), .B(n1332), .Z(n1330) );
  XOR U4918 ( .A(DB[2288]), .B(DB[2273]), .Z(n1332) );
  AND U4919 ( .A(n418), .B(n1333), .Z(n1331) );
  XOR U4920 ( .A(n1334), .B(n1335), .Z(n1333) );
  XOR U4921 ( .A(DB[2273]), .B(DB[2258]), .Z(n1335) );
  AND U4922 ( .A(n422), .B(n1336), .Z(n1334) );
  XOR U4923 ( .A(n1337), .B(n1338), .Z(n1336) );
  XOR U4924 ( .A(DB[2258]), .B(DB[2243]), .Z(n1338) );
  AND U4925 ( .A(n426), .B(n1339), .Z(n1337) );
  XOR U4926 ( .A(n1340), .B(n1341), .Z(n1339) );
  XOR U4927 ( .A(DB[2243]), .B(DB[2228]), .Z(n1341) );
  AND U4928 ( .A(n430), .B(n1342), .Z(n1340) );
  XOR U4929 ( .A(n1343), .B(n1344), .Z(n1342) );
  XOR U4930 ( .A(DB[2228]), .B(DB[2213]), .Z(n1344) );
  AND U4931 ( .A(n434), .B(n1345), .Z(n1343) );
  XOR U4932 ( .A(n1346), .B(n1347), .Z(n1345) );
  XOR U4933 ( .A(DB[2213]), .B(DB[2198]), .Z(n1347) );
  AND U4934 ( .A(n438), .B(n1348), .Z(n1346) );
  XOR U4935 ( .A(n1349), .B(n1350), .Z(n1348) );
  XOR U4936 ( .A(DB[2198]), .B(DB[2183]), .Z(n1350) );
  AND U4937 ( .A(n442), .B(n1351), .Z(n1349) );
  XOR U4938 ( .A(n1352), .B(n1353), .Z(n1351) );
  XOR U4939 ( .A(DB[2183]), .B(DB[2168]), .Z(n1353) );
  AND U4940 ( .A(n446), .B(n1354), .Z(n1352) );
  XOR U4941 ( .A(n1355), .B(n1356), .Z(n1354) );
  XOR U4942 ( .A(DB[2168]), .B(DB[2153]), .Z(n1356) );
  AND U4943 ( .A(n450), .B(n1357), .Z(n1355) );
  XOR U4944 ( .A(n1358), .B(n1359), .Z(n1357) );
  XOR U4945 ( .A(DB[2153]), .B(DB[2138]), .Z(n1359) );
  AND U4946 ( .A(n454), .B(n1360), .Z(n1358) );
  XOR U4947 ( .A(n1361), .B(n1362), .Z(n1360) );
  XOR U4948 ( .A(DB[2138]), .B(DB[2123]), .Z(n1362) );
  AND U4949 ( .A(n458), .B(n1363), .Z(n1361) );
  XOR U4950 ( .A(n1364), .B(n1365), .Z(n1363) );
  XOR U4951 ( .A(DB[2123]), .B(DB[2108]), .Z(n1365) );
  AND U4952 ( .A(n462), .B(n1366), .Z(n1364) );
  XOR U4953 ( .A(n1367), .B(n1368), .Z(n1366) );
  XOR U4954 ( .A(DB[2108]), .B(DB[2093]), .Z(n1368) );
  AND U4955 ( .A(n466), .B(n1369), .Z(n1367) );
  XOR U4956 ( .A(n1370), .B(n1371), .Z(n1369) );
  XOR U4957 ( .A(DB[2093]), .B(DB[2078]), .Z(n1371) );
  AND U4958 ( .A(n470), .B(n1372), .Z(n1370) );
  XOR U4959 ( .A(n1373), .B(n1374), .Z(n1372) );
  XOR U4960 ( .A(DB[2078]), .B(DB[2063]), .Z(n1374) );
  AND U4961 ( .A(n474), .B(n1375), .Z(n1373) );
  XOR U4962 ( .A(n1376), .B(n1377), .Z(n1375) );
  XOR U4963 ( .A(DB[2063]), .B(DB[2048]), .Z(n1377) );
  AND U4964 ( .A(n478), .B(n1378), .Z(n1376) );
  XOR U4965 ( .A(n1379), .B(n1380), .Z(n1378) );
  XOR U4966 ( .A(DB[2048]), .B(DB[2033]), .Z(n1380) );
  AND U4967 ( .A(n482), .B(n1381), .Z(n1379) );
  XOR U4968 ( .A(n1382), .B(n1383), .Z(n1381) );
  XOR U4969 ( .A(DB[2033]), .B(DB[2018]), .Z(n1383) );
  AND U4970 ( .A(n486), .B(n1384), .Z(n1382) );
  XOR U4971 ( .A(n1385), .B(n1386), .Z(n1384) );
  XOR U4972 ( .A(DB[2018]), .B(DB[2003]), .Z(n1386) );
  AND U4973 ( .A(n490), .B(n1387), .Z(n1385) );
  XOR U4974 ( .A(n1388), .B(n1389), .Z(n1387) );
  XOR U4975 ( .A(DB[2003]), .B(DB[1988]), .Z(n1389) );
  AND U4976 ( .A(n494), .B(n1390), .Z(n1388) );
  XOR U4977 ( .A(n1391), .B(n1392), .Z(n1390) );
  XOR U4978 ( .A(DB[1988]), .B(DB[1973]), .Z(n1392) );
  AND U4979 ( .A(n498), .B(n1393), .Z(n1391) );
  XOR U4980 ( .A(n1394), .B(n1395), .Z(n1393) );
  XOR U4981 ( .A(DB[1973]), .B(DB[1958]), .Z(n1395) );
  AND U4982 ( .A(n502), .B(n1396), .Z(n1394) );
  XOR U4983 ( .A(n1397), .B(n1398), .Z(n1396) );
  XOR U4984 ( .A(DB[1958]), .B(DB[1943]), .Z(n1398) );
  AND U4985 ( .A(n506), .B(n1399), .Z(n1397) );
  XOR U4986 ( .A(n1400), .B(n1401), .Z(n1399) );
  XOR U4987 ( .A(DB[1943]), .B(DB[1928]), .Z(n1401) );
  AND U4988 ( .A(n510), .B(n1402), .Z(n1400) );
  XOR U4989 ( .A(n1403), .B(n1404), .Z(n1402) );
  XOR U4990 ( .A(DB[1928]), .B(DB[1913]), .Z(n1404) );
  AND U4991 ( .A(n514), .B(n1405), .Z(n1403) );
  XOR U4992 ( .A(n1406), .B(n1407), .Z(n1405) );
  XOR U4993 ( .A(DB[1913]), .B(DB[1898]), .Z(n1407) );
  AND U4994 ( .A(n518), .B(n1408), .Z(n1406) );
  XOR U4995 ( .A(n1409), .B(n1410), .Z(n1408) );
  XOR U4996 ( .A(DB[1898]), .B(DB[1883]), .Z(n1410) );
  AND U4997 ( .A(n522), .B(n1411), .Z(n1409) );
  XOR U4998 ( .A(n1412), .B(n1413), .Z(n1411) );
  XOR U4999 ( .A(DB[1883]), .B(DB[1868]), .Z(n1413) );
  AND U5000 ( .A(n526), .B(n1414), .Z(n1412) );
  XOR U5001 ( .A(n1415), .B(n1416), .Z(n1414) );
  XOR U5002 ( .A(DB[1868]), .B(DB[1853]), .Z(n1416) );
  AND U5003 ( .A(n530), .B(n1417), .Z(n1415) );
  XOR U5004 ( .A(n1418), .B(n1419), .Z(n1417) );
  XOR U5005 ( .A(DB[1853]), .B(DB[1838]), .Z(n1419) );
  AND U5006 ( .A(n534), .B(n1420), .Z(n1418) );
  XOR U5007 ( .A(n1421), .B(n1422), .Z(n1420) );
  XOR U5008 ( .A(DB[1838]), .B(DB[1823]), .Z(n1422) );
  AND U5009 ( .A(n538), .B(n1423), .Z(n1421) );
  XOR U5010 ( .A(n1424), .B(n1425), .Z(n1423) );
  XOR U5011 ( .A(DB[1823]), .B(DB[1808]), .Z(n1425) );
  AND U5012 ( .A(n542), .B(n1426), .Z(n1424) );
  XOR U5013 ( .A(n1427), .B(n1428), .Z(n1426) );
  XOR U5014 ( .A(DB[1808]), .B(DB[1793]), .Z(n1428) );
  AND U5015 ( .A(n546), .B(n1429), .Z(n1427) );
  XOR U5016 ( .A(n1430), .B(n1431), .Z(n1429) );
  XOR U5017 ( .A(DB[1793]), .B(DB[1778]), .Z(n1431) );
  AND U5018 ( .A(n550), .B(n1432), .Z(n1430) );
  XOR U5019 ( .A(n1433), .B(n1434), .Z(n1432) );
  XOR U5020 ( .A(DB[1778]), .B(DB[1763]), .Z(n1434) );
  AND U5021 ( .A(n554), .B(n1435), .Z(n1433) );
  XOR U5022 ( .A(n1436), .B(n1437), .Z(n1435) );
  XOR U5023 ( .A(DB[1763]), .B(DB[1748]), .Z(n1437) );
  AND U5024 ( .A(n558), .B(n1438), .Z(n1436) );
  XOR U5025 ( .A(n1439), .B(n1440), .Z(n1438) );
  XOR U5026 ( .A(DB[1748]), .B(DB[1733]), .Z(n1440) );
  AND U5027 ( .A(n562), .B(n1441), .Z(n1439) );
  XOR U5028 ( .A(n1442), .B(n1443), .Z(n1441) );
  XOR U5029 ( .A(DB[1733]), .B(DB[1718]), .Z(n1443) );
  AND U5030 ( .A(n566), .B(n1444), .Z(n1442) );
  XOR U5031 ( .A(n1445), .B(n1446), .Z(n1444) );
  XOR U5032 ( .A(DB[1718]), .B(DB[1703]), .Z(n1446) );
  AND U5033 ( .A(n570), .B(n1447), .Z(n1445) );
  XOR U5034 ( .A(n1448), .B(n1449), .Z(n1447) );
  XOR U5035 ( .A(DB[1703]), .B(DB[1688]), .Z(n1449) );
  AND U5036 ( .A(n574), .B(n1450), .Z(n1448) );
  XOR U5037 ( .A(n1451), .B(n1452), .Z(n1450) );
  XOR U5038 ( .A(DB[1688]), .B(DB[1673]), .Z(n1452) );
  AND U5039 ( .A(n578), .B(n1453), .Z(n1451) );
  XOR U5040 ( .A(n1454), .B(n1455), .Z(n1453) );
  XOR U5041 ( .A(DB[1673]), .B(DB[1658]), .Z(n1455) );
  AND U5042 ( .A(n582), .B(n1456), .Z(n1454) );
  XOR U5043 ( .A(n1457), .B(n1458), .Z(n1456) );
  XOR U5044 ( .A(DB[1658]), .B(DB[1643]), .Z(n1458) );
  AND U5045 ( .A(n586), .B(n1459), .Z(n1457) );
  XOR U5046 ( .A(n1460), .B(n1461), .Z(n1459) );
  XOR U5047 ( .A(DB[1643]), .B(DB[1628]), .Z(n1461) );
  AND U5048 ( .A(n590), .B(n1462), .Z(n1460) );
  XOR U5049 ( .A(n1463), .B(n1464), .Z(n1462) );
  XOR U5050 ( .A(DB[1628]), .B(DB[1613]), .Z(n1464) );
  AND U5051 ( .A(n594), .B(n1465), .Z(n1463) );
  XOR U5052 ( .A(n1466), .B(n1467), .Z(n1465) );
  XOR U5053 ( .A(DB[1613]), .B(DB[1598]), .Z(n1467) );
  AND U5054 ( .A(n598), .B(n1468), .Z(n1466) );
  XOR U5055 ( .A(n1469), .B(n1470), .Z(n1468) );
  XOR U5056 ( .A(DB[1598]), .B(DB[1583]), .Z(n1470) );
  AND U5057 ( .A(n602), .B(n1471), .Z(n1469) );
  XOR U5058 ( .A(n1472), .B(n1473), .Z(n1471) );
  XOR U5059 ( .A(DB[1583]), .B(DB[1568]), .Z(n1473) );
  AND U5060 ( .A(n606), .B(n1474), .Z(n1472) );
  XOR U5061 ( .A(n1475), .B(n1476), .Z(n1474) );
  XOR U5062 ( .A(DB[1568]), .B(DB[1553]), .Z(n1476) );
  AND U5063 ( .A(n610), .B(n1477), .Z(n1475) );
  XOR U5064 ( .A(n1478), .B(n1479), .Z(n1477) );
  XOR U5065 ( .A(DB[1553]), .B(DB[1538]), .Z(n1479) );
  AND U5066 ( .A(n614), .B(n1480), .Z(n1478) );
  XOR U5067 ( .A(n1481), .B(n1482), .Z(n1480) );
  XOR U5068 ( .A(DB[1538]), .B(DB[1523]), .Z(n1482) );
  AND U5069 ( .A(n618), .B(n1483), .Z(n1481) );
  XOR U5070 ( .A(n1484), .B(n1485), .Z(n1483) );
  XOR U5071 ( .A(DB[1523]), .B(DB[1508]), .Z(n1485) );
  AND U5072 ( .A(n622), .B(n1486), .Z(n1484) );
  XOR U5073 ( .A(n1487), .B(n1488), .Z(n1486) );
  XOR U5074 ( .A(DB[1508]), .B(DB[1493]), .Z(n1488) );
  AND U5075 ( .A(n626), .B(n1489), .Z(n1487) );
  XOR U5076 ( .A(n1490), .B(n1491), .Z(n1489) );
  XOR U5077 ( .A(DB[1493]), .B(DB[1478]), .Z(n1491) );
  AND U5078 ( .A(n630), .B(n1492), .Z(n1490) );
  XOR U5079 ( .A(n1493), .B(n1494), .Z(n1492) );
  XOR U5080 ( .A(DB[1478]), .B(DB[1463]), .Z(n1494) );
  AND U5081 ( .A(n634), .B(n1495), .Z(n1493) );
  XOR U5082 ( .A(n1496), .B(n1497), .Z(n1495) );
  XOR U5083 ( .A(DB[1463]), .B(DB[1448]), .Z(n1497) );
  AND U5084 ( .A(n638), .B(n1498), .Z(n1496) );
  XOR U5085 ( .A(n1499), .B(n1500), .Z(n1498) );
  XOR U5086 ( .A(DB[1448]), .B(DB[1433]), .Z(n1500) );
  AND U5087 ( .A(n642), .B(n1501), .Z(n1499) );
  XOR U5088 ( .A(n1502), .B(n1503), .Z(n1501) );
  XOR U5089 ( .A(DB[1433]), .B(DB[1418]), .Z(n1503) );
  AND U5090 ( .A(n646), .B(n1504), .Z(n1502) );
  XOR U5091 ( .A(n1505), .B(n1506), .Z(n1504) );
  XOR U5092 ( .A(DB[1418]), .B(DB[1403]), .Z(n1506) );
  AND U5093 ( .A(n650), .B(n1507), .Z(n1505) );
  XOR U5094 ( .A(n1508), .B(n1509), .Z(n1507) );
  XOR U5095 ( .A(DB[1403]), .B(DB[1388]), .Z(n1509) );
  AND U5096 ( .A(n654), .B(n1510), .Z(n1508) );
  XOR U5097 ( .A(n1511), .B(n1512), .Z(n1510) );
  XOR U5098 ( .A(DB[1388]), .B(DB[1373]), .Z(n1512) );
  AND U5099 ( .A(n658), .B(n1513), .Z(n1511) );
  XOR U5100 ( .A(n1514), .B(n1515), .Z(n1513) );
  XOR U5101 ( .A(DB[1373]), .B(DB[1358]), .Z(n1515) );
  AND U5102 ( .A(n662), .B(n1516), .Z(n1514) );
  XOR U5103 ( .A(n1517), .B(n1518), .Z(n1516) );
  XOR U5104 ( .A(DB[1358]), .B(DB[1343]), .Z(n1518) );
  AND U5105 ( .A(n666), .B(n1519), .Z(n1517) );
  XOR U5106 ( .A(n1520), .B(n1521), .Z(n1519) );
  XOR U5107 ( .A(DB[1343]), .B(DB[1328]), .Z(n1521) );
  AND U5108 ( .A(n670), .B(n1522), .Z(n1520) );
  XOR U5109 ( .A(n1523), .B(n1524), .Z(n1522) );
  XOR U5110 ( .A(DB[1328]), .B(DB[1313]), .Z(n1524) );
  AND U5111 ( .A(n674), .B(n1525), .Z(n1523) );
  XOR U5112 ( .A(n1526), .B(n1527), .Z(n1525) );
  XOR U5113 ( .A(DB[1313]), .B(DB[1298]), .Z(n1527) );
  AND U5114 ( .A(n678), .B(n1528), .Z(n1526) );
  XOR U5115 ( .A(n1529), .B(n1530), .Z(n1528) );
  XOR U5116 ( .A(DB[1298]), .B(DB[1283]), .Z(n1530) );
  AND U5117 ( .A(n682), .B(n1531), .Z(n1529) );
  XOR U5118 ( .A(n1532), .B(n1533), .Z(n1531) );
  XOR U5119 ( .A(DB[1283]), .B(DB[1268]), .Z(n1533) );
  AND U5120 ( .A(n686), .B(n1534), .Z(n1532) );
  XOR U5121 ( .A(n1535), .B(n1536), .Z(n1534) );
  XOR U5122 ( .A(DB[1268]), .B(DB[1253]), .Z(n1536) );
  AND U5123 ( .A(n690), .B(n1537), .Z(n1535) );
  XOR U5124 ( .A(n1538), .B(n1539), .Z(n1537) );
  XOR U5125 ( .A(DB[1253]), .B(DB[1238]), .Z(n1539) );
  AND U5126 ( .A(n694), .B(n1540), .Z(n1538) );
  XOR U5127 ( .A(n1541), .B(n1542), .Z(n1540) );
  XOR U5128 ( .A(DB[1238]), .B(DB[1223]), .Z(n1542) );
  AND U5129 ( .A(n698), .B(n1543), .Z(n1541) );
  XOR U5130 ( .A(n1544), .B(n1545), .Z(n1543) );
  XOR U5131 ( .A(DB[1223]), .B(DB[1208]), .Z(n1545) );
  AND U5132 ( .A(n702), .B(n1546), .Z(n1544) );
  XOR U5133 ( .A(n1547), .B(n1548), .Z(n1546) );
  XOR U5134 ( .A(DB[1208]), .B(DB[1193]), .Z(n1548) );
  AND U5135 ( .A(n706), .B(n1549), .Z(n1547) );
  XOR U5136 ( .A(n1550), .B(n1551), .Z(n1549) );
  XOR U5137 ( .A(DB[1193]), .B(DB[1178]), .Z(n1551) );
  AND U5138 ( .A(n710), .B(n1552), .Z(n1550) );
  XOR U5139 ( .A(n1553), .B(n1554), .Z(n1552) );
  XOR U5140 ( .A(DB[1178]), .B(DB[1163]), .Z(n1554) );
  AND U5141 ( .A(n714), .B(n1555), .Z(n1553) );
  XOR U5142 ( .A(n1556), .B(n1557), .Z(n1555) );
  XOR U5143 ( .A(DB[1163]), .B(DB[1148]), .Z(n1557) );
  AND U5144 ( .A(n718), .B(n1558), .Z(n1556) );
  XOR U5145 ( .A(n1559), .B(n1560), .Z(n1558) );
  XOR U5146 ( .A(DB[1148]), .B(DB[1133]), .Z(n1560) );
  AND U5147 ( .A(n722), .B(n1561), .Z(n1559) );
  XOR U5148 ( .A(n1562), .B(n1563), .Z(n1561) );
  XOR U5149 ( .A(DB[1133]), .B(DB[1118]), .Z(n1563) );
  AND U5150 ( .A(n726), .B(n1564), .Z(n1562) );
  XOR U5151 ( .A(n1565), .B(n1566), .Z(n1564) );
  XOR U5152 ( .A(DB[1118]), .B(DB[1103]), .Z(n1566) );
  AND U5153 ( .A(n730), .B(n1567), .Z(n1565) );
  XOR U5154 ( .A(n1568), .B(n1569), .Z(n1567) );
  XOR U5155 ( .A(DB[1103]), .B(DB[1088]), .Z(n1569) );
  AND U5156 ( .A(n734), .B(n1570), .Z(n1568) );
  XOR U5157 ( .A(n1571), .B(n1572), .Z(n1570) );
  XOR U5158 ( .A(DB[1088]), .B(DB[1073]), .Z(n1572) );
  AND U5159 ( .A(n738), .B(n1573), .Z(n1571) );
  XOR U5160 ( .A(n1574), .B(n1575), .Z(n1573) );
  XOR U5161 ( .A(DB[1073]), .B(DB[1058]), .Z(n1575) );
  AND U5162 ( .A(n742), .B(n1576), .Z(n1574) );
  XOR U5163 ( .A(n1577), .B(n1578), .Z(n1576) );
  XOR U5164 ( .A(DB[1058]), .B(DB[1043]), .Z(n1578) );
  AND U5165 ( .A(n746), .B(n1579), .Z(n1577) );
  XOR U5166 ( .A(n1580), .B(n1581), .Z(n1579) );
  XOR U5167 ( .A(DB[1043]), .B(DB[1028]), .Z(n1581) );
  AND U5168 ( .A(n750), .B(n1582), .Z(n1580) );
  XOR U5169 ( .A(n1583), .B(n1584), .Z(n1582) );
  XOR U5170 ( .A(DB[1028]), .B(DB[1013]), .Z(n1584) );
  AND U5171 ( .A(n754), .B(n1585), .Z(n1583) );
  XOR U5172 ( .A(n1586), .B(n1587), .Z(n1585) );
  XOR U5173 ( .A(DB[998]), .B(DB[1013]), .Z(n1587) );
  AND U5174 ( .A(n758), .B(n1588), .Z(n1586) );
  XOR U5175 ( .A(n1589), .B(n1590), .Z(n1588) );
  XOR U5176 ( .A(DB[998]), .B(DB[983]), .Z(n1590) );
  AND U5177 ( .A(n762), .B(n1591), .Z(n1589) );
  XOR U5178 ( .A(n1592), .B(n1593), .Z(n1591) );
  XOR U5179 ( .A(DB[983]), .B(DB[968]), .Z(n1593) );
  AND U5180 ( .A(n766), .B(n1594), .Z(n1592) );
  XOR U5181 ( .A(n1595), .B(n1596), .Z(n1594) );
  XOR U5182 ( .A(DB[968]), .B(DB[953]), .Z(n1596) );
  AND U5183 ( .A(n770), .B(n1597), .Z(n1595) );
  XOR U5184 ( .A(n1598), .B(n1599), .Z(n1597) );
  XOR U5185 ( .A(DB[953]), .B(DB[938]), .Z(n1599) );
  AND U5186 ( .A(n774), .B(n1600), .Z(n1598) );
  XOR U5187 ( .A(n1601), .B(n1602), .Z(n1600) );
  XOR U5188 ( .A(DB[938]), .B(DB[923]), .Z(n1602) );
  AND U5189 ( .A(n778), .B(n1603), .Z(n1601) );
  XOR U5190 ( .A(n1604), .B(n1605), .Z(n1603) );
  XOR U5191 ( .A(DB[923]), .B(DB[908]), .Z(n1605) );
  AND U5192 ( .A(n782), .B(n1606), .Z(n1604) );
  XOR U5193 ( .A(n1607), .B(n1608), .Z(n1606) );
  XOR U5194 ( .A(DB[908]), .B(DB[893]), .Z(n1608) );
  AND U5195 ( .A(n786), .B(n1609), .Z(n1607) );
  XOR U5196 ( .A(n1610), .B(n1611), .Z(n1609) );
  XOR U5197 ( .A(DB[893]), .B(DB[878]), .Z(n1611) );
  AND U5198 ( .A(n790), .B(n1612), .Z(n1610) );
  XOR U5199 ( .A(n1613), .B(n1614), .Z(n1612) );
  XOR U5200 ( .A(DB[878]), .B(DB[863]), .Z(n1614) );
  AND U5201 ( .A(n794), .B(n1615), .Z(n1613) );
  XOR U5202 ( .A(n1616), .B(n1617), .Z(n1615) );
  XOR U5203 ( .A(DB[863]), .B(DB[848]), .Z(n1617) );
  AND U5204 ( .A(n798), .B(n1618), .Z(n1616) );
  XOR U5205 ( .A(n1619), .B(n1620), .Z(n1618) );
  XOR U5206 ( .A(DB[848]), .B(DB[833]), .Z(n1620) );
  AND U5207 ( .A(n802), .B(n1621), .Z(n1619) );
  XOR U5208 ( .A(n1622), .B(n1623), .Z(n1621) );
  XOR U5209 ( .A(DB[833]), .B(DB[818]), .Z(n1623) );
  AND U5210 ( .A(n806), .B(n1624), .Z(n1622) );
  XOR U5211 ( .A(n1625), .B(n1626), .Z(n1624) );
  XOR U5212 ( .A(DB[818]), .B(DB[803]), .Z(n1626) );
  AND U5213 ( .A(n810), .B(n1627), .Z(n1625) );
  XOR U5214 ( .A(n1628), .B(n1629), .Z(n1627) );
  XOR U5215 ( .A(DB[803]), .B(DB[788]), .Z(n1629) );
  AND U5216 ( .A(n814), .B(n1630), .Z(n1628) );
  XOR U5217 ( .A(n1631), .B(n1632), .Z(n1630) );
  XOR U5218 ( .A(DB[788]), .B(DB[773]), .Z(n1632) );
  AND U5219 ( .A(n818), .B(n1633), .Z(n1631) );
  XOR U5220 ( .A(n1634), .B(n1635), .Z(n1633) );
  XOR U5221 ( .A(DB[773]), .B(DB[758]), .Z(n1635) );
  AND U5222 ( .A(n822), .B(n1636), .Z(n1634) );
  XOR U5223 ( .A(n1637), .B(n1638), .Z(n1636) );
  XOR U5224 ( .A(DB[758]), .B(DB[743]), .Z(n1638) );
  AND U5225 ( .A(n826), .B(n1639), .Z(n1637) );
  XOR U5226 ( .A(n1640), .B(n1641), .Z(n1639) );
  XOR U5227 ( .A(DB[743]), .B(DB[728]), .Z(n1641) );
  AND U5228 ( .A(n830), .B(n1642), .Z(n1640) );
  XOR U5229 ( .A(n1643), .B(n1644), .Z(n1642) );
  XOR U5230 ( .A(DB[728]), .B(DB[713]), .Z(n1644) );
  AND U5231 ( .A(n834), .B(n1645), .Z(n1643) );
  XOR U5232 ( .A(n1646), .B(n1647), .Z(n1645) );
  XOR U5233 ( .A(DB[713]), .B(DB[698]), .Z(n1647) );
  AND U5234 ( .A(n838), .B(n1648), .Z(n1646) );
  XOR U5235 ( .A(n1649), .B(n1650), .Z(n1648) );
  XOR U5236 ( .A(DB[698]), .B(DB[683]), .Z(n1650) );
  AND U5237 ( .A(n842), .B(n1651), .Z(n1649) );
  XOR U5238 ( .A(n1652), .B(n1653), .Z(n1651) );
  XOR U5239 ( .A(DB[683]), .B(DB[668]), .Z(n1653) );
  AND U5240 ( .A(n846), .B(n1654), .Z(n1652) );
  XOR U5241 ( .A(n1655), .B(n1656), .Z(n1654) );
  XOR U5242 ( .A(DB[668]), .B(DB[653]), .Z(n1656) );
  AND U5243 ( .A(n850), .B(n1657), .Z(n1655) );
  XOR U5244 ( .A(n1658), .B(n1659), .Z(n1657) );
  XOR U5245 ( .A(DB[653]), .B(DB[638]), .Z(n1659) );
  AND U5246 ( .A(n854), .B(n1660), .Z(n1658) );
  XOR U5247 ( .A(n1661), .B(n1662), .Z(n1660) );
  XOR U5248 ( .A(DB[638]), .B(DB[623]), .Z(n1662) );
  AND U5249 ( .A(n858), .B(n1663), .Z(n1661) );
  XOR U5250 ( .A(n1664), .B(n1665), .Z(n1663) );
  XOR U5251 ( .A(DB[623]), .B(DB[608]), .Z(n1665) );
  AND U5252 ( .A(n862), .B(n1666), .Z(n1664) );
  XOR U5253 ( .A(n1667), .B(n1668), .Z(n1666) );
  XOR U5254 ( .A(DB[608]), .B(DB[593]), .Z(n1668) );
  AND U5255 ( .A(n866), .B(n1669), .Z(n1667) );
  XOR U5256 ( .A(n1670), .B(n1671), .Z(n1669) );
  XOR U5257 ( .A(DB[593]), .B(DB[578]), .Z(n1671) );
  AND U5258 ( .A(n870), .B(n1672), .Z(n1670) );
  XOR U5259 ( .A(n1673), .B(n1674), .Z(n1672) );
  XOR U5260 ( .A(DB[578]), .B(DB[563]), .Z(n1674) );
  AND U5261 ( .A(n874), .B(n1675), .Z(n1673) );
  XOR U5262 ( .A(n1676), .B(n1677), .Z(n1675) );
  XOR U5263 ( .A(DB[563]), .B(DB[548]), .Z(n1677) );
  AND U5264 ( .A(n878), .B(n1678), .Z(n1676) );
  XOR U5265 ( .A(n1679), .B(n1680), .Z(n1678) );
  XOR U5266 ( .A(DB[548]), .B(DB[533]), .Z(n1680) );
  AND U5267 ( .A(n882), .B(n1681), .Z(n1679) );
  XOR U5268 ( .A(n1682), .B(n1683), .Z(n1681) );
  XOR U5269 ( .A(DB[533]), .B(DB[518]), .Z(n1683) );
  AND U5270 ( .A(n886), .B(n1684), .Z(n1682) );
  XOR U5271 ( .A(n1685), .B(n1686), .Z(n1684) );
  XOR U5272 ( .A(DB[518]), .B(DB[503]), .Z(n1686) );
  AND U5273 ( .A(n890), .B(n1687), .Z(n1685) );
  XOR U5274 ( .A(n1688), .B(n1689), .Z(n1687) );
  XOR U5275 ( .A(DB[503]), .B(DB[488]), .Z(n1689) );
  AND U5276 ( .A(n894), .B(n1690), .Z(n1688) );
  XOR U5277 ( .A(n1691), .B(n1692), .Z(n1690) );
  XOR U5278 ( .A(DB[488]), .B(DB[473]), .Z(n1692) );
  AND U5279 ( .A(n898), .B(n1693), .Z(n1691) );
  XOR U5280 ( .A(n1694), .B(n1695), .Z(n1693) );
  XOR U5281 ( .A(DB[473]), .B(DB[458]), .Z(n1695) );
  AND U5282 ( .A(n902), .B(n1696), .Z(n1694) );
  XOR U5283 ( .A(n1697), .B(n1698), .Z(n1696) );
  XOR U5284 ( .A(DB[458]), .B(DB[443]), .Z(n1698) );
  AND U5285 ( .A(n906), .B(n1699), .Z(n1697) );
  XOR U5286 ( .A(n1700), .B(n1701), .Z(n1699) );
  XOR U5287 ( .A(DB[443]), .B(DB[428]), .Z(n1701) );
  AND U5288 ( .A(n910), .B(n1702), .Z(n1700) );
  XOR U5289 ( .A(n1703), .B(n1704), .Z(n1702) );
  XOR U5290 ( .A(DB[428]), .B(DB[413]), .Z(n1704) );
  AND U5291 ( .A(n914), .B(n1705), .Z(n1703) );
  XOR U5292 ( .A(n1706), .B(n1707), .Z(n1705) );
  XOR U5293 ( .A(DB[413]), .B(DB[398]), .Z(n1707) );
  AND U5294 ( .A(n918), .B(n1708), .Z(n1706) );
  XOR U5295 ( .A(n1709), .B(n1710), .Z(n1708) );
  XOR U5296 ( .A(DB[398]), .B(DB[383]), .Z(n1710) );
  AND U5297 ( .A(n922), .B(n1711), .Z(n1709) );
  XOR U5298 ( .A(n1712), .B(n1713), .Z(n1711) );
  XOR U5299 ( .A(DB[383]), .B(DB[368]), .Z(n1713) );
  AND U5300 ( .A(n926), .B(n1714), .Z(n1712) );
  XOR U5301 ( .A(n1715), .B(n1716), .Z(n1714) );
  XOR U5302 ( .A(DB[368]), .B(DB[353]), .Z(n1716) );
  AND U5303 ( .A(n930), .B(n1717), .Z(n1715) );
  XOR U5304 ( .A(n1718), .B(n1719), .Z(n1717) );
  XOR U5305 ( .A(DB[353]), .B(DB[338]), .Z(n1719) );
  AND U5306 ( .A(n934), .B(n1720), .Z(n1718) );
  XOR U5307 ( .A(n1721), .B(n1722), .Z(n1720) );
  XOR U5308 ( .A(DB[338]), .B(DB[323]), .Z(n1722) );
  AND U5309 ( .A(n938), .B(n1723), .Z(n1721) );
  XOR U5310 ( .A(n1724), .B(n1725), .Z(n1723) );
  XOR U5311 ( .A(DB[323]), .B(DB[308]), .Z(n1725) );
  AND U5312 ( .A(n942), .B(n1726), .Z(n1724) );
  XOR U5313 ( .A(n1727), .B(n1728), .Z(n1726) );
  XOR U5314 ( .A(DB[308]), .B(DB[293]), .Z(n1728) );
  AND U5315 ( .A(n946), .B(n1729), .Z(n1727) );
  XOR U5316 ( .A(n1730), .B(n1731), .Z(n1729) );
  XOR U5317 ( .A(DB[293]), .B(DB[278]), .Z(n1731) );
  AND U5318 ( .A(n950), .B(n1732), .Z(n1730) );
  XOR U5319 ( .A(n1733), .B(n1734), .Z(n1732) );
  XOR U5320 ( .A(DB[278]), .B(DB[263]), .Z(n1734) );
  AND U5321 ( .A(n954), .B(n1735), .Z(n1733) );
  XOR U5322 ( .A(n1736), .B(n1737), .Z(n1735) );
  XOR U5323 ( .A(DB[263]), .B(DB[248]), .Z(n1737) );
  AND U5324 ( .A(n958), .B(n1738), .Z(n1736) );
  XOR U5325 ( .A(n1739), .B(n1740), .Z(n1738) );
  XOR U5326 ( .A(DB[248]), .B(DB[233]), .Z(n1740) );
  AND U5327 ( .A(n962), .B(n1741), .Z(n1739) );
  XOR U5328 ( .A(n1742), .B(n1743), .Z(n1741) );
  XOR U5329 ( .A(DB[233]), .B(DB[218]), .Z(n1743) );
  AND U5330 ( .A(n966), .B(n1744), .Z(n1742) );
  XOR U5331 ( .A(n1745), .B(n1746), .Z(n1744) );
  XOR U5332 ( .A(DB[218]), .B(DB[203]), .Z(n1746) );
  AND U5333 ( .A(n970), .B(n1747), .Z(n1745) );
  XOR U5334 ( .A(n1748), .B(n1749), .Z(n1747) );
  XOR U5335 ( .A(DB[203]), .B(DB[188]), .Z(n1749) );
  AND U5336 ( .A(n974), .B(n1750), .Z(n1748) );
  XOR U5337 ( .A(n1751), .B(n1752), .Z(n1750) );
  XOR U5338 ( .A(DB[188]), .B(DB[173]), .Z(n1752) );
  AND U5339 ( .A(n978), .B(n1753), .Z(n1751) );
  XOR U5340 ( .A(n1754), .B(n1755), .Z(n1753) );
  XOR U5341 ( .A(DB[173]), .B(DB[158]), .Z(n1755) );
  AND U5342 ( .A(n982), .B(n1756), .Z(n1754) );
  XOR U5343 ( .A(n1757), .B(n1758), .Z(n1756) );
  XOR U5344 ( .A(DB[158]), .B(DB[143]), .Z(n1758) );
  AND U5345 ( .A(n986), .B(n1759), .Z(n1757) );
  XOR U5346 ( .A(n1760), .B(n1761), .Z(n1759) );
  XOR U5347 ( .A(DB[143]), .B(DB[128]), .Z(n1761) );
  AND U5348 ( .A(n990), .B(n1762), .Z(n1760) );
  XOR U5349 ( .A(n1763), .B(n1764), .Z(n1762) );
  XOR U5350 ( .A(DB[128]), .B(DB[113]), .Z(n1764) );
  AND U5351 ( .A(n994), .B(n1765), .Z(n1763) );
  XOR U5352 ( .A(n1766), .B(n1767), .Z(n1765) );
  XOR U5353 ( .A(DB[98]), .B(DB[113]), .Z(n1767) );
  AND U5354 ( .A(n998), .B(n1768), .Z(n1766) );
  XOR U5355 ( .A(n1769), .B(n1770), .Z(n1768) );
  XOR U5356 ( .A(DB[98]), .B(DB[83]), .Z(n1770) );
  AND U5357 ( .A(n1002), .B(n1771), .Z(n1769) );
  XOR U5358 ( .A(n1772), .B(n1773), .Z(n1771) );
  XOR U5359 ( .A(DB[83]), .B(DB[68]), .Z(n1773) );
  AND U5360 ( .A(n1006), .B(n1774), .Z(n1772) );
  XOR U5361 ( .A(n1775), .B(n1776), .Z(n1774) );
  XOR U5362 ( .A(DB[68]), .B(DB[53]), .Z(n1776) );
  AND U5363 ( .A(n1010), .B(n1777), .Z(n1775) );
  XOR U5364 ( .A(n1778), .B(n1779), .Z(n1777) );
  XOR U5365 ( .A(DB[53]), .B(DB[38]), .Z(n1779) );
  AND U5366 ( .A(n1014), .B(n1780), .Z(n1778) );
  XOR U5367 ( .A(n1781), .B(n1782), .Z(n1780) );
  XOR U5368 ( .A(DB[38]), .B(DB[23]), .Z(n1782) );
  AND U5369 ( .A(n1018), .B(n1783), .Z(n1781) );
  XOR U5370 ( .A(DB[8]), .B(DB[23]), .Z(n1783) );
  XOR U5371 ( .A(DB[3832]), .B(n1784), .Z(min_val_out[7]) );
  AND U5372 ( .A(n2), .B(n1785), .Z(n1784) );
  XOR U5373 ( .A(n1786), .B(n1787), .Z(n1785) );
  XOR U5374 ( .A(DB[3832]), .B(DB[3817]), .Z(n1787) );
  AND U5375 ( .A(n6), .B(n1788), .Z(n1786) );
  XOR U5376 ( .A(n1789), .B(n1790), .Z(n1788) );
  XOR U5377 ( .A(DB[3817]), .B(DB[3802]), .Z(n1790) );
  AND U5378 ( .A(n10), .B(n1791), .Z(n1789) );
  XOR U5379 ( .A(n1792), .B(n1793), .Z(n1791) );
  XOR U5380 ( .A(DB[3802]), .B(DB[3787]), .Z(n1793) );
  AND U5381 ( .A(n14), .B(n1794), .Z(n1792) );
  XOR U5382 ( .A(n1795), .B(n1796), .Z(n1794) );
  XOR U5383 ( .A(DB[3787]), .B(DB[3772]), .Z(n1796) );
  AND U5384 ( .A(n18), .B(n1797), .Z(n1795) );
  XOR U5385 ( .A(n1798), .B(n1799), .Z(n1797) );
  XOR U5386 ( .A(DB[3772]), .B(DB[3757]), .Z(n1799) );
  AND U5387 ( .A(n22), .B(n1800), .Z(n1798) );
  XOR U5388 ( .A(n1801), .B(n1802), .Z(n1800) );
  XOR U5389 ( .A(DB[3757]), .B(DB[3742]), .Z(n1802) );
  AND U5390 ( .A(n26), .B(n1803), .Z(n1801) );
  XOR U5391 ( .A(n1804), .B(n1805), .Z(n1803) );
  XOR U5392 ( .A(DB[3742]), .B(DB[3727]), .Z(n1805) );
  AND U5393 ( .A(n30), .B(n1806), .Z(n1804) );
  XOR U5394 ( .A(n1807), .B(n1808), .Z(n1806) );
  XOR U5395 ( .A(DB[3727]), .B(DB[3712]), .Z(n1808) );
  AND U5396 ( .A(n34), .B(n1809), .Z(n1807) );
  XOR U5397 ( .A(n1810), .B(n1811), .Z(n1809) );
  XOR U5398 ( .A(DB[3712]), .B(DB[3697]), .Z(n1811) );
  AND U5399 ( .A(n38), .B(n1812), .Z(n1810) );
  XOR U5400 ( .A(n1813), .B(n1814), .Z(n1812) );
  XOR U5401 ( .A(DB[3697]), .B(DB[3682]), .Z(n1814) );
  AND U5402 ( .A(n42), .B(n1815), .Z(n1813) );
  XOR U5403 ( .A(n1816), .B(n1817), .Z(n1815) );
  XOR U5404 ( .A(DB[3682]), .B(DB[3667]), .Z(n1817) );
  AND U5405 ( .A(n46), .B(n1818), .Z(n1816) );
  XOR U5406 ( .A(n1819), .B(n1820), .Z(n1818) );
  XOR U5407 ( .A(DB[3667]), .B(DB[3652]), .Z(n1820) );
  AND U5408 ( .A(n50), .B(n1821), .Z(n1819) );
  XOR U5409 ( .A(n1822), .B(n1823), .Z(n1821) );
  XOR U5410 ( .A(DB[3652]), .B(DB[3637]), .Z(n1823) );
  AND U5411 ( .A(n54), .B(n1824), .Z(n1822) );
  XOR U5412 ( .A(n1825), .B(n1826), .Z(n1824) );
  XOR U5413 ( .A(DB[3637]), .B(DB[3622]), .Z(n1826) );
  AND U5414 ( .A(n58), .B(n1827), .Z(n1825) );
  XOR U5415 ( .A(n1828), .B(n1829), .Z(n1827) );
  XOR U5416 ( .A(DB[3622]), .B(DB[3607]), .Z(n1829) );
  AND U5417 ( .A(n62), .B(n1830), .Z(n1828) );
  XOR U5418 ( .A(n1831), .B(n1832), .Z(n1830) );
  XOR U5419 ( .A(DB[3607]), .B(DB[3592]), .Z(n1832) );
  AND U5420 ( .A(n66), .B(n1833), .Z(n1831) );
  XOR U5421 ( .A(n1834), .B(n1835), .Z(n1833) );
  XOR U5422 ( .A(DB[3592]), .B(DB[3577]), .Z(n1835) );
  AND U5423 ( .A(n70), .B(n1836), .Z(n1834) );
  XOR U5424 ( .A(n1837), .B(n1838), .Z(n1836) );
  XOR U5425 ( .A(DB[3577]), .B(DB[3562]), .Z(n1838) );
  AND U5426 ( .A(n74), .B(n1839), .Z(n1837) );
  XOR U5427 ( .A(n1840), .B(n1841), .Z(n1839) );
  XOR U5428 ( .A(DB[3562]), .B(DB[3547]), .Z(n1841) );
  AND U5429 ( .A(n78), .B(n1842), .Z(n1840) );
  XOR U5430 ( .A(n1843), .B(n1844), .Z(n1842) );
  XOR U5431 ( .A(DB[3547]), .B(DB[3532]), .Z(n1844) );
  AND U5432 ( .A(n82), .B(n1845), .Z(n1843) );
  XOR U5433 ( .A(n1846), .B(n1847), .Z(n1845) );
  XOR U5434 ( .A(DB[3532]), .B(DB[3517]), .Z(n1847) );
  AND U5435 ( .A(n86), .B(n1848), .Z(n1846) );
  XOR U5436 ( .A(n1849), .B(n1850), .Z(n1848) );
  XOR U5437 ( .A(DB[3517]), .B(DB[3502]), .Z(n1850) );
  AND U5438 ( .A(n90), .B(n1851), .Z(n1849) );
  XOR U5439 ( .A(n1852), .B(n1853), .Z(n1851) );
  XOR U5440 ( .A(DB[3502]), .B(DB[3487]), .Z(n1853) );
  AND U5441 ( .A(n94), .B(n1854), .Z(n1852) );
  XOR U5442 ( .A(n1855), .B(n1856), .Z(n1854) );
  XOR U5443 ( .A(DB[3487]), .B(DB[3472]), .Z(n1856) );
  AND U5444 ( .A(n98), .B(n1857), .Z(n1855) );
  XOR U5445 ( .A(n1858), .B(n1859), .Z(n1857) );
  XOR U5446 ( .A(DB[3472]), .B(DB[3457]), .Z(n1859) );
  AND U5447 ( .A(n102), .B(n1860), .Z(n1858) );
  XOR U5448 ( .A(n1861), .B(n1862), .Z(n1860) );
  XOR U5449 ( .A(DB[3457]), .B(DB[3442]), .Z(n1862) );
  AND U5450 ( .A(n106), .B(n1863), .Z(n1861) );
  XOR U5451 ( .A(n1864), .B(n1865), .Z(n1863) );
  XOR U5452 ( .A(DB[3442]), .B(DB[3427]), .Z(n1865) );
  AND U5453 ( .A(n110), .B(n1866), .Z(n1864) );
  XOR U5454 ( .A(n1867), .B(n1868), .Z(n1866) );
  XOR U5455 ( .A(DB[3427]), .B(DB[3412]), .Z(n1868) );
  AND U5456 ( .A(n114), .B(n1869), .Z(n1867) );
  XOR U5457 ( .A(n1870), .B(n1871), .Z(n1869) );
  XOR U5458 ( .A(DB[3412]), .B(DB[3397]), .Z(n1871) );
  AND U5459 ( .A(n118), .B(n1872), .Z(n1870) );
  XOR U5460 ( .A(n1873), .B(n1874), .Z(n1872) );
  XOR U5461 ( .A(DB[3397]), .B(DB[3382]), .Z(n1874) );
  AND U5462 ( .A(n122), .B(n1875), .Z(n1873) );
  XOR U5463 ( .A(n1876), .B(n1877), .Z(n1875) );
  XOR U5464 ( .A(DB[3382]), .B(DB[3367]), .Z(n1877) );
  AND U5465 ( .A(n126), .B(n1878), .Z(n1876) );
  XOR U5466 ( .A(n1879), .B(n1880), .Z(n1878) );
  XOR U5467 ( .A(DB[3367]), .B(DB[3352]), .Z(n1880) );
  AND U5468 ( .A(n130), .B(n1881), .Z(n1879) );
  XOR U5469 ( .A(n1882), .B(n1883), .Z(n1881) );
  XOR U5470 ( .A(DB[3352]), .B(DB[3337]), .Z(n1883) );
  AND U5471 ( .A(n134), .B(n1884), .Z(n1882) );
  XOR U5472 ( .A(n1885), .B(n1886), .Z(n1884) );
  XOR U5473 ( .A(DB[3337]), .B(DB[3322]), .Z(n1886) );
  AND U5474 ( .A(n138), .B(n1887), .Z(n1885) );
  XOR U5475 ( .A(n1888), .B(n1889), .Z(n1887) );
  XOR U5476 ( .A(DB[3322]), .B(DB[3307]), .Z(n1889) );
  AND U5477 ( .A(n142), .B(n1890), .Z(n1888) );
  XOR U5478 ( .A(n1891), .B(n1892), .Z(n1890) );
  XOR U5479 ( .A(DB[3307]), .B(DB[3292]), .Z(n1892) );
  AND U5480 ( .A(n146), .B(n1893), .Z(n1891) );
  XOR U5481 ( .A(n1894), .B(n1895), .Z(n1893) );
  XOR U5482 ( .A(DB[3292]), .B(DB[3277]), .Z(n1895) );
  AND U5483 ( .A(n150), .B(n1896), .Z(n1894) );
  XOR U5484 ( .A(n1897), .B(n1898), .Z(n1896) );
  XOR U5485 ( .A(DB[3277]), .B(DB[3262]), .Z(n1898) );
  AND U5486 ( .A(n154), .B(n1899), .Z(n1897) );
  XOR U5487 ( .A(n1900), .B(n1901), .Z(n1899) );
  XOR U5488 ( .A(DB[3262]), .B(DB[3247]), .Z(n1901) );
  AND U5489 ( .A(n158), .B(n1902), .Z(n1900) );
  XOR U5490 ( .A(n1903), .B(n1904), .Z(n1902) );
  XOR U5491 ( .A(DB[3247]), .B(DB[3232]), .Z(n1904) );
  AND U5492 ( .A(n162), .B(n1905), .Z(n1903) );
  XOR U5493 ( .A(n1906), .B(n1907), .Z(n1905) );
  XOR U5494 ( .A(DB[3232]), .B(DB[3217]), .Z(n1907) );
  AND U5495 ( .A(n166), .B(n1908), .Z(n1906) );
  XOR U5496 ( .A(n1909), .B(n1910), .Z(n1908) );
  XOR U5497 ( .A(DB[3217]), .B(DB[3202]), .Z(n1910) );
  AND U5498 ( .A(n170), .B(n1911), .Z(n1909) );
  XOR U5499 ( .A(n1912), .B(n1913), .Z(n1911) );
  XOR U5500 ( .A(DB[3202]), .B(DB[3187]), .Z(n1913) );
  AND U5501 ( .A(n174), .B(n1914), .Z(n1912) );
  XOR U5502 ( .A(n1915), .B(n1916), .Z(n1914) );
  XOR U5503 ( .A(DB[3187]), .B(DB[3172]), .Z(n1916) );
  AND U5504 ( .A(n178), .B(n1917), .Z(n1915) );
  XOR U5505 ( .A(n1918), .B(n1919), .Z(n1917) );
  XOR U5506 ( .A(DB[3172]), .B(DB[3157]), .Z(n1919) );
  AND U5507 ( .A(n182), .B(n1920), .Z(n1918) );
  XOR U5508 ( .A(n1921), .B(n1922), .Z(n1920) );
  XOR U5509 ( .A(DB[3157]), .B(DB[3142]), .Z(n1922) );
  AND U5510 ( .A(n186), .B(n1923), .Z(n1921) );
  XOR U5511 ( .A(n1924), .B(n1925), .Z(n1923) );
  XOR U5512 ( .A(DB[3142]), .B(DB[3127]), .Z(n1925) );
  AND U5513 ( .A(n190), .B(n1926), .Z(n1924) );
  XOR U5514 ( .A(n1927), .B(n1928), .Z(n1926) );
  XOR U5515 ( .A(DB[3127]), .B(DB[3112]), .Z(n1928) );
  AND U5516 ( .A(n194), .B(n1929), .Z(n1927) );
  XOR U5517 ( .A(n1930), .B(n1931), .Z(n1929) );
  XOR U5518 ( .A(DB[3112]), .B(DB[3097]), .Z(n1931) );
  AND U5519 ( .A(n198), .B(n1932), .Z(n1930) );
  XOR U5520 ( .A(n1933), .B(n1934), .Z(n1932) );
  XOR U5521 ( .A(DB[3097]), .B(DB[3082]), .Z(n1934) );
  AND U5522 ( .A(n202), .B(n1935), .Z(n1933) );
  XOR U5523 ( .A(n1936), .B(n1937), .Z(n1935) );
  XOR U5524 ( .A(DB[3082]), .B(DB[3067]), .Z(n1937) );
  AND U5525 ( .A(n206), .B(n1938), .Z(n1936) );
  XOR U5526 ( .A(n1939), .B(n1940), .Z(n1938) );
  XOR U5527 ( .A(DB[3067]), .B(DB[3052]), .Z(n1940) );
  AND U5528 ( .A(n210), .B(n1941), .Z(n1939) );
  XOR U5529 ( .A(n1942), .B(n1943), .Z(n1941) );
  XOR U5530 ( .A(DB[3052]), .B(DB[3037]), .Z(n1943) );
  AND U5531 ( .A(n214), .B(n1944), .Z(n1942) );
  XOR U5532 ( .A(n1945), .B(n1946), .Z(n1944) );
  XOR U5533 ( .A(DB[3037]), .B(DB[3022]), .Z(n1946) );
  AND U5534 ( .A(n218), .B(n1947), .Z(n1945) );
  XOR U5535 ( .A(n1948), .B(n1949), .Z(n1947) );
  XOR U5536 ( .A(DB[3022]), .B(DB[3007]), .Z(n1949) );
  AND U5537 ( .A(n222), .B(n1950), .Z(n1948) );
  XOR U5538 ( .A(n1951), .B(n1952), .Z(n1950) );
  XOR U5539 ( .A(DB[3007]), .B(DB[2992]), .Z(n1952) );
  AND U5540 ( .A(n226), .B(n1953), .Z(n1951) );
  XOR U5541 ( .A(n1954), .B(n1955), .Z(n1953) );
  XOR U5542 ( .A(DB[2992]), .B(DB[2977]), .Z(n1955) );
  AND U5543 ( .A(n230), .B(n1956), .Z(n1954) );
  XOR U5544 ( .A(n1957), .B(n1958), .Z(n1956) );
  XOR U5545 ( .A(DB[2977]), .B(DB[2962]), .Z(n1958) );
  AND U5546 ( .A(n234), .B(n1959), .Z(n1957) );
  XOR U5547 ( .A(n1960), .B(n1961), .Z(n1959) );
  XOR U5548 ( .A(DB[2962]), .B(DB[2947]), .Z(n1961) );
  AND U5549 ( .A(n238), .B(n1962), .Z(n1960) );
  XOR U5550 ( .A(n1963), .B(n1964), .Z(n1962) );
  XOR U5551 ( .A(DB[2947]), .B(DB[2932]), .Z(n1964) );
  AND U5552 ( .A(n242), .B(n1965), .Z(n1963) );
  XOR U5553 ( .A(n1966), .B(n1967), .Z(n1965) );
  XOR U5554 ( .A(DB[2932]), .B(DB[2917]), .Z(n1967) );
  AND U5555 ( .A(n246), .B(n1968), .Z(n1966) );
  XOR U5556 ( .A(n1969), .B(n1970), .Z(n1968) );
  XOR U5557 ( .A(DB[2917]), .B(DB[2902]), .Z(n1970) );
  AND U5558 ( .A(n250), .B(n1971), .Z(n1969) );
  XOR U5559 ( .A(n1972), .B(n1973), .Z(n1971) );
  XOR U5560 ( .A(DB[2902]), .B(DB[2887]), .Z(n1973) );
  AND U5561 ( .A(n254), .B(n1974), .Z(n1972) );
  XOR U5562 ( .A(n1975), .B(n1976), .Z(n1974) );
  XOR U5563 ( .A(DB[2887]), .B(DB[2872]), .Z(n1976) );
  AND U5564 ( .A(n258), .B(n1977), .Z(n1975) );
  XOR U5565 ( .A(n1978), .B(n1979), .Z(n1977) );
  XOR U5566 ( .A(DB[2872]), .B(DB[2857]), .Z(n1979) );
  AND U5567 ( .A(n262), .B(n1980), .Z(n1978) );
  XOR U5568 ( .A(n1981), .B(n1982), .Z(n1980) );
  XOR U5569 ( .A(DB[2857]), .B(DB[2842]), .Z(n1982) );
  AND U5570 ( .A(n266), .B(n1983), .Z(n1981) );
  XOR U5571 ( .A(n1984), .B(n1985), .Z(n1983) );
  XOR U5572 ( .A(DB[2842]), .B(DB[2827]), .Z(n1985) );
  AND U5573 ( .A(n270), .B(n1986), .Z(n1984) );
  XOR U5574 ( .A(n1987), .B(n1988), .Z(n1986) );
  XOR U5575 ( .A(DB[2827]), .B(DB[2812]), .Z(n1988) );
  AND U5576 ( .A(n274), .B(n1989), .Z(n1987) );
  XOR U5577 ( .A(n1990), .B(n1991), .Z(n1989) );
  XOR U5578 ( .A(DB[2812]), .B(DB[2797]), .Z(n1991) );
  AND U5579 ( .A(n278), .B(n1992), .Z(n1990) );
  XOR U5580 ( .A(n1993), .B(n1994), .Z(n1992) );
  XOR U5581 ( .A(DB[2797]), .B(DB[2782]), .Z(n1994) );
  AND U5582 ( .A(n282), .B(n1995), .Z(n1993) );
  XOR U5583 ( .A(n1996), .B(n1997), .Z(n1995) );
  XOR U5584 ( .A(DB[2782]), .B(DB[2767]), .Z(n1997) );
  AND U5585 ( .A(n286), .B(n1998), .Z(n1996) );
  XOR U5586 ( .A(n1999), .B(n2000), .Z(n1998) );
  XOR U5587 ( .A(DB[2767]), .B(DB[2752]), .Z(n2000) );
  AND U5588 ( .A(n290), .B(n2001), .Z(n1999) );
  XOR U5589 ( .A(n2002), .B(n2003), .Z(n2001) );
  XOR U5590 ( .A(DB[2752]), .B(DB[2737]), .Z(n2003) );
  AND U5591 ( .A(n294), .B(n2004), .Z(n2002) );
  XOR U5592 ( .A(n2005), .B(n2006), .Z(n2004) );
  XOR U5593 ( .A(DB[2737]), .B(DB[2722]), .Z(n2006) );
  AND U5594 ( .A(n298), .B(n2007), .Z(n2005) );
  XOR U5595 ( .A(n2008), .B(n2009), .Z(n2007) );
  XOR U5596 ( .A(DB[2722]), .B(DB[2707]), .Z(n2009) );
  AND U5597 ( .A(n302), .B(n2010), .Z(n2008) );
  XOR U5598 ( .A(n2011), .B(n2012), .Z(n2010) );
  XOR U5599 ( .A(DB[2707]), .B(DB[2692]), .Z(n2012) );
  AND U5600 ( .A(n306), .B(n2013), .Z(n2011) );
  XOR U5601 ( .A(n2014), .B(n2015), .Z(n2013) );
  XOR U5602 ( .A(DB[2692]), .B(DB[2677]), .Z(n2015) );
  AND U5603 ( .A(n310), .B(n2016), .Z(n2014) );
  XOR U5604 ( .A(n2017), .B(n2018), .Z(n2016) );
  XOR U5605 ( .A(DB[2677]), .B(DB[2662]), .Z(n2018) );
  AND U5606 ( .A(n314), .B(n2019), .Z(n2017) );
  XOR U5607 ( .A(n2020), .B(n2021), .Z(n2019) );
  XOR U5608 ( .A(DB[2662]), .B(DB[2647]), .Z(n2021) );
  AND U5609 ( .A(n318), .B(n2022), .Z(n2020) );
  XOR U5610 ( .A(n2023), .B(n2024), .Z(n2022) );
  XOR U5611 ( .A(DB[2647]), .B(DB[2632]), .Z(n2024) );
  AND U5612 ( .A(n322), .B(n2025), .Z(n2023) );
  XOR U5613 ( .A(n2026), .B(n2027), .Z(n2025) );
  XOR U5614 ( .A(DB[2632]), .B(DB[2617]), .Z(n2027) );
  AND U5615 ( .A(n326), .B(n2028), .Z(n2026) );
  XOR U5616 ( .A(n2029), .B(n2030), .Z(n2028) );
  XOR U5617 ( .A(DB[2617]), .B(DB[2602]), .Z(n2030) );
  AND U5618 ( .A(n330), .B(n2031), .Z(n2029) );
  XOR U5619 ( .A(n2032), .B(n2033), .Z(n2031) );
  XOR U5620 ( .A(DB[2602]), .B(DB[2587]), .Z(n2033) );
  AND U5621 ( .A(n334), .B(n2034), .Z(n2032) );
  XOR U5622 ( .A(n2035), .B(n2036), .Z(n2034) );
  XOR U5623 ( .A(DB[2587]), .B(DB[2572]), .Z(n2036) );
  AND U5624 ( .A(n338), .B(n2037), .Z(n2035) );
  XOR U5625 ( .A(n2038), .B(n2039), .Z(n2037) );
  XOR U5626 ( .A(DB[2572]), .B(DB[2557]), .Z(n2039) );
  AND U5627 ( .A(n342), .B(n2040), .Z(n2038) );
  XOR U5628 ( .A(n2041), .B(n2042), .Z(n2040) );
  XOR U5629 ( .A(DB[2557]), .B(DB[2542]), .Z(n2042) );
  AND U5630 ( .A(n346), .B(n2043), .Z(n2041) );
  XOR U5631 ( .A(n2044), .B(n2045), .Z(n2043) );
  XOR U5632 ( .A(DB[2542]), .B(DB[2527]), .Z(n2045) );
  AND U5633 ( .A(n350), .B(n2046), .Z(n2044) );
  XOR U5634 ( .A(n2047), .B(n2048), .Z(n2046) );
  XOR U5635 ( .A(DB[2527]), .B(DB[2512]), .Z(n2048) );
  AND U5636 ( .A(n354), .B(n2049), .Z(n2047) );
  XOR U5637 ( .A(n2050), .B(n2051), .Z(n2049) );
  XOR U5638 ( .A(DB[2512]), .B(DB[2497]), .Z(n2051) );
  AND U5639 ( .A(n358), .B(n2052), .Z(n2050) );
  XOR U5640 ( .A(n2053), .B(n2054), .Z(n2052) );
  XOR U5641 ( .A(DB[2497]), .B(DB[2482]), .Z(n2054) );
  AND U5642 ( .A(n362), .B(n2055), .Z(n2053) );
  XOR U5643 ( .A(n2056), .B(n2057), .Z(n2055) );
  XOR U5644 ( .A(DB[2482]), .B(DB[2467]), .Z(n2057) );
  AND U5645 ( .A(n366), .B(n2058), .Z(n2056) );
  XOR U5646 ( .A(n2059), .B(n2060), .Z(n2058) );
  XOR U5647 ( .A(DB[2467]), .B(DB[2452]), .Z(n2060) );
  AND U5648 ( .A(n370), .B(n2061), .Z(n2059) );
  XOR U5649 ( .A(n2062), .B(n2063), .Z(n2061) );
  XOR U5650 ( .A(DB[2452]), .B(DB[2437]), .Z(n2063) );
  AND U5651 ( .A(n374), .B(n2064), .Z(n2062) );
  XOR U5652 ( .A(n2065), .B(n2066), .Z(n2064) );
  XOR U5653 ( .A(DB[2437]), .B(DB[2422]), .Z(n2066) );
  AND U5654 ( .A(n378), .B(n2067), .Z(n2065) );
  XOR U5655 ( .A(n2068), .B(n2069), .Z(n2067) );
  XOR U5656 ( .A(DB[2422]), .B(DB[2407]), .Z(n2069) );
  AND U5657 ( .A(n382), .B(n2070), .Z(n2068) );
  XOR U5658 ( .A(n2071), .B(n2072), .Z(n2070) );
  XOR U5659 ( .A(DB[2407]), .B(DB[2392]), .Z(n2072) );
  AND U5660 ( .A(n386), .B(n2073), .Z(n2071) );
  XOR U5661 ( .A(n2074), .B(n2075), .Z(n2073) );
  XOR U5662 ( .A(DB[2392]), .B(DB[2377]), .Z(n2075) );
  AND U5663 ( .A(n390), .B(n2076), .Z(n2074) );
  XOR U5664 ( .A(n2077), .B(n2078), .Z(n2076) );
  XOR U5665 ( .A(DB[2377]), .B(DB[2362]), .Z(n2078) );
  AND U5666 ( .A(n394), .B(n2079), .Z(n2077) );
  XOR U5667 ( .A(n2080), .B(n2081), .Z(n2079) );
  XOR U5668 ( .A(DB[2362]), .B(DB[2347]), .Z(n2081) );
  AND U5669 ( .A(n398), .B(n2082), .Z(n2080) );
  XOR U5670 ( .A(n2083), .B(n2084), .Z(n2082) );
  XOR U5671 ( .A(DB[2347]), .B(DB[2332]), .Z(n2084) );
  AND U5672 ( .A(n402), .B(n2085), .Z(n2083) );
  XOR U5673 ( .A(n2086), .B(n2087), .Z(n2085) );
  XOR U5674 ( .A(DB[2332]), .B(DB[2317]), .Z(n2087) );
  AND U5675 ( .A(n406), .B(n2088), .Z(n2086) );
  XOR U5676 ( .A(n2089), .B(n2090), .Z(n2088) );
  XOR U5677 ( .A(DB[2317]), .B(DB[2302]), .Z(n2090) );
  AND U5678 ( .A(n410), .B(n2091), .Z(n2089) );
  XOR U5679 ( .A(n2092), .B(n2093), .Z(n2091) );
  XOR U5680 ( .A(DB[2302]), .B(DB[2287]), .Z(n2093) );
  AND U5681 ( .A(n414), .B(n2094), .Z(n2092) );
  XOR U5682 ( .A(n2095), .B(n2096), .Z(n2094) );
  XOR U5683 ( .A(DB[2287]), .B(DB[2272]), .Z(n2096) );
  AND U5684 ( .A(n418), .B(n2097), .Z(n2095) );
  XOR U5685 ( .A(n2098), .B(n2099), .Z(n2097) );
  XOR U5686 ( .A(DB[2272]), .B(DB[2257]), .Z(n2099) );
  AND U5687 ( .A(n422), .B(n2100), .Z(n2098) );
  XOR U5688 ( .A(n2101), .B(n2102), .Z(n2100) );
  XOR U5689 ( .A(DB[2257]), .B(DB[2242]), .Z(n2102) );
  AND U5690 ( .A(n426), .B(n2103), .Z(n2101) );
  XOR U5691 ( .A(n2104), .B(n2105), .Z(n2103) );
  XOR U5692 ( .A(DB[2242]), .B(DB[2227]), .Z(n2105) );
  AND U5693 ( .A(n430), .B(n2106), .Z(n2104) );
  XOR U5694 ( .A(n2107), .B(n2108), .Z(n2106) );
  XOR U5695 ( .A(DB[2227]), .B(DB[2212]), .Z(n2108) );
  AND U5696 ( .A(n434), .B(n2109), .Z(n2107) );
  XOR U5697 ( .A(n2110), .B(n2111), .Z(n2109) );
  XOR U5698 ( .A(DB[2212]), .B(DB[2197]), .Z(n2111) );
  AND U5699 ( .A(n438), .B(n2112), .Z(n2110) );
  XOR U5700 ( .A(n2113), .B(n2114), .Z(n2112) );
  XOR U5701 ( .A(DB[2197]), .B(DB[2182]), .Z(n2114) );
  AND U5702 ( .A(n442), .B(n2115), .Z(n2113) );
  XOR U5703 ( .A(n2116), .B(n2117), .Z(n2115) );
  XOR U5704 ( .A(DB[2182]), .B(DB[2167]), .Z(n2117) );
  AND U5705 ( .A(n446), .B(n2118), .Z(n2116) );
  XOR U5706 ( .A(n2119), .B(n2120), .Z(n2118) );
  XOR U5707 ( .A(DB[2167]), .B(DB[2152]), .Z(n2120) );
  AND U5708 ( .A(n450), .B(n2121), .Z(n2119) );
  XOR U5709 ( .A(n2122), .B(n2123), .Z(n2121) );
  XOR U5710 ( .A(DB[2152]), .B(DB[2137]), .Z(n2123) );
  AND U5711 ( .A(n454), .B(n2124), .Z(n2122) );
  XOR U5712 ( .A(n2125), .B(n2126), .Z(n2124) );
  XOR U5713 ( .A(DB[2137]), .B(DB[2122]), .Z(n2126) );
  AND U5714 ( .A(n458), .B(n2127), .Z(n2125) );
  XOR U5715 ( .A(n2128), .B(n2129), .Z(n2127) );
  XOR U5716 ( .A(DB[2122]), .B(DB[2107]), .Z(n2129) );
  AND U5717 ( .A(n462), .B(n2130), .Z(n2128) );
  XOR U5718 ( .A(n2131), .B(n2132), .Z(n2130) );
  XOR U5719 ( .A(DB[2107]), .B(DB[2092]), .Z(n2132) );
  AND U5720 ( .A(n466), .B(n2133), .Z(n2131) );
  XOR U5721 ( .A(n2134), .B(n2135), .Z(n2133) );
  XOR U5722 ( .A(DB[2092]), .B(DB[2077]), .Z(n2135) );
  AND U5723 ( .A(n470), .B(n2136), .Z(n2134) );
  XOR U5724 ( .A(n2137), .B(n2138), .Z(n2136) );
  XOR U5725 ( .A(DB[2077]), .B(DB[2062]), .Z(n2138) );
  AND U5726 ( .A(n474), .B(n2139), .Z(n2137) );
  XOR U5727 ( .A(n2140), .B(n2141), .Z(n2139) );
  XOR U5728 ( .A(DB[2062]), .B(DB[2047]), .Z(n2141) );
  AND U5729 ( .A(n478), .B(n2142), .Z(n2140) );
  XOR U5730 ( .A(n2143), .B(n2144), .Z(n2142) );
  XOR U5731 ( .A(DB[2047]), .B(DB[2032]), .Z(n2144) );
  AND U5732 ( .A(n482), .B(n2145), .Z(n2143) );
  XOR U5733 ( .A(n2146), .B(n2147), .Z(n2145) );
  XOR U5734 ( .A(DB[2032]), .B(DB[2017]), .Z(n2147) );
  AND U5735 ( .A(n486), .B(n2148), .Z(n2146) );
  XOR U5736 ( .A(n2149), .B(n2150), .Z(n2148) );
  XOR U5737 ( .A(DB[2017]), .B(DB[2002]), .Z(n2150) );
  AND U5738 ( .A(n490), .B(n2151), .Z(n2149) );
  XOR U5739 ( .A(n2152), .B(n2153), .Z(n2151) );
  XOR U5740 ( .A(DB[2002]), .B(DB[1987]), .Z(n2153) );
  AND U5741 ( .A(n494), .B(n2154), .Z(n2152) );
  XOR U5742 ( .A(n2155), .B(n2156), .Z(n2154) );
  XOR U5743 ( .A(DB[1987]), .B(DB[1972]), .Z(n2156) );
  AND U5744 ( .A(n498), .B(n2157), .Z(n2155) );
  XOR U5745 ( .A(n2158), .B(n2159), .Z(n2157) );
  XOR U5746 ( .A(DB[1972]), .B(DB[1957]), .Z(n2159) );
  AND U5747 ( .A(n502), .B(n2160), .Z(n2158) );
  XOR U5748 ( .A(n2161), .B(n2162), .Z(n2160) );
  XOR U5749 ( .A(DB[1957]), .B(DB[1942]), .Z(n2162) );
  AND U5750 ( .A(n506), .B(n2163), .Z(n2161) );
  XOR U5751 ( .A(n2164), .B(n2165), .Z(n2163) );
  XOR U5752 ( .A(DB[1942]), .B(DB[1927]), .Z(n2165) );
  AND U5753 ( .A(n510), .B(n2166), .Z(n2164) );
  XOR U5754 ( .A(n2167), .B(n2168), .Z(n2166) );
  XOR U5755 ( .A(DB[1927]), .B(DB[1912]), .Z(n2168) );
  AND U5756 ( .A(n514), .B(n2169), .Z(n2167) );
  XOR U5757 ( .A(n2170), .B(n2171), .Z(n2169) );
  XOR U5758 ( .A(DB[1912]), .B(DB[1897]), .Z(n2171) );
  AND U5759 ( .A(n518), .B(n2172), .Z(n2170) );
  XOR U5760 ( .A(n2173), .B(n2174), .Z(n2172) );
  XOR U5761 ( .A(DB[1897]), .B(DB[1882]), .Z(n2174) );
  AND U5762 ( .A(n522), .B(n2175), .Z(n2173) );
  XOR U5763 ( .A(n2176), .B(n2177), .Z(n2175) );
  XOR U5764 ( .A(DB[1882]), .B(DB[1867]), .Z(n2177) );
  AND U5765 ( .A(n526), .B(n2178), .Z(n2176) );
  XOR U5766 ( .A(n2179), .B(n2180), .Z(n2178) );
  XOR U5767 ( .A(DB[1867]), .B(DB[1852]), .Z(n2180) );
  AND U5768 ( .A(n530), .B(n2181), .Z(n2179) );
  XOR U5769 ( .A(n2182), .B(n2183), .Z(n2181) );
  XOR U5770 ( .A(DB[1852]), .B(DB[1837]), .Z(n2183) );
  AND U5771 ( .A(n534), .B(n2184), .Z(n2182) );
  XOR U5772 ( .A(n2185), .B(n2186), .Z(n2184) );
  XOR U5773 ( .A(DB[1837]), .B(DB[1822]), .Z(n2186) );
  AND U5774 ( .A(n538), .B(n2187), .Z(n2185) );
  XOR U5775 ( .A(n2188), .B(n2189), .Z(n2187) );
  XOR U5776 ( .A(DB[1822]), .B(DB[1807]), .Z(n2189) );
  AND U5777 ( .A(n542), .B(n2190), .Z(n2188) );
  XOR U5778 ( .A(n2191), .B(n2192), .Z(n2190) );
  XOR U5779 ( .A(DB[1807]), .B(DB[1792]), .Z(n2192) );
  AND U5780 ( .A(n546), .B(n2193), .Z(n2191) );
  XOR U5781 ( .A(n2194), .B(n2195), .Z(n2193) );
  XOR U5782 ( .A(DB[1792]), .B(DB[1777]), .Z(n2195) );
  AND U5783 ( .A(n550), .B(n2196), .Z(n2194) );
  XOR U5784 ( .A(n2197), .B(n2198), .Z(n2196) );
  XOR U5785 ( .A(DB[1777]), .B(DB[1762]), .Z(n2198) );
  AND U5786 ( .A(n554), .B(n2199), .Z(n2197) );
  XOR U5787 ( .A(n2200), .B(n2201), .Z(n2199) );
  XOR U5788 ( .A(DB[1762]), .B(DB[1747]), .Z(n2201) );
  AND U5789 ( .A(n558), .B(n2202), .Z(n2200) );
  XOR U5790 ( .A(n2203), .B(n2204), .Z(n2202) );
  XOR U5791 ( .A(DB[1747]), .B(DB[1732]), .Z(n2204) );
  AND U5792 ( .A(n562), .B(n2205), .Z(n2203) );
  XOR U5793 ( .A(n2206), .B(n2207), .Z(n2205) );
  XOR U5794 ( .A(DB[1732]), .B(DB[1717]), .Z(n2207) );
  AND U5795 ( .A(n566), .B(n2208), .Z(n2206) );
  XOR U5796 ( .A(n2209), .B(n2210), .Z(n2208) );
  XOR U5797 ( .A(DB[1717]), .B(DB[1702]), .Z(n2210) );
  AND U5798 ( .A(n570), .B(n2211), .Z(n2209) );
  XOR U5799 ( .A(n2212), .B(n2213), .Z(n2211) );
  XOR U5800 ( .A(DB[1702]), .B(DB[1687]), .Z(n2213) );
  AND U5801 ( .A(n574), .B(n2214), .Z(n2212) );
  XOR U5802 ( .A(n2215), .B(n2216), .Z(n2214) );
  XOR U5803 ( .A(DB[1687]), .B(DB[1672]), .Z(n2216) );
  AND U5804 ( .A(n578), .B(n2217), .Z(n2215) );
  XOR U5805 ( .A(n2218), .B(n2219), .Z(n2217) );
  XOR U5806 ( .A(DB[1672]), .B(DB[1657]), .Z(n2219) );
  AND U5807 ( .A(n582), .B(n2220), .Z(n2218) );
  XOR U5808 ( .A(n2221), .B(n2222), .Z(n2220) );
  XOR U5809 ( .A(DB[1657]), .B(DB[1642]), .Z(n2222) );
  AND U5810 ( .A(n586), .B(n2223), .Z(n2221) );
  XOR U5811 ( .A(n2224), .B(n2225), .Z(n2223) );
  XOR U5812 ( .A(DB[1642]), .B(DB[1627]), .Z(n2225) );
  AND U5813 ( .A(n590), .B(n2226), .Z(n2224) );
  XOR U5814 ( .A(n2227), .B(n2228), .Z(n2226) );
  XOR U5815 ( .A(DB[1627]), .B(DB[1612]), .Z(n2228) );
  AND U5816 ( .A(n594), .B(n2229), .Z(n2227) );
  XOR U5817 ( .A(n2230), .B(n2231), .Z(n2229) );
  XOR U5818 ( .A(DB[1612]), .B(DB[1597]), .Z(n2231) );
  AND U5819 ( .A(n598), .B(n2232), .Z(n2230) );
  XOR U5820 ( .A(n2233), .B(n2234), .Z(n2232) );
  XOR U5821 ( .A(DB[1597]), .B(DB[1582]), .Z(n2234) );
  AND U5822 ( .A(n602), .B(n2235), .Z(n2233) );
  XOR U5823 ( .A(n2236), .B(n2237), .Z(n2235) );
  XOR U5824 ( .A(DB[1582]), .B(DB[1567]), .Z(n2237) );
  AND U5825 ( .A(n606), .B(n2238), .Z(n2236) );
  XOR U5826 ( .A(n2239), .B(n2240), .Z(n2238) );
  XOR U5827 ( .A(DB[1567]), .B(DB[1552]), .Z(n2240) );
  AND U5828 ( .A(n610), .B(n2241), .Z(n2239) );
  XOR U5829 ( .A(n2242), .B(n2243), .Z(n2241) );
  XOR U5830 ( .A(DB[1552]), .B(DB[1537]), .Z(n2243) );
  AND U5831 ( .A(n614), .B(n2244), .Z(n2242) );
  XOR U5832 ( .A(n2245), .B(n2246), .Z(n2244) );
  XOR U5833 ( .A(DB[1537]), .B(DB[1522]), .Z(n2246) );
  AND U5834 ( .A(n618), .B(n2247), .Z(n2245) );
  XOR U5835 ( .A(n2248), .B(n2249), .Z(n2247) );
  XOR U5836 ( .A(DB[1522]), .B(DB[1507]), .Z(n2249) );
  AND U5837 ( .A(n622), .B(n2250), .Z(n2248) );
  XOR U5838 ( .A(n2251), .B(n2252), .Z(n2250) );
  XOR U5839 ( .A(DB[1507]), .B(DB[1492]), .Z(n2252) );
  AND U5840 ( .A(n626), .B(n2253), .Z(n2251) );
  XOR U5841 ( .A(n2254), .B(n2255), .Z(n2253) );
  XOR U5842 ( .A(DB[1492]), .B(DB[1477]), .Z(n2255) );
  AND U5843 ( .A(n630), .B(n2256), .Z(n2254) );
  XOR U5844 ( .A(n2257), .B(n2258), .Z(n2256) );
  XOR U5845 ( .A(DB[1477]), .B(DB[1462]), .Z(n2258) );
  AND U5846 ( .A(n634), .B(n2259), .Z(n2257) );
  XOR U5847 ( .A(n2260), .B(n2261), .Z(n2259) );
  XOR U5848 ( .A(DB[1462]), .B(DB[1447]), .Z(n2261) );
  AND U5849 ( .A(n638), .B(n2262), .Z(n2260) );
  XOR U5850 ( .A(n2263), .B(n2264), .Z(n2262) );
  XOR U5851 ( .A(DB[1447]), .B(DB[1432]), .Z(n2264) );
  AND U5852 ( .A(n642), .B(n2265), .Z(n2263) );
  XOR U5853 ( .A(n2266), .B(n2267), .Z(n2265) );
  XOR U5854 ( .A(DB[1432]), .B(DB[1417]), .Z(n2267) );
  AND U5855 ( .A(n646), .B(n2268), .Z(n2266) );
  XOR U5856 ( .A(n2269), .B(n2270), .Z(n2268) );
  XOR U5857 ( .A(DB[1417]), .B(DB[1402]), .Z(n2270) );
  AND U5858 ( .A(n650), .B(n2271), .Z(n2269) );
  XOR U5859 ( .A(n2272), .B(n2273), .Z(n2271) );
  XOR U5860 ( .A(DB[1402]), .B(DB[1387]), .Z(n2273) );
  AND U5861 ( .A(n654), .B(n2274), .Z(n2272) );
  XOR U5862 ( .A(n2275), .B(n2276), .Z(n2274) );
  XOR U5863 ( .A(DB[1387]), .B(DB[1372]), .Z(n2276) );
  AND U5864 ( .A(n658), .B(n2277), .Z(n2275) );
  XOR U5865 ( .A(n2278), .B(n2279), .Z(n2277) );
  XOR U5866 ( .A(DB[1372]), .B(DB[1357]), .Z(n2279) );
  AND U5867 ( .A(n662), .B(n2280), .Z(n2278) );
  XOR U5868 ( .A(n2281), .B(n2282), .Z(n2280) );
  XOR U5869 ( .A(DB[1357]), .B(DB[1342]), .Z(n2282) );
  AND U5870 ( .A(n666), .B(n2283), .Z(n2281) );
  XOR U5871 ( .A(n2284), .B(n2285), .Z(n2283) );
  XOR U5872 ( .A(DB[1342]), .B(DB[1327]), .Z(n2285) );
  AND U5873 ( .A(n670), .B(n2286), .Z(n2284) );
  XOR U5874 ( .A(n2287), .B(n2288), .Z(n2286) );
  XOR U5875 ( .A(DB[1327]), .B(DB[1312]), .Z(n2288) );
  AND U5876 ( .A(n674), .B(n2289), .Z(n2287) );
  XOR U5877 ( .A(n2290), .B(n2291), .Z(n2289) );
  XOR U5878 ( .A(DB[1312]), .B(DB[1297]), .Z(n2291) );
  AND U5879 ( .A(n678), .B(n2292), .Z(n2290) );
  XOR U5880 ( .A(n2293), .B(n2294), .Z(n2292) );
  XOR U5881 ( .A(DB[1297]), .B(DB[1282]), .Z(n2294) );
  AND U5882 ( .A(n682), .B(n2295), .Z(n2293) );
  XOR U5883 ( .A(n2296), .B(n2297), .Z(n2295) );
  XOR U5884 ( .A(DB[1282]), .B(DB[1267]), .Z(n2297) );
  AND U5885 ( .A(n686), .B(n2298), .Z(n2296) );
  XOR U5886 ( .A(n2299), .B(n2300), .Z(n2298) );
  XOR U5887 ( .A(DB[1267]), .B(DB[1252]), .Z(n2300) );
  AND U5888 ( .A(n690), .B(n2301), .Z(n2299) );
  XOR U5889 ( .A(n2302), .B(n2303), .Z(n2301) );
  XOR U5890 ( .A(DB[1252]), .B(DB[1237]), .Z(n2303) );
  AND U5891 ( .A(n694), .B(n2304), .Z(n2302) );
  XOR U5892 ( .A(n2305), .B(n2306), .Z(n2304) );
  XOR U5893 ( .A(DB[1237]), .B(DB[1222]), .Z(n2306) );
  AND U5894 ( .A(n698), .B(n2307), .Z(n2305) );
  XOR U5895 ( .A(n2308), .B(n2309), .Z(n2307) );
  XOR U5896 ( .A(DB[1222]), .B(DB[1207]), .Z(n2309) );
  AND U5897 ( .A(n702), .B(n2310), .Z(n2308) );
  XOR U5898 ( .A(n2311), .B(n2312), .Z(n2310) );
  XOR U5899 ( .A(DB[1207]), .B(DB[1192]), .Z(n2312) );
  AND U5900 ( .A(n706), .B(n2313), .Z(n2311) );
  XOR U5901 ( .A(n2314), .B(n2315), .Z(n2313) );
  XOR U5902 ( .A(DB[1192]), .B(DB[1177]), .Z(n2315) );
  AND U5903 ( .A(n710), .B(n2316), .Z(n2314) );
  XOR U5904 ( .A(n2317), .B(n2318), .Z(n2316) );
  XOR U5905 ( .A(DB[1177]), .B(DB[1162]), .Z(n2318) );
  AND U5906 ( .A(n714), .B(n2319), .Z(n2317) );
  XOR U5907 ( .A(n2320), .B(n2321), .Z(n2319) );
  XOR U5908 ( .A(DB[1162]), .B(DB[1147]), .Z(n2321) );
  AND U5909 ( .A(n718), .B(n2322), .Z(n2320) );
  XOR U5910 ( .A(n2323), .B(n2324), .Z(n2322) );
  XOR U5911 ( .A(DB[1147]), .B(DB[1132]), .Z(n2324) );
  AND U5912 ( .A(n722), .B(n2325), .Z(n2323) );
  XOR U5913 ( .A(n2326), .B(n2327), .Z(n2325) );
  XOR U5914 ( .A(DB[1132]), .B(DB[1117]), .Z(n2327) );
  AND U5915 ( .A(n726), .B(n2328), .Z(n2326) );
  XOR U5916 ( .A(n2329), .B(n2330), .Z(n2328) );
  XOR U5917 ( .A(DB[1117]), .B(DB[1102]), .Z(n2330) );
  AND U5918 ( .A(n730), .B(n2331), .Z(n2329) );
  XOR U5919 ( .A(n2332), .B(n2333), .Z(n2331) );
  XOR U5920 ( .A(DB[1102]), .B(DB[1087]), .Z(n2333) );
  AND U5921 ( .A(n734), .B(n2334), .Z(n2332) );
  XOR U5922 ( .A(n2335), .B(n2336), .Z(n2334) );
  XOR U5923 ( .A(DB[1087]), .B(DB[1072]), .Z(n2336) );
  AND U5924 ( .A(n738), .B(n2337), .Z(n2335) );
  XOR U5925 ( .A(n2338), .B(n2339), .Z(n2337) );
  XOR U5926 ( .A(DB[1072]), .B(DB[1057]), .Z(n2339) );
  AND U5927 ( .A(n742), .B(n2340), .Z(n2338) );
  XOR U5928 ( .A(n2341), .B(n2342), .Z(n2340) );
  XOR U5929 ( .A(DB[1057]), .B(DB[1042]), .Z(n2342) );
  AND U5930 ( .A(n746), .B(n2343), .Z(n2341) );
  XOR U5931 ( .A(n2344), .B(n2345), .Z(n2343) );
  XOR U5932 ( .A(DB[1042]), .B(DB[1027]), .Z(n2345) );
  AND U5933 ( .A(n750), .B(n2346), .Z(n2344) );
  XOR U5934 ( .A(n2347), .B(n2348), .Z(n2346) );
  XOR U5935 ( .A(DB[1027]), .B(DB[1012]), .Z(n2348) );
  AND U5936 ( .A(n754), .B(n2349), .Z(n2347) );
  XOR U5937 ( .A(n2350), .B(n2351), .Z(n2349) );
  XOR U5938 ( .A(DB[997]), .B(DB[1012]), .Z(n2351) );
  AND U5939 ( .A(n758), .B(n2352), .Z(n2350) );
  XOR U5940 ( .A(n2353), .B(n2354), .Z(n2352) );
  XOR U5941 ( .A(DB[997]), .B(DB[982]), .Z(n2354) );
  AND U5942 ( .A(n762), .B(n2355), .Z(n2353) );
  XOR U5943 ( .A(n2356), .B(n2357), .Z(n2355) );
  XOR U5944 ( .A(DB[982]), .B(DB[967]), .Z(n2357) );
  AND U5945 ( .A(n766), .B(n2358), .Z(n2356) );
  XOR U5946 ( .A(n2359), .B(n2360), .Z(n2358) );
  XOR U5947 ( .A(DB[967]), .B(DB[952]), .Z(n2360) );
  AND U5948 ( .A(n770), .B(n2361), .Z(n2359) );
  XOR U5949 ( .A(n2362), .B(n2363), .Z(n2361) );
  XOR U5950 ( .A(DB[952]), .B(DB[937]), .Z(n2363) );
  AND U5951 ( .A(n774), .B(n2364), .Z(n2362) );
  XOR U5952 ( .A(n2365), .B(n2366), .Z(n2364) );
  XOR U5953 ( .A(DB[937]), .B(DB[922]), .Z(n2366) );
  AND U5954 ( .A(n778), .B(n2367), .Z(n2365) );
  XOR U5955 ( .A(n2368), .B(n2369), .Z(n2367) );
  XOR U5956 ( .A(DB[922]), .B(DB[907]), .Z(n2369) );
  AND U5957 ( .A(n782), .B(n2370), .Z(n2368) );
  XOR U5958 ( .A(n2371), .B(n2372), .Z(n2370) );
  XOR U5959 ( .A(DB[907]), .B(DB[892]), .Z(n2372) );
  AND U5960 ( .A(n786), .B(n2373), .Z(n2371) );
  XOR U5961 ( .A(n2374), .B(n2375), .Z(n2373) );
  XOR U5962 ( .A(DB[892]), .B(DB[877]), .Z(n2375) );
  AND U5963 ( .A(n790), .B(n2376), .Z(n2374) );
  XOR U5964 ( .A(n2377), .B(n2378), .Z(n2376) );
  XOR U5965 ( .A(DB[877]), .B(DB[862]), .Z(n2378) );
  AND U5966 ( .A(n794), .B(n2379), .Z(n2377) );
  XOR U5967 ( .A(n2380), .B(n2381), .Z(n2379) );
  XOR U5968 ( .A(DB[862]), .B(DB[847]), .Z(n2381) );
  AND U5969 ( .A(n798), .B(n2382), .Z(n2380) );
  XOR U5970 ( .A(n2383), .B(n2384), .Z(n2382) );
  XOR U5971 ( .A(DB[847]), .B(DB[832]), .Z(n2384) );
  AND U5972 ( .A(n802), .B(n2385), .Z(n2383) );
  XOR U5973 ( .A(n2386), .B(n2387), .Z(n2385) );
  XOR U5974 ( .A(DB[832]), .B(DB[817]), .Z(n2387) );
  AND U5975 ( .A(n806), .B(n2388), .Z(n2386) );
  XOR U5976 ( .A(n2389), .B(n2390), .Z(n2388) );
  XOR U5977 ( .A(DB[817]), .B(DB[802]), .Z(n2390) );
  AND U5978 ( .A(n810), .B(n2391), .Z(n2389) );
  XOR U5979 ( .A(n2392), .B(n2393), .Z(n2391) );
  XOR U5980 ( .A(DB[802]), .B(DB[787]), .Z(n2393) );
  AND U5981 ( .A(n814), .B(n2394), .Z(n2392) );
  XOR U5982 ( .A(n2395), .B(n2396), .Z(n2394) );
  XOR U5983 ( .A(DB[787]), .B(DB[772]), .Z(n2396) );
  AND U5984 ( .A(n818), .B(n2397), .Z(n2395) );
  XOR U5985 ( .A(n2398), .B(n2399), .Z(n2397) );
  XOR U5986 ( .A(DB[772]), .B(DB[757]), .Z(n2399) );
  AND U5987 ( .A(n822), .B(n2400), .Z(n2398) );
  XOR U5988 ( .A(n2401), .B(n2402), .Z(n2400) );
  XOR U5989 ( .A(DB[757]), .B(DB[742]), .Z(n2402) );
  AND U5990 ( .A(n826), .B(n2403), .Z(n2401) );
  XOR U5991 ( .A(n2404), .B(n2405), .Z(n2403) );
  XOR U5992 ( .A(DB[742]), .B(DB[727]), .Z(n2405) );
  AND U5993 ( .A(n830), .B(n2406), .Z(n2404) );
  XOR U5994 ( .A(n2407), .B(n2408), .Z(n2406) );
  XOR U5995 ( .A(DB[727]), .B(DB[712]), .Z(n2408) );
  AND U5996 ( .A(n834), .B(n2409), .Z(n2407) );
  XOR U5997 ( .A(n2410), .B(n2411), .Z(n2409) );
  XOR U5998 ( .A(DB[712]), .B(DB[697]), .Z(n2411) );
  AND U5999 ( .A(n838), .B(n2412), .Z(n2410) );
  XOR U6000 ( .A(n2413), .B(n2414), .Z(n2412) );
  XOR U6001 ( .A(DB[697]), .B(DB[682]), .Z(n2414) );
  AND U6002 ( .A(n842), .B(n2415), .Z(n2413) );
  XOR U6003 ( .A(n2416), .B(n2417), .Z(n2415) );
  XOR U6004 ( .A(DB[682]), .B(DB[667]), .Z(n2417) );
  AND U6005 ( .A(n846), .B(n2418), .Z(n2416) );
  XOR U6006 ( .A(n2419), .B(n2420), .Z(n2418) );
  XOR U6007 ( .A(DB[667]), .B(DB[652]), .Z(n2420) );
  AND U6008 ( .A(n850), .B(n2421), .Z(n2419) );
  XOR U6009 ( .A(n2422), .B(n2423), .Z(n2421) );
  XOR U6010 ( .A(DB[652]), .B(DB[637]), .Z(n2423) );
  AND U6011 ( .A(n854), .B(n2424), .Z(n2422) );
  XOR U6012 ( .A(n2425), .B(n2426), .Z(n2424) );
  XOR U6013 ( .A(DB[637]), .B(DB[622]), .Z(n2426) );
  AND U6014 ( .A(n858), .B(n2427), .Z(n2425) );
  XOR U6015 ( .A(n2428), .B(n2429), .Z(n2427) );
  XOR U6016 ( .A(DB[622]), .B(DB[607]), .Z(n2429) );
  AND U6017 ( .A(n862), .B(n2430), .Z(n2428) );
  XOR U6018 ( .A(n2431), .B(n2432), .Z(n2430) );
  XOR U6019 ( .A(DB[607]), .B(DB[592]), .Z(n2432) );
  AND U6020 ( .A(n866), .B(n2433), .Z(n2431) );
  XOR U6021 ( .A(n2434), .B(n2435), .Z(n2433) );
  XOR U6022 ( .A(DB[592]), .B(DB[577]), .Z(n2435) );
  AND U6023 ( .A(n870), .B(n2436), .Z(n2434) );
  XOR U6024 ( .A(n2437), .B(n2438), .Z(n2436) );
  XOR U6025 ( .A(DB[577]), .B(DB[562]), .Z(n2438) );
  AND U6026 ( .A(n874), .B(n2439), .Z(n2437) );
  XOR U6027 ( .A(n2440), .B(n2441), .Z(n2439) );
  XOR U6028 ( .A(DB[562]), .B(DB[547]), .Z(n2441) );
  AND U6029 ( .A(n878), .B(n2442), .Z(n2440) );
  XOR U6030 ( .A(n2443), .B(n2444), .Z(n2442) );
  XOR U6031 ( .A(DB[547]), .B(DB[532]), .Z(n2444) );
  AND U6032 ( .A(n882), .B(n2445), .Z(n2443) );
  XOR U6033 ( .A(n2446), .B(n2447), .Z(n2445) );
  XOR U6034 ( .A(DB[532]), .B(DB[517]), .Z(n2447) );
  AND U6035 ( .A(n886), .B(n2448), .Z(n2446) );
  XOR U6036 ( .A(n2449), .B(n2450), .Z(n2448) );
  XOR U6037 ( .A(DB[517]), .B(DB[502]), .Z(n2450) );
  AND U6038 ( .A(n890), .B(n2451), .Z(n2449) );
  XOR U6039 ( .A(n2452), .B(n2453), .Z(n2451) );
  XOR U6040 ( .A(DB[502]), .B(DB[487]), .Z(n2453) );
  AND U6041 ( .A(n894), .B(n2454), .Z(n2452) );
  XOR U6042 ( .A(n2455), .B(n2456), .Z(n2454) );
  XOR U6043 ( .A(DB[487]), .B(DB[472]), .Z(n2456) );
  AND U6044 ( .A(n898), .B(n2457), .Z(n2455) );
  XOR U6045 ( .A(n2458), .B(n2459), .Z(n2457) );
  XOR U6046 ( .A(DB[472]), .B(DB[457]), .Z(n2459) );
  AND U6047 ( .A(n902), .B(n2460), .Z(n2458) );
  XOR U6048 ( .A(n2461), .B(n2462), .Z(n2460) );
  XOR U6049 ( .A(DB[457]), .B(DB[442]), .Z(n2462) );
  AND U6050 ( .A(n906), .B(n2463), .Z(n2461) );
  XOR U6051 ( .A(n2464), .B(n2465), .Z(n2463) );
  XOR U6052 ( .A(DB[442]), .B(DB[427]), .Z(n2465) );
  AND U6053 ( .A(n910), .B(n2466), .Z(n2464) );
  XOR U6054 ( .A(n2467), .B(n2468), .Z(n2466) );
  XOR U6055 ( .A(DB[427]), .B(DB[412]), .Z(n2468) );
  AND U6056 ( .A(n914), .B(n2469), .Z(n2467) );
  XOR U6057 ( .A(n2470), .B(n2471), .Z(n2469) );
  XOR U6058 ( .A(DB[412]), .B(DB[397]), .Z(n2471) );
  AND U6059 ( .A(n918), .B(n2472), .Z(n2470) );
  XOR U6060 ( .A(n2473), .B(n2474), .Z(n2472) );
  XOR U6061 ( .A(DB[397]), .B(DB[382]), .Z(n2474) );
  AND U6062 ( .A(n922), .B(n2475), .Z(n2473) );
  XOR U6063 ( .A(n2476), .B(n2477), .Z(n2475) );
  XOR U6064 ( .A(DB[382]), .B(DB[367]), .Z(n2477) );
  AND U6065 ( .A(n926), .B(n2478), .Z(n2476) );
  XOR U6066 ( .A(n2479), .B(n2480), .Z(n2478) );
  XOR U6067 ( .A(DB[367]), .B(DB[352]), .Z(n2480) );
  AND U6068 ( .A(n930), .B(n2481), .Z(n2479) );
  XOR U6069 ( .A(n2482), .B(n2483), .Z(n2481) );
  XOR U6070 ( .A(DB[352]), .B(DB[337]), .Z(n2483) );
  AND U6071 ( .A(n934), .B(n2484), .Z(n2482) );
  XOR U6072 ( .A(n2485), .B(n2486), .Z(n2484) );
  XOR U6073 ( .A(DB[337]), .B(DB[322]), .Z(n2486) );
  AND U6074 ( .A(n938), .B(n2487), .Z(n2485) );
  XOR U6075 ( .A(n2488), .B(n2489), .Z(n2487) );
  XOR U6076 ( .A(DB[322]), .B(DB[307]), .Z(n2489) );
  AND U6077 ( .A(n942), .B(n2490), .Z(n2488) );
  XOR U6078 ( .A(n2491), .B(n2492), .Z(n2490) );
  XOR U6079 ( .A(DB[307]), .B(DB[292]), .Z(n2492) );
  AND U6080 ( .A(n946), .B(n2493), .Z(n2491) );
  XOR U6081 ( .A(n2494), .B(n2495), .Z(n2493) );
  XOR U6082 ( .A(DB[292]), .B(DB[277]), .Z(n2495) );
  AND U6083 ( .A(n950), .B(n2496), .Z(n2494) );
  XOR U6084 ( .A(n2497), .B(n2498), .Z(n2496) );
  XOR U6085 ( .A(DB[277]), .B(DB[262]), .Z(n2498) );
  AND U6086 ( .A(n954), .B(n2499), .Z(n2497) );
  XOR U6087 ( .A(n2500), .B(n2501), .Z(n2499) );
  XOR U6088 ( .A(DB[262]), .B(DB[247]), .Z(n2501) );
  AND U6089 ( .A(n958), .B(n2502), .Z(n2500) );
  XOR U6090 ( .A(n2503), .B(n2504), .Z(n2502) );
  XOR U6091 ( .A(DB[247]), .B(DB[232]), .Z(n2504) );
  AND U6092 ( .A(n962), .B(n2505), .Z(n2503) );
  XOR U6093 ( .A(n2506), .B(n2507), .Z(n2505) );
  XOR U6094 ( .A(DB[232]), .B(DB[217]), .Z(n2507) );
  AND U6095 ( .A(n966), .B(n2508), .Z(n2506) );
  XOR U6096 ( .A(n2509), .B(n2510), .Z(n2508) );
  XOR U6097 ( .A(DB[217]), .B(DB[202]), .Z(n2510) );
  AND U6098 ( .A(n970), .B(n2511), .Z(n2509) );
  XOR U6099 ( .A(n2512), .B(n2513), .Z(n2511) );
  XOR U6100 ( .A(DB[202]), .B(DB[187]), .Z(n2513) );
  AND U6101 ( .A(n974), .B(n2514), .Z(n2512) );
  XOR U6102 ( .A(n2515), .B(n2516), .Z(n2514) );
  XOR U6103 ( .A(DB[187]), .B(DB[172]), .Z(n2516) );
  AND U6104 ( .A(n978), .B(n2517), .Z(n2515) );
  XOR U6105 ( .A(n2518), .B(n2519), .Z(n2517) );
  XOR U6106 ( .A(DB[172]), .B(DB[157]), .Z(n2519) );
  AND U6107 ( .A(n982), .B(n2520), .Z(n2518) );
  XOR U6108 ( .A(n2521), .B(n2522), .Z(n2520) );
  XOR U6109 ( .A(DB[157]), .B(DB[142]), .Z(n2522) );
  AND U6110 ( .A(n986), .B(n2523), .Z(n2521) );
  XOR U6111 ( .A(n2524), .B(n2525), .Z(n2523) );
  XOR U6112 ( .A(DB[142]), .B(DB[127]), .Z(n2525) );
  AND U6113 ( .A(n990), .B(n2526), .Z(n2524) );
  XOR U6114 ( .A(n2527), .B(n2528), .Z(n2526) );
  XOR U6115 ( .A(DB[127]), .B(DB[112]), .Z(n2528) );
  AND U6116 ( .A(n994), .B(n2529), .Z(n2527) );
  XOR U6117 ( .A(n2530), .B(n2531), .Z(n2529) );
  XOR U6118 ( .A(DB[97]), .B(DB[112]), .Z(n2531) );
  AND U6119 ( .A(n998), .B(n2532), .Z(n2530) );
  XOR U6120 ( .A(n2533), .B(n2534), .Z(n2532) );
  XOR U6121 ( .A(DB[97]), .B(DB[82]), .Z(n2534) );
  AND U6122 ( .A(n1002), .B(n2535), .Z(n2533) );
  XOR U6123 ( .A(n2536), .B(n2537), .Z(n2535) );
  XOR U6124 ( .A(DB[82]), .B(DB[67]), .Z(n2537) );
  AND U6125 ( .A(n1006), .B(n2538), .Z(n2536) );
  XOR U6126 ( .A(n2539), .B(n2540), .Z(n2538) );
  XOR U6127 ( .A(DB[67]), .B(DB[52]), .Z(n2540) );
  AND U6128 ( .A(n1010), .B(n2541), .Z(n2539) );
  XOR U6129 ( .A(n2542), .B(n2543), .Z(n2541) );
  XOR U6130 ( .A(DB[52]), .B(DB[37]), .Z(n2543) );
  AND U6131 ( .A(n1014), .B(n2544), .Z(n2542) );
  XOR U6132 ( .A(n2545), .B(n2546), .Z(n2544) );
  XOR U6133 ( .A(DB[37]), .B(DB[22]), .Z(n2546) );
  AND U6134 ( .A(n1018), .B(n2547), .Z(n2545) );
  XOR U6135 ( .A(DB[7]), .B(DB[22]), .Z(n2547) );
  XOR U6136 ( .A(DB[3831]), .B(n2548), .Z(min_val_out[6]) );
  AND U6137 ( .A(n2), .B(n2549), .Z(n2548) );
  XOR U6138 ( .A(n2550), .B(n2551), .Z(n2549) );
  XOR U6139 ( .A(DB[3831]), .B(DB[3816]), .Z(n2551) );
  AND U6140 ( .A(n6), .B(n2552), .Z(n2550) );
  XOR U6141 ( .A(n2553), .B(n2554), .Z(n2552) );
  XOR U6142 ( .A(DB[3816]), .B(DB[3801]), .Z(n2554) );
  AND U6143 ( .A(n10), .B(n2555), .Z(n2553) );
  XOR U6144 ( .A(n2556), .B(n2557), .Z(n2555) );
  XOR U6145 ( .A(DB[3801]), .B(DB[3786]), .Z(n2557) );
  AND U6146 ( .A(n14), .B(n2558), .Z(n2556) );
  XOR U6147 ( .A(n2559), .B(n2560), .Z(n2558) );
  XOR U6148 ( .A(DB[3786]), .B(DB[3771]), .Z(n2560) );
  AND U6149 ( .A(n18), .B(n2561), .Z(n2559) );
  XOR U6150 ( .A(n2562), .B(n2563), .Z(n2561) );
  XOR U6151 ( .A(DB[3771]), .B(DB[3756]), .Z(n2563) );
  AND U6152 ( .A(n22), .B(n2564), .Z(n2562) );
  XOR U6153 ( .A(n2565), .B(n2566), .Z(n2564) );
  XOR U6154 ( .A(DB[3756]), .B(DB[3741]), .Z(n2566) );
  AND U6155 ( .A(n26), .B(n2567), .Z(n2565) );
  XOR U6156 ( .A(n2568), .B(n2569), .Z(n2567) );
  XOR U6157 ( .A(DB[3741]), .B(DB[3726]), .Z(n2569) );
  AND U6158 ( .A(n30), .B(n2570), .Z(n2568) );
  XOR U6159 ( .A(n2571), .B(n2572), .Z(n2570) );
  XOR U6160 ( .A(DB[3726]), .B(DB[3711]), .Z(n2572) );
  AND U6161 ( .A(n34), .B(n2573), .Z(n2571) );
  XOR U6162 ( .A(n2574), .B(n2575), .Z(n2573) );
  XOR U6163 ( .A(DB[3711]), .B(DB[3696]), .Z(n2575) );
  AND U6164 ( .A(n38), .B(n2576), .Z(n2574) );
  XOR U6165 ( .A(n2577), .B(n2578), .Z(n2576) );
  XOR U6166 ( .A(DB[3696]), .B(DB[3681]), .Z(n2578) );
  AND U6167 ( .A(n42), .B(n2579), .Z(n2577) );
  XOR U6168 ( .A(n2580), .B(n2581), .Z(n2579) );
  XOR U6169 ( .A(DB[3681]), .B(DB[3666]), .Z(n2581) );
  AND U6170 ( .A(n46), .B(n2582), .Z(n2580) );
  XOR U6171 ( .A(n2583), .B(n2584), .Z(n2582) );
  XOR U6172 ( .A(DB[3666]), .B(DB[3651]), .Z(n2584) );
  AND U6173 ( .A(n50), .B(n2585), .Z(n2583) );
  XOR U6174 ( .A(n2586), .B(n2587), .Z(n2585) );
  XOR U6175 ( .A(DB[3651]), .B(DB[3636]), .Z(n2587) );
  AND U6176 ( .A(n54), .B(n2588), .Z(n2586) );
  XOR U6177 ( .A(n2589), .B(n2590), .Z(n2588) );
  XOR U6178 ( .A(DB[3636]), .B(DB[3621]), .Z(n2590) );
  AND U6179 ( .A(n58), .B(n2591), .Z(n2589) );
  XOR U6180 ( .A(n2592), .B(n2593), .Z(n2591) );
  XOR U6181 ( .A(DB[3621]), .B(DB[3606]), .Z(n2593) );
  AND U6182 ( .A(n62), .B(n2594), .Z(n2592) );
  XOR U6183 ( .A(n2595), .B(n2596), .Z(n2594) );
  XOR U6184 ( .A(DB[3606]), .B(DB[3591]), .Z(n2596) );
  AND U6185 ( .A(n66), .B(n2597), .Z(n2595) );
  XOR U6186 ( .A(n2598), .B(n2599), .Z(n2597) );
  XOR U6187 ( .A(DB[3591]), .B(DB[3576]), .Z(n2599) );
  AND U6188 ( .A(n70), .B(n2600), .Z(n2598) );
  XOR U6189 ( .A(n2601), .B(n2602), .Z(n2600) );
  XOR U6190 ( .A(DB[3576]), .B(DB[3561]), .Z(n2602) );
  AND U6191 ( .A(n74), .B(n2603), .Z(n2601) );
  XOR U6192 ( .A(n2604), .B(n2605), .Z(n2603) );
  XOR U6193 ( .A(DB[3561]), .B(DB[3546]), .Z(n2605) );
  AND U6194 ( .A(n78), .B(n2606), .Z(n2604) );
  XOR U6195 ( .A(n2607), .B(n2608), .Z(n2606) );
  XOR U6196 ( .A(DB[3546]), .B(DB[3531]), .Z(n2608) );
  AND U6197 ( .A(n82), .B(n2609), .Z(n2607) );
  XOR U6198 ( .A(n2610), .B(n2611), .Z(n2609) );
  XOR U6199 ( .A(DB[3531]), .B(DB[3516]), .Z(n2611) );
  AND U6200 ( .A(n86), .B(n2612), .Z(n2610) );
  XOR U6201 ( .A(n2613), .B(n2614), .Z(n2612) );
  XOR U6202 ( .A(DB[3516]), .B(DB[3501]), .Z(n2614) );
  AND U6203 ( .A(n90), .B(n2615), .Z(n2613) );
  XOR U6204 ( .A(n2616), .B(n2617), .Z(n2615) );
  XOR U6205 ( .A(DB[3501]), .B(DB[3486]), .Z(n2617) );
  AND U6206 ( .A(n94), .B(n2618), .Z(n2616) );
  XOR U6207 ( .A(n2619), .B(n2620), .Z(n2618) );
  XOR U6208 ( .A(DB[3486]), .B(DB[3471]), .Z(n2620) );
  AND U6209 ( .A(n98), .B(n2621), .Z(n2619) );
  XOR U6210 ( .A(n2622), .B(n2623), .Z(n2621) );
  XOR U6211 ( .A(DB[3471]), .B(DB[3456]), .Z(n2623) );
  AND U6212 ( .A(n102), .B(n2624), .Z(n2622) );
  XOR U6213 ( .A(n2625), .B(n2626), .Z(n2624) );
  XOR U6214 ( .A(DB[3456]), .B(DB[3441]), .Z(n2626) );
  AND U6215 ( .A(n106), .B(n2627), .Z(n2625) );
  XOR U6216 ( .A(n2628), .B(n2629), .Z(n2627) );
  XOR U6217 ( .A(DB[3441]), .B(DB[3426]), .Z(n2629) );
  AND U6218 ( .A(n110), .B(n2630), .Z(n2628) );
  XOR U6219 ( .A(n2631), .B(n2632), .Z(n2630) );
  XOR U6220 ( .A(DB[3426]), .B(DB[3411]), .Z(n2632) );
  AND U6221 ( .A(n114), .B(n2633), .Z(n2631) );
  XOR U6222 ( .A(n2634), .B(n2635), .Z(n2633) );
  XOR U6223 ( .A(DB[3411]), .B(DB[3396]), .Z(n2635) );
  AND U6224 ( .A(n118), .B(n2636), .Z(n2634) );
  XOR U6225 ( .A(n2637), .B(n2638), .Z(n2636) );
  XOR U6226 ( .A(DB[3396]), .B(DB[3381]), .Z(n2638) );
  AND U6227 ( .A(n122), .B(n2639), .Z(n2637) );
  XOR U6228 ( .A(n2640), .B(n2641), .Z(n2639) );
  XOR U6229 ( .A(DB[3381]), .B(DB[3366]), .Z(n2641) );
  AND U6230 ( .A(n126), .B(n2642), .Z(n2640) );
  XOR U6231 ( .A(n2643), .B(n2644), .Z(n2642) );
  XOR U6232 ( .A(DB[3366]), .B(DB[3351]), .Z(n2644) );
  AND U6233 ( .A(n130), .B(n2645), .Z(n2643) );
  XOR U6234 ( .A(n2646), .B(n2647), .Z(n2645) );
  XOR U6235 ( .A(DB[3351]), .B(DB[3336]), .Z(n2647) );
  AND U6236 ( .A(n134), .B(n2648), .Z(n2646) );
  XOR U6237 ( .A(n2649), .B(n2650), .Z(n2648) );
  XOR U6238 ( .A(DB[3336]), .B(DB[3321]), .Z(n2650) );
  AND U6239 ( .A(n138), .B(n2651), .Z(n2649) );
  XOR U6240 ( .A(n2652), .B(n2653), .Z(n2651) );
  XOR U6241 ( .A(DB[3321]), .B(DB[3306]), .Z(n2653) );
  AND U6242 ( .A(n142), .B(n2654), .Z(n2652) );
  XOR U6243 ( .A(n2655), .B(n2656), .Z(n2654) );
  XOR U6244 ( .A(DB[3306]), .B(DB[3291]), .Z(n2656) );
  AND U6245 ( .A(n146), .B(n2657), .Z(n2655) );
  XOR U6246 ( .A(n2658), .B(n2659), .Z(n2657) );
  XOR U6247 ( .A(DB[3291]), .B(DB[3276]), .Z(n2659) );
  AND U6248 ( .A(n150), .B(n2660), .Z(n2658) );
  XOR U6249 ( .A(n2661), .B(n2662), .Z(n2660) );
  XOR U6250 ( .A(DB[3276]), .B(DB[3261]), .Z(n2662) );
  AND U6251 ( .A(n154), .B(n2663), .Z(n2661) );
  XOR U6252 ( .A(n2664), .B(n2665), .Z(n2663) );
  XOR U6253 ( .A(DB[3261]), .B(DB[3246]), .Z(n2665) );
  AND U6254 ( .A(n158), .B(n2666), .Z(n2664) );
  XOR U6255 ( .A(n2667), .B(n2668), .Z(n2666) );
  XOR U6256 ( .A(DB[3246]), .B(DB[3231]), .Z(n2668) );
  AND U6257 ( .A(n162), .B(n2669), .Z(n2667) );
  XOR U6258 ( .A(n2670), .B(n2671), .Z(n2669) );
  XOR U6259 ( .A(DB[3231]), .B(DB[3216]), .Z(n2671) );
  AND U6260 ( .A(n166), .B(n2672), .Z(n2670) );
  XOR U6261 ( .A(n2673), .B(n2674), .Z(n2672) );
  XOR U6262 ( .A(DB[3216]), .B(DB[3201]), .Z(n2674) );
  AND U6263 ( .A(n170), .B(n2675), .Z(n2673) );
  XOR U6264 ( .A(n2676), .B(n2677), .Z(n2675) );
  XOR U6265 ( .A(DB[3201]), .B(DB[3186]), .Z(n2677) );
  AND U6266 ( .A(n174), .B(n2678), .Z(n2676) );
  XOR U6267 ( .A(n2679), .B(n2680), .Z(n2678) );
  XOR U6268 ( .A(DB[3186]), .B(DB[3171]), .Z(n2680) );
  AND U6269 ( .A(n178), .B(n2681), .Z(n2679) );
  XOR U6270 ( .A(n2682), .B(n2683), .Z(n2681) );
  XOR U6271 ( .A(DB[3171]), .B(DB[3156]), .Z(n2683) );
  AND U6272 ( .A(n182), .B(n2684), .Z(n2682) );
  XOR U6273 ( .A(n2685), .B(n2686), .Z(n2684) );
  XOR U6274 ( .A(DB[3156]), .B(DB[3141]), .Z(n2686) );
  AND U6275 ( .A(n186), .B(n2687), .Z(n2685) );
  XOR U6276 ( .A(n2688), .B(n2689), .Z(n2687) );
  XOR U6277 ( .A(DB[3141]), .B(DB[3126]), .Z(n2689) );
  AND U6278 ( .A(n190), .B(n2690), .Z(n2688) );
  XOR U6279 ( .A(n2691), .B(n2692), .Z(n2690) );
  XOR U6280 ( .A(DB[3126]), .B(DB[3111]), .Z(n2692) );
  AND U6281 ( .A(n194), .B(n2693), .Z(n2691) );
  XOR U6282 ( .A(n2694), .B(n2695), .Z(n2693) );
  XOR U6283 ( .A(DB[3111]), .B(DB[3096]), .Z(n2695) );
  AND U6284 ( .A(n198), .B(n2696), .Z(n2694) );
  XOR U6285 ( .A(n2697), .B(n2698), .Z(n2696) );
  XOR U6286 ( .A(DB[3096]), .B(DB[3081]), .Z(n2698) );
  AND U6287 ( .A(n202), .B(n2699), .Z(n2697) );
  XOR U6288 ( .A(n2700), .B(n2701), .Z(n2699) );
  XOR U6289 ( .A(DB[3081]), .B(DB[3066]), .Z(n2701) );
  AND U6290 ( .A(n206), .B(n2702), .Z(n2700) );
  XOR U6291 ( .A(n2703), .B(n2704), .Z(n2702) );
  XOR U6292 ( .A(DB[3066]), .B(DB[3051]), .Z(n2704) );
  AND U6293 ( .A(n210), .B(n2705), .Z(n2703) );
  XOR U6294 ( .A(n2706), .B(n2707), .Z(n2705) );
  XOR U6295 ( .A(DB[3051]), .B(DB[3036]), .Z(n2707) );
  AND U6296 ( .A(n214), .B(n2708), .Z(n2706) );
  XOR U6297 ( .A(n2709), .B(n2710), .Z(n2708) );
  XOR U6298 ( .A(DB[3036]), .B(DB[3021]), .Z(n2710) );
  AND U6299 ( .A(n218), .B(n2711), .Z(n2709) );
  XOR U6300 ( .A(n2712), .B(n2713), .Z(n2711) );
  XOR U6301 ( .A(DB[3021]), .B(DB[3006]), .Z(n2713) );
  AND U6302 ( .A(n222), .B(n2714), .Z(n2712) );
  XOR U6303 ( .A(n2715), .B(n2716), .Z(n2714) );
  XOR U6304 ( .A(DB[3006]), .B(DB[2991]), .Z(n2716) );
  AND U6305 ( .A(n226), .B(n2717), .Z(n2715) );
  XOR U6306 ( .A(n2718), .B(n2719), .Z(n2717) );
  XOR U6307 ( .A(DB[2991]), .B(DB[2976]), .Z(n2719) );
  AND U6308 ( .A(n230), .B(n2720), .Z(n2718) );
  XOR U6309 ( .A(n2721), .B(n2722), .Z(n2720) );
  XOR U6310 ( .A(DB[2976]), .B(DB[2961]), .Z(n2722) );
  AND U6311 ( .A(n234), .B(n2723), .Z(n2721) );
  XOR U6312 ( .A(n2724), .B(n2725), .Z(n2723) );
  XOR U6313 ( .A(DB[2961]), .B(DB[2946]), .Z(n2725) );
  AND U6314 ( .A(n238), .B(n2726), .Z(n2724) );
  XOR U6315 ( .A(n2727), .B(n2728), .Z(n2726) );
  XOR U6316 ( .A(DB[2946]), .B(DB[2931]), .Z(n2728) );
  AND U6317 ( .A(n242), .B(n2729), .Z(n2727) );
  XOR U6318 ( .A(n2730), .B(n2731), .Z(n2729) );
  XOR U6319 ( .A(DB[2931]), .B(DB[2916]), .Z(n2731) );
  AND U6320 ( .A(n246), .B(n2732), .Z(n2730) );
  XOR U6321 ( .A(n2733), .B(n2734), .Z(n2732) );
  XOR U6322 ( .A(DB[2916]), .B(DB[2901]), .Z(n2734) );
  AND U6323 ( .A(n250), .B(n2735), .Z(n2733) );
  XOR U6324 ( .A(n2736), .B(n2737), .Z(n2735) );
  XOR U6325 ( .A(DB[2901]), .B(DB[2886]), .Z(n2737) );
  AND U6326 ( .A(n254), .B(n2738), .Z(n2736) );
  XOR U6327 ( .A(n2739), .B(n2740), .Z(n2738) );
  XOR U6328 ( .A(DB[2886]), .B(DB[2871]), .Z(n2740) );
  AND U6329 ( .A(n258), .B(n2741), .Z(n2739) );
  XOR U6330 ( .A(n2742), .B(n2743), .Z(n2741) );
  XOR U6331 ( .A(DB[2871]), .B(DB[2856]), .Z(n2743) );
  AND U6332 ( .A(n262), .B(n2744), .Z(n2742) );
  XOR U6333 ( .A(n2745), .B(n2746), .Z(n2744) );
  XOR U6334 ( .A(DB[2856]), .B(DB[2841]), .Z(n2746) );
  AND U6335 ( .A(n266), .B(n2747), .Z(n2745) );
  XOR U6336 ( .A(n2748), .B(n2749), .Z(n2747) );
  XOR U6337 ( .A(DB[2841]), .B(DB[2826]), .Z(n2749) );
  AND U6338 ( .A(n270), .B(n2750), .Z(n2748) );
  XOR U6339 ( .A(n2751), .B(n2752), .Z(n2750) );
  XOR U6340 ( .A(DB[2826]), .B(DB[2811]), .Z(n2752) );
  AND U6341 ( .A(n274), .B(n2753), .Z(n2751) );
  XOR U6342 ( .A(n2754), .B(n2755), .Z(n2753) );
  XOR U6343 ( .A(DB[2811]), .B(DB[2796]), .Z(n2755) );
  AND U6344 ( .A(n278), .B(n2756), .Z(n2754) );
  XOR U6345 ( .A(n2757), .B(n2758), .Z(n2756) );
  XOR U6346 ( .A(DB[2796]), .B(DB[2781]), .Z(n2758) );
  AND U6347 ( .A(n282), .B(n2759), .Z(n2757) );
  XOR U6348 ( .A(n2760), .B(n2761), .Z(n2759) );
  XOR U6349 ( .A(DB[2781]), .B(DB[2766]), .Z(n2761) );
  AND U6350 ( .A(n286), .B(n2762), .Z(n2760) );
  XOR U6351 ( .A(n2763), .B(n2764), .Z(n2762) );
  XOR U6352 ( .A(DB[2766]), .B(DB[2751]), .Z(n2764) );
  AND U6353 ( .A(n290), .B(n2765), .Z(n2763) );
  XOR U6354 ( .A(n2766), .B(n2767), .Z(n2765) );
  XOR U6355 ( .A(DB[2751]), .B(DB[2736]), .Z(n2767) );
  AND U6356 ( .A(n294), .B(n2768), .Z(n2766) );
  XOR U6357 ( .A(n2769), .B(n2770), .Z(n2768) );
  XOR U6358 ( .A(DB[2736]), .B(DB[2721]), .Z(n2770) );
  AND U6359 ( .A(n298), .B(n2771), .Z(n2769) );
  XOR U6360 ( .A(n2772), .B(n2773), .Z(n2771) );
  XOR U6361 ( .A(DB[2721]), .B(DB[2706]), .Z(n2773) );
  AND U6362 ( .A(n302), .B(n2774), .Z(n2772) );
  XOR U6363 ( .A(n2775), .B(n2776), .Z(n2774) );
  XOR U6364 ( .A(DB[2706]), .B(DB[2691]), .Z(n2776) );
  AND U6365 ( .A(n306), .B(n2777), .Z(n2775) );
  XOR U6366 ( .A(n2778), .B(n2779), .Z(n2777) );
  XOR U6367 ( .A(DB[2691]), .B(DB[2676]), .Z(n2779) );
  AND U6368 ( .A(n310), .B(n2780), .Z(n2778) );
  XOR U6369 ( .A(n2781), .B(n2782), .Z(n2780) );
  XOR U6370 ( .A(DB[2676]), .B(DB[2661]), .Z(n2782) );
  AND U6371 ( .A(n314), .B(n2783), .Z(n2781) );
  XOR U6372 ( .A(n2784), .B(n2785), .Z(n2783) );
  XOR U6373 ( .A(DB[2661]), .B(DB[2646]), .Z(n2785) );
  AND U6374 ( .A(n318), .B(n2786), .Z(n2784) );
  XOR U6375 ( .A(n2787), .B(n2788), .Z(n2786) );
  XOR U6376 ( .A(DB[2646]), .B(DB[2631]), .Z(n2788) );
  AND U6377 ( .A(n322), .B(n2789), .Z(n2787) );
  XOR U6378 ( .A(n2790), .B(n2791), .Z(n2789) );
  XOR U6379 ( .A(DB[2631]), .B(DB[2616]), .Z(n2791) );
  AND U6380 ( .A(n326), .B(n2792), .Z(n2790) );
  XOR U6381 ( .A(n2793), .B(n2794), .Z(n2792) );
  XOR U6382 ( .A(DB[2616]), .B(DB[2601]), .Z(n2794) );
  AND U6383 ( .A(n330), .B(n2795), .Z(n2793) );
  XOR U6384 ( .A(n2796), .B(n2797), .Z(n2795) );
  XOR U6385 ( .A(DB[2601]), .B(DB[2586]), .Z(n2797) );
  AND U6386 ( .A(n334), .B(n2798), .Z(n2796) );
  XOR U6387 ( .A(n2799), .B(n2800), .Z(n2798) );
  XOR U6388 ( .A(DB[2586]), .B(DB[2571]), .Z(n2800) );
  AND U6389 ( .A(n338), .B(n2801), .Z(n2799) );
  XOR U6390 ( .A(n2802), .B(n2803), .Z(n2801) );
  XOR U6391 ( .A(DB[2571]), .B(DB[2556]), .Z(n2803) );
  AND U6392 ( .A(n342), .B(n2804), .Z(n2802) );
  XOR U6393 ( .A(n2805), .B(n2806), .Z(n2804) );
  XOR U6394 ( .A(DB[2556]), .B(DB[2541]), .Z(n2806) );
  AND U6395 ( .A(n346), .B(n2807), .Z(n2805) );
  XOR U6396 ( .A(n2808), .B(n2809), .Z(n2807) );
  XOR U6397 ( .A(DB[2541]), .B(DB[2526]), .Z(n2809) );
  AND U6398 ( .A(n350), .B(n2810), .Z(n2808) );
  XOR U6399 ( .A(n2811), .B(n2812), .Z(n2810) );
  XOR U6400 ( .A(DB[2526]), .B(DB[2511]), .Z(n2812) );
  AND U6401 ( .A(n354), .B(n2813), .Z(n2811) );
  XOR U6402 ( .A(n2814), .B(n2815), .Z(n2813) );
  XOR U6403 ( .A(DB[2511]), .B(DB[2496]), .Z(n2815) );
  AND U6404 ( .A(n358), .B(n2816), .Z(n2814) );
  XOR U6405 ( .A(n2817), .B(n2818), .Z(n2816) );
  XOR U6406 ( .A(DB[2496]), .B(DB[2481]), .Z(n2818) );
  AND U6407 ( .A(n362), .B(n2819), .Z(n2817) );
  XOR U6408 ( .A(n2820), .B(n2821), .Z(n2819) );
  XOR U6409 ( .A(DB[2481]), .B(DB[2466]), .Z(n2821) );
  AND U6410 ( .A(n366), .B(n2822), .Z(n2820) );
  XOR U6411 ( .A(n2823), .B(n2824), .Z(n2822) );
  XOR U6412 ( .A(DB[2466]), .B(DB[2451]), .Z(n2824) );
  AND U6413 ( .A(n370), .B(n2825), .Z(n2823) );
  XOR U6414 ( .A(n2826), .B(n2827), .Z(n2825) );
  XOR U6415 ( .A(DB[2451]), .B(DB[2436]), .Z(n2827) );
  AND U6416 ( .A(n374), .B(n2828), .Z(n2826) );
  XOR U6417 ( .A(n2829), .B(n2830), .Z(n2828) );
  XOR U6418 ( .A(DB[2436]), .B(DB[2421]), .Z(n2830) );
  AND U6419 ( .A(n378), .B(n2831), .Z(n2829) );
  XOR U6420 ( .A(n2832), .B(n2833), .Z(n2831) );
  XOR U6421 ( .A(DB[2421]), .B(DB[2406]), .Z(n2833) );
  AND U6422 ( .A(n382), .B(n2834), .Z(n2832) );
  XOR U6423 ( .A(n2835), .B(n2836), .Z(n2834) );
  XOR U6424 ( .A(DB[2406]), .B(DB[2391]), .Z(n2836) );
  AND U6425 ( .A(n386), .B(n2837), .Z(n2835) );
  XOR U6426 ( .A(n2838), .B(n2839), .Z(n2837) );
  XOR U6427 ( .A(DB[2391]), .B(DB[2376]), .Z(n2839) );
  AND U6428 ( .A(n390), .B(n2840), .Z(n2838) );
  XOR U6429 ( .A(n2841), .B(n2842), .Z(n2840) );
  XOR U6430 ( .A(DB[2376]), .B(DB[2361]), .Z(n2842) );
  AND U6431 ( .A(n394), .B(n2843), .Z(n2841) );
  XOR U6432 ( .A(n2844), .B(n2845), .Z(n2843) );
  XOR U6433 ( .A(DB[2361]), .B(DB[2346]), .Z(n2845) );
  AND U6434 ( .A(n398), .B(n2846), .Z(n2844) );
  XOR U6435 ( .A(n2847), .B(n2848), .Z(n2846) );
  XOR U6436 ( .A(DB[2346]), .B(DB[2331]), .Z(n2848) );
  AND U6437 ( .A(n402), .B(n2849), .Z(n2847) );
  XOR U6438 ( .A(n2850), .B(n2851), .Z(n2849) );
  XOR U6439 ( .A(DB[2331]), .B(DB[2316]), .Z(n2851) );
  AND U6440 ( .A(n406), .B(n2852), .Z(n2850) );
  XOR U6441 ( .A(n2853), .B(n2854), .Z(n2852) );
  XOR U6442 ( .A(DB[2316]), .B(DB[2301]), .Z(n2854) );
  AND U6443 ( .A(n410), .B(n2855), .Z(n2853) );
  XOR U6444 ( .A(n2856), .B(n2857), .Z(n2855) );
  XOR U6445 ( .A(DB[2301]), .B(DB[2286]), .Z(n2857) );
  AND U6446 ( .A(n414), .B(n2858), .Z(n2856) );
  XOR U6447 ( .A(n2859), .B(n2860), .Z(n2858) );
  XOR U6448 ( .A(DB[2286]), .B(DB[2271]), .Z(n2860) );
  AND U6449 ( .A(n418), .B(n2861), .Z(n2859) );
  XOR U6450 ( .A(n2862), .B(n2863), .Z(n2861) );
  XOR U6451 ( .A(DB[2271]), .B(DB[2256]), .Z(n2863) );
  AND U6452 ( .A(n422), .B(n2864), .Z(n2862) );
  XOR U6453 ( .A(n2865), .B(n2866), .Z(n2864) );
  XOR U6454 ( .A(DB[2256]), .B(DB[2241]), .Z(n2866) );
  AND U6455 ( .A(n426), .B(n2867), .Z(n2865) );
  XOR U6456 ( .A(n2868), .B(n2869), .Z(n2867) );
  XOR U6457 ( .A(DB[2241]), .B(DB[2226]), .Z(n2869) );
  AND U6458 ( .A(n430), .B(n2870), .Z(n2868) );
  XOR U6459 ( .A(n2871), .B(n2872), .Z(n2870) );
  XOR U6460 ( .A(DB[2226]), .B(DB[2211]), .Z(n2872) );
  AND U6461 ( .A(n434), .B(n2873), .Z(n2871) );
  XOR U6462 ( .A(n2874), .B(n2875), .Z(n2873) );
  XOR U6463 ( .A(DB[2211]), .B(DB[2196]), .Z(n2875) );
  AND U6464 ( .A(n438), .B(n2876), .Z(n2874) );
  XOR U6465 ( .A(n2877), .B(n2878), .Z(n2876) );
  XOR U6466 ( .A(DB[2196]), .B(DB[2181]), .Z(n2878) );
  AND U6467 ( .A(n442), .B(n2879), .Z(n2877) );
  XOR U6468 ( .A(n2880), .B(n2881), .Z(n2879) );
  XOR U6469 ( .A(DB[2181]), .B(DB[2166]), .Z(n2881) );
  AND U6470 ( .A(n446), .B(n2882), .Z(n2880) );
  XOR U6471 ( .A(n2883), .B(n2884), .Z(n2882) );
  XOR U6472 ( .A(DB[2166]), .B(DB[2151]), .Z(n2884) );
  AND U6473 ( .A(n450), .B(n2885), .Z(n2883) );
  XOR U6474 ( .A(n2886), .B(n2887), .Z(n2885) );
  XOR U6475 ( .A(DB[2151]), .B(DB[2136]), .Z(n2887) );
  AND U6476 ( .A(n454), .B(n2888), .Z(n2886) );
  XOR U6477 ( .A(n2889), .B(n2890), .Z(n2888) );
  XOR U6478 ( .A(DB[2136]), .B(DB[2121]), .Z(n2890) );
  AND U6479 ( .A(n458), .B(n2891), .Z(n2889) );
  XOR U6480 ( .A(n2892), .B(n2893), .Z(n2891) );
  XOR U6481 ( .A(DB[2121]), .B(DB[2106]), .Z(n2893) );
  AND U6482 ( .A(n462), .B(n2894), .Z(n2892) );
  XOR U6483 ( .A(n2895), .B(n2896), .Z(n2894) );
  XOR U6484 ( .A(DB[2106]), .B(DB[2091]), .Z(n2896) );
  AND U6485 ( .A(n466), .B(n2897), .Z(n2895) );
  XOR U6486 ( .A(n2898), .B(n2899), .Z(n2897) );
  XOR U6487 ( .A(DB[2091]), .B(DB[2076]), .Z(n2899) );
  AND U6488 ( .A(n470), .B(n2900), .Z(n2898) );
  XOR U6489 ( .A(n2901), .B(n2902), .Z(n2900) );
  XOR U6490 ( .A(DB[2076]), .B(DB[2061]), .Z(n2902) );
  AND U6491 ( .A(n474), .B(n2903), .Z(n2901) );
  XOR U6492 ( .A(n2904), .B(n2905), .Z(n2903) );
  XOR U6493 ( .A(DB[2061]), .B(DB[2046]), .Z(n2905) );
  AND U6494 ( .A(n478), .B(n2906), .Z(n2904) );
  XOR U6495 ( .A(n2907), .B(n2908), .Z(n2906) );
  XOR U6496 ( .A(DB[2046]), .B(DB[2031]), .Z(n2908) );
  AND U6497 ( .A(n482), .B(n2909), .Z(n2907) );
  XOR U6498 ( .A(n2910), .B(n2911), .Z(n2909) );
  XOR U6499 ( .A(DB[2031]), .B(DB[2016]), .Z(n2911) );
  AND U6500 ( .A(n486), .B(n2912), .Z(n2910) );
  XOR U6501 ( .A(n2913), .B(n2914), .Z(n2912) );
  XOR U6502 ( .A(DB[2016]), .B(DB[2001]), .Z(n2914) );
  AND U6503 ( .A(n490), .B(n2915), .Z(n2913) );
  XOR U6504 ( .A(n2916), .B(n2917), .Z(n2915) );
  XOR U6505 ( .A(DB[2001]), .B(DB[1986]), .Z(n2917) );
  AND U6506 ( .A(n494), .B(n2918), .Z(n2916) );
  XOR U6507 ( .A(n2919), .B(n2920), .Z(n2918) );
  XOR U6508 ( .A(DB[1986]), .B(DB[1971]), .Z(n2920) );
  AND U6509 ( .A(n498), .B(n2921), .Z(n2919) );
  XOR U6510 ( .A(n2922), .B(n2923), .Z(n2921) );
  XOR U6511 ( .A(DB[1971]), .B(DB[1956]), .Z(n2923) );
  AND U6512 ( .A(n502), .B(n2924), .Z(n2922) );
  XOR U6513 ( .A(n2925), .B(n2926), .Z(n2924) );
  XOR U6514 ( .A(DB[1956]), .B(DB[1941]), .Z(n2926) );
  AND U6515 ( .A(n506), .B(n2927), .Z(n2925) );
  XOR U6516 ( .A(n2928), .B(n2929), .Z(n2927) );
  XOR U6517 ( .A(DB[1941]), .B(DB[1926]), .Z(n2929) );
  AND U6518 ( .A(n510), .B(n2930), .Z(n2928) );
  XOR U6519 ( .A(n2931), .B(n2932), .Z(n2930) );
  XOR U6520 ( .A(DB[1926]), .B(DB[1911]), .Z(n2932) );
  AND U6521 ( .A(n514), .B(n2933), .Z(n2931) );
  XOR U6522 ( .A(n2934), .B(n2935), .Z(n2933) );
  XOR U6523 ( .A(DB[1911]), .B(DB[1896]), .Z(n2935) );
  AND U6524 ( .A(n518), .B(n2936), .Z(n2934) );
  XOR U6525 ( .A(n2937), .B(n2938), .Z(n2936) );
  XOR U6526 ( .A(DB[1896]), .B(DB[1881]), .Z(n2938) );
  AND U6527 ( .A(n522), .B(n2939), .Z(n2937) );
  XOR U6528 ( .A(n2940), .B(n2941), .Z(n2939) );
  XOR U6529 ( .A(DB[1881]), .B(DB[1866]), .Z(n2941) );
  AND U6530 ( .A(n526), .B(n2942), .Z(n2940) );
  XOR U6531 ( .A(n2943), .B(n2944), .Z(n2942) );
  XOR U6532 ( .A(DB[1866]), .B(DB[1851]), .Z(n2944) );
  AND U6533 ( .A(n530), .B(n2945), .Z(n2943) );
  XOR U6534 ( .A(n2946), .B(n2947), .Z(n2945) );
  XOR U6535 ( .A(DB[1851]), .B(DB[1836]), .Z(n2947) );
  AND U6536 ( .A(n534), .B(n2948), .Z(n2946) );
  XOR U6537 ( .A(n2949), .B(n2950), .Z(n2948) );
  XOR U6538 ( .A(DB[1836]), .B(DB[1821]), .Z(n2950) );
  AND U6539 ( .A(n538), .B(n2951), .Z(n2949) );
  XOR U6540 ( .A(n2952), .B(n2953), .Z(n2951) );
  XOR U6541 ( .A(DB[1821]), .B(DB[1806]), .Z(n2953) );
  AND U6542 ( .A(n542), .B(n2954), .Z(n2952) );
  XOR U6543 ( .A(n2955), .B(n2956), .Z(n2954) );
  XOR U6544 ( .A(DB[1806]), .B(DB[1791]), .Z(n2956) );
  AND U6545 ( .A(n546), .B(n2957), .Z(n2955) );
  XOR U6546 ( .A(n2958), .B(n2959), .Z(n2957) );
  XOR U6547 ( .A(DB[1791]), .B(DB[1776]), .Z(n2959) );
  AND U6548 ( .A(n550), .B(n2960), .Z(n2958) );
  XOR U6549 ( .A(n2961), .B(n2962), .Z(n2960) );
  XOR U6550 ( .A(DB[1776]), .B(DB[1761]), .Z(n2962) );
  AND U6551 ( .A(n554), .B(n2963), .Z(n2961) );
  XOR U6552 ( .A(n2964), .B(n2965), .Z(n2963) );
  XOR U6553 ( .A(DB[1761]), .B(DB[1746]), .Z(n2965) );
  AND U6554 ( .A(n558), .B(n2966), .Z(n2964) );
  XOR U6555 ( .A(n2967), .B(n2968), .Z(n2966) );
  XOR U6556 ( .A(DB[1746]), .B(DB[1731]), .Z(n2968) );
  AND U6557 ( .A(n562), .B(n2969), .Z(n2967) );
  XOR U6558 ( .A(n2970), .B(n2971), .Z(n2969) );
  XOR U6559 ( .A(DB[1731]), .B(DB[1716]), .Z(n2971) );
  AND U6560 ( .A(n566), .B(n2972), .Z(n2970) );
  XOR U6561 ( .A(n2973), .B(n2974), .Z(n2972) );
  XOR U6562 ( .A(DB[1716]), .B(DB[1701]), .Z(n2974) );
  AND U6563 ( .A(n570), .B(n2975), .Z(n2973) );
  XOR U6564 ( .A(n2976), .B(n2977), .Z(n2975) );
  XOR U6565 ( .A(DB[1701]), .B(DB[1686]), .Z(n2977) );
  AND U6566 ( .A(n574), .B(n2978), .Z(n2976) );
  XOR U6567 ( .A(n2979), .B(n2980), .Z(n2978) );
  XOR U6568 ( .A(DB[1686]), .B(DB[1671]), .Z(n2980) );
  AND U6569 ( .A(n578), .B(n2981), .Z(n2979) );
  XOR U6570 ( .A(n2982), .B(n2983), .Z(n2981) );
  XOR U6571 ( .A(DB[1671]), .B(DB[1656]), .Z(n2983) );
  AND U6572 ( .A(n582), .B(n2984), .Z(n2982) );
  XOR U6573 ( .A(n2985), .B(n2986), .Z(n2984) );
  XOR U6574 ( .A(DB[1656]), .B(DB[1641]), .Z(n2986) );
  AND U6575 ( .A(n586), .B(n2987), .Z(n2985) );
  XOR U6576 ( .A(n2988), .B(n2989), .Z(n2987) );
  XOR U6577 ( .A(DB[1641]), .B(DB[1626]), .Z(n2989) );
  AND U6578 ( .A(n590), .B(n2990), .Z(n2988) );
  XOR U6579 ( .A(n2991), .B(n2992), .Z(n2990) );
  XOR U6580 ( .A(DB[1626]), .B(DB[1611]), .Z(n2992) );
  AND U6581 ( .A(n594), .B(n2993), .Z(n2991) );
  XOR U6582 ( .A(n2994), .B(n2995), .Z(n2993) );
  XOR U6583 ( .A(DB[1611]), .B(DB[1596]), .Z(n2995) );
  AND U6584 ( .A(n598), .B(n2996), .Z(n2994) );
  XOR U6585 ( .A(n2997), .B(n2998), .Z(n2996) );
  XOR U6586 ( .A(DB[1596]), .B(DB[1581]), .Z(n2998) );
  AND U6587 ( .A(n602), .B(n2999), .Z(n2997) );
  XOR U6588 ( .A(n3000), .B(n3001), .Z(n2999) );
  XOR U6589 ( .A(DB[1581]), .B(DB[1566]), .Z(n3001) );
  AND U6590 ( .A(n606), .B(n3002), .Z(n3000) );
  XOR U6591 ( .A(n3003), .B(n3004), .Z(n3002) );
  XOR U6592 ( .A(DB[1566]), .B(DB[1551]), .Z(n3004) );
  AND U6593 ( .A(n610), .B(n3005), .Z(n3003) );
  XOR U6594 ( .A(n3006), .B(n3007), .Z(n3005) );
  XOR U6595 ( .A(DB[1551]), .B(DB[1536]), .Z(n3007) );
  AND U6596 ( .A(n614), .B(n3008), .Z(n3006) );
  XOR U6597 ( .A(n3009), .B(n3010), .Z(n3008) );
  XOR U6598 ( .A(DB[1536]), .B(DB[1521]), .Z(n3010) );
  AND U6599 ( .A(n618), .B(n3011), .Z(n3009) );
  XOR U6600 ( .A(n3012), .B(n3013), .Z(n3011) );
  XOR U6601 ( .A(DB[1521]), .B(DB[1506]), .Z(n3013) );
  AND U6602 ( .A(n622), .B(n3014), .Z(n3012) );
  XOR U6603 ( .A(n3015), .B(n3016), .Z(n3014) );
  XOR U6604 ( .A(DB[1506]), .B(DB[1491]), .Z(n3016) );
  AND U6605 ( .A(n626), .B(n3017), .Z(n3015) );
  XOR U6606 ( .A(n3018), .B(n3019), .Z(n3017) );
  XOR U6607 ( .A(DB[1491]), .B(DB[1476]), .Z(n3019) );
  AND U6608 ( .A(n630), .B(n3020), .Z(n3018) );
  XOR U6609 ( .A(n3021), .B(n3022), .Z(n3020) );
  XOR U6610 ( .A(DB[1476]), .B(DB[1461]), .Z(n3022) );
  AND U6611 ( .A(n634), .B(n3023), .Z(n3021) );
  XOR U6612 ( .A(n3024), .B(n3025), .Z(n3023) );
  XOR U6613 ( .A(DB[1461]), .B(DB[1446]), .Z(n3025) );
  AND U6614 ( .A(n638), .B(n3026), .Z(n3024) );
  XOR U6615 ( .A(n3027), .B(n3028), .Z(n3026) );
  XOR U6616 ( .A(DB[1446]), .B(DB[1431]), .Z(n3028) );
  AND U6617 ( .A(n642), .B(n3029), .Z(n3027) );
  XOR U6618 ( .A(n3030), .B(n3031), .Z(n3029) );
  XOR U6619 ( .A(DB[1431]), .B(DB[1416]), .Z(n3031) );
  AND U6620 ( .A(n646), .B(n3032), .Z(n3030) );
  XOR U6621 ( .A(n3033), .B(n3034), .Z(n3032) );
  XOR U6622 ( .A(DB[1416]), .B(DB[1401]), .Z(n3034) );
  AND U6623 ( .A(n650), .B(n3035), .Z(n3033) );
  XOR U6624 ( .A(n3036), .B(n3037), .Z(n3035) );
  XOR U6625 ( .A(DB[1401]), .B(DB[1386]), .Z(n3037) );
  AND U6626 ( .A(n654), .B(n3038), .Z(n3036) );
  XOR U6627 ( .A(n3039), .B(n3040), .Z(n3038) );
  XOR U6628 ( .A(DB[1386]), .B(DB[1371]), .Z(n3040) );
  AND U6629 ( .A(n658), .B(n3041), .Z(n3039) );
  XOR U6630 ( .A(n3042), .B(n3043), .Z(n3041) );
  XOR U6631 ( .A(DB[1371]), .B(DB[1356]), .Z(n3043) );
  AND U6632 ( .A(n662), .B(n3044), .Z(n3042) );
  XOR U6633 ( .A(n3045), .B(n3046), .Z(n3044) );
  XOR U6634 ( .A(DB[1356]), .B(DB[1341]), .Z(n3046) );
  AND U6635 ( .A(n666), .B(n3047), .Z(n3045) );
  XOR U6636 ( .A(n3048), .B(n3049), .Z(n3047) );
  XOR U6637 ( .A(DB[1341]), .B(DB[1326]), .Z(n3049) );
  AND U6638 ( .A(n670), .B(n3050), .Z(n3048) );
  XOR U6639 ( .A(n3051), .B(n3052), .Z(n3050) );
  XOR U6640 ( .A(DB[1326]), .B(DB[1311]), .Z(n3052) );
  AND U6641 ( .A(n674), .B(n3053), .Z(n3051) );
  XOR U6642 ( .A(n3054), .B(n3055), .Z(n3053) );
  XOR U6643 ( .A(DB[1311]), .B(DB[1296]), .Z(n3055) );
  AND U6644 ( .A(n678), .B(n3056), .Z(n3054) );
  XOR U6645 ( .A(n3057), .B(n3058), .Z(n3056) );
  XOR U6646 ( .A(DB[1296]), .B(DB[1281]), .Z(n3058) );
  AND U6647 ( .A(n682), .B(n3059), .Z(n3057) );
  XOR U6648 ( .A(n3060), .B(n3061), .Z(n3059) );
  XOR U6649 ( .A(DB[1281]), .B(DB[1266]), .Z(n3061) );
  AND U6650 ( .A(n686), .B(n3062), .Z(n3060) );
  XOR U6651 ( .A(n3063), .B(n3064), .Z(n3062) );
  XOR U6652 ( .A(DB[1266]), .B(DB[1251]), .Z(n3064) );
  AND U6653 ( .A(n690), .B(n3065), .Z(n3063) );
  XOR U6654 ( .A(n3066), .B(n3067), .Z(n3065) );
  XOR U6655 ( .A(DB[1251]), .B(DB[1236]), .Z(n3067) );
  AND U6656 ( .A(n694), .B(n3068), .Z(n3066) );
  XOR U6657 ( .A(n3069), .B(n3070), .Z(n3068) );
  XOR U6658 ( .A(DB[1236]), .B(DB[1221]), .Z(n3070) );
  AND U6659 ( .A(n698), .B(n3071), .Z(n3069) );
  XOR U6660 ( .A(n3072), .B(n3073), .Z(n3071) );
  XOR U6661 ( .A(DB[1221]), .B(DB[1206]), .Z(n3073) );
  AND U6662 ( .A(n702), .B(n3074), .Z(n3072) );
  XOR U6663 ( .A(n3075), .B(n3076), .Z(n3074) );
  XOR U6664 ( .A(DB[1206]), .B(DB[1191]), .Z(n3076) );
  AND U6665 ( .A(n706), .B(n3077), .Z(n3075) );
  XOR U6666 ( .A(n3078), .B(n3079), .Z(n3077) );
  XOR U6667 ( .A(DB[1191]), .B(DB[1176]), .Z(n3079) );
  AND U6668 ( .A(n710), .B(n3080), .Z(n3078) );
  XOR U6669 ( .A(n3081), .B(n3082), .Z(n3080) );
  XOR U6670 ( .A(DB[1176]), .B(DB[1161]), .Z(n3082) );
  AND U6671 ( .A(n714), .B(n3083), .Z(n3081) );
  XOR U6672 ( .A(n3084), .B(n3085), .Z(n3083) );
  XOR U6673 ( .A(DB[1161]), .B(DB[1146]), .Z(n3085) );
  AND U6674 ( .A(n718), .B(n3086), .Z(n3084) );
  XOR U6675 ( .A(n3087), .B(n3088), .Z(n3086) );
  XOR U6676 ( .A(DB[1146]), .B(DB[1131]), .Z(n3088) );
  AND U6677 ( .A(n722), .B(n3089), .Z(n3087) );
  XOR U6678 ( .A(n3090), .B(n3091), .Z(n3089) );
  XOR U6679 ( .A(DB[1131]), .B(DB[1116]), .Z(n3091) );
  AND U6680 ( .A(n726), .B(n3092), .Z(n3090) );
  XOR U6681 ( .A(n3093), .B(n3094), .Z(n3092) );
  XOR U6682 ( .A(DB[1116]), .B(DB[1101]), .Z(n3094) );
  AND U6683 ( .A(n730), .B(n3095), .Z(n3093) );
  XOR U6684 ( .A(n3096), .B(n3097), .Z(n3095) );
  XOR U6685 ( .A(DB[1101]), .B(DB[1086]), .Z(n3097) );
  AND U6686 ( .A(n734), .B(n3098), .Z(n3096) );
  XOR U6687 ( .A(n3099), .B(n3100), .Z(n3098) );
  XOR U6688 ( .A(DB[1086]), .B(DB[1071]), .Z(n3100) );
  AND U6689 ( .A(n738), .B(n3101), .Z(n3099) );
  XOR U6690 ( .A(n3102), .B(n3103), .Z(n3101) );
  XOR U6691 ( .A(DB[1071]), .B(DB[1056]), .Z(n3103) );
  AND U6692 ( .A(n742), .B(n3104), .Z(n3102) );
  XOR U6693 ( .A(n3105), .B(n3106), .Z(n3104) );
  XOR U6694 ( .A(DB[1056]), .B(DB[1041]), .Z(n3106) );
  AND U6695 ( .A(n746), .B(n3107), .Z(n3105) );
  XOR U6696 ( .A(n3108), .B(n3109), .Z(n3107) );
  XOR U6697 ( .A(DB[1041]), .B(DB[1026]), .Z(n3109) );
  AND U6698 ( .A(n750), .B(n3110), .Z(n3108) );
  XOR U6699 ( .A(n3111), .B(n3112), .Z(n3110) );
  XOR U6700 ( .A(DB[1026]), .B(DB[1011]), .Z(n3112) );
  AND U6701 ( .A(n754), .B(n3113), .Z(n3111) );
  XOR U6702 ( .A(n3114), .B(n3115), .Z(n3113) );
  XOR U6703 ( .A(DB[996]), .B(DB[1011]), .Z(n3115) );
  AND U6704 ( .A(n758), .B(n3116), .Z(n3114) );
  XOR U6705 ( .A(n3117), .B(n3118), .Z(n3116) );
  XOR U6706 ( .A(DB[996]), .B(DB[981]), .Z(n3118) );
  AND U6707 ( .A(n762), .B(n3119), .Z(n3117) );
  XOR U6708 ( .A(n3120), .B(n3121), .Z(n3119) );
  XOR U6709 ( .A(DB[981]), .B(DB[966]), .Z(n3121) );
  AND U6710 ( .A(n766), .B(n3122), .Z(n3120) );
  XOR U6711 ( .A(n3123), .B(n3124), .Z(n3122) );
  XOR U6712 ( .A(DB[966]), .B(DB[951]), .Z(n3124) );
  AND U6713 ( .A(n770), .B(n3125), .Z(n3123) );
  XOR U6714 ( .A(n3126), .B(n3127), .Z(n3125) );
  XOR U6715 ( .A(DB[951]), .B(DB[936]), .Z(n3127) );
  AND U6716 ( .A(n774), .B(n3128), .Z(n3126) );
  XOR U6717 ( .A(n3129), .B(n3130), .Z(n3128) );
  XOR U6718 ( .A(DB[936]), .B(DB[921]), .Z(n3130) );
  AND U6719 ( .A(n778), .B(n3131), .Z(n3129) );
  XOR U6720 ( .A(n3132), .B(n3133), .Z(n3131) );
  XOR U6721 ( .A(DB[921]), .B(DB[906]), .Z(n3133) );
  AND U6722 ( .A(n782), .B(n3134), .Z(n3132) );
  XOR U6723 ( .A(n3135), .B(n3136), .Z(n3134) );
  XOR U6724 ( .A(DB[906]), .B(DB[891]), .Z(n3136) );
  AND U6725 ( .A(n786), .B(n3137), .Z(n3135) );
  XOR U6726 ( .A(n3138), .B(n3139), .Z(n3137) );
  XOR U6727 ( .A(DB[891]), .B(DB[876]), .Z(n3139) );
  AND U6728 ( .A(n790), .B(n3140), .Z(n3138) );
  XOR U6729 ( .A(n3141), .B(n3142), .Z(n3140) );
  XOR U6730 ( .A(DB[876]), .B(DB[861]), .Z(n3142) );
  AND U6731 ( .A(n794), .B(n3143), .Z(n3141) );
  XOR U6732 ( .A(n3144), .B(n3145), .Z(n3143) );
  XOR U6733 ( .A(DB[861]), .B(DB[846]), .Z(n3145) );
  AND U6734 ( .A(n798), .B(n3146), .Z(n3144) );
  XOR U6735 ( .A(n3147), .B(n3148), .Z(n3146) );
  XOR U6736 ( .A(DB[846]), .B(DB[831]), .Z(n3148) );
  AND U6737 ( .A(n802), .B(n3149), .Z(n3147) );
  XOR U6738 ( .A(n3150), .B(n3151), .Z(n3149) );
  XOR U6739 ( .A(DB[831]), .B(DB[816]), .Z(n3151) );
  AND U6740 ( .A(n806), .B(n3152), .Z(n3150) );
  XOR U6741 ( .A(n3153), .B(n3154), .Z(n3152) );
  XOR U6742 ( .A(DB[816]), .B(DB[801]), .Z(n3154) );
  AND U6743 ( .A(n810), .B(n3155), .Z(n3153) );
  XOR U6744 ( .A(n3156), .B(n3157), .Z(n3155) );
  XOR U6745 ( .A(DB[801]), .B(DB[786]), .Z(n3157) );
  AND U6746 ( .A(n814), .B(n3158), .Z(n3156) );
  XOR U6747 ( .A(n3159), .B(n3160), .Z(n3158) );
  XOR U6748 ( .A(DB[786]), .B(DB[771]), .Z(n3160) );
  AND U6749 ( .A(n818), .B(n3161), .Z(n3159) );
  XOR U6750 ( .A(n3162), .B(n3163), .Z(n3161) );
  XOR U6751 ( .A(DB[771]), .B(DB[756]), .Z(n3163) );
  AND U6752 ( .A(n822), .B(n3164), .Z(n3162) );
  XOR U6753 ( .A(n3165), .B(n3166), .Z(n3164) );
  XOR U6754 ( .A(DB[756]), .B(DB[741]), .Z(n3166) );
  AND U6755 ( .A(n826), .B(n3167), .Z(n3165) );
  XOR U6756 ( .A(n3168), .B(n3169), .Z(n3167) );
  XOR U6757 ( .A(DB[741]), .B(DB[726]), .Z(n3169) );
  AND U6758 ( .A(n830), .B(n3170), .Z(n3168) );
  XOR U6759 ( .A(n3171), .B(n3172), .Z(n3170) );
  XOR U6760 ( .A(DB[726]), .B(DB[711]), .Z(n3172) );
  AND U6761 ( .A(n834), .B(n3173), .Z(n3171) );
  XOR U6762 ( .A(n3174), .B(n3175), .Z(n3173) );
  XOR U6763 ( .A(DB[711]), .B(DB[696]), .Z(n3175) );
  AND U6764 ( .A(n838), .B(n3176), .Z(n3174) );
  XOR U6765 ( .A(n3177), .B(n3178), .Z(n3176) );
  XOR U6766 ( .A(DB[696]), .B(DB[681]), .Z(n3178) );
  AND U6767 ( .A(n842), .B(n3179), .Z(n3177) );
  XOR U6768 ( .A(n3180), .B(n3181), .Z(n3179) );
  XOR U6769 ( .A(DB[681]), .B(DB[666]), .Z(n3181) );
  AND U6770 ( .A(n846), .B(n3182), .Z(n3180) );
  XOR U6771 ( .A(n3183), .B(n3184), .Z(n3182) );
  XOR U6772 ( .A(DB[666]), .B(DB[651]), .Z(n3184) );
  AND U6773 ( .A(n850), .B(n3185), .Z(n3183) );
  XOR U6774 ( .A(n3186), .B(n3187), .Z(n3185) );
  XOR U6775 ( .A(DB[651]), .B(DB[636]), .Z(n3187) );
  AND U6776 ( .A(n854), .B(n3188), .Z(n3186) );
  XOR U6777 ( .A(n3189), .B(n3190), .Z(n3188) );
  XOR U6778 ( .A(DB[636]), .B(DB[621]), .Z(n3190) );
  AND U6779 ( .A(n858), .B(n3191), .Z(n3189) );
  XOR U6780 ( .A(n3192), .B(n3193), .Z(n3191) );
  XOR U6781 ( .A(DB[621]), .B(DB[606]), .Z(n3193) );
  AND U6782 ( .A(n862), .B(n3194), .Z(n3192) );
  XOR U6783 ( .A(n3195), .B(n3196), .Z(n3194) );
  XOR U6784 ( .A(DB[606]), .B(DB[591]), .Z(n3196) );
  AND U6785 ( .A(n866), .B(n3197), .Z(n3195) );
  XOR U6786 ( .A(n3198), .B(n3199), .Z(n3197) );
  XOR U6787 ( .A(DB[591]), .B(DB[576]), .Z(n3199) );
  AND U6788 ( .A(n870), .B(n3200), .Z(n3198) );
  XOR U6789 ( .A(n3201), .B(n3202), .Z(n3200) );
  XOR U6790 ( .A(DB[576]), .B(DB[561]), .Z(n3202) );
  AND U6791 ( .A(n874), .B(n3203), .Z(n3201) );
  XOR U6792 ( .A(n3204), .B(n3205), .Z(n3203) );
  XOR U6793 ( .A(DB[561]), .B(DB[546]), .Z(n3205) );
  AND U6794 ( .A(n878), .B(n3206), .Z(n3204) );
  XOR U6795 ( .A(n3207), .B(n3208), .Z(n3206) );
  XOR U6796 ( .A(DB[546]), .B(DB[531]), .Z(n3208) );
  AND U6797 ( .A(n882), .B(n3209), .Z(n3207) );
  XOR U6798 ( .A(n3210), .B(n3211), .Z(n3209) );
  XOR U6799 ( .A(DB[531]), .B(DB[516]), .Z(n3211) );
  AND U6800 ( .A(n886), .B(n3212), .Z(n3210) );
  XOR U6801 ( .A(n3213), .B(n3214), .Z(n3212) );
  XOR U6802 ( .A(DB[516]), .B(DB[501]), .Z(n3214) );
  AND U6803 ( .A(n890), .B(n3215), .Z(n3213) );
  XOR U6804 ( .A(n3216), .B(n3217), .Z(n3215) );
  XOR U6805 ( .A(DB[501]), .B(DB[486]), .Z(n3217) );
  AND U6806 ( .A(n894), .B(n3218), .Z(n3216) );
  XOR U6807 ( .A(n3219), .B(n3220), .Z(n3218) );
  XOR U6808 ( .A(DB[486]), .B(DB[471]), .Z(n3220) );
  AND U6809 ( .A(n898), .B(n3221), .Z(n3219) );
  XOR U6810 ( .A(n3222), .B(n3223), .Z(n3221) );
  XOR U6811 ( .A(DB[471]), .B(DB[456]), .Z(n3223) );
  AND U6812 ( .A(n902), .B(n3224), .Z(n3222) );
  XOR U6813 ( .A(n3225), .B(n3226), .Z(n3224) );
  XOR U6814 ( .A(DB[456]), .B(DB[441]), .Z(n3226) );
  AND U6815 ( .A(n906), .B(n3227), .Z(n3225) );
  XOR U6816 ( .A(n3228), .B(n3229), .Z(n3227) );
  XOR U6817 ( .A(DB[441]), .B(DB[426]), .Z(n3229) );
  AND U6818 ( .A(n910), .B(n3230), .Z(n3228) );
  XOR U6819 ( .A(n3231), .B(n3232), .Z(n3230) );
  XOR U6820 ( .A(DB[426]), .B(DB[411]), .Z(n3232) );
  AND U6821 ( .A(n914), .B(n3233), .Z(n3231) );
  XOR U6822 ( .A(n3234), .B(n3235), .Z(n3233) );
  XOR U6823 ( .A(DB[411]), .B(DB[396]), .Z(n3235) );
  AND U6824 ( .A(n918), .B(n3236), .Z(n3234) );
  XOR U6825 ( .A(n3237), .B(n3238), .Z(n3236) );
  XOR U6826 ( .A(DB[396]), .B(DB[381]), .Z(n3238) );
  AND U6827 ( .A(n922), .B(n3239), .Z(n3237) );
  XOR U6828 ( .A(n3240), .B(n3241), .Z(n3239) );
  XOR U6829 ( .A(DB[381]), .B(DB[366]), .Z(n3241) );
  AND U6830 ( .A(n926), .B(n3242), .Z(n3240) );
  XOR U6831 ( .A(n3243), .B(n3244), .Z(n3242) );
  XOR U6832 ( .A(DB[366]), .B(DB[351]), .Z(n3244) );
  AND U6833 ( .A(n930), .B(n3245), .Z(n3243) );
  XOR U6834 ( .A(n3246), .B(n3247), .Z(n3245) );
  XOR U6835 ( .A(DB[351]), .B(DB[336]), .Z(n3247) );
  AND U6836 ( .A(n934), .B(n3248), .Z(n3246) );
  XOR U6837 ( .A(n3249), .B(n3250), .Z(n3248) );
  XOR U6838 ( .A(DB[336]), .B(DB[321]), .Z(n3250) );
  AND U6839 ( .A(n938), .B(n3251), .Z(n3249) );
  XOR U6840 ( .A(n3252), .B(n3253), .Z(n3251) );
  XOR U6841 ( .A(DB[321]), .B(DB[306]), .Z(n3253) );
  AND U6842 ( .A(n942), .B(n3254), .Z(n3252) );
  XOR U6843 ( .A(n3255), .B(n3256), .Z(n3254) );
  XOR U6844 ( .A(DB[306]), .B(DB[291]), .Z(n3256) );
  AND U6845 ( .A(n946), .B(n3257), .Z(n3255) );
  XOR U6846 ( .A(n3258), .B(n3259), .Z(n3257) );
  XOR U6847 ( .A(DB[291]), .B(DB[276]), .Z(n3259) );
  AND U6848 ( .A(n950), .B(n3260), .Z(n3258) );
  XOR U6849 ( .A(n3261), .B(n3262), .Z(n3260) );
  XOR U6850 ( .A(DB[276]), .B(DB[261]), .Z(n3262) );
  AND U6851 ( .A(n954), .B(n3263), .Z(n3261) );
  XOR U6852 ( .A(n3264), .B(n3265), .Z(n3263) );
  XOR U6853 ( .A(DB[261]), .B(DB[246]), .Z(n3265) );
  AND U6854 ( .A(n958), .B(n3266), .Z(n3264) );
  XOR U6855 ( .A(n3267), .B(n3268), .Z(n3266) );
  XOR U6856 ( .A(DB[246]), .B(DB[231]), .Z(n3268) );
  AND U6857 ( .A(n962), .B(n3269), .Z(n3267) );
  XOR U6858 ( .A(n3270), .B(n3271), .Z(n3269) );
  XOR U6859 ( .A(DB[231]), .B(DB[216]), .Z(n3271) );
  AND U6860 ( .A(n966), .B(n3272), .Z(n3270) );
  XOR U6861 ( .A(n3273), .B(n3274), .Z(n3272) );
  XOR U6862 ( .A(DB[216]), .B(DB[201]), .Z(n3274) );
  AND U6863 ( .A(n970), .B(n3275), .Z(n3273) );
  XOR U6864 ( .A(n3276), .B(n3277), .Z(n3275) );
  XOR U6865 ( .A(DB[201]), .B(DB[186]), .Z(n3277) );
  AND U6866 ( .A(n974), .B(n3278), .Z(n3276) );
  XOR U6867 ( .A(n3279), .B(n3280), .Z(n3278) );
  XOR U6868 ( .A(DB[186]), .B(DB[171]), .Z(n3280) );
  AND U6869 ( .A(n978), .B(n3281), .Z(n3279) );
  XOR U6870 ( .A(n3282), .B(n3283), .Z(n3281) );
  XOR U6871 ( .A(DB[171]), .B(DB[156]), .Z(n3283) );
  AND U6872 ( .A(n982), .B(n3284), .Z(n3282) );
  XOR U6873 ( .A(n3285), .B(n3286), .Z(n3284) );
  XOR U6874 ( .A(DB[156]), .B(DB[141]), .Z(n3286) );
  AND U6875 ( .A(n986), .B(n3287), .Z(n3285) );
  XOR U6876 ( .A(n3288), .B(n3289), .Z(n3287) );
  XOR U6877 ( .A(DB[141]), .B(DB[126]), .Z(n3289) );
  AND U6878 ( .A(n990), .B(n3290), .Z(n3288) );
  XOR U6879 ( .A(n3291), .B(n3292), .Z(n3290) );
  XOR U6880 ( .A(DB[126]), .B(DB[111]), .Z(n3292) );
  AND U6881 ( .A(n994), .B(n3293), .Z(n3291) );
  XOR U6882 ( .A(n3294), .B(n3295), .Z(n3293) );
  XOR U6883 ( .A(DB[96]), .B(DB[111]), .Z(n3295) );
  AND U6884 ( .A(n998), .B(n3296), .Z(n3294) );
  XOR U6885 ( .A(n3297), .B(n3298), .Z(n3296) );
  XOR U6886 ( .A(DB[96]), .B(DB[81]), .Z(n3298) );
  AND U6887 ( .A(n1002), .B(n3299), .Z(n3297) );
  XOR U6888 ( .A(n3300), .B(n3301), .Z(n3299) );
  XOR U6889 ( .A(DB[81]), .B(DB[66]), .Z(n3301) );
  AND U6890 ( .A(n1006), .B(n3302), .Z(n3300) );
  XOR U6891 ( .A(n3303), .B(n3304), .Z(n3302) );
  XOR U6892 ( .A(DB[66]), .B(DB[51]), .Z(n3304) );
  AND U6893 ( .A(n1010), .B(n3305), .Z(n3303) );
  XOR U6894 ( .A(n3306), .B(n3307), .Z(n3305) );
  XOR U6895 ( .A(DB[51]), .B(DB[36]), .Z(n3307) );
  AND U6896 ( .A(n1014), .B(n3308), .Z(n3306) );
  XOR U6897 ( .A(n3309), .B(n3310), .Z(n3308) );
  XOR U6898 ( .A(DB[36]), .B(DB[21]), .Z(n3310) );
  AND U6899 ( .A(n1018), .B(n3311), .Z(n3309) );
  XOR U6900 ( .A(DB[6]), .B(DB[21]), .Z(n3311) );
  XOR U6901 ( .A(DB[3830]), .B(n3312), .Z(min_val_out[5]) );
  AND U6902 ( .A(n2), .B(n3313), .Z(n3312) );
  XOR U6903 ( .A(n3314), .B(n3315), .Z(n3313) );
  XOR U6904 ( .A(DB[3830]), .B(DB[3815]), .Z(n3315) );
  AND U6905 ( .A(n6), .B(n3316), .Z(n3314) );
  XOR U6906 ( .A(n3317), .B(n3318), .Z(n3316) );
  XOR U6907 ( .A(DB[3815]), .B(DB[3800]), .Z(n3318) );
  AND U6908 ( .A(n10), .B(n3319), .Z(n3317) );
  XOR U6909 ( .A(n3320), .B(n3321), .Z(n3319) );
  XOR U6910 ( .A(DB[3800]), .B(DB[3785]), .Z(n3321) );
  AND U6911 ( .A(n14), .B(n3322), .Z(n3320) );
  XOR U6912 ( .A(n3323), .B(n3324), .Z(n3322) );
  XOR U6913 ( .A(DB[3785]), .B(DB[3770]), .Z(n3324) );
  AND U6914 ( .A(n18), .B(n3325), .Z(n3323) );
  XOR U6915 ( .A(n3326), .B(n3327), .Z(n3325) );
  XOR U6916 ( .A(DB[3770]), .B(DB[3755]), .Z(n3327) );
  AND U6917 ( .A(n22), .B(n3328), .Z(n3326) );
  XOR U6918 ( .A(n3329), .B(n3330), .Z(n3328) );
  XOR U6919 ( .A(DB[3755]), .B(DB[3740]), .Z(n3330) );
  AND U6920 ( .A(n26), .B(n3331), .Z(n3329) );
  XOR U6921 ( .A(n3332), .B(n3333), .Z(n3331) );
  XOR U6922 ( .A(DB[3740]), .B(DB[3725]), .Z(n3333) );
  AND U6923 ( .A(n30), .B(n3334), .Z(n3332) );
  XOR U6924 ( .A(n3335), .B(n3336), .Z(n3334) );
  XOR U6925 ( .A(DB[3725]), .B(DB[3710]), .Z(n3336) );
  AND U6926 ( .A(n34), .B(n3337), .Z(n3335) );
  XOR U6927 ( .A(n3338), .B(n3339), .Z(n3337) );
  XOR U6928 ( .A(DB[3710]), .B(DB[3695]), .Z(n3339) );
  AND U6929 ( .A(n38), .B(n3340), .Z(n3338) );
  XOR U6930 ( .A(n3341), .B(n3342), .Z(n3340) );
  XOR U6931 ( .A(DB[3695]), .B(DB[3680]), .Z(n3342) );
  AND U6932 ( .A(n42), .B(n3343), .Z(n3341) );
  XOR U6933 ( .A(n3344), .B(n3345), .Z(n3343) );
  XOR U6934 ( .A(DB[3680]), .B(DB[3665]), .Z(n3345) );
  AND U6935 ( .A(n46), .B(n3346), .Z(n3344) );
  XOR U6936 ( .A(n3347), .B(n3348), .Z(n3346) );
  XOR U6937 ( .A(DB[3665]), .B(DB[3650]), .Z(n3348) );
  AND U6938 ( .A(n50), .B(n3349), .Z(n3347) );
  XOR U6939 ( .A(n3350), .B(n3351), .Z(n3349) );
  XOR U6940 ( .A(DB[3650]), .B(DB[3635]), .Z(n3351) );
  AND U6941 ( .A(n54), .B(n3352), .Z(n3350) );
  XOR U6942 ( .A(n3353), .B(n3354), .Z(n3352) );
  XOR U6943 ( .A(DB[3635]), .B(DB[3620]), .Z(n3354) );
  AND U6944 ( .A(n58), .B(n3355), .Z(n3353) );
  XOR U6945 ( .A(n3356), .B(n3357), .Z(n3355) );
  XOR U6946 ( .A(DB[3620]), .B(DB[3605]), .Z(n3357) );
  AND U6947 ( .A(n62), .B(n3358), .Z(n3356) );
  XOR U6948 ( .A(n3359), .B(n3360), .Z(n3358) );
  XOR U6949 ( .A(DB[3605]), .B(DB[3590]), .Z(n3360) );
  AND U6950 ( .A(n66), .B(n3361), .Z(n3359) );
  XOR U6951 ( .A(n3362), .B(n3363), .Z(n3361) );
  XOR U6952 ( .A(DB[3590]), .B(DB[3575]), .Z(n3363) );
  AND U6953 ( .A(n70), .B(n3364), .Z(n3362) );
  XOR U6954 ( .A(n3365), .B(n3366), .Z(n3364) );
  XOR U6955 ( .A(DB[3575]), .B(DB[3560]), .Z(n3366) );
  AND U6956 ( .A(n74), .B(n3367), .Z(n3365) );
  XOR U6957 ( .A(n3368), .B(n3369), .Z(n3367) );
  XOR U6958 ( .A(DB[3560]), .B(DB[3545]), .Z(n3369) );
  AND U6959 ( .A(n78), .B(n3370), .Z(n3368) );
  XOR U6960 ( .A(n3371), .B(n3372), .Z(n3370) );
  XOR U6961 ( .A(DB[3545]), .B(DB[3530]), .Z(n3372) );
  AND U6962 ( .A(n82), .B(n3373), .Z(n3371) );
  XOR U6963 ( .A(n3374), .B(n3375), .Z(n3373) );
  XOR U6964 ( .A(DB[3530]), .B(DB[3515]), .Z(n3375) );
  AND U6965 ( .A(n86), .B(n3376), .Z(n3374) );
  XOR U6966 ( .A(n3377), .B(n3378), .Z(n3376) );
  XOR U6967 ( .A(DB[3515]), .B(DB[3500]), .Z(n3378) );
  AND U6968 ( .A(n90), .B(n3379), .Z(n3377) );
  XOR U6969 ( .A(n3380), .B(n3381), .Z(n3379) );
  XOR U6970 ( .A(DB[3500]), .B(DB[3485]), .Z(n3381) );
  AND U6971 ( .A(n94), .B(n3382), .Z(n3380) );
  XOR U6972 ( .A(n3383), .B(n3384), .Z(n3382) );
  XOR U6973 ( .A(DB[3485]), .B(DB[3470]), .Z(n3384) );
  AND U6974 ( .A(n98), .B(n3385), .Z(n3383) );
  XOR U6975 ( .A(n3386), .B(n3387), .Z(n3385) );
  XOR U6976 ( .A(DB[3470]), .B(DB[3455]), .Z(n3387) );
  AND U6977 ( .A(n102), .B(n3388), .Z(n3386) );
  XOR U6978 ( .A(n3389), .B(n3390), .Z(n3388) );
  XOR U6979 ( .A(DB[3455]), .B(DB[3440]), .Z(n3390) );
  AND U6980 ( .A(n106), .B(n3391), .Z(n3389) );
  XOR U6981 ( .A(n3392), .B(n3393), .Z(n3391) );
  XOR U6982 ( .A(DB[3440]), .B(DB[3425]), .Z(n3393) );
  AND U6983 ( .A(n110), .B(n3394), .Z(n3392) );
  XOR U6984 ( .A(n3395), .B(n3396), .Z(n3394) );
  XOR U6985 ( .A(DB[3425]), .B(DB[3410]), .Z(n3396) );
  AND U6986 ( .A(n114), .B(n3397), .Z(n3395) );
  XOR U6987 ( .A(n3398), .B(n3399), .Z(n3397) );
  XOR U6988 ( .A(DB[3410]), .B(DB[3395]), .Z(n3399) );
  AND U6989 ( .A(n118), .B(n3400), .Z(n3398) );
  XOR U6990 ( .A(n3401), .B(n3402), .Z(n3400) );
  XOR U6991 ( .A(DB[3395]), .B(DB[3380]), .Z(n3402) );
  AND U6992 ( .A(n122), .B(n3403), .Z(n3401) );
  XOR U6993 ( .A(n3404), .B(n3405), .Z(n3403) );
  XOR U6994 ( .A(DB[3380]), .B(DB[3365]), .Z(n3405) );
  AND U6995 ( .A(n126), .B(n3406), .Z(n3404) );
  XOR U6996 ( .A(n3407), .B(n3408), .Z(n3406) );
  XOR U6997 ( .A(DB[3365]), .B(DB[3350]), .Z(n3408) );
  AND U6998 ( .A(n130), .B(n3409), .Z(n3407) );
  XOR U6999 ( .A(n3410), .B(n3411), .Z(n3409) );
  XOR U7000 ( .A(DB[3350]), .B(DB[3335]), .Z(n3411) );
  AND U7001 ( .A(n134), .B(n3412), .Z(n3410) );
  XOR U7002 ( .A(n3413), .B(n3414), .Z(n3412) );
  XOR U7003 ( .A(DB[3335]), .B(DB[3320]), .Z(n3414) );
  AND U7004 ( .A(n138), .B(n3415), .Z(n3413) );
  XOR U7005 ( .A(n3416), .B(n3417), .Z(n3415) );
  XOR U7006 ( .A(DB[3320]), .B(DB[3305]), .Z(n3417) );
  AND U7007 ( .A(n142), .B(n3418), .Z(n3416) );
  XOR U7008 ( .A(n3419), .B(n3420), .Z(n3418) );
  XOR U7009 ( .A(DB[3305]), .B(DB[3290]), .Z(n3420) );
  AND U7010 ( .A(n146), .B(n3421), .Z(n3419) );
  XOR U7011 ( .A(n3422), .B(n3423), .Z(n3421) );
  XOR U7012 ( .A(DB[3290]), .B(DB[3275]), .Z(n3423) );
  AND U7013 ( .A(n150), .B(n3424), .Z(n3422) );
  XOR U7014 ( .A(n3425), .B(n3426), .Z(n3424) );
  XOR U7015 ( .A(DB[3275]), .B(DB[3260]), .Z(n3426) );
  AND U7016 ( .A(n154), .B(n3427), .Z(n3425) );
  XOR U7017 ( .A(n3428), .B(n3429), .Z(n3427) );
  XOR U7018 ( .A(DB[3260]), .B(DB[3245]), .Z(n3429) );
  AND U7019 ( .A(n158), .B(n3430), .Z(n3428) );
  XOR U7020 ( .A(n3431), .B(n3432), .Z(n3430) );
  XOR U7021 ( .A(DB[3245]), .B(DB[3230]), .Z(n3432) );
  AND U7022 ( .A(n162), .B(n3433), .Z(n3431) );
  XOR U7023 ( .A(n3434), .B(n3435), .Z(n3433) );
  XOR U7024 ( .A(DB[3230]), .B(DB[3215]), .Z(n3435) );
  AND U7025 ( .A(n166), .B(n3436), .Z(n3434) );
  XOR U7026 ( .A(n3437), .B(n3438), .Z(n3436) );
  XOR U7027 ( .A(DB[3215]), .B(DB[3200]), .Z(n3438) );
  AND U7028 ( .A(n170), .B(n3439), .Z(n3437) );
  XOR U7029 ( .A(n3440), .B(n3441), .Z(n3439) );
  XOR U7030 ( .A(DB[3200]), .B(DB[3185]), .Z(n3441) );
  AND U7031 ( .A(n174), .B(n3442), .Z(n3440) );
  XOR U7032 ( .A(n3443), .B(n3444), .Z(n3442) );
  XOR U7033 ( .A(DB[3185]), .B(DB[3170]), .Z(n3444) );
  AND U7034 ( .A(n178), .B(n3445), .Z(n3443) );
  XOR U7035 ( .A(n3446), .B(n3447), .Z(n3445) );
  XOR U7036 ( .A(DB[3170]), .B(DB[3155]), .Z(n3447) );
  AND U7037 ( .A(n182), .B(n3448), .Z(n3446) );
  XOR U7038 ( .A(n3449), .B(n3450), .Z(n3448) );
  XOR U7039 ( .A(DB[3155]), .B(DB[3140]), .Z(n3450) );
  AND U7040 ( .A(n186), .B(n3451), .Z(n3449) );
  XOR U7041 ( .A(n3452), .B(n3453), .Z(n3451) );
  XOR U7042 ( .A(DB[3140]), .B(DB[3125]), .Z(n3453) );
  AND U7043 ( .A(n190), .B(n3454), .Z(n3452) );
  XOR U7044 ( .A(n3455), .B(n3456), .Z(n3454) );
  XOR U7045 ( .A(DB[3125]), .B(DB[3110]), .Z(n3456) );
  AND U7046 ( .A(n194), .B(n3457), .Z(n3455) );
  XOR U7047 ( .A(n3458), .B(n3459), .Z(n3457) );
  XOR U7048 ( .A(DB[3110]), .B(DB[3095]), .Z(n3459) );
  AND U7049 ( .A(n198), .B(n3460), .Z(n3458) );
  XOR U7050 ( .A(n3461), .B(n3462), .Z(n3460) );
  XOR U7051 ( .A(DB[3095]), .B(DB[3080]), .Z(n3462) );
  AND U7052 ( .A(n202), .B(n3463), .Z(n3461) );
  XOR U7053 ( .A(n3464), .B(n3465), .Z(n3463) );
  XOR U7054 ( .A(DB[3080]), .B(DB[3065]), .Z(n3465) );
  AND U7055 ( .A(n206), .B(n3466), .Z(n3464) );
  XOR U7056 ( .A(n3467), .B(n3468), .Z(n3466) );
  XOR U7057 ( .A(DB[3065]), .B(DB[3050]), .Z(n3468) );
  AND U7058 ( .A(n210), .B(n3469), .Z(n3467) );
  XOR U7059 ( .A(n3470), .B(n3471), .Z(n3469) );
  XOR U7060 ( .A(DB[3050]), .B(DB[3035]), .Z(n3471) );
  AND U7061 ( .A(n214), .B(n3472), .Z(n3470) );
  XOR U7062 ( .A(n3473), .B(n3474), .Z(n3472) );
  XOR U7063 ( .A(DB[3035]), .B(DB[3020]), .Z(n3474) );
  AND U7064 ( .A(n218), .B(n3475), .Z(n3473) );
  XOR U7065 ( .A(n3476), .B(n3477), .Z(n3475) );
  XOR U7066 ( .A(DB[3020]), .B(DB[3005]), .Z(n3477) );
  AND U7067 ( .A(n222), .B(n3478), .Z(n3476) );
  XOR U7068 ( .A(n3479), .B(n3480), .Z(n3478) );
  XOR U7069 ( .A(DB[3005]), .B(DB[2990]), .Z(n3480) );
  AND U7070 ( .A(n226), .B(n3481), .Z(n3479) );
  XOR U7071 ( .A(n3482), .B(n3483), .Z(n3481) );
  XOR U7072 ( .A(DB[2990]), .B(DB[2975]), .Z(n3483) );
  AND U7073 ( .A(n230), .B(n3484), .Z(n3482) );
  XOR U7074 ( .A(n3485), .B(n3486), .Z(n3484) );
  XOR U7075 ( .A(DB[2975]), .B(DB[2960]), .Z(n3486) );
  AND U7076 ( .A(n234), .B(n3487), .Z(n3485) );
  XOR U7077 ( .A(n3488), .B(n3489), .Z(n3487) );
  XOR U7078 ( .A(DB[2960]), .B(DB[2945]), .Z(n3489) );
  AND U7079 ( .A(n238), .B(n3490), .Z(n3488) );
  XOR U7080 ( .A(n3491), .B(n3492), .Z(n3490) );
  XOR U7081 ( .A(DB[2945]), .B(DB[2930]), .Z(n3492) );
  AND U7082 ( .A(n242), .B(n3493), .Z(n3491) );
  XOR U7083 ( .A(n3494), .B(n3495), .Z(n3493) );
  XOR U7084 ( .A(DB[2930]), .B(DB[2915]), .Z(n3495) );
  AND U7085 ( .A(n246), .B(n3496), .Z(n3494) );
  XOR U7086 ( .A(n3497), .B(n3498), .Z(n3496) );
  XOR U7087 ( .A(DB[2915]), .B(DB[2900]), .Z(n3498) );
  AND U7088 ( .A(n250), .B(n3499), .Z(n3497) );
  XOR U7089 ( .A(n3500), .B(n3501), .Z(n3499) );
  XOR U7090 ( .A(DB[2900]), .B(DB[2885]), .Z(n3501) );
  AND U7091 ( .A(n254), .B(n3502), .Z(n3500) );
  XOR U7092 ( .A(n3503), .B(n3504), .Z(n3502) );
  XOR U7093 ( .A(DB[2885]), .B(DB[2870]), .Z(n3504) );
  AND U7094 ( .A(n258), .B(n3505), .Z(n3503) );
  XOR U7095 ( .A(n3506), .B(n3507), .Z(n3505) );
  XOR U7096 ( .A(DB[2870]), .B(DB[2855]), .Z(n3507) );
  AND U7097 ( .A(n262), .B(n3508), .Z(n3506) );
  XOR U7098 ( .A(n3509), .B(n3510), .Z(n3508) );
  XOR U7099 ( .A(DB[2855]), .B(DB[2840]), .Z(n3510) );
  AND U7100 ( .A(n266), .B(n3511), .Z(n3509) );
  XOR U7101 ( .A(n3512), .B(n3513), .Z(n3511) );
  XOR U7102 ( .A(DB[2840]), .B(DB[2825]), .Z(n3513) );
  AND U7103 ( .A(n270), .B(n3514), .Z(n3512) );
  XOR U7104 ( .A(n3515), .B(n3516), .Z(n3514) );
  XOR U7105 ( .A(DB[2825]), .B(DB[2810]), .Z(n3516) );
  AND U7106 ( .A(n274), .B(n3517), .Z(n3515) );
  XOR U7107 ( .A(n3518), .B(n3519), .Z(n3517) );
  XOR U7108 ( .A(DB[2810]), .B(DB[2795]), .Z(n3519) );
  AND U7109 ( .A(n278), .B(n3520), .Z(n3518) );
  XOR U7110 ( .A(n3521), .B(n3522), .Z(n3520) );
  XOR U7111 ( .A(DB[2795]), .B(DB[2780]), .Z(n3522) );
  AND U7112 ( .A(n282), .B(n3523), .Z(n3521) );
  XOR U7113 ( .A(n3524), .B(n3525), .Z(n3523) );
  XOR U7114 ( .A(DB[2780]), .B(DB[2765]), .Z(n3525) );
  AND U7115 ( .A(n286), .B(n3526), .Z(n3524) );
  XOR U7116 ( .A(n3527), .B(n3528), .Z(n3526) );
  XOR U7117 ( .A(DB[2765]), .B(DB[2750]), .Z(n3528) );
  AND U7118 ( .A(n290), .B(n3529), .Z(n3527) );
  XOR U7119 ( .A(n3530), .B(n3531), .Z(n3529) );
  XOR U7120 ( .A(DB[2750]), .B(DB[2735]), .Z(n3531) );
  AND U7121 ( .A(n294), .B(n3532), .Z(n3530) );
  XOR U7122 ( .A(n3533), .B(n3534), .Z(n3532) );
  XOR U7123 ( .A(DB[2735]), .B(DB[2720]), .Z(n3534) );
  AND U7124 ( .A(n298), .B(n3535), .Z(n3533) );
  XOR U7125 ( .A(n3536), .B(n3537), .Z(n3535) );
  XOR U7126 ( .A(DB[2720]), .B(DB[2705]), .Z(n3537) );
  AND U7127 ( .A(n302), .B(n3538), .Z(n3536) );
  XOR U7128 ( .A(n3539), .B(n3540), .Z(n3538) );
  XOR U7129 ( .A(DB[2705]), .B(DB[2690]), .Z(n3540) );
  AND U7130 ( .A(n306), .B(n3541), .Z(n3539) );
  XOR U7131 ( .A(n3542), .B(n3543), .Z(n3541) );
  XOR U7132 ( .A(DB[2690]), .B(DB[2675]), .Z(n3543) );
  AND U7133 ( .A(n310), .B(n3544), .Z(n3542) );
  XOR U7134 ( .A(n3545), .B(n3546), .Z(n3544) );
  XOR U7135 ( .A(DB[2675]), .B(DB[2660]), .Z(n3546) );
  AND U7136 ( .A(n314), .B(n3547), .Z(n3545) );
  XOR U7137 ( .A(n3548), .B(n3549), .Z(n3547) );
  XOR U7138 ( .A(DB[2660]), .B(DB[2645]), .Z(n3549) );
  AND U7139 ( .A(n318), .B(n3550), .Z(n3548) );
  XOR U7140 ( .A(n3551), .B(n3552), .Z(n3550) );
  XOR U7141 ( .A(DB[2645]), .B(DB[2630]), .Z(n3552) );
  AND U7142 ( .A(n322), .B(n3553), .Z(n3551) );
  XOR U7143 ( .A(n3554), .B(n3555), .Z(n3553) );
  XOR U7144 ( .A(DB[2630]), .B(DB[2615]), .Z(n3555) );
  AND U7145 ( .A(n326), .B(n3556), .Z(n3554) );
  XOR U7146 ( .A(n3557), .B(n3558), .Z(n3556) );
  XOR U7147 ( .A(DB[2615]), .B(DB[2600]), .Z(n3558) );
  AND U7148 ( .A(n330), .B(n3559), .Z(n3557) );
  XOR U7149 ( .A(n3560), .B(n3561), .Z(n3559) );
  XOR U7150 ( .A(DB[2600]), .B(DB[2585]), .Z(n3561) );
  AND U7151 ( .A(n334), .B(n3562), .Z(n3560) );
  XOR U7152 ( .A(n3563), .B(n3564), .Z(n3562) );
  XOR U7153 ( .A(DB[2585]), .B(DB[2570]), .Z(n3564) );
  AND U7154 ( .A(n338), .B(n3565), .Z(n3563) );
  XOR U7155 ( .A(n3566), .B(n3567), .Z(n3565) );
  XOR U7156 ( .A(DB[2570]), .B(DB[2555]), .Z(n3567) );
  AND U7157 ( .A(n342), .B(n3568), .Z(n3566) );
  XOR U7158 ( .A(n3569), .B(n3570), .Z(n3568) );
  XOR U7159 ( .A(DB[2555]), .B(DB[2540]), .Z(n3570) );
  AND U7160 ( .A(n346), .B(n3571), .Z(n3569) );
  XOR U7161 ( .A(n3572), .B(n3573), .Z(n3571) );
  XOR U7162 ( .A(DB[2540]), .B(DB[2525]), .Z(n3573) );
  AND U7163 ( .A(n350), .B(n3574), .Z(n3572) );
  XOR U7164 ( .A(n3575), .B(n3576), .Z(n3574) );
  XOR U7165 ( .A(DB[2525]), .B(DB[2510]), .Z(n3576) );
  AND U7166 ( .A(n354), .B(n3577), .Z(n3575) );
  XOR U7167 ( .A(n3578), .B(n3579), .Z(n3577) );
  XOR U7168 ( .A(DB[2510]), .B(DB[2495]), .Z(n3579) );
  AND U7169 ( .A(n358), .B(n3580), .Z(n3578) );
  XOR U7170 ( .A(n3581), .B(n3582), .Z(n3580) );
  XOR U7171 ( .A(DB[2495]), .B(DB[2480]), .Z(n3582) );
  AND U7172 ( .A(n362), .B(n3583), .Z(n3581) );
  XOR U7173 ( .A(n3584), .B(n3585), .Z(n3583) );
  XOR U7174 ( .A(DB[2480]), .B(DB[2465]), .Z(n3585) );
  AND U7175 ( .A(n366), .B(n3586), .Z(n3584) );
  XOR U7176 ( .A(n3587), .B(n3588), .Z(n3586) );
  XOR U7177 ( .A(DB[2465]), .B(DB[2450]), .Z(n3588) );
  AND U7178 ( .A(n370), .B(n3589), .Z(n3587) );
  XOR U7179 ( .A(n3590), .B(n3591), .Z(n3589) );
  XOR U7180 ( .A(DB[2450]), .B(DB[2435]), .Z(n3591) );
  AND U7181 ( .A(n374), .B(n3592), .Z(n3590) );
  XOR U7182 ( .A(n3593), .B(n3594), .Z(n3592) );
  XOR U7183 ( .A(DB[2435]), .B(DB[2420]), .Z(n3594) );
  AND U7184 ( .A(n378), .B(n3595), .Z(n3593) );
  XOR U7185 ( .A(n3596), .B(n3597), .Z(n3595) );
  XOR U7186 ( .A(DB[2420]), .B(DB[2405]), .Z(n3597) );
  AND U7187 ( .A(n382), .B(n3598), .Z(n3596) );
  XOR U7188 ( .A(n3599), .B(n3600), .Z(n3598) );
  XOR U7189 ( .A(DB[2405]), .B(DB[2390]), .Z(n3600) );
  AND U7190 ( .A(n386), .B(n3601), .Z(n3599) );
  XOR U7191 ( .A(n3602), .B(n3603), .Z(n3601) );
  XOR U7192 ( .A(DB[2390]), .B(DB[2375]), .Z(n3603) );
  AND U7193 ( .A(n390), .B(n3604), .Z(n3602) );
  XOR U7194 ( .A(n3605), .B(n3606), .Z(n3604) );
  XOR U7195 ( .A(DB[2375]), .B(DB[2360]), .Z(n3606) );
  AND U7196 ( .A(n394), .B(n3607), .Z(n3605) );
  XOR U7197 ( .A(n3608), .B(n3609), .Z(n3607) );
  XOR U7198 ( .A(DB[2360]), .B(DB[2345]), .Z(n3609) );
  AND U7199 ( .A(n398), .B(n3610), .Z(n3608) );
  XOR U7200 ( .A(n3611), .B(n3612), .Z(n3610) );
  XOR U7201 ( .A(DB[2345]), .B(DB[2330]), .Z(n3612) );
  AND U7202 ( .A(n402), .B(n3613), .Z(n3611) );
  XOR U7203 ( .A(n3614), .B(n3615), .Z(n3613) );
  XOR U7204 ( .A(DB[2330]), .B(DB[2315]), .Z(n3615) );
  AND U7205 ( .A(n406), .B(n3616), .Z(n3614) );
  XOR U7206 ( .A(n3617), .B(n3618), .Z(n3616) );
  XOR U7207 ( .A(DB[2315]), .B(DB[2300]), .Z(n3618) );
  AND U7208 ( .A(n410), .B(n3619), .Z(n3617) );
  XOR U7209 ( .A(n3620), .B(n3621), .Z(n3619) );
  XOR U7210 ( .A(DB[2300]), .B(DB[2285]), .Z(n3621) );
  AND U7211 ( .A(n414), .B(n3622), .Z(n3620) );
  XOR U7212 ( .A(n3623), .B(n3624), .Z(n3622) );
  XOR U7213 ( .A(DB[2285]), .B(DB[2270]), .Z(n3624) );
  AND U7214 ( .A(n418), .B(n3625), .Z(n3623) );
  XOR U7215 ( .A(n3626), .B(n3627), .Z(n3625) );
  XOR U7216 ( .A(DB[2270]), .B(DB[2255]), .Z(n3627) );
  AND U7217 ( .A(n422), .B(n3628), .Z(n3626) );
  XOR U7218 ( .A(n3629), .B(n3630), .Z(n3628) );
  XOR U7219 ( .A(DB[2255]), .B(DB[2240]), .Z(n3630) );
  AND U7220 ( .A(n426), .B(n3631), .Z(n3629) );
  XOR U7221 ( .A(n3632), .B(n3633), .Z(n3631) );
  XOR U7222 ( .A(DB[2240]), .B(DB[2225]), .Z(n3633) );
  AND U7223 ( .A(n430), .B(n3634), .Z(n3632) );
  XOR U7224 ( .A(n3635), .B(n3636), .Z(n3634) );
  XOR U7225 ( .A(DB[2225]), .B(DB[2210]), .Z(n3636) );
  AND U7226 ( .A(n434), .B(n3637), .Z(n3635) );
  XOR U7227 ( .A(n3638), .B(n3639), .Z(n3637) );
  XOR U7228 ( .A(DB[2210]), .B(DB[2195]), .Z(n3639) );
  AND U7229 ( .A(n438), .B(n3640), .Z(n3638) );
  XOR U7230 ( .A(n3641), .B(n3642), .Z(n3640) );
  XOR U7231 ( .A(DB[2195]), .B(DB[2180]), .Z(n3642) );
  AND U7232 ( .A(n442), .B(n3643), .Z(n3641) );
  XOR U7233 ( .A(n3644), .B(n3645), .Z(n3643) );
  XOR U7234 ( .A(DB[2180]), .B(DB[2165]), .Z(n3645) );
  AND U7235 ( .A(n446), .B(n3646), .Z(n3644) );
  XOR U7236 ( .A(n3647), .B(n3648), .Z(n3646) );
  XOR U7237 ( .A(DB[2165]), .B(DB[2150]), .Z(n3648) );
  AND U7238 ( .A(n450), .B(n3649), .Z(n3647) );
  XOR U7239 ( .A(n3650), .B(n3651), .Z(n3649) );
  XOR U7240 ( .A(DB[2150]), .B(DB[2135]), .Z(n3651) );
  AND U7241 ( .A(n454), .B(n3652), .Z(n3650) );
  XOR U7242 ( .A(n3653), .B(n3654), .Z(n3652) );
  XOR U7243 ( .A(DB[2135]), .B(DB[2120]), .Z(n3654) );
  AND U7244 ( .A(n458), .B(n3655), .Z(n3653) );
  XOR U7245 ( .A(n3656), .B(n3657), .Z(n3655) );
  XOR U7246 ( .A(DB[2120]), .B(DB[2105]), .Z(n3657) );
  AND U7247 ( .A(n462), .B(n3658), .Z(n3656) );
  XOR U7248 ( .A(n3659), .B(n3660), .Z(n3658) );
  XOR U7249 ( .A(DB[2105]), .B(DB[2090]), .Z(n3660) );
  AND U7250 ( .A(n466), .B(n3661), .Z(n3659) );
  XOR U7251 ( .A(n3662), .B(n3663), .Z(n3661) );
  XOR U7252 ( .A(DB[2090]), .B(DB[2075]), .Z(n3663) );
  AND U7253 ( .A(n470), .B(n3664), .Z(n3662) );
  XOR U7254 ( .A(n3665), .B(n3666), .Z(n3664) );
  XOR U7255 ( .A(DB[2075]), .B(DB[2060]), .Z(n3666) );
  AND U7256 ( .A(n474), .B(n3667), .Z(n3665) );
  XOR U7257 ( .A(n3668), .B(n3669), .Z(n3667) );
  XOR U7258 ( .A(DB[2060]), .B(DB[2045]), .Z(n3669) );
  AND U7259 ( .A(n478), .B(n3670), .Z(n3668) );
  XOR U7260 ( .A(n3671), .B(n3672), .Z(n3670) );
  XOR U7261 ( .A(DB[2045]), .B(DB[2030]), .Z(n3672) );
  AND U7262 ( .A(n482), .B(n3673), .Z(n3671) );
  XOR U7263 ( .A(n3674), .B(n3675), .Z(n3673) );
  XOR U7264 ( .A(DB[2030]), .B(DB[2015]), .Z(n3675) );
  AND U7265 ( .A(n486), .B(n3676), .Z(n3674) );
  XOR U7266 ( .A(n3677), .B(n3678), .Z(n3676) );
  XOR U7267 ( .A(DB[2015]), .B(DB[2000]), .Z(n3678) );
  AND U7268 ( .A(n490), .B(n3679), .Z(n3677) );
  XOR U7269 ( .A(n3680), .B(n3681), .Z(n3679) );
  XOR U7270 ( .A(DB[2000]), .B(DB[1985]), .Z(n3681) );
  AND U7271 ( .A(n494), .B(n3682), .Z(n3680) );
  XOR U7272 ( .A(n3683), .B(n3684), .Z(n3682) );
  XOR U7273 ( .A(DB[1985]), .B(DB[1970]), .Z(n3684) );
  AND U7274 ( .A(n498), .B(n3685), .Z(n3683) );
  XOR U7275 ( .A(n3686), .B(n3687), .Z(n3685) );
  XOR U7276 ( .A(DB[1970]), .B(DB[1955]), .Z(n3687) );
  AND U7277 ( .A(n502), .B(n3688), .Z(n3686) );
  XOR U7278 ( .A(n3689), .B(n3690), .Z(n3688) );
  XOR U7279 ( .A(DB[1955]), .B(DB[1940]), .Z(n3690) );
  AND U7280 ( .A(n506), .B(n3691), .Z(n3689) );
  XOR U7281 ( .A(n3692), .B(n3693), .Z(n3691) );
  XOR U7282 ( .A(DB[1940]), .B(DB[1925]), .Z(n3693) );
  AND U7283 ( .A(n510), .B(n3694), .Z(n3692) );
  XOR U7284 ( .A(n3695), .B(n3696), .Z(n3694) );
  XOR U7285 ( .A(DB[1925]), .B(DB[1910]), .Z(n3696) );
  AND U7286 ( .A(n514), .B(n3697), .Z(n3695) );
  XOR U7287 ( .A(n3698), .B(n3699), .Z(n3697) );
  XOR U7288 ( .A(DB[1910]), .B(DB[1895]), .Z(n3699) );
  AND U7289 ( .A(n518), .B(n3700), .Z(n3698) );
  XOR U7290 ( .A(n3701), .B(n3702), .Z(n3700) );
  XOR U7291 ( .A(DB[1895]), .B(DB[1880]), .Z(n3702) );
  AND U7292 ( .A(n522), .B(n3703), .Z(n3701) );
  XOR U7293 ( .A(n3704), .B(n3705), .Z(n3703) );
  XOR U7294 ( .A(DB[1880]), .B(DB[1865]), .Z(n3705) );
  AND U7295 ( .A(n526), .B(n3706), .Z(n3704) );
  XOR U7296 ( .A(n3707), .B(n3708), .Z(n3706) );
  XOR U7297 ( .A(DB[1865]), .B(DB[1850]), .Z(n3708) );
  AND U7298 ( .A(n530), .B(n3709), .Z(n3707) );
  XOR U7299 ( .A(n3710), .B(n3711), .Z(n3709) );
  XOR U7300 ( .A(DB[1850]), .B(DB[1835]), .Z(n3711) );
  AND U7301 ( .A(n534), .B(n3712), .Z(n3710) );
  XOR U7302 ( .A(n3713), .B(n3714), .Z(n3712) );
  XOR U7303 ( .A(DB[1835]), .B(DB[1820]), .Z(n3714) );
  AND U7304 ( .A(n538), .B(n3715), .Z(n3713) );
  XOR U7305 ( .A(n3716), .B(n3717), .Z(n3715) );
  XOR U7306 ( .A(DB[1820]), .B(DB[1805]), .Z(n3717) );
  AND U7307 ( .A(n542), .B(n3718), .Z(n3716) );
  XOR U7308 ( .A(n3719), .B(n3720), .Z(n3718) );
  XOR U7309 ( .A(DB[1805]), .B(DB[1790]), .Z(n3720) );
  AND U7310 ( .A(n546), .B(n3721), .Z(n3719) );
  XOR U7311 ( .A(n3722), .B(n3723), .Z(n3721) );
  XOR U7312 ( .A(DB[1790]), .B(DB[1775]), .Z(n3723) );
  AND U7313 ( .A(n550), .B(n3724), .Z(n3722) );
  XOR U7314 ( .A(n3725), .B(n3726), .Z(n3724) );
  XOR U7315 ( .A(DB[1775]), .B(DB[1760]), .Z(n3726) );
  AND U7316 ( .A(n554), .B(n3727), .Z(n3725) );
  XOR U7317 ( .A(n3728), .B(n3729), .Z(n3727) );
  XOR U7318 ( .A(DB[1760]), .B(DB[1745]), .Z(n3729) );
  AND U7319 ( .A(n558), .B(n3730), .Z(n3728) );
  XOR U7320 ( .A(n3731), .B(n3732), .Z(n3730) );
  XOR U7321 ( .A(DB[1745]), .B(DB[1730]), .Z(n3732) );
  AND U7322 ( .A(n562), .B(n3733), .Z(n3731) );
  XOR U7323 ( .A(n3734), .B(n3735), .Z(n3733) );
  XOR U7324 ( .A(DB[1730]), .B(DB[1715]), .Z(n3735) );
  AND U7325 ( .A(n566), .B(n3736), .Z(n3734) );
  XOR U7326 ( .A(n3737), .B(n3738), .Z(n3736) );
  XOR U7327 ( .A(DB[1715]), .B(DB[1700]), .Z(n3738) );
  AND U7328 ( .A(n570), .B(n3739), .Z(n3737) );
  XOR U7329 ( .A(n3740), .B(n3741), .Z(n3739) );
  XOR U7330 ( .A(DB[1700]), .B(DB[1685]), .Z(n3741) );
  AND U7331 ( .A(n574), .B(n3742), .Z(n3740) );
  XOR U7332 ( .A(n3743), .B(n3744), .Z(n3742) );
  XOR U7333 ( .A(DB[1685]), .B(DB[1670]), .Z(n3744) );
  AND U7334 ( .A(n578), .B(n3745), .Z(n3743) );
  XOR U7335 ( .A(n3746), .B(n3747), .Z(n3745) );
  XOR U7336 ( .A(DB[1670]), .B(DB[1655]), .Z(n3747) );
  AND U7337 ( .A(n582), .B(n3748), .Z(n3746) );
  XOR U7338 ( .A(n3749), .B(n3750), .Z(n3748) );
  XOR U7339 ( .A(DB[1655]), .B(DB[1640]), .Z(n3750) );
  AND U7340 ( .A(n586), .B(n3751), .Z(n3749) );
  XOR U7341 ( .A(n3752), .B(n3753), .Z(n3751) );
  XOR U7342 ( .A(DB[1640]), .B(DB[1625]), .Z(n3753) );
  AND U7343 ( .A(n590), .B(n3754), .Z(n3752) );
  XOR U7344 ( .A(n3755), .B(n3756), .Z(n3754) );
  XOR U7345 ( .A(DB[1625]), .B(DB[1610]), .Z(n3756) );
  AND U7346 ( .A(n594), .B(n3757), .Z(n3755) );
  XOR U7347 ( .A(n3758), .B(n3759), .Z(n3757) );
  XOR U7348 ( .A(DB[1610]), .B(DB[1595]), .Z(n3759) );
  AND U7349 ( .A(n598), .B(n3760), .Z(n3758) );
  XOR U7350 ( .A(n3761), .B(n3762), .Z(n3760) );
  XOR U7351 ( .A(DB[1595]), .B(DB[1580]), .Z(n3762) );
  AND U7352 ( .A(n602), .B(n3763), .Z(n3761) );
  XOR U7353 ( .A(n3764), .B(n3765), .Z(n3763) );
  XOR U7354 ( .A(DB[1580]), .B(DB[1565]), .Z(n3765) );
  AND U7355 ( .A(n606), .B(n3766), .Z(n3764) );
  XOR U7356 ( .A(n3767), .B(n3768), .Z(n3766) );
  XOR U7357 ( .A(DB[1565]), .B(DB[1550]), .Z(n3768) );
  AND U7358 ( .A(n610), .B(n3769), .Z(n3767) );
  XOR U7359 ( .A(n3770), .B(n3771), .Z(n3769) );
  XOR U7360 ( .A(DB[1550]), .B(DB[1535]), .Z(n3771) );
  AND U7361 ( .A(n614), .B(n3772), .Z(n3770) );
  XOR U7362 ( .A(n3773), .B(n3774), .Z(n3772) );
  XOR U7363 ( .A(DB[1535]), .B(DB[1520]), .Z(n3774) );
  AND U7364 ( .A(n618), .B(n3775), .Z(n3773) );
  XOR U7365 ( .A(n3776), .B(n3777), .Z(n3775) );
  XOR U7366 ( .A(DB[1520]), .B(DB[1505]), .Z(n3777) );
  AND U7367 ( .A(n622), .B(n3778), .Z(n3776) );
  XOR U7368 ( .A(n3779), .B(n3780), .Z(n3778) );
  XOR U7369 ( .A(DB[1505]), .B(DB[1490]), .Z(n3780) );
  AND U7370 ( .A(n626), .B(n3781), .Z(n3779) );
  XOR U7371 ( .A(n3782), .B(n3783), .Z(n3781) );
  XOR U7372 ( .A(DB[1490]), .B(DB[1475]), .Z(n3783) );
  AND U7373 ( .A(n630), .B(n3784), .Z(n3782) );
  XOR U7374 ( .A(n3785), .B(n3786), .Z(n3784) );
  XOR U7375 ( .A(DB[1475]), .B(DB[1460]), .Z(n3786) );
  AND U7376 ( .A(n634), .B(n3787), .Z(n3785) );
  XOR U7377 ( .A(n3788), .B(n3789), .Z(n3787) );
  XOR U7378 ( .A(DB[1460]), .B(DB[1445]), .Z(n3789) );
  AND U7379 ( .A(n638), .B(n3790), .Z(n3788) );
  XOR U7380 ( .A(n3791), .B(n3792), .Z(n3790) );
  XOR U7381 ( .A(DB[1445]), .B(DB[1430]), .Z(n3792) );
  AND U7382 ( .A(n642), .B(n3793), .Z(n3791) );
  XOR U7383 ( .A(n3794), .B(n3795), .Z(n3793) );
  XOR U7384 ( .A(DB[1430]), .B(DB[1415]), .Z(n3795) );
  AND U7385 ( .A(n646), .B(n3796), .Z(n3794) );
  XOR U7386 ( .A(n3797), .B(n3798), .Z(n3796) );
  XOR U7387 ( .A(DB[1415]), .B(DB[1400]), .Z(n3798) );
  AND U7388 ( .A(n650), .B(n3799), .Z(n3797) );
  XOR U7389 ( .A(n3800), .B(n3801), .Z(n3799) );
  XOR U7390 ( .A(DB[1400]), .B(DB[1385]), .Z(n3801) );
  AND U7391 ( .A(n654), .B(n3802), .Z(n3800) );
  XOR U7392 ( .A(n3803), .B(n3804), .Z(n3802) );
  XOR U7393 ( .A(DB[1385]), .B(DB[1370]), .Z(n3804) );
  AND U7394 ( .A(n658), .B(n3805), .Z(n3803) );
  XOR U7395 ( .A(n3806), .B(n3807), .Z(n3805) );
  XOR U7396 ( .A(DB[1370]), .B(DB[1355]), .Z(n3807) );
  AND U7397 ( .A(n662), .B(n3808), .Z(n3806) );
  XOR U7398 ( .A(n3809), .B(n3810), .Z(n3808) );
  XOR U7399 ( .A(DB[1355]), .B(DB[1340]), .Z(n3810) );
  AND U7400 ( .A(n666), .B(n3811), .Z(n3809) );
  XOR U7401 ( .A(n3812), .B(n3813), .Z(n3811) );
  XOR U7402 ( .A(DB[1340]), .B(DB[1325]), .Z(n3813) );
  AND U7403 ( .A(n670), .B(n3814), .Z(n3812) );
  XOR U7404 ( .A(n3815), .B(n3816), .Z(n3814) );
  XOR U7405 ( .A(DB[1325]), .B(DB[1310]), .Z(n3816) );
  AND U7406 ( .A(n674), .B(n3817), .Z(n3815) );
  XOR U7407 ( .A(n3818), .B(n3819), .Z(n3817) );
  XOR U7408 ( .A(DB[1310]), .B(DB[1295]), .Z(n3819) );
  AND U7409 ( .A(n678), .B(n3820), .Z(n3818) );
  XOR U7410 ( .A(n3821), .B(n3822), .Z(n3820) );
  XOR U7411 ( .A(DB[1295]), .B(DB[1280]), .Z(n3822) );
  AND U7412 ( .A(n682), .B(n3823), .Z(n3821) );
  XOR U7413 ( .A(n3824), .B(n3825), .Z(n3823) );
  XOR U7414 ( .A(DB[1280]), .B(DB[1265]), .Z(n3825) );
  AND U7415 ( .A(n686), .B(n3826), .Z(n3824) );
  XOR U7416 ( .A(n3827), .B(n3828), .Z(n3826) );
  XOR U7417 ( .A(DB[1265]), .B(DB[1250]), .Z(n3828) );
  AND U7418 ( .A(n690), .B(n3829), .Z(n3827) );
  XOR U7419 ( .A(n3830), .B(n3831), .Z(n3829) );
  XOR U7420 ( .A(DB[1250]), .B(DB[1235]), .Z(n3831) );
  AND U7421 ( .A(n694), .B(n3832), .Z(n3830) );
  XOR U7422 ( .A(n3833), .B(n3834), .Z(n3832) );
  XOR U7423 ( .A(DB[1235]), .B(DB[1220]), .Z(n3834) );
  AND U7424 ( .A(n698), .B(n3835), .Z(n3833) );
  XOR U7425 ( .A(n3836), .B(n3837), .Z(n3835) );
  XOR U7426 ( .A(DB[1220]), .B(DB[1205]), .Z(n3837) );
  AND U7427 ( .A(n702), .B(n3838), .Z(n3836) );
  XOR U7428 ( .A(n3839), .B(n3840), .Z(n3838) );
  XOR U7429 ( .A(DB[1205]), .B(DB[1190]), .Z(n3840) );
  AND U7430 ( .A(n706), .B(n3841), .Z(n3839) );
  XOR U7431 ( .A(n3842), .B(n3843), .Z(n3841) );
  XOR U7432 ( .A(DB[1190]), .B(DB[1175]), .Z(n3843) );
  AND U7433 ( .A(n710), .B(n3844), .Z(n3842) );
  XOR U7434 ( .A(n3845), .B(n3846), .Z(n3844) );
  XOR U7435 ( .A(DB[1175]), .B(DB[1160]), .Z(n3846) );
  AND U7436 ( .A(n714), .B(n3847), .Z(n3845) );
  XOR U7437 ( .A(n3848), .B(n3849), .Z(n3847) );
  XOR U7438 ( .A(DB[1160]), .B(DB[1145]), .Z(n3849) );
  AND U7439 ( .A(n718), .B(n3850), .Z(n3848) );
  XOR U7440 ( .A(n3851), .B(n3852), .Z(n3850) );
  XOR U7441 ( .A(DB[1145]), .B(DB[1130]), .Z(n3852) );
  AND U7442 ( .A(n722), .B(n3853), .Z(n3851) );
  XOR U7443 ( .A(n3854), .B(n3855), .Z(n3853) );
  XOR U7444 ( .A(DB[1130]), .B(DB[1115]), .Z(n3855) );
  AND U7445 ( .A(n726), .B(n3856), .Z(n3854) );
  XOR U7446 ( .A(n3857), .B(n3858), .Z(n3856) );
  XOR U7447 ( .A(DB[1115]), .B(DB[1100]), .Z(n3858) );
  AND U7448 ( .A(n730), .B(n3859), .Z(n3857) );
  XOR U7449 ( .A(n3860), .B(n3861), .Z(n3859) );
  XOR U7450 ( .A(DB[1100]), .B(DB[1085]), .Z(n3861) );
  AND U7451 ( .A(n734), .B(n3862), .Z(n3860) );
  XOR U7452 ( .A(n3863), .B(n3864), .Z(n3862) );
  XOR U7453 ( .A(DB[1085]), .B(DB[1070]), .Z(n3864) );
  AND U7454 ( .A(n738), .B(n3865), .Z(n3863) );
  XOR U7455 ( .A(n3866), .B(n3867), .Z(n3865) );
  XOR U7456 ( .A(DB[1070]), .B(DB[1055]), .Z(n3867) );
  AND U7457 ( .A(n742), .B(n3868), .Z(n3866) );
  XOR U7458 ( .A(n3869), .B(n3870), .Z(n3868) );
  XOR U7459 ( .A(DB[1055]), .B(DB[1040]), .Z(n3870) );
  AND U7460 ( .A(n746), .B(n3871), .Z(n3869) );
  XOR U7461 ( .A(n3872), .B(n3873), .Z(n3871) );
  XOR U7462 ( .A(DB[1040]), .B(DB[1025]), .Z(n3873) );
  AND U7463 ( .A(n750), .B(n3874), .Z(n3872) );
  XOR U7464 ( .A(n3875), .B(n3876), .Z(n3874) );
  XOR U7465 ( .A(DB[1025]), .B(DB[1010]), .Z(n3876) );
  AND U7466 ( .A(n754), .B(n3877), .Z(n3875) );
  XOR U7467 ( .A(n3878), .B(n3879), .Z(n3877) );
  XOR U7468 ( .A(DB[995]), .B(DB[1010]), .Z(n3879) );
  AND U7469 ( .A(n758), .B(n3880), .Z(n3878) );
  XOR U7470 ( .A(n3881), .B(n3882), .Z(n3880) );
  XOR U7471 ( .A(DB[995]), .B(DB[980]), .Z(n3882) );
  AND U7472 ( .A(n762), .B(n3883), .Z(n3881) );
  XOR U7473 ( .A(n3884), .B(n3885), .Z(n3883) );
  XOR U7474 ( .A(DB[980]), .B(DB[965]), .Z(n3885) );
  AND U7475 ( .A(n766), .B(n3886), .Z(n3884) );
  XOR U7476 ( .A(n3887), .B(n3888), .Z(n3886) );
  XOR U7477 ( .A(DB[965]), .B(DB[950]), .Z(n3888) );
  AND U7478 ( .A(n770), .B(n3889), .Z(n3887) );
  XOR U7479 ( .A(n3890), .B(n3891), .Z(n3889) );
  XOR U7480 ( .A(DB[950]), .B(DB[935]), .Z(n3891) );
  AND U7481 ( .A(n774), .B(n3892), .Z(n3890) );
  XOR U7482 ( .A(n3893), .B(n3894), .Z(n3892) );
  XOR U7483 ( .A(DB[935]), .B(DB[920]), .Z(n3894) );
  AND U7484 ( .A(n778), .B(n3895), .Z(n3893) );
  XOR U7485 ( .A(n3896), .B(n3897), .Z(n3895) );
  XOR U7486 ( .A(DB[920]), .B(DB[905]), .Z(n3897) );
  AND U7487 ( .A(n782), .B(n3898), .Z(n3896) );
  XOR U7488 ( .A(n3899), .B(n3900), .Z(n3898) );
  XOR U7489 ( .A(DB[905]), .B(DB[890]), .Z(n3900) );
  AND U7490 ( .A(n786), .B(n3901), .Z(n3899) );
  XOR U7491 ( .A(n3902), .B(n3903), .Z(n3901) );
  XOR U7492 ( .A(DB[890]), .B(DB[875]), .Z(n3903) );
  AND U7493 ( .A(n790), .B(n3904), .Z(n3902) );
  XOR U7494 ( .A(n3905), .B(n3906), .Z(n3904) );
  XOR U7495 ( .A(DB[875]), .B(DB[860]), .Z(n3906) );
  AND U7496 ( .A(n794), .B(n3907), .Z(n3905) );
  XOR U7497 ( .A(n3908), .B(n3909), .Z(n3907) );
  XOR U7498 ( .A(DB[860]), .B(DB[845]), .Z(n3909) );
  AND U7499 ( .A(n798), .B(n3910), .Z(n3908) );
  XOR U7500 ( .A(n3911), .B(n3912), .Z(n3910) );
  XOR U7501 ( .A(DB[845]), .B(DB[830]), .Z(n3912) );
  AND U7502 ( .A(n802), .B(n3913), .Z(n3911) );
  XOR U7503 ( .A(n3914), .B(n3915), .Z(n3913) );
  XOR U7504 ( .A(DB[830]), .B(DB[815]), .Z(n3915) );
  AND U7505 ( .A(n806), .B(n3916), .Z(n3914) );
  XOR U7506 ( .A(n3917), .B(n3918), .Z(n3916) );
  XOR U7507 ( .A(DB[815]), .B(DB[800]), .Z(n3918) );
  AND U7508 ( .A(n810), .B(n3919), .Z(n3917) );
  XOR U7509 ( .A(n3920), .B(n3921), .Z(n3919) );
  XOR U7510 ( .A(DB[800]), .B(DB[785]), .Z(n3921) );
  AND U7511 ( .A(n814), .B(n3922), .Z(n3920) );
  XOR U7512 ( .A(n3923), .B(n3924), .Z(n3922) );
  XOR U7513 ( .A(DB[785]), .B(DB[770]), .Z(n3924) );
  AND U7514 ( .A(n818), .B(n3925), .Z(n3923) );
  XOR U7515 ( .A(n3926), .B(n3927), .Z(n3925) );
  XOR U7516 ( .A(DB[770]), .B(DB[755]), .Z(n3927) );
  AND U7517 ( .A(n822), .B(n3928), .Z(n3926) );
  XOR U7518 ( .A(n3929), .B(n3930), .Z(n3928) );
  XOR U7519 ( .A(DB[755]), .B(DB[740]), .Z(n3930) );
  AND U7520 ( .A(n826), .B(n3931), .Z(n3929) );
  XOR U7521 ( .A(n3932), .B(n3933), .Z(n3931) );
  XOR U7522 ( .A(DB[740]), .B(DB[725]), .Z(n3933) );
  AND U7523 ( .A(n830), .B(n3934), .Z(n3932) );
  XOR U7524 ( .A(n3935), .B(n3936), .Z(n3934) );
  XOR U7525 ( .A(DB[725]), .B(DB[710]), .Z(n3936) );
  AND U7526 ( .A(n834), .B(n3937), .Z(n3935) );
  XOR U7527 ( .A(n3938), .B(n3939), .Z(n3937) );
  XOR U7528 ( .A(DB[710]), .B(DB[695]), .Z(n3939) );
  AND U7529 ( .A(n838), .B(n3940), .Z(n3938) );
  XOR U7530 ( .A(n3941), .B(n3942), .Z(n3940) );
  XOR U7531 ( .A(DB[695]), .B(DB[680]), .Z(n3942) );
  AND U7532 ( .A(n842), .B(n3943), .Z(n3941) );
  XOR U7533 ( .A(n3944), .B(n3945), .Z(n3943) );
  XOR U7534 ( .A(DB[680]), .B(DB[665]), .Z(n3945) );
  AND U7535 ( .A(n846), .B(n3946), .Z(n3944) );
  XOR U7536 ( .A(n3947), .B(n3948), .Z(n3946) );
  XOR U7537 ( .A(DB[665]), .B(DB[650]), .Z(n3948) );
  AND U7538 ( .A(n850), .B(n3949), .Z(n3947) );
  XOR U7539 ( .A(n3950), .B(n3951), .Z(n3949) );
  XOR U7540 ( .A(DB[650]), .B(DB[635]), .Z(n3951) );
  AND U7541 ( .A(n854), .B(n3952), .Z(n3950) );
  XOR U7542 ( .A(n3953), .B(n3954), .Z(n3952) );
  XOR U7543 ( .A(DB[635]), .B(DB[620]), .Z(n3954) );
  AND U7544 ( .A(n858), .B(n3955), .Z(n3953) );
  XOR U7545 ( .A(n3956), .B(n3957), .Z(n3955) );
  XOR U7546 ( .A(DB[620]), .B(DB[605]), .Z(n3957) );
  AND U7547 ( .A(n862), .B(n3958), .Z(n3956) );
  XOR U7548 ( .A(n3959), .B(n3960), .Z(n3958) );
  XOR U7549 ( .A(DB[605]), .B(DB[590]), .Z(n3960) );
  AND U7550 ( .A(n866), .B(n3961), .Z(n3959) );
  XOR U7551 ( .A(n3962), .B(n3963), .Z(n3961) );
  XOR U7552 ( .A(DB[590]), .B(DB[575]), .Z(n3963) );
  AND U7553 ( .A(n870), .B(n3964), .Z(n3962) );
  XOR U7554 ( .A(n3965), .B(n3966), .Z(n3964) );
  XOR U7555 ( .A(DB[575]), .B(DB[560]), .Z(n3966) );
  AND U7556 ( .A(n874), .B(n3967), .Z(n3965) );
  XOR U7557 ( .A(n3968), .B(n3969), .Z(n3967) );
  XOR U7558 ( .A(DB[560]), .B(DB[545]), .Z(n3969) );
  AND U7559 ( .A(n878), .B(n3970), .Z(n3968) );
  XOR U7560 ( .A(n3971), .B(n3972), .Z(n3970) );
  XOR U7561 ( .A(DB[545]), .B(DB[530]), .Z(n3972) );
  AND U7562 ( .A(n882), .B(n3973), .Z(n3971) );
  XOR U7563 ( .A(n3974), .B(n3975), .Z(n3973) );
  XOR U7564 ( .A(DB[530]), .B(DB[515]), .Z(n3975) );
  AND U7565 ( .A(n886), .B(n3976), .Z(n3974) );
  XOR U7566 ( .A(n3977), .B(n3978), .Z(n3976) );
  XOR U7567 ( .A(DB[515]), .B(DB[500]), .Z(n3978) );
  AND U7568 ( .A(n890), .B(n3979), .Z(n3977) );
  XOR U7569 ( .A(n3980), .B(n3981), .Z(n3979) );
  XOR U7570 ( .A(DB[500]), .B(DB[485]), .Z(n3981) );
  AND U7571 ( .A(n894), .B(n3982), .Z(n3980) );
  XOR U7572 ( .A(n3983), .B(n3984), .Z(n3982) );
  XOR U7573 ( .A(DB[485]), .B(DB[470]), .Z(n3984) );
  AND U7574 ( .A(n898), .B(n3985), .Z(n3983) );
  XOR U7575 ( .A(n3986), .B(n3987), .Z(n3985) );
  XOR U7576 ( .A(DB[470]), .B(DB[455]), .Z(n3987) );
  AND U7577 ( .A(n902), .B(n3988), .Z(n3986) );
  XOR U7578 ( .A(n3989), .B(n3990), .Z(n3988) );
  XOR U7579 ( .A(DB[455]), .B(DB[440]), .Z(n3990) );
  AND U7580 ( .A(n906), .B(n3991), .Z(n3989) );
  XOR U7581 ( .A(n3992), .B(n3993), .Z(n3991) );
  XOR U7582 ( .A(DB[440]), .B(DB[425]), .Z(n3993) );
  AND U7583 ( .A(n910), .B(n3994), .Z(n3992) );
  XOR U7584 ( .A(n3995), .B(n3996), .Z(n3994) );
  XOR U7585 ( .A(DB[425]), .B(DB[410]), .Z(n3996) );
  AND U7586 ( .A(n914), .B(n3997), .Z(n3995) );
  XOR U7587 ( .A(n3998), .B(n3999), .Z(n3997) );
  XOR U7588 ( .A(DB[410]), .B(DB[395]), .Z(n3999) );
  AND U7589 ( .A(n918), .B(n4000), .Z(n3998) );
  XOR U7590 ( .A(n4001), .B(n4002), .Z(n4000) );
  XOR U7591 ( .A(DB[395]), .B(DB[380]), .Z(n4002) );
  AND U7592 ( .A(n922), .B(n4003), .Z(n4001) );
  XOR U7593 ( .A(n4004), .B(n4005), .Z(n4003) );
  XOR U7594 ( .A(DB[380]), .B(DB[365]), .Z(n4005) );
  AND U7595 ( .A(n926), .B(n4006), .Z(n4004) );
  XOR U7596 ( .A(n4007), .B(n4008), .Z(n4006) );
  XOR U7597 ( .A(DB[365]), .B(DB[350]), .Z(n4008) );
  AND U7598 ( .A(n930), .B(n4009), .Z(n4007) );
  XOR U7599 ( .A(n4010), .B(n4011), .Z(n4009) );
  XOR U7600 ( .A(DB[350]), .B(DB[335]), .Z(n4011) );
  AND U7601 ( .A(n934), .B(n4012), .Z(n4010) );
  XOR U7602 ( .A(n4013), .B(n4014), .Z(n4012) );
  XOR U7603 ( .A(DB[335]), .B(DB[320]), .Z(n4014) );
  AND U7604 ( .A(n938), .B(n4015), .Z(n4013) );
  XOR U7605 ( .A(n4016), .B(n4017), .Z(n4015) );
  XOR U7606 ( .A(DB[320]), .B(DB[305]), .Z(n4017) );
  AND U7607 ( .A(n942), .B(n4018), .Z(n4016) );
  XOR U7608 ( .A(n4019), .B(n4020), .Z(n4018) );
  XOR U7609 ( .A(DB[305]), .B(DB[290]), .Z(n4020) );
  AND U7610 ( .A(n946), .B(n4021), .Z(n4019) );
  XOR U7611 ( .A(n4022), .B(n4023), .Z(n4021) );
  XOR U7612 ( .A(DB[290]), .B(DB[275]), .Z(n4023) );
  AND U7613 ( .A(n950), .B(n4024), .Z(n4022) );
  XOR U7614 ( .A(n4025), .B(n4026), .Z(n4024) );
  XOR U7615 ( .A(DB[275]), .B(DB[260]), .Z(n4026) );
  AND U7616 ( .A(n954), .B(n4027), .Z(n4025) );
  XOR U7617 ( .A(n4028), .B(n4029), .Z(n4027) );
  XOR U7618 ( .A(DB[260]), .B(DB[245]), .Z(n4029) );
  AND U7619 ( .A(n958), .B(n4030), .Z(n4028) );
  XOR U7620 ( .A(n4031), .B(n4032), .Z(n4030) );
  XOR U7621 ( .A(DB[245]), .B(DB[230]), .Z(n4032) );
  AND U7622 ( .A(n962), .B(n4033), .Z(n4031) );
  XOR U7623 ( .A(n4034), .B(n4035), .Z(n4033) );
  XOR U7624 ( .A(DB[230]), .B(DB[215]), .Z(n4035) );
  AND U7625 ( .A(n966), .B(n4036), .Z(n4034) );
  XOR U7626 ( .A(n4037), .B(n4038), .Z(n4036) );
  XOR U7627 ( .A(DB[215]), .B(DB[200]), .Z(n4038) );
  AND U7628 ( .A(n970), .B(n4039), .Z(n4037) );
  XOR U7629 ( .A(n4040), .B(n4041), .Z(n4039) );
  XOR U7630 ( .A(DB[200]), .B(DB[185]), .Z(n4041) );
  AND U7631 ( .A(n974), .B(n4042), .Z(n4040) );
  XOR U7632 ( .A(n4043), .B(n4044), .Z(n4042) );
  XOR U7633 ( .A(DB[185]), .B(DB[170]), .Z(n4044) );
  AND U7634 ( .A(n978), .B(n4045), .Z(n4043) );
  XOR U7635 ( .A(n4046), .B(n4047), .Z(n4045) );
  XOR U7636 ( .A(DB[170]), .B(DB[155]), .Z(n4047) );
  AND U7637 ( .A(n982), .B(n4048), .Z(n4046) );
  XOR U7638 ( .A(n4049), .B(n4050), .Z(n4048) );
  XOR U7639 ( .A(DB[155]), .B(DB[140]), .Z(n4050) );
  AND U7640 ( .A(n986), .B(n4051), .Z(n4049) );
  XOR U7641 ( .A(n4052), .B(n4053), .Z(n4051) );
  XOR U7642 ( .A(DB[140]), .B(DB[125]), .Z(n4053) );
  AND U7643 ( .A(n990), .B(n4054), .Z(n4052) );
  XOR U7644 ( .A(n4055), .B(n4056), .Z(n4054) );
  XOR U7645 ( .A(DB[125]), .B(DB[110]), .Z(n4056) );
  AND U7646 ( .A(n994), .B(n4057), .Z(n4055) );
  XOR U7647 ( .A(n4058), .B(n4059), .Z(n4057) );
  XOR U7648 ( .A(DB[95]), .B(DB[110]), .Z(n4059) );
  AND U7649 ( .A(n998), .B(n4060), .Z(n4058) );
  XOR U7650 ( .A(n4061), .B(n4062), .Z(n4060) );
  XOR U7651 ( .A(DB[95]), .B(DB[80]), .Z(n4062) );
  AND U7652 ( .A(n1002), .B(n4063), .Z(n4061) );
  XOR U7653 ( .A(n4064), .B(n4065), .Z(n4063) );
  XOR U7654 ( .A(DB[80]), .B(DB[65]), .Z(n4065) );
  AND U7655 ( .A(n1006), .B(n4066), .Z(n4064) );
  XOR U7656 ( .A(n4067), .B(n4068), .Z(n4066) );
  XOR U7657 ( .A(DB[65]), .B(DB[50]), .Z(n4068) );
  AND U7658 ( .A(n1010), .B(n4069), .Z(n4067) );
  XOR U7659 ( .A(n4070), .B(n4071), .Z(n4069) );
  XOR U7660 ( .A(DB[50]), .B(DB[35]), .Z(n4071) );
  AND U7661 ( .A(n1014), .B(n4072), .Z(n4070) );
  XOR U7662 ( .A(n4073), .B(n4074), .Z(n4072) );
  XOR U7663 ( .A(DB[35]), .B(DB[20]), .Z(n4074) );
  AND U7664 ( .A(n1018), .B(n4075), .Z(n4073) );
  XOR U7665 ( .A(DB[5]), .B(DB[20]), .Z(n4075) );
  XOR U7666 ( .A(DB[3829]), .B(n4076), .Z(min_val_out[4]) );
  AND U7667 ( .A(n2), .B(n4077), .Z(n4076) );
  XOR U7668 ( .A(n4078), .B(n4079), .Z(n4077) );
  XOR U7669 ( .A(DB[3829]), .B(DB[3814]), .Z(n4079) );
  AND U7670 ( .A(n6), .B(n4080), .Z(n4078) );
  XOR U7671 ( .A(n4081), .B(n4082), .Z(n4080) );
  XOR U7672 ( .A(DB[3814]), .B(DB[3799]), .Z(n4082) );
  AND U7673 ( .A(n10), .B(n4083), .Z(n4081) );
  XOR U7674 ( .A(n4084), .B(n4085), .Z(n4083) );
  XOR U7675 ( .A(DB[3799]), .B(DB[3784]), .Z(n4085) );
  AND U7676 ( .A(n14), .B(n4086), .Z(n4084) );
  XOR U7677 ( .A(n4087), .B(n4088), .Z(n4086) );
  XOR U7678 ( .A(DB[3784]), .B(DB[3769]), .Z(n4088) );
  AND U7679 ( .A(n18), .B(n4089), .Z(n4087) );
  XOR U7680 ( .A(n4090), .B(n4091), .Z(n4089) );
  XOR U7681 ( .A(DB[3769]), .B(DB[3754]), .Z(n4091) );
  AND U7682 ( .A(n22), .B(n4092), .Z(n4090) );
  XOR U7683 ( .A(n4093), .B(n4094), .Z(n4092) );
  XOR U7684 ( .A(DB[3754]), .B(DB[3739]), .Z(n4094) );
  AND U7685 ( .A(n26), .B(n4095), .Z(n4093) );
  XOR U7686 ( .A(n4096), .B(n4097), .Z(n4095) );
  XOR U7687 ( .A(DB[3739]), .B(DB[3724]), .Z(n4097) );
  AND U7688 ( .A(n30), .B(n4098), .Z(n4096) );
  XOR U7689 ( .A(n4099), .B(n4100), .Z(n4098) );
  XOR U7690 ( .A(DB[3724]), .B(DB[3709]), .Z(n4100) );
  AND U7691 ( .A(n34), .B(n4101), .Z(n4099) );
  XOR U7692 ( .A(n4102), .B(n4103), .Z(n4101) );
  XOR U7693 ( .A(DB[3709]), .B(DB[3694]), .Z(n4103) );
  AND U7694 ( .A(n38), .B(n4104), .Z(n4102) );
  XOR U7695 ( .A(n4105), .B(n4106), .Z(n4104) );
  XOR U7696 ( .A(DB[3694]), .B(DB[3679]), .Z(n4106) );
  AND U7697 ( .A(n42), .B(n4107), .Z(n4105) );
  XOR U7698 ( .A(n4108), .B(n4109), .Z(n4107) );
  XOR U7699 ( .A(DB[3679]), .B(DB[3664]), .Z(n4109) );
  AND U7700 ( .A(n46), .B(n4110), .Z(n4108) );
  XOR U7701 ( .A(n4111), .B(n4112), .Z(n4110) );
  XOR U7702 ( .A(DB[3664]), .B(DB[3649]), .Z(n4112) );
  AND U7703 ( .A(n50), .B(n4113), .Z(n4111) );
  XOR U7704 ( .A(n4114), .B(n4115), .Z(n4113) );
  XOR U7705 ( .A(DB[3649]), .B(DB[3634]), .Z(n4115) );
  AND U7706 ( .A(n54), .B(n4116), .Z(n4114) );
  XOR U7707 ( .A(n4117), .B(n4118), .Z(n4116) );
  XOR U7708 ( .A(DB[3634]), .B(DB[3619]), .Z(n4118) );
  AND U7709 ( .A(n58), .B(n4119), .Z(n4117) );
  XOR U7710 ( .A(n4120), .B(n4121), .Z(n4119) );
  XOR U7711 ( .A(DB[3619]), .B(DB[3604]), .Z(n4121) );
  AND U7712 ( .A(n62), .B(n4122), .Z(n4120) );
  XOR U7713 ( .A(n4123), .B(n4124), .Z(n4122) );
  XOR U7714 ( .A(DB[3604]), .B(DB[3589]), .Z(n4124) );
  AND U7715 ( .A(n66), .B(n4125), .Z(n4123) );
  XOR U7716 ( .A(n4126), .B(n4127), .Z(n4125) );
  XOR U7717 ( .A(DB[3589]), .B(DB[3574]), .Z(n4127) );
  AND U7718 ( .A(n70), .B(n4128), .Z(n4126) );
  XOR U7719 ( .A(n4129), .B(n4130), .Z(n4128) );
  XOR U7720 ( .A(DB[3574]), .B(DB[3559]), .Z(n4130) );
  AND U7721 ( .A(n74), .B(n4131), .Z(n4129) );
  XOR U7722 ( .A(n4132), .B(n4133), .Z(n4131) );
  XOR U7723 ( .A(DB[3559]), .B(DB[3544]), .Z(n4133) );
  AND U7724 ( .A(n78), .B(n4134), .Z(n4132) );
  XOR U7725 ( .A(n4135), .B(n4136), .Z(n4134) );
  XOR U7726 ( .A(DB[3544]), .B(DB[3529]), .Z(n4136) );
  AND U7727 ( .A(n82), .B(n4137), .Z(n4135) );
  XOR U7728 ( .A(n4138), .B(n4139), .Z(n4137) );
  XOR U7729 ( .A(DB[3529]), .B(DB[3514]), .Z(n4139) );
  AND U7730 ( .A(n86), .B(n4140), .Z(n4138) );
  XOR U7731 ( .A(n4141), .B(n4142), .Z(n4140) );
  XOR U7732 ( .A(DB[3514]), .B(DB[3499]), .Z(n4142) );
  AND U7733 ( .A(n90), .B(n4143), .Z(n4141) );
  XOR U7734 ( .A(n4144), .B(n4145), .Z(n4143) );
  XOR U7735 ( .A(DB[3499]), .B(DB[3484]), .Z(n4145) );
  AND U7736 ( .A(n94), .B(n4146), .Z(n4144) );
  XOR U7737 ( .A(n4147), .B(n4148), .Z(n4146) );
  XOR U7738 ( .A(DB[3484]), .B(DB[3469]), .Z(n4148) );
  AND U7739 ( .A(n98), .B(n4149), .Z(n4147) );
  XOR U7740 ( .A(n4150), .B(n4151), .Z(n4149) );
  XOR U7741 ( .A(DB[3469]), .B(DB[3454]), .Z(n4151) );
  AND U7742 ( .A(n102), .B(n4152), .Z(n4150) );
  XOR U7743 ( .A(n4153), .B(n4154), .Z(n4152) );
  XOR U7744 ( .A(DB[3454]), .B(DB[3439]), .Z(n4154) );
  AND U7745 ( .A(n106), .B(n4155), .Z(n4153) );
  XOR U7746 ( .A(n4156), .B(n4157), .Z(n4155) );
  XOR U7747 ( .A(DB[3439]), .B(DB[3424]), .Z(n4157) );
  AND U7748 ( .A(n110), .B(n4158), .Z(n4156) );
  XOR U7749 ( .A(n4159), .B(n4160), .Z(n4158) );
  XOR U7750 ( .A(DB[3424]), .B(DB[3409]), .Z(n4160) );
  AND U7751 ( .A(n114), .B(n4161), .Z(n4159) );
  XOR U7752 ( .A(n4162), .B(n4163), .Z(n4161) );
  XOR U7753 ( .A(DB[3409]), .B(DB[3394]), .Z(n4163) );
  AND U7754 ( .A(n118), .B(n4164), .Z(n4162) );
  XOR U7755 ( .A(n4165), .B(n4166), .Z(n4164) );
  XOR U7756 ( .A(DB[3394]), .B(DB[3379]), .Z(n4166) );
  AND U7757 ( .A(n122), .B(n4167), .Z(n4165) );
  XOR U7758 ( .A(n4168), .B(n4169), .Z(n4167) );
  XOR U7759 ( .A(DB[3379]), .B(DB[3364]), .Z(n4169) );
  AND U7760 ( .A(n126), .B(n4170), .Z(n4168) );
  XOR U7761 ( .A(n4171), .B(n4172), .Z(n4170) );
  XOR U7762 ( .A(DB[3364]), .B(DB[3349]), .Z(n4172) );
  AND U7763 ( .A(n130), .B(n4173), .Z(n4171) );
  XOR U7764 ( .A(n4174), .B(n4175), .Z(n4173) );
  XOR U7765 ( .A(DB[3349]), .B(DB[3334]), .Z(n4175) );
  AND U7766 ( .A(n134), .B(n4176), .Z(n4174) );
  XOR U7767 ( .A(n4177), .B(n4178), .Z(n4176) );
  XOR U7768 ( .A(DB[3334]), .B(DB[3319]), .Z(n4178) );
  AND U7769 ( .A(n138), .B(n4179), .Z(n4177) );
  XOR U7770 ( .A(n4180), .B(n4181), .Z(n4179) );
  XOR U7771 ( .A(DB[3319]), .B(DB[3304]), .Z(n4181) );
  AND U7772 ( .A(n142), .B(n4182), .Z(n4180) );
  XOR U7773 ( .A(n4183), .B(n4184), .Z(n4182) );
  XOR U7774 ( .A(DB[3304]), .B(DB[3289]), .Z(n4184) );
  AND U7775 ( .A(n146), .B(n4185), .Z(n4183) );
  XOR U7776 ( .A(n4186), .B(n4187), .Z(n4185) );
  XOR U7777 ( .A(DB[3289]), .B(DB[3274]), .Z(n4187) );
  AND U7778 ( .A(n150), .B(n4188), .Z(n4186) );
  XOR U7779 ( .A(n4189), .B(n4190), .Z(n4188) );
  XOR U7780 ( .A(DB[3274]), .B(DB[3259]), .Z(n4190) );
  AND U7781 ( .A(n154), .B(n4191), .Z(n4189) );
  XOR U7782 ( .A(n4192), .B(n4193), .Z(n4191) );
  XOR U7783 ( .A(DB[3259]), .B(DB[3244]), .Z(n4193) );
  AND U7784 ( .A(n158), .B(n4194), .Z(n4192) );
  XOR U7785 ( .A(n4195), .B(n4196), .Z(n4194) );
  XOR U7786 ( .A(DB[3244]), .B(DB[3229]), .Z(n4196) );
  AND U7787 ( .A(n162), .B(n4197), .Z(n4195) );
  XOR U7788 ( .A(n4198), .B(n4199), .Z(n4197) );
  XOR U7789 ( .A(DB[3229]), .B(DB[3214]), .Z(n4199) );
  AND U7790 ( .A(n166), .B(n4200), .Z(n4198) );
  XOR U7791 ( .A(n4201), .B(n4202), .Z(n4200) );
  XOR U7792 ( .A(DB[3214]), .B(DB[3199]), .Z(n4202) );
  AND U7793 ( .A(n170), .B(n4203), .Z(n4201) );
  XOR U7794 ( .A(n4204), .B(n4205), .Z(n4203) );
  XOR U7795 ( .A(DB[3199]), .B(DB[3184]), .Z(n4205) );
  AND U7796 ( .A(n174), .B(n4206), .Z(n4204) );
  XOR U7797 ( .A(n4207), .B(n4208), .Z(n4206) );
  XOR U7798 ( .A(DB[3184]), .B(DB[3169]), .Z(n4208) );
  AND U7799 ( .A(n178), .B(n4209), .Z(n4207) );
  XOR U7800 ( .A(n4210), .B(n4211), .Z(n4209) );
  XOR U7801 ( .A(DB[3169]), .B(DB[3154]), .Z(n4211) );
  AND U7802 ( .A(n182), .B(n4212), .Z(n4210) );
  XOR U7803 ( .A(n4213), .B(n4214), .Z(n4212) );
  XOR U7804 ( .A(DB[3154]), .B(DB[3139]), .Z(n4214) );
  AND U7805 ( .A(n186), .B(n4215), .Z(n4213) );
  XOR U7806 ( .A(n4216), .B(n4217), .Z(n4215) );
  XOR U7807 ( .A(DB[3139]), .B(DB[3124]), .Z(n4217) );
  AND U7808 ( .A(n190), .B(n4218), .Z(n4216) );
  XOR U7809 ( .A(n4219), .B(n4220), .Z(n4218) );
  XOR U7810 ( .A(DB[3124]), .B(DB[3109]), .Z(n4220) );
  AND U7811 ( .A(n194), .B(n4221), .Z(n4219) );
  XOR U7812 ( .A(n4222), .B(n4223), .Z(n4221) );
  XOR U7813 ( .A(DB[3109]), .B(DB[3094]), .Z(n4223) );
  AND U7814 ( .A(n198), .B(n4224), .Z(n4222) );
  XOR U7815 ( .A(n4225), .B(n4226), .Z(n4224) );
  XOR U7816 ( .A(DB[3094]), .B(DB[3079]), .Z(n4226) );
  AND U7817 ( .A(n202), .B(n4227), .Z(n4225) );
  XOR U7818 ( .A(n4228), .B(n4229), .Z(n4227) );
  XOR U7819 ( .A(DB[3079]), .B(DB[3064]), .Z(n4229) );
  AND U7820 ( .A(n206), .B(n4230), .Z(n4228) );
  XOR U7821 ( .A(n4231), .B(n4232), .Z(n4230) );
  XOR U7822 ( .A(DB[3064]), .B(DB[3049]), .Z(n4232) );
  AND U7823 ( .A(n210), .B(n4233), .Z(n4231) );
  XOR U7824 ( .A(n4234), .B(n4235), .Z(n4233) );
  XOR U7825 ( .A(DB[3049]), .B(DB[3034]), .Z(n4235) );
  AND U7826 ( .A(n214), .B(n4236), .Z(n4234) );
  XOR U7827 ( .A(n4237), .B(n4238), .Z(n4236) );
  XOR U7828 ( .A(DB[3034]), .B(DB[3019]), .Z(n4238) );
  AND U7829 ( .A(n218), .B(n4239), .Z(n4237) );
  XOR U7830 ( .A(n4240), .B(n4241), .Z(n4239) );
  XOR U7831 ( .A(DB[3019]), .B(DB[3004]), .Z(n4241) );
  AND U7832 ( .A(n222), .B(n4242), .Z(n4240) );
  XOR U7833 ( .A(n4243), .B(n4244), .Z(n4242) );
  XOR U7834 ( .A(DB[3004]), .B(DB[2989]), .Z(n4244) );
  AND U7835 ( .A(n226), .B(n4245), .Z(n4243) );
  XOR U7836 ( .A(n4246), .B(n4247), .Z(n4245) );
  XOR U7837 ( .A(DB[2989]), .B(DB[2974]), .Z(n4247) );
  AND U7838 ( .A(n230), .B(n4248), .Z(n4246) );
  XOR U7839 ( .A(n4249), .B(n4250), .Z(n4248) );
  XOR U7840 ( .A(DB[2974]), .B(DB[2959]), .Z(n4250) );
  AND U7841 ( .A(n234), .B(n4251), .Z(n4249) );
  XOR U7842 ( .A(n4252), .B(n4253), .Z(n4251) );
  XOR U7843 ( .A(DB[2959]), .B(DB[2944]), .Z(n4253) );
  AND U7844 ( .A(n238), .B(n4254), .Z(n4252) );
  XOR U7845 ( .A(n4255), .B(n4256), .Z(n4254) );
  XOR U7846 ( .A(DB[2944]), .B(DB[2929]), .Z(n4256) );
  AND U7847 ( .A(n242), .B(n4257), .Z(n4255) );
  XOR U7848 ( .A(n4258), .B(n4259), .Z(n4257) );
  XOR U7849 ( .A(DB[2929]), .B(DB[2914]), .Z(n4259) );
  AND U7850 ( .A(n246), .B(n4260), .Z(n4258) );
  XOR U7851 ( .A(n4261), .B(n4262), .Z(n4260) );
  XOR U7852 ( .A(DB[2914]), .B(DB[2899]), .Z(n4262) );
  AND U7853 ( .A(n250), .B(n4263), .Z(n4261) );
  XOR U7854 ( .A(n4264), .B(n4265), .Z(n4263) );
  XOR U7855 ( .A(DB[2899]), .B(DB[2884]), .Z(n4265) );
  AND U7856 ( .A(n254), .B(n4266), .Z(n4264) );
  XOR U7857 ( .A(n4267), .B(n4268), .Z(n4266) );
  XOR U7858 ( .A(DB[2884]), .B(DB[2869]), .Z(n4268) );
  AND U7859 ( .A(n258), .B(n4269), .Z(n4267) );
  XOR U7860 ( .A(n4270), .B(n4271), .Z(n4269) );
  XOR U7861 ( .A(DB[2869]), .B(DB[2854]), .Z(n4271) );
  AND U7862 ( .A(n262), .B(n4272), .Z(n4270) );
  XOR U7863 ( .A(n4273), .B(n4274), .Z(n4272) );
  XOR U7864 ( .A(DB[2854]), .B(DB[2839]), .Z(n4274) );
  AND U7865 ( .A(n266), .B(n4275), .Z(n4273) );
  XOR U7866 ( .A(n4276), .B(n4277), .Z(n4275) );
  XOR U7867 ( .A(DB[2839]), .B(DB[2824]), .Z(n4277) );
  AND U7868 ( .A(n270), .B(n4278), .Z(n4276) );
  XOR U7869 ( .A(n4279), .B(n4280), .Z(n4278) );
  XOR U7870 ( .A(DB[2824]), .B(DB[2809]), .Z(n4280) );
  AND U7871 ( .A(n274), .B(n4281), .Z(n4279) );
  XOR U7872 ( .A(n4282), .B(n4283), .Z(n4281) );
  XOR U7873 ( .A(DB[2809]), .B(DB[2794]), .Z(n4283) );
  AND U7874 ( .A(n278), .B(n4284), .Z(n4282) );
  XOR U7875 ( .A(n4285), .B(n4286), .Z(n4284) );
  XOR U7876 ( .A(DB[2794]), .B(DB[2779]), .Z(n4286) );
  AND U7877 ( .A(n282), .B(n4287), .Z(n4285) );
  XOR U7878 ( .A(n4288), .B(n4289), .Z(n4287) );
  XOR U7879 ( .A(DB[2779]), .B(DB[2764]), .Z(n4289) );
  AND U7880 ( .A(n286), .B(n4290), .Z(n4288) );
  XOR U7881 ( .A(n4291), .B(n4292), .Z(n4290) );
  XOR U7882 ( .A(DB[2764]), .B(DB[2749]), .Z(n4292) );
  AND U7883 ( .A(n290), .B(n4293), .Z(n4291) );
  XOR U7884 ( .A(n4294), .B(n4295), .Z(n4293) );
  XOR U7885 ( .A(DB[2749]), .B(DB[2734]), .Z(n4295) );
  AND U7886 ( .A(n294), .B(n4296), .Z(n4294) );
  XOR U7887 ( .A(n4297), .B(n4298), .Z(n4296) );
  XOR U7888 ( .A(DB[2734]), .B(DB[2719]), .Z(n4298) );
  AND U7889 ( .A(n298), .B(n4299), .Z(n4297) );
  XOR U7890 ( .A(n4300), .B(n4301), .Z(n4299) );
  XOR U7891 ( .A(DB[2719]), .B(DB[2704]), .Z(n4301) );
  AND U7892 ( .A(n302), .B(n4302), .Z(n4300) );
  XOR U7893 ( .A(n4303), .B(n4304), .Z(n4302) );
  XOR U7894 ( .A(DB[2704]), .B(DB[2689]), .Z(n4304) );
  AND U7895 ( .A(n306), .B(n4305), .Z(n4303) );
  XOR U7896 ( .A(n4306), .B(n4307), .Z(n4305) );
  XOR U7897 ( .A(DB[2689]), .B(DB[2674]), .Z(n4307) );
  AND U7898 ( .A(n310), .B(n4308), .Z(n4306) );
  XOR U7899 ( .A(n4309), .B(n4310), .Z(n4308) );
  XOR U7900 ( .A(DB[2674]), .B(DB[2659]), .Z(n4310) );
  AND U7901 ( .A(n314), .B(n4311), .Z(n4309) );
  XOR U7902 ( .A(n4312), .B(n4313), .Z(n4311) );
  XOR U7903 ( .A(DB[2659]), .B(DB[2644]), .Z(n4313) );
  AND U7904 ( .A(n318), .B(n4314), .Z(n4312) );
  XOR U7905 ( .A(n4315), .B(n4316), .Z(n4314) );
  XOR U7906 ( .A(DB[2644]), .B(DB[2629]), .Z(n4316) );
  AND U7907 ( .A(n322), .B(n4317), .Z(n4315) );
  XOR U7908 ( .A(n4318), .B(n4319), .Z(n4317) );
  XOR U7909 ( .A(DB[2629]), .B(DB[2614]), .Z(n4319) );
  AND U7910 ( .A(n326), .B(n4320), .Z(n4318) );
  XOR U7911 ( .A(n4321), .B(n4322), .Z(n4320) );
  XOR U7912 ( .A(DB[2614]), .B(DB[2599]), .Z(n4322) );
  AND U7913 ( .A(n330), .B(n4323), .Z(n4321) );
  XOR U7914 ( .A(n4324), .B(n4325), .Z(n4323) );
  XOR U7915 ( .A(DB[2599]), .B(DB[2584]), .Z(n4325) );
  AND U7916 ( .A(n334), .B(n4326), .Z(n4324) );
  XOR U7917 ( .A(n4327), .B(n4328), .Z(n4326) );
  XOR U7918 ( .A(DB[2584]), .B(DB[2569]), .Z(n4328) );
  AND U7919 ( .A(n338), .B(n4329), .Z(n4327) );
  XOR U7920 ( .A(n4330), .B(n4331), .Z(n4329) );
  XOR U7921 ( .A(DB[2569]), .B(DB[2554]), .Z(n4331) );
  AND U7922 ( .A(n342), .B(n4332), .Z(n4330) );
  XOR U7923 ( .A(n4333), .B(n4334), .Z(n4332) );
  XOR U7924 ( .A(DB[2554]), .B(DB[2539]), .Z(n4334) );
  AND U7925 ( .A(n346), .B(n4335), .Z(n4333) );
  XOR U7926 ( .A(n4336), .B(n4337), .Z(n4335) );
  XOR U7927 ( .A(DB[2539]), .B(DB[2524]), .Z(n4337) );
  AND U7928 ( .A(n350), .B(n4338), .Z(n4336) );
  XOR U7929 ( .A(n4339), .B(n4340), .Z(n4338) );
  XOR U7930 ( .A(DB[2524]), .B(DB[2509]), .Z(n4340) );
  AND U7931 ( .A(n354), .B(n4341), .Z(n4339) );
  XOR U7932 ( .A(n4342), .B(n4343), .Z(n4341) );
  XOR U7933 ( .A(DB[2509]), .B(DB[2494]), .Z(n4343) );
  AND U7934 ( .A(n358), .B(n4344), .Z(n4342) );
  XOR U7935 ( .A(n4345), .B(n4346), .Z(n4344) );
  XOR U7936 ( .A(DB[2494]), .B(DB[2479]), .Z(n4346) );
  AND U7937 ( .A(n362), .B(n4347), .Z(n4345) );
  XOR U7938 ( .A(n4348), .B(n4349), .Z(n4347) );
  XOR U7939 ( .A(DB[2479]), .B(DB[2464]), .Z(n4349) );
  AND U7940 ( .A(n366), .B(n4350), .Z(n4348) );
  XOR U7941 ( .A(n4351), .B(n4352), .Z(n4350) );
  XOR U7942 ( .A(DB[2464]), .B(DB[2449]), .Z(n4352) );
  AND U7943 ( .A(n370), .B(n4353), .Z(n4351) );
  XOR U7944 ( .A(n4354), .B(n4355), .Z(n4353) );
  XOR U7945 ( .A(DB[2449]), .B(DB[2434]), .Z(n4355) );
  AND U7946 ( .A(n374), .B(n4356), .Z(n4354) );
  XOR U7947 ( .A(n4357), .B(n4358), .Z(n4356) );
  XOR U7948 ( .A(DB[2434]), .B(DB[2419]), .Z(n4358) );
  AND U7949 ( .A(n378), .B(n4359), .Z(n4357) );
  XOR U7950 ( .A(n4360), .B(n4361), .Z(n4359) );
  XOR U7951 ( .A(DB[2419]), .B(DB[2404]), .Z(n4361) );
  AND U7952 ( .A(n382), .B(n4362), .Z(n4360) );
  XOR U7953 ( .A(n4363), .B(n4364), .Z(n4362) );
  XOR U7954 ( .A(DB[2404]), .B(DB[2389]), .Z(n4364) );
  AND U7955 ( .A(n386), .B(n4365), .Z(n4363) );
  XOR U7956 ( .A(n4366), .B(n4367), .Z(n4365) );
  XOR U7957 ( .A(DB[2389]), .B(DB[2374]), .Z(n4367) );
  AND U7958 ( .A(n390), .B(n4368), .Z(n4366) );
  XOR U7959 ( .A(n4369), .B(n4370), .Z(n4368) );
  XOR U7960 ( .A(DB[2374]), .B(DB[2359]), .Z(n4370) );
  AND U7961 ( .A(n394), .B(n4371), .Z(n4369) );
  XOR U7962 ( .A(n4372), .B(n4373), .Z(n4371) );
  XOR U7963 ( .A(DB[2359]), .B(DB[2344]), .Z(n4373) );
  AND U7964 ( .A(n398), .B(n4374), .Z(n4372) );
  XOR U7965 ( .A(n4375), .B(n4376), .Z(n4374) );
  XOR U7966 ( .A(DB[2344]), .B(DB[2329]), .Z(n4376) );
  AND U7967 ( .A(n402), .B(n4377), .Z(n4375) );
  XOR U7968 ( .A(n4378), .B(n4379), .Z(n4377) );
  XOR U7969 ( .A(DB[2329]), .B(DB[2314]), .Z(n4379) );
  AND U7970 ( .A(n406), .B(n4380), .Z(n4378) );
  XOR U7971 ( .A(n4381), .B(n4382), .Z(n4380) );
  XOR U7972 ( .A(DB[2314]), .B(DB[2299]), .Z(n4382) );
  AND U7973 ( .A(n410), .B(n4383), .Z(n4381) );
  XOR U7974 ( .A(n4384), .B(n4385), .Z(n4383) );
  XOR U7975 ( .A(DB[2299]), .B(DB[2284]), .Z(n4385) );
  AND U7976 ( .A(n414), .B(n4386), .Z(n4384) );
  XOR U7977 ( .A(n4387), .B(n4388), .Z(n4386) );
  XOR U7978 ( .A(DB[2284]), .B(DB[2269]), .Z(n4388) );
  AND U7979 ( .A(n418), .B(n4389), .Z(n4387) );
  XOR U7980 ( .A(n4390), .B(n4391), .Z(n4389) );
  XOR U7981 ( .A(DB[2269]), .B(DB[2254]), .Z(n4391) );
  AND U7982 ( .A(n422), .B(n4392), .Z(n4390) );
  XOR U7983 ( .A(n4393), .B(n4394), .Z(n4392) );
  XOR U7984 ( .A(DB[2254]), .B(DB[2239]), .Z(n4394) );
  AND U7985 ( .A(n426), .B(n4395), .Z(n4393) );
  XOR U7986 ( .A(n4396), .B(n4397), .Z(n4395) );
  XOR U7987 ( .A(DB[2239]), .B(DB[2224]), .Z(n4397) );
  AND U7988 ( .A(n430), .B(n4398), .Z(n4396) );
  XOR U7989 ( .A(n4399), .B(n4400), .Z(n4398) );
  XOR U7990 ( .A(DB[2224]), .B(DB[2209]), .Z(n4400) );
  AND U7991 ( .A(n434), .B(n4401), .Z(n4399) );
  XOR U7992 ( .A(n4402), .B(n4403), .Z(n4401) );
  XOR U7993 ( .A(DB[2209]), .B(DB[2194]), .Z(n4403) );
  AND U7994 ( .A(n438), .B(n4404), .Z(n4402) );
  XOR U7995 ( .A(n4405), .B(n4406), .Z(n4404) );
  XOR U7996 ( .A(DB[2194]), .B(DB[2179]), .Z(n4406) );
  AND U7997 ( .A(n442), .B(n4407), .Z(n4405) );
  XOR U7998 ( .A(n4408), .B(n4409), .Z(n4407) );
  XOR U7999 ( .A(DB[2179]), .B(DB[2164]), .Z(n4409) );
  AND U8000 ( .A(n446), .B(n4410), .Z(n4408) );
  XOR U8001 ( .A(n4411), .B(n4412), .Z(n4410) );
  XOR U8002 ( .A(DB[2164]), .B(DB[2149]), .Z(n4412) );
  AND U8003 ( .A(n450), .B(n4413), .Z(n4411) );
  XOR U8004 ( .A(n4414), .B(n4415), .Z(n4413) );
  XOR U8005 ( .A(DB[2149]), .B(DB[2134]), .Z(n4415) );
  AND U8006 ( .A(n454), .B(n4416), .Z(n4414) );
  XOR U8007 ( .A(n4417), .B(n4418), .Z(n4416) );
  XOR U8008 ( .A(DB[2134]), .B(DB[2119]), .Z(n4418) );
  AND U8009 ( .A(n458), .B(n4419), .Z(n4417) );
  XOR U8010 ( .A(n4420), .B(n4421), .Z(n4419) );
  XOR U8011 ( .A(DB[2119]), .B(DB[2104]), .Z(n4421) );
  AND U8012 ( .A(n462), .B(n4422), .Z(n4420) );
  XOR U8013 ( .A(n4423), .B(n4424), .Z(n4422) );
  XOR U8014 ( .A(DB[2104]), .B(DB[2089]), .Z(n4424) );
  AND U8015 ( .A(n466), .B(n4425), .Z(n4423) );
  XOR U8016 ( .A(n4426), .B(n4427), .Z(n4425) );
  XOR U8017 ( .A(DB[2089]), .B(DB[2074]), .Z(n4427) );
  AND U8018 ( .A(n470), .B(n4428), .Z(n4426) );
  XOR U8019 ( .A(n4429), .B(n4430), .Z(n4428) );
  XOR U8020 ( .A(DB[2074]), .B(DB[2059]), .Z(n4430) );
  AND U8021 ( .A(n474), .B(n4431), .Z(n4429) );
  XOR U8022 ( .A(n4432), .B(n4433), .Z(n4431) );
  XOR U8023 ( .A(DB[2059]), .B(DB[2044]), .Z(n4433) );
  AND U8024 ( .A(n478), .B(n4434), .Z(n4432) );
  XOR U8025 ( .A(n4435), .B(n4436), .Z(n4434) );
  XOR U8026 ( .A(DB[2044]), .B(DB[2029]), .Z(n4436) );
  AND U8027 ( .A(n482), .B(n4437), .Z(n4435) );
  XOR U8028 ( .A(n4438), .B(n4439), .Z(n4437) );
  XOR U8029 ( .A(DB[2029]), .B(DB[2014]), .Z(n4439) );
  AND U8030 ( .A(n486), .B(n4440), .Z(n4438) );
  XOR U8031 ( .A(n4441), .B(n4442), .Z(n4440) );
  XOR U8032 ( .A(DB[2014]), .B(DB[1999]), .Z(n4442) );
  AND U8033 ( .A(n490), .B(n4443), .Z(n4441) );
  XOR U8034 ( .A(n4444), .B(n4445), .Z(n4443) );
  XOR U8035 ( .A(DB[1999]), .B(DB[1984]), .Z(n4445) );
  AND U8036 ( .A(n494), .B(n4446), .Z(n4444) );
  XOR U8037 ( .A(n4447), .B(n4448), .Z(n4446) );
  XOR U8038 ( .A(DB[1984]), .B(DB[1969]), .Z(n4448) );
  AND U8039 ( .A(n498), .B(n4449), .Z(n4447) );
  XOR U8040 ( .A(n4450), .B(n4451), .Z(n4449) );
  XOR U8041 ( .A(DB[1969]), .B(DB[1954]), .Z(n4451) );
  AND U8042 ( .A(n502), .B(n4452), .Z(n4450) );
  XOR U8043 ( .A(n4453), .B(n4454), .Z(n4452) );
  XOR U8044 ( .A(DB[1954]), .B(DB[1939]), .Z(n4454) );
  AND U8045 ( .A(n506), .B(n4455), .Z(n4453) );
  XOR U8046 ( .A(n4456), .B(n4457), .Z(n4455) );
  XOR U8047 ( .A(DB[1939]), .B(DB[1924]), .Z(n4457) );
  AND U8048 ( .A(n510), .B(n4458), .Z(n4456) );
  XOR U8049 ( .A(n4459), .B(n4460), .Z(n4458) );
  XOR U8050 ( .A(DB[1924]), .B(DB[1909]), .Z(n4460) );
  AND U8051 ( .A(n514), .B(n4461), .Z(n4459) );
  XOR U8052 ( .A(n4462), .B(n4463), .Z(n4461) );
  XOR U8053 ( .A(DB[1909]), .B(DB[1894]), .Z(n4463) );
  AND U8054 ( .A(n518), .B(n4464), .Z(n4462) );
  XOR U8055 ( .A(n4465), .B(n4466), .Z(n4464) );
  XOR U8056 ( .A(DB[1894]), .B(DB[1879]), .Z(n4466) );
  AND U8057 ( .A(n522), .B(n4467), .Z(n4465) );
  XOR U8058 ( .A(n4468), .B(n4469), .Z(n4467) );
  XOR U8059 ( .A(DB[1879]), .B(DB[1864]), .Z(n4469) );
  AND U8060 ( .A(n526), .B(n4470), .Z(n4468) );
  XOR U8061 ( .A(n4471), .B(n4472), .Z(n4470) );
  XOR U8062 ( .A(DB[1864]), .B(DB[1849]), .Z(n4472) );
  AND U8063 ( .A(n530), .B(n4473), .Z(n4471) );
  XOR U8064 ( .A(n4474), .B(n4475), .Z(n4473) );
  XOR U8065 ( .A(DB[1849]), .B(DB[1834]), .Z(n4475) );
  AND U8066 ( .A(n534), .B(n4476), .Z(n4474) );
  XOR U8067 ( .A(n4477), .B(n4478), .Z(n4476) );
  XOR U8068 ( .A(DB[1834]), .B(DB[1819]), .Z(n4478) );
  AND U8069 ( .A(n538), .B(n4479), .Z(n4477) );
  XOR U8070 ( .A(n4480), .B(n4481), .Z(n4479) );
  XOR U8071 ( .A(DB[1819]), .B(DB[1804]), .Z(n4481) );
  AND U8072 ( .A(n542), .B(n4482), .Z(n4480) );
  XOR U8073 ( .A(n4483), .B(n4484), .Z(n4482) );
  XOR U8074 ( .A(DB[1804]), .B(DB[1789]), .Z(n4484) );
  AND U8075 ( .A(n546), .B(n4485), .Z(n4483) );
  XOR U8076 ( .A(n4486), .B(n4487), .Z(n4485) );
  XOR U8077 ( .A(DB[1789]), .B(DB[1774]), .Z(n4487) );
  AND U8078 ( .A(n550), .B(n4488), .Z(n4486) );
  XOR U8079 ( .A(n4489), .B(n4490), .Z(n4488) );
  XOR U8080 ( .A(DB[1774]), .B(DB[1759]), .Z(n4490) );
  AND U8081 ( .A(n554), .B(n4491), .Z(n4489) );
  XOR U8082 ( .A(n4492), .B(n4493), .Z(n4491) );
  XOR U8083 ( .A(DB[1759]), .B(DB[1744]), .Z(n4493) );
  AND U8084 ( .A(n558), .B(n4494), .Z(n4492) );
  XOR U8085 ( .A(n4495), .B(n4496), .Z(n4494) );
  XOR U8086 ( .A(DB[1744]), .B(DB[1729]), .Z(n4496) );
  AND U8087 ( .A(n562), .B(n4497), .Z(n4495) );
  XOR U8088 ( .A(n4498), .B(n4499), .Z(n4497) );
  XOR U8089 ( .A(DB[1729]), .B(DB[1714]), .Z(n4499) );
  AND U8090 ( .A(n566), .B(n4500), .Z(n4498) );
  XOR U8091 ( .A(n4501), .B(n4502), .Z(n4500) );
  XOR U8092 ( .A(DB[1714]), .B(DB[1699]), .Z(n4502) );
  AND U8093 ( .A(n570), .B(n4503), .Z(n4501) );
  XOR U8094 ( .A(n4504), .B(n4505), .Z(n4503) );
  XOR U8095 ( .A(DB[1699]), .B(DB[1684]), .Z(n4505) );
  AND U8096 ( .A(n574), .B(n4506), .Z(n4504) );
  XOR U8097 ( .A(n4507), .B(n4508), .Z(n4506) );
  XOR U8098 ( .A(DB[1684]), .B(DB[1669]), .Z(n4508) );
  AND U8099 ( .A(n578), .B(n4509), .Z(n4507) );
  XOR U8100 ( .A(n4510), .B(n4511), .Z(n4509) );
  XOR U8101 ( .A(DB[1669]), .B(DB[1654]), .Z(n4511) );
  AND U8102 ( .A(n582), .B(n4512), .Z(n4510) );
  XOR U8103 ( .A(n4513), .B(n4514), .Z(n4512) );
  XOR U8104 ( .A(DB[1654]), .B(DB[1639]), .Z(n4514) );
  AND U8105 ( .A(n586), .B(n4515), .Z(n4513) );
  XOR U8106 ( .A(n4516), .B(n4517), .Z(n4515) );
  XOR U8107 ( .A(DB[1639]), .B(DB[1624]), .Z(n4517) );
  AND U8108 ( .A(n590), .B(n4518), .Z(n4516) );
  XOR U8109 ( .A(n4519), .B(n4520), .Z(n4518) );
  XOR U8110 ( .A(DB[1624]), .B(DB[1609]), .Z(n4520) );
  AND U8111 ( .A(n594), .B(n4521), .Z(n4519) );
  XOR U8112 ( .A(n4522), .B(n4523), .Z(n4521) );
  XOR U8113 ( .A(DB[1609]), .B(DB[1594]), .Z(n4523) );
  AND U8114 ( .A(n598), .B(n4524), .Z(n4522) );
  XOR U8115 ( .A(n4525), .B(n4526), .Z(n4524) );
  XOR U8116 ( .A(DB[1594]), .B(DB[1579]), .Z(n4526) );
  AND U8117 ( .A(n602), .B(n4527), .Z(n4525) );
  XOR U8118 ( .A(n4528), .B(n4529), .Z(n4527) );
  XOR U8119 ( .A(DB[1579]), .B(DB[1564]), .Z(n4529) );
  AND U8120 ( .A(n606), .B(n4530), .Z(n4528) );
  XOR U8121 ( .A(n4531), .B(n4532), .Z(n4530) );
  XOR U8122 ( .A(DB[1564]), .B(DB[1549]), .Z(n4532) );
  AND U8123 ( .A(n610), .B(n4533), .Z(n4531) );
  XOR U8124 ( .A(n4534), .B(n4535), .Z(n4533) );
  XOR U8125 ( .A(DB[1549]), .B(DB[1534]), .Z(n4535) );
  AND U8126 ( .A(n614), .B(n4536), .Z(n4534) );
  XOR U8127 ( .A(n4537), .B(n4538), .Z(n4536) );
  XOR U8128 ( .A(DB[1534]), .B(DB[1519]), .Z(n4538) );
  AND U8129 ( .A(n618), .B(n4539), .Z(n4537) );
  XOR U8130 ( .A(n4540), .B(n4541), .Z(n4539) );
  XOR U8131 ( .A(DB[1519]), .B(DB[1504]), .Z(n4541) );
  AND U8132 ( .A(n622), .B(n4542), .Z(n4540) );
  XOR U8133 ( .A(n4543), .B(n4544), .Z(n4542) );
  XOR U8134 ( .A(DB[1504]), .B(DB[1489]), .Z(n4544) );
  AND U8135 ( .A(n626), .B(n4545), .Z(n4543) );
  XOR U8136 ( .A(n4546), .B(n4547), .Z(n4545) );
  XOR U8137 ( .A(DB[1489]), .B(DB[1474]), .Z(n4547) );
  AND U8138 ( .A(n630), .B(n4548), .Z(n4546) );
  XOR U8139 ( .A(n4549), .B(n4550), .Z(n4548) );
  XOR U8140 ( .A(DB[1474]), .B(DB[1459]), .Z(n4550) );
  AND U8141 ( .A(n634), .B(n4551), .Z(n4549) );
  XOR U8142 ( .A(n4552), .B(n4553), .Z(n4551) );
  XOR U8143 ( .A(DB[1459]), .B(DB[1444]), .Z(n4553) );
  AND U8144 ( .A(n638), .B(n4554), .Z(n4552) );
  XOR U8145 ( .A(n4555), .B(n4556), .Z(n4554) );
  XOR U8146 ( .A(DB[1444]), .B(DB[1429]), .Z(n4556) );
  AND U8147 ( .A(n642), .B(n4557), .Z(n4555) );
  XOR U8148 ( .A(n4558), .B(n4559), .Z(n4557) );
  XOR U8149 ( .A(DB[1429]), .B(DB[1414]), .Z(n4559) );
  AND U8150 ( .A(n646), .B(n4560), .Z(n4558) );
  XOR U8151 ( .A(n4561), .B(n4562), .Z(n4560) );
  XOR U8152 ( .A(DB[1414]), .B(DB[1399]), .Z(n4562) );
  AND U8153 ( .A(n650), .B(n4563), .Z(n4561) );
  XOR U8154 ( .A(n4564), .B(n4565), .Z(n4563) );
  XOR U8155 ( .A(DB[1399]), .B(DB[1384]), .Z(n4565) );
  AND U8156 ( .A(n654), .B(n4566), .Z(n4564) );
  XOR U8157 ( .A(n4567), .B(n4568), .Z(n4566) );
  XOR U8158 ( .A(DB[1384]), .B(DB[1369]), .Z(n4568) );
  AND U8159 ( .A(n658), .B(n4569), .Z(n4567) );
  XOR U8160 ( .A(n4570), .B(n4571), .Z(n4569) );
  XOR U8161 ( .A(DB[1369]), .B(DB[1354]), .Z(n4571) );
  AND U8162 ( .A(n662), .B(n4572), .Z(n4570) );
  XOR U8163 ( .A(n4573), .B(n4574), .Z(n4572) );
  XOR U8164 ( .A(DB[1354]), .B(DB[1339]), .Z(n4574) );
  AND U8165 ( .A(n666), .B(n4575), .Z(n4573) );
  XOR U8166 ( .A(n4576), .B(n4577), .Z(n4575) );
  XOR U8167 ( .A(DB[1339]), .B(DB[1324]), .Z(n4577) );
  AND U8168 ( .A(n670), .B(n4578), .Z(n4576) );
  XOR U8169 ( .A(n4579), .B(n4580), .Z(n4578) );
  XOR U8170 ( .A(DB[1324]), .B(DB[1309]), .Z(n4580) );
  AND U8171 ( .A(n674), .B(n4581), .Z(n4579) );
  XOR U8172 ( .A(n4582), .B(n4583), .Z(n4581) );
  XOR U8173 ( .A(DB[1309]), .B(DB[1294]), .Z(n4583) );
  AND U8174 ( .A(n678), .B(n4584), .Z(n4582) );
  XOR U8175 ( .A(n4585), .B(n4586), .Z(n4584) );
  XOR U8176 ( .A(DB[1294]), .B(DB[1279]), .Z(n4586) );
  AND U8177 ( .A(n682), .B(n4587), .Z(n4585) );
  XOR U8178 ( .A(n4588), .B(n4589), .Z(n4587) );
  XOR U8179 ( .A(DB[1279]), .B(DB[1264]), .Z(n4589) );
  AND U8180 ( .A(n686), .B(n4590), .Z(n4588) );
  XOR U8181 ( .A(n4591), .B(n4592), .Z(n4590) );
  XOR U8182 ( .A(DB[1264]), .B(DB[1249]), .Z(n4592) );
  AND U8183 ( .A(n690), .B(n4593), .Z(n4591) );
  XOR U8184 ( .A(n4594), .B(n4595), .Z(n4593) );
  XOR U8185 ( .A(DB[1249]), .B(DB[1234]), .Z(n4595) );
  AND U8186 ( .A(n694), .B(n4596), .Z(n4594) );
  XOR U8187 ( .A(n4597), .B(n4598), .Z(n4596) );
  XOR U8188 ( .A(DB[1234]), .B(DB[1219]), .Z(n4598) );
  AND U8189 ( .A(n698), .B(n4599), .Z(n4597) );
  XOR U8190 ( .A(n4600), .B(n4601), .Z(n4599) );
  XOR U8191 ( .A(DB[1219]), .B(DB[1204]), .Z(n4601) );
  AND U8192 ( .A(n702), .B(n4602), .Z(n4600) );
  XOR U8193 ( .A(n4603), .B(n4604), .Z(n4602) );
  XOR U8194 ( .A(DB[1204]), .B(DB[1189]), .Z(n4604) );
  AND U8195 ( .A(n706), .B(n4605), .Z(n4603) );
  XOR U8196 ( .A(n4606), .B(n4607), .Z(n4605) );
  XOR U8197 ( .A(DB[1189]), .B(DB[1174]), .Z(n4607) );
  AND U8198 ( .A(n710), .B(n4608), .Z(n4606) );
  XOR U8199 ( .A(n4609), .B(n4610), .Z(n4608) );
  XOR U8200 ( .A(DB[1174]), .B(DB[1159]), .Z(n4610) );
  AND U8201 ( .A(n714), .B(n4611), .Z(n4609) );
  XOR U8202 ( .A(n4612), .B(n4613), .Z(n4611) );
  XOR U8203 ( .A(DB[1159]), .B(DB[1144]), .Z(n4613) );
  AND U8204 ( .A(n718), .B(n4614), .Z(n4612) );
  XOR U8205 ( .A(n4615), .B(n4616), .Z(n4614) );
  XOR U8206 ( .A(DB[1144]), .B(DB[1129]), .Z(n4616) );
  AND U8207 ( .A(n722), .B(n4617), .Z(n4615) );
  XOR U8208 ( .A(n4618), .B(n4619), .Z(n4617) );
  XOR U8209 ( .A(DB[1129]), .B(DB[1114]), .Z(n4619) );
  AND U8210 ( .A(n726), .B(n4620), .Z(n4618) );
  XOR U8211 ( .A(n4621), .B(n4622), .Z(n4620) );
  XOR U8212 ( .A(DB[1114]), .B(DB[1099]), .Z(n4622) );
  AND U8213 ( .A(n730), .B(n4623), .Z(n4621) );
  XOR U8214 ( .A(n4624), .B(n4625), .Z(n4623) );
  XOR U8215 ( .A(DB[1099]), .B(DB[1084]), .Z(n4625) );
  AND U8216 ( .A(n734), .B(n4626), .Z(n4624) );
  XOR U8217 ( .A(n4627), .B(n4628), .Z(n4626) );
  XOR U8218 ( .A(DB[1084]), .B(DB[1069]), .Z(n4628) );
  AND U8219 ( .A(n738), .B(n4629), .Z(n4627) );
  XOR U8220 ( .A(n4630), .B(n4631), .Z(n4629) );
  XOR U8221 ( .A(DB[1069]), .B(DB[1054]), .Z(n4631) );
  AND U8222 ( .A(n742), .B(n4632), .Z(n4630) );
  XOR U8223 ( .A(n4633), .B(n4634), .Z(n4632) );
  XOR U8224 ( .A(DB[1054]), .B(DB[1039]), .Z(n4634) );
  AND U8225 ( .A(n746), .B(n4635), .Z(n4633) );
  XOR U8226 ( .A(n4636), .B(n4637), .Z(n4635) );
  XOR U8227 ( .A(DB[1039]), .B(DB[1024]), .Z(n4637) );
  AND U8228 ( .A(n750), .B(n4638), .Z(n4636) );
  XOR U8229 ( .A(n4639), .B(n4640), .Z(n4638) );
  XOR U8230 ( .A(DB[1024]), .B(DB[1009]), .Z(n4640) );
  AND U8231 ( .A(n754), .B(n4641), .Z(n4639) );
  XOR U8232 ( .A(n4642), .B(n4643), .Z(n4641) );
  XOR U8233 ( .A(DB[994]), .B(DB[1009]), .Z(n4643) );
  AND U8234 ( .A(n758), .B(n4644), .Z(n4642) );
  XOR U8235 ( .A(n4645), .B(n4646), .Z(n4644) );
  XOR U8236 ( .A(DB[994]), .B(DB[979]), .Z(n4646) );
  AND U8237 ( .A(n762), .B(n4647), .Z(n4645) );
  XOR U8238 ( .A(n4648), .B(n4649), .Z(n4647) );
  XOR U8239 ( .A(DB[979]), .B(DB[964]), .Z(n4649) );
  AND U8240 ( .A(n766), .B(n4650), .Z(n4648) );
  XOR U8241 ( .A(n4651), .B(n4652), .Z(n4650) );
  XOR U8242 ( .A(DB[964]), .B(DB[949]), .Z(n4652) );
  AND U8243 ( .A(n770), .B(n4653), .Z(n4651) );
  XOR U8244 ( .A(n4654), .B(n4655), .Z(n4653) );
  XOR U8245 ( .A(DB[949]), .B(DB[934]), .Z(n4655) );
  AND U8246 ( .A(n774), .B(n4656), .Z(n4654) );
  XOR U8247 ( .A(n4657), .B(n4658), .Z(n4656) );
  XOR U8248 ( .A(DB[934]), .B(DB[919]), .Z(n4658) );
  AND U8249 ( .A(n778), .B(n4659), .Z(n4657) );
  XOR U8250 ( .A(n4660), .B(n4661), .Z(n4659) );
  XOR U8251 ( .A(DB[919]), .B(DB[904]), .Z(n4661) );
  AND U8252 ( .A(n782), .B(n4662), .Z(n4660) );
  XOR U8253 ( .A(n4663), .B(n4664), .Z(n4662) );
  XOR U8254 ( .A(DB[904]), .B(DB[889]), .Z(n4664) );
  AND U8255 ( .A(n786), .B(n4665), .Z(n4663) );
  XOR U8256 ( .A(n4666), .B(n4667), .Z(n4665) );
  XOR U8257 ( .A(DB[889]), .B(DB[874]), .Z(n4667) );
  AND U8258 ( .A(n790), .B(n4668), .Z(n4666) );
  XOR U8259 ( .A(n4669), .B(n4670), .Z(n4668) );
  XOR U8260 ( .A(DB[874]), .B(DB[859]), .Z(n4670) );
  AND U8261 ( .A(n794), .B(n4671), .Z(n4669) );
  XOR U8262 ( .A(n4672), .B(n4673), .Z(n4671) );
  XOR U8263 ( .A(DB[859]), .B(DB[844]), .Z(n4673) );
  AND U8264 ( .A(n798), .B(n4674), .Z(n4672) );
  XOR U8265 ( .A(n4675), .B(n4676), .Z(n4674) );
  XOR U8266 ( .A(DB[844]), .B(DB[829]), .Z(n4676) );
  AND U8267 ( .A(n802), .B(n4677), .Z(n4675) );
  XOR U8268 ( .A(n4678), .B(n4679), .Z(n4677) );
  XOR U8269 ( .A(DB[829]), .B(DB[814]), .Z(n4679) );
  AND U8270 ( .A(n806), .B(n4680), .Z(n4678) );
  XOR U8271 ( .A(n4681), .B(n4682), .Z(n4680) );
  XOR U8272 ( .A(DB[814]), .B(DB[799]), .Z(n4682) );
  AND U8273 ( .A(n810), .B(n4683), .Z(n4681) );
  XOR U8274 ( .A(n4684), .B(n4685), .Z(n4683) );
  XOR U8275 ( .A(DB[799]), .B(DB[784]), .Z(n4685) );
  AND U8276 ( .A(n814), .B(n4686), .Z(n4684) );
  XOR U8277 ( .A(n4687), .B(n4688), .Z(n4686) );
  XOR U8278 ( .A(DB[784]), .B(DB[769]), .Z(n4688) );
  AND U8279 ( .A(n818), .B(n4689), .Z(n4687) );
  XOR U8280 ( .A(n4690), .B(n4691), .Z(n4689) );
  XOR U8281 ( .A(DB[769]), .B(DB[754]), .Z(n4691) );
  AND U8282 ( .A(n822), .B(n4692), .Z(n4690) );
  XOR U8283 ( .A(n4693), .B(n4694), .Z(n4692) );
  XOR U8284 ( .A(DB[754]), .B(DB[739]), .Z(n4694) );
  AND U8285 ( .A(n826), .B(n4695), .Z(n4693) );
  XOR U8286 ( .A(n4696), .B(n4697), .Z(n4695) );
  XOR U8287 ( .A(DB[739]), .B(DB[724]), .Z(n4697) );
  AND U8288 ( .A(n830), .B(n4698), .Z(n4696) );
  XOR U8289 ( .A(n4699), .B(n4700), .Z(n4698) );
  XOR U8290 ( .A(DB[724]), .B(DB[709]), .Z(n4700) );
  AND U8291 ( .A(n834), .B(n4701), .Z(n4699) );
  XOR U8292 ( .A(n4702), .B(n4703), .Z(n4701) );
  XOR U8293 ( .A(DB[709]), .B(DB[694]), .Z(n4703) );
  AND U8294 ( .A(n838), .B(n4704), .Z(n4702) );
  XOR U8295 ( .A(n4705), .B(n4706), .Z(n4704) );
  XOR U8296 ( .A(DB[694]), .B(DB[679]), .Z(n4706) );
  AND U8297 ( .A(n842), .B(n4707), .Z(n4705) );
  XOR U8298 ( .A(n4708), .B(n4709), .Z(n4707) );
  XOR U8299 ( .A(DB[679]), .B(DB[664]), .Z(n4709) );
  AND U8300 ( .A(n846), .B(n4710), .Z(n4708) );
  XOR U8301 ( .A(n4711), .B(n4712), .Z(n4710) );
  XOR U8302 ( .A(DB[664]), .B(DB[649]), .Z(n4712) );
  AND U8303 ( .A(n850), .B(n4713), .Z(n4711) );
  XOR U8304 ( .A(n4714), .B(n4715), .Z(n4713) );
  XOR U8305 ( .A(DB[649]), .B(DB[634]), .Z(n4715) );
  AND U8306 ( .A(n854), .B(n4716), .Z(n4714) );
  XOR U8307 ( .A(n4717), .B(n4718), .Z(n4716) );
  XOR U8308 ( .A(DB[634]), .B(DB[619]), .Z(n4718) );
  AND U8309 ( .A(n858), .B(n4719), .Z(n4717) );
  XOR U8310 ( .A(n4720), .B(n4721), .Z(n4719) );
  XOR U8311 ( .A(DB[619]), .B(DB[604]), .Z(n4721) );
  AND U8312 ( .A(n862), .B(n4722), .Z(n4720) );
  XOR U8313 ( .A(n4723), .B(n4724), .Z(n4722) );
  XOR U8314 ( .A(DB[604]), .B(DB[589]), .Z(n4724) );
  AND U8315 ( .A(n866), .B(n4725), .Z(n4723) );
  XOR U8316 ( .A(n4726), .B(n4727), .Z(n4725) );
  XOR U8317 ( .A(DB[589]), .B(DB[574]), .Z(n4727) );
  AND U8318 ( .A(n870), .B(n4728), .Z(n4726) );
  XOR U8319 ( .A(n4729), .B(n4730), .Z(n4728) );
  XOR U8320 ( .A(DB[574]), .B(DB[559]), .Z(n4730) );
  AND U8321 ( .A(n874), .B(n4731), .Z(n4729) );
  XOR U8322 ( .A(n4732), .B(n4733), .Z(n4731) );
  XOR U8323 ( .A(DB[559]), .B(DB[544]), .Z(n4733) );
  AND U8324 ( .A(n878), .B(n4734), .Z(n4732) );
  XOR U8325 ( .A(n4735), .B(n4736), .Z(n4734) );
  XOR U8326 ( .A(DB[544]), .B(DB[529]), .Z(n4736) );
  AND U8327 ( .A(n882), .B(n4737), .Z(n4735) );
  XOR U8328 ( .A(n4738), .B(n4739), .Z(n4737) );
  XOR U8329 ( .A(DB[529]), .B(DB[514]), .Z(n4739) );
  AND U8330 ( .A(n886), .B(n4740), .Z(n4738) );
  XOR U8331 ( .A(n4741), .B(n4742), .Z(n4740) );
  XOR U8332 ( .A(DB[514]), .B(DB[499]), .Z(n4742) );
  AND U8333 ( .A(n890), .B(n4743), .Z(n4741) );
  XOR U8334 ( .A(n4744), .B(n4745), .Z(n4743) );
  XOR U8335 ( .A(DB[499]), .B(DB[484]), .Z(n4745) );
  AND U8336 ( .A(n894), .B(n4746), .Z(n4744) );
  XOR U8337 ( .A(n4747), .B(n4748), .Z(n4746) );
  XOR U8338 ( .A(DB[484]), .B(DB[469]), .Z(n4748) );
  AND U8339 ( .A(n898), .B(n4749), .Z(n4747) );
  XOR U8340 ( .A(n4750), .B(n4751), .Z(n4749) );
  XOR U8341 ( .A(DB[469]), .B(DB[454]), .Z(n4751) );
  AND U8342 ( .A(n902), .B(n4752), .Z(n4750) );
  XOR U8343 ( .A(n4753), .B(n4754), .Z(n4752) );
  XOR U8344 ( .A(DB[454]), .B(DB[439]), .Z(n4754) );
  AND U8345 ( .A(n906), .B(n4755), .Z(n4753) );
  XOR U8346 ( .A(n4756), .B(n4757), .Z(n4755) );
  XOR U8347 ( .A(DB[439]), .B(DB[424]), .Z(n4757) );
  AND U8348 ( .A(n910), .B(n4758), .Z(n4756) );
  XOR U8349 ( .A(n4759), .B(n4760), .Z(n4758) );
  XOR U8350 ( .A(DB[424]), .B(DB[409]), .Z(n4760) );
  AND U8351 ( .A(n914), .B(n4761), .Z(n4759) );
  XOR U8352 ( .A(n4762), .B(n4763), .Z(n4761) );
  XOR U8353 ( .A(DB[409]), .B(DB[394]), .Z(n4763) );
  AND U8354 ( .A(n918), .B(n4764), .Z(n4762) );
  XOR U8355 ( .A(n4765), .B(n4766), .Z(n4764) );
  XOR U8356 ( .A(DB[394]), .B(DB[379]), .Z(n4766) );
  AND U8357 ( .A(n922), .B(n4767), .Z(n4765) );
  XOR U8358 ( .A(n4768), .B(n4769), .Z(n4767) );
  XOR U8359 ( .A(DB[379]), .B(DB[364]), .Z(n4769) );
  AND U8360 ( .A(n926), .B(n4770), .Z(n4768) );
  XOR U8361 ( .A(n4771), .B(n4772), .Z(n4770) );
  XOR U8362 ( .A(DB[364]), .B(DB[349]), .Z(n4772) );
  AND U8363 ( .A(n930), .B(n4773), .Z(n4771) );
  XOR U8364 ( .A(n4774), .B(n4775), .Z(n4773) );
  XOR U8365 ( .A(DB[349]), .B(DB[334]), .Z(n4775) );
  AND U8366 ( .A(n934), .B(n4776), .Z(n4774) );
  XOR U8367 ( .A(n4777), .B(n4778), .Z(n4776) );
  XOR U8368 ( .A(DB[334]), .B(DB[319]), .Z(n4778) );
  AND U8369 ( .A(n938), .B(n4779), .Z(n4777) );
  XOR U8370 ( .A(n4780), .B(n4781), .Z(n4779) );
  XOR U8371 ( .A(DB[319]), .B(DB[304]), .Z(n4781) );
  AND U8372 ( .A(n942), .B(n4782), .Z(n4780) );
  XOR U8373 ( .A(n4783), .B(n4784), .Z(n4782) );
  XOR U8374 ( .A(DB[304]), .B(DB[289]), .Z(n4784) );
  AND U8375 ( .A(n946), .B(n4785), .Z(n4783) );
  XOR U8376 ( .A(n4786), .B(n4787), .Z(n4785) );
  XOR U8377 ( .A(DB[289]), .B(DB[274]), .Z(n4787) );
  AND U8378 ( .A(n950), .B(n4788), .Z(n4786) );
  XOR U8379 ( .A(n4789), .B(n4790), .Z(n4788) );
  XOR U8380 ( .A(DB[274]), .B(DB[259]), .Z(n4790) );
  AND U8381 ( .A(n954), .B(n4791), .Z(n4789) );
  XOR U8382 ( .A(n4792), .B(n4793), .Z(n4791) );
  XOR U8383 ( .A(DB[259]), .B(DB[244]), .Z(n4793) );
  AND U8384 ( .A(n958), .B(n4794), .Z(n4792) );
  XOR U8385 ( .A(n4795), .B(n4796), .Z(n4794) );
  XOR U8386 ( .A(DB[244]), .B(DB[229]), .Z(n4796) );
  AND U8387 ( .A(n962), .B(n4797), .Z(n4795) );
  XOR U8388 ( .A(n4798), .B(n4799), .Z(n4797) );
  XOR U8389 ( .A(DB[229]), .B(DB[214]), .Z(n4799) );
  AND U8390 ( .A(n966), .B(n4800), .Z(n4798) );
  XOR U8391 ( .A(n4801), .B(n4802), .Z(n4800) );
  XOR U8392 ( .A(DB[214]), .B(DB[199]), .Z(n4802) );
  AND U8393 ( .A(n970), .B(n4803), .Z(n4801) );
  XOR U8394 ( .A(n4804), .B(n4805), .Z(n4803) );
  XOR U8395 ( .A(DB[199]), .B(DB[184]), .Z(n4805) );
  AND U8396 ( .A(n974), .B(n4806), .Z(n4804) );
  XOR U8397 ( .A(n4807), .B(n4808), .Z(n4806) );
  XOR U8398 ( .A(DB[184]), .B(DB[169]), .Z(n4808) );
  AND U8399 ( .A(n978), .B(n4809), .Z(n4807) );
  XOR U8400 ( .A(n4810), .B(n4811), .Z(n4809) );
  XOR U8401 ( .A(DB[169]), .B(DB[154]), .Z(n4811) );
  AND U8402 ( .A(n982), .B(n4812), .Z(n4810) );
  XOR U8403 ( .A(n4813), .B(n4814), .Z(n4812) );
  XOR U8404 ( .A(DB[154]), .B(DB[139]), .Z(n4814) );
  AND U8405 ( .A(n986), .B(n4815), .Z(n4813) );
  XOR U8406 ( .A(n4816), .B(n4817), .Z(n4815) );
  XOR U8407 ( .A(DB[139]), .B(DB[124]), .Z(n4817) );
  AND U8408 ( .A(n990), .B(n4818), .Z(n4816) );
  XOR U8409 ( .A(n4819), .B(n4820), .Z(n4818) );
  XOR U8410 ( .A(DB[124]), .B(DB[109]), .Z(n4820) );
  AND U8411 ( .A(n994), .B(n4821), .Z(n4819) );
  XOR U8412 ( .A(n4822), .B(n4823), .Z(n4821) );
  XOR U8413 ( .A(DB[94]), .B(DB[109]), .Z(n4823) );
  AND U8414 ( .A(n998), .B(n4824), .Z(n4822) );
  XOR U8415 ( .A(n4825), .B(n4826), .Z(n4824) );
  XOR U8416 ( .A(DB[94]), .B(DB[79]), .Z(n4826) );
  AND U8417 ( .A(n1002), .B(n4827), .Z(n4825) );
  XOR U8418 ( .A(n4828), .B(n4829), .Z(n4827) );
  XOR U8419 ( .A(DB[79]), .B(DB[64]), .Z(n4829) );
  AND U8420 ( .A(n1006), .B(n4830), .Z(n4828) );
  XOR U8421 ( .A(n4831), .B(n4832), .Z(n4830) );
  XOR U8422 ( .A(DB[64]), .B(DB[49]), .Z(n4832) );
  AND U8423 ( .A(n1010), .B(n4833), .Z(n4831) );
  XOR U8424 ( .A(n4834), .B(n4835), .Z(n4833) );
  XOR U8425 ( .A(DB[49]), .B(DB[34]), .Z(n4835) );
  AND U8426 ( .A(n1014), .B(n4836), .Z(n4834) );
  XOR U8427 ( .A(n4837), .B(n4838), .Z(n4836) );
  XOR U8428 ( .A(DB[34]), .B(DB[19]), .Z(n4838) );
  AND U8429 ( .A(n1018), .B(n4839), .Z(n4837) );
  XOR U8430 ( .A(DB[4]), .B(DB[19]), .Z(n4839) );
  XOR U8431 ( .A(DB[3828]), .B(n4840), .Z(min_val_out[3]) );
  AND U8432 ( .A(n2), .B(n4841), .Z(n4840) );
  XOR U8433 ( .A(n4842), .B(n4843), .Z(n4841) );
  XOR U8434 ( .A(DB[3828]), .B(DB[3813]), .Z(n4843) );
  AND U8435 ( .A(n6), .B(n4844), .Z(n4842) );
  XOR U8436 ( .A(n4845), .B(n4846), .Z(n4844) );
  XOR U8437 ( .A(DB[3813]), .B(DB[3798]), .Z(n4846) );
  AND U8438 ( .A(n10), .B(n4847), .Z(n4845) );
  XOR U8439 ( .A(n4848), .B(n4849), .Z(n4847) );
  XOR U8440 ( .A(DB[3798]), .B(DB[3783]), .Z(n4849) );
  AND U8441 ( .A(n14), .B(n4850), .Z(n4848) );
  XOR U8442 ( .A(n4851), .B(n4852), .Z(n4850) );
  XOR U8443 ( .A(DB[3783]), .B(DB[3768]), .Z(n4852) );
  AND U8444 ( .A(n18), .B(n4853), .Z(n4851) );
  XOR U8445 ( .A(n4854), .B(n4855), .Z(n4853) );
  XOR U8446 ( .A(DB[3768]), .B(DB[3753]), .Z(n4855) );
  AND U8447 ( .A(n22), .B(n4856), .Z(n4854) );
  XOR U8448 ( .A(n4857), .B(n4858), .Z(n4856) );
  XOR U8449 ( .A(DB[3753]), .B(DB[3738]), .Z(n4858) );
  AND U8450 ( .A(n26), .B(n4859), .Z(n4857) );
  XOR U8451 ( .A(n4860), .B(n4861), .Z(n4859) );
  XOR U8452 ( .A(DB[3738]), .B(DB[3723]), .Z(n4861) );
  AND U8453 ( .A(n30), .B(n4862), .Z(n4860) );
  XOR U8454 ( .A(n4863), .B(n4864), .Z(n4862) );
  XOR U8455 ( .A(DB[3723]), .B(DB[3708]), .Z(n4864) );
  AND U8456 ( .A(n34), .B(n4865), .Z(n4863) );
  XOR U8457 ( .A(n4866), .B(n4867), .Z(n4865) );
  XOR U8458 ( .A(DB[3708]), .B(DB[3693]), .Z(n4867) );
  AND U8459 ( .A(n38), .B(n4868), .Z(n4866) );
  XOR U8460 ( .A(n4869), .B(n4870), .Z(n4868) );
  XOR U8461 ( .A(DB[3693]), .B(DB[3678]), .Z(n4870) );
  AND U8462 ( .A(n42), .B(n4871), .Z(n4869) );
  XOR U8463 ( .A(n4872), .B(n4873), .Z(n4871) );
  XOR U8464 ( .A(DB[3678]), .B(DB[3663]), .Z(n4873) );
  AND U8465 ( .A(n46), .B(n4874), .Z(n4872) );
  XOR U8466 ( .A(n4875), .B(n4876), .Z(n4874) );
  XOR U8467 ( .A(DB[3663]), .B(DB[3648]), .Z(n4876) );
  AND U8468 ( .A(n50), .B(n4877), .Z(n4875) );
  XOR U8469 ( .A(n4878), .B(n4879), .Z(n4877) );
  XOR U8470 ( .A(DB[3648]), .B(DB[3633]), .Z(n4879) );
  AND U8471 ( .A(n54), .B(n4880), .Z(n4878) );
  XOR U8472 ( .A(n4881), .B(n4882), .Z(n4880) );
  XOR U8473 ( .A(DB[3633]), .B(DB[3618]), .Z(n4882) );
  AND U8474 ( .A(n58), .B(n4883), .Z(n4881) );
  XOR U8475 ( .A(n4884), .B(n4885), .Z(n4883) );
  XOR U8476 ( .A(DB[3618]), .B(DB[3603]), .Z(n4885) );
  AND U8477 ( .A(n62), .B(n4886), .Z(n4884) );
  XOR U8478 ( .A(n4887), .B(n4888), .Z(n4886) );
  XOR U8479 ( .A(DB[3603]), .B(DB[3588]), .Z(n4888) );
  AND U8480 ( .A(n66), .B(n4889), .Z(n4887) );
  XOR U8481 ( .A(n4890), .B(n4891), .Z(n4889) );
  XOR U8482 ( .A(DB[3588]), .B(DB[3573]), .Z(n4891) );
  AND U8483 ( .A(n70), .B(n4892), .Z(n4890) );
  XOR U8484 ( .A(n4893), .B(n4894), .Z(n4892) );
  XOR U8485 ( .A(DB[3573]), .B(DB[3558]), .Z(n4894) );
  AND U8486 ( .A(n74), .B(n4895), .Z(n4893) );
  XOR U8487 ( .A(n4896), .B(n4897), .Z(n4895) );
  XOR U8488 ( .A(DB[3558]), .B(DB[3543]), .Z(n4897) );
  AND U8489 ( .A(n78), .B(n4898), .Z(n4896) );
  XOR U8490 ( .A(n4899), .B(n4900), .Z(n4898) );
  XOR U8491 ( .A(DB[3543]), .B(DB[3528]), .Z(n4900) );
  AND U8492 ( .A(n82), .B(n4901), .Z(n4899) );
  XOR U8493 ( .A(n4902), .B(n4903), .Z(n4901) );
  XOR U8494 ( .A(DB[3528]), .B(DB[3513]), .Z(n4903) );
  AND U8495 ( .A(n86), .B(n4904), .Z(n4902) );
  XOR U8496 ( .A(n4905), .B(n4906), .Z(n4904) );
  XOR U8497 ( .A(DB[3513]), .B(DB[3498]), .Z(n4906) );
  AND U8498 ( .A(n90), .B(n4907), .Z(n4905) );
  XOR U8499 ( .A(n4908), .B(n4909), .Z(n4907) );
  XOR U8500 ( .A(DB[3498]), .B(DB[3483]), .Z(n4909) );
  AND U8501 ( .A(n94), .B(n4910), .Z(n4908) );
  XOR U8502 ( .A(n4911), .B(n4912), .Z(n4910) );
  XOR U8503 ( .A(DB[3483]), .B(DB[3468]), .Z(n4912) );
  AND U8504 ( .A(n98), .B(n4913), .Z(n4911) );
  XOR U8505 ( .A(n4914), .B(n4915), .Z(n4913) );
  XOR U8506 ( .A(DB[3468]), .B(DB[3453]), .Z(n4915) );
  AND U8507 ( .A(n102), .B(n4916), .Z(n4914) );
  XOR U8508 ( .A(n4917), .B(n4918), .Z(n4916) );
  XOR U8509 ( .A(DB[3453]), .B(DB[3438]), .Z(n4918) );
  AND U8510 ( .A(n106), .B(n4919), .Z(n4917) );
  XOR U8511 ( .A(n4920), .B(n4921), .Z(n4919) );
  XOR U8512 ( .A(DB[3438]), .B(DB[3423]), .Z(n4921) );
  AND U8513 ( .A(n110), .B(n4922), .Z(n4920) );
  XOR U8514 ( .A(n4923), .B(n4924), .Z(n4922) );
  XOR U8515 ( .A(DB[3423]), .B(DB[3408]), .Z(n4924) );
  AND U8516 ( .A(n114), .B(n4925), .Z(n4923) );
  XOR U8517 ( .A(n4926), .B(n4927), .Z(n4925) );
  XOR U8518 ( .A(DB[3408]), .B(DB[3393]), .Z(n4927) );
  AND U8519 ( .A(n118), .B(n4928), .Z(n4926) );
  XOR U8520 ( .A(n4929), .B(n4930), .Z(n4928) );
  XOR U8521 ( .A(DB[3393]), .B(DB[3378]), .Z(n4930) );
  AND U8522 ( .A(n122), .B(n4931), .Z(n4929) );
  XOR U8523 ( .A(n4932), .B(n4933), .Z(n4931) );
  XOR U8524 ( .A(DB[3378]), .B(DB[3363]), .Z(n4933) );
  AND U8525 ( .A(n126), .B(n4934), .Z(n4932) );
  XOR U8526 ( .A(n4935), .B(n4936), .Z(n4934) );
  XOR U8527 ( .A(DB[3363]), .B(DB[3348]), .Z(n4936) );
  AND U8528 ( .A(n130), .B(n4937), .Z(n4935) );
  XOR U8529 ( .A(n4938), .B(n4939), .Z(n4937) );
  XOR U8530 ( .A(DB[3348]), .B(DB[3333]), .Z(n4939) );
  AND U8531 ( .A(n134), .B(n4940), .Z(n4938) );
  XOR U8532 ( .A(n4941), .B(n4942), .Z(n4940) );
  XOR U8533 ( .A(DB[3333]), .B(DB[3318]), .Z(n4942) );
  AND U8534 ( .A(n138), .B(n4943), .Z(n4941) );
  XOR U8535 ( .A(n4944), .B(n4945), .Z(n4943) );
  XOR U8536 ( .A(DB[3318]), .B(DB[3303]), .Z(n4945) );
  AND U8537 ( .A(n142), .B(n4946), .Z(n4944) );
  XOR U8538 ( .A(n4947), .B(n4948), .Z(n4946) );
  XOR U8539 ( .A(DB[3303]), .B(DB[3288]), .Z(n4948) );
  AND U8540 ( .A(n146), .B(n4949), .Z(n4947) );
  XOR U8541 ( .A(n4950), .B(n4951), .Z(n4949) );
  XOR U8542 ( .A(DB[3288]), .B(DB[3273]), .Z(n4951) );
  AND U8543 ( .A(n150), .B(n4952), .Z(n4950) );
  XOR U8544 ( .A(n4953), .B(n4954), .Z(n4952) );
  XOR U8545 ( .A(DB[3273]), .B(DB[3258]), .Z(n4954) );
  AND U8546 ( .A(n154), .B(n4955), .Z(n4953) );
  XOR U8547 ( .A(n4956), .B(n4957), .Z(n4955) );
  XOR U8548 ( .A(DB[3258]), .B(DB[3243]), .Z(n4957) );
  AND U8549 ( .A(n158), .B(n4958), .Z(n4956) );
  XOR U8550 ( .A(n4959), .B(n4960), .Z(n4958) );
  XOR U8551 ( .A(DB[3243]), .B(DB[3228]), .Z(n4960) );
  AND U8552 ( .A(n162), .B(n4961), .Z(n4959) );
  XOR U8553 ( .A(n4962), .B(n4963), .Z(n4961) );
  XOR U8554 ( .A(DB[3228]), .B(DB[3213]), .Z(n4963) );
  AND U8555 ( .A(n166), .B(n4964), .Z(n4962) );
  XOR U8556 ( .A(n4965), .B(n4966), .Z(n4964) );
  XOR U8557 ( .A(DB[3213]), .B(DB[3198]), .Z(n4966) );
  AND U8558 ( .A(n170), .B(n4967), .Z(n4965) );
  XOR U8559 ( .A(n4968), .B(n4969), .Z(n4967) );
  XOR U8560 ( .A(DB[3198]), .B(DB[3183]), .Z(n4969) );
  AND U8561 ( .A(n174), .B(n4970), .Z(n4968) );
  XOR U8562 ( .A(n4971), .B(n4972), .Z(n4970) );
  XOR U8563 ( .A(DB[3183]), .B(DB[3168]), .Z(n4972) );
  AND U8564 ( .A(n178), .B(n4973), .Z(n4971) );
  XOR U8565 ( .A(n4974), .B(n4975), .Z(n4973) );
  XOR U8566 ( .A(DB[3168]), .B(DB[3153]), .Z(n4975) );
  AND U8567 ( .A(n182), .B(n4976), .Z(n4974) );
  XOR U8568 ( .A(n4977), .B(n4978), .Z(n4976) );
  XOR U8569 ( .A(DB[3153]), .B(DB[3138]), .Z(n4978) );
  AND U8570 ( .A(n186), .B(n4979), .Z(n4977) );
  XOR U8571 ( .A(n4980), .B(n4981), .Z(n4979) );
  XOR U8572 ( .A(DB[3138]), .B(DB[3123]), .Z(n4981) );
  AND U8573 ( .A(n190), .B(n4982), .Z(n4980) );
  XOR U8574 ( .A(n4983), .B(n4984), .Z(n4982) );
  XOR U8575 ( .A(DB[3123]), .B(DB[3108]), .Z(n4984) );
  AND U8576 ( .A(n194), .B(n4985), .Z(n4983) );
  XOR U8577 ( .A(n4986), .B(n4987), .Z(n4985) );
  XOR U8578 ( .A(DB[3108]), .B(DB[3093]), .Z(n4987) );
  AND U8579 ( .A(n198), .B(n4988), .Z(n4986) );
  XOR U8580 ( .A(n4989), .B(n4990), .Z(n4988) );
  XOR U8581 ( .A(DB[3093]), .B(DB[3078]), .Z(n4990) );
  AND U8582 ( .A(n202), .B(n4991), .Z(n4989) );
  XOR U8583 ( .A(n4992), .B(n4993), .Z(n4991) );
  XOR U8584 ( .A(DB[3078]), .B(DB[3063]), .Z(n4993) );
  AND U8585 ( .A(n206), .B(n4994), .Z(n4992) );
  XOR U8586 ( .A(n4995), .B(n4996), .Z(n4994) );
  XOR U8587 ( .A(DB[3063]), .B(DB[3048]), .Z(n4996) );
  AND U8588 ( .A(n210), .B(n4997), .Z(n4995) );
  XOR U8589 ( .A(n4998), .B(n4999), .Z(n4997) );
  XOR U8590 ( .A(DB[3048]), .B(DB[3033]), .Z(n4999) );
  AND U8591 ( .A(n214), .B(n5000), .Z(n4998) );
  XOR U8592 ( .A(n5001), .B(n5002), .Z(n5000) );
  XOR U8593 ( .A(DB[3033]), .B(DB[3018]), .Z(n5002) );
  AND U8594 ( .A(n218), .B(n5003), .Z(n5001) );
  XOR U8595 ( .A(n5004), .B(n5005), .Z(n5003) );
  XOR U8596 ( .A(DB[3018]), .B(DB[3003]), .Z(n5005) );
  AND U8597 ( .A(n222), .B(n5006), .Z(n5004) );
  XOR U8598 ( .A(n5007), .B(n5008), .Z(n5006) );
  XOR U8599 ( .A(DB[3003]), .B(DB[2988]), .Z(n5008) );
  AND U8600 ( .A(n226), .B(n5009), .Z(n5007) );
  XOR U8601 ( .A(n5010), .B(n5011), .Z(n5009) );
  XOR U8602 ( .A(DB[2988]), .B(DB[2973]), .Z(n5011) );
  AND U8603 ( .A(n230), .B(n5012), .Z(n5010) );
  XOR U8604 ( .A(n5013), .B(n5014), .Z(n5012) );
  XOR U8605 ( .A(DB[2973]), .B(DB[2958]), .Z(n5014) );
  AND U8606 ( .A(n234), .B(n5015), .Z(n5013) );
  XOR U8607 ( .A(n5016), .B(n5017), .Z(n5015) );
  XOR U8608 ( .A(DB[2958]), .B(DB[2943]), .Z(n5017) );
  AND U8609 ( .A(n238), .B(n5018), .Z(n5016) );
  XOR U8610 ( .A(n5019), .B(n5020), .Z(n5018) );
  XOR U8611 ( .A(DB[2943]), .B(DB[2928]), .Z(n5020) );
  AND U8612 ( .A(n242), .B(n5021), .Z(n5019) );
  XOR U8613 ( .A(n5022), .B(n5023), .Z(n5021) );
  XOR U8614 ( .A(DB[2928]), .B(DB[2913]), .Z(n5023) );
  AND U8615 ( .A(n246), .B(n5024), .Z(n5022) );
  XOR U8616 ( .A(n5025), .B(n5026), .Z(n5024) );
  XOR U8617 ( .A(DB[2913]), .B(DB[2898]), .Z(n5026) );
  AND U8618 ( .A(n250), .B(n5027), .Z(n5025) );
  XOR U8619 ( .A(n5028), .B(n5029), .Z(n5027) );
  XOR U8620 ( .A(DB[2898]), .B(DB[2883]), .Z(n5029) );
  AND U8621 ( .A(n254), .B(n5030), .Z(n5028) );
  XOR U8622 ( .A(n5031), .B(n5032), .Z(n5030) );
  XOR U8623 ( .A(DB[2883]), .B(DB[2868]), .Z(n5032) );
  AND U8624 ( .A(n258), .B(n5033), .Z(n5031) );
  XOR U8625 ( .A(n5034), .B(n5035), .Z(n5033) );
  XOR U8626 ( .A(DB[2868]), .B(DB[2853]), .Z(n5035) );
  AND U8627 ( .A(n262), .B(n5036), .Z(n5034) );
  XOR U8628 ( .A(n5037), .B(n5038), .Z(n5036) );
  XOR U8629 ( .A(DB[2853]), .B(DB[2838]), .Z(n5038) );
  AND U8630 ( .A(n266), .B(n5039), .Z(n5037) );
  XOR U8631 ( .A(n5040), .B(n5041), .Z(n5039) );
  XOR U8632 ( .A(DB[2838]), .B(DB[2823]), .Z(n5041) );
  AND U8633 ( .A(n270), .B(n5042), .Z(n5040) );
  XOR U8634 ( .A(n5043), .B(n5044), .Z(n5042) );
  XOR U8635 ( .A(DB[2823]), .B(DB[2808]), .Z(n5044) );
  AND U8636 ( .A(n274), .B(n5045), .Z(n5043) );
  XOR U8637 ( .A(n5046), .B(n5047), .Z(n5045) );
  XOR U8638 ( .A(DB[2808]), .B(DB[2793]), .Z(n5047) );
  AND U8639 ( .A(n278), .B(n5048), .Z(n5046) );
  XOR U8640 ( .A(n5049), .B(n5050), .Z(n5048) );
  XOR U8641 ( .A(DB[2793]), .B(DB[2778]), .Z(n5050) );
  AND U8642 ( .A(n282), .B(n5051), .Z(n5049) );
  XOR U8643 ( .A(n5052), .B(n5053), .Z(n5051) );
  XOR U8644 ( .A(DB[2778]), .B(DB[2763]), .Z(n5053) );
  AND U8645 ( .A(n286), .B(n5054), .Z(n5052) );
  XOR U8646 ( .A(n5055), .B(n5056), .Z(n5054) );
  XOR U8647 ( .A(DB[2763]), .B(DB[2748]), .Z(n5056) );
  AND U8648 ( .A(n290), .B(n5057), .Z(n5055) );
  XOR U8649 ( .A(n5058), .B(n5059), .Z(n5057) );
  XOR U8650 ( .A(DB[2748]), .B(DB[2733]), .Z(n5059) );
  AND U8651 ( .A(n294), .B(n5060), .Z(n5058) );
  XOR U8652 ( .A(n5061), .B(n5062), .Z(n5060) );
  XOR U8653 ( .A(DB[2733]), .B(DB[2718]), .Z(n5062) );
  AND U8654 ( .A(n298), .B(n5063), .Z(n5061) );
  XOR U8655 ( .A(n5064), .B(n5065), .Z(n5063) );
  XOR U8656 ( .A(DB[2718]), .B(DB[2703]), .Z(n5065) );
  AND U8657 ( .A(n302), .B(n5066), .Z(n5064) );
  XOR U8658 ( .A(n5067), .B(n5068), .Z(n5066) );
  XOR U8659 ( .A(DB[2703]), .B(DB[2688]), .Z(n5068) );
  AND U8660 ( .A(n306), .B(n5069), .Z(n5067) );
  XOR U8661 ( .A(n5070), .B(n5071), .Z(n5069) );
  XOR U8662 ( .A(DB[2688]), .B(DB[2673]), .Z(n5071) );
  AND U8663 ( .A(n310), .B(n5072), .Z(n5070) );
  XOR U8664 ( .A(n5073), .B(n5074), .Z(n5072) );
  XOR U8665 ( .A(DB[2673]), .B(DB[2658]), .Z(n5074) );
  AND U8666 ( .A(n314), .B(n5075), .Z(n5073) );
  XOR U8667 ( .A(n5076), .B(n5077), .Z(n5075) );
  XOR U8668 ( .A(DB[2658]), .B(DB[2643]), .Z(n5077) );
  AND U8669 ( .A(n318), .B(n5078), .Z(n5076) );
  XOR U8670 ( .A(n5079), .B(n5080), .Z(n5078) );
  XOR U8671 ( .A(DB[2643]), .B(DB[2628]), .Z(n5080) );
  AND U8672 ( .A(n322), .B(n5081), .Z(n5079) );
  XOR U8673 ( .A(n5082), .B(n5083), .Z(n5081) );
  XOR U8674 ( .A(DB[2628]), .B(DB[2613]), .Z(n5083) );
  AND U8675 ( .A(n326), .B(n5084), .Z(n5082) );
  XOR U8676 ( .A(n5085), .B(n5086), .Z(n5084) );
  XOR U8677 ( .A(DB[2613]), .B(DB[2598]), .Z(n5086) );
  AND U8678 ( .A(n330), .B(n5087), .Z(n5085) );
  XOR U8679 ( .A(n5088), .B(n5089), .Z(n5087) );
  XOR U8680 ( .A(DB[2598]), .B(DB[2583]), .Z(n5089) );
  AND U8681 ( .A(n334), .B(n5090), .Z(n5088) );
  XOR U8682 ( .A(n5091), .B(n5092), .Z(n5090) );
  XOR U8683 ( .A(DB[2583]), .B(DB[2568]), .Z(n5092) );
  AND U8684 ( .A(n338), .B(n5093), .Z(n5091) );
  XOR U8685 ( .A(n5094), .B(n5095), .Z(n5093) );
  XOR U8686 ( .A(DB[2568]), .B(DB[2553]), .Z(n5095) );
  AND U8687 ( .A(n342), .B(n5096), .Z(n5094) );
  XOR U8688 ( .A(n5097), .B(n5098), .Z(n5096) );
  XOR U8689 ( .A(DB[2553]), .B(DB[2538]), .Z(n5098) );
  AND U8690 ( .A(n346), .B(n5099), .Z(n5097) );
  XOR U8691 ( .A(n5100), .B(n5101), .Z(n5099) );
  XOR U8692 ( .A(DB[2538]), .B(DB[2523]), .Z(n5101) );
  AND U8693 ( .A(n350), .B(n5102), .Z(n5100) );
  XOR U8694 ( .A(n5103), .B(n5104), .Z(n5102) );
  XOR U8695 ( .A(DB[2523]), .B(DB[2508]), .Z(n5104) );
  AND U8696 ( .A(n354), .B(n5105), .Z(n5103) );
  XOR U8697 ( .A(n5106), .B(n5107), .Z(n5105) );
  XOR U8698 ( .A(DB[2508]), .B(DB[2493]), .Z(n5107) );
  AND U8699 ( .A(n358), .B(n5108), .Z(n5106) );
  XOR U8700 ( .A(n5109), .B(n5110), .Z(n5108) );
  XOR U8701 ( .A(DB[2493]), .B(DB[2478]), .Z(n5110) );
  AND U8702 ( .A(n362), .B(n5111), .Z(n5109) );
  XOR U8703 ( .A(n5112), .B(n5113), .Z(n5111) );
  XOR U8704 ( .A(DB[2478]), .B(DB[2463]), .Z(n5113) );
  AND U8705 ( .A(n366), .B(n5114), .Z(n5112) );
  XOR U8706 ( .A(n5115), .B(n5116), .Z(n5114) );
  XOR U8707 ( .A(DB[2463]), .B(DB[2448]), .Z(n5116) );
  AND U8708 ( .A(n370), .B(n5117), .Z(n5115) );
  XOR U8709 ( .A(n5118), .B(n5119), .Z(n5117) );
  XOR U8710 ( .A(DB[2448]), .B(DB[2433]), .Z(n5119) );
  AND U8711 ( .A(n374), .B(n5120), .Z(n5118) );
  XOR U8712 ( .A(n5121), .B(n5122), .Z(n5120) );
  XOR U8713 ( .A(DB[2433]), .B(DB[2418]), .Z(n5122) );
  AND U8714 ( .A(n378), .B(n5123), .Z(n5121) );
  XOR U8715 ( .A(n5124), .B(n5125), .Z(n5123) );
  XOR U8716 ( .A(DB[2418]), .B(DB[2403]), .Z(n5125) );
  AND U8717 ( .A(n382), .B(n5126), .Z(n5124) );
  XOR U8718 ( .A(n5127), .B(n5128), .Z(n5126) );
  XOR U8719 ( .A(DB[2403]), .B(DB[2388]), .Z(n5128) );
  AND U8720 ( .A(n386), .B(n5129), .Z(n5127) );
  XOR U8721 ( .A(n5130), .B(n5131), .Z(n5129) );
  XOR U8722 ( .A(DB[2388]), .B(DB[2373]), .Z(n5131) );
  AND U8723 ( .A(n390), .B(n5132), .Z(n5130) );
  XOR U8724 ( .A(n5133), .B(n5134), .Z(n5132) );
  XOR U8725 ( .A(DB[2373]), .B(DB[2358]), .Z(n5134) );
  AND U8726 ( .A(n394), .B(n5135), .Z(n5133) );
  XOR U8727 ( .A(n5136), .B(n5137), .Z(n5135) );
  XOR U8728 ( .A(DB[2358]), .B(DB[2343]), .Z(n5137) );
  AND U8729 ( .A(n398), .B(n5138), .Z(n5136) );
  XOR U8730 ( .A(n5139), .B(n5140), .Z(n5138) );
  XOR U8731 ( .A(DB[2343]), .B(DB[2328]), .Z(n5140) );
  AND U8732 ( .A(n402), .B(n5141), .Z(n5139) );
  XOR U8733 ( .A(n5142), .B(n5143), .Z(n5141) );
  XOR U8734 ( .A(DB[2328]), .B(DB[2313]), .Z(n5143) );
  AND U8735 ( .A(n406), .B(n5144), .Z(n5142) );
  XOR U8736 ( .A(n5145), .B(n5146), .Z(n5144) );
  XOR U8737 ( .A(DB[2313]), .B(DB[2298]), .Z(n5146) );
  AND U8738 ( .A(n410), .B(n5147), .Z(n5145) );
  XOR U8739 ( .A(n5148), .B(n5149), .Z(n5147) );
  XOR U8740 ( .A(DB[2298]), .B(DB[2283]), .Z(n5149) );
  AND U8741 ( .A(n414), .B(n5150), .Z(n5148) );
  XOR U8742 ( .A(n5151), .B(n5152), .Z(n5150) );
  XOR U8743 ( .A(DB[2283]), .B(DB[2268]), .Z(n5152) );
  AND U8744 ( .A(n418), .B(n5153), .Z(n5151) );
  XOR U8745 ( .A(n5154), .B(n5155), .Z(n5153) );
  XOR U8746 ( .A(DB[2268]), .B(DB[2253]), .Z(n5155) );
  AND U8747 ( .A(n422), .B(n5156), .Z(n5154) );
  XOR U8748 ( .A(n5157), .B(n5158), .Z(n5156) );
  XOR U8749 ( .A(DB[2253]), .B(DB[2238]), .Z(n5158) );
  AND U8750 ( .A(n426), .B(n5159), .Z(n5157) );
  XOR U8751 ( .A(n5160), .B(n5161), .Z(n5159) );
  XOR U8752 ( .A(DB[2238]), .B(DB[2223]), .Z(n5161) );
  AND U8753 ( .A(n430), .B(n5162), .Z(n5160) );
  XOR U8754 ( .A(n5163), .B(n5164), .Z(n5162) );
  XOR U8755 ( .A(DB[2223]), .B(DB[2208]), .Z(n5164) );
  AND U8756 ( .A(n434), .B(n5165), .Z(n5163) );
  XOR U8757 ( .A(n5166), .B(n5167), .Z(n5165) );
  XOR U8758 ( .A(DB[2208]), .B(DB[2193]), .Z(n5167) );
  AND U8759 ( .A(n438), .B(n5168), .Z(n5166) );
  XOR U8760 ( .A(n5169), .B(n5170), .Z(n5168) );
  XOR U8761 ( .A(DB[2193]), .B(DB[2178]), .Z(n5170) );
  AND U8762 ( .A(n442), .B(n5171), .Z(n5169) );
  XOR U8763 ( .A(n5172), .B(n5173), .Z(n5171) );
  XOR U8764 ( .A(DB[2178]), .B(DB[2163]), .Z(n5173) );
  AND U8765 ( .A(n446), .B(n5174), .Z(n5172) );
  XOR U8766 ( .A(n5175), .B(n5176), .Z(n5174) );
  XOR U8767 ( .A(DB[2163]), .B(DB[2148]), .Z(n5176) );
  AND U8768 ( .A(n450), .B(n5177), .Z(n5175) );
  XOR U8769 ( .A(n5178), .B(n5179), .Z(n5177) );
  XOR U8770 ( .A(DB[2148]), .B(DB[2133]), .Z(n5179) );
  AND U8771 ( .A(n454), .B(n5180), .Z(n5178) );
  XOR U8772 ( .A(n5181), .B(n5182), .Z(n5180) );
  XOR U8773 ( .A(DB[2133]), .B(DB[2118]), .Z(n5182) );
  AND U8774 ( .A(n458), .B(n5183), .Z(n5181) );
  XOR U8775 ( .A(n5184), .B(n5185), .Z(n5183) );
  XOR U8776 ( .A(DB[2118]), .B(DB[2103]), .Z(n5185) );
  AND U8777 ( .A(n462), .B(n5186), .Z(n5184) );
  XOR U8778 ( .A(n5187), .B(n5188), .Z(n5186) );
  XOR U8779 ( .A(DB[2103]), .B(DB[2088]), .Z(n5188) );
  AND U8780 ( .A(n466), .B(n5189), .Z(n5187) );
  XOR U8781 ( .A(n5190), .B(n5191), .Z(n5189) );
  XOR U8782 ( .A(DB[2088]), .B(DB[2073]), .Z(n5191) );
  AND U8783 ( .A(n470), .B(n5192), .Z(n5190) );
  XOR U8784 ( .A(n5193), .B(n5194), .Z(n5192) );
  XOR U8785 ( .A(DB[2073]), .B(DB[2058]), .Z(n5194) );
  AND U8786 ( .A(n474), .B(n5195), .Z(n5193) );
  XOR U8787 ( .A(n5196), .B(n5197), .Z(n5195) );
  XOR U8788 ( .A(DB[2058]), .B(DB[2043]), .Z(n5197) );
  AND U8789 ( .A(n478), .B(n5198), .Z(n5196) );
  XOR U8790 ( .A(n5199), .B(n5200), .Z(n5198) );
  XOR U8791 ( .A(DB[2043]), .B(DB[2028]), .Z(n5200) );
  AND U8792 ( .A(n482), .B(n5201), .Z(n5199) );
  XOR U8793 ( .A(n5202), .B(n5203), .Z(n5201) );
  XOR U8794 ( .A(DB[2028]), .B(DB[2013]), .Z(n5203) );
  AND U8795 ( .A(n486), .B(n5204), .Z(n5202) );
  XOR U8796 ( .A(n5205), .B(n5206), .Z(n5204) );
  XOR U8797 ( .A(DB[2013]), .B(DB[1998]), .Z(n5206) );
  AND U8798 ( .A(n490), .B(n5207), .Z(n5205) );
  XOR U8799 ( .A(n5208), .B(n5209), .Z(n5207) );
  XOR U8800 ( .A(DB[1998]), .B(DB[1983]), .Z(n5209) );
  AND U8801 ( .A(n494), .B(n5210), .Z(n5208) );
  XOR U8802 ( .A(n5211), .B(n5212), .Z(n5210) );
  XOR U8803 ( .A(DB[1983]), .B(DB[1968]), .Z(n5212) );
  AND U8804 ( .A(n498), .B(n5213), .Z(n5211) );
  XOR U8805 ( .A(n5214), .B(n5215), .Z(n5213) );
  XOR U8806 ( .A(DB[1968]), .B(DB[1953]), .Z(n5215) );
  AND U8807 ( .A(n502), .B(n5216), .Z(n5214) );
  XOR U8808 ( .A(n5217), .B(n5218), .Z(n5216) );
  XOR U8809 ( .A(DB[1953]), .B(DB[1938]), .Z(n5218) );
  AND U8810 ( .A(n506), .B(n5219), .Z(n5217) );
  XOR U8811 ( .A(n5220), .B(n5221), .Z(n5219) );
  XOR U8812 ( .A(DB[1938]), .B(DB[1923]), .Z(n5221) );
  AND U8813 ( .A(n510), .B(n5222), .Z(n5220) );
  XOR U8814 ( .A(n5223), .B(n5224), .Z(n5222) );
  XOR U8815 ( .A(DB[1923]), .B(DB[1908]), .Z(n5224) );
  AND U8816 ( .A(n514), .B(n5225), .Z(n5223) );
  XOR U8817 ( .A(n5226), .B(n5227), .Z(n5225) );
  XOR U8818 ( .A(DB[1908]), .B(DB[1893]), .Z(n5227) );
  AND U8819 ( .A(n518), .B(n5228), .Z(n5226) );
  XOR U8820 ( .A(n5229), .B(n5230), .Z(n5228) );
  XOR U8821 ( .A(DB[1893]), .B(DB[1878]), .Z(n5230) );
  AND U8822 ( .A(n522), .B(n5231), .Z(n5229) );
  XOR U8823 ( .A(n5232), .B(n5233), .Z(n5231) );
  XOR U8824 ( .A(DB[1878]), .B(DB[1863]), .Z(n5233) );
  AND U8825 ( .A(n526), .B(n5234), .Z(n5232) );
  XOR U8826 ( .A(n5235), .B(n5236), .Z(n5234) );
  XOR U8827 ( .A(DB[1863]), .B(DB[1848]), .Z(n5236) );
  AND U8828 ( .A(n530), .B(n5237), .Z(n5235) );
  XOR U8829 ( .A(n5238), .B(n5239), .Z(n5237) );
  XOR U8830 ( .A(DB[1848]), .B(DB[1833]), .Z(n5239) );
  AND U8831 ( .A(n534), .B(n5240), .Z(n5238) );
  XOR U8832 ( .A(n5241), .B(n5242), .Z(n5240) );
  XOR U8833 ( .A(DB[1833]), .B(DB[1818]), .Z(n5242) );
  AND U8834 ( .A(n538), .B(n5243), .Z(n5241) );
  XOR U8835 ( .A(n5244), .B(n5245), .Z(n5243) );
  XOR U8836 ( .A(DB[1818]), .B(DB[1803]), .Z(n5245) );
  AND U8837 ( .A(n542), .B(n5246), .Z(n5244) );
  XOR U8838 ( .A(n5247), .B(n5248), .Z(n5246) );
  XOR U8839 ( .A(DB[1803]), .B(DB[1788]), .Z(n5248) );
  AND U8840 ( .A(n546), .B(n5249), .Z(n5247) );
  XOR U8841 ( .A(n5250), .B(n5251), .Z(n5249) );
  XOR U8842 ( .A(DB[1788]), .B(DB[1773]), .Z(n5251) );
  AND U8843 ( .A(n550), .B(n5252), .Z(n5250) );
  XOR U8844 ( .A(n5253), .B(n5254), .Z(n5252) );
  XOR U8845 ( .A(DB[1773]), .B(DB[1758]), .Z(n5254) );
  AND U8846 ( .A(n554), .B(n5255), .Z(n5253) );
  XOR U8847 ( .A(n5256), .B(n5257), .Z(n5255) );
  XOR U8848 ( .A(DB[1758]), .B(DB[1743]), .Z(n5257) );
  AND U8849 ( .A(n558), .B(n5258), .Z(n5256) );
  XOR U8850 ( .A(n5259), .B(n5260), .Z(n5258) );
  XOR U8851 ( .A(DB[1743]), .B(DB[1728]), .Z(n5260) );
  AND U8852 ( .A(n562), .B(n5261), .Z(n5259) );
  XOR U8853 ( .A(n5262), .B(n5263), .Z(n5261) );
  XOR U8854 ( .A(DB[1728]), .B(DB[1713]), .Z(n5263) );
  AND U8855 ( .A(n566), .B(n5264), .Z(n5262) );
  XOR U8856 ( .A(n5265), .B(n5266), .Z(n5264) );
  XOR U8857 ( .A(DB[1713]), .B(DB[1698]), .Z(n5266) );
  AND U8858 ( .A(n570), .B(n5267), .Z(n5265) );
  XOR U8859 ( .A(n5268), .B(n5269), .Z(n5267) );
  XOR U8860 ( .A(DB[1698]), .B(DB[1683]), .Z(n5269) );
  AND U8861 ( .A(n574), .B(n5270), .Z(n5268) );
  XOR U8862 ( .A(n5271), .B(n5272), .Z(n5270) );
  XOR U8863 ( .A(DB[1683]), .B(DB[1668]), .Z(n5272) );
  AND U8864 ( .A(n578), .B(n5273), .Z(n5271) );
  XOR U8865 ( .A(n5274), .B(n5275), .Z(n5273) );
  XOR U8866 ( .A(DB[1668]), .B(DB[1653]), .Z(n5275) );
  AND U8867 ( .A(n582), .B(n5276), .Z(n5274) );
  XOR U8868 ( .A(n5277), .B(n5278), .Z(n5276) );
  XOR U8869 ( .A(DB[1653]), .B(DB[1638]), .Z(n5278) );
  AND U8870 ( .A(n586), .B(n5279), .Z(n5277) );
  XOR U8871 ( .A(n5280), .B(n5281), .Z(n5279) );
  XOR U8872 ( .A(DB[1638]), .B(DB[1623]), .Z(n5281) );
  AND U8873 ( .A(n590), .B(n5282), .Z(n5280) );
  XOR U8874 ( .A(n5283), .B(n5284), .Z(n5282) );
  XOR U8875 ( .A(DB[1623]), .B(DB[1608]), .Z(n5284) );
  AND U8876 ( .A(n594), .B(n5285), .Z(n5283) );
  XOR U8877 ( .A(n5286), .B(n5287), .Z(n5285) );
  XOR U8878 ( .A(DB[1608]), .B(DB[1593]), .Z(n5287) );
  AND U8879 ( .A(n598), .B(n5288), .Z(n5286) );
  XOR U8880 ( .A(n5289), .B(n5290), .Z(n5288) );
  XOR U8881 ( .A(DB[1593]), .B(DB[1578]), .Z(n5290) );
  AND U8882 ( .A(n602), .B(n5291), .Z(n5289) );
  XOR U8883 ( .A(n5292), .B(n5293), .Z(n5291) );
  XOR U8884 ( .A(DB[1578]), .B(DB[1563]), .Z(n5293) );
  AND U8885 ( .A(n606), .B(n5294), .Z(n5292) );
  XOR U8886 ( .A(n5295), .B(n5296), .Z(n5294) );
  XOR U8887 ( .A(DB[1563]), .B(DB[1548]), .Z(n5296) );
  AND U8888 ( .A(n610), .B(n5297), .Z(n5295) );
  XOR U8889 ( .A(n5298), .B(n5299), .Z(n5297) );
  XOR U8890 ( .A(DB[1548]), .B(DB[1533]), .Z(n5299) );
  AND U8891 ( .A(n614), .B(n5300), .Z(n5298) );
  XOR U8892 ( .A(n5301), .B(n5302), .Z(n5300) );
  XOR U8893 ( .A(DB[1533]), .B(DB[1518]), .Z(n5302) );
  AND U8894 ( .A(n618), .B(n5303), .Z(n5301) );
  XOR U8895 ( .A(n5304), .B(n5305), .Z(n5303) );
  XOR U8896 ( .A(DB[1518]), .B(DB[1503]), .Z(n5305) );
  AND U8897 ( .A(n622), .B(n5306), .Z(n5304) );
  XOR U8898 ( .A(n5307), .B(n5308), .Z(n5306) );
  XOR U8899 ( .A(DB[1503]), .B(DB[1488]), .Z(n5308) );
  AND U8900 ( .A(n626), .B(n5309), .Z(n5307) );
  XOR U8901 ( .A(n5310), .B(n5311), .Z(n5309) );
  XOR U8902 ( .A(DB[1488]), .B(DB[1473]), .Z(n5311) );
  AND U8903 ( .A(n630), .B(n5312), .Z(n5310) );
  XOR U8904 ( .A(n5313), .B(n5314), .Z(n5312) );
  XOR U8905 ( .A(DB[1473]), .B(DB[1458]), .Z(n5314) );
  AND U8906 ( .A(n634), .B(n5315), .Z(n5313) );
  XOR U8907 ( .A(n5316), .B(n5317), .Z(n5315) );
  XOR U8908 ( .A(DB[1458]), .B(DB[1443]), .Z(n5317) );
  AND U8909 ( .A(n638), .B(n5318), .Z(n5316) );
  XOR U8910 ( .A(n5319), .B(n5320), .Z(n5318) );
  XOR U8911 ( .A(DB[1443]), .B(DB[1428]), .Z(n5320) );
  AND U8912 ( .A(n642), .B(n5321), .Z(n5319) );
  XOR U8913 ( .A(n5322), .B(n5323), .Z(n5321) );
  XOR U8914 ( .A(DB[1428]), .B(DB[1413]), .Z(n5323) );
  AND U8915 ( .A(n646), .B(n5324), .Z(n5322) );
  XOR U8916 ( .A(n5325), .B(n5326), .Z(n5324) );
  XOR U8917 ( .A(DB[1413]), .B(DB[1398]), .Z(n5326) );
  AND U8918 ( .A(n650), .B(n5327), .Z(n5325) );
  XOR U8919 ( .A(n5328), .B(n5329), .Z(n5327) );
  XOR U8920 ( .A(DB[1398]), .B(DB[1383]), .Z(n5329) );
  AND U8921 ( .A(n654), .B(n5330), .Z(n5328) );
  XOR U8922 ( .A(n5331), .B(n5332), .Z(n5330) );
  XOR U8923 ( .A(DB[1383]), .B(DB[1368]), .Z(n5332) );
  AND U8924 ( .A(n658), .B(n5333), .Z(n5331) );
  XOR U8925 ( .A(n5334), .B(n5335), .Z(n5333) );
  XOR U8926 ( .A(DB[1368]), .B(DB[1353]), .Z(n5335) );
  AND U8927 ( .A(n662), .B(n5336), .Z(n5334) );
  XOR U8928 ( .A(n5337), .B(n5338), .Z(n5336) );
  XOR U8929 ( .A(DB[1353]), .B(DB[1338]), .Z(n5338) );
  AND U8930 ( .A(n666), .B(n5339), .Z(n5337) );
  XOR U8931 ( .A(n5340), .B(n5341), .Z(n5339) );
  XOR U8932 ( .A(DB[1338]), .B(DB[1323]), .Z(n5341) );
  AND U8933 ( .A(n670), .B(n5342), .Z(n5340) );
  XOR U8934 ( .A(n5343), .B(n5344), .Z(n5342) );
  XOR U8935 ( .A(DB[1323]), .B(DB[1308]), .Z(n5344) );
  AND U8936 ( .A(n674), .B(n5345), .Z(n5343) );
  XOR U8937 ( .A(n5346), .B(n5347), .Z(n5345) );
  XOR U8938 ( .A(DB[1308]), .B(DB[1293]), .Z(n5347) );
  AND U8939 ( .A(n678), .B(n5348), .Z(n5346) );
  XOR U8940 ( .A(n5349), .B(n5350), .Z(n5348) );
  XOR U8941 ( .A(DB[1293]), .B(DB[1278]), .Z(n5350) );
  AND U8942 ( .A(n682), .B(n5351), .Z(n5349) );
  XOR U8943 ( .A(n5352), .B(n5353), .Z(n5351) );
  XOR U8944 ( .A(DB[1278]), .B(DB[1263]), .Z(n5353) );
  AND U8945 ( .A(n686), .B(n5354), .Z(n5352) );
  XOR U8946 ( .A(n5355), .B(n5356), .Z(n5354) );
  XOR U8947 ( .A(DB[1263]), .B(DB[1248]), .Z(n5356) );
  AND U8948 ( .A(n690), .B(n5357), .Z(n5355) );
  XOR U8949 ( .A(n5358), .B(n5359), .Z(n5357) );
  XOR U8950 ( .A(DB[1248]), .B(DB[1233]), .Z(n5359) );
  AND U8951 ( .A(n694), .B(n5360), .Z(n5358) );
  XOR U8952 ( .A(n5361), .B(n5362), .Z(n5360) );
  XOR U8953 ( .A(DB[1233]), .B(DB[1218]), .Z(n5362) );
  AND U8954 ( .A(n698), .B(n5363), .Z(n5361) );
  XOR U8955 ( .A(n5364), .B(n5365), .Z(n5363) );
  XOR U8956 ( .A(DB[1218]), .B(DB[1203]), .Z(n5365) );
  AND U8957 ( .A(n702), .B(n5366), .Z(n5364) );
  XOR U8958 ( .A(n5367), .B(n5368), .Z(n5366) );
  XOR U8959 ( .A(DB[1203]), .B(DB[1188]), .Z(n5368) );
  AND U8960 ( .A(n706), .B(n5369), .Z(n5367) );
  XOR U8961 ( .A(n5370), .B(n5371), .Z(n5369) );
  XOR U8962 ( .A(DB[1188]), .B(DB[1173]), .Z(n5371) );
  AND U8963 ( .A(n710), .B(n5372), .Z(n5370) );
  XOR U8964 ( .A(n5373), .B(n5374), .Z(n5372) );
  XOR U8965 ( .A(DB[1173]), .B(DB[1158]), .Z(n5374) );
  AND U8966 ( .A(n714), .B(n5375), .Z(n5373) );
  XOR U8967 ( .A(n5376), .B(n5377), .Z(n5375) );
  XOR U8968 ( .A(DB[1158]), .B(DB[1143]), .Z(n5377) );
  AND U8969 ( .A(n718), .B(n5378), .Z(n5376) );
  XOR U8970 ( .A(n5379), .B(n5380), .Z(n5378) );
  XOR U8971 ( .A(DB[1143]), .B(DB[1128]), .Z(n5380) );
  AND U8972 ( .A(n722), .B(n5381), .Z(n5379) );
  XOR U8973 ( .A(n5382), .B(n5383), .Z(n5381) );
  XOR U8974 ( .A(DB[1128]), .B(DB[1113]), .Z(n5383) );
  AND U8975 ( .A(n726), .B(n5384), .Z(n5382) );
  XOR U8976 ( .A(n5385), .B(n5386), .Z(n5384) );
  XOR U8977 ( .A(DB[1113]), .B(DB[1098]), .Z(n5386) );
  AND U8978 ( .A(n730), .B(n5387), .Z(n5385) );
  XOR U8979 ( .A(n5388), .B(n5389), .Z(n5387) );
  XOR U8980 ( .A(DB[1098]), .B(DB[1083]), .Z(n5389) );
  AND U8981 ( .A(n734), .B(n5390), .Z(n5388) );
  XOR U8982 ( .A(n5391), .B(n5392), .Z(n5390) );
  XOR U8983 ( .A(DB[1083]), .B(DB[1068]), .Z(n5392) );
  AND U8984 ( .A(n738), .B(n5393), .Z(n5391) );
  XOR U8985 ( .A(n5394), .B(n5395), .Z(n5393) );
  XOR U8986 ( .A(DB[1068]), .B(DB[1053]), .Z(n5395) );
  AND U8987 ( .A(n742), .B(n5396), .Z(n5394) );
  XOR U8988 ( .A(n5397), .B(n5398), .Z(n5396) );
  XOR U8989 ( .A(DB[1053]), .B(DB[1038]), .Z(n5398) );
  AND U8990 ( .A(n746), .B(n5399), .Z(n5397) );
  XOR U8991 ( .A(n5400), .B(n5401), .Z(n5399) );
  XOR U8992 ( .A(DB[1038]), .B(DB[1023]), .Z(n5401) );
  AND U8993 ( .A(n750), .B(n5402), .Z(n5400) );
  XOR U8994 ( .A(n5403), .B(n5404), .Z(n5402) );
  XOR U8995 ( .A(DB[1023]), .B(DB[1008]), .Z(n5404) );
  AND U8996 ( .A(n754), .B(n5405), .Z(n5403) );
  XOR U8997 ( .A(n5406), .B(n5407), .Z(n5405) );
  XOR U8998 ( .A(DB[993]), .B(DB[1008]), .Z(n5407) );
  AND U8999 ( .A(n758), .B(n5408), .Z(n5406) );
  XOR U9000 ( .A(n5409), .B(n5410), .Z(n5408) );
  XOR U9001 ( .A(DB[993]), .B(DB[978]), .Z(n5410) );
  AND U9002 ( .A(n762), .B(n5411), .Z(n5409) );
  XOR U9003 ( .A(n5412), .B(n5413), .Z(n5411) );
  XOR U9004 ( .A(DB[978]), .B(DB[963]), .Z(n5413) );
  AND U9005 ( .A(n766), .B(n5414), .Z(n5412) );
  XOR U9006 ( .A(n5415), .B(n5416), .Z(n5414) );
  XOR U9007 ( .A(DB[963]), .B(DB[948]), .Z(n5416) );
  AND U9008 ( .A(n770), .B(n5417), .Z(n5415) );
  XOR U9009 ( .A(n5418), .B(n5419), .Z(n5417) );
  XOR U9010 ( .A(DB[948]), .B(DB[933]), .Z(n5419) );
  AND U9011 ( .A(n774), .B(n5420), .Z(n5418) );
  XOR U9012 ( .A(n5421), .B(n5422), .Z(n5420) );
  XOR U9013 ( .A(DB[933]), .B(DB[918]), .Z(n5422) );
  AND U9014 ( .A(n778), .B(n5423), .Z(n5421) );
  XOR U9015 ( .A(n5424), .B(n5425), .Z(n5423) );
  XOR U9016 ( .A(DB[918]), .B(DB[903]), .Z(n5425) );
  AND U9017 ( .A(n782), .B(n5426), .Z(n5424) );
  XOR U9018 ( .A(n5427), .B(n5428), .Z(n5426) );
  XOR U9019 ( .A(DB[903]), .B(DB[888]), .Z(n5428) );
  AND U9020 ( .A(n786), .B(n5429), .Z(n5427) );
  XOR U9021 ( .A(n5430), .B(n5431), .Z(n5429) );
  XOR U9022 ( .A(DB[888]), .B(DB[873]), .Z(n5431) );
  AND U9023 ( .A(n790), .B(n5432), .Z(n5430) );
  XOR U9024 ( .A(n5433), .B(n5434), .Z(n5432) );
  XOR U9025 ( .A(DB[873]), .B(DB[858]), .Z(n5434) );
  AND U9026 ( .A(n794), .B(n5435), .Z(n5433) );
  XOR U9027 ( .A(n5436), .B(n5437), .Z(n5435) );
  XOR U9028 ( .A(DB[858]), .B(DB[843]), .Z(n5437) );
  AND U9029 ( .A(n798), .B(n5438), .Z(n5436) );
  XOR U9030 ( .A(n5439), .B(n5440), .Z(n5438) );
  XOR U9031 ( .A(DB[843]), .B(DB[828]), .Z(n5440) );
  AND U9032 ( .A(n802), .B(n5441), .Z(n5439) );
  XOR U9033 ( .A(n5442), .B(n5443), .Z(n5441) );
  XOR U9034 ( .A(DB[828]), .B(DB[813]), .Z(n5443) );
  AND U9035 ( .A(n806), .B(n5444), .Z(n5442) );
  XOR U9036 ( .A(n5445), .B(n5446), .Z(n5444) );
  XOR U9037 ( .A(DB[813]), .B(DB[798]), .Z(n5446) );
  AND U9038 ( .A(n810), .B(n5447), .Z(n5445) );
  XOR U9039 ( .A(n5448), .B(n5449), .Z(n5447) );
  XOR U9040 ( .A(DB[798]), .B(DB[783]), .Z(n5449) );
  AND U9041 ( .A(n814), .B(n5450), .Z(n5448) );
  XOR U9042 ( .A(n5451), .B(n5452), .Z(n5450) );
  XOR U9043 ( .A(DB[783]), .B(DB[768]), .Z(n5452) );
  AND U9044 ( .A(n818), .B(n5453), .Z(n5451) );
  XOR U9045 ( .A(n5454), .B(n5455), .Z(n5453) );
  XOR U9046 ( .A(DB[768]), .B(DB[753]), .Z(n5455) );
  AND U9047 ( .A(n822), .B(n5456), .Z(n5454) );
  XOR U9048 ( .A(n5457), .B(n5458), .Z(n5456) );
  XOR U9049 ( .A(DB[753]), .B(DB[738]), .Z(n5458) );
  AND U9050 ( .A(n826), .B(n5459), .Z(n5457) );
  XOR U9051 ( .A(n5460), .B(n5461), .Z(n5459) );
  XOR U9052 ( .A(DB[738]), .B(DB[723]), .Z(n5461) );
  AND U9053 ( .A(n830), .B(n5462), .Z(n5460) );
  XOR U9054 ( .A(n5463), .B(n5464), .Z(n5462) );
  XOR U9055 ( .A(DB[723]), .B(DB[708]), .Z(n5464) );
  AND U9056 ( .A(n834), .B(n5465), .Z(n5463) );
  XOR U9057 ( .A(n5466), .B(n5467), .Z(n5465) );
  XOR U9058 ( .A(DB[708]), .B(DB[693]), .Z(n5467) );
  AND U9059 ( .A(n838), .B(n5468), .Z(n5466) );
  XOR U9060 ( .A(n5469), .B(n5470), .Z(n5468) );
  XOR U9061 ( .A(DB[693]), .B(DB[678]), .Z(n5470) );
  AND U9062 ( .A(n842), .B(n5471), .Z(n5469) );
  XOR U9063 ( .A(n5472), .B(n5473), .Z(n5471) );
  XOR U9064 ( .A(DB[678]), .B(DB[663]), .Z(n5473) );
  AND U9065 ( .A(n846), .B(n5474), .Z(n5472) );
  XOR U9066 ( .A(n5475), .B(n5476), .Z(n5474) );
  XOR U9067 ( .A(DB[663]), .B(DB[648]), .Z(n5476) );
  AND U9068 ( .A(n850), .B(n5477), .Z(n5475) );
  XOR U9069 ( .A(n5478), .B(n5479), .Z(n5477) );
  XOR U9070 ( .A(DB[648]), .B(DB[633]), .Z(n5479) );
  AND U9071 ( .A(n854), .B(n5480), .Z(n5478) );
  XOR U9072 ( .A(n5481), .B(n5482), .Z(n5480) );
  XOR U9073 ( .A(DB[633]), .B(DB[618]), .Z(n5482) );
  AND U9074 ( .A(n858), .B(n5483), .Z(n5481) );
  XOR U9075 ( .A(n5484), .B(n5485), .Z(n5483) );
  XOR U9076 ( .A(DB[618]), .B(DB[603]), .Z(n5485) );
  AND U9077 ( .A(n862), .B(n5486), .Z(n5484) );
  XOR U9078 ( .A(n5487), .B(n5488), .Z(n5486) );
  XOR U9079 ( .A(DB[603]), .B(DB[588]), .Z(n5488) );
  AND U9080 ( .A(n866), .B(n5489), .Z(n5487) );
  XOR U9081 ( .A(n5490), .B(n5491), .Z(n5489) );
  XOR U9082 ( .A(DB[588]), .B(DB[573]), .Z(n5491) );
  AND U9083 ( .A(n870), .B(n5492), .Z(n5490) );
  XOR U9084 ( .A(n5493), .B(n5494), .Z(n5492) );
  XOR U9085 ( .A(DB[573]), .B(DB[558]), .Z(n5494) );
  AND U9086 ( .A(n874), .B(n5495), .Z(n5493) );
  XOR U9087 ( .A(n5496), .B(n5497), .Z(n5495) );
  XOR U9088 ( .A(DB[558]), .B(DB[543]), .Z(n5497) );
  AND U9089 ( .A(n878), .B(n5498), .Z(n5496) );
  XOR U9090 ( .A(n5499), .B(n5500), .Z(n5498) );
  XOR U9091 ( .A(DB[543]), .B(DB[528]), .Z(n5500) );
  AND U9092 ( .A(n882), .B(n5501), .Z(n5499) );
  XOR U9093 ( .A(n5502), .B(n5503), .Z(n5501) );
  XOR U9094 ( .A(DB[528]), .B(DB[513]), .Z(n5503) );
  AND U9095 ( .A(n886), .B(n5504), .Z(n5502) );
  XOR U9096 ( .A(n5505), .B(n5506), .Z(n5504) );
  XOR U9097 ( .A(DB[513]), .B(DB[498]), .Z(n5506) );
  AND U9098 ( .A(n890), .B(n5507), .Z(n5505) );
  XOR U9099 ( .A(n5508), .B(n5509), .Z(n5507) );
  XOR U9100 ( .A(DB[498]), .B(DB[483]), .Z(n5509) );
  AND U9101 ( .A(n894), .B(n5510), .Z(n5508) );
  XOR U9102 ( .A(n5511), .B(n5512), .Z(n5510) );
  XOR U9103 ( .A(DB[483]), .B(DB[468]), .Z(n5512) );
  AND U9104 ( .A(n898), .B(n5513), .Z(n5511) );
  XOR U9105 ( .A(n5514), .B(n5515), .Z(n5513) );
  XOR U9106 ( .A(DB[468]), .B(DB[453]), .Z(n5515) );
  AND U9107 ( .A(n902), .B(n5516), .Z(n5514) );
  XOR U9108 ( .A(n5517), .B(n5518), .Z(n5516) );
  XOR U9109 ( .A(DB[453]), .B(DB[438]), .Z(n5518) );
  AND U9110 ( .A(n906), .B(n5519), .Z(n5517) );
  XOR U9111 ( .A(n5520), .B(n5521), .Z(n5519) );
  XOR U9112 ( .A(DB[438]), .B(DB[423]), .Z(n5521) );
  AND U9113 ( .A(n910), .B(n5522), .Z(n5520) );
  XOR U9114 ( .A(n5523), .B(n5524), .Z(n5522) );
  XOR U9115 ( .A(DB[423]), .B(DB[408]), .Z(n5524) );
  AND U9116 ( .A(n914), .B(n5525), .Z(n5523) );
  XOR U9117 ( .A(n5526), .B(n5527), .Z(n5525) );
  XOR U9118 ( .A(DB[408]), .B(DB[393]), .Z(n5527) );
  AND U9119 ( .A(n918), .B(n5528), .Z(n5526) );
  XOR U9120 ( .A(n5529), .B(n5530), .Z(n5528) );
  XOR U9121 ( .A(DB[393]), .B(DB[378]), .Z(n5530) );
  AND U9122 ( .A(n922), .B(n5531), .Z(n5529) );
  XOR U9123 ( .A(n5532), .B(n5533), .Z(n5531) );
  XOR U9124 ( .A(DB[378]), .B(DB[363]), .Z(n5533) );
  AND U9125 ( .A(n926), .B(n5534), .Z(n5532) );
  XOR U9126 ( .A(n5535), .B(n5536), .Z(n5534) );
  XOR U9127 ( .A(DB[363]), .B(DB[348]), .Z(n5536) );
  AND U9128 ( .A(n930), .B(n5537), .Z(n5535) );
  XOR U9129 ( .A(n5538), .B(n5539), .Z(n5537) );
  XOR U9130 ( .A(DB[348]), .B(DB[333]), .Z(n5539) );
  AND U9131 ( .A(n934), .B(n5540), .Z(n5538) );
  XOR U9132 ( .A(n5541), .B(n5542), .Z(n5540) );
  XOR U9133 ( .A(DB[333]), .B(DB[318]), .Z(n5542) );
  AND U9134 ( .A(n938), .B(n5543), .Z(n5541) );
  XOR U9135 ( .A(n5544), .B(n5545), .Z(n5543) );
  XOR U9136 ( .A(DB[318]), .B(DB[303]), .Z(n5545) );
  AND U9137 ( .A(n942), .B(n5546), .Z(n5544) );
  XOR U9138 ( .A(n5547), .B(n5548), .Z(n5546) );
  XOR U9139 ( .A(DB[303]), .B(DB[288]), .Z(n5548) );
  AND U9140 ( .A(n946), .B(n5549), .Z(n5547) );
  XOR U9141 ( .A(n5550), .B(n5551), .Z(n5549) );
  XOR U9142 ( .A(DB[288]), .B(DB[273]), .Z(n5551) );
  AND U9143 ( .A(n950), .B(n5552), .Z(n5550) );
  XOR U9144 ( .A(n5553), .B(n5554), .Z(n5552) );
  XOR U9145 ( .A(DB[273]), .B(DB[258]), .Z(n5554) );
  AND U9146 ( .A(n954), .B(n5555), .Z(n5553) );
  XOR U9147 ( .A(n5556), .B(n5557), .Z(n5555) );
  XOR U9148 ( .A(DB[258]), .B(DB[243]), .Z(n5557) );
  AND U9149 ( .A(n958), .B(n5558), .Z(n5556) );
  XOR U9150 ( .A(n5559), .B(n5560), .Z(n5558) );
  XOR U9151 ( .A(DB[243]), .B(DB[228]), .Z(n5560) );
  AND U9152 ( .A(n962), .B(n5561), .Z(n5559) );
  XOR U9153 ( .A(n5562), .B(n5563), .Z(n5561) );
  XOR U9154 ( .A(DB[228]), .B(DB[213]), .Z(n5563) );
  AND U9155 ( .A(n966), .B(n5564), .Z(n5562) );
  XOR U9156 ( .A(n5565), .B(n5566), .Z(n5564) );
  XOR U9157 ( .A(DB[213]), .B(DB[198]), .Z(n5566) );
  AND U9158 ( .A(n970), .B(n5567), .Z(n5565) );
  XOR U9159 ( .A(n5568), .B(n5569), .Z(n5567) );
  XOR U9160 ( .A(DB[198]), .B(DB[183]), .Z(n5569) );
  AND U9161 ( .A(n974), .B(n5570), .Z(n5568) );
  XOR U9162 ( .A(n5571), .B(n5572), .Z(n5570) );
  XOR U9163 ( .A(DB[183]), .B(DB[168]), .Z(n5572) );
  AND U9164 ( .A(n978), .B(n5573), .Z(n5571) );
  XOR U9165 ( .A(n5574), .B(n5575), .Z(n5573) );
  XOR U9166 ( .A(DB[168]), .B(DB[153]), .Z(n5575) );
  AND U9167 ( .A(n982), .B(n5576), .Z(n5574) );
  XOR U9168 ( .A(n5577), .B(n5578), .Z(n5576) );
  XOR U9169 ( .A(DB[153]), .B(DB[138]), .Z(n5578) );
  AND U9170 ( .A(n986), .B(n5579), .Z(n5577) );
  XOR U9171 ( .A(n5580), .B(n5581), .Z(n5579) );
  XOR U9172 ( .A(DB[138]), .B(DB[123]), .Z(n5581) );
  AND U9173 ( .A(n990), .B(n5582), .Z(n5580) );
  XOR U9174 ( .A(n5583), .B(n5584), .Z(n5582) );
  XOR U9175 ( .A(DB[123]), .B(DB[108]), .Z(n5584) );
  AND U9176 ( .A(n994), .B(n5585), .Z(n5583) );
  XOR U9177 ( .A(n5586), .B(n5587), .Z(n5585) );
  XOR U9178 ( .A(DB[93]), .B(DB[108]), .Z(n5587) );
  AND U9179 ( .A(n998), .B(n5588), .Z(n5586) );
  XOR U9180 ( .A(n5589), .B(n5590), .Z(n5588) );
  XOR U9181 ( .A(DB[93]), .B(DB[78]), .Z(n5590) );
  AND U9182 ( .A(n1002), .B(n5591), .Z(n5589) );
  XOR U9183 ( .A(n5592), .B(n5593), .Z(n5591) );
  XOR U9184 ( .A(DB[78]), .B(DB[63]), .Z(n5593) );
  AND U9185 ( .A(n1006), .B(n5594), .Z(n5592) );
  XOR U9186 ( .A(n5595), .B(n5596), .Z(n5594) );
  XOR U9187 ( .A(DB[63]), .B(DB[48]), .Z(n5596) );
  AND U9188 ( .A(n1010), .B(n5597), .Z(n5595) );
  XOR U9189 ( .A(n5598), .B(n5599), .Z(n5597) );
  XOR U9190 ( .A(DB[48]), .B(DB[33]), .Z(n5599) );
  AND U9191 ( .A(n1014), .B(n5600), .Z(n5598) );
  XOR U9192 ( .A(n5601), .B(n5602), .Z(n5600) );
  XOR U9193 ( .A(DB[33]), .B(DB[18]), .Z(n5602) );
  AND U9194 ( .A(n1018), .B(n5603), .Z(n5601) );
  XOR U9195 ( .A(DB[3]), .B(DB[18]), .Z(n5603) );
  XOR U9196 ( .A(DB[3827]), .B(n5604), .Z(min_val_out[2]) );
  AND U9197 ( .A(n2), .B(n5605), .Z(n5604) );
  XOR U9198 ( .A(n5606), .B(n5607), .Z(n5605) );
  XOR U9199 ( .A(DB[3827]), .B(DB[3812]), .Z(n5607) );
  AND U9200 ( .A(n6), .B(n5608), .Z(n5606) );
  XOR U9201 ( .A(n5609), .B(n5610), .Z(n5608) );
  XOR U9202 ( .A(DB[3812]), .B(DB[3797]), .Z(n5610) );
  AND U9203 ( .A(n10), .B(n5611), .Z(n5609) );
  XOR U9204 ( .A(n5612), .B(n5613), .Z(n5611) );
  XOR U9205 ( .A(DB[3797]), .B(DB[3782]), .Z(n5613) );
  AND U9206 ( .A(n14), .B(n5614), .Z(n5612) );
  XOR U9207 ( .A(n5615), .B(n5616), .Z(n5614) );
  XOR U9208 ( .A(DB[3782]), .B(DB[3767]), .Z(n5616) );
  AND U9209 ( .A(n18), .B(n5617), .Z(n5615) );
  XOR U9210 ( .A(n5618), .B(n5619), .Z(n5617) );
  XOR U9211 ( .A(DB[3767]), .B(DB[3752]), .Z(n5619) );
  AND U9212 ( .A(n22), .B(n5620), .Z(n5618) );
  XOR U9213 ( .A(n5621), .B(n5622), .Z(n5620) );
  XOR U9214 ( .A(DB[3752]), .B(DB[3737]), .Z(n5622) );
  AND U9215 ( .A(n26), .B(n5623), .Z(n5621) );
  XOR U9216 ( .A(n5624), .B(n5625), .Z(n5623) );
  XOR U9217 ( .A(DB[3737]), .B(DB[3722]), .Z(n5625) );
  AND U9218 ( .A(n30), .B(n5626), .Z(n5624) );
  XOR U9219 ( .A(n5627), .B(n5628), .Z(n5626) );
  XOR U9220 ( .A(DB[3722]), .B(DB[3707]), .Z(n5628) );
  AND U9221 ( .A(n34), .B(n5629), .Z(n5627) );
  XOR U9222 ( .A(n5630), .B(n5631), .Z(n5629) );
  XOR U9223 ( .A(DB[3707]), .B(DB[3692]), .Z(n5631) );
  AND U9224 ( .A(n38), .B(n5632), .Z(n5630) );
  XOR U9225 ( .A(n5633), .B(n5634), .Z(n5632) );
  XOR U9226 ( .A(DB[3692]), .B(DB[3677]), .Z(n5634) );
  AND U9227 ( .A(n42), .B(n5635), .Z(n5633) );
  XOR U9228 ( .A(n5636), .B(n5637), .Z(n5635) );
  XOR U9229 ( .A(DB[3677]), .B(DB[3662]), .Z(n5637) );
  AND U9230 ( .A(n46), .B(n5638), .Z(n5636) );
  XOR U9231 ( .A(n5639), .B(n5640), .Z(n5638) );
  XOR U9232 ( .A(DB[3662]), .B(DB[3647]), .Z(n5640) );
  AND U9233 ( .A(n50), .B(n5641), .Z(n5639) );
  XOR U9234 ( .A(n5642), .B(n5643), .Z(n5641) );
  XOR U9235 ( .A(DB[3647]), .B(DB[3632]), .Z(n5643) );
  AND U9236 ( .A(n54), .B(n5644), .Z(n5642) );
  XOR U9237 ( .A(n5645), .B(n5646), .Z(n5644) );
  XOR U9238 ( .A(DB[3632]), .B(DB[3617]), .Z(n5646) );
  AND U9239 ( .A(n58), .B(n5647), .Z(n5645) );
  XOR U9240 ( .A(n5648), .B(n5649), .Z(n5647) );
  XOR U9241 ( .A(DB[3617]), .B(DB[3602]), .Z(n5649) );
  AND U9242 ( .A(n62), .B(n5650), .Z(n5648) );
  XOR U9243 ( .A(n5651), .B(n5652), .Z(n5650) );
  XOR U9244 ( .A(DB[3602]), .B(DB[3587]), .Z(n5652) );
  AND U9245 ( .A(n66), .B(n5653), .Z(n5651) );
  XOR U9246 ( .A(n5654), .B(n5655), .Z(n5653) );
  XOR U9247 ( .A(DB[3587]), .B(DB[3572]), .Z(n5655) );
  AND U9248 ( .A(n70), .B(n5656), .Z(n5654) );
  XOR U9249 ( .A(n5657), .B(n5658), .Z(n5656) );
  XOR U9250 ( .A(DB[3572]), .B(DB[3557]), .Z(n5658) );
  AND U9251 ( .A(n74), .B(n5659), .Z(n5657) );
  XOR U9252 ( .A(n5660), .B(n5661), .Z(n5659) );
  XOR U9253 ( .A(DB[3557]), .B(DB[3542]), .Z(n5661) );
  AND U9254 ( .A(n78), .B(n5662), .Z(n5660) );
  XOR U9255 ( .A(n5663), .B(n5664), .Z(n5662) );
  XOR U9256 ( .A(DB[3542]), .B(DB[3527]), .Z(n5664) );
  AND U9257 ( .A(n82), .B(n5665), .Z(n5663) );
  XOR U9258 ( .A(n5666), .B(n5667), .Z(n5665) );
  XOR U9259 ( .A(DB[3527]), .B(DB[3512]), .Z(n5667) );
  AND U9260 ( .A(n86), .B(n5668), .Z(n5666) );
  XOR U9261 ( .A(n5669), .B(n5670), .Z(n5668) );
  XOR U9262 ( .A(DB[3512]), .B(DB[3497]), .Z(n5670) );
  AND U9263 ( .A(n90), .B(n5671), .Z(n5669) );
  XOR U9264 ( .A(n5672), .B(n5673), .Z(n5671) );
  XOR U9265 ( .A(DB[3497]), .B(DB[3482]), .Z(n5673) );
  AND U9266 ( .A(n94), .B(n5674), .Z(n5672) );
  XOR U9267 ( .A(n5675), .B(n5676), .Z(n5674) );
  XOR U9268 ( .A(DB[3482]), .B(DB[3467]), .Z(n5676) );
  AND U9269 ( .A(n98), .B(n5677), .Z(n5675) );
  XOR U9270 ( .A(n5678), .B(n5679), .Z(n5677) );
  XOR U9271 ( .A(DB[3467]), .B(DB[3452]), .Z(n5679) );
  AND U9272 ( .A(n102), .B(n5680), .Z(n5678) );
  XOR U9273 ( .A(n5681), .B(n5682), .Z(n5680) );
  XOR U9274 ( .A(DB[3452]), .B(DB[3437]), .Z(n5682) );
  AND U9275 ( .A(n106), .B(n5683), .Z(n5681) );
  XOR U9276 ( .A(n5684), .B(n5685), .Z(n5683) );
  XOR U9277 ( .A(DB[3437]), .B(DB[3422]), .Z(n5685) );
  AND U9278 ( .A(n110), .B(n5686), .Z(n5684) );
  XOR U9279 ( .A(n5687), .B(n5688), .Z(n5686) );
  XOR U9280 ( .A(DB[3422]), .B(DB[3407]), .Z(n5688) );
  AND U9281 ( .A(n114), .B(n5689), .Z(n5687) );
  XOR U9282 ( .A(n5690), .B(n5691), .Z(n5689) );
  XOR U9283 ( .A(DB[3407]), .B(DB[3392]), .Z(n5691) );
  AND U9284 ( .A(n118), .B(n5692), .Z(n5690) );
  XOR U9285 ( .A(n5693), .B(n5694), .Z(n5692) );
  XOR U9286 ( .A(DB[3392]), .B(DB[3377]), .Z(n5694) );
  AND U9287 ( .A(n122), .B(n5695), .Z(n5693) );
  XOR U9288 ( .A(n5696), .B(n5697), .Z(n5695) );
  XOR U9289 ( .A(DB[3377]), .B(DB[3362]), .Z(n5697) );
  AND U9290 ( .A(n126), .B(n5698), .Z(n5696) );
  XOR U9291 ( .A(n5699), .B(n5700), .Z(n5698) );
  XOR U9292 ( .A(DB[3362]), .B(DB[3347]), .Z(n5700) );
  AND U9293 ( .A(n130), .B(n5701), .Z(n5699) );
  XOR U9294 ( .A(n5702), .B(n5703), .Z(n5701) );
  XOR U9295 ( .A(DB[3347]), .B(DB[3332]), .Z(n5703) );
  AND U9296 ( .A(n134), .B(n5704), .Z(n5702) );
  XOR U9297 ( .A(n5705), .B(n5706), .Z(n5704) );
  XOR U9298 ( .A(DB[3332]), .B(DB[3317]), .Z(n5706) );
  AND U9299 ( .A(n138), .B(n5707), .Z(n5705) );
  XOR U9300 ( .A(n5708), .B(n5709), .Z(n5707) );
  XOR U9301 ( .A(DB[3317]), .B(DB[3302]), .Z(n5709) );
  AND U9302 ( .A(n142), .B(n5710), .Z(n5708) );
  XOR U9303 ( .A(n5711), .B(n5712), .Z(n5710) );
  XOR U9304 ( .A(DB[3302]), .B(DB[3287]), .Z(n5712) );
  AND U9305 ( .A(n146), .B(n5713), .Z(n5711) );
  XOR U9306 ( .A(n5714), .B(n5715), .Z(n5713) );
  XOR U9307 ( .A(DB[3287]), .B(DB[3272]), .Z(n5715) );
  AND U9308 ( .A(n150), .B(n5716), .Z(n5714) );
  XOR U9309 ( .A(n5717), .B(n5718), .Z(n5716) );
  XOR U9310 ( .A(DB[3272]), .B(DB[3257]), .Z(n5718) );
  AND U9311 ( .A(n154), .B(n5719), .Z(n5717) );
  XOR U9312 ( .A(n5720), .B(n5721), .Z(n5719) );
  XOR U9313 ( .A(DB[3257]), .B(DB[3242]), .Z(n5721) );
  AND U9314 ( .A(n158), .B(n5722), .Z(n5720) );
  XOR U9315 ( .A(n5723), .B(n5724), .Z(n5722) );
  XOR U9316 ( .A(DB[3242]), .B(DB[3227]), .Z(n5724) );
  AND U9317 ( .A(n162), .B(n5725), .Z(n5723) );
  XOR U9318 ( .A(n5726), .B(n5727), .Z(n5725) );
  XOR U9319 ( .A(DB[3227]), .B(DB[3212]), .Z(n5727) );
  AND U9320 ( .A(n166), .B(n5728), .Z(n5726) );
  XOR U9321 ( .A(n5729), .B(n5730), .Z(n5728) );
  XOR U9322 ( .A(DB[3212]), .B(DB[3197]), .Z(n5730) );
  AND U9323 ( .A(n170), .B(n5731), .Z(n5729) );
  XOR U9324 ( .A(n5732), .B(n5733), .Z(n5731) );
  XOR U9325 ( .A(DB[3197]), .B(DB[3182]), .Z(n5733) );
  AND U9326 ( .A(n174), .B(n5734), .Z(n5732) );
  XOR U9327 ( .A(n5735), .B(n5736), .Z(n5734) );
  XOR U9328 ( .A(DB[3182]), .B(DB[3167]), .Z(n5736) );
  AND U9329 ( .A(n178), .B(n5737), .Z(n5735) );
  XOR U9330 ( .A(n5738), .B(n5739), .Z(n5737) );
  XOR U9331 ( .A(DB[3167]), .B(DB[3152]), .Z(n5739) );
  AND U9332 ( .A(n182), .B(n5740), .Z(n5738) );
  XOR U9333 ( .A(n5741), .B(n5742), .Z(n5740) );
  XOR U9334 ( .A(DB[3152]), .B(DB[3137]), .Z(n5742) );
  AND U9335 ( .A(n186), .B(n5743), .Z(n5741) );
  XOR U9336 ( .A(n5744), .B(n5745), .Z(n5743) );
  XOR U9337 ( .A(DB[3137]), .B(DB[3122]), .Z(n5745) );
  AND U9338 ( .A(n190), .B(n5746), .Z(n5744) );
  XOR U9339 ( .A(n5747), .B(n5748), .Z(n5746) );
  XOR U9340 ( .A(DB[3122]), .B(DB[3107]), .Z(n5748) );
  AND U9341 ( .A(n194), .B(n5749), .Z(n5747) );
  XOR U9342 ( .A(n5750), .B(n5751), .Z(n5749) );
  XOR U9343 ( .A(DB[3107]), .B(DB[3092]), .Z(n5751) );
  AND U9344 ( .A(n198), .B(n5752), .Z(n5750) );
  XOR U9345 ( .A(n5753), .B(n5754), .Z(n5752) );
  XOR U9346 ( .A(DB[3092]), .B(DB[3077]), .Z(n5754) );
  AND U9347 ( .A(n202), .B(n5755), .Z(n5753) );
  XOR U9348 ( .A(n5756), .B(n5757), .Z(n5755) );
  XOR U9349 ( .A(DB[3077]), .B(DB[3062]), .Z(n5757) );
  AND U9350 ( .A(n206), .B(n5758), .Z(n5756) );
  XOR U9351 ( .A(n5759), .B(n5760), .Z(n5758) );
  XOR U9352 ( .A(DB[3062]), .B(DB[3047]), .Z(n5760) );
  AND U9353 ( .A(n210), .B(n5761), .Z(n5759) );
  XOR U9354 ( .A(n5762), .B(n5763), .Z(n5761) );
  XOR U9355 ( .A(DB[3047]), .B(DB[3032]), .Z(n5763) );
  AND U9356 ( .A(n214), .B(n5764), .Z(n5762) );
  XOR U9357 ( .A(n5765), .B(n5766), .Z(n5764) );
  XOR U9358 ( .A(DB[3032]), .B(DB[3017]), .Z(n5766) );
  AND U9359 ( .A(n218), .B(n5767), .Z(n5765) );
  XOR U9360 ( .A(n5768), .B(n5769), .Z(n5767) );
  XOR U9361 ( .A(DB[3017]), .B(DB[3002]), .Z(n5769) );
  AND U9362 ( .A(n222), .B(n5770), .Z(n5768) );
  XOR U9363 ( .A(n5771), .B(n5772), .Z(n5770) );
  XOR U9364 ( .A(DB[3002]), .B(DB[2987]), .Z(n5772) );
  AND U9365 ( .A(n226), .B(n5773), .Z(n5771) );
  XOR U9366 ( .A(n5774), .B(n5775), .Z(n5773) );
  XOR U9367 ( .A(DB[2987]), .B(DB[2972]), .Z(n5775) );
  AND U9368 ( .A(n230), .B(n5776), .Z(n5774) );
  XOR U9369 ( .A(n5777), .B(n5778), .Z(n5776) );
  XOR U9370 ( .A(DB[2972]), .B(DB[2957]), .Z(n5778) );
  AND U9371 ( .A(n234), .B(n5779), .Z(n5777) );
  XOR U9372 ( .A(n5780), .B(n5781), .Z(n5779) );
  XOR U9373 ( .A(DB[2957]), .B(DB[2942]), .Z(n5781) );
  AND U9374 ( .A(n238), .B(n5782), .Z(n5780) );
  XOR U9375 ( .A(n5783), .B(n5784), .Z(n5782) );
  XOR U9376 ( .A(DB[2942]), .B(DB[2927]), .Z(n5784) );
  AND U9377 ( .A(n242), .B(n5785), .Z(n5783) );
  XOR U9378 ( .A(n5786), .B(n5787), .Z(n5785) );
  XOR U9379 ( .A(DB[2927]), .B(DB[2912]), .Z(n5787) );
  AND U9380 ( .A(n246), .B(n5788), .Z(n5786) );
  XOR U9381 ( .A(n5789), .B(n5790), .Z(n5788) );
  XOR U9382 ( .A(DB[2912]), .B(DB[2897]), .Z(n5790) );
  AND U9383 ( .A(n250), .B(n5791), .Z(n5789) );
  XOR U9384 ( .A(n5792), .B(n5793), .Z(n5791) );
  XOR U9385 ( .A(DB[2897]), .B(DB[2882]), .Z(n5793) );
  AND U9386 ( .A(n254), .B(n5794), .Z(n5792) );
  XOR U9387 ( .A(n5795), .B(n5796), .Z(n5794) );
  XOR U9388 ( .A(DB[2882]), .B(DB[2867]), .Z(n5796) );
  AND U9389 ( .A(n258), .B(n5797), .Z(n5795) );
  XOR U9390 ( .A(n5798), .B(n5799), .Z(n5797) );
  XOR U9391 ( .A(DB[2867]), .B(DB[2852]), .Z(n5799) );
  AND U9392 ( .A(n262), .B(n5800), .Z(n5798) );
  XOR U9393 ( .A(n5801), .B(n5802), .Z(n5800) );
  XOR U9394 ( .A(DB[2852]), .B(DB[2837]), .Z(n5802) );
  AND U9395 ( .A(n266), .B(n5803), .Z(n5801) );
  XOR U9396 ( .A(n5804), .B(n5805), .Z(n5803) );
  XOR U9397 ( .A(DB[2837]), .B(DB[2822]), .Z(n5805) );
  AND U9398 ( .A(n270), .B(n5806), .Z(n5804) );
  XOR U9399 ( .A(n5807), .B(n5808), .Z(n5806) );
  XOR U9400 ( .A(DB[2822]), .B(DB[2807]), .Z(n5808) );
  AND U9401 ( .A(n274), .B(n5809), .Z(n5807) );
  XOR U9402 ( .A(n5810), .B(n5811), .Z(n5809) );
  XOR U9403 ( .A(DB[2807]), .B(DB[2792]), .Z(n5811) );
  AND U9404 ( .A(n278), .B(n5812), .Z(n5810) );
  XOR U9405 ( .A(n5813), .B(n5814), .Z(n5812) );
  XOR U9406 ( .A(DB[2792]), .B(DB[2777]), .Z(n5814) );
  AND U9407 ( .A(n282), .B(n5815), .Z(n5813) );
  XOR U9408 ( .A(n5816), .B(n5817), .Z(n5815) );
  XOR U9409 ( .A(DB[2777]), .B(DB[2762]), .Z(n5817) );
  AND U9410 ( .A(n286), .B(n5818), .Z(n5816) );
  XOR U9411 ( .A(n5819), .B(n5820), .Z(n5818) );
  XOR U9412 ( .A(DB[2762]), .B(DB[2747]), .Z(n5820) );
  AND U9413 ( .A(n290), .B(n5821), .Z(n5819) );
  XOR U9414 ( .A(n5822), .B(n5823), .Z(n5821) );
  XOR U9415 ( .A(DB[2747]), .B(DB[2732]), .Z(n5823) );
  AND U9416 ( .A(n294), .B(n5824), .Z(n5822) );
  XOR U9417 ( .A(n5825), .B(n5826), .Z(n5824) );
  XOR U9418 ( .A(DB[2732]), .B(DB[2717]), .Z(n5826) );
  AND U9419 ( .A(n298), .B(n5827), .Z(n5825) );
  XOR U9420 ( .A(n5828), .B(n5829), .Z(n5827) );
  XOR U9421 ( .A(DB[2717]), .B(DB[2702]), .Z(n5829) );
  AND U9422 ( .A(n302), .B(n5830), .Z(n5828) );
  XOR U9423 ( .A(n5831), .B(n5832), .Z(n5830) );
  XOR U9424 ( .A(DB[2702]), .B(DB[2687]), .Z(n5832) );
  AND U9425 ( .A(n306), .B(n5833), .Z(n5831) );
  XOR U9426 ( .A(n5834), .B(n5835), .Z(n5833) );
  XOR U9427 ( .A(DB[2687]), .B(DB[2672]), .Z(n5835) );
  AND U9428 ( .A(n310), .B(n5836), .Z(n5834) );
  XOR U9429 ( .A(n5837), .B(n5838), .Z(n5836) );
  XOR U9430 ( .A(DB[2672]), .B(DB[2657]), .Z(n5838) );
  AND U9431 ( .A(n314), .B(n5839), .Z(n5837) );
  XOR U9432 ( .A(n5840), .B(n5841), .Z(n5839) );
  XOR U9433 ( .A(DB[2657]), .B(DB[2642]), .Z(n5841) );
  AND U9434 ( .A(n318), .B(n5842), .Z(n5840) );
  XOR U9435 ( .A(n5843), .B(n5844), .Z(n5842) );
  XOR U9436 ( .A(DB[2642]), .B(DB[2627]), .Z(n5844) );
  AND U9437 ( .A(n322), .B(n5845), .Z(n5843) );
  XOR U9438 ( .A(n5846), .B(n5847), .Z(n5845) );
  XOR U9439 ( .A(DB[2627]), .B(DB[2612]), .Z(n5847) );
  AND U9440 ( .A(n326), .B(n5848), .Z(n5846) );
  XOR U9441 ( .A(n5849), .B(n5850), .Z(n5848) );
  XOR U9442 ( .A(DB[2612]), .B(DB[2597]), .Z(n5850) );
  AND U9443 ( .A(n330), .B(n5851), .Z(n5849) );
  XOR U9444 ( .A(n5852), .B(n5853), .Z(n5851) );
  XOR U9445 ( .A(DB[2597]), .B(DB[2582]), .Z(n5853) );
  AND U9446 ( .A(n334), .B(n5854), .Z(n5852) );
  XOR U9447 ( .A(n5855), .B(n5856), .Z(n5854) );
  XOR U9448 ( .A(DB[2582]), .B(DB[2567]), .Z(n5856) );
  AND U9449 ( .A(n338), .B(n5857), .Z(n5855) );
  XOR U9450 ( .A(n5858), .B(n5859), .Z(n5857) );
  XOR U9451 ( .A(DB[2567]), .B(DB[2552]), .Z(n5859) );
  AND U9452 ( .A(n342), .B(n5860), .Z(n5858) );
  XOR U9453 ( .A(n5861), .B(n5862), .Z(n5860) );
  XOR U9454 ( .A(DB[2552]), .B(DB[2537]), .Z(n5862) );
  AND U9455 ( .A(n346), .B(n5863), .Z(n5861) );
  XOR U9456 ( .A(n5864), .B(n5865), .Z(n5863) );
  XOR U9457 ( .A(DB[2537]), .B(DB[2522]), .Z(n5865) );
  AND U9458 ( .A(n350), .B(n5866), .Z(n5864) );
  XOR U9459 ( .A(n5867), .B(n5868), .Z(n5866) );
  XOR U9460 ( .A(DB[2522]), .B(DB[2507]), .Z(n5868) );
  AND U9461 ( .A(n354), .B(n5869), .Z(n5867) );
  XOR U9462 ( .A(n5870), .B(n5871), .Z(n5869) );
  XOR U9463 ( .A(DB[2507]), .B(DB[2492]), .Z(n5871) );
  AND U9464 ( .A(n358), .B(n5872), .Z(n5870) );
  XOR U9465 ( .A(n5873), .B(n5874), .Z(n5872) );
  XOR U9466 ( .A(DB[2492]), .B(DB[2477]), .Z(n5874) );
  AND U9467 ( .A(n362), .B(n5875), .Z(n5873) );
  XOR U9468 ( .A(n5876), .B(n5877), .Z(n5875) );
  XOR U9469 ( .A(DB[2477]), .B(DB[2462]), .Z(n5877) );
  AND U9470 ( .A(n366), .B(n5878), .Z(n5876) );
  XOR U9471 ( .A(n5879), .B(n5880), .Z(n5878) );
  XOR U9472 ( .A(DB[2462]), .B(DB[2447]), .Z(n5880) );
  AND U9473 ( .A(n370), .B(n5881), .Z(n5879) );
  XOR U9474 ( .A(n5882), .B(n5883), .Z(n5881) );
  XOR U9475 ( .A(DB[2447]), .B(DB[2432]), .Z(n5883) );
  AND U9476 ( .A(n374), .B(n5884), .Z(n5882) );
  XOR U9477 ( .A(n5885), .B(n5886), .Z(n5884) );
  XOR U9478 ( .A(DB[2432]), .B(DB[2417]), .Z(n5886) );
  AND U9479 ( .A(n378), .B(n5887), .Z(n5885) );
  XOR U9480 ( .A(n5888), .B(n5889), .Z(n5887) );
  XOR U9481 ( .A(DB[2417]), .B(DB[2402]), .Z(n5889) );
  AND U9482 ( .A(n382), .B(n5890), .Z(n5888) );
  XOR U9483 ( .A(n5891), .B(n5892), .Z(n5890) );
  XOR U9484 ( .A(DB[2402]), .B(DB[2387]), .Z(n5892) );
  AND U9485 ( .A(n386), .B(n5893), .Z(n5891) );
  XOR U9486 ( .A(n5894), .B(n5895), .Z(n5893) );
  XOR U9487 ( .A(DB[2387]), .B(DB[2372]), .Z(n5895) );
  AND U9488 ( .A(n390), .B(n5896), .Z(n5894) );
  XOR U9489 ( .A(n5897), .B(n5898), .Z(n5896) );
  XOR U9490 ( .A(DB[2372]), .B(DB[2357]), .Z(n5898) );
  AND U9491 ( .A(n394), .B(n5899), .Z(n5897) );
  XOR U9492 ( .A(n5900), .B(n5901), .Z(n5899) );
  XOR U9493 ( .A(DB[2357]), .B(DB[2342]), .Z(n5901) );
  AND U9494 ( .A(n398), .B(n5902), .Z(n5900) );
  XOR U9495 ( .A(n5903), .B(n5904), .Z(n5902) );
  XOR U9496 ( .A(DB[2342]), .B(DB[2327]), .Z(n5904) );
  AND U9497 ( .A(n402), .B(n5905), .Z(n5903) );
  XOR U9498 ( .A(n5906), .B(n5907), .Z(n5905) );
  XOR U9499 ( .A(DB[2327]), .B(DB[2312]), .Z(n5907) );
  AND U9500 ( .A(n406), .B(n5908), .Z(n5906) );
  XOR U9501 ( .A(n5909), .B(n5910), .Z(n5908) );
  XOR U9502 ( .A(DB[2312]), .B(DB[2297]), .Z(n5910) );
  AND U9503 ( .A(n410), .B(n5911), .Z(n5909) );
  XOR U9504 ( .A(n5912), .B(n5913), .Z(n5911) );
  XOR U9505 ( .A(DB[2297]), .B(DB[2282]), .Z(n5913) );
  AND U9506 ( .A(n414), .B(n5914), .Z(n5912) );
  XOR U9507 ( .A(n5915), .B(n5916), .Z(n5914) );
  XOR U9508 ( .A(DB[2282]), .B(DB[2267]), .Z(n5916) );
  AND U9509 ( .A(n418), .B(n5917), .Z(n5915) );
  XOR U9510 ( .A(n5918), .B(n5919), .Z(n5917) );
  XOR U9511 ( .A(DB[2267]), .B(DB[2252]), .Z(n5919) );
  AND U9512 ( .A(n422), .B(n5920), .Z(n5918) );
  XOR U9513 ( .A(n5921), .B(n5922), .Z(n5920) );
  XOR U9514 ( .A(DB[2252]), .B(DB[2237]), .Z(n5922) );
  AND U9515 ( .A(n426), .B(n5923), .Z(n5921) );
  XOR U9516 ( .A(n5924), .B(n5925), .Z(n5923) );
  XOR U9517 ( .A(DB[2237]), .B(DB[2222]), .Z(n5925) );
  AND U9518 ( .A(n430), .B(n5926), .Z(n5924) );
  XOR U9519 ( .A(n5927), .B(n5928), .Z(n5926) );
  XOR U9520 ( .A(DB[2222]), .B(DB[2207]), .Z(n5928) );
  AND U9521 ( .A(n434), .B(n5929), .Z(n5927) );
  XOR U9522 ( .A(n5930), .B(n5931), .Z(n5929) );
  XOR U9523 ( .A(DB[2207]), .B(DB[2192]), .Z(n5931) );
  AND U9524 ( .A(n438), .B(n5932), .Z(n5930) );
  XOR U9525 ( .A(n5933), .B(n5934), .Z(n5932) );
  XOR U9526 ( .A(DB[2192]), .B(DB[2177]), .Z(n5934) );
  AND U9527 ( .A(n442), .B(n5935), .Z(n5933) );
  XOR U9528 ( .A(n5936), .B(n5937), .Z(n5935) );
  XOR U9529 ( .A(DB[2177]), .B(DB[2162]), .Z(n5937) );
  AND U9530 ( .A(n446), .B(n5938), .Z(n5936) );
  XOR U9531 ( .A(n5939), .B(n5940), .Z(n5938) );
  XOR U9532 ( .A(DB[2162]), .B(DB[2147]), .Z(n5940) );
  AND U9533 ( .A(n450), .B(n5941), .Z(n5939) );
  XOR U9534 ( .A(n5942), .B(n5943), .Z(n5941) );
  XOR U9535 ( .A(DB[2147]), .B(DB[2132]), .Z(n5943) );
  AND U9536 ( .A(n454), .B(n5944), .Z(n5942) );
  XOR U9537 ( .A(n5945), .B(n5946), .Z(n5944) );
  XOR U9538 ( .A(DB[2132]), .B(DB[2117]), .Z(n5946) );
  AND U9539 ( .A(n458), .B(n5947), .Z(n5945) );
  XOR U9540 ( .A(n5948), .B(n5949), .Z(n5947) );
  XOR U9541 ( .A(DB[2117]), .B(DB[2102]), .Z(n5949) );
  AND U9542 ( .A(n462), .B(n5950), .Z(n5948) );
  XOR U9543 ( .A(n5951), .B(n5952), .Z(n5950) );
  XOR U9544 ( .A(DB[2102]), .B(DB[2087]), .Z(n5952) );
  AND U9545 ( .A(n466), .B(n5953), .Z(n5951) );
  XOR U9546 ( .A(n5954), .B(n5955), .Z(n5953) );
  XOR U9547 ( .A(DB[2087]), .B(DB[2072]), .Z(n5955) );
  AND U9548 ( .A(n470), .B(n5956), .Z(n5954) );
  XOR U9549 ( .A(n5957), .B(n5958), .Z(n5956) );
  XOR U9550 ( .A(DB[2072]), .B(DB[2057]), .Z(n5958) );
  AND U9551 ( .A(n474), .B(n5959), .Z(n5957) );
  XOR U9552 ( .A(n5960), .B(n5961), .Z(n5959) );
  XOR U9553 ( .A(DB[2057]), .B(DB[2042]), .Z(n5961) );
  AND U9554 ( .A(n478), .B(n5962), .Z(n5960) );
  XOR U9555 ( .A(n5963), .B(n5964), .Z(n5962) );
  XOR U9556 ( .A(DB[2042]), .B(DB[2027]), .Z(n5964) );
  AND U9557 ( .A(n482), .B(n5965), .Z(n5963) );
  XOR U9558 ( .A(n5966), .B(n5967), .Z(n5965) );
  XOR U9559 ( .A(DB[2027]), .B(DB[2012]), .Z(n5967) );
  AND U9560 ( .A(n486), .B(n5968), .Z(n5966) );
  XOR U9561 ( .A(n5969), .B(n5970), .Z(n5968) );
  XOR U9562 ( .A(DB[2012]), .B(DB[1997]), .Z(n5970) );
  AND U9563 ( .A(n490), .B(n5971), .Z(n5969) );
  XOR U9564 ( .A(n5972), .B(n5973), .Z(n5971) );
  XOR U9565 ( .A(DB[1997]), .B(DB[1982]), .Z(n5973) );
  AND U9566 ( .A(n494), .B(n5974), .Z(n5972) );
  XOR U9567 ( .A(n5975), .B(n5976), .Z(n5974) );
  XOR U9568 ( .A(DB[1982]), .B(DB[1967]), .Z(n5976) );
  AND U9569 ( .A(n498), .B(n5977), .Z(n5975) );
  XOR U9570 ( .A(n5978), .B(n5979), .Z(n5977) );
  XOR U9571 ( .A(DB[1967]), .B(DB[1952]), .Z(n5979) );
  AND U9572 ( .A(n502), .B(n5980), .Z(n5978) );
  XOR U9573 ( .A(n5981), .B(n5982), .Z(n5980) );
  XOR U9574 ( .A(DB[1952]), .B(DB[1937]), .Z(n5982) );
  AND U9575 ( .A(n506), .B(n5983), .Z(n5981) );
  XOR U9576 ( .A(n5984), .B(n5985), .Z(n5983) );
  XOR U9577 ( .A(DB[1937]), .B(DB[1922]), .Z(n5985) );
  AND U9578 ( .A(n510), .B(n5986), .Z(n5984) );
  XOR U9579 ( .A(n5987), .B(n5988), .Z(n5986) );
  XOR U9580 ( .A(DB[1922]), .B(DB[1907]), .Z(n5988) );
  AND U9581 ( .A(n514), .B(n5989), .Z(n5987) );
  XOR U9582 ( .A(n5990), .B(n5991), .Z(n5989) );
  XOR U9583 ( .A(DB[1907]), .B(DB[1892]), .Z(n5991) );
  AND U9584 ( .A(n518), .B(n5992), .Z(n5990) );
  XOR U9585 ( .A(n5993), .B(n5994), .Z(n5992) );
  XOR U9586 ( .A(DB[1892]), .B(DB[1877]), .Z(n5994) );
  AND U9587 ( .A(n522), .B(n5995), .Z(n5993) );
  XOR U9588 ( .A(n5996), .B(n5997), .Z(n5995) );
  XOR U9589 ( .A(DB[1877]), .B(DB[1862]), .Z(n5997) );
  AND U9590 ( .A(n526), .B(n5998), .Z(n5996) );
  XOR U9591 ( .A(n5999), .B(n6000), .Z(n5998) );
  XOR U9592 ( .A(DB[1862]), .B(DB[1847]), .Z(n6000) );
  AND U9593 ( .A(n530), .B(n6001), .Z(n5999) );
  XOR U9594 ( .A(n6002), .B(n6003), .Z(n6001) );
  XOR U9595 ( .A(DB[1847]), .B(DB[1832]), .Z(n6003) );
  AND U9596 ( .A(n534), .B(n6004), .Z(n6002) );
  XOR U9597 ( .A(n6005), .B(n6006), .Z(n6004) );
  XOR U9598 ( .A(DB[1832]), .B(DB[1817]), .Z(n6006) );
  AND U9599 ( .A(n538), .B(n6007), .Z(n6005) );
  XOR U9600 ( .A(n6008), .B(n6009), .Z(n6007) );
  XOR U9601 ( .A(DB[1817]), .B(DB[1802]), .Z(n6009) );
  AND U9602 ( .A(n542), .B(n6010), .Z(n6008) );
  XOR U9603 ( .A(n6011), .B(n6012), .Z(n6010) );
  XOR U9604 ( .A(DB[1802]), .B(DB[1787]), .Z(n6012) );
  AND U9605 ( .A(n546), .B(n6013), .Z(n6011) );
  XOR U9606 ( .A(n6014), .B(n6015), .Z(n6013) );
  XOR U9607 ( .A(DB[1787]), .B(DB[1772]), .Z(n6015) );
  AND U9608 ( .A(n550), .B(n6016), .Z(n6014) );
  XOR U9609 ( .A(n6017), .B(n6018), .Z(n6016) );
  XOR U9610 ( .A(DB[1772]), .B(DB[1757]), .Z(n6018) );
  AND U9611 ( .A(n554), .B(n6019), .Z(n6017) );
  XOR U9612 ( .A(n6020), .B(n6021), .Z(n6019) );
  XOR U9613 ( .A(DB[1757]), .B(DB[1742]), .Z(n6021) );
  AND U9614 ( .A(n558), .B(n6022), .Z(n6020) );
  XOR U9615 ( .A(n6023), .B(n6024), .Z(n6022) );
  XOR U9616 ( .A(DB[1742]), .B(DB[1727]), .Z(n6024) );
  AND U9617 ( .A(n562), .B(n6025), .Z(n6023) );
  XOR U9618 ( .A(n6026), .B(n6027), .Z(n6025) );
  XOR U9619 ( .A(DB[1727]), .B(DB[1712]), .Z(n6027) );
  AND U9620 ( .A(n566), .B(n6028), .Z(n6026) );
  XOR U9621 ( .A(n6029), .B(n6030), .Z(n6028) );
  XOR U9622 ( .A(DB[1712]), .B(DB[1697]), .Z(n6030) );
  AND U9623 ( .A(n570), .B(n6031), .Z(n6029) );
  XOR U9624 ( .A(n6032), .B(n6033), .Z(n6031) );
  XOR U9625 ( .A(DB[1697]), .B(DB[1682]), .Z(n6033) );
  AND U9626 ( .A(n574), .B(n6034), .Z(n6032) );
  XOR U9627 ( .A(n6035), .B(n6036), .Z(n6034) );
  XOR U9628 ( .A(DB[1682]), .B(DB[1667]), .Z(n6036) );
  AND U9629 ( .A(n578), .B(n6037), .Z(n6035) );
  XOR U9630 ( .A(n6038), .B(n6039), .Z(n6037) );
  XOR U9631 ( .A(DB[1667]), .B(DB[1652]), .Z(n6039) );
  AND U9632 ( .A(n582), .B(n6040), .Z(n6038) );
  XOR U9633 ( .A(n6041), .B(n6042), .Z(n6040) );
  XOR U9634 ( .A(DB[1652]), .B(DB[1637]), .Z(n6042) );
  AND U9635 ( .A(n586), .B(n6043), .Z(n6041) );
  XOR U9636 ( .A(n6044), .B(n6045), .Z(n6043) );
  XOR U9637 ( .A(DB[1637]), .B(DB[1622]), .Z(n6045) );
  AND U9638 ( .A(n590), .B(n6046), .Z(n6044) );
  XOR U9639 ( .A(n6047), .B(n6048), .Z(n6046) );
  XOR U9640 ( .A(DB[1622]), .B(DB[1607]), .Z(n6048) );
  AND U9641 ( .A(n594), .B(n6049), .Z(n6047) );
  XOR U9642 ( .A(n6050), .B(n6051), .Z(n6049) );
  XOR U9643 ( .A(DB[1607]), .B(DB[1592]), .Z(n6051) );
  AND U9644 ( .A(n598), .B(n6052), .Z(n6050) );
  XOR U9645 ( .A(n6053), .B(n6054), .Z(n6052) );
  XOR U9646 ( .A(DB[1592]), .B(DB[1577]), .Z(n6054) );
  AND U9647 ( .A(n602), .B(n6055), .Z(n6053) );
  XOR U9648 ( .A(n6056), .B(n6057), .Z(n6055) );
  XOR U9649 ( .A(DB[1577]), .B(DB[1562]), .Z(n6057) );
  AND U9650 ( .A(n606), .B(n6058), .Z(n6056) );
  XOR U9651 ( .A(n6059), .B(n6060), .Z(n6058) );
  XOR U9652 ( .A(DB[1562]), .B(DB[1547]), .Z(n6060) );
  AND U9653 ( .A(n610), .B(n6061), .Z(n6059) );
  XOR U9654 ( .A(n6062), .B(n6063), .Z(n6061) );
  XOR U9655 ( .A(DB[1547]), .B(DB[1532]), .Z(n6063) );
  AND U9656 ( .A(n614), .B(n6064), .Z(n6062) );
  XOR U9657 ( .A(n6065), .B(n6066), .Z(n6064) );
  XOR U9658 ( .A(DB[1532]), .B(DB[1517]), .Z(n6066) );
  AND U9659 ( .A(n618), .B(n6067), .Z(n6065) );
  XOR U9660 ( .A(n6068), .B(n6069), .Z(n6067) );
  XOR U9661 ( .A(DB[1517]), .B(DB[1502]), .Z(n6069) );
  AND U9662 ( .A(n622), .B(n6070), .Z(n6068) );
  XOR U9663 ( .A(n6071), .B(n6072), .Z(n6070) );
  XOR U9664 ( .A(DB[1502]), .B(DB[1487]), .Z(n6072) );
  AND U9665 ( .A(n626), .B(n6073), .Z(n6071) );
  XOR U9666 ( .A(n6074), .B(n6075), .Z(n6073) );
  XOR U9667 ( .A(DB[1487]), .B(DB[1472]), .Z(n6075) );
  AND U9668 ( .A(n630), .B(n6076), .Z(n6074) );
  XOR U9669 ( .A(n6077), .B(n6078), .Z(n6076) );
  XOR U9670 ( .A(DB[1472]), .B(DB[1457]), .Z(n6078) );
  AND U9671 ( .A(n634), .B(n6079), .Z(n6077) );
  XOR U9672 ( .A(n6080), .B(n6081), .Z(n6079) );
  XOR U9673 ( .A(DB[1457]), .B(DB[1442]), .Z(n6081) );
  AND U9674 ( .A(n638), .B(n6082), .Z(n6080) );
  XOR U9675 ( .A(n6083), .B(n6084), .Z(n6082) );
  XOR U9676 ( .A(DB[1442]), .B(DB[1427]), .Z(n6084) );
  AND U9677 ( .A(n642), .B(n6085), .Z(n6083) );
  XOR U9678 ( .A(n6086), .B(n6087), .Z(n6085) );
  XOR U9679 ( .A(DB[1427]), .B(DB[1412]), .Z(n6087) );
  AND U9680 ( .A(n646), .B(n6088), .Z(n6086) );
  XOR U9681 ( .A(n6089), .B(n6090), .Z(n6088) );
  XOR U9682 ( .A(DB[1412]), .B(DB[1397]), .Z(n6090) );
  AND U9683 ( .A(n650), .B(n6091), .Z(n6089) );
  XOR U9684 ( .A(n6092), .B(n6093), .Z(n6091) );
  XOR U9685 ( .A(DB[1397]), .B(DB[1382]), .Z(n6093) );
  AND U9686 ( .A(n654), .B(n6094), .Z(n6092) );
  XOR U9687 ( .A(n6095), .B(n6096), .Z(n6094) );
  XOR U9688 ( .A(DB[1382]), .B(DB[1367]), .Z(n6096) );
  AND U9689 ( .A(n658), .B(n6097), .Z(n6095) );
  XOR U9690 ( .A(n6098), .B(n6099), .Z(n6097) );
  XOR U9691 ( .A(DB[1367]), .B(DB[1352]), .Z(n6099) );
  AND U9692 ( .A(n662), .B(n6100), .Z(n6098) );
  XOR U9693 ( .A(n6101), .B(n6102), .Z(n6100) );
  XOR U9694 ( .A(DB[1352]), .B(DB[1337]), .Z(n6102) );
  AND U9695 ( .A(n666), .B(n6103), .Z(n6101) );
  XOR U9696 ( .A(n6104), .B(n6105), .Z(n6103) );
  XOR U9697 ( .A(DB[1337]), .B(DB[1322]), .Z(n6105) );
  AND U9698 ( .A(n670), .B(n6106), .Z(n6104) );
  XOR U9699 ( .A(n6107), .B(n6108), .Z(n6106) );
  XOR U9700 ( .A(DB[1322]), .B(DB[1307]), .Z(n6108) );
  AND U9701 ( .A(n674), .B(n6109), .Z(n6107) );
  XOR U9702 ( .A(n6110), .B(n6111), .Z(n6109) );
  XOR U9703 ( .A(DB[1307]), .B(DB[1292]), .Z(n6111) );
  AND U9704 ( .A(n678), .B(n6112), .Z(n6110) );
  XOR U9705 ( .A(n6113), .B(n6114), .Z(n6112) );
  XOR U9706 ( .A(DB[1292]), .B(DB[1277]), .Z(n6114) );
  AND U9707 ( .A(n682), .B(n6115), .Z(n6113) );
  XOR U9708 ( .A(n6116), .B(n6117), .Z(n6115) );
  XOR U9709 ( .A(DB[1277]), .B(DB[1262]), .Z(n6117) );
  AND U9710 ( .A(n686), .B(n6118), .Z(n6116) );
  XOR U9711 ( .A(n6119), .B(n6120), .Z(n6118) );
  XOR U9712 ( .A(DB[1262]), .B(DB[1247]), .Z(n6120) );
  AND U9713 ( .A(n690), .B(n6121), .Z(n6119) );
  XOR U9714 ( .A(n6122), .B(n6123), .Z(n6121) );
  XOR U9715 ( .A(DB[1247]), .B(DB[1232]), .Z(n6123) );
  AND U9716 ( .A(n694), .B(n6124), .Z(n6122) );
  XOR U9717 ( .A(n6125), .B(n6126), .Z(n6124) );
  XOR U9718 ( .A(DB[1232]), .B(DB[1217]), .Z(n6126) );
  AND U9719 ( .A(n698), .B(n6127), .Z(n6125) );
  XOR U9720 ( .A(n6128), .B(n6129), .Z(n6127) );
  XOR U9721 ( .A(DB[1217]), .B(DB[1202]), .Z(n6129) );
  AND U9722 ( .A(n702), .B(n6130), .Z(n6128) );
  XOR U9723 ( .A(n6131), .B(n6132), .Z(n6130) );
  XOR U9724 ( .A(DB[1202]), .B(DB[1187]), .Z(n6132) );
  AND U9725 ( .A(n706), .B(n6133), .Z(n6131) );
  XOR U9726 ( .A(n6134), .B(n6135), .Z(n6133) );
  XOR U9727 ( .A(DB[1187]), .B(DB[1172]), .Z(n6135) );
  AND U9728 ( .A(n710), .B(n6136), .Z(n6134) );
  XOR U9729 ( .A(n6137), .B(n6138), .Z(n6136) );
  XOR U9730 ( .A(DB[1172]), .B(DB[1157]), .Z(n6138) );
  AND U9731 ( .A(n714), .B(n6139), .Z(n6137) );
  XOR U9732 ( .A(n6140), .B(n6141), .Z(n6139) );
  XOR U9733 ( .A(DB[1157]), .B(DB[1142]), .Z(n6141) );
  AND U9734 ( .A(n718), .B(n6142), .Z(n6140) );
  XOR U9735 ( .A(n6143), .B(n6144), .Z(n6142) );
  XOR U9736 ( .A(DB[1142]), .B(DB[1127]), .Z(n6144) );
  AND U9737 ( .A(n722), .B(n6145), .Z(n6143) );
  XOR U9738 ( .A(n6146), .B(n6147), .Z(n6145) );
  XOR U9739 ( .A(DB[1127]), .B(DB[1112]), .Z(n6147) );
  AND U9740 ( .A(n726), .B(n6148), .Z(n6146) );
  XOR U9741 ( .A(n6149), .B(n6150), .Z(n6148) );
  XOR U9742 ( .A(DB[1112]), .B(DB[1097]), .Z(n6150) );
  AND U9743 ( .A(n730), .B(n6151), .Z(n6149) );
  XOR U9744 ( .A(n6152), .B(n6153), .Z(n6151) );
  XOR U9745 ( .A(DB[1097]), .B(DB[1082]), .Z(n6153) );
  AND U9746 ( .A(n734), .B(n6154), .Z(n6152) );
  XOR U9747 ( .A(n6155), .B(n6156), .Z(n6154) );
  XOR U9748 ( .A(DB[1082]), .B(DB[1067]), .Z(n6156) );
  AND U9749 ( .A(n738), .B(n6157), .Z(n6155) );
  XOR U9750 ( .A(n6158), .B(n6159), .Z(n6157) );
  XOR U9751 ( .A(DB[1067]), .B(DB[1052]), .Z(n6159) );
  AND U9752 ( .A(n742), .B(n6160), .Z(n6158) );
  XOR U9753 ( .A(n6161), .B(n6162), .Z(n6160) );
  XOR U9754 ( .A(DB[1052]), .B(DB[1037]), .Z(n6162) );
  AND U9755 ( .A(n746), .B(n6163), .Z(n6161) );
  XOR U9756 ( .A(n6164), .B(n6165), .Z(n6163) );
  XOR U9757 ( .A(DB[1037]), .B(DB[1022]), .Z(n6165) );
  AND U9758 ( .A(n750), .B(n6166), .Z(n6164) );
  XOR U9759 ( .A(n6167), .B(n6168), .Z(n6166) );
  XOR U9760 ( .A(DB[1022]), .B(DB[1007]), .Z(n6168) );
  AND U9761 ( .A(n754), .B(n6169), .Z(n6167) );
  XOR U9762 ( .A(n6170), .B(n6171), .Z(n6169) );
  XOR U9763 ( .A(DB[992]), .B(DB[1007]), .Z(n6171) );
  AND U9764 ( .A(n758), .B(n6172), .Z(n6170) );
  XOR U9765 ( .A(n6173), .B(n6174), .Z(n6172) );
  XOR U9766 ( .A(DB[992]), .B(DB[977]), .Z(n6174) );
  AND U9767 ( .A(n762), .B(n6175), .Z(n6173) );
  XOR U9768 ( .A(n6176), .B(n6177), .Z(n6175) );
  XOR U9769 ( .A(DB[977]), .B(DB[962]), .Z(n6177) );
  AND U9770 ( .A(n766), .B(n6178), .Z(n6176) );
  XOR U9771 ( .A(n6179), .B(n6180), .Z(n6178) );
  XOR U9772 ( .A(DB[962]), .B(DB[947]), .Z(n6180) );
  AND U9773 ( .A(n770), .B(n6181), .Z(n6179) );
  XOR U9774 ( .A(n6182), .B(n6183), .Z(n6181) );
  XOR U9775 ( .A(DB[947]), .B(DB[932]), .Z(n6183) );
  AND U9776 ( .A(n774), .B(n6184), .Z(n6182) );
  XOR U9777 ( .A(n6185), .B(n6186), .Z(n6184) );
  XOR U9778 ( .A(DB[932]), .B(DB[917]), .Z(n6186) );
  AND U9779 ( .A(n778), .B(n6187), .Z(n6185) );
  XOR U9780 ( .A(n6188), .B(n6189), .Z(n6187) );
  XOR U9781 ( .A(DB[917]), .B(DB[902]), .Z(n6189) );
  AND U9782 ( .A(n782), .B(n6190), .Z(n6188) );
  XOR U9783 ( .A(n6191), .B(n6192), .Z(n6190) );
  XOR U9784 ( .A(DB[902]), .B(DB[887]), .Z(n6192) );
  AND U9785 ( .A(n786), .B(n6193), .Z(n6191) );
  XOR U9786 ( .A(n6194), .B(n6195), .Z(n6193) );
  XOR U9787 ( .A(DB[887]), .B(DB[872]), .Z(n6195) );
  AND U9788 ( .A(n790), .B(n6196), .Z(n6194) );
  XOR U9789 ( .A(n6197), .B(n6198), .Z(n6196) );
  XOR U9790 ( .A(DB[872]), .B(DB[857]), .Z(n6198) );
  AND U9791 ( .A(n794), .B(n6199), .Z(n6197) );
  XOR U9792 ( .A(n6200), .B(n6201), .Z(n6199) );
  XOR U9793 ( .A(DB[857]), .B(DB[842]), .Z(n6201) );
  AND U9794 ( .A(n798), .B(n6202), .Z(n6200) );
  XOR U9795 ( .A(n6203), .B(n6204), .Z(n6202) );
  XOR U9796 ( .A(DB[842]), .B(DB[827]), .Z(n6204) );
  AND U9797 ( .A(n802), .B(n6205), .Z(n6203) );
  XOR U9798 ( .A(n6206), .B(n6207), .Z(n6205) );
  XOR U9799 ( .A(DB[827]), .B(DB[812]), .Z(n6207) );
  AND U9800 ( .A(n806), .B(n6208), .Z(n6206) );
  XOR U9801 ( .A(n6209), .B(n6210), .Z(n6208) );
  XOR U9802 ( .A(DB[812]), .B(DB[797]), .Z(n6210) );
  AND U9803 ( .A(n810), .B(n6211), .Z(n6209) );
  XOR U9804 ( .A(n6212), .B(n6213), .Z(n6211) );
  XOR U9805 ( .A(DB[797]), .B(DB[782]), .Z(n6213) );
  AND U9806 ( .A(n814), .B(n6214), .Z(n6212) );
  XOR U9807 ( .A(n6215), .B(n6216), .Z(n6214) );
  XOR U9808 ( .A(DB[782]), .B(DB[767]), .Z(n6216) );
  AND U9809 ( .A(n818), .B(n6217), .Z(n6215) );
  XOR U9810 ( .A(n6218), .B(n6219), .Z(n6217) );
  XOR U9811 ( .A(DB[767]), .B(DB[752]), .Z(n6219) );
  AND U9812 ( .A(n822), .B(n6220), .Z(n6218) );
  XOR U9813 ( .A(n6221), .B(n6222), .Z(n6220) );
  XOR U9814 ( .A(DB[752]), .B(DB[737]), .Z(n6222) );
  AND U9815 ( .A(n826), .B(n6223), .Z(n6221) );
  XOR U9816 ( .A(n6224), .B(n6225), .Z(n6223) );
  XOR U9817 ( .A(DB[737]), .B(DB[722]), .Z(n6225) );
  AND U9818 ( .A(n830), .B(n6226), .Z(n6224) );
  XOR U9819 ( .A(n6227), .B(n6228), .Z(n6226) );
  XOR U9820 ( .A(DB[722]), .B(DB[707]), .Z(n6228) );
  AND U9821 ( .A(n834), .B(n6229), .Z(n6227) );
  XOR U9822 ( .A(n6230), .B(n6231), .Z(n6229) );
  XOR U9823 ( .A(DB[707]), .B(DB[692]), .Z(n6231) );
  AND U9824 ( .A(n838), .B(n6232), .Z(n6230) );
  XOR U9825 ( .A(n6233), .B(n6234), .Z(n6232) );
  XOR U9826 ( .A(DB[692]), .B(DB[677]), .Z(n6234) );
  AND U9827 ( .A(n842), .B(n6235), .Z(n6233) );
  XOR U9828 ( .A(n6236), .B(n6237), .Z(n6235) );
  XOR U9829 ( .A(DB[677]), .B(DB[662]), .Z(n6237) );
  AND U9830 ( .A(n846), .B(n6238), .Z(n6236) );
  XOR U9831 ( .A(n6239), .B(n6240), .Z(n6238) );
  XOR U9832 ( .A(DB[662]), .B(DB[647]), .Z(n6240) );
  AND U9833 ( .A(n850), .B(n6241), .Z(n6239) );
  XOR U9834 ( .A(n6242), .B(n6243), .Z(n6241) );
  XOR U9835 ( .A(DB[647]), .B(DB[632]), .Z(n6243) );
  AND U9836 ( .A(n854), .B(n6244), .Z(n6242) );
  XOR U9837 ( .A(n6245), .B(n6246), .Z(n6244) );
  XOR U9838 ( .A(DB[632]), .B(DB[617]), .Z(n6246) );
  AND U9839 ( .A(n858), .B(n6247), .Z(n6245) );
  XOR U9840 ( .A(n6248), .B(n6249), .Z(n6247) );
  XOR U9841 ( .A(DB[617]), .B(DB[602]), .Z(n6249) );
  AND U9842 ( .A(n862), .B(n6250), .Z(n6248) );
  XOR U9843 ( .A(n6251), .B(n6252), .Z(n6250) );
  XOR U9844 ( .A(DB[602]), .B(DB[587]), .Z(n6252) );
  AND U9845 ( .A(n866), .B(n6253), .Z(n6251) );
  XOR U9846 ( .A(n6254), .B(n6255), .Z(n6253) );
  XOR U9847 ( .A(DB[587]), .B(DB[572]), .Z(n6255) );
  AND U9848 ( .A(n870), .B(n6256), .Z(n6254) );
  XOR U9849 ( .A(n6257), .B(n6258), .Z(n6256) );
  XOR U9850 ( .A(DB[572]), .B(DB[557]), .Z(n6258) );
  AND U9851 ( .A(n874), .B(n6259), .Z(n6257) );
  XOR U9852 ( .A(n6260), .B(n6261), .Z(n6259) );
  XOR U9853 ( .A(DB[557]), .B(DB[542]), .Z(n6261) );
  AND U9854 ( .A(n878), .B(n6262), .Z(n6260) );
  XOR U9855 ( .A(n6263), .B(n6264), .Z(n6262) );
  XOR U9856 ( .A(DB[542]), .B(DB[527]), .Z(n6264) );
  AND U9857 ( .A(n882), .B(n6265), .Z(n6263) );
  XOR U9858 ( .A(n6266), .B(n6267), .Z(n6265) );
  XOR U9859 ( .A(DB[527]), .B(DB[512]), .Z(n6267) );
  AND U9860 ( .A(n886), .B(n6268), .Z(n6266) );
  XOR U9861 ( .A(n6269), .B(n6270), .Z(n6268) );
  XOR U9862 ( .A(DB[512]), .B(DB[497]), .Z(n6270) );
  AND U9863 ( .A(n890), .B(n6271), .Z(n6269) );
  XOR U9864 ( .A(n6272), .B(n6273), .Z(n6271) );
  XOR U9865 ( .A(DB[497]), .B(DB[482]), .Z(n6273) );
  AND U9866 ( .A(n894), .B(n6274), .Z(n6272) );
  XOR U9867 ( .A(n6275), .B(n6276), .Z(n6274) );
  XOR U9868 ( .A(DB[482]), .B(DB[467]), .Z(n6276) );
  AND U9869 ( .A(n898), .B(n6277), .Z(n6275) );
  XOR U9870 ( .A(n6278), .B(n6279), .Z(n6277) );
  XOR U9871 ( .A(DB[467]), .B(DB[452]), .Z(n6279) );
  AND U9872 ( .A(n902), .B(n6280), .Z(n6278) );
  XOR U9873 ( .A(n6281), .B(n6282), .Z(n6280) );
  XOR U9874 ( .A(DB[452]), .B(DB[437]), .Z(n6282) );
  AND U9875 ( .A(n906), .B(n6283), .Z(n6281) );
  XOR U9876 ( .A(n6284), .B(n6285), .Z(n6283) );
  XOR U9877 ( .A(DB[437]), .B(DB[422]), .Z(n6285) );
  AND U9878 ( .A(n910), .B(n6286), .Z(n6284) );
  XOR U9879 ( .A(n6287), .B(n6288), .Z(n6286) );
  XOR U9880 ( .A(DB[422]), .B(DB[407]), .Z(n6288) );
  AND U9881 ( .A(n914), .B(n6289), .Z(n6287) );
  XOR U9882 ( .A(n6290), .B(n6291), .Z(n6289) );
  XOR U9883 ( .A(DB[407]), .B(DB[392]), .Z(n6291) );
  AND U9884 ( .A(n918), .B(n6292), .Z(n6290) );
  XOR U9885 ( .A(n6293), .B(n6294), .Z(n6292) );
  XOR U9886 ( .A(DB[392]), .B(DB[377]), .Z(n6294) );
  AND U9887 ( .A(n922), .B(n6295), .Z(n6293) );
  XOR U9888 ( .A(n6296), .B(n6297), .Z(n6295) );
  XOR U9889 ( .A(DB[377]), .B(DB[362]), .Z(n6297) );
  AND U9890 ( .A(n926), .B(n6298), .Z(n6296) );
  XOR U9891 ( .A(n6299), .B(n6300), .Z(n6298) );
  XOR U9892 ( .A(DB[362]), .B(DB[347]), .Z(n6300) );
  AND U9893 ( .A(n930), .B(n6301), .Z(n6299) );
  XOR U9894 ( .A(n6302), .B(n6303), .Z(n6301) );
  XOR U9895 ( .A(DB[347]), .B(DB[332]), .Z(n6303) );
  AND U9896 ( .A(n934), .B(n6304), .Z(n6302) );
  XOR U9897 ( .A(n6305), .B(n6306), .Z(n6304) );
  XOR U9898 ( .A(DB[332]), .B(DB[317]), .Z(n6306) );
  AND U9899 ( .A(n938), .B(n6307), .Z(n6305) );
  XOR U9900 ( .A(n6308), .B(n6309), .Z(n6307) );
  XOR U9901 ( .A(DB[317]), .B(DB[302]), .Z(n6309) );
  AND U9902 ( .A(n942), .B(n6310), .Z(n6308) );
  XOR U9903 ( .A(n6311), .B(n6312), .Z(n6310) );
  XOR U9904 ( .A(DB[302]), .B(DB[287]), .Z(n6312) );
  AND U9905 ( .A(n946), .B(n6313), .Z(n6311) );
  XOR U9906 ( .A(n6314), .B(n6315), .Z(n6313) );
  XOR U9907 ( .A(DB[287]), .B(DB[272]), .Z(n6315) );
  AND U9908 ( .A(n950), .B(n6316), .Z(n6314) );
  XOR U9909 ( .A(n6317), .B(n6318), .Z(n6316) );
  XOR U9910 ( .A(DB[272]), .B(DB[257]), .Z(n6318) );
  AND U9911 ( .A(n954), .B(n6319), .Z(n6317) );
  XOR U9912 ( .A(n6320), .B(n6321), .Z(n6319) );
  XOR U9913 ( .A(DB[257]), .B(DB[242]), .Z(n6321) );
  AND U9914 ( .A(n958), .B(n6322), .Z(n6320) );
  XOR U9915 ( .A(n6323), .B(n6324), .Z(n6322) );
  XOR U9916 ( .A(DB[242]), .B(DB[227]), .Z(n6324) );
  AND U9917 ( .A(n962), .B(n6325), .Z(n6323) );
  XOR U9918 ( .A(n6326), .B(n6327), .Z(n6325) );
  XOR U9919 ( .A(DB[227]), .B(DB[212]), .Z(n6327) );
  AND U9920 ( .A(n966), .B(n6328), .Z(n6326) );
  XOR U9921 ( .A(n6329), .B(n6330), .Z(n6328) );
  XOR U9922 ( .A(DB[212]), .B(DB[197]), .Z(n6330) );
  AND U9923 ( .A(n970), .B(n6331), .Z(n6329) );
  XOR U9924 ( .A(n6332), .B(n6333), .Z(n6331) );
  XOR U9925 ( .A(DB[197]), .B(DB[182]), .Z(n6333) );
  AND U9926 ( .A(n974), .B(n6334), .Z(n6332) );
  XOR U9927 ( .A(n6335), .B(n6336), .Z(n6334) );
  XOR U9928 ( .A(DB[182]), .B(DB[167]), .Z(n6336) );
  AND U9929 ( .A(n978), .B(n6337), .Z(n6335) );
  XOR U9930 ( .A(n6338), .B(n6339), .Z(n6337) );
  XOR U9931 ( .A(DB[167]), .B(DB[152]), .Z(n6339) );
  AND U9932 ( .A(n982), .B(n6340), .Z(n6338) );
  XOR U9933 ( .A(n6341), .B(n6342), .Z(n6340) );
  XOR U9934 ( .A(DB[152]), .B(DB[137]), .Z(n6342) );
  AND U9935 ( .A(n986), .B(n6343), .Z(n6341) );
  XOR U9936 ( .A(n6344), .B(n6345), .Z(n6343) );
  XOR U9937 ( .A(DB[137]), .B(DB[122]), .Z(n6345) );
  AND U9938 ( .A(n990), .B(n6346), .Z(n6344) );
  XOR U9939 ( .A(n6347), .B(n6348), .Z(n6346) );
  XOR U9940 ( .A(DB[122]), .B(DB[107]), .Z(n6348) );
  AND U9941 ( .A(n994), .B(n6349), .Z(n6347) );
  XOR U9942 ( .A(n6350), .B(n6351), .Z(n6349) );
  XOR U9943 ( .A(DB[92]), .B(DB[107]), .Z(n6351) );
  AND U9944 ( .A(n998), .B(n6352), .Z(n6350) );
  XOR U9945 ( .A(n6353), .B(n6354), .Z(n6352) );
  XOR U9946 ( .A(DB[92]), .B(DB[77]), .Z(n6354) );
  AND U9947 ( .A(n1002), .B(n6355), .Z(n6353) );
  XOR U9948 ( .A(n6356), .B(n6357), .Z(n6355) );
  XOR U9949 ( .A(DB[77]), .B(DB[62]), .Z(n6357) );
  AND U9950 ( .A(n1006), .B(n6358), .Z(n6356) );
  XOR U9951 ( .A(n6359), .B(n6360), .Z(n6358) );
  XOR U9952 ( .A(DB[62]), .B(DB[47]), .Z(n6360) );
  AND U9953 ( .A(n1010), .B(n6361), .Z(n6359) );
  XOR U9954 ( .A(n6362), .B(n6363), .Z(n6361) );
  XOR U9955 ( .A(DB[47]), .B(DB[32]), .Z(n6363) );
  AND U9956 ( .A(n1014), .B(n6364), .Z(n6362) );
  XOR U9957 ( .A(n6365), .B(n6366), .Z(n6364) );
  XOR U9958 ( .A(DB[32]), .B(DB[17]), .Z(n6366) );
  AND U9959 ( .A(n1018), .B(n6367), .Z(n6365) );
  XOR U9960 ( .A(DB[2]), .B(DB[17]), .Z(n6367) );
  XOR U9961 ( .A(DB[3826]), .B(n6368), .Z(min_val_out[1]) );
  AND U9962 ( .A(n2), .B(n6369), .Z(n6368) );
  XOR U9963 ( .A(n6370), .B(n6371), .Z(n6369) );
  XOR U9964 ( .A(DB[3826]), .B(DB[3811]), .Z(n6371) );
  AND U9965 ( .A(n6), .B(n6372), .Z(n6370) );
  XOR U9966 ( .A(n6373), .B(n6374), .Z(n6372) );
  XOR U9967 ( .A(DB[3811]), .B(DB[3796]), .Z(n6374) );
  AND U9968 ( .A(n10), .B(n6375), .Z(n6373) );
  XOR U9969 ( .A(n6376), .B(n6377), .Z(n6375) );
  XOR U9970 ( .A(DB[3796]), .B(DB[3781]), .Z(n6377) );
  AND U9971 ( .A(n14), .B(n6378), .Z(n6376) );
  XOR U9972 ( .A(n6379), .B(n6380), .Z(n6378) );
  XOR U9973 ( .A(DB[3781]), .B(DB[3766]), .Z(n6380) );
  AND U9974 ( .A(n18), .B(n6381), .Z(n6379) );
  XOR U9975 ( .A(n6382), .B(n6383), .Z(n6381) );
  XOR U9976 ( .A(DB[3766]), .B(DB[3751]), .Z(n6383) );
  AND U9977 ( .A(n22), .B(n6384), .Z(n6382) );
  XOR U9978 ( .A(n6385), .B(n6386), .Z(n6384) );
  XOR U9979 ( .A(DB[3751]), .B(DB[3736]), .Z(n6386) );
  AND U9980 ( .A(n26), .B(n6387), .Z(n6385) );
  XOR U9981 ( .A(n6388), .B(n6389), .Z(n6387) );
  XOR U9982 ( .A(DB[3736]), .B(DB[3721]), .Z(n6389) );
  AND U9983 ( .A(n30), .B(n6390), .Z(n6388) );
  XOR U9984 ( .A(n6391), .B(n6392), .Z(n6390) );
  XOR U9985 ( .A(DB[3721]), .B(DB[3706]), .Z(n6392) );
  AND U9986 ( .A(n34), .B(n6393), .Z(n6391) );
  XOR U9987 ( .A(n6394), .B(n6395), .Z(n6393) );
  XOR U9988 ( .A(DB[3706]), .B(DB[3691]), .Z(n6395) );
  AND U9989 ( .A(n38), .B(n6396), .Z(n6394) );
  XOR U9990 ( .A(n6397), .B(n6398), .Z(n6396) );
  XOR U9991 ( .A(DB[3691]), .B(DB[3676]), .Z(n6398) );
  AND U9992 ( .A(n42), .B(n6399), .Z(n6397) );
  XOR U9993 ( .A(n6400), .B(n6401), .Z(n6399) );
  XOR U9994 ( .A(DB[3676]), .B(DB[3661]), .Z(n6401) );
  AND U9995 ( .A(n46), .B(n6402), .Z(n6400) );
  XOR U9996 ( .A(n6403), .B(n6404), .Z(n6402) );
  XOR U9997 ( .A(DB[3661]), .B(DB[3646]), .Z(n6404) );
  AND U9998 ( .A(n50), .B(n6405), .Z(n6403) );
  XOR U9999 ( .A(n6406), .B(n6407), .Z(n6405) );
  XOR U10000 ( .A(DB[3646]), .B(DB[3631]), .Z(n6407) );
  AND U10001 ( .A(n54), .B(n6408), .Z(n6406) );
  XOR U10002 ( .A(n6409), .B(n6410), .Z(n6408) );
  XOR U10003 ( .A(DB[3631]), .B(DB[3616]), .Z(n6410) );
  AND U10004 ( .A(n58), .B(n6411), .Z(n6409) );
  XOR U10005 ( .A(n6412), .B(n6413), .Z(n6411) );
  XOR U10006 ( .A(DB[3616]), .B(DB[3601]), .Z(n6413) );
  AND U10007 ( .A(n62), .B(n6414), .Z(n6412) );
  XOR U10008 ( .A(n6415), .B(n6416), .Z(n6414) );
  XOR U10009 ( .A(DB[3601]), .B(DB[3586]), .Z(n6416) );
  AND U10010 ( .A(n66), .B(n6417), .Z(n6415) );
  XOR U10011 ( .A(n6418), .B(n6419), .Z(n6417) );
  XOR U10012 ( .A(DB[3586]), .B(DB[3571]), .Z(n6419) );
  AND U10013 ( .A(n70), .B(n6420), .Z(n6418) );
  XOR U10014 ( .A(n6421), .B(n6422), .Z(n6420) );
  XOR U10015 ( .A(DB[3571]), .B(DB[3556]), .Z(n6422) );
  AND U10016 ( .A(n74), .B(n6423), .Z(n6421) );
  XOR U10017 ( .A(n6424), .B(n6425), .Z(n6423) );
  XOR U10018 ( .A(DB[3556]), .B(DB[3541]), .Z(n6425) );
  AND U10019 ( .A(n78), .B(n6426), .Z(n6424) );
  XOR U10020 ( .A(n6427), .B(n6428), .Z(n6426) );
  XOR U10021 ( .A(DB[3541]), .B(DB[3526]), .Z(n6428) );
  AND U10022 ( .A(n82), .B(n6429), .Z(n6427) );
  XOR U10023 ( .A(n6430), .B(n6431), .Z(n6429) );
  XOR U10024 ( .A(DB[3526]), .B(DB[3511]), .Z(n6431) );
  AND U10025 ( .A(n86), .B(n6432), .Z(n6430) );
  XOR U10026 ( .A(n6433), .B(n6434), .Z(n6432) );
  XOR U10027 ( .A(DB[3511]), .B(DB[3496]), .Z(n6434) );
  AND U10028 ( .A(n90), .B(n6435), .Z(n6433) );
  XOR U10029 ( .A(n6436), .B(n6437), .Z(n6435) );
  XOR U10030 ( .A(DB[3496]), .B(DB[3481]), .Z(n6437) );
  AND U10031 ( .A(n94), .B(n6438), .Z(n6436) );
  XOR U10032 ( .A(n6439), .B(n6440), .Z(n6438) );
  XOR U10033 ( .A(DB[3481]), .B(DB[3466]), .Z(n6440) );
  AND U10034 ( .A(n98), .B(n6441), .Z(n6439) );
  XOR U10035 ( .A(n6442), .B(n6443), .Z(n6441) );
  XOR U10036 ( .A(DB[3466]), .B(DB[3451]), .Z(n6443) );
  AND U10037 ( .A(n102), .B(n6444), .Z(n6442) );
  XOR U10038 ( .A(n6445), .B(n6446), .Z(n6444) );
  XOR U10039 ( .A(DB[3451]), .B(DB[3436]), .Z(n6446) );
  AND U10040 ( .A(n106), .B(n6447), .Z(n6445) );
  XOR U10041 ( .A(n6448), .B(n6449), .Z(n6447) );
  XOR U10042 ( .A(DB[3436]), .B(DB[3421]), .Z(n6449) );
  AND U10043 ( .A(n110), .B(n6450), .Z(n6448) );
  XOR U10044 ( .A(n6451), .B(n6452), .Z(n6450) );
  XOR U10045 ( .A(DB[3421]), .B(DB[3406]), .Z(n6452) );
  AND U10046 ( .A(n114), .B(n6453), .Z(n6451) );
  XOR U10047 ( .A(n6454), .B(n6455), .Z(n6453) );
  XOR U10048 ( .A(DB[3406]), .B(DB[3391]), .Z(n6455) );
  AND U10049 ( .A(n118), .B(n6456), .Z(n6454) );
  XOR U10050 ( .A(n6457), .B(n6458), .Z(n6456) );
  XOR U10051 ( .A(DB[3391]), .B(DB[3376]), .Z(n6458) );
  AND U10052 ( .A(n122), .B(n6459), .Z(n6457) );
  XOR U10053 ( .A(n6460), .B(n6461), .Z(n6459) );
  XOR U10054 ( .A(DB[3376]), .B(DB[3361]), .Z(n6461) );
  AND U10055 ( .A(n126), .B(n6462), .Z(n6460) );
  XOR U10056 ( .A(n6463), .B(n6464), .Z(n6462) );
  XOR U10057 ( .A(DB[3361]), .B(DB[3346]), .Z(n6464) );
  AND U10058 ( .A(n130), .B(n6465), .Z(n6463) );
  XOR U10059 ( .A(n6466), .B(n6467), .Z(n6465) );
  XOR U10060 ( .A(DB[3346]), .B(DB[3331]), .Z(n6467) );
  AND U10061 ( .A(n134), .B(n6468), .Z(n6466) );
  XOR U10062 ( .A(n6469), .B(n6470), .Z(n6468) );
  XOR U10063 ( .A(DB[3331]), .B(DB[3316]), .Z(n6470) );
  AND U10064 ( .A(n138), .B(n6471), .Z(n6469) );
  XOR U10065 ( .A(n6472), .B(n6473), .Z(n6471) );
  XOR U10066 ( .A(DB[3316]), .B(DB[3301]), .Z(n6473) );
  AND U10067 ( .A(n142), .B(n6474), .Z(n6472) );
  XOR U10068 ( .A(n6475), .B(n6476), .Z(n6474) );
  XOR U10069 ( .A(DB[3301]), .B(DB[3286]), .Z(n6476) );
  AND U10070 ( .A(n146), .B(n6477), .Z(n6475) );
  XOR U10071 ( .A(n6478), .B(n6479), .Z(n6477) );
  XOR U10072 ( .A(DB[3286]), .B(DB[3271]), .Z(n6479) );
  AND U10073 ( .A(n150), .B(n6480), .Z(n6478) );
  XOR U10074 ( .A(n6481), .B(n6482), .Z(n6480) );
  XOR U10075 ( .A(DB[3271]), .B(DB[3256]), .Z(n6482) );
  AND U10076 ( .A(n154), .B(n6483), .Z(n6481) );
  XOR U10077 ( .A(n6484), .B(n6485), .Z(n6483) );
  XOR U10078 ( .A(DB[3256]), .B(DB[3241]), .Z(n6485) );
  AND U10079 ( .A(n158), .B(n6486), .Z(n6484) );
  XOR U10080 ( .A(n6487), .B(n6488), .Z(n6486) );
  XOR U10081 ( .A(DB[3241]), .B(DB[3226]), .Z(n6488) );
  AND U10082 ( .A(n162), .B(n6489), .Z(n6487) );
  XOR U10083 ( .A(n6490), .B(n6491), .Z(n6489) );
  XOR U10084 ( .A(DB[3226]), .B(DB[3211]), .Z(n6491) );
  AND U10085 ( .A(n166), .B(n6492), .Z(n6490) );
  XOR U10086 ( .A(n6493), .B(n6494), .Z(n6492) );
  XOR U10087 ( .A(DB[3211]), .B(DB[3196]), .Z(n6494) );
  AND U10088 ( .A(n170), .B(n6495), .Z(n6493) );
  XOR U10089 ( .A(n6496), .B(n6497), .Z(n6495) );
  XOR U10090 ( .A(DB[3196]), .B(DB[3181]), .Z(n6497) );
  AND U10091 ( .A(n174), .B(n6498), .Z(n6496) );
  XOR U10092 ( .A(n6499), .B(n6500), .Z(n6498) );
  XOR U10093 ( .A(DB[3181]), .B(DB[3166]), .Z(n6500) );
  AND U10094 ( .A(n178), .B(n6501), .Z(n6499) );
  XOR U10095 ( .A(n6502), .B(n6503), .Z(n6501) );
  XOR U10096 ( .A(DB[3166]), .B(DB[3151]), .Z(n6503) );
  AND U10097 ( .A(n182), .B(n6504), .Z(n6502) );
  XOR U10098 ( .A(n6505), .B(n6506), .Z(n6504) );
  XOR U10099 ( .A(DB[3151]), .B(DB[3136]), .Z(n6506) );
  AND U10100 ( .A(n186), .B(n6507), .Z(n6505) );
  XOR U10101 ( .A(n6508), .B(n6509), .Z(n6507) );
  XOR U10102 ( .A(DB[3136]), .B(DB[3121]), .Z(n6509) );
  AND U10103 ( .A(n190), .B(n6510), .Z(n6508) );
  XOR U10104 ( .A(n6511), .B(n6512), .Z(n6510) );
  XOR U10105 ( .A(DB[3121]), .B(DB[3106]), .Z(n6512) );
  AND U10106 ( .A(n194), .B(n6513), .Z(n6511) );
  XOR U10107 ( .A(n6514), .B(n6515), .Z(n6513) );
  XOR U10108 ( .A(DB[3106]), .B(DB[3091]), .Z(n6515) );
  AND U10109 ( .A(n198), .B(n6516), .Z(n6514) );
  XOR U10110 ( .A(n6517), .B(n6518), .Z(n6516) );
  XOR U10111 ( .A(DB[3091]), .B(DB[3076]), .Z(n6518) );
  AND U10112 ( .A(n202), .B(n6519), .Z(n6517) );
  XOR U10113 ( .A(n6520), .B(n6521), .Z(n6519) );
  XOR U10114 ( .A(DB[3076]), .B(DB[3061]), .Z(n6521) );
  AND U10115 ( .A(n206), .B(n6522), .Z(n6520) );
  XOR U10116 ( .A(n6523), .B(n6524), .Z(n6522) );
  XOR U10117 ( .A(DB[3061]), .B(DB[3046]), .Z(n6524) );
  AND U10118 ( .A(n210), .B(n6525), .Z(n6523) );
  XOR U10119 ( .A(n6526), .B(n6527), .Z(n6525) );
  XOR U10120 ( .A(DB[3046]), .B(DB[3031]), .Z(n6527) );
  AND U10121 ( .A(n214), .B(n6528), .Z(n6526) );
  XOR U10122 ( .A(n6529), .B(n6530), .Z(n6528) );
  XOR U10123 ( .A(DB[3031]), .B(DB[3016]), .Z(n6530) );
  AND U10124 ( .A(n218), .B(n6531), .Z(n6529) );
  XOR U10125 ( .A(n6532), .B(n6533), .Z(n6531) );
  XOR U10126 ( .A(DB[3016]), .B(DB[3001]), .Z(n6533) );
  AND U10127 ( .A(n222), .B(n6534), .Z(n6532) );
  XOR U10128 ( .A(n6535), .B(n6536), .Z(n6534) );
  XOR U10129 ( .A(DB[3001]), .B(DB[2986]), .Z(n6536) );
  AND U10130 ( .A(n226), .B(n6537), .Z(n6535) );
  XOR U10131 ( .A(n6538), .B(n6539), .Z(n6537) );
  XOR U10132 ( .A(DB[2986]), .B(DB[2971]), .Z(n6539) );
  AND U10133 ( .A(n230), .B(n6540), .Z(n6538) );
  XOR U10134 ( .A(n6541), .B(n6542), .Z(n6540) );
  XOR U10135 ( .A(DB[2971]), .B(DB[2956]), .Z(n6542) );
  AND U10136 ( .A(n234), .B(n6543), .Z(n6541) );
  XOR U10137 ( .A(n6544), .B(n6545), .Z(n6543) );
  XOR U10138 ( .A(DB[2956]), .B(DB[2941]), .Z(n6545) );
  AND U10139 ( .A(n238), .B(n6546), .Z(n6544) );
  XOR U10140 ( .A(n6547), .B(n6548), .Z(n6546) );
  XOR U10141 ( .A(DB[2941]), .B(DB[2926]), .Z(n6548) );
  AND U10142 ( .A(n242), .B(n6549), .Z(n6547) );
  XOR U10143 ( .A(n6550), .B(n6551), .Z(n6549) );
  XOR U10144 ( .A(DB[2926]), .B(DB[2911]), .Z(n6551) );
  AND U10145 ( .A(n246), .B(n6552), .Z(n6550) );
  XOR U10146 ( .A(n6553), .B(n6554), .Z(n6552) );
  XOR U10147 ( .A(DB[2911]), .B(DB[2896]), .Z(n6554) );
  AND U10148 ( .A(n250), .B(n6555), .Z(n6553) );
  XOR U10149 ( .A(n6556), .B(n6557), .Z(n6555) );
  XOR U10150 ( .A(DB[2896]), .B(DB[2881]), .Z(n6557) );
  AND U10151 ( .A(n254), .B(n6558), .Z(n6556) );
  XOR U10152 ( .A(n6559), .B(n6560), .Z(n6558) );
  XOR U10153 ( .A(DB[2881]), .B(DB[2866]), .Z(n6560) );
  AND U10154 ( .A(n258), .B(n6561), .Z(n6559) );
  XOR U10155 ( .A(n6562), .B(n6563), .Z(n6561) );
  XOR U10156 ( .A(DB[2866]), .B(DB[2851]), .Z(n6563) );
  AND U10157 ( .A(n262), .B(n6564), .Z(n6562) );
  XOR U10158 ( .A(n6565), .B(n6566), .Z(n6564) );
  XOR U10159 ( .A(DB[2851]), .B(DB[2836]), .Z(n6566) );
  AND U10160 ( .A(n266), .B(n6567), .Z(n6565) );
  XOR U10161 ( .A(n6568), .B(n6569), .Z(n6567) );
  XOR U10162 ( .A(DB[2836]), .B(DB[2821]), .Z(n6569) );
  AND U10163 ( .A(n270), .B(n6570), .Z(n6568) );
  XOR U10164 ( .A(n6571), .B(n6572), .Z(n6570) );
  XOR U10165 ( .A(DB[2821]), .B(DB[2806]), .Z(n6572) );
  AND U10166 ( .A(n274), .B(n6573), .Z(n6571) );
  XOR U10167 ( .A(n6574), .B(n6575), .Z(n6573) );
  XOR U10168 ( .A(DB[2806]), .B(DB[2791]), .Z(n6575) );
  AND U10169 ( .A(n278), .B(n6576), .Z(n6574) );
  XOR U10170 ( .A(n6577), .B(n6578), .Z(n6576) );
  XOR U10171 ( .A(DB[2791]), .B(DB[2776]), .Z(n6578) );
  AND U10172 ( .A(n282), .B(n6579), .Z(n6577) );
  XOR U10173 ( .A(n6580), .B(n6581), .Z(n6579) );
  XOR U10174 ( .A(DB[2776]), .B(DB[2761]), .Z(n6581) );
  AND U10175 ( .A(n286), .B(n6582), .Z(n6580) );
  XOR U10176 ( .A(n6583), .B(n6584), .Z(n6582) );
  XOR U10177 ( .A(DB[2761]), .B(DB[2746]), .Z(n6584) );
  AND U10178 ( .A(n290), .B(n6585), .Z(n6583) );
  XOR U10179 ( .A(n6586), .B(n6587), .Z(n6585) );
  XOR U10180 ( .A(DB[2746]), .B(DB[2731]), .Z(n6587) );
  AND U10181 ( .A(n294), .B(n6588), .Z(n6586) );
  XOR U10182 ( .A(n6589), .B(n6590), .Z(n6588) );
  XOR U10183 ( .A(DB[2731]), .B(DB[2716]), .Z(n6590) );
  AND U10184 ( .A(n298), .B(n6591), .Z(n6589) );
  XOR U10185 ( .A(n6592), .B(n6593), .Z(n6591) );
  XOR U10186 ( .A(DB[2716]), .B(DB[2701]), .Z(n6593) );
  AND U10187 ( .A(n302), .B(n6594), .Z(n6592) );
  XOR U10188 ( .A(n6595), .B(n6596), .Z(n6594) );
  XOR U10189 ( .A(DB[2701]), .B(DB[2686]), .Z(n6596) );
  AND U10190 ( .A(n306), .B(n6597), .Z(n6595) );
  XOR U10191 ( .A(n6598), .B(n6599), .Z(n6597) );
  XOR U10192 ( .A(DB[2686]), .B(DB[2671]), .Z(n6599) );
  AND U10193 ( .A(n310), .B(n6600), .Z(n6598) );
  XOR U10194 ( .A(n6601), .B(n6602), .Z(n6600) );
  XOR U10195 ( .A(DB[2671]), .B(DB[2656]), .Z(n6602) );
  AND U10196 ( .A(n314), .B(n6603), .Z(n6601) );
  XOR U10197 ( .A(n6604), .B(n6605), .Z(n6603) );
  XOR U10198 ( .A(DB[2656]), .B(DB[2641]), .Z(n6605) );
  AND U10199 ( .A(n318), .B(n6606), .Z(n6604) );
  XOR U10200 ( .A(n6607), .B(n6608), .Z(n6606) );
  XOR U10201 ( .A(DB[2641]), .B(DB[2626]), .Z(n6608) );
  AND U10202 ( .A(n322), .B(n6609), .Z(n6607) );
  XOR U10203 ( .A(n6610), .B(n6611), .Z(n6609) );
  XOR U10204 ( .A(DB[2626]), .B(DB[2611]), .Z(n6611) );
  AND U10205 ( .A(n326), .B(n6612), .Z(n6610) );
  XOR U10206 ( .A(n6613), .B(n6614), .Z(n6612) );
  XOR U10207 ( .A(DB[2611]), .B(DB[2596]), .Z(n6614) );
  AND U10208 ( .A(n330), .B(n6615), .Z(n6613) );
  XOR U10209 ( .A(n6616), .B(n6617), .Z(n6615) );
  XOR U10210 ( .A(DB[2596]), .B(DB[2581]), .Z(n6617) );
  AND U10211 ( .A(n334), .B(n6618), .Z(n6616) );
  XOR U10212 ( .A(n6619), .B(n6620), .Z(n6618) );
  XOR U10213 ( .A(DB[2581]), .B(DB[2566]), .Z(n6620) );
  AND U10214 ( .A(n338), .B(n6621), .Z(n6619) );
  XOR U10215 ( .A(n6622), .B(n6623), .Z(n6621) );
  XOR U10216 ( .A(DB[2566]), .B(DB[2551]), .Z(n6623) );
  AND U10217 ( .A(n342), .B(n6624), .Z(n6622) );
  XOR U10218 ( .A(n6625), .B(n6626), .Z(n6624) );
  XOR U10219 ( .A(DB[2551]), .B(DB[2536]), .Z(n6626) );
  AND U10220 ( .A(n346), .B(n6627), .Z(n6625) );
  XOR U10221 ( .A(n6628), .B(n6629), .Z(n6627) );
  XOR U10222 ( .A(DB[2536]), .B(DB[2521]), .Z(n6629) );
  AND U10223 ( .A(n350), .B(n6630), .Z(n6628) );
  XOR U10224 ( .A(n6631), .B(n6632), .Z(n6630) );
  XOR U10225 ( .A(DB[2521]), .B(DB[2506]), .Z(n6632) );
  AND U10226 ( .A(n354), .B(n6633), .Z(n6631) );
  XOR U10227 ( .A(n6634), .B(n6635), .Z(n6633) );
  XOR U10228 ( .A(DB[2506]), .B(DB[2491]), .Z(n6635) );
  AND U10229 ( .A(n358), .B(n6636), .Z(n6634) );
  XOR U10230 ( .A(n6637), .B(n6638), .Z(n6636) );
  XOR U10231 ( .A(DB[2491]), .B(DB[2476]), .Z(n6638) );
  AND U10232 ( .A(n362), .B(n6639), .Z(n6637) );
  XOR U10233 ( .A(n6640), .B(n6641), .Z(n6639) );
  XOR U10234 ( .A(DB[2476]), .B(DB[2461]), .Z(n6641) );
  AND U10235 ( .A(n366), .B(n6642), .Z(n6640) );
  XOR U10236 ( .A(n6643), .B(n6644), .Z(n6642) );
  XOR U10237 ( .A(DB[2461]), .B(DB[2446]), .Z(n6644) );
  AND U10238 ( .A(n370), .B(n6645), .Z(n6643) );
  XOR U10239 ( .A(n6646), .B(n6647), .Z(n6645) );
  XOR U10240 ( .A(DB[2446]), .B(DB[2431]), .Z(n6647) );
  AND U10241 ( .A(n374), .B(n6648), .Z(n6646) );
  XOR U10242 ( .A(n6649), .B(n6650), .Z(n6648) );
  XOR U10243 ( .A(DB[2431]), .B(DB[2416]), .Z(n6650) );
  AND U10244 ( .A(n378), .B(n6651), .Z(n6649) );
  XOR U10245 ( .A(n6652), .B(n6653), .Z(n6651) );
  XOR U10246 ( .A(DB[2416]), .B(DB[2401]), .Z(n6653) );
  AND U10247 ( .A(n382), .B(n6654), .Z(n6652) );
  XOR U10248 ( .A(n6655), .B(n6656), .Z(n6654) );
  XOR U10249 ( .A(DB[2401]), .B(DB[2386]), .Z(n6656) );
  AND U10250 ( .A(n386), .B(n6657), .Z(n6655) );
  XOR U10251 ( .A(n6658), .B(n6659), .Z(n6657) );
  XOR U10252 ( .A(DB[2386]), .B(DB[2371]), .Z(n6659) );
  AND U10253 ( .A(n390), .B(n6660), .Z(n6658) );
  XOR U10254 ( .A(n6661), .B(n6662), .Z(n6660) );
  XOR U10255 ( .A(DB[2371]), .B(DB[2356]), .Z(n6662) );
  AND U10256 ( .A(n394), .B(n6663), .Z(n6661) );
  XOR U10257 ( .A(n6664), .B(n6665), .Z(n6663) );
  XOR U10258 ( .A(DB[2356]), .B(DB[2341]), .Z(n6665) );
  AND U10259 ( .A(n398), .B(n6666), .Z(n6664) );
  XOR U10260 ( .A(n6667), .B(n6668), .Z(n6666) );
  XOR U10261 ( .A(DB[2341]), .B(DB[2326]), .Z(n6668) );
  AND U10262 ( .A(n402), .B(n6669), .Z(n6667) );
  XOR U10263 ( .A(n6670), .B(n6671), .Z(n6669) );
  XOR U10264 ( .A(DB[2326]), .B(DB[2311]), .Z(n6671) );
  AND U10265 ( .A(n406), .B(n6672), .Z(n6670) );
  XOR U10266 ( .A(n6673), .B(n6674), .Z(n6672) );
  XOR U10267 ( .A(DB[2311]), .B(DB[2296]), .Z(n6674) );
  AND U10268 ( .A(n410), .B(n6675), .Z(n6673) );
  XOR U10269 ( .A(n6676), .B(n6677), .Z(n6675) );
  XOR U10270 ( .A(DB[2296]), .B(DB[2281]), .Z(n6677) );
  AND U10271 ( .A(n414), .B(n6678), .Z(n6676) );
  XOR U10272 ( .A(n6679), .B(n6680), .Z(n6678) );
  XOR U10273 ( .A(DB[2281]), .B(DB[2266]), .Z(n6680) );
  AND U10274 ( .A(n418), .B(n6681), .Z(n6679) );
  XOR U10275 ( .A(n6682), .B(n6683), .Z(n6681) );
  XOR U10276 ( .A(DB[2266]), .B(DB[2251]), .Z(n6683) );
  AND U10277 ( .A(n422), .B(n6684), .Z(n6682) );
  XOR U10278 ( .A(n6685), .B(n6686), .Z(n6684) );
  XOR U10279 ( .A(DB[2251]), .B(DB[2236]), .Z(n6686) );
  AND U10280 ( .A(n426), .B(n6687), .Z(n6685) );
  XOR U10281 ( .A(n6688), .B(n6689), .Z(n6687) );
  XOR U10282 ( .A(DB[2236]), .B(DB[2221]), .Z(n6689) );
  AND U10283 ( .A(n430), .B(n6690), .Z(n6688) );
  XOR U10284 ( .A(n6691), .B(n6692), .Z(n6690) );
  XOR U10285 ( .A(DB[2221]), .B(DB[2206]), .Z(n6692) );
  AND U10286 ( .A(n434), .B(n6693), .Z(n6691) );
  XOR U10287 ( .A(n6694), .B(n6695), .Z(n6693) );
  XOR U10288 ( .A(DB[2206]), .B(DB[2191]), .Z(n6695) );
  AND U10289 ( .A(n438), .B(n6696), .Z(n6694) );
  XOR U10290 ( .A(n6697), .B(n6698), .Z(n6696) );
  XOR U10291 ( .A(DB[2191]), .B(DB[2176]), .Z(n6698) );
  AND U10292 ( .A(n442), .B(n6699), .Z(n6697) );
  XOR U10293 ( .A(n6700), .B(n6701), .Z(n6699) );
  XOR U10294 ( .A(DB[2176]), .B(DB[2161]), .Z(n6701) );
  AND U10295 ( .A(n446), .B(n6702), .Z(n6700) );
  XOR U10296 ( .A(n6703), .B(n6704), .Z(n6702) );
  XOR U10297 ( .A(DB[2161]), .B(DB[2146]), .Z(n6704) );
  AND U10298 ( .A(n450), .B(n6705), .Z(n6703) );
  XOR U10299 ( .A(n6706), .B(n6707), .Z(n6705) );
  XOR U10300 ( .A(DB[2146]), .B(DB[2131]), .Z(n6707) );
  AND U10301 ( .A(n454), .B(n6708), .Z(n6706) );
  XOR U10302 ( .A(n6709), .B(n6710), .Z(n6708) );
  XOR U10303 ( .A(DB[2131]), .B(DB[2116]), .Z(n6710) );
  AND U10304 ( .A(n458), .B(n6711), .Z(n6709) );
  XOR U10305 ( .A(n6712), .B(n6713), .Z(n6711) );
  XOR U10306 ( .A(DB[2116]), .B(DB[2101]), .Z(n6713) );
  AND U10307 ( .A(n462), .B(n6714), .Z(n6712) );
  XOR U10308 ( .A(n6715), .B(n6716), .Z(n6714) );
  XOR U10309 ( .A(DB[2101]), .B(DB[2086]), .Z(n6716) );
  AND U10310 ( .A(n466), .B(n6717), .Z(n6715) );
  XOR U10311 ( .A(n6718), .B(n6719), .Z(n6717) );
  XOR U10312 ( .A(DB[2086]), .B(DB[2071]), .Z(n6719) );
  AND U10313 ( .A(n470), .B(n6720), .Z(n6718) );
  XOR U10314 ( .A(n6721), .B(n6722), .Z(n6720) );
  XOR U10315 ( .A(DB[2071]), .B(DB[2056]), .Z(n6722) );
  AND U10316 ( .A(n474), .B(n6723), .Z(n6721) );
  XOR U10317 ( .A(n6724), .B(n6725), .Z(n6723) );
  XOR U10318 ( .A(DB[2056]), .B(DB[2041]), .Z(n6725) );
  AND U10319 ( .A(n478), .B(n6726), .Z(n6724) );
  XOR U10320 ( .A(n6727), .B(n6728), .Z(n6726) );
  XOR U10321 ( .A(DB[2041]), .B(DB[2026]), .Z(n6728) );
  AND U10322 ( .A(n482), .B(n6729), .Z(n6727) );
  XOR U10323 ( .A(n6730), .B(n6731), .Z(n6729) );
  XOR U10324 ( .A(DB[2026]), .B(DB[2011]), .Z(n6731) );
  AND U10325 ( .A(n486), .B(n6732), .Z(n6730) );
  XOR U10326 ( .A(n6733), .B(n6734), .Z(n6732) );
  XOR U10327 ( .A(DB[2011]), .B(DB[1996]), .Z(n6734) );
  AND U10328 ( .A(n490), .B(n6735), .Z(n6733) );
  XOR U10329 ( .A(n6736), .B(n6737), .Z(n6735) );
  XOR U10330 ( .A(DB[1996]), .B(DB[1981]), .Z(n6737) );
  AND U10331 ( .A(n494), .B(n6738), .Z(n6736) );
  XOR U10332 ( .A(n6739), .B(n6740), .Z(n6738) );
  XOR U10333 ( .A(DB[1981]), .B(DB[1966]), .Z(n6740) );
  AND U10334 ( .A(n498), .B(n6741), .Z(n6739) );
  XOR U10335 ( .A(n6742), .B(n6743), .Z(n6741) );
  XOR U10336 ( .A(DB[1966]), .B(DB[1951]), .Z(n6743) );
  AND U10337 ( .A(n502), .B(n6744), .Z(n6742) );
  XOR U10338 ( .A(n6745), .B(n6746), .Z(n6744) );
  XOR U10339 ( .A(DB[1951]), .B(DB[1936]), .Z(n6746) );
  AND U10340 ( .A(n506), .B(n6747), .Z(n6745) );
  XOR U10341 ( .A(n6748), .B(n6749), .Z(n6747) );
  XOR U10342 ( .A(DB[1936]), .B(DB[1921]), .Z(n6749) );
  AND U10343 ( .A(n510), .B(n6750), .Z(n6748) );
  XOR U10344 ( .A(n6751), .B(n6752), .Z(n6750) );
  XOR U10345 ( .A(DB[1921]), .B(DB[1906]), .Z(n6752) );
  AND U10346 ( .A(n514), .B(n6753), .Z(n6751) );
  XOR U10347 ( .A(n6754), .B(n6755), .Z(n6753) );
  XOR U10348 ( .A(DB[1906]), .B(DB[1891]), .Z(n6755) );
  AND U10349 ( .A(n518), .B(n6756), .Z(n6754) );
  XOR U10350 ( .A(n6757), .B(n6758), .Z(n6756) );
  XOR U10351 ( .A(DB[1891]), .B(DB[1876]), .Z(n6758) );
  AND U10352 ( .A(n522), .B(n6759), .Z(n6757) );
  XOR U10353 ( .A(n6760), .B(n6761), .Z(n6759) );
  XOR U10354 ( .A(DB[1876]), .B(DB[1861]), .Z(n6761) );
  AND U10355 ( .A(n526), .B(n6762), .Z(n6760) );
  XOR U10356 ( .A(n6763), .B(n6764), .Z(n6762) );
  XOR U10357 ( .A(DB[1861]), .B(DB[1846]), .Z(n6764) );
  AND U10358 ( .A(n530), .B(n6765), .Z(n6763) );
  XOR U10359 ( .A(n6766), .B(n6767), .Z(n6765) );
  XOR U10360 ( .A(DB[1846]), .B(DB[1831]), .Z(n6767) );
  AND U10361 ( .A(n534), .B(n6768), .Z(n6766) );
  XOR U10362 ( .A(n6769), .B(n6770), .Z(n6768) );
  XOR U10363 ( .A(DB[1831]), .B(DB[1816]), .Z(n6770) );
  AND U10364 ( .A(n538), .B(n6771), .Z(n6769) );
  XOR U10365 ( .A(n6772), .B(n6773), .Z(n6771) );
  XOR U10366 ( .A(DB[1816]), .B(DB[1801]), .Z(n6773) );
  AND U10367 ( .A(n542), .B(n6774), .Z(n6772) );
  XOR U10368 ( .A(n6775), .B(n6776), .Z(n6774) );
  XOR U10369 ( .A(DB[1801]), .B(DB[1786]), .Z(n6776) );
  AND U10370 ( .A(n546), .B(n6777), .Z(n6775) );
  XOR U10371 ( .A(n6778), .B(n6779), .Z(n6777) );
  XOR U10372 ( .A(DB[1786]), .B(DB[1771]), .Z(n6779) );
  AND U10373 ( .A(n550), .B(n6780), .Z(n6778) );
  XOR U10374 ( .A(n6781), .B(n6782), .Z(n6780) );
  XOR U10375 ( .A(DB[1771]), .B(DB[1756]), .Z(n6782) );
  AND U10376 ( .A(n554), .B(n6783), .Z(n6781) );
  XOR U10377 ( .A(n6784), .B(n6785), .Z(n6783) );
  XOR U10378 ( .A(DB[1756]), .B(DB[1741]), .Z(n6785) );
  AND U10379 ( .A(n558), .B(n6786), .Z(n6784) );
  XOR U10380 ( .A(n6787), .B(n6788), .Z(n6786) );
  XOR U10381 ( .A(DB[1741]), .B(DB[1726]), .Z(n6788) );
  AND U10382 ( .A(n562), .B(n6789), .Z(n6787) );
  XOR U10383 ( .A(n6790), .B(n6791), .Z(n6789) );
  XOR U10384 ( .A(DB[1726]), .B(DB[1711]), .Z(n6791) );
  AND U10385 ( .A(n566), .B(n6792), .Z(n6790) );
  XOR U10386 ( .A(n6793), .B(n6794), .Z(n6792) );
  XOR U10387 ( .A(DB[1711]), .B(DB[1696]), .Z(n6794) );
  AND U10388 ( .A(n570), .B(n6795), .Z(n6793) );
  XOR U10389 ( .A(n6796), .B(n6797), .Z(n6795) );
  XOR U10390 ( .A(DB[1696]), .B(DB[1681]), .Z(n6797) );
  AND U10391 ( .A(n574), .B(n6798), .Z(n6796) );
  XOR U10392 ( .A(n6799), .B(n6800), .Z(n6798) );
  XOR U10393 ( .A(DB[1681]), .B(DB[1666]), .Z(n6800) );
  AND U10394 ( .A(n578), .B(n6801), .Z(n6799) );
  XOR U10395 ( .A(n6802), .B(n6803), .Z(n6801) );
  XOR U10396 ( .A(DB[1666]), .B(DB[1651]), .Z(n6803) );
  AND U10397 ( .A(n582), .B(n6804), .Z(n6802) );
  XOR U10398 ( .A(n6805), .B(n6806), .Z(n6804) );
  XOR U10399 ( .A(DB[1651]), .B(DB[1636]), .Z(n6806) );
  AND U10400 ( .A(n586), .B(n6807), .Z(n6805) );
  XOR U10401 ( .A(n6808), .B(n6809), .Z(n6807) );
  XOR U10402 ( .A(DB[1636]), .B(DB[1621]), .Z(n6809) );
  AND U10403 ( .A(n590), .B(n6810), .Z(n6808) );
  XOR U10404 ( .A(n6811), .B(n6812), .Z(n6810) );
  XOR U10405 ( .A(DB[1621]), .B(DB[1606]), .Z(n6812) );
  AND U10406 ( .A(n594), .B(n6813), .Z(n6811) );
  XOR U10407 ( .A(n6814), .B(n6815), .Z(n6813) );
  XOR U10408 ( .A(DB[1606]), .B(DB[1591]), .Z(n6815) );
  AND U10409 ( .A(n598), .B(n6816), .Z(n6814) );
  XOR U10410 ( .A(n6817), .B(n6818), .Z(n6816) );
  XOR U10411 ( .A(DB[1591]), .B(DB[1576]), .Z(n6818) );
  AND U10412 ( .A(n602), .B(n6819), .Z(n6817) );
  XOR U10413 ( .A(n6820), .B(n6821), .Z(n6819) );
  XOR U10414 ( .A(DB[1576]), .B(DB[1561]), .Z(n6821) );
  AND U10415 ( .A(n606), .B(n6822), .Z(n6820) );
  XOR U10416 ( .A(n6823), .B(n6824), .Z(n6822) );
  XOR U10417 ( .A(DB[1561]), .B(DB[1546]), .Z(n6824) );
  AND U10418 ( .A(n610), .B(n6825), .Z(n6823) );
  XOR U10419 ( .A(n6826), .B(n6827), .Z(n6825) );
  XOR U10420 ( .A(DB[1546]), .B(DB[1531]), .Z(n6827) );
  AND U10421 ( .A(n614), .B(n6828), .Z(n6826) );
  XOR U10422 ( .A(n6829), .B(n6830), .Z(n6828) );
  XOR U10423 ( .A(DB[1531]), .B(DB[1516]), .Z(n6830) );
  AND U10424 ( .A(n618), .B(n6831), .Z(n6829) );
  XOR U10425 ( .A(n6832), .B(n6833), .Z(n6831) );
  XOR U10426 ( .A(DB[1516]), .B(DB[1501]), .Z(n6833) );
  AND U10427 ( .A(n622), .B(n6834), .Z(n6832) );
  XOR U10428 ( .A(n6835), .B(n6836), .Z(n6834) );
  XOR U10429 ( .A(DB[1501]), .B(DB[1486]), .Z(n6836) );
  AND U10430 ( .A(n626), .B(n6837), .Z(n6835) );
  XOR U10431 ( .A(n6838), .B(n6839), .Z(n6837) );
  XOR U10432 ( .A(DB[1486]), .B(DB[1471]), .Z(n6839) );
  AND U10433 ( .A(n630), .B(n6840), .Z(n6838) );
  XOR U10434 ( .A(n6841), .B(n6842), .Z(n6840) );
  XOR U10435 ( .A(DB[1471]), .B(DB[1456]), .Z(n6842) );
  AND U10436 ( .A(n634), .B(n6843), .Z(n6841) );
  XOR U10437 ( .A(n6844), .B(n6845), .Z(n6843) );
  XOR U10438 ( .A(DB[1456]), .B(DB[1441]), .Z(n6845) );
  AND U10439 ( .A(n638), .B(n6846), .Z(n6844) );
  XOR U10440 ( .A(n6847), .B(n6848), .Z(n6846) );
  XOR U10441 ( .A(DB[1441]), .B(DB[1426]), .Z(n6848) );
  AND U10442 ( .A(n642), .B(n6849), .Z(n6847) );
  XOR U10443 ( .A(n6850), .B(n6851), .Z(n6849) );
  XOR U10444 ( .A(DB[1426]), .B(DB[1411]), .Z(n6851) );
  AND U10445 ( .A(n646), .B(n6852), .Z(n6850) );
  XOR U10446 ( .A(n6853), .B(n6854), .Z(n6852) );
  XOR U10447 ( .A(DB[1411]), .B(DB[1396]), .Z(n6854) );
  AND U10448 ( .A(n650), .B(n6855), .Z(n6853) );
  XOR U10449 ( .A(n6856), .B(n6857), .Z(n6855) );
  XOR U10450 ( .A(DB[1396]), .B(DB[1381]), .Z(n6857) );
  AND U10451 ( .A(n654), .B(n6858), .Z(n6856) );
  XOR U10452 ( .A(n6859), .B(n6860), .Z(n6858) );
  XOR U10453 ( .A(DB[1381]), .B(DB[1366]), .Z(n6860) );
  AND U10454 ( .A(n658), .B(n6861), .Z(n6859) );
  XOR U10455 ( .A(n6862), .B(n6863), .Z(n6861) );
  XOR U10456 ( .A(DB[1366]), .B(DB[1351]), .Z(n6863) );
  AND U10457 ( .A(n662), .B(n6864), .Z(n6862) );
  XOR U10458 ( .A(n6865), .B(n6866), .Z(n6864) );
  XOR U10459 ( .A(DB[1351]), .B(DB[1336]), .Z(n6866) );
  AND U10460 ( .A(n666), .B(n6867), .Z(n6865) );
  XOR U10461 ( .A(n6868), .B(n6869), .Z(n6867) );
  XOR U10462 ( .A(DB[1336]), .B(DB[1321]), .Z(n6869) );
  AND U10463 ( .A(n670), .B(n6870), .Z(n6868) );
  XOR U10464 ( .A(n6871), .B(n6872), .Z(n6870) );
  XOR U10465 ( .A(DB[1321]), .B(DB[1306]), .Z(n6872) );
  AND U10466 ( .A(n674), .B(n6873), .Z(n6871) );
  XOR U10467 ( .A(n6874), .B(n6875), .Z(n6873) );
  XOR U10468 ( .A(DB[1306]), .B(DB[1291]), .Z(n6875) );
  AND U10469 ( .A(n678), .B(n6876), .Z(n6874) );
  XOR U10470 ( .A(n6877), .B(n6878), .Z(n6876) );
  XOR U10471 ( .A(DB[1291]), .B(DB[1276]), .Z(n6878) );
  AND U10472 ( .A(n682), .B(n6879), .Z(n6877) );
  XOR U10473 ( .A(n6880), .B(n6881), .Z(n6879) );
  XOR U10474 ( .A(DB[1276]), .B(DB[1261]), .Z(n6881) );
  AND U10475 ( .A(n686), .B(n6882), .Z(n6880) );
  XOR U10476 ( .A(n6883), .B(n6884), .Z(n6882) );
  XOR U10477 ( .A(DB[1261]), .B(DB[1246]), .Z(n6884) );
  AND U10478 ( .A(n690), .B(n6885), .Z(n6883) );
  XOR U10479 ( .A(n6886), .B(n6887), .Z(n6885) );
  XOR U10480 ( .A(DB[1246]), .B(DB[1231]), .Z(n6887) );
  AND U10481 ( .A(n694), .B(n6888), .Z(n6886) );
  XOR U10482 ( .A(n6889), .B(n6890), .Z(n6888) );
  XOR U10483 ( .A(DB[1231]), .B(DB[1216]), .Z(n6890) );
  AND U10484 ( .A(n698), .B(n6891), .Z(n6889) );
  XOR U10485 ( .A(n6892), .B(n6893), .Z(n6891) );
  XOR U10486 ( .A(DB[1216]), .B(DB[1201]), .Z(n6893) );
  AND U10487 ( .A(n702), .B(n6894), .Z(n6892) );
  XOR U10488 ( .A(n6895), .B(n6896), .Z(n6894) );
  XOR U10489 ( .A(DB[1201]), .B(DB[1186]), .Z(n6896) );
  AND U10490 ( .A(n706), .B(n6897), .Z(n6895) );
  XOR U10491 ( .A(n6898), .B(n6899), .Z(n6897) );
  XOR U10492 ( .A(DB[1186]), .B(DB[1171]), .Z(n6899) );
  AND U10493 ( .A(n710), .B(n6900), .Z(n6898) );
  XOR U10494 ( .A(n6901), .B(n6902), .Z(n6900) );
  XOR U10495 ( .A(DB[1171]), .B(DB[1156]), .Z(n6902) );
  AND U10496 ( .A(n714), .B(n6903), .Z(n6901) );
  XOR U10497 ( .A(n6904), .B(n6905), .Z(n6903) );
  XOR U10498 ( .A(DB[1156]), .B(DB[1141]), .Z(n6905) );
  AND U10499 ( .A(n718), .B(n6906), .Z(n6904) );
  XOR U10500 ( .A(n6907), .B(n6908), .Z(n6906) );
  XOR U10501 ( .A(DB[1141]), .B(DB[1126]), .Z(n6908) );
  AND U10502 ( .A(n722), .B(n6909), .Z(n6907) );
  XOR U10503 ( .A(n6910), .B(n6911), .Z(n6909) );
  XOR U10504 ( .A(DB[1126]), .B(DB[1111]), .Z(n6911) );
  AND U10505 ( .A(n726), .B(n6912), .Z(n6910) );
  XOR U10506 ( .A(n6913), .B(n6914), .Z(n6912) );
  XOR U10507 ( .A(DB[1111]), .B(DB[1096]), .Z(n6914) );
  AND U10508 ( .A(n730), .B(n6915), .Z(n6913) );
  XOR U10509 ( .A(n6916), .B(n6917), .Z(n6915) );
  XOR U10510 ( .A(DB[1096]), .B(DB[1081]), .Z(n6917) );
  AND U10511 ( .A(n734), .B(n6918), .Z(n6916) );
  XOR U10512 ( .A(n6919), .B(n6920), .Z(n6918) );
  XOR U10513 ( .A(DB[1081]), .B(DB[1066]), .Z(n6920) );
  AND U10514 ( .A(n738), .B(n6921), .Z(n6919) );
  XOR U10515 ( .A(n6922), .B(n6923), .Z(n6921) );
  XOR U10516 ( .A(DB[1066]), .B(DB[1051]), .Z(n6923) );
  AND U10517 ( .A(n742), .B(n6924), .Z(n6922) );
  XOR U10518 ( .A(n6925), .B(n6926), .Z(n6924) );
  XOR U10519 ( .A(DB[1051]), .B(DB[1036]), .Z(n6926) );
  AND U10520 ( .A(n746), .B(n6927), .Z(n6925) );
  XOR U10521 ( .A(n6928), .B(n6929), .Z(n6927) );
  XOR U10522 ( .A(DB[1036]), .B(DB[1021]), .Z(n6929) );
  AND U10523 ( .A(n750), .B(n6930), .Z(n6928) );
  XOR U10524 ( .A(n6931), .B(n6932), .Z(n6930) );
  XOR U10525 ( .A(DB[1021]), .B(DB[1006]), .Z(n6932) );
  AND U10526 ( .A(n754), .B(n6933), .Z(n6931) );
  XOR U10527 ( .A(n6934), .B(n6935), .Z(n6933) );
  XOR U10528 ( .A(DB[991]), .B(DB[1006]), .Z(n6935) );
  AND U10529 ( .A(n758), .B(n6936), .Z(n6934) );
  XOR U10530 ( .A(n6937), .B(n6938), .Z(n6936) );
  XOR U10531 ( .A(DB[991]), .B(DB[976]), .Z(n6938) );
  AND U10532 ( .A(n762), .B(n6939), .Z(n6937) );
  XOR U10533 ( .A(n6940), .B(n6941), .Z(n6939) );
  XOR U10534 ( .A(DB[976]), .B(DB[961]), .Z(n6941) );
  AND U10535 ( .A(n766), .B(n6942), .Z(n6940) );
  XOR U10536 ( .A(n6943), .B(n6944), .Z(n6942) );
  XOR U10537 ( .A(DB[961]), .B(DB[946]), .Z(n6944) );
  AND U10538 ( .A(n770), .B(n6945), .Z(n6943) );
  XOR U10539 ( .A(n6946), .B(n6947), .Z(n6945) );
  XOR U10540 ( .A(DB[946]), .B(DB[931]), .Z(n6947) );
  AND U10541 ( .A(n774), .B(n6948), .Z(n6946) );
  XOR U10542 ( .A(n6949), .B(n6950), .Z(n6948) );
  XOR U10543 ( .A(DB[931]), .B(DB[916]), .Z(n6950) );
  AND U10544 ( .A(n778), .B(n6951), .Z(n6949) );
  XOR U10545 ( .A(n6952), .B(n6953), .Z(n6951) );
  XOR U10546 ( .A(DB[916]), .B(DB[901]), .Z(n6953) );
  AND U10547 ( .A(n782), .B(n6954), .Z(n6952) );
  XOR U10548 ( .A(n6955), .B(n6956), .Z(n6954) );
  XOR U10549 ( .A(DB[901]), .B(DB[886]), .Z(n6956) );
  AND U10550 ( .A(n786), .B(n6957), .Z(n6955) );
  XOR U10551 ( .A(n6958), .B(n6959), .Z(n6957) );
  XOR U10552 ( .A(DB[886]), .B(DB[871]), .Z(n6959) );
  AND U10553 ( .A(n790), .B(n6960), .Z(n6958) );
  XOR U10554 ( .A(n6961), .B(n6962), .Z(n6960) );
  XOR U10555 ( .A(DB[871]), .B(DB[856]), .Z(n6962) );
  AND U10556 ( .A(n794), .B(n6963), .Z(n6961) );
  XOR U10557 ( .A(n6964), .B(n6965), .Z(n6963) );
  XOR U10558 ( .A(DB[856]), .B(DB[841]), .Z(n6965) );
  AND U10559 ( .A(n798), .B(n6966), .Z(n6964) );
  XOR U10560 ( .A(n6967), .B(n6968), .Z(n6966) );
  XOR U10561 ( .A(DB[841]), .B(DB[826]), .Z(n6968) );
  AND U10562 ( .A(n802), .B(n6969), .Z(n6967) );
  XOR U10563 ( .A(n6970), .B(n6971), .Z(n6969) );
  XOR U10564 ( .A(DB[826]), .B(DB[811]), .Z(n6971) );
  AND U10565 ( .A(n806), .B(n6972), .Z(n6970) );
  XOR U10566 ( .A(n6973), .B(n6974), .Z(n6972) );
  XOR U10567 ( .A(DB[811]), .B(DB[796]), .Z(n6974) );
  AND U10568 ( .A(n810), .B(n6975), .Z(n6973) );
  XOR U10569 ( .A(n6976), .B(n6977), .Z(n6975) );
  XOR U10570 ( .A(DB[796]), .B(DB[781]), .Z(n6977) );
  AND U10571 ( .A(n814), .B(n6978), .Z(n6976) );
  XOR U10572 ( .A(n6979), .B(n6980), .Z(n6978) );
  XOR U10573 ( .A(DB[781]), .B(DB[766]), .Z(n6980) );
  AND U10574 ( .A(n818), .B(n6981), .Z(n6979) );
  XOR U10575 ( .A(n6982), .B(n6983), .Z(n6981) );
  XOR U10576 ( .A(DB[766]), .B(DB[751]), .Z(n6983) );
  AND U10577 ( .A(n822), .B(n6984), .Z(n6982) );
  XOR U10578 ( .A(n6985), .B(n6986), .Z(n6984) );
  XOR U10579 ( .A(DB[751]), .B(DB[736]), .Z(n6986) );
  AND U10580 ( .A(n826), .B(n6987), .Z(n6985) );
  XOR U10581 ( .A(n6988), .B(n6989), .Z(n6987) );
  XOR U10582 ( .A(DB[736]), .B(DB[721]), .Z(n6989) );
  AND U10583 ( .A(n830), .B(n6990), .Z(n6988) );
  XOR U10584 ( .A(n6991), .B(n6992), .Z(n6990) );
  XOR U10585 ( .A(DB[721]), .B(DB[706]), .Z(n6992) );
  AND U10586 ( .A(n834), .B(n6993), .Z(n6991) );
  XOR U10587 ( .A(n6994), .B(n6995), .Z(n6993) );
  XOR U10588 ( .A(DB[706]), .B(DB[691]), .Z(n6995) );
  AND U10589 ( .A(n838), .B(n6996), .Z(n6994) );
  XOR U10590 ( .A(n6997), .B(n6998), .Z(n6996) );
  XOR U10591 ( .A(DB[691]), .B(DB[676]), .Z(n6998) );
  AND U10592 ( .A(n842), .B(n6999), .Z(n6997) );
  XOR U10593 ( .A(n7000), .B(n7001), .Z(n6999) );
  XOR U10594 ( .A(DB[676]), .B(DB[661]), .Z(n7001) );
  AND U10595 ( .A(n846), .B(n7002), .Z(n7000) );
  XOR U10596 ( .A(n7003), .B(n7004), .Z(n7002) );
  XOR U10597 ( .A(DB[661]), .B(DB[646]), .Z(n7004) );
  AND U10598 ( .A(n850), .B(n7005), .Z(n7003) );
  XOR U10599 ( .A(n7006), .B(n7007), .Z(n7005) );
  XOR U10600 ( .A(DB[646]), .B(DB[631]), .Z(n7007) );
  AND U10601 ( .A(n854), .B(n7008), .Z(n7006) );
  XOR U10602 ( .A(n7009), .B(n7010), .Z(n7008) );
  XOR U10603 ( .A(DB[631]), .B(DB[616]), .Z(n7010) );
  AND U10604 ( .A(n858), .B(n7011), .Z(n7009) );
  XOR U10605 ( .A(n7012), .B(n7013), .Z(n7011) );
  XOR U10606 ( .A(DB[616]), .B(DB[601]), .Z(n7013) );
  AND U10607 ( .A(n862), .B(n7014), .Z(n7012) );
  XOR U10608 ( .A(n7015), .B(n7016), .Z(n7014) );
  XOR U10609 ( .A(DB[601]), .B(DB[586]), .Z(n7016) );
  AND U10610 ( .A(n866), .B(n7017), .Z(n7015) );
  XOR U10611 ( .A(n7018), .B(n7019), .Z(n7017) );
  XOR U10612 ( .A(DB[586]), .B(DB[571]), .Z(n7019) );
  AND U10613 ( .A(n870), .B(n7020), .Z(n7018) );
  XOR U10614 ( .A(n7021), .B(n7022), .Z(n7020) );
  XOR U10615 ( .A(DB[571]), .B(DB[556]), .Z(n7022) );
  AND U10616 ( .A(n874), .B(n7023), .Z(n7021) );
  XOR U10617 ( .A(n7024), .B(n7025), .Z(n7023) );
  XOR U10618 ( .A(DB[556]), .B(DB[541]), .Z(n7025) );
  AND U10619 ( .A(n878), .B(n7026), .Z(n7024) );
  XOR U10620 ( .A(n7027), .B(n7028), .Z(n7026) );
  XOR U10621 ( .A(DB[541]), .B(DB[526]), .Z(n7028) );
  AND U10622 ( .A(n882), .B(n7029), .Z(n7027) );
  XOR U10623 ( .A(n7030), .B(n7031), .Z(n7029) );
  XOR U10624 ( .A(DB[526]), .B(DB[511]), .Z(n7031) );
  AND U10625 ( .A(n886), .B(n7032), .Z(n7030) );
  XOR U10626 ( .A(n7033), .B(n7034), .Z(n7032) );
  XOR U10627 ( .A(DB[511]), .B(DB[496]), .Z(n7034) );
  AND U10628 ( .A(n890), .B(n7035), .Z(n7033) );
  XOR U10629 ( .A(n7036), .B(n7037), .Z(n7035) );
  XOR U10630 ( .A(DB[496]), .B(DB[481]), .Z(n7037) );
  AND U10631 ( .A(n894), .B(n7038), .Z(n7036) );
  XOR U10632 ( .A(n7039), .B(n7040), .Z(n7038) );
  XOR U10633 ( .A(DB[481]), .B(DB[466]), .Z(n7040) );
  AND U10634 ( .A(n898), .B(n7041), .Z(n7039) );
  XOR U10635 ( .A(n7042), .B(n7043), .Z(n7041) );
  XOR U10636 ( .A(DB[466]), .B(DB[451]), .Z(n7043) );
  AND U10637 ( .A(n902), .B(n7044), .Z(n7042) );
  XOR U10638 ( .A(n7045), .B(n7046), .Z(n7044) );
  XOR U10639 ( .A(DB[451]), .B(DB[436]), .Z(n7046) );
  AND U10640 ( .A(n906), .B(n7047), .Z(n7045) );
  XOR U10641 ( .A(n7048), .B(n7049), .Z(n7047) );
  XOR U10642 ( .A(DB[436]), .B(DB[421]), .Z(n7049) );
  AND U10643 ( .A(n910), .B(n7050), .Z(n7048) );
  XOR U10644 ( .A(n7051), .B(n7052), .Z(n7050) );
  XOR U10645 ( .A(DB[421]), .B(DB[406]), .Z(n7052) );
  AND U10646 ( .A(n914), .B(n7053), .Z(n7051) );
  XOR U10647 ( .A(n7054), .B(n7055), .Z(n7053) );
  XOR U10648 ( .A(DB[406]), .B(DB[391]), .Z(n7055) );
  AND U10649 ( .A(n918), .B(n7056), .Z(n7054) );
  XOR U10650 ( .A(n7057), .B(n7058), .Z(n7056) );
  XOR U10651 ( .A(DB[391]), .B(DB[376]), .Z(n7058) );
  AND U10652 ( .A(n922), .B(n7059), .Z(n7057) );
  XOR U10653 ( .A(n7060), .B(n7061), .Z(n7059) );
  XOR U10654 ( .A(DB[376]), .B(DB[361]), .Z(n7061) );
  AND U10655 ( .A(n926), .B(n7062), .Z(n7060) );
  XOR U10656 ( .A(n7063), .B(n7064), .Z(n7062) );
  XOR U10657 ( .A(DB[361]), .B(DB[346]), .Z(n7064) );
  AND U10658 ( .A(n930), .B(n7065), .Z(n7063) );
  XOR U10659 ( .A(n7066), .B(n7067), .Z(n7065) );
  XOR U10660 ( .A(DB[346]), .B(DB[331]), .Z(n7067) );
  AND U10661 ( .A(n934), .B(n7068), .Z(n7066) );
  XOR U10662 ( .A(n7069), .B(n7070), .Z(n7068) );
  XOR U10663 ( .A(DB[331]), .B(DB[316]), .Z(n7070) );
  AND U10664 ( .A(n938), .B(n7071), .Z(n7069) );
  XOR U10665 ( .A(n7072), .B(n7073), .Z(n7071) );
  XOR U10666 ( .A(DB[316]), .B(DB[301]), .Z(n7073) );
  AND U10667 ( .A(n942), .B(n7074), .Z(n7072) );
  XOR U10668 ( .A(n7075), .B(n7076), .Z(n7074) );
  XOR U10669 ( .A(DB[301]), .B(DB[286]), .Z(n7076) );
  AND U10670 ( .A(n946), .B(n7077), .Z(n7075) );
  XOR U10671 ( .A(n7078), .B(n7079), .Z(n7077) );
  XOR U10672 ( .A(DB[286]), .B(DB[271]), .Z(n7079) );
  AND U10673 ( .A(n950), .B(n7080), .Z(n7078) );
  XOR U10674 ( .A(n7081), .B(n7082), .Z(n7080) );
  XOR U10675 ( .A(DB[271]), .B(DB[256]), .Z(n7082) );
  AND U10676 ( .A(n954), .B(n7083), .Z(n7081) );
  XOR U10677 ( .A(n7084), .B(n7085), .Z(n7083) );
  XOR U10678 ( .A(DB[256]), .B(DB[241]), .Z(n7085) );
  AND U10679 ( .A(n958), .B(n7086), .Z(n7084) );
  XOR U10680 ( .A(n7087), .B(n7088), .Z(n7086) );
  XOR U10681 ( .A(DB[241]), .B(DB[226]), .Z(n7088) );
  AND U10682 ( .A(n962), .B(n7089), .Z(n7087) );
  XOR U10683 ( .A(n7090), .B(n7091), .Z(n7089) );
  XOR U10684 ( .A(DB[226]), .B(DB[211]), .Z(n7091) );
  AND U10685 ( .A(n966), .B(n7092), .Z(n7090) );
  XOR U10686 ( .A(n7093), .B(n7094), .Z(n7092) );
  XOR U10687 ( .A(DB[211]), .B(DB[196]), .Z(n7094) );
  AND U10688 ( .A(n970), .B(n7095), .Z(n7093) );
  XOR U10689 ( .A(n7096), .B(n7097), .Z(n7095) );
  XOR U10690 ( .A(DB[196]), .B(DB[181]), .Z(n7097) );
  AND U10691 ( .A(n974), .B(n7098), .Z(n7096) );
  XOR U10692 ( .A(n7099), .B(n7100), .Z(n7098) );
  XOR U10693 ( .A(DB[181]), .B(DB[166]), .Z(n7100) );
  AND U10694 ( .A(n978), .B(n7101), .Z(n7099) );
  XOR U10695 ( .A(n7102), .B(n7103), .Z(n7101) );
  XOR U10696 ( .A(DB[166]), .B(DB[151]), .Z(n7103) );
  AND U10697 ( .A(n982), .B(n7104), .Z(n7102) );
  XOR U10698 ( .A(n7105), .B(n7106), .Z(n7104) );
  XOR U10699 ( .A(DB[151]), .B(DB[136]), .Z(n7106) );
  AND U10700 ( .A(n986), .B(n7107), .Z(n7105) );
  XOR U10701 ( .A(n7108), .B(n7109), .Z(n7107) );
  XOR U10702 ( .A(DB[136]), .B(DB[121]), .Z(n7109) );
  AND U10703 ( .A(n990), .B(n7110), .Z(n7108) );
  XOR U10704 ( .A(n7111), .B(n7112), .Z(n7110) );
  XOR U10705 ( .A(DB[121]), .B(DB[106]), .Z(n7112) );
  AND U10706 ( .A(n994), .B(n7113), .Z(n7111) );
  XOR U10707 ( .A(n7114), .B(n7115), .Z(n7113) );
  XOR U10708 ( .A(DB[91]), .B(DB[106]), .Z(n7115) );
  AND U10709 ( .A(n998), .B(n7116), .Z(n7114) );
  XOR U10710 ( .A(n7117), .B(n7118), .Z(n7116) );
  XOR U10711 ( .A(DB[91]), .B(DB[76]), .Z(n7118) );
  AND U10712 ( .A(n1002), .B(n7119), .Z(n7117) );
  XOR U10713 ( .A(n7120), .B(n7121), .Z(n7119) );
  XOR U10714 ( .A(DB[76]), .B(DB[61]), .Z(n7121) );
  AND U10715 ( .A(n1006), .B(n7122), .Z(n7120) );
  XOR U10716 ( .A(n7123), .B(n7124), .Z(n7122) );
  XOR U10717 ( .A(DB[61]), .B(DB[46]), .Z(n7124) );
  AND U10718 ( .A(n1010), .B(n7125), .Z(n7123) );
  XOR U10719 ( .A(n7126), .B(n7127), .Z(n7125) );
  XOR U10720 ( .A(DB[46]), .B(DB[31]), .Z(n7127) );
  AND U10721 ( .A(n1014), .B(n7128), .Z(n7126) );
  XOR U10722 ( .A(n7129), .B(n7130), .Z(n7128) );
  XOR U10723 ( .A(DB[31]), .B(DB[16]), .Z(n7130) );
  AND U10724 ( .A(n1018), .B(n7131), .Z(n7129) );
  XOR U10725 ( .A(DB[1]), .B(DB[16]), .Z(n7131) );
  XOR U10726 ( .A(DB[3839]), .B(n7132), .Z(min_val_out[14]) );
  AND U10727 ( .A(n2), .B(n7133), .Z(n7132) );
  XOR U10728 ( .A(n7134), .B(n7135), .Z(n7133) );
  XOR U10729 ( .A(DB[3839]), .B(DB[3824]), .Z(n7135) );
  AND U10730 ( .A(n6), .B(n7136), .Z(n7134) );
  XOR U10731 ( .A(n7137), .B(n7138), .Z(n7136) );
  XOR U10732 ( .A(DB[3824]), .B(DB[3809]), .Z(n7138) );
  AND U10733 ( .A(n10), .B(n7139), .Z(n7137) );
  XOR U10734 ( .A(n7140), .B(n7141), .Z(n7139) );
  XOR U10735 ( .A(DB[3809]), .B(DB[3794]), .Z(n7141) );
  AND U10736 ( .A(n14), .B(n7142), .Z(n7140) );
  XOR U10737 ( .A(n7143), .B(n7144), .Z(n7142) );
  XOR U10738 ( .A(DB[3794]), .B(DB[3779]), .Z(n7144) );
  AND U10739 ( .A(n18), .B(n7145), .Z(n7143) );
  XOR U10740 ( .A(n7146), .B(n7147), .Z(n7145) );
  XOR U10741 ( .A(DB[3779]), .B(DB[3764]), .Z(n7147) );
  AND U10742 ( .A(n22), .B(n7148), .Z(n7146) );
  XOR U10743 ( .A(n7149), .B(n7150), .Z(n7148) );
  XOR U10744 ( .A(DB[3764]), .B(DB[3749]), .Z(n7150) );
  AND U10745 ( .A(n26), .B(n7151), .Z(n7149) );
  XOR U10746 ( .A(n7152), .B(n7153), .Z(n7151) );
  XOR U10747 ( .A(DB[3749]), .B(DB[3734]), .Z(n7153) );
  AND U10748 ( .A(n30), .B(n7154), .Z(n7152) );
  XOR U10749 ( .A(n7155), .B(n7156), .Z(n7154) );
  XOR U10750 ( .A(DB[3734]), .B(DB[3719]), .Z(n7156) );
  AND U10751 ( .A(n34), .B(n7157), .Z(n7155) );
  XOR U10752 ( .A(n7158), .B(n7159), .Z(n7157) );
  XOR U10753 ( .A(DB[3719]), .B(DB[3704]), .Z(n7159) );
  AND U10754 ( .A(n38), .B(n7160), .Z(n7158) );
  XOR U10755 ( .A(n7161), .B(n7162), .Z(n7160) );
  XOR U10756 ( .A(DB[3704]), .B(DB[3689]), .Z(n7162) );
  AND U10757 ( .A(n42), .B(n7163), .Z(n7161) );
  XOR U10758 ( .A(n7164), .B(n7165), .Z(n7163) );
  XOR U10759 ( .A(DB[3689]), .B(DB[3674]), .Z(n7165) );
  AND U10760 ( .A(n46), .B(n7166), .Z(n7164) );
  XOR U10761 ( .A(n7167), .B(n7168), .Z(n7166) );
  XOR U10762 ( .A(DB[3674]), .B(DB[3659]), .Z(n7168) );
  AND U10763 ( .A(n50), .B(n7169), .Z(n7167) );
  XOR U10764 ( .A(n7170), .B(n7171), .Z(n7169) );
  XOR U10765 ( .A(DB[3659]), .B(DB[3644]), .Z(n7171) );
  AND U10766 ( .A(n54), .B(n7172), .Z(n7170) );
  XOR U10767 ( .A(n7173), .B(n7174), .Z(n7172) );
  XOR U10768 ( .A(DB[3644]), .B(DB[3629]), .Z(n7174) );
  AND U10769 ( .A(n58), .B(n7175), .Z(n7173) );
  XOR U10770 ( .A(n7176), .B(n7177), .Z(n7175) );
  XOR U10771 ( .A(DB[3629]), .B(DB[3614]), .Z(n7177) );
  AND U10772 ( .A(n62), .B(n7178), .Z(n7176) );
  XOR U10773 ( .A(n7179), .B(n7180), .Z(n7178) );
  XOR U10774 ( .A(DB[3614]), .B(DB[3599]), .Z(n7180) );
  AND U10775 ( .A(n66), .B(n7181), .Z(n7179) );
  XOR U10776 ( .A(n7182), .B(n7183), .Z(n7181) );
  XOR U10777 ( .A(DB[3599]), .B(DB[3584]), .Z(n7183) );
  AND U10778 ( .A(n70), .B(n7184), .Z(n7182) );
  XOR U10779 ( .A(n7185), .B(n7186), .Z(n7184) );
  XOR U10780 ( .A(DB[3584]), .B(DB[3569]), .Z(n7186) );
  AND U10781 ( .A(n74), .B(n7187), .Z(n7185) );
  XOR U10782 ( .A(n7188), .B(n7189), .Z(n7187) );
  XOR U10783 ( .A(DB[3569]), .B(DB[3554]), .Z(n7189) );
  AND U10784 ( .A(n78), .B(n7190), .Z(n7188) );
  XOR U10785 ( .A(n7191), .B(n7192), .Z(n7190) );
  XOR U10786 ( .A(DB[3554]), .B(DB[3539]), .Z(n7192) );
  AND U10787 ( .A(n82), .B(n7193), .Z(n7191) );
  XOR U10788 ( .A(n7194), .B(n7195), .Z(n7193) );
  XOR U10789 ( .A(DB[3539]), .B(DB[3524]), .Z(n7195) );
  AND U10790 ( .A(n86), .B(n7196), .Z(n7194) );
  XOR U10791 ( .A(n7197), .B(n7198), .Z(n7196) );
  XOR U10792 ( .A(DB[3524]), .B(DB[3509]), .Z(n7198) );
  AND U10793 ( .A(n90), .B(n7199), .Z(n7197) );
  XOR U10794 ( .A(n7200), .B(n7201), .Z(n7199) );
  XOR U10795 ( .A(DB[3509]), .B(DB[3494]), .Z(n7201) );
  AND U10796 ( .A(n94), .B(n7202), .Z(n7200) );
  XOR U10797 ( .A(n7203), .B(n7204), .Z(n7202) );
  XOR U10798 ( .A(DB[3494]), .B(DB[3479]), .Z(n7204) );
  AND U10799 ( .A(n98), .B(n7205), .Z(n7203) );
  XOR U10800 ( .A(n7206), .B(n7207), .Z(n7205) );
  XOR U10801 ( .A(DB[3479]), .B(DB[3464]), .Z(n7207) );
  AND U10802 ( .A(n102), .B(n7208), .Z(n7206) );
  XOR U10803 ( .A(n7209), .B(n7210), .Z(n7208) );
  XOR U10804 ( .A(DB[3464]), .B(DB[3449]), .Z(n7210) );
  AND U10805 ( .A(n106), .B(n7211), .Z(n7209) );
  XOR U10806 ( .A(n7212), .B(n7213), .Z(n7211) );
  XOR U10807 ( .A(DB[3449]), .B(DB[3434]), .Z(n7213) );
  AND U10808 ( .A(n110), .B(n7214), .Z(n7212) );
  XOR U10809 ( .A(n7215), .B(n7216), .Z(n7214) );
  XOR U10810 ( .A(DB[3434]), .B(DB[3419]), .Z(n7216) );
  AND U10811 ( .A(n114), .B(n7217), .Z(n7215) );
  XOR U10812 ( .A(n7218), .B(n7219), .Z(n7217) );
  XOR U10813 ( .A(DB[3419]), .B(DB[3404]), .Z(n7219) );
  AND U10814 ( .A(n118), .B(n7220), .Z(n7218) );
  XOR U10815 ( .A(n7221), .B(n7222), .Z(n7220) );
  XOR U10816 ( .A(DB[3404]), .B(DB[3389]), .Z(n7222) );
  AND U10817 ( .A(n122), .B(n7223), .Z(n7221) );
  XOR U10818 ( .A(n7224), .B(n7225), .Z(n7223) );
  XOR U10819 ( .A(DB[3389]), .B(DB[3374]), .Z(n7225) );
  AND U10820 ( .A(n126), .B(n7226), .Z(n7224) );
  XOR U10821 ( .A(n7227), .B(n7228), .Z(n7226) );
  XOR U10822 ( .A(DB[3374]), .B(DB[3359]), .Z(n7228) );
  AND U10823 ( .A(n130), .B(n7229), .Z(n7227) );
  XOR U10824 ( .A(n7230), .B(n7231), .Z(n7229) );
  XOR U10825 ( .A(DB[3359]), .B(DB[3344]), .Z(n7231) );
  AND U10826 ( .A(n134), .B(n7232), .Z(n7230) );
  XOR U10827 ( .A(n7233), .B(n7234), .Z(n7232) );
  XOR U10828 ( .A(DB[3344]), .B(DB[3329]), .Z(n7234) );
  AND U10829 ( .A(n138), .B(n7235), .Z(n7233) );
  XOR U10830 ( .A(n7236), .B(n7237), .Z(n7235) );
  XOR U10831 ( .A(DB[3329]), .B(DB[3314]), .Z(n7237) );
  AND U10832 ( .A(n142), .B(n7238), .Z(n7236) );
  XOR U10833 ( .A(n7239), .B(n7240), .Z(n7238) );
  XOR U10834 ( .A(DB[3314]), .B(DB[3299]), .Z(n7240) );
  AND U10835 ( .A(n146), .B(n7241), .Z(n7239) );
  XOR U10836 ( .A(n7242), .B(n7243), .Z(n7241) );
  XOR U10837 ( .A(DB[3299]), .B(DB[3284]), .Z(n7243) );
  AND U10838 ( .A(n150), .B(n7244), .Z(n7242) );
  XOR U10839 ( .A(n7245), .B(n7246), .Z(n7244) );
  XOR U10840 ( .A(DB[3284]), .B(DB[3269]), .Z(n7246) );
  AND U10841 ( .A(n154), .B(n7247), .Z(n7245) );
  XOR U10842 ( .A(n7248), .B(n7249), .Z(n7247) );
  XOR U10843 ( .A(DB[3269]), .B(DB[3254]), .Z(n7249) );
  AND U10844 ( .A(n158), .B(n7250), .Z(n7248) );
  XOR U10845 ( .A(n7251), .B(n7252), .Z(n7250) );
  XOR U10846 ( .A(DB[3254]), .B(DB[3239]), .Z(n7252) );
  AND U10847 ( .A(n162), .B(n7253), .Z(n7251) );
  XOR U10848 ( .A(n7254), .B(n7255), .Z(n7253) );
  XOR U10849 ( .A(DB[3239]), .B(DB[3224]), .Z(n7255) );
  AND U10850 ( .A(n166), .B(n7256), .Z(n7254) );
  XOR U10851 ( .A(n7257), .B(n7258), .Z(n7256) );
  XOR U10852 ( .A(DB[3224]), .B(DB[3209]), .Z(n7258) );
  AND U10853 ( .A(n170), .B(n7259), .Z(n7257) );
  XOR U10854 ( .A(n7260), .B(n7261), .Z(n7259) );
  XOR U10855 ( .A(DB[3209]), .B(DB[3194]), .Z(n7261) );
  AND U10856 ( .A(n174), .B(n7262), .Z(n7260) );
  XOR U10857 ( .A(n7263), .B(n7264), .Z(n7262) );
  XOR U10858 ( .A(DB[3194]), .B(DB[3179]), .Z(n7264) );
  AND U10859 ( .A(n178), .B(n7265), .Z(n7263) );
  XOR U10860 ( .A(n7266), .B(n7267), .Z(n7265) );
  XOR U10861 ( .A(DB[3179]), .B(DB[3164]), .Z(n7267) );
  AND U10862 ( .A(n182), .B(n7268), .Z(n7266) );
  XOR U10863 ( .A(n7269), .B(n7270), .Z(n7268) );
  XOR U10864 ( .A(DB[3164]), .B(DB[3149]), .Z(n7270) );
  AND U10865 ( .A(n186), .B(n7271), .Z(n7269) );
  XOR U10866 ( .A(n7272), .B(n7273), .Z(n7271) );
  XOR U10867 ( .A(DB[3149]), .B(DB[3134]), .Z(n7273) );
  AND U10868 ( .A(n190), .B(n7274), .Z(n7272) );
  XOR U10869 ( .A(n7275), .B(n7276), .Z(n7274) );
  XOR U10870 ( .A(DB[3134]), .B(DB[3119]), .Z(n7276) );
  AND U10871 ( .A(n194), .B(n7277), .Z(n7275) );
  XOR U10872 ( .A(n7278), .B(n7279), .Z(n7277) );
  XOR U10873 ( .A(DB[3119]), .B(DB[3104]), .Z(n7279) );
  AND U10874 ( .A(n198), .B(n7280), .Z(n7278) );
  XOR U10875 ( .A(n7281), .B(n7282), .Z(n7280) );
  XOR U10876 ( .A(DB[3104]), .B(DB[3089]), .Z(n7282) );
  AND U10877 ( .A(n202), .B(n7283), .Z(n7281) );
  XOR U10878 ( .A(n7284), .B(n7285), .Z(n7283) );
  XOR U10879 ( .A(DB[3089]), .B(DB[3074]), .Z(n7285) );
  AND U10880 ( .A(n206), .B(n7286), .Z(n7284) );
  XOR U10881 ( .A(n7287), .B(n7288), .Z(n7286) );
  XOR U10882 ( .A(DB[3074]), .B(DB[3059]), .Z(n7288) );
  AND U10883 ( .A(n210), .B(n7289), .Z(n7287) );
  XOR U10884 ( .A(n7290), .B(n7291), .Z(n7289) );
  XOR U10885 ( .A(DB[3059]), .B(DB[3044]), .Z(n7291) );
  AND U10886 ( .A(n214), .B(n7292), .Z(n7290) );
  XOR U10887 ( .A(n7293), .B(n7294), .Z(n7292) );
  XOR U10888 ( .A(DB[3044]), .B(DB[3029]), .Z(n7294) );
  AND U10889 ( .A(n218), .B(n7295), .Z(n7293) );
  XOR U10890 ( .A(n7296), .B(n7297), .Z(n7295) );
  XOR U10891 ( .A(DB[3029]), .B(DB[3014]), .Z(n7297) );
  AND U10892 ( .A(n222), .B(n7298), .Z(n7296) );
  XOR U10893 ( .A(n7299), .B(n7300), .Z(n7298) );
  XOR U10894 ( .A(DB[3014]), .B(DB[2999]), .Z(n7300) );
  AND U10895 ( .A(n226), .B(n7301), .Z(n7299) );
  XOR U10896 ( .A(n7302), .B(n7303), .Z(n7301) );
  XOR U10897 ( .A(DB[2999]), .B(DB[2984]), .Z(n7303) );
  AND U10898 ( .A(n230), .B(n7304), .Z(n7302) );
  XOR U10899 ( .A(n7305), .B(n7306), .Z(n7304) );
  XOR U10900 ( .A(DB[2984]), .B(DB[2969]), .Z(n7306) );
  AND U10901 ( .A(n234), .B(n7307), .Z(n7305) );
  XOR U10902 ( .A(n7308), .B(n7309), .Z(n7307) );
  XOR U10903 ( .A(DB[2969]), .B(DB[2954]), .Z(n7309) );
  AND U10904 ( .A(n238), .B(n7310), .Z(n7308) );
  XOR U10905 ( .A(n7311), .B(n7312), .Z(n7310) );
  XOR U10906 ( .A(DB[2954]), .B(DB[2939]), .Z(n7312) );
  AND U10907 ( .A(n242), .B(n7313), .Z(n7311) );
  XOR U10908 ( .A(n7314), .B(n7315), .Z(n7313) );
  XOR U10909 ( .A(DB[2939]), .B(DB[2924]), .Z(n7315) );
  AND U10910 ( .A(n246), .B(n7316), .Z(n7314) );
  XOR U10911 ( .A(n7317), .B(n7318), .Z(n7316) );
  XOR U10912 ( .A(DB[2924]), .B(DB[2909]), .Z(n7318) );
  AND U10913 ( .A(n250), .B(n7319), .Z(n7317) );
  XOR U10914 ( .A(n7320), .B(n7321), .Z(n7319) );
  XOR U10915 ( .A(DB[2909]), .B(DB[2894]), .Z(n7321) );
  AND U10916 ( .A(n254), .B(n7322), .Z(n7320) );
  XOR U10917 ( .A(n7323), .B(n7324), .Z(n7322) );
  XOR U10918 ( .A(DB[2894]), .B(DB[2879]), .Z(n7324) );
  AND U10919 ( .A(n258), .B(n7325), .Z(n7323) );
  XOR U10920 ( .A(n7326), .B(n7327), .Z(n7325) );
  XOR U10921 ( .A(DB[2879]), .B(DB[2864]), .Z(n7327) );
  AND U10922 ( .A(n262), .B(n7328), .Z(n7326) );
  XOR U10923 ( .A(n7329), .B(n7330), .Z(n7328) );
  XOR U10924 ( .A(DB[2864]), .B(DB[2849]), .Z(n7330) );
  AND U10925 ( .A(n266), .B(n7331), .Z(n7329) );
  XOR U10926 ( .A(n7332), .B(n7333), .Z(n7331) );
  XOR U10927 ( .A(DB[2849]), .B(DB[2834]), .Z(n7333) );
  AND U10928 ( .A(n270), .B(n7334), .Z(n7332) );
  XOR U10929 ( .A(n7335), .B(n7336), .Z(n7334) );
  XOR U10930 ( .A(DB[2834]), .B(DB[2819]), .Z(n7336) );
  AND U10931 ( .A(n274), .B(n7337), .Z(n7335) );
  XOR U10932 ( .A(n7338), .B(n7339), .Z(n7337) );
  XOR U10933 ( .A(DB[2819]), .B(DB[2804]), .Z(n7339) );
  AND U10934 ( .A(n278), .B(n7340), .Z(n7338) );
  XOR U10935 ( .A(n7341), .B(n7342), .Z(n7340) );
  XOR U10936 ( .A(DB[2804]), .B(DB[2789]), .Z(n7342) );
  AND U10937 ( .A(n282), .B(n7343), .Z(n7341) );
  XOR U10938 ( .A(n7344), .B(n7345), .Z(n7343) );
  XOR U10939 ( .A(DB[2789]), .B(DB[2774]), .Z(n7345) );
  AND U10940 ( .A(n286), .B(n7346), .Z(n7344) );
  XOR U10941 ( .A(n7347), .B(n7348), .Z(n7346) );
  XOR U10942 ( .A(DB[2774]), .B(DB[2759]), .Z(n7348) );
  AND U10943 ( .A(n290), .B(n7349), .Z(n7347) );
  XOR U10944 ( .A(n7350), .B(n7351), .Z(n7349) );
  XOR U10945 ( .A(DB[2759]), .B(DB[2744]), .Z(n7351) );
  AND U10946 ( .A(n294), .B(n7352), .Z(n7350) );
  XOR U10947 ( .A(n7353), .B(n7354), .Z(n7352) );
  XOR U10948 ( .A(DB[2744]), .B(DB[2729]), .Z(n7354) );
  AND U10949 ( .A(n298), .B(n7355), .Z(n7353) );
  XOR U10950 ( .A(n7356), .B(n7357), .Z(n7355) );
  XOR U10951 ( .A(DB[2729]), .B(DB[2714]), .Z(n7357) );
  AND U10952 ( .A(n302), .B(n7358), .Z(n7356) );
  XOR U10953 ( .A(n7359), .B(n7360), .Z(n7358) );
  XOR U10954 ( .A(DB[2714]), .B(DB[2699]), .Z(n7360) );
  AND U10955 ( .A(n306), .B(n7361), .Z(n7359) );
  XOR U10956 ( .A(n7362), .B(n7363), .Z(n7361) );
  XOR U10957 ( .A(DB[2699]), .B(DB[2684]), .Z(n7363) );
  AND U10958 ( .A(n310), .B(n7364), .Z(n7362) );
  XOR U10959 ( .A(n7365), .B(n7366), .Z(n7364) );
  XOR U10960 ( .A(DB[2684]), .B(DB[2669]), .Z(n7366) );
  AND U10961 ( .A(n314), .B(n7367), .Z(n7365) );
  XOR U10962 ( .A(n7368), .B(n7369), .Z(n7367) );
  XOR U10963 ( .A(DB[2669]), .B(DB[2654]), .Z(n7369) );
  AND U10964 ( .A(n318), .B(n7370), .Z(n7368) );
  XOR U10965 ( .A(n7371), .B(n7372), .Z(n7370) );
  XOR U10966 ( .A(DB[2654]), .B(DB[2639]), .Z(n7372) );
  AND U10967 ( .A(n322), .B(n7373), .Z(n7371) );
  XOR U10968 ( .A(n7374), .B(n7375), .Z(n7373) );
  XOR U10969 ( .A(DB[2639]), .B(DB[2624]), .Z(n7375) );
  AND U10970 ( .A(n326), .B(n7376), .Z(n7374) );
  XOR U10971 ( .A(n7377), .B(n7378), .Z(n7376) );
  XOR U10972 ( .A(DB[2624]), .B(DB[2609]), .Z(n7378) );
  AND U10973 ( .A(n330), .B(n7379), .Z(n7377) );
  XOR U10974 ( .A(n7380), .B(n7381), .Z(n7379) );
  XOR U10975 ( .A(DB[2609]), .B(DB[2594]), .Z(n7381) );
  AND U10976 ( .A(n334), .B(n7382), .Z(n7380) );
  XOR U10977 ( .A(n7383), .B(n7384), .Z(n7382) );
  XOR U10978 ( .A(DB[2594]), .B(DB[2579]), .Z(n7384) );
  AND U10979 ( .A(n338), .B(n7385), .Z(n7383) );
  XOR U10980 ( .A(n7386), .B(n7387), .Z(n7385) );
  XOR U10981 ( .A(DB[2579]), .B(DB[2564]), .Z(n7387) );
  AND U10982 ( .A(n342), .B(n7388), .Z(n7386) );
  XOR U10983 ( .A(n7389), .B(n7390), .Z(n7388) );
  XOR U10984 ( .A(DB[2564]), .B(DB[2549]), .Z(n7390) );
  AND U10985 ( .A(n346), .B(n7391), .Z(n7389) );
  XOR U10986 ( .A(n7392), .B(n7393), .Z(n7391) );
  XOR U10987 ( .A(DB[2549]), .B(DB[2534]), .Z(n7393) );
  AND U10988 ( .A(n350), .B(n7394), .Z(n7392) );
  XOR U10989 ( .A(n7395), .B(n7396), .Z(n7394) );
  XOR U10990 ( .A(DB[2534]), .B(DB[2519]), .Z(n7396) );
  AND U10991 ( .A(n354), .B(n7397), .Z(n7395) );
  XOR U10992 ( .A(n7398), .B(n7399), .Z(n7397) );
  XOR U10993 ( .A(DB[2519]), .B(DB[2504]), .Z(n7399) );
  AND U10994 ( .A(n358), .B(n7400), .Z(n7398) );
  XOR U10995 ( .A(n7401), .B(n7402), .Z(n7400) );
  XOR U10996 ( .A(DB[2504]), .B(DB[2489]), .Z(n7402) );
  AND U10997 ( .A(n362), .B(n7403), .Z(n7401) );
  XOR U10998 ( .A(n7404), .B(n7405), .Z(n7403) );
  XOR U10999 ( .A(DB[2489]), .B(DB[2474]), .Z(n7405) );
  AND U11000 ( .A(n366), .B(n7406), .Z(n7404) );
  XOR U11001 ( .A(n7407), .B(n7408), .Z(n7406) );
  XOR U11002 ( .A(DB[2474]), .B(DB[2459]), .Z(n7408) );
  AND U11003 ( .A(n370), .B(n7409), .Z(n7407) );
  XOR U11004 ( .A(n7410), .B(n7411), .Z(n7409) );
  XOR U11005 ( .A(DB[2459]), .B(DB[2444]), .Z(n7411) );
  AND U11006 ( .A(n374), .B(n7412), .Z(n7410) );
  XOR U11007 ( .A(n7413), .B(n7414), .Z(n7412) );
  XOR U11008 ( .A(DB[2444]), .B(DB[2429]), .Z(n7414) );
  AND U11009 ( .A(n378), .B(n7415), .Z(n7413) );
  XOR U11010 ( .A(n7416), .B(n7417), .Z(n7415) );
  XOR U11011 ( .A(DB[2429]), .B(DB[2414]), .Z(n7417) );
  AND U11012 ( .A(n382), .B(n7418), .Z(n7416) );
  XOR U11013 ( .A(n7419), .B(n7420), .Z(n7418) );
  XOR U11014 ( .A(DB[2414]), .B(DB[2399]), .Z(n7420) );
  AND U11015 ( .A(n386), .B(n7421), .Z(n7419) );
  XOR U11016 ( .A(n7422), .B(n7423), .Z(n7421) );
  XOR U11017 ( .A(DB[2399]), .B(DB[2384]), .Z(n7423) );
  AND U11018 ( .A(n390), .B(n7424), .Z(n7422) );
  XOR U11019 ( .A(n7425), .B(n7426), .Z(n7424) );
  XOR U11020 ( .A(DB[2384]), .B(DB[2369]), .Z(n7426) );
  AND U11021 ( .A(n394), .B(n7427), .Z(n7425) );
  XOR U11022 ( .A(n7428), .B(n7429), .Z(n7427) );
  XOR U11023 ( .A(DB[2369]), .B(DB[2354]), .Z(n7429) );
  AND U11024 ( .A(n398), .B(n7430), .Z(n7428) );
  XOR U11025 ( .A(n7431), .B(n7432), .Z(n7430) );
  XOR U11026 ( .A(DB[2354]), .B(DB[2339]), .Z(n7432) );
  AND U11027 ( .A(n402), .B(n7433), .Z(n7431) );
  XOR U11028 ( .A(n7434), .B(n7435), .Z(n7433) );
  XOR U11029 ( .A(DB[2339]), .B(DB[2324]), .Z(n7435) );
  AND U11030 ( .A(n406), .B(n7436), .Z(n7434) );
  XOR U11031 ( .A(n7437), .B(n7438), .Z(n7436) );
  XOR U11032 ( .A(DB[2324]), .B(DB[2309]), .Z(n7438) );
  AND U11033 ( .A(n410), .B(n7439), .Z(n7437) );
  XOR U11034 ( .A(n7440), .B(n7441), .Z(n7439) );
  XOR U11035 ( .A(DB[2309]), .B(DB[2294]), .Z(n7441) );
  AND U11036 ( .A(n414), .B(n7442), .Z(n7440) );
  XOR U11037 ( .A(n7443), .B(n7444), .Z(n7442) );
  XOR U11038 ( .A(DB[2294]), .B(DB[2279]), .Z(n7444) );
  AND U11039 ( .A(n418), .B(n7445), .Z(n7443) );
  XOR U11040 ( .A(n7446), .B(n7447), .Z(n7445) );
  XOR U11041 ( .A(DB[2279]), .B(DB[2264]), .Z(n7447) );
  AND U11042 ( .A(n422), .B(n7448), .Z(n7446) );
  XOR U11043 ( .A(n7449), .B(n7450), .Z(n7448) );
  XOR U11044 ( .A(DB[2264]), .B(DB[2249]), .Z(n7450) );
  AND U11045 ( .A(n426), .B(n7451), .Z(n7449) );
  XOR U11046 ( .A(n7452), .B(n7453), .Z(n7451) );
  XOR U11047 ( .A(DB[2249]), .B(DB[2234]), .Z(n7453) );
  AND U11048 ( .A(n430), .B(n7454), .Z(n7452) );
  XOR U11049 ( .A(n7455), .B(n7456), .Z(n7454) );
  XOR U11050 ( .A(DB[2234]), .B(DB[2219]), .Z(n7456) );
  AND U11051 ( .A(n434), .B(n7457), .Z(n7455) );
  XOR U11052 ( .A(n7458), .B(n7459), .Z(n7457) );
  XOR U11053 ( .A(DB[2219]), .B(DB[2204]), .Z(n7459) );
  AND U11054 ( .A(n438), .B(n7460), .Z(n7458) );
  XOR U11055 ( .A(n7461), .B(n7462), .Z(n7460) );
  XOR U11056 ( .A(DB[2204]), .B(DB[2189]), .Z(n7462) );
  AND U11057 ( .A(n442), .B(n7463), .Z(n7461) );
  XOR U11058 ( .A(n7464), .B(n7465), .Z(n7463) );
  XOR U11059 ( .A(DB[2189]), .B(DB[2174]), .Z(n7465) );
  AND U11060 ( .A(n446), .B(n7466), .Z(n7464) );
  XOR U11061 ( .A(n7467), .B(n7468), .Z(n7466) );
  XOR U11062 ( .A(DB[2174]), .B(DB[2159]), .Z(n7468) );
  AND U11063 ( .A(n450), .B(n7469), .Z(n7467) );
  XOR U11064 ( .A(n7470), .B(n7471), .Z(n7469) );
  XOR U11065 ( .A(DB[2159]), .B(DB[2144]), .Z(n7471) );
  AND U11066 ( .A(n454), .B(n7472), .Z(n7470) );
  XOR U11067 ( .A(n7473), .B(n7474), .Z(n7472) );
  XOR U11068 ( .A(DB[2144]), .B(DB[2129]), .Z(n7474) );
  AND U11069 ( .A(n458), .B(n7475), .Z(n7473) );
  XOR U11070 ( .A(n7476), .B(n7477), .Z(n7475) );
  XOR U11071 ( .A(DB[2129]), .B(DB[2114]), .Z(n7477) );
  AND U11072 ( .A(n462), .B(n7478), .Z(n7476) );
  XOR U11073 ( .A(n7479), .B(n7480), .Z(n7478) );
  XOR U11074 ( .A(DB[2114]), .B(DB[2099]), .Z(n7480) );
  AND U11075 ( .A(n466), .B(n7481), .Z(n7479) );
  XOR U11076 ( .A(n7482), .B(n7483), .Z(n7481) );
  XOR U11077 ( .A(DB[2099]), .B(DB[2084]), .Z(n7483) );
  AND U11078 ( .A(n470), .B(n7484), .Z(n7482) );
  XOR U11079 ( .A(n7485), .B(n7486), .Z(n7484) );
  XOR U11080 ( .A(DB[2084]), .B(DB[2069]), .Z(n7486) );
  AND U11081 ( .A(n474), .B(n7487), .Z(n7485) );
  XOR U11082 ( .A(n7488), .B(n7489), .Z(n7487) );
  XOR U11083 ( .A(DB[2069]), .B(DB[2054]), .Z(n7489) );
  AND U11084 ( .A(n478), .B(n7490), .Z(n7488) );
  XOR U11085 ( .A(n7491), .B(n7492), .Z(n7490) );
  XOR U11086 ( .A(DB[2054]), .B(DB[2039]), .Z(n7492) );
  AND U11087 ( .A(n482), .B(n7493), .Z(n7491) );
  XOR U11088 ( .A(n7494), .B(n7495), .Z(n7493) );
  XOR U11089 ( .A(DB[2039]), .B(DB[2024]), .Z(n7495) );
  AND U11090 ( .A(n486), .B(n7496), .Z(n7494) );
  XOR U11091 ( .A(n7497), .B(n7498), .Z(n7496) );
  XOR U11092 ( .A(DB[2024]), .B(DB[2009]), .Z(n7498) );
  AND U11093 ( .A(n490), .B(n7499), .Z(n7497) );
  XOR U11094 ( .A(n7500), .B(n7501), .Z(n7499) );
  XOR U11095 ( .A(DB[2009]), .B(DB[1994]), .Z(n7501) );
  AND U11096 ( .A(n494), .B(n7502), .Z(n7500) );
  XOR U11097 ( .A(n7503), .B(n7504), .Z(n7502) );
  XOR U11098 ( .A(DB[1994]), .B(DB[1979]), .Z(n7504) );
  AND U11099 ( .A(n498), .B(n7505), .Z(n7503) );
  XOR U11100 ( .A(n7506), .B(n7507), .Z(n7505) );
  XOR U11101 ( .A(DB[1979]), .B(DB[1964]), .Z(n7507) );
  AND U11102 ( .A(n502), .B(n7508), .Z(n7506) );
  XOR U11103 ( .A(n7509), .B(n7510), .Z(n7508) );
  XOR U11104 ( .A(DB[1964]), .B(DB[1949]), .Z(n7510) );
  AND U11105 ( .A(n506), .B(n7511), .Z(n7509) );
  XOR U11106 ( .A(n7512), .B(n7513), .Z(n7511) );
  XOR U11107 ( .A(DB[1949]), .B(DB[1934]), .Z(n7513) );
  AND U11108 ( .A(n510), .B(n7514), .Z(n7512) );
  XOR U11109 ( .A(n7515), .B(n7516), .Z(n7514) );
  XOR U11110 ( .A(DB[1934]), .B(DB[1919]), .Z(n7516) );
  AND U11111 ( .A(n514), .B(n7517), .Z(n7515) );
  XOR U11112 ( .A(n7518), .B(n7519), .Z(n7517) );
  XOR U11113 ( .A(DB[1919]), .B(DB[1904]), .Z(n7519) );
  AND U11114 ( .A(n518), .B(n7520), .Z(n7518) );
  XOR U11115 ( .A(n7521), .B(n7522), .Z(n7520) );
  XOR U11116 ( .A(DB[1904]), .B(DB[1889]), .Z(n7522) );
  AND U11117 ( .A(n522), .B(n7523), .Z(n7521) );
  XOR U11118 ( .A(n7524), .B(n7525), .Z(n7523) );
  XOR U11119 ( .A(DB[1889]), .B(DB[1874]), .Z(n7525) );
  AND U11120 ( .A(n526), .B(n7526), .Z(n7524) );
  XOR U11121 ( .A(n7527), .B(n7528), .Z(n7526) );
  XOR U11122 ( .A(DB[1874]), .B(DB[1859]), .Z(n7528) );
  AND U11123 ( .A(n530), .B(n7529), .Z(n7527) );
  XOR U11124 ( .A(n7530), .B(n7531), .Z(n7529) );
  XOR U11125 ( .A(DB[1859]), .B(DB[1844]), .Z(n7531) );
  AND U11126 ( .A(n534), .B(n7532), .Z(n7530) );
  XOR U11127 ( .A(n7533), .B(n7534), .Z(n7532) );
  XOR U11128 ( .A(DB[1844]), .B(DB[1829]), .Z(n7534) );
  AND U11129 ( .A(n538), .B(n7535), .Z(n7533) );
  XOR U11130 ( .A(n7536), .B(n7537), .Z(n7535) );
  XOR U11131 ( .A(DB[1829]), .B(DB[1814]), .Z(n7537) );
  AND U11132 ( .A(n542), .B(n7538), .Z(n7536) );
  XOR U11133 ( .A(n7539), .B(n7540), .Z(n7538) );
  XOR U11134 ( .A(DB[1814]), .B(DB[1799]), .Z(n7540) );
  AND U11135 ( .A(n546), .B(n7541), .Z(n7539) );
  XOR U11136 ( .A(n7542), .B(n7543), .Z(n7541) );
  XOR U11137 ( .A(DB[1799]), .B(DB[1784]), .Z(n7543) );
  AND U11138 ( .A(n550), .B(n7544), .Z(n7542) );
  XOR U11139 ( .A(n7545), .B(n7546), .Z(n7544) );
  XOR U11140 ( .A(DB[1784]), .B(DB[1769]), .Z(n7546) );
  AND U11141 ( .A(n554), .B(n7547), .Z(n7545) );
  XOR U11142 ( .A(n7548), .B(n7549), .Z(n7547) );
  XOR U11143 ( .A(DB[1769]), .B(DB[1754]), .Z(n7549) );
  AND U11144 ( .A(n558), .B(n7550), .Z(n7548) );
  XOR U11145 ( .A(n7551), .B(n7552), .Z(n7550) );
  XOR U11146 ( .A(DB[1754]), .B(DB[1739]), .Z(n7552) );
  AND U11147 ( .A(n562), .B(n7553), .Z(n7551) );
  XOR U11148 ( .A(n7554), .B(n7555), .Z(n7553) );
  XOR U11149 ( .A(DB[1739]), .B(DB[1724]), .Z(n7555) );
  AND U11150 ( .A(n566), .B(n7556), .Z(n7554) );
  XOR U11151 ( .A(n7557), .B(n7558), .Z(n7556) );
  XOR U11152 ( .A(DB[1724]), .B(DB[1709]), .Z(n7558) );
  AND U11153 ( .A(n570), .B(n7559), .Z(n7557) );
  XOR U11154 ( .A(n7560), .B(n7561), .Z(n7559) );
  XOR U11155 ( .A(DB[1709]), .B(DB[1694]), .Z(n7561) );
  AND U11156 ( .A(n574), .B(n7562), .Z(n7560) );
  XOR U11157 ( .A(n7563), .B(n7564), .Z(n7562) );
  XOR U11158 ( .A(DB[1694]), .B(DB[1679]), .Z(n7564) );
  AND U11159 ( .A(n578), .B(n7565), .Z(n7563) );
  XOR U11160 ( .A(n7566), .B(n7567), .Z(n7565) );
  XOR U11161 ( .A(DB[1679]), .B(DB[1664]), .Z(n7567) );
  AND U11162 ( .A(n582), .B(n7568), .Z(n7566) );
  XOR U11163 ( .A(n7569), .B(n7570), .Z(n7568) );
  XOR U11164 ( .A(DB[1664]), .B(DB[1649]), .Z(n7570) );
  AND U11165 ( .A(n586), .B(n7571), .Z(n7569) );
  XOR U11166 ( .A(n7572), .B(n7573), .Z(n7571) );
  XOR U11167 ( .A(DB[1649]), .B(DB[1634]), .Z(n7573) );
  AND U11168 ( .A(n590), .B(n7574), .Z(n7572) );
  XOR U11169 ( .A(n7575), .B(n7576), .Z(n7574) );
  XOR U11170 ( .A(DB[1634]), .B(DB[1619]), .Z(n7576) );
  AND U11171 ( .A(n594), .B(n7577), .Z(n7575) );
  XOR U11172 ( .A(n7578), .B(n7579), .Z(n7577) );
  XOR U11173 ( .A(DB[1619]), .B(DB[1604]), .Z(n7579) );
  AND U11174 ( .A(n598), .B(n7580), .Z(n7578) );
  XOR U11175 ( .A(n7581), .B(n7582), .Z(n7580) );
  XOR U11176 ( .A(DB[1604]), .B(DB[1589]), .Z(n7582) );
  AND U11177 ( .A(n602), .B(n7583), .Z(n7581) );
  XOR U11178 ( .A(n7584), .B(n7585), .Z(n7583) );
  XOR U11179 ( .A(DB[1589]), .B(DB[1574]), .Z(n7585) );
  AND U11180 ( .A(n606), .B(n7586), .Z(n7584) );
  XOR U11181 ( .A(n7587), .B(n7588), .Z(n7586) );
  XOR U11182 ( .A(DB[1574]), .B(DB[1559]), .Z(n7588) );
  AND U11183 ( .A(n610), .B(n7589), .Z(n7587) );
  XOR U11184 ( .A(n7590), .B(n7591), .Z(n7589) );
  XOR U11185 ( .A(DB[1559]), .B(DB[1544]), .Z(n7591) );
  AND U11186 ( .A(n614), .B(n7592), .Z(n7590) );
  XOR U11187 ( .A(n7593), .B(n7594), .Z(n7592) );
  XOR U11188 ( .A(DB[1544]), .B(DB[1529]), .Z(n7594) );
  AND U11189 ( .A(n618), .B(n7595), .Z(n7593) );
  XOR U11190 ( .A(n7596), .B(n7597), .Z(n7595) );
  XOR U11191 ( .A(DB[1529]), .B(DB[1514]), .Z(n7597) );
  AND U11192 ( .A(n622), .B(n7598), .Z(n7596) );
  XOR U11193 ( .A(n7599), .B(n7600), .Z(n7598) );
  XOR U11194 ( .A(DB[1514]), .B(DB[1499]), .Z(n7600) );
  AND U11195 ( .A(n626), .B(n7601), .Z(n7599) );
  XOR U11196 ( .A(n7602), .B(n7603), .Z(n7601) );
  XOR U11197 ( .A(DB[1499]), .B(DB[1484]), .Z(n7603) );
  AND U11198 ( .A(n630), .B(n7604), .Z(n7602) );
  XOR U11199 ( .A(n7605), .B(n7606), .Z(n7604) );
  XOR U11200 ( .A(DB[1484]), .B(DB[1469]), .Z(n7606) );
  AND U11201 ( .A(n634), .B(n7607), .Z(n7605) );
  XOR U11202 ( .A(n7608), .B(n7609), .Z(n7607) );
  XOR U11203 ( .A(DB[1469]), .B(DB[1454]), .Z(n7609) );
  AND U11204 ( .A(n638), .B(n7610), .Z(n7608) );
  XOR U11205 ( .A(n7611), .B(n7612), .Z(n7610) );
  XOR U11206 ( .A(DB[1454]), .B(DB[1439]), .Z(n7612) );
  AND U11207 ( .A(n642), .B(n7613), .Z(n7611) );
  XOR U11208 ( .A(n7614), .B(n7615), .Z(n7613) );
  XOR U11209 ( .A(DB[1439]), .B(DB[1424]), .Z(n7615) );
  AND U11210 ( .A(n646), .B(n7616), .Z(n7614) );
  XOR U11211 ( .A(n7617), .B(n7618), .Z(n7616) );
  XOR U11212 ( .A(DB[1424]), .B(DB[1409]), .Z(n7618) );
  AND U11213 ( .A(n650), .B(n7619), .Z(n7617) );
  XOR U11214 ( .A(n7620), .B(n7621), .Z(n7619) );
  XOR U11215 ( .A(DB[1409]), .B(DB[1394]), .Z(n7621) );
  AND U11216 ( .A(n654), .B(n7622), .Z(n7620) );
  XOR U11217 ( .A(n7623), .B(n7624), .Z(n7622) );
  XOR U11218 ( .A(DB[1394]), .B(DB[1379]), .Z(n7624) );
  AND U11219 ( .A(n658), .B(n7625), .Z(n7623) );
  XOR U11220 ( .A(n7626), .B(n7627), .Z(n7625) );
  XOR U11221 ( .A(DB[1379]), .B(DB[1364]), .Z(n7627) );
  AND U11222 ( .A(n662), .B(n7628), .Z(n7626) );
  XOR U11223 ( .A(n7629), .B(n7630), .Z(n7628) );
  XOR U11224 ( .A(DB[1364]), .B(DB[1349]), .Z(n7630) );
  AND U11225 ( .A(n666), .B(n7631), .Z(n7629) );
  XOR U11226 ( .A(n7632), .B(n7633), .Z(n7631) );
  XOR U11227 ( .A(DB[1349]), .B(DB[1334]), .Z(n7633) );
  AND U11228 ( .A(n670), .B(n7634), .Z(n7632) );
  XOR U11229 ( .A(n7635), .B(n7636), .Z(n7634) );
  XOR U11230 ( .A(DB[1334]), .B(DB[1319]), .Z(n7636) );
  AND U11231 ( .A(n674), .B(n7637), .Z(n7635) );
  XOR U11232 ( .A(n7638), .B(n7639), .Z(n7637) );
  XOR U11233 ( .A(DB[1319]), .B(DB[1304]), .Z(n7639) );
  AND U11234 ( .A(n678), .B(n7640), .Z(n7638) );
  XOR U11235 ( .A(n7641), .B(n7642), .Z(n7640) );
  XOR U11236 ( .A(DB[1304]), .B(DB[1289]), .Z(n7642) );
  AND U11237 ( .A(n682), .B(n7643), .Z(n7641) );
  XOR U11238 ( .A(n7644), .B(n7645), .Z(n7643) );
  XOR U11239 ( .A(DB[1289]), .B(DB[1274]), .Z(n7645) );
  AND U11240 ( .A(n686), .B(n7646), .Z(n7644) );
  XOR U11241 ( .A(n7647), .B(n7648), .Z(n7646) );
  XOR U11242 ( .A(DB[1274]), .B(DB[1259]), .Z(n7648) );
  AND U11243 ( .A(n690), .B(n7649), .Z(n7647) );
  XOR U11244 ( .A(n7650), .B(n7651), .Z(n7649) );
  XOR U11245 ( .A(DB[1259]), .B(DB[1244]), .Z(n7651) );
  AND U11246 ( .A(n694), .B(n7652), .Z(n7650) );
  XOR U11247 ( .A(n7653), .B(n7654), .Z(n7652) );
  XOR U11248 ( .A(DB[1244]), .B(DB[1229]), .Z(n7654) );
  AND U11249 ( .A(n698), .B(n7655), .Z(n7653) );
  XOR U11250 ( .A(n7656), .B(n7657), .Z(n7655) );
  XOR U11251 ( .A(DB[1229]), .B(DB[1214]), .Z(n7657) );
  AND U11252 ( .A(n702), .B(n7658), .Z(n7656) );
  XOR U11253 ( .A(n7659), .B(n7660), .Z(n7658) );
  XOR U11254 ( .A(DB[1214]), .B(DB[1199]), .Z(n7660) );
  AND U11255 ( .A(n706), .B(n7661), .Z(n7659) );
  XOR U11256 ( .A(n7662), .B(n7663), .Z(n7661) );
  XOR U11257 ( .A(DB[1199]), .B(DB[1184]), .Z(n7663) );
  AND U11258 ( .A(n710), .B(n7664), .Z(n7662) );
  XOR U11259 ( .A(n7665), .B(n7666), .Z(n7664) );
  XOR U11260 ( .A(DB[1184]), .B(DB[1169]), .Z(n7666) );
  AND U11261 ( .A(n714), .B(n7667), .Z(n7665) );
  XOR U11262 ( .A(n7668), .B(n7669), .Z(n7667) );
  XOR U11263 ( .A(DB[1169]), .B(DB[1154]), .Z(n7669) );
  AND U11264 ( .A(n718), .B(n7670), .Z(n7668) );
  XOR U11265 ( .A(n7671), .B(n7672), .Z(n7670) );
  XOR U11266 ( .A(DB[1154]), .B(DB[1139]), .Z(n7672) );
  AND U11267 ( .A(n722), .B(n7673), .Z(n7671) );
  XOR U11268 ( .A(n7674), .B(n7675), .Z(n7673) );
  XOR U11269 ( .A(DB[1139]), .B(DB[1124]), .Z(n7675) );
  AND U11270 ( .A(n726), .B(n7676), .Z(n7674) );
  XOR U11271 ( .A(n7677), .B(n7678), .Z(n7676) );
  XOR U11272 ( .A(DB[1124]), .B(DB[1109]), .Z(n7678) );
  AND U11273 ( .A(n730), .B(n7679), .Z(n7677) );
  XOR U11274 ( .A(n7680), .B(n7681), .Z(n7679) );
  XOR U11275 ( .A(DB[1109]), .B(DB[1094]), .Z(n7681) );
  AND U11276 ( .A(n734), .B(n7682), .Z(n7680) );
  XOR U11277 ( .A(n7683), .B(n7684), .Z(n7682) );
  XOR U11278 ( .A(DB[1094]), .B(DB[1079]), .Z(n7684) );
  AND U11279 ( .A(n738), .B(n7685), .Z(n7683) );
  XOR U11280 ( .A(n7686), .B(n7687), .Z(n7685) );
  XOR U11281 ( .A(DB[1079]), .B(DB[1064]), .Z(n7687) );
  AND U11282 ( .A(n742), .B(n7688), .Z(n7686) );
  XOR U11283 ( .A(n7689), .B(n7690), .Z(n7688) );
  XOR U11284 ( .A(DB[1064]), .B(DB[1049]), .Z(n7690) );
  AND U11285 ( .A(n746), .B(n7691), .Z(n7689) );
  XOR U11286 ( .A(n7692), .B(n7693), .Z(n7691) );
  XOR U11287 ( .A(DB[1049]), .B(DB[1034]), .Z(n7693) );
  AND U11288 ( .A(n750), .B(n7694), .Z(n7692) );
  XOR U11289 ( .A(n7695), .B(n7696), .Z(n7694) );
  XOR U11290 ( .A(DB[1034]), .B(DB[1019]), .Z(n7696) );
  AND U11291 ( .A(n754), .B(n7697), .Z(n7695) );
  XOR U11292 ( .A(n7698), .B(n7699), .Z(n7697) );
  XOR U11293 ( .A(DB[1019]), .B(DB[1004]), .Z(n7699) );
  AND U11294 ( .A(n758), .B(n7700), .Z(n7698) );
  XOR U11295 ( .A(n7701), .B(n7702), .Z(n7700) );
  XOR U11296 ( .A(DB[989]), .B(DB[1004]), .Z(n7702) );
  AND U11297 ( .A(n762), .B(n7703), .Z(n7701) );
  XOR U11298 ( .A(n7704), .B(n7705), .Z(n7703) );
  XOR U11299 ( .A(DB[989]), .B(DB[974]), .Z(n7705) );
  AND U11300 ( .A(n766), .B(n7706), .Z(n7704) );
  XOR U11301 ( .A(n7707), .B(n7708), .Z(n7706) );
  XOR U11302 ( .A(DB[974]), .B(DB[959]), .Z(n7708) );
  AND U11303 ( .A(n770), .B(n7709), .Z(n7707) );
  XOR U11304 ( .A(n7710), .B(n7711), .Z(n7709) );
  XOR U11305 ( .A(DB[959]), .B(DB[944]), .Z(n7711) );
  AND U11306 ( .A(n774), .B(n7712), .Z(n7710) );
  XOR U11307 ( .A(n7713), .B(n7714), .Z(n7712) );
  XOR U11308 ( .A(DB[944]), .B(DB[929]), .Z(n7714) );
  AND U11309 ( .A(n778), .B(n7715), .Z(n7713) );
  XOR U11310 ( .A(n7716), .B(n7717), .Z(n7715) );
  XOR U11311 ( .A(DB[929]), .B(DB[914]), .Z(n7717) );
  AND U11312 ( .A(n782), .B(n7718), .Z(n7716) );
  XOR U11313 ( .A(n7719), .B(n7720), .Z(n7718) );
  XOR U11314 ( .A(DB[914]), .B(DB[899]), .Z(n7720) );
  AND U11315 ( .A(n786), .B(n7721), .Z(n7719) );
  XOR U11316 ( .A(n7722), .B(n7723), .Z(n7721) );
  XOR U11317 ( .A(DB[899]), .B(DB[884]), .Z(n7723) );
  AND U11318 ( .A(n790), .B(n7724), .Z(n7722) );
  XOR U11319 ( .A(n7725), .B(n7726), .Z(n7724) );
  XOR U11320 ( .A(DB[884]), .B(DB[869]), .Z(n7726) );
  AND U11321 ( .A(n794), .B(n7727), .Z(n7725) );
  XOR U11322 ( .A(n7728), .B(n7729), .Z(n7727) );
  XOR U11323 ( .A(DB[869]), .B(DB[854]), .Z(n7729) );
  AND U11324 ( .A(n798), .B(n7730), .Z(n7728) );
  XOR U11325 ( .A(n7731), .B(n7732), .Z(n7730) );
  XOR U11326 ( .A(DB[854]), .B(DB[839]), .Z(n7732) );
  AND U11327 ( .A(n802), .B(n7733), .Z(n7731) );
  XOR U11328 ( .A(n7734), .B(n7735), .Z(n7733) );
  XOR U11329 ( .A(DB[839]), .B(DB[824]), .Z(n7735) );
  AND U11330 ( .A(n806), .B(n7736), .Z(n7734) );
  XOR U11331 ( .A(n7737), .B(n7738), .Z(n7736) );
  XOR U11332 ( .A(DB[824]), .B(DB[809]), .Z(n7738) );
  AND U11333 ( .A(n810), .B(n7739), .Z(n7737) );
  XOR U11334 ( .A(n7740), .B(n7741), .Z(n7739) );
  XOR U11335 ( .A(DB[809]), .B(DB[794]), .Z(n7741) );
  AND U11336 ( .A(n814), .B(n7742), .Z(n7740) );
  XOR U11337 ( .A(n7743), .B(n7744), .Z(n7742) );
  XOR U11338 ( .A(DB[794]), .B(DB[779]), .Z(n7744) );
  AND U11339 ( .A(n818), .B(n7745), .Z(n7743) );
  XOR U11340 ( .A(n7746), .B(n7747), .Z(n7745) );
  XOR U11341 ( .A(DB[779]), .B(DB[764]), .Z(n7747) );
  AND U11342 ( .A(n822), .B(n7748), .Z(n7746) );
  XOR U11343 ( .A(n7749), .B(n7750), .Z(n7748) );
  XOR U11344 ( .A(DB[764]), .B(DB[749]), .Z(n7750) );
  AND U11345 ( .A(n826), .B(n7751), .Z(n7749) );
  XOR U11346 ( .A(n7752), .B(n7753), .Z(n7751) );
  XOR U11347 ( .A(DB[749]), .B(DB[734]), .Z(n7753) );
  AND U11348 ( .A(n830), .B(n7754), .Z(n7752) );
  XOR U11349 ( .A(n7755), .B(n7756), .Z(n7754) );
  XOR U11350 ( .A(DB[734]), .B(DB[719]), .Z(n7756) );
  AND U11351 ( .A(n834), .B(n7757), .Z(n7755) );
  XOR U11352 ( .A(n7758), .B(n7759), .Z(n7757) );
  XOR U11353 ( .A(DB[719]), .B(DB[704]), .Z(n7759) );
  AND U11354 ( .A(n838), .B(n7760), .Z(n7758) );
  XOR U11355 ( .A(n7761), .B(n7762), .Z(n7760) );
  XOR U11356 ( .A(DB[704]), .B(DB[689]), .Z(n7762) );
  AND U11357 ( .A(n842), .B(n7763), .Z(n7761) );
  XOR U11358 ( .A(n7764), .B(n7765), .Z(n7763) );
  XOR U11359 ( .A(DB[689]), .B(DB[674]), .Z(n7765) );
  AND U11360 ( .A(n846), .B(n7766), .Z(n7764) );
  XOR U11361 ( .A(n7767), .B(n7768), .Z(n7766) );
  XOR U11362 ( .A(DB[674]), .B(DB[659]), .Z(n7768) );
  AND U11363 ( .A(n850), .B(n7769), .Z(n7767) );
  XOR U11364 ( .A(n7770), .B(n7771), .Z(n7769) );
  XOR U11365 ( .A(DB[659]), .B(DB[644]), .Z(n7771) );
  AND U11366 ( .A(n854), .B(n7772), .Z(n7770) );
  XOR U11367 ( .A(n7773), .B(n7774), .Z(n7772) );
  XOR U11368 ( .A(DB[644]), .B(DB[629]), .Z(n7774) );
  AND U11369 ( .A(n858), .B(n7775), .Z(n7773) );
  XOR U11370 ( .A(n7776), .B(n7777), .Z(n7775) );
  XOR U11371 ( .A(DB[629]), .B(DB[614]), .Z(n7777) );
  AND U11372 ( .A(n862), .B(n7778), .Z(n7776) );
  XOR U11373 ( .A(n7779), .B(n7780), .Z(n7778) );
  XOR U11374 ( .A(DB[614]), .B(DB[599]), .Z(n7780) );
  AND U11375 ( .A(n866), .B(n7781), .Z(n7779) );
  XOR U11376 ( .A(n7782), .B(n7783), .Z(n7781) );
  XOR U11377 ( .A(DB[599]), .B(DB[584]), .Z(n7783) );
  AND U11378 ( .A(n870), .B(n7784), .Z(n7782) );
  XOR U11379 ( .A(n7785), .B(n7786), .Z(n7784) );
  XOR U11380 ( .A(DB[584]), .B(DB[569]), .Z(n7786) );
  AND U11381 ( .A(n874), .B(n7787), .Z(n7785) );
  XOR U11382 ( .A(n7788), .B(n7789), .Z(n7787) );
  XOR U11383 ( .A(DB[569]), .B(DB[554]), .Z(n7789) );
  AND U11384 ( .A(n878), .B(n7790), .Z(n7788) );
  XOR U11385 ( .A(n7791), .B(n7792), .Z(n7790) );
  XOR U11386 ( .A(DB[554]), .B(DB[539]), .Z(n7792) );
  AND U11387 ( .A(n882), .B(n7793), .Z(n7791) );
  XOR U11388 ( .A(n7794), .B(n7795), .Z(n7793) );
  XOR U11389 ( .A(DB[539]), .B(DB[524]), .Z(n7795) );
  AND U11390 ( .A(n886), .B(n7796), .Z(n7794) );
  XOR U11391 ( .A(n7797), .B(n7798), .Z(n7796) );
  XOR U11392 ( .A(DB[524]), .B(DB[509]), .Z(n7798) );
  AND U11393 ( .A(n890), .B(n7799), .Z(n7797) );
  XOR U11394 ( .A(n7800), .B(n7801), .Z(n7799) );
  XOR U11395 ( .A(DB[509]), .B(DB[494]), .Z(n7801) );
  AND U11396 ( .A(n894), .B(n7802), .Z(n7800) );
  XOR U11397 ( .A(n7803), .B(n7804), .Z(n7802) );
  XOR U11398 ( .A(DB[494]), .B(DB[479]), .Z(n7804) );
  AND U11399 ( .A(n898), .B(n7805), .Z(n7803) );
  XOR U11400 ( .A(n7806), .B(n7807), .Z(n7805) );
  XOR U11401 ( .A(DB[479]), .B(DB[464]), .Z(n7807) );
  AND U11402 ( .A(n902), .B(n7808), .Z(n7806) );
  XOR U11403 ( .A(n7809), .B(n7810), .Z(n7808) );
  XOR U11404 ( .A(DB[464]), .B(DB[449]), .Z(n7810) );
  AND U11405 ( .A(n906), .B(n7811), .Z(n7809) );
  XOR U11406 ( .A(n7812), .B(n7813), .Z(n7811) );
  XOR U11407 ( .A(DB[449]), .B(DB[434]), .Z(n7813) );
  AND U11408 ( .A(n910), .B(n7814), .Z(n7812) );
  XOR U11409 ( .A(n7815), .B(n7816), .Z(n7814) );
  XOR U11410 ( .A(DB[434]), .B(DB[419]), .Z(n7816) );
  AND U11411 ( .A(n914), .B(n7817), .Z(n7815) );
  XOR U11412 ( .A(n7818), .B(n7819), .Z(n7817) );
  XOR U11413 ( .A(DB[419]), .B(DB[404]), .Z(n7819) );
  AND U11414 ( .A(n918), .B(n7820), .Z(n7818) );
  XOR U11415 ( .A(n7821), .B(n7822), .Z(n7820) );
  XOR U11416 ( .A(DB[404]), .B(DB[389]), .Z(n7822) );
  AND U11417 ( .A(n922), .B(n7823), .Z(n7821) );
  XOR U11418 ( .A(n7824), .B(n7825), .Z(n7823) );
  XOR U11419 ( .A(DB[389]), .B(DB[374]), .Z(n7825) );
  AND U11420 ( .A(n926), .B(n7826), .Z(n7824) );
  XOR U11421 ( .A(n7827), .B(n7828), .Z(n7826) );
  XOR U11422 ( .A(DB[374]), .B(DB[359]), .Z(n7828) );
  AND U11423 ( .A(n930), .B(n7829), .Z(n7827) );
  XOR U11424 ( .A(n7830), .B(n7831), .Z(n7829) );
  XOR U11425 ( .A(DB[359]), .B(DB[344]), .Z(n7831) );
  AND U11426 ( .A(n934), .B(n7832), .Z(n7830) );
  XOR U11427 ( .A(n7833), .B(n7834), .Z(n7832) );
  XOR U11428 ( .A(DB[344]), .B(DB[329]), .Z(n7834) );
  AND U11429 ( .A(n938), .B(n7835), .Z(n7833) );
  XOR U11430 ( .A(n7836), .B(n7837), .Z(n7835) );
  XOR U11431 ( .A(DB[329]), .B(DB[314]), .Z(n7837) );
  AND U11432 ( .A(n942), .B(n7838), .Z(n7836) );
  XOR U11433 ( .A(n7839), .B(n7840), .Z(n7838) );
  XOR U11434 ( .A(DB[314]), .B(DB[299]), .Z(n7840) );
  AND U11435 ( .A(n946), .B(n7841), .Z(n7839) );
  XOR U11436 ( .A(n7842), .B(n7843), .Z(n7841) );
  XOR U11437 ( .A(DB[299]), .B(DB[284]), .Z(n7843) );
  AND U11438 ( .A(n950), .B(n7844), .Z(n7842) );
  XOR U11439 ( .A(n7845), .B(n7846), .Z(n7844) );
  XOR U11440 ( .A(DB[284]), .B(DB[269]), .Z(n7846) );
  AND U11441 ( .A(n954), .B(n7847), .Z(n7845) );
  XOR U11442 ( .A(n7848), .B(n7849), .Z(n7847) );
  XOR U11443 ( .A(DB[269]), .B(DB[254]), .Z(n7849) );
  AND U11444 ( .A(n958), .B(n7850), .Z(n7848) );
  XOR U11445 ( .A(n7851), .B(n7852), .Z(n7850) );
  XOR U11446 ( .A(DB[254]), .B(DB[239]), .Z(n7852) );
  AND U11447 ( .A(n962), .B(n7853), .Z(n7851) );
  XOR U11448 ( .A(n7854), .B(n7855), .Z(n7853) );
  XOR U11449 ( .A(DB[239]), .B(DB[224]), .Z(n7855) );
  AND U11450 ( .A(n966), .B(n7856), .Z(n7854) );
  XOR U11451 ( .A(n7857), .B(n7858), .Z(n7856) );
  XOR U11452 ( .A(DB[224]), .B(DB[209]), .Z(n7858) );
  AND U11453 ( .A(n970), .B(n7859), .Z(n7857) );
  XOR U11454 ( .A(n7860), .B(n7861), .Z(n7859) );
  XOR U11455 ( .A(DB[209]), .B(DB[194]), .Z(n7861) );
  AND U11456 ( .A(n974), .B(n7862), .Z(n7860) );
  XOR U11457 ( .A(n7863), .B(n7864), .Z(n7862) );
  XOR U11458 ( .A(DB[194]), .B(DB[179]), .Z(n7864) );
  AND U11459 ( .A(n978), .B(n7865), .Z(n7863) );
  XOR U11460 ( .A(n7866), .B(n7867), .Z(n7865) );
  XOR U11461 ( .A(DB[179]), .B(DB[164]), .Z(n7867) );
  AND U11462 ( .A(n982), .B(n7868), .Z(n7866) );
  XOR U11463 ( .A(n7869), .B(n7870), .Z(n7868) );
  XOR U11464 ( .A(DB[164]), .B(DB[149]), .Z(n7870) );
  AND U11465 ( .A(n986), .B(n7871), .Z(n7869) );
  XOR U11466 ( .A(n7872), .B(n7873), .Z(n7871) );
  XOR U11467 ( .A(DB[149]), .B(DB[134]), .Z(n7873) );
  AND U11468 ( .A(n990), .B(n7874), .Z(n7872) );
  XOR U11469 ( .A(n7875), .B(n7876), .Z(n7874) );
  XOR U11470 ( .A(DB[134]), .B(DB[119]), .Z(n7876) );
  AND U11471 ( .A(n994), .B(n7877), .Z(n7875) );
  XOR U11472 ( .A(n7878), .B(n7879), .Z(n7877) );
  XOR U11473 ( .A(DB[119]), .B(DB[104]), .Z(n7879) );
  AND U11474 ( .A(n998), .B(n7880), .Z(n7878) );
  XOR U11475 ( .A(n7881), .B(n7882), .Z(n7880) );
  XOR U11476 ( .A(DB[89]), .B(DB[104]), .Z(n7882) );
  AND U11477 ( .A(n1002), .B(n7883), .Z(n7881) );
  XOR U11478 ( .A(n7884), .B(n7885), .Z(n7883) );
  XOR U11479 ( .A(DB[89]), .B(DB[74]), .Z(n7885) );
  AND U11480 ( .A(n1006), .B(n7886), .Z(n7884) );
  XOR U11481 ( .A(n7887), .B(n7888), .Z(n7886) );
  XOR U11482 ( .A(DB[74]), .B(DB[59]), .Z(n7888) );
  AND U11483 ( .A(n1010), .B(n7889), .Z(n7887) );
  XOR U11484 ( .A(n7890), .B(n7891), .Z(n7889) );
  XOR U11485 ( .A(DB[59]), .B(DB[44]), .Z(n7891) );
  AND U11486 ( .A(n1014), .B(n7892), .Z(n7890) );
  XOR U11487 ( .A(n7893), .B(n7894), .Z(n7892) );
  XOR U11488 ( .A(DB[44]), .B(DB[29]), .Z(n7894) );
  AND U11489 ( .A(n1018), .B(n7895), .Z(n7893) );
  XOR U11490 ( .A(DB[29]), .B(DB[14]), .Z(n7895) );
  XOR U11491 ( .A(DB[3838]), .B(n7896), .Z(min_val_out[13]) );
  AND U11492 ( .A(n2), .B(n7897), .Z(n7896) );
  XOR U11493 ( .A(n7898), .B(n7899), .Z(n7897) );
  XOR U11494 ( .A(DB[3838]), .B(DB[3823]), .Z(n7899) );
  AND U11495 ( .A(n6), .B(n7900), .Z(n7898) );
  XOR U11496 ( .A(n7901), .B(n7902), .Z(n7900) );
  XOR U11497 ( .A(DB[3823]), .B(DB[3808]), .Z(n7902) );
  AND U11498 ( .A(n10), .B(n7903), .Z(n7901) );
  XOR U11499 ( .A(n7904), .B(n7905), .Z(n7903) );
  XOR U11500 ( .A(DB[3808]), .B(DB[3793]), .Z(n7905) );
  AND U11501 ( .A(n14), .B(n7906), .Z(n7904) );
  XOR U11502 ( .A(n7907), .B(n7908), .Z(n7906) );
  XOR U11503 ( .A(DB[3793]), .B(DB[3778]), .Z(n7908) );
  AND U11504 ( .A(n18), .B(n7909), .Z(n7907) );
  XOR U11505 ( .A(n7910), .B(n7911), .Z(n7909) );
  XOR U11506 ( .A(DB[3778]), .B(DB[3763]), .Z(n7911) );
  AND U11507 ( .A(n22), .B(n7912), .Z(n7910) );
  XOR U11508 ( .A(n7913), .B(n7914), .Z(n7912) );
  XOR U11509 ( .A(DB[3763]), .B(DB[3748]), .Z(n7914) );
  AND U11510 ( .A(n26), .B(n7915), .Z(n7913) );
  XOR U11511 ( .A(n7916), .B(n7917), .Z(n7915) );
  XOR U11512 ( .A(DB[3748]), .B(DB[3733]), .Z(n7917) );
  AND U11513 ( .A(n30), .B(n7918), .Z(n7916) );
  XOR U11514 ( .A(n7919), .B(n7920), .Z(n7918) );
  XOR U11515 ( .A(DB[3733]), .B(DB[3718]), .Z(n7920) );
  AND U11516 ( .A(n34), .B(n7921), .Z(n7919) );
  XOR U11517 ( .A(n7922), .B(n7923), .Z(n7921) );
  XOR U11518 ( .A(DB[3718]), .B(DB[3703]), .Z(n7923) );
  AND U11519 ( .A(n38), .B(n7924), .Z(n7922) );
  XOR U11520 ( .A(n7925), .B(n7926), .Z(n7924) );
  XOR U11521 ( .A(DB[3703]), .B(DB[3688]), .Z(n7926) );
  AND U11522 ( .A(n42), .B(n7927), .Z(n7925) );
  XOR U11523 ( .A(n7928), .B(n7929), .Z(n7927) );
  XOR U11524 ( .A(DB[3688]), .B(DB[3673]), .Z(n7929) );
  AND U11525 ( .A(n46), .B(n7930), .Z(n7928) );
  XOR U11526 ( .A(n7931), .B(n7932), .Z(n7930) );
  XOR U11527 ( .A(DB[3673]), .B(DB[3658]), .Z(n7932) );
  AND U11528 ( .A(n50), .B(n7933), .Z(n7931) );
  XOR U11529 ( .A(n7934), .B(n7935), .Z(n7933) );
  XOR U11530 ( .A(DB[3658]), .B(DB[3643]), .Z(n7935) );
  AND U11531 ( .A(n54), .B(n7936), .Z(n7934) );
  XOR U11532 ( .A(n7937), .B(n7938), .Z(n7936) );
  XOR U11533 ( .A(DB[3643]), .B(DB[3628]), .Z(n7938) );
  AND U11534 ( .A(n58), .B(n7939), .Z(n7937) );
  XOR U11535 ( .A(n7940), .B(n7941), .Z(n7939) );
  XOR U11536 ( .A(DB[3628]), .B(DB[3613]), .Z(n7941) );
  AND U11537 ( .A(n62), .B(n7942), .Z(n7940) );
  XOR U11538 ( .A(n7943), .B(n7944), .Z(n7942) );
  XOR U11539 ( .A(DB[3613]), .B(DB[3598]), .Z(n7944) );
  AND U11540 ( .A(n66), .B(n7945), .Z(n7943) );
  XOR U11541 ( .A(n7946), .B(n7947), .Z(n7945) );
  XOR U11542 ( .A(DB[3598]), .B(DB[3583]), .Z(n7947) );
  AND U11543 ( .A(n70), .B(n7948), .Z(n7946) );
  XOR U11544 ( .A(n7949), .B(n7950), .Z(n7948) );
  XOR U11545 ( .A(DB[3583]), .B(DB[3568]), .Z(n7950) );
  AND U11546 ( .A(n74), .B(n7951), .Z(n7949) );
  XOR U11547 ( .A(n7952), .B(n7953), .Z(n7951) );
  XOR U11548 ( .A(DB[3568]), .B(DB[3553]), .Z(n7953) );
  AND U11549 ( .A(n78), .B(n7954), .Z(n7952) );
  XOR U11550 ( .A(n7955), .B(n7956), .Z(n7954) );
  XOR U11551 ( .A(DB[3553]), .B(DB[3538]), .Z(n7956) );
  AND U11552 ( .A(n82), .B(n7957), .Z(n7955) );
  XOR U11553 ( .A(n7958), .B(n7959), .Z(n7957) );
  XOR U11554 ( .A(DB[3538]), .B(DB[3523]), .Z(n7959) );
  AND U11555 ( .A(n86), .B(n7960), .Z(n7958) );
  XOR U11556 ( .A(n7961), .B(n7962), .Z(n7960) );
  XOR U11557 ( .A(DB[3523]), .B(DB[3508]), .Z(n7962) );
  AND U11558 ( .A(n90), .B(n7963), .Z(n7961) );
  XOR U11559 ( .A(n7964), .B(n7965), .Z(n7963) );
  XOR U11560 ( .A(DB[3508]), .B(DB[3493]), .Z(n7965) );
  AND U11561 ( .A(n94), .B(n7966), .Z(n7964) );
  XOR U11562 ( .A(n7967), .B(n7968), .Z(n7966) );
  XOR U11563 ( .A(DB[3493]), .B(DB[3478]), .Z(n7968) );
  AND U11564 ( .A(n98), .B(n7969), .Z(n7967) );
  XOR U11565 ( .A(n7970), .B(n7971), .Z(n7969) );
  XOR U11566 ( .A(DB[3478]), .B(DB[3463]), .Z(n7971) );
  AND U11567 ( .A(n102), .B(n7972), .Z(n7970) );
  XOR U11568 ( .A(n7973), .B(n7974), .Z(n7972) );
  XOR U11569 ( .A(DB[3463]), .B(DB[3448]), .Z(n7974) );
  AND U11570 ( .A(n106), .B(n7975), .Z(n7973) );
  XOR U11571 ( .A(n7976), .B(n7977), .Z(n7975) );
  XOR U11572 ( .A(DB[3448]), .B(DB[3433]), .Z(n7977) );
  AND U11573 ( .A(n110), .B(n7978), .Z(n7976) );
  XOR U11574 ( .A(n7979), .B(n7980), .Z(n7978) );
  XOR U11575 ( .A(DB[3433]), .B(DB[3418]), .Z(n7980) );
  AND U11576 ( .A(n114), .B(n7981), .Z(n7979) );
  XOR U11577 ( .A(n7982), .B(n7983), .Z(n7981) );
  XOR U11578 ( .A(DB[3418]), .B(DB[3403]), .Z(n7983) );
  AND U11579 ( .A(n118), .B(n7984), .Z(n7982) );
  XOR U11580 ( .A(n7985), .B(n7986), .Z(n7984) );
  XOR U11581 ( .A(DB[3403]), .B(DB[3388]), .Z(n7986) );
  AND U11582 ( .A(n122), .B(n7987), .Z(n7985) );
  XOR U11583 ( .A(n7988), .B(n7989), .Z(n7987) );
  XOR U11584 ( .A(DB[3388]), .B(DB[3373]), .Z(n7989) );
  AND U11585 ( .A(n126), .B(n7990), .Z(n7988) );
  XOR U11586 ( .A(n7991), .B(n7992), .Z(n7990) );
  XOR U11587 ( .A(DB[3373]), .B(DB[3358]), .Z(n7992) );
  AND U11588 ( .A(n130), .B(n7993), .Z(n7991) );
  XOR U11589 ( .A(n7994), .B(n7995), .Z(n7993) );
  XOR U11590 ( .A(DB[3358]), .B(DB[3343]), .Z(n7995) );
  AND U11591 ( .A(n134), .B(n7996), .Z(n7994) );
  XOR U11592 ( .A(n7997), .B(n7998), .Z(n7996) );
  XOR U11593 ( .A(DB[3343]), .B(DB[3328]), .Z(n7998) );
  AND U11594 ( .A(n138), .B(n7999), .Z(n7997) );
  XOR U11595 ( .A(n8000), .B(n8001), .Z(n7999) );
  XOR U11596 ( .A(DB[3328]), .B(DB[3313]), .Z(n8001) );
  AND U11597 ( .A(n142), .B(n8002), .Z(n8000) );
  XOR U11598 ( .A(n8003), .B(n8004), .Z(n8002) );
  XOR U11599 ( .A(DB[3313]), .B(DB[3298]), .Z(n8004) );
  AND U11600 ( .A(n146), .B(n8005), .Z(n8003) );
  XOR U11601 ( .A(n8006), .B(n8007), .Z(n8005) );
  XOR U11602 ( .A(DB[3298]), .B(DB[3283]), .Z(n8007) );
  AND U11603 ( .A(n150), .B(n8008), .Z(n8006) );
  XOR U11604 ( .A(n8009), .B(n8010), .Z(n8008) );
  XOR U11605 ( .A(DB[3283]), .B(DB[3268]), .Z(n8010) );
  AND U11606 ( .A(n154), .B(n8011), .Z(n8009) );
  XOR U11607 ( .A(n8012), .B(n8013), .Z(n8011) );
  XOR U11608 ( .A(DB[3268]), .B(DB[3253]), .Z(n8013) );
  AND U11609 ( .A(n158), .B(n8014), .Z(n8012) );
  XOR U11610 ( .A(n8015), .B(n8016), .Z(n8014) );
  XOR U11611 ( .A(DB[3253]), .B(DB[3238]), .Z(n8016) );
  AND U11612 ( .A(n162), .B(n8017), .Z(n8015) );
  XOR U11613 ( .A(n8018), .B(n8019), .Z(n8017) );
  XOR U11614 ( .A(DB[3238]), .B(DB[3223]), .Z(n8019) );
  AND U11615 ( .A(n166), .B(n8020), .Z(n8018) );
  XOR U11616 ( .A(n8021), .B(n8022), .Z(n8020) );
  XOR U11617 ( .A(DB[3223]), .B(DB[3208]), .Z(n8022) );
  AND U11618 ( .A(n170), .B(n8023), .Z(n8021) );
  XOR U11619 ( .A(n8024), .B(n8025), .Z(n8023) );
  XOR U11620 ( .A(DB[3208]), .B(DB[3193]), .Z(n8025) );
  AND U11621 ( .A(n174), .B(n8026), .Z(n8024) );
  XOR U11622 ( .A(n8027), .B(n8028), .Z(n8026) );
  XOR U11623 ( .A(DB[3193]), .B(DB[3178]), .Z(n8028) );
  AND U11624 ( .A(n178), .B(n8029), .Z(n8027) );
  XOR U11625 ( .A(n8030), .B(n8031), .Z(n8029) );
  XOR U11626 ( .A(DB[3178]), .B(DB[3163]), .Z(n8031) );
  AND U11627 ( .A(n182), .B(n8032), .Z(n8030) );
  XOR U11628 ( .A(n8033), .B(n8034), .Z(n8032) );
  XOR U11629 ( .A(DB[3163]), .B(DB[3148]), .Z(n8034) );
  AND U11630 ( .A(n186), .B(n8035), .Z(n8033) );
  XOR U11631 ( .A(n8036), .B(n8037), .Z(n8035) );
  XOR U11632 ( .A(DB[3148]), .B(DB[3133]), .Z(n8037) );
  AND U11633 ( .A(n190), .B(n8038), .Z(n8036) );
  XOR U11634 ( .A(n8039), .B(n8040), .Z(n8038) );
  XOR U11635 ( .A(DB[3133]), .B(DB[3118]), .Z(n8040) );
  AND U11636 ( .A(n194), .B(n8041), .Z(n8039) );
  XOR U11637 ( .A(n8042), .B(n8043), .Z(n8041) );
  XOR U11638 ( .A(DB[3118]), .B(DB[3103]), .Z(n8043) );
  AND U11639 ( .A(n198), .B(n8044), .Z(n8042) );
  XOR U11640 ( .A(n8045), .B(n8046), .Z(n8044) );
  XOR U11641 ( .A(DB[3103]), .B(DB[3088]), .Z(n8046) );
  AND U11642 ( .A(n202), .B(n8047), .Z(n8045) );
  XOR U11643 ( .A(n8048), .B(n8049), .Z(n8047) );
  XOR U11644 ( .A(DB[3088]), .B(DB[3073]), .Z(n8049) );
  AND U11645 ( .A(n206), .B(n8050), .Z(n8048) );
  XOR U11646 ( .A(n8051), .B(n8052), .Z(n8050) );
  XOR U11647 ( .A(DB[3073]), .B(DB[3058]), .Z(n8052) );
  AND U11648 ( .A(n210), .B(n8053), .Z(n8051) );
  XOR U11649 ( .A(n8054), .B(n8055), .Z(n8053) );
  XOR U11650 ( .A(DB[3058]), .B(DB[3043]), .Z(n8055) );
  AND U11651 ( .A(n214), .B(n8056), .Z(n8054) );
  XOR U11652 ( .A(n8057), .B(n8058), .Z(n8056) );
  XOR U11653 ( .A(DB[3043]), .B(DB[3028]), .Z(n8058) );
  AND U11654 ( .A(n218), .B(n8059), .Z(n8057) );
  XOR U11655 ( .A(n8060), .B(n8061), .Z(n8059) );
  XOR U11656 ( .A(DB[3028]), .B(DB[3013]), .Z(n8061) );
  AND U11657 ( .A(n222), .B(n8062), .Z(n8060) );
  XOR U11658 ( .A(n8063), .B(n8064), .Z(n8062) );
  XOR U11659 ( .A(DB[3013]), .B(DB[2998]), .Z(n8064) );
  AND U11660 ( .A(n226), .B(n8065), .Z(n8063) );
  XOR U11661 ( .A(n8066), .B(n8067), .Z(n8065) );
  XOR U11662 ( .A(DB[2998]), .B(DB[2983]), .Z(n8067) );
  AND U11663 ( .A(n230), .B(n8068), .Z(n8066) );
  XOR U11664 ( .A(n8069), .B(n8070), .Z(n8068) );
  XOR U11665 ( .A(DB[2983]), .B(DB[2968]), .Z(n8070) );
  AND U11666 ( .A(n234), .B(n8071), .Z(n8069) );
  XOR U11667 ( .A(n8072), .B(n8073), .Z(n8071) );
  XOR U11668 ( .A(DB[2968]), .B(DB[2953]), .Z(n8073) );
  AND U11669 ( .A(n238), .B(n8074), .Z(n8072) );
  XOR U11670 ( .A(n8075), .B(n8076), .Z(n8074) );
  XOR U11671 ( .A(DB[2953]), .B(DB[2938]), .Z(n8076) );
  AND U11672 ( .A(n242), .B(n8077), .Z(n8075) );
  XOR U11673 ( .A(n8078), .B(n8079), .Z(n8077) );
  XOR U11674 ( .A(DB[2938]), .B(DB[2923]), .Z(n8079) );
  AND U11675 ( .A(n246), .B(n8080), .Z(n8078) );
  XOR U11676 ( .A(n8081), .B(n8082), .Z(n8080) );
  XOR U11677 ( .A(DB[2923]), .B(DB[2908]), .Z(n8082) );
  AND U11678 ( .A(n250), .B(n8083), .Z(n8081) );
  XOR U11679 ( .A(n8084), .B(n8085), .Z(n8083) );
  XOR U11680 ( .A(DB[2908]), .B(DB[2893]), .Z(n8085) );
  AND U11681 ( .A(n254), .B(n8086), .Z(n8084) );
  XOR U11682 ( .A(n8087), .B(n8088), .Z(n8086) );
  XOR U11683 ( .A(DB[2893]), .B(DB[2878]), .Z(n8088) );
  AND U11684 ( .A(n258), .B(n8089), .Z(n8087) );
  XOR U11685 ( .A(n8090), .B(n8091), .Z(n8089) );
  XOR U11686 ( .A(DB[2878]), .B(DB[2863]), .Z(n8091) );
  AND U11687 ( .A(n262), .B(n8092), .Z(n8090) );
  XOR U11688 ( .A(n8093), .B(n8094), .Z(n8092) );
  XOR U11689 ( .A(DB[2863]), .B(DB[2848]), .Z(n8094) );
  AND U11690 ( .A(n266), .B(n8095), .Z(n8093) );
  XOR U11691 ( .A(n8096), .B(n8097), .Z(n8095) );
  XOR U11692 ( .A(DB[2848]), .B(DB[2833]), .Z(n8097) );
  AND U11693 ( .A(n270), .B(n8098), .Z(n8096) );
  XOR U11694 ( .A(n8099), .B(n8100), .Z(n8098) );
  XOR U11695 ( .A(DB[2833]), .B(DB[2818]), .Z(n8100) );
  AND U11696 ( .A(n274), .B(n8101), .Z(n8099) );
  XOR U11697 ( .A(n8102), .B(n8103), .Z(n8101) );
  XOR U11698 ( .A(DB[2818]), .B(DB[2803]), .Z(n8103) );
  AND U11699 ( .A(n278), .B(n8104), .Z(n8102) );
  XOR U11700 ( .A(n8105), .B(n8106), .Z(n8104) );
  XOR U11701 ( .A(DB[2803]), .B(DB[2788]), .Z(n8106) );
  AND U11702 ( .A(n282), .B(n8107), .Z(n8105) );
  XOR U11703 ( .A(n8108), .B(n8109), .Z(n8107) );
  XOR U11704 ( .A(DB[2788]), .B(DB[2773]), .Z(n8109) );
  AND U11705 ( .A(n286), .B(n8110), .Z(n8108) );
  XOR U11706 ( .A(n8111), .B(n8112), .Z(n8110) );
  XOR U11707 ( .A(DB[2773]), .B(DB[2758]), .Z(n8112) );
  AND U11708 ( .A(n290), .B(n8113), .Z(n8111) );
  XOR U11709 ( .A(n8114), .B(n8115), .Z(n8113) );
  XOR U11710 ( .A(DB[2758]), .B(DB[2743]), .Z(n8115) );
  AND U11711 ( .A(n294), .B(n8116), .Z(n8114) );
  XOR U11712 ( .A(n8117), .B(n8118), .Z(n8116) );
  XOR U11713 ( .A(DB[2743]), .B(DB[2728]), .Z(n8118) );
  AND U11714 ( .A(n298), .B(n8119), .Z(n8117) );
  XOR U11715 ( .A(n8120), .B(n8121), .Z(n8119) );
  XOR U11716 ( .A(DB[2728]), .B(DB[2713]), .Z(n8121) );
  AND U11717 ( .A(n302), .B(n8122), .Z(n8120) );
  XOR U11718 ( .A(n8123), .B(n8124), .Z(n8122) );
  XOR U11719 ( .A(DB[2713]), .B(DB[2698]), .Z(n8124) );
  AND U11720 ( .A(n306), .B(n8125), .Z(n8123) );
  XOR U11721 ( .A(n8126), .B(n8127), .Z(n8125) );
  XOR U11722 ( .A(DB[2698]), .B(DB[2683]), .Z(n8127) );
  AND U11723 ( .A(n310), .B(n8128), .Z(n8126) );
  XOR U11724 ( .A(n8129), .B(n8130), .Z(n8128) );
  XOR U11725 ( .A(DB[2683]), .B(DB[2668]), .Z(n8130) );
  AND U11726 ( .A(n314), .B(n8131), .Z(n8129) );
  XOR U11727 ( .A(n8132), .B(n8133), .Z(n8131) );
  XOR U11728 ( .A(DB[2668]), .B(DB[2653]), .Z(n8133) );
  AND U11729 ( .A(n318), .B(n8134), .Z(n8132) );
  XOR U11730 ( .A(n8135), .B(n8136), .Z(n8134) );
  XOR U11731 ( .A(DB[2653]), .B(DB[2638]), .Z(n8136) );
  AND U11732 ( .A(n322), .B(n8137), .Z(n8135) );
  XOR U11733 ( .A(n8138), .B(n8139), .Z(n8137) );
  XOR U11734 ( .A(DB[2638]), .B(DB[2623]), .Z(n8139) );
  AND U11735 ( .A(n326), .B(n8140), .Z(n8138) );
  XOR U11736 ( .A(n8141), .B(n8142), .Z(n8140) );
  XOR U11737 ( .A(DB[2623]), .B(DB[2608]), .Z(n8142) );
  AND U11738 ( .A(n330), .B(n8143), .Z(n8141) );
  XOR U11739 ( .A(n8144), .B(n8145), .Z(n8143) );
  XOR U11740 ( .A(DB[2608]), .B(DB[2593]), .Z(n8145) );
  AND U11741 ( .A(n334), .B(n8146), .Z(n8144) );
  XOR U11742 ( .A(n8147), .B(n8148), .Z(n8146) );
  XOR U11743 ( .A(DB[2593]), .B(DB[2578]), .Z(n8148) );
  AND U11744 ( .A(n338), .B(n8149), .Z(n8147) );
  XOR U11745 ( .A(n8150), .B(n8151), .Z(n8149) );
  XOR U11746 ( .A(DB[2578]), .B(DB[2563]), .Z(n8151) );
  AND U11747 ( .A(n342), .B(n8152), .Z(n8150) );
  XOR U11748 ( .A(n8153), .B(n8154), .Z(n8152) );
  XOR U11749 ( .A(DB[2563]), .B(DB[2548]), .Z(n8154) );
  AND U11750 ( .A(n346), .B(n8155), .Z(n8153) );
  XOR U11751 ( .A(n8156), .B(n8157), .Z(n8155) );
  XOR U11752 ( .A(DB[2548]), .B(DB[2533]), .Z(n8157) );
  AND U11753 ( .A(n350), .B(n8158), .Z(n8156) );
  XOR U11754 ( .A(n8159), .B(n8160), .Z(n8158) );
  XOR U11755 ( .A(DB[2533]), .B(DB[2518]), .Z(n8160) );
  AND U11756 ( .A(n354), .B(n8161), .Z(n8159) );
  XOR U11757 ( .A(n8162), .B(n8163), .Z(n8161) );
  XOR U11758 ( .A(DB[2518]), .B(DB[2503]), .Z(n8163) );
  AND U11759 ( .A(n358), .B(n8164), .Z(n8162) );
  XOR U11760 ( .A(n8165), .B(n8166), .Z(n8164) );
  XOR U11761 ( .A(DB[2503]), .B(DB[2488]), .Z(n8166) );
  AND U11762 ( .A(n362), .B(n8167), .Z(n8165) );
  XOR U11763 ( .A(n8168), .B(n8169), .Z(n8167) );
  XOR U11764 ( .A(DB[2488]), .B(DB[2473]), .Z(n8169) );
  AND U11765 ( .A(n366), .B(n8170), .Z(n8168) );
  XOR U11766 ( .A(n8171), .B(n8172), .Z(n8170) );
  XOR U11767 ( .A(DB[2473]), .B(DB[2458]), .Z(n8172) );
  AND U11768 ( .A(n370), .B(n8173), .Z(n8171) );
  XOR U11769 ( .A(n8174), .B(n8175), .Z(n8173) );
  XOR U11770 ( .A(DB[2458]), .B(DB[2443]), .Z(n8175) );
  AND U11771 ( .A(n374), .B(n8176), .Z(n8174) );
  XOR U11772 ( .A(n8177), .B(n8178), .Z(n8176) );
  XOR U11773 ( .A(DB[2443]), .B(DB[2428]), .Z(n8178) );
  AND U11774 ( .A(n378), .B(n8179), .Z(n8177) );
  XOR U11775 ( .A(n8180), .B(n8181), .Z(n8179) );
  XOR U11776 ( .A(DB[2428]), .B(DB[2413]), .Z(n8181) );
  AND U11777 ( .A(n382), .B(n8182), .Z(n8180) );
  XOR U11778 ( .A(n8183), .B(n8184), .Z(n8182) );
  XOR U11779 ( .A(DB[2413]), .B(DB[2398]), .Z(n8184) );
  AND U11780 ( .A(n386), .B(n8185), .Z(n8183) );
  XOR U11781 ( .A(n8186), .B(n8187), .Z(n8185) );
  XOR U11782 ( .A(DB[2398]), .B(DB[2383]), .Z(n8187) );
  AND U11783 ( .A(n390), .B(n8188), .Z(n8186) );
  XOR U11784 ( .A(n8189), .B(n8190), .Z(n8188) );
  XOR U11785 ( .A(DB[2383]), .B(DB[2368]), .Z(n8190) );
  AND U11786 ( .A(n394), .B(n8191), .Z(n8189) );
  XOR U11787 ( .A(n8192), .B(n8193), .Z(n8191) );
  XOR U11788 ( .A(DB[2368]), .B(DB[2353]), .Z(n8193) );
  AND U11789 ( .A(n398), .B(n8194), .Z(n8192) );
  XOR U11790 ( .A(n8195), .B(n8196), .Z(n8194) );
  XOR U11791 ( .A(DB[2353]), .B(DB[2338]), .Z(n8196) );
  AND U11792 ( .A(n402), .B(n8197), .Z(n8195) );
  XOR U11793 ( .A(n8198), .B(n8199), .Z(n8197) );
  XOR U11794 ( .A(DB[2338]), .B(DB[2323]), .Z(n8199) );
  AND U11795 ( .A(n406), .B(n8200), .Z(n8198) );
  XOR U11796 ( .A(n8201), .B(n8202), .Z(n8200) );
  XOR U11797 ( .A(DB[2323]), .B(DB[2308]), .Z(n8202) );
  AND U11798 ( .A(n410), .B(n8203), .Z(n8201) );
  XOR U11799 ( .A(n8204), .B(n8205), .Z(n8203) );
  XOR U11800 ( .A(DB[2308]), .B(DB[2293]), .Z(n8205) );
  AND U11801 ( .A(n414), .B(n8206), .Z(n8204) );
  XOR U11802 ( .A(n8207), .B(n8208), .Z(n8206) );
  XOR U11803 ( .A(DB[2293]), .B(DB[2278]), .Z(n8208) );
  AND U11804 ( .A(n418), .B(n8209), .Z(n8207) );
  XOR U11805 ( .A(n8210), .B(n8211), .Z(n8209) );
  XOR U11806 ( .A(DB[2278]), .B(DB[2263]), .Z(n8211) );
  AND U11807 ( .A(n422), .B(n8212), .Z(n8210) );
  XOR U11808 ( .A(n8213), .B(n8214), .Z(n8212) );
  XOR U11809 ( .A(DB[2263]), .B(DB[2248]), .Z(n8214) );
  AND U11810 ( .A(n426), .B(n8215), .Z(n8213) );
  XOR U11811 ( .A(n8216), .B(n8217), .Z(n8215) );
  XOR U11812 ( .A(DB[2248]), .B(DB[2233]), .Z(n8217) );
  AND U11813 ( .A(n430), .B(n8218), .Z(n8216) );
  XOR U11814 ( .A(n8219), .B(n8220), .Z(n8218) );
  XOR U11815 ( .A(DB[2233]), .B(DB[2218]), .Z(n8220) );
  AND U11816 ( .A(n434), .B(n8221), .Z(n8219) );
  XOR U11817 ( .A(n8222), .B(n8223), .Z(n8221) );
  XOR U11818 ( .A(DB[2218]), .B(DB[2203]), .Z(n8223) );
  AND U11819 ( .A(n438), .B(n8224), .Z(n8222) );
  XOR U11820 ( .A(n8225), .B(n8226), .Z(n8224) );
  XOR U11821 ( .A(DB[2203]), .B(DB[2188]), .Z(n8226) );
  AND U11822 ( .A(n442), .B(n8227), .Z(n8225) );
  XOR U11823 ( .A(n8228), .B(n8229), .Z(n8227) );
  XOR U11824 ( .A(DB[2188]), .B(DB[2173]), .Z(n8229) );
  AND U11825 ( .A(n446), .B(n8230), .Z(n8228) );
  XOR U11826 ( .A(n8231), .B(n8232), .Z(n8230) );
  XOR U11827 ( .A(DB[2173]), .B(DB[2158]), .Z(n8232) );
  AND U11828 ( .A(n450), .B(n8233), .Z(n8231) );
  XOR U11829 ( .A(n8234), .B(n8235), .Z(n8233) );
  XOR U11830 ( .A(DB[2158]), .B(DB[2143]), .Z(n8235) );
  AND U11831 ( .A(n454), .B(n8236), .Z(n8234) );
  XOR U11832 ( .A(n8237), .B(n8238), .Z(n8236) );
  XOR U11833 ( .A(DB[2143]), .B(DB[2128]), .Z(n8238) );
  AND U11834 ( .A(n458), .B(n8239), .Z(n8237) );
  XOR U11835 ( .A(n8240), .B(n8241), .Z(n8239) );
  XOR U11836 ( .A(DB[2128]), .B(DB[2113]), .Z(n8241) );
  AND U11837 ( .A(n462), .B(n8242), .Z(n8240) );
  XOR U11838 ( .A(n8243), .B(n8244), .Z(n8242) );
  XOR U11839 ( .A(DB[2113]), .B(DB[2098]), .Z(n8244) );
  AND U11840 ( .A(n466), .B(n8245), .Z(n8243) );
  XOR U11841 ( .A(n8246), .B(n8247), .Z(n8245) );
  XOR U11842 ( .A(DB[2098]), .B(DB[2083]), .Z(n8247) );
  AND U11843 ( .A(n470), .B(n8248), .Z(n8246) );
  XOR U11844 ( .A(n8249), .B(n8250), .Z(n8248) );
  XOR U11845 ( .A(DB[2083]), .B(DB[2068]), .Z(n8250) );
  AND U11846 ( .A(n474), .B(n8251), .Z(n8249) );
  XOR U11847 ( .A(n8252), .B(n8253), .Z(n8251) );
  XOR U11848 ( .A(DB[2068]), .B(DB[2053]), .Z(n8253) );
  AND U11849 ( .A(n478), .B(n8254), .Z(n8252) );
  XOR U11850 ( .A(n8255), .B(n8256), .Z(n8254) );
  XOR U11851 ( .A(DB[2053]), .B(DB[2038]), .Z(n8256) );
  AND U11852 ( .A(n482), .B(n8257), .Z(n8255) );
  XOR U11853 ( .A(n8258), .B(n8259), .Z(n8257) );
  XOR U11854 ( .A(DB[2038]), .B(DB[2023]), .Z(n8259) );
  AND U11855 ( .A(n486), .B(n8260), .Z(n8258) );
  XOR U11856 ( .A(n8261), .B(n8262), .Z(n8260) );
  XOR U11857 ( .A(DB[2023]), .B(DB[2008]), .Z(n8262) );
  AND U11858 ( .A(n490), .B(n8263), .Z(n8261) );
  XOR U11859 ( .A(n8264), .B(n8265), .Z(n8263) );
  XOR U11860 ( .A(DB[2008]), .B(DB[1993]), .Z(n8265) );
  AND U11861 ( .A(n494), .B(n8266), .Z(n8264) );
  XOR U11862 ( .A(n8267), .B(n8268), .Z(n8266) );
  XOR U11863 ( .A(DB[1993]), .B(DB[1978]), .Z(n8268) );
  AND U11864 ( .A(n498), .B(n8269), .Z(n8267) );
  XOR U11865 ( .A(n8270), .B(n8271), .Z(n8269) );
  XOR U11866 ( .A(DB[1978]), .B(DB[1963]), .Z(n8271) );
  AND U11867 ( .A(n502), .B(n8272), .Z(n8270) );
  XOR U11868 ( .A(n8273), .B(n8274), .Z(n8272) );
  XOR U11869 ( .A(DB[1963]), .B(DB[1948]), .Z(n8274) );
  AND U11870 ( .A(n506), .B(n8275), .Z(n8273) );
  XOR U11871 ( .A(n8276), .B(n8277), .Z(n8275) );
  XOR U11872 ( .A(DB[1948]), .B(DB[1933]), .Z(n8277) );
  AND U11873 ( .A(n510), .B(n8278), .Z(n8276) );
  XOR U11874 ( .A(n8279), .B(n8280), .Z(n8278) );
  XOR U11875 ( .A(DB[1933]), .B(DB[1918]), .Z(n8280) );
  AND U11876 ( .A(n514), .B(n8281), .Z(n8279) );
  XOR U11877 ( .A(n8282), .B(n8283), .Z(n8281) );
  XOR U11878 ( .A(DB[1918]), .B(DB[1903]), .Z(n8283) );
  AND U11879 ( .A(n518), .B(n8284), .Z(n8282) );
  XOR U11880 ( .A(n8285), .B(n8286), .Z(n8284) );
  XOR U11881 ( .A(DB[1903]), .B(DB[1888]), .Z(n8286) );
  AND U11882 ( .A(n522), .B(n8287), .Z(n8285) );
  XOR U11883 ( .A(n8288), .B(n8289), .Z(n8287) );
  XOR U11884 ( .A(DB[1888]), .B(DB[1873]), .Z(n8289) );
  AND U11885 ( .A(n526), .B(n8290), .Z(n8288) );
  XOR U11886 ( .A(n8291), .B(n8292), .Z(n8290) );
  XOR U11887 ( .A(DB[1873]), .B(DB[1858]), .Z(n8292) );
  AND U11888 ( .A(n530), .B(n8293), .Z(n8291) );
  XOR U11889 ( .A(n8294), .B(n8295), .Z(n8293) );
  XOR U11890 ( .A(DB[1858]), .B(DB[1843]), .Z(n8295) );
  AND U11891 ( .A(n534), .B(n8296), .Z(n8294) );
  XOR U11892 ( .A(n8297), .B(n8298), .Z(n8296) );
  XOR U11893 ( .A(DB[1843]), .B(DB[1828]), .Z(n8298) );
  AND U11894 ( .A(n538), .B(n8299), .Z(n8297) );
  XOR U11895 ( .A(n8300), .B(n8301), .Z(n8299) );
  XOR U11896 ( .A(DB[1828]), .B(DB[1813]), .Z(n8301) );
  AND U11897 ( .A(n542), .B(n8302), .Z(n8300) );
  XOR U11898 ( .A(n8303), .B(n8304), .Z(n8302) );
  XOR U11899 ( .A(DB[1813]), .B(DB[1798]), .Z(n8304) );
  AND U11900 ( .A(n546), .B(n8305), .Z(n8303) );
  XOR U11901 ( .A(n8306), .B(n8307), .Z(n8305) );
  XOR U11902 ( .A(DB[1798]), .B(DB[1783]), .Z(n8307) );
  AND U11903 ( .A(n550), .B(n8308), .Z(n8306) );
  XOR U11904 ( .A(n8309), .B(n8310), .Z(n8308) );
  XOR U11905 ( .A(DB[1783]), .B(DB[1768]), .Z(n8310) );
  AND U11906 ( .A(n554), .B(n8311), .Z(n8309) );
  XOR U11907 ( .A(n8312), .B(n8313), .Z(n8311) );
  XOR U11908 ( .A(DB[1768]), .B(DB[1753]), .Z(n8313) );
  AND U11909 ( .A(n558), .B(n8314), .Z(n8312) );
  XOR U11910 ( .A(n8315), .B(n8316), .Z(n8314) );
  XOR U11911 ( .A(DB[1753]), .B(DB[1738]), .Z(n8316) );
  AND U11912 ( .A(n562), .B(n8317), .Z(n8315) );
  XOR U11913 ( .A(n8318), .B(n8319), .Z(n8317) );
  XOR U11914 ( .A(DB[1738]), .B(DB[1723]), .Z(n8319) );
  AND U11915 ( .A(n566), .B(n8320), .Z(n8318) );
  XOR U11916 ( .A(n8321), .B(n8322), .Z(n8320) );
  XOR U11917 ( .A(DB[1723]), .B(DB[1708]), .Z(n8322) );
  AND U11918 ( .A(n570), .B(n8323), .Z(n8321) );
  XOR U11919 ( .A(n8324), .B(n8325), .Z(n8323) );
  XOR U11920 ( .A(DB[1708]), .B(DB[1693]), .Z(n8325) );
  AND U11921 ( .A(n574), .B(n8326), .Z(n8324) );
  XOR U11922 ( .A(n8327), .B(n8328), .Z(n8326) );
  XOR U11923 ( .A(DB[1693]), .B(DB[1678]), .Z(n8328) );
  AND U11924 ( .A(n578), .B(n8329), .Z(n8327) );
  XOR U11925 ( .A(n8330), .B(n8331), .Z(n8329) );
  XOR U11926 ( .A(DB[1678]), .B(DB[1663]), .Z(n8331) );
  AND U11927 ( .A(n582), .B(n8332), .Z(n8330) );
  XOR U11928 ( .A(n8333), .B(n8334), .Z(n8332) );
  XOR U11929 ( .A(DB[1663]), .B(DB[1648]), .Z(n8334) );
  AND U11930 ( .A(n586), .B(n8335), .Z(n8333) );
  XOR U11931 ( .A(n8336), .B(n8337), .Z(n8335) );
  XOR U11932 ( .A(DB[1648]), .B(DB[1633]), .Z(n8337) );
  AND U11933 ( .A(n590), .B(n8338), .Z(n8336) );
  XOR U11934 ( .A(n8339), .B(n8340), .Z(n8338) );
  XOR U11935 ( .A(DB[1633]), .B(DB[1618]), .Z(n8340) );
  AND U11936 ( .A(n594), .B(n8341), .Z(n8339) );
  XOR U11937 ( .A(n8342), .B(n8343), .Z(n8341) );
  XOR U11938 ( .A(DB[1618]), .B(DB[1603]), .Z(n8343) );
  AND U11939 ( .A(n598), .B(n8344), .Z(n8342) );
  XOR U11940 ( .A(n8345), .B(n8346), .Z(n8344) );
  XOR U11941 ( .A(DB[1603]), .B(DB[1588]), .Z(n8346) );
  AND U11942 ( .A(n602), .B(n8347), .Z(n8345) );
  XOR U11943 ( .A(n8348), .B(n8349), .Z(n8347) );
  XOR U11944 ( .A(DB[1588]), .B(DB[1573]), .Z(n8349) );
  AND U11945 ( .A(n606), .B(n8350), .Z(n8348) );
  XOR U11946 ( .A(n8351), .B(n8352), .Z(n8350) );
  XOR U11947 ( .A(DB[1573]), .B(DB[1558]), .Z(n8352) );
  AND U11948 ( .A(n610), .B(n8353), .Z(n8351) );
  XOR U11949 ( .A(n8354), .B(n8355), .Z(n8353) );
  XOR U11950 ( .A(DB[1558]), .B(DB[1543]), .Z(n8355) );
  AND U11951 ( .A(n614), .B(n8356), .Z(n8354) );
  XOR U11952 ( .A(n8357), .B(n8358), .Z(n8356) );
  XOR U11953 ( .A(DB[1543]), .B(DB[1528]), .Z(n8358) );
  AND U11954 ( .A(n618), .B(n8359), .Z(n8357) );
  XOR U11955 ( .A(n8360), .B(n8361), .Z(n8359) );
  XOR U11956 ( .A(DB[1528]), .B(DB[1513]), .Z(n8361) );
  AND U11957 ( .A(n622), .B(n8362), .Z(n8360) );
  XOR U11958 ( .A(n8363), .B(n8364), .Z(n8362) );
  XOR U11959 ( .A(DB[1513]), .B(DB[1498]), .Z(n8364) );
  AND U11960 ( .A(n626), .B(n8365), .Z(n8363) );
  XOR U11961 ( .A(n8366), .B(n8367), .Z(n8365) );
  XOR U11962 ( .A(DB[1498]), .B(DB[1483]), .Z(n8367) );
  AND U11963 ( .A(n630), .B(n8368), .Z(n8366) );
  XOR U11964 ( .A(n8369), .B(n8370), .Z(n8368) );
  XOR U11965 ( .A(DB[1483]), .B(DB[1468]), .Z(n8370) );
  AND U11966 ( .A(n634), .B(n8371), .Z(n8369) );
  XOR U11967 ( .A(n8372), .B(n8373), .Z(n8371) );
  XOR U11968 ( .A(DB[1468]), .B(DB[1453]), .Z(n8373) );
  AND U11969 ( .A(n638), .B(n8374), .Z(n8372) );
  XOR U11970 ( .A(n8375), .B(n8376), .Z(n8374) );
  XOR U11971 ( .A(DB[1453]), .B(DB[1438]), .Z(n8376) );
  AND U11972 ( .A(n642), .B(n8377), .Z(n8375) );
  XOR U11973 ( .A(n8378), .B(n8379), .Z(n8377) );
  XOR U11974 ( .A(DB[1438]), .B(DB[1423]), .Z(n8379) );
  AND U11975 ( .A(n646), .B(n8380), .Z(n8378) );
  XOR U11976 ( .A(n8381), .B(n8382), .Z(n8380) );
  XOR U11977 ( .A(DB[1423]), .B(DB[1408]), .Z(n8382) );
  AND U11978 ( .A(n650), .B(n8383), .Z(n8381) );
  XOR U11979 ( .A(n8384), .B(n8385), .Z(n8383) );
  XOR U11980 ( .A(DB[1408]), .B(DB[1393]), .Z(n8385) );
  AND U11981 ( .A(n654), .B(n8386), .Z(n8384) );
  XOR U11982 ( .A(n8387), .B(n8388), .Z(n8386) );
  XOR U11983 ( .A(DB[1393]), .B(DB[1378]), .Z(n8388) );
  AND U11984 ( .A(n658), .B(n8389), .Z(n8387) );
  XOR U11985 ( .A(n8390), .B(n8391), .Z(n8389) );
  XOR U11986 ( .A(DB[1378]), .B(DB[1363]), .Z(n8391) );
  AND U11987 ( .A(n662), .B(n8392), .Z(n8390) );
  XOR U11988 ( .A(n8393), .B(n8394), .Z(n8392) );
  XOR U11989 ( .A(DB[1363]), .B(DB[1348]), .Z(n8394) );
  AND U11990 ( .A(n666), .B(n8395), .Z(n8393) );
  XOR U11991 ( .A(n8396), .B(n8397), .Z(n8395) );
  XOR U11992 ( .A(DB[1348]), .B(DB[1333]), .Z(n8397) );
  AND U11993 ( .A(n670), .B(n8398), .Z(n8396) );
  XOR U11994 ( .A(n8399), .B(n8400), .Z(n8398) );
  XOR U11995 ( .A(DB[1333]), .B(DB[1318]), .Z(n8400) );
  AND U11996 ( .A(n674), .B(n8401), .Z(n8399) );
  XOR U11997 ( .A(n8402), .B(n8403), .Z(n8401) );
  XOR U11998 ( .A(DB[1318]), .B(DB[1303]), .Z(n8403) );
  AND U11999 ( .A(n678), .B(n8404), .Z(n8402) );
  XOR U12000 ( .A(n8405), .B(n8406), .Z(n8404) );
  XOR U12001 ( .A(DB[1303]), .B(DB[1288]), .Z(n8406) );
  AND U12002 ( .A(n682), .B(n8407), .Z(n8405) );
  XOR U12003 ( .A(n8408), .B(n8409), .Z(n8407) );
  XOR U12004 ( .A(DB[1288]), .B(DB[1273]), .Z(n8409) );
  AND U12005 ( .A(n686), .B(n8410), .Z(n8408) );
  XOR U12006 ( .A(n8411), .B(n8412), .Z(n8410) );
  XOR U12007 ( .A(DB[1273]), .B(DB[1258]), .Z(n8412) );
  AND U12008 ( .A(n690), .B(n8413), .Z(n8411) );
  XOR U12009 ( .A(n8414), .B(n8415), .Z(n8413) );
  XOR U12010 ( .A(DB[1258]), .B(DB[1243]), .Z(n8415) );
  AND U12011 ( .A(n694), .B(n8416), .Z(n8414) );
  XOR U12012 ( .A(n8417), .B(n8418), .Z(n8416) );
  XOR U12013 ( .A(DB[1243]), .B(DB[1228]), .Z(n8418) );
  AND U12014 ( .A(n698), .B(n8419), .Z(n8417) );
  XOR U12015 ( .A(n8420), .B(n8421), .Z(n8419) );
  XOR U12016 ( .A(DB[1228]), .B(DB[1213]), .Z(n8421) );
  AND U12017 ( .A(n702), .B(n8422), .Z(n8420) );
  XOR U12018 ( .A(n8423), .B(n8424), .Z(n8422) );
  XOR U12019 ( .A(DB[1213]), .B(DB[1198]), .Z(n8424) );
  AND U12020 ( .A(n706), .B(n8425), .Z(n8423) );
  XOR U12021 ( .A(n8426), .B(n8427), .Z(n8425) );
  XOR U12022 ( .A(DB[1198]), .B(DB[1183]), .Z(n8427) );
  AND U12023 ( .A(n710), .B(n8428), .Z(n8426) );
  XOR U12024 ( .A(n8429), .B(n8430), .Z(n8428) );
  XOR U12025 ( .A(DB[1183]), .B(DB[1168]), .Z(n8430) );
  AND U12026 ( .A(n714), .B(n8431), .Z(n8429) );
  XOR U12027 ( .A(n8432), .B(n8433), .Z(n8431) );
  XOR U12028 ( .A(DB[1168]), .B(DB[1153]), .Z(n8433) );
  AND U12029 ( .A(n718), .B(n8434), .Z(n8432) );
  XOR U12030 ( .A(n8435), .B(n8436), .Z(n8434) );
  XOR U12031 ( .A(DB[1153]), .B(DB[1138]), .Z(n8436) );
  AND U12032 ( .A(n722), .B(n8437), .Z(n8435) );
  XOR U12033 ( .A(n8438), .B(n8439), .Z(n8437) );
  XOR U12034 ( .A(DB[1138]), .B(DB[1123]), .Z(n8439) );
  AND U12035 ( .A(n726), .B(n8440), .Z(n8438) );
  XOR U12036 ( .A(n8441), .B(n8442), .Z(n8440) );
  XOR U12037 ( .A(DB[1123]), .B(DB[1108]), .Z(n8442) );
  AND U12038 ( .A(n730), .B(n8443), .Z(n8441) );
  XOR U12039 ( .A(n8444), .B(n8445), .Z(n8443) );
  XOR U12040 ( .A(DB[1108]), .B(DB[1093]), .Z(n8445) );
  AND U12041 ( .A(n734), .B(n8446), .Z(n8444) );
  XOR U12042 ( .A(n8447), .B(n8448), .Z(n8446) );
  XOR U12043 ( .A(DB[1093]), .B(DB[1078]), .Z(n8448) );
  AND U12044 ( .A(n738), .B(n8449), .Z(n8447) );
  XOR U12045 ( .A(n8450), .B(n8451), .Z(n8449) );
  XOR U12046 ( .A(DB[1078]), .B(DB[1063]), .Z(n8451) );
  AND U12047 ( .A(n742), .B(n8452), .Z(n8450) );
  XOR U12048 ( .A(n8453), .B(n8454), .Z(n8452) );
  XOR U12049 ( .A(DB[1063]), .B(DB[1048]), .Z(n8454) );
  AND U12050 ( .A(n746), .B(n8455), .Z(n8453) );
  XOR U12051 ( .A(n8456), .B(n8457), .Z(n8455) );
  XOR U12052 ( .A(DB[1048]), .B(DB[1033]), .Z(n8457) );
  AND U12053 ( .A(n750), .B(n8458), .Z(n8456) );
  XOR U12054 ( .A(n8459), .B(n8460), .Z(n8458) );
  XOR U12055 ( .A(DB[1033]), .B(DB[1018]), .Z(n8460) );
  AND U12056 ( .A(n754), .B(n8461), .Z(n8459) );
  XOR U12057 ( .A(n8462), .B(n8463), .Z(n8461) );
  XOR U12058 ( .A(DB[1018]), .B(DB[1003]), .Z(n8463) );
  AND U12059 ( .A(n758), .B(n8464), .Z(n8462) );
  XOR U12060 ( .A(n8465), .B(n8466), .Z(n8464) );
  XOR U12061 ( .A(DB[988]), .B(DB[1003]), .Z(n8466) );
  AND U12062 ( .A(n762), .B(n8467), .Z(n8465) );
  XOR U12063 ( .A(n8468), .B(n8469), .Z(n8467) );
  XOR U12064 ( .A(DB[988]), .B(DB[973]), .Z(n8469) );
  AND U12065 ( .A(n766), .B(n8470), .Z(n8468) );
  XOR U12066 ( .A(n8471), .B(n8472), .Z(n8470) );
  XOR U12067 ( .A(DB[973]), .B(DB[958]), .Z(n8472) );
  AND U12068 ( .A(n770), .B(n8473), .Z(n8471) );
  XOR U12069 ( .A(n8474), .B(n8475), .Z(n8473) );
  XOR U12070 ( .A(DB[958]), .B(DB[943]), .Z(n8475) );
  AND U12071 ( .A(n774), .B(n8476), .Z(n8474) );
  XOR U12072 ( .A(n8477), .B(n8478), .Z(n8476) );
  XOR U12073 ( .A(DB[943]), .B(DB[928]), .Z(n8478) );
  AND U12074 ( .A(n778), .B(n8479), .Z(n8477) );
  XOR U12075 ( .A(n8480), .B(n8481), .Z(n8479) );
  XOR U12076 ( .A(DB[928]), .B(DB[913]), .Z(n8481) );
  AND U12077 ( .A(n782), .B(n8482), .Z(n8480) );
  XOR U12078 ( .A(n8483), .B(n8484), .Z(n8482) );
  XOR U12079 ( .A(DB[913]), .B(DB[898]), .Z(n8484) );
  AND U12080 ( .A(n786), .B(n8485), .Z(n8483) );
  XOR U12081 ( .A(n8486), .B(n8487), .Z(n8485) );
  XOR U12082 ( .A(DB[898]), .B(DB[883]), .Z(n8487) );
  AND U12083 ( .A(n790), .B(n8488), .Z(n8486) );
  XOR U12084 ( .A(n8489), .B(n8490), .Z(n8488) );
  XOR U12085 ( .A(DB[883]), .B(DB[868]), .Z(n8490) );
  AND U12086 ( .A(n794), .B(n8491), .Z(n8489) );
  XOR U12087 ( .A(n8492), .B(n8493), .Z(n8491) );
  XOR U12088 ( .A(DB[868]), .B(DB[853]), .Z(n8493) );
  AND U12089 ( .A(n798), .B(n8494), .Z(n8492) );
  XOR U12090 ( .A(n8495), .B(n8496), .Z(n8494) );
  XOR U12091 ( .A(DB[853]), .B(DB[838]), .Z(n8496) );
  AND U12092 ( .A(n802), .B(n8497), .Z(n8495) );
  XOR U12093 ( .A(n8498), .B(n8499), .Z(n8497) );
  XOR U12094 ( .A(DB[838]), .B(DB[823]), .Z(n8499) );
  AND U12095 ( .A(n806), .B(n8500), .Z(n8498) );
  XOR U12096 ( .A(n8501), .B(n8502), .Z(n8500) );
  XOR U12097 ( .A(DB[823]), .B(DB[808]), .Z(n8502) );
  AND U12098 ( .A(n810), .B(n8503), .Z(n8501) );
  XOR U12099 ( .A(n8504), .B(n8505), .Z(n8503) );
  XOR U12100 ( .A(DB[808]), .B(DB[793]), .Z(n8505) );
  AND U12101 ( .A(n814), .B(n8506), .Z(n8504) );
  XOR U12102 ( .A(n8507), .B(n8508), .Z(n8506) );
  XOR U12103 ( .A(DB[793]), .B(DB[778]), .Z(n8508) );
  AND U12104 ( .A(n818), .B(n8509), .Z(n8507) );
  XOR U12105 ( .A(n8510), .B(n8511), .Z(n8509) );
  XOR U12106 ( .A(DB[778]), .B(DB[763]), .Z(n8511) );
  AND U12107 ( .A(n822), .B(n8512), .Z(n8510) );
  XOR U12108 ( .A(n8513), .B(n8514), .Z(n8512) );
  XOR U12109 ( .A(DB[763]), .B(DB[748]), .Z(n8514) );
  AND U12110 ( .A(n826), .B(n8515), .Z(n8513) );
  XOR U12111 ( .A(n8516), .B(n8517), .Z(n8515) );
  XOR U12112 ( .A(DB[748]), .B(DB[733]), .Z(n8517) );
  AND U12113 ( .A(n830), .B(n8518), .Z(n8516) );
  XOR U12114 ( .A(n8519), .B(n8520), .Z(n8518) );
  XOR U12115 ( .A(DB[733]), .B(DB[718]), .Z(n8520) );
  AND U12116 ( .A(n834), .B(n8521), .Z(n8519) );
  XOR U12117 ( .A(n8522), .B(n8523), .Z(n8521) );
  XOR U12118 ( .A(DB[718]), .B(DB[703]), .Z(n8523) );
  AND U12119 ( .A(n838), .B(n8524), .Z(n8522) );
  XOR U12120 ( .A(n8525), .B(n8526), .Z(n8524) );
  XOR U12121 ( .A(DB[703]), .B(DB[688]), .Z(n8526) );
  AND U12122 ( .A(n842), .B(n8527), .Z(n8525) );
  XOR U12123 ( .A(n8528), .B(n8529), .Z(n8527) );
  XOR U12124 ( .A(DB[688]), .B(DB[673]), .Z(n8529) );
  AND U12125 ( .A(n846), .B(n8530), .Z(n8528) );
  XOR U12126 ( .A(n8531), .B(n8532), .Z(n8530) );
  XOR U12127 ( .A(DB[673]), .B(DB[658]), .Z(n8532) );
  AND U12128 ( .A(n850), .B(n8533), .Z(n8531) );
  XOR U12129 ( .A(n8534), .B(n8535), .Z(n8533) );
  XOR U12130 ( .A(DB[658]), .B(DB[643]), .Z(n8535) );
  AND U12131 ( .A(n854), .B(n8536), .Z(n8534) );
  XOR U12132 ( .A(n8537), .B(n8538), .Z(n8536) );
  XOR U12133 ( .A(DB[643]), .B(DB[628]), .Z(n8538) );
  AND U12134 ( .A(n858), .B(n8539), .Z(n8537) );
  XOR U12135 ( .A(n8540), .B(n8541), .Z(n8539) );
  XOR U12136 ( .A(DB[628]), .B(DB[613]), .Z(n8541) );
  AND U12137 ( .A(n862), .B(n8542), .Z(n8540) );
  XOR U12138 ( .A(n8543), .B(n8544), .Z(n8542) );
  XOR U12139 ( .A(DB[613]), .B(DB[598]), .Z(n8544) );
  AND U12140 ( .A(n866), .B(n8545), .Z(n8543) );
  XOR U12141 ( .A(n8546), .B(n8547), .Z(n8545) );
  XOR U12142 ( .A(DB[598]), .B(DB[583]), .Z(n8547) );
  AND U12143 ( .A(n870), .B(n8548), .Z(n8546) );
  XOR U12144 ( .A(n8549), .B(n8550), .Z(n8548) );
  XOR U12145 ( .A(DB[583]), .B(DB[568]), .Z(n8550) );
  AND U12146 ( .A(n874), .B(n8551), .Z(n8549) );
  XOR U12147 ( .A(n8552), .B(n8553), .Z(n8551) );
  XOR U12148 ( .A(DB[568]), .B(DB[553]), .Z(n8553) );
  AND U12149 ( .A(n878), .B(n8554), .Z(n8552) );
  XOR U12150 ( .A(n8555), .B(n8556), .Z(n8554) );
  XOR U12151 ( .A(DB[553]), .B(DB[538]), .Z(n8556) );
  AND U12152 ( .A(n882), .B(n8557), .Z(n8555) );
  XOR U12153 ( .A(n8558), .B(n8559), .Z(n8557) );
  XOR U12154 ( .A(DB[538]), .B(DB[523]), .Z(n8559) );
  AND U12155 ( .A(n886), .B(n8560), .Z(n8558) );
  XOR U12156 ( .A(n8561), .B(n8562), .Z(n8560) );
  XOR U12157 ( .A(DB[523]), .B(DB[508]), .Z(n8562) );
  AND U12158 ( .A(n890), .B(n8563), .Z(n8561) );
  XOR U12159 ( .A(n8564), .B(n8565), .Z(n8563) );
  XOR U12160 ( .A(DB[508]), .B(DB[493]), .Z(n8565) );
  AND U12161 ( .A(n894), .B(n8566), .Z(n8564) );
  XOR U12162 ( .A(n8567), .B(n8568), .Z(n8566) );
  XOR U12163 ( .A(DB[493]), .B(DB[478]), .Z(n8568) );
  AND U12164 ( .A(n898), .B(n8569), .Z(n8567) );
  XOR U12165 ( .A(n8570), .B(n8571), .Z(n8569) );
  XOR U12166 ( .A(DB[478]), .B(DB[463]), .Z(n8571) );
  AND U12167 ( .A(n902), .B(n8572), .Z(n8570) );
  XOR U12168 ( .A(n8573), .B(n8574), .Z(n8572) );
  XOR U12169 ( .A(DB[463]), .B(DB[448]), .Z(n8574) );
  AND U12170 ( .A(n906), .B(n8575), .Z(n8573) );
  XOR U12171 ( .A(n8576), .B(n8577), .Z(n8575) );
  XOR U12172 ( .A(DB[448]), .B(DB[433]), .Z(n8577) );
  AND U12173 ( .A(n910), .B(n8578), .Z(n8576) );
  XOR U12174 ( .A(n8579), .B(n8580), .Z(n8578) );
  XOR U12175 ( .A(DB[433]), .B(DB[418]), .Z(n8580) );
  AND U12176 ( .A(n914), .B(n8581), .Z(n8579) );
  XOR U12177 ( .A(n8582), .B(n8583), .Z(n8581) );
  XOR U12178 ( .A(DB[418]), .B(DB[403]), .Z(n8583) );
  AND U12179 ( .A(n918), .B(n8584), .Z(n8582) );
  XOR U12180 ( .A(n8585), .B(n8586), .Z(n8584) );
  XOR U12181 ( .A(DB[403]), .B(DB[388]), .Z(n8586) );
  AND U12182 ( .A(n922), .B(n8587), .Z(n8585) );
  XOR U12183 ( .A(n8588), .B(n8589), .Z(n8587) );
  XOR U12184 ( .A(DB[388]), .B(DB[373]), .Z(n8589) );
  AND U12185 ( .A(n926), .B(n8590), .Z(n8588) );
  XOR U12186 ( .A(n8591), .B(n8592), .Z(n8590) );
  XOR U12187 ( .A(DB[373]), .B(DB[358]), .Z(n8592) );
  AND U12188 ( .A(n930), .B(n8593), .Z(n8591) );
  XOR U12189 ( .A(n8594), .B(n8595), .Z(n8593) );
  XOR U12190 ( .A(DB[358]), .B(DB[343]), .Z(n8595) );
  AND U12191 ( .A(n934), .B(n8596), .Z(n8594) );
  XOR U12192 ( .A(n8597), .B(n8598), .Z(n8596) );
  XOR U12193 ( .A(DB[343]), .B(DB[328]), .Z(n8598) );
  AND U12194 ( .A(n938), .B(n8599), .Z(n8597) );
  XOR U12195 ( .A(n8600), .B(n8601), .Z(n8599) );
  XOR U12196 ( .A(DB[328]), .B(DB[313]), .Z(n8601) );
  AND U12197 ( .A(n942), .B(n8602), .Z(n8600) );
  XOR U12198 ( .A(n8603), .B(n8604), .Z(n8602) );
  XOR U12199 ( .A(DB[313]), .B(DB[298]), .Z(n8604) );
  AND U12200 ( .A(n946), .B(n8605), .Z(n8603) );
  XOR U12201 ( .A(n8606), .B(n8607), .Z(n8605) );
  XOR U12202 ( .A(DB[298]), .B(DB[283]), .Z(n8607) );
  AND U12203 ( .A(n950), .B(n8608), .Z(n8606) );
  XOR U12204 ( .A(n8609), .B(n8610), .Z(n8608) );
  XOR U12205 ( .A(DB[283]), .B(DB[268]), .Z(n8610) );
  AND U12206 ( .A(n954), .B(n8611), .Z(n8609) );
  XOR U12207 ( .A(n8612), .B(n8613), .Z(n8611) );
  XOR U12208 ( .A(DB[268]), .B(DB[253]), .Z(n8613) );
  AND U12209 ( .A(n958), .B(n8614), .Z(n8612) );
  XOR U12210 ( .A(n8615), .B(n8616), .Z(n8614) );
  XOR U12211 ( .A(DB[253]), .B(DB[238]), .Z(n8616) );
  AND U12212 ( .A(n962), .B(n8617), .Z(n8615) );
  XOR U12213 ( .A(n8618), .B(n8619), .Z(n8617) );
  XOR U12214 ( .A(DB[238]), .B(DB[223]), .Z(n8619) );
  AND U12215 ( .A(n966), .B(n8620), .Z(n8618) );
  XOR U12216 ( .A(n8621), .B(n8622), .Z(n8620) );
  XOR U12217 ( .A(DB[223]), .B(DB[208]), .Z(n8622) );
  AND U12218 ( .A(n970), .B(n8623), .Z(n8621) );
  XOR U12219 ( .A(n8624), .B(n8625), .Z(n8623) );
  XOR U12220 ( .A(DB[208]), .B(DB[193]), .Z(n8625) );
  AND U12221 ( .A(n974), .B(n8626), .Z(n8624) );
  XOR U12222 ( .A(n8627), .B(n8628), .Z(n8626) );
  XOR U12223 ( .A(DB[193]), .B(DB[178]), .Z(n8628) );
  AND U12224 ( .A(n978), .B(n8629), .Z(n8627) );
  XOR U12225 ( .A(n8630), .B(n8631), .Z(n8629) );
  XOR U12226 ( .A(DB[178]), .B(DB[163]), .Z(n8631) );
  AND U12227 ( .A(n982), .B(n8632), .Z(n8630) );
  XOR U12228 ( .A(n8633), .B(n8634), .Z(n8632) );
  XOR U12229 ( .A(DB[163]), .B(DB[148]), .Z(n8634) );
  AND U12230 ( .A(n986), .B(n8635), .Z(n8633) );
  XOR U12231 ( .A(n8636), .B(n8637), .Z(n8635) );
  XOR U12232 ( .A(DB[148]), .B(DB[133]), .Z(n8637) );
  AND U12233 ( .A(n990), .B(n8638), .Z(n8636) );
  XOR U12234 ( .A(n8639), .B(n8640), .Z(n8638) );
  XOR U12235 ( .A(DB[133]), .B(DB[118]), .Z(n8640) );
  AND U12236 ( .A(n994), .B(n8641), .Z(n8639) );
  XOR U12237 ( .A(n8642), .B(n8643), .Z(n8641) );
  XOR U12238 ( .A(DB[118]), .B(DB[103]), .Z(n8643) );
  AND U12239 ( .A(n998), .B(n8644), .Z(n8642) );
  XOR U12240 ( .A(n8645), .B(n8646), .Z(n8644) );
  XOR U12241 ( .A(DB[88]), .B(DB[103]), .Z(n8646) );
  AND U12242 ( .A(n1002), .B(n8647), .Z(n8645) );
  XOR U12243 ( .A(n8648), .B(n8649), .Z(n8647) );
  XOR U12244 ( .A(DB[88]), .B(DB[73]), .Z(n8649) );
  AND U12245 ( .A(n1006), .B(n8650), .Z(n8648) );
  XOR U12246 ( .A(n8651), .B(n8652), .Z(n8650) );
  XOR U12247 ( .A(DB[73]), .B(DB[58]), .Z(n8652) );
  AND U12248 ( .A(n1010), .B(n8653), .Z(n8651) );
  XOR U12249 ( .A(n8654), .B(n8655), .Z(n8653) );
  XOR U12250 ( .A(DB[58]), .B(DB[43]), .Z(n8655) );
  AND U12251 ( .A(n1014), .B(n8656), .Z(n8654) );
  XOR U12252 ( .A(n8657), .B(n8658), .Z(n8656) );
  XOR U12253 ( .A(DB[43]), .B(DB[28]), .Z(n8658) );
  AND U12254 ( .A(n1018), .B(n8659), .Z(n8657) );
  XOR U12255 ( .A(DB[28]), .B(DB[13]), .Z(n8659) );
  XOR U12256 ( .A(DB[3837]), .B(n8660), .Z(min_val_out[12]) );
  AND U12257 ( .A(n2), .B(n8661), .Z(n8660) );
  XOR U12258 ( .A(n8662), .B(n8663), .Z(n8661) );
  XOR U12259 ( .A(n8664), .B(n8665), .Z(n8663) );
  IV U12260 ( .A(DB[3837]), .Z(n8664) );
  AND U12261 ( .A(n6), .B(n8666), .Z(n8662) );
  XOR U12262 ( .A(n8667), .B(n8668), .Z(n8666) );
  XOR U12263 ( .A(DB[3822]), .B(DB[3807]), .Z(n8668) );
  AND U12264 ( .A(n10), .B(n8669), .Z(n8667) );
  XOR U12265 ( .A(n8670), .B(n8671), .Z(n8669) );
  XOR U12266 ( .A(DB[3807]), .B(DB[3792]), .Z(n8671) );
  AND U12267 ( .A(n14), .B(n8672), .Z(n8670) );
  XOR U12268 ( .A(n8673), .B(n8674), .Z(n8672) );
  XOR U12269 ( .A(DB[3792]), .B(DB[3777]), .Z(n8674) );
  AND U12270 ( .A(n18), .B(n8675), .Z(n8673) );
  XOR U12271 ( .A(n8676), .B(n8677), .Z(n8675) );
  XOR U12272 ( .A(DB[3777]), .B(DB[3762]), .Z(n8677) );
  AND U12273 ( .A(n22), .B(n8678), .Z(n8676) );
  XOR U12274 ( .A(n8679), .B(n8680), .Z(n8678) );
  XOR U12275 ( .A(DB[3762]), .B(DB[3747]), .Z(n8680) );
  AND U12276 ( .A(n26), .B(n8681), .Z(n8679) );
  XOR U12277 ( .A(n8682), .B(n8683), .Z(n8681) );
  XOR U12278 ( .A(DB[3747]), .B(DB[3732]), .Z(n8683) );
  AND U12279 ( .A(n30), .B(n8684), .Z(n8682) );
  XOR U12280 ( .A(n8685), .B(n8686), .Z(n8684) );
  XOR U12281 ( .A(DB[3732]), .B(DB[3717]), .Z(n8686) );
  AND U12282 ( .A(n34), .B(n8687), .Z(n8685) );
  XOR U12283 ( .A(n8688), .B(n8689), .Z(n8687) );
  XOR U12284 ( .A(DB[3717]), .B(DB[3702]), .Z(n8689) );
  AND U12285 ( .A(n38), .B(n8690), .Z(n8688) );
  XOR U12286 ( .A(n8691), .B(n8692), .Z(n8690) );
  XOR U12287 ( .A(DB[3702]), .B(DB[3687]), .Z(n8692) );
  AND U12288 ( .A(n42), .B(n8693), .Z(n8691) );
  XOR U12289 ( .A(n8694), .B(n8695), .Z(n8693) );
  XOR U12290 ( .A(DB[3687]), .B(DB[3672]), .Z(n8695) );
  AND U12291 ( .A(n46), .B(n8696), .Z(n8694) );
  XOR U12292 ( .A(n8697), .B(n8698), .Z(n8696) );
  XOR U12293 ( .A(DB[3672]), .B(DB[3657]), .Z(n8698) );
  AND U12294 ( .A(n50), .B(n8699), .Z(n8697) );
  XOR U12295 ( .A(n8700), .B(n8701), .Z(n8699) );
  XOR U12296 ( .A(DB[3657]), .B(DB[3642]), .Z(n8701) );
  AND U12297 ( .A(n54), .B(n8702), .Z(n8700) );
  XOR U12298 ( .A(n8703), .B(n8704), .Z(n8702) );
  XOR U12299 ( .A(DB[3642]), .B(DB[3627]), .Z(n8704) );
  AND U12300 ( .A(n58), .B(n8705), .Z(n8703) );
  XOR U12301 ( .A(n8706), .B(n8707), .Z(n8705) );
  XOR U12302 ( .A(DB[3627]), .B(DB[3612]), .Z(n8707) );
  AND U12303 ( .A(n62), .B(n8708), .Z(n8706) );
  XOR U12304 ( .A(n8709), .B(n8710), .Z(n8708) );
  XOR U12305 ( .A(DB[3612]), .B(DB[3597]), .Z(n8710) );
  AND U12306 ( .A(n66), .B(n8711), .Z(n8709) );
  XOR U12307 ( .A(n8712), .B(n8713), .Z(n8711) );
  XOR U12308 ( .A(DB[3597]), .B(DB[3582]), .Z(n8713) );
  AND U12309 ( .A(n70), .B(n8714), .Z(n8712) );
  XOR U12310 ( .A(n8715), .B(n8716), .Z(n8714) );
  XOR U12311 ( .A(DB[3582]), .B(DB[3567]), .Z(n8716) );
  AND U12312 ( .A(n74), .B(n8717), .Z(n8715) );
  XOR U12313 ( .A(n8718), .B(n8719), .Z(n8717) );
  XOR U12314 ( .A(DB[3567]), .B(DB[3552]), .Z(n8719) );
  AND U12315 ( .A(n78), .B(n8720), .Z(n8718) );
  XOR U12316 ( .A(n8721), .B(n8722), .Z(n8720) );
  XOR U12317 ( .A(DB[3552]), .B(DB[3537]), .Z(n8722) );
  AND U12318 ( .A(n82), .B(n8723), .Z(n8721) );
  XOR U12319 ( .A(n8724), .B(n8725), .Z(n8723) );
  XOR U12320 ( .A(DB[3537]), .B(DB[3522]), .Z(n8725) );
  AND U12321 ( .A(n86), .B(n8726), .Z(n8724) );
  XOR U12322 ( .A(n8727), .B(n8728), .Z(n8726) );
  XOR U12323 ( .A(DB[3522]), .B(DB[3507]), .Z(n8728) );
  AND U12324 ( .A(n90), .B(n8729), .Z(n8727) );
  XOR U12325 ( .A(n8730), .B(n8731), .Z(n8729) );
  XOR U12326 ( .A(DB[3507]), .B(DB[3492]), .Z(n8731) );
  AND U12327 ( .A(n94), .B(n8732), .Z(n8730) );
  XOR U12328 ( .A(n8733), .B(n8734), .Z(n8732) );
  XOR U12329 ( .A(DB[3492]), .B(DB[3477]), .Z(n8734) );
  AND U12330 ( .A(n98), .B(n8735), .Z(n8733) );
  XOR U12331 ( .A(n8736), .B(n8737), .Z(n8735) );
  XOR U12332 ( .A(DB[3477]), .B(DB[3462]), .Z(n8737) );
  AND U12333 ( .A(n102), .B(n8738), .Z(n8736) );
  XOR U12334 ( .A(n8739), .B(n8740), .Z(n8738) );
  XOR U12335 ( .A(DB[3462]), .B(DB[3447]), .Z(n8740) );
  AND U12336 ( .A(n106), .B(n8741), .Z(n8739) );
  XOR U12337 ( .A(n8742), .B(n8743), .Z(n8741) );
  XOR U12338 ( .A(DB[3447]), .B(DB[3432]), .Z(n8743) );
  AND U12339 ( .A(n110), .B(n8744), .Z(n8742) );
  XOR U12340 ( .A(n8745), .B(n8746), .Z(n8744) );
  XOR U12341 ( .A(DB[3432]), .B(DB[3417]), .Z(n8746) );
  AND U12342 ( .A(n114), .B(n8747), .Z(n8745) );
  XOR U12343 ( .A(n8748), .B(n8749), .Z(n8747) );
  XOR U12344 ( .A(DB[3417]), .B(DB[3402]), .Z(n8749) );
  AND U12345 ( .A(n118), .B(n8750), .Z(n8748) );
  XOR U12346 ( .A(n8751), .B(n8752), .Z(n8750) );
  XOR U12347 ( .A(DB[3402]), .B(DB[3387]), .Z(n8752) );
  AND U12348 ( .A(n122), .B(n8753), .Z(n8751) );
  XOR U12349 ( .A(n8754), .B(n8755), .Z(n8753) );
  XOR U12350 ( .A(DB[3387]), .B(DB[3372]), .Z(n8755) );
  AND U12351 ( .A(n126), .B(n8756), .Z(n8754) );
  XOR U12352 ( .A(n8757), .B(n8758), .Z(n8756) );
  XOR U12353 ( .A(DB[3372]), .B(DB[3357]), .Z(n8758) );
  AND U12354 ( .A(n130), .B(n8759), .Z(n8757) );
  XOR U12355 ( .A(n8760), .B(n8761), .Z(n8759) );
  XOR U12356 ( .A(DB[3357]), .B(DB[3342]), .Z(n8761) );
  AND U12357 ( .A(n134), .B(n8762), .Z(n8760) );
  XOR U12358 ( .A(n8763), .B(n8764), .Z(n8762) );
  XOR U12359 ( .A(DB[3342]), .B(DB[3327]), .Z(n8764) );
  AND U12360 ( .A(n138), .B(n8765), .Z(n8763) );
  XOR U12361 ( .A(n8766), .B(n8767), .Z(n8765) );
  XOR U12362 ( .A(DB[3327]), .B(DB[3312]), .Z(n8767) );
  AND U12363 ( .A(n142), .B(n8768), .Z(n8766) );
  XOR U12364 ( .A(n8769), .B(n8770), .Z(n8768) );
  XOR U12365 ( .A(DB[3312]), .B(DB[3297]), .Z(n8770) );
  AND U12366 ( .A(n146), .B(n8771), .Z(n8769) );
  XOR U12367 ( .A(n8772), .B(n8773), .Z(n8771) );
  XOR U12368 ( .A(DB[3297]), .B(DB[3282]), .Z(n8773) );
  AND U12369 ( .A(n150), .B(n8774), .Z(n8772) );
  XOR U12370 ( .A(n8775), .B(n8776), .Z(n8774) );
  XOR U12371 ( .A(DB[3282]), .B(DB[3267]), .Z(n8776) );
  AND U12372 ( .A(n154), .B(n8777), .Z(n8775) );
  XOR U12373 ( .A(n8778), .B(n8779), .Z(n8777) );
  XOR U12374 ( .A(DB[3267]), .B(DB[3252]), .Z(n8779) );
  AND U12375 ( .A(n158), .B(n8780), .Z(n8778) );
  XOR U12376 ( .A(n8781), .B(n8782), .Z(n8780) );
  XOR U12377 ( .A(DB[3252]), .B(DB[3237]), .Z(n8782) );
  AND U12378 ( .A(n162), .B(n8783), .Z(n8781) );
  XOR U12379 ( .A(n8784), .B(n8785), .Z(n8783) );
  XOR U12380 ( .A(DB[3237]), .B(DB[3222]), .Z(n8785) );
  AND U12381 ( .A(n166), .B(n8786), .Z(n8784) );
  XOR U12382 ( .A(n8787), .B(n8788), .Z(n8786) );
  XOR U12383 ( .A(DB[3222]), .B(DB[3207]), .Z(n8788) );
  AND U12384 ( .A(n170), .B(n8789), .Z(n8787) );
  XOR U12385 ( .A(n8790), .B(n8791), .Z(n8789) );
  XOR U12386 ( .A(DB[3207]), .B(DB[3192]), .Z(n8791) );
  AND U12387 ( .A(n174), .B(n8792), .Z(n8790) );
  XOR U12388 ( .A(n8793), .B(n8794), .Z(n8792) );
  XOR U12389 ( .A(DB[3192]), .B(DB[3177]), .Z(n8794) );
  AND U12390 ( .A(n178), .B(n8795), .Z(n8793) );
  XOR U12391 ( .A(n8796), .B(n8797), .Z(n8795) );
  XOR U12392 ( .A(DB[3177]), .B(DB[3162]), .Z(n8797) );
  AND U12393 ( .A(n182), .B(n8798), .Z(n8796) );
  XOR U12394 ( .A(n8799), .B(n8800), .Z(n8798) );
  XOR U12395 ( .A(DB[3162]), .B(DB[3147]), .Z(n8800) );
  AND U12396 ( .A(n186), .B(n8801), .Z(n8799) );
  XOR U12397 ( .A(n8802), .B(n8803), .Z(n8801) );
  XOR U12398 ( .A(DB[3147]), .B(DB[3132]), .Z(n8803) );
  AND U12399 ( .A(n190), .B(n8804), .Z(n8802) );
  XOR U12400 ( .A(n8805), .B(n8806), .Z(n8804) );
  XOR U12401 ( .A(DB[3132]), .B(DB[3117]), .Z(n8806) );
  AND U12402 ( .A(n194), .B(n8807), .Z(n8805) );
  XOR U12403 ( .A(n8808), .B(n8809), .Z(n8807) );
  XOR U12404 ( .A(DB[3117]), .B(DB[3102]), .Z(n8809) );
  AND U12405 ( .A(n198), .B(n8810), .Z(n8808) );
  XOR U12406 ( .A(n8811), .B(n8812), .Z(n8810) );
  XOR U12407 ( .A(DB[3102]), .B(DB[3087]), .Z(n8812) );
  AND U12408 ( .A(n202), .B(n8813), .Z(n8811) );
  XOR U12409 ( .A(n8814), .B(n8815), .Z(n8813) );
  XOR U12410 ( .A(DB[3087]), .B(DB[3072]), .Z(n8815) );
  AND U12411 ( .A(n206), .B(n8816), .Z(n8814) );
  XOR U12412 ( .A(n8817), .B(n8818), .Z(n8816) );
  XOR U12413 ( .A(DB[3072]), .B(DB[3057]), .Z(n8818) );
  AND U12414 ( .A(n210), .B(n8819), .Z(n8817) );
  XOR U12415 ( .A(n8820), .B(n8821), .Z(n8819) );
  XOR U12416 ( .A(DB[3057]), .B(DB[3042]), .Z(n8821) );
  AND U12417 ( .A(n214), .B(n8822), .Z(n8820) );
  XOR U12418 ( .A(n8823), .B(n8824), .Z(n8822) );
  XOR U12419 ( .A(DB[3042]), .B(DB[3027]), .Z(n8824) );
  AND U12420 ( .A(n218), .B(n8825), .Z(n8823) );
  XOR U12421 ( .A(n8826), .B(n8827), .Z(n8825) );
  XOR U12422 ( .A(DB[3027]), .B(DB[3012]), .Z(n8827) );
  AND U12423 ( .A(n222), .B(n8828), .Z(n8826) );
  XOR U12424 ( .A(n8829), .B(n8830), .Z(n8828) );
  XOR U12425 ( .A(DB[3012]), .B(DB[2997]), .Z(n8830) );
  AND U12426 ( .A(n226), .B(n8831), .Z(n8829) );
  XOR U12427 ( .A(n8832), .B(n8833), .Z(n8831) );
  XOR U12428 ( .A(DB[2997]), .B(DB[2982]), .Z(n8833) );
  AND U12429 ( .A(n230), .B(n8834), .Z(n8832) );
  XOR U12430 ( .A(n8835), .B(n8836), .Z(n8834) );
  XOR U12431 ( .A(DB[2982]), .B(DB[2967]), .Z(n8836) );
  AND U12432 ( .A(n234), .B(n8837), .Z(n8835) );
  XOR U12433 ( .A(n8838), .B(n8839), .Z(n8837) );
  XOR U12434 ( .A(DB[2967]), .B(DB[2952]), .Z(n8839) );
  AND U12435 ( .A(n238), .B(n8840), .Z(n8838) );
  XOR U12436 ( .A(n8841), .B(n8842), .Z(n8840) );
  XOR U12437 ( .A(DB[2952]), .B(DB[2937]), .Z(n8842) );
  AND U12438 ( .A(n242), .B(n8843), .Z(n8841) );
  XOR U12439 ( .A(n8844), .B(n8845), .Z(n8843) );
  XOR U12440 ( .A(DB[2937]), .B(DB[2922]), .Z(n8845) );
  AND U12441 ( .A(n246), .B(n8846), .Z(n8844) );
  XOR U12442 ( .A(n8847), .B(n8848), .Z(n8846) );
  XOR U12443 ( .A(DB[2922]), .B(DB[2907]), .Z(n8848) );
  AND U12444 ( .A(n250), .B(n8849), .Z(n8847) );
  XOR U12445 ( .A(n8850), .B(n8851), .Z(n8849) );
  XOR U12446 ( .A(DB[2907]), .B(DB[2892]), .Z(n8851) );
  AND U12447 ( .A(n254), .B(n8852), .Z(n8850) );
  XOR U12448 ( .A(n8853), .B(n8854), .Z(n8852) );
  XOR U12449 ( .A(DB[2892]), .B(DB[2877]), .Z(n8854) );
  AND U12450 ( .A(n258), .B(n8855), .Z(n8853) );
  XOR U12451 ( .A(n8856), .B(n8857), .Z(n8855) );
  XOR U12452 ( .A(DB[2877]), .B(DB[2862]), .Z(n8857) );
  AND U12453 ( .A(n262), .B(n8858), .Z(n8856) );
  XOR U12454 ( .A(n8859), .B(n8860), .Z(n8858) );
  XOR U12455 ( .A(DB[2862]), .B(DB[2847]), .Z(n8860) );
  AND U12456 ( .A(n266), .B(n8861), .Z(n8859) );
  XOR U12457 ( .A(n8862), .B(n8863), .Z(n8861) );
  XOR U12458 ( .A(DB[2847]), .B(DB[2832]), .Z(n8863) );
  AND U12459 ( .A(n270), .B(n8864), .Z(n8862) );
  XOR U12460 ( .A(n8865), .B(n8866), .Z(n8864) );
  XOR U12461 ( .A(DB[2832]), .B(DB[2817]), .Z(n8866) );
  AND U12462 ( .A(n274), .B(n8867), .Z(n8865) );
  XOR U12463 ( .A(n8868), .B(n8869), .Z(n8867) );
  XOR U12464 ( .A(DB[2817]), .B(DB[2802]), .Z(n8869) );
  AND U12465 ( .A(n278), .B(n8870), .Z(n8868) );
  XOR U12466 ( .A(n8871), .B(n8872), .Z(n8870) );
  XOR U12467 ( .A(DB[2802]), .B(DB[2787]), .Z(n8872) );
  AND U12468 ( .A(n282), .B(n8873), .Z(n8871) );
  XOR U12469 ( .A(n8874), .B(n8875), .Z(n8873) );
  XOR U12470 ( .A(DB[2787]), .B(DB[2772]), .Z(n8875) );
  AND U12471 ( .A(n286), .B(n8876), .Z(n8874) );
  XOR U12472 ( .A(n8877), .B(n8878), .Z(n8876) );
  XOR U12473 ( .A(DB[2772]), .B(DB[2757]), .Z(n8878) );
  AND U12474 ( .A(n290), .B(n8879), .Z(n8877) );
  XOR U12475 ( .A(n8880), .B(n8881), .Z(n8879) );
  XOR U12476 ( .A(DB[2757]), .B(DB[2742]), .Z(n8881) );
  AND U12477 ( .A(n294), .B(n8882), .Z(n8880) );
  XOR U12478 ( .A(n8883), .B(n8884), .Z(n8882) );
  XOR U12479 ( .A(DB[2742]), .B(DB[2727]), .Z(n8884) );
  AND U12480 ( .A(n298), .B(n8885), .Z(n8883) );
  XOR U12481 ( .A(n8886), .B(n8887), .Z(n8885) );
  XOR U12482 ( .A(DB[2727]), .B(DB[2712]), .Z(n8887) );
  AND U12483 ( .A(n302), .B(n8888), .Z(n8886) );
  XOR U12484 ( .A(n8889), .B(n8890), .Z(n8888) );
  XOR U12485 ( .A(DB[2712]), .B(DB[2697]), .Z(n8890) );
  AND U12486 ( .A(n306), .B(n8891), .Z(n8889) );
  XOR U12487 ( .A(n8892), .B(n8893), .Z(n8891) );
  XOR U12488 ( .A(DB[2697]), .B(DB[2682]), .Z(n8893) );
  AND U12489 ( .A(n310), .B(n8894), .Z(n8892) );
  XOR U12490 ( .A(n8895), .B(n8896), .Z(n8894) );
  XOR U12491 ( .A(DB[2682]), .B(DB[2667]), .Z(n8896) );
  AND U12492 ( .A(n314), .B(n8897), .Z(n8895) );
  XOR U12493 ( .A(n8898), .B(n8899), .Z(n8897) );
  XOR U12494 ( .A(DB[2667]), .B(DB[2652]), .Z(n8899) );
  AND U12495 ( .A(n318), .B(n8900), .Z(n8898) );
  XOR U12496 ( .A(n8901), .B(n8902), .Z(n8900) );
  XOR U12497 ( .A(DB[2652]), .B(DB[2637]), .Z(n8902) );
  AND U12498 ( .A(n322), .B(n8903), .Z(n8901) );
  XOR U12499 ( .A(n8904), .B(n8905), .Z(n8903) );
  XOR U12500 ( .A(DB[2637]), .B(DB[2622]), .Z(n8905) );
  AND U12501 ( .A(n326), .B(n8906), .Z(n8904) );
  XOR U12502 ( .A(n8907), .B(n8908), .Z(n8906) );
  XOR U12503 ( .A(DB[2622]), .B(DB[2607]), .Z(n8908) );
  AND U12504 ( .A(n330), .B(n8909), .Z(n8907) );
  XOR U12505 ( .A(n8910), .B(n8911), .Z(n8909) );
  XOR U12506 ( .A(DB[2607]), .B(DB[2592]), .Z(n8911) );
  AND U12507 ( .A(n334), .B(n8912), .Z(n8910) );
  XOR U12508 ( .A(n8913), .B(n8914), .Z(n8912) );
  XOR U12509 ( .A(DB[2592]), .B(DB[2577]), .Z(n8914) );
  AND U12510 ( .A(n338), .B(n8915), .Z(n8913) );
  XOR U12511 ( .A(n8916), .B(n8917), .Z(n8915) );
  XOR U12512 ( .A(DB[2577]), .B(DB[2562]), .Z(n8917) );
  AND U12513 ( .A(n342), .B(n8918), .Z(n8916) );
  XOR U12514 ( .A(n8919), .B(n8920), .Z(n8918) );
  XOR U12515 ( .A(DB[2562]), .B(DB[2547]), .Z(n8920) );
  AND U12516 ( .A(n346), .B(n8921), .Z(n8919) );
  XOR U12517 ( .A(n8922), .B(n8923), .Z(n8921) );
  XOR U12518 ( .A(DB[2547]), .B(DB[2532]), .Z(n8923) );
  AND U12519 ( .A(n350), .B(n8924), .Z(n8922) );
  XOR U12520 ( .A(n8925), .B(n8926), .Z(n8924) );
  XOR U12521 ( .A(DB[2532]), .B(DB[2517]), .Z(n8926) );
  AND U12522 ( .A(n354), .B(n8927), .Z(n8925) );
  XOR U12523 ( .A(n8928), .B(n8929), .Z(n8927) );
  XOR U12524 ( .A(DB[2517]), .B(DB[2502]), .Z(n8929) );
  AND U12525 ( .A(n358), .B(n8930), .Z(n8928) );
  XOR U12526 ( .A(n8931), .B(n8932), .Z(n8930) );
  XOR U12527 ( .A(DB[2502]), .B(DB[2487]), .Z(n8932) );
  AND U12528 ( .A(n362), .B(n8933), .Z(n8931) );
  XOR U12529 ( .A(n8934), .B(n8935), .Z(n8933) );
  XOR U12530 ( .A(DB[2487]), .B(DB[2472]), .Z(n8935) );
  AND U12531 ( .A(n366), .B(n8936), .Z(n8934) );
  XOR U12532 ( .A(n8937), .B(n8938), .Z(n8936) );
  XOR U12533 ( .A(DB[2472]), .B(DB[2457]), .Z(n8938) );
  AND U12534 ( .A(n370), .B(n8939), .Z(n8937) );
  XOR U12535 ( .A(n8940), .B(n8941), .Z(n8939) );
  XOR U12536 ( .A(DB[2457]), .B(DB[2442]), .Z(n8941) );
  AND U12537 ( .A(n374), .B(n8942), .Z(n8940) );
  XOR U12538 ( .A(n8943), .B(n8944), .Z(n8942) );
  XOR U12539 ( .A(DB[2442]), .B(DB[2427]), .Z(n8944) );
  AND U12540 ( .A(n378), .B(n8945), .Z(n8943) );
  XOR U12541 ( .A(n8946), .B(n8947), .Z(n8945) );
  XOR U12542 ( .A(DB[2427]), .B(DB[2412]), .Z(n8947) );
  AND U12543 ( .A(n382), .B(n8948), .Z(n8946) );
  XOR U12544 ( .A(n8949), .B(n8950), .Z(n8948) );
  XOR U12545 ( .A(DB[2412]), .B(DB[2397]), .Z(n8950) );
  AND U12546 ( .A(n386), .B(n8951), .Z(n8949) );
  XOR U12547 ( .A(n8952), .B(n8953), .Z(n8951) );
  XOR U12548 ( .A(DB[2397]), .B(DB[2382]), .Z(n8953) );
  AND U12549 ( .A(n390), .B(n8954), .Z(n8952) );
  XOR U12550 ( .A(n8955), .B(n8956), .Z(n8954) );
  XOR U12551 ( .A(DB[2382]), .B(DB[2367]), .Z(n8956) );
  AND U12552 ( .A(n394), .B(n8957), .Z(n8955) );
  XOR U12553 ( .A(n8958), .B(n8959), .Z(n8957) );
  XOR U12554 ( .A(DB[2367]), .B(DB[2352]), .Z(n8959) );
  AND U12555 ( .A(n398), .B(n8960), .Z(n8958) );
  XOR U12556 ( .A(n8961), .B(n8962), .Z(n8960) );
  XOR U12557 ( .A(DB[2352]), .B(DB[2337]), .Z(n8962) );
  AND U12558 ( .A(n402), .B(n8963), .Z(n8961) );
  XOR U12559 ( .A(n8964), .B(n8965), .Z(n8963) );
  XOR U12560 ( .A(DB[2337]), .B(DB[2322]), .Z(n8965) );
  AND U12561 ( .A(n406), .B(n8966), .Z(n8964) );
  XOR U12562 ( .A(n8967), .B(n8968), .Z(n8966) );
  XOR U12563 ( .A(DB[2322]), .B(DB[2307]), .Z(n8968) );
  AND U12564 ( .A(n410), .B(n8969), .Z(n8967) );
  XOR U12565 ( .A(n8970), .B(n8971), .Z(n8969) );
  XOR U12566 ( .A(DB[2307]), .B(DB[2292]), .Z(n8971) );
  AND U12567 ( .A(n414), .B(n8972), .Z(n8970) );
  XOR U12568 ( .A(n8973), .B(n8974), .Z(n8972) );
  XOR U12569 ( .A(DB[2292]), .B(DB[2277]), .Z(n8974) );
  AND U12570 ( .A(n418), .B(n8975), .Z(n8973) );
  XOR U12571 ( .A(n8976), .B(n8977), .Z(n8975) );
  XOR U12572 ( .A(DB[2277]), .B(DB[2262]), .Z(n8977) );
  AND U12573 ( .A(n422), .B(n8978), .Z(n8976) );
  XOR U12574 ( .A(n8979), .B(n8980), .Z(n8978) );
  XOR U12575 ( .A(DB[2262]), .B(DB[2247]), .Z(n8980) );
  AND U12576 ( .A(n426), .B(n8981), .Z(n8979) );
  XOR U12577 ( .A(n8982), .B(n8983), .Z(n8981) );
  XOR U12578 ( .A(DB[2247]), .B(DB[2232]), .Z(n8983) );
  AND U12579 ( .A(n430), .B(n8984), .Z(n8982) );
  XOR U12580 ( .A(n8985), .B(n8986), .Z(n8984) );
  XOR U12581 ( .A(DB[2232]), .B(DB[2217]), .Z(n8986) );
  AND U12582 ( .A(n434), .B(n8987), .Z(n8985) );
  XOR U12583 ( .A(n8988), .B(n8989), .Z(n8987) );
  XOR U12584 ( .A(DB[2217]), .B(DB[2202]), .Z(n8989) );
  AND U12585 ( .A(n438), .B(n8990), .Z(n8988) );
  XOR U12586 ( .A(n8991), .B(n8992), .Z(n8990) );
  XOR U12587 ( .A(DB[2202]), .B(DB[2187]), .Z(n8992) );
  AND U12588 ( .A(n442), .B(n8993), .Z(n8991) );
  XOR U12589 ( .A(n8994), .B(n8995), .Z(n8993) );
  XOR U12590 ( .A(DB[2187]), .B(DB[2172]), .Z(n8995) );
  AND U12591 ( .A(n446), .B(n8996), .Z(n8994) );
  XOR U12592 ( .A(n8997), .B(n8998), .Z(n8996) );
  XOR U12593 ( .A(DB[2172]), .B(DB[2157]), .Z(n8998) );
  AND U12594 ( .A(n450), .B(n8999), .Z(n8997) );
  XOR U12595 ( .A(n9000), .B(n9001), .Z(n8999) );
  XOR U12596 ( .A(DB[2157]), .B(DB[2142]), .Z(n9001) );
  AND U12597 ( .A(n454), .B(n9002), .Z(n9000) );
  XOR U12598 ( .A(n9003), .B(n9004), .Z(n9002) );
  XOR U12599 ( .A(DB[2142]), .B(DB[2127]), .Z(n9004) );
  AND U12600 ( .A(n458), .B(n9005), .Z(n9003) );
  XOR U12601 ( .A(n9006), .B(n9007), .Z(n9005) );
  XOR U12602 ( .A(DB[2127]), .B(DB[2112]), .Z(n9007) );
  AND U12603 ( .A(n462), .B(n9008), .Z(n9006) );
  XOR U12604 ( .A(n9009), .B(n9010), .Z(n9008) );
  XOR U12605 ( .A(DB[2112]), .B(DB[2097]), .Z(n9010) );
  AND U12606 ( .A(n466), .B(n9011), .Z(n9009) );
  XOR U12607 ( .A(n9012), .B(n9013), .Z(n9011) );
  XOR U12608 ( .A(DB[2097]), .B(DB[2082]), .Z(n9013) );
  AND U12609 ( .A(n470), .B(n9014), .Z(n9012) );
  XOR U12610 ( .A(n9015), .B(n9016), .Z(n9014) );
  XOR U12611 ( .A(DB[2082]), .B(DB[2067]), .Z(n9016) );
  AND U12612 ( .A(n474), .B(n9017), .Z(n9015) );
  XOR U12613 ( .A(n9018), .B(n9019), .Z(n9017) );
  XOR U12614 ( .A(DB[2067]), .B(DB[2052]), .Z(n9019) );
  AND U12615 ( .A(n478), .B(n9020), .Z(n9018) );
  XOR U12616 ( .A(n9021), .B(n9022), .Z(n9020) );
  XOR U12617 ( .A(DB[2052]), .B(DB[2037]), .Z(n9022) );
  AND U12618 ( .A(n482), .B(n9023), .Z(n9021) );
  XOR U12619 ( .A(n9024), .B(n9025), .Z(n9023) );
  XOR U12620 ( .A(DB[2037]), .B(DB[2022]), .Z(n9025) );
  AND U12621 ( .A(n486), .B(n9026), .Z(n9024) );
  XOR U12622 ( .A(n9027), .B(n9028), .Z(n9026) );
  XOR U12623 ( .A(DB[2022]), .B(DB[2007]), .Z(n9028) );
  AND U12624 ( .A(n490), .B(n9029), .Z(n9027) );
  XOR U12625 ( .A(n9030), .B(n9031), .Z(n9029) );
  XOR U12626 ( .A(DB[2007]), .B(DB[1992]), .Z(n9031) );
  AND U12627 ( .A(n494), .B(n9032), .Z(n9030) );
  XOR U12628 ( .A(n9033), .B(n9034), .Z(n9032) );
  XOR U12629 ( .A(DB[1992]), .B(DB[1977]), .Z(n9034) );
  AND U12630 ( .A(n498), .B(n9035), .Z(n9033) );
  XOR U12631 ( .A(n9036), .B(n9037), .Z(n9035) );
  XOR U12632 ( .A(DB[1977]), .B(DB[1962]), .Z(n9037) );
  AND U12633 ( .A(n502), .B(n9038), .Z(n9036) );
  XOR U12634 ( .A(n9039), .B(n9040), .Z(n9038) );
  XOR U12635 ( .A(DB[1962]), .B(DB[1947]), .Z(n9040) );
  AND U12636 ( .A(n506), .B(n9041), .Z(n9039) );
  XOR U12637 ( .A(n9042), .B(n9043), .Z(n9041) );
  XOR U12638 ( .A(DB[1947]), .B(DB[1932]), .Z(n9043) );
  AND U12639 ( .A(n510), .B(n9044), .Z(n9042) );
  XOR U12640 ( .A(n9045), .B(n9046), .Z(n9044) );
  XOR U12641 ( .A(DB[1932]), .B(DB[1917]), .Z(n9046) );
  AND U12642 ( .A(n514), .B(n9047), .Z(n9045) );
  XOR U12643 ( .A(n9048), .B(n9049), .Z(n9047) );
  XOR U12644 ( .A(DB[1917]), .B(DB[1902]), .Z(n9049) );
  AND U12645 ( .A(n518), .B(n9050), .Z(n9048) );
  XOR U12646 ( .A(n9051), .B(n9052), .Z(n9050) );
  XOR U12647 ( .A(DB[1902]), .B(DB[1887]), .Z(n9052) );
  AND U12648 ( .A(n522), .B(n9053), .Z(n9051) );
  XOR U12649 ( .A(n9054), .B(n9055), .Z(n9053) );
  XOR U12650 ( .A(DB[1887]), .B(DB[1872]), .Z(n9055) );
  AND U12651 ( .A(n526), .B(n9056), .Z(n9054) );
  XOR U12652 ( .A(n9057), .B(n9058), .Z(n9056) );
  XOR U12653 ( .A(DB[1872]), .B(DB[1857]), .Z(n9058) );
  AND U12654 ( .A(n530), .B(n9059), .Z(n9057) );
  XOR U12655 ( .A(n9060), .B(n9061), .Z(n9059) );
  XOR U12656 ( .A(DB[1857]), .B(DB[1842]), .Z(n9061) );
  AND U12657 ( .A(n534), .B(n9062), .Z(n9060) );
  XOR U12658 ( .A(n9063), .B(n9064), .Z(n9062) );
  XOR U12659 ( .A(DB[1842]), .B(DB[1827]), .Z(n9064) );
  AND U12660 ( .A(n538), .B(n9065), .Z(n9063) );
  XOR U12661 ( .A(n9066), .B(n9067), .Z(n9065) );
  XOR U12662 ( .A(DB[1827]), .B(DB[1812]), .Z(n9067) );
  AND U12663 ( .A(n542), .B(n9068), .Z(n9066) );
  XOR U12664 ( .A(n9069), .B(n9070), .Z(n9068) );
  XOR U12665 ( .A(DB[1812]), .B(DB[1797]), .Z(n9070) );
  AND U12666 ( .A(n546), .B(n9071), .Z(n9069) );
  XOR U12667 ( .A(n9072), .B(n9073), .Z(n9071) );
  XOR U12668 ( .A(DB[1797]), .B(DB[1782]), .Z(n9073) );
  AND U12669 ( .A(n550), .B(n9074), .Z(n9072) );
  XOR U12670 ( .A(n9075), .B(n9076), .Z(n9074) );
  XOR U12671 ( .A(DB[1782]), .B(DB[1767]), .Z(n9076) );
  AND U12672 ( .A(n554), .B(n9077), .Z(n9075) );
  XOR U12673 ( .A(n9078), .B(n9079), .Z(n9077) );
  XOR U12674 ( .A(DB[1767]), .B(DB[1752]), .Z(n9079) );
  AND U12675 ( .A(n558), .B(n9080), .Z(n9078) );
  XOR U12676 ( .A(n9081), .B(n9082), .Z(n9080) );
  XOR U12677 ( .A(DB[1752]), .B(DB[1737]), .Z(n9082) );
  AND U12678 ( .A(n562), .B(n9083), .Z(n9081) );
  XOR U12679 ( .A(n9084), .B(n9085), .Z(n9083) );
  XOR U12680 ( .A(DB[1737]), .B(DB[1722]), .Z(n9085) );
  AND U12681 ( .A(n566), .B(n9086), .Z(n9084) );
  XOR U12682 ( .A(n9087), .B(n9088), .Z(n9086) );
  XOR U12683 ( .A(DB[1722]), .B(DB[1707]), .Z(n9088) );
  AND U12684 ( .A(n570), .B(n9089), .Z(n9087) );
  XOR U12685 ( .A(n9090), .B(n9091), .Z(n9089) );
  XOR U12686 ( .A(DB[1707]), .B(DB[1692]), .Z(n9091) );
  AND U12687 ( .A(n574), .B(n9092), .Z(n9090) );
  XOR U12688 ( .A(n9093), .B(n9094), .Z(n9092) );
  XOR U12689 ( .A(DB[1692]), .B(DB[1677]), .Z(n9094) );
  AND U12690 ( .A(n578), .B(n9095), .Z(n9093) );
  XOR U12691 ( .A(n9096), .B(n9097), .Z(n9095) );
  XOR U12692 ( .A(DB[1677]), .B(DB[1662]), .Z(n9097) );
  AND U12693 ( .A(n582), .B(n9098), .Z(n9096) );
  XOR U12694 ( .A(n9099), .B(n9100), .Z(n9098) );
  XOR U12695 ( .A(DB[1662]), .B(DB[1647]), .Z(n9100) );
  AND U12696 ( .A(n586), .B(n9101), .Z(n9099) );
  XOR U12697 ( .A(n9102), .B(n9103), .Z(n9101) );
  XOR U12698 ( .A(DB[1647]), .B(DB[1632]), .Z(n9103) );
  AND U12699 ( .A(n590), .B(n9104), .Z(n9102) );
  XOR U12700 ( .A(n9105), .B(n9106), .Z(n9104) );
  XOR U12701 ( .A(DB[1632]), .B(DB[1617]), .Z(n9106) );
  AND U12702 ( .A(n594), .B(n9107), .Z(n9105) );
  XOR U12703 ( .A(n9108), .B(n9109), .Z(n9107) );
  XOR U12704 ( .A(DB[1617]), .B(DB[1602]), .Z(n9109) );
  AND U12705 ( .A(n598), .B(n9110), .Z(n9108) );
  XOR U12706 ( .A(n9111), .B(n9112), .Z(n9110) );
  XOR U12707 ( .A(DB[1602]), .B(DB[1587]), .Z(n9112) );
  AND U12708 ( .A(n602), .B(n9113), .Z(n9111) );
  XOR U12709 ( .A(n9114), .B(n9115), .Z(n9113) );
  XOR U12710 ( .A(DB[1587]), .B(DB[1572]), .Z(n9115) );
  AND U12711 ( .A(n606), .B(n9116), .Z(n9114) );
  XOR U12712 ( .A(n9117), .B(n9118), .Z(n9116) );
  XOR U12713 ( .A(DB[1572]), .B(DB[1557]), .Z(n9118) );
  AND U12714 ( .A(n610), .B(n9119), .Z(n9117) );
  XOR U12715 ( .A(n9120), .B(n9121), .Z(n9119) );
  XOR U12716 ( .A(DB[1557]), .B(DB[1542]), .Z(n9121) );
  AND U12717 ( .A(n614), .B(n9122), .Z(n9120) );
  XOR U12718 ( .A(n9123), .B(n9124), .Z(n9122) );
  XOR U12719 ( .A(DB[1542]), .B(DB[1527]), .Z(n9124) );
  AND U12720 ( .A(n618), .B(n9125), .Z(n9123) );
  XOR U12721 ( .A(n9126), .B(n9127), .Z(n9125) );
  XOR U12722 ( .A(DB[1527]), .B(DB[1512]), .Z(n9127) );
  AND U12723 ( .A(n622), .B(n9128), .Z(n9126) );
  XOR U12724 ( .A(n9129), .B(n9130), .Z(n9128) );
  XOR U12725 ( .A(DB[1512]), .B(DB[1497]), .Z(n9130) );
  AND U12726 ( .A(n626), .B(n9131), .Z(n9129) );
  XOR U12727 ( .A(n9132), .B(n9133), .Z(n9131) );
  XOR U12728 ( .A(DB[1497]), .B(DB[1482]), .Z(n9133) );
  AND U12729 ( .A(n630), .B(n9134), .Z(n9132) );
  XOR U12730 ( .A(n9135), .B(n9136), .Z(n9134) );
  XOR U12731 ( .A(DB[1482]), .B(DB[1467]), .Z(n9136) );
  AND U12732 ( .A(n634), .B(n9137), .Z(n9135) );
  XOR U12733 ( .A(n9138), .B(n9139), .Z(n9137) );
  XOR U12734 ( .A(DB[1467]), .B(DB[1452]), .Z(n9139) );
  AND U12735 ( .A(n638), .B(n9140), .Z(n9138) );
  XOR U12736 ( .A(n9141), .B(n9142), .Z(n9140) );
  XOR U12737 ( .A(DB[1452]), .B(DB[1437]), .Z(n9142) );
  AND U12738 ( .A(n642), .B(n9143), .Z(n9141) );
  XOR U12739 ( .A(n9144), .B(n9145), .Z(n9143) );
  XOR U12740 ( .A(DB[1437]), .B(DB[1422]), .Z(n9145) );
  AND U12741 ( .A(n646), .B(n9146), .Z(n9144) );
  XOR U12742 ( .A(n9147), .B(n9148), .Z(n9146) );
  XOR U12743 ( .A(DB[1422]), .B(DB[1407]), .Z(n9148) );
  AND U12744 ( .A(n650), .B(n9149), .Z(n9147) );
  XOR U12745 ( .A(n9150), .B(n9151), .Z(n9149) );
  XOR U12746 ( .A(DB[1407]), .B(DB[1392]), .Z(n9151) );
  AND U12747 ( .A(n654), .B(n9152), .Z(n9150) );
  XOR U12748 ( .A(n9153), .B(n9154), .Z(n9152) );
  XOR U12749 ( .A(DB[1392]), .B(DB[1377]), .Z(n9154) );
  AND U12750 ( .A(n658), .B(n9155), .Z(n9153) );
  XOR U12751 ( .A(n9156), .B(n9157), .Z(n9155) );
  XOR U12752 ( .A(DB[1377]), .B(DB[1362]), .Z(n9157) );
  AND U12753 ( .A(n662), .B(n9158), .Z(n9156) );
  XOR U12754 ( .A(n9159), .B(n9160), .Z(n9158) );
  XOR U12755 ( .A(DB[1362]), .B(DB[1347]), .Z(n9160) );
  AND U12756 ( .A(n666), .B(n9161), .Z(n9159) );
  XOR U12757 ( .A(n9162), .B(n9163), .Z(n9161) );
  XOR U12758 ( .A(DB[1347]), .B(DB[1332]), .Z(n9163) );
  AND U12759 ( .A(n670), .B(n9164), .Z(n9162) );
  XOR U12760 ( .A(n9165), .B(n9166), .Z(n9164) );
  XOR U12761 ( .A(DB[1332]), .B(DB[1317]), .Z(n9166) );
  AND U12762 ( .A(n674), .B(n9167), .Z(n9165) );
  XOR U12763 ( .A(n9168), .B(n9169), .Z(n9167) );
  XOR U12764 ( .A(DB[1317]), .B(DB[1302]), .Z(n9169) );
  AND U12765 ( .A(n678), .B(n9170), .Z(n9168) );
  XOR U12766 ( .A(n9171), .B(n9172), .Z(n9170) );
  XOR U12767 ( .A(DB[1302]), .B(DB[1287]), .Z(n9172) );
  AND U12768 ( .A(n682), .B(n9173), .Z(n9171) );
  XOR U12769 ( .A(n9174), .B(n9175), .Z(n9173) );
  XOR U12770 ( .A(DB[1287]), .B(DB[1272]), .Z(n9175) );
  AND U12771 ( .A(n686), .B(n9176), .Z(n9174) );
  XOR U12772 ( .A(n9177), .B(n9178), .Z(n9176) );
  XOR U12773 ( .A(DB[1272]), .B(DB[1257]), .Z(n9178) );
  AND U12774 ( .A(n690), .B(n9179), .Z(n9177) );
  XOR U12775 ( .A(n9180), .B(n9181), .Z(n9179) );
  XOR U12776 ( .A(DB[1257]), .B(DB[1242]), .Z(n9181) );
  AND U12777 ( .A(n694), .B(n9182), .Z(n9180) );
  XOR U12778 ( .A(n9183), .B(n9184), .Z(n9182) );
  XOR U12779 ( .A(DB[1242]), .B(DB[1227]), .Z(n9184) );
  AND U12780 ( .A(n698), .B(n9185), .Z(n9183) );
  XOR U12781 ( .A(n9186), .B(n9187), .Z(n9185) );
  XOR U12782 ( .A(DB[1227]), .B(DB[1212]), .Z(n9187) );
  AND U12783 ( .A(n702), .B(n9188), .Z(n9186) );
  XOR U12784 ( .A(n9189), .B(n9190), .Z(n9188) );
  XOR U12785 ( .A(DB[1212]), .B(DB[1197]), .Z(n9190) );
  AND U12786 ( .A(n706), .B(n9191), .Z(n9189) );
  XOR U12787 ( .A(n9192), .B(n9193), .Z(n9191) );
  XOR U12788 ( .A(DB[1197]), .B(DB[1182]), .Z(n9193) );
  AND U12789 ( .A(n710), .B(n9194), .Z(n9192) );
  XOR U12790 ( .A(n9195), .B(n9196), .Z(n9194) );
  XOR U12791 ( .A(DB[1182]), .B(DB[1167]), .Z(n9196) );
  AND U12792 ( .A(n714), .B(n9197), .Z(n9195) );
  XOR U12793 ( .A(n9198), .B(n9199), .Z(n9197) );
  XOR U12794 ( .A(DB[1167]), .B(DB[1152]), .Z(n9199) );
  AND U12795 ( .A(n718), .B(n9200), .Z(n9198) );
  XOR U12796 ( .A(n9201), .B(n9202), .Z(n9200) );
  XOR U12797 ( .A(DB[1152]), .B(DB[1137]), .Z(n9202) );
  AND U12798 ( .A(n722), .B(n9203), .Z(n9201) );
  XOR U12799 ( .A(n9204), .B(n9205), .Z(n9203) );
  XOR U12800 ( .A(DB[1137]), .B(DB[1122]), .Z(n9205) );
  AND U12801 ( .A(n726), .B(n9206), .Z(n9204) );
  XOR U12802 ( .A(n9207), .B(n9208), .Z(n9206) );
  XOR U12803 ( .A(DB[1122]), .B(DB[1107]), .Z(n9208) );
  AND U12804 ( .A(n730), .B(n9209), .Z(n9207) );
  XOR U12805 ( .A(n9210), .B(n9211), .Z(n9209) );
  XOR U12806 ( .A(DB[1107]), .B(DB[1092]), .Z(n9211) );
  AND U12807 ( .A(n734), .B(n9212), .Z(n9210) );
  XOR U12808 ( .A(n9213), .B(n9214), .Z(n9212) );
  XOR U12809 ( .A(DB[1092]), .B(DB[1077]), .Z(n9214) );
  AND U12810 ( .A(n738), .B(n9215), .Z(n9213) );
  XOR U12811 ( .A(n9216), .B(n9217), .Z(n9215) );
  XOR U12812 ( .A(DB[1077]), .B(DB[1062]), .Z(n9217) );
  AND U12813 ( .A(n742), .B(n9218), .Z(n9216) );
  XOR U12814 ( .A(n9219), .B(n9220), .Z(n9218) );
  XOR U12815 ( .A(DB[1062]), .B(DB[1047]), .Z(n9220) );
  AND U12816 ( .A(n746), .B(n9221), .Z(n9219) );
  XOR U12817 ( .A(n9222), .B(n9223), .Z(n9221) );
  XOR U12818 ( .A(DB[1047]), .B(DB[1032]), .Z(n9223) );
  AND U12819 ( .A(n750), .B(n9224), .Z(n9222) );
  XOR U12820 ( .A(n9225), .B(n9226), .Z(n9224) );
  XOR U12821 ( .A(DB[1032]), .B(DB[1017]), .Z(n9226) );
  AND U12822 ( .A(n754), .B(n9227), .Z(n9225) );
  XOR U12823 ( .A(n9228), .B(n9229), .Z(n9227) );
  XOR U12824 ( .A(DB[1017]), .B(DB[1002]), .Z(n9229) );
  AND U12825 ( .A(n758), .B(n9230), .Z(n9228) );
  XOR U12826 ( .A(n9231), .B(n9232), .Z(n9230) );
  XOR U12827 ( .A(DB[987]), .B(DB[1002]), .Z(n9232) );
  AND U12828 ( .A(n762), .B(n9233), .Z(n9231) );
  XOR U12829 ( .A(n9234), .B(n9235), .Z(n9233) );
  XOR U12830 ( .A(DB[987]), .B(DB[972]), .Z(n9235) );
  AND U12831 ( .A(n766), .B(n9236), .Z(n9234) );
  XOR U12832 ( .A(n9237), .B(n9238), .Z(n9236) );
  XOR U12833 ( .A(DB[972]), .B(DB[957]), .Z(n9238) );
  AND U12834 ( .A(n770), .B(n9239), .Z(n9237) );
  XOR U12835 ( .A(n9240), .B(n9241), .Z(n9239) );
  XOR U12836 ( .A(DB[957]), .B(DB[942]), .Z(n9241) );
  AND U12837 ( .A(n774), .B(n9242), .Z(n9240) );
  XOR U12838 ( .A(n9243), .B(n9244), .Z(n9242) );
  XOR U12839 ( .A(DB[942]), .B(DB[927]), .Z(n9244) );
  AND U12840 ( .A(n778), .B(n9245), .Z(n9243) );
  XOR U12841 ( .A(n9246), .B(n9247), .Z(n9245) );
  XOR U12842 ( .A(DB[927]), .B(DB[912]), .Z(n9247) );
  AND U12843 ( .A(n782), .B(n9248), .Z(n9246) );
  XOR U12844 ( .A(n9249), .B(n9250), .Z(n9248) );
  XOR U12845 ( .A(DB[912]), .B(DB[897]), .Z(n9250) );
  AND U12846 ( .A(n786), .B(n9251), .Z(n9249) );
  XOR U12847 ( .A(n9252), .B(n9253), .Z(n9251) );
  XOR U12848 ( .A(DB[897]), .B(DB[882]), .Z(n9253) );
  AND U12849 ( .A(n790), .B(n9254), .Z(n9252) );
  XOR U12850 ( .A(n9255), .B(n9256), .Z(n9254) );
  XOR U12851 ( .A(DB[882]), .B(DB[867]), .Z(n9256) );
  AND U12852 ( .A(n794), .B(n9257), .Z(n9255) );
  XOR U12853 ( .A(n9258), .B(n9259), .Z(n9257) );
  XOR U12854 ( .A(DB[867]), .B(DB[852]), .Z(n9259) );
  AND U12855 ( .A(n798), .B(n9260), .Z(n9258) );
  XOR U12856 ( .A(n9261), .B(n9262), .Z(n9260) );
  XOR U12857 ( .A(DB[852]), .B(DB[837]), .Z(n9262) );
  AND U12858 ( .A(n802), .B(n9263), .Z(n9261) );
  XOR U12859 ( .A(n9264), .B(n9265), .Z(n9263) );
  XOR U12860 ( .A(DB[837]), .B(DB[822]), .Z(n9265) );
  AND U12861 ( .A(n806), .B(n9266), .Z(n9264) );
  XOR U12862 ( .A(n9267), .B(n9268), .Z(n9266) );
  XOR U12863 ( .A(DB[822]), .B(DB[807]), .Z(n9268) );
  AND U12864 ( .A(n810), .B(n9269), .Z(n9267) );
  XOR U12865 ( .A(n9270), .B(n9271), .Z(n9269) );
  XOR U12866 ( .A(DB[807]), .B(DB[792]), .Z(n9271) );
  AND U12867 ( .A(n814), .B(n9272), .Z(n9270) );
  XOR U12868 ( .A(n9273), .B(n9274), .Z(n9272) );
  XOR U12869 ( .A(DB[792]), .B(DB[777]), .Z(n9274) );
  AND U12870 ( .A(n818), .B(n9275), .Z(n9273) );
  XOR U12871 ( .A(n9276), .B(n9277), .Z(n9275) );
  XOR U12872 ( .A(DB[777]), .B(DB[762]), .Z(n9277) );
  AND U12873 ( .A(n822), .B(n9278), .Z(n9276) );
  XOR U12874 ( .A(n9279), .B(n9280), .Z(n9278) );
  XOR U12875 ( .A(DB[762]), .B(DB[747]), .Z(n9280) );
  AND U12876 ( .A(n826), .B(n9281), .Z(n9279) );
  XOR U12877 ( .A(n9282), .B(n9283), .Z(n9281) );
  XOR U12878 ( .A(DB[747]), .B(DB[732]), .Z(n9283) );
  AND U12879 ( .A(n830), .B(n9284), .Z(n9282) );
  XOR U12880 ( .A(n9285), .B(n9286), .Z(n9284) );
  XOR U12881 ( .A(DB[732]), .B(DB[717]), .Z(n9286) );
  AND U12882 ( .A(n834), .B(n9287), .Z(n9285) );
  XOR U12883 ( .A(n9288), .B(n9289), .Z(n9287) );
  XOR U12884 ( .A(DB[717]), .B(DB[702]), .Z(n9289) );
  AND U12885 ( .A(n838), .B(n9290), .Z(n9288) );
  XOR U12886 ( .A(n9291), .B(n9292), .Z(n9290) );
  XOR U12887 ( .A(DB[702]), .B(DB[687]), .Z(n9292) );
  AND U12888 ( .A(n842), .B(n9293), .Z(n9291) );
  XOR U12889 ( .A(n9294), .B(n9295), .Z(n9293) );
  XOR U12890 ( .A(DB[687]), .B(DB[672]), .Z(n9295) );
  AND U12891 ( .A(n846), .B(n9296), .Z(n9294) );
  XOR U12892 ( .A(n9297), .B(n9298), .Z(n9296) );
  XOR U12893 ( .A(DB[672]), .B(DB[657]), .Z(n9298) );
  AND U12894 ( .A(n850), .B(n9299), .Z(n9297) );
  XOR U12895 ( .A(n9300), .B(n9301), .Z(n9299) );
  XOR U12896 ( .A(DB[657]), .B(DB[642]), .Z(n9301) );
  AND U12897 ( .A(n854), .B(n9302), .Z(n9300) );
  XOR U12898 ( .A(n9303), .B(n9304), .Z(n9302) );
  XOR U12899 ( .A(DB[642]), .B(DB[627]), .Z(n9304) );
  AND U12900 ( .A(n858), .B(n9305), .Z(n9303) );
  XOR U12901 ( .A(n9306), .B(n9307), .Z(n9305) );
  XOR U12902 ( .A(DB[627]), .B(DB[612]), .Z(n9307) );
  AND U12903 ( .A(n862), .B(n9308), .Z(n9306) );
  XOR U12904 ( .A(n9309), .B(n9310), .Z(n9308) );
  XOR U12905 ( .A(DB[612]), .B(DB[597]), .Z(n9310) );
  AND U12906 ( .A(n866), .B(n9311), .Z(n9309) );
  XOR U12907 ( .A(n9312), .B(n9313), .Z(n9311) );
  XOR U12908 ( .A(DB[597]), .B(DB[582]), .Z(n9313) );
  AND U12909 ( .A(n870), .B(n9314), .Z(n9312) );
  XOR U12910 ( .A(n9315), .B(n9316), .Z(n9314) );
  XOR U12911 ( .A(DB[582]), .B(DB[567]), .Z(n9316) );
  AND U12912 ( .A(n874), .B(n9317), .Z(n9315) );
  XOR U12913 ( .A(n9318), .B(n9319), .Z(n9317) );
  XOR U12914 ( .A(DB[567]), .B(DB[552]), .Z(n9319) );
  AND U12915 ( .A(n878), .B(n9320), .Z(n9318) );
  XOR U12916 ( .A(n9321), .B(n9322), .Z(n9320) );
  XOR U12917 ( .A(DB[552]), .B(DB[537]), .Z(n9322) );
  AND U12918 ( .A(n882), .B(n9323), .Z(n9321) );
  XOR U12919 ( .A(n9324), .B(n9325), .Z(n9323) );
  XOR U12920 ( .A(DB[537]), .B(DB[522]), .Z(n9325) );
  AND U12921 ( .A(n886), .B(n9326), .Z(n9324) );
  XOR U12922 ( .A(n9327), .B(n9328), .Z(n9326) );
  XOR U12923 ( .A(DB[522]), .B(DB[507]), .Z(n9328) );
  AND U12924 ( .A(n890), .B(n9329), .Z(n9327) );
  XOR U12925 ( .A(n9330), .B(n9331), .Z(n9329) );
  XOR U12926 ( .A(DB[507]), .B(DB[492]), .Z(n9331) );
  AND U12927 ( .A(n894), .B(n9332), .Z(n9330) );
  XOR U12928 ( .A(n9333), .B(n9334), .Z(n9332) );
  XOR U12929 ( .A(DB[492]), .B(DB[477]), .Z(n9334) );
  AND U12930 ( .A(n898), .B(n9335), .Z(n9333) );
  XOR U12931 ( .A(n9336), .B(n9337), .Z(n9335) );
  XOR U12932 ( .A(DB[477]), .B(DB[462]), .Z(n9337) );
  AND U12933 ( .A(n902), .B(n9338), .Z(n9336) );
  XOR U12934 ( .A(n9339), .B(n9340), .Z(n9338) );
  XOR U12935 ( .A(DB[462]), .B(DB[447]), .Z(n9340) );
  AND U12936 ( .A(n906), .B(n9341), .Z(n9339) );
  XOR U12937 ( .A(n9342), .B(n9343), .Z(n9341) );
  XOR U12938 ( .A(DB[447]), .B(DB[432]), .Z(n9343) );
  AND U12939 ( .A(n910), .B(n9344), .Z(n9342) );
  XOR U12940 ( .A(n9345), .B(n9346), .Z(n9344) );
  XOR U12941 ( .A(DB[432]), .B(DB[417]), .Z(n9346) );
  AND U12942 ( .A(n914), .B(n9347), .Z(n9345) );
  XOR U12943 ( .A(n9348), .B(n9349), .Z(n9347) );
  XOR U12944 ( .A(DB[417]), .B(DB[402]), .Z(n9349) );
  AND U12945 ( .A(n918), .B(n9350), .Z(n9348) );
  XOR U12946 ( .A(n9351), .B(n9352), .Z(n9350) );
  XOR U12947 ( .A(DB[402]), .B(DB[387]), .Z(n9352) );
  AND U12948 ( .A(n922), .B(n9353), .Z(n9351) );
  XOR U12949 ( .A(n9354), .B(n9355), .Z(n9353) );
  XOR U12950 ( .A(DB[387]), .B(DB[372]), .Z(n9355) );
  AND U12951 ( .A(n926), .B(n9356), .Z(n9354) );
  XOR U12952 ( .A(n9357), .B(n9358), .Z(n9356) );
  XOR U12953 ( .A(DB[372]), .B(DB[357]), .Z(n9358) );
  AND U12954 ( .A(n930), .B(n9359), .Z(n9357) );
  XOR U12955 ( .A(n9360), .B(n9361), .Z(n9359) );
  XOR U12956 ( .A(DB[357]), .B(DB[342]), .Z(n9361) );
  AND U12957 ( .A(n934), .B(n9362), .Z(n9360) );
  XOR U12958 ( .A(n9363), .B(n9364), .Z(n9362) );
  XOR U12959 ( .A(DB[342]), .B(DB[327]), .Z(n9364) );
  AND U12960 ( .A(n938), .B(n9365), .Z(n9363) );
  XOR U12961 ( .A(n9366), .B(n9367), .Z(n9365) );
  XOR U12962 ( .A(DB[327]), .B(DB[312]), .Z(n9367) );
  AND U12963 ( .A(n942), .B(n9368), .Z(n9366) );
  XOR U12964 ( .A(n9369), .B(n9370), .Z(n9368) );
  XOR U12965 ( .A(DB[312]), .B(DB[297]), .Z(n9370) );
  AND U12966 ( .A(n946), .B(n9371), .Z(n9369) );
  XOR U12967 ( .A(n9372), .B(n9373), .Z(n9371) );
  XOR U12968 ( .A(DB[297]), .B(DB[282]), .Z(n9373) );
  AND U12969 ( .A(n950), .B(n9374), .Z(n9372) );
  XOR U12970 ( .A(n9375), .B(n9376), .Z(n9374) );
  XOR U12971 ( .A(DB[282]), .B(DB[267]), .Z(n9376) );
  AND U12972 ( .A(n954), .B(n9377), .Z(n9375) );
  XOR U12973 ( .A(n9378), .B(n9379), .Z(n9377) );
  XOR U12974 ( .A(DB[267]), .B(DB[252]), .Z(n9379) );
  AND U12975 ( .A(n958), .B(n9380), .Z(n9378) );
  XOR U12976 ( .A(n9381), .B(n9382), .Z(n9380) );
  XOR U12977 ( .A(DB[252]), .B(DB[237]), .Z(n9382) );
  AND U12978 ( .A(n962), .B(n9383), .Z(n9381) );
  XOR U12979 ( .A(n9384), .B(n9385), .Z(n9383) );
  XOR U12980 ( .A(DB[237]), .B(DB[222]), .Z(n9385) );
  AND U12981 ( .A(n966), .B(n9386), .Z(n9384) );
  XOR U12982 ( .A(n9387), .B(n9388), .Z(n9386) );
  XOR U12983 ( .A(DB[222]), .B(DB[207]), .Z(n9388) );
  AND U12984 ( .A(n970), .B(n9389), .Z(n9387) );
  XOR U12985 ( .A(n9390), .B(n9391), .Z(n9389) );
  XOR U12986 ( .A(DB[207]), .B(DB[192]), .Z(n9391) );
  AND U12987 ( .A(n974), .B(n9392), .Z(n9390) );
  XOR U12988 ( .A(n9393), .B(n9394), .Z(n9392) );
  XOR U12989 ( .A(DB[192]), .B(DB[177]), .Z(n9394) );
  AND U12990 ( .A(n978), .B(n9395), .Z(n9393) );
  XOR U12991 ( .A(n9396), .B(n9397), .Z(n9395) );
  XOR U12992 ( .A(DB[177]), .B(DB[162]), .Z(n9397) );
  AND U12993 ( .A(n982), .B(n9398), .Z(n9396) );
  XOR U12994 ( .A(n9399), .B(n9400), .Z(n9398) );
  XOR U12995 ( .A(DB[162]), .B(DB[147]), .Z(n9400) );
  AND U12996 ( .A(n986), .B(n9401), .Z(n9399) );
  XOR U12997 ( .A(n9402), .B(n9403), .Z(n9401) );
  XOR U12998 ( .A(DB[147]), .B(DB[132]), .Z(n9403) );
  AND U12999 ( .A(n990), .B(n9404), .Z(n9402) );
  XOR U13000 ( .A(n9405), .B(n9406), .Z(n9404) );
  XOR U13001 ( .A(DB[132]), .B(DB[117]), .Z(n9406) );
  AND U13002 ( .A(n994), .B(n9407), .Z(n9405) );
  XOR U13003 ( .A(n9408), .B(n9409), .Z(n9407) );
  XOR U13004 ( .A(DB[117]), .B(DB[102]), .Z(n9409) );
  AND U13005 ( .A(n998), .B(n9410), .Z(n9408) );
  XOR U13006 ( .A(n9411), .B(n9412), .Z(n9410) );
  XOR U13007 ( .A(DB[87]), .B(DB[102]), .Z(n9412) );
  AND U13008 ( .A(n1002), .B(n9413), .Z(n9411) );
  XOR U13009 ( .A(n9414), .B(n9415), .Z(n9413) );
  XOR U13010 ( .A(DB[87]), .B(DB[72]), .Z(n9415) );
  AND U13011 ( .A(n1006), .B(n9416), .Z(n9414) );
  XOR U13012 ( .A(n9417), .B(n9418), .Z(n9416) );
  XOR U13013 ( .A(DB[72]), .B(DB[57]), .Z(n9418) );
  AND U13014 ( .A(n1010), .B(n9419), .Z(n9417) );
  XOR U13015 ( .A(n9420), .B(n9421), .Z(n9419) );
  XOR U13016 ( .A(DB[57]), .B(DB[42]), .Z(n9421) );
  AND U13017 ( .A(n1014), .B(n9422), .Z(n9420) );
  XOR U13018 ( .A(n9423), .B(n9424), .Z(n9422) );
  XOR U13019 ( .A(DB[42]), .B(DB[27]), .Z(n9424) );
  AND U13020 ( .A(n1018), .B(n9425), .Z(n9423) );
  XOR U13021 ( .A(DB[27]), .B(DB[12]), .Z(n9425) );
  XOR U13022 ( .A(DB[3836]), .B(n9426), .Z(min_val_out[11]) );
  AND U13023 ( .A(n2), .B(n9427), .Z(n9426) );
  XOR U13024 ( .A(n9428), .B(n9429), .Z(n9427) );
  XOR U13025 ( .A(n9430), .B(n9431), .Z(n9429) );
  IV U13026 ( .A(DB[3836]), .Z(n9430) );
  AND U13027 ( .A(n6), .B(n9432), .Z(n9428) );
  XOR U13028 ( .A(n9433), .B(n9434), .Z(n9432) );
  XOR U13029 ( .A(DB[3821]), .B(DB[3806]), .Z(n9434) );
  AND U13030 ( .A(n10), .B(n9435), .Z(n9433) );
  XOR U13031 ( .A(n9436), .B(n9437), .Z(n9435) );
  XOR U13032 ( .A(DB[3806]), .B(DB[3791]), .Z(n9437) );
  AND U13033 ( .A(n14), .B(n9438), .Z(n9436) );
  XOR U13034 ( .A(n9439), .B(n9440), .Z(n9438) );
  XOR U13035 ( .A(DB[3791]), .B(DB[3776]), .Z(n9440) );
  AND U13036 ( .A(n18), .B(n9441), .Z(n9439) );
  XOR U13037 ( .A(n9442), .B(n9443), .Z(n9441) );
  XOR U13038 ( .A(DB[3776]), .B(DB[3761]), .Z(n9443) );
  AND U13039 ( .A(n22), .B(n9444), .Z(n9442) );
  XOR U13040 ( .A(n9445), .B(n9446), .Z(n9444) );
  XOR U13041 ( .A(DB[3761]), .B(DB[3746]), .Z(n9446) );
  AND U13042 ( .A(n26), .B(n9447), .Z(n9445) );
  XOR U13043 ( .A(n9448), .B(n9449), .Z(n9447) );
  XOR U13044 ( .A(DB[3746]), .B(DB[3731]), .Z(n9449) );
  AND U13045 ( .A(n30), .B(n9450), .Z(n9448) );
  XOR U13046 ( .A(n9451), .B(n9452), .Z(n9450) );
  XOR U13047 ( .A(DB[3731]), .B(DB[3716]), .Z(n9452) );
  AND U13048 ( .A(n34), .B(n9453), .Z(n9451) );
  XOR U13049 ( .A(n9454), .B(n9455), .Z(n9453) );
  XOR U13050 ( .A(DB[3716]), .B(DB[3701]), .Z(n9455) );
  AND U13051 ( .A(n38), .B(n9456), .Z(n9454) );
  XOR U13052 ( .A(n9457), .B(n9458), .Z(n9456) );
  XOR U13053 ( .A(DB[3701]), .B(DB[3686]), .Z(n9458) );
  AND U13054 ( .A(n42), .B(n9459), .Z(n9457) );
  XOR U13055 ( .A(n9460), .B(n9461), .Z(n9459) );
  XOR U13056 ( .A(DB[3686]), .B(DB[3671]), .Z(n9461) );
  AND U13057 ( .A(n46), .B(n9462), .Z(n9460) );
  XOR U13058 ( .A(n9463), .B(n9464), .Z(n9462) );
  XOR U13059 ( .A(DB[3671]), .B(DB[3656]), .Z(n9464) );
  AND U13060 ( .A(n50), .B(n9465), .Z(n9463) );
  XOR U13061 ( .A(n9466), .B(n9467), .Z(n9465) );
  XOR U13062 ( .A(DB[3656]), .B(DB[3641]), .Z(n9467) );
  AND U13063 ( .A(n54), .B(n9468), .Z(n9466) );
  XOR U13064 ( .A(n9469), .B(n9470), .Z(n9468) );
  XOR U13065 ( .A(DB[3641]), .B(DB[3626]), .Z(n9470) );
  AND U13066 ( .A(n58), .B(n9471), .Z(n9469) );
  XOR U13067 ( .A(n9472), .B(n9473), .Z(n9471) );
  XOR U13068 ( .A(DB[3626]), .B(DB[3611]), .Z(n9473) );
  AND U13069 ( .A(n62), .B(n9474), .Z(n9472) );
  XOR U13070 ( .A(n9475), .B(n9476), .Z(n9474) );
  XOR U13071 ( .A(DB[3611]), .B(DB[3596]), .Z(n9476) );
  AND U13072 ( .A(n66), .B(n9477), .Z(n9475) );
  XOR U13073 ( .A(n9478), .B(n9479), .Z(n9477) );
  XOR U13074 ( .A(DB[3596]), .B(DB[3581]), .Z(n9479) );
  AND U13075 ( .A(n70), .B(n9480), .Z(n9478) );
  XOR U13076 ( .A(n9481), .B(n9482), .Z(n9480) );
  XOR U13077 ( .A(DB[3581]), .B(DB[3566]), .Z(n9482) );
  AND U13078 ( .A(n74), .B(n9483), .Z(n9481) );
  XOR U13079 ( .A(n9484), .B(n9485), .Z(n9483) );
  XOR U13080 ( .A(DB[3566]), .B(DB[3551]), .Z(n9485) );
  AND U13081 ( .A(n78), .B(n9486), .Z(n9484) );
  XOR U13082 ( .A(n9487), .B(n9488), .Z(n9486) );
  XOR U13083 ( .A(DB[3551]), .B(DB[3536]), .Z(n9488) );
  AND U13084 ( .A(n82), .B(n9489), .Z(n9487) );
  XOR U13085 ( .A(n9490), .B(n9491), .Z(n9489) );
  XOR U13086 ( .A(DB[3536]), .B(DB[3521]), .Z(n9491) );
  AND U13087 ( .A(n86), .B(n9492), .Z(n9490) );
  XOR U13088 ( .A(n9493), .B(n9494), .Z(n9492) );
  XOR U13089 ( .A(DB[3521]), .B(DB[3506]), .Z(n9494) );
  AND U13090 ( .A(n90), .B(n9495), .Z(n9493) );
  XOR U13091 ( .A(n9496), .B(n9497), .Z(n9495) );
  XOR U13092 ( .A(DB[3506]), .B(DB[3491]), .Z(n9497) );
  AND U13093 ( .A(n94), .B(n9498), .Z(n9496) );
  XOR U13094 ( .A(n9499), .B(n9500), .Z(n9498) );
  XOR U13095 ( .A(DB[3491]), .B(DB[3476]), .Z(n9500) );
  AND U13096 ( .A(n98), .B(n9501), .Z(n9499) );
  XOR U13097 ( .A(n9502), .B(n9503), .Z(n9501) );
  XOR U13098 ( .A(DB[3476]), .B(DB[3461]), .Z(n9503) );
  AND U13099 ( .A(n102), .B(n9504), .Z(n9502) );
  XOR U13100 ( .A(n9505), .B(n9506), .Z(n9504) );
  XOR U13101 ( .A(DB[3461]), .B(DB[3446]), .Z(n9506) );
  AND U13102 ( .A(n106), .B(n9507), .Z(n9505) );
  XOR U13103 ( .A(n9508), .B(n9509), .Z(n9507) );
  XOR U13104 ( .A(DB[3446]), .B(DB[3431]), .Z(n9509) );
  AND U13105 ( .A(n110), .B(n9510), .Z(n9508) );
  XOR U13106 ( .A(n9511), .B(n9512), .Z(n9510) );
  XOR U13107 ( .A(DB[3431]), .B(DB[3416]), .Z(n9512) );
  AND U13108 ( .A(n114), .B(n9513), .Z(n9511) );
  XOR U13109 ( .A(n9514), .B(n9515), .Z(n9513) );
  XOR U13110 ( .A(DB[3416]), .B(DB[3401]), .Z(n9515) );
  AND U13111 ( .A(n118), .B(n9516), .Z(n9514) );
  XOR U13112 ( .A(n9517), .B(n9518), .Z(n9516) );
  XOR U13113 ( .A(DB[3401]), .B(DB[3386]), .Z(n9518) );
  AND U13114 ( .A(n122), .B(n9519), .Z(n9517) );
  XOR U13115 ( .A(n9520), .B(n9521), .Z(n9519) );
  XOR U13116 ( .A(DB[3386]), .B(DB[3371]), .Z(n9521) );
  AND U13117 ( .A(n126), .B(n9522), .Z(n9520) );
  XOR U13118 ( .A(n9523), .B(n9524), .Z(n9522) );
  XOR U13119 ( .A(DB[3371]), .B(DB[3356]), .Z(n9524) );
  AND U13120 ( .A(n130), .B(n9525), .Z(n9523) );
  XOR U13121 ( .A(n9526), .B(n9527), .Z(n9525) );
  XOR U13122 ( .A(DB[3356]), .B(DB[3341]), .Z(n9527) );
  AND U13123 ( .A(n134), .B(n9528), .Z(n9526) );
  XOR U13124 ( .A(n9529), .B(n9530), .Z(n9528) );
  XOR U13125 ( .A(DB[3341]), .B(DB[3326]), .Z(n9530) );
  AND U13126 ( .A(n138), .B(n9531), .Z(n9529) );
  XOR U13127 ( .A(n9532), .B(n9533), .Z(n9531) );
  XOR U13128 ( .A(DB[3326]), .B(DB[3311]), .Z(n9533) );
  AND U13129 ( .A(n142), .B(n9534), .Z(n9532) );
  XOR U13130 ( .A(n9535), .B(n9536), .Z(n9534) );
  XOR U13131 ( .A(DB[3311]), .B(DB[3296]), .Z(n9536) );
  AND U13132 ( .A(n146), .B(n9537), .Z(n9535) );
  XOR U13133 ( .A(n9538), .B(n9539), .Z(n9537) );
  XOR U13134 ( .A(DB[3296]), .B(DB[3281]), .Z(n9539) );
  AND U13135 ( .A(n150), .B(n9540), .Z(n9538) );
  XOR U13136 ( .A(n9541), .B(n9542), .Z(n9540) );
  XOR U13137 ( .A(DB[3281]), .B(DB[3266]), .Z(n9542) );
  AND U13138 ( .A(n154), .B(n9543), .Z(n9541) );
  XOR U13139 ( .A(n9544), .B(n9545), .Z(n9543) );
  XOR U13140 ( .A(DB[3266]), .B(DB[3251]), .Z(n9545) );
  AND U13141 ( .A(n158), .B(n9546), .Z(n9544) );
  XOR U13142 ( .A(n9547), .B(n9548), .Z(n9546) );
  XOR U13143 ( .A(DB[3251]), .B(DB[3236]), .Z(n9548) );
  AND U13144 ( .A(n162), .B(n9549), .Z(n9547) );
  XOR U13145 ( .A(n9550), .B(n9551), .Z(n9549) );
  XOR U13146 ( .A(DB[3236]), .B(DB[3221]), .Z(n9551) );
  AND U13147 ( .A(n166), .B(n9552), .Z(n9550) );
  XOR U13148 ( .A(n9553), .B(n9554), .Z(n9552) );
  XOR U13149 ( .A(DB[3221]), .B(DB[3206]), .Z(n9554) );
  AND U13150 ( .A(n170), .B(n9555), .Z(n9553) );
  XOR U13151 ( .A(n9556), .B(n9557), .Z(n9555) );
  XOR U13152 ( .A(DB[3206]), .B(DB[3191]), .Z(n9557) );
  AND U13153 ( .A(n174), .B(n9558), .Z(n9556) );
  XOR U13154 ( .A(n9559), .B(n9560), .Z(n9558) );
  XOR U13155 ( .A(DB[3191]), .B(DB[3176]), .Z(n9560) );
  AND U13156 ( .A(n178), .B(n9561), .Z(n9559) );
  XOR U13157 ( .A(n9562), .B(n9563), .Z(n9561) );
  XOR U13158 ( .A(DB[3176]), .B(DB[3161]), .Z(n9563) );
  AND U13159 ( .A(n182), .B(n9564), .Z(n9562) );
  XOR U13160 ( .A(n9565), .B(n9566), .Z(n9564) );
  XOR U13161 ( .A(DB[3161]), .B(DB[3146]), .Z(n9566) );
  AND U13162 ( .A(n186), .B(n9567), .Z(n9565) );
  XOR U13163 ( .A(n9568), .B(n9569), .Z(n9567) );
  XOR U13164 ( .A(DB[3146]), .B(DB[3131]), .Z(n9569) );
  AND U13165 ( .A(n190), .B(n9570), .Z(n9568) );
  XOR U13166 ( .A(n9571), .B(n9572), .Z(n9570) );
  XOR U13167 ( .A(DB[3131]), .B(DB[3116]), .Z(n9572) );
  AND U13168 ( .A(n194), .B(n9573), .Z(n9571) );
  XOR U13169 ( .A(n9574), .B(n9575), .Z(n9573) );
  XOR U13170 ( .A(DB[3116]), .B(DB[3101]), .Z(n9575) );
  AND U13171 ( .A(n198), .B(n9576), .Z(n9574) );
  XOR U13172 ( .A(n9577), .B(n9578), .Z(n9576) );
  XOR U13173 ( .A(DB[3101]), .B(DB[3086]), .Z(n9578) );
  AND U13174 ( .A(n202), .B(n9579), .Z(n9577) );
  XOR U13175 ( .A(n9580), .B(n9581), .Z(n9579) );
  XOR U13176 ( .A(DB[3086]), .B(DB[3071]), .Z(n9581) );
  AND U13177 ( .A(n206), .B(n9582), .Z(n9580) );
  XOR U13178 ( .A(n9583), .B(n9584), .Z(n9582) );
  XOR U13179 ( .A(DB[3071]), .B(DB[3056]), .Z(n9584) );
  AND U13180 ( .A(n210), .B(n9585), .Z(n9583) );
  XOR U13181 ( .A(n9586), .B(n9587), .Z(n9585) );
  XOR U13182 ( .A(DB[3056]), .B(DB[3041]), .Z(n9587) );
  AND U13183 ( .A(n214), .B(n9588), .Z(n9586) );
  XOR U13184 ( .A(n9589), .B(n9590), .Z(n9588) );
  XOR U13185 ( .A(DB[3041]), .B(DB[3026]), .Z(n9590) );
  AND U13186 ( .A(n218), .B(n9591), .Z(n9589) );
  XOR U13187 ( .A(n9592), .B(n9593), .Z(n9591) );
  XOR U13188 ( .A(DB[3026]), .B(DB[3011]), .Z(n9593) );
  AND U13189 ( .A(n222), .B(n9594), .Z(n9592) );
  XOR U13190 ( .A(n9595), .B(n9596), .Z(n9594) );
  XOR U13191 ( .A(DB[3011]), .B(DB[2996]), .Z(n9596) );
  AND U13192 ( .A(n226), .B(n9597), .Z(n9595) );
  XOR U13193 ( .A(n9598), .B(n9599), .Z(n9597) );
  XOR U13194 ( .A(DB[2996]), .B(DB[2981]), .Z(n9599) );
  AND U13195 ( .A(n230), .B(n9600), .Z(n9598) );
  XOR U13196 ( .A(n9601), .B(n9602), .Z(n9600) );
  XOR U13197 ( .A(DB[2981]), .B(DB[2966]), .Z(n9602) );
  AND U13198 ( .A(n234), .B(n9603), .Z(n9601) );
  XOR U13199 ( .A(n9604), .B(n9605), .Z(n9603) );
  XOR U13200 ( .A(DB[2966]), .B(DB[2951]), .Z(n9605) );
  AND U13201 ( .A(n238), .B(n9606), .Z(n9604) );
  XOR U13202 ( .A(n9607), .B(n9608), .Z(n9606) );
  XOR U13203 ( .A(DB[2951]), .B(DB[2936]), .Z(n9608) );
  AND U13204 ( .A(n242), .B(n9609), .Z(n9607) );
  XOR U13205 ( .A(n9610), .B(n9611), .Z(n9609) );
  XOR U13206 ( .A(DB[2936]), .B(DB[2921]), .Z(n9611) );
  AND U13207 ( .A(n246), .B(n9612), .Z(n9610) );
  XOR U13208 ( .A(n9613), .B(n9614), .Z(n9612) );
  XOR U13209 ( .A(DB[2921]), .B(DB[2906]), .Z(n9614) );
  AND U13210 ( .A(n250), .B(n9615), .Z(n9613) );
  XOR U13211 ( .A(n9616), .B(n9617), .Z(n9615) );
  XOR U13212 ( .A(DB[2906]), .B(DB[2891]), .Z(n9617) );
  AND U13213 ( .A(n254), .B(n9618), .Z(n9616) );
  XOR U13214 ( .A(n9619), .B(n9620), .Z(n9618) );
  XOR U13215 ( .A(DB[2891]), .B(DB[2876]), .Z(n9620) );
  AND U13216 ( .A(n258), .B(n9621), .Z(n9619) );
  XOR U13217 ( .A(n9622), .B(n9623), .Z(n9621) );
  XOR U13218 ( .A(DB[2876]), .B(DB[2861]), .Z(n9623) );
  AND U13219 ( .A(n262), .B(n9624), .Z(n9622) );
  XOR U13220 ( .A(n9625), .B(n9626), .Z(n9624) );
  XOR U13221 ( .A(DB[2861]), .B(DB[2846]), .Z(n9626) );
  AND U13222 ( .A(n266), .B(n9627), .Z(n9625) );
  XOR U13223 ( .A(n9628), .B(n9629), .Z(n9627) );
  XOR U13224 ( .A(DB[2846]), .B(DB[2831]), .Z(n9629) );
  AND U13225 ( .A(n270), .B(n9630), .Z(n9628) );
  XOR U13226 ( .A(n9631), .B(n9632), .Z(n9630) );
  XOR U13227 ( .A(DB[2831]), .B(DB[2816]), .Z(n9632) );
  AND U13228 ( .A(n274), .B(n9633), .Z(n9631) );
  XOR U13229 ( .A(n9634), .B(n9635), .Z(n9633) );
  XOR U13230 ( .A(DB[2816]), .B(DB[2801]), .Z(n9635) );
  AND U13231 ( .A(n278), .B(n9636), .Z(n9634) );
  XOR U13232 ( .A(n9637), .B(n9638), .Z(n9636) );
  XOR U13233 ( .A(DB[2801]), .B(DB[2786]), .Z(n9638) );
  AND U13234 ( .A(n282), .B(n9639), .Z(n9637) );
  XOR U13235 ( .A(n9640), .B(n9641), .Z(n9639) );
  XOR U13236 ( .A(DB[2786]), .B(DB[2771]), .Z(n9641) );
  AND U13237 ( .A(n286), .B(n9642), .Z(n9640) );
  XOR U13238 ( .A(n9643), .B(n9644), .Z(n9642) );
  XOR U13239 ( .A(DB[2771]), .B(DB[2756]), .Z(n9644) );
  AND U13240 ( .A(n290), .B(n9645), .Z(n9643) );
  XOR U13241 ( .A(n9646), .B(n9647), .Z(n9645) );
  XOR U13242 ( .A(DB[2756]), .B(DB[2741]), .Z(n9647) );
  AND U13243 ( .A(n294), .B(n9648), .Z(n9646) );
  XOR U13244 ( .A(n9649), .B(n9650), .Z(n9648) );
  XOR U13245 ( .A(DB[2741]), .B(DB[2726]), .Z(n9650) );
  AND U13246 ( .A(n298), .B(n9651), .Z(n9649) );
  XOR U13247 ( .A(n9652), .B(n9653), .Z(n9651) );
  XOR U13248 ( .A(DB[2726]), .B(DB[2711]), .Z(n9653) );
  AND U13249 ( .A(n302), .B(n9654), .Z(n9652) );
  XOR U13250 ( .A(n9655), .B(n9656), .Z(n9654) );
  XOR U13251 ( .A(DB[2711]), .B(DB[2696]), .Z(n9656) );
  AND U13252 ( .A(n306), .B(n9657), .Z(n9655) );
  XOR U13253 ( .A(n9658), .B(n9659), .Z(n9657) );
  XOR U13254 ( .A(DB[2696]), .B(DB[2681]), .Z(n9659) );
  AND U13255 ( .A(n310), .B(n9660), .Z(n9658) );
  XOR U13256 ( .A(n9661), .B(n9662), .Z(n9660) );
  XOR U13257 ( .A(DB[2681]), .B(DB[2666]), .Z(n9662) );
  AND U13258 ( .A(n314), .B(n9663), .Z(n9661) );
  XOR U13259 ( .A(n9664), .B(n9665), .Z(n9663) );
  XOR U13260 ( .A(DB[2666]), .B(DB[2651]), .Z(n9665) );
  AND U13261 ( .A(n318), .B(n9666), .Z(n9664) );
  XOR U13262 ( .A(n9667), .B(n9668), .Z(n9666) );
  XOR U13263 ( .A(DB[2651]), .B(DB[2636]), .Z(n9668) );
  AND U13264 ( .A(n322), .B(n9669), .Z(n9667) );
  XOR U13265 ( .A(n9670), .B(n9671), .Z(n9669) );
  XOR U13266 ( .A(DB[2636]), .B(DB[2621]), .Z(n9671) );
  AND U13267 ( .A(n326), .B(n9672), .Z(n9670) );
  XOR U13268 ( .A(n9673), .B(n9674), .Z(n9672) );
  XOR U13269 ( .A(DB[2621]), .B(DB[2606]), .Z(n9674) );
  AND U13270 ( .A(n330), .B(n9675), .Z(n9673) );
  XOR U13271 ( .A(n9676), .B(n9677), .Z(n9675) );
  XOR U13272 ( .A(DB[2606]), .B(DB[2591]), .Z(n9677) );
  AND U13273 ( .A(n334), .B(n9678), .Z(n9676) );
  XOR U13274 ( .A(n9679), .B(n9680), .Z(n9678) );
  XOR U13275 ( .A(DB[2591]), .B(DB[2576]), .Z(n9680) );
  AND U13276 ( .A(n338), .B(n9681), .Z(n9679) );
  XOR U13277 ( .A(n9682), .B(n9683), .Z(n9681) );
  XOR U13278 ( .A(DB[2576]), .B(DB[2561]), .Z(n9683) );
  AND U13279 ( .A(n342), .B(n9684), .Z(n9682) );
  XOR U13280 ( .A(n9685), .B(n9686), .Z(n9684) );
  XOR U13281 ( .A(DB[2561]), .B(DB[2546]), .Z(n9686) );
  AND U13282 ( .A(n346), .B(n9687), .Z(n9685) );
  XOR U13283 ( .A(n9688), .B(n9689), .Z(n9687) );
  XOR U13284 ( .A(DB[2546]), .B(DB[2531]), .Z(n9689) );
  AND U13285 ( .A(n350), .B(n9690), .Z(n9688) );
  XOR U13286 ( .A(n9691), .B(n9692), .Z(n9690) );
  XOR U13287 ( .A(DB[2531]), .B(DB[2516]), .Z(n9692) );
  AND U13288 ( .A(n354), .B(n9693), .Z(n9691) );
  XOR U13289 ( .A(n9694), .B(n9695), .Z(n9693) );
  XOR U13290 ( .A(DB[2516]), .B(DB[2501]), .Z(n9695) );
  AND U13291 ( .A(n358), .B(n9696), .Z(n9694) );
  XOR U13292 ( .A(n9697), .B(n9698), .Z(n9696) );
  XOR U13293 ( .A(DB[2501]), .B(DB[2486]), .Z(n9698) );
  AND U13294 ( .A(n362), .B(n9699), .Z(n9697) );
  XOR U13295 ( .A(n9700), .B(n9701), .Z(n9699) );
  XOR U13296 ( .A(DB[2486]), .B(DB[2471]), .Z(n9701) );
  AND U13297 ( .A(n366), .B(n9702), .Z(n9700) );
  XOR U13298 ( .A(n9703), .B(n9704), .Z(n9702) );
  XOR U13299 ( .A(DB[2471]), .B(DB[2456]), .Z(n9704) );
  AND U13300 ( .A(n370), .B(n9705), .Z(n9703) );
  XOR U13301 ( .A(n9706), .B(n9707), .Z(n9705) );
  XOR U13302 ( .A(DB[2456]), .B(DB[2441]), .Z(n9707) );
  AND U13303 ( .A(n374), .B(n9708), .Z(n9706) );
  XOR U13304 ( .A(n9709), .B(n9710), .Z(n9708) );
  XOR U13305 ( .A(DB[2441]), .B(DB[2426]), .Z(n9710) );
  AND U13306 ( .A(n378), .B(n9711), .Z(n9709) );
  XOR U13307 ( .A(n9712), .B(n9713), .Z(n9711) );
  XOR U13308 ( .A(DB[2426]), .B(DB[2411]), .Z(n9713) );
  AND U13309 ( .A(n382), .B(n9714), .Z(n9712) );
  XOR U13310 ( .A(n9715), .B(n9716), .Z(n9714) );
  XOR U13311 ( .A(DB[2411]), .B(DB[2396]), .Z(n9716) );
  AND U13312 ( .A(n386), .B(n9717), .Z(n9715) );
  XOR U13313 ( .A(n9718), .B(n9719), .Z(n9717) );
  XOR U13314 ( .A(DB[2396]), .B(DB[2381]), .Z(n9719) );
  AND U13315 ( .A(n390), .B(n9720), .Z(n9718) );
  XOR U13316 ( .A(n9721), .B(n9722), .Z(n9720) );
  XOR U13317 ( .A(DB[2381]), .B(DB[2366]), .Z(n9722) );
  AND U13318 ( .A(n394), .B(n9723), .Z(n9721) );
  XOR U13319 ( .A(n9724), .B(n9725), .Z(n9723) );
  XOR U13320 ( .A(DB[2366]), .B(DB[2351]), .Z(n9725) );
  AND U13321 ( .A(n398), .B(n9726), .Z(n9724) );
  XOR U13322 ( .A(n9727), .B(n9728), .Z(n9726) );
  XOR U13323 ( .A(DB[2351]), .B(DB[2336]), .Z(n9728) );
  AND U13324 ( .A(n402), .B(n9729), .Z(n9727) );
  XOR U13325 ( .A(n9730), .B(n9731), .Z(n9729) );
  XOR U13326 ( .A(DB[2336]), .B(DB[2321]), .Z(n9731) );
  AND U13327 ( .A(n406), .B(n9732), .Z(n9730) );
  XOR U13328 ( .A(n9733), .B(n9734), .Z(n9732) );
  XOR U13329 ( .A(DB[2321]), .B(DB[2306]), .Z(n9734) );
  AND U13330 ( .A(n410), .B(n9735), .Z(n9733) );
  XOR U13331 ( .A(n9736), .B(n9737), .Z(n9735) );
  XOR U13332 ( .A(DB[2306]), .B(DB[2291]), .Z(n9737) );
  AND U13333 ( .A(n414), .B(n9738), .Z(n9736) );
  XOR U13334 ( .A(n9739), .B(n9740), .Z(n9738) );
  XOR U13335 ( .A(DB[2291]), .B(DB[2276]), .Z(n9740) );
  AND U13336 ( .A(n418), .B(n9741), .Z(n9739) );
  XOR U13337 ( .A(n9742), .B(n9743), .Z(n9741) );
  XOR U13338 ( .A(DB[2276]), .B(DB[2261]), .Z(n9743) );
  AND U13339 ( .A(n422), .B(n9744), .Z(n9742) );
  XOR U13340 ( .A(n9745), .B(n9746), .Z(n9744) );
  XOR U13341 ( .A(DB[2261]), .B(DB[2246]), .Z(n9746) );
  AND U13342 ( .A(n426), .B(n9747), .Z(n9745) );
  XOR U13343 ( .A(n9748), .B(n9749), .Z(n9747) );
  XOR U13344 ( .A(DB[2246]), .B(DB[2231]), .Z(n9749) );
  AND U13345 ( .A(n430), .B(n9750), .Z(n9748) );
  XOR U13346 ( .A(n9751), .B(n9752), .Z(n9750) );
  XOR U13347 ( .A(DB[2231]), .B(DB[2216]), .Z(n9752) );
  AND U13348 ( .A(n434), .B(n9753), .Z(n9751) );
  XOR U13349 ( .A(n9754), .B(n9755), .Z(n9753) );
  XOR U13350 ( .A(DB[2216]), .B(DB[2201]), .Z(n9755) );
  AND U13351 ( .A(n438), .B(n9756), .Z(n9754) );
  XOR U13352 ( .A(n9757), .B(n9758), .Z(n9756) );
  XOR U13353 ( .A(DB[2201]), .B(DB[2186]), .Z(n9758) );
  AND U13354 ( .A(n442), .B(n9759), .Z(n9757) );
  XOR U13355 ( .A(n9760), .B(n9761), .Z(n9759) );
  XOR U13356 ( .A(DB[2186]), .B(DB[2171]), .Z(n9761) );
  AND U13357 ( .A(n446), .B(n9762), .Z(n9760) );
  XOR U13358 ( .A(n9763), .B(n9764), .Z(n9762) );
  XOR U13359 ( .A(DB[2171]), .B(DB[2156]), .Z(n9764) );
  AND U13360 ( .A(n450), .B(n9765), .Z(n9763) );
  XOR U13361 ( .A(n9766), .B(n9767), .Z(n9765) );
  XOR U13362 ( .A(DB[2156]), .B(DB[2141]), .Z(n9767) );
  AND U13363 ( .A(n454), .B(n9768), .Z(n9766) );
  XOR U13364 ( .A(n9769), .B(n9770), .Z(n9768) );
  XOR U13365 ( .A(DB[2141]), .B(DB[2126]), .Z(n9770) );
  AND U13366 ( .A(n458), .B(n9771), .Z(n9769) );
  XOR U13367 ( .A(n9772), .B(n9773), .Z(n9771) );
  XOR U13368 ( .A(DB[2126]), .B(DB[2111]), .Z(n9773) );
  AND U13369 ( .A(n462), .B(n9774), .Z(n9772) );
  XOR U13370 ( .A(n9775), .B(n9776), .Z(n9774) );
  XOR U13371 ( .A(DB[2111]), .B(DB[2096]), .Z(n9776) );
  AND U13372 ( .A(n466), .B(n9777), .Z(n9775) );
  XOR U13373 ( .A(n9778), .B(n9779), .Z(n9777) );
  XOR U13374 ( .A(DB[2096]), .B(DB[2081]), .Z(n9779) );
  AND U13375 ( .A(n470), .B(n9780), .Z(n9778) );
  XOR U13376 ( .A(n9781), .B(n9782), .Z(n9780) );
  XOR U13377 ( .A(DB[2081]), .B(DB[2066]), .Z(n9782) );
  AND U13378 ( .A(n474), .B(n9783), .Z(n9781) );
  XOR U13379 ( .A(n9784), .B(n9785), .Z(n9783) );
  XOR U13380 ( .A(DB[2066]), .B(DB[2051]), .Z(n9785) );
  AND U13381 ( .A(n478), .B(n9786), .Z(n9784) );
  XOR U13382 ( .A(n9787), .B(n9788), .Z(n9786) );
  XOR U13383 ( .A(DB[2051]), .B(DB[2036]), .Z(n9788) );
  AND U13384 ( .A(n482), .B(n9789), .Z(n9787) );
  XOR U13385 ( .A(n9790), .B(n9791), .Z(n9789) );
  XOR U13386 ( .A(DB[2036]), .B(DB[2021]), .Z(n9791) );
  AND U13387 ( .A(n486), .B(n9792), .Z(n9790) );
  XOR U13388 ( .A(n9793), .B(n9794), .Z(n9792) );
  XOR U13389 ( .A(DB[2021]), .B(DB[2006]), .Z(n9794) );
  AND U13390 ( .A(n490), .B(n9795), .Z(n9793) );
  XOR U13391 ( .A(n9796), .B(n9797), .Z(n9795) );
  XOR U13392 ( .A(DB[2006]), .B(DB[1991]), .Z(n9797) );
  AND U13393 ( .A(n494), .B(n9798), .Z(n9796) );
  XOR U13394 ( .A(n9799), .B(n9800), .Z(n9798) );
  XOR U13395 ( .A(DB[1991]), .B(DB[1976]), .Z(n9800) );
  AND U13396 ( .A(n498), .B(n9801), .Z(n9799) );
  XOR U13397 ( .A(n9802), .B(n9803), .Z(n9801) );
  XOR U13398 ( .A(DB[1976]), .B(DB[1961]), .Z(n9803) );
  AND U13399 ( .A(n502), .B(n9804), .Z(n9802) );
  XOR U13400 ( .A(n9805), .B(n9806), .Z(n9804) );
  XOR U13401 ( .A(DB[1961]), .B(DB[1946]), .Z(n9806) );
  AND U13402 ( .A(n506), .B(n9807), .Z(n9805) );
  XOR U13403 ( .A(n9808), .B(n9809), .Z(n9807) );
  XOR U13404 ( .A(DB[1946]), .B(DB[1931]), .Z(n9809) );
  AND U13405 ( .A(n510), .B(n9810), .Z(n9808) );
  XOR U13406 ( .A(n9811), .B(n9812), .Z(n9810) );
  XOR U13407 ( .A(DB[1931]), .B(DB[1916]), .Z(n9812) );
  AND U13408 ( .A(n514), .B(n9813), .Z(n9811) );
  XOR U13409 ( .A(n9814), .B(n9815), .Z(n9813) );
  XOR U13410 ( .A(DB[1916]), .B(DB[1901]), .Z(n9815) );
  AND U13411 ( .A(n518), .B(n9816), .Z(n9814) );
  XOR U13412 ( .A(n9817), .B(n9818), .Z(n9816) );
  XOR U13413 ( .A(DB[1901]), .B(DB[1886]), .Z(n9818) );
  AND U13414 ( .A(n522), .B(n9819), .Z(n9817) );
  XOR U13415 ( .A(n9820), .B(n9821), .Z(n9819) );
  XOR U13416 ( .A(DB[1886]), .B(DB[1871]), .Z(n9821) );
  AND U13417 ( .A(n526), .B(n9822), .Z(n9820) );
  XOR U13418 ( .A(n9823), .B(n9824), .Z(n9822) );
  XOR U13419 ( .A(DB[1871]), .B(DB[1856]), .Z(n9824) );
  AND U13420 ( .A(n530), .B(n9825), .Z(n9823) );
  XOR U13421 ( .A(n9826), .B(n9827), .Z(n9825) );
  XOR U13422 ( .A(DB[1856]), .B(DB[1841]), .Z(n9827) );
  AND U13423 ( .A(n534), .B(n9828), .Z(n9826) );
  XOR U13424 ( .A(n9829), .B(n9830), .Z(n9828) );
  XOR U13425 ( .A(DB[1841]), .B(DB[1826]), .Z(n9830) );
  AND U13426 ( .A(n538), .B(n9831), .Z(n9829) );
  XOR U13427 ( .A(n9832), .B(n9833), .Z(n9831) );
  XOR U13428 ( .A(DB[1826]), .B(DB[1811]), .Z(n9833) );
  AND U13429 ( .A(n542), .B(n9834), .Z(n9832) );
  XOR U13430 ( .A(n9835), .B(n9836), .Z(n9834) );
  XOR U13431 ( .A(DB[1811]), .B(DB[1796]), .Z(n9836) );
  AND U13432 ( .A(n546), .B(n9837), .Z(n9835) );
  XOR U13433 ( .A(n9838), .B(n9839), .Z(n9837) );
  XOR U13434 ( .A(DB[1796]), .B(DB[1781]), .Z(n9839) );
  AND U13435 ( .A(n550), .B(n9840), .Z(n9838) );
  XOR U13436 ( .A(n9841), .B(n9842), .Z(n9840) );
  XOR U13437 ( .A(DB[1781]), .B(DB[1766]), .Z(n9842) );
  AND U13438 ( .A(n554), .B(n9843), .Z(n9841) );
  XOR U13439 ( .A(n9844), .B(n9845), .Z(n9843) );
  XOR U13440 ( .A(DB[1766]), .B(DB[1751]), .Z(n9845) );
  AND U13441 ( .A(n558), .B(n9846), .Z(n9844) );
  XOR U13442 ( .A(n9847), .B(n9848), .Z(n9846) );
  XOR U13443 ( .A(DB[1751]), .B(DB[1736]), .Z(n9848) );
  AND U13444 ( .A(n562), .B(n9849), .Z(n9847) );
  XOR U13445 ( .A(n9850), .B(n9851), .Z(n9849) );
  XOR U13446 ( .A(DB[1736]), .B(DB[1721]), .Z(n9851) );
  AND U13447 ( .A(n566), .B(n9852), .Z(n9850) );
  XOR U13448 ( .A(n9853), .B(n9854), .Z(n9852) );
  XOR U13449 ( .A(DB[1721]), .B(DB[1706]), .Z(n9854) );
  AND U13450 ( .A(n570), .B(n9855), .Z(n9853) );
  XOR U13451 ( .A(n9856), .B(n9857), .Z(n9855) );
  XOR U13452 ( .A(DB[1706]), .B(DB[1691]), .Z(n9857) );
  AND U13453 ( .A(n574), .B(n9858), .Z(n9856) );
  XOR U13454 ( .A(n9859), .B(n9860), .Z(n9858) );
  XOR U13455 ( .A(DB[1691]), .B(DB[1676]), .Z(n9860) );
  AND U13456 ( .A(n578), .B(n9861), .Z(n9859) );
  XOR U13457 ( .A(n9862), .B(n9863), .Z(n9861) );
  XOR U13458 ( .A(DB[1676]), .B(DB[1661]), .Z(n9863) );
  AND U13459 ( .A(n582), .B(n9864), .Z(n9862) );
  XOR U13460 ( .A(n9865), .B(n9866), .Z(n9864) );
  XOR U13461 ( .A(DB[1661]), .B(DB[1646]), .Z(n9866) );
  AND U13462 ( .A(n586), .B(n9867), .Z(n9865) );
  XOR U13463 ( .A(n9868), .B(n9869), .Z(n9867) );
  XOR U13464 ( .A(DB[1646]), .B(DB[1631]), .Z(n9869) );
  AND U13465 ( .A(n590), .B(n9870), .Z(n9868) );
  XOR U13466 ( .A(n9871), .B(n9872), .Z(n9870) );
  XOR U13467 ( .A(DB[1631]), .B(DB[1616]), .Z(n9872) );
  AND U13468 ( .A(n594), .B(n9873), .Z(n9871) );
  XOR U13469 ( .A(n9874), .B(n9875), .Z(n9873) );
  XOR U13470 ( .A(DB[1616]), .B(DB[1601]), .Z(n9875) );
  AND U13471 ( .A(n598), .B(n9876), .Z(n9874) );
  XOR U13472 ( .A(n9877), .B(n9878), .Z(n9876) );
  XOR U13473 ( .A(DB[1601]), .B(DB[1586]), .Z(n9878) );
  AND U13474 ( .A(n602), .B(n9879), .Z(n9877) );
  XOR U13475 ( .A(n9880), .B(n9881), .Z(n9879) );
  XOR U13476 ( .A(DB[1586]), .B(DB[1571]), .Z(n9881) );
  AND U13477 ( .A(n606), .B(n9882), .Z(n9880) );
  XOR U13478 ( .A(n9883), .B(n9884), .Z(n9882) );
  XOR U13479 ( .A(DB[1571]), .B(DB[1556]), .Z(n9884) );
  AND U13480 ( .A(n610), .B(n9885), .Z(n9883) );
  XOR U13481 ( .A(n9886), .B(n9887), .Z(n9885) );
  XOR U13482 ( .A(DB[1556]), .B(DB[1541]), .Z(n9887) );
  AND U13483 ( .A(n614), .B(n9888), .Z(n9886) );
  XOR U13484 ( .A(n9889), .B(n9890), .Z(n9888) );
  XOR U13485 ( .A(DB[1541]), .B(DB[1526]), .Z(n9890) );
  AND U13486 ( .A(n618), .B(n9891), .Z(n9889) );
  XOR U13487 ( .A(n9892), .B(n9893), .Z(n9891) );
  XOR U13488 ( .A(DB[1526]), .B(DB[1511]), .Z(n9893) );
  AND U13489 ( .A(n622), .B(n9894), .Z(n9892) );
  XOR U13490 ( .A(n9895), .B(n9896), .Z(n9894) );
  XOR U13491 ( .A(DB[1511]), .B(DB[1496]), .Z(n9896) );
  AND U13492 ( .A(n626), .B(n9897), .Z(n9895) );
  XOR U13493 ( .A(n9898), .B(n9899), .Z(n9897) );
  XOR U13494 ( .A(DB[1496]), .B(DB[1481]), .Z(n9899) );
  AND U13495 ( .A(n630), .B(n9900), .Z(n9898) );
  XOR U13496 ( .A(n9901), .B(n9902), .Z(n9900) );
  XOR U13497 ( .A(DB[1481]), .B(DB[1466]), .Z(n9902) );
  AND U13498 ( .A(n634), .B(n9903), .Z(n9901) );
  XOR U13499 ( .A(n9904), .B(n9905), .Z(n9903) );
  XOR U13500 ( .A(DB[1466]), .B(DB[1451]), .Z(n9905) );
  AND U13501 ( .A(n638), .B(n9906), .Z(n9904) );
  XOR U13502 ( .A(n9907), .B(n9908), .Z(n9906) );
  XOR U13503 ( .A(DB[1451]), .B(DB[1436]), .Z(n9908) );
  AND U13504 ( .A(n642), .B(n9909), .Z(n9907) );
  XOR U13505 ( .A(n9910), .B(n9911), .Z(n9909) );
  XOR U13506 ( .A(DB[1436]), .B(DB[1421]), .Z(n9911) );
  AND U13507 ( .A(n646), .B(n9912), .Z(n9910) );
  XOR U13508 ( .A(n9913), .B(n9914), .Z(n9912) );
  XOR U13509 ( .A(DB[1421]), .B(DB[1406]), .Z(n9914) );
  AND U13510 ( .A(n650), .B(n9915), .Z(n9913) );
  XOR U13511 ( .A(n9916), .B(n9917), .Z(n9915) );
  XOR U13512 ( .A(DB[1406]), .B(DB[1391]), .Z(n9917) );
  AND U13513 ( .A(n654), .B(n9918), .Z(n9916) );
  XOR U13514 ( .A(n9919), .B(n9920), .Z(n9918) );
  XOR U13515 ( .A(DB[1391]), .B(DB[1376]), .Z(n9920) );
  AND U13516 ( .A(n658), .B(n9921), .Z(n9919) );
  XOR U13517 ( .A(n9922), .B(n9923), .Z(n9921) );
  XOR U13518 ( .A(DB[1376]), .B(DB[1361]), .Z(n9923) );
  AND U13519 ( .A(n662), .B(n9924), .Z(n9922) );
  XOR U13520 ( .A(n9925), .B(n9926), .Z(n9924) );
  XOR U13521 ( .A(DB[1361]), .B(DB[1346]), .Z(n9926) );
  AND U13522 ( .A(n666), .B(n9927), .Z(n9925) );
  XOR U13523 ( .A(n9928), .B(n9929), .Z(n9927) );
  XOR U13524 ( .A(DB[1346]), .B(DB[1331]), .Z(n9929) );
  AND U13525 ( .A(n670), .B(n9930), .Z(n9928) );
  XOR U13526 ( .A(n9931), .B(n9932), .Z(n9930) );
  XOR U13527 ( .A(DB[1331]), .B(DB[1316]), .Z(n9932) );
  AND U13528 ( .A(n674), .B(n9933), .Z(n9931) );
  XOR U13529 ( .A(n9934), .B(n9935), .Z(n9933) );
  XOR U13530 ( .A(DB[1316]), .B(DB[1301]), .Z(n9935) );
  AND U13531 ( .A(n678), .B(n9936), .Z(n9934) );
  XOR U13532 ( .A(n9937), .B(n9938), .Z(n9936) );
  XOR U13533 ( .A(DB[1301]), .B(DB[1286]), .Z(n9938) );
  AND U13534 ( .A(n682), .B(n9939), .Z(n9937) );
  XOR U13535 ( .A(n9940), .B(n9941), .Z(n9939) );
  XOR U13536 ( .A(DB[1286]), .B(DB[1271]), .Z(n9941) );
  AND U13537 ( .A(n686), .B(n9942), .Z(n9940) );
  XOR U13538 ( .A(n9943), .B(n9944), .Z(n9942) );
  XOR U13539 ( .A(DB[1271]), .B(DB[1256]), .Z(n9944) );
  AND U13540 ( .A(n690), .B(n9945), .Z(n9943) );
  XOR U13541 ( .A(n9946), .B(n9947), .Z(n9945) );
  XOR U13542 ( .A(DB[1256]), .B(DB[1241]), .Z(n9947) );
  AND U13543 ( .A(n694), .B(n9948), .Z(n9946) );
  XOR U13544 ( .A(n9949), .B(n9950), .Z(n9948) );
  XOR U13545 ( .A(DB[1241]), .B(DB[1226]), .Z(n9950) );
  AND U13546 ( .A(n698), .B(n9951), .Z(n9949) );
  XOR U13547 ( .A(n9952), .B(n9953), .Z(n9951) );
  XOR U13548 ( .A(DB[1226]), .B(DB[1211]), .Z(n9953) );
  AND U13549 ( .A(n702), .B(n9954), .Z(n9952) );
  XOR U13550 ( .A(n9955), .B(n9956), .Z(n9954) );
  XOR U13551 ( .A(DB[1211]), .B(DB[1196]), .Z(n9956) );
  AND U13552 ( .A(n706), .B(n9957), .Z(n9955) );
  XOR U13553 ( .A(n9958), .B(n9959), .Z(n9957) );
  XOR U13554 ( .A(DB[1196]), .B(DB[1181]), .Z(n9959) );
  AND U13555 ( .A(n710), .B(n9960), .Z(n9958) );
  XOR U13556 ( .A(n9961), .B(n9962), .Z(n9960) );
  XOR U13557 ( .A(DB[1181]), .B(DB[1166]), .Z(n9962) );
  AND U13558 ( .A(n714), .B(n9963), .Z(n9961) );
  XOR U13559 ( .A(n9964), .B(n9965), .Z(n9963) );
  XOR U13560 ( .A(DB[1166]), .B(DB[1151]), .Z(n9965) );
  AND U13561 ( .A(n718), .B(n9966), .Z(n9964) );
  XOR U13562 ( .A(n9967), .B(n9968), .Z(n9966) );
  XOR U13563 ( .A(DB[1151]), .B(DB[1136]), .Z(n9968) );
  AND U13564 ( .A(n722), .B(n9969), .Z(n9967) );
  XOR U13565 ( .A(n9970), .B(n9971), .Z(n9969) );
  XOR U13566 ( .A(DB[1136]), .B(DB[1121]), .Z(n9971) );
  AND U13567 ( .A(n726), .B(n9972), .Z(n9970) );
  XOR U13568 ( .A(n9973), .B(n9974), .Z(n9972) );
  XOR U13569 ( .A(DB[1121]), .B(DB[1106]), .Z(n9974) );
  AND U13570 ( .A(n730), .B(n9975), .Z(n9973) );
  XOR U13571 ( .A(n9976), .B(n9977), .Z(n9975) );
  XOR U13572 ( .A(DB[1106]), .B(DB[1091]), .Z(n9977) );
  AND U13573 ( .A(n734), .B(n9978), .Z(n9976) );
  XOR U13574 ( .A(n9979), .B(n9980), .Z(n9978) );
  XOR U13575 ( .A(DB[1091]), .B(DB[1076]), .Z(n9980) );
  AND U13576 ( .A(n738), .B(n9981), .Z(n9979) );
  XOR U13577 ( .A(n9982), .B(n9983), .Z(n9981) );
  XOR U13578 ( .A(DB[1076]), .B(DB[1061]), .Z(n9983) );
  AND U13579 ( .A(n742), .B(n9984), .Z(n9982) );
  XOR U13580 ( .A(n9985), .B(n9986), .Z(n9984) );
  XOR U13581 ( .A(DB[1061]), .B(DB[1046]), .Z(n9986) );
  AND U13582 ( .A(n746), .B(n9987), .Z(n9985) );
  XOR U13583 ( .A(n9988), .B(n9989), .Z(n9987) );
  XOR U13584 ( .A(DB[1046]), .B(DB[1031]), .Z(n9989) );
  AND U13585 ( .A(n750), .B(n9990), .Z(n9988) );
  XOR U13586 ( .A(n9991), .B(n9992), .Z(n9990) );
  XOR U13587 ( .A(DB[1031]), .B(DB[1016]), .Z(n9992) );
  AND U13588 ( .A(n754), .B(n9993), .Z(n9991) );
  XOR U13589 ( .A(n9994), .B(n9995), .Z(n9993) );
  XOR U13590 ( .A(DB[1016]), .B(DB[1001]), .Z(n9995) );
  AND U13591 ( .A(n758), .B(n9996), .Z(n9994) );
  XOR U13592 ( .A(n9997), .B(n9998), .Z(n9996) );
  XOR U13593 ( .A(DB[986]), .B(DB[1001]), .Z(n9998) );
  AND U13594 ( .A(n762), .B(n9999), .Z(n9997) );
  XOR U13595 ( .A(n10000), .B(n10001), .Z(n9999) );
  XOR U13596 ( .A(DB[986]), .B(DB[971]), .Z(n10001) );
  AND U13597 ( .A(n766), .B(n10002), .Z(n10000) );
  XOR U13598 ( .A(n10003), .B(n10004), .Z(n10002) );
  XOR U13599 ( .A(DB[971]), .B(DB[956]), .Z(n10004) );
  AND U13600 ( .A(n770), .B(n10005), .Z(n10003) );
  XOR U13601 ( .A(n10006), .B(n10007), .Z(n10005) );
  XOR U13602 ( .A(DB[956]), .B(DB[941]), .Z(n10007) );
  AND U13603 ( .A(n774), .B(n10008), .Z(n10006) );
  XOR U13604 ( .A(n10009), .B(n10010), .Z(n10008) );
  XOR U13605 ( .A(DB[941]), .B(DB[926]), .Z(n10010) );
  AND U13606 ( .A(n778), .B(n10011), .Z(n10009) );
  XOR U13607 ( .A(n10012), .B(n10013), .Z(n10011) );
  XOR U13608 ( .A(DB[926]), .B(DB[911]), .Z(n10013) );
  AND U13609 ( .A(n782), .B(n10014), .Z(n10012) );
  XOR U13610 ( .A(n10015), .B(n10016), .Z(n10014) );
  XOR U13611 ( .A(DB[911]), .B(DB[896]), .Z(n10016) );
  AND U13612 ( .A(n786), .B(n10017), .Z(n10015) );
  XOR U13613 ( .A(n10018), .B(n10019), .Z(n10017) );
  XOR U13614 ( .A(DB[896]), .B(DB[881]), .Z(n10019) );
  AND U13615 ( .A(n790), .B(n10020), .Z(n10018) );
  XOR U13616 ( .A(n10021), .B(n10022), .Z(n10020) );
  XOR U13617 ( .A(DB[881]), .B(DB[866]), .Z(n10022) );
  AND U13618 ( .A(n794), .B(n10023), .Z(n10021) );
  XOR U13619 ( .A(n10024), .B(n10025), .Z(n10023) );
  XOR U13620 ( .A(DB[866]), .B(DB[851]), .Z(n10025) );
  AND U13621 ( .A(n798), .B(n10026), .Z(n10024) );
  XOR U13622 ( .A(n10027), .B(n10028), .Z(n10026) );
  XOR U13623 ( .A(DB[851]), .B(DB[836]), .Z(n10028) );
  AND U13624 ( .A(n802), .B(n10029), .Z(n10027) );
  XOR U13625 ( .A(n10030), .B(n10031), .Z(n10029) );
  XOR U13626 ( .A(DB[836]), .B(DB[821]), .Z(n10031) );
  AND U13627 ( .A(n806), .B(n10032), .Z(n10030) );
  XOR U13628 ( .A(n10033), .B(n10034), .Z(n10032) );
  XOR U13629 ( .A(DB[821]), .B(DB[806]), .Z(n10034) );
  AND U13630 ( .A(n810), .B(n10035), .Z(n10033) );
  XOR U13631 ( .A(n10036), .B(n10037), .Z(n10035) );
  XOR U13632 ( .A(DB[806]), .B(DB[791]), .Z(n10037) );
  AND U13633 ( .A(n814), .B(n10038), .Z(n10036) );
  XOR U13634 ( .A(n10039), .B(n10040), .Z(n10038) );
  XOR U13635 ( .A(DB[791]), .B(DB[776]), .Z(n10040) );
  AND U13636 ( .A(n818), .B(n10041), .Z(n10039) );
  XOR U13637 ( .A(n10042), .B(n10043), .Z(n10041) );
  XOR U13638 ( .A(DB[776]), .B(DB[761]), .Z(n10043) );
  AND U13639 ( .A(n822), .B(n10044), .Z(n10042) );
  XOR U13640 ( .A(n10045), .B(n10046), .Z(n10044) );
  XOR U13641 ( .A(DB[761]), .B(DB[746]), .Z(n10046) );
  AND U13642 ( .A(n826), .B(n10047), .Z(n10045) );
  XOR U13643 ( .A(n10048), .B(n10049), .Z(n10047) );
  XOR U13644 ( .A(DB[746]), .B(DB[731]), .Z(n10049) );
  AND U13645 ( .A(n830), .B(n10050), .Z(n10048) );
  XOR U13646 ( .A(n10051), .B(n10052), .Z(n10050) );
  XOR U13647 ( .A(DB[731]), .B(DB[716]), .Z(n10052) );
  AND U13648 ( .A(n834), .B(n10053), .Z(n10051) );
  XOR U13649 ( .A(n10054), .B(n10055), .Z(n10053) );
  XOR U13650 ( .A(DB[716]), .B(DB[701]), .Z(n10055) );
  AND U13651 ( .A(n838), .B(n10056), .Z(n10054) );
  XOR U13652 ( .A(n10057), .B(n10058), .Z(n10056) );
  XOR U13653 ( .A(DB[701]), .B(DB[686]), .Z(n10058) );
  AND U13654 ( .A(n842), .B(n10059), .Z(n10057) );
  XOR U13655 ( .A(n10060), .B(n10061), .Z(n10059) );
  XOR U13656 ( .A(DB[686]), .B(DB[671]), .Z(n10061) );
  AND U13657 ( .A(n846), .B(n10062), .Z(n10060) );
  XOR U13658 ( .A(n10063), .B(n10064), .Z(n10062) );
  XOR U13659 ( .A(DB[671]), .B(DB[656]), .Z(n10064) );
  AND U13660 ( .A(n850), .B(n10065), .Z(n10063) );
  XOR U13661 ( .A(n10066), .B(n10067), .Z(n10065) );
  XOR U13662 ( .A(DB[656]), .B(DB[641]), .Z(n10067) );
  AND U13663 ( .A(n854), .B(n10068), .Z(n10066) );
  XOR U13664 ( .A(n10069), .B(n10070), .Z(n10068) );
  XOR U13665 ( .A(DB[641]), .B(DB[626]), .Z(n10070) );
  AND U13666 ( .A(n858), .B(n10071), .Z(n10069) );
  XOR U13667 ( .A(n10072), .B(n10073), .Z(n10071) );
  XOR U13668 ( .A(DB[626]), .B(DB[611]), .Z(n10073) );
  AND U13669 ( .A(n862), .B(n10074), .Z(n10072) );
  XOR U13670 ( .A(n10075), .B(n10076), .Z(n10074) );
  XOR U13671 ( .A(DB[611]), .B(DB[596]), .Z(n10076) );
  AND U13672 ( .A(n866), .B(n10077), .Z(n10075) );
  XOR U13673 ( .A(n10078), .B(n10079), .Z(n10077) );
  XOR U13674 ( .A(DB[596]), .B(DB[581]), .Z(n10079) );
  AND U13675 ( .A(n870), .B(n10080), .Z(n10078) );
  XOR U13676 ( .A(n10081), .B(n10082), .Z(n10080) );
  XOR U13677 ( .A(DB[581]), .B(DB[566]), .Z(n10082) );
  AND U13678 ( .A(n874), .B(n10083), .Z(n10081) );
  XOR U13679 ( .A(n10084), .B(n10085), .Z(n10083) );
  XOR U13680 ( .A(DB[566]), .B(DB[551]), .Z(n10085) );
  AND U13681 ( .A(n878), .B(n10086), .Z(n10084) );
  XOR U13682 ( .A(n10087), .B(n10088), .Z(n10086) );
  XOR U13683 ( .A(DB[551]), .B(DB[536]), .Z(n10088) );
  AND U13684 ( .A(n882), .B(n10089), .Z(n10087) );
  XOR U13685 ( .A(n10090), .B(n10091), .Z(n10089) );
  XOR U13686 ( .A(DB[536]), .B(DB[521]), .Z(n10091) );
  AND U13687 ( .A(n886), .B(n10092), .Z(n10090) );
  XOR U13688 ( .A(n10093), .B(n10094), .Z(n10092) );
  XOR U13689 ( .A(DB[521]), .B(DB[506]), .Z(n10094) );
  AND U13690 ( .A(n890), .B(n10095), .Z(n10093) );
  XOR U13691 ( .A(n10096), .B(n10097), .Z(n10095) );
  XOR U13692 ( .A(DB[506]), .B(DB[491]), .Z(n10097) );
  AND U13693 ( .A(n894), .B(n10098), .Z(n10096) );
  XOR U13694 ( .A(n10099), .B(n10100), .Z(n10098) );
  XOR U13695 ( .A(DB[491]), .B(DB[476]), .Z(n10100) );
  AND U13696 ( .A(n898), .B(n10101), .Z(n10099) );
  XOR U13697 ( .A(n10102), .B(n10103), .Z(n10101) );
  XOR U13698 ( .A(DB[476]), .B(DB[461]), .Z(n10103) );
  AND U13699 ( .A(n902), .B(n10104), .Z(n10102) );
  XOR U13700 ( .A(n10105), .B(n10106), .Z(n10104) );
  XOR U13701 ( .A(DB[461]), .B(DB[446]), .Z(n10106) );
  AND U13702 ( .A(n906), .B(n10107), .Z(n10105) );
  XOR U13703 ( .A(n10108), .B(n10109), .Z(n10107) );
  XOR U13704 ( .A(DB[446]), .B(DB[431]), .Z(n10109) );
  AND U13705 ( .A(n910), .B(n10110), .Z(n10108) );
  XOR U13706 ( .A(n10111), .B(n10112), .Z(n10110) );
  XOR U13707 ( .A(DB[431]), .B(DB[416]), .Z(n10112) );
  AND U13708 ( .A(n914), .B(n10113), .Z(n10111) );
  XOR U13709 ( .A(n10114), .B(n10115), .Z(n10113) );
  XOR U13710 ( .A(DB[416]), .B(DB[401]), .Z(n10115) );
  AND U13711 ( .A(n918), .B(n10116), .Z(n10114) );
  XOR U13712 ( .A(n10117), .B(n10118), .Z(n10116) );
  XOR U13713 ( .A(DB[401]), .B(DB[386]), .Z(n10118) );
  AND U13714 ( .A(n922), .B(n10119), .Z(n10117) );
  XOR U13715 ( .A(n10120), .B(n10121), .Z(n10119) );
  XOR U13716 ( .A(DB[386]), .B(DB[371]), .Z(n10121) );
  AND U13717 ( .A(n926), .B(n10122), .Z(n10120) );
  XOR U13718 ( .A(n10123), .B(n10124), .Z(n10122) );
  XOR U13719 ( .A(DB[371]), .B(DB[356]), .Z(n10124) );
  AND U13720 ( .A(n930), .B(n10125), .Z(n10123) );
  XOR U13721 ( .A(n10126), .B(n10127), .Z(n10125) );
  XOR U13722 ( .A(DB[356]), .B(DB[341]), .Z(n10127) );
  AND U13723 ( .A(n934), .B(n10128), .Z(n10126) );
  XOR U13724 ( .A(n10129), .B(n10130), .Z(n10128) );
  XOR U13725 ( .A(DB[341]), .B(DB[326]), .Z(n10130) );
  AND U13726 ( .A(n938), .B(n10131), .Z(n10129) );
  XOR U13727 ( .A(n10132), .B(n10133), .Z(n10131) );
  XOR U13728 ( .A(DB[326]), .B(DB[311]), .Z(n10133) );
  AND U13729 ( .A(n942), .B(n10134), .Z(n10132) );
  XOR U13730 ( .A(n10135), .B(n10136), .Z(n10134) );
  XOR U13731 ( .A(DB[311]), .B(DB[296]), .Z(n10136) );
  AND U13732 ( .A(n946), .B(n10137), .Z(n10135) );
  XOR U13733 ( .A(n10138), .B(n10139), .Z(n10137) );
  XOR U13734 ( .A(DB[296]), .B(DB[281]), .Z(n10139) );
  AND U13735 ( .A(n950), .B(n10140), .Z(n10138) );
  XOR U13736 ( .A(n10141), .B(n10142), .Z(n10140) );
  XOR U13737 ( .A(DB[281]), .B(DB[266]), .Z(n10142) );
  AND U13738 ( .A(n954), .B(n10143), .Z(n10141) );
  XOR U13739 ( .A(n10144), .B(n10145), .Z(n10143) );
  XOR U13740 ( .A(DB[266]), .B(DB[251]), .Z(n10145) );
  AND U13741 ( .A(n958), .B(n10146), .Z(n10144) );
  XOR U13742 ( .A(n10147), .B(n10148), .Z(n10146) );
  XOR U13743 ( .A(DB[251]), .B(DB[236]), .Z(n10148) );
  AND U13744 ( .A(n962), .B(n10149), .Z(n10147) );
  XOR U13745 ( .A(n10150), .B(n10151), .Z(n10149) );
  XOR U13746 ( .A(DB[236]), .B(DB[221]), .Z(n10151) );
  AND U13747 ( .A(n966), .B(n10152), .Z(n10150) );
  XOR U13748 ( .A(n10153), .B(n10154), .Z(n10152) );
  XOR U13749 ( .A(DB[221]), .B(DB[206]), .Z(n10154) );
  AND U13750 ( .A(n970), .B(n10155), .Z(n10153) );
  XOR U13751 ( .A(n10156), .B(n10157), .Z(n10155) );
  XOR U13752 ( .A(DB[206]), .B(DB[191]), .Z(n10157) );
  AND U13753 ( .A(n974), .B(n10158), .Z(n10156) );
  XOR U13754 ( .A(n10159), .B(n10160), .Z(n10158) );
  XOR U13755 ( .A(DB[191]), .B(DB[176]), .Z(n10160) );
  AND U13756 ( .A(n978), .B(n10161), .Z(n10159) );
  XOR U13757 ( .A(n10162), .B(n10163), .Z(n10161) );
  XOR U13758 ( .A(DB[176]), .B(DB[161]), .Z(n10163) );
  AND U13759 ( .A(n982), .B(n10164), .Z(n10162) );
  XOR U13760 ( .A(n10165), .B(n10166), .Z(n10164) );
  XOR U13761 ( .A(DB[161]), .B(DB[146]), .Z(n10166) );
  AND U13762 ( .A(n986), .B(n10167), .Z(n10165) );
  XOR U13763 ( .A(n10168), .B(n10169), .Z(n10167) );
  XOR U13764 ( .A(DB[146]), .B(DB[131]), .Z(n10169) );
  AND U13765 ( .A(n990), .B(n10170), .Z(n10168) );
  XOR U13766 ( .A(n10171), .B(n10172), .Z(n10170) );
  XOR U13767 ( .A(DB[131]), .B(DB[116]), .Z(n10172) );
  AND U13768 ( .A(n994), .B(n10173), .Z(n10171) );
  XOR U13769 ( .A(n10174), .B(n10175), .Z(n10173) );
  XOR U13770 ( .A(DB[116]), .B(DB[101]), .Z(n10175) );
  AND U13771 ( .A(n998), .B(n10176), .Z(n10174) );
  XOR U13772 ( .A(n10177), .B(n10178), .Z(n10176) );
  XOR U13773 ( .A(DB[86]), .B(DB[101]), .Z(n10178) );
  AND U13774 ( .A(n1002), .B(n10179), .Z(n10177) );
  XOR U13775 ( .A(n10180), .B(n10181), .Z(n10179) );
  XOR U13776 ( .A(DB[86]), .B(DB[71]), .Z(n10181) );
  AND U13777 ( .A(n1006), .B(n10182), .Z(n10180) );
  XOR U13778 ( .A(n10183), .B(n10184), .Z(n10182) );
  XOR U13779 ( .A(DB[71]), .B(DB[56]), .Z(n10184) );
  AND U13780 ( .A(n1010), .B(n10185), .Z(n10183) );
  XOR U13781 ( .A(n10186), .B(n10187), .Z(n10185) );
  XOR U13782 ( .A(DB[56]), .B(DB[41]), .Z(n10187) );
  AND U13783 ( .A(n1014), .B(n10188), .Z(n10186) );
  XOR U13784 ( .A(n10189), .B(n10190), .Z(n10188) );
  XOR U13785 ( .A(DB[41]), .B(DB[26]), .Z(n10190) );
  AND U13786 ( .A(n1018), .B(n10191), .Z(n10189) );
  XOR U13787 ( .A(DB[26]), .B(DB[11]), .Z(n10191) );
  XOR U13788 ( .A(DB[3835]), .B(n10192), .Z(min_val_out[10]) );
  AND U13789 ( .A(n2), .B(n10193), .Z(n10192) );
  XOR U13790 ( .A(n10194), .B(n10195), .Z(n10193) );
  XOR U13791 ( .A(DB[3835]), .B(DB[3820]), .Z(n10195) );
  AND U13792 ( .A(n6), .B(n10196), .Z(n10194) );
  XOR U13793 ( .A(n10197), .B(n10198), .Z(n10196) );
  XOR U13794 ( .A(DB[3820]), .B(DB[3805]), .Z(n10198) );
  AND U13795 ( .A(n10), .B(n10199), .Z(n10197) );
  XOR U13796 ( .A(n10200), .B(n10201), .Z(n10199) );
  XOR U13797 ( .A(DB[3805]), .B(DB[3790]), .Z(n10201) );
  AND U13798 ( .A(n14), .B(n10202), .Z(n10200) );
  XOR U13799 ( .A(n10203), .B(n10204), .Z(n10202) );
  XOR U13800 ( .A(DB[3790]), .B(DB[3775]), .Z(n10204) );
  AND U13801 ( .A(n18), .B(n10205), .Z(n10203) );
  XOR U13802 ( .A(n10206), .B(n10207), .Z(n10205) );
  XOR U13803 ( .A(DB[3775]), .B(DB[3760]), .Z(n10207) );
  AND U13804 ( .A(n22), .B(n10208), .Z(n10206) );
  XOR U13805 ( .A(n10209), .B(n10210), .Z(n10208) );
  XOR U13806 ( .A(DB[3760]), .B(DB[3745]), .Z(n10210) );
  AND U13807 ( .A(n26), .B(n10211), .Z(n10209) );
  XOR U13808 ( .A(n10212), .B(n10213), .Z(n10211) );
  XOR U13809 ( .A(DB[3745]), .B(DB[3730]), .Z(n10213) );
  AND U13810 ( .A(n30), .B(n10214), .Z(n10212) );
  XOR U13811 ( .A(n10215), .B(n10216), .Z(n10214) );
  XOR U13812 ( .A(DB[3730]), .B(DB[3715]), .Z(n10216) );
  AND U13813 ( .A(n34), .B(n10217), .Z(n10215) );
  XOR U13814 ( .A(n10218), .B(n10219), .Z(n10217) );
  XOR U13815 ( .A(DB[3715]), .B(DB[3700]), .Z(n10219) );
  AND U13816 ( .A(n38), .B(n10220), .Z(n10218) );
  XOR U13817 ( .A(n10221), .B(n10222), .Z(n10220) );
  XOR U13818 ( .A(DB[3700]), .B(DB[3685]), .Z(n10222) );
  AND U13819 ( .A(n42), .B(n10223), .Z(n10221) );
  XOR U13820 ( .A(n10224), .B(n10225), .Z(n10223) );
  XOR U13821 ( .A(DB[3685]), .B(DB[3670]), .Z(n10225) );
  AND U13822 ( .A(n46), .B(n10226), .Z(n10224) );
  XOR U13823 ( .A(n10227), .B(n10228), .Z(n10226) );
  XOR U13824 ( .A(DB[3670]), .B(DB[3655]), .Z(n10228) );
  AND U13825 ( .A(n50), .B(n10229), .Z(n10227) );
  XOR U13826 ( .A(n10230), .B(n10231), .Z(n10229) );
  XOR U13827 ( .A(DB[3655]), .B(DB[3640]), .Z(n10231) );
  AND U13828 ( .A(n54), .B(n10232), .Z(n10230) );
  XOR U13829 ( .A(n10233), .B(n10234), .Z(n10232) );
  XOR U13830 ( .A(DB[3640]), .B(DB[3625]), .Z(n10234) );
  AND U13831 ( .A(n58), .B(n10235), .Z(n10233) );
  XOR U13832 ( .A(n10236), .B(n10237), .Z(n10235) );
  XOR U13833 ( .A(DB[3625]), .B(DB[3610]), .Z(n10237) );
  AND U13834 ( .A(n62), .B(n10238), .Z(n10236) );
  XOR U13835 ( .A(n10239), .B(n10240), .Z(n10238) );
  XOR U13836 ( .A(DB[3610]), .B(DB[3595]), .Z(n10240) );
  AND U13837 ( .A(n66), .B(n10241), .Z(n10239) );
  XOR U13838 ( .A(n10242), .B(n10243), .Z(n10241) );
  XOR U13839 ( .A(DB[3595]), .B(DB[3580]), .Z(n10243) );
  AND U13840 ( .A(n70), .B(n10244), .Z(n10242) );
  XOR U13841 ( .A(n10245), .B(n10246), .Z(n10244) );
  XOR U13842 ( .A(DB[3580]), .B(DB[3565]), .Z(n10246) );
  AND U13843 ( .A(n74), .B(n10247), .Z(n10245) );
  XOR U13844 ( .A(n10248), .B(n10249), .Z(n10247) );
  XOR U13845 ( .A(DB[3565]), .B(DB[3550]), .Z(n10249) );
  AND U13846 ( .A(n78), .B(n10250), .Z(n10248) );
  XOR U13847 ( .A(n10251), .B(n10252), .Z(n10250) );
  XOR U13848 ( .A(DB[3550]), .B(DB[3535]), .Z(n10252) );
  AND U13849 ( .A(n82), .B(n10253), .Z(n10251) );
  XOR U13850 ( .A(n10254), .B(n10255), .Z(n10253) );
  XOR U13851 ( .A(DB[3535]), .B(DB[3520]), .Z(n10255) );
  AND U13852 ( .A(n86), .B(n10256), .Z(n10254) );
  XOR U13853 ( .A(n10257), .B(n10258), .Z(n10256) );
  XOR U13854 ( .A(DB[3520]), .B(DB[3505]), .Z(n10258) );
  AND U13855 ( .A(n90), .B(n10259), .Z(n10257) );
  XOR U13856 ( .A(n10260), .B(n10261), .Z(n10259) );
  XOR U13857 ( .A(DB[3505]), .B(DB[3490]), .Z(n10261) );
  AND U13858 ( .A(n94), .B(n10262), .Z(n10260) );
  XOR U13859 ( .A(n10263), .B(n10264), .Z(n10262) );
  XOR U13860 ( .A(DB[3490]), .B(DB[3475]), .Z(n10264) );
  AND U13861 ( .A(n98), .B(n10265), .Z(n10263) );
  XOR U13862 ( .A(n10266), .B(n10267), .Z(n10265) );
  XOR U13863 ( .A(DB[3475]), .B(DB[3460]), .Z(n10267) );
  AND U13864 ( .A(n102), .B(n10268), .Z(n10266) );
  XOR U13865 ( .A(n10269), .B(n10270), .Z(n10268) );
  XOR U13866 ( .A(DB[3460]), .B(DB[3445]), .Z(n10270) );
  AND U13867 ( .A(n106), .B(n10271), .Z(n10269) );
  XOR U13868 ( .A(n10272), .B(n10273), .Z(n10271) );
  XOR U13869 ( .A(DB[3445]), .B(DB[3430]), .Z(n10273) );
  AND U13870 ( .A(n110), .B(n10274), .Z(n10272) );
  XOR U13871 ( .A(n10275), .B(n10276), .Z(n10274) );
  XOR U13872 ( .A(DB[3430]), .B(DB[3415]), .Z(n10276) );
  AND U13873 ( .A(n114), .B(n10277), .Z(n10275) );
  XOR U13874 ( .A(n10278), .B(n10279), .Z(n10277) );
  XOR U13875 ( .A(DB[3415]), .B(DB[3400]), .Z(n10279) );
  AND U13876 ( .A(n118), .B(n10280), .Z(n10278) );
  XOR U13877 ( .A(n10281), .B(n10282), .Z(n10280) );
  XOR U13878 ( .A(DB[3400]), .B(DB[3385]), .Z(n10282) );
  AND U13879 ( .A(n122), .B(n10283), .Z(n10281) );
  XOR U13880 ( .A(n10284), .B(n10285), .Z(n10283) );
  XOR U13881 ( .A(DB[3385]), .B(DB[3370]), .Z(n10285) );
  AND U13882 ( .A(n126), .B(n10286), .Z(n10284) );
  XOR U13883 ( .A(n10287), .B(n10288), .Z(n10286) );
  XOR U13884 ( .A(DB[3370]), .B(DB[3355]), .Z(n10288) );
  AND U13885 ( .A(n130), .B(n10289), .Z(n10287) );
  XOR U13886 ( .A(n10290), .B(n10291), .Z(n10289) );
  XOR U13887 ( .A(DB[3355]), .B(DB[3340]), .Z(n10291) );
  AND U13888 ( .A(n134), .B(n10292), .Z(n10290) );
  XOR U13889 ( .A(n10293), .B(n10294), .Z(n10292) );
  XOR U13890 ( .A(DB[3340]), .B(DB[3325]), .Z(n10294) );
  AND U13891 ( .A(n138), .B(n10295), .Z(n10293) );
  XOR U13892 ( .A(n10296), .B(n10297), .Z(n10295) );
  XOR U13893 ( .A(DB[3325]), .B(DB[3310]), .Z(n10297) );
  AND U13894 ( .A(n142), .B(n10298), .Z(n10296) );
  XOR U13895 ( .A(n10299), .B(n10300), .Z(n10298) );
  XOR U13896 ( .A(DB[3310]), .B(DB[3295]), .Z(n10300) );
  AND U13897 ( .A(n146), .B(n10301), .Z(n10299) );
  XOR U13898 ( .A(n10302), .B(n10303), .Z(n10301) );
  XOR U13899 ( .A(DB[3295]), .B(DB[3280]), .Z(n10303) );
  AND U13900 ( .A(n150), .B(n10304), .Z(n10302) );
  XOR U13901 ( .A(n10305), .B(n10306), .Z(n10304) );
  XOR U13902 ( .A(DB[3280]), .B(DB[3265]), .Z(n10306) );
  AND U13903 ( .A(n154), .B(n10307), .Z(n10305) );
  XOR U13904 ( .A(n10308), .B(n10309), .Z(n10307) );
  XOR U13905 ( .A(DB[3265]), .B(DB[3250]), .Z(n10309) );
  AND U13906 ( .A(n158), .B(n10310), .Z(n10308) );
  XOR U13907 ( .A(n10311), .B(n10312), .Z(n10310) );
  XOR U13908 ( .A(DB[3250]), .B(DB[3235]), .Z(n10312) );
  AND U13909 ( .A(n162), .B(n10313), .Z(n10311) );
  XOR U13910 ( .A(n10314), .B(n10315), .Z(n10313) );
  XOR U13911 ( .A(DB[3235]), .B(DB[3220]), .Z(n10315) );
  AND U13912 ( .A(n166), .B(n10316), .Z(n10314) );
  XOR U13913 ( .A(n10317), .B(n10318), .Z(n10316) );
  XOR U13914 ( .A(DB[3220]), .B(DB[3205]), .Z(n10318) );
  AND U13915 ( .A(n170), .B(n10319), .Z(n10317) );
  XOR U13916 ( .A(n10320), .B(n10321), .Z(n10319) );
  XOR U13917 ( .A(DB[3205]), .B(DB[3190]), .Z(n10321) );
  AND U13918 ( .A(n174), .B(n10322), .Z(n10320) );
  XOR U13919 ( .A(n10323), .B(n10324), .Z(n10322) );
  XOR U13920 ( .A(DB[3190]), .B(DB[3175]), .Z(n10324) );
  AND U13921 ( .A(n178), .B(n10325), .Z(n10323) );
  XOR U13922 ( .A(n10326), .B(n10327), .Z(n10325) );
  XOR U13923 ( .A(DB[3175]), .B(DB[3160]), .Z(n10327) );
  AND U13924 ( .A(n182), .B(n10328), .Z(n10326) );
  XOR U13925 ( .A(n10329), .B(n10330), .Z(n10328) );
  XOR U13926 ( .A(DB[3160]), .B(DB[3145]), .Z(n10330) );
  AND U13927 ( .A(n186), .B(n10331), .Z(n10329) );
  XOR U13928 ( .A(n10332), .B(n10333), .Z(n10331) );
  XOR U13929 ( .A(DB[3145]), .B(DB[3130]), .Z(n10333) );
  AND U13930 ( .A(n190), .B(n10334), .Z(n10332) );
  XOR U13931 ( .A(n10335), .B(n10336), .Z(n10334) );
  XOR U13932 ( .A(DB[3130]), .B(DB[3115]), .Z(n10336) );
  AND U13933 ( .A(n194), .B(n10337), .Z(n10335) );
  XOR U13934 ( .A(n10338), .B(n10339), .Z(n10337) );
  XOR U13935 ( .A(DB[3115]), .B(DB[3100]), .Z(n10339) );
  AND U13936 ( .A(n198), .B(n10340), .Z(n10338) );
  XOR U13937 ( .A(n10341), .B(n10342), .Z(n10340) );
  XOR U13938 ( .A(DB[3100]), .B(DB[3085]), .Z(n10342) );
  AND U13939 ( .A(n202), .B(n10343), .Z(n10341) );
  XOR U13940 ( .A(n10344), .B(n10345), .Z(n10343) );
  XOR U13941 ( .A(DB[3085]), .B(DB[3070]), .Z(n10345) );
  AND U13942 ( .A(n206), .B(n10346), .Z(n10344) );
  XOR U13943 ( .A(n10347), .B(n10348), .Z(n10346) );
  XOR U13944 ( .A(DB[3070]), .B(DB[3055]), .Z(n10348) );
  AND U13945 ( .A(n210), .B(n10349), .Z(n10347) );
  XOR U13946 ( .A(n10350), .B(n10351), .Z(n10349) );
  XOR U13947 ( .A(DB[3055]), .B(DB[3040]), .Z(n10351) );
  AND U13948 ( .A(n214), .B(n10352), .Z(n10350) );
  XOR U13949 ( .A(n10353), .B(n10354), .Z(n10352) );
  XOR U13950 ( .A(DB[3040]), .B(DB[3025]), .Z(n10354) );
  AND U13951 ( .A(n218), .B(n10355), .Z(n10353) );
  XOR U13952 ( .A(n10356), .B(n10357), .Z(n10355) );
  XOR U13953 ( .A(DB[3025]), .B(DB[3010]), .Z(n10357) );
  AND U13954 ( .A(n222), .B(n10358), .Z(n10356) );
  XOR U13955 ( .A(n10359), .B(n10360), .Z(n10358) );
  XOR U13956 ( .A(DB[3010]), .B(DB[2995]), .Z(n10360) );
  AND U13957 ( .A(n226), .B(n10361), .Z(n10359) );
  XOR U13958 ( .A(n10362), .B(n10363), .Z(n10361) );
  XOR U13959 ( .A(DB[2995]), .B(DB[2980]), .Z(n10363) );
  AND U13960 ( .A(n230), .B(n10364), .Z(n10362) );
  XOR U13961 ( .A(n10365), .B(n10366), .Z(n10364) );
  XOR U13962 ( .A(DB[2980]), .B(DB[2965]), .Z(n10366) );
  AND U13963 ( .A(n234), .B(n10367), .Z(n10365) );
  XOR U13964 ( .A(n10368), .B(n10369), .Z(n10367) );
  XOR U13965 ( .A(DB[2965]), .B(DB[2950]), .Z(n10369) );
  AND U13966 ( .A(n238), .B(n10370), .Z(n10368) );
  XOR U13967 ( .A(n10371), .B(n10372), .Z(n10370) );
  XOR U13968 ( .A(DB[2950]), .B(DB[2935]), .Z(n10372) );
  AND U13969 ( .A(n242), .B(n10373), .Z(n10371) );
  XOR U13970 ( .A(n10374), .B(n10375), .Z(n10373) );
  XOR U13971 ( .A(DB[2935]), .B(DB[2920]), .Z(n10375) );
  AND U13972 ( .A(n246), .B(n10376), .Z(n10374) );
  XOR U13973 ( .A(n10377), .B(n10378), .Z(n10376) );
  XOR U13974 ( .A(DB[2920]), .B(DB[2905]), .Z(n10378) );
  AND U13975 ( .A(n250), .B(n10379), .Z(n10377) );
  XOR U13976 ( .A(n10380), .B(n10381), .Z(n10379) );
  XOR U13977 ( .A(DB[2905]), .B(DB[2890]), .Z(n10381) );
  AND U13978 ( .A(n254), .B(n10382), .Z(n10380) );
  XOR U13979 ( .A(n10383), .B(n10384), .Z(n10382) );
  XOR U13980 ( .A(DB[2890]), .B(DB[2875]), .Z(n10384) );
  AND U13981 ( .A(n258), .B(n10385), .Z(n10383) );
  XOR U13982 ( .A(n10386), .B(n10387), .Z(n10385) );
  XOR U13983 ( .A(DB[2875]), .B(DB[2860]), .Z(n10387) );
  AND U13984 ( .A(n262), .B(n10388), .Z(n10386) );
  XOR U13985 ( .A(n10389), .B(n10390), .Z(n10388) );
  XOR U13986 ( .A(DB[2860]), .B(DB[2845]), .Z(n10390) );
  AND U13987 ( .A(n266), .B(n10391), .Z(n10389) );
  XOR U13988 ( .A(n10392), .B(n10393), .Z(n10391) );
  XOR U13989 ( .A(DB[2845]), .B(DB[2830]), .Z(n10393) );
  AND U13990 ( .A(n270), .B(n10394), .Z(n10392) );
  XOR U13991 ( .A(n10395), .B(n10396), .Z(n10394) );
  XOR U13992 ( .A(DB[2830]), .B(DB[2815]), .Z(n10396) );
  AND U13993 ( .A(n274), .B(n10397), .Z(n10395) );
  XOR U13994 ( .A(n10398), .B(n10399), .Z(n10397) );
  XOR U13995 ( .A(DB[2815]), .B(DB[2800]), .Z(n10399) );
  AND U13996 ( .A(n278), .B(n10400), .Z(n10398) );
  XOR U13997 ( .A(n10401), .B(n10402), .Z(n10400) );
  XOR U13998 ( .A(DB[2800]), .B(DB[2785]), .Z(n10402) );
  AND U13999 ( .A(n282), .B(n10403), .Z(n10401) );
  XOR U14000 ( .A(n10404), .B(n10405), .Z(n10403) );
  XOR U14001 ( .A(DB[2785]), .B(DB[2770]), .Z(n10405) );
  AND U14002 ( .A(n286), .B(n10406), .Z(n10404) );
  XOR U14003 ( .A(n10407), .B(n10408), .Z(n10406) );
  XOR U14004 ( .A(DB[2770]), .B(DB[2755]), .Z(n10408) );
  AND U14005 ( .A(n290), .B(n10409), .Z(n10407) );
  XOR U14006 ( .A(n10410), .B(n10411), .Z(n10409) );
  XOR U14007 ( .A(DB[2755]), .B(DB[2740]), .Z(n10411) );
  AND U14008 ( .A(n294), .B(n10412), .Z(n10410) );
  XOR U14009 ( .A(n10413), .B(n10414), .Z(n10412) );
  XOR U14010 ( .A(DB[2740]), .B(DB[2725]), .Z(n10414) );
  AND U14011 ( .A(n298), .B(n10415), .Z(n10413) );
  XOR U14012 ( .A(n10416), .B(n10417), .Z(n10415) );
  XOR U14013 ( .A(DB[2725]), .B(DB[2710]), .Z(n10417) );
  AND U14014 ( .A(n302), .B(n10418), .Z(n10416) );
  XOR U14015 ( .A(n10419), .B(n10420), .Z(n10418) );
  XOR U14016 ( .A(DB[2710]), .B(DB[2695]), .Z(n10420) );
  AND U14017 ( .A(n306), .B(n10421), .Z(n10419) );
  XOR U14018 ( .A(n10422), .B(n10423), .Z(n10421) );
  XOR U14019 ( .A(DB[2695]), .B(DB[2680]), .Z(n10423) );
  AND U14020 ( .A(n310), .B(n10424), .Z(n10422) );
  XOR U14021 ( .A(n10425), .B(n10426), .Z(n10424) );
  XOR U14022 ( .A(DB[2680]), .B(DB[2665]), .Z(n10426) );
  AND U14023 ( .A(n314), .B(n10427), .Z(n10425) );
  XOR U14024 ( .A(n10428), .B(n10429), .Z(n10427) );
  XOR U14025 ( .A(DB[2665]), .B(DB[2650]), .Z(n10429) );
  AND U14026 ( .A(n318), .B(n10430), .Z(n10428) );
  XOR U14027 ( .A(n10431), .B(n10432), .Z(n10430) );
  XOR U14028 ( .A(DB[2650]), .B(DB[2635]), .Z(n10432) );
  AND U14029 ( .A(n322), .B(n10433), .Z(n10431) );
  XOR U14030 ( .A(n10434), .B(n10435), .Z(n10433) );
  XOR U14031 ( .A(DB[2635]), .B(DB[2620]), .Z(n10435) );
  AND U14032 ( .A(n326), .B(n10436), .Z(n10434) );
  XOR U14033 ( .A(n10437), .B(n10438), .Z(n10436) );
  XOR U14034 ( .A(DB[2620]), .B(DB[2605]), .Z(n10438) );
  AND U14035 ( .A(n330), .B(n10439), .Z(n10437) );
  XOR U14036 ( .A(n10440), .B(n10441), .Z(n10439) );
  XOR U14037 ( .A(DB[2605]), .B(DB[2590]), .Z(n10441) );
  AND U14038 ( .A(n334), .B(n10442), .Z(n10440) );
  XOR U14039 ( .A(n10443), .B(n10444), .Z(n10442) );
  XOR U14040 ( .A(DB[2590]), .B(DB[2575]), .Z(n10444) );
  AND U14041 ( .A(n338), .B(n10445), .Z(n10443) );
  XOR U14042 ( .A(n10446), .B(n10447), .Z(n10445) );
  XOR U14043 ( .A(DB[2575]), .B(DB[2560]), .Z(n10447) );
  AND U14044 ( .A(n342), .B(n10448), .Z(n10446) );
  XOR U14045 ( .A(n10449), .B(n10450), .Z(n10448) );
  XOR U14046 ( .A(DB[2560]), .B(DB[2545]), .Z(n10450) );
  AND U14047 ( .A(n346), .B(n10451), .Z(n10449) );
  XOR U14048 ( .A(n10452), .B(n10453), .Z(n10451) );
  XOR U14049 ( .A(DB[2545]), .B(DB[2530]), .Z(n10453) );
  AND U14050 ( .A(n350), .B(n10454), .Z(n10452) );
  XOR U14051 ( .A(n10455), .B(n10456), .Z(n10454) );
  XOR U14052 ( .A(DB[2530]), .B(DB[2515]), .Z(n10456) );
  AND U14053 ( .A(n354), .B(n10457), .Z(n10455) );
  XOR U14054 ( .A(n10458), .B(n10459), .Z(n10457) );
  XOR U14055 ( .A(DB[2515]), .B(DB[2500]), .Z(n10459) );
  AND U14056 ( .A(n358), .B(n10460), .Z(n10458) );
  XOR U14057 ( .A(n10461), .B(n10462), .Z(n10460) );
  XOR U14058 ( .A(DB[2500]), .B(DB[2485]), .Z(n10462) );
  AND U14059 ( .A(n362), .B(n10463), .Z(n10461) );
  XOR U14060 ( .A(n10464), .B(n10465), .Z(n10463) );
  XOR U14061 ( .A(DB[2485]), .B(DB[2470]), .Z(n10465) );
  AND U14062 ( .A(n366), .B(n10466), .Z(n10464) );
  XOR U14063 ( .A(n10467), .B(n10468), .Z(n10466) );
  XOR U14064 ( .A(DB[2470]), .B(DB[2455]), .Z(n10468) );
  AND U14065 ( .A(n370), .B(n10469), .Z(n10467) );
  XOR U14066 ( .A(n10470), .B(n10471), .Z(n10469) );
  XOR U14067 ( .A(DB[2455]), .B(DB[2440]), .Z(n10471) );
  AND U14068 ( .A(n374), .B(n10472), .Z(n10470) );
  XOR U14069 ( .A(n10473), .B(n10474), .Z(n10472) );
  XOR U14070 ( .A(DB[2440]), .B(DB[2425]), .Z(n10474) );
  AND U14071 ( .A(n378), .B(n10475), .Z(n10473) );
  XOR U14072 ( .A(n10476), .B(n10477), .Z(n10475) );
  XOR U14073 ( .A(DB[2425]), .B(DB[2410]), .Z(n10477) );
  AND U14074 ( .A(n382), .B(n10478), .Z(n10476) );
  XOR U14075 ( .A(n10479), .B(n10480), .Z(n10478) );
  XOR U14076 ( .A(DB[2410]), .B(DB[2395]), .Z(n10480) );
  AND U14077 ( .A(n386), .B(n10481), .Z(n10479) );
  XOR U14078 ( .A(n10482), .B(n10483), .Z(n10481) );
  XOR U14079 ( .A(DB[2395]), .B(DB[2380]), .Z(n10483) );
  AND U14080 ( .A(n390), .B(n10484), .Z(n10482) );
  XOR U14081 ( .A(n10485), .B(n10486), .Z(n10484) );
  XOR U14082 ( .A(DB[2380]), .B(DB[2365]), .Z(n10486) );
  AND U14083 ( .A(n394), .B(n10487), .Z(n10485) );
  XOR U14084 ( .A(n10488), .B(n10489), .Z(n10487) );
  XOR U14085 ( .A(DB[2365]), .B(DB[2350]), .Z(n10489) );
  AND U14086 ( .A(n398), .B(n10490), .Z(n10488) );
  XOR U14087 ( .A(n10491), .B(n10492), .Z(n10490) );
  XOR U14088 ( .A(DB[2350]), .B(DB[2335]), .Z(n10492) );
  AND U14089 ( .A(n402), .B(n10493), .Z(n10491) );
  XOR U14090 ( .A(n10494), .B(n10495), .Z(n10493) );
  XOR U14091 ( .A(DB[2335]), .B(DB[2320]), .Z(n10495) );
  AND U14092 ( .A(n406), .B(n10496), .Z(n10494) );
  XOR U14093 ( .A(n10497), .B(n10498), .Z(n10496) );
  XOR U14094 ( .A(DB[2320]), .B(DB[2305]), .Z(n10498) );
  AND U14095 ( .A(n410), .B(n10499), .Z(n10497) );
  XOR U14096 ( .A(n10500), .B(n10501), .Z(n10499) );
  XOR U14097 ( .A(DB[2305]), .B(DB[2290]), .Z(n10501) );
  AND U14098 ( .A(n414), .B(n10502), .Z(n10500) );
  XOR U14099 ( .A(n10503), .B(n10504), .Z(n10502) );
  XOR U14100 ( .A(DB[2290]), .B(DB[2275]), .Z(n10504) );
  AND U14101 ( .A(n418), .B(n10505), .Z(n10503) );
  XOR U14102 ( .A(n10506), .B(n10507), .Z(n10505) );
  XOR U14103 ( .A(DB[2275]), .B(DB[2260]), .Z(n10507) );
  AND U14104 ( .A(n422), .B(n10508), .Z(n10506) );
  XOR U14105 ( .A(n10509), .B(n10510), .Z(n10508) );
  XOR U14106 ( .A(DB[2260]), .B(DB[2245]), .Z(n10510) );
  AND U14107 ( .A(n426), .B(n10511), .Z(n10509) );
  XOR U14108 ( .A(n10512), .B(n10513), .Z(n10511) );
  XOR U14109 ( .A(DB[2245]), .B(DB[2230]), .Z(n10513) );
  AND U14110 ( .A(n430), .B(n10514), .Z(n10512) );
  XOR U14111 ( .A(n10515), .B(n10516), .Z(n10514) );
  XOR U14112 ( .A(DB[2230]), .B(DB[2215]), .Z(n10516) );
  AND U14113 ( .A(n434), .B(n10517), .Z(n10515) );
  XOR U14114 ( .A(n10518), .B(n10519), .Z(n10517) );
  XOR U14115 ( .A(DB[2215]), .B(DB[2200]), .Z(n10519) );
  AND U14116 ( .A(n438), .B(n10520), .Z(n10518) );
  XOR U14117 ( .A(n10521), .B(n10522), .Z(n10520) );
  XOR U14118 ( .A(DB[2200]), .B(DB[2185]), .Z(n10522) );
  AND U14119 ( .A(n442), .B(n10523), .Z(n10521) );
  XOR U14120 ( .A(n10524), .B(n10525), .Z(n10523) );
  XOR U14121 ( .A(DB[2185]), .B(DB[2170]), .Z(n10525) );
  AND U14122 ( .A(n446), .B(n10526), .Z(n10524) );
  XOR U14123 ( .A(n10527), .B(n10528), .Z(n10526) );
  XOR U14124 ( .A(DB[2170]), .B(DB[2155]), .Z(n10528) );
  AND U14125 ( .A(n450), .B(n10529), .Z(n10527) );
  XOR U14126 ( .A(n10530), .B(n10531), .Z(n10529) );
  XOR U14127 ( .A(DB[2155]), .B(DB[2140]), .Z(n10531) );
  AND U14128 ( .A(n454), .B(n10532), .Z(n10530) );
  XOR U14129 ( .A(n10533), .B(n10534), .Z(n10532) );
  XOR U14130 ( .A(DB[2140]), .B(DB[2125]), .Z(n10534) );
  AND U14131 ( .A(n458), .B(n10535), .Z(n10533) );
  XOR U14132 ( .A(n10536), .B(n10537), .Z(n10535) );
  XOR U14133 ( .A(DB[2125]), .B(DB[2110]), .Z(n10537) );
  AND U14134 ( .A(n462), .B(n10538), .Z(n10536) );
  XOR U14135 ( .A(n10539), .B(n10540), .Z(n10538) );
  XOR U14136 ( .A(DB[2110]), .B(DB[2095]), .Z(n10540) );
  AND U14137 ( .A(n466), .B(n10541), .Z(n10539) );
  XOR U14138 ( .A(n10542), .B(n10543), .Z(n10541) );
  XOR U14139 ( .A(DB[2095]), .B(DB[2080]), .Z(n10543) );
  AND U14140 ( .A(n470), .B(n10544), .Z(n10542) );
  XOR U14141 ( .A(n10545), .B(n10546), .Z(n10544) );
  XOR U14142 ( .A(DB[2080]), .B(DB[2065]), .Z(n10546) );
  AND U14143 ( .A(n474), .B(n10547), .Z(n10545) );
  XOR U14144 ( .A(n10548), .B(n10549), .Z(n10547) );
  XOR U14145 ( .A(DB[2065]), .B(DB[2050]), .Z(n10549) );
  AND U14146 ( .A(n478), .B(n10550), .Z(n10548) );
  XOR U14147 ( .A(n10551), .B(n10552), .Z(n10550) );
  XOR U14148 ( .A(DB[2050]), .B(DB[2035]), .Z(n10552) );
  AND U14149 ( .A(n482), .B(n10553), .Z(n10551) );
  XOR U14150 ( .A(n10554), .B(n10555), .Z(n10553) );
  XOR U14151 ( .A(DB[2035]), .B(DB[2020]), .Z(n10555) );
  AND U14152 ( .A(n486), .B(n10556), .Z(n10554) );
  XOR U14153 ( .A(n10557), .B(n10558), .Z(n10556) );
  XOR U14154 ( .A(DB[2020]), .B(DB[2005]), .Z(n10558) );
  AND U14155 ( .A(n490), .B(n10559), .Z(n10557) );
  XOR U14156 ( .A(n10560), .B(n10561), .Z(n10559) );
  XOR U14157 ( .A(DB[2005]), .B(DB[1990]), .Z(n10561) );
  AND U14158 ( .A(n494), .B(n10562), .Z(n10560) );
  XOR U14159 ( .A(n10563), .B(n10564), .Z(n10562) );
  XOR U14160 ( .A(DB[1990]), .B(DB[1975]), .Z(n10564) );
  AND U14161 ( .A(n498), .B(n10565), .Z(n10563) );
  XOR U14162 ( .A(n10566), .B(n10567), .Z(n10565) );
  XOR U14163 ( .A(DB[1975]), .B(DB[1960]), .Z(n10567) );
  AND U14164 ( .A(n502), .B(n10568), .Z(n10566) );
  XOR U14165 ( .A(n10569), .B(n10570), .Z(n10568) );
  XOR U14166 ( .A(DB[1960]), .B(DB[1945]), .Z(n10570) );
  AND U14167 ( .A(n506), .B(n10571), .Z(n10569) );
  XOR U14168 ( .A(n10572), .B(n10573), .Z(n10571) );
  XOR U14169 ( .A(DB[1945]), .B(DB[1930]), .Z(n10573) );
  AND U14170 ( .A(n510), .B(n10574), .Z(n10572) );
  XOR U14171 ( .A(n10575), .B(n10576), .Z(n10574) );
  XOR U14172 ( .A(DB[1930]), .B(DB[1915]), .Z(n10576) );
  AND U14173 ( .A(n514), .B(n10577), .Z(n10575) );
  XOR U14174 ( .A(n10578), .B(n10579), .Z(n10577) );
  XOR U14175 ( .A(DB[1915]), .B(DB[1900]), .Z(n10579) );
  AND U14176 ( .A(n518), .B(n10580), .Z(n10578) );
  XOR U14177 ( .A(n10581), .B(n10582), .Z(n10580) );
  XOR U14178 ( .A(DB[1900]), .B(DB[1885]), .Z(n10582) );
  AND U14179 ( .A(n522), .B(n10583), .Z(n10581) );
  XOR U14180 ( .A(n10584), .B(n10585), .Z(n10583) );
  XOR U14181 ( .A(DB[1885]), .B(DB[1870]), .Z(n10585) );
  AND U14182 ( .A(n526), .B(n10586), .Z(n10584) );
  XOR U14183 ( .A(n10587), .B(n10588), .Z(n10586) );
  XOR U14184 ( .A(DB[1870]), .B(DB[1855]), .Z(n10588) );
  AND U14185 ( .A(n530), .B(n10589), .Z(n10587) );
  XOR U14186 ( .A(n10590), .B(n10591), .Z(n10589) );
  XOR U14187 ( .A(DB[1855]), .B(DB[1840]), .Z(n10591) );
  AND U14188 ( .A(n534), .B(n10592), .Z(n10590) );
  XOR U14189 ( .A(n10593), .B(n10594), .Z(n10592) );
  XOR U14190 ( .A(DB[1840]), .B(DB[1825]), .Z(n10594) );
  AND U14191 ( .A(n538), .B(n10595), .Z(n10593) );
  XOR U14192 ( .A(n10596), .B(n10597), .Z(n10595) );
  XOR U14193 ( .A(DB[1825]), .B(DB[1810]), .Z(n10597) );
  AND U14194 ( .A(n542), .B(n10598), .Z(n10596) );
  XOR U14195 ( .A(n10599), .B(n10600), .Z(n10598) );
  XOR U14196 ( .A(DB[1810]), .B(DB[1795]), .Z(n10600) );
  AND U14197 ( .A(n546), .B(n10601), .Z(n10599) );
  XOR U14198 ( .A(n10602), .B(n10603), .Z(n10601) );
  XOR U14199 ( .A(DB[1795]), .B(DB[1780]), .Z(n10603) );
  AND U14200 ( .A(n550), .B(n10604), .Z(n10602) );
  XOR U14201 ( .A(n10605), .B(n10606), .Z(n10604) );
  XOR U14202 ( .A(DB[1780]), .B(DB[1765]), .Z(n10606) );
  AND U14203 ( .A(n554), .B(n10607), .Z(n10605) );
  XOR U14204 ( .A(n10608), .B(n10609), .Z(n10607) );
  XOR U14205 ( .A(DB[1765]), .B(DB[1750]), .Z(n10609) );
  AND U14206 ( .A(n558), .B(n10610), .Z(n10608) );
  XOR U14207 ( .A(n10611), .B(n10612), .Z(n10610) );
  XOR U14208 ( .A(DB[1750]), .B(DB[1735]), .Z(n10612) );
  AND U14209 ( .A(n562), .B(n10613), .Z(n10611) );
  XOR U14210 ( .A(n10614), .B(n10615), .Z(n10613) );
  XOR U14211 ( .A(DB[1735]), .B(DB[1720]), .Z(n10615) );
  AND U14212 ( .A(n566), .B(n10616), .Z(n10614) );
  XOR U14213 ( .A(n10617), .B(n10618), .Z(n10616) );
  XOR U14214 ( .A(DB[1720]), .B(DB[1705]), .Z(n10618) );
  AND U14215 ( .A(n570), .B(n10619), .Z(n10617) );
  XOR U14216 ( .A(n10620), .B(n10621), .Z(n10619) );
  XOR U14217 ( .A(DB[1705]), .B(DB[1690]), .Z(n10621) );
  AND U14218 ( .A(n574), .B(n10622), .Z(n10620) );
  XOR U14219 ( .A(n10623), .B(n10624), .Z(n10622) );
  XOR U14220 ( .A(DB[1690]), .B(DB[1675]), .Z(n10624) );
  AND U14221 ( .A(n578), .B(n10625), .Z(n10623) );
  XOR U14222 ( .A(n10626), .B(n10627), .Z(n10625) );
  XOR U14223 ( .A(DB[1675]), .B(DB[1660]), .Z(n10627) );
  AND U14224 ( .A(n582), .B(n10628), .Z(n10626) );
  XOR U14225 ( .A(n10629), .B(n10630), .Z(n10628) );
  XOR U14226 ( .A(DB[1660]), .B(DB[1645]), .Z(n10630) );
  AND U14227 ( .A(n586), .B(n10631), .Z(n10629) );
  XOR U14228 ( .A(n10632), .B(n10633), .Z(n10631) );
  XOR U14229 ( .A(DB[1645]), .B(DB[1630]), .Z(n10633) );
  AND U14230 ( .A(n590), .B(n10634), .Z(n10632) );
  XOR U14231 ( .A(n10635), .B(n10636), .Z(n10634) );
  XOR U14232 ( .A(DB[1630]), .B(DB[1615]), .Z(n10636) );
  AND U14233 ( .A(n594), .B(n10637), .Z(n10635) );
  XOR U14234 ( .A(n10638), .B(n10639), .Z(n10637) );
  XOR U14235 ( .A(DB[1615]), .B(DB[1600]), .Z(n10639) );
  AND U14236 ( .A(n598), .B(n10640), .Z(n10638) );
  XOR U14237 ( .A(n10641), .B(n10642), .Z(n10640) );
  XOR U14238 ( .A(DB[1600]), .B(DB[1585]), .Z(n10642) );
  AND U14239 ( .A(n602), .B(n10643), .Z(n10641) );
  XOR U14240 ( .A(n10644), .B(n10645), .Z(n10643) );
  XOR U14241 ( .A(DB[1585]), .B(DB[1570]), .Z(n10645) );
  AND U14242 ( .A(n606), .B(n10646), .Z(n10644) );
  XOR U14243 ( .A(n10647), .B(n10648), .Z(n10646) );
  XOR U14244 ( .A(DB[1570]), .B(DB[1555]), .Z(n10648) );
  AND U14245 ( .A(n610), .B(n10649), .Z(n10647) );
  XOR U14246 ( .A(n10650), .B(n10651), .Z(n10649) );
  XOR U14247 ( .A(DB[1555]), .B(DB[1540]), .Z(n10651) );
  AND U14248 ( .A(n614), .B(n10652), .Z(n10650) );
  XOR U14249 ( .A(n10653), .B(n10654), .Z(n10652) );
  XOR U14250 ( .A(DB[1540]), .B(DB[1525]), .Z(n10654) );
  AND U14251 ( .A(n618), .B(n10655), .Z(n10653) );
  XOR U14252 ( .A(n10656), .B(n10657), .Z(n10655) );
  XOR U14253 ( .A(DB[1525]), .B(DB[1510]), .Z(n10657) );
  AND U14254 ( .A(n622), .B(n10658), .Z(n10656) );
  XOR U14255 ( .A(n10659), .B(n10660), .Z(n10658) );
  XOR U14256 ( .A(DB[1510]), .B(DB[1495]), .Z(n10660) );
  AND U14257 ( .A(n626), .B(n10661), .Z(n10659) );
  XOR U14258 ( .A(n10662), .B(n10663), .Z(n10661) );
  XOR U14259 ( .A(DB[1495]), .B(DB[1480]), .Z(n10663) );
  AND U14260 ( .A(n630), .B(n10664), .Z(n10662) );
  XOR U14261 ( .A(n10665), .B(n10666), .Z(n10664) );
  XOR U14262 ( .A(DB[1480]), .B(DB[1465]), .Z(n10666) );
  AND U14263 ( .A(n634), .B(n10667), .Z(n10665) );
  XOR U14264 ( .A(n10668), .B(n10669), .Z(n10667) );
  XOR U14265 ( .A(DB[1465]), .B(DB[1450]), .Z(n10669) );
  AND U14266 ( .A(n638), .B(n10670), .Z(n10668) );
  XOR U14267 ( .A(n10671), .B(n10672), .Z(n10670) );
  XOR U14268 ( .A(DB[1450]), .B(DB[1435]), .Z(n10672) );
  AND U14269 ( .A(n642), .B(n10673), .Z(n10671) );
  XOR U14270 ( .A(n10674), .B(n10675), .Z(n10673) );
  XOR U14271 ( .A(DB[1435]), .B(DB[1420]), .Z(n10675) );
  AND U14272 ( .A(n646), .B(n10676), .Z(n10674) );
  XOR U14273 ( .A(n10677), .B(n10678), .Z(n10676) );
  XOR U14274 ( .A(DB[1420]), .B(DB[1405]), .Z(n10678) );
  AND U14275 ( .A(n650), .B(n10679), .Z(n10677) );
  XOR U14276 ( .A(n10680), .B(n10681), .Z(n10679) );
  XOR U14277 ( .A(DB[1405]), .B(DB[1390]), .Z(n10681) );
  AND U14278 ( .A(n654), .B(n10682), .Z(n10680) );
  XOR U14279 ( .A(n10683), .B(n10684), .Z(n10682) );
  XOR U14280 ( .A(DB[1390]), .B(DB[1375]), .Z(n10684) );
  AND U14281 ( .A(n658), .B(n10685), .Z(n10683) );
  XOR U14282 ( .A(n10686), .B(n10687), .Z(n10685) );
  XOR U14283 ( .A(DB[1375]), .B(DB[1360]), .Z(n10687) );
  AND U14284 ( .A(n662), .B(n10688), .Z(n10686) );
  XOR U14285 ( .A(n10689), .B(n10690), .Z(n10688) );
  XOR U14286 ( .A(DB[1360]), .B(DB[1345]), .Z(n10690) );
  AND U14287 ( .A(n666), .B(n10691), .Z(n10689) );
  XOR U14288 ( .A(n10692), .B(n10693), .Z(n10691) );
  XOR U14289 ( .A(DB[1345]), .B(DB[1330]), .Z(n10693) );
  AND U14290 ( .A(n670), .B(n10694), .Z(n10692) );
  XOR U14291 ( .A(n10695), .B(n10696), .Z(n10694) );
  XOR U14292 ( .A(DB[1330]), .B(DB[1315]), .Z(n10696) );
  AND U14293 ( .A(n674), .B(n10697), .Z(n10695) );
  XOR U14294 ( .A(n10698), .B(n10699), .Z(n10697) );
  XOR U14295 ( .A(DB[1315]), .B(DB[1300]), .Z(n10699) );
  AND U14296 ( .A(n678), .B(n10700), .Z(n10698) );
  XOR U14297 ( .A(n10701), .B(n10702), .Z(n10700) );
  XOR U14298 ( .A(DB[1300]), .B(DB[1285]), .Z(n10702) );
  AND U14299 ( .A(n682), .B(n10703), .Z(n10701) );
  XOR U14300 ( .A(n10704), .B(n10705), .Z(n10703) );
  XOR U14301 ( .A(DB[1285]), .B(DB[1270]), .Z(n10705) );
  AND U14302 ( .A(n686), .B(n10706), .Z(n10704) );
  XOR U14303 ( .A(n10707), .B(n10708), .Z(n10706) );
  XOR U14304 ( .A(DB[1270]), .B(DB[1255]), .Z(n10708) );
  AND U14305 ( .A(n690), .B(n10709), .Z(n10707) );
  XOR U14306 ( .A(n10710), .B(n10711), .Z(n10709) );
  XOR U14307 ( .A(DB[1255]), .B(DB[1240]), .Z(n10711) );
  AND U14308 ( .A(n694), .B(n10712), .Z(n10710) );
  XOR U14309 ( .A(n10713), .B(n10714), .Z(n10712) );
  XOR U14310 ( .A(DB[1240]), .B(DB[1225]), .Z(n10714) );
  AND U14311 ( .A(n698), .B(n10715), .Z(n10713) );
  XOR U14312 ( .A(n10716), .B(n10717), .Z(n10715) );
  XOR U14313 ( .A(DB[1225]), .B(DB[1210]), .Z(n10717) );
  AND U14314 ( .A(n702), .B(n10718), .Z(n10716) );
  XOR U14315 ( .A(n10719), .B(n10720), .Z(n10718) );
  XOR U14316 ( .A(DB[1210]), .B(DB[1195]), .Z(n10720) );
  AND U14317 ( .A(n706), .B(n10721), .Z(n10719) );
  XOR U14318 ( .A(n10722), .B(n10723), .Z(n10721) );
  XOR U14319 ( .A(DB[1195]), .B(DB[1180]), .Z(n10723) );
  AND U14320 ( .A(n710), .B(n10724), .Z(n10722) );
  XOR U14321 ( .A(n10725), .B(n10726), .Z(n10724) );
  XOR U14322 ( .A(DB[1180]), .B(DB[1165]), .Z(n10726) );
  AND U14323 ( .A(n714), .B(n10727), .Z(n10725) );
  XOR U14324 ( .A(n10728), .B(n10729), .Z(n10727) );
  XOR U14325 ( .A(DB[1165]), .B(DB[1150]), .Z(n10729) );
  AND U14326 ( .A(n718), .B(n10730), .Z(n10728) );
  XOR U14327 ( .A(n10731), .B(n10732), .Z(n10730) );
  XOR U14328 ( .A(DB[1150]), .B(DB[1135]), .Z(n10732) );
  AND U14329 ( .A(n722), .B(n10733), .Z(n10731) );
  XOR U14330 ( .A(n10734), .B(n10735), .Z(n10733) );
  XOR U14331 ( .A(DB[1135]), .B(DB[1120]), .Z(n10735) );
  AND U14332 ( .A(n726), .B(n10736), .Z(n10734) );
  XOR U14333 ( .A(n10737), .B(n10738), .Z(n10736) );
  XOR U14334 ( .A(DB[1120]), .B(DB[1105]), .Z(n10738) );
  AND U14335 ( .A(n730), .B(n10739), .Z(n10737) );
  XOR U14336 ( .A(n10740), .B(n10741), .Z(n10739) );
  XOR U14337 ( .A(DB[1105]), .B(DB[1090]), .Z(n10741) );
  AND U14338 ( .A(n734), .B(n10742), .Z(n10740) );
  XOR U14339 ( .A(n10743), .B(n10744), .Z(n10742) );
  XOR U14340 ( .A(DB[1090]), .B(DB[1075]), .Z(n10744) );
  AND U14341 ( .A(n738), .B(n10745), .Z(n10743) );
  XOR U14342 ( .A(n10746), .B(n10747), .Z(n10745) );
  XOR U14343 ( .A(DB[1075]), .B(DB[1060]), .Z(n10747) );
  AND U14344 ( .A(n742), .B(n10748), .Z(n10746) );
  XOR U14345 ( .A(n10749), .B(n10750), .Z(n10748) );
  XOR U14346 ( .A(DB[1060]), .B(DB[1045]), .Z(n10750) );
  AND U14347 ( .A(n746), .B(n10751), .Z(n10749) );
  XOR U14348 ( .A(n10752), .B(n10753), .Z(n10751) );
  XOR U14349 ( .A(DB[1045]), .B(DB[1030]), .Z(n10753) );
  AND U14350 ( .A(n750), .B(n10754), .Z(n10752) );
  XOR U14351 ( .A(n10755), .B(n10756), .Z(n10754) );
  XOR U14352 ( .A(DB[1030]), .B(DB[1015]), .Z(n10756) );
  AND U14353 ( .A(n754), .B(n10757), .Z(n10755) );
  XOR U14354 ( .A(n10758), .B(n10759), .Z(n10757) );
  XOR U14355 ( .A(DB[1015]), .B(DB[1000]), .Z(n10759) );
  AND U14356 ( .A(n758), .B(n10760), .Z(n10758) );
  XOR U14357 ( .A(n10761), .B(n10762), .Z(n10760) );
  XOR U14358 ( .A(DB[985]), .B(DB[1000]), .Z(n10762) );
  AND U14359 ( .A(n762), .B(n10763), .Z(n10761) );
  XOR U14360 ( .A(n10764), .B(n10765), .Z(n10763) );
  XOR U14361 ( .A(DB[985]), .B(DB[970]), .Z(n10765) );
  AND U14362 ( .A(n766), .B(n10766), .Z(n10764) );
  XOR U14363 ( .A(n10767), .B(n10768), .Z(n10766) );
  XOR U14364 ( .A(DB[970]), .B(DB[955]), .Z(n10768) );
  AND U14365 ( .A(n770), .B(n10769), .Z(n10767) );
  XOR U14366 ( .A(n10770), .B(n10771), .Z(n10769) );
  XOR U14367 ( .A(DB[955]), .B(DB[940]), .Z(n10771) );
  AND U14368 ( .A(n774), .B(n10772), .Z(n10770) );
  XOR U14369 ( .A(n10773), .B(n10774), .Z(n10772) );
  XOR U14370 ( .A(DB[940]), .B(DB[925]), .Z(n10774) );
  AND U14371 ( .A(n778), .B(n10775), .Z(n10773) );
  XOR U14372 ( .A(n10776), .B(n10777), .Z(n10775) );
  XOR U14373 ( .A(DB[925]), .B(DB[910]), .Z(n10777) );
  AND U14374 ( .A(n782), .B(n10778), .Z(n10776) );
  XOR U14375 ( .A(n10779), .B(n10780), .Z(n10778) );
  XOR U14376 ( .A(DB[910]), .B(DB[895]), .Z(n10780) );
  AND U14377 ( .A(n786), .B(n10781), .Z(n10779) );
  XOR U14378 ( .A(n10782), .B(n10783), .Z(n10781) );
  XOR U14379 ( .A(DB[895]), .B(DB[880]), .Z(n10783) );
  AND U14380 ( .A(n790), .B(n10784), .Z(n10782) );
  XOR U14381 ( .A(n10785), .B(n10786), .Z(n10784) );
  XOR U14382 ( .A(DB[880]), .B(DB[865]), .Z(n10786) );
  AND U14383 ( .A(n794), .B(n10787), .Z(n10785) );
  XOR U14384 ( .A(n10788), .B(n10789), .Z(n10787) );
  XOR U14385 ( .A(DB[865]), .B(DB[850]), .Z(n10789) );
  AND U14386 ( .A(n798), .B(n10790), .Z(n10788) );
  XOR U14387 ( .A(n10791), .B(n10792), .Z(n10790) );
  XOR U14388 ( .A(DB[850]), .B(DB[835]), .Z(n10792) );
  AND U14389 ( .A(n802), .B(n10793), .Z(n10791) );
  XOR U14390 ( .A(n10794), .B(n10795), .Z(n10793) );
  XOR U14391 ( .A(DB[835]), .B(DB[820]), .Z(n10795) );
  AND U14392 ( .A(n806), .B(n10796), .Z(n10794) );
  XOR U14393 ( .A(n10797), .B(n10798), .Z(n10796) );
  XOR U14394 ( .A(DB[820]), .B(DB[805]), .Z(n10798) );
  AND U14395 ( .A(n810), .B(n10799), .Z(n10797) );
  XOR U14396 ( .A(n10800), .B(n10801), .Z(n10799) );
  XOR U14397 ( .A(DB[805]), .B(DB[790]), .Z(n10801) );
  AND U14398 ( .A(n814), .B(n10802), .Z(n10800) );
  XOR U14399 ( .A(n10803), .B(n10804), .Z(n10802) );
  XOR U14400 ( .A(DB[790]), .B(DB[775]), .Z(n10804) );
  AND U14401 ( .A(n818), .B(n10805), .Z(n10803) );
  XOR U14402 ( .A(n10806), .B(n10807), .Z(n10805) );
  XOR U14403 ( .A(DB[775]), .B(DB[760]), .Z(n10807) );
  AND U14404 ( .A(n822), .B(n10808), .Z(n10806) );
  XOR U14405 ( .A(n10809), .B(n10810), .Z(n10808) );
  XOR U14406 ( .A(DB[760]), .B(DB[745]), .Z(n10810) );
  AND U14407 ( .A(n826), .B(n10811), .Z(n10809) );
  XOR U14408 ( .A(n10812), .B(n10813), .Z(n10811) );
  XOR U14409 ( .A(DB[745]), .B(DB[730]), .Z(n10813) );
  AND U14410 ( .A(n830), .B(n10814), .Z(n10812) );
  XOR U14411 ( .A(n10815), .B(n10816), .Z(n10814) );
  XOR U14412 ( .A(DB[730]), .B(DB[715]), .Z(n10816) );
  AND U14413 ( .A(n834), .B(n10817), .Z(n10815) );
  XOR U14414 ( .A(n10818), .B(n10819), .Z(n10817) );
  XOR U14415 ( .A(DB[715]), .B(DB[700]), .Z(n10819) );
  AND U14416 ( .A(n838), .B(n10820), .Z(n10818) );
  XOR U14417 ( .A(n10821), .B(n10822), .Z(n10820) );
  XOR U14418 ( .A(DB[700]), .B(DB[685]), .Z(n10822) );
  AND U14419 ( .A(n842), .B(n10823), .Z(n10821) );
  XOR U14420 ( .A(n10824), .B(n10825), .Z(n10823) );
  XOR U14421 ( .A(DB[685]), .B(DB[670]), .Z(n10825) );
  AND U14422 ( .A(n846), .B(n10826), .Z(n10824) );
  XOR U14423 ( .A(n10827), .B(n10828), .Z(n10826) );
  XOR U14424 ( .A(DB[670]), .B(DB[655]), .Z(n10828) );
  AND U14425 ( .A(n850), .B(n10829), .Z(n10827) );
  XOR U14426 ( .A(n10830), .B(n10831), .Z(n10829) );
  XOR U14427 ( .A(DB[655]), .B(DB[640]), .Z(n10831) );
  AND U14428 ( .A(n854), .B(n10832), .Z(n10830) );
  XOR U14429 ( .A(n10833), .B(n10834), .Z(n10832) );
  XOR U14430 ( .A(DB[640]), .B(DB[625]), .Z(n10834) );
  AND U14431 ( .A(n858), .B(n10835), .Z(n10833) );
  XOR U14432 ( .A(n10836), .B(n10837), .Z(n10835) );
  XOR U14433 ( .A(DB[625]), .B(DB[610]), .Z(n10837) );
  AND U14434 ( .A(n862), .B(n10838), .Z(n10836) );
  XOR U14435 ( .A(n10839), .B(n10840), .Z(n10838) );
  XOR U14436 ( .A(DB[610]), .B(DB[595]), .Z(n10840) );
  AND U14437 ( .A(n866), .B(n10841), .Z(n10839) );
  XOR U14438 ( .A(n10842), .B(n10843), .Z(n10841) );
  XOR U14439 ( .A(DB[595]), .B(DB[580]), .Z(n10843) );
  AND U14440 ( .A(n870), .B(n10844), .Z(n10842) );
  XOR U14441 ( .A(n10845), .B(n10846), .Z(n10844) );
  XOR U14442 ( .A(DB[580]), .B(DB[565]), .Z(n10846) );
  AND U14443 ( .A(n874), .B(n10847), .Z(n10845) );
  XOR U14444 ( .A(n10848), .B(n10849), .Z(n10847) );
  XOR U14445 ( .A(DB[565]), .B(DB[550]), .Z(n10849) );
  AND U14446 ( .A(n878), .B(n10850), .Z(n10848) );
  XOR U14447 ( .A(n10851), .B(n10852), .Z(n10850) );
  XOR U14448 ( .A(DB[550]), .B(DB[535]), .Z(n10852) );
  AND U14449 ( .A(n882), .B(n10853), .Z(n10851) );
  XOR U14450 ( .A(n10854), .B(n10855), .Z(n10853) );
  XOR U14451 ( .A(DB[535]), .B(DB[520]), .Z(n10855) );
  AND U14452 ( .A(n886), .B(n10856), .Z(n10854) );
  XOR U14453 ( .A(n10857), .B(n10858), .Z(n10856) );
  XOR U14454 ( .A(DB[520]), .B(DB[505]), .Z(n10858) );
  AND U14455 ( .A(n890), .B(n10859), .Z(n10857) );
  XOR U14456 ( .A(n10860), .B(n10861), .Z(n10859) );
  XOR U14457 ( .A(DB[505]), .B(DB[490]), .Z(n10861) );
  AND U14458 ( .A(n894), .B(n10862), .Z(n10860) );
  XOR U14459 ( .A(n10863), .B(n10864), .Z(n10862) );
  XOR U14460 ( .A(DB[490]), .B(DB[475]), .Z(n10864) );
  AND U14461 ( .A(n898), .B(n10865), .Z(n10863) );
  XOR U14462 ( .A(n10866), .B(n10867), .Z(n10865) );
  XOR U14463 ( .A(DB[475]), .B(DB[460]), .Z(n10867) );
  AND U14464 ( .A(n902), .B(n10868), .Z(n10866) );
  XOR U14465 ( .A(n10869), .B(n10870), .Z(n10868) );
  XOR U14466 ( .A(DB[460]), .B(DB[445]), .Z(n10870) );
  AND U14467 ( .A(n906), .B(n10871), .Z(n10869) );
  XOR U14468 ( .A(n10872), .B(n10873), .Z(n10871) );
  XOR U14469 ( .A(DB[445]), .B(DB[430]), .Z(n10873) );
  AND U14470 ( .A(n910), .B(n10874), .Z(n10872) );
  XOR U14471 ( .A(n10875), .B(n10876), .Z(n10874) );
  XOR U14472 ( .A(DB[430]), .B(DB[415]), .Z(n10876) );
  AND U14473 ( .A(n914), .B(n10877), .Z(n10875) );
  XOR U14474 ( .A(n10878), .B(n10879), .Z(n10877) );
  XOR U14475 ( .A(DB[415]), .B(DB[400]), .Z(n10879) );
  AND U14476 ( .A(n918), .B(n10880), .Z(n10878) );
  XOR U14477 ( .A(n10881), .B(n10882), .Z(n10880) );
  XOR U14478 ( .A(DB[400]), .B(DB[385]), .Z(n10882) );
  AND U14479 ( .A(n922), .B(n10883), .Z(n10881) );
  XOR U14480 ( .A(n10884), .B(n10885), .Z(n10883) );
  XOR U14481 ( .A(DB[385]), .B(DB[370]), .Z(n10885) );
  AND U14482 ( .A(n926), .B(n10886), .Z(n10884) );
  XOR U14483 ( .A(n10887), .B(n10888), .Z(n10886) );
  XOR U14484 ( .A(DB[370]), .B(DB[355]), .Z(n10888) );
  AND U14485 ( .A(n930), .B(n10889), .Z(n10887) );
  XOR U14486 ( .A(n10890), .B(n10891), .Z(n10889) );
  XOR U14487 ( .A(DB[355]), .B(DB[340]), .Z(n10891) );
  AND U14488 ( .A(n934), .B(n10892), .Z(n10890) );
  XOR U14489 ( .A(n10893), .B(n10894), .Z(n10892) );
  XOR U14490 ( .A(DB[340]), .B(DB[325]), .Z(n10894) );
  AND U14491 ( .A(n938), .B(n10895), .Z(n10893) );
  XOR U14492 ( .A(n10896), .B(n10897), .Z(n10895) );
  XOR U14493 ( .A(DB[325]), .B(DB[310]), .Z(n10897) );
  AND U14494 ( .A(n942), .B(n10898), .Z(n10896) );
  XOR U14495 ( .A(n10899), .B(n10900), .Z(n10898) );
  XOR U14496 ( .A(DB[310]), .B(DB[295]), .Z(n10900) );
  AND U14497 ( .A(n946), .B(n10901), .Z(n10899) );
  XOR U14498 ( .A(n10902), .B(n10903), .Z(n10901) );
  XOR U14499 ( .A(DB[295]), .B(DB[280]), .Z(n10903) );
  AND U14500 ( .A(n950), .B(n10904), .Z(n10902) );
  XOR U14501 ( .A(n10905), .B(n10906), .Z(n10904) );
  XOR U14502 ( .A(DB[280]), .B(DB[265]), .Z(n10906) );
  AND U14503 ( .A(n954), .B(n10907), .Z(n10905) );
  XOR U14504 ( .A(n10908), .B(n10909), .Z(n10907) );
  XOR U14505 ( .A(DB[265]), .B(DB[250]), .Z(n10909) );
  AND U14506 ( .A(n958), .B(n10910), .Z(n10908) );
  XOR U14507 ( .A(n10911), .B(n10912), .Z(n10910) );
  XOR U14508 ( .A(DB[250]), .B(DB[235]), .Z(n10912) );
  AND U14509 ( .A(n962), .B(n10913), .Z(n10911) );
  XOR U14510 ( .A(n10914), .B(n10915), .Z(n10913) );
  XOR U14511 ( .A(DB[235]), .B(DB[220]), .Z(n10915) );
  AND U14512 ( .A(n966), .B(n10916), .Z(n10914) );
  XOR U14513 ( .A(n10917), .B(n10918), .Z(n10916) );
  XOR U14514 ( .A(DB[220]), .B(DB[205]), .Z(n10918) );
  AND U14515 ( .A(n970), .B(n10919), .Z(n10917) );
  XOR U14516 ( .A(n10920), .B(n10921), .Z(n10919) );
  XOR U14517 ( .A(DB[205]), .B(DB[190]), .Z(n10921) );
  AND U14518 ( .A(n974), .B(n10922), .Z(n10920) );
  XOR U14519 ( .A(n10923), .B(n10924), .Z(n10922) );
  XOR U14520 ( .A(DB[190]), .B(DB[175]), .Z(n10924) );
  AND U14521 ( .A(n978), .B(n10925), .Z(n10923) );
  XOR U14522 ( .A(n10926), .B(n10927), .Z(n10925) );
  XOR U14523 ( .A(DB[175]), .B(DB[160]), .Z(n10927) );
  AND U14524 ( .A(n982), .B(n10928), .Z(n10926) );
  XOR U14525 ( .A(n10929), .B(n10930), .Z(n10928) );
  XOR U14526 ( .A(DB[160]), .B(DB[145]), .Z(n10930) );
  AND U14527 ( .A(n986), .B(n10931), .Z(n10929) );
  XOR U14528 ( .A(n10932), .B(n10933), .Z(n10931) );
  XOR U14529 ( .A(DB[145]), .B(DB[130]), .Z(n10933) );
  AND U14530 ( .A(n990), .B(n10934), .Z(n10932) );
  XOR U14531 ( .A(n10935), .B(n10936), .Z(n10934) );
  XOR U14532 ( .A(DB[130]), .B(DB[115]), .Z(n10936) );
  AND U14533 ( .A(n994), .B(n10937), .Z(n10935) );
  XOR U14534 ( .A(n10938), .B(n10939), .Z(n10937) );
  XOR U14535 ( .A(DB[115]), .B(DB[100]), .Z(n10939) );
  AND U14536 ( .A(n998), .B(n10940), .Z(n10938) );
  XOR U14537 ( .A(n10941), .B(n10942), .Z(n10940) );
  XOR U14538 ( .A(DB[85]), .B(DB[100]), .Z(n10942) );
  AND U14539 ( .A(n1002), .B(n10943), .Z(n10941) );
  XOR U14540 ( .A(n10944), .B(n10945), .Z(n10943) );
  XOR U14541 ( .A(DB[85]), .B(DB[70]), .Z(n10945) );
  AND U14542 ( .A(n1006), .B(n10946), .Z(n10944) );
  XOR U14543 ( .A(n10947), .B(n10948), .Z(n10946) );
  XOR U14544 ( .A(DB[70]), .B(DB[55]), .Z(n10948) );
  AND U14545 ( .A(n1010), .B(n10949), .Z(n10947) );
  XOR U14546 ( .A(n10950), .B(n10951), .Z(n10949) );
  XOR U14547 ( .A(DB[55]), .B(DB[40]), .Z(n10951) );
  AND U14548 ( .A(n1014), .B(n10952), .Z(n10950) );
  XOR U14549 ( .A(n10953), .B(n10954), .Z(n10952) );
  XOR U14550 ( .A(DB[40]), .B(DB[25]), .Z(n10954) );
  AND U14551 ( .A(n1018), .B(n10955), .Z(n10953) );
  XOR U14552 ( .A(DB[25]), .B(DB[10]), .Z(n10955) );
  XOR U14553 ( .A(DB[3825]), .B(n10956), .Z(min_val_out[0]) );
  AND U14554 ( .A(n2), .B(n10957), .Z(n10956) );
  XOR U14555 ( .A(n10958), .B(n10959), .Z(n10957) );
  XOR U14556 ( .A(DB[3825]), .B(DB[3810]), .Z(n10959) );
  AND U14557 ( .A(n6), .B(n10960), .Z(n10958) );
  XOR U14558 ( .A(n10961), .B(n10962), .Z(n10960) );
  XOR U14559 ( .A(DB[3810]), .B(DB[3795]), .Z(n10962) );
  AND U14560 ( .A(n10), .B(n10963), .Z(n10961) );
  XOR U14561 ( .A(n10964), .B(n10965), .Z(n10963) );
  XOR U14562 ( .A(DB[3795]), .B(DB[3780]), .Z(n10965) );
  AND U14563 ( .A(n14), .B(n10966), .Z(n10964) );
  XOR U14564 ( .A(n10967), .B(n10968), .Z(n10966) );
  XOR U14565 ( .A(DB[3780]), .B(DB[3765]), .Z(n10968) );
  AND U14566 ( .A(n18), .B(n10969), .Z(n10967) );
  XOR U14567 ( .A(n10970), .B(n10971), .Z(n10969) );
  XOR U14568 ( .A(DB[3765]), .B(DB[3750]), .Z(n10971) );
  AND U14569 ( .A(n22), .B(n10972), .Z(n10970) );
  XOR U14570 ( .A(n10973), .B(n10974), .Z(n10972) );
  XOR U14571 ( .A(DB[3750]), .B(DB[3735]), .Z(n10974) );
  AND U14572 ( .A(n26), .B(n10975), .Z(n10973) );
  XOR U14573 ( .A(n10976), .B(n10977), .Z(n10975) );
  XOR U14574 ( .A(DB[3735]), .B(DB[3720]), .Z(n10977) );
  AND U14575 ( .A(n30), .B(n10978), .Z(n10976) );
  XOR U14576 ( .A(n10979), .B(n10980), .Z(n10978) );
  XOR U14577 ( .A(DB[3720]), .B(DB[3705]), .Z(n10980) );
  AND U14578 ( .A(n34), .B(n10981), .Z(n10979) );
  XOR U14579 ( .A(n10982), .B(n10983), .Z(n10981) );
  XOR U14580 ( .A(DB[3705]), .B(DB[3690]), .Z(n10983) );
  AND U14581 ( .A(n38), .B(n10984), .Z(n10982) );
  XOR U14582 ( .A(n10985), .B(n10986), .Z(n10984) );
  XOR U14583 ( .A(DB[3690]), .B(DB[3675]), .Z(n10986) );
  AND U14584 ( .A(n42), .B(n10987), .Z(n10985) );
  XOR U14585 ( .A(n10988), .B(n10989), .Z(n10987) );
  XOR U14586 ( .A(DB[3675]), .B(DB[3660]), .Z(n10989) );
  AND U14587 ( .A(n46), .B(n10990), .Z(n10988) );
  XOR U14588 ( .A(n10991), .B(n10992), .Z(n10990) );
  XOR U14589 ( .A(DB[3660]), .B(DB[3645]), .Z(n10992) );
  AND U14590 ( .A(n50), .B(n10993), .Z(n10991) );
  XOR U14591 ( .A(n10994), .B(n10995), .Z(n10993) );
  XOR U14592 ( .A(DB[3645]), .B(DB[3630]), .Z(n10995) );
  AND U14593 ( .A(n54), .B(n10996), .Z(n10994) );
  XOR U14594 ( .A(n10997), .B(n10998), .Z(n10996) );
  XOR U14595 ( .A(DB[3630]), .B(DB[3615]), .Z(n10998) );
  AND U14596 ( .A(n58), .B(n10999), .Z(n10997) );
  XOR U14597 ( .A(n11000), .B(n11001), .Z(n10999) );
  XOR U14598 ( .A(DB[3615]), .B(DB[3600]), .Z(n11001) );
  AND U14599 ( .A(n62), .B(n11002), .Z(n11000) );
  XOR U14600 ( .A(n11003), .B(n11004), .Z(n11002) );
  XOR U14601 ( .A(DB[3600]), .B(DB[3585]), .Z(n11004) );
  AND U14602 ( .A(n66), .B(n11005), .Z(n11003) );
  XOR U14603 ( .A(n11006), .B(n11007), .Z(n11005) );
  XOR U14604 ( .A(DB[3585]), .B(DB[3570]), .Z(n11007) );
  AND U14605 ( .A(n70), .B(n11008), .Z(n11006) );
  XOR U14606 ( .A(n11009), .B(n11010), .Z(n11008) );
  XOR U14607 ( .A(DB[3570]), .B(DB[3555]), .Z(n11010) );
  AND U14608 ( .A(n74), .B(n11011), .Z(n11009) );
  XOR U14609 ( .A(n11012), .B(n11013), .Z(n11011) );
  XOR U14610 ( .A(DB[3555]), .B(DB[3540]), .Z(n11013) );
  AND U14611 ( .A(n78), .B(n11014), .Z(n11012) );
  XOR U14612 ( .A(n11015), .B(n11016), .Z(n11014) );
  XOR U14613 ( .A(DB[3540]), .B(DB[3525]), .Z(n11016) );
  AND U14614 ( .A(n82), .B(n11017), .Z(n11015) );
  XOR U14615 ( .A(n11018), .B(n11019), .Z(n11017) );
  XOR U14616 ( .A(DB[3525]), .B(DB[3510]), .Z(n11019) );
  AND U14617 ( .A(n86), .B(n11020), .Z(n11018) );
  XOR U14618 ( .A(n11021), .B(n11022), .Z(n11020) );
  XOR U14619 ( .A(DB[3510]), .B(DB[3495]), .Z(n11022) );
  AND U14620 ( .A(n90), .B(n11023), .Z(n11021) );
  XOR U14621 ( .A(n11024), .B(n11025), .Z(n11023) );
  XOR U14622 ( .A(DB[3495]), .B(DB[3480]), .Z(n11025) );
  AND U14623 ( .A(n94), .B(n11026), .Z(n11024) );
  XOR U14624 ( .A(n11027), .B(n11028), .Z(n11026) );
  XOR U14625 ( .A(DB[3480]), .B(DB[3465]), .Z(n11028) );
  AND U14626 ( .A(n98), .B(n11029), .Z(n11027) );
  XOR U14627 ( .A(n11030), .B(n11031), .Z(n11029) );
  XOR U14628 ( .A(DB[3465]), .B(DB[3450]), .Z(n11031) );
  AND U14629 ( .A(n102), .B(n11032), .Z(n11030) );
  XOR U14630 ( .A(n11033), .B(n11034), .Z(n11032) );
  XOR U14631 ( .A(DB[3450]), .B(DB[3435]), .Z(n11034) );
  AND U14632 ( .A(n106), .B(n11035), .Z(n11033) );
  XOR U14633 ( .A(n11036), .B(n11037), .Z(n11035) );
  XOR U14634 ( .A(DB[3435]), .B(DB[3420]), .Z(n11037) );
  AND U14635 ( .A(n110), .B(n11038), .Z(n11036) );
  XOR U14636 ( .A(n11039), .B(n11040), .Z(n11038) );
  XOR U14637 ( .A(DB[3420]), .B(DB[3405]), .Z(n11040) );
  AND U14638 ( .A(n114), .B(n11041), .Z(n11039) );
  XOR U14639 ( .A(n11042), .B(n11043), .Z(n11041) );
  XOR U14640 ( .A(DB[3405]), .B(DB[3390]), .Z(n11043) );
  AND U14641 ( .A(n118), .B(n11044), .Z(n11042) );
  XOR U14642 ( .A(n11045), .B(n11046), .Z(n11044) );
  XOR U14643 ( .A(DB[3390]), .B(DB[3375]), .Z(n11046) );
  AND U14644 ( .A(n122), .B(n11047), .Z(n11045) );
  XOR U14645 ( .A(n11048), .B(n11049), .Z(n11047) );
  XOR U14646 ( .A(DB[3375]), .B(DB[3360]), .Z(n11049) );
  AND U14647 ( .A(n126), .B(n11050), .Z(n11048) );
  XOR U14648 ( .A(n11051), .B(n11052), .Z(n11050) );
  XOR U14649 ( .A(DB[3360]), .B(DB[3345]), .Z(n11052) );
  AND U14650 ( .A(n130), .B(n11053), .Z(n11051) );
  XOR U14651 ( .A(n11054), .B(n11055), .Z(n11053) );
  XOR U14652 ( .A(DB[3345]), .B(DB[3330]), .Z(n11055) );
  AND U14653 ( .A(n134), .B(n11056), .Z(n11054) );
  XOR U14654 ( .A(n11057), .B(n11058), .Z(n11056) );
  XOR U14655 ( .A(DB[3330]), .B(DB[3315]), .Z(n11058) );
  AND U14656 ( .A(n138), .B(n11059), .Z(n11057) );
  XOR U14657 ( .A(n11060), .B(n11061), .Z(n11059) );
  XOR U14658 ( .A(DB[3315]), .B(DB[3300]), .Z(n11061) );
  AND U14659 ( .A(n142), .B(n11062), .Z(n11060) );
  XOR U14660 ( .A(n11063), .B(n11064), .Z(n11062) );
  XOR U14661 ( .A(DB[3300]), .B(DB[3285]), .Z(n11064) );
  AND U14662 ( .A(n146), .B(n11065), .Z(n11063) );
  XOR U14663 ( .A(n11066), .B(n11067), .Z(n11065) );
  XOR U14664 ( .A(DB[3285]), .B(DB[3270]), .Z(n11067) );
  AND U14665 ( .A(n150), .B(n11068), .Z(n11066) );
  XOR U14666 ( .A(n11069), .B(n11070), .Z(n11068) );
  XOR U14667 ( .A(DB[3270]), .B(DB[3255]), .Z(n11070) );
  AND U14668 ( .A(n154), .B(n11071), .Z(n11069) );
  XOR U14669 ( .A(n11072), .B(n11073), .Z(n11071) );
  XOR U14670 ( .A(DB[3255]), .B(DB[3240]), .Z(n11073) );
  AND U14671 ( .A(n158), .B(n11074), .Z(n11072) );
  XOR U14672 ( .A(n11075), .B(n11076), .Z(n11074) );
  XOR U14673 ( .A(DB[3240]), .B(DB[3225]), .Z(n11076) );
  AND U14674 ( .A(n162), .B(n11077), .Z(n11075) );
  XOR U14675 ( .A(n11078), .B(n11079), .Z(n11077) );
  XOR U14676 ( .A(DB[3225]), .B(DB[3210]), .Z(n11079) );
  AND U14677 ( .A(n166), .B(n11080), .Z(n11078) );
  XOR U14678 ( .A(n11081), .B(n11082), .Z(n11080) );
  XOR U14679 ( .A(DB[3210]), .B(DB[3195]), .Z(n11082) );
  AND U14680 ( .A(n170), .B(n11083), .Z(n11081) );
  XOR U14681 ( .A(n11084), .B(n11085), .Z(n11083) );
  XOR U14682 ( .A(DB[3195]), .B(DB[3180]), .Z(n11085) );
  AND U14683 ( .A(n174), .B(n11086), .Z(n11084) );
  XOR U14684 ( .A(n11087), .B(n11088), .Z(n11086) );
  XOR U14685 ( .A(DB[3180]), .B(DB[3165]), .Z(n11088) );
  AND U14686 ( .A(n178), .B(n11089), .Z(n11087) );
  XOR U14687 ( .A(n11090), .B(n11091), .Z(n11089) );
  XOR U14688 ( .A(DB[3165]), .B(DB[3150]), .Z(n11091) );
  AND U14689 ( .A(n182), .B(n11092), .Z(n11090) );
  XOR U14690 ( .A(n11093), .B(n11094), .Z(n11092) );
  XOR U14691 ( .A(DB[3150]), .B(DB[3135]), .Z(n11094) );
  AND U14692 ( .A(n186), .B(n11095), .Z(n11093) );
  XOR U14693 ( .A(n11096), .B(n11097), .Z(n11095) );
  XOR U14694 ( .A(DB[3135]), .B(DB[3120]), .Z(n11097) );
  AND U14695 ( .A(n190), .B(n11098), .Z(n11096) );
  XOR U14696 ( .A(n11099), .B(n11100), .Z(n11098) );
  XOR U14697 ( .A(DB[3120]), .B(DB[3105]), .Z(n11100) );
  AND U14698 ( .A(n194), .B(n11101), .Z(n11099) );
  XOR U14699 ( .A(n11102), .B(n11103), .Z(n11101) );
  XOR U14700 ( .A(DB[3105]), .B(DB[3090]), .Z(n11103) );
  AND U14701 ( .A(n198), .B(n11104), .Z(n11102) );
  XOR U14702 ( .A(n11105), .B(n11106), .Z(n11104) );
  XOR U14703 ( .A(DB[3090]), .B(DB[3075]), .Z(n11106) );
  AND U14704 ( .A(n202), .B(n11107), .Z(n11105) );
  XOR U14705 ( .A(n11108), .B(n11109), .Z(n11107) );
  XOR U14706 ( .A(DB[3075]), .B(DB[3060]), .Z(n11109) );
  AND U14707 ( .A(n206), .B(n11110), .Z(n11108) );
  XOR U14708 ( .A(n11111), .B(n11112), .Z(n11110) );
  XOR U14709 ( .A(DB[3060]), .B(DB[3045]), .Z(n11112) );
  AND U14710 ( .A(n210), .B(n11113), .Z(n11111) );
  XOR U14711 ( .A(n11114), .B(n11115), .Z(n11113) );
  XOR U14712 ( .A(DB[3045]), .B(DB[3030]), .Z(n11115) );
  AND U14713 ( .A(n214), .B(n11116), .Z(n11114) );
  XOR U14714 ( .A(n11117), .B(n11118), .Z(n11116) );
  XOR U14715 ( .A(DB[3030]), .B(DB[3015]), .Z(n11118) );
  AND U14716 ( .A(n218), .B(n11119), .Z(n11117) );
  XOR U14717 ( .A(n11120), .B(n11121), .Z(n11119) );
  XOR U14718 ( .A(DB[3015]), .B(DB[3000]), .Z(n11121) );
  AND U14719 ( .A(n222), .B(n11122), .Z(n11120) );
  XOR U14720 ( .A(n11123), .B(n11124), .Z(n11122) );
  XOR U14721 ( .A(DB[3000]), .B(DB[2985]), .Z(n11124) );
  AND U14722 ( .A(n226), .B(n11125), .Z(n11123) );
  XOR U14723 ( .A(n11126), .B(n11127), .Z(n11125) );
  XOR U14724 ( .A(DB[2985]), .B(DB[2970]), .Z(n11127) );
  AND U14725 ( .A(n230), .B(n11128), .Z(n11126) );
  XOR U14726 ( .A(n11129), .B(n11130), .Z(n11128) );
  XOR U14727 ( .A(DB[2970]), .B(DB[2955]), .Z(n11130) );
  AND U14728 ( .A(n234), .B(n11131), .Z(n11129) );
  XOR U14729 ( .A(n11132), .B(n11133), .Z(n11131) );
  XOR U14730 ( .A(DB[2955]), .B(DB[2940]), .Z(n11133) );
  AND U14731 ( .A(n238), .B(n11134), .Z(n11132) );
  XOR U14732 ( .A(n11135), .B(n11136), .Z(n11134) );
  XOR U14733 ( .A(DB[2940]), .B(DB[2925]), .Z(n11136) );
  AND U14734 ( .A(n242), .B(n11137), .Z(n11135) );
  XOR U14735 ( .A(n11138), .B(n11139), .Z(n11137) );
  XOR U14736 ( .A(DB[2925]), .B(DB[2910]), .Z(n11139) );
  AND U14737 ( .A(n246), .B(n11140), .Z(n11138) );
  XOR U14738 ( .A(n11141), .B(n11142), .Z(n11140) );
  XOR U14739 ( .A(DB[2910]), .B(DB[2895]), .Z(n11142) );
  AND U14740 ( .A(n250), .B(n11143), .Z(n11141) );
  XOR U14741 ( .A(n11144), .B(n11145), .Z(n11143) );
  XOR U14742 ( .A(DB[2895]), .B(DB[2880]), .Z(n11145) );
  AND U14743 ( .A(n254), .B(n11146), .Z(n11144) );
  XOR U14744 ( .A(n11147), .B(n11148), .Z(n11146) );
  XOR U14745 ( .A(DB[2880]), .B(DB[2865]), .Z(n11148) );
  AND U14746 ( .A(n258), .B(n11149), .Z(n11147) );
  XOR U14747 ( .A(n11150), .B(n11151), .Z(n11149) );
  XOR U14748 ( .A(DB[2865]), .B(DB[2850]), .Z(n11151) );
  AND U14749 ( .A(n262), .B(n11152), .Z(n11150) );
  XOR U14750 ( .A(n11153), .B(n11154), .Z(n11152) );
  XOR U14751 ( .A(DB[2850]), .B(DB[2835]), .Z(n11154) );
  AND U14752 ( .A(n266), .B(n11155), .Z(n11153) );
  XOR U14753 ( .A(n11156), .B(n11157), .Z(n11155) );
  XOR U14754 ( .A(DB[2835]), .B(DB[2820]), .Z(n11157) );
  AND U14755 ( .A(n270), .B(n11158), .Z(n11156) );
  XOR U14756 ( .A(n11159), .B(n11160), .Z(n11158) );
  XOR U14757 ( .A(DB[2820]), .B(DB[2805]), .Z(n11160) );
  AND U14758 ( .A(n274), .B(n11161), .Z(n11159) );
  XOR U14759 ( .A(n11162), .B(n11163), .Z(n11161) );
  XOR U14760 ( .A(DB[2805]), .B(DB[2790]), .Z(n11163) );
  AND U14761 ( .A(n278), .B(n11164), .Z(n11162) );
  XOR U14762 ( .A(n11165), .B(n11166), .Z(n11164) );
  XOR U14763 ( .A(DB[2790]), .B(DB[2775]), .Z(n11166) );
  AND U14764 ( .A(n282), .B(n11167), .Z(n11165) );
  XOR U14765 ( .A(n11168), .B(n11169), .Z(n11167) );
  XOR U14766 ( .A(DB[2775]), .B(DB[2760]), .Z(n11169) );
  AND U14767 ( .A(n286), .B(n11170), .Z(n11168) );
  XOR U14768 ( .A(n11171), .B(n11172), .Z(n11170) );
  XOR U14769 ( .A(DB[2760]), .B(DB[2745]), .Z(n11172) );
  AND U14770 ( .A(n290), .B(n11173), .Z(n11171) );
  XOR U14771 ( .A(n11174), .B(n11175), .Z(n11173) );
  XOR U14772 ( .A(DB[2745]), .B(DB[2730]), .Z(n11175) );
  AND U14773 ( .A(n294), .B(n11176), .Z(n11174) );
  XOR U14774 ( .A(n11177), .B(n11178), .Z(n11176) );
  XOR U14775 ( .A(DB[2730]), .B(DB[2715]), .Z(n11178) );
  AND U14776 ( .A(n298), .B(n11179), .Z(n11177) );
  XOR U14777 ( .A(n11180), .B(n11181), .Z(n11179) );
  XOR U14778 ( .A(DB[2715]), .B(DB[2700]), .Z(n11181) );
  AND U14779 ( .A(n302), .B(n11182), .Z(n11180) );
  XOR U14780 ( .A(n11183), .B(n11184), .Z(n11182) );
  XOR U14781 ( .A(DB[2700]), .B(DB[2685]), .Z(n11184) );
  AND U14782 ( .A(n306), .B(n11185), .Z(n11183) );
  XOR U14783 ( .A(n11186), .B(n11187), .Z(n11185) );
  XOR U14784 ( .A(DB[2685]), .B(DB[2670]), .Z(n11187) );
  AND U14785 ( .A(n310), .B(n11188), .Z(n11186) );
  XOR U14786 ( .A(n11189), .B(n11190), .Z(n11188) );
  XOR U14787 ( .A(DB[2670]), .B(DB[2655]), .Z(n11190) );
  AND U14788 ( .A(n314), .B(n11191), .Z(n11189) );
  XOR U14789 ( .A(n11192), .B(n11193), .Z(n11191) );
  XOR U14790 ( .A(DB[2655]), .B(DB[2640]), .Z(n11193) );
  AND U14791 ( .A(n318), .B(n11194), .Z(n11192) );
  XOR U14792 ( .A(n11195), .B(n11196), .Z(n11194) );
  XOR U14793 ( .A(DB[2640]), .B(DB[2625]), .Z(n11196) );
  AND U14794 ( .A(n322), .B(n11197), .Z(n11195) );
  XOR U14795 ( .A(n11198), .B(n11199), .Z(n11197) );
  XOR U14796 ( .A(DB[2625]), .B(DB[2610]), .Z(n11199) );
  AND U14797 ( .A(n326), .B(n11200), .Z(n11198) );
  XOR U14798 ( .A(n11201), .B(n11202), .Z(n11200) );
  XOR U14799 ( .A(DB[2610]), .B(DB[2595]), .Z(n11202) );
  AND U14800 ( .A(n330), .B(n11203), .Z(n11201) );
  XOR U14801 ( .A(n11204), .B(n11205), .Z(n11203) );
  XOR U14802 ( .A(DB[2595]), .B(DB[2580]), .Z(n11205) );
  AND U14803 ( .A(n334), .B(n11206), .Z(n11204) );
  XOR U14804 ( .A(n11207), .B(n11208), .Z(n11206) );
  XOR U14805 ( .A(DB[2580]), .B(DB[2565]), .Z(n11208) );
  AND U14806 ( .A(n338), .B(n11209), .Z(n11207) );
  XOR U14807 ( .A(n11210), .B(n11211), .Z(n11209) );
  XOR U14808 ( .A(DB[2565]), .B(DB[2550]), .Z(n11211) );
  AND U14809 ( .A(n342), .B(n11212), .Z(n11210) );
  XOR U14810 ( .A(n11213), .B(n11214), .Z(n11212) );
  XOR U14811 ( .A(DB[2550]), .B(DB[2535]), .Z(n11214) );
  AND U14812 ( .A(n346), .B(n11215), .Z(n11213) );
  XOR U14813 ( .A(n11216), .B(n11217), .Z(n11215) );
  XOR U14814 ( .A(DB[2535]), .B(DB[2520]), .Z(n11217) );
  AND U14815 ( .A(n350), .B(n11218), .Z(n11216) );
  XOR U14816 ( .A(n11219), .B(n11220), .Z(n11218) );
  XOR U14817 ( .A(DB[2520]), .B(DB[2505]), .Z(n11220) );
  AND U14818 ( .A(n354), .B(n11221), .Z(n11219) );
  XOR U14819 ( .A(n11222), .B(n11223), .Z(n11221) );
  XOR U14820 ( .A(DB[2505]), .B(DB[2490]), .Z(n11223) );
  AND U14821 ( .A(n358), .B(n11224), .Z(n11222) );
  XOR U14822 ( .A(n11225), .B(n11226), .Z(n11224) );
  XOR U14823 ( .A(DB[2490]), .B(DB[2475]), .Z(n11226) );
  AND U14824 ( .A(n362), .B(n11227), .Z(n11225) );
  XOR U14825 ( .A(n11228), .B(n11229), .Z(n11227) );
  XOR U14826 ( .A(DB[2475]), .B(DB[2460]), .Z(n11229) );
  AND U14827 ( .A(n366), .B(n11230), .Z(n11228) );
  XOR U14828 ( .A(n11231), .B(n11232), .Z(n11230) );
  XOR U14829 ( .A(DB[2460]), .B(DB[2445]), .Z(n11232) );
  AND U14830 ( .A(n370), .B(n11233), .Z(n11231) );
  XOR U14831 ( .A(n11234), .B(n11235), .Z(n11233) );
  XOR U14832 ( .A(DB[2445]), .B(DB[2430]), .Z(n11235) );
  AND U14833 ( .A(n374), .B(n11236), .Z(n11234) );
  XOR U14834 ( .A(n11237), .B(n11238), .Z(n11236) );
  XOR U14835 ( .A(DB[2430]), .B(DB[2415]), .Z(n11238) );
  AND U14836 ( .A(n378), .B(n11239), .Z(n11237) );
  XOR U14837 ( .A(n11240), .B(n11241), .Z(n11239) );
  XOR U14838 ( .A(DB[2415]), .B(DB[2400]), .Z(n11241) );
  AND U14839 ( .A(n382), .B(n11242), .Z(n11240) );
  XOR U14840 ( .A(n11243), .B(n11244), .Z(n11242) );
  XOR U14841 ( .A(DB[2400]), .B(DB[2385]), .Z(n11244) );
  AND U14842 ( .A(n386), .B(n11245), .Z(n11243) );
  XOR U14843 ( .A(n11246), .B(n11247), .Z(n11245) );
  XOR U14844 ( .A(DB[2385]), .B(DB[2370]), .Z(n11247) );
  AND U14845 ( .A(n390), .B(n11248), .Z(n11246) );
  XOR U14846 ( .A(n11249), .B(n11250), .Z(n11248) );
  XOR U14847 ( .A(DB[2370]), .B(DB[2355]), .Z(n11250) );
  AND U14848 ( .A(n394), .B(n11251), .Z(n11249) );
  XOR U14849 ( .A(n11252), .B(n11253), .Z(n11251) );
  XOR U14850 ( .A(DB[2355]), .B(DB[2340]), .Z(n11253) );
  AND U14851 ( .A(n398), .B(n11254), .Z(n11252) );
  XOR U14852 ( .A(n11255), .B(n11256), .Z(n11254) );
  XOR U14853 ( .A(DB[2340]), .B(DB[2325]), .Z(n11256) );
  AND U14854 ( .A(n402), .B(n11257), .Z(n11255) );
  XOR U14855 ( .A(n11258), .B(n11259), .Z(n11257) );
  XOR U14856 ( .A(DB[2325]), .B(DB[2310]), .Z(n11259) );
  AND U14857 ( .A(n406), .B(n11260), .Z(n11258) );
  XOR U14858 ( .A(n11261), .B(n11262), .Z(n11260) );
  XOR U14859 ( .A(DB[2310]), .B(DB[2295]), .Z(n11262) );
  AND U14860 ( .A(n410), .B(n11263), .Z(n11261) );
  XOR U14861 ( .A(n11264), .B(n11265), .Z(n11263) );
  XOR U14862 ( .A(DB[2295]), .B(DB[2280]), .Z(n11265) );
  AND U14863 ( .A(n414), .B(n11266), .Z(n11264) );
  XOR U14864 ( .A(n11267), .B(n11268), .Z(n11266) );
  XOR U14865 ( .A(DB[2280]), .B(DB[2265]), .Z(n11268) );
  AND U14866 ( .A(n418), .B(n11269), .Z(n11267) );
  XOR U14867 ( .A(n11270), .B(n11271), .Z(n11269) );
  XOR U14868 ( .A(DB[2265]), .B(DB[2250]), .Z(n11271) );
  AND U14869 ( .A(n422), .B(n11272), .Z(n11270) );
  XOR U14870 ( .A(n11273), .B(n11274), .Z(n11272) );
  XOR U14871 ( .A(DB[2250]), .B(DB[2235]), .Z(n11274) );
  AND U14872 ( .A(n426), .B(n11275), .Z(n11273) );
  XOR U14873 ( .A(n11276), .B(n11277), .Z(n11275) );
  XOR U14874 ( .A(DB[2235]), .B(DB[2220]), .Z(n11277) );
  AND U14875 ( .A(n430), .B(n11278), .Z(n11276) );
  XOR U14876 ( .A(n11279), .B(n11280), .Z(n11278) );
  XOR U14877 ( .A(DB[2220]), .B(DB[2205]), .Z(n11280) );
  AND U14878 ( .A(n434), .B(n11281), .Z(n11279) );
  XOR U14879 ( .A(n11282), .B(n11283), .Z(n11281) );
  XOR U14880 ( .A(DB[2205]), .B(DB[2190]), .Z(n11283) );
  AND U14881 ( .A(n438), .B(n11284), .Z(n11282) );
  XOR U14882 ( .A(n11285), .B(n11286), .Z(n11284) );
  XOR U14883 ( .A(DB[2190]), .B(DB[2175]), .Z(n11286) );
  AND U14884 ( .A(n442), .B(n11287), .Z(n11285) );
  XOR U14885 ( .A(n11288), .B(n11289), .Z(n11287) );
  XOR U14886 ( .A(DB[2175]), .B(DB[2160]), .Z(n11289) );
  AND U14887 ( .A(n446), .B(n11290), .Z(n11288) );
  XOR U14888 ( .A(n11291), .B(n11292), .Z(n11290) );
  XOR U14889 ( .A(DB[2160]), .B(DB[2145]), .Z(n11292) );
  AND U14890 ( .A(n450), .B(n11293), .Z(n11291) );
  XOR U14891 ( .A(n11294), .B(n11295), .Z(n11293) );
  XOR U14892 ( .A(DB[2145]), .B(DB[2130]), .Z(n11295) );
  AND U14893 ( .A(n454), .B(n11296), .Z(n11294) );
  XOR U14894 ( .A(n11297), .B(n11298), .Z(n11296) );
  XOR U14895 ( .A(DB[2130]), .B(DB[2115]), .Z(n11298) );
  AND U14896 ( .A(n458), .B(n11299), .Z(n11297) );
  XOR U14897 ( .A(n11300), .B(n11301), .Z(n11299) );
  XOR U14898 ( .A(DB[2115]), .B(DB[2100]), .Z(n11301) );
  AND U14899 ( .A(n462), .B(n11302), .Z(n11300) );
  XOR U14900 ( .A(n11303), .B(n11304), .Z(n11302) );
  XOR U14901 ( .A(DB[2100]), .B(DB[2085]), .Z(n11304) );
  AND U14902 ( .A(n466), .B(n11305), .Z(n11303) );
  XOR U14903 ( .A(n11306), .B(n11307), .Z(n11305) );
  XOR U14904 ( .A(DB[2085]), .B(DB[2070]), .Z(n11307) );
  AND U14905 ( .A(n470), .B(n11308), .Z(n11306) );
  XOR U14906 ( .A(n11309), .B(n11310), .Z(n11308) );
  XOR U14907 ( .A(DB[2070]), .B(DB[2055]), .Z(n11310) );
  AND U14908 ( .A(n474), .B(n11311), .Z(n11309) );
  XOR U14909 ( .A(n11312), .B(n11313), .Z(n11311) );
  XOR U14910 ( .A(DB[2055]), .B(DB[2040]), .Z(n11313) );
  AND U14911 ( .A(n478), .B(n11314), .Z(n11312) );
  XOR U14912 ( .A(n11315), .B(n11316), .Z(n11314) );
  XOR U14913 ( .A(DB[2040]), .B(DB[2025]), .Z(n11316) );
  AND U14914 ( .A(n482), .B(n11317), .Z(n11315) );
  XOR U14915 ( .A(n11318), .B(n11319), .Z(n11317) );
  XOR U14916 ( .A(DB[2025]), .B(DB[2010]), .Z(n11319) );
  AND U14917 ( .A(n486), .B(n11320), .Z(n11318) );
  XOR U14918 ( .A(n11321), .B(n11322), .Z(n11320) );
  XOR U14919 ( .A(DB[2010]), .B(DB[1995]), .Z(n11322) );
  AND U14920 ( .A(n490), .B(n11323), .Z(n11321) );
  XOR U14921 ( .A(n11324), .B(n11325), .Z(n11323) );
  XOR U14922 ( .A(DB[1995]), .B(DB[1980]), .Z(n11325) );
  AND U14923 ( .A(n494), .B(n11326), .Z(n11324) );
  XOR U14924 ( .A(n11327), .B(n11328), .Z(n11326) );
  XOR U14925 ( .A(DB[1980]), .B(DB[1965]), .Z(n11328) );
  AND U14926 ( .A(n498), .B(n11329), .Z(n11327) );
  XOR U14927 ( .A(n11330), .B(n11331), .Z(n11329) );
  XOR U14928 ( .A(DB[1965]), .B(DB[1950]), .Z(n11331) );
  AND U14929 ( .A(n502), .B(n11332), .Z(n11330) );
  XOR U14930 ( .A(n11333), .B(n11334), .Z(n11332) );
  XOR U14931 ( .A(DB[1950]), .B(DB[1935]), .Z(n11334) );
  AND U14932 ( .A(n506), .B(n11335), .Z(n11333) );
  XOR U14933 ( .A(n11336), .B(n11337), .Z(n11335) );
  XOR U14934 ( .A(DB[1935]), .B(DB[1920]), .Z(n11337) );
  AND U14935 ( .A(n510), .B(n11338), .Z(n11336) );
  XOR U14936 ( .A(n11339), .B(n11340), .Z(n11338) );
  XOR U14937 ( .A(DB[1920]), .B(DB[1905]), .Z(n11340) );
  AND U14938 ( .A(n514), .B(n11341), .Z(n11339) );
  XOR U14939 ( .A(n11342), .B(n11343), .Z(n11341) );
  XOR U14940 ( .A(DB[1905]), .B(DB[1890]), .Z(n11343) );
  AND U14941 ( .A(n518), .B(n11344), .Z(n11342) );
  XOR U14942 ( .A(n11345), .B(n11346), .Z(n11344) );
  XOR U14943 ( .A(DB[1890]), .B(DB[1875]), .Z(n11346) );
  AND U14944 ( .A(n522), .B(n11347), .Z(n11345) );
  XOR U14945 ( .A(n11348), .B(n11349), .Z(n11347) );
  XOR U14946 ( .A(DB[1875]), .B(DB[1860]), .Z(n11349) );
  AND U14947 ( .A(n526), .B(n11350), .Z(n11348) );
  XOR U14948 ( .A(n11351), .B(n11352), .Z(n11350) );
  XOR U14949 ( .A(DB[1860]), .B(DB[1845]), .Z(n11352) );
  AND U14950 ( .A(n530), .B(n11353), .Z(n11351) );
  XOR U14951 ( .A(n11354), .B(n11355), .Z(n11353) );
  XOR U14952 ( .A(DB[1845]), .B(DB[1830]), .Z(n11355) );
  AND U14953 ( .A(n534), .B(n11356), .Z(n11354) );
  XOR U14954 ( .A(n11357), .B(n11358), .Z(n11356) );
  XOR U14955 ( .A(DB[1830]), .B(DB[1815]), .Z(n11358) );
  AND U14956 ( .A(n538), .B(n11359), .Z(n11357) );
  XOR U14957 ( .A(n11360), .B(n11361), .Z(n11359) );
  XOR U14958 ( .A(DB[1815]), .B(DB[1800]), .Z(n11361) );
  AND U14959 ( .A(n542), .B(n11362), .Z(n11360) );
  XOR U14960 ( .A(n11363), .B(n11364), .Z(n11362) );
  XOR U14961 ( .A(DB[1800]), .B(DB[1785]), .Z(n11364) );
  AND U14962 ( .A(n546), .B(n11365), .Z(n11363) );
  XOR U14963 ( .A(n11366), .B(n11367), .Z(n11365) );
  XOR U14964 ( .A(DB[1785]), .B(DB[1770]), .Z(n11367) );
  AND U14965 ( .A(n550), .B(n11368), .Z(n11366) );
  XOR U14966 ( .A(n11369), .B(n11370), .Z(n11368) );
  XOR U14967 ( .A(DB[1770]), .B(DB[1755]), .Z(n11370) );
  AND U14968 ( .A(n554), .B(n11371), .Z(n11369) );
  XOR U14969 ( .A(n11372), .B(n11373), .Z(n11371) );
  XOR U14970 ( .A(DB[1755]), .B(DB[1740]), .Z(n11373) );
  AND U14971 ( .A(n558), .B(n11374), .Z(n11372) );
  XOR U14972 ( .A(n11375), .B(n11376), .Z(n11374) );
  XOR U14973 ( .A(DB[1740]), .B(DB[1725]), .Z(n11376) );
  AND U14974 ( .A(n562), .B(n11377), .Z(n11375) );
  XOR U14975 ( .A(n11378), .B(n11379), .Z(n11377) );
  XOR U14976 ( .A(DB[1725]), .B(DB[1710]), .Z(n11379) );
  AND U14977 ( .A(n566), .B(n11380), .Z(n11378) );
  XOR U14978 ( .A(n11381), .B(n11382), .Z(n11380) );
  XOR U14979 ( .A(DB[1710]), .B(DB[1695]), .Z(n11382) );
  AND U14980 ( .A(n570), .B(n11383), .Z(n11381) );
  XOR U14981 ( .A(n11384), .B(n11385), .Z(n11383) );
  XOR U14982 ( .A(DB[1695]), .B(DB[1680]), .Z(n11385) );
  AND U14983 ( .A(n574), .B(n11386), .Z(n11384) );
  XOR U14984 ( .A(n11387), .B(n11388), .Z(n11386) );
  XOR U14985 ( .A(DB[1680]), .B(DB[1665]), .Z(n11388) );
  AND U14986 ( .A(n578), .B(n11389), .Z(n11387) );
  XOR U14987 ( .A(n11390), .B(n11391), .Z(n11389) );
  XOR U14988 ( .A(DB[1665]), .B(DB[1650]), .Z(n11391) );
  AND U14989 ( .A(n582), .B(n11392), .Z(n11390) );
  XOR U14990 ( .A(n11393), .B(n11394), .Z(n11392) );
  XOR U14991 ( .A(DB[1650]), .B(DB[1635]), .Z(n11394) );
  AND U14992 ( .A(n586), .B(n11395), .Z(n11393) );
  XOR U14993 ( .A(n11396), .B(n11397), .Z(n11395) );
  XOR U14994 ( .A(DB[1635]), .B(DB[1620]), .Z(n11397) );
  AND U14995 ( .A(n590), .B(n11398), .Z(n11396) );
  XOR U14996 ( .A(n11399), .B(n11400), .Z(n11398) );
  XOR U14997 ( .A(DB[1620]), .B(DB[1605]), .Z(n11400) );
  AND U14998 ( .A(n594), .B(n11401), .Z(n11399) );
  XOR U14999 ( .A(n11402), .B(n11403), .Z(n11401) );
  XOR U15000 ( .A(DB[1605]), .B(DB[1590]), .Z(n11403) );
  AND U15001 ( .A(n598), .B(n11404), .Z(n11402) );
  XOR U15002 ( .A(n11405), .B(n11406), .Z(n11404) );
  XOR U15003 ( .A(DB[1590]), .B(DB[1575]), .Z(n11406) );
  AND U15004 ( .A(n602), .B(n11407), .Z(n11405) );
  XOR U15005 ( .A(n11408), .B(n11409), .Z(n11407) );
  XOR U15006 ( .A(DB[1575]), .B(DB[1560]), .Z(n11409) );
  AND U15007 ( .A(n606), .B(n11410), .Z(n11408) );
  XOR U15008 ( .A(n11411), .B(n11412), .Z(n11410) );
  XOR U15009 ( .A(DB[1560]), .B(DB[1545]), .Z(n11412) );
  AND U15010 ( .A(n610), .B(n11413), .Z(n11411) );
  XOR U15011 ( .A(n11414), .B(n11415), .Z(n11413) );
  XOR U15012 ( .A(DB[1545]), .B(DB[1530]), .Z(n11415) );
  AND U15013 ( .A(n614), .B(n11416), .Z(n11414) );
  XOR U15014 ( .A(n11417), .B(n11418), .Z(n11416) );
  XOR U15015 ( .A(DB[1530]), .B(DB[1515]), .Z(n11418) );
  AND U15016 ( .A(n618), .B(n11419), .Z(n11417) );
  XOR U15017 ( .A(n11420), .B(n11421), .Z(n11419) );
  XOR U15018 ( .A(DB[1515]), .B(DB[1500]), .Z(n11421) );
  AND U15019 ( .A(n622), .B(n11422), .Z(n11420) );
  XOR U15020 ( .A(n11423), .B(n11424), .Z(n11422) );
  XOR U15021 ( .A(DB[1500]), .B(DB[1485]), .Z(n11424) );
  AND U15022 ( .A(n626), .B(n11425), .Z(n11423) );
  XOR U15023 ( .A(n11426), .B(n11427), .Z(n11425) );
  XOR U15024 ( .A(DB[1485]), .B(DB[1470]), .Z(n11427) );
  AND U15025 ( .A(n630), .B(n11428), .Z(n11426) );
  XOR U15026 ( .A(n11429), .B(n11430), .Z(n11428) );
  XOR U15027 ( .A(DB[1470]), .B(DB[1455]), .Z(n11430) );
  AND U15028 ( .A(n634), .B(n11431), .Z(n11429) );
  XOR U15029 ( .A(n11432), .B(n11433), .Z(n11431) );
  XOR U15030 ( .A(DB[1455]), .B(DB[1440]), .Z(n11433) );
  AND U15031 ( .A(n638), .B(n11434), .Z(n11432) );
  XOR U15032 ( .A(n11435), .B(n11436), .Z(n11434) );
  XOR U15033 ( .A(DB[1440]), .B(DB[1425]), .Z(n11436) );
  AND U15034 ( .A(n642), .B(n11437), .Z(n11435) );
  XOR U15035 ( .A(n11438), .B(n11439), .Z(n11437) );
  XOR U15036 ( .A(DB[1425]), .B(DB[1410]), .Z(n11439) );
  AND U15037 ( .A(n646), .B(n11440), .Z(n11438) );
  XOR U15038 ( .A(n11441), .B(n11442), .Z(n11440) );
  XOR U15039 ( .A(DB[1410]), .B(DB[1395]), .Z(n11442) );
  AND U15040 ( .A(n650), .B(n11443), .Z(n11441) );
  XOR U15041 ( .A(n11444), .B(n11445), .Z(n11443) );
  XOR U15042 ( .A(DB[1395]), .B(DB[1380]), .Z(n11445) );
  AND U15043 ( .A(n654), .B(n11446), .Z(n11444) );
  XOR U15044 ( .A(n11447), .B(n11448), .Z(n11446) );
  XOR U15045 ( .A(DB[1380]), .B(DB[1365]), .Z(n11448) );
  AND U15046 ( .A(n658), .B(n11449), .Z(n11447) );
  XOR U15047 ( .A(n11450), .B(n11451), .Z(n11449) );
  XOR U15048 ( .A(DB[1365]), .B(DB[1350]), .Z(n11451) );
  AND U15049 ( .A(n662), .B(n11452), .Z(n11450) );
  XOR U15050 ( .A(n11453), .B(n11454), .Z(n11452) );
  XOR U15051 ( .A(DB[1350]), .B(DB[1335]), .Z(n11454) );
  AND U15052 ( .A(n666), .B(n11455), .Z(n11453) );
  XOR U15053 ( .A(n11456), .B(n11457), .Z(n11455) );
  XOR U15054 ( .A(DB[1335]), .B(DB[1320]), .Z(n11457) );
  AND U15055 ( .A(n670), .B(n11458), .Z(n11456) );
  XOR U15056 ( .A(n11459), .B(n11460), .Z(n11458) );
  XOR U15057 ( .A(DB[1320]), .B(DB[1305]), .Z(n11460) );
  AND U15058 ( .A(n674), .B(n11461), .Z(n11459) );
  XOR U15059 ( .A(n11462), .B(n11463), .Z(n11461) );
  XOR U15060 ( .A(DB[1305]), .B(DB[1290]), .Z(n11463) );
  AND U15061 ( .A(n678), .B(n11464), .Z(n11462) );
  XOR U15062 ( .A(n11465), .B(n11466), .Z(n11464) );
  XOR U15063 ( .A(DB[1290]), .B(DB[1275]), .Z(n11466) );
  AND U15064 ( .A(n682), .B(n11467), .Z(n11465) );
  XOR U15065 ( .A(n11468), .B(n11469), .Z(n11467) );
  XOR U15066 ( .A(DB[1275]), .B(DB[1260]), .Z(n11469) );
  AND U15067 ( .A(n686), .B(n11470), .Z(n11468) );
  XOR U15068 ( .A(n11471), .B(n11472), .Z(n11470) );
  XOR U15069 ( .A(DB[1260]), .B(DB[1245]), .Z(n11472) );
  AND U15070 ( .A(n690), .B(n11473), .Z(n11471) );
  XOR U15071 ( .A(n11474), .B(n11475), .Z(n11473) );
  XOR U15072 ( .A(DB[1245]), .B(DB[1230]), .Z(n11475) );
  AND U15073 ( .A(n694), .B(n11476), .Z(n11474) );
  XOR U15074 ( .A(n11477), .B(n11478), .Z(n11476) );
  XOR U15075 ( .A(DB[1230]), .B(DB[1215]), .Z(n11478) );
  AND U15076 ( .A(n698), .B(n11479), .Z(n11477) );
  XOR U15077 ( .A(n11480), .B(n11481), .Z(n11479) );
  XOR U15078 ( .A(DB[1215]), .B(DB[1200]), .Z(n11481) );
  AND U15079 ( .A(n702), .B(n11482), .Z(n11480) );
  XOR U15080 ( .A(n11483), .B(n11484), .Z(n11482) );
  XOR U15081 ( .A(DB[1200]), .B(DB[1185]), .Z(n11484) );
  AND U15082 ( .A(n706), .B(n11485), .Z(n11483) );
  XOR U15083 ( .A(n11486), .B(n11487), .Z(n11485) );
  XOR U15084 ( .A(DB[1185]), .B(DB[1170]), .Z(n11487) );
  AND U15085 ( .A(n710), .B(n11488), .Z(n11486) );
  XOR U15086 ( .A(n11489), .B(n11490), .Z(n11488) );
  XOR U15087 ( .A(DB[1170]), .B(DB[1155]), .Z(n11490) );
  AND U15088 ( .A(n714), .B(n11491), .Z(n11489) );
  XOR U15089 ( .A(n11492), .B(n11493), .Z(n11491) );
  XOR U15090 ( .A(DB[1155]), .B(DB[1140]), .Z(n11493) );
  AND U15091 ( .A(n718), .B(n11494), .Z(n11492) );
  XOR U15092 ( .A(n11495), .B(n11496), .Z(n11494) );
  XOR U15093 ( .A(DB[1140]), .B(DB[1125]), .Z(n11496) );
  AND U15094 ( .A(n722), .B(n11497), .Z(n11495) );
  XOR U15095 ( .A(n11498), .B(n11499), .Z(n11497) );
  XOR U15096 ( .A(DB[1125]), .B(DB[1110]), .Z(n11499) );
  AND U15097 ( .A(n726), .B(n11500), .Z(n11498) );
  XOR U15098 ( .A(n11501), .B(n11502), .Z(n11500) );
  XOR U15099 ( .A(DB[1110]), .B(DB[1095]), .Z(n11502) );
  AND U15100 ( .A(n730), .B(n11503), .Z(n11501) );
  XOR U15101 ( .A(n11504), .B(n11505), .Z(n11503) );
  XOR U15102 ( .A(DB[1095]), .B(DB[1080]), .Z(n11505) );
  AND U15103 ( .A(n734), .B(n11506), .Z(n11504) );
  XOR U15104 ( .A(n11507), .B(n11508), .Z(n11506) );
  XOR U15105 ( .A(DB[1080]), .B(DB[1065]), .Z(n11508) );
  AND U15106 ( .A(n738), .B(n11509), .Z(n11507) );
  XOR U15107 ( .A(n11510), .B(n11511), .Z(n11509) );
  XOR U15108 ( .A(DB[1065]), .B(DB[1050]), .Z(n11511) );
  AND U15109 ( .A(n742), .B(n11512), .Z(n11510) );
  XOR U15110 ( .A(n11513), .B(n11514), .Z(n11512) );
  XOR U15111 ( .A(DB[1050]), .B(DB[1035]), .Z(n11514) );
  AND U15112 ( .A(n746), .B(n11515), .Z(n11513) );
  XOR U15113 ( .A(n11516), .B(n11517), .Z(n11515) );
  XOR U15114 ( .A(DB[1035]), .B(DB[1020]), .Z(n11517) );
  AND U15115 ( .A(n750), .B(n11518), .Z(n11516) );
  XOR U15116 ( .A(n11519), .B(n11520), .Z(n11518) );
  XOR U15117 ( .A(DB[1020]), .B(DB[1005]), .Z(n11520) );
  AND U15118 ( .A(n754), .B(n11521), .Z(n11519) );
  XOR U15119 ( .A(n11522), .B(n11523), .Z(n11521) );
  XOR U15120 ( .A(DB[990]), .B(DB[1005]), .Z(n11523) );
  AND U15121 ( .A(n758), .B(n11524), .Z(n11522) );
  XOR U15122 ( .A(n11525), .B(n11526), .Z(n11524) );
  XOR U15123 ( .A(DB[990]), .B(DB[975]), .Z(n11526) );
  AND U15124 ( .A(n762), .B(n11527), .Z(n11525) );
  XOR U15125 ( .A(n11528), .B(n11529), .Z(n11527) );
  XOR U15126 ( .A(DB[975]), .B(DB[960]), .Z(n11529) );
  AND U15127 ( .A(n766), .B(n11530), .Z(n11528) );
  XOR U15128 ( .A(n11531), .B(n11532), .Z(n11530) );
  XOR U15129 ( .A(DB[960]), .B(DB[945]), .Z(n11532) );
  AND U15130 ( .A(n770), .B(n11533), .Z(n11531) );
  XOR U15131 ( .A(n11534), .B(n11535), .Z(n11533) );
  XOR U15132 ( .A(DB[945]), .B(DB[930]), .Z(n11535) );
  AND U15133 ( .A(n774), .B(n11536), .Z(n11534) );
  XOR U15134 ( .A(n11537), .B(n11538), .Z(n11536) );
  XOR U15135 ( .A(DB[930]), .B(DB[915]), .Z(n11538) );
  AND U15136 ( .A(n778), .B(n11539), .Z(n11537) );
  XOR U15137 ( .A(n11540), .B(n11541), .Z(n11539) );
  XOR U15138 ( .A(DB[915]), .B(DB[900]), .Z(n11541) );
  AND U15139 ( .A(n782), .B(n11542), .Z(n11540) );
  XOR U15140 ( .A(n11543), .B(n11544), .Z(n11542) );
  XOR U15141 ( .A(DB[900]), .B(DB[885]), .Z(n11544) );
  AND U15142 ( .A(n786), .B(n11545), .Z(n11543) );
  XOR U15143 ( .A(n11546), .B(n11547), .Z(n11545) );
  XOR U15144 ( .A(DB[885]), .B(DB[870]), .Z(n11547) );
  AND U15145 ( .A(n790), .B(n11548), .Z(n11546) );
  XOR U15146 ( .A(n11549), .B(n11550), .Z(n11548) );
  XOR U15147 ( .A(DB[870]), .B(DB[855]), .Z(n11550) );
  AND U15148 ( .A(n794), .B(n11551), .Z(n11549) );
  XOR U15149 ( .A(n11552), .B(n11553), .Z(n11551) );
  XOR U15150 ( .A(DB[855]), .B(DB[840]), .Z(n11553) );
  AND U15151 ( .A(n798), .B(n11554), .Z(n11552) );
  XOR U15152 ( .A(n11555), .B(n11556), .Z(n11554) );
  XOR U15153 ( .A(DB[840]), .B(DB[825]), .Z(n11556) );
  AND U15154 ( .A(n802), .B(n11557), .Z(n11555) );
  XOR U15155 ( .A(n11558), .B(n11559), .Z(n11557) );
  XOR U15156 ( .A(DB[825]), .B(DB[810]), .Z(n11559) );
  AND U15157 ( .A(n806), .B(n11560), .Z(n11558) );
  XOR U15158 ( .A(n11561), .B(n11562), .Z(n11560) );
  XOR U15159 ( .A(DB[810]), .B(DB[795]), .Z(n11562) );
  AND U15160 ( .A(n810), .B(n11563), .Z(n11561) );
  XOR U15161 ( .A(n11564), .B(n11565), .Z(n11563) );
  XOR U15162 ( .A(DB[795]), .B(DB[780]), .Z(n11565) );
  AND U15163 ( .A(n814), .B(n11566), .Z(n11564) );
  XOR U15164 ( .A(n11567), .B(n11568), .Z(n11566) );
  XOR U15165 ( .A(DB[780]), .B(DB[765]), .Z(n11568) );
  AND U15166 ( .A(n818), .B(n11569), .Z(n11567) );
  XOR U15167 ( .A(n11570), .B(n11571), .Z(n11569) );
  XOR U15168 ( .A(DB[765]), .B(DB[750]), .Z(n11571) );
  AND U15169 ( .A(n822), .B(n11572), .Z(n11570) );
  XOR U15170 ( .A(n11573), .B(n11574), .Z(n11572) );
  XOR U15171 ( .A(DB[750]), .B(DB[735]), .Z(n11574) );
  AND U15172 ( .A(n826), .B(n11575), .Z(n11573) );
  XOR U15173 ( .A(n11576), .B(n11577), .Z(n11575) );
  XOR U15174 ( .A(DB[735]), .B(DB[720]), .Z(n11577) );
  AND U15175 ( .A(n830), .B(n11578), .Z(n11576) );
  XOR U15176 ( .A(n11579), .B(n11580), .Z(n11578) );
  XOR U15177 ( .A(DB[720]), .B(DB[705]), .Z(n11580) );
  AND U15178 ( .A(n834), .B(n11581), .Z(n11579) );
  XOR U15179 ( .A(n11582), .B(n11583), .Z(n11581) );
  XOR U15180 ( .A(DB[705]), .B(DB[690]), .Z(n11583) );
  AND U15181 ( .A(n838), .B(n11584), .Z(n11582) );
  XOR U15182 ( .A(n11585), .B(n11586), .Z(n11584) );
  XOR U15183 ( .A(DB[690]), .B(DB[675]), .Z(n11586) );
  AND U15184 ( .A(n842), .B(n11587), .Z(n11585) );
  XOR U15185 ( .A(n11588), .B(n11589), .Z(n11587) );
  XOR U15186 ( .A(DB[675]), .B(DB[660]), .Z(n11589) );
  AND U15187 ( .A(n846), .B(n11590), .Z(n11588) );
  XOR U15188 ( .A(n11591), .B(n11592), .Z(n11590) );
  XOR U15189 ( .A(DB[660]), .B(DB[645]), .Z(n11592) );
  AND U15190 ( .A(n850), .B(n11593), .Z(n11591) );
  XOR U15191 ( .A(n11594), .B(n11595), .Z(n11593) );
  XOR U15192 ( .A(DB[645]), .B(DB[630]), .Z(n11595) );
  AND U15193 ( .A(n854), .B(n11596), .Z(n11594) );
  XOR U15194 ( .A(n11597), .B(n11598), .Z(n11596) );
  XOR U15195 ( .A(DB[630]), .B(DB[615]), .Z(n11598) );
  AND U15196 ( .A(n858), .B(n11599), .Z(n11597) );
  XOR U15197 ( .A(n11600), .B(n11601), .Z(n11599) );
  XOR U15198 ( .A(DB[615]), .B(DB[600]), .Z(n11601) );
  AND U15199 ( .A(n862), .B(n11602), .Z(n11600) );
  XOR U15200 ( .A(n11603), .B(n11604), .Z(n11602) );
  XOR U15201 ( .A(DB[600]), .B(DB[585]), .Z(n11604) );
  AND U15202 ( .A(n866), .B(n11605), .Z(n11603) );
  XOR U15203 ( .A(n11606), .B(n11607), .Z(n11605) );
  XOR U15204 ( .A(DB[585]), .B(DB[570]), .Z(n11607) );
  AND U15205 ( .A(n870), .B(n11608), .Z(n11606) );
  XOR U15206 ( .A(n11609), .B(n11610), .Z(n11608) );
  XOR U15207 ( .A(DB[570]), .B(DB[555]), .Z(n11610) );
  AND U15208 ( .A(n874), .B(n11611), .Z(n11609) );
  XOR U15209 ( .A(n11612), .B(n11613), .Z(n11611) );
  XOR U15210 ( .A(DB[555]), .B(DB[540]), .Z(n11613) );
  AND U15211 ( .A(n878), .B(n11614), .Z(n11612) );
  XOR U15212 ( .A(n11615), .B(n11616), .Z(n11614) );
  XOR U15213 ( .A(DB[540]), .B(DB[525]), .Z(n11616) );
  AND U15214 ( .A(n882), .B(n11617), .Z(n11615) );
  XOR U15215 ( .A(n11618), .B(n11619), .Z(n11617) );
  XOR U15216 ( .A(DB[525]), .B(DB[510]), .Z(n11619) );
  AND U15217 ( .A(n886), .B(n11620), .Z(n11618) );
  XOR U15218 ( .A(n11621), .B(n11622), .Z(n11620) );
  XOR U15219 ( .A(DB[510]), .B(DB[495]), .Z(n11622) );
  AND U15220 ( .A(n890), .B(n11623), .Z(n11621) );
  XOR U15221 ( .A(n11624), .B(n11625), .Z(n11623) );
  XOR U15222 ( .A(DB[495]), .B(DB[480]), .Z(n11625) );
  AND U15223 ( .A(n894), .B(n11626), .Z(n11624) );
  XOR U15224 ( .A(n11627), .B(n11628), .Z(n11626) );
  XOR U15225 ( .A(DB[480]), .B(DB[465]), .Z(n11628) );
  AND U15226 ( .A(n898), .B(n11629), .Z(n11627) );
  XOR U15227 ( .A(n11630), .B(n11631), .Z(n11629) );
  XOR U15228 ( .A(DB[465]), .B(DB[450]), .Z(n11631) );
  AND U15229 ( .A(n902), .B(n11632), .Z(n11630) );
  XOR U15230 ( .A(n11633), .B(n11634), .Z(n11632) );
  XOR U15231 ( .A(DB[450]), .B(DB[435]), .Z(n11634) );
  AND U15232 ( .A(n906), .B(n11635), .Z(n11633) );
  XOR U15233 ( .A(n11636), .B(n11637), .Z(n11635) );
  XOR U15234 ( .A(DB[435]), .B(DB[420]), .Z(n11637) );
  AND U15235 ( .A(n910), .B(n11638), .Z(n11636) );
  XOR U15236 ( .A(n11639), .B(n11640), .Z(n11638) );
  XOR U15237 ( .A(DB[420]), .B(DB[405]), .Z(n11640) );
  AND U15238 ( .A(n914), .B(n11641), .Z(n11639) );
  XOR U15239 ( .A(n11642), .B(n11643), .Z(n11641) );
  XOR U15240 ( .A(DB[405]), .B(DB[390]), .Z(n11643) );
  AND U15241 ( .A(n918), .B(n11644), .Z(n11642) );
  XOR U15242 ( .A(n11645), .B(n11646), .Z(n11644) );
  XOR U15243 ( .A(DB[390]), .B(DB[375]), .Z(n11646) );
  AND U15244 ( .A(n922), .B(n11647), .Z(n11645) );
  XOR U15245 ( .A(n11648), .B(n11649), .Z(n11647) );
  XOR U15246 ( .A(DB[375]), .B(DB[360]), .Z(n11649) );
  AND U15247 ( .A(n926), .B(n11650), .Z(n11648) );
  XOR U15248 ( .A(n11651), .B(n11652), .Z(n11650) );
  XOR U15249 ( .A(DB[360]), .B(DB[345]), .Z(n11652) );
  AND U15250 ( .A(n930), .B(n11653), .Z(n11651) );
  XOR U15251 ( .A(n11654), .B(n11655), .Z(n11653) );
  XOR U15252 ( .A(DB[345]), .B(DB[330]), .Z(n11655) );
  AND U15253 ( .A(n934), .B(n11656), .Z(n11654) );
  XOR U15254 ( .A(n11657), .B(n11658), .Z(n11656) );
  XOR U15255 ( .A(DB[330]), .B(DB[315]), .Z(n11658) );
  AND U15256 ( .A(n938), .B(n11659), .Z(n11657) );
  XOR U15257 ( .A(n11660), .B(n11661), .Z(n11659) );
  XOR U15258 ( .A(DB[315]), .B(DB[300]), .Z(n11661) );
  AND U15259 ( .A(n942), .B(n11662), .Z(n11660) );
  XOR U15260 ( .A(n11663), .B(n11664), .Z(n11662) );
  XOR U15261 ( .A(DB[300]), .B(DB[285]), .Z(n11664) );
  AND U15262 ( .A(n946), .B(n11665), .Z(n11663) );
  XOR U15263 ( .A(n11666), .B(n11667), .Z(n11665) );
  XOR U15264 ( .A(DB[285]), .B(DB[270]), .Z(n11667) );
  AND U15265 ( .A(n950), .B(n11668), .Z(n11666) );
  XOR U15266 ( .A(n11669), .B(n11670), .Z(n11668) );
  XOR U15267 ( .A(DB[270]), .B(DB[255]), .Z(n11670) );
  AND U15268 ( .A(n954), .B(n11671), .Z(n11669) );
  XOR U15269 ( .A(n11672), .B(n11673), .Z(n11671) );
  XOR U15270 ( .A(DB[255]), .B(DB[240]), .Z(n11673) );
  AND U15271 ( .A(n958), .B(n11674), .Z(n11672) );
  XOR U15272 ( .A(n11675), .B(n11676), .Z(n11674) );
  XOR U15273 ( .A(DB[240]), .B(DB[225]), .Z(n11676) );
  AND U15274 ( .A(n962), .B(n11677), .Z(n11675) );
  XOR U15275 ( .A(n11678), .B(n11679), .Z(n11677) );
  XOR U15276 ( .A(DB[225]), .B(DB[210]), .Z(n11679) );
  AND U15277 ( .A(n966), .B(n11680), .Z(n11678) );
  XOR U15278 ( .A(n11681), .B(n11682), .Z(n11680) );
  XOR U15279 ( .A(DB[210]), .B(DB[195]), .Z(n11682) );
  AND U15280 ( .A(n970), .B(n11683), .Z(n11681) );
  XOR U15281 ( .A(n11684), .B(n11685), .Z(n11683) );
  XOR U15282 ( .A(DB[195]), .B(DB[180]), .Z(n11685) );
  AND U15283 ( .A(n974), .B(n11686), .Z(n11684) );
  XOR U15284 ( .A(n11687), .B(n11688), .Z(n11686) );
  XOR U15285 ( .A(DB[180]), .B(DB[165]), .Z(n11688) );
  AND U15286 ( .A(n978), .B(n11689), .Z(n11687) );
  XOR U15287 ( .A(n11690), .B(n11691), .Z(n11689) );
  XOR U15288 ( .A(DB[165]), .B(DB[150]), .Z(n11691) );
  AND U15289 ( .A(n982), .B(n11692), .Z(n11690) );
  XOR U15290 ( .A(n11693), .B(n11694), .Z(n11692) );
  XOR U15291 ( .A(DB[150]), .B(DB[135]), .Z(n11694) );
  AND U15292 ( .A(n986), .B(n11695), .Z(n11693) );
  XOR U15293 ( .A(n11696), .B(n11697), .Z(n11695) );
  XOR U15294 ( .A(DB[135]), .B(DB[120]), .Z(n11697) );
  AND U15295 ( .A(n990), .B(n11698), .Z(n11696) );
  XOR U15296 ( .A(n11699), .B(n11700), .Z(n11698) );
  XOR U15297 ( .A(DB[120]), .B(DB[105]), .Z(n11700) );
  AND U15298 ( .A(n994), .B(n11701), .Z(n11699) );
  XOR U15299 ( .A(n11702), .B(n11703), .Z(n11701) );
  XOR U15300 ( .A(DB[90]), .B(DB[105]), .Z(n11703) );
  AND U15301 ( .A(n998), .B(n11704), .Z(n11702) );
  XOR U15302 ( .A(n11705), .B(n11706), .Z(n11704) );
  XOR U15303 ( .A(DB[90]), .B(DB[75]), .Z(n11706) );
  AND U15304 ( .A(n1002), .B(n11707), .Z(n11705) );
  XOR U15305 ( .A(n11708), .B(n11709), .Z(n11707) );
  XOR U15306 ( .A(DB[75]), .B(DB[60]), .Z(n11709) );
  AND U15307 ( .A(n1006), .B(n11710), .Z(n11708) );
  XOR U15308 ( .A(n11711), .B(n11712), .Z(n11710) );
  XOR U15309 ( .A(DB[60]), .B(DB[45]), .Z(n11712) );
  AND U15310 ( .A(n1010), .B(n11713), .Z(n11711) );
  XOR U15311 ( .A(n11714), .B(n11715), .Z(n11713) );
  XOR U15312 ( .A(DB[45]), .B(DB[30]), .Z(n11715) );
  AND U15313 ( .A(n1014), .B(n11716), .Z(n11714) );
  XOR U15314 ( .A(n11717), .B(n11718), .Z(n11716) );
  XOR U15315 ( .A(DB[30]), .B(DB[15]), .Z(n11718) );
  AND U15316 ( .A(n1018), .B(n11719), .Z(n11717) );
  XOR U15317 ( .A(DB[15]), .B(DB[0]), .Z(n11719) );
  XNOR U15318 ( .A(n11720), .B(n11721), .Z(n2) );
  AND U15319 ( .A(n11722), .B(n11723), .Z(n11720) );
  XOR U15320 ( .A(n11721), .B(n11724), .Z(n11723) );
  XOR U15321 ( .A(n11725), .B(n11726), .Z(n11724) );
  AND U15322 ( .A(n11727), .B(n11728), .Z(n11725) );
  XNOR U15323 ( .A(n11729), .B(n11730), .Z(n11728) );
  XOR U15324 ( .A(n11721), .B(n11731), .Z(n11722) );
  XNOR U15325 ( .A(n11732), .B(n11733), .Z(n11731) );
  AND U15326 ( .A(n6), .B(n11734), .Z(n11732) );
  XOR U15327 ( .A(n11735), .B(n11733), .Z(n11734) );
  XNOR U15328 ( .A(n11736), .B(n11737), .Z(n11721) );
  AND U15329 ( .A(n11738), .B(n11739), .Z(n11736) );
  XOR U15330 ( .A(n11727), .B(n11740), .Z(n11739) );
  XNOR U15331 ( .A(n11737), .B(n11729), .Z(n11740) );
  XNOR U15332 ( .A(n11741), .B(n11742), .Z(n11729) );
  ANDN U15333 ( .B(n11743), .A(n11744), .Z(n11741) );
  XOR U15334 ( .A(n11742), .B(n11745), .Z(n11743) );
  XNOR U15335 ( .A(n11726), .B(n11746), .Z(n11727) );
  XNOR U15336 ( .A(n11747), .B(n11748), .Z(n11746) );
  ANDN U15337 ( .B(n11749), .A(n11750), .Z(n11747) );
  XNOR U15338 ( .A(n11751), .B(n11752), .Z(n11749) );
  IV U15339 ( .A(n11730), .Z(n11726) );
  XOR U15340 ( .A(n11753), .B(n11754), .Z(n11730) );
  AND U15341 ( .A(n11755), .B(n11756), .Z(n11753) );
  XOR U15342 ( .A(n11757), .B(n11754), .Z(n11756) );
  XNOR U15343 ( .A(n11737), .B(n11758), .Z(n11738) );
  XOR U15344 ( .A(n11759), .B(n11760), .Z(n11758) );
  AND U15345 ( .A(n6), .B(n11761), .Z(n11759) );
  XNOR U15346 ( .A(n11762), .B(n11760), .Z(n11761) );
  XNOR U15347 ( .A(n11763), .B(n11764), .Z(n11737) );
  NAND U15348 ( .A(n11765), .B(n11766), .Z(n11764) );
  XOR U15349 ( .A(n11755), .B(n11767), .Z(n11766) );
  XOR U15350 ( .A(n11763), .B(n11757), .Z(n11767) );
  XOR U15351 ( .A(n11768), .B(n11745), .Z(n11757) );
  XNOR U15352 ( .A(n11769), .B(n11770), .Z(n11745) );
  ANDN U15353 ( .B(n11771), .A(n11772), .Z(n11769) );
  XNOR U15354 ( .A(n11770), .B(n11773), .Z(n11771) );
  IV U15355 ( .A(n11744), .Z(n11768) );
  XOR U15356 ( .A(n11774), .B(n11775), .Z(n11744) );
  XNOR U15357 ( .A(n11776), .B(n11777), .Z(n11775) );
  ANDN U15358 ( .B(n11778), .A(n11779), .Z(n11776) );
  XNOR U15359 ( .A(n11780), .B(n11781), .Z(n11778) );
  IV U15360 ( .A(n11777), .Z(n11781) );
  IV U15361 ( .A(n11742), .Z(n11774) );
  XNOR U15362 ( .A(n11782), .B(n11783), .Z(n11742) );
  ANDN U15363 ( .B(n11784), .A(n11785), .Z(n11782) );
  XNOR U15364 ( .A(n11783), .B(n11786), .Z(n11784) );
  XNOR U15365 ( .A(n11787), .B(n11788), .Z(n11755) );
  XNOR U15366 ( .A(n11751), .B(n11789), .Z(n11788) );
  IV U15367 ( .A(n11754), .Z(n11789) );
  XNOR U15368 ( .A(n11790), .B(n11791), .Z(n11754) );
  AND U15369 ( .A(n11792), .B(n11793), .Z(n11790) );
  XNOR U15370 ( .A(n11791), .B(n11794), .Z(n11793) );
  XOR U15371 ( .A(n11795), .B(n11796), .Z(n11751) );
  ANDN U15372 ( .B(n11797), .A(n11798), .Z(n11795) );
  XNOR U15373 ( .A(n11796), .B(n11799), .Z(n11797) );
  IV U15374 ( .A(n11750), .Z(n11787) );
  XOR U15375 ( .A(n11748), .B(n11800), .Z(n11750) );
  XNOR U15376 ( .A(n11801), .B(n11802), .Z(n11800) );
  ANDN U15377 ( .B(n11803), .A(n11804), .Z(n11801) );
  XNOR U15378 ( .A(n11805), .B(n11806), .Z(n11803) );
  IV U15379 ( .A(n11802), .Z(n11806) );
  IV U15380 ( .A(n11752), .Z(n11748) );
  XNOR U15381 ( .A(n11807), .B(n11808), .Z(n11752) );
  ANDN U15382 ( .B(n11809), .A(n11810), .Z(n11807) );
  XNOR U15383 ( .A(n11811), .B(n11808), .Z(n11809) );
  XOR U15384 ( .A(n11812), .B(n11813), .Z(n11765) );
  XNOR U15385 ( .A(n11763), .B(n11814), .Z(n11813) );
  NAND U15386 ( .A(n11815), .B(n6), .Z(n11814) );
  XOR U15387 ( .A(n11816), .B(n11812), .Z(n11815) );
  NAND U15388 ( .A(n11817), .B(n11818), .Z(n11763) );
  XNOR U15389 ( .A(n11792), .B(n11794), .Z(n11818) );
  XOR U15390 ( .A(n11819), .B(n11786), .Z(n11794) );
  XOR U15391 ( .A(n11820), .B(n11773), .Z(n11786) );
  XNOR U15392 ( .A(q[14]), .B(DB[3839]), .Z(n11773) );
  IV U15393 ( .A(n11772), .Z(n11820) );
  XOR U15394 ( .A(n11770), .B(n11821), .Z(n11772) );
  XNOR U15395 ( .A(q[13]), .B(DB[3838]), .Z(n11821) );
  XOR U15396 ( .A(q[12]), .B(DB[3837]), .Z(n11770) );
  IV U15397 ( .A(n11785), .Z(n11819) );
  XOR U15398 ( .A(n11822), .B(n11823), .Z(n11785) );
  XNOR U15399 ( .A(n11780), .B(n11783), .Z(n11823) );
  XOR U15400 ( .A(q[8]), .B(DB[3833]), .Z(n11783) );
  XOR U15401 ( .A(q[11]), .B(DB[3836]), .Z(n11780) );
  IV U15402 ( .A(n11779), .Z(n11822) );
  XOR U15403 ( .A(n11777), .B(n11824), .Z(n11779) );
  XNOR U15404 ( .A(q[10]), .B(DB[3835]), .Z(n11824) );
  XOR U15405 ( .A(q[9]), .B(DB[3834]), .Z(n11777) );
  XNOR U15406 ( .A(n11825), .B(n11826), .Z(n11792) );
  XOR U15407 ( .A(n11811), .B(n11791), .Z(n11826) );
  XOR U15408 ( .A(q[0]), .B(DB[3825]), .Z(n11791) );
  XOR U15409 ( .A(n11827), .B(n11799), .Z(n11811) );
  XNOR U15410 ( .A(q[7]), .B(DB[3832]), .Z(n11799) );
  IV U15411 ( .A(n11798), .Z(n11827) );
  XOR U15412 ( .A(n11796), .B(n11828), .Z(n11798) );
  XNOR U15413 ( .A(q[6]), .B(DB[3831]), .Z(n11828) );
  XOR U15414 ( .A(q[5]), .B(DB[3830]), .Z(n11796) );
  IV U15415 ( .A(n11810), .Z(n11825) );
  XOR U15416 ( .A(n11829), .B(n11830), .Z(n11810) );
  XNOR U15417 ( .A(n11805), .B(n11808), .Z(n11830) );
  XOR U15418 ( .A(q[1]), .B(DB[3826]), .Z(n11808) );
  XOR U15419 ( .A(q[4]), .B(DB[3829]), .Z(n11805) );
  IV U15420 ( .A(n11804), .Z(n11829) );
  XOR U15421 ( .A(n11802), .B(n11831), .Z(n11804) );
  XNOR U15422 ( .A(q[3]), .B(DB[3828]), .Z(n11831) );
  XOR U15423 ( .A(q[2]), .B(DB[3827]), .Z(n11802) );
  XOR U15424 ( .A(n11832), .B(n11833), .Z(n11817) );
  AND U15425 ( .A(n6), .B(n11834), .Z(n11832) );
  XOR U15426 ( .A(n11833), .B(n11835), .Z(n11834) );
  XNOR U15427 ( .A(n11836), .B(n11837), .Z(n6) );
  AND U15428 ( .A(n11838), .B(n11839), .Z(n11836) );
  XOR U15429 ( .A(n11837), .B(n11733), .Z(n11839) );
  XNOR U15430 ( .A(n11840), .B(n11841), .Z(n11733) );
  ANDN U15431 ( .B(n11842), .A(n11843), .Z(n11840) );
  XOR U15432 ( .A(n11841), .B(n11844), .Z(n11842) );
  XNOR U15433 ( .A(n11837), .B(n11735), .Z(n11838) );
  XOR U15434 ( .A(n11845), .B(n11846), .Z(n11735) );
  AND U15435 ( .A(n10), .B(n11847), .Z(n11845) );
  XOR U15436 ( .A(n11848), .B(n11846), .Z(n11847) );
  XNOR U15437 ( .A(n11849), .B(n11850), .Z(n11837) );
  AND U15438 ( .A(n11851), .B(n11852), .Z(n11849) );
  XOR U15439 ( .A(n11850), .B(n11760), .Z(n11852) );
  XOR U15440 ( .A(n11853), .B(n11844), .Z(n11760) );
  XNOR U15441 ( .A(n11854), .B(n11855), .Z(n11844) );
  ANDN U15442 ( .B(n11856), .A(n11857), .Z(n11854) );
  XOR U15443 ( .A(n11858), .B(n11859), .Z(n11856) );
  IV U15444 ( .A(n11843), .Z(n11853) );
  XOR U15445 ( .A(n11860), .B(n11861), .Z(n11843) );
  XNOR U15446 ( .A(n11862), .B(n11863), .Z(n11861) );
  ANDN U15447 ( .B(n11864), .A(n11865), .Z(n11862) );
  XNOR U15448 ( .A(n11866), .B(n11867), .Z(n11864) );
  IV U15449 ( .A(n11841), .Z(n11860) );
  XOR U15450 ( .A(n11868), .B(n11869), .Z(n11841) );
  ANDN U15451 ( .B(n11870), .A(n11871), .Z(n11868) );
  XOR U15452 ( .A(n11869), .B(n11872), .Z(n11870) );
  XOR U15453 ( .A(n11850), .B(n11762), .Z(n11851) );
  XOR U15454 ( .A(n11873), .B(n11874), .Z(n11762) );
  AND U15455 ( .A(n10), .B(n11875), .Z(n11873) );
  XOR U15456 ( .A(n11876), .B(n11874), .Z(n11875) );
  XNOR U15457 ( .A(n11877), .B(n11878), .Z(n11850) );
  NAND U15458 ( .A(n11879), .B(n11880), .Z(n11878) );
  XOR U15459 ( .A(n11881), .B(n11812), .Z(n11880) );
  XNOR U15460 ( .A(n11882), .B(n11872), .Z(n11812) );
  XOR U15461 ( .A(n11883), .B(n11859), .Z(n11872) );
  XOR U15462 ( .A(n11884), .B(n11885), .Z(n11859) );
  ANDN U15463 ( .B(n11886), .A(n11887), .Z(n11884) );
  XOR U15464 ( .A(n11885), .B(n11888), .Z(n11886) );
  IV U15465 ( .A(n11857), .Z(n11883) );
  XOR U15466 ( .A(n11855), .B(n11889), .Z(n11857) );
  XOR U15467 ( .A(n11890), .B(n11891), .Z(n11889) );
  ANDN U15468 ( .B(n11892), .A(n11893), .Z(n11890) );
  XOR U15469 ( .A(n11894), .B(n11891), .Z(n11892) );
  IV U15470 ( .A(n11858), .Z(n11855) );
  XOR U15471 ( .A(n11895), .B(n11896), .Z(n11858) );
  ANDN U15472 ( .B(n11897), .A(n11898), .Z(n11895) );
  XOR U15473 ( .A(n11896), .B(n11899), .Z(n11897) );
  IV U15474 ( .A(n11871), .Z(n11882) );
  XOR U15475 ( .A(n11900), .B(n11901), .Z(n11871) );
  XNOR U15476 ( .A(n11866), .B(n11902), .Z(n11901) );
  IV U15477 ( .A(n11869), .Z(n11902) );
  XOR U15478 ( .A(n11903), .B(n11904), .Z(n11869) );
  ANDN U15479 ( .B(n11905), .A(n11906), .Z(n11903) );
  XOR U15480 ( .A(n11904), .B(n11907), .Z(n11905) );
  XNOR U15481 ( .A(n11908), .B(n11909), .Z(n11866) );
  ANDN U15482 ( .B(n11910), .A(n11911), .Z(n11908) );
  XOR U15483 ( .A(n11909), .B(n11912), .Z(n11910) );
  IV U15484 ( .A(n11865), .Z(n11900) );
  XOR U15485 ( .A(n11863), .B(n11913), .Z(n11865) );
  XOR U15486 ( .A(n11914), .B(n11915), .Z(n11913) );
  ANDN U15487 ( .B(n11916), .A(n11917), .Z(n11914) );
  XOR U15488 ( .A(n11918), .B(n11915), .Z(n11916) );
  IV U15489 ( .A(n11867), .Z(n11863) );
  XOR U15490 ( .A(n11919), .B(n11920), .Z(n11867) );
  ANDN U15491 ( .B(n11921), .A(n11922), .Z(n11919) );
  XOR U15492 ( .A(n11923), .B(n11920), .Z(n11921) );
  IV U15493 ( .A(n11877), .Z(n11881) );
  XOR U15494 ( .A(n11877), .B(n11816), .Z(n11879) );
  XOR U15495 ( .A(n11924), .B(n11925), .Z(n11816) );
  AND U15496 ( .A(n10), .B(n11926), .Z(n11924) );
  XOR U15497 ( .A(n11927), .B(n11925), .Z(n11926) );
  NANDN U15498 ( .A(n11833), .B(n11835), .Z(n11877) );
  XOR U15499 ( .A(n11928), .B(n11929), .Z(n11835) );
  AND U15500 ( .A(n10), .B(n11930), .Z(n11928) );
  XOR U15501 ( .A(n11929), .B(n11931), .Z(n11930) );
  XNOR U15502 ( .A(n11932), .B(n11933), .Z(n10) );
  AND U15503 ( .A(n11934), .B(n11935), .Z(n11932) );
  XOR U15504 ( .A(n11933), .B(n11846), .Z(n11935) );
  XNOR U15505 ( .A(n11936), .B(n11937), .Z(n11846) );
  ANDN U15506 ( .B(n11938), .A(n11939), .Z(n11936) );
  XOR U15507 ( .A(n11937), .B(n11940), .Z(n11938) );
  XNOR U15508 ( .A(n11933), .B(n11848), .Z(n11934) );
  XOR U15509 ( .A(n11941), .B(n11942), .Z(n11848) );
  AND U15510 ( .A(n14), .B(n11943), .Z(n11941) );
  XOR U15511 ( .A(n11944), .B(n11942), .Z(n11943) );
  XNOR U15512 ( .A(n11945), .B(n11946), .Z(n11933) );
  AND U15513 ( .A(n11947), .B(n11948), .Z(n11945) );
  XNOR U15514 ( .A(n11946), .B(n11874), .Z(n11948) );
  XOR U15515 ( .A(n11939), .B(n11940), .Z(n11874) );
  XNOR U15516 ( .A(n11949), .B(n11950), .Z(n11940) );
  ANDN U15517 ( .B(n11951), .A(n11952), .Z(n11949) );
  XOR U15518 ( .A(n11953), .B(n11954), .Z(n11951) );
  XOR U15519 ( .A(n11955), .B(n11956), .Z(n11939) );
  XNOR U15520 ( .A(n11957), .B(n11958), .Z(n11956) );
  ANDN U15521 ( .B(n11959), .A(n11960), .Z(n11957) );
  XNOR U15522 ( .A(n11961), .B(n11962), .Z(n11959) );
  IV U15523 ( .A(n11937), .Z(n11955) );
  XOR U15524 ( .A(n11963), .B(n11964), .Z(n11937) );
  ANDN U15525 ( .B(n11965), .A(n11966), .Z(n11963) );
  XOR U15526 ( .A(n11964), .B(n11967), .Z(n11965) );
  XOR U15527 ( .A(n11946), .B(n11876), .Z(n11947) );
  XOR U15528 ( .A(n11968), .B(n11969), .Z(n11876) );
  AND U15529 ( .A(n14), .B(n11970), .Z(n11968) );
  XOR U15530 ( .A(n11971), .B(n11969), .Z(n11970) );
  XNOR U15531 ( .A(n11972), .B(n11973), .Z(n11946) );
  NAND U15532 ( .A(n11974), .B(n11975), .Z(n11973) );
  XOR U15533 ( .A(n11976), .B(n11925), .Z(n11975) );
  XOR U15534 ( .A(n11966), .B(n11967), .Z(n11925) );
  XOR U15535 ( .A(n11977), .B(n11954), .Z(n11967) );
  XOR U15536 ( .A(n11978), .B(n11979), .Z(n11954) );
  ANDN U15537 ( .B(n11980), .A(n11981), .Z(n11978) );
  XOR U15538 ( .A(n11979), .B(n11982), .Z(n11980) );
  IV U15539 ( .A(n11952), .Z(n11977) );
  XOR U15540 ( .A(n11950), .B(n11983), .Z(n11952) );
  XOR U15541 ( .A(n11984), .B(n11985), .Z(n11983) );
  ANDN U15542 ( .B(n11986), .A(n11987), .Z(n11984) );
  XOR U15543 ( .A(n11988), .B(n11985), .Z(n11986) );
  IV U15544 ( .A(n11953), .Z(n11950) );
  XOR U15545 ( .A(n11989), .B(n11990), .Z(n11953) );
  ANDN U15546 ( .B(n11991), .A(n11992), .Z(n11989) );
  XOR U15547 ( .A(n11990), .B(n11993), .Z(n11991) );
  XOR U15548 ( .A(n11994), .B(n11995), .Z(n11966) );
  XNOR U15549 ( .A(n11961), .B(n11996), .Z(n11995) );
  IV U15550 ( .A(n11964), .Z(n11996) );
  XOR U15551 ( .A(n11997), .B(n11998), .Z(n11964) );
  ANDN U15552 ( .B(n11999), .A(n12000), .Z(n11997) );
  XOR U15553 ( .A(n11998), .B(n12001), .Z(n11999) );
  XNOR U15554 ( .A(n12002), .B(n12003), .Z(n11961) );
  ANDN U15555 ( .B(n12004), .A(n12005), .Z(n12002) );
  XOR U15556 ( .A(n12003), .B(n12006), .Z(n12004) );
  IV U15557 ( .A(n11960), .Z(n11994) );
  XOR U15558 ( .A(n11958), .B(n12007), .Z(n11960) );
  XOR U15559 ( .A(n12008), .B(n12009), .Z(n12007) );
  ANDN U15560 ( .B(n12010), .A(n12011), .Z(n12008) );
  XOR U15561 ( .A(n12012), .B(n12009), .Z(n12010) );
  IV U15562 ( .A(n11962), .Z(n11958) );
  XOR U15563 ( .A(n12013), .B(n12014), .Z(n11962) );
  ANDN U15564 ( .B(n12015), .A(n12016), .Z(n12013) );
  XOR U15565 ( .A(n12017), .B(n12014), .Z(n12015) );
  IV U15566 ( .A(n11972), .Z(n11976) );
  XOR U15567 ( .A(n11972), .B(n11927), .Z(n11974) );
  XOR U15568 ( .A(n12018), .B(n12019), .Z(n11927) );
  AND U15569 ( .A(n14), .B(n12020), .Z(n12018) );
  XOR U15570 ( .A(n12021), .B(n12019), .Z(n12020) );
  NANDN U15571 ( .A(n11929), .B(n11931), .Z(n11972) );
  XOR U15572 ( .A(n12022), .B(n12023), .Z(n11931) );
  AND U15573 ( .A(n14), .B(n12024), .Z(n12022) );
  XOR U15574 ( .A(n12023), .B(n12025), .Z(n12024) );
  XNOR U15575 ( .A(n12026), .B(n12027), .Z(n14) );
  AND U15576 ( .A(n12028), .B(n12029), .Z(n12026) );
  XOR U15577 ( .A(n12027), .B(n11942), .Z(n12029) );
  XNOR U15578 ( .A(n12030), .B(n12031), .Z(n11942) );
  ANDN U15579 ( .B(n12032), .A(n12033), .Z(n12030) );
  XOR U15580 ( .A(n12031), .B(n12034), .Z(n12032) );
  XNOR U15581 ( .A(n12027), .B(n11944), .Z(n12028) );
  XOR U15582 ( .A(n12035), .B(n12036), .Z(n11944) );
  AND U15583 ( .A(n18), .B(n12037), .Z(n12035) );
  XOR U15584 ( .A(n12038), .B(n12036), .Z(n12037) );
  XNOR U15585 ( .A(n12039), .B(n12040), .Z(n12027) );
  AND U15586 ( .A(n12041), .B(n12042), .Z(n12039) );
  XNOR U15587 ( .A(n12040), .B(n11969), .Z(n12042) );
  XOR U15588 ( .A(n12033), .B(n12034), .Z(n11969) );
  XNOR U15589 ( .A(n12043), .B(n12044), .Z(n12034) );
  ANDN U15590 ( .B(n12045), .A(n12046), .Z(n12043) );
  XOR U15591 ( .A(n12047), .B(n12048), .Z(n12045) );
  XOR U15592 ( .A(n12049), .B(n12050), .Z(n12033) );
  XNOR U15593 ( .A(n12051), .B(n12052), .Z(n12050) );
  ANDN U15594 ( .B(n12053), .A(n12054), .Z(n12051) );
  XNOR U15595 ( .A(n12055), .B(n12056), .Z(n12053) );
  IV U15596 ( .A(n12031), .Z(n12049) );
  XOR U15597 ( .A(n12057), .B(n12058), .Z(n12031) );
  ANDN U15598 ( .B(n12059), .A(n12060), .Z(n12057) );
  XOR U15599 ( .A(n12058), .B(n12061), .Z(n12059) );
  XOR U15600 ( .A(n12040), .B(n11971), .Z(n12041) );
  XOR U15601 ( .A(n12062), .B(n12063), .Z(n11971) );
  AND U15602 ( .A(n18), .B(n12064), .Z(n12062) );
  XOR U15603 ( .A(n12065), .B(n12063), .Z(n12064) );
  XNOR U15604 ( .A(n12066), .B(n12067), .Z(n12040) );
  NAND U15605 ( .A(n12068), .B(n12069), .Z(n12067) );
  XOR U15606 ( .A(n12070), .B(n12019), .Z(n12069) );
  XOR U15607 ( .A(n12060), .B(n12061), .Z(n12019) );
  XOR U15608 ( .A(n12071), .B(n12048), .Z(n12061) );
  XOR U15609 ( .A(n12072), .B(n12073), .Z(n12048) );
  ANDN U15610 ( .B(n12074), .A(n12075), .Z(n12072) );
  XOR U15611 ( .A(n12073), .B(n12076), .Z(n12074) );
  IV U15612 ( .A(n12046), .Z(n12071) );
  XOR U15613 ( .A(n12044), .B(n12077), .Z(n12046) );
  XOR U15614 ( .A(n12078), .B(n12079), .Z(n12077) );
  ANDN U15615 ( .B(n12080), .A(n12081), .Z(n12078) );
  XOR U15616 ( .A(n12082), .B(n12079), .Z(n12080) );
  IV U15617 ( .A(n12047), .Z(n12044) );
  XOR U15618 ( .A(n12083), .B(n12084), .Z(n12047) );
  ANDN U15619 ( .B(n12085), .A(n12086), .Z(n12083) );
  XOR U15620 ( .A(n12084), .B(n12087), .Z(n12085) );
  XOR U15621 ( .A(n12088), .B(n12089), .Z(n12060) );
  XNOR U15622 ( .A(n12055), .B(n12090), .Z(n12089) );
  IV U15623 ( .A(n12058), .Z(n12090) );
  XOR U15624 ( .A(n12091), .B(n12092), .Z(n12058) );
  ANDN U15625 ( .B(n12093), .A(n12094), .Z(n12091) );
  XOR U15626 ( .A(n12092), .B(n12095), .Z(n12093) );
  XNOR U15627 ( .A(n12096), .B(n12097), .Z(n12055) );
  ANDN U15628 ( .B(n12098), .A(n12099), .Z(n12096) );
  XOR U15629 ( .A(n12097), .B(n12100), .Z(n12098) );
  IV U15630 ( .A(n12054), .Z(n12088) );
  XOR U15631 ( .A(n12052), .B(n12101), .Z(n12054) );
  XOR U15632 ( .A(n12102), .B(n12103), .Z(n12101) );
  ANDN U15633 ( .B(n12104), .A(n12105), .Z(n12102) );
  XOR U15634 ( .A(n12106), .B(n12103), .Z(n12104) );
  IV U15635 ( .A(n12056), .Z(n12052) );
  XOR U15636 ( .A(n12107), .B(n12108), .Z(n12056) );
  ANDN U15637 ( .B(n12109), .A(n12110), .Z(n12107) );
  XOR U15638 ( .A(n12111), .B(n12108), .Z(n12109) );
  IV U15639 ( .A(n12066), .Z(n12070) );
  XOR U15640 ( .A(n12066), .B(n12021), .Z(n12068) );
  XOR U15641 ( .A(n12112), .B(n12113), .Z(n12021) );
  AND U15642 ( .A(n18), .B(n12114), .Z(n12112) );
  XOR U15643 ( .A(n12115), .B(n12113), .Z(n12114) );
  NANDN U15644 ( .A(n12023), .B(n12025), .Z(n12066) );
  XOR U15645 ( .A(n12116), .B(n12117), .Z(n12025) );
  AND U15646 ( .A(n18), .B(n12118), .Z(n12116) );
  XOR U15647 ( .A(n12117), .B(n12119), .Z(n12118) );
  XNOR U15648 ( .A(n12120), .B(n12121), .Z(n18) );
  AND U15649 ( .A(n12122), .B(n12123), .Z(n12120) );
  XOR U15650 ( .A(n12121), .B(n12036), .Z(n12123) );
  XNOR U15651 ( .A(n12124), .B(n12125), .Z(n12036) );
  ANDN U15652 ( .B(n12126), .A(n12127), .Z(n12124) );
  XOR U15653 ( .A(n12125), .B(n12128), .Z(n12126) );
  XNOR U15654 ( .A(n12121), .B(n12038), .Z(n12122) );
  XOR U15655 ( .A(n12129), .B(n12130), .Z(n12038) );
  AND U15656 ( .A(n22), .B(n12131), .Z(n12129) );
  XOR U15657 ( .A(n12132), .B(n12130), .Z(n12131) );
  XNOR U15658 ( .A(n12133), .B(n12134), .Z(n12121) );
  AND U15659 ( .A(n12135), .B(n12136), .Z(n12133) );
  XNOR U15660 ( .A(n12134), .B(n12063), .Z(n12136) );
  XOR U15661 ( .A(n12127), .B(n12128), .Z(n12063) );
  XNOR U15662 ( .A(n12137), .B(n12138), .Z(n12128) );
  ANDN U15663 ( .B(n12139), .A(n12140), .Z(n12137) );
  XOR U15664 ( .A(n12141), .B(n12142), .Z(n12139) );
  XOR U15665 ( .A(n12143), .B(n12144), .Z(n12127) );
  XNOR U15666 ( .A(n12145), .B(n12146), .Z(n12144) );
  ANDN U15667 ( .B(n12147), .A(n12148), .Z(n12145) );
  XNOR U15668 ( .A(n12149), .B(n12150), .Z(n12147) );
  IV U15669 ( .A(n12125), .Z(n12143) );
  XOR U15670 ( .A(n12151), .B(n12152), .Z(n12125) );
  ANDN U15671 ( .B(n12153), .A(n12154), .Z(n12151) );
  XOR U15672 ( .A(n12152), .B(n12155), .Z(n12153) );
  XOR U15673 ( .A(n12134), .B(n12065), .Z(n12135) );
  XOR U15674 ( .A(n12156), .B(n12157), .Z(n12065) );
  AND U15675 ( .A(n22), .B(n12158), .Z(n12156) );
  XOR U15676 ( .A(n12159), .B(n12157), .Z(n12158) );
  XNOR U15677 ( .A(n12160), .B(n12161), .Z(n12134) );
  NAND U15678 ( .A(n12162), .B(n12163), .Z(n12161) );
  XOR U15679 ( .A(n12164), .B(n12113), .Z(n12163) );
  XOR U15680 ( .A(n12154), .B(n12155), .Z(n12113) );
  XOR U15681 ( .A(n12165), .B(n12142), .Z(n12155) );
  XOR U15682 ( .A(n12166), .B(n12167), .Z(n12142) );
  ANDN U15683 ( .B(n12168), .A(n12169), .Z(n12166) );
  XOR U15684 ( .A(n12167), .B(n12170), .Z(n12168) );
  IV U15685 ( .A(n12140), .Z(n12165) );
  XOR U15686 ( .A(n12138), .B(n12171), .Z(n12140) );
  XOR U15687 ( .A(n12172), .B(n12173), .Z(n12171) );
  ANDN U15688 ( .B(n12174), .A(n12175), .Z(n12172) );
  XOR U15689 ( .A(n12176), .B(n12173), .Z(n12174) );
  IV U15690 ( .A(n12141), .Z(n12138) );
  XOR U15691 ( .A(n12177), .B(n12178), .Z(n12141) );
  ANDN U15692 ( .B(n12179), .A(n12180), .Z(n12177) );
  XOR U15693 ( .A(n12178), .B(n12181), .Z(n12179) );
  XOR U15694 ( .A(n12182), .B(n12183), .Z(n12154) );
  XNOR U15695 ( .A(n12149), .B(n12184), .Z(n12183) );
  IV U15696 ( .A(n12152), .Z(n12184) );
  XOR U15697 ( .A(n12185), .B(n12186), .Z(n12152) );
  ANDN U15698 ( .B(n12187), .A(n12188), .Z(n12185) );
  XOR U15699 ( .A(n12186), .B(n12189), .Z(n12187) );
  XNOR U15700 ( .A(n12190), .B(n12191), .Z(n12149) );
  ANDN U15701 ( .B(n12192), .A(n12193), .Z(n12190) );
  XOR U15702 ( .A(n12191), .B(n12194), .Z(n12192) );
  IV U15703 ( .A(n12148), .Z(n12182) );
  XOR U15704 ( .A(n12146), .B(n12195), .Z(n12148) );
  XOR U15705 ( .A(n12196), .B(n12197), .Z(n12195) );
  ANDN U15706 ( .B(n12198), .A(n12199), .Z(n12196) );
  XOR U15707 ( .A(n12200), .B(n12197), .Z(n12198) );
  IV U15708 ( .A(n12150), .Z(n12146) );
  XOR U15709 ( .A(n12201), .B(n12202), .Z(n12150) );
  ANDN U15710 ( .B(n12203), .A(n12204), .Z(n12201) );
  XOR U15711 ( .A(n12205), .B(n12202), .Z(n12203) );
  IV U15712 ( .A(n12160), .Z(n12164) );
  XOR U15713 ( .A(n12160), .B(n12115), .Z(n12162) );
  XOR U15714 ( .A(n12206), .B(n12207), .Z(n12115) );
  AND U15715 ( .A(n22), .B(n12208), .Z(n12206) );
  XOR U15716 ( .A(n12209), .B(n12207), .Z(n12208) );
  NANDN U15717 ( .A(n12117), .B(n12119), .Z(n12160) );
  XOR U15718 ( .A(n12210), .B(n12211), .Z(n12119) );
  AND U15719 ( .A(n22), .B(n12212), .Z(n12210) );
  XOR U15720 ( .A(n12211), .B(n12213), .Z(n12212) );
  XNOR U15721 ( .A(n12214), .B(n12215), .Z(n22) );
  AND U15722 ( .A(n12216), .B(n12217), .Z(n12214) );
  XOR U15723 ( .A(n12215), .B(n12130), .Z(n12217) );
  XNOR U15724 ( .A(n12218), .B(n12219), .Z(n12130) );
  ANDN U15725 ( .B(n12220), .A(n12221), .Z(n12218) );
  XOR U15726 ( .A(n12219), .B(n12222), .Z(n12220) );
  XNOR U15727 ( .A(n12215), .B(n12132), .Z(n12216) );
  XOR U15728 ( .A(n12223), .B(n12224), .Z(n12132) );
  AND U15729 ( .A(n26), .B(n12225), .Z(n12223) );
  XOR U15730 ( .A(n12226), .B(n12224), .Z(n12225) );
  XNOR U15731 ( .A(n12227), .B(n12228), .Z(n12215) );
  AND U15732 ( .A(n12229), .B(n12230), .Z(n12227) );
  XNOR U15733 ( .A(n12228), .B(n12157), .Z(n12230) );
  XOR U15734 ( .A(n12221), .B(n12222), .Z(n12157) );
  XNOR U15735 ( .A(n12231), .B(n12232), .Z(n12222) );
  ANDN U15736 ( .B(n12233), .A(n12234), .Z(n12231) );
  XOR U15737 ( .A(n12235), .B(n12236), .Z(n12233) );
  XOR U15738 ( .A(n12237), .B(n12238), .Z(n12221) );
  XNOR U15739 ( .A(n12239), .B(n12240), .Z(n12238) );
  ANDN U15740 ( .B(n12241), .A(n12242), .Z(n12239) );
  XNOR U15741 ( .A(n12243), .B(n12244), .Z(n12241) );
  IV U15742 ( .A(n12219), .Z(n12237) );
  XOR U15743 ( .A(n12245), .B(n12246), .Z(n12219) );
  ANDN U15744 ( .B(n12247), .A(n12248), .Z(n12245) );
  XOR U15745 ( .A(n12246), .B(n12249), .Z(n12247) );
  XOR U15746 ( .A(n12228), .B(n12159), .Z(n12229) );
  XOR U15747 ( .A(n12250), .B(n12251), .Z(n12159) );
  AND U15748 ( .A(n26), .B(n12252), .Z(n12250) );
  XOR U15749 ( .A(n12253), .B(n12251), .Z(n12252) );
  XNOR U15750 ( .A(n12254), .B(n12255), .Z(n12228) );
  NAND U15751 ( .A(n12256), .B(n12257), .Z(n12255) );
  XOR U15752 ( .A(n12258), .B(n12207), .Z(n12257) );
  XOR U15753 ( .A(n12248), .B(n12249), .Z(n12207) );
  XOR U15754 ( .A(n12259), .B(n12236), .Z(n12249) );
  XOR U15755 ( .A(n12260), .B(n12261), .Z(n12236) );
  ANDN U15756 ( .B(n12262), .A(n12263), .Z(n12260) );
  XOR U15757 ( .A(n12261), .B(n12264), .Z(n12262) );
  IV U15758 ( .A(n12234), .Z(n12259) );
  XOR U15759 ( .A(n12232), .B(n12265), .Z(n12234) );
  XOR U15760 ( .A(n12266), .B(n12267), .Z(n12265) );
  ANDN U15761 ( .B(n12268), .A(n12269), .Z(n12266) );
  XOR U15762 ( .A(n12270), .B(n12267), .Z(n12268) );
  IV U15763 ( .A(n12235), .Z(n12232) );
  XOR U15764 ( .A(n12271), .B(n12272), .Z(n12235) );
  ANDN U15765 ( .B(n12273), .A(n12274), .Z(n12271) );
  XOR U15766 ( .A(n12272), .B(n12275), .Z(n12273) );
  XOR U15767 ( .A(n12276), .B(n12277), .Z(n12248) );
  XNOR U15768 ( .A(n12243), .B(n12278), .Z(n12277) );
  IV U15769 ( .A(n12246), .Z(n12278) );
  XOR U15770 ( .A(n12279), .B(n12280), .Z(n12246) );
  ANDN U15771 ( .B(n12281), .A(n12282), .Z(n12279) );
  XOR U15772 ( .A(n12280), .B(n12283), .Z(n12281) );
  XNOR U15773 ( .A(n12284), .B(n12285), .Z(n12243) );
  ANDN U15774 ( .B(n12286), .A(n12287), .Z(n12284) );
  XOR U15775 ( .A(n12285), .B(n12288), .Z(n12286) );
  IV U15776 ( .A(n12242), .Z(n12276) );
  XOR U15777 ( .A(n12240), .B(n12289), .Z(n12242) );
  XOR U15778 ( .A(n12290), .B(n12291), .Z(n12289) );
  ANDN U15779 ( .B(n12292), .A(n12293), .Z(n12290) );
  XOR U15780 ( .A(n12294), .B(n12291), .Z(n12292) );
  IV U15781 ( .A(n12244), .Z(n12240) );
  XOR U15782 ( .A(n12295), .B(n12296), .Z(n12244) );
  ANDN U15783 ( .B(n12297), .A(n12298), .Z(n12295) );
  XOR U15784 ( .A(n12299), .B(n12296), .Z(n12297) );
  IV U15785 ( .A(n12254), .Z(n12258) );
  XOR U15786 ( .A(n12254), .B(n12209), .Z(n12256) );
  XOR U15787 ( .A(n12300), .B(n12301), .Z(n12209) );
  AND U15788 ( .A(n26), .B(n12302), .Z(n12300) );
  XOR U15789 ( .A(n12303), .B(n12301), .Z(n12302) );
  NANDN U15790 ( .A(n12211), .B(n12213), .Z(n12254) );
  XOR U15791 ( .A(n12304), .B(n12305), .Z(n12213) );
  AND U15792 ( .A(n26), .B(n12306), .Z(n12304) );
  XOR U15793 ( .A(n12305), .B(n12307), .Z(n12306) );
  XNOR U15794 ( .A(n12308), .B(n12309), .Z(n26) );
  AND U15795 ( .A(n12310), .B(n12311), .Z(n12308) );
  XOR U15796 ( .A(n12309), .B(n12224), .Z(n12311) );
  XNOR U15797 ( .A(n12312), .B(n12313), .Z(n12224) );
  ANDN U15798 ( .B(n12314), .A(n12315), .Z(n12312) );
  XOR U15799 ( .A(n12313), .B(n12316), .Z(n12314) );
  XNOR U15800 ( .A(n12309), .B(n12226), .Z(n12310) );
  XOR U15801 ( .A(n12317), .B(n12318), .Z(n12226) );
  AND U15802 ( .A(n30), .B(n12319), .Z(n12317) );
  XOR U15803 ( .A(n12320), .B(n12318), .Z(n12319) );
  XNOR U15804 ( .A(n12321), .B(n12322), .Z(n12309) );
  AND U15805 ( .A(n12323), .B(n12324), .Z(n12321) );
  XNOR U15806 ( .A(n12322), .B(n12251), .Z(n12324) );
  XOR U15807 ( .A(n12315), .B(n12316), .Z(n12251) );
  XNOR U15808 ( .A(n12325), .B(n12326), .Z(n12316) );
  ANDN U15809 ( .B(n12327), .A(n12328), .Z(n12325) );
  XOR U15810 ( .A(n12329), .B(n12330), .Z(n12327) );
  XOR U15811 ( .A(n12331), .B(n12332), .Z(n12315) );
  XNOR U15812 ( .A(n12333), .B(n12334), .Z(n12332) );
  ANDN U15813 ( .B(n12335), .A(n12336), .Z(n12333) );
  XNOR U15814 ( .A(n12337), .B(n12338), .Z(n12335) );
  IV U15815 ( .A(n12313), .Z(n12331) );
  XOR U15816 ( .A(n12339), .B(n12340), .Z(n12313) );
  ANDN U15817 ( .B(n12341), .A(n12342), .Z(n12339) );
  XOR U15818 ( .A(n12340), .B(n12343), .Z(n12341) );
  XOR U15819 ( .A(n12322), .B(n12253), .Z(n12323) );
  XOR U15820 ( .A(n12344), .B(n12345), .Z(n12253) );
  AND U15821 ( .A(n30), .B(n12346), .Z(n12344) );
  XOR U15822 ( .A(n12347), .B(n12345), .Z(n12346) );
  XNOR U15823 ( .A(n12348), .B(n12349), .Z(n12322) );
  NAND U15824 ( .A(n12350), .B(n12351), .Z(n12349) );
  XOR U15825 ( .A(n12352), .B(n12301), .Z(n12351) );
  XOR U15826 ( .A(n12342), .B(n12343), .Z(n12301) );
  XOR U15827 ( .A(n12353), .B(n12330), .Z(n12343) );
  XOR U15828 ( .A(n12354), .B(n12355), .Z(n12330) );
  ANDN U15829 ( .B(n12356), .A(n12357), .Z(n12354) );
  XOR U15830 ( .A(n12355), .B(n12358), .Z(n12356) );
  IV U15831 ( .A(n12328), .Z(n12353) );
  XOR U15832 ( .A(n12326), .B(n12359), .Z(n12328) );
  XOR U15833 ( .A(n12360), .B(n12361), .Z(n12359) );
  ANDN U15834 ( .B(n12362), .A(n12363), .Z(n12360) );
  XOR U15835 ( .A(n12364), .B(n12361), .Z(n12362) );
  IV U15836 ( .A(n12329), .Z(n12326) );
  XOR U15837 ( .A(n12365), .B(n12366), .Z(n12329) );
  ANDN U15838 ( .B(n12367), .A(n12368), .Z(n12365) );
  XOR U15839 ( .A(n12366), .B(n12369), .Z(n12367) );
  XOR U15840 ( .A(n12370), .B(n12371), .Z(n12342) );
  XNOR U15841 ( .A(n12337), .B(n12372), .Z(n12371) );
  IV U15842 ( .A(n12340), .Z(n12372) );
  XOR U15843 ( .A(n12373), .B(n12374), .Z(n12340) );
  ANDN U15844 ( .B(n12375), .A(n12376), .Z(n12373) );
  XOR U15845 ( .A(n12374), .B(n12377), .Z(n12375) );
  XNOR U15846 ( .A(n12378), .B(n12379), .Z(n12337) );
  ANDN U15847 ( .B(n12380), .A(n12381), .Z(n12378) );
  XOR U15848 ( .A(n12379), .B(n12382), .Z(n12380) );
  IV U15849 ( .A(n12336), .Z(n12370) );
  XOR U15850 ( .A(n12334), .B(n12383), .Z(n12336) );
  XOR U15851 ( .A(n12384), .B(n12385), .Z(n12383) );
  ANDN U15852 ( .B(n12386), .A(n12387), .Z(n12384) );
  XOR U15853 ( .A(n12388), .B(n12385), .Z(n12386) );
  IV U15854 ( .A(n12338), .Z(n12334) );
  XOR U15855 ( .A(n12389), .B(n12390), .Z(n12338) );
  ANDN U15856 ( .B(n12391), .A(n12392), .Z(n12389) );
  XOR U15857 ( .A(n12393), .B(n12390), .Z(n12391) );
  IV U15858 ( .A(n12348), .Z(n12352) );
  XOR U15859 ( .A(n12348), .B(n12303), .Z(n12350) );
  XOR U15860 ( .A(n12394), .B(n12395), .Z(n12303) );
  AND U15861 ( .A(n30), .B(n12396), .Z(n12394) );
  XOR U15862 ( .A(n12397), .B(n12395), .Z(n12396) );
  NANDN U15863 ( .A(n12305), .B(n12307), .Z(n12348) );
  XOR U15864 ( .A(n12398), .B(n12399), .Z(n12307) );
  AND U15865 ( .A(n30), .B(n12400), .Z(n12398) );
  XOR U15866 ( .A(n12399), .B(n12401), .Z(n12400) );
  XNOR U15867 ( .A(n12402), .B(n12403), .Z(n30) );
  AND U15868 ( .A(n12404), .B(n12405), .Z(n12402) );
  XOR U15869 ( .A(n12403), .B(n12318), .Z(n12405) );
  XNOR U15870 ( .A(n12406), .B(n12407), .Z(n12318) );
  ANDN U15871 ( .B(n12408), .A(n12409), .Z(n12406) );
  XOR U15872 ( .A(n12407), .B(n12410), .Z(n12408) );
  XNOR U15873 ( .A(n12403), .B(n12320), .Z(n12404) );
  XOR U15874 ( .A(n12411), .B(n12412), .Z(n12320) );
  AND U15875 ( .A(n34), .B(n12413), .Z(n12411) );
  XOR U15876 ( .A(n12414), .B(n12412), .Z(n12413) );
  XNOR U15877 ( .A(n12415), .B(n12416), .Z(n12403) );
  AND U15878 ( .A(n12417), .B(n12418), .Z(n12415) );
  XNOR U15879 ( .A(n12416), .B(n12345), .Z(n12418) );
  XOR U15880 ( .A(n12409), .B(n12410), .Z(n12345) );
  XNOR U15881 ( .A(n12419), .B(n12420), .Z(n12410) );
  ANDN U15882 ( .B(n12421), .A(n12422), .Z(n12419) );
  XOR U15883 ( .A(n12423), .B(n12424), .Z(n12421) );
  XOR U15884 ( .A(n12425), .B(n12426), .Z(n12409) );
  XNOR U15885 ( .A(n12427), .B(n12428), .Z(n12426) );
  ANDN U15886 ( .B(n12429), .A(n12430), .Z(n12427) );
  XNOR U15887 ( .A(n12431), .B(n12432), .Z(n12429) );
  IV U15888 ( .A(n12407), .Z(n12425) );
  XOR U15889 ( .A(n12433), .B(n12434), .Z(n12407) );
  ANDN U15890 ( .B(n12435), .A(n12436), .Z(n12433) );
  XOR U15891 ( .A(n12434), .B(n12437), .Z(n12435) );
  XOR U15892 ( .A(n12416), .B(n12347), .Z(n12417) );
  XOR U15893 ( .A(n12438), .B(n12439), .Z(n12347) );
  AND U15894 ( .A(n34), .B(n12440), .Z(n12438) );
  XOR U15895 ( .A(n12441), .B(n12439), .Z(n12440) );
  XNOR U15896 ( .A(n12442), .B(n12443), .Z(n12416) );
  NAND U15897 ( .A(n12444), .B(n12445), .Z(n12443) );
  XOR U15898 ( .A(n12446), .B(n12395), .Z(n12445) );
  XOR U15899 ( .A(n12436), .B(n12437), .Z(n12395) );
  XOR U15900 ( .A(n12447), .B(n12424), .Z(n12437) );
  XOR U15901 ( .A(n12448), .B(n12449), .Z(n12424) );
  ANDN U15902 ( .B(n12450), .A(n12451), .Z(n12448) );
  XOR U15903 ( .A(n12449), .B(n12452), .Z(n12450) );
  IV U15904 ( .A(n12422), .Z(n12447) );
  XOR U15905 ( .A(n12420), .B(n12453), .Z(n12422) );
  XOR U15906 ( .A(n12454), .B(n12455), .Z(n12453) );
  ANDN U15907 ( .B(n12456), .A(n12457), .Z(n12454) );
  XOR U15908 ( .A(n12458), .B(n12455), .Z(n12456) );
  IV U15909 ( .A(n12423), .Z(n12420) );
  XOR U15910 ( .A(n12459), .B(n12460), .Z(n12423) );
  ANDN U15911 ( .B(n12461), .A(n12462), .Z(n12459) );
  XOR U15912 ( .A(n12460), .B(n12463), .Z(n12461) );
  XOR U15913 ( .A(n12464), .B(n12465), .Z(n12436) );
  XNOR U15914 ( .A(n12431), .B(n12466), .Z(n12465) );
  IV U15915 ( .A(n12434), .Z(n12466) );
  XOR U15916 ( .A(n12467), .B(n12468), .Z(n12434) );
  ANDN U15917 ( .B(n12469), .A(n12470), .Z(n12467) );
  XOR U15918 ( .A(n12468), .B(n12471), .Z(n12469) );
  XNOR U15919 ( .A(n12472), .B(n12473), .Z(n12431) );
  ANDN U15920 ( .B(n12474), .A(n12475), .Z(n12472) );
  XOR U15921 ( .A(n12473), .B(n12476), .Z(n12474) );
  IV U15922 ( .A(n12430), .Z(n12464) );
  XOR U15923 ( .A(n12428), .B(n12477), .Z(n12430) );
  XOR U15924 ( .A(n12478), .B(n12479), .Z(n12477) );
  ANDN U15925 ( .B(n12480), .A(n12481), .Z(n12478) );
  XOR U15926 ( .A(n12482), .B(n12479), .Z(n12480) );
  IV U15927 ( .A(n12432), .Z(n12428) );
  XOR U15928 ( .A(n12483), .B(n12484), .Z(n12432) );
  ANDN U15929 ( .B(n12485), .A(n12486), .Z(n12483) );
  XOR U15930 ( .A(n12487), .B(n12484), .Z(n12485) );
  IV U15931 ( .A(n12442), .Z(n12446) );
  XOR U15932 ( .A(n12442), .B(n12397), .Z(n12444) );
  XOR U15933 ( .A(n12488), .B(n12489), .Z(n12397) );
  AND U15934 ( .A(n34), .B(n12490), .Z(n12488) );
  XOR U15935 ( .A(n12491), .B(n12489), .Z(n12490) );
  NANDN U15936 ( .A(n12399), .B(n12401), .Z(n12442) );
  XOR U15937 ( .A(n12492), .B(n12493), .Z(n12401) );
  AND U15938 ( .A(n34), .B(n12494), .Z(n12492) );
  XOR U15939 ( .A(n12493), .B(n12495), .Z(n12494) );
  XNOR U15940 ( .A(n12496), .B(n12497), .Z(n34) );
  AND U15941 ( .A(n12498), .B(n12499), .Z(n12496) );
  XOR U15942 ( .A(n12497), .B(n12412), .Z(n12499) );
  XNOR U15943 ( .A(n12500), .B(n12501), .Z(n12412) );
  ANDN U15944 ( .B(n12502), .A(n12503), .Z(n12500) );
  XOR U15945 ( .A(n12501), .B(n12504), .Z(n12502) );
  XNOR U15946 ( .A(n12497), .B(n12414), .Z(n12498) );
  XOR U15947 ( .A(n12505), .B(n12506), .Z(n12414) );
  AND U15948 ( .A(n38), .B(n12507), .Z(n12505) );
  XOR U15949 ( .A(n12508), .B(n12506), .Z(n12507) );
  XNOR U15950 ( .A(n12509), .B(n12510), .Z(n12497) );
  AND U15951 ( .A(n12511), .B(n12512), .Z(n12509) );
  XNOR U15952 ( .A(n12510), .B(n12439), .Z(n12512) );
  XOR U15953 ( .A(n12503), .B(n12504), .Z(n12439) );
  XNOR U15954 ( .A(n12513), .B(n12514), .Z(n12504) );
  ANDN U15955 ( .B(n12515), .A(n12516), .Z(n12513) );
  XOR U15956 ( .A(n12517), .B(n12518), .Z(n12515) );
  XOR U15957 ( .A(n12519), .B(n12520), .Z(n12503) );
  XNOR U15958 ( .A(n12521), .B(n12522), .Z(n12520) );
  ANDN U15959 ( .B(n12523), .A(n12524), .Z(n12521) );
  XNOR U15960 ( .A(n12525), .B(n12526), .Z(n12523) );
  IV U15961 ( .A(n12501), .Z(n12519) );
  XOR U15962 ( .A(n12527), .B(n12528), .Z(n12501) );
  ANDN U15963 ( .B(n12529), .A(n12530), .Z(n12527) );
  XOR U15964 ( .A(n12528), .B(n12531), .Z(n12529) );
  XOR U15965 ( .A(n12510), .B(n12441), .Z(n12511) );
  XOR U15966 ( .A(n12532), .B(n12533), .Z(n12441) );
  AND U15967 ( .A(n38), .B(n12534), .Z(n12532) );
  XOR U15968 ( .A(n12535), .B(n12533), .Z(n12534) );
  XNOR U15969 ( .A(n12536), .B(n12537), .Z(n12510) );
  NAND U15970 ( .A(n12538), .B(n12539), .Z(n12537) );
  XOR U15971 ( .A(n12540), .B(n12489), .Z(n12539) );
  XOR U15972 ( .A(n12530), .B(n12531), .Z(n12489) );
  XOR U15973 ( .A(n12541), .B(n12518), .Z(n12531) );
  XOR U15974 ( .A(n12542), .B(n12543), .Z(n12518) );
  ANDN U15975 ( .B(n12544), .A(n12545), .Z(n12542) );
  XOR U15976 ( .A(n12543), .B(n12546), .Z(n12544) );
  IV U15977 ( .A(n12516), .Z(n12541) );
  XOR U15978 ( .A(n12514), .B(n12547), .Z(n12516) );
  XOR U15979 ( .A(n12548), .B(n12549), .Z(n12547) );
  ANDN U15980 ( .B(n12550), .A(n12551), .Z(n12548) );
  XOR U15981 ( .A(n12552), .B(n12549), .Z(n12550) );
  IV U15982 ( .A(n12517), .Z(n12514) );
  XOR U15983 ( .A(n12553), .B(n12554), .Z(n12517) );
  ANDN U15984 ( .B(n12555), .A(n12556), .Z(n12553) );
  XOR U15985 ( .A(n12554), .B(n12557), .Z(n12555) );
  XOR U15986 ( .A(n12558), .B(n12559), .Z(n12530) );
  XNOR U15987 ( .A(n12525), .B(n12560), .Z(n12559) );
  IV U15988 ( .A(n12528), .Z(n12560) );
  XOR U15989 ( .A(n12561), .B(n12562), .Z(n12528) );
  ANDN U15990 ( .B(n12563), .A(n12564), .Z(n12561) );
  XOR U15991 ( .A(n12562), .B(n12565), .Z(n12563) );
  XNOR U15992 ( .A(n12566), .B(n12567), .Z(n12525) );
  ANDN U15993 ( .B(n12568), .A(n12569), .Z(n12566) );
  XOR U15994 ( .A(n12567), .B(n12570), .Z(n12568) );
  IV U15995 ( .A(n12524), .Z(n12558) );
  XOR U15996 ( .A(n12522), .B(n12571), .Z(n12524) );
  XOR U15997 ( .A(n12572), .B(n12573), .Z(n12571) );
  ANDN U15998 ( .B(n12574), .A(n12575), .Z(n12572) );
  XOR U15999 ( .A(n12576), .B(n12573), .Z(n12574) );
  IV U16000 ( .A(n12526), .Z(n12522) );
  XOR U16001 ( .A(n12577), .B(n12578), .Z(n12526) );
  ANDN U16002 ( .B(n12579), .A(n12580), .Z(n12577) );
  XOR U16003 ( .A(n12581), .B(n12578), .Z(n12579) );
  IV U16004 ( .A(n12536), .Z(n12540) );
  XOR U16005 ( .A(n12536), .B(n12491), .Z(n12538) );
  XOR U16006 ( .A(n12582), .B(n12583), .Z(n12491) );
  AND U16007 ( .A(n38), .B(n12584), .Z(n12582) );
  XOR U16008 ( .A(n12585), .B(n12583), .Z(n12584) );
  NANDN U16009 ( .A(n12493), .B(n12495), .Z(n12536) );
  XOR U16010 ( .A(n12586), .B(n12587), .Z(n12495) );
  AND U16011 ( .A(n38), .B(n12588), .Z(n12586) );
  XOR U16012 ( .A(n12587), .B(n12589), .Z(n12588) );
  XNOR U16013 ( .A(n12590), .B(n12591), .Z(n38) );
  AND U16014 ( .A(n12592), .B(n12593), .Z(n12590) );
  XOR U16015 ( .A(n12591), .B(n12506), .Z(n12593) );
  XNOR U16016 ( .A(n12594), .B(n12595), .Z(n12506) );
  ANDN U16017 ( .B(n12596), .A(n12597), .Z(n12594) );
  XOR U16018 ( .A(n12595), .B(n12598), .Z(n12596) );
  XNOR U16019 ( .A(n12591), .B(n12508), .Z(n12592) );
  XOR U16020 ( .A(n12599), .B(n12600), .Z(n12508) );
  AND U16021 ( .A(n42), .B(n12601), .Z(n12599) );
  XOR U16022 ( .A(n12602), .B(n12600), .Z(n12601) );
  XNOR U16023 ( .A(n12603), .B(n12604), .Z(n12591) );
  AND U16024 ( .A(n12605), .B(n12606), .Z(n12603) );
  XNOR U16025 ( .A(n12604), .B(n12533), .Z(n12606) );
  XOR U16026 ( .A(n12597), .B(n12598), .Z(n12533) );
  XNOR U16027 ( .A(n12607), .B(n12608), .Z(n12598) );
  ANDN U16028 ( .B(n12609), .A(n12610), .Z(n12607) );
  XOR U16029 ( .A(n12611), .B(n12612), .Z(n12609) );
  XOR U16030 ( .A(n12613), .B(n12614), .Z(n12597) );
  XNOR U16031 ( .A(n12615), .B(n12616), .Z(n12614) );
  ANDN U16032 ( .B(n12617), .A(n12618), .Z(n12615) );
  XNOR U16033 ( .A(n12619), .B(n12620), .Z(n12617) );
  IV U16034 ( .A(n12595), .Z(n12613) );
  XOR U16035 ( .A(n12621), .B(n12622), .Z(n12595) );
  ANDN U16036 ( .B(n12623), .A(n12624), .Z(n12621) );
  XOR U16037 ( .A(n12622), .B(n12625), .Z(n12623) );
  XOR U16038 ( .A(n12604), .B(n12535), .Z(n12605) );
  XOR U16039 ( .A(n12626), .B(n12627), .Z(n12535) );
  AND U16040 ( .A(n42), .B(n12628), .Z(n12626) );
  XOR U16041 ( .A(n12629), .B(n12627), .Z(n12628) );
  XNOR U16042 ( .A(n12630), .B(n12631), .Z(n12604) );
  NAND U16043 ( .A(n12632), .B(n12633), .Z(n12631) );
  XOR U16044 ( .A(n12634), .B(n12583), .Z(n12633) );
  XOR U16045 ( .A(n12624), .B(n12625), .Z(n12583) );
  XOR U16046 ( .A(n12635), .B(n12612), .Z(n12625) );
  XOR U16047 ( .A(n12636), .B(n12637), .Z(n12612) );
  ANDN U16048 ( .B(n12638), .A(n12639), .Z(n12636) );
  XOR U16049 ( .A(n12637), .B(n12640), .Z(n12638) );
  IV U16050 ( .A(n12610), .Z(n12635) );
  XOR U16051 ( .A(n12608), .B(n12641), .Z(n12610) );
  XOR U16052 ( .A(n12642), .B(n12643), .Z(n12641) );
  ANDN U16053 ( .B(n12644), .A(n12645), .Z(n12642) );
  XOR U16054 ( .A(n12646), .B(n12643), .Z(n12644) );
  IV U16055 ( .A(n12611), .Z(n12608) );
  XOR U16056 ( .A(n12647), .B(n12648), .Z(n12611) );
  ANDN U16057 ( .B(n12649), .A(n12650), .Z(n12647) );
  XOR U16058 ( .A(n12648), .B(n12651), .Z(n12649) );
  XOR U16059 ( .A(n12652), .B(n12653), .Z(n12624) );
  XNOR U16060 ( .A(n12619), .B(n12654), .Z(n12653) );
  IV U16061 ( .A(n12622), .Z(n12654) );
  XOR U16062 ( .A(n12655), .B(n12656), .Z(n12622) );
  ANDN U16063 ( .B(n12657), .A(n12658), .Z(n12655) );
  XOR U16064 ( .A(n12656), .B(n12659), .Z(n12657) );
  XNOR U16065 ( .A(n12660), .B(n12661), .Z(n12619) );
  ANDN U16066 ( .B(n12662), .A(n12663), .Z(n12660) );
  XOR U16067 ( .A(n12661), .B(n12664), .Z(n12662) );
  IV U16068 ( .A(n12618), .Z(n12652) );
  XOR U16069 ( .A(n12616), .B(n12665), .Z(n12618) );
  XOR U16070 ( .A(n12666), .B(n12667), .Z(n12665) );
  ANDN U16071 ( .B(n12668), .A(n12669), .Z(n12666) );
  XOR U16072 ( .A(n12670), .B(n12667), .Z(n12668) );
  IV U16073 ( .A(n12620), .Z(n12616) );
  XOR U16074 ( .A(n12671), .B(n12672), .Z(n12620) );
  ANDN U16075 ( .B(n12673), .A(n12674), .Z(n12671) );
  XOR U16076 ( .A(n12675), .B(n12672), .Z(n12673) );
  IV U16077 ( .A(n12630), .Z(n12634) );
  XOR U16078 ( .A(n12630), .B(n12585), .Z(n12632) );
  XOR U16079 ( .A(n12676), .B(n12677), .Z(n12585) );
  AND U16080 ( .A(n42), .B(n12678), .Z(n12676) );
  XOR U16081 ( .A(n12679), .B(n12677), .Z(n12678) );
  NANDN U16082 ( .A(n12587), .B(n12589), .Z(n12630) );
  XOR U16083 ( .A(n12680), .B(n12681), .Z(n12589) );
  AND U16084 ( .A(n42), .B(n12682), .Z(n12680) );
  XOR U16085 ( .A(n12681), .B(n12683), .Z(n12682) );
  XNOR U16086 ( .A(n12684), .B(n12685), .Z(n42) );
  AND U16087 ( .A(n12686), .B(n12687), .Z(n12684) );
  XOR U16088 ( .A(n12685), .B(n12600), .Z(n12687) );
  XNOR U16089 ( .A(n12688), .B(n12689), .Z(n12600) );
  ANDN U16090 ( .B(n12690), .A(n12691), .Z(n12688) );
  XOR U16091 ( .A(n12689), .B(n12692), .Z(n12690) );
  XNOR U16092 ( .A(n12685), .B(n12602), .Z(n12686) );
  XOR U16093 ( .A(n12693), .B(n12694), .Z(n12602) );
  AND U16094 ( .A(n46), .B(n12695), .Z(n12693) );
  XOR U16095 ( .A(n12696), .B(n12694), .Z(n12695) );
  XNOR U16096 ( .A(n12697), .B(n12698), .Z(n12685) );
  AND U16097 ( .A(n12699), .B(n12700), .Z(n12697) );
  XNOR U16098 ( .A(n12698), .B(n12627), .Z(n12700) );
  XOR U16099 ( .A(n12691), .B(n12692), .Z(n12627) );
  XNOR U16100 ( .A(n12701), .B(n12702), .Z(n12692) );
  ANDN U16101 ( .B(n12703), .A(n12704), .Z(n12701) );
  XOR U16102 ( .A(n12705), .B(n12706), .Z(n12703) );
  XOR U16103 ( .A(n12707), .B(n12708), .Z(n12691) );
  XNOR U16104 ( .A(n12709), .B(n12710), .Z(n12708) );
  ANDN U16105 ( .B(n12711), .A(n12712), .Z(n12709) );
  XNOR U16106 ( .A(n12713), .B(n12714), .Z(n12711) );
  IV U16107 ( .A(n12689), .Z(n12707) );
  XOR U16108 ( .A(n12715), .B(n12716), .Z(n12689) );
  ANDN U16109 ( .B(n12717), .A(n12718), .Z(n12715) );
  XOR U16110 ( .A(n12716), .B(n12719), .Z(n12717) );
  XOR U16111 ( .A(n12698), .B(n12629), .Z(n12699) );
  XOR U16112 ( .A(n12720), .B(n12721), .Z(n12629) );
  AND U16113 ( .A(n46), .B(n12722), .Z(n12720) );
  XOR U16114 ( .A(n12723), .B(n12721), .Z(n12722) );
  XNOR U16115 ( .A(n12724), .B(n12725), .Z(n12698) );
  NAND U16116 ( .A(n12726), .B(n12727), .Z(n12725) );
  XOR U16117 ( .A(n12728), .B(n12677), .Z(n12727) );
  XOR U16118 ( .A(n12718), .B(n12719), .Z(n12677) );
  XOR U16119 ( .A(n12729), .B(n12706), .Z(n12719) );
  XOR U16120 ( .A(n12730), .B(n12731), .Z(n12706) );
  ANDN U16121 ( .B(n12732), .A(n12733), .Z(n12730) );
  XOR U16122 ( .A(n12731), .B(n12734), .Z(n12732) );
  IV U16123 ( .A(n12704), .Z(n12729) );
  XOR U16124 ( .A(n12702), .B(n12735), .Z(n12704) );
  XOR U16125 ( .A(n12736), .B(n12737), .Z(n12735) );
  ANDN U16126 ( .B(n12738), .A(n12739), .Z(n12736) );
  XOR U16127 ( .A(n12740), .B(n12737), .Z(n12738) );
  IV U16128 ( .A(n12705), .Z(n12702) );
  XOR U16129 ( .A(n12741), .B(n12742), .Z(n12705) );
  ANDN U16130 ( .B(n12743), .A(n12744), .Z(n12741) );
  XOR U16131 ( .A(n12742), .B(n12745), .Z(n12743) );
  XOR U16132 ( .A(n12746), .B(n12747), .Z(n12718) );
  XNOR U16133 ( .A(n12713), .B(n12748), .Z(n12747) );
  IV U16134 ( .A(n12716), .Z(n12748) );
  XOR U16135 ( .A(n12749), .B(n12750), .Z(n12716) );
  ANDN U16136 ( .B(n12751), .A(n12752), .Z(n12749) );
  XOR U16137 ( .A(n12750), .B(n12753), .Z(n12751) );
  XNOR U16138 ( .A(n12754), .B(n12755), .Z(n12713) );
  ANDN U16139 ( .B(n12756), .A(n12757), .Z(n12754) );
  XOR U16140 ( .A(n12755), .B(n12758), .Z(n12756) );
  IV U16141 ( .A(n12712), .Z(n12746) );
  XOR U16142 ( .A(n12710), .B(n12759), .Z(n12712) );
  XOR U16143 ( .A(n12760), .B(n12761), .Z(n12759) );
  ANDN U16144 ( .B(n12762), .A(n12763), .Z(n12760) );
  XOR U16145 ( .A(n12764), .B(n12761), .Z(n12762) );
  IV U16146 ( .A(n12714), .Z(n12710) );
  XOR U16147 ( .A(n12765), .B(n12766), .Z(n12714) );
  ANDN U16148 ( .B(n12767), .A(n12768), .Z(n12765) );
  XOR U16149 ( .A(n12769), .B(n12766), .Z(n12767) );
  IV U16150 ( .A(n12724), .Z(n12728) );
  XOR U16151 ( .A(n12724), .B(n12679), .Z(n12726) );
  XOR U16152 ( .A(n12770), .B(n12771), .Z(n12679) );
  AND U16153 ( .A(n46), .B(n12772), .Z(n12770) );
  XOR U16154 ( .A(n12773), .B(n12771), .Z(n12772) );
  NANDN U16155 ( .A(n12681), .B(n12683), .Z(n12724) );
  XOR U16156 ( .A(n12774), .B(n12775), .Z(n12683) );
  AND U16157 ( .A(n46), .B(n12776), .Z(n12774) );
  XOR U16158 ( .A(n12775), .B(n12777), .Z(n12776) );
  XNOR U16159 ( .A(n12778), .B(n12779), .Z(n46) );
  AND U16160 ( .A(n12780), .B(n12781), .Z(n12778) );
  XOR U16161 ( .A(n12779), .B(n12694), .Z(n12781) );
  XNOR U16162 ( .A(n12782), .B(n12783), .Z(n12694) );
  ANDN U16163 ( .B(n12784), .A(n12785), .Z(n12782) );
  XOR U16164 ( .A(n12783), .B(n12786), .Z(n12784) );
  XNOR U16165 ( .A(n12779), .B(n12696), .Z(n12780) );
  XOR U16166 ( .A(n12787), .B(n12788), .Z(n12696) );
  AND U16167 ( .A(n50), .B(n12789), .Z(n12787) );
  XOR U16168 ( .A(n12790), .B(n12788), .Z(n12789) );
  XNOR U16169 ( .A(n12791), .B(n12792), .Z(n12779) );
  AND U16170 ( .A(n12793), .B(n12794), .Z(n12791) );
  XNOR U16171 ( .A(n12792), .B(n12721), .Z(n12794) );
  XOR U16172 ( .A(n12785), .B(n12786), .Z(n12721) );
  XNOR U16173 ( .A(n12795), .B(n12796), .Z(n12786) );
  ANDN U16174 ( .B(n12797), .A(n12798), .Z(n12795) );
  XOR U16175 ( .A(n12799), .B(n12800), .Z(n12797) );
  XOR U16176 ( .A(n12801), .B(n12802), .Z(n12785) );
  XNOR U16177 ( .A(n12803), .B(n12804), .Z(n12802) );
  ANDN U16178 ( .B(n12805), .A(n12806), .Z(n12803) );
  XNOR U16179 ( .A(n12807), .B(n12808), .Z(n12805) );
  IV U16180 ( .A(n12783), .Z(n12801) );
  XOR U16181 ( .A(n12809), .B(n12810), .Z(n12783) );
  ANDN U16182 ( .B(n12811), .A(n12812), .Z(n12809) );
  XOR U16183 ( .A(n12810), .B(n12813), .Z(n12811) );
  XOR U16184 ( .A(n12792), .B(n12723), .Z(n12793) );
  XOR U16185 ( .A(n12814), .B(n12815), .Z(n12723) );
  AND U16186 ( .A(n50), .B(n12816), .Z(n12814) );
  XOR U16187 ( .A(n12817), .B(n12815), .Z(n12816) );
  XNOR U16188 ( .A(n12818), .B(n12819), .Z(n12792) );
  NAND U16189 ( .A(n12820), .B(n12821), .Z(n12819) );
  XOR U16190 ( .A(n12822), .B(n12771), .Z(n12821) );
  XOR U16191 ( .A(n12812), .B(n12813), .Z(n12771) );
  XOR U16192 ( .A(n12823), .B(n12800), .Z(n12813) );
  XOR U16193 ( .A(n12824), .B(n12825), .Z(n12800) );
  ANDN U16194 ( .B(n12826), .A(n12827), .Z(n12824) );
  XOR U16195 ( .A(n12825), .B(n12828), .Z(n12826) );
  IV U16196 ( .A(n12798), .Z(n12823) );
  XOR U16197 ( .A(n12796), .B(n12829), .Z(n12798) );
  XOR U16198 ( .A(n12830), .B(n12831), .Z(n12829) );
  ANDN U16199 ( .B(n12832), .A(n12833), .Z(n12830) );
  XOR U16200 ( .A(n12834), .B(n12831), .Z(n12832) );
  IV U16201 ( .A(n12799), .Z(n12796) );
  XOR U16202 ( .A(n12835), .B(n12836), .Z(n12799) );
  ANDN U16203 ( .B(n12837), .A(n12838), .Z(n12835) );
  XOR U16204 ( .A(n12836), .B(n12839), .Z(n12837) );
  XOR U16205 ( .A(n12840), .B(n12841), .Z(n12812) );
  XNOR U16206 ( .A(n12807), .B(n12842), .Z(n12841) );
  IV U16207 ( .A(n12810), .Z(n12842) );
  XOR U16208 ( .A(n12843), .B(n12844), .Z(n12810) );
  ANDN U16209 ( .B(n12845), .A(n12846), .Z(n12843) );
  XOR U16210 ( .A(n12844), .B(n12847), .Z(n12845) );
  XNOR U16211 ( .A(n12848), .B(n12849), .Z(n12807) );
  ANDN U16212 ( .B(n12850), .A(n12851), .Z(n12848) );
  XOR U16213 ( .A(n12849), .B(n12852), .Z(n12850) );
  IV U16214 ( .A(n12806), .Z(n12840) );
  XOR U16215 ( .A(n12804), .B(n12853), .Z(n12806) );
  XOR U16216 ( .A(n12854), .B(n12855), .Z(n12853) );
  ANDN U16217 ( .B(n12856), .A(n12857), .Z(n12854) );
  XOR U16218 ( .A(n12858), .B(n12855), .Z(n12856) );
  IV U16219 ( .A(n12808), .Z(n12804) );
  XOR U16220 ( .A(n12859), .B(n12860), .Z(n12808) );
  ANDN U16221 ( .B(n12861), .A(n12862), .Z(n12859) );
  XOR U16222 ( .A(n12863), .B(n12860), .Z(n12861) );
  IV U16223 ( .A(n12818), .Z(n12822) );
  XOR U16224 ( .A(n12818), .B(n12773), .Z(n12820) );
  XOR U16225 ( .A(n12864), .B(n12865), .Z(n12773) );
  AND U16226 ( .A(n50), .B(n12866), .Z(n12864) );
  XOR U16227 ( .A(n12867), .B(n12865), .Z(n12866) );
  NANDN U16228 ( .A(n12775), .B(n12777), .Z(n12818) );
  XOR U16229 ( .A(n12868), .B(n12869), .Z(n12777) );
  AND U16230 ( .A(n50), .B(n12870), .Z(n12868) );
  XOR U16231 ( .A(n12869), .B(n12871), .Z(n12870) );
  XNOR U16232 ( .A(n12872), .B(n12873), .Z(n50) );
  AND U16233 ( .A(n12874), .B(n12875), .Z(n12872) );
  XOR U16234 ( .A(n12873), .B(n12788), .Z(n12875) );
  XNOR U16235 ( .A(n12876), .B(n12877), .Z(n12788) );
  ANDN U16236 ( .B(n12878), .A(n12879), .Z(n12876) );
  XOR U16237 ( .A(n12877), .B(n12880), .Z(n12878) );
  XNOR U16238 ( .A(n12873), .B(n12790), .Z(n12874) );
  XOR U16239 ( .A(n12881), .B(n12882), .Z(n12790) );
  AND U16240 ( .A(n54), .B(n12883), .Z(n12881) );
  XOR U16241 ( .A(n12884), .B(n12882), .Z(n12883) );
  XNOR U16242 ( .A(n12885), .B(n12886), .Z(n12873) );
  AND U16243 ( .A(n12887), .B(n12888), .Z(n12885) );
  XNOR U16244 ( .A(n12886), .B(n12815), .Z(n12888) );
  XOR U16245 ( .A(n12879), .B(n12880), .Z(n12815) );
  XNOR U16246 ( .A(n12889), .B(n12890), .Z(n12880) );
  ANDN U16247 ( .B(n12891), .A(n12892), .Z(n12889) );
  XOR U16248 ( .A(n12893), .B(n12894), .Z(n12891) );
  XOR U16249 ( .A(n12895), .B(n12896), .Z(n12879) );
  XNOR U16250 ( .A(n12897), .B(n12898), .Z(n12896) );
  ANDN U16251 ( .B(n12899), .A(n12900), .Z(n12897) );
  XNOR U16252 ( .A(n12901), .B(n12902), .Z(n12899) );
  IV U16253 ( .A(n12877), .Z(n12895) );
  XOR U16254 ( .A(n12903), .B(n12904), .Z(n12877) );
  ANDN U16255 ( .B(n12905), .A(n12906), .Z(n12903) );
  XOR U16256 ( .A(n12904), .B(n12907), .Z(n12905) );
  XOR U16257 ( .A(n12886), .B(n12817), .Z(n12887) );
  XOR U16258 ( .A(n12908), .B(n12909), .Z(n12817) );
  AND U16259 ( .A(n54), .B(n12910), .Z(n12908) );
  XOR U16260 ( .A(n12911), .B(n12909), .Z(n12910) );
  XNOR U16261 ( .A(n12912), .B(n12913), .Z(n12886) );
  NAND U16262 ( .A(n12914), .B(n12915), .Z(n12913) );
  XOR U16263 ( .A(n12916), .B(n12865), .Z(n12915) );
  XOR U16264 ( .A(n12906), .B(n12907), .Z(n12865) );
  XOR U16265 ( .A(n12917), .B(n12894), .Z(n12907) );
  XOR U16266 ( .A(n12918), .B(n12919), .Z(n12894) );
  ANDN U16267 ( .B(n12920), .A(n12921), .Z(n12918) );
  XOR U16268 ( .A(n12919), .B(n12922), .Z(n12920) );
  IV U16269 ( .A(n12892), .Z(n12917) );
  XOR U16270 ( .A(n12890), .B(n12923), .Z(n12892) );
  XOR U16271 ( .A(n12924), .B(n12925), .Z(n12923) );
  ANDN U16272 ( .B(n12926), .A(n12927), .Z(n12924) );
  XOR U16273 ( .A(n12928), .B(n12925), .Z(n12926) );
  IV U16274 ( .A(n12893), .Z(n12890) );
  XOR U16275 ( .A(n12929), .B(n12930), .Z(n12893) );
  ANDN U16276 ( .B(n12931), .A(n12932), .Z(n12929) );
  XOR U16277 ( .A(n12930), .B(n12933), .Z(n12931) );
  XOR U16278 ( .A(n12934), .B(n12935), .Z(n12906) );
  XNOR U16279 ( .A(n12901), .B(n12936), .Z(n12935) );
  IV U16280 ( .A(n12904), .Z(n12936) );
  XOR U16281 ( .A(n12937), .B(n12938), .Z(n12904) );
  ANDN U16282 ( .B(n12939), .A(n12940), .Z(n12937) );
  XOR U16283 ( .A(n12938), .B(n12941), .Z(n12939) );
  XNOR U16284 ( .A(n12942), .B(n12943), .Z(n12901) );
  ANDN U16285 ( .B(n12944), .A(n12945), .Z(n12942) );
  XOR U16286 ( .A(n12943), .B(n12946), .Z(n12944) );
  IV U16287 ( .A(n12900), .Z(n12934) );
  XOR U16288 ( .A(n12898), .B(n12947), .Z(n12900) );
  XOR U16289 ( .A(n12948), .B(n12949), .Z(n12947) );
  ANDN U16290 ( .B(n12950), .A(n12951), .Z(n12948) );
  XOR U16291 ( .A(n12952), .B(n12949), .Z(n12950) );
  IV U16292 ( .A(n12902), .Z(n12898) );
  XOR U16293 ( .A(n12953), .B(n12954), .Z(n12902) );
  ANDN U16294 ( .B(n12955), .A(n12956), .Z(n12953) );
  XOR U16295 ( .A(n12957), .B(n12954), .Z(n12955) );
  IV U16296 ( .A(n12912), .Z(n12916) );
  XOR U16297 ( .A(n12912), .B(n12867), .Z(n12914) );
  XOR U16298 ( .A(n12958), .B(n12959), .Z(n12867) );
  AND U16299 ( .A(n54), .B(n12960), .Z(n12958) );
  XOR U16300 ( .A(n12961), .B(n12959), .Z(n12960) );
  NANDN U16301 ( .A(n12869), .B(n12871), .Z(n12912) );
  XOR U16302 ( .A(n12962), .B(n12963), .Z(n12871) );
  AND U16303 ( .A(n54), .B(n12964), .Z(n12962) );
  XOR U16304 ( .A(n12963), .B(n12965), .Z(n12964) );
  XNOR U16305 ( .A(n12966), .B(n12967), .Z(n54) );
  AND U16306 ( .A(n12968), .B(n12969), .Z(n12966) );
  XOR U16307 ( .A(n12967), .B(n12882), .Z(n12969) );
  XNOR U16308 ( .A(n12970), .B(n12971), .Z(n12882) );
  ANDN U16309 ( .B(n12972), .A(n12973), .Z(n12970) );
  XOR U16310 ( .A(n12971), .B(n12974), .Z(n12972) );
  XNOR U16311 ( .A(n12967), .B(n12884), .Z(n12968) );
  XOR U16312 ( .A(n12975), .B(n12976), .Z(n12884) );
  AND U16313 ( .A(n58), .B(n12977), .Z(n12975) );
  XOR U16314 ( .A(n12978), .B(n12976), .Z(n12977) );
  XNOR U16315 ( .A(n12979), .B(n12980), .Z(n12967) );
  AND U16316 ( .A(n12981), .B(n12982), .Z(n12979) );
  XNOR U16317 ( .A(n12980), .B(n12909), .Z(n12982) );
  XOR U16318 ( .A(n12973), .B(n12974), .Z(n12909) );
  XNOR U16319 ( .A(n12983), .B(n12984), .Z(n12974) );
  ANDN U16320 ( .B(n12985), .A(n12986), .Z(n12983) );
  XOR U16321 ( .A(n12987), .B(n12988), .Z(n12985) );
  XOR U16322 ( .A(n12989), .B(n12990), .Z(n12973) );
  XNOR U16323 ( .A(n12991), .B(n12992), .Z(n12990) );
  ANDN U16324 ( .B(n12993), .A(n12994), .Z(n12991) );
  XNOR U16325 ( .A(n12995), .B(n12996), .Z(n12993) );
  IV U16326 ( .A(n12971), .Z(n12989) );
  XOR U16327 ( .A(n12997), .B(n12998), .Z(n12971) );
  ANDN U16328 ( .B(n12999), .A(n13000), .Z(n12997) );
  XOR U16329 ( .A(n12998), .B(n13001), .Z(n12999) );
  XOR U16330 ( .A(n12980), .B(n12911), .Z(n12981) );
  XOR U16331 ( .A(n13002), .B(n13003), .Z(n12911) );
  AND U16332 ( .A(n58), .B(n13004), .Z(n13002) );
  XOR U16333 ( .A(n13005), .B(n13003), .Z(n13004) );
  XNOR U16334 ( .A(n13006), .B(n13007), .Z(n12980) );
  NAND U16335 ( .A(n13008), .B(n13009), .Z(n13007) );
  XOR U16336 ( .A(n13010), .B(n12959), .Z(n13009) );
  XOR U16337 ( .A(n13000), .B(n13001), .Z(n12959) );
  XOR U16338 ( .A(n13011), .B(n12988), .Z(n13001) );
  XOR U16339 ( .A(n13012), .B(n13013), .Z(n12988) );
  ANDN U16340 ( .B(n13014), .A(n13015), .Z(n13012) );
  XOR U16341 ( .A(n13013), .B(n13016), .Z(n13014) );
  IV U16342 ( .A(n12986), .Z(n13011) );
  XOR U16343 ( .A(n12984), .B(n13017), .Z(n12986) );
  XOR U16344 ( .A(n13018), .B(n13019), .Z(n13017) );
  ANDN U16345 ( .B(n13020), .A(n13021), .Z(n13018) );
  XOR U16346 ( .A(n13022), .B(n13019), .Z(n13020) );
  IV U16347 ( .A(n12987), .Z(n12984) );
  XOR U16348 ( .A(n13023), .B(n13024), .Z(n12987) );
  ANDN U16349 ( .B(n13025), .A(n13026), .Z(n13023) );
  XOR U16350 ( .A(n13024), .B(n13027), .Z(n13025) );
  XOR U16351 ( .A(n13028), .B(n13029), .Z(n13000) );
  XNOR U16352 ( .A(n12995), .B(n13030), .Z(n13029) );
  IV U16353 ( .A(n12998), .Z(n13030) );
  XOR U16354 ( .A(n13031), .B(n13032), .Z(n12998) );
  ANDN U16355 ( .B(n13033), .A(n13034), .Z(n13031) );
  XOR U16356 ( .A(n13032), .B(n13035), .Z(n13033) );
  XNOR U16357 ( .A(n13036), .B(n13037), .Z(n12995) );
  ANDN U16358 ( .B(n13038), .A(n13039), .Z(n13036) );
  XOR U16359 ( .A(n13037), .B(n13040), .Z(n13038) );
  IV U16360 ( .A(n12994), .Z(n13028) );
  XOR U16361 ( .A(n12992), .B(n13041), .Z(n12994) );
  XOR U16362 ( .A(n13042), .B(n13043), .Z(n13041) );
  ANDN U16363 ( .B(n13044), .A(n13045), .Z(n13042) );
  XOR U16364 ( .A(n13046), .B(n13043), .Z(n13044) );
  IV U16365 ( .A(n12996), .Z(n12992) );
  XOR U16366 ( .A(n13047), .B(n13048), .Z(n12996) );
  ANDN U16367 ( .B(n13049), .A(n13050), .Z(n13047) );
  XOR U16368 ( .A(n13051), .B(n13048), .Z(n13049) );
  IV U16369 ( .A(n13006), .Z(n13010) );
  XOR U16370 ( .A(n13006), .B(n12961), .Z(n13008) );
  XOR U16371 ( .A(n13052), .B(n13053), .Z(n12961) );
  AND U16372 ( .A(n58), .B(n13054), .Z(n13052) );
  XOR U16373 ( .A(n13055), .B(n13053), .Z(n13054) );
  NANDN U16374 ( .A(n12963), .B(n12965), .Z(n13006) );
  XOR U16375 ( .A(n13056), .B(n13057), .Z(n12965) );
  AND U16376 ( .A(n58), .B(n13058), .Z(n13056) );
  XOR U16377 ( .A(n13057), .B(n13059), .Z(n13058) );
  XNOR U16378 ( .A(n13060), .B(n13061), .Z(n58) );
  AND U16379 ( .A(n13062), .B(n13063), .Z(n13060) );
  XOR U16380 ( .A(n13061), .B(n12976), .Z(n13063) );
  XNOR U16381 ( .A(n13064), .B(n13065), .Z(n12976) );
  ANDN U16382 ( .B(n13066), .A(n13067), .Z(n13064) );
  XOR U16383 ( .A(n13065), .B(n13068), .Z(n13066) );
  XNOR U16384 ( .A(n13061), .B(n12978), .Z(n13062) );
  XOR U16385 ( .A(n13069), .B(n13070), .Z(n12978) );
  AND U16386 ( .A(n62), .B(n13071), .Z(n13069) );
  XOR U16387 ( .A(n13072), .B(n13070), .Z(n13071) );
  XNOR U16388 ( .A(n13073), .B(n13074), .Z(n13061) );
  AND U16389 ( .A(n13075), .B(n13076), .Z(n13073) );
  XNOR U16390 ( .A(n13074), .B(n13003), .Z(n13076) );
  XOR U16391 ( .A(n13067), .B(n13068), .Z(n13003) );
  XNOR U16392 ( .A(n13077), .B(n13078), .Z(n13068) );
  ANDN U16393 ( .B(n13079), .A(n13080), .Z(n13077) );
  XOR U16394 ( .A(n13081), .B(n13082), .Z(n13079) );
  XOR U16395 ( .A(n13083), .B(n13084), .Z(n13067) );
  XNOR U16396 ( .A(n13085), .B(n13086), .Z(n13084) );
  ANDN U16397 ( .B(n13087), .A(n13088), .Z(n13085) );
  XNOR U16398 ( .A(n13089), .B(n13090), .Z(n13087) );
  IV U16399 ( .A(n13065), .Z(n13083) );
  XOR U16400 ( .A(n13091), .B(n13092), .Z(n13065) );
  ANDN U16401 ( .B(n13093), .A(n13094), .Z(n13091) );
  XOR U16402 ( .A(n13092), .B(n13095), .Z(n13093) );
  XOR U16403 ( .A(n13074), .B(n13005), .Z(n13075) );
  XOR U16404 ( .A(n13096), .B(n13097), .Z(n13005) );
  AND U16405 ( .A(n62), .B(n13098), .Z(n13096) );
  XOR U16406 ( .A(n13099), .B(n13097), .Z(n13098) );
  XNOR U16407 ( .A(n13100), .B(n13101), .Z(n13074) );
  NAND U16408 ( .A(n13102), .B(n13103), .Z(n13101) );
  XOR U16409 ( .A(n13104), .B(n13053), .Z(n13103) );
  XOR U16410 ( .A(n13094), .B(n13095), .Z(n13053) );
  XOR U16411 ( .A(n13105), .B(n13082), .Z(n13095) );
  XOR U16412 ( .A(n13106), .B(n13107), .Z(n13082) );
  ANDN U16413 ( .B(n13108), .A(n13109), .Z(n13106) );
  XOR U16414 ( .A(n13107), .B(n13110), .Z(n13108) );
  IV U16415 ( .A(n13080), .Z(n13105) );
  XOR U16416 ( .A(n13078), .B(n13111), .Z(n13080) );
  XOR U16417 ( .A(n13112), .B(n13113), .Z(n13111) );
  ANDN U16418 ( .B(n13114), .A(n13115), .Z(n13112) );
  XOR U16419 ( .A(n13116), .B(n13113), .Z(n13114) );
  IV U16420 ( .A(n13081), .Z(n13078) );
  XOR U16421 ( .A(n13117), .B(n13118), .Z(n13081) );
  ANDN U16422 ( .B(n13119), .A(n13120), .Z(n13117) );
  XOR U16423 ( .A(n13118), .B(n13121), .Z(n13119) );
  XOR U16424 ( .A(n13122), .B(n13123), .Z(n13094) );
  XNOR U16425 ( .A(n13089), .B(n13124), .Z(n13123) );
  IV U16426 ( .A(n13092), .Z(n13124) );
  XOR U16427 ( .A(n13125), .B(n13126), .Z(n13092) );
  ANDN U16428 ( .B(n13127), .A(n13128), .Z(n13125) );
  XOR U16429 ( .A(n13126), .B(n13129), .Z(n13127) );
  XNOR U16430 ( .A(n13130), .B(n13131), .Z(n13089) );
  ANDN U16431 ( .B(n13132), .A(n13133), .Z(n13130) );
  XOR U16432 ( .A(n13131), .B(n13134), .Z(n13132) );
  IV U16433 ( .A(n13088), .Z(n13122) );
  XOR U16434 ( .A(n13086), .B(n13135), .Z(n13088) );
  XOR U16435 ( .A(n13136), .B(n13137), .Z(n13135) );
  ANDN U16436 ( .B(n13138), .A(n13139), .Z(n13136) );
  XOR U16437 ( .A(n13140), .B(n13137), .Z(n13138) );
  IV U16438 ( .A(n13090), .Z(n13086) );
  XOR U16439 ( .A(n13141), .B(n13142), .Z(n13090) );
  ANDN U16440 ( .B(n13143), .A(n13144), .Z(n13141) );
  XOR U16441 ( .A(n13145), .B(n13142), .Z(n13143) );
  IV U16442 ( .A(n13100), .Z(n13104) );
  XOR U16443 ( .A(n13100), .B(n13055), .Z(n13102) );
  XOR U16444 ( .A(n13146), .B(n13147), .Z(n13055) );
  AND U16445 ( .A(n62), .B(n13148), .Z(n13146) );
  XOR U16446 ( .A(n13149), .B(n13147), .Z(n13148) );
  NANDN U16447 ( .A(n13057), .B(n13059), .Z(n13100) );
  XOR U16448 ( .A(n13150), .B(n13151), .Z(n13059) );
  AND U16449 ( .A(n62), .B(n13152), .Z(n13150) );
  XOR U16450 ( .A(n13151), .B(n13153), .Z(n13152) );
  XNOR U16451 ( .A(n13154), .B(n13155), .Z(n62) );
  AND U16452 ( .A(n13156), .B(n13157), .Z(n13154) );
  XOR U16453 ( .A(n13155), .B(n13070), .Z(n13157) );
  XNOR U16454 ( .A(n13158), .B(n13159), .Z(n13070) );
  ANDN U16455 ( .B(n13160), .A(n13161), .Z(n13158) );
  XOR U16456 ( .A(n13159), .B(n13162), .Z(n13160) );
  XNOR U16457 ( .A(n13155), .B(n13072), .Z(n13156) );
  XOR U16458 ( .A(n13163), .B(n13164), .Z(n13072) );
  AND U16459 ( .A(n66), .B(n13165), .Z(n13163) );
  XOR U16460 ( .A(n13166), .B(n13164), .Z(n13165) );
  XNOR U16461 ( .A(n13167), .B(n13168), .Z(n13155) );
  AND U16462 ( .A(n13169), .B(n13170), .Z(n13167) );
  XNOR U16463 ( .A(n13168), .B(n13097), .Z(n13170) );
  XOR U16464 ( .A(n13161), .B(n13162), .Z(n13097) );
  XNOR U16465 ( .A(n13171), .B(n13172), .Z(n13162) );
  ANDN U16466 ( .B(n13173), .A(n13174), .Z(n13171) );
  XOR U16467 ( .A(n13175), .B(n13176), .Z(n13173) );
  XOR U16468 ( .A(n13177), .B(n13178), .Z(n13161) );
  XNOR U16469 ( .A(n13179), .B(n13180), .Z(n13178) );
  ANDN U16470 ( .B(n13181), .A(n13182), .Z(n13179) );
  XNOR U16471 ( .A(n13183), .B(n13184), .Z(n13181) );
  IV U16472 ( .A(n13159), .Z(n13177) );
  XOR U16473 ( .A(n13185), .B(n13186), .Z(n13159) );
  ANDN U16474 ( .B(n13187), .A(n13188), .Z(n13185) );
  XOR U16475 ( .A(n13186), .B(n13189), .Z(n13187) );
  XOR U16476 ( .A(n13168), .B(n13099), .Z(n13169) );
  XOR U16477 ( .A(n13190), .B(n13191), .Z(n13099) );
  AND U16478 ( .A(n66), .B(n13192), .Z(n13190) );
  XOR U16479 ( .A(n13193), .B(n13191), .Z(n13192) );
  XNOR U16480 ( .A(n13194), .B(n13195), .Z(n13168) );
  NAND U16481 ( .A(n13196), .B(n13197), .Z(n13195) );
  XOR U16482 ( .A(n13198), .B(n13147), .Z(n13197) );
  XOR U16483 ( .A(n13188), .B(n13189), .Z(n13147) );
  XOR U16484 ( .A(n13199), .B(n13176), .Z(n13189) );
  XOR U16485 ( .A(n13200), .B(n13201), .Z(n13176) );
  ANDN U16486 ( .B(n13202), .A(n13203), .Z(n13200) );
  XOR U16487 ( .A(n13201), .B(n13204), .Z(n13202) );
  IV U16488 ( .A(n13174), .Z(n13199) );
  XOR U16489 ( .A(n13172), .B(n13205), .Z(n13174) );
  XOR U16490 ( .A(n13206), .B(n13207), .Z(n13205) );
  ANDN U16491 ( .B(n13208), .A(n13209), .Z(n13206) );
  XOR U16492 ( .A(n13210), .B(n13207), .Z(n13208) );
  IV U16493 ( .A(n13175), .Z(n13172) );
  XOR U16494 ( .A(n13211), .B(n13212), .Z(n13175) );
  ANDN U16495 ( .B(n13213), .A(n13214), .Z(n13211) );
  XOR U16496 ( .A(n13212), .B(n13215), .Z(n13213) );
  XOR U16497 ( .A(n13216), .B(n13217), .Z(n13188) );
  XNOR U16498 ( .A(n13183), .B(n13218), .Z(n13217) );
  IV U16499 ( .A(n13186), .Z(n13218) );
  XOR U16500 ( .A(n13219), .B(n13220), .Z(n13186) );
  ANDN U16501 ( .B(n13221), .A(n13222), .Z(n13219) );
  XOR U16502 ( .A(n13220), .B(n13223), .Z(n13221) );
  XNOR U16503 ( .A(n13224), .B(n13225), .Z(n13183) );
  ANDN U16504 ( .B(n13226), .A(n13227), .Z(n13224) );
  XOR U16505 ( .A(n13225), .B(n13228), .Z(n13226) );
  IV U16506 ( .A(n13182), .Z(n13216) );
  XOR U16507 ( .A(n13180), .B(n13229), .Z(n13182) );
  XOR U16508 ( .A(n13230), .B(n13231), .Z(n13229) );
  ANDN U16509 ( .B(n13232), .A(n13233), .Z(n13230) );
  XOR U16510 ( .A(n13234), .B(n13231), .Z(n13232) );
  IV U16511 ( .A(n13184), .Z(n13180) );
  XOR U16512 ( .A(n13235), .B(n13236), .Z(n13184) );
  ANDN U16513 ( .B(n13237), .A(n13238), .Z(n13235) );
  XOR U16514 ( .A(n13239), .B(n13236), .Z(n13237) );
  IV U16515 ( .A(n13194), .Z(n13198) );
  XOR U16516 ( .A(n13194), .B(n13149), .Z(n13196) );
  XOR U16517 ( .A(n13240), .B(n13241), .Z(n13149) );
  AND U16518 ( .A(n66), .B(n13242), .Z(n13240) );
  XOR U16519 ( .A(n13243), .B(n13241), .Z(n13242) );
  NANDN U16520 ( .A(n13151), .B(n13153), .Z(n13194) );
  XOR U16521 ( .A(n13244), .B(n13245), .Z(n13153) );
  AND U16522 ( .A(n66), .B(n13246), .Z(n13244) );
  XOR U16523 ( .A(n13245), .B(n13247), .Z(n13246) );
  XNOR U16524 ( .A(n13248), .B(n13249), .Z(n66) );
  AND U16525 ( .A(n13250), .B(n13251), .Z(n13248) );
  XOR U16526 ( .A(n13249), .B(n13164), .Z(n13251) );
  XNOR U16527 ( .A(n13252), .B(n13253), .Z(n13164) );
  ANDN U16528 ( .B(n13254), .A(n13255), .Z(n13252) );
  XOR U16529 ( .A(n13253), .B(n13256), .Z(n13254) );
  XNOR U16530 ( .A(n13249), .B(n13166), .Z(n13250) );
  XOR U16531 ( .A(n13257), .B(n13258), .Z(n13166) );
  AND U16532 ( .A(n70), .B(n13259), .Z(n13257) );
  XOR U16533 ( .A(n13260), .B(n13258), .Z(n13259) );
  XNOR U16534 ( .A(n13261), .B(n13262), .Z(n13249) );
  AND U16535 ( .A(n13263), .B(n13264), .Z(n13261) );
  XNOR U16536 ( .A(n13262), .B(n13191), .Z(n13264) );
  XOR U16537 ( .A(n13255), .B(n13256), .Z(n13191) );
  XNOR U16538 ( .A(n13265), .B(n13266), .Z(n13256) );
  ANDN U16539 ( .B(n13267), .A(n13268), .Z(n13265) );
  XOR U16540 ( .A(n13269), .B(n13270), .Z(n13267) );
  XOR U16541 ( .A(n13271), .B(n13272), .Z(n13255) );
  XNOR U16542 ( .A(n13273), .B(n13274), .Z(n13272) );
  ANDN U16543 ( .B(n13275), .A(n13276), .Z(n13273) );
  XNOR U16544 ( .A(n13277), .B(n13278), .Z(n13275) );
  IV U16545 ( .A(n13253), .Z(n13271) );
  XOR U16546 ( .A(n13279), .B(n13280), .Z(n13253) );
  ANDN U16547 ( .B(n13281), .A(n13282), .Z(n13279) );
  XOR U16548 ( .A(n13280), .B(n13283), .Z(n13281) );
  XOR U16549 ( .A(n13262), .B(n13193), .Z(n13263) );
  XOR U16550 ( .A(n13284), .B(n13285), .Z(n13193) );
  AND U16551 ( .A(n70), .B(n13286), .Z(n13284) );
  XOR U16552 ( .A(n13287), .B(n13285), .Z(n13286) );
  XNOR U16553 ( .A(n13288), .B(n13289), .Z(n13262) );
  NAND U16554 ( .A(n13290), .B(n13291), .Z(n13289) );
  XOR U16555 ( .A(n13292), .B(n13241), .Z(n13291) );
  XOR U16556 ( .A(n13282), .B(n13283), .Z(n13241) );
  XOR U16557 ( .A(n13293), .B(n13270), .Z(n13283) );
  XOR U16558 ( .A(n13294), .B(n13295), .Z(n13270) );
  ANDN U16559 ( .B(n13296), .A(n13297), .Z(n13294) );
  XOR U16560 ( .A(n13295), .B(n13298), .Z(n13296) );
  IV U16561 ( .A(n13268), .Z(n13293) );
  XOR U16562 ( .A(n13266), .B(n13299), .Z(n13268) );
  XOR U16563 ( .A(n13300), .B(n13301), .Z(n13299) );
  ANDN U16564 ( .B(n13302), .A(n13303), .Z(n13300) );
  XOR U16565 ( .A(n13304), .B(n13301), .Z(n13302) );
  IV U16566 ( .A(n13269), .Z(n13266) );
  XOR U16567 ( .A(n13305), .B(n13306), .Z(n13269) );
  ANDN U16568 ( .B(n13307), .A(n13308), .Z(n13305) );
  XOR U16569 ( .A(n13306), .B(n13309), .Z(n13307) );
  XOR U16570 ( .A(n13310), .B(n13311), .Z(n13282) );
  XNOR U16571 ( .A(n13277), .B(n13312), .Z(n13311) );
  IV U16572 ( .A(n13280), .Z(n13312) );
  XOR U16573 ( .A(n13313), .B(n13314), .Z(n13280) );
  ANDN U16574 ( .B(n13315), .A(n13316), .Z(n13313) );
  XOR U16575 ( .A(n13314), .B(n13317), .Z(n13315) );
  XNOR U16576 ( .A(n13318), .B(n13319), .Z(n13277) );
  ANDN U16577 ( .B(n13320), .A(n13321), .Z(n13318) );
  XOR U16578 ( .A(n13319), .B(n13322), .Z(n13320) );
  IV U16579 ( .A(n13276), .Z(n13310) );
  XOR U16580 ( .A(n13274), .B(n13323), .Z(n13276) );
  XOR U16581 ( .A(n13324), .B(n13325), .Z(n13323) );
  ANDN U16582 ( .B(n13326), .A(n13327), .Z(n13324) );
  XOR U16583 ( .A(n13328), .B(n13325), .Z(n13326) );
  IV U16584 ( .A(n13278), .Z(n13274) );
  XOR U16585 ( .A(n13329), .B(n13330), .Z(n13278) );
  ANDN U16586 ( .B(n13331), .A(n13332), .Z(n13329) );
  XOR U16587 ( .A(n13333), .B(n13330), .Z(n13331) );
  IV U16588 ( .A(n13288), .Z(n13292) );
  XOR U16589 ( .A(n13288), .B(n13243), .Z(n13290) );
  XOR U16590 ( .A(n13334), .B(n13335), .Z(n13243) );
  AND U16591 ( .A(n70), .B(n13336), .Z(n13334) );
  XOR U16592 ( .A(n13337), .B(n13335), .Z(n13336) );
  NANDN U16593 ( .A(n13245), .B(n13247), .Z(n13288) );
  XOR U16594 ( .A(n13338), .B(n13339), .Z(n13247) );
  AND U16595 ( .A(n70), .B(n13340), .Z(n13338) );
  XOR U16596 ( .A(n13339), .B(n13341), .Z(n13340) );
  XNOR U16597 ( .A(n13342), .B(n13343), .Z(n70) );
  AND U16598 ( .A(n13344), .B(n13345), .Z(n13342) );
  XOR U16599 ( .A(n13343), .B(n13258), .Z(n13345) );
  XNOR U16600 ( .A(n13346), .B(n13347), .Z(n13258) );
  ANDN U16601 ( .B(n13348), .A(n13349), .Z(n13346) );
  XOR U16602 ( .A(n13347), .B(n13350), .Z(n13348) );
  XNOR U16603 ( .A(n13343), .B(n13260), .Z(n13344) );
  XOR U16604 ( .A(n13351), .B(n13352), .Z(n13260) );
  AND U16605 ( .A(n74), .B(n13353), .Z(n13351) );
  XOR U16606 ( .A(n13354), .B(n13352), .Z(n13353) );
  XNOR U16607 ( .A(n13355), .B(n13356), .Z(n13343) );
  AND U16608 ( .A(n13357), .B(n13358), .Z(n13355) );
  XNOR U16609 ( .A(n13356), .B(n13285), .Z(n13358) );
  XOR U16610 ( .A(n13349), .B(n13350), .Z(n13285) );
  XNOR U16611 ( .A(n13359), .B(n13360), .Z(n13350) );
  ANDN U16612 ( .B(n13361), .A(n13362), .Z(n13359) );
  XOR U16613 ( .A(n13363), .B(n13364), .Z(n13361) );
  XOR U16614 ( .A(n13365), .B(n13366), .Z(n13349) );
  XNOR U16615 ( .A(n13367), .B(n13368), .Z(n13366) );
  ANDN U16616 ( .B(n13369), .A(n13370), .Z(n13367) );
  XNOR U16617 ( .A(n13371), .B(n13372), .Z(n13369) );
  IV U16618 ( .A(n13347), .Z(n13365) );
  XOR U16619 ( .A(n13373), .B(n13374), .Z(n13347) );
  ANDN U16620 ( .B(n13375), .A(n13376), .Z(n13373) );
  XOR U16621 ( .A(n13374), .B(n13377), .Z(n13375) );
  XOR U16622 ( .A(n13356), .B(n13287), .Z(n13357) );
  XOR U16623 ( .A(n13378), .B(n13379), .Z(n13287) );
  AND U16624 ( .A(n74), .B(n13380), .Z(n13378) );
  XOR U16625 ( .A(n13381), .B(n13379), .Z(n13380) );
  XNOR U16626 ( .A(n13382), .B(n13383), .Z(n13356) );
  NAND U16627 ( .A(n13384), .B(n13385), .Z(n13383) );
  XOR U16628 ( .A(n13386), .B(n13335), .Z(n13385) );
  XOR U16629 ( .A(n13376), .B(n13377), .Z(n13335) );
  XOR U16630 ( .A(n13387), .B(n13364), .Z(n13377) );
  XOR U16631 ( .A(n13388), .B(n13389), .Z(n13364) );
  ANDN U16632 ( .B(n13390), .A(n13391), .Z(n13388) );
  XOR U16633 ( .A(n13389), .B(n13392), .Z(n13390) );
  IV U16634 ( .A(n13362), .Z(n13387) );
  XOR U16635 ( .A(n13360), .B(n13393), .Z(n13362) );
  XOR U16636 ( .A(n13394), .B(n13395), .Z(n13393) );
  ANDN U16637 ( .B(n13396), .A(n13397), .Z(n13394) );
  XOR U16638 ( .A(n13398), .B(n13395), .Z(n13396) );
  IV U16639 ( .A(n13363), .Z(n13360) );
  XOR U16640 ( .A(n13399), .B(n13400), .Z(n13363) );
  ANDN U16641 ( .B(n13401), .A(n13402), .Z(n13399) );
  XOR U16642 ( .A(n13400), .B(n13403), .Z(n13401) );
  XOR U16643 ( .A(n13404), .B(n13405), .Z(n13376) );
  XNOR U16644 ( .A(n13371), .B(n13406), .Z(n13405) );
  IV U16645 ( .A(n13374), .Z(n13406) );
  XOR U16646 ( .A(n13407), .B(n13408), .Z(n13374) );
  ANDN U16647 ( .B(n13409), .A(n13410), .Z(n13407) );
  XOR U16648 ( .A(n13408), .B(n13411), .Z(n13409) );
  XNOR U16649 ( .A(n13412), .B(n13413), .Z(n13371) );
  ANDN U16650 ( .B(n13414), .A(n13415), .Z(n13412) );
  XOR U16651 ( .A(n13413), .B(n13416), .Z(n13414) );
  IV U16652 ( .A(n13370), .Z(n13404) );
  XOR U16653 ( .A(n13368), .B(n13417), .Z(n13370) );
  XOR U16654 ( .A(n13418), .B(n13419), .Z(n13417) );
  ANDN U16655 ( .B(n13420), .A(n13421), .Z(n13418) );
  XOR U16656 ( .A(n13422), .B(n13419), .Z(n13420) );
  IV U16657 ( .A(n13372), .Z(n13368) );
  XOR U16658 ( .A(n13423), .B(n13424), .Z(n13372) );
  ANDN U16659 ( .B(n13425), .A(n13426), .Z(n13423) );
  XOR U16660 ( .A(n13427), .B(n13424), .Z(n13425) );
  IV U16661 ( .A(n13382), .Z(n13386) );
  XOR U16662 ( .A(n13382), .B(n13337), .Z(n13384) );
  XOR U16663 ( .A(n13428), .B(n13429), .Z(n13337) );
  AND U16664 ( .A(n74), .B(n13430), .Z(n13428) );
  XOR U16665 ( .A(n13431), .B(n13429), .Z(n13430) );
  NANDN U16666 ( .A(n13339), .B(n13341), .Z(n13382) );
  XOR U16667 ( .A(n13432), .B(n13433), .Z(n13341) );
  AND U16668 ( .A(n74), .B(n13434), .Z(n13432) );
  XOR U16669 ( .A(n13433), .B(n13435), .Z(n13434) );
  XNOR U16670 ( .A(n13436), .B(n13437), .Z(n74) );
  AND U16671 ( .A(n13438), .B(n13439), .Z(n13436) );
  XOR U16672 ( .A(n13437), .B(n13352), .Z(n13439) );
  XNOR U16673 ( .A(n13440), .B(n13441), .Z(n13352) );
  ANDN U16674 ( .B(n13442), .A(n13443), .Z(n13440) );
  XOR U16675 ( .A(n13441), .B(n13444), .Z(n13442) );
  XNOR U16676 ( .A(n13437), .B(n13354), .Z(n13438) );
  XOR U16677 ( .A(n13445), .B(n13446), .Z(n13354) );
  AND U16678 ( .A(n78), .B(n13447), .Z(n13445) );
  XOR U16679 ( .A(n13448), .B(n13446), .Z(n13447) );
  XNOR U16680 ( .A(n13449), .B(n13450), .Z(n13437) );
  AND U16681 ( .A(n13451), .B(n13452), .Z(n13449) );
  XNOR U16682 ( .A(n13450), .B(n13379), .Z(n13452) );
  XOR U16683 ( .A(n13443), .B(n13444), .Z(n13379) );
  XNOR U16684 ( .A(n13453), .B(n13454), .Z(n13444) );
  ANDN U16685 ( .B(n13455), .A(n13456), .Z(n13453) );
  XOR U16686 ( .A(n13457), .B(n13458), .Z(n13455) );
  XOR U16687 ( .A(n13459), .B(n13460), .Z(n13443) );
  XNOR U16688 ( .A(n13461), .B(n13462), .Z(n13460) );
  ANDN U16689 ( .B(n13463), .A(n13464), .Z(n13461) );
  XNOR U16690 ( .A(n13465), .B(n13466), .Z(n13463) );
  IV U16691 ( .A(n13441), .Z(n13459) );
  XOR U16692 ( .A(n13467), .B(n13468), .Z(n13441) );
  ANDN U16693 ( .B(n13469), .A(n13470), .Z(n13467) );
  XOR U16694 ( .A(n13468), .B(n13471), .Z(n13469) );
  XOR U16695 ( .A(n13450), .B(n13381), .Z(n13451) );
  XOR U16696 ( .A(n13472), .B(n13473), .Z(n13381) );
  AND U16697 ( .A(n78), .B(n13474), .Z(n13472) );
  XOR U16698 ( .A(n13475), .B(n13473), .Z(n13474) );
  XNOR U16699 ( .A(n13476), .B(n13477), .Z(n13450) );
  NAND U16700 ( .A(n13478), .B(n13479), .Z(n13477) );
  XOR U16701 ( .A(n13480), .B(n13429), .Z(n13479) );
  XOR U16702 ( .A(n13470), .B(n13471), .Z(n13429) );
  XOR U16703 ( .A(n13481), .B(n13458), .Z(n13471) );
  XOR U16704 ( .A(n13482), .B(n13483), .Z(n13458) );
  ANDN U16705 ( .B(n13484), .A(n13485), .Z(n13482) );
  XOR U16706 ( .A(n13483), .B(n13486), .Z(n13484) );
  IV U16707 ( .A(n13456), .Z(n13481) );
  XOR U16708 ( .A(n13454), .B(n13487), .Z(n13456) );
  XOR U16709 ( .A(n13488), .B(n13489), .Z(n13487) );
  ANDN U16710 ( .B(n13490), .A(n13491), .Z(n13488) );
  XOR U16711 ( .A(n13492), .B(n13489), .Z(n13490) );
  IV U16712 ( .A(n13457), .Z(n13454) );
  XOR U16713 ( .A(n13493), .B(n13494), .Z(n13457) );
  ANDN U16714 ( .B(n13495), .A(n13496), .Z(n13493) );
  XOR U16715 ( .A(n13494), .B(n13497), .Z(n13495) );
  XOR U16716 ( .A(n13498), .B(n13499), .Z(n13470) );
  XNOR U16717 ( .A(n13465), .B(n13500), .Z(n13499) );
  IV U16718 ( .A(n13468), .Z(n13500) );
  XOR U16719 ( .A(n13501), .B(n13502), .Z(n13468) );
  ANDN U16720 ( .B(n13503), .A(n13504), .Z(n13501) );
  XOR U16721 ( .A(n13502), .B(n13505), .Z(n13503) );
  XNOR U16722 ( .A(n13506), .B(n13507), .Z(n13465) );
  ANDN U16723 ( .B(n13508), .A(n13509), .Z(n13506) );
  XOR U16724 ( .A(n13507), .B(n13510), .Z(n13508) );
  IV U16725 ( .A(n13464), .Z(n13498) );
  XOR U16726 ( .A(n13462), .B(n13511), .Z(n13464) );
  XOR U16727 ( .A(n13512), .B(n13513), .Z(n13511) );
  ANDN U16728 ( .B(n13514), .A(n13515), .Z(n13512) );
  XOR U16729 ( .A(n13516), .B(n13513), .Z(n13514) );
  IV U16730 ( .A(n13466), .Z(n13462) );
  XOR U16731 ( .A(n13517), .B(n13518), .Z(n13466) );
  ANDN U16732 ( .B(n13519), .A(n13520), .Z(n13517) );
  XOR U16733 ( .A(n13521), .B(n13518), .Z(n13519) );
  IV U16734 ( .A(n13476), .Z(n13480) );
  XOR U16735 ( .A(n13476), .B(n13431), .Z(n13478) );
  XOR U16736 ( .A(n13522), .B(n13523), .Z(n13431) );
  AND U16737 ( .A(n78), .B(n13524), .Z(n13522) );
  XOR U16738 ( .A(n13525), .B(n13523), .Z(n13524) );
  NANDN U16739 ( .A(n13433), .B(n13435), .Z(n13476) );
  XOR U16740 ( .A(n13526), .B(n13527), .Z(n13435) );
  AND U16741 ( .A(n78), .B(n13528), .Z(n13526) );
  XOR U16742 ( .A(n13527), .B(n13529), .Z(n13528) );
  XNOR U16743 ( .A(n13530), .B(n13531), .Z(n78) );
  AND U16744 ( .A(n13532), .B(n13533), .Z(n13530) );
  XOR U16745 ( .A(n13531), .B(n13446), .Z(n13533) );
  XNOR U16746 ( .A(n13534), .B(n13535), .Z(n13446) );
  ANDN U16747 ( .B(n13536), .A(n13537), .Z(n13534) );
  XOR U16748 ( .A(n13535), .B(n13538), .Z(n13536) );
  XNOR U16749 ( .A(n13531), .B(n13448), .Z(n13532) );
  XOR U16750 ( .A(n13539), .B(n13540), .Z(n13448) );
  AND U16751 ( .A(n82), .B(n13541), .Z(n13539) );
  XOR U16752 ( .A(n13542), .B(n13540), .Z(n13541) );
  XNOR U16753 ( .A(n13543), .B(n13544), .Z(n13531) );
  AND U16754 ( .A(n13545), .B(n13546), .Z(n13543) );
  XNOR U16755 ( .A(n13544), .B(n13473), .Z(n13546) );
  XOR U16756 ( .A(n13537), .B(n13538), .Z(n13473) );
  XNOR U16757 ( .A(n13547), .B(n13548), .Z(n13538) );
  ANDN U16758 ( .B(n13549), .A(n13550), .Z(n13547) );
  XOR U16759 ( .A(n13551), .B(n13552), .Z(n13549) );
  XOR U16760 ( .A(n13553), .B(n13554), .Z(n13537) );
  XNOR U16761 ( .A(n13555), .B(n13556), .Z(n13554) );
  ANDN U16762 ( .B(n13557), .A(n13558), .Z(n13555) );
  XNOR U16763 ( .A(n13559), .B(n13560), .Z(n13557) );
  IV U16764 ( .A(n13535), .Z(n13553) );
  XOR U16765 ( .A(n13561), .B(n13562), .Z(n13535) );
  ANDN U16766 ( .B(n13563), .A(n13564), .Z(n13561) );
  XOR U16767 ( .A(n13562), .B(n13565), .Z(n13563) );
  XOR U16768 ( .A(n13544), .B(n13475), .Z(n13545) );
  XOR U16769 ( .A(n13566), .B(n13567), .Z(n13475) );
  AND U16770 ( .A(n82), .B(n13568), .Z(n13566) );
  XOR U16771 ( .A(n13569), .B(n13567), .Z(n13568) );
  XNOR U16772 ( .A(n13570), .B(n13571), .Z(n13544) );
  NAND U16773 ( .A(n13572), .B(n13573), .Z(n13571) );
  XOR U16774 ( .A(n13574), .B(n13523), .Z(n13573) );
  XOR U16775 ( .A(n13564), .B(n13565), .Z(n13523) );
  XOR U16776 ( .A(n13575), .B(n13552), .Z(n13565) );
  XOR U16777 ( .A(n13576), .B(n13577), .Z(n13552) );
  ANDN U16778 ( .B(n13578), .A(n13579), .Z(n13576) );
  XOR U16779 ( .A(n13577), .B(n13580), .Z(n13578) );
  IV U16780 ( .A(n13550), .Z(n13575) );
  XOR U16781 ( .A(n13548), .B(n13581), .Z(n13550) );
  XOR U16782 ( .A(n13582), .B(n13583), .Z(n13581) );
  ANDN U16783 ( .B(n13584), .A(n13585), .Z(n13582) );
  XOR U16784 ( .A(n13586), .B(n13583), .Z(n13584) );
  IV U16785 ( .A(n13551), .Z(n13548) );
  XOR U16786 ( .A(n13587), .B(n13588), .Z(n13551) );
  ANDN U16787 ( .B(n13589), .A(n13590), .Z(n13587) );
  XOR U16788 ( .A(n13588), .B(n13591), .Z(n13589) );
  XOR U16789 ( .A(n13592), .B(n13593), .Z(n13564) );
  XNOR U16790 ( .A(n13559), .B(n13594), .Z(n13593) );
  IV U16791 ( .A(n13562), .Z(n13594) );
  XOR U16792 ( .A(n13595), .B(n13596), .Z(n13562) );
  ANDN U16793 ( .B(n13597), .A(n13598), .Z(n13595) );
  XOR U16794 ( .A(n13596), .B(n13599), .Z(n13597) );
  XNOR U16795 ( .A(n13600), .B(n13601), .Z(n13559) );
  ANDN U16796 ( .B(n13602), .A(n13603), .Z(n13600) );
  XOR U16797 ( .A(n13601), .B(n13604), .Z(n13602) );
  IV U16798 ( .A(n13558), .Z(n13592) );
  XOR U16799 ( .A(n13556), .B(n13605), .Z(n13558) );
  XOR U16800 ( .A(n13606), .B(n13607), .Z(n13605) );
  ANDN U16801 ( .B(n13608), .A(n13609), .Z(n13606) );
  XOR U16802 ( .A(n13610), .B(n13607), .Z(n13608) );
  IV U16803 ( .A(n13560), .Z(n13556) );
  XOR U16804 ( .A(n13611), .B(n13612), .Z(n13560) );
  ANDN U16805 ( .B(n13613), .A(n13614), .Z(n13611) );
  XOR U16806 ( .A(n13615), .B(n13612), .Z(n13613) );
  IV U16807 ( .A(n13570), .Z(n13574) );
  XOR U16808 ( .A(n13570), .B(n13525), .Z(n13572) );
  XOR U16809 ( .A(n13616), .B(n13617), .Z(n13525) );
  AND U16810 ( .A(n82), .B(n13618), .Z(n13616) );
  XOR U16811 ( .A(n13619), .B(n13617), .Z(n13618) );
  NANDN U16812 ( .A(n13527), .B(n13529), .Z(n13570) );
  XOR U16813 ( .A(n13620), .B(n13621), .Z(n13529) );
  AND U16814 ( .A(n82), .B(n13622), .Z(n13620) );
  XOR U16815 ( .A(n13621), .B(n13623), .Z(n13622) );
  XNOR U16816 ( .A(n13624), .B(n13625), .Z(n82) );
  AND U16817 ( .A(n13626), .B(n13627), .Z(n13624) );
  XOR U16818 ( .A(n13625), .B(n13540), .Z(n13627) );
  XNOR U16819 ( .A(n13628), .B(n13629), .Z(n13540) );
  ANDN U16820 ( .B(n13630), .A(n13631), .Z(n13628) );
  XOR U16821 ( .A(n13629), .B(n13632), .Z(n13630) );
  XNOR U16822 ( .A(n13625), .B(n13542), .Z(n13626) );
  XOR U16823 ( .A(n13633), .B(n13634), .Z(n13542) );
  AND U16824 ( .A(n86), .B(n13635), .Z(n13633) );
  XOR U16825 ( .A(n13636), .B(n13634), .Z(n13635) );
  XNOR U16826 ( .A(n13637), .B(n13638), .Z(n13625) );
  AND U16827 ( .A(n13639), .B(n13640), .Z(n13637) );
  XNOR U16828 ( .A(n13638), .B(n13567), .Z(n13640) );
  XOR U16829 ( .A(n13631), .B(n13632), .Z(n13567) );
  XNOR U16830 ( .A(n13641), .B(n13642), .Z(n13632) );
  ANDN U16831 ( .B(n13643), .A(n13644), .Z(n13641) );
  XOR U16832 ( .A(n13645), .B(n13646), .Z(n13643) );
  XOR U16833 ( .A(n13647), .B(n13648), .Z(n13631) );
  XNOR U16834 ( .A(n13649), .B(n13650), .Z(n13648) );
  ANDN U16835 ( .B(n13651), .A(n13652), .Z(n13649) );
  XNOR U16836 ( .A(n13653), .B(n13654), .Z(n13651) );
  IV U16837 ( .A(n13629), .Z(n13647) );
  XOR U16838 ( .A(n13655), .B(n13656), .Z(n13629) );
  ANDN U16839 ( .B(n13657), .A(n13658), .Z(n13655) );
  XOR U16840 ( .A(n13656), .B(n13659), .Z(n13657) );
  XOR U16841 ( .A(n13638), .B(n13569), .Z(n13639) );
  XOR U16842 ( .A(n13660), .B(n13661), .Z(n13569) );
  AND U16843 ( .A(n86), .B(n13662), .Z(n13660) );
  XOR U16844 ( .A(n13663), .B(n13661), .Z(n13662) );
  XNOR U16845 ( .A(n13664), .B(n13665), .Z(n13638) );
  NAND U16846 ( .A(n13666), .B(n13667), .Z(n13665) );
  XOR U16847 ( .A(n13668), .B(n13617), .Z(n13667) );
  XOR U16848 ( .A(n13658), .B(n13659), .Z(n13617) );
  XOR U16849 ( .A(n13669), .B(n13646), .Z(n13659) );
  XOR U16850 ( .A(n13670), .B(n13671), .Z(n13646) );
  ANDN U16851 ( .B(n13672), .A(n13673), .Z(n13670) );
  XOR U16852 ( .A(n13671), .B(n13674), .Z(n13672) );
  IV U16853 ( .A(n13644), .Z(n13669) );
  XOR U16854 ( .A(n13642), .B(n13675), .Z(n13644) );
  XOR U16855 ( .A(n13676), .B(n13677), .Z(n13675) );
  ANDN U16856 ( .B(n13678), .A(n13679), .Z(n13676) );
  XOR U16857 ( .A(n13680), .B(n13677), .Z(n13678) );
  IV U16858 ( .A(n13645), .Z(n13642) );
  XOR U16859 ( .A(n13681), .B(n13682), .Z(n13645) );
  ANDN U16860 ( .B(n13683), .A(n13684), .Z(n13681) );
  XOR U16861 ( .A(n13682), .B(n13685), .Z(n13683) );
  XOR U16862 ( .A(n13686), .B(n13687), .Z(n13658) );
  XNOR U16863 ( .A(n13653), .B(n13688), .Z(n13687) );
  IV U16864 ( .A(n13656), .Z(n13688) );
  XOR U16865 ( .A(n13689), .B(n13690), .Z(n13656) );
  ANDN U16866 ( .B(n13691), .A(n13692), .Z(n13689) );
  XOR U16867 ( .A(n13690), .B(n13693), .Z(n13691) );
  XNOR U16868 ( .A(n13694), .B(n13695), .Z(n13653) );
  ANDN U16869 ( .B(n13696), .A(n13697), .Z(n13694) );
  XOR U16870 ( .A(n13695), .B(n13698), .Z(n13696) );
  IV U16871 ( .A(n13652), .Z(n13686) );
  XOR U16872 ( .A(n13650), .B(n13699), .Z(n13652) );
  XOR U16873 ( .A(n13700), .B(n13701), .Z(n13699) );
  ANDN U16874 ( .B(n13702), .A(n13703), .Z(n13700) );
  XOR U16875 ( .A(n13704), .B(n13701), .Z(n13702) );
  IV U16876 ( .A(n13654), .Z(n13650) );
  XOR U16877 ( .A(n13705), .B(n13706), .Z(n13654) );
  ANDN U16878 ( .B(n13707), .A(n13708), .Z(n13705) );
  XOR U16879 ( .A(n13709), .B(n13706), .Z(n13707) );
  IV U16880 ( .A(n13664), .Z(n13668) );
  XOR U16881 ( .A(n13664), .B(n13619), .Z(n13666) );
  XOR U16882 ( .A(n13710), .B(n13711), .Z(n13619) );
  AND U16883 ( .A(n86), .B(n13712), .Z(n13710) );
  XOR U16884 ( .A(n13713), .B(n13711), .Z(n13712) );
  NANDN U16885 ( .A(n13621), .B(n13623), .Z(n13664) );
  XOR U16886 ( .A(n13714), .B(n13715), .Z(n13623) );
  AND U16887 ( .A(n86), .B(n13716), .Z(n13714) );
  XOR U16888 ( .A(n13715), .B(n13717), .Z(n13716) );
  XNOR U16889 ( .A(n13718), .B(n13719), .Z(n86) );
  AND U16890 ( .A(n13720), .B(n13721), .Z(n13718) );
  XOR U16891 ( .A(n13719), .B(n13634), .Z(n13721) );
  XNOR U16892 ( .A(n13722), .B(n13723), .Z(n13634) );
  ANDN U16893 ( .B(n13724), .A(n13725), .Z(n13722) );
  XOR U16894 ( .A(n13723), .B(n13726), .Z(n13724) );
  XNOR U16895 ( .A(n13719), .B(n13636), .Z(n13720) );
  XOR U16896 ( .A(n13727), .B(n13728), .Z(n13636) );
  AND U16897 ( .A(n90), .B(n13729), .Z(n13727) );
  XOR U16898 ( .A(n13730), .B(n13728), .Z(n13729) );
  XNOR U16899 ( .A(n13731), .B(n13732), .Z(n13719) );
  AND U16900 ( .A(n13733), .B(n13734), .Z(n13731) );
  XNOR U16901 ( .A(n13732), .B(n13661), .Z(n13734) );
  XOR U16902 ( .A(n13725), .B(n13726), .Z(n13661) );
  XNOR U16903 ( .A(n13735), .B(n13736), .Z(n13726) );
  ANDN U16904 ( .B(n13737), .A(n13738), .Z(n13735) );
  XOR U16905 ( .A(n13739), .B(n13740), .Z(n13737) );
  XOR U16906 ( .A(n13741), .B(n13742), .Z(n13725) );
  XNOR U16907 ( .A(n13743), .B(n13744), .Z(n13742) );
  ANDN U16908 ( .B(n13745), .A(n13746), .Z(n13743) );
  XNOR U16909 ( .A(n13747), .B(n13748), .Z(n13745) );
  IV U16910 ( .A(n13723), .Z(n13741) );
  XOR U16911 ( .A(n13749), .B(n13750), .Z(n13723) );
  ANDN U16912 ( .B(n13751), .A(n13752), .Z(n13749) );
  XOR U16913 ( .A(n13750), .B(n13753), .Z(n13751) );
  XOR U16914 ( .A(n13732), .B(n13663), .Z(n13733) );
  XOR U16915 ( .A(n13754), .B(n13755), .Z(n13663) );
  AND U16916 ( .A(n90), .B(n13756), .Z(n13754) );
  XOR U16917 ( .A(n13757), .B(n13755), .Z(n13756) );
  XNOR U16918 ( .A(n13758), .B(n13759), .Z(n13732) );
  NAND U16919 ( .A(n13760), .B(n13761), .Z(n13759) );
  XOR U16920 ( .A(n13762), .B(n13711), .Z(n13761) );
  XOR U16921 ( .A(n13752), .B(n13753), .Z(n13711) );
  XOR U16922 ( .A(n13763), .B(n13740), .Z(n13753) );
  XOR U16923 ( .A(n13764), .B(n13765), .Z(n13740) );
  ANDN U16924 ( .B(n13766), .A(n13767), .Z(n13764) );
  XOR U16925 ( .A(n13765), .B(n13768), .Z(n13766) );
  IV U16926 ( .A(n13738), .Z(n13763) );
  XOR U16927 ( .A(n13736), .B(n13769), .Z(n13738) );
  XOR U16928 ( .A(n13770), .B(n13771), .Z(n13769) );
  ANDN U16929 ( .B(n13772), .A(n13773), .Z(n13770) );
  XOR U16930 ( .A(n13774), .B(n13771), .Z(n13772) );
  IV U16931 ( .A(n13739), .Z(n13736) );
  XOR U16932 ( .A(n13775), .B(n13776), .Z(n13739) );
  ANDN U16933 ( .B(n13777), .A(n13778), .Z(n13775) );
  XOR U16934 ( .A(n13776), .B(n13779), .Z(n13777) );
  XOR U16935 ( .A(n13780), .B(n13781), .Z(n13752) );
  XNOR U16936 ( .A(n13747), .B(n13782), .Z(n13781) );
  IV U16937 ( .A(n13750), .Z(n13782) );
  XOR U16938 ( .A(n13783), .B(n13784), .Z(n13750) );
  ANDN U16939 ( .B(n13785), .A(n13786), .Z(n13783) );
  XOR U16940 ( .A(n13784), .B(n13787), .Z(n13785) );
  XNOR U16941 ( .A(n13788), .B(n13789), .Z(n13747) );
  ANDN U16942 ( .B(n13790), .A(n13791), .Z(n13788) );
  XOR U16943 ( .A(n13789), .B(n13792), .Z(n13790) );
  IV U16944 ( .A(n13746), .Z(n13780) );
  XOR U16945 ( .A(n13744), .B(n13793), .Z(n13746) );
  XOR U16946 ( .A(n13794), .B(n13795), .Z(n13793) );
  ANDN U16947 ( .B(n13796), .A(n13797), .Z(n13794) );
  XOR U16948 ( .A(n13798), .B(n13795), .Z(n13796) );
  IV U16949 ( .A(n13748), .Z(n13744) );
  XOR U16950 ( .A(n13799), .B(n13800), .Z(n13748) );
  ANDN U16951 ( .B(n13801), .A(n13802), .Z(n13799) );
  XOR U16952 ( .A(n13803), .B(n13800), .Z(n13801) );
  IV U16953 ( .A(n13758), .Z(n13762) );
  XOR U16954 ( .A(n13758), .B(n13713), .Z(n13760) );
  XOR U16955 ( .A(n13804), .B(n13805), .Z(n13713) );
  AND U16956 ( .A(n90), .B(n13806), .Z(n13804) );
  XOR U16957 ( .A(n13807), .B(n13805), .Z(n13806) );
  NANDN U16958 ( .A(n13715), .B(n13717), .Z(n13758) );
  XOR U16959 ( .A(n13808), .B(n13809), .Z(n13717) );
  AND U16960 ( .A(n90), .B(n13810), .Z(n13808) );
  XOR U16961 ( .A(n13809), .B(n13811), .Z(n13810) );
  XNOR U16962 ( .A(n13812), .B(n13813), .Z(n90) );
  AND U16963 ( .A(n13814), .B(n13815), .Z(n13812) );
  XOR U16964 ( .A(n13813), .B(n13728), .Z(n13815) );
  XNOR U16965 ( .A(n13816), .B(n13817), .Z(n13728) );
  ANDN U16966 ( .B(n13818), .A(n13819), .Z(n13816) );
  XOR U16967 ( .A(n13817), .B(n13820), .Z(n13818) );
  XNOR U16968 ( .A(n13813), .B(n13730), .Z(n13814) );
  XOR U16969 ( .A(n13821), .B(n13822), .Z(n13730) );
  AND U16970 ( .A(n94), .B(n13823), .Z(n13821) );
  XOR U16971 ( .A(n13824), .B(n13822), .Z(n13823) );
  XNOR U16972 ( .A(n13825), .B(n13826), .Z(n13813) );
  AND U16973 ( .A(n13827), .B(n13828), .Z(n13825) );
  XNOR U16974 ( .A(n13826), .B(n13755), .Z(n13828) );
  XOR U16975 ( .A(n13819), .B(n13820), .Z(n13755) );
  XNOR U16976 ( .A(n13829), .B(n13830), .Z(n13820) );
  ANDN U16977 ( .B(n13831), .A(n13832), .Z(n13829) );
  XOR U16978 ( .A(n13833), .B(n13834), .Z(n13831) );
  XOR U16979 ( .A(n13835), .B(n13836), .Z(n13819) );
  XNOR U16980 ( .A(n13837), .B(n13838), .Z(n13836) );
  ANDN U16981 ( .B(n13839), .A(n13840), .Z(n13837) );
  XNOR U16982 ( .A(n13841), .B(n13842), .Z(n13839) );
  IV U16983 ( .A(n13817), .Z(n13835) );
  XOR U16984 ( .A(n13843), .B(n13844), .Z(n13817) );
  ANDN U16985 ( .B(n13845), .A(n13846), .Z(n13843) );
  XOR U16986 ( .A(n13844), .B(n13847), .Z(n13845) );
  XOR U16987 ( .A(n13826), .B(n13757), .Z(n13827) );
  XOR U16988 ( .A(n13848), .B(n13849), .Z(n13757) );
  AND U16989 ( .A(n94), .B(n13850), .Z(n13848) );
  XOR U16990 ( .A(n13851), .B(n13849), .Z(n13850) );
  XNOR U16991 ( .A(n13852), .B(n13853), .Z(n13826) );
  NAND U16992 ( .A(n13854), .B(n13855), .Z(n13853) );
  XOR U16993 ( .A(n13856), .B(n13805), .Z(n13855) );
  XOR U16994 ( .A(n13846), .B(n13847), .Z(n13805) );
  XOR U16995 ( .A(n13857), .B(n13834), .Z(n13847) );
  XOR U16996 ( .A(n13858), .B(n13859), .Z(n13834) );
  ANDN U16997 ( .B(n13860), .A(n13861), .Z(n13858) );
  XOR U16998 ( .A(n13859), .B(n13862), .Z(n13860) );
  IV U16999 ( .A(n13832), .Z(n13857) );
  XOR U17000 ( .A(n13830), .B(n13863), .Z(n13832) );
  XOR U17001 ( .A(n13864), .B(n13865), .Z(n13863) );
  ANDN U17002 ( .B(n13866), .A(n13867), .Z(n13864) );
  XOR U17003 ( .A(n13868), .B(n13865), .Z(n13866) );
  IV U17004 ( .A(n13833), .Z(n13830) );
  XOR U17005 ( .A(n13869), .B(n13870), .Z(n13833) );
  ANDN U17006 ( .B(n13871), .A(n13872), .Z(n13869) );
  XOR U17007 ( .A(n13870), .B(n13873), .Z(n13871) );
  XOR U17008 ( .A(n13874), .B(n13875), .Z(n13846) );
  XNOR U17009 ( .A(n13841), .B(n13876), .Z(n13875) );
  IV U17010 ( .A(n13844), .Z(n13876) );
  XOR U17011 ( .A(n13877), .B(n13878), .Z(n13844) );
  ANDN U17012 ( .B(n13879), .A(n13880), .Z(n13877) );
  XOR U17013 ( .A(n13878), .B(n13881), .Z(n13879) );
  XNOR U17014 ( .A(n13882), .B(n13883), .Z(n13841) );
  ANDN U17015 ( .B(n13884), .A(n13885), .Z(n13882) );
  XOR U17016 ( .A(n13883), .B(n13886), .Z(n13884) );
  IV U17017 ( .A(n13840), .Z(n13874) );
  XOR U17018 ( .A(n13838), .B(n13887), .Z(n13840) );
  XOR U17019 ( .A(n13888), .B(n13889), .Z(n13887) );
  ANDN U17020 ( .B(n13890), .A(n13891), .Z(n13888) );
  XOR U17021 ( .A(n13892), .B(n13889), .Z(n13890) );
  IV U17022 ( .A(n13842), .Z(n13838) );
  XOR U17023 ( .A(n13893), .B(n13894), .Z(n13842) );
  ANDN U17024 ( .B(n13895), .A(n13896), .Z(n13893) );
  XOR U17025 ( .A(n13897), .B(n13894), .Z(n13895) );
  IV U17026 ( .A(n13852), .Z(n13856) );
  XOR U17027 ( .A(n13852), .B(n13807), .Z(n13854) );
  XOR U17028 ( .A(n13898), .B(n13899), .Z(n13807) );
  AND U17029 ( .A(n94), .B(n13900), .Z(n13898) );
  XOR U17030 ( .A(n13901), .B(n13899), .Z(n13900) );
  NANDN U17031 ( .A(n13809), .B(n13811), .Z(n13852) );
  XOR U17032 ( .A(n13902), .B(n13903), .Z(n13811) );
  AND U17033 ( .A(n94), .B(n13904), .Z(n13902) );
  XOR U17034 ( .A(n13903), .B(n13905), .Z(n13904) );
  XNOR U17035 ( .A(n13906), .B(n13907), .Z(n94) );
  AND U17036 ( .A(n13908), .B(n13909), .Z(n13906) );
  XOR U17037 ( .A(n13907), .B(n13822), .Z(n13909) );
  XNOR U17038 ( .A(n13910), .B(n13911), .Z(n13822) );
  ANDN U17039 ( .B(n13912), .A(n13913), .Z(n13910) );
  XOR U17040 ( .A(n13911), .B(n13914), .Z(n13912) );
  XNOR U17041 ( .A(n13907), .B(n13824), .Z(n13908) );
  XOR U17042 ( .A(n13915), .B(n13916), .Z(n13824) );
  AND U17043 ( .A(n98), .B(n13917), .Z(n13915) );
  XOR U17044 ( .A(n13918), .B(n13916), .Z(n13917) );
  XNOR U17045 ( .A(n13919), .B(n13920), .Z(n13907) );
  AND U17046 ( .A(n13921), .B(n13922), .Z(n13919) );
  XNOR U17047 ( .A(n13920), .B(n13849), .Z(n13922) );
  XOR U17048 ( .A(n13913), .B(n13914), .Z(n13849) );
  XNOR U17049 ( .A(n13923), .B(n13924), .Z(n13914) );
  ANDN U17050 ( .B(n13925), .A(n13926), .Z(n13923) );
  XOR U17051 ( .A(n13927), .B(n13928), .Z(n13925) );
  XOR U17052 ( .A(n13929), .B(n13930), .Z(n13913) );
  XNOR U17053 ( .A(n13931), .B(n13932), .Z(n13930) );
  ANDN U17054 ( .B(n13933), .A(n13934), .Z(n13931) );
  XNOR U17055 ( .A(n13935), .B(n13936), .Z(n13933) );
  IV U17056 ( .A(n13911), .Z(n13929) );
  XOR U17057 ( .A(n13937), .B(n13938), .Z(n13911) );
  ANDN U17058 ( .B(n13939), .A(n13940), .Z(n13937) );
  XOR U17059 ( .A(n13938), .B(n13941), .Z(n13939) );
  XOR U17060 ( .A(n13920), .B(n13851), .Z(n13921) );
  XOR U17061 ( .A(n13942), .B(n13943), .Z(n13851) );
  AND U17062 ( .A(n98), .B(n13944), .Z(n13942) );
  XOR U17063 ( .A(n13945), .B(n13943), .Z(n13944) );
  XNOR U17064 ( .A(n13946), .B(n13947), .Z(n13920) );
  NAND U17065 ( .A(n13948), .B(n13949), .Z(n13947) );
  XOR U17066 ( .A(n13950), .B(n13899), .Z(n13949) );
  XOR U17067 ( .A(n13940), .B(n13941), .Z(n13899) );
  XOR U17068 ( .A(n13951), .B(n13928), .Z(n13941) );
  XOR U17069 ( .A(n13952), .B(n13953), .Z(n13928) );
  ANDN U17070 ( .B(n13954), .A(n13955), .Z(n13952) );
  XOR U17071 ( .A(n13953), .B(n13956), .Z(n13954) );
  IV U17072 ( .A(n13926), .Z(n13951) );
  XOR U17073 ( .A(n13924), .B(n13957), .Z(n13926) );
  XOR U17074 ( .A(n13958), .B(n13959), .Z(n13957) );
  ANDN U17075 ( .B(n13960), .A(n13961), .Z(n13958) );
  XOR U17076 ( .A(n13962), .B(n13959), .Z(n13960) );
  IV U17077 ( .A(n13927), .Z(n13924) );
  XOR U17078 ( .A(n13963), .B(n13964), .Z(n13927) );
  ANDN U17079 ( .B(n13965), .A(n13966), .Z(n13963) );
  XOR U17080 ( .A(n13964), .B(n13967), .Z(n13965) );
  XOR U17081 ( .A(n13968), .B(n13969), .Z(n13940) );
  XNOR U17082 ( .A(n13935), .B(n13970), .Z(n13969) );
  IV U17083 ( .A(n13938), .Z(n13970) );
  XOR U17084 ( .A(n13971), .B(n13972), .Z(n13938) );
  ANDN U17085 ( .B(n13973), .A(n13974), .Z(n13971) );
  XOR U17086 ( .A(n13972), .B(n13975), .Z(n13973) );
  XNOR U17087 ( .A(n13976), .B(n13977), .Z(n13935) );
  ANDN U17088 ( .B(n13978), .A(n13979), .Z(n13976) );
  XOR U17089 ( .A(n13977), .B(n13980), .Z(n13978) );
  IV U17090 ( .A(n13934), .Z(n13968) );
  XOR U17091 ( .A(n13932), .B(n13981), .Z(n13934) );
  XOR U17092 ( .A(n13982), .B(n13983), .Z(n13981) );
  ANDN U17093 ( .B(n13984), .A(n13985), .Z(n13982) );
  XOR U17094 ( .A(n13986), .B(n13983), .Z(n13984) );
  IV U17095 ( .A(n13936), .Z(n13932) );
  XOR U17096 ( .A(n13987), .B(n13988), .Z(n13936) );
  ANDN U17097 ( .B(n13989), .A(n13990), .Z(n13987) );
  XOR U17098 ( .A(n13991), .B(n13988), .Z(n13989) );
  IV U17099 ( .A(n13946), .Z(n13950) );
  XOR U17100 ( .A(n13946), .B(n13901), .Z(n13948) );
  XOR U17101 ( .A(n13992), .B(n13993), .Z(n13901) );
  AND U17102 ( .A(n98), .B(n13994), .Z(n13992) );
  XOR U17103 ( .A(n13995), .B(n13993), .Z(n13994) );
  NANDN U17104 ( .A(n13903), .B(n13905), .Z(n13946) );
  XOR U17105 ( .A(n13996), .B(n13997), .Z(n13905) );
  AND U17106 ( .A(n98), .B(n13998), .Z(n13996) );
  XOR U17107 ( .A(n13997), .B(n13999), .Z(n13998) );
  XNOR U17108 ( .A(n14000), .B(n14001), .Z(n98) );
  AND U17109 ( .A(n14002), .B(n14003), .Z(n14000) );
  XOR U17110 ( .A(n14001), .B(n13916), .Z(n14003) );
  XNOR U17111 ( .A(n14004), .B(n14005), .Z(n13916) );
  ANDN U17112 ( .B(n14006), .A(n14007), .Z(n14004) );
  XOR U17113 ( .A(n14005), .B(n14008), .Z(n14006) );
  XNOR U17114 ( .A(n14001), .B(n13918), .Z(n14002) );
  XOR U17115 ( .A(n14009), .B(n14010), .Z(n13918) );
  AND U17116 ( .A(n102), .B(n14011), .Z(n14009) );
  XOR U17117 ( .A(n14012), .B(n14010), .Z(n14011) );
  XNOR U17118 ( .A(n14013), .B(n14014), .Z(n14001) );
  AND U17119 ( .A(n14015), .B(n14016), .Z(n14013) );
  XNOR U17120 ( .A(n14014), .B(n13943), .Z(n14016) );
  XOR U17121 ( .A(n14007), .B(n14008), .Z(n13943) );
  XNOR U17122 ( .A(n14017), .B(n14018), .Z(n14008) );
  ANDN U17123 ( .B(n14019), .A(n14020), .Z(n14017) );
  XOR U17124 ( .A(n14021), .B(n14022), .Z(n14019) );
  XOR U17125 ( .A(n14023), .B(n14024), .Z(n14007) );
  XNOR U17126 ( .A(n14025), .B(n14026), .Z(n14024) );
  ANDN U17127 ( .B(n14027), .A(n14028), .Z(n14025) );
  XNOR U17128 ( .A(n14029), .B(n14030), .Z(n14027) );
  IV U17129 ( .A(n14005), .Z(n14023) );
  XOR U17130 ( .A(n14031), .B(n14032), .Z(n14005) );
  ANDN U17131 ( .B(n14033), .A(n14034), .Z(n14031) );
  XOR U17132 ( .A(n14032), .B(n14035), .Z(n14033) );
  XOR U17133 ( .A(n14014), .B(n13945), .Z(n14015) );
  XOR U17134 ( .A(n14036), .B(n14037), .Z(n13945) );
  AND U17135 ( .A(n102), .B(n14038), .Z(n14036) );
  XOR U17136 ( .A(n14039), .B(n14037), .Z(n14038) );
  XNOR U17137 ( .A(n14040), .B(n14041), .Z(n14014) );
  NAND U17138 ( .A(n14042), .B(n14043), .Z(n14041) );
  XOR U17139 ( .A(n14044), .B(n13993), .Z(n14043) );
  XOR U17140 ( .A(n14034), .B(n14035), .Z(n13993) );
  XOR U17141 ( .A(n14045), .B(n14022), .Z(n14035) );
  XOR U17142 ( .A(n14046), .B(n14047), .Z(n14022) );
  ANDN U17143 ( .B(n14048), .A(n14049), .Z(n14046) );
  XOR U17144 ( .A(n14047), .B(n14050), .Z(n14048) );
  IV U17145 ( .A(n14020), .Z(n14045) );
  XOR U17146 ( .A(n14018), .B(n14051), .Z(n14020) );
  XOR U17147 ( .A(n14052), .B(n14053), .Z(n14051) );
  ANDN U17148 ( .B(n14054), .A(n14055), .Z(n14052) );
  XOR U17149 ( .A(n14056), .B(n14053), .Z(n14054) );
  IV U17150 ( .A(n14021), .Z(n14018) );
  XOR U17151 ( .A(n14057), .B(n14058), .Z(n14021) );
  ANDN U17152 ( .B(n14059), .A(n14060), .Z(n14057) );
  XOR U17153 ( .A(n14058), .B(n14061), .Z(n14059) );
  XOR U17154 ( .A(n14062), .B(n14063), .Z(n14034) );
  XNOR U17155 ( .A(n14029), .B(n14064), .Z(n14063) );
  IV U17156 ( .A(n14032), .Z(n14064) );
  XOR U17157 ( .A(n14065), .B(n14066), .Z(n14032) );
  ANDN U17158 ( .B(n14067), .A(n14068), .Z(n14065) );
  XOR U17159 ( .A(n14066), .B(n14069), .Z(n14067) );
  XNOR U17160 ( .A(n14070), .B(n14071), .Z(n14029) );
  ANDN U17161 ( .B(n14072), .A(n14073), .Z(n14070) );
  XOR U17162 ( .A(n14071), .B(n14074), .Z(n14072) );
  IV U17163 ( .A(n14028), .Z(n14062) );
  XOR U17164 ( .A(n14026), .B(n14075), .Z(n14028) );
  XOR U17165 ( .A(n14076), .B(n14077), .Z(n14075) );
  ANDN U17166 ( .B(n14078), .A(n14079), .Z(n14076) );
  XOR U17167 ( .A(n14080), .B(n14077), .Z(n14078) );
  IV U17168 ( .A(n14030), .Z(n14026) );
  XOR U17169 ( .A(n14081), .B(n14082), .Z(n14030) );
  ANDN U17170 ( .B(n14083), .A(n14084), .Z(n14081) );
  XOR U17171 ( .A(n14085), .B(n14082), .Z(n14083) );
  IV U17172 ( .A(n14040), .Z(n14044) );
  XOR U17173 ( .A(n14040), .B(n13995), .Z(n14042) );
  XOR U17174 ( .A(n14086), .B(n14087), .Z(n13995) );
  AND U17175 ( .A(n102), .B(n14088), .Z(n14086) );
  XOR U17176 ( .A(n14089), .B(n14087), .Z(n14088) );
  NANDN U17177 ( .A(n13997), .B(n13999), .Z(n14040) );
  XOR U17178 ( .A(n14090), .B(n14091), .Z(n13999) );
  AND U17179 ( .A(n102), .B(n14092), .Z(n14090) );
  XOR U17180 ( .A(n14091), .B(n14093), .Z(n14092) );
  XNOR U17181 ( .A(n14094), .B(n14095), .Z(n102) );
  AND U17182 ( .A(n14096), .B(n14097), .Z(n14094) );
  XOR U17183 ( .A(n14095), .B(n14010), .Z(n14097) );
  XNOR U17184 ( .A(n14098), .B(n14099), .Z(n14010) );
  ANDN U17185 ( .B(n14100), .A(n14101), .Z(n14098) );
  XOR U17186 ( .A(n14099), .B(n14102), .Z(n14100) );
  XNOR U17187 ( .A(n14095), .B(n14012), .Z(n14096) );
  XOR U17188 ( .A(n14103), .B(n14104), .Z(n14012) );
  AND U17189 ( .A(n106), .B(n14105), .Z(n14103) );
  XOR U17190 ( .A(n14106), .B(n14104), .Z(n14105) );
  XNOR U17191 ( .A(n14107), .B(n14108), .Z(n14095) );
  AND U17192 ( .A(n14109), .B(n14110), .Z(n14107) );
  XNOR U17193 ( .A(n14108), .B(n14037), .Z(n14110) );
  XOR U17194 ( .A(n14101), .B(n14102), .Z(n14037) );
  XNOR U17195 ( .A(n14111), .B(n14112), .Z(n14102) );
  ANDN U17196 ( .B(n14113), .A(n14114), .Z(n14111) );
  XOR U17197 ( .A(n14115), .B(n14116), .Z(n14113) );
  XOR U17198 ( .A(n14117), .B(n14118), .Z(n14101) );
  XNOR U17199 ( .A(n14119), .B(n14120), .Z(n14118) );
  ANDN U17200 ( .B(n14121), .A(n14122), .Z(n14119) );
  XNOR U17201 ( .A(n14123), .B(n14124), .Z(n14121) );
  IV U17202 ( .A(n14099), .Z(n14117) );
  XOR U17203 ( .A(n14125), .B(n14126), .Z(n14099) );
  ANDN U17204 ( .B(n14127), .A(n14128), .Z(n14125) );
  XOR U17205 ( .A(n14126), .B(n14129), .Z(n14127) );
  XOR U17206 ( .A(n14108), .B(n14039), .Z(n14109) );
  XOR U17207 ( .A(n14130), .B(n14131), .Z(n14039) );
  AND U17208 ( .A(n106), .B(n14132), .Z(n14130) );
  XOR U17209 ( .A(n14133), .B(n14131), .Z(n14132) );
  XNOR U17210 ( .A(n14134), .B(n14135), .Z(n14108) );
  NAND U17211 ( .A(n14136), .B(n14137), .Z(n14135) );
  XOR U17212 ( .A(n14138), .B(n14087), .Z(n14137) );
  XOR U17213 ( .A(n14128), .B(n14129), .Z(n14087) );
  XOR U17214 ( .A(n14139), .B(n14116), .Z(n14129) );
  XOR U17215 ( .A(n14140), .B(n14141), .Z(n14116) );
  ANDN U17216 ( .B(n14142), .A(n14143), .Z(n14140) );
  XOR U17217 ( .A(n14141), .B(n14144), .Z(n14142) );
  IV U17218 ( .A(n14114), .Z(n14139) );
  XOR U17219 ( .A(n14112), .B(n14145), .Z(n14114) );
  XOR U17220 ( .A(n14146), .B(n14147), .Z(n14145) );
  ANDN U17221 ( .B(n14148), .A(n14149), .Z(n14146) );
  XOR U17222 ( .A(n14150), .B(n14147), .Z(n14148) );
  IV U17223 ( .A(n14115), .Z(n14112) );
  XOR U17224 ( .A(n14151), .B(n14152), .Z(n14115) );
  ANDN U17225 ( .B(n14153), .A(n14154), .Z(n14151) );
  XOR U17226 ( .A(n14152), .B(n14155), .Z(n14153) );
  XOR U17227 ( .A(n14156), .B(n14157), .Z(n14128) );
  XNOR U17228 ( .A(n14123), .B(n14158), .Z(n14157) );
  IV U17229 ( .A(n14126), .Z(n14158) );
  XOR U17230 ( .A(n14159), .B(n14160), .Z(n14126) );
  ANDN U17231 ( .B(n14161), .A(n14162), .Z(n14159) );
  XOR U17232 ( .A(n14160), .B(n14163), .Z(n14161) );
  XNOR U17233 ( .A(n14164), .B(n14165), .Z(n14123) );
  ANDN U17234 ( .B(n14166), .A(n14167), .Z(n14164) );
  XOR U17235 ( .A(n14165), .B(n14168), .Z(n14166) );
  IV U17236 ( .A(n14122), .Z(n14156) );
  XOR U17237 ( .A(n14120), .B(n14169), .Z(n14122) );
  XOR U17238 ( .A(n14170), .B(n14171), .Z(n14169) );
  ANDN U17239 ( .B(n14172), .A(n14173), .Z(n14170) );
  XOR U17240 ( .A(n14174), .B(n14171), .Z(n14172) );
  IV U17241 ( .A(n14124), .Z(n14120) );
  XOR U17242 ( .A(n14175), .B(n14176), .Z(n14124) );
  ANDN U17243 ( .B(n14177), .A(n14178), .Z(n14175) );
  XOR U17244 ( .A(n14179), .B(n14176), .Z(n14177) );
  IV U17245 ( .A(n14134), .Z(n14138) );
  XOR U17246 ( .A(n14134), .B(n14089), .Z(n14136) );
  XOR U17247 ( .A(n14180), .B(n14181), .Z(n14089) );
  AND U17248 ( .A(n106), .B(n14182), .Z(n14180) );
  XOR U17249 ( .A(n14183), .B(n14181), .Z(n14182) );
  NANDN U17250 ( .A(n14091), .B(n14093), .Z(n14134) );
  XOR U17251 ( .A(n14184), .B(n14185), .Z(n14093) );
  AND U17252 ( .A(n106), .B(n14186), .Z(n14184) );
  XOR U17253 ( .A(n14185), .B(n14187), .Z(n14186) );
  XNOR U17254 ( .A(n14188), .B(n14189), .Z(n106) );
  AND U17255 ( .A(n14190), .B(n14191), .Z(n14188) );
  XOR U17256 ( .A(n14189), .B(n14104), .Z(n14191) );
  XNOR U17257 ( .A(n14192), .B(n14193), .Z(n14104) );
  ANDN U17258 ( .B(n14194), .A(n14195), .Z(n14192) );
  XOR U17259 ( .A(n14193), .B(n14196), .Z(n14194) );
  XNOR U17260 ( .A(n14189), .B(n14106), .Z(n14190) );
  XOR U17261 ( .A(n14197), .B(n14198), .Z(n14106) );
  AND U17262 ( .A(n110), .B(n14199), .Z(n14197) );
  XOR U17263 ( .A(n14200), .B(n14198), .Z(n14199) );
  XNOR U17264 ( .A(n14201), .B(n14202), .Z(n14189) );
  AND U17265 ( .A(n14203), .B(n14204), .Z(n14201) );
  XNOR U17266 ( .A(n14202), .B(n14131), .Z(n14204) );
  XOR U17267 ( .A(n14195), .B(n14196), .Z(n14131) );
  XNOR U17268 ( .A(n14205), .B(n14206), .Z(n14196) );
  ANDN U17269 ( .B(n14207), .A(n14208), .Z(n14205) );
  XOR U17270 ( .A(n14209), .B(n14210), .Z(n14207) );
  XOR U17271 ( .A(n14211), .B(n14212), .Z(n14195) );
  XNOR U17272 ( .A(n14213), .B(n14214), .Z(n14212) );
  ANDN U17273 ( .B(n14215), .A(n14216), .Z(n14213) );
  XNOR U17274 ( .A(n14217), .B(n14218), .Z(n14215) );
  IV U17275 ( .A(n14193), .Z(n14211) );
  XOR U17276 ( .A(n14219), .B(n14220), .Z(n14193) );
  ANDN U17277 ( .B(n14221), .A(n14222), .Z(n14219) );
  XOR U17278 ( .A(n14220), .B(n14223), .Z(n14221) );
  XOR U17279 ( .A(n14202), .B(n14133), .Z(n14203) );
  XOR U17280 ( .A(n14224), .B(n14225), .Z(n14133) );
  AND U17281 ( .A(n110), .B(n14226), .Z(n14224) );
  XOR U17282 ( .A(n14227), .B(n14225), .Z(n14226) );
  XNOR U17283 ( .A(n14228), .B(n14229), .Z(n14202) );
  NAND U17284 ( .A(n14230), .B(n14231), .Z(n14229) );
  XOR U17285 ( .A(n14232), .B(n14181), .Z(n14231) );
  XOR U17286 ( .A(n14222), .B(n14223), .Z(n14181) );
  XOR U17287 ( .A(n14233), .B(n14210), .Z(n14223) );
  XOR U17288 ( .A(n14234), .B(n14235), .Z(n14210) );
  ANDN U17289 ( .B(n14236), .A(n14237), .Z(n14234) );
  XOR U17290 ( .A(n14235), .B(n14238), .Z(n14236) );
  IV U17291 ( .A(n14208), .Z(n14233) );
  XOR U17292 ( .A(n14206), .B(n14239), .Z(n14208) );
  XOR U17293 ( .A(n14240), .B(n14241), .Z(n14239) );
  ANDN U17294 ( .B(n14242), .A(n14243), .Z(n14240) );
  XOR U17295 ( .A(n14244), .B(n14241), .Z(n14242) );
  IV U17296 ( .A(n14209), .Z(n14206) );
  XOR U17297 ( .A(n14245), .B(n14246), .Z(n14209) );
  ANDN U17298 ( .B(n14247), .A(n14248), .Z(n14245) );
  XOR U17299 ( .A(n14246), .B(n14249), .Z(n14247) );
  XOR U17300 ( .A(n14250), .B(n14251), .Z(n14222) );
  XNOR U17301 ( .A(n14217), .B(n14252), .Z(n14251) );
  IV U17302 ( .A(n14220), .Z(n14252) );
  XOR U17303 ( .A(n14253), .B(n14254), .Z(n14220) );
  ANDN U17304 ( .B(n14255), .A(n14256), .Z(n14253) );
  XOR U17305 ( .A(n14254), .B(n14257), .Z(n14255) );
  XNOR U17306 ( .A(n14258), .B(n14259), .Z(n14217) );
  ANDN U17307 ( .B(n14260), .A(n14261), .Z(n14258) );
  XOR U17308 ( .A(n14259), .B(n14262), .Z(n14260) );
  IV U17309 ( .A(n14216), .Z(n14250) );
  XOR U17310 ( .A(n14214), .B(n14263), .Z(n14216) );
  XOR U17311 ( .A(n14264), .B(n14265), .Z(n14263) );
  ANDN U17312 ( .B(n14266), .A(n14267), .Z(n14264) );
  XOR U17313 ( .A(n14268), .B(n14265), .Z(n14266) );
  IV U17314 ( .A(n14218), .Z(n14214) );
  XOR U17315 ( .A(n14269), .B(n14270), .Z(n14218) );
  ANDN U17316 ( .B(n14271), .A(n14272), .Z(n14269) );
  XOR U17317 ( .A(n14273), .B(n14270), .Z(n14271) );
  IV U17318 ( .A(n14228), .Z(n14232) );
  XOR U17319 ( .A(n14228), .B(n14183), .Z(n14230) );
  XOR U17320 ( .A(n14274), .B(n14275), .Z(n14183) );
  AND U17321 ( .A(n110), .B(n14276), .Z(n14274) );
  XOR U17322 ( .A(n14277), .B(n14275), .Z(n14276) );
  NANDN U17323 ( .A(n14185), .B(n14187), .Z(n14228) );
  XOR U17324 ( .A(n14278), .B(n14279), .Z(n14187) );
  AND U17325 ( .A(n110), .B(n14280), .Z(n14278) );
  XOR U17326 ( .A(n14279), .B(n14281), .Z(n14280) );
  XNOR U17327 ( .A(n14282), .B(n14283), .Z(n110) );
  AND U17328 ( .A(n14284), .B(n14285), .Z(n14282) );
  XOR U17329 ( .A(n14283), .B(n14198), .Z(n14285) );
  XNOR U17330 ( .A(n14286), .B(n14287), .Z(n14198) );
  ANDN U17331 ( .B(n14288), .A(n14289), .Z(n14286) );
  XOR U17332 ( .A(n14287), .B(n14290), .Z(n14288) );
  XNOR U17333 ( .A(n14283), .B(n14200), .Z(n14284) );
  XOR U17334 ( .A(n14291), .B(n14292), .Z(n14200) );
  AND U17335 ( .A(n114), .B(n14293), .Z(n14291) );
  XOR U17336 ( .A(n14294), .B(n14292), .Z(n14293) );
  XNOR U17337 ( .A(n14295), .B(n14296), .Z(n14283) );
  AND U17338 ( .A(n14297), .B(n14298), .Z(n14295) );
  XNOR U17339 ( .A(n14296), .B(n14225), .Z(n14298) );
  XOR U17340 ( .A(n14289), .B(n14290), .Z(n14225) );
  XNOR U17341 ( .A(n14299), .B(n14300), .Z(n14290) );
  ANDN U17342 ( .B(n14301), .A(n14302), .Z(n14299) );
  XOR U17343 ( .A(n14303), .B(n14304), .Z(n14301) );
  XOR U17344 ( .A(n14305), .B(n14306), .Z(n14289) );
  XNOR U17345 ( .A(n14307), .B(n14308), .Z(n14306) );
  ANDN U17346 ( .B(n14309), .A(n14310), .Z(n14307) );
  XNOR U17347 ( .A(n14311), .B(n14312), .Z(n14309) );
  IV U17348 ( .A(n14287), .Z(n14305) );
  XOR U17349 ( .A(n14313), .B(n14314), .Z(n14287) );
  ANDN U17350 ( .B(n14315), .A(n14316), .Z(n14313) );
  XOR U17351 ( .A(n14314), .B(n14317), .Z(n14315) );
  XOR U17352 ( .A(n14296), .B(n14227), .Z(n14297) );
  XOR U17353 ( .A(n14318), .B(n14319), .Z(n14227) );
  AND U17354 ( .A(n114), .B(n14320), .Z(n14318) );
  XOR U17355 ( .A(n14321), .B(n14319), .Z(n14320) );
  XNOR U17356 ( .A(n14322), .B(n14323), .Z(n14296) );
  NAND U17357 ( .A(n14324), .B(n14325), .Z(n14323) );
  XOR U17358 ( .A(n14326), .B(n14275), .Z(n14325) );
  XOR U17359 ( .A(n14316), .B(n14317), .Z(n14275) );
  XOR U17360 ( .A(n14327), .B(n14304), .Z(n14317) );
  XOR U17361 ( .A(n14328), .B(n14329), .Z(n14304) );
  ANDN U17362 ( .B(n14330), .A(n14331), .Z(n14328) );
  XOR U17363 ( .A(n14329), .B(n14332), .Z(n14330) );
  IV U17364 ( .A(n14302), .Z(n14327) );
  XOR U17365 ( .A(n14300), .B(n14333), .Z(n14302) );
  XOR U17366 ( .A(n14334), .B(n14335), .Z(n14333) );
  ANDN U17367 ( .B(n14336), .A(n14337), .Z(n14334) );
  XOR U17368 ( .A(n14338), .B(n14335), .Z(n14336) );
  IV U17369 ( .A(n14303), .Z(n14300) );
  XOR U17370 ( .A(n14339), .B(n14340), .Z(n14303) );
  ANDN U17371 ( .B(n14341), .A(n14342), .Z(n14339) );
  XOR U17372 ( .A(n14340), .B(n14343), .Z(n14341) );
  XOR U17373 ( .A(n14344), .B(n14345), .Z(n14316) );
  XNOR U17374 ( .A(n14311), .B(n14346), .Z(n14345) );
  IV U17375 ( .A(n14314), .Z(n14346) );
  XOR U17376 ( .A(n14347), .B(n14348), .Z(n14314) );
  ANDN U17377 ( .B(n14349), .A(n14350), .Z(n14347) );
  XOR U17378 ( .A(n14348), .B(n14351), .Z(n14349) );
  XNOR U17379 ( .A(n14352), .B(n14353), .Z(n14311) );
  ANDN U17380 ( .B(n14354), .A(n14355), .Z(n14352) );
  XOR U17381 ( .A(n14353), .B(n14356), .Z(n14354) );
  IV U17382 ( .A(n14310), .Z(n14344) );
  XOR U17383 ( .A(n14308), .B(n14357), .Z(n14310) );
  XOR U17384 ( .A(n14358), .B(n14359), .Z(n14357) );
  ANDN U17385 ( .B(n14360), .A(n14361), .Z(n14358) );
  XOR U17386 ( .A(n14362), .B(n14359), .Z(n14360) );
  IV U17387 ( .A(n14312), .Z(n14308) );
  XOR U17388 ( .A(n14363), .B(n14364), .Z(n14312) );
  ANDN U17389 ( .B(n14365), .A(n14366), .Z(n14363) );
  XOR U17390 ( .A(n14367), .B(n14364), .Z(n14365) );
  IV U17391 ( .A(n14322), .Z(n14326) );
  XOR U17392 ( .A(n14322), .B(n14277), .Z(n14324) );
  XOR U17393 ( .A(n14368), .B(n14369), .Z(n14277) );
  AND U17394 ( .A(n114), .B(n14370), .Z(n14368) );
  XOR U17395 ( .A(n14371), .B(n14369), .Z(n14370) );
  NANDN U17396 ( .A(n14279), .B(n14281), .Z(n14322) );
  XOR U17397 ( .A(n14372), .B(n14373), .Z(n14281) );
  AND U17398 ( .A(n114), .B(n14374), .Z(n14372) );
  XOR U17399 ( .A(n14373), .B(n14375), .Z(n14374) );
  XNOR U17400 ( .A(n14376), .B(n14377), .Z(n114) );
  AND U17401 ( .A(n14378), .B(n14379), .Z(n14376) );
  XOR U17402 ( .A(n14377), .B(n14292), .Z(n14379) );
  XNOR U17403 ( .A(n14380), .B(n14381), .Z(n14292) );
  ANDN U17404 ( .B(n14382), .A(n14383), .Z(n14380) );
  XOR U17405 ( .A(n14381), .B(n14384), .Z(n14382) );
  XNOR U17406 ( .A(n14377), .B(n14294), .Z(n14378) );
  XOR U17407 ( .A(n14385), .B(n14386), .Z(n14294) );
  AND U17408 ( .A(n118), .B(n14387), .Z(n14385) );
  XOR U17409 ( .A(n14388), .B(n14386), .Z(n14387) );
  XNOR U17410 ( .A(n14389), .B(n14390), .Z(n14377) );
  AND U17411 ( .A(n14391), .B(n14392), .Z(n14389) );
  XNOR U17412 ( .A(n14390), .B(n14319), .Z(n14392) );
  XOR U17413 ( .A(n14383), .B(n14384), .Z(n14319) );
  XNOR U17414 ( .A(n14393), .B(n14394), .Z(n14384) );
  ANDN U17415 ( .B(n14395), .A(n14396), .Z(n14393) );
  XOR U17416 ( .A(n14397), .B(n14398), .Z(n14395) );
  XOR U17417 ( .A(n14399), .B(n14400), .Z(n14383) );
  XNOR U17418 ( .A(n14401), .B(n14402), .Z(n14400) );
  ANDN U17419 ( .B(n14403), .A(n14404), .Z(n14401) );
  XNOR U17420 ( .A(n14405), .B(n14406), .Z(n14403) );
  IV U17421 ( .A(n14381), .Z(n14399) );
  XOR U17422 ( .A(n14407), .B(n14408), .Z(n14381) );
  ANDN U17423 ( .B(n14409), .A(n14410), .Z(n14407) );
  XOR U17424 ( .A(n14408), .B(n14411), .Z(n14409) );
  XOR U17425 ( .A(n14390), .B(n14321), .Z(n14391) );
  XOR U17426 ( .A(n14412), .B(n14413), .Z(n14321) );
  AND U17427 ( .A(n118), .B(n14414), .Z(n14412) );
  XOR U17428 ( .A(n14415), .B(n14413), .Z(n14414) );
  XNOR U17429 ( .A(n14416), .B(n14417), .Z(n14390) );
  NAND U17430 ( .A(n14418), .B(n14419), .Z(n14417) );
  XOR U17431 ( .A(n14420), .B(n14369), .Z(n14419) );
  XOR U17432 ( .A(n14410), .B(n14411), .Z(n14369) );
  XOR U17433 ( .A(n14421), .B(n14398), .Z(n14411) );
  XOR U17434 ( .A(n14422), .B(n14423), .Z(n14398) );
  ANDN U17435 ( .B(n14424), .A(n14425), .Z(n14422) );
  XOR U17436 ( .A(n14423), .B(n14426), .Z(n14424) );
  IV U17437 ( .A(n14396), .Z(n14421) );
  XOR U17438 ( .A(n14394), .B(n14427), .Z(n14396) );
  XOR U17439 ( .A(n14428), .B(n14429), .Z(n14427) );
  ANDN U17440 ( .B(n14430), .A(n14431), .Z(n14428) );
  XOR U17441 ( .A(n14432), .B(n14429), .Z(n14430) );
  IV U17442 ( .A(n14397), .Z(n14394) );
  XOR U17443 ( .A(n14433), .B(n14434), .Z(n14397) );
  ANDN U17444 ( .B(n14435), .A(n14436), .Z(n14433) );
  XOR U17445 ( .A(n14434), .B(n14437), .Z(n14435) );
  XOR U17446 ( .A(n14438), .B(n14439), .Z(n14410) );
  XNOR U17447 ( .A(n14405), .B(n14440), .Z(n14439) );
  IV U17448 ( .A(n14408), .Z(n14440) );
  XOR U17449 ( .A(n14441), .B(n14442), .Z(n14408) );
  ANDN U17450 ( .B(n14443), .A(n14444), .Z(n14441) );
  XOR U17451 ( .A(n14442), .B(n14445), .Z(n14443) );
  XNOR U17452 ( .A(n14446), .B(n14447), .Z(n14405) );
  ANDN U17453 ( .B(n14448), .A(n14449), .Z(n14446) );
  XOR U17454 ( .A(n14447), .B(n14450), .Z(n14448) );
  IV U17455 ( .A(n14404), .Z(n14438) );
  XOR U17456 ( .A(n14402), .B(n14451), .Z(n14404) );
  XOR U17457 ( .A(n14452), .B(n14453), .Z(n14451) );
  ANDN U17458 ( .B(n14454), .A(n14455), .Z(n14452) );
  XOR U17459 ( .A(n14456), .B(n14453), .Z(n14454) );
  IV U17460 ( .A(n14406), .Z(n14402) );
  XOR U17461 ( .A(n14457), .B(n14458), .Z(n14406) );
  ANDN U17462 ( .B(n14459), .A(n14460), .Z(n14457) );
  XOR U17463 ( .A(n14461), .B(n14458), .Z(n14459) );
  IV U17464 ( .A(n14416), .Z(n14420) );
  XOR U17465 ( .A(n14416), .B(n14371), .Z(n14418) );
  XOR U17466 ( .A(n14462), .B(n14463), .Z(n14371) );
  AND U17467 ( .A(n118), .B(n14464), .Z(n14462) );
  XOR U17468 ( .A(n14465), .B(n14463), .Z(n14464) );
  NANDN U17469 ( .A(n14373), .B(n14375), .Z(n14416) );
  XOR U17470 ( .A(n14466), .B(n14467), .Z(n14375) );
  AND U17471 ( .A(n118), .B(n14468), .Z(n14466) );
  XOR U17472 ( .A(n14467), .B(n14469), .Z(n14468) );
  XNOR U17473 ( .A(n14470), .B(n14471), .Z(n118) );
  AND U17474 ( .A(n14472), .B(n14473), .Z(n14470) );
  XOR U17475 ( .A(n14471), .B(n14386), .Z(n14473) );
  XNOR U17476 ( .A(n14474), .B(n14475), .Z(n14386) );
  ANDN U17477 ( .B(n14476), .A(n14477), .Z(n14474) );
  XOR U17478 ( .A(n14475), .B(n14478), .Z(n14476) );
  XNOR U17479 ( .A(n14471), .B(n14388), .Z(n14472) );
  XOR U17480 ( .A(n14479), .B(n14480), .Z(n14388) );
  AND U17481 ( .A(n122), .B(n14481), .Z(n14479) );
  XOR U17482 ( .A(n14482), .B(n14480), .Z(n14481) );
  XNOR U17483 ( .A(n14483), .B(n14484), .Z(n14471) );
  AND U17484 ( .A(n14485), .B(n14486), .Z(n14483) );
  XNOR U17485 ( .A(n14484), .B(n14413), .Z(n14486) );
  XOR U17486 ( .A(n14477), .B(n14478), .Z(n14413) );
  XNOR U17487 ( .A(n14487), .B(n14488), .Z(n14478) );
  ANDN U17488 ( .B(n14489), .A(n14490), .Z(n14487) );
  XOR U17489 ( .A(n14491), .B(n14492), .Z(n14489) );
  XOR U17490 ( .A(n14493), .B(n14494), .Z(n14477) );
  XNOR U17491 ( .A(n14495), .B(n14496), .Z(n14494) );
  ANDN U17492 ( .B(n14497), .A(n14498), .Z(n14495) );
  XNOR U17493 ( .A(n14499), .B(n14500), .Z(n14497) );
  IV U17494 ( .A(n14475), .Z(n14493) );
  XOR U17495 ( .A(n14501), .B(n14502), .Z(n14475) );
  ANDN U17496 ( .B(n14503), .A(n14504), .Z(n14501) );
  XOR U17497 ( .A(n14502), .B(n14505), .Z(n14503) );
  XOR U17498 ( .A(n14484), .B(n14415), .Z(n14485) );
  XOR U17499 ( .A(n14506), .B(n14507), .Z(n14415) );
  AND U17500 ( .A(n122), .B(n14508), .Z(n14506) );
  XOR U17501 ( .A(n14509), .B(n14507), .Z(n14508) );
  XNOR U17502 ( .A(n14510), .B(n14511), .Z(n14484) );
  NAND U17503 ( .A(n14512), .B(n14513), .Z(n14511) );
  XOR U17504 ( .A(n14514), .B(n14463), .Z(n14513) );
  XOR U17505 ( .A(n14504), .B(n14505), .Z(n14463) );
  XOR U17506 ( .A(n14515), .B(n14492), .Z(n14505) );
  XOR U17507 ( .A(n14516), .B(n14517), .Z(n14492) );
  ANDN U17508 ( .B(n14518), .A(n14519), .Z(n14516) );
  XOR U17509 ( .A(n14517), .B(n14520), .Z(n14518) );
  IV U17510 ( .A(n14490), .Z(n14515) );
  XOR U17511 ( .A(n14488), .B(n14521), .Z(n14490) );
  XOR U17512 ( .A(n14522), .B(n14523), .Z(n14521) );
  ANDN U17513 ( .B(n14524), .A(n14525), .Z(n14522) );
  XOR U17514 ( .A(n14526), .B(n14523), .Z(n14524) );
  IV U17515 ( .A(n14491), .Z(n14488) );
  XOR U17516 ( .A(n14527), .B(n14528), .Z(n14491) );
  ANDN U17517 ( .B(n14529), .A(n14530), .Z(n14527) );
  XOR U17518 ( .A(n14528), .B(n14531), .Z(n14529) );
  XOR U17519 ( .A(n14532), .B(n14533), .Z(n14504) );
  XNOR U17520 ( .A(n14499), .B(n14534), .Z(n14533) );
  IV U17521 ( .A(n14502), .Z(n14534) );
  XOR U17522 ( .A(n14535), .B(n14536), .Z(n14502) );
  ANDN U17523 ( .B(n14537), .A(n14538), .Z(n14535) );
  XOR U17524 ( .A(n14536), .B(n14539), .Z(n14537) );
  XNOR U17525 ( .A(n14540), .B(n14541), .Z(n14499) );
  ANDN U17526 ( .B(n14542), .A(n14543), .Z(n14540) );
  XOR U17527 ( .A(n14541), .B(n14544), .Z(n14542) );
  IV U17528 ( .A(n14498), .Z(n14532) );
  XOR U17529 ( .A(n14496), .B(n14545), .Z(n14498) );
  XOR U17530 ( .A(n14546), .B(n14547), .Z(n14545) );
  ANDN U17531 ( .B(n14548), .A(n14549), .Z(n14546) );
  XOR U17532 ( .A(n14550), .B(n14547), .Z(n14548) );
  IV U17533 ( .A(n14500), .Z(n14496) );
  XOR U17534 ( .A(n14551), .B(n14552), .Z(n14500) );
  ANDN U17535 ( .B(n14553), .A(n14554), .Z(n14551) );
  XOR U17536 ( .A(n14555), .B(n14552), .Z(n14553) );
  IV U17537 ( .A(n14510), .Z(n14514) );
  XOR U17538 ( .A(n14510), .B(n14465), .Z(n14512) );
  XOR U17539 ( .A(n14556), .B(n14557), .Z(n14465) );
  AND U17540 ( .A(n122), .B(n14558), .Z(n14556) );
  XOR U17541 ( .A(n14559), .B(n14557), .Z(n14558) );
  NANDN U17542 ( .A(n14467), .B(n14469), .Z(n14510) );
  XOR U17543 ( .A(n14560), .B(n14561), .Z(n14469) );
  AND U17544 ( .A(n122), .B(n14562), .Z(n14560) );
  XOR U17545 ( .A(n14561), .B(n14563), .Z(n14562) );
  XNOR U17546 ( .A(n14564), .B(n14565), .Z(n122) );
  AND U17547 ( .A(n14566), .B(n14567), .Z(n14564) );
  XOR U17548 ( .A(n14565), .B(n14480), .Z(n14567) );
  XNOR U17549 ( .A(n14568), .B(n14569), .Z(n14480) );
  ANDN U17550 ( .B(n14570), .A(n14571), .Z(n14568) );
  XOR U17551 ( .A(n14569), .B(n14572), .Z(n14570) );
  XNOR U17552 ( .A(n14565), .B(n14482), .Z(n14566) );
  XOR U17553 ( .A(n14573), .B(n14574), .Z(n14482) );
  AND U17554 ( .A(n126), .B(n14575), .Z(n14573) );
  XOR U17555 ( .A(n14576), .B(n14574), .Z(n14575) );
  XNOR U17556 ( .A(n14577), .B(n14578), .Z(n14565) );
  AND U17557 ( .A(n14579), .B(n14580), .Z(n14577) );
  XNOR U17558 ( .A(n14578), .B(n14507), .Z(n14580) );
  XOR U17559 ( .A(n14571), .B(n14572), .Z(n14507) );
  XNOR U17560 ( .A(n14581), .B(n14582), .Z(n14572) );
  ANDN U17561 ( .B(n14583), .A(n14584), .Z(n14581) );
  XOR U17562 ( .A(n14585), .B(n14586), .Z(n14583) );
  XOR U17563 ( .A(n14587), .B(n14588), .Z(n14571) );
  XNOR U17564 ( .A(n14589), .B(n14590), .Z(n14588) );
  ANDN U17565 ( .B(n14591), .A(n14592), .Z(n14589) );
  XNOR U17566 ( .A(n14593), .B(n14594), .Z(n14591) );
  IV U17567 ( .A(n14569), .Z(n14587) );
  XOR U17568 ( .A(n14595), .B(n14596), .Z(n14569) );
  ANDN U17569 ( .B(n14597), .A(n14598), .Z(n14595) );
  XOR U17570 ( .A(n14596), .B(n14599), .Z(n14597) );
  XOR U17571 ( .A(n14578), .B(n14509), .Z(n14579) );
  XOR U17572 ( .A(n14600), .B(n14601), .Z(n14509) );
  AND U17573 ( .A(n126), .B(n14602), .Z(n14600) );
  XOR U17574 ( .A(n14603), .B(n14601), .Z(n14602) );
  XNOR U17575 ( .A(n14604), .B(n14605), .Z(n14578) );
  NAND U17576 ( .A(n14606), .B(n14607), .Z(n14605) );
  XOR U17577 ( .A(n14608), .B(n14557), .Z(n14607) );
  XOR U17578 ( .A(n14598), .B(n14599), .Z(n14557) );
  XOR U17579 ( .A(n14609), .B(n14586), .Z(n14599) );
  XOR U17580 ( .A(n14610), .B(n14611), .Z(n14586) );
  ANDN U17581 ( .B(n14612), .A(n14613), .Z(n14610) );
  XOR U17582 ( .A(n14611), .B(n14614), .Z(n14612) );
  IV U17583 ( .A(n14584), .Z(n14609) );
  XOR U17584 ( .A(n14582), .B(n14615), .Z(n14584) );
  XOR U17585 ( .A(n14616), .B(n14617), .Z(n14615) );
  ANDN U17586 ( .B(n14618), .A(n14619), .Z(n14616) );
  XOR U17587 ( .A(n14620), .B(n14617), .Z(n14618) );
  IV U17588 ( .A(n14585), .Z(n14582) );
  XOR U17589 ( .A(n14621), .B(n14622), .Z(n14585) );
  ANDN U17590 ( .B(n14623), .A(n14624), .Z(n14621) );
  XOR U17591 ( .A(n14622), .B(n14625), .Z(n14623) );
  XOR U17592 ( .A(n14626), .B(n14627), .Z(n14598) );
  XNOR U17593 ( .A(n14593), .B(n14628), .Z(n14627) );
  IV U17594 ( .A(n14596), .Z(n14628) );
  XOR U17595 ( .A(n14629), .B(n14630), .Z(n14596) );
  ANDN U17596 ( .B(n14631), .A(n14632), .Z(n14629) );
  XOR U17597 ( .A(n14630), .B(n14633), .Z(n14631) );
  XNOR U17598 ( .A(n14634), .B(n14635), .Z(n14593) );
  ANDN U17599 ( .B(n14636), .A(n14637), .Z(n14634) );
  XOR U17600 ( .A(n14635), .B(n14638), .Z(n14636) );
  IV U17601 ( .A(n14592), .Z(n14626) );
  XOR U17602 ( .A(n14590), .B(n14639), .Z(n14592) );
  XOR U17603 ( .A(n14640), .B(n14641), .Z(n14639) );
  ANDN U17604 ( .B(n14642), .A(n14643), .Z(n14640) );
  XOR U17605 ( .A(n14644), .B(n14641), .Z(n14642) );
  IV U17606 ( .A(n14594), .Z(n14590) );
  XOR U17607 ( .A(n14645), .B(n14646), .Z(n14594) );
  ANDN U17608 ( .B(n14647), .A(n14648), .Z(n14645) );
  XOR U17609 ( .A(n14649), .B(n14646), .Z(n14647) );
  IV U17610 ( .A(n14604), .Z(n14608) );
  XOR U17611 ( .A(n14604), .B(n14559), .Z(n14606) );
  XOR U17612 ( .A(n14650), .B(n14651), .Z(n14559) );
  AND U17613 ( .A(n126), .B(n14652), .Z(n14650) );
  XOR U17614 ( .A(n14653), .B(n14651), .Z(n14652) );
  NANDN U17615 ( .A(n14561), .B(n14563), .Z(n14604) );
  XOR U17616 ( .A(n14654), .B(n14655), .Z(n14563) );
  AND U17617 ( .A(n126), .B(n14656), .Z(n14654) );
  XOR U17618 ( .A(n14655), .B(n14657), .Z(n14656) );
  XNOR U17619 ( .A(n14658), .B(n14659), .Z(n126) );
  AND U17620 ( .A(n14660), .B(n14661), .Z(n14658) );
  XOR U17621 ( .A(n14659), .B(n14574), .Z(n14661) );
  XNOR U17622 ( .A(n14662), .B(n14663), .Z(n14574) );
  ANDN U17623 ( .B(n14664), .A(n14665), .Z(n14662) );
  XOR U17624 ( .A(n14663), .B(n14666), .Z(n14664) );
  XNOR U17625 ( .A(n14659), .B(n14576), .Z(n14660) );
  XOR U17626 ( .A(n14667), .B(n14668), .Z(n14576) );
  AND U17627 ( .A(n130), .B(n14669), .Z(n14667) );
  XOR U17628 ( .A(n14670), .B(n14668), .Z(n14669) );
  XNOR U17629 ( .A(n14671), .B(n14672), .Z(n14659) );
  AND U17630 ( .A(n14673), .B(n14674), .Z(n14671) );
  XNOR U17631 ( .A(n14672), .B(n14601), .Z(n14674) );
  XOR U17632 ( .A(n14665), .B(n14666), .Z(n14601) );
  XNOR U17633 ( .A(n14675), .B(n14676), .Z(n14666) );
  ANDN U17634 ( .B(n14677), .A(n14678), .Z(n14675) );
  XOR U17635 ( .A(n14679), .B(n14680), .Z(n14677) );
  XOR U17636 ( .A(n14681), .B(n14682), .Z(n14665) );
  XNOR U17637 ( .A(n14683), .B(n14684), .Z(n14682) );
  ANDN U17638 ( .B(n14685), .A(n14686), .Z(n14683) );
  XNOR U17639 ( .A(n14687), .B(n14688), .Z(n14685) );
  IV U17640 ( .A(n14663), .Z(n14681) );
  XOR U17641 ( .A(n14689), .B(n14690), .Z(n14663) );
  ANDN U17642 ( .B(n14691), .A(n14692), .Z(n14689) );
  XOR U17643 ( .A(n14690), .B(n14693), .Z(n14691) );
  XOR U17644 ( .A(n14672), .B(n14603), .Z(n14673) );
  XOR U17645 ( .A(n14694), .B(n14695), .Z(n14603) );
  AND U17646 ( .A(n130), .B(n14696), .Z(n14694) );
  XOR U17647 ( .A(n14697), .B(n14695), .Z(n14696) );
  XNOR U17648 ( .A(n14698), .B(n14699), .Z(n14672) );
  NAND U17649 ( .A(n14700), .B(n14701), .Z(n14699) );
  XOR U17650 ( .A(n14702), .B(n14651), .Z(n14701) );
  XOR U17651 ( .A(n14692), .B(n14693), .Z(n14651) );
  XOR U17652 ( .A(n14703), .B(n14680), .Z(n14693) );
  XOR U17653 ( .A(n14704), .B(n14705), .Z(n14680) );
  ANDN U17654 ( .B(n14706), .A(n14707), .Z(n14704) );
  XOR U17655 ( .A(n14705), .B(n14708), .Z(n14706) );
  IV U17656 ( .A(n14678), .Z(n14703) );
  XOR U17657 ( .A(n14676), .B(n14709), .Z(n14678) );
  XOR U17658 ( .A(n14710), .B(n14711), .Z(n14709) );
  ANDN U17659 ( .B(n14712), .A(n14713), .Z(n14710) );
  XOR U17660 ( .A(n14714), .B(n14711), .Z(n14712) );
  IV U17661 ( .A(n14679), .Z(n14676) );
  XOR U17662 ( .A(n14715), .B(n14716), .Z(n14679) );
  ANDN U17663 ( .B(n14717), .A(n14718), .Z(n14715) );
  XOR U17664 ( .A(n14716), .B(n14719), .Z(n14717) );
  XOR U17665 ( .A(n14720), .B(n14721), .Z(n14692) );
  XNOR U17666 ( .A(n14687), .B(n14722), .Z(n14721) );
  IV U17667 ( .A(n14690), .Z(n14722) );
  XOR U17668 ( .A(n14723), .B(n14724), .Z(n14690) );
  ANDN U17669 ( .B(n14725), .A(n14726), .Z(n14723) );
  XOR U17670 ( .A(n14724), .B(n14727), .Z(n14725) );
  XNOR U17671 ( .A(n14728), .B(n14729), .Z(n14687) );
  ANDN U17672 ( .B(n14730), .A(n14731), .Z(n14728) );
  XOR U17673 ( .A(n14729), .B(n14732), .Z(n14730) );
  IV U17674 ( .A(n14686), .Z(n14720) );
  XOR U17675 ( .A(n14684), .B(n14733), .Z(n14686) );
  XOR U17676 ( .A(n14734), .B(n14735), .Z(n14733) );
  ANDN U17677 ( .B(n14736), .A(n14737), .Z(n14734) );
  XOR U17678 ( .A(n14738), .B(n14735), .Z(n14736) );
  IV U17679 ( .A(n14688), .Z(n14684) );
  XOR U17680 ( .A(n14739), .B(n14740), .Z(n14688) );
  ANDN U17681 ( .B(n14741), .A(n14742), .Z(n14739) );
  XOR U17682 ( .A(n14743), .B(n14740), .Z(n14741) );
  IV U17683 ( .A(n14698), .Z(n14702) );
  XOR U17684 ( .A(n14698), .B(n14653), .Z(n14700) );
  XOR U17685 ( .A(n14744), .B(n14745), .Z(n14653) );
  AND U17686 ( .A(n130), .B(n14746), .Z(n14744) );
  XOR U17687 ( .A(n14747), .B(n14745), .Z(n14746) );
  NANDN U17688 ( .A(n14655), .B(n14657), .Z(n14698) );
  XOR U17689 ( .A(n14748), .B(n14749), .Z(n14657) );
  AND U17690 ( .A(n130), .B(n14750), .Z(n14748) );
  XOR U17691 ( .A(n14749), .B(n14751), .Z(n14750) );
  XNOR U17692 ( .A(n14752), .B(n14753), .Z(n130) );
  AND U17693 ( .A(n14754), .B(n14755), .Z(n14752) );
  XOR U17694 ( .A(n14753), .B(n14668), .Z(n14755) );
  XNOR U17695 ( .A(n14756), .B(n14757), .Z(n14668) );
  ANDN U17696 ( .B(n14758), .A(n14759), .Z(n14756) );
  XOR U17697 ( .A(n14757), .B(n14760), .Z(n14758) );
  XNOR U17698 ( .A(n14753), .B(n14670), .Z(n14754) );
  XOR U17699 ( .A(n14761), .B(n14762), .Z(n14670) );
  AND U17700 ( .A(n134), .B(n14763), .Z(n14761) );
  XOR U17701 ( .A(n14764), .B(n14762), .Z(n14763) );
  XNOR U17702 ( .A(n14765), .B(n14766), .Z(n14753) );
  AND U17703 ( .A(n14767), .B(n14768), .Z(n14765) );
  XNOR U17704 ( .A(n14766), .B(n14695), .Z(n14768) );
  XOR U17705 ( .A(n14759), .B(n14760), .Z(n14695) );
  XNOR U17706 ( .A(n14769), .B(n14770), .Z(n14760) );
  ANDN U17707 ( .B(n14771), .A(n14772), .Z(n14769) );
  XOR U17708 ( .A(n14773), .B(n14774), .Z(n14771) );
  XOR U17709 ( .A(n14775), .B(n14776), .Z(n14759) );
  XNOR U17710 ( .A(n14777), .B(n14778), .Z(n14776) );
  ANDN U17711 ( .B(n14779), .A(n14780), .Z(n14777) );
  XNOR U17712 ( .A(n14781), .B(n14782), .Z(n14779) );
  IV U17713 ( .A(n14757), .Z(n14775) );
  XOR U17714 ( .A(n14783), .B(n14784), .Z(n14757) );
  ANDN U17715 ( .B(n14785), .A(n14786), .Z(n14783) );
  XOR U17716 ( .A(n14784), .B(n14787), .Z(n14785) );
  XOR U17717 ( .A(n14766), .B(n14697), .Z(n14767) );
  XOR U17718 ( .A(n14788), .B(n14789), .Z(n14697) );
  AND U17719 ( .A(n134), .B(n14790), .Z(n14788) );
  XOR U17720 ( .A(n14791), .B(n14789), .Z(n14790) );
  XNOR U17721 ( .A(n14792), .B(n14793), .Z(n14766) );
  NAND U17722 ( .A(n14794), .B(n14795), .Z(n14793) );
  XOR U17723 ( .A(n14796), .B(n14745), .Z(n14795) );
  XOR U17724 ( .A(n14786), .B(n14787), .Z(n14745) );
  XOR U17725 ( .A(n14797), .B(n14774), .Z(n14787) );
  XOR U17726 ( .A(n14798), .B(n14799), .Z(n14774) );
  ANDN U17727 ( .B(n14800), .A(n14801), .Z(n14798) );
  XOR U17728 ( .A(n14799), .B(n14802), .Z(n14800) );
  IV U17729 ( .A(n14772), .Z(n14797) );
  XOR U17730 ( .A(n14770), .B(n14803), .Z(n14772) );
  XOR U17731 ( .A(n14804), .B(n14805), .Z(n14803) );
  ANDN U17732 ( .B(n14806), .A(n14807), .Z(n14804) );
  XOR U17733 ( .A(n14808), .B(n14805), .Z(n14806) );
  IV U17734 ( .A(n14773), .Z(n14770) );
  XOR U17735 ( .A(n14809), .B(n14810), .Z(n14773) );
  ANDN U17736 ( .B(n14811), .A(n14812), .Z(n14809) );
  XOR U17737 ( .A(n14810), .B(n14813), .Z(n14811) );
  XOR U17738 ( .A(n14814), .B(n14815), .Z(n14786) );
  XNOR U17739 ( .A(n14781), .B(n14816), .Z(n14815) );
  IV U17740 ( .A(n14784), .Z(n14816) );
  XOR U17741 ( .A(n14817), .B(n14818), .Z(n14784) );
  ANDN U17742 ( .B(n14819), .A(n14820), .Z(n14817) );
  XOR U17743 ( .A(n14818), .B(n14821), .Z(n14819) );
  XNOR U17744 ( .A(n14822), .B(n14823), .Z(n14781) );
  ANDN U17745 ( .B(n14824), .A(n14825), .Z(n14822) );
  XOR U17746 ( .A(n14823), .B(n14826), .Z(n14824) );
  IV U17747 ( .A(n14780), .Z(n14814) );
  XOR U17748 ( .A(n14778), .B(n14827), .Z(n14780) );
  XOR U17749 ( .A(n14828), .B(n14829), .Z(n14827) );
  ANDN U17750 ( .B(n14830), .A(n14831), .Z(n14828) );
  XOR U17751 ( .A(n14832), .B(n14829), .Z(n14830) );
  IV U17752 ( .A(n14782), .Z(n14778) );
  XOR U17753 ( .A(n14833), .B(n14834), .Z(n14782) );
  ANDN U17754 ( .B(n14835), .A(n14836), .Z(n14833) );
  XOR U17755 ( .A(n14837), .B(n14834), .Z(n14835) );
  IV U17756 ( .A(n14792), .Z(n14796) );
  XOR U17757 ( .A(n14792), .B(n14747), .Z(n14794) );
  XOR U17758 ( .A(n14838), .B(n14839), .Z(n14747) );
  AND U17759 ( .A(n134), .B(n14840), .Z(n14838) );
  XOR U17760 ( .A(n14841), .B(n14839), .Z(n14840) );
  NANDN U17761 ( .A(n14749), .B(n14751), .Z(n14792) );
  XOR U17762 ( .A(n14842), .B(n14843), .Z(n14751) );
  AND U17763 ( .A(n134), .B(n14844), .Z(n14842) );
  XOR U17764 ( .A(n14843), .B(n14845), .Z(n14844) );
  XNOR U17765 ( .A(n14846), .B(n14847), .Z(n134) );
  AND U17766 ( .A(n14848), .B(n14849), .Z(n14846) );
  XOR U17767 ( .A(n14847), .B(n14762), .Z(n14849) );
  XNOR U17768 ( .A(n14850), .B(n14851), .Z(n14762) );
  ANDN U17769 ( .B(n14852), .A(n14853), .Z(n14850) );
  XOR U17770 ( .A(n14851), .B(n14854), .Z(n14852) );
  XNOR U17771 ( .A(n14847), .B(n14764), .Z(n14848) );
  XOR U17772 ( .A(n14855), .B(n14856), .Z(n14764) );
  AND U17773 ( .A(n138), .B(n14857), .Z(n14855) );
  XOR U17774 ( .A(n14858), .B(n14856), .Z(n14857) );
  XNOR U17775 ( .A(n14859), .B(n14860), .Z(n14847) );
  AND U17776 ( .A(n14861), .B(n14862), .Z(n14859) );
  XNOR U17777 ( .A(n14860), .B(n14789), .Z(n14862) );
  XOR U17778 ( .A(n14853), .B(n14854), .Z(n14789) );
  XNOR U17779 ( .A(n14863), .B(n14864), .Z(n14854) );
  ANDN U17780 ( .B(n14865), .A(n14866), .Z(n14863) );
  XOR U17781 ( .A(n14867), .B(n14868), .Z(n14865) );
  XOR U17782 ( .A(n14869), .B(n14870), .Z(n14853) );
  XNOR U17783 ( .A(n14871), .B(n14872), .Z(n14870) );
  ANDN U17784 ( .B(n14873), .A(n14874), .Z(n14871) );
  XNOR U17785 ( .A(n14875), .B(n14876), .Z(n14873) );
  IV U17786 ( .A(n14851), .Z(n14869) );
  XOR U17787 ( .A(n14877), .B(n14878), .Z(n14851) );
  ANDN U17788 ( .B(n14879), .A(n14880), .Z(n14877) );
  XOR U17789 ( .A(n14878), .B(n14881), .Z(n14879) );
  XOR U17790 ( .A(n14860), .B(n14791), .Z(n14861) );
  XOR U17791 ( .A(n14882), .B(n14883), .Z(n14791) );
  AND U17792 ( .A(n138), .B(n14884), .Z(n14882) );
  XOR U17793 ( .A(n14885), .B(n14883), .Z(n14884) );
  XNOR U17794 ( .A(n14886), .B(n14887), .Z(n14860) );
  NAND U17795 ( .A(n14888), .B(n14889), .Z(n14887) );
  XOR U17796 ( .A(n14890), .B(n14839), .Z(n14889) );
  XOR U17797 ( .A(n14880), .B(n14881), .Z(n14839) );
  XOR U17798 ( .A(n14891), .B(n14868), .Z(n14881) );
  XOR U17799 ( .A(n14892), .B(n14893), .Z(n14868) );
  ANDN U17800 ( .B(n14894), .A(n14895), .Z(n14892) );
  XOR U17801 ( .A(n14893), .B(n14896), .Z(n14894) );
  IV U17802 ( .A(n14866), .Z(n14891) );
  XOR U17803 ( .A(n14864), .B(n14897), .Z(n14866) );
  XOR U17804 ( .A(n14898), .B(n14899), .Z(n14897) );
  ANDN U17805 ( .B(n14900), .A(n14901), .Z(n14898) );
  XOR U17806 ( .A(n14902), .B(n14899), .Z(n14900) );
  IV U17807 ( .A(n14867), .Z(n14864) );
  XOR U17808 ( .A(n14903), .B(n14904), .Z(n14867) );
  ANDN U17809 ( .B(n14905), .A(n14906), .Z(n14903) );
  XOR U17810 ( .A(n14904), .B(n14907), .Z(n14905) );
  XOR U17811 ( .A(n14908), .B(n14909), .Z(n14880) );
  XNOR U17812 ( .A(n14875), .B(n14910), .Z(n14909) );
  IV U17813 ( .A(n14878), .Z(n14910) );
  XOR U17814 ( .A(n14911), .B(n14912), .Z(n14878) );
  ANDN U17815 ( .B(n14913), .A(n14914), .Z(n14911) );
  XOR U17816 ( .A(n14912), .B(n14915), .Z(n14913) );
  XNOR U17817 ( .A(n14916), .B(n14917), .Z(n14875) );
  ANDN U17818 ( .B(n14918), .A(n14919), .Z(n14916) );
  XOR U17819 ( .A(n14917), .B(n14920), .Z(n14918) );
  IV U17820 ( .A(n14874), .Z(n14908) );
  XOR U17821 ( .A(n14872), .B(n14921), .Z(n14874) );
  XOR U17822 ( .A(n14922), .B(n14923), .Z(n14921) );
  ANDN U17823 ( .B(n14924), .A(n14925), .Z(n14922) );
  XOR U17824 ( .A(n14926), .B(n14923), .Z(n14924) );
  IV U17825 ( .A(n14876), .Z(n14872) );
  XOR U17826 ( .A(n14927), .B(n14928), .Z(n14876) );
  ANDN U17827 ( .B(n14929), .A(n14930), .Z(n14927) );
  XOR U17828 ( .A(n14931), .B(n14928), .Z(n14929) );
  IV U17829 ( .A(n14886), .Z(n14890) );
  XOR U17830 ( .A(n14886), .B(n14841), .Z(n14888) );
  XOR U17831 ( .A(n14932), .B(n14933), .Z(n14841) );
  AND U17832 ( .A(n138), .B(n14934), .Z(n14932) );
  XOR U17833 ( .A(n14935), .B(n14933), .Z(n14934) );
  NANDN U17834 ( .A(n14843), .B(n14845), .Z(n14886) );
  XOR U17835 ( .A(n14936), .B(n14937), .Z(n14845) );
  AND U17836 ( .A(n138), .B(n14938), .Z(n14936) );
  XOR U17837 ( .A(n14937), .B(n14939), .Z(n14938) );
  XNOR U17838 ( .A(n14940), .B(n14941), .Z(n138) );
  AND U17839 ( .A(n14942), .B(n14943), .Z(n14940) );
  XOR U17840 ( .A(n14941), .B(n14856), .Z(n14943) );
  XNOR U17841 ( .A(n14944), .B(n14945), .Z(n14856) );
  ANDN U17842 ( .B(n14946), .A(n14947), .Z(n14944) );
  XOR U17843 ( .A(n14945), .B(n14948), .Z(n14946) );
  XNOR U17844 ( .A(n14941), .B(n14858), .Z(n14942) );
  XOR U17845 ( .A(n14949), .B(n14950), .Z(n14858) );
  AND U17846 ( .A(n142), .B(n14951), .Z(n14949) );
  XOR U17847 ( .A(n14952), .B(n14950), .Z(n14951) );
  XNOR U17848 ( .A(n14953), .B(n14954), .Z(n14941) );
  AND U17849 ( .A(n14955), .B(n14956), .Z(n14953) );
  XNOR U17850 ( .A(n14954), .B(n14883), .Z(n14956) );
  XOR U17851 ( .A(n14947), .B(n14948), .Z(n14883) );
  XNOR U17852 ( .A(n14957), .B(n14958), .Z(n14948) );
  ANDN U17853 ( .B(n14959), .A(n14960), .Z(n14957) );
  XOR U17854 ( .A(n14961), .B(n14962), .Z(n14959) );
  XOR U17855 ( .A(n14963), .B(n14964), .Z(n14947) );
  XNOR U17856 ( .A(n14965), .B(n14966), .Z(n14964) );
  ANDN U17857 ( .B(n14967), .A(n14968), .Z(n14965) );
  XNOR U17858 ( .A(n14969), .B(n14970), .Z(n14967) );
  IV U17859 ( .A(n14945), .Z(n14963) );
  XOR U17860 ( .A(n14971), .B(n14972), .Z(n14945) );
  ANDN U17861 ( .B(n14973), .A(n14974), .Z(n14971) );
  XOR U17862 ( .A(n14972), .B(n14975), .Z(n14973) );
  XOR U17863 ( .A(n14954), .B(n14885), .Z(n14955) );
  XOR U17864 ( .A(n14976), .B(n14977), .Z(n14885) );
  AND U17865 ( .A(n142), .B(n14978), .Z(n14976) );
  XOR U17866 ( .A(n14979), .B(n14977), .Z(n14978) );
  XNOR U17867 ( .A(n14980), .B(n14981), .Z(n14954) );
  NAND U17868 ( .A(n14982), .B(n14983), .Z(n14981) );
  XOR U17869 ( .A(n14984), .B(n14933), .Z(n14983) );
  XOR U17870 ( .A(n14974), .B(n14975), .Z(n14933) );
  XOR U17871 ( .A(n14985), .B(n14962), .Z(n14975) );
  XOR U17872 ( .A(n14986), .B(n14987), .Z(n14962) );
  ANDN U17873 ( .B(n14988), .A(n14989), .Z(n14986) );
  XOR U17874 ( .A(n14987), .B(n14990), .Z(n14988) );
  IV U17875 ( .A(n14960), .Z(n14985) );
  XOR U17876 ( .A(n14958), .B(n14991), .Z(n14960) );
  XOR U17877 ( .A(n14992), .B(n14993), .Z(n14991) );
  ANDN U17878 ( .B(n14994), .A(n14995), .Z(n14992) );
  XOR U17879 ( .A(n14996), .B(n14993), .Z(n14994) );
  IV U17880 ( .A(n14961), .Z(n14958) );
  XOR U17881 ( .A(n14997), .B(n14998), .Z(n14961) );
  ANDN U17882 ( .B(n14999), .A(n15000), .Z(n14997) );
  XOR U17883 ( .A(n14998), .B(n15001), .Z(n14999) );
  XOR U17884 ( .A(n15002), .B(n15003), .Z(n14974) );
  XNOR U17885 ( .A(n14969), .B(n15004), .Z(n15003) );
  IV U17886 ( .A(n14972), .Z(n15004) );
  XOR U17887 ( .A(n15005), .B(n15006), .Z(n14972) );
  ANDN U17888 ( .B(n15007), .A(n15008), .Z(n15005) );
  XOR U17889 ( .A(n15006), .B(n15009), .Z(n15007) );
  XNOR U17890 ( .A(n15010), .B(n15011), .Z(n14969) );
  ANDN U17891 ( .B(n15012), .A(n15013), .Z(n15010) );
  XOR U17892 ( .A(n15011), .B(n15014), .Z(n15012) );
  IV U17893 ( .A(n14968), .Z(n15002) );
  XOR U17894 ( .A(n14966), .B(n15015), .Z(n14968) );
  XOR U17895 ( .A(n15016), .B(n15017), .Z(n15015) );
  ANDN U17896 ( .B(n15018), .A(n15019), .Z(n15016) );
  XOR U17897 ( .A(n15020), .B(n15017), .Z(n15018) );
  IV U17898 ( .A(n14970), .Z(n14966) );
  XOR U17899 ( .A(n15021), .B(n15022), .Z(n14970) );
  ANDN U17900 ( .B(n15023), .A(n15024), .Z(n15021) );
  XOR U17901 ( .A(n15025), .B(n15022), .Z(n15023) );
  IV U17902 ( .A(n14980), .Z(n14984) );
  XOR U17903 ( .A(n14980), .B(n14935), .Z(n14982) );
  XOR U17904 ( .A(n15026), .B(n15027), .Z(n14935) );
  AND U17905 ( .A(n142), .B(n15028), .Z(n15026) );
  XOR U17906 ( .A(n15029), .B(n15027), .Z(n15028) );
  NANDN U17907 ( .A(n14937), .B(n14939), .Z(n14980) );
  XOR U17908 ( .A(n15030), .B(n15031), .Z(n14939) );
  AND U17909 ( .A(n142), .B(n15032), .Z(n15030) );
  XOR U17910 ( .A(n15031), .B(n15033), .Z(n15032) );
  XNOR U17911 ( .A(n15034), .B(n15035), .Z(n142) );
  AND U17912 ( .A(n15036), .B(n15037), .Z(n15034) );
  XOR U17913 ( .A(n15035), .B(n14950), .Z(n15037) );
  XNOR U17914 ( .A(n15038), .B(n15039), .Z(n14950) );
  ANDN U17915 ( .B(n15040), .A(n15041), .Z(n15038) );
  XOR U17916 ( .A(n15039), .B(n15042), .Z(n15040) );
  XNOR U17917 ( .A(n15035), .B(n14952), .Z(n15036) );
  XOR U17918 ( .A(n15043), .B(n15044), .Z(n14952) );
  AND U17919 ( .A(n146), .B(n15045), .Z(n15043) );
  XOR U17920 ( .A(n15046), .B(n15044), .Z(n15045) );
  XNOR U17921 ( .A(n15047), .B(n15048), .Z(n15035) );
  AND U17922 ( .A(n15049), .B(n15050), .Z(n15047) );
  XNOR U17923 ( .A(n15048), .B(n14977), .Z(n15050) );
  XOR U17924 ( .A(n15041), .B(n15042), .Z(n14977) );
  XNOR U17925 ( .A(n15051), .B(n15052), .Z(n15042) );
  ANDN U17926 ( .B(n15053), .A(n15054), .Z(n15051) );
  XOR U17927 ( .A(n15055), .B(n15056), .Z(n15053) );
  XOR U17928 ( .A(n15057), .B(n15058), .Z(n15041) );
  XNOR U17929 ( .A(n15059), .B(n15060), .Z(n15058) );
  ANDN U17930 ( .B(n15061), .A(n15062), .Z(n15059) );
  XNOR U17931 ( .A(n15063), .B(n15064), .Z(n15061) );
  IV U17932 ( .A(n15039), .Z(n15057) );
  XOR U17933 ( .A(n15065), .B(n15066), .Z(n15039) );
  ANDN U17934 ( .B(n15067), .A(n15068), .Z(n15065) );
  XOR U17935 ( .A(n15066), .B(n15069), .Z(n15067) );
  XOR U17936 ( .A(n15048), .B(n14979), .Z(n15049) );
  XOR U17937 ( .A(n15070), .B(n15071), .Z(n14979) );
  AND U17938 ( .A(n146), .B(n15072), .Z(n15070) );
  XOR U17939 ( .A(n15073), .B(n15071), .Z(n15072) );
  XNOR U17940 ( .A(n15074), .B(n15075), .Z(n15048) );
  NAND U17941 ( .A(n15076), .B(n15077), .Z(n15075) );
  XOR U17942 ( .A(n15078), .B(n15027), .Z(n15077) );
  XOR U17943 ( .A(n15068), .B(n15069), .Z(n15027) );
  XOR U17944 ( .A(n15079), .B(n15056), .Z(n15069) );
  XOR U17945 ( .A(n15080), .B(n15081), .Z(n15056) );
  ANDN U17946 ( .B(n15082), .A(n15083), .Z(n15080) );
  XOR U17947 ( .A(n15081), .B(n15084), .Z(n15082) );
  IV U17948 ( .A(n15054), .Z(n15079) );
  XOR U17949 ( .A(n15052), .B(n15085), .Z(n15054) );
  XOR U17950 ( .A(n15086), .B(n15087), .Z(n15085) );
  ANDN U17951 ( .B(n15088), .A(n15089), .Z(n15086) );
  XOR U17952 ( .A(n15090), .B(n15087), .Z(n15088) );
  IV U17953 ( .A(n15055), .Z(n15052) );
  XOR U17954 ( .A(n15091), .B(n15092), .Z(n15055) );
  ANDN U17955 ( .B(n15093), .A(n15094), .Z(n15091) );
  XOR U17956 ( .A(n15092), .B(n15095), .Z(n15093) );
  XOR U17957 ( .A(n15096), .B(n15097), .Z(n15068) );
  XNOR U17958 ( .A(n15063), .B(n15098), .Z(n15097) );
  IV U17959 ( .A(n15066), .Z(n15098) );
  XOR U17960 ( .A(n15099), .B(n15100), .Z(n15066) );
  ANDN U17961 ( .B(n15101), .A(n15102), .Z(n15099) );
  XOR U17962 ( .A(n15100), .B(n15103), .Z(n15101) );
  XNOR U17963 ( .A(n15104), .B(n15105), .Z(n15063) );
  ANDN U17964 ( .B(n15106), .A(n15107), .Z(n15104) );
  XOR U17965 ( .A(n15105), .B(n15108), .Z(n15106) );
  IV U17966 ( .A(n15062), .Z(n15096) );
  XOR U17967 ( .A(n15060), .B(n15109), .Z(n15062) );
  XOR U17968 ( .A(n15110), .B(n15111), .Z(n15109) );
  ANDN U17969 ( .B(n15112), .A(n15113), .Z(n15110) );
  XOR U17970 ( .A(n15114), .B(n15111), .Z(n15112) );
  IV U17971 ( .A(n15064), .Z(n15060) );
  XOR U17972 ( .A(n15115), .B(n15116), .Z(n15064) );
  ANDN U17973 ( .B(n15117), .A(n15118), .Z(n15115) );
  XOR U17974 ( .A(n15119), .B(n15116), .Z(n15117) );
  IV U17975 ( .A(n15074), .Z(n15078) );
  XOR U17976 ( .A(n15074), .B(n15029), .Z(n15076) );
  XOR U17977 ( .A(n15120), .B(n15121), .Z(n15029) );
  AND U17978 ( .A(n146), .B(n15122), .Z(n15120) );
  XOR U17979 ( .A(n15123), .B(n15121), .Z(n15122) );
  NANDN U17980 ( .A(n15031), .B(n15033), .Z(n15074) );
  XOR U17981 ( .A(n15124), .B(n15125), .Z(n15033) );
  AND U17982 ( .A(n146), .B(n15126), .Z(n15124) );
  XOR U17983 ( .A(n15125), .B(n15127), .Z(n15126) );
  XNOR U17984 ( .A(n15128), .B(n15129), .Z(n146) );
  AND U17985 ( .A(n15130), .B(n15131), .Z(n15128) );
  XOR U17986 ( .A(n15129), .B(n15044), .Z(n15131) );
  XNOR U17987 ( .A(n15132), .B(n15133), .Z(n15044) );
  ANDN U17988 ( .B(n15134), .A(n15135), .Z(n15132) );
  XOR U17989 ( .A(n15133), .B(n15136), .Z(n15134) );
  XNOR U17990 ( .A(n15129), .B(n15046), .Z(n15130) );
  XOR U17991 ( .A(n15137), .B(n15138), .Z(n15046) );
  AND U17992 ( .A(n150), .B(n15139), .Z(n15137) );
  XOR U17993 ( .A(n15140), .B(n15138), .Z(n15139) );
  XNOR U17994 ( .A(n15141), .B(n15142), .Z(n15129) );
  AND U17995 ( .A(n15143), .B(n15144), .Z(n15141) );
  XNOR U17996 ( .A(n15142), .B(n15071), .Z(n15144) );
  XOR U17997 ( .A(n15135), .B(n15136), .Z(n15071) );
  XNOR U17998 ( .A(n15145), .B(n15146), .Z(n15136) );
  ANDN U17999 ( .B(n15147), .A(n15148), .Z(n15145) );
  XOR U18000 ( .A(n15149), .B(n15150), .Z(n15147) );
  XOR U18001 ( .A(n15151), .B(n15152), .Z(n15135) );
  XNOR U18002 ( .A(n15153), .B(n15154), .Z(n15152) );
  ANDN U18003 ( .B(n15155), .A(n15156), .Z(n15153) );
  XNOR U18004 ( .A(n15157), .B(n15158), .Z(n15155) );
  IV U18005 ( .A(n15133), .Z(n15151) );
  XOR U18006 ( .A(n15159), .B(n15160), .Z(n15133) );
  ANDN U18007 ( .B(n15161), .A(n15162), .Z(n15159) );
  XOR U18008 ( .A(n15160), .B(n15163), .Z(n15161) );
  XOR U18009 ( .A(n15142), .B(n15073), .Z(n15143) );
  XOR U18010 ( .A(n15164), .B(n15165), .Z(n15073) );
  AND U18011 ( .A(n150), .B(n15166), .Z(n15164) );
  XOR U18012 ( .A(n15167), .B(n15165), .Z(n15166) );
  XNOR U18013 ( .A(n15168), .B(n15169), .Z(n15142) );
  NAND U18014 ( .A(n15170), .B(n15171), .Z(n15169) );
  XOR U18015 ( .A(n15172), .B(n15121), .Z(n15171) );
  XOR U18016 ( .A(n15162), .B(n15163), .Z(n15121) );
  XOR U18017 ( .A(n15173), .B(n15150), .Z(n15163) );
  XOR U18018 ( .A(n15174), .B(n15175), .Z(n15150) );
  ANDN U18019 ( .B(n15176), .A(n15177), .Z(n15174) );
  XOR U18020 ( .A(n15175), .B(n15178), .Z(n15176) );
  IV U18021 ( .A(n15148), .Z(n15173) );
  XOR U18022 ( .A(n15146), .B(n15179), .Z(n15148) );
  XOR U18023 ( .A(n15180), .B(n15181), .Z(n15179) );
  ANDN U18024 ( .B(n15182), .A(n15183), .Z(n15180) );
  XOR U18025 ( .A(n15184), .B(n15181), .Z(n15182) );
  IV U18026 ( .A(n15149), .Z(n15146) );
  XOR U18027 ( .A(n15185), .B(n15186), .Z(n15149) );
  ANDN U18028 ( .B(n15187), .A(n15188), .Z(n15185) );
  XOR U18029 ( .A(n15186), .B(n15189), .Z(n15187) );
  XOR U18030 ( .A(n15190), .B(n15191), .Z(n15162) );
  XNOR U18031 ( .A(n15157), .B(n15192), .Z(n15191) );
  IV U18032 ( .A(n15160), .Z(n15192) );
  XOR U18033 ( .A(n15193), .B(n15194), .Z(n15160) );
  ANDN U18034 ( .B(n15195), .A(n15196), .Z(n15193) );
  XOR U18035 ( .A(n15194), .B(n15197), .Z(n15195) );
  XNOR U18036 ( .A(n15198), .B(n15199), .Z(n15157) );
  ANDN U18037 ( .B(n15200), .A(n15201), .Z(n15198) );
  XOR U18038 ( .A(n15199), .B(n15202), .Z(n15200) );
  IV U18039 ( .A(n15156), .Z(n15190) );
  XOR U18040 ( .A(n15154), .B(n15203), .Z(n15156) );
  XOR U18041 ( .A(n15204), .B(n15205), .Z(n15203) );
  ANDN U18042 ( .B(n15206), .A(n15207), .Z(n15204) );
  XOR U18043 ( .A(n15208), .B(n15205), .Z(n15206) );
  IV U18044 ( .A(n15158), .Z(n15154) );
  XOR U18045 ( .A(n15209), .B(n15210), .Z(n15158) );
  ANDN U18046 ( .B(n15211), .A(n15212), .Z(n15209) );
  XOR U18047 ( .A(n15213), .B(n15210), .Z(n15211) );
  IV U18048 ( .A(n15168), .Z(n15172) );
  XOR U18049 ( .A(n15168), .B(n15123), .Z(n15170) );
  XOR U18050 ( .A(n15214), .B(n15215), .Z(n15123) );
  AND U18051 ( .A(n150), .B(n15216), .Z(n15214) );
  XOR U18052 ( .A(n15217), .B(n15215), .Z(n15216) );
  NANDN U18053 ( .A(n15125), .B(n15127), .Z(n15168) );
  XOR U18054 ( .A(n15218), .B(n15219), .Z(n15127) );
  AND U18055 ( .A(n150), .B(n15220), .Z(n15218) );
  XOR U18056 ( .A(n15219), .B(n15221), .Z(n15220) );
  XNOR U18057 ( .A(n15222), .B(n15223), .Z(n150) );
  AND U18058 ( .A(n15224), .B(n15225), .Z(n15222) );
  XOR U18059 ( .A(n15223), .B(n15138), .Z(n15225) );
  XNOR U18060 ( .A(n15226), .B(n15227), .Z(n15138) );
  ANDN U18061 ( .B(n15228), .A(n15229), .Z(n15226) );
  XOR U18062 ( .A(n15227), .B(n15230), .Z(n15228) );
  XNOR U18063 ( .A(n15223), .B(n15140), .Z(n15224) );
  XOR U18064 ( .A(n15231), .B(n15232), .Z(n15140) );
  AND U18065 ( .A(n154), .B(n15233), .Z(n15231) );
  XOR U18066 ( .A(n15234), .B(n15232), .Z(n15233) );
  XNOR U18067 ( .A(n15235), .B(n15236), .Z(n15223) );
  AND U18068 ( .A(n15237), .B(n15238), .Z(n15235) );
  XNOR U18069 ( .A(n15236), .B(n15165), .Z(n15238) );
  XOR U18070 ( .A(n15229), .B(n15230), .Z(n15165) );
  XNOR U18071 ( .A(n15239), .B(n15240), .Z(n15230) );
  ANDN U18072 ( .B(n15241), .A(n15242), .Z(n15239) );
  XOR U18073 ( .A(n15243), .B(n15244), .Z(n15241) );
  XOR U18074 ( .A(n15245), .B(n15246), .Z(n15229) );
  XNOR U18075 ( .A(n15247), .B(n15248), .Z(n15246) );
  ANDN U18076 ( .B(n15249), .A(n15250), .Z(n15247) );
  XNOR U18077 ( .A(n15251), .B(n15252), .Z(n15249) );
  IV U18078 ( .A(n15227), .Z(n15245) );
  XOR U18079 ( .A(n15253), .B(n15254), .Z(n15227) );
  ANDN U18080 ( .B(n15255), .A(n15256), .Z(n15253) );
  XOR U18081 ( .A(n15254), .B(n15257), .Z(n15255) );
  XOR U18082 ( .A(n15236), .B(n15167), .Z(n15237) );
  XOR U18083 ( .A(n15258), .B(n15259), .Z(n15167) );
  AND U18084 ( .A(n154), .B(n15260), .Z(n15258) );
  XOR U18085 ( .A(n15261), .B(n15259), .Z(n15260) );
  XNOR U18086 ( .A(n15262), .B(n15263), .Z(n15236) );
  NAND U18087 ( .A(n15264), .B(n15265), .Z(n15263) );
  XOR U18088 ( .A(n15266), .B(n15215), .Z(n15265) );
  XOR U18089 ( .A(n15256), .B(n15257), .Z(n15215) );
  XOR U18090 ( .A(n15267), .B(n15244), .Z(n15257) );
  XOR U18091 ( .A(n15268), .B(n15269), .Z(n15244) );
  ANDN U18092 ( .B(n15270), .A(n15271), .Z(n15268) );
  XOR U18093 ( .A(n15269), .B(n15272), .Z(n15270) );
  IV U18094 ( .A(n15242), .Z(n15267) );
  XOR U18095 ( .A(n15240), .B(n15273), .Z(n15242) );
  XOR U18096 ( .A(n15274), .B(n15275), .Z(n15273) );
  ANDN U18097 ( .B(n15276), .A(n15277), .Z(n15274) );
  XOR U18098 ( .A(n15278), .B(n15275), .Z(n15276) );
  IV U18099 ( .A(n15243), .Z(n15240) );
  XOR U18100 ( .A(n15279), .B(n15280), .Z(n15243) );
  ANDN U18101 ( .B(n15281), .A(n15282), .Z(n15279) );
  XOR U18102 ( .A(n15280), .B(n15283), .Z(n15281) );
  XOR U18103 ( .A(n15284), .B(n15285), .Z(n15256) );
  XNOR U18104 ( .A(n15251), .B(n15286), .Z(n15285) );
  IV U18105 ( .A(n15254), .Z(n15286) );
  XOR U18106 ( .A(n15287), .B(n15288), .Z(n15254) );
  ANDN U18107 ( .B(n15289), .A(n15290), .Z(n15287) );
  XOR U18108 ( .A(n15288), .B(n15291), .Z(n15289) );
  XNOR U18109 ( .A(n15292), .B(n15293), .Z(n15251) );
  ANDN U18110 ( .B(n15294), .A(n15295), .Z(n15292) );
  XOR U18111 ( .A(n15293), .B(n15296), .Z(n15294) );
  IV U18112 ( .A(n15250), .Z(n15284) );
  XOR U18113 ( .A(n15248), .B(n15297), .Z(n15250) );
  XOR U18114 ( .A(n15298), .B(n15299), .Z(n15297) );
  ANDN U18115 ( .B(n15300), .A(n15301), .Z(n15298) );
  XOR U18116 ( .A(n15302), .B(n15299), .Z(n15300) );
  IV U18117 ( .A(n15252), .Z(n15248) );
  XOR U18118 ( .A(n15303), .B(n15304), .Z(n15252) );
  ANDN U18119 ( .B(n15305), .A(n15306), .Z(n15303) );
  XOR U18120 ( .A(n15307), .B(n15304), .Z(n15305) );
  IV U18121 ( .A(n15262), .Z(n15266) );
  XOR U18122 ( .A(n15262), .B(n15217), .Z(n15264) );
  XOR U18123 ( .A(n15308), .B(n15309), .Z(n15217) );
  AND U18124 ( .A(n154), .B(n15310), .Z(n15308) );
  XOR U18125 ( .A(n15311), .B(n15309), .Z(n15310) );
  NANDN U18126 ( .A(n15219), .B(n15221), .Z(n15262) );
  XOR U18127 ( .A(n15312), .B(n15313), .Z(n15221) );
  AND U18128 ( .A(n154), .B(n15314), .Z(n15312) );
  XOR U18129 ( .A(n15313), .B(n15315), .Z(n15314) );
  XNOR U18130 ( .A(n15316), .B(n15317), .Z(n154) );
  AND U18131 ( .A(n15318), .B(n15319), .Z(n15316) );
  XOR U18132 ( .A(n15317), .B(n15232), .Z(n15319) );
  XNOR U18133 ( .A(n15320), .B(n15321), .Z(n15232) );
  ANDN U18134 ( .B(n15322), .A(n15323), .Z(n15320) );
  XOR U18135 ( .A(n15321), .B(n15324), .Z(n15322) );
  XNOR U18136 ( .A(n15317), .B(n15234), .Z(n15318) );
  XOR U18137 ( .A(n15325), .B(n15326), .Z(n15234) );
  AND U18138 ( .A(n158), .B(n15327), .Z(n15325) );
  XOR U18139 ( .A(n15328), .B(n15326), .Z(n15327) );
  XNOR U18140 ( .A(n15329), .B(n15330), .Z(n15317) );
  AND U18141 ( .A(n15331), .B(n15332), .Z(n15329) );
  XNOR U18142 ( .A(n15330), .B(n15259), .Z(n15332) );
  XOR U18143 ( .A(n15323), .B(n15324), .Z(n15259) );
  XNOR U18144 ( .A(n15333), .B(n15334), .Z(n15324) );
  ANDN U18145 ( .B(n15335), .A(n15336), .Z(n15333) );
  XOR U18146 ( .A(n15337), .B(n15338), .Z(n15335) );
  XOR U18147 ( .A(n15339), .B(n15340), .Z(n15323) );
  XNOR U18148 ( .A(n15341), .B(n15342), .Z(n15340) );
  ANDN U18149 ( .B(n15343), .A(n15344), .Z(n15341) );
  XNOR U18150 ( .A(n15345), .B(n15346), .Z(n15343) );
  IV U18151 ( .A(n15321), .Z(n15339) );
  XOR U18152 ( .A(n15347), .B(n15348), .Z(n15321) );
  ANDN U18153 ( .B(n15349), .A(n15350), .Z(n15347) );
  XOR U18154 ( .A(n15348), .B(n15351), .Z(n15349) );
  XOR U18155 ( .A(n15330), .B(n15261), .Z(n15331) );
  XOR U18156 ( .A(n15352), .B(n15353), .Z(n15261) );
  AND U18157 ( .A(n158), .B(n15354), .Z(n15352) );
  XOR U18158 ( .A(n15355), .B(n15353), .Z(n15354) );
  XNOR U18159 ( .A(n15356), .B(n15357), .Z(n15330) );
  NAND U18160 ( .A(n15358), .B(n15359), .Z(n15357) );
  XOR U18161 ( .A(n15360), .B(n15309), .Z(n15359) );
  XOR U18162 ( .A(n15350), .B(n15351), .Z(n15309) );
  XOR U18163 ( .A(n15361), .B(n15338), .Z(n15351) );
  XOR U18164 ( .A(n15362), .B(n15363), .Z(n15338) );
  ANDN U18165 ( .B(n15364), .A(n15365), .Z(n15362) );
  XOR U18166 ( .A(n15363), .B(n15366), .Z(n15364) );
  IV U18167 ( .A(n15336), .Z(n15361) );
  XOR U18168 ( .A(n15334), .B(n15367), .Z(n15336) );
  XOR U18169 ( .A(n15368), .B(n15369), .Z(n15367) );
  ANDN U18170 ( .B(n15370), .A(n15371), .Z(n15368) );
  XOR U18171 ( .A(n15372), .B(n15369), .Z(n15370) );
  IV U18172 ( .A(n15337), .Z(n15334) );
  XOR U18173 ( .A(n15373), .B(n15374), .Z(n15337) );
  ANDN U18174 ( .B(n15375), .A(n15376), .Z(n15373) );
  XOR U18175 ( .A(n15374), .B(n15377), .Z(n15375) );
  XOR U18176 ( .A(n15378), .B(n15379), .Z(n15350) );
  XNOR U18177 ( .A(n15345), .B(n15380), .Z(n15379) );
  IV U18178 ( .A(n15348), .Z(n15380) );
  XOR U18179 ( .A(n15381), .B(n15382), .Z(n15348) );
  ANDN U18180 ( .B(n15383), .A(n15384), .Z(n15381) );
  XOR U18181 ( .A(n15382), .B(n15385), .Z(n15383) );
  XNOR U18182 ( .A(n15386), .B(n15387), .Z(n15345) );
  ANDN U18183 ( .B(n15388), .A(n15389), .Z(n15386) );
  XOR U18184 ( .A(n15387), .B(n15390), .Z(n15388) );
  IV U18185 ( .A(n15344), .Z(n15378) );
  XOR U18186 ( .A(n15342), .B(n15391), .Z(n15344) );
  XOR U18187 ( .A(n15392), .B(n15393), .Z(n15391) );
  ANDN U18188 ( .B(n15394), .A(n15395), .Z(n15392) );
  XOR U18189 ( .A(n15396), .B(n15393), .Z(n15394) );
  IV U18190 ( .A(n15346), .Z(n15342) );
  XOR U18191 ( .A(n15397), .B(n15398), .Z(n15346) );
  ANDN U18192 ( .B(n15399), .A(n15400), .Z(n15397) );
  XOR U18193 ( .A(n15401), .B(n15398), .Z(n15399) );
  IV U18194 ( .A(n15356), .Z(n15360) );
  XOR U18195 ( .A(n15356), .B(n15311), .Z(n15358) );
  XOR U18196 ( .A(n15402), .B(n15403), .Z(n15311) );
  AND U18197 ( .A(n158), .B(n15404), .Z(n15402) );
  XOR U18198 ( .A(n15405), .B(n15403), .Z(n15404) );
  NANDN U18199 ( .A(n15313), .B(n15315), .Z(n15356) );
  XOR U18200 ( .A(n15406), .B(n15407), .Z(n15315) );
  AND U18201 ( .A(n158), .B(n15408), .Z(n15406) );
  XOR U18202 ( .A(n15407), .B(n15409), .Z(n15408) );
  XNOR U18203 ( .A(n15410), .B(n15411), .Z(n158) );
  AND U18204 ( .A(n15412), .B(n15413), .Z(n15410) );
  XOR U18205 ( .A(n15411), .B(n15326), .Z(n15413) );
  XNOR U18206 ( .A(n15414), .B(n15415), .Z(n15326) );
  ANDN U18207 ( .B(n15416), .A(n15417), .Z(n15414) );
  XOR U18208 ( .A(n15415), .B(n15418), .Z(n15416) );
  XNOR U18209 ( .A(n15411), .B(n15328), .Z(n15412) );
  XOR U18210 ( .A(n15419), .B(n15420), .Z(n15328) );
  AND U18211 ( .A(n162), .B(n15421), .Z(n15419) );
  XOR U18212 ( .A(n15422), .B(n15420), .Z(n15421) );
  XNOR U18213 ( .A(n15423), .B(n15424), .Z(n15411) );
  AND U18214 ( .A(n15425), .B(n15426), .Z(n15423) );
  XNOR U18215 ( .A(n15424), .B(n15353), .Z(n15426) );
  XOR U18216 ( .A(n15417), .B(n15418), .Z(n15353) );
  XNOR U18217 ( .A(n15427), .B(n15428), .Z(n15418) );
  ANDN U18218 ( .B(n15429), .A(n15430), .Z(n15427) );
  XOR U18219 ( .A(n15431), .B(n15432), .Z(n15429) );
  XOR U18220 ( .A(n15433), .B(n15434), .Z(n15417) );
  XNOR U18221 ( .A(n15435), .B(n15436), .Z(n15434) );
  ANDN U18222 ( .B(n15437), .A(n15438), .Z(n15435) );
  XNOR U18223 ( .A(n15439), .B(n15440), .Z(n15437) );
  IV U18224 ( .A(n15415), .Z(n15433) );
  XOR U18225 ( .A(n15441), .B(n15442), .Z(n15415) );
  ANDN U18226 ( .B(n15443), .A(n15444), .Z(n15441) );
  XOR U18227 ( .A(n15442), .B(n15445), .Z(n15443) );
  XOR U18228 ( .A(n15424), .B(n15355), .Z(n15425) );
  XOR U18229 ( .A(n15446), .B(n15447), .Z(n15355) );
  AND U18230 ( .A(n162), .B(n15448), .Z(n15446) );
  XOR U18231 ( .A(n15449), .B(n15447), .Z(n15448) );
  XNOR U18232 ( .A(n15450), .B(n15451), .Z(n15424) );
  NAND U18233 ( .A(n15452), .B(n15453), .Z(n15451) );
  XOR U18234 ( .A(n15454), .B(n15403), .Z(n15453) );
  XOR U18235 ( .A(n15444), .B(n15445), .Z(n15403) );
  XOR U18236 ( .A(n15455), .B(n15432), .Z(n15445) );
  XOR U18237 ( .A(n15456), .B(n15457), .Z(n15432) );
  ANDN U18238 ( .B(n15458), .A(n15459), .Z(n15456) );
  XOR U18239 ( .A(n15457), .B(n15460), .Z(n15458) );
  IV U18240 ( .A(n15430), .Z(n15455) );
  XOR U18241 ( .A(n15428), .B(n15461), .Z(n15430) );
  XOR U18242 ( .A(n15462), .B(n15463), .Z(n15461) );
  ANDN U18243 ( .B(n15464), .A(n15465), .Z(n15462) );
  XOR U18244 ( .A(n15466), .B(n15463), .Z(n15464) );
  IV U18245 ( .A(n15431), .Z(n15428) );
  XOR U18246 ( .A(n15467), .B(n15468), .Z(n15431) );
  ANDN U18247 ( .B(n15469), .A(n15470), .Z(n15467) );
  XOR U18248 ( .A(n15468), .B(n15471), .Z(n15469) );
  XOR U18249 ( .A(n15472), .B(n15473), .Z(n15444) );
  XNOR U18250 ( .A(n15439), .B(n15474), .Z(n15473) );
  IV U18251 ( .A(n15442), .Z(n15474) );
  XOR U18252 ( .A(n15475), .B(n15476), .Z(n15442) );
  ANDN U18253 ( .B(n15477), .A(n15478), .Z(n15475) );
  XOR U18254 ( .A(n15476), .B(n15479), .Z(n15477) );
  XNOR U18255 ( .A(n15480), .B(n15481), .Z(n15439) );
  ANDN U18256 ( .B(n15482), .A(n15483), .Z(n15480) );
  XOR U18257 ( .A(n15481), .B(n15484), .Z(n15482) );
  IV U18258 ( .A(n15438), .Z(n15472) );
  XOR U18259 ( .A(n15436), .B(n15485), .Z(n15438) );
  XOR U18260 ( .A(n15486), .B(n15487), .Z(n15485) );
  ANDN U18261 ( .B(n15488), .A(n15489), .Z(n15486) );
  XOR U18262 ( .A(n15490), .B(n15487), .Z(n15488) );
  IV U18263 ( .A(n15440), .Z(n15436) );
  XOR U18264 ( .A(n15491), .B(n15492), .Z(n15440) );
  ANDN U18265 ( .B(n15493), .A(n15494), .Z(n15491) );
  XOR U18266 ( .A(n15495), .B(n15492), .Z(n15493) );
  IV U18267 ( .A(n15450), .Z(n15454) );
  XOR U18268 ( .A(n15450), .B(n15405), .Z(n15452) );
  XOR U18269 ( .A(n15496), .B(n15497), .Z(n15405) );
  AND U18270 ( .A(n162), .B(n15498), .Z(n15496) );
  XOR U18271 ( .A(n15499), .B(n15497), .Z(n15498) );
  NANDN U18272 ( .A(n15407), .B(n15409), .Z(n15450) );
  XOR U18273 ( .A(n15500), .B(n15501), .Z(n15409) );
  AND U18274 ( .A(n162), .B(n15502), .Z(n15500) );
  XOR U18275 ( .A(n15501), .B(n15503), .Z(n15502) );
  XNOR U18276 ( .A(n15504), .B(n15505), .Z(n162) );
  AND U18277 ( .A(n15506), .B(n15507), .Z(n15504) );
  XOR U18278 ( .A(n15505), .B(n15420), .Z(n15507) );
  XNOR U18279 ( .A(n15508), .B(n15509), .Z(n15420) );
  ANDN U18280 ( .B(n15510), .A(n15511), .Z(n15508) );
  XOR U18281 ( .A(n15509), .B(n15512), .Z(n15510) );
  XNOR U18282 ( .A(n15505), .B(n15422), .Z(n15506) );
  XOR U18283 ( .A(n15513), .B(n15514), .Z(n15422) );
  AND U18284 ( .A(n166), .B(n15515), .Z(n15513) );
  XOR U18285 ( .A(n15516), .B(n15514), .Z(n15515) );
  XNOR U18286 ( .A(n15517), .B(n15518), .Z(n15505) );
  AND U18287 ( .A(n15519), .B(n15520), .Z(n15517) );
  XNOR U18288 ( .A(n15518), .B(n15447), .Z(n15520) );
  XOR U18289 ( .A(n15511), .B(n15512), .Z(n15447) );
  XNOR U18290 ( .A(n15521), .B(n15522), .Z(n15512) );
  ANDN U18291 ( .B(n15523), .A(n15524), .Z(n15521) );
  XOR U18292 ( .A(n15525), .B(n15526), .Z(n15523) );
  XOR U18293 ( .A(n15527), .B(n15528), .Z(n15511) );
  XNOR U18294 ( .A(n15529), .B(n15530), .Z(n15528) );
  ANDN U18295 ( .B(n15531), .A(n15532), .Z(n15529) );
  XNOR U18296 ( .A(n15533), .B(n15534), .Z(n15531) );
  IV U18297 ( .A(n15509), .Z(n15527) );
  XOR U18298 ( .A(n15535), .B(n15536), .Z(n15509) );
  ANDN U18299 ( .B(n15537), .A(n15538), .Z(n15535) );
  XOR U18300 ( .A(n15536), .B(n15539), .Z(n15537) );
  XOR U18301 ( .A(n15518), .B(n15449), .Z(n15519) );
  XOR U18302 ( .A(n15540), .B(n15541), .Z(n15449) );
  AND U18303 ( .A(n166), .B(n15542), .Z(n15540) );
  XOR U18304 ( .A(n15543), .B(n15541), .Z(n15542) );
  XNOR U18305 ( .A(n15544), .B(n15545), .Z(n15518) );
  NAND U18306 ( .A(n15546), .B(n15547), .Z(n15545) );
  XOR U18307 ( .A(n15548), .B(n15497), .Z(n15547) );
  XOR U18308 ( .A(n15538), .B(n15539), .Z(n15497) );
  XOR U18309 ( .A(n15549), .B(n15526), .Z(n15539) );
  XOR U18310 ( .A(n15550), .B(n15551), .Z(n15526) );
  ANDN U18311 ( .B(n15552), .A(n15553), .Z(n15550) );
  XOR U18312 ( .A(n15551), .B(n15554), .Z(n15552) );
  IV U18313 ( .A(n15524), .Z(n15549) );
  XOR U18314 ( .A(n15522), .B(n15555), .Z(n15524) );
  XOR U18315 ( .A(n15556), .B(n15557), .Z(n15555) );
  ANDN U18316 ( .B(n15558), .A(n15559), .Z(n15556) );
  XOR U18317 ( .A(n15560), .B(n15557), .Z(n15558) );
  IV U18318 ( .A(n15525), .Z(n15522) );
  XOR U18319 ( .A(n15561), .B(n15562), .Z(n15525) );
  ANDN U18320 ( .B(n15563), .A(n15564), .Z(n15561) );
  XOR U18321 ( .A(n15562), .B(n15565), .Z(n15563) );
  XOR U18322 ( .A(n15566), .B(n15567), .Z(n15538) );
  XNOR U18323 ( .A(n15533), .B(n15568), .Z(n15567) );
  IV U18324 ( .A(n15536), .Z(n15568) );
  XOR U18325 ( .A(n15569), .B(n15570), .Z(n15536) );
  ANDN U18326 ( .B(n15571), .A(n15572), .Z(n15569) );
  XOR U18327 ( .A(n15570), .B(n15573), .Z(n15571) );
  XNOR U18328 ( .A(n15574), .B(n15575), .Z(n15533) );
  ANDN U18329 ( .B(n15576), .A(n15577), .Z(n15574) );
  XOR U18330 ( .A(n15575), .B(n15578), .Z(n15576) );
  IV U18331 ( .A(n15532), .Z(n15566) );
  XOR U18332 ( .A(n15530), .B(n15579), .Z(n15532) );
  XOR U18333 ( .A(n15580), .B(n15581), .Z(n15579) );
  ANDN U18334 ( .B(n15582), .A(n15583), .Z(n15580) );
  XOR U18335 ( .A(n15584), .B(n15581), .Z(n15582) );
  IV U18336 ( .A(n15534), .Z(n15530) );
  XOR U18337 ( .A(n15585), .B(n15586), .Z(n15534) );
  ANDN U18338 ( .B(n15587), .A(n15588), .Z(n15585) );
  XOR U18339 ( .A(n15589), .B(n15586), .Z(n15587) );
  IV U18340 ( .A(n15544), .Z(n15548) );
  XOR U18341 ( .A(n15544), .B(n15499), .Z(n15546) );
  XOR U18342 ( .A(n15590), .B(n15591), .Z(n15499) );
  AND U18343 ( .A(n166), .B(n15592), .Z(n15590) );
  XOR U18344 ( .A(n15593), .B(n15591), .Z(n15592) );
  NANDN U18345 ( .A(n15501), .B(n15503), .Z(n15544) );
  XOR U18346 ( .A(n15594), .B(n15595), .Z(n15503) );
  AND U18347 ( .A(n166), .B(n15596), .Z(n15594) );
  XOR U18348 ( .A(n15595), .B(n15597), .Z(n15596) );
  XNOR U18349 ( .A(n15598), .B(n15599), .Z(n166) );
  AND U18350 ( .A(n15600), .B(n15601), .Z(n15598) );
  XOR U18351 ( .A(n15599), .B(n15514), .Z(n15601) );
  XNOR U18352 ( .A(n15602), .B(n15603), .Z(n15514) );
  ANDN U18353 ( .B(n15604), .A(n15605), .Z(n15602) );
  XOR U18354 ( .A(n15603), .B(n15606), .Z(n15604) );
  XNOR U18355 ( .A(n15599), .B(n15516), .Z(n15600) );
  XOR U18356 ( .A(n15607), .B(n15608), .Z(n15516) );
  AND U18357 ( .A(n170), .B(n15609), .Z(n15607) );
  XOR U18358 ( .A(n15610), .B(n15608), .Z(n15609) );
  XNOR U18359 ( .A(n15611), .B(n15612), .Z(n15599) );
  AND U18360 ( .A(n15613), .B(n15614), .Z(n15611) );
  XNOR U18361 ( .A(n15612), .B(n15541), .Z(n15614) );
  XOR U18362 ( .A(n15605), .B(n15606), .Z(n15541) );
  XNOR U18363 ( .A(n15615), .B(n15616), .Z(n15606) );
  ANDN U18364 ( .B(n15617), .A(n15618), .Z(n15615) );
  XOR U18365 ( .A(n15619), .B(n15620), .Z(n15617) );
  XOR U18366 ( .A(n15621), .B(n15622), .Z(n15605) );
  XNOR U18367 ( .A(n15623), .B(n15624), .Z(n15622) );
  ANDN U18368 ( .B(n15625), .A(n15626), .Z(n15623) );
  XNOR U18369 ( .A(n15627), .B(n15628), .Z(n15625) );
  IV U18370 ( .A(n15603), .Z(n15621) );
  XOR U18371 ( .A(n15629), .B(n15630), .Z(n15603) );
  ANDN U18372 ( .B(n15631), .A(n15632), .Z(n15629) );
  XOR U18373 ( .A(n15630), .B(n15633), .Z(n15631) );
  XOR U18374 ( .A(n15612), .B(n15543), .Z(n15613) );
  XOR U18375 ( .A(n15634), .B(n15635), .Z(n15543) );
  AND U18376 ( .A(n170), .B(n15636), .Z(n15634) );
  XOR U18377 ( .A(n15637), .B(n15635), .Z(n15636) );
  XNOR U18378 ( .A(n15638), .B(n15639), .Z(n15612) );
  NAND U18379 ( .A(n15640), .B(n15641), .Z(n15639) );
  XOR U18380 ( .A(n15642), .B(n15591), .Z(n15641) );
  XOR U18381 ( .A(n15632), .B(n15633), .Z(n15591) );
  XOR U18382 ( .A(n15643), .B(n15620), .Z(n15633) );
  XOR U18383 ( .A(n15644), .B(n15645), .Z(n15620) );
  ANDN U18384 ( .B(n15646), .A(n15647), .Z(n15644) );
  XOR U18385 ( .A(n15645), .B(n15648), .Z(n15646) );
  IV U18386 ( .A(n15618), .Z(n15643) );
  XOR U18387 ( .A(n15616), .B(n15649), .Z(n15618) );
  XOR U18388 ( .A(n15650), .B(n15651), .Z(n15649) );
  ANDN U18389 ( .B(n15652), .A(n15653), .Z(n15650) );
  XOR U18390 ( .A(n15654), .B(n15651), .Z(n15652) );
  IV U18391 ( .A(n15619), .Z(n15616) );
  XOR U18392 ( .A(n15655), .B(n15656), .Z(n15619) );
  ANDN U18393 ( .B(n15657), .A(n15658), .Z(n15655) );
  XOR U18394 ( .A(n15656), .B(n15659), .Z(n15657) );
  XOR U18395 ( .A(n15660), .B(n15661), .Z(n15632) );
  XNOR U18396 ( .A(n15627), .B(n15662), .Z(n15661) );
  IV U18397 ( .A(n15630), .Z(n15662) );
  XOR U18398 ( .A(n15663), .B(n15664), .Z(n15630) );
  ANDN U18399 ( .B(n15665), .A(n15666), .Z(n15663) );
  XOR U18400 ( .A(n15664), .B(n15667), .Z(n15665) );
  XNOR U18401 ( .A(n15668), .B(n15669), .Z(n15627) );
  ANDN U18402 ( .B(n15670), .A(n15671), .Z(n15668) );
  XOR U18403 ( .A(n15669), .B(n15672), .Z(n15670) );
  IV U18404 ( .A(n15626), .Z(n15660) );
  XOR U18405 ( .A(n15624), .B(n15673), .Z(n15626) );
  XOR U18406 ( .A(n15674), .B(n15675), .Z(n15673) );
  ANDN U18407 ( .B(n15676), .A(n15677), .Z(n15674) );
  XOR U18408 ( .A(n15678), .B(n15675), .Z(n15676) );
  IV U18409 ( .A(n15628), .Z(n15624) );
  XOR U18410 ( .A(n15679), .B(n15680), .Z(n15628) );
  ANDN U18411 ( .B(n15681), .A(n15682), .Z(n15679) );
  XOR U18412 ( .A(n15683), .B(n15680), .Z(n15681) );
  IV U18413 ( .A(n15638), .Z(n15642) );
  XOR U18414 ( .A(n15638), .B(n15593), .Z(n15640) );
  XOR U18415 ( .A(n15684), .B(n15685), .Z(n15593) );
  AND U18416 ( .A(n170), .B(n15686), .Z(n15684) );
  XOR U18417 ( .A(n15687), .B(n15685), .Z(n15686) );
  NANDN U18418 ( .A(n15595), .B(n15597), .Z(n15638) );
  XOR U18419 ( .A(n15688), .B(n15689), .Z(n15597) );
  AND U18420 ( .A(n170), .B(n15690), .Z(n15688) );
  XOR U18421 ( .A(n15689), .B(n15691), .Z(n15690) );
  XNOR U18422 ( .A(n15692), .B(n15693), .Z(n170) );
  AND U18423 ( .A(n15694), .B(n15695), .Z(n15692) );
  XOR U18424 ( .A(n15693), .B(n15608), .Z(n15695) );
  XNOR U18425 ( .A(n15696), .B(n15697), .Z(n15608) );
  ANDN U18426 ( .B(n15698), .A(n15699), .Z(n15696) );
  XOR U18427 ( .A(n15697), .B(n15700), .Z(n15698) );
  XNOR U18428 ( .A(n15693), .B(n15610), .Z(n15694) );
  XOR U18429 ( .A(n15701), .B(n15702), .Z(n15610) );
  AND U18430 ( .A(n174), .B(n15703), .Z(n15701) );
  XOR U18431 ( .A(n15704), .B(n15702), .Z(n15703) );
  XNOR U18432 ( .A(n15705), .B(n15706), .Z(n15693) );
  AND U18433 ( .A(n15707), .B(n15708), .Z(n15705) );
  XNOR U18434 ( .A(n15706), .B(n15635), .Z(n15708) );
  XOR U18435 ( .A(n15699), .B(n15700), .Z(n15635) );
  XNOR U18436 ( .A(n15709), .B(n15710), .Z(n15700) );
  ANDN U18437 ( .B(n15711), .A(n15712), .Z(n15709) );
  XOR U18438 ( .A(n15713), .B(n15714), .Z(n15711) );
  XOR U18439 ( .A(n15715), .B(n15716), .Z(n15699) );
  XNOR U18440 ( .A(n15717), .B(n15718), .Z(n15716) );
  ANDN U18441 ( .B(n15719), .A(n15720), .Z(n15717) );
  XNOR U18442 ( .A(n15721), .B(n15722), .Z(n15719) );
  IV U18443 ( .A(n15697), .Z(n15715) );
  XOR U18444 ( .A(n15723), .B(n15724), .Z(n15697) );
  ANDN U18445 ( .B(n15725), .A(n15726), .Z(n15723) );
  XOR U18446 ( .A(n15724), .B(n15727), .Z(n15725) );
  XOR U18447 ( .A(n15706), .B(n15637), .Z(n15707) );
  XOR U18448 ( .A(n15728), .B(n15729), .Z(n15637) );
  AND U18449 ( .A(n174), .B(n15730), .Z(n15728) );
  XOR U18450 ( .A(n15731), .B(n15729), .Z(n15730) );
  XNOR U18451 ( .A(n15732), .B(n15733), .Z(n15706) );
  NAND U18452 ( .A(n15734), .B(n15735), .Z(n15733) );
  XOR U18453 ( .A(n15736), .B(n15685), .Z(n15735) );
  XOR U18454 ( .A(n15726), .B(n15727), .Z(n15685) );
  XOR U18455 ( .A(n15737), .B(n15714), .Z(n15727) );
  XOR U18456 ( .A(n15738), .B(n15739), .Z(n15714) );
  ANDN U18457 ( .B(n15740), .A(n15741), .Z(n15738) );
  XOR U18458 ( .A(n15739), .B(n15742), .Z(n15740) );
  IV U18459 ( .A(n15712), .Z(n15737) );
  XOR U18460 ( .A(n15710), .B(n15743), .Z(n15712) );
  XOR U18461 ( .A(n15744), .B(n15745), .Z(n15743) );
  ANDN U18462 ( .B(n15746), .A(n15747), .Z(n15744) );
  XOR U18463 ( .A(n15748), .B(n15745), .Z(n15746) );
  IV U18464 ( .A(n15713), .Z(n15710) );
  XOR U18465 ( .A(n15749), .B(n15750), .Z(n15713) );
  ANDN U18466 ( .B(n15751), .A(n15752), .Z(n15749) );
  XOR U18467 ( .A(n15750), .B(n15753), .Z(n15751) );
  XOR U18468 ( .A(n15754), .B(n15755), .Z(n15726) );
  XNOR U18469 ( .A(n15721), .B(n15756), .Z(n15755) );
  IV U18470 ( .A(n15724), .Z(n15756) );
  XOR U18471 ( .A(n15757), .B(n15758), .Z(n15724) );
  ANDN U18472 ( .B(n15759), .A(n15760), .Z(n15757) );
  XOR U18473 ( .A(n15758), .B(n15761), .Z(n15759) );
  XNOR U18474 ( .A(n15762), .B(n15763), .Z(n15721) );
  ANDN U18475 ( .B(n15764), .A(n15765), .Z(n15762) );
  XOR U18476 ( .A(n15763), .B(n15766), .Z(n15764) );
  IV U18477 ( .A(n15720), .Z(n15754) );
  XOR U18478 ( .A(n15718), .B(n15767), .Z(n15720) );
  XOR U18479 ( .A(n15768), .B(n15769), .Z(n15767) );
  ANDN U18480 ( .B(n15770), .A(n15771), .Z(n15768) );
  XOR U18481 ( .A(n15772), .B(n15769), .Z(n15770) );
  IV U18482 ( .A(n15722), .Z(n15718) );
  XOR U18483 ( .A(n15773), .B(n15774), .Z(n15722) );
  ANDN U18484 ( .B(n15775), .A(n15776), .Z(n15773) );
  XOR U18485 ( .A(n15777), .B(n15774), .Z(n15775) );
  IV U18486 ( .A(n15732), .Z(n15736) );
  XOR U18487 ( .A(n15732), .B(n15687), .Z(n15734) );
  XOR U18488 ( .A(n15778), .B(n15779), .Z(n15687) );
  AND U18489 ( .A(n174), .B(n15780), .Z(n15778) );
  XOR U18490 ( .A(n15781), .B(n15779), .Z(n15780) );
  NANDN U18491 ( .A(n15689), .B(n15691), .Z(n15732) );
  XOR U18492 ( .A(n15782), .B(n15783), .Z(n15691) );
  AND U18493 ( .A(n174), .B(n15784), .Z(n15782) );
  XOR U18494 ( .A(n15783), .B(n15785), .Z(n15784) );
  XNOR U18495 ( .A(n15786), .B(n15787), .Z(n174) );
  AND U18496 ( .A(n15788), .B(n15789), .Z(n15786) );
  XOR U18497 ( .A(n15787), .B(n15702), .Z(n15789) );
  XNOR U18498 ( .A(n15790), .B(n15791), .Z(n15702) );
  ANDN U18499 ( .B(n15792), .A(n15793), .Z(n15790) );
  XOR U18500 ( .A(n15791), .B(n15794), .Z(n15792) );
  XNOR U18501 ( .A(n15787), .B(n15704), .Z(n15788) );
  XOR U18502 ( .A(n15795), .B(n15796), .Z(n15704) );
  AND U18503 ( .A(n178), .B(n15797), .Z(n15795) );
  XOR U18504 ( .A(n15798), .B(n15796), .Z(n15797) );
  XNOR U18505 ( .A(n15799), .B(n15800), .Z(n15787) );
  AND U18506 ( .A(n15801), .B(n15802), .Z(n15799) );
  XNOR U18507 ( .A(n15800), .B(n15729), .Z(n15802) );
  XOR U18508 ( .A(n15793), .B(n15794), .Z(n15729) );
  XNOR U18509 ( .A(n15803), .B(n15804), .Z(n15794) );
  ANDN U18510 ( .B(n15805), .A(n15806), .Z(n15803) );
  XOR U18511 ( .A(n15807), .B(n15808), .Z(n15805) );
  XOR U18512 ( .A(n15809), .B(n15810), .Z(n15793) );
  XNOR U18513 ( .A(n15811), .B(n15812), .Z(n15810) );
  ANDN U18514 ( .B(n15813), .A(n15814), .Z(n15811) );
  XNOR U18515 ( .A(n15815), .B(n15816), .Z(n15813) );
  IV U18516 ( .A(n15791), .Z(n15809) );
  XOR U18517 ( .A(n15817), .B(n15818), .Z(n15791) );
  ANDN U18518 ( .B(n15819), .A(n15820), .Z(n15817) );
  XOR U18519 ( .A(n15818), .B(n15821), .Z(n15819) );
  XOR U18520 ( .A(n15800), .B(n15731), .Z(n15801) );
  XOR U18521 ( .A(n15822), .B(n15823), .Z(n15731) );
  AND U18522 ( .A(n178), .B(n15824), .Z(n15822) );
  XOR U18523 ( .A(n15825), .B(n15823), .Z(n15824) );
  XNOR U18524 ( .A(n15826), .B(n15827), .Z(n15800) );
  NAND U18525 ( .A(n15828), .B(n15829), .Z(n15827) );
  XOR U18526 ( .A(n15830), .B(n15779), .Z(n15829) );
  XOR U18527 ( .A(n15820), .B(n15821), .Z(n15779) );
  XOR U18528 ( .A(n15831), .B(n15808), .Z(n15821) );
  XOR U18529 ( .A(n15832), .B(n15833), .Z(n15808) );
  ANDN U18530 ( .B(n15834), .A(n15835), .Z(n15832) );
  XOR U18531 ( .A(n15833), .B(n15836), .Z(n15834) );
  IV U18532 ( .A(n15806), .Z(n15831) );
  XOR U18533 ( .A(n15804), .B(n15837), .Z(n15806) );
  XOR U18534 ( .A(n15838), .B(n15839), .Z(n15837) );
  ANDN U18535 ( .B(n15840), .A(n15841), .Z(n15838) );
  XOR U18536 ( .A(n15842), .B(n15839), .Z(n15840) );
  IV U18537 ( .A(n15807), .Z(n15804) );
  XOR U18538 ( .A(n15843), .B(n15844), .Z(n15807) );
  ANDN U18539 ( .B(n15845), .A(n15846), .Z(n15843) );
  XOR U18540 ( .A(n15844), .B(n15847), .Z(n15845) );
  XOR U18541 ( .A(n15848), .B(n15849), .Z(n15820) );
  XNOR U18542 ( .A(n15815), .B(n15850), .Z(n15849) );
  IV U18543 ( .A(n15818), .Z(n15850) );
  XOR U18544 ( .A(n15851), .B(n15852), .Z(n15818) );
  ANDN U18545 ( .B(n15853), .A(n15854), .Z(n15851) );
  XOR U18546 ( .A(n15852), .B(n15855), .Z(n15853) );
  XNOR U18547 ( .A(n15856), .B(n15857), .Z(n15815) );
  ANDN U18548 ( .B(n15858), .A(n15859), .Z(n15856) );
  XOR U18549 ( .A(n15857), .B(n15860), .Z(n15858) );
  IV U18550 ( .A(n15814), .Z(n15848) );
  XOR U18551 ( .A(n15812), .B(n15861), .Z(n15814) );
  XOR U18552 ( .A(n15862), .B(n15863), .Z(n15861) );
  ANDN U18553 ( .B(n15864), .A(n15865), .Z(n15862) );
  XOR U18554 ( .A(n15866), .B(n15863), .Z(n15864) );
  IV U18555 ( .A(n15816), .Z(n15812) );
  XOR U18556 ( .A(n15867), .B(n15868), .Z(n15816) );
  ANDN U18557 ( .B(n15869), .A(n15870), .Z(n15867) );
  XOR U18558 ( .A(n15871), .B(n15868), .Z(n15869) );
  IV U18559 ( .A(n15826), .Z(n15830) );
  XOR U18560 ( .A(n15826), .B(n15781), .Z(n15828) );
  XOR U18561 ( .A(n15872), .B(n15873), .Z(n15781) );
  AND U18562 ( .A(n178), .B(n15874), .Z(n15872) );
  XOR U18563 ( .A(n15875), .B(n15873), .Z(n15874) );
  NANDN U18564 ( .A(n15783), .B(n15785), .Z(n15826) );
  XOR U18565 ( .A(n15876), .B(n15877), .Z(n15785) );
  AND U18566 ( .A(n178), .B(n15878), .Z(n15876) );
  XOR U18567 ( .A(n15877), .B(n15879), .Z(n15878) );
  XNOR U18568 ( .A(n15880), .B(n15881), .Z(n178) );
  AND U18569 ( .A(n15882), .B(n15883), .Z(n15880) );
  XOR U18570 ( .A(n15881), .B(n15796), .Z(n15883) );
  XNOR U18571 ( .A(n15884), .B(n15885), .Z(n15796) );
  ANDN U18572 ( .B(n15886), .A(n15887), .Z(n15884) );
  XOR U18573 ( .A(n15885), .B(n15888), .Z(n15886) );
  XNOR U18574 ( .A(n15881), .B(n15798), .Z(n15882) );
  XOR U18575 ( .A(n15889), .B(n15890), .Z(n15798) );
  AND U18576 ( .A(n182), .B(n15891), .Z(n15889) );
  XOR U18577 ( .A(n15892), .B(n15890), .Z(n15891) );
  XNOR U18578 ( .A(n15893), .B(n15894), .Z(n15881) );
  AND U18579 ( .A(n15895), .B(n15896), .Z(n15893) );
  XNOR U18580 ( .A(n15894), .B(n15823), .Z(n15896) );
  XOR U18581 ( .A(n15887), .B(n15888), .Z(n15823) );
  XNOR U18582 ( .A(n15897), .B(n15898), .Z(n15888) );
  ANDN U18583 ( .B(n15899), .A(n15900), .Z(n15897) );
  XOR U18584 ( .A(n15901), .B(n15902), .Z(n15899) );
  XOR U18585 ( .A(n15903), .B(n15904), .Z(n15887) );
  XNOR U18586 ( .A(n15905), .B(n15906), .Z(n15904) );
  ANDN U18587 ( .B(n15907), .A(n15908), .Z(n15905) );
  XNOR U18588 ( .A(n15909), .B(n15910), .Z(n15907) );
  IV U18589 ( .A(n15885), .Z(n15903) );
  XOR U18590 ( .A(n15911), .B(n15912), .Z(n15885) );
  ANDN U18591 ( .B(n15913), .A(n15914), .Z(n15911) );
  XOR U18592 ( .A(n15912), .B(n15915), .Z(n15913) );
  XOR U18593 ( .A(n15894), .B(n15825), .Z(n15895) );
  XOR U18594 ( .A(n15916), .B(n15917), .Z(n15825) );
  AND U18595 ( .A(n182), .B(n15918), .Z(n15916) );
  XOR U18596 ( .A(n15919), .B(n15917), .Z(n15918) );
  XNOR U18597 ( .A(n15920), .B(n15921), .Z(n15894) );
  NAND U18598 ( .A(n15922), .B(n15923), .Z(n15921) );
  XOR U18599 ( .A(n15924), .B(n15873), .Z(n15923) );
  XOR U18600 ( .A(n15914), .B(n15915), .Z(n15873) );
  XOR U18601 ( .A(n15925), .B(n15902), .Z(n15915) );
  XOR U18602 ( .A(n15926), .B(n15927), .Z(n15902) );
  ANDN U18603 ( .B(n15928), .A(n15929), .Z(n15926) );
  XOR U18604 ( .A(n15927), .B(n15930), .Z(n15928) );
  IV U18605 ( .A(n15900), .Z(n15925) );
  XOR U18606 ( .A(n15898), .B(n15931), .Z(n15900) );
  XOR U18607 ( .A(n15932), .B(n15933), .Z(n15931) );
  ANDN U18608 ( .B(n15934), .A(n15935), .Z(n15932) );
  XOR U18609 ( .A(n15936), .B(n15933), .Z(n15934) );
  IV U18610 ( .A(n15901), .Z(n15898) );
  XOR U18611 ( .A(n15937), .B(n15938), .Z(n15901) );
  ANDN U18612 ( .B(n15939), .A(n15940), .Z(n15937) );
  XOR U18613 ( .A(n15938), .B(n15941), .Z(n15939) );
  XOR U18614 ( .A(n15942), .B(n15943), .Z(n15914) );
  XNOR U18615 ( .A(n15909), .B(n15944), .Z(n15943) );
  IV U18616 ( .A(n15912), .Z(n15944) );
  XOR U18617 ( .A(n15945), .B(n15946), .Z(n15912) );
  ANDN U18618 ( .B(n15947), .A(n15948), .Z(n15945) );
  XOR U18619 ( .A(n15946), .B(n15949), .Z(n15947) );
  XNOR U18620 ( .A(n15950), .B(n15951), .Z(n15909) );
  ANDN U18621 ( .B(n15952), .A(n15953), .Z(n15950) );
  XOR U18622 ( .A(n15951), .B(n15954), .Z(n15952) );
  IV U18623 ( .A(n15908), .Z(n15942) );
  XOR U18624 ( .A(n15906), .B(n15955), .Z(n15908) );
  XOR U18625 ( .A(n15956), .B(n15957), .Z(n15955) );
  ANDN U18626 ( .B(n15958), .A(n15959), .Z(n15956) );
  XOR U18627 ( .A(n15960), .B(n15957), .Z(n15958) );
  IV U18628 ( .A(n15910), .Z(n15906) );
  XOR U18629 ( .A(n15961), .B(n15962), .Z(n15910) );
  ANDN U18630 ( .B(n15963), .A(n15964), .Z(n15961) );
  XOR U18631 ( .A(n15965), .B(n15962), .Z(n15963) );
  IV U18632 ( .A(n15920), .Z(n15924) );
  XOR U18633 ( .A(n15920), .B(n15875), .Z(n15922) );
  XOR U18634 ( .A(n15966), .B(n15967), .Z(n15875) );
  AND U18635 ( .A(n182), .B(n15968), .Z(n15966) );
  XOR U18636 ( .A(n15969), .B(n15967), .Z(n15968) );
  NANDN U18637 ( .A(n15877), .B(n15879), .Z(n15920) );
  XOR U18638 ( .A(n15970), .B(n15971), .Z(n15879) );
  AND U18639 ( .A(n182), .B(n15972), .Z(n15970) );
  XOR U18640 ( .A(n15971), .B(n15973), .Z(n15972) );
  XNOR U18641 ( .A(n15974), .B(n15975), .Z(n182) );
  AND U18642 ( .A(n15976), .B(n15977), .Z(n15974) );
  XOR U18643 ( .A(n15975), .B(n15890), .Z(n15977) );
  XNOR U18644 ( .A(n15978), .B(n15979), .Z(n15890) );
  ANDN U18645 ( .B(n15980), .A(n15981), .Z(n15978) );
  XOR U18646 ( .A(n15979), .B(n15982), .Z(n15980) );
  XNOR U18647 ( .A(n15975), .B(n15892), .Z(n15976) );
  XOR U18648 ( .A(n15983), .B(n15984), .Z(n15892) );
  AND U18649 ( .A(n186), .B(n15985), .Z(n15983) );
  XOR U18650 ( .A(n15986), .B(n15984), .Z(n15985) );
  XNOR U18651 ( .A(n15987), .B(n15988), .Z(n15975) );
  AND U18652 ( .A(n15989), .B(n15990), .Z(n15987) );
  XNOR U18653 ( .A(n15988), .B(n15917), .Z(n15990) );
  XOR U18654 ( .A(n15981), .B(n15982), .Z(n15917) );
  XNOR U18655 ( .A(n15991), .B(n15992), .Z(n15982) );
  ANDN U18656 ( .B(n15993), .A(n15994), .Z(n15991) );
  XOR U18657 ( .A(n15995), .B(n15996), .Z(n15993) );
  XOR U18658 ( .A(n15997), .B(n15998), .Z(n15981) );
  XNOR U18659 ( .A(n15999), .B(n16000), .Z(n15998) );
  ANDN U18660 ( .B(n16001), .A(n16002), .Z(n15999) );
  XNOR U18661 ( .A(n16003), .B(n16004), .Z(n16001) );
  IV U18662 ( .A(n15979), .Z(n15997) );
  XOR U18663 ( .A(n16005), .B(n16006), .Z(n15979) );
  ANDN U18664 ( .B(n16007), .A(n16008), .Z(n16005) );
  XOR U18665 ( .A(n16006), .B(n16009), .Z(n16007) );
  XOR U18666 ( .A(n15988), .B(n15919), .Z(n15989) );
  XOR U18667 ( .A(n16010), .B(n16011), .Z(n15919) );
  AND U18668 ( .A(n186), .B(n16012), .Z(n16010) );
  XOR U18669 ( .A(n16013), .B(n16011), .Z(n16012) );
  XNOR U18670 ( .A(n16014), .B(n16015), .Z(n15988) );
  NAND U18671 ( .A(n16016), .B(n16017), .Z(n16015) );
  XOR U18672 ( .A(n16018), .B(n15967), .Z(n16017) );
  XOR U18673 ( .A(n16008), .B(n16009), .Z(n15967) );
  XOR U18674 ( .A(n16019), .B(n15996), .Z(n16009) );
  XOR U18675 ( .A(n16020), .B(n16021), .Z(n15996) );
  ANDN U18676 ( .B(n16022), .A(n16023), .Z(n16020) );
  XOR U18677 ( .A(n16021), .B(n16024), .Z(n16022) );
  IV U18678 ( .A(n15994), .Z(n16019) );
  XOR U18679 ( .A(n15992), .B(n16025), .Z(n15994) );
  XOR U18680 ( .A(n16026), .B(n16027), .Z(n16025) );
  ANDN U18681 ( .B(n16028), .A(n16029), .Z(n16026) );
  XOR U18682 ( .A(n16030), .B(n16027), .Z(n16028) );
  IV U18683 ( .A(n15995), .Z(n15992) );
  XOR U18684 ( .A(n16031), .B(n16032), .Z(n15995) );
  ANDN U18685 ( .B(n16033), .A(n16034), .Z(n16031) );
  XOR U18686 ( .A(n16032), .B(n16035), .Z(n16033) );
  XOR U18687 ( .A(n16036), .B(n16037), .Z(n16008) );
  XNOR U18688 ( .A(n16003), .B(n16038), .Z(n16037) );
  IV U18689 ( .A(n16006), .Z(n16038) );
  XOR U18690 ( .A(n16039), .B(n16040), .Z(n16006) );
  ANDN U18691 ( .B(n16041), .A(n16042), .Z(n16039) );
  XOR U18692 ( .A(n16040), .B(n16043), .Z(n16041) );
  XNOR U18693 ( .A(n16044), .B(n16045), .Z(n16003) );
  ANDN U18694 ( .B(n16046), .A(n16047), .Z(n16044) );
  XOR U18695 ( .A(n16045), .B(n16048), .Z(n16046) );
  IV U18696 ( .A(n16002), .Z(n16036) );
  XOR U18697 ( .A(n16000), .B(n16049), .Z(n16002) );
  XOR U18698 ( .A(n16050), .B(n16051), .Z(n16049) );
  ANDN U18699 ( .B(n16052), .A(n16053), .Z(n16050) );
  XOR U18700 ( .A(n16054), .B(n16051), .Z(n16052) );
  IV U18701 ( .A(n16004), .Z(n16000) );
  XOR U18702 ( .A(n16055), .B(n16056), .Z(n16004) );
  ANDN U18703 ( .B(n16057), .A(n16058), .Z(n16055) );
  XOR U18704 ( .A(n16059), .B(n16056), .Z(n16057) );
  IV U18705 ( .A(n16014), .Z(n16018) );
  XOR U18706 ( .A(n16014), .B(n15969), .Z(n16016) );
  XOR U18707 ( .A(n16060), .B(n16061), .Z(n15969) );
  AND U18708 ( .A(n186), .B(n16062), .Z(n16060) );
  XOR U18709 ( .A(n16063), .B(n16061), .Z(n16062) );
  NANDN U18710 ( .A(n15971), .B(n15973), .Z(n16014) );
  XOR U18711 ( .A(n16064), .B(n16065), .Z(n15973) );
  AND U18712 ( .A(n186), .B(n16066), .Z(n16064) );
  XOR U18713 ( .A(n16065), .B(n16067), .Z(n16066) );
  XNOR U18714 ( .A(n16068), .B(n16069), .Z(n186) );
  AND U18715 ( .A(n16070), .B(n16071), .Z(n16068) );
  XOR U18716 ( .A(n16069), .B(n15984), .Z(n16071) );
  XNOR U18717 ( .A(n16072), .B(n16073), .Z(n15984) );
  ANDN U18718 ( .B(n16074), .A(n16075), .Z(n16072) );
  XOR U18719 ( .A(n16073), .B(n16076), .Z(n16074) );
  XNOR U18720 ( .A(n16069), .B(n15986), .Z(n16070) );
  XOR U18721 ( .A(n16077), .B(n16078), .Z(n15986) );
  AND U18722 ( .A(n190), .B(n16079), .Z(n16077) );
  XOR U18723 ( .A(n16080), .B(n16078), .Z(n16079) );
  XNOR U18724 ( .A(n16081), .B(n16082), .Z(n16069) );
  AND U18725 ( .A(n16083), .B(n16084), .Z(n16081) );
  XNOR U18726 ( .A(n16082), .B(n16011), .Z(n16084) );
  XOR U18727 ( .A(n16075), .B(n16076), .Z(n16011) );
  XNOR U18728 ( .A(n16085), .B(n16086), .Z(n16076) );
  ANDN U18729 ( .B(n16087), .A(n16088), .Z(n16085) );
  XOR U18730 ( .A(n16089), .B(n16090), .Z(n16087) );
  XOR U18731 ( .A(n16091), .B(n16092), .Z(n16075) );
  XNOR U18732 ( .A(n16093), .B(n16094), .Z(n16092) );
  ANDN U18733 ( .B(n16095), .A(n16096), .Z(n16093) );
  XNOR U18734 ( .A(n16097), .B(n16098), .Z(n16095) );
  IV U18735 ( .A(n16073), .Z(n16091) );
  XOR U18736 ( .A(n16099), .B(n16100), .Z(n16073) );
  ANDN U18737 ( .B(n16101), .A(n16102), .Z(n16099) );
  XOR U18738 ( .A(n16100), .B(n16103), .Z(n16101) );
  XOR U18739 ( .A(n16082), .B(n16013), .Z(n16083) );
  XOR U18740 ( .A(n16104), .B(n16105), .Z(n16013) );
  AND U18741 ( .A(n190), .B(n16106), .Z(n16104) );
  XOR U18742 ( .A(n16107), .B(n16105), .Z(n16106) );
  XNOR U18743 ( .A(n16108), .B(n16109), .Z(n16082) );
  NAND U18744 ( .A(n16110), .B(n16111), .Z(n16109) );
  XOR U18745 ( .A(n16112), .B(n16061), .Z(n16111) );
  XOR U18746 ( .A(n16102), .B(n16103), .Z(n16061) );
  XOR U18747 ( .A(n16113), .B(n16090), .Z(n16103) );
  XOR U18748 ( .A(n16114), .B(n16115), .Z(n16090) );
  ANDN U18749 ( .B(n16116), .A(n16117), .Z(n16114) );
  XOR U18750 ( .A(n16115), .B(n16118), .Z(n16116) );
  IV U18751 ( .A(n16088), .Z(n16113) );
  XOR U18752 ( .A(n16086), .B(n16119), .Z(n16088) );
  XOR U18753 ( .A(n16120), .B(n16121), .Z(n16119) );
  ANDN U18754 ( .B(n16122), .A(n16123), .Z(n16120) );
  XOR U18755 ( .A(n16124), .B(n16121), .Z(n16122) );
  IV U18756 ( .A(n16089), .Z(n16086) );
  XOR U18757 ( .A(n16125), .B(n16126), .Z(n16089) );
  ANDN U18758 ( .B(n16127), .A(n16128), .Z(n16125) );
  XOR U18759 ( .A(n16126), .B(n16129), .Z(n16127) );
  XOR U18760 ( .A(n16130), .B(n16131), .Z(n16102) );
  XNOR U18761 ( .A(n16097), .B(n16132), .Z(n16131) );
  IV U18762 ( .A(n16100), .Z(n16132) );
  XOR U18763 ( .A(n16133), .B(n16134), .Z(n16100) );
  ANDN U18764 ( .B(n16135), .A(n16136), .Z(n16133) );
  XOR U18765 ( .A(n16134), .B(n16137), .Z(n16135) );
  XNOR U18766 ( .A(n16138), .B(n16139), .Z(n16097) );
  ANDN U18767 ( .B(n16140), .A(n16141), .Z(n16138) );
  XOR U18768 ( .A(n16139), .B(n16142), .Z(n16140) );
  IV U18769 ( .A(n16096), .Z(n16130) );
  XOR U18770 ( .A(n16094), .B(n16143), .Z(n16096) );
  XOR U18771 ( .A(n16144), .B(n16145), .Z(n16143) );
  ANDN U18772 ( .B(n16146), .A(n16147), .Z(n16144) );
  XOR U18773 ( .A(n16148), .B(n16145), .Z(n16146) );
  IV U18774 ( .A(n16098), .Z(n16094) );
  XOR U18775 ( .A(n16149), .B(n16150), .Z(n16098) );
  ANDN U18776 ( .B(n16151), .A(n16152), .Z(n16149) );
  XOR U18777 ( .A(n16153), .B(n16150), .Z(n16151) );
  IV U18778 ( .A(n16108), .Z(n16112) );
  XOR U18779 ( .A(n16108), .B(n16063), .Z(n16110) );
  XOR U18780 ( .A(n16154), .B(n16155), .Z(n16063) );
  AND U18781 ( .A(n190), .B(n16156), .Z(n16154) );
  XOR U18782 ( .A(n16157), .B(n16155), .Z(n16156) );
  NANDN U18783 ( .A(n16065), .B(n16067), .Z(n16108) );
  XOR U18784 ( .A(n16158), .B(n16159), .Z(n16067) );
  AND U18785 ( .A(n190), .B(n16160), .Z(n16158) );
  XOR U18786 ( .A(n16159), .B(n16161), .Z(n16160) );
  XNOR U18787 ( .A(n16162), .B(n16163), .Z(n190) );
  AND U18788 ( .A(n16164), .B(n16165), .Z(n16162) );
  XOR U18789 ( .A(n16163), .B(n16078), .Z(n16165) );
  XNOR U18790 ( .A(n16166), .B(n16167), .Z(n16078) );
  ANDN U18791 ( .B(n16168), .A(n16169), .Z(n16166) );
  XOR U18792 ( .A(n16167), .B(n16170), .Z(n16168) );
  XNOR U18793 ( .A(n16163), .B(n16080), .Z(n16164) );
  XOR U18794 ( .A(n16171), .B(n16172), .Z(n16080) );
  AND U18795 ( .A(n194), .B(n16173), .Z(n16171) );
  XOR U18796 ( .A(n16174), .B(n16172), .Z(n16173) );
  XNOR U18797 ( .A(n16175), .B(n16176), .Z(n16163) );
  AND U18798 ( .A(n16177), .B(n16178), .Z(n16175) );
  XNOR U18799 ( .A(n16176), .B(n16105), .Z(n16178) );
  XOR U18800 ( .A(n16169), .B(n16170), .Z(n16105) );
  XNOR U18801 ( .A(n16179), .B(n16180), .Z(n16170) );
  ANDN U18802 ( .B(n16181), .A(n16182), .Z(n16179) );
  XOR U18803 ( .A(n16183), .B(n16184), .Z(n16181) );
  XOR U18804 ( .A(n16185), .B(n16186), .Z(n16169) );
  XNOR U18805 ( .A(n16187), .B(n16188), .Z(n16186) );
  ANDN U18806 ( .B(n16189), .A(n16190), .Z(n16187) );
  XNOR U18807 ( .A(n16191), .B(n16192), .Z(n16189) );
  IV U18808 ( .A(n16167), .Z(n16185) );
  XOR U18809 ( .A(n16193), .B(n16194), .Z(n16167) );
  ANDN U18810 ( .B(n16195), .A(n16196), .Z(n16193) );
  XOR U18811 ( .A(n16194), .B(n16197), .Z(n16195) );
  XOR U18812 ( .A(n16176), .B(n16107), .Z(n16177) );
  XOR U18813 ( .A(n16198), .B(n16199), .Z(n16107) );
  AND U18814 ( .A(n194), .B(n16200), .Z(n16198) );
  XOR U18815 ( .A(n16201), .B(n16199), .Z(n16200) );
  XNOR U18816 ( .A(n16202), .B(n16203), .Z(n16176) );
  NAND U18817 ( .A(n16204), .B(n16205), .Z(n16203) );
  XOR U18818 ( .A(n16206), .B(n16155), .Z(n16205) );
  XOR U18819 ( .A(n16196), .B(n16197), .Z(n16155) );
  XOR U18820 ( .A(n16207), .B(n16184), .Z(n16197) );
  XOR U18821 ( .A(n16208), .B(n16209), .Z(n16184) );
  ANDN U18822 ( .B(n16210), .A(n16211), .Z(n16208) );
  XOR U18823 ( .A(n16209), .B(n16212), .Z(n16210) );
  IV U18824 ( .A(n16182), .Z(n16207) );
  XOR U18825 ( .A(n16180), .B(n16213), .Z(n16182) );
  XOR U18826 ( .A(n16214), .B(n16215), .Z(n16213) );
  ANDN U18827 ( .B(n16216), .A(n16217), .Z(n16214) );
  XOR U18828 ( .A(n16218), .B(n16215), .Z(n16216) );
  IV U18829 ( .A(n16183), .Z(n16180) );
  XOR U18830 ( .A(n16219), .B(n16220), .Z(n16183) );
  ANDN U18831 ( .B(n16221), .A(n16222), .Z(n16219) );
  XOR U18832 ( .A(n16220), .B(n16223), .Z(n16221) );
  XOR U18833 ( .A(n16224), .B(n16225), .Z(n16196) );
  XNOR U18834 ( .A(n16191), .B(n16226), .Z(n16225) );
  IV U18835 ( .A(n16194), .Z(n16226) );
  XOR U18836 ( .A(n16227), .B(n16228), .Z(n16194) );
  ANDN U18837 ( .B(n16229), .A(n16230), .Z(n16227) );
  XOR U18838 ( .A(n16228), .B(n16231), .Z(n16229) );
  XNOR U18839 ( .A(n16232), .B(n16233), .Z(n16191) );
  ANDN U18840 ( .B(n16234), .A(n16235), .Z(n16232) );
  XOR U18841 ( .A(n16233), .B(n16236), .Z(n16234) );
  IV U18842 ( .A(n16190), .Z(n16224) );
  XOR U18843 ( .A(n16188), .B(n16237), .Z(n16190) );
  XOR U18844 ( .A(n16238), .B(n16239), .Z(n16237) );
  ANDN U18845 ( .B(n16240), .A(n16241), .Z(n16238) );
  XOR U18846 ( .A(n16242), .B(n16239), .Z(n16240) );
  IV U18847 ( .A(n16192), .Z(n16188) );
  XOR U18848 ( .A(n16243), .B(n16244), .Z(n16192) );
  ANDN U18849 ( .B(n16245), .A(n16246), .Z(n16243) );
  XOR U18850 ( .A(n16247), .B(n16244), .Z(n16245) );
  IV U18851 ( .A(n16202), .Z(n16206) );
  XOR U18852 ( .A(n16202), .B(n16157), .Z(n16204) );
  XOR U18853 ( .A(n16248), .B(n16249), .Z(n16157) );
  AND U18854 ( .A(n194), .B(n16250), .Z(n16248) );
  XOR U18855 ( .A(n16251), .B(n16249), .Z(n16250) );
  NANDN U18856 ( .A(n16159), .B(n16161), .Z(n16202) );
  XOR U18857 ( .A(n16252), .B(n16253), .Z(n16161) );
  AND U18858 ( .A(n194), .B(n16254), .Z(n16252) );
  XOR U18859 ( .A(n16253), .B(n16255), .Z(n16254) );
  XNOR U18860 ( .A(n16256), .B(n16257), .Z(n194) );
  AND U18861 ( .A(n16258), .B(n16259), .Z(n16256) );
  XOR U18862 ( .A(n16257), .B(n16172), .Z(n16259) );
  XNOR U18863 ( .A(n16260), .B(n16261), .Z(n16172) );
  ANDN U18864 ( .B(n16262), .A(n16263), .Z(n16260) );
  XOR U18865 ( .A(n16261), .B(n16264), .Z(n16262) );
  XNOR U18866 ( .A(n16257), .B(n16174), .Z(n16258) );
  XOR U18867 ( .A(n16265), .B(n16266), .Z(n16174) );
  AND U18868 ( .A(n198), .B(n16267), .Z(n16265) );
  XOR U18869 ( .A(n16268), .B(n16266), .Z(n16267) );
  XNOR U18870 ( .A(n16269), .B(n16270), .Z(n16257) );
  AND U18871 ( .A(n16271), .B(n16272), .Z(n16269) );
  XNOR U18872 ( .A(n16270), .B(n16199), .Z(n16272) );
  XOR U18873 ( .A(n16263), .B(n16264), .Z(n16199) );
  XNOR U18874 ( .A(n16273), .B(n16274), .Z(n16264) );
  ANDN U18875 ( .B(n16275), .A(n16276), .Z(n16273) );
  XOR U18876 ( .A(n16277), .B(n16278), .Z(n16275) );
  XOR U18877 ( .A(n16279), .B(n16280), .Z(n16263) );
  XNOR U18878 ( .A(n16281), .B(n16282), .Z(n16280) );
  ANDN U18879 ( .B(n16283), .A(n16284), .Z(n16281) );
  XNOR U18880 ( .A(n16285), .B(n16286), .Z(n16283) );
  IV U18881 ( .A(n16261), .Z(n16279) );
  XOR U18882 ( .A(n16287), .B(n16288), .Z(n16261) );
  ANDN U18883 ( .B(n16289), .A(n16290), .Z(n16287) );
  XOR U18884 ( .A(n16288), .B(n16291), .Z(n16289) );
  XOR U18885 ( .A(n16270), .B(n16201), .Z(n16271) );
  XOR U18886 ( .A(n16292), .B(n16293), .Z(n16201) );
  AND U18887 ( .A(n198), .B(n16294), .Z(n16292) );
  XOR U18888 ( .A(n16295), .B(n16293), .Z(n16294) );
  XNOR U18889 ( .A(n16296), .B(n16297), .Z(n16270) );
  NAND U18890 ( .A(n16298), .B(n16299), .Z(n16297) );
  XOR U18891 ( .A(n16300), .B(n16249), .Z(n16299) );
  XOR U18892 ( .A(n16290), .B(n16291), .Z(n16249) );
  XOR U18893 ( .A(n16301), .B(n16278), .Z(n16291) );
  XOR U18894 ( .A(n16302), .B(n16303), .Z(n16278) );
  ANDN U18895 ( .B(n16304), .A(n16305), .Z(n16302) );
  XOR U18896 ( .A(n16303), .B(n16306), .Z(n16304) );
  IV U18897 ( .A(n16276), .Z(n16301) );
  XOR U18898 ( .A(n16274), .B(n16307), .Z(n16276) );
  XOR U18899 ( .A(n16308), .B(n16309), .Z(n16307) );
  ANDN U18900 ( .B(n16310), .A(n16311), .Z(n16308) );
  XOR U18901 ( .A(n16312), .B(n16309), .Z(n16310) );
  IV U18902 ( .A(n16277), .Z(n16274) );
  XOR U18903 ( .A(n16313), .B(n16314), .Z(n16277) );
  ANDN U18904 ( .B(n16315), .A(n16316), .Z(n16313) );
  XOR U18905 ( .A(n16314), .B(n16317), .Z(n16315) );
  XOR U18906 ( .A(n16318), .B(n16319), .Z(n16290) );
  XNOR U18907 ( .A(n16285), .B(n16320), .Z(n16319) );
  IV U18908 ( .A(n16288), .Z(n16320) );
  XOR U18909 ( .A(n16321), .B(n16322), .Z(n16288) );
  ANDN U18910 ( .B(n16323), .A(n16324), .Z(n16321) );
  XOR U18911 ( .A(n16322), .B(n16325), .Z(n16323) );
  XNOR U18912 ( .A(n16326), .B(n16327), .Z(n16285) );
  ANDN U18913 ( .B(n16328), .A(n16329), .Z(n16326) );
  XOR U18914 ( .A(n16327), .B(n16330), .Z(n16328) );
  IV U18915 ( .A(n16284), .Z(n16318) );
  XOR U18916 ( .A(n16282), .B(n16331), .Z(n16284) );
  XOR U18917 ( .A(n16332), .B(n16333), .Z(n16331) );
  ANDN U18918 ( .B(n16334), .A(n16335), .Z(n16332) );
  XOR U18919 ( .A(n16336), .B(n16333), .Z(n16334) );
  IV U18920 ( .A(n16286), .Z(n16282) );
  XOR U18921 ( .A(n16337), .B(n16338), .Z(n16286) );
  ANDN U18922 ( .B(n16339), .A(n16340), .Z(n16337) );
  XOR U18923 ( .A(n16341), .B(n16338), .Z(n16339) );
  IV U18924 ( .A(n16296), .Z(n16300) );
  XOR U18925 ( .A(n16296), .B(n16251), .Z(n16298) );
  XOR U18926 ( .A(n16342), .B(n16343), .Z(n16251) );
  AND U18927 ( .A(n198), .B(n16344), .Z(n16342) );
  XOR U18928 ( .A(n16345), .B(n16343), .Z(n16344) );
  NANDN U18929 ( .A(n16253), .B(n16255), .Z(n16296) );
  XOR U18930 ( .A(n16346), .B(n16347), .Z(n16255) );
  AND U18931 ( .A(n198), .B(n16348), .Z(n16346) );
  XOR U18932 ( .A(n16347), .B(n16349), .Z(n16348) );
  XNOR U18933 ( .A(n16350), .B(n16351), .Z(n198) );
  AND U18934 ( .A(n16352), .B(n16353), .Z(n16350) );
  XOR U18935 ( .A(n16351), .B(n16266), .Z(n16353) );
  XNOR U18936 ( .A(n16354), .B(n16355), .Z(n16266) );
  ANDN U18937 ( .B(n16356), .A(n16357), .Z(n16354) );
  XOR U18938 ( .A(n16355), .B(n16358), .Z(n16356) );
  XNOR U18939 ( .A(n16351), .B(n16268), .Z(n16352) );
  XOR U18940 ( .A(n16359), .B(n16360), .Z(n16268) );
  AND U18941 ( .A(n202), .B(n16361), .Z(n16359) );
  XOR U18942 ( .A(n16362), .B(n16360), .Z(n16361) );
  XNOR U18943 ( .A(n16363), .B(n16364), .Z(n16351) );
  AND U18944 ( .A(n16365), .B(n16366), .Z(n16363) );
  XNOR U18945 ( .A(n16364), .B(n16293), .Z(n16366) );
  XOR U18946 ( .A(n16357), .B(n16358), .Z(n16293) );
  XNOR U18947 ( .A(n16367), .B(n16368), .Z(n16358) );
  ANDN U18948 ( .B(n16369), .A(n16370), .Z(n16367) );
  XOR U18949 ( .A(n16371), .B(n16372), .Z(n16369) );
  XOR U18950 ( .A(n16373), .B(n16374), .Z(n16357) );
  XNOR U18951 ( .A(n16375), .B(n16376), .Z(n16374) );
  ANDN U18952 ( .B(n16377), .A(n16378), .Z(n16375) );
  XNOR U18953 ( .A(n16379), .B(n16380), .Z(n16377) );
  IV U18954 ( .A(n16355), .Z(n16373) );
  XOR U18955 ( .A(n16381), .B(n16382), .Z(n16355) );
  ANDN U18956 ( .B(n16383), .A(n16384), .Z(n16381) );
  XOR U18957 ( .A(n16382), .B(n16385), .Z(n16383) );
  XOR U18958 ( .A(n16364), .B(n16295), .Z(n16365) );
  XOR U18959 ( .A(n16386), .B(n16387), .Z(n16295) );
  AND U18960 ( .A(n202), .B(n16388), .Z(n16386) );
  XOR U18961 ( .A(n16389), .B(n16387), .Z(n16388) );
  XNOR U18962 ( .A(n16390), .B(n16391), .Z(n16364) );
  NAND U18963 ( .A(n16392), .B(n16393), .Z(n16391) );
  XOR U18964 ( .A(n16394), .B(n16343), .Z(n16393) );
  XOR U18965 ( .A(n16384), .B(n16385), .Z(n16343) );
  XOR U18966 ( .A(n16395), .B(n16372), .Z(n16385) );
  XOR U18967 ( .A(n16396), .B(n16397), .Z(n16372) );
  ANDN U18968 ( .B(n16398), .A(n16399), .Z(n16396) );
  XOR U18969 ( .A(n16397), .B(n16400), .Z(n16398) );
  IV U18970 ( .A(n16370), .Z(n16395) );
  XOR U18971 ( .A(n16368), .B(n16401), .Z(n16370) );
  XOR U18972 ( .A(n16402), .B(n16403), .Z(n16401) );
  ANDN U18973 ( .B(n16404), .A(n16405), .Z(n16402) );
  XOR U18974 ( .A(n16406), .B(n16403), .Z(n16404) );
  IV U18975 ( .A(n16371), .Z(n16368) );
  XOR U18976 ( .A(n16407), .B(n16408), .Z(n16371) );
  ANDN U18977 ( .B(n16409), .A(n16410), .Z(n16407) );
  XOR U18978 ( .A(n16408), .B(n16411), .Z(n16409) );
  XOR U18979 ( .A(n16412), .B(n16413), .Z(n16384) );
  XNOR U18980 ( .A(n16379), .B(n16414), .Z(n16413) );
  IV U18981 ( .A(n16382), .Z(n16414) );
  XOR U18982 ( .A(n16415), .B(n16416), .Z(n16382) );
  ANDN U18983 ( .B(n16417), .A(n16418), .Z(n16415) );
  XOR U18984 ( .A(n16416), .B(n16419), .Z(n16417) );
  XNOR U18985 ( .A(n16420), .B(n16421), .Z(n16379) );
  ANDN U18986 ( .B(n16422), .A(n16423), .Z(n16420) );
  XOR U18987 ( .A(n16421), .B(n16424), .Z(n16422) );
  IV U18988 ( .A(n16378), .Z(n16412) );
  XOR U18989 ( .A(n16376), .B(n16425), .Z(n16378) );
  XOR U18990 ( .A(n16426), .B(n16427), .Z(n16425) );
  ANDN U18991 ( .B(n16428), .A(n16429), .Z(n16426) );
  XOR U18992 ( .A(n16430), .B(n16427), .Z(n16428) );
  IV U18993 ( .A(n16380), .Z(n16376) );
  XOR U18994 ( .A(n16431), .B(n16432), .Z(n16380) );
  ANDN U18995 ( .B(n16433), .A(n16434), .Z(n16431) );
  XOR U18996 ( .A(n16435), .B(n16432), .Z(n16433) );
  IV U18997 ( .A(n16390), .Z(n16394) );
  XOR U18998 ( .A(n16390), .B(n16345), .Z(n16392) );
  XOR U18999 ( .A(n16436), .B(n16437), .Z(n16345) );
  AND U19000 ( .A(n202), .B(n16438), .Z(n16436) );
  XOR U19001 ( .A(n16439), .B(n16437), .Z(n16438) );
  NANDN U19002 ( .A(n16347), .B(n16349), .Z(n16390) );
  XOR U19003 ( .A(n16440), .B(n16441), .Z(n16349) );
  AND U19004 ( .A(n202), .B(n16442), .Z(n16440) );
  XOR U19005 ( .A(n16441), .B(n16443), .Z(n16442) );
  XNOR U19006 ( .A(n16444), .B(n16445), .Z(n202) );
  AND U19007 ( .A(n16446), .B(n16447), .Z(n16444) );
  XOR U19008 ( .A(n16445), .B(n16360), .Z(n16447) );
  XNOR U19009 ( .A(n16448), .B(n16449), .Z(n16360) );
  ANDN U19010 ( .B(n16450), .A(n16451), .Z(n16448) );
  XOR U19011 ( .A(n16449), .B(n16452), .Z(n16450) );
  XNOR U19012 ( .A(n16445), .B(n16362), .Z(n16446) );
  XOR U19013 ( .A(n16453), .B(n16454), .Z(n16362) );
  AND U19014 ( .A(n206), .B(n16455), .Z(n16453) );
  XOR U19015 ( .A(n16456), .B(n16454), .Z(n16455) );
  XNOR U19016 ( .A(n16457), .B(n16458), .Z(n16445) );
  AND U19017 ( .A(n16459), .B(n16460), .Z(n16457) );
  XNOR U19018 ( .A(n16458), .B(n16387), .Z(n16460) );
  XOR U19019 ( .A(n16451), .B(n16452), .Z(n16387) );
  XNOR U19020 ( .A(n16461), .B(n16462), .Z(n16452) );
  ANDN U19021 ( .B(n16463), .A(n16464), .Z(n16461) );
  XOR U19022 ( .A(n16465), .B(n16466), .Z(n16463) );
  XOR U19023 ( .A(n16467), .B(n16468), .Z(n16451) );
  XNOR U19024 ( .A(n16469), .B(n16470), .Z(n16468) );
  ANDN U19025 ( .B(n16471), .A(n16472), .Z(n16469) );
  XNOR U19026 ( .A(n16473), .B(n16474), .Z(n16471) );
  IV U19027 ( .A(n16449), .Z(n16467) );
  XOR U19028 ( .A(n16475), .B(n16476), .Z(n16449) );
  ANDN U19029 ( .B(n16477), .A(n16478), .Z(n16475) );
  XOR U19030 ( .A(n16476), .B(n16479), .Z(n16477) );
  XOR U19031 ( .A(n16458), .B(n16389), .Z(n16459) );
  XOR U19032 ( .A(n16480), .B(n16481), .Z(n16389) );
  AND U19033 ( .A(n206), .B(n16482), .Z(n16480) );
  XOR U19034 ( .A(n16483), .B(n16481), .Z(n16482) );
  XNOR U19035 ( .A(n16484), .B(n16485), .Z(n16458) );
  NAND U19036 ( .A(n16486), .B(n16487), .Z(n16485) );
  XOR U19037 ( .A(n16488), .B(n16437), .Z(n16487) );
  XOR U19038 ( .A(n16478), .B(n16479), .Z(n16437) );
  XOR U19039 ( .A(n16489), .B(n16466), .Z(n16479) );
  XOR U19040 ( .A(n16490), .B(n16491), .Z(n16466) );
  ANDN U19041 ( .B(n16492), .A(n16493), .Z(n16490) );
  XOR U19042 ( .A(n16491), .B(n16494), .Z(n16492) );
  IV U19043 ( .A(n16464), .Z(n16489) );
  XOR U19044 ( .A(n16462), .B(n16495), .Z(n16464) );
  XOR U19045 ( .A(n16496), .B(n16497), .Z(n16495) );
  ANDN U19046 ( .B(n16498), .A(n16499), .Z(n16496) );
  XOR U19047 ( .A(n16500), .B(n16497), .Z(n16498) );
  IV U19048 ( .A(n16465), .Z(n16462) );
  XOR U19049 ( .A(n16501), .B(n16502), .Z(n16465) );
  ANDN U19050 ( .B(n16503), .A(n16504), .Z(n16501) );
  XOR U19051 ( .A(n16502), .B(n16505), .Z(n16503) );
  XOR U19052 ( .A(n16506), .B(n16507), .Z(n16478) );
  XNOR U19053 ( .A(n16473), .B(n16508), .Z(n16507) );
  IV U19054 ( .A(n16476), .Z(n16508) );
  XOR U19055 ( .A(n16509), .B(n16510), .Z(n16476) );
  ANDN U19056 ( .B(n16511), .A(n16512), .Z(n16509) );
  XOR U19057 ( .A(n16510), .B(n16513), .Z(n16511) );
  XNOR U19058 ( .A(n16514), .B(n16515), .Z(n16473) );
  ANDN U19059 ( .B(n16516), .A(n16517), .Z(n16514) );
  XOR U19060 ( .A(n16515), .B(n16518), .Z(n16516) );
  IV U19061 ( .A(n16472), .Z(n16506) );
  XOR U19062 ( .A(n16470), .B(n16519), .Z(n16472) );
  XOR U19063 ( .A(n16520), .B(n16521), .Z(n16519) );
  ANDN U19064 ( .B(n16522), .A(n16523), .Z(n16520) );
  XOR U19065 ( .A(n16524), .B(n16521), .Z(n16522) );
  IV U19066 ( .A(n16474), .Z(n16470) );
  XOR U19067 ( .A(n16525), .B(n16526), .Z(n16474) );
  ANDN U19068 ( .B(n16527), .A(n16528), .Z(n16525) );
  XOR U19069 ( .A(n16529), .B(n16526), .Z(n16527) );
  IV U19070 ( .A(n16484), .Z(n16488) );
  XOR U19071 ( .A(n16484), .B(n16439), .Z(n16486) );
  XOR U19072 ( .A(n16530), .B(n16531), .Z(n16439) );
  AND U19073 ( .A(n206), .B(n16532), .Z(n16530) );
  XOR U19074 ( .A(n16533), .B(n16531), .Z(n16532) );
  NANDN U19075 ( .A(n16441), .B(n16443), .Z(n16484) );
  XOR U19076 ( .A(n16534), .B(n16535), .Z(n16443) );
  AND U19077 ( .A(n206), .B(n16536), .Z(n16534) );
  XOR U19078 ( .A(n16535), .B(n16537), .Z(n16536) );
  XNOR U19079 ( .A(n16538), .B(n16539), .Z(n206) );
  AND U19080 ( .A(n16540), .B(n16541), .Z(n16538) );
  XOR U19081 ( .A(n16539), .B(n16454), .Z(n16541) );
  XNOR U19082 ( .A(n16542), .B(n16543), .Z(n16454) );
  ANDN U19083 ( .B(n16544), .A(n16545), .Z(n16542) );
  XOR U19084 ( .A(n16543), .B(n16546), .Z(n16544) );
  XNOR U19085 ( .A(n16539), .B(n16456), .Z(n16540) );
  XOR U19086 ( .A(n16547), .B(n16548), .Z(n16456) );
  AND U19087 ( .A(n210), .B(n16549), .Z(n16547) );
  XOR U19088 ( .A(n16550), .B(n16548), .Z(n16549) );
  XNOR U19089 ( .A(n16551), .B(n16552), .Z(n16539) );
  AND U19090 ( .A(n16553), .B(n16554), .Z(n16551) );
  XNOR U19091 ( .A(n16552), .B(n16481), .Z(n16554) );
  XOR U19092 ( .A(n16545), .B(n16546), .Z(n16481) );
  XNOR U19093 ( .A(n16555), .B(n16556), .Z(n16546) );
  ANDN U19094 ( .B(n16557), .A(n16558), .Z(n16555) );
  XOR U19095 ( .A(n16559), .B(n16560), .Z(n16557) );
  XOR U19096 ( .A(n16561), .B(n16562), .Z(n16545) );
  XNOR U19097 ( .A(n16563), .B(n16564), .Z(n16562) );
  ANDN U19098 ( .B(n16565), .A(n16566), .Z(n16563) );
  XNOR U19099 ( .A(n16567), .B(n16568), .Z(n16565) );
  IV U19100 ( .A(n16543), .Z(n16561) );
  XOR U19101 ( .A(n16569), .B(n16570), .Z(n16543) );
  ANDN U19102 ( .B(n16571), .A(n16572), .Z(n16569) );
  XOR U19103 ( .A(n16570), .B(n16573), .Z(n16571) );
  XOR U19104 ( .A(n16552), .B(n16483), .Z(n16553) );
  XOR U19105 ( .A(n16574), .B(n16575), .Z(n16483) );
  AND U19106 ( .A(n210), .B(n16576), .Z(n16574) );
  XOR U19107 ( .A(n16577), .B(n16575), .Z(n16576) );
  XNOR U19108 ( .A(n16578), .B(n16579), .Z(n16552) );
  NAND U19109 ( .A(n16580), .B(n16581), .Z(n16579) );
  XOR U19110 ( .A(n16582), .B(n16531), .Z(n16581) );
  XOR U19111 ( .A(n16572), .B(n16573), .Z(n16531) );
  XOR U19112 ( .A(n16583), .B(n16560), .Z(n16573) );
  XOR U19113 ( .A(n16584), .B(n16585), .Z(n16560) );
  ANDN U19114 ( .B(n16586), .A(n16587), .Z(n16584) );
  XOR U19115 ( .A(n16585), .B(n16588), .Z(n16586) );
  IV U19116 ( .A(n16558), .Z(n16583) );
  XOR U19117 ( .A(n16556), .B(n16589), .Z(n16558) );
  XOR U19118 ( .A(n16590), .B(n16591), .Z(n16589) );
  ANDN U19119 ( .B(n16592), .A(n16593), .Z(n16590) );
  XOR U19120 ( .A(n16594), .B(n16591), .Z(n16592) );
  IV U19121 ( .A(n16559), .Z(n16556) );
  XOR U19122 ( .A(n16595), .B(n16596), .Z(n16559) );
  ANDN U19123 ( .B(n16597), .A(n16598), .Z(n16595) );
  XOR U19124 ( .A(n16596), .B(n16599), .Z(n16597) );
  XOR U19125 ( .A(n16600), .B(n16601), .Z(n16572) );
  XNOR U19126 ( .A(n16567), .B(n16602), .Z(n16601) );
  IV U19127 ( .A(n16570), .Z(n16602) );
  XOR U19128 ( .A(n16603), .B(n16604), .Z(n16570) );
  ANDN U19129 ( .B(n16605), .A(n16606), .Z(n16603) );
  XOR U19130 ( .A(n16604), .B(n16607), .Z(n16605) );
  XNOR U19131 ( .A(n16608), .B(n16609), .Z(n16567) );
  ANDN U19132 ( .B(n16610), .A(n16611), .Z(n16608) );
  XOR U19133 ( .A(n16609), .B(n16612), .Z(n16610) );
  IV U19134 ( .A(n16566), .Z(n16600) );
  XOR U19135 ( .A(n16564), .B(n16613), .Z(n16566) );
  XOR U19136 ( .A(n16614), .B(n16615), .Z(n16613) );
  ANDN U19137 ( .B(n16616), .A(n16617), .Z(n16614) );
  XOR U19138 ( .A(n16618), .B(n16615), .Z(n16616) );
  IV U19139 ( .A(n16568), .Z(n16564) );
  XOR U19140 ( .A(n16619), .B(n16620), .Z(n16568) );
  ANDN U19141 ( .B(n16621), .A(n16622), .Z(n16619) );
  XOR U19142 ( .A(n16623), .B(n16620), .Z(n16621) );
  IV U19143 ( .A(n16578), .Z(n16582) );
  XOR U19144 ( .A(n16578), .B(n16533), .Z(n16580) );
  XOR U19145 ( .A(n16624), .B(n16625), .Z(n16533) );
  AND U19146 ( .A(n210), .B(n16626), .Z(n16624) );
  XOR U19147 ( .A(n16627), .B(n16625), .Z(n16626) );
  NANDN U19148 ( .A(n16535), .B(n16537), .Z(n16578) );
  XOR U19149 ( .A(n16628), .B(n16629), .Z(n16537) );
  AND U19150 ( .A(n210), .B(n16630), .Z(n16628) );
  XOR U19151 ( .A(n16629), .B(n16631), .Z(n16630) );
  XNOR U19152 ( .A(n16632), .B(n16633), .Z(n210) );
  AND U19153 ( .A(n16634), .B(n16635), .Z(n16632) );
  XOR U19154 ( .A(n16633), .B(n16548), .Z(n16635) );
  XNOR U19155 ( .A(n16636), .B(n16637), .Z(n16548) );
  ANDN U19156 ( .B(n16638), .A(n16639), .Z(n16636) );
  XOR U19157 ( .A(n16637), .B(n16640), .Z(n16638) );
  XNOR U19158 ( .A(n16633), .B(n16550), .Z(n16634) );
  XOR U19159 ( .A(n16641), .B(n16642), .Z(n16550) );
  AND U19160 ( .A(n214), .B(n16643), .Z(n16641) );
  XOR U19161 ( .A(n16644), .B(n16642), .Z(n16643) );
  XNOR U19162 ( .A(n16645), .B(n16646), .Z(n16633) );
  AND U19163 ( .A(n16647), .B(n16648), .Z(n16645) );
  XNOR U19164 ( .A(n16646), .B(n16575), .Z(n16648) );
  XOR U19165 ( .A(n16639), .B(n16640), .Z(n16575) );
  XNOR U19166 ( .A(n16649), .B(n16650), .Z(n16640) );
  ANDN U19167 ( .B(n16651), .A(n16652), .Z(n16649) );
  XOR U19168 ( .A(n16653), .B(n16654), .Z(n16651) );
  XOR U19169 ( .A(n16655), .B(n16656), .Z(n16639) );
  XNOR U19170 ( .A(n16657), .B(n16658), .Z(n16656) );
  ANDN U19171 ( .B(n16659), .A(n16660), .Z(n16657) );
  XNOR U19172 ( .A(n16661), .B(n16662), .Z(n16659) );
  IV U19173 ( .A(n16637), .Z(n16655) );
  XOR U19174 ( .A(n16663), .B(n16664), .Z(n16637) );
  ANDN U19175 ( .B(n16665), .A(n16666), .Z(n16663) );
  XOR U19176 ( .A(n16664), .B(n16667), .Z(n16665) );
  XOR U19177 ( .A(n16646), .B(n16577), .Z(n16647) );
  XOR U19178 ( .A(n16668), .B(n16669), .Z(n16577) );
  AND U19179 ( .A(n214), .B(n16670), .Z(n16668) );
  XOR U19180 ( .A(n16671), .B(n16669), .Z(n16670) );
  XNOR U19181 ( .A(n16672), .B(n16673), .Z(n16646) );
  NAND U19182 ( .A(n16674), .B(n16675), .Z(n16673) );
  XOR U19183 ( .A(n16676), .B(n16625), .Z(n16675) );
  XOR U19184 ( .A(n16666), .B(n16667), .Z(n16625) );
  XOR U19185 ( .A(n16677), .B(n16654), .Z(n16667) );
  XOR U19186 ( .A(n16678), .B(n16679), .Z(n16654) );
  ANDN U19187 ( .B(n16680), .A(n16681), .Z(n16678) );
  XOR U19188 ( .A(n16679), .B(n16682), .Z(n16680) );
  IV U19189 ( .A(n16652), .Z(n16677) );
  XOR U19190 ( .A(n16650), .B(n16683), .Z(n16652) );
  XOR U19191 ( .A(n16684), .B(n16685), .Z(n16683) );
  ANDN U19192 ( .B(n16686), .A(n16687), .Z(n16684) );
  XOR U19193 ( .A(n16688), .B(n16685), .Z(n16686) );
  IV U19194 ( .A(n16653), .Z(n16650) );
  XOR U19195 ( .A(n16689), .B(n16690), .Z(n16653) );
  ANDN U19196 ( .B(n16691), .A(n16692), .Z(n16689) );
  XOR U19197 ( .A(n16690), .B(n16693), .Z(n16691) );
  XOR U19198 ( .A(n16694), .B(n16695), .Z(n16666) );
  XNOR U19199 ( .A(n16661), .B(n16696), .Z(n16695) );
  IV U19200 ( .A(n16664), .Z(n16696) );
  XOR U19201 ( .A(n16697), .B(n16698), .Z(n16664) );
  ANDN U19202 ( .B(n16699), .A(n16700), .Z(n16697) );
  XOR U19203 ( .A(n16698), .B(n16701), .Z(n16699) );
  XNOR U19204 ( .A(n16702), .B(n16703), .Z(n16661) );
  ANDN U19205 ( .B(n16704), .A(n16705), .Z(n16702) );
  XOR U19206 ( .A(n16703), .B(n16706), .Z(n16704) );
  IV U19207 ( .A(n16660), .Z(n16694) );
  XOR U19208 ( .A(n16658), .B(n16707), .Z(n16660) );
  XOR U19209 ( .A(n16708), .B(n16709), .Z(n16707) );
  ANDN U19210 ( .B(n16710), .A(n16711), .Z(n16708) );
  XOR U19211 ( .A(n16712), .B(n16709), .Z(n16710) );
  IV U19212 ( .A(n16662), .Z(n16658) );
  XOR U19213 ( .A(n16713), .B(n16714), .Z(n16662) );
  ANDN U19214 ( .B(n16715), .A(n16716), .Z(n16713) );
  XOR U19215 ( .A(n16717), .B(n16714), .Z(n16715) );
  IV U19216 ( .A(n16672), .Z(n16676) );
  XOR U19217 ( .A(n16672), .B(n16627), .Z(n16674) );
  XOR U19218 ( .A(n16718), .B(n16719), .Z(n16627) );
  AND U19219 ( .A(n214), .B(n16720), .Z(n16718) );
  XOR U19220 ( .A(n16721), .B(n16719), .Z(n16720) );
  NANDN U19221 ( .A(n16629), .B(n16631), .Z(n16672) );
  XOR U19222 ( .A(n16722), .B(n16723), .Z(n16631) );
  AND U19223 ( .A(n214), .B(n16724), .Z(n16722) );
  XOR U19224 ( .A(n16723), .B(n16725), .Z(n16724) );
  XNOR U19225 ( .A(n16726), .B(n16727), .Z(n214) );
  AND U19226 ( .A(n16728), .B(n16729), .Z(n16726) );
  XOR U19227 ( .A(n16727), .B(n16642), .Z(n16729) );
  XNOR U19228 ( .A(n16730), .B(n16731), .Z(n16642) );
  ANDN U19229 ( .B(n16732), .A(n16733), .Z(n16730) );
  XOR U19230 ( .A(n16731), .B(n16734), .Z(n16732) );
  XNOR U19231 ( .A(n16727), .B(n16644), .Z(n16728) );
  XOR U19232 ( .A(n16735), .B(n16736), .Z(n16644) );
  AND U19233 ( .A(n218), .B(n16737), .Z(n16735) );
  XOR U19234 ( .A(n16738), .B(n16736), .Z(n16737) );
  XNOR U19235 ( .A(n16739), .B(n16740), .Z(n16727) );
  AND U19236 ( .A(n16741), .B(n16742), .Z(n16739) );
  XNOR U19237 ( .A(n16740), .B(n16669), .Z(n16742) );
  XOR U19238 ( .A(n16733), .B(n16734), .Z(n16669) );
  XNOR U19239 ( .A(n16743), .B(n16744), .Z(n16734) );
  ANDN U19240 ( .B(n16745), .A(n16746), .Z(n16743) );
  XOR U19241 ( .A(n16747), .B(n16748), .Z(n16745) );
  XOR U19242 ( .A(n16749), .B(n16750), .Z(n16733) );
  XNOR U19243 ( .A(n16751), .B(n16752), .Z(n16750) );
  ANDN U19244 ( .B(n16753), .A(n16754), .Z(n16751) );
  XNOR U19245 ( .A(n16755), .B(n16756), .Z(n16753) );
  IV U19246 ( .A(n16731), .Z(n16749) );
  XOR U19247 ( .A(n16757), .B(n16758), .Z(n16731) );
  ANDN U19248 ( .B(n16759), .A(n16760), .Z(n16757) );
  XOR U19249 ( .A(n16758), .B(n16761), .Z(n16759) );
  XOR U19250 ( .A(n16740), .B(n16671), .Z(n16741) );
  XOR U19251 ( .A(n16762), .B(n16763), .Z(n16671) );
  AND U19252 ( .A(n218), .B(n16764), .Z(n16762) );
  XOR U19253 ( .A(n16765), .B(n16763), .Z(n16764) );
  XNOR U19254 ( .A(n16766), .B(n16767), .Z(n16740) );
  NAND U19255 ( .A(n16768), .B(n16769), .Z(n16767) );
  XOR U19256 ( .A(n16770), .B(n16719), .Z(n16769) );
  XOR U19257 ( .A(n16760), .B(n16761), .Z(n16719) );
  XOR U19258 ( .A(n16771), .B(n16748), .Z(n16761) );
  XOR U19259 ( .A(n16772), .B(n16773), .Z(n16748) );
  ANDN U19260 ( .B(n16774), .A(n16775), .Z(n16772) );
  XOR U19261 ( .A(n16773), .B(n16776), .Z(n16774) );
  IV U19262 ( .A(n16746), .Z(n16771) );
  XOR U19263 ( .A(n16744), .B(n16777), .Z(n16746) );
  XOR U19264 ( .A(n16778), .B(n16779), .Z(n16777) );
  ANDN U19265 ( .B(n16780), .A(n16781), .Z(n16778) );
  XOR U19266 ( .A(n16782), .B(n16779), .Z(n16780) );
  IV U19267 ( .A(n16747), .Z(n16744) );
  XOR U19268 ( .A(n16783), .B(n16784), .Z(n16747) );
  ANDN U19269 ( .B(n16785), .A(n16786), .Z(n16783) );
  XOR U19270 ( .A(n16784), .B(n16787), .Z(n16785) );
  XOR U19271 ( .A(n16788), .B(n16789), .Z(n16760) );
  XNOR U19272 ( .A(n16755), .B(n16790), .Z(n16789) );
  IV U19273 ( .A(n16758), .Z(n16790) );
  XOR U19274 ( .A(n16791), .B(n16792), .Z(n16758) );
  ANDN U19275 ( .B(n16793), .A(n16794), .Z(n16791) );
  XOR U19276 ( .A(n16792), .B(n16795), .Z(n16793) );
  XNOR U19277 ( .A(n16796), .B(n16797), .Z(n16755) );
  ANDN U19278 ( .B(n16798), .A(n16799), .Z(n16796) );
  XOR U19279 ( .A(n16797), .B(n16800), .Z(n16798) );
  IV U19280 ( .A(n16754), .Z(n16788) );
  XOR U19281 ( .A(n16752), .B(n16801), .Z(n16754) );
  XOR U19282 ( .A(n16802), .B(n16803), .Z(n16801) );
  ANDN U19283 ( .B(n16804), .A(n16805), .Z(n16802) );
  XOR U19284 ( .A(n16806), .B(n16803), .Z(n16804) );
  IV U19285 ( .A(n16756), .Z(n16752) );
  XOR U19286 ( .A(n16807), .B(n16808), .Z(n16756) );
  ANDN U19287 ( .B(n16809), .A(n16810), .Z(n16807) );
  XOR U19288 ( .A(n16811), .B(n16808), .Z(n16809) );
  IV U19289 ( .A(n16766), .Z(n16770) );
  XOR U19290 ( .A(n16766), .B(n16721), .Z(n16768) );
  XOR U19291 ( .A(n16812), .B(n16813), .Z(n16721) );
  AND U19292 ( .A(n218), .B(n16814), .Z(n16812) );
  XOR U19293 ( .A(n16815), .B(n16813), .Z(n16814) );
  NANDN U19294 ( .A(n16723), .B(n16725), .Z(n16766) );
  XOR U19295 ( .A(n16816), .B(n16817), .Z(n16725) );
  AND U19296 ( .A(n218), .B(n16818), .Z(n16816) );
  XOR U19297 ( .A(n16817), .B(n16819), .Z(n16818) );
  XNOR U19298 ( .A(n16820), .B(n16821), .Z(n218) );
  AND U19299 ( .A(n16822), .B(n16823), .Z(n16820) );
  XOR U19300 ( .A(n16821), .B(n16736), .Z(n16823) );
  XNOR U19301 ( .A(n16824), .B(n16825), .Z(n16736) );
  ANDN U19302 ( .B(n16826), .A(n16827), .Z(n16824) );
  XOR U19303 ( .A(n16825), .B(n16828), .Z(n16826) );
  XNOR U19304 ( .A(n16821), .B(n16738), .Z(n16822) );
  XOR U19305 ( .A(n16829), .B(n16830), .Z(n16738) );
  AND U19306 ( .A(n222), .B(n16831), .Z(n16829) );
  XOR U19307 ( .A(n16832), .B(n16830), .Z(n16831) );
  XNOR U19308 ( .A(n16833), .B(n16834), .Z(n16821) );
  AND U19309 ( .A(n16835), .B(n16836), .Z(n16833) );
  XNOR U19310 ( .A(n16834), .B(n16763), .Z(n16836) );
  XOR U19311 ( .A(n16827), .B(n16828), .Z(n16763) );
  XNOR U19312 ( .A(n16837), .B(n16838), .Z(n16828) );
  ANDN U19313 ( .B(n16839), .A(n16840), .Z(n16837) );
  XOR U19314 ( .A(n16841), .B(n16842), .Z(n16839) );
  XOR U19315 ( .A(n16843), .B(n16844), .Z(n16827) );
  XNOR U19316 ( .A(n16845), .B(n16846), .Z(n16844) );
  ANDN U19317 ( .B(n16847), .A(n16848), .Z(n16845) );
  XNOR U19318 ( .A(n16849), .B(n16850), .Z(n16847) );
  IV U19319 ( .A(n16825), .Z(n16843) );
  XOR U19320 ( .A(n16851), .B(n16852), .Z(n16825) );
  ANDN U19321 ( .B(n16853), .A(n16854), .Z(n16851) );
  XOR U19322 ( .A(n16852), .B(n16855), .Z(n16853) );
  XOR U19323 ( .A(n16834), .B(n16765), .Z(n16835) );
  XOR U19324 ( .A(n16856), .B(n16857), .Z(n16765) );
  AND U19325 ( .A(n222), .B(n16858), .Z(n16856) );
  XOR U19326 ( .A(n16859), .B(n16857), .Z(n16858) );
  XNOR U19327 ( .A(n16860), .B(n16861), .Z(n16834) );
  NAND U19328 ( .A(n16862), .B(n16863), .Z(n16861) );
  XOR U19329 ( .A(n16864), .B(n16813), .Z(n16863) );
  XOR U19330 ( .A(n16854), .B(n16855), .Z(n16813) );
  XOR U19331 ( .A(n16865), .B(n16842), .Z(n16855) );
  XOR U19332 ( .A(n16866), .B(n16867), .Z(n16842) );
  ANDN U19333 ( .B(n16868), .A(n16869), .Z(n16866) );
  XOR U19334 ( .A(n16867), .B(n16870), .Z(n16868) );
  IV U19335 ( .A(n16840), .Z(n16865) );
  XOR U19336 ( .A(n16838), .B(n16871), .Z(n16840) );
  XOR U19337 ( .A(n16872), .B(n16873), .Z(n16871) );
  ANDN U19338 ( .B(n16874), .A(n16875), .Z(n16872) );
  XOR U19339 ( .A(n16876), .B(n16873), .Z(n16874) );
  IV U19340 ( .A(n16841), .Z(n16838) );
  XOR U19341 ( .A(n16877), .B(n16878), .Z(n16841) );
  ANDN U19342 ( .B(n16879), .A(n16880), .Z(n16877) );
  XOR U19343 ( .A(n16878), .B(n16881), .Z(n16879) );
  XOR U19344 ( .A(n16882), .B(n16883), .Z(n16854) );
  XNOR U19345 ( .A(n16849), .B(n16884), .Z(n16883) );
  IV U19346 ( .A(n16852), .Z(n16884) );
  XOR U19347 ( .A(n16885), .B(n16886), .Z(n16852) );
  ANDN U19348 ( .B(n16887), .A(n16888), .Z(n16885) );
  XOR U19349 ( .A(n16886), .B(n16889), .Z(n16887) );
  XNOR U19350 ( .A(n16890), .B(n16891), .Z(n16849) );
  ANDN U19351 ( .B(n16892), .A(n16893), .Z(n16890) );
  XOR U19352 ( .A(n16891), .B(n16894), .Z(n16892) );
  IV U19353 ( .A(n16848), .Z(n16882) );
  XOR U19354 ( .A(n16846), .B(n16895), .Z(n16848) );
  XOR U19355 ( .A(n16896), .B(n16897), .Z(n16895) );
  ANDN U19356 ( .B(n16898), .A(n16899), .Z(n16896) );
  XOR U19357 ( .A(n16900), .B(n16897), .Z(n16898) );
  IV U19358 ( .A(n16850), .Z(n16846) );
  XOR U19359 ( .A(n16901), .B(n16902), .Z(n16850) );
  ANDN U19360 ( .B(n16903), .A(n16904), .Z(n16901) );
  XOR U19361 ( .A(n16905), .B(n16902), .Z(n16903) );
  IV U19362 ( .A(n16860), .Z(n16864) );
  XOR U19363 ( .A(n16860), .B(n16815), .Z(n16862) );
  XOR U19364 ( .A(n16906), .B(n16907), .Z(n16815) );
  AND U19365 ( .A(n222), .B(n16908), .Z(n16906) );
  XOR U19366 ( .A(n16909), .B(n16907), .Z(n16908) );
  NANDN U19367 ( .A(n16817), .B(n16819), .Z(n16860) );
  XOR U19368 ( .A(n16910), .B(n16911), .Z(n16819) );
  AND U19369 ( .A(n222), .B(n16912), .Z(n16910) );
  XOR U19370 ( .A(n16911), .B(n16913), .Z(n16912) );
  XNOR U19371 ( .A(n16914), .B(n16915), .Z(n222) );
  AND U19372 ( .A(n16916), .B(n16917), .Z(n16914) );
  XOR U19373 ( .A(n16915), .B(n16830), .Z(n16917) );
  XNOR U19374 ( .A(n16918), .B(n16919), .Z(n16830) );
  ANDN U19375 ( .B(n16920), .A(n16921), .Z(n16918) );
  XOR U19376 ( .A(n16919), .B(n16922), .Z(n16920) );
  XNOR U19377 ( .A(n16915), .B(n16832), .Z(n16916) );
  XOR U19378 ( .A(n16923), .B(n16924), .Z(n16832) );
  AND U19379 ( .A(n226), .B(n16925), .Z(n16923) );
  XOR U19380 ( .A(n16926), .B(n16924), .Z(n16925) );
  XNOR U19381 ( .A(n16927), .B(n16928), .Z(n16915) );
  AND U19382 ( .A(n16929), .B(n16930), .Z(n16927) );
  XNOR U19383 ( .A(n16928), .B(n16857), .Z(n16930) );
  XOR U19384 ( .A(n16921), .B(n16922), .Z(n16857) );
  XNOR U19385 ( .A(n16931), .B(n16932), .Z(n16922) );
  ANDN U19386 ( .B(n16933), .A(n16934), .Z(n16931) );
  XOR U19387 ( .A(n16935), .B(n16936), .Z(n16933) );
  XOR U19388 ( .A(n16937), .B(n16938), .Z(n16921) );
  XNOR U19389 ( .A(n16939), .B(n16940), .Z(n16938) );
  ANDN U19390 ( .B(n16941), .A(n16942), .Z(n16939) );
  XNOR U19391 ( .A(n16943), .B(n16944), .Z(n16941) );
  IV U19392 ( .A(n16919), .Z(n16937) );
  XOR U19393 ( .A(n16945), .B(n16946), .Z(n16919) );
  ANDN U19394 ( .B(n16947), .A(n16948), .Z(n16945) );
  XOR U19395 ( .A(n16946), .B(n16949), .Z(n16947) );
  XOR U19396 ( .A(n16928), .B(n16859), .Z(n16929) );
  XOR U19397 ( .A(n16950), .B(n16951), .Z(n16859) );
  AND U19398 ( .A(n226), .B(n16952), .Z(n16950) );
  XOR U19399 ( .A(n16953), .B(n16951), .Z(n16952) );
  XNOR U19400 ( .A(n16954), .B(n16955), .Z(n16928) );
  NAND U19401 ( .A(n16956), .B(n16957), .Z(n16955) );
  XOR U19402 ( .A(n16958), .B(n16907), .Z(n16957) );
  XOR U19403 ( .A(n16948), .B(n16949), .Z(n16907) );
  XOR U19404 ( .A(n16959), .B(n16936), .Z(n16949) );
  XOR U19405 ( .A(n16960), .B(n16961), .Z(n16936) );
  ANDN U19406 ( .B(n16962), .A(n16963), .Z(n16960) );
  XOR U19407 ( .A(n16961), .B(n16964), .Z(n16962) );
  IV U19408 ( .A(n16934), .Z(n16959) );
  XOR U19409 ( .A(n16932), .B(n16965), .Z(n16934) );
  XOR U19410 ( .A(n16966), .B(n16967), .Z(n16965) );
  ANDN U19411 ( .B(n16968), .A(n16969), .Z(n16966) );
  XOR U19412 ( .A(n16970), .B(n16967), .Z(n16968) );
  IV U19413 ( .A(n16935), .Z(n16932) );
  XOR U19414 ( .A(n16971), .B(n16972), .Z(n16935) );
  ANDN U19415 ( .B(n16973), .A(n16974), .Z(n16971) );
  XOR U19416 ( .A(n16972), .B(n16975), .Z(n16973) );
  XOR U19417 ( .A(n16976), .B(n16977), .Z(n16948) );
  XNOR U19418 ( .A(n16943), .B(n16978), .Z(n16977) );
  IV U19419 ( .A(n16946), .Z(n16978) );
  XOR U19420 ( .A(n16979), .B(n16980), .Z(n16946) );
  ANDN U19421 ( .B(n16981), .A(n16982), .Z(n16979) );
  XOR U19422 ( .A(n16980), .B(n16983), .Z(n16981) );
  XNOR U19423 ( .A(n16984), .B(n16985), .Z(n16943) );
  ANDN U19424 ( .B(n16986), .A(n16987), .Z(n16984) );
  XOR U19425 ( .A(n16985), .B(n16988), .Z(n16986) );
  IV U19426 ( .A(n16942), .Z(n16976) );
  XOR U19427 ( .A(n16940), .B(n16989), .Z(n16942) );
  XOR U19428 ( .A(n16990), .B(n16991), .Z(n16989) );
  ANDN U19429 ( .B(n16992), .A(n16993), .Z(n16990) );
  XOR U19430 ( .A(n16994), .B(n16991), .Z(n16992) );
  IV U19431 ( .A(n16944), .Z(n16940) );
  XOR U19432 ( .A(n16995), .B(n16996), .Z(n16944) );
  ANDN U19433 ( .B(n16997), .A(n16998), .Z(n16995) );
  XOR U19434 ( .A(n16999), .B(n16996), .Z(n16997) );
  IV U19435 ( .A(n16954), .Z(n16958) );
  XOR U19436 ( .A(n16954), .B(n16909), .Z(n16956) );
  XOR U19437 ( .A(n17000), .B(n17001), .Z(n16909) );
  AND U19438 ( .A(n226), .B(n17002), .Z(n17000) );
  XOR U19439 ( .A(n17003), .B(n17001), .Z(n17002) );
  NANDN U19440 ( .A(n16911), .B(n16913), .Z(n16954) );
  XOR U19441 ( .A(n17004), .B(n17005), .Z(n16913) );
  AND U19442 ( .A(n226), .B(n17006), .Z(n17004) );
  XOR U19443 ( .A(n17005), .B(n17007), .Z(n17006) );
  XNOR U19444 ( .A(n17008), .B(n17009), .Z(n226) );
  AND U19445 ( .A(n17010), .B(n17011), .Z(n17008) );
  XOR U19446 ( .A(n17009), .B(n16924), .Z(n17011) );
  XNOR U19447 ( .A(n17012), .B(n17013), .Z(n16924) );
  ANDN U19448 ( .B(n17014), .A(n17015), .Z(n17012) );
  XOR U19449 ( .A(n17013), .B(n17016), .Z(n17014) );
  XNOR U19450 ( .A(n17009), .B(n16926), .Z(n17010) );
  XOR U19451 ( .A(n17017), .B(n17018), .Z(n16926) );
  AND U19452 ( .A(n230), .B(n17019), .Z(n17017) );
  XOR U19453 ( .A(n17020), .B(n17018), .Z(n17019) );
  XNOR U19454 ( .A(n17021), .B(n17022), .Z(n17009) );
  AND U19455 ( .A(n17023), .B(n17024), .Z(n17021) );
  XNOR U19456 ( .A(n17022), .B(n16951), .Z(n17024) );
  XOR U19457 ( .A(n17015), .B(n17016), .Z(n16951) );
  XNOR U19458 ( .A(n17025), .B(n17026), .Z(n17016) );
  ANDN U19459 ( .B(n17027), .A(n17028), .Z(n17025) );
  XOR U19460 ( .A(n17029), .B(n17030), .Z(n17027) );
  XOR U19461 ( .A(n17031), .B(n17032), .Z(n17015) );
  XNOR U19462 ( .A(n17033), .B(n17034), .Z(n17032) );
  ANDN U19463 ( .B(n17035), .A(n17036), .Z(n17033) );
  XNOR U19464 ( .A(n17037), .B(n17038), .Z(n17035) );
  IV U19465 ( .A(n17013), .Z(n17031) );
  XOR U19466 ( .A(n17039), .B(n17040), .Z(n17013) );
  ANDN U19467 ( .B(n17041), .A(n17042), .Z(n17039) );
  XOR U19468 ( .A(n17040), .B(n17043), .Z(n17041) );
  XOR U19469 ( .A(n17022), .B(n16953), .Z(n17023) );
  XOR U19470 ( .A(n17044), .B(n17045), .Z(n16953) );
  AND U19471 ( .A(n230), .B(n17046), .Z(n17044) );
  XOR U19472 ( .A(n17047), .B(n17045), .Z(n17046) );
  XNOR U19473 ( .A(n17048), .B(n17049), .Z(n17022) );
  NAND U19474 ( .A(n17050), .B(n17051), .Z(n17049) );
  XOR U19475 ( .A(n17052), .B(n17001), .Z(n17051) );
  XOR U19476 ( .A(n17042), .B(n17043), .Z(n17001) );
  XOR U19477 ( .A(n17053), .B(n17030), .Z(n17043) );
  XOR U19478 ( .A(n17054), .B(n17055), .Z(n17030) );
  ANDN U19479 ( .B(n17056), .A(n17057), .Z(n17054) );
  XOR U19480 ( .A(n17055), .B(n17058), .Z(n17056) );
  IV U19481 ( .A(n17028), .Z(n17053) );
  XOR U19482 ( .A(n17026), .B(n17059), .Z(n17028) );
  XOR U19483 ( .A(n17060), .B(n17061), .Z(n17059) );
  ANDN U19484 ( .B(n17062), .A(n17063), .Z(n17060) );
  XOR U19485 ( .A(n17064), .B(n17061), .Z(n17062) );
  IV U19486 ( .A(n17029), .Z(n17026) );
  XOR U19487 ( .A(n17065), .B(n17066), .Z(n17029) );
  ANDN U19488 ( .B(n17067), .A(n17068), .Z(n17065) );
  XOR U19489 ( .A(n17066), .B(n17069), .Z(n17067) );
  XOR U19490 ( .A(n17070), .B(n17071), .Z(n17042) );
  XNOR U19491 ( .A(n17037), .B(n17072), .Z(n17071) );
  IV U19492 ( .A(n17040), .Z(n17072) );
  XOR U19493 ( .A(n17073), .B(n17074), .Z(n17040) );
  ANDN U19494 ( .B(n17075), .A(n17076), .Z(n17073) );
  XOR U19495 ( .A(n17074), .B(n17077), .Z(n17075) );
  XNOR U19496 ( .A(n17078), .B(n17079), .Z(n17037) );
  ANDN U19497 ( .B(n17080), .A(n17081), .Z(n17078) );
  XOR U19498 ( .A(n17079), .B(n17082), .Z(n17080) );
  IV U19499 ( .A(n17036), .Z(n17070) );
  XOR U19500 ( .A(n17034), .B(n17083), .Z(n17036) );
  XOR U19501 ( .A(n17084), .B(n17085), .Z(n17083) );
  ANDN U19502 ( .B(n17086), .A(n17087), .Z(n17084) );
  XOR U19503 ( .A(n17088), .B(n17085), .Z(n17086) );
  IV U19504 ( .A(n17038), .Z(n17034) );
  XOR U19505 ( .A(n17089), .B(n17090), .Z(n17038) );
  ANDN U19506 ( .B(n17091), .A(n17092), .Z(n17089) );
  XOR U19507 ( .A(n17093), .B(n17090), .Z(n17091) );
  IV U19508 ( .A(n17048), .Z(n17052) );
  XOR U19509 ( .A(n17048), .B(n17003), .Z(n17050) );
  XOR U19510 ( .A(n17094), .B(n17095), .Z(n17003) );
  AND U19511 ( .A(n230), .B(n17096), .Z(n17094) );
  XOR U19512 ( .A(n17097), .B(n17095), .Z(n17096) );
  NANDN U19513 ( .A(n17005), .B(n17007), .Z(n17048) );
  XOR U19514 ( .A(n17098), .B(n17099), .Z(n17007) );
  AND U19515 ( .A(n230), .B(n17100), .Z(n17098) );
  XOR U19516 ( .A(n17099), .B(n17101), .Z(n17100) );
  XNOR U19517 ( .A(n17102), .B(n17103), .Z(n230) );
  AND U19518 ( .A(n17104), .B(n17105), .Z(n17102) );
  XOR U19519 ( .A(n17103), .B(n17018), .Z(n17105) );
  XNOR U19520 ( .A(n17106), .B(n17107), .Z(n17018) );
  ANDN U19521 ( .B(n17108), .A(n17109), .Z(n17106) );
  XOR U19522 ( .A(n17107), .B(n17110), .Z(n17108) );
  XNOR U19523 ( .A(n17103), .B(n17020), .Z(n17104) );
  XOR U19524 ( .A(n17111), .B(n17112), .Z(n17020) );
  AND U19525 ( .A(n234), .B(n17113), .Z(n17111) );
  XOR U19526 ( .A(n17114), .B(n17112), .Z(n17113) );
  XNOR U19527 ( .A(n17115), .B(n17116), .Z(n17103) );
  AND U19528 ( .A(n17117), .B(n17118), .Z(n17115) );
  XNOR U19529 ( .A(n17116), .B(n17045), .Z(n17118) );
  XOR U19530 ( .A(n17109), .B(n17110), .Z(n17045) );
  XNOR U19531 ( .A(n17119), .B(n17120), .Z(n17110) );
  ANDN U19532 ( .B(n17121), .A(n17122), .Z(n17119) );
  XOR U19533 ( .A(n17123), .B(n17124), .Z(n17121) );
  XOR U19534 ( .A(n17125), .B(n17126), .Z(n17109) );
  XNOR U19535 ( .A(n17127), .B(n17128), .Z(n17126) );
  ANDN U19536 ( .B(n17129), .A(n17130), .Z(n17127) );
  XNOR U19537 ( .A(n17131), .B(n17132), .Z(n17129) );
  IV U19538 ( .A(n17107), .Z(n17125) );
  XOR U19539 ( .A(n17133), .B(n17134), .Z(n17107) );
  ANDN U19540 ( .B(n17135), .A(n17136), .Z(n17133) );
  XOR U19541 ( .A(n17134), .B(n17137), .Z(n17135) );
  XOR U19542 ( .A(n17116), .B(n17047), .Z(n17117) );
  XOR U19543 ( .A(n17138), .B(n17139), .Z(n17047) );
  AND U19544 ( .A(n234), .B(n17140), .Z(n17138) );
  XOR U19545 ( .A(n17141), .B(n17139), .Z(n17140) );
  XNOR U19546 ( .A(n17142), .B(n17143), .Z(n17116) );
  NAND U19547 ( .A(n17144), .B(n17145), .Z(n17143) );
  XOR U19548 ( .A(n17146), .B(n17095), .Z(n17145) );
  XOR U19549 ( .A(n17136), .B(n17137), .Z(n17095) );
  XOR U19550 ( .A(n17147), .B(n17124), .Z(n17137) );
  XOR U19551 ( .A(n17148), .B(n17149), .Z(n17124) );
  ANDN U19552 ( .B(n17150), .A(n17151), .Z(n17148) );
  XOR U19553 ( .A(n17149), .B(n17152), .Z(n17150) );
  IV U19554 ( .A(n17122), .Z(n17147) );
  XOR U19555 ( .A(n17120), .B(n17153), .Z(n17122) );
  XOR U19556 ( .A(n17154), .B(n17155), .Z(n17153) );
  ANDN U19557 ( .B(n17156), .A(n17157), .Z(n17154) );
  XOR U19558 ( .A(n17158), .B(n17155), .Z(n17156) );
  IV U19559 ( .A(n17123), .Z(n17120) );
  XOR U19560 ( .A(n17159), .B(n17160), .Z(n17123) );
  ANDN U19561 ( .B(n17161), .A(n17162), .Z(n17159) );
  XOR U19562 ( .A(n17160), .B(n17163), .Z(n17161) );
  XOR U19563 ( .A(n17164), .B(n17165), .Z(n17136) );
  XNOR U19564 ( .A(n17131), .B(n17166), .Z(n17165) );
  IV U19565 ( .A(n17134), .Z(n17166) );
  XOR U19566 ( .A(n17167), .B(n17168), .Z(n17134) );
  ANDN U19567 ( .B(n17169), .A(n17170), .Z(n17167) );
  XOR U19568 ( .A(n17168), .B(n17171), .Z(n17169) );
  XNOR U19569 ( .A(n17172), .B(n17173), .Z(n17131) );
  ANDN U19570 ( .B(n17174), .A(n17175), .Z(n17172) );
  XOR U19571 ( .A(n17173), .B(n17176), .Z(n17174) );
  IV U19572 ( .A(n17130), .Z(n17164) );
  XOR U19573 ( .A(n17128), .B(n17177), .Z(n17130) );
  XOR U19574 ( .A(n17178), .B(n17179), .Z(n17177) );
  ANDN U19575 ( .B(n17180), .A(n17181), .Z(n17178) );
  XOR U19576 ( .A(n17182), .B(n17179), .Z(n17180) );
  IV U19577 ( .A(n17132), .Z(n17128) );
  XOR U19578 ( .A(n17183), .B(n17184), .Z(n17132) );
  ANDN U19579 ( .B(n17185), .A(n17186), .Z(n17183) );
  XOR U19580 ( .A(n17187), .B(n17184), .Z(n17185) );
  IV U19581 ( .A(n17142), .Z(n17146) );
  XOR U19582 ( .A(n17142), .B(n17097), .Z(n17144) );
  XOR U19583 ( .A(n17188), .B(n17189), .Z(n17097) );
  AND U19584 ( .A(n234), .B(n17190), .Z(n17188) );
  XOR U19585 ( .A(n17191), .B(n17189), .Z(n17190) );
  NANDN U19586 ( .A(n17099), .B(n17101), .Z(n17142) );
  XOR U19587 ( .A(n17192), .B(n17193), .Z(n17101) );
  AND U19588 ( .A(n234), .B(n17194), .Z(n17192) );
  XOR U19589 ( .A(n17193), .B(n17195), .Z(n17194) );
  XNOR U19590 ( .A(n17196), .B(n17197), .Z(n234) );
  AND U19591 ( .A(n17198), .B(n17199), .Z(n17196) );
  XOR U19592 ( .A(n17197), .B(n17112), .Z(n17199) );
  XNOR U19593 ( .A(n17200), .B(n17201), .Z(n17112) );
  ANDN U19594 ( .B(n17202), .A(n17203), .Z(n17200) );
  XOR U19595 ( .A(n17201), .B(n17204), .Z(n17202) );
  XNOR U19596 ( .A(n17197), .B(n17114), .Z(n17198) );
  XOR U19597 ( .A(n17205), .B(n17206), .Z(n17114) );
  AND U19598 ( .A(n238), .B(n17207), .Z(n17205) );
  XOR U19599 ( .A(n17208), .B(n17206), .Z(n17207) );
  XNOR U19600 ( .A(n17209), .B(n17210), .Z(n17197) );
  AND U19601 ( .A(n17211), .B(n17212), .Z(n17209) );
  XNOR U19602 ( .A(n17210), .B(n17139), .Z(n17212) );
  XOR U19603 ( .A(n17203), .B(n17204), .Z(n17139) );
  XNOR U19604 ( .A(n17213), .B(n17214), .Z(n17204) );
  ANDN U19605 ( .B(n17215), .A(n17216), .Z(n17213) );
  XOR U19606 ( .A(n17217), .B(n17218), .Z(n17215) );
  XOR U19607 ( .A(n17219), .B(n17220), .Z(n17203) );
  XNOR U19608 ( .A(n17221), .B(n17222), .Z(n17220) );
  ANDN U19609 ( .B(n17223), .A(n17224), .Z(n17221) );
  XNOR U19610 ( .A(n17225), .B(n17226), .Z(n17223) );
  IV U19611 ( .A(n17201), .Z(n17219) );
  XOR U19612 ( .A(n17227), .B(n17228), .Z(n17201) );
  ANDN U19613 ( .B(n17229), .A(n17230), .Z(n17227) );
  XOR U19614 ( .A(n17228), .B(n17231), .Z(n17229) );
  XOR U19615 ( .A(n17210), .B(n17141), .Z(n17211) );
  XOR U19616 ( .A(n17232), .B(n17233), .Z(n17141) );
  AND U19617 ( .A(n238), .B(n17234), .Z(n17232) );
  XOR U19618 ( .A(n17235), .B(n17233), .Z(n17234) );
  XNOR U19619 ( .A(n17236), .B(n17237), .Z(n17210) );
  NAND U19620 ( .A(n17238), .B(n17239), .Z(n17237) );
  XOR U19621 ( .A(n17240), .B(n17189), .Z(n17239) );
  XOR U19622 ( .A(n17230), .B(n17231), .Z(n17189) );
  XOR U19623 ( .A(n17241), .B(n17218), .Z(n17231) );
  XOR U19624 ( .A(n17242), .B(n17243), .Z(n17218) );
  ANDN U19625 ( .B(n17244), .A(n17245), .Z(n17242) );
  XOR U19626 ( .A(n17243), .B(n17246), .Z(n17244) );
  IV U19627 ( .A(n17216), .Z(n17241) );
  XOR U19628 ( .A(n17214), .B(n17247), .Z(n17216) );
  XOR U19629 ( .A(n17248), .B(n17249), .Z(n17247) );
  ANDN U19630 ( .B(n17250), .A(n17251), .Z(n17248) );
  XOR U19631 ( .A(n17252), .B(n17249), .Z(n17250) );
  IV U19632 ( .A(n17217), .Z(n17214) );
  XOR U19633 ( .A(n17253), .B(n17254), .Z(n17217) );
  ANDN U19634 ( .B(n17255), .A(n17256), .Z(n17253) );
  XOR U19635 ( .A(n17254), .B(n17257), .Z(n17255) );
  XOR U19636 ( .A(n17258), .B(n17259), .Z(n17230) );
  XNOR U19637 ( .A(n17225), .B(n17260), .Z(n17259) );
  IV U19638 ( .A(n17228), .Z(n17260) );
  XOR U19639 ( .A(n17261), .B(n17262), .Z(n17228) );
  ANDN U19640 ( .B(n17263), .A(n17264), .Z(n17261) );
  XOR U19641 ( .A(n17262), .B(n17265), .Z(n17263) );
  XNOR U19642 ( .A(n17266), .B(n17267), .Z(n17225) );
  ANDN U19643 ( .B(n17268), .A(n17269), .Z(n17266) );
  XOR U19644 ( .A(n17267), .B(n17270), .Z(n17268) );
  IV U19645 ( .A(n17224), .Z(n17258) );
  XOR U19646 ( .A(n17222), .B(n17271), .Z(n17224) );
  XOR U19647 ( .A(n17272), .B(n17273), .Z(n17271) );
  ANDN U19648 ( .B(n17274), .A(n17275), .Z(n17272) );
  XOR U19649 ( .A(n17276), .B(n17273), .Z(n17274) );
  IV U19650 ( .A(n17226), .Z(n17222) );
  XOR U19651 ( .A(n17277), .B(n17278), .Z(n17226) );
  ANDN U19652 ( .B(n17279), .A(n17280), .Z(n17277) );
  XOR U19653 ( .A(n17281), .B(n17278), .Z(n17279) );
  IV U19654 ( .A(n17236), .Z(n17240) );
  XOR U19655 ( .A(n17236), .B(n17191), .Z(n17238) );
  XOR U19656 ( .A(n17282), .B(n17283), .Z(n17191) );
  AND U19657 ( .A(n238), .B(n17284), .Z(n17282) );
  XOR U19658 ( .A(n17285), .B(n17283), .Z(n17284) );
  NANDN U19659 ( .A(n17193), .B(n17195), .Z(n17236) );
  XOR U19660 ( .A(n17286), .B(n17287), .Z(n17195) );
  AND U19661 ( .A(n238), .B(n17288), .Z(n17286) );
  XOR U19662 ( .A(n17287), .B(n17289), .Z(n17288) );
  XNOR U19663 ( .A(n17290), .B(n17291), .Z(n238) );
  AND U19664 ( .A(n17292), .B(n17293), .Z(n17290) );
  XOR U19665 ( .A(n17291), .B(n17206), .Z(n17293) );
  XNOR U19666 ( .A(n17294), .B(n17295), .Z(n17206) );
  ANDN U19667 ( .B(n17296), .A(n17297), .Z(n17294) );
  XOR U19668 ( .A(n17295), .B(n17298), .Z(n17296) );
  XNOR U19669 ( .A(n17291), .B(n17208), .Z(n17292) );
  XOR U19670 ( .A(n17299), .B(n17300), .Z(n17208) );
  AND U19671 ( .A(n242), .B(n17301), .Z(n17299) );
  XOR U19672 ( .A(n17302), .B(n17300), .Z(n17301) );
  XNOR U19673 ( .A(n17303), .B(n17304), .Z(n17291) );
  AND U19674 ( .A(n17305), .B(n17306), .Z(n17303) );
  XNOR U19675 ( .A(n17304), .B(n17233), .Z(n17306) );
  XOR U19676 ( .A(n17297), .B(n17298), .Z(n17233) );
  XNOR U19677 ( .A(n17307), .B(n17308), .Z(n17298) );
  ANDN U19678 ( .B(n17309), .A(n17310), .Z(n17307) );
  XOR U19679 ( .A(n17311), .B(n17312), .Z(n17309) );
  XOR U19680 ( .A(n17313), .B(n17314), .Z(n17297) );
  XNOR U19681 ( .A(n17315), .B(n17316), .Z(n17314) );
  ANDN U19682 ( .B(n17317), .A(n17318), .Z(n17315) );
  XNOR U19683 ( .A(n17319), .B(n17320), .Z(n17317) );
  IV U19684 ( .A(n17295), .Z(n17313) );
  XOR U19685 ( .A(n17321), .B(n17322), .Z(n17295) );
  ANDN U19686 ( .B(n17323), .A(n17324), .Z(n17321) );
  XOR U19687 ( .A(n17322), .B(n17325), .Z(n17323) );
  XOR U19688 ( .A(n17304), .B(n17235), .Z(n17305) );
  XOR U19689 ( .A(n17326), .B(n17327), .Z(n17235) );
  AND U19690 ( .A(n242), .B(n17328), .Z(n17326) );
  XOR U19691 ( .A(n17329), .B(n17327), .Z(n17328) );
  XNOR U19692 ( .A(n17330), .B(n17331), .Z(n17304) );
  NAND U19693 ( .A(n17332), .B(n17333), .Z(n17331) );
  XOR U19694 ( .A(n17334), .B(n17283), .Z(n17333) );
  XOR U19695 ( .A(n17324), .B(n17325), .Z(n17283) );
  XOR U19696 ( .A(n17335), .B(n17312), .Z(n17325) );
  XOR U19697 ( .A(n17336), .B(n17337), .Z(n17312) );
  ANDN U19698 ( .B(n17338), .A(n17339), .Z(n17336) );
  XOR U19699 ( .A(n17337), .B(n17340), .Z(n17338) );
  IV U19700 ( .A(n17310), .Z(n17335) );
  XOR U19701 ( .A(n17308), .B(n17341), .Z(n17310) );
  XOR U19702 ( .A(n17342), .B(n17343), .Z(n17341) );
  ANDN U19703 ( .B(n17344), .A(n17345), .Z(n17342) );
  XOR U19704 ( .A(n17346), .B(n17343), .Z(n17344) );
  IV U19705 ( .A(n17311), .Z(n17308) );
  XOR U19706 ( .A(n17347), .B(n17348), .Z(n17311) );
  ANDN U19707 ( .B(n17349), .A(n17350), .Z(n17347) );
  XOR U19708 ( .A(n17348), .B(n17351), .Z(n17349) );
  XOR U19709 ( .A(n17352), .B(n17353), .Z(n17324) );
  XNOR U19710 ( .A(n17319), .B(n17354), .Z(n17353) );
  IV U19711 ( .A(n17322), .Z(n17354) );
  XOR U19712 ( .A(n17355), .B(n17356), .Z(n17322) );
  ANDN U19713 ( .B(n17357), .A(n17358), .Z(n17355) );
  XOR U19714 ( .A(n17356), .B(n17359), .Z(n17357) );
  XNOR U19715 ( .A(n17360), .B(n17361), .Z(n17319) );
  ANDN U19716 ( .B(n17362), .A(n17363), .Z(n17360) );
  XOR U19717 ( .A(n17361), .B(n17364), .Z(n17362) );
  IV U19718 ( .A(n17318), .Z(n17352) );
  XOR U19719 ( .A(n17316), .B(n17365), .Z(n17318) );
  XOR U19720 ( .A(n17366), .B(n17367), .Z(n17365) );
  ANDN U19721 ( .B(n17368), .A(n17369), .Z(n17366) );
  XOR U19722 ( .A(n17370), .B(n17367), .Z(n17368) );
  IV U19723 ( .A(n17320), .Z(n17316) );
  XOR U19724 ( .A(n17371), .B(n17372), .Z(n17320) );
  ANDN U19725 ( .B(n17373), .A(n17374), .Z(n17371) );
  XOR U19726 ( .A(n17375), .B(n17372), .Z(n17373) );
  IV U19727 ( .A(n17330), .Z(n17334) );
  XOR U19728 ( .A(n17330), .B(n17285), .Z(n17332) );
  XOR U19729 ( .A(n17376), .B(n17377), .Z(n17285) );
  AND U19730 ( .A(n242), .B(n17378), .Z(n17376) );
  XOR U19731 ( .A(n17379), .B(n17377), .Z(n17378) );
  NANDN U19732 ( .A(n17287), .B(n17289), .Z(n17330) );
  XOR U19733 ( .A(n17380), .B(n17381), .Z(n17289) );
  AND U19734 ( .A(n242), .B(n17382), .Z(n17380) );
  XOR U19735 ( .A(n17381), .B(n17383), .Z(n17382) );
  XNOR U19736 ( .A(n17384), .B(n17385), .Z(n242) );
  AND U19737 ( .A(n17386), .B(n17387), .Z(n17384) );
  XOR U19738 ( .A(n17385), .B(n17300), .Z(n17387) );
  XNOR U19739 ( .A(n17388), .B(n17389), .Z(n17300) );
  ANDN U19740 ( .B(n17390), .A(n17391), .Z(n17388) );
  XOR U19741 ( .A(n17389), .B(n17392), .Z(n17390) );
  XNOR U19742 ( .A(n17385), .B(n17302), .Z(n17386) );
  XOR U19743 ( .A(n17393), .B(n17394), .Z(n17302) );
  AND U19744 ( .A(n246), .B(n17395), .Z(n17393) );
  XOR U19745 ( .A(n17396), .B(n17394), .Z(n17395) );
  XNOR U19746 ( .A(n17397), .B(n17398), .Z(n17385) );
  AND U19747 ( .A(n17399), .B(n17400), .Z(n17397) );
  XNOR U19748 ( .A(n17398), .B(n17327), .Z(n17400) );
  XOR U19749 ( .A(n17391), .B(n17392), .Z(n17327) );
  XNOR U19750 ( .A(n17401), .B(n17402), .Z(n17392) );
  ANDN U19751 ( .B(n17403), .A(n17404), .Z(n17401) );
  XOR U19752 ( .A(n17405), .B(n17406), .Z(n17403) );
  XOR U19753 ( .A(n17407), .B(n17408), .Z(n17391) );
  XNOR U19754 ( .A(n17409), .B(n17410), .Z(n17408) );
  ANDN U19755 ( .B(n17411), .A(n17412), .Z(n17409) );
  XNOR U19756 ( .A(n17413), .B(n17414), .Z(n17411) );
  IV U19757 ( .A(n17389), .Z(n17407) );
  XOR U19758 ( .A(n17415), .B(n17416), .Z(n17389) );
  ANDN U19759 ( .B(n17417), .A(n17418), .Z(n17415) );
  XOR U19760 ( .A(n17416), .B(n17419), .Z(n17417) );
  XOR U19761 ( .A(n17398), .B(n17329), .Z(n17399) );
  XOR U19762 ( .A(n17420), .B(n17421), .Z(n17329) );
  AND U19763 ( .A(n246), .B(n17422), .Z(n17420) );
  XOR U19764 ( .A(n17423), .B(n17421), .Z(n17422) );
  XNOR U19765 ( .A(n17424), .B(n17425), .Z(n17398) );
  NAND U19766 ( .A(n17426), .B(n17427), .Z(n17425) );
  XOR U19767 ( .A(n17428), .B(n17377), .Z(n17427) );
  XOR U19768 ( .A(n17418), .B(n17419), .Z(n17377) );
  XOR U19769 ( .A(n17429), .B(n17406), .Z(n17419) );
  XOR U19770 ( .A(n17430), .B(n17431), .Z(n17406) );
  ANDN U19771 ( .B(n17432), .A(n17433), .Z(n17430) );
  XOR U19772 ( .A(n17431), .B(n17434), .Z(n17432) );
  IV U19773 ( .A(n17404), .Z(n17429) );
  XOR U19774 ( .A(n17402), .B(n17435), .Z(n17404) );
  XOR U19775 ( .A(n17436), .B(n17437), .Z(n17435) );
  ANDN U19776 ( .B(n17438), .A(n17439), .Z(n17436) );
  XOR U19777 ( .A(n17440), .B(n17437), .Z(n17438) );
  IV U19778 ( .A(n17405), .Z(n17402) );
  XOR U19779 ( .A(n17441), .B(n17442), .Z(n17405) );
  ANDN U19780 ( .B(n17443), .A(n17444), .Z(n17441) );
  XOR U19781 ( .A(n17442), .B(n17445), .Z(n17443) );
  XOR U19782 ( .A(n17446), .B(n17447), .Z(n17418) );
  XNOR U19783 ( .A(n17413), .B(n17448), .Z(n17447) );
  IV U19784 ( .A(n17416), .Z(n17448) );
  XOR U19785 ( .A(n17449), .B(n17450), .Z(n17416) );
  ANDN U19786 ( .B(n17451), .A(n17452), .Z(n17449) );
  XOR U19787 ( .A(n17450), .B(n17453), .Z(n17451) );
  XNOR U19788 ( .A(n17454), .B(n17455), .Z(n17413) );
  ANDN U19789 ( .B(n17456), .A(n17457), .Z(n17454) );
  XOR U19790 ( .A(n17455), .B(n17458), .Z(n17456) );
  IV U19791 ( .A(n17412), .Z(n17446) );
  XOR U19792 ( .A(n17410), .B(n17459), .Z(n17412) );
  XOR U19793 ( .A(n17460), .B(n17461), .Z(n17459) );
  ANDN U19794 ( .B(n17462), .A(n17463), .Z(n17460) );
  XOR U19795 ( .A(n17464), .B(n17461), .Z(n17462) );
  IV U19796 ( .A(n17414), .Z(n17410) );
  XOR U19797 ( .A(n17465), .B(n17466), .Z(n17414) );
  ANDN U19798 ( .B(n17467), .A(n17468), .Z(n17465) );
  XOR U19799 ( .A(n17469), .B(n17466), .Z(n17467) );
  IV U19800 ( .A(n17424), .Z(n17428) );
  XOR U19801 ( .A(n17424), .B(n17379), .Z(n17426) );
  XOR U19802 ( .A(n17470), .B(n17471), .Z(n17379) );
  AND U19803 ( .A(n246), .B(n17472), .Z(n17470) );
  XOR U19804 ( .A(n17473), .B(n17471), .Z(n17472) );
  NANDN U19805 ( .A(n17381), .B(n17383), .Z(n17424) );
  XOR U19806 ( .A(n17474), .B(n17475), .Z(n17383) );
  AND U19807 ( .A(n246), .B(n17476), .Z(n17474) );
  XOR U19808 ( .A(n17475), .B(n17477), .Z(n17476) );
  XNOR U19809 ( .A(n17478), .B(n17479), .Z(n246) );
  AND U19810 ( .A(n17480), .B(n17481), .Z(n17478) );
  XOR U19811 ( .A(n17479), .B(n17394), .Z(n17481) );
  XNOR U19812 ( .A(n17482), .B(n17483), .Z(n17394) );
  ANDN U19813 ( .B(n17484), .A(n17485), .Z(n17482) );
  XOR U19814 ( .A(n17483), .B(n17486), .Z(n17484) );
  XNOR U19815 ( .A(n17479), .B(n17396), .Z(n17480) );
  XOR U19816 ( .A(n17487), .B(n17488), .Z(n17396) );
  AND U19817 ( .A(n250), .B(n17489), .Z(n17487) );
  XOR U19818 ( .A(n17490), .B(n17488), .Z(n17489) );
  XNOR U19819 ( .A(n17491), .B(n17492), .Z(n17479) );
  AND U19820 ( .A(n17493), .B(n17494), .Z(n17491) );
  XNOR U19821 ( .A(n17492), .B(n17421), .Z(n17494) );
  XOR U19822 ( .A(n17485), .B(n17486), .Z(n17421) );
  XNOR U19823 ( .A(n17495), .B(n17496), .Z(n17486) );
  ANDN U19824 ( .B(n17497), .A(n17498), .Z(n17495) );
  XOR U19825 ( .A(n17499), .B(n17500), .Z(n17497) );
  XOR U19826 ( .A(n17501), .B(n17502), .Z(n17485) );
  XNOR U19827 ( .A(n17503), .B(n17504), .Z(n17502) );
  ANDN U19828 ( .B(n17505), .A(n17506), .Z(n17503) );
  XNOR U19829 ( .A(n17507), .B(n17508), .Z(n17505) );
  IV U19830 ( .A(n17483), .Z(n17501) );
  XOR U19831 ( .A(n17509), .B(n17510), .Z(n17483) );
  ANDN U19832 ( .B(n17511), .A(n17512), .Z(n17509) );
  XOR U19833 ( .A(n17510), .B(n17513), .Z(n17511) );
  XOR U19834 ( .A(n17492), .B(n17423), .Z(n17493) );
  XOR U19835 ( .A(n17514), .B(n17515), .Z(n17423) );
  AND U19836 ( .A(n250), .B(n17516), .Z(n17514) );
  XOR U19837 ( .A(n17517), .B(n17515), .Z(n17516) );
  XNOR U19838 ( .A(n17518), .B(n17519), .Z(n17492) );
  NAND U19839 ( .A(n17520), .B(n17521), .Z(n17519) );
  XOR U19840 ( .A(n17522), .B(n17471), .Z(n17521) );
  XOR U19841 ( .A(n17512), .B(n17513), .Z(n17471) );
  XOR U19842 ( .A(n17523), .B(n17500), .Z(n17513) );
  XOR U19843 ( .A(n17524), .B(n17525), .Z(n17500) );
  ANDN U19844 ( .B(n17526), .A(n17527), .Z(n17524) );
  XOR U19845 ( .A(n17525), .B(n17528), .Z(n17526) );
  IV U19846 ( .A(n17498), .Z(n17523) );
  XOR U19847 ( .A(n17496), .B(n17529), .Z(n17498) );
  XOR U19848 ( .A(n17530), .B(n17531), .Z(n17529) );
  ANDN U19849 ( .B(n17532), .A(n17533), .Z(n17530) );
  XOR U19850 ( .A(n17534), .B(n17531), .Z(n17532) );
  IV U19851 ( .A(n17499), .Z(n17496) );
  XOR U19852 ( .A(n17535), .B(n17536), .Z(n17499) );
  ANDN U19853 ( .B(n17537), .A(n17538), .Z(n17535) );
  XOR U19854 ( .A(n17536), .B(n17539), .Z(n17537) );
  XOR U19855 ( .A(n17540), .B(n17541), .Z(n17512) );
  XNOR U19856 ( .A(n17507), .B(n17542), .Z(n17541) );
  IV U19857 ( .A(n17510), .Z(n17542) );
  XOR U19858 ( .A(n17543), .B(n17544), .Z(n17510) );
  ANDN U19859 ( .B(n17545), .A(n17546), .Z(n17543) );
  XOR U19860 ( .A(n17544), .B(n17547), .Z(n17545) );
  XNOR U19861 ( .A(n17548), .B(n17549), .Z(n17507) );
  ANDN U19862 ( .B(n17550), .A(n17551), .Z(n17548) );
  XOR U19863 ( .A(n17549), .B(n17552), .Z(n17550) );
  IV U19864 ( .A(n17506), .Z(n17540) );
  XOR U19865 ( .A(n17504), .B(n17553), .Z(n17506) );
  XOR U19866 ( .A(n17554), .B(n17555), .Z(n17553) );
  ANDN U19867 ( .B(n17556), .A(n17557), .Z(n17554) );
  XOR U19868 ( .A(n17558), .B(n17555), .Z(n17556) );
  IV U19869 ( .A(n17508), .Z(n17504) );
  XOR U19870 ( .A(n17559), .B(n17560), .Z(n17508) );
  ANDN U19871 ( .B(n17561), .A(n17562), .Z(n17559) );
  XOR U19872 ( .A(n17563), .B(n17560), .Z(n17561) );
  IV U19873 ( .A(n17518), .Z(n17522) );
  XOR U19874 ( .A(n17518), .B(n17473), .Z(n17520) );
  XOR U19875 ( .A(n17564), .B(n17565), .Z(n17473) );
  AND U19876 ( .A(n250), .B(n17566), .Z(n17564) );
  XOR U19877 ( .A(n17567), .B(n17565), .Z(n17566) );
  NANDN U19878 ( .A(n17475), .B(n17477), .Z(n17518) );
  XOR U19879 ( .A(n17568), .B(n17569), .Z(n17477) );
  AND U19880 ( .A(n250), .B(n17570), .Z(n17568) );
  XOR U19881 ( .A(n17569), .B(n17571), .Z(n17570) );
  XNOR U19882 ( .A(n17572), .B(n17573), .Z(n250) );
  AND U19883 ( .A(n17574), .B(n17575), .Z(n17572) );
  XOR U19884 ( .A(n17573), .B(n17488), .Z(n17575) );
  XNOR U19885 ( .A(n17576), .B(n17577), .Z(n17488) );
  ANDN U19886 ( .B(n17578), .A(n17579), .Z(n17576) );
  XOR U19887 ( .A(n17577), .B(n17580), .Z(n17578) );
  XNOR U19888 ( .A(n17573), .B(n17490), .Z(n17574) );
  XOR U19889 ( .A(n17581), .B(n17582), .Z(n17490) );
  AND U19890 ( .A(n254), .B(n17583), .Z(n17581) );
  XOR U19891 ( .A(n17584), .B(n17582), .Z(n17583) );
  XNOR U19892 ( .A(n17585), .B(n17586), .Z(n17573) );
  AND U19893 ( .A(n17587), .B(n17588), .Z(n17585) );
  XNOR U19894 ( .A(n17586), .B(n17515), .Z(n17588) );
  XOR U19895 ( .A(n17579), .B(n17580), .Z(n17515) );
  XNOR U19896 ( .A(n17589), .B(n17590), .Z(n17580) );
  ANDN U19897 ( .B(n17591), .A(n17592), .Z(n17589) );
  XOR U19898 ( .A(n17593), .B(n17594), .Z(n17591) );
  XOR U19899 ( .A(n17595), .B(n17596), .Z(n17579) );
  XNOR U19900 ( .A(n17597), .B(n17598), .Z(n17596) );
  ANDN U19901 ( .B(n17599), .A(n17600), .Z(n17597) );
  XNOR U19902 ( .A(n17601), .B(n17602), .Z(n17599) );
  IV U19903 ( .A(n17577), .Z(n17595) );
  XOR U19904 ( .A(n17603), .B(n17604), .Z(n17577) );
  ANDN U19905 ( .B(n17605), .A(n17606), .Z(n17603) );
  XOR U19906 ( .A(n17604), .B(n17607), .Z(n17605) );
  XOR U19907 ( .A(n17586), .B(n17517), .Z(n17587) );
  XOR U19908 ( .A(n17608), .B(n17609), .Z(n17517) );
  AND U19909 ( .A(n254), .B(n17610), .Z(n17608) );
  XOR U19910 ( .A(n17611), .B(n17609), .Z(n17610) );
  XNOR U19911 ( .A(n17612), .B(n17613), .Z(n17586) );
  NAND U19912 ( .A(n17614), .B(n17615), .Z(n17613) );
  XOR U19913 ( .A(n17616), .B(n17565), .Z(n17615) );
  XOR U19914 ( .A(n17606), .B(n17607), .Z(n17565) );
  XOR U19915 ( .A(n17617), .B(n17594), .Z(n17607) );
  XOR U19916 ( .A(n17618), .B(n17619), .Z(n17594) );
  ANDN U19917 ( .B(n17620), .A(n17621), .Z(n17618) );
  XOR U19918 ( .A(n17619), .B(n17622), .Z(n17620) );
  IV U19919 ( .A(n17592), .Z(n17617) );
  XOR U19920 ( .A(n17590), .B(n17623), .Z(n17592) );
  XOR U19921 ( .A(n17624), .B(n17625), .Z(n17623) );
  ANDN U19922 ( .B(n17626), .A(n17627), .Z(n17624) );
  XOR U19923 ( .A(n17628), .B(n17625), .Z(n17626) );
  IV U19924 ( .A(n17593), .Z(n17590) );
  XOR U19925 ( .A(n17629), .B(n17630), .Z(n17593) );
  ANDN U19926 ( .B(n17631), .A(n17632), .Z(n17629) );
  XOR U19927 ( .A(n17630), .B(n17633), .Z(n17631) );
  XOR U19928 ( .A(n17634), .B(n17635), .Z(n17606) );
  XNOR U19929 ( .A(n17601), .B(n17636), .Z(n17635) );
  IV U19930 ( .A(n17604), .Z(n17636) );
  XOR U19931 ( .A(n17637), .B(n17638), .Z(n17604) );
  ANDN U19932 ( .B(n17639), .A(n17640), .Z(n17637) );
  XOR U19933 ( .A(n17638), .B(n17641), .Z(n17639) );
  XNOR U19934 ( .A(n17642), .B(n17643), .Z(n17601) );
  ANDN U19935 ( .B(n17644), .A(n17645), .Z(n17642) );
  XOR U19936 ( .A(n17643), .B(n17646), .Z(n17644) );
  IV U19937 ( .A(n17600), .Z(n17634) );
  XOR U19938 ( .A(n17598), .B(n17647), .Z(n17600) );
  XOR U19939 ( .A(n17648), .B(n17649), .Z(n17647) );
  ANDN U19940 ( .B(n17650), .A(n17651), .Z(n17648) );
  XOR U19941 ( .A(n17652), .B(n17649), .Z(n17650) );
  IV U19942 ( .A(n17602), .Z(n17598) );
  XOR U19943 ( .A(n17653), .B(n17654), .Z(n17602) );
  ANDN U19944 ( .B(n17655), .A(n17656), .Z(n17653) );
  XOR U19945 ( .A(n17657), .B(n17654), .Z(n17655) );
  IV U19946 ( .A(n17612), .Z(n17616) );
  XOR U19947 ( .A(n17612), .B(n17567), .Z(n17614) );
  XOR U19948 ( .A(n17658), .B(n17659), .Z(n17567) );
  AND U19949 ( .A(n254), .B(n17660), .Z(n17658) );
  XOR U19950 ( .A(n17661), .B(n17659), .Z(n17660) );
  NANDN U19951 ( .A(n17569), .B(n17571), .Z(n17612) );
  XOR U19952 ( .A(n17662), .B(n17663), .Z(n17571) );
  AND U19953 ( .A(n254), .B(n17664), .Z(n17662) );
  XOR U19954 ( .A(n17663), .B(n17665), .Z(n17664) );
  XNOR U19955 ( .A(n17666), .B(n17667), .Z(n254) );
  AND U19956 ( .A(n17668), .B(n17669), .Z(n17666) );
  XOR U19957 ( .A(n17667), .B(n17582), .Z(n17669) );
  XNOR U19958 ( .A(n17670), .B(n17671), .Z(n17582) );
  ANDN U19959 ( .B(n17672), .A(n17673), .Z(n17670) );
  XOR U19960 ( .A(n17671), .B(n17674), .Z(n17672) );
  XNOR U19961 ( .A(n17667), .B(n17584), .Z(n17668) );
  XOR U19962 ( .A(n17675), .B(n17676), .Z(n17584) );
  AND U19963 ( .A(n258), .B(n17677), .Z(n17675) );
  XOR U19964 ( .A(n17678), .B(n17676), .Z(n17677) );
  XNOR U19965 ( .A(n17679), .B(n17680), .Z(n17667) );
  AND U19966 ( .A(n17681), .B(n17682), .Z(n17679) );
  XNOR U19967 ( .A(n17680), .B(n17609), .Z(n17682) );
  XOR U19968 ( .A(n17673), .B(n17674), .Z(n17609) );
  XNOR U19969 ( .A(n17683), .B(n17684), .Z(n17674) );
  ANDN U19970 ( .B(n17685), .A(n17686), .Z(n17683) );
  XOR U19971 ( .A(n17687), .B(n17688), .Z(n17685) );
  XOR U19972 ( .A(n17689), .B(n17690), .Z(n17673) );
  XNOR U19973 ( .A(n17691), .B(n17692), .Z(n17690) );
  ANDN U19974 ( .B(n17693), .A(n17694), .Z(n17691) );
  XNOR U19975 ( .A(n17695), .B(n17696), .Z(n17693) );
  IV U19976 ( .A(n17671), .Z(n17689) );
  XOR U19977 ( .A(n17697), .B(n17698), .Z(n17671) );
  ANDN U19978 ( .B(n17699), .A(n17700), .Z(n17697) );
  XOR U19979 ( .A(n17698), .B(n17701), .Z(n17699) );
  XOR U19980 ( .A(n17680), .B(n17611), .Z(n17681) );
  XOR U19981 ( .A(n17702), .B(n17703), .Z(n17611) );
  AND U19982 ( .A(n258), .B(n17704), .Z(n17702) );
  XOR U19983 ( .A(n17705), .B(n17703), .Z(n17704) );
  XNOR U19984 ( .A(n17706), .B(n17707), .Z(n17680) );
  NAND U19985 ( .A(n17708), .B(n17709), .Z(n17707) );
  XOR U19986 ( .A(n17710), .B(n17659), .Z(n17709) );
  XOR U19987 ( .A(n17700), .B(n17701), .Z(n17659) );
  XOR U19988 ( .A(n17711), .B(n17688), .Z(n17701) );
  XOR U19989 ( .A(n17712), .B(n17713), .Z(n17688) );
  ANDN U19990 ( .B(n17714), .A(n17715), .Z(n17712) );
  XOR U19991 ( .A(n17713), .B(n17716), .Z(n17714) );
  IV U19992 ( .A(n17686), .Z(n17711) );
  XOR U19993 ( .A(n17684), .B(n17717), .Z(n17686) );
  XOR U19994 ( .A(n17718), .B(n17719), .Z(n17717) );
  ANDN U19995 ( .B(n17720), .A(n17721), .Z(n17718) );
  XOR U19996 ( .A(n17722), .B(n17719), .Z(n17720) );
  IV U19997 ( .A(n17687), .Z(n17684) );
  XOR U19998 ( .A(n17723), .B(n17724), .Z(n17687) );
  ANDN U19999 ( .B(n17725), .A(n17726), .Z(n17723) );
  XOR U20000 ( .A(n17724), .B(n17727), .Z(n17725) );
  XOR U20001 ( .A(n17728), .B(n17729), .Z(n17700) );
  XNOR U20002 ( .A(n17695), .B(n17730), .Z(n17729) );
  IV U20003 ( .A(n17698), .Z(n17730) );
  XOR U20004 ( .A(n17731), .B(n17732), .Z(n17698) );
  ANDN U20005 ( .B(n17733), .A(n17734), .Z(n17731) );
  XOR U20006 ( .A(n17732), .B(n17735), .Z(n17733) );
  XNOR U20007 ( .A(n17736), .B(n17737), .Z(n17695) );
  ANDN U20008 ( .B(n17738), .A(n17739), .Z(n17736) );
  XOR U20009 ( .A(n17737), .B(n17740), .Z(n17738) );
  IV U20010 ( .A(n17694), .Z(n17728) );
  XOR U20011 ( .A(n17692), .B(n17741), .Z(n17694) );
  XOR U20012 ( .A(n17742), .B(n17743), .Z(n17741) );
  ANDN U20013 ( .B(n17744), .A(n17745), .Z(n17742) );
  XOR U20014 ( .A(n17746), .B(n17743), .Z(n17744) );
  IV U20015 ( .A(n17696), .Z(n17692) );
  XOR U20016 ( .A(n17747), .B(n17748), .Z(n17696) );
  ANDN U20017 ( .B(n17749), .A(n17750), .Z(n17747) );
  XOR U20018 ( .A(n17751), .B(n17748), .Z(n17749) );
  IV U20019 ( .A(n17706), .Z(n17710) );
  XOR U20020 ( .A(n17706), .B(n17661), .Z(n17708) );
  XOR U20021 ( .A(n17752), .B(n17753), .Z(n17661) );
  AND U20022 ( .A(n258), .B(n17754), .Z(n17752) );
  XOR U20023 ( .A(n17755), .B(n17753), .Z(n17754) );
  NANDN U20024 ( .A(n17663), .B(n17665), .Z(n17706) );
  XOR U20025 ( .A(n17756), .B(n17757), .Z(n17665) );
  AND U20026 ( .A(n258), .B(n17758), .Z(n17756) );
  XOR U20027 ( .A(n17757), .B(n17759), .Z(n17758) );
  XNOR U20028 ( .A(n17760), .B(n17761), .Z(n258) );
  AND U20029 ( .A(n17762), .B(n17763), .Z(n17760) );
  XOR U20030 ( .A(n17761), .B(n17676), .Z(n17763) );
  XNOR U20031 ( .A(n17764), .B(n17765), .Z(n17676) );
  ANDN U20032 ( .B(n17766), .A(n17767), .Z(n17764) );
  XOR U20033 ( .A(n17765), .B(n17768), .Z(n17766) );
  XNOR U20034 ( .A(n17761), .B(n17678), .Z(n17762) );
  XOR U20035 ( .A(n17769), .B(n17770), .Z(n17678) );
  AND U20036 ( .A(n262), .B(n17771), .Z(n17769) );
  XOR U20037 ( .A(n17772), .B(n17770), .Z(n17771) );
  XNOR U20038 ( .A(n17773), .B(n17774), .Z(n17761) );
  AND U20039 ( .A(n17775), .B(n17776), .Z(n17773) );
  XNOR U20040 ( .A(n17774), .B(n17703), .Z(n17776) );
  XOR U20041 ( .A(n17767), .B(n17768), .Z(n17703) );
  XNOR U20042 ( .A(n17777), .B(n17778), .Z(n17768) );
  ANDN U20043 ( .B(n17779), .A(n17780), .Z(n17777) );
  XOR U20044 ( .A(n17781), .B(n17782), .Z(n17779) );
  XOR U20045 ( .A(n17783), .B(n17784), .Z(n17767) );
  XNOR U20046 ( .A(n17785), .B(n17786), .Z(n17784) );
  ANDN U20047 ( .B(n17787), .A(n17788), .Z(n17785) );
  XNOR U20048 ( .A(n17789), .B(n17790), .Z(n17787) );
  IV U20049 ( .A(n17765), .Z(n17783) );
  XOR U20050 ( .A(n17791), .B(n17792), .Z(n17765) );
  ANDN U20051 ( .B(n17793), .A(n17794), .Z(n17791) );
  XOR U20052 ( .A(n17792), .B(n17795), .Z(n17793) );
  XOR U20053 ( .A(n17774), .B(n17705), .Z(n17775) );
  XOR U20054 ( .A(n17796), .B(n17797), .Z(n17705) );
  AND U20055 ( .A(n262), .B(n17798), .Z(n17796) );
  XOR U20056 ( .A(n17799), .B(n17797), .Z(n17798) );
  XNOR U20057 ( .A(n17800), .B(n17801), .Z(n17774) );
  NAND U20058 ( .A(n17802), .B(n17803), .Z(n17801) );
  XOR U20059 ( .A(n17804), .B(n17753), .Z(n17803) );
  XOR U20060 ( .A(n17794), .B(n17795), .Z(n17753) );
  XOR U20061 ( .A(n17805), .B(n17782), .Z(n17795) );
  XOR U20062 ( .A(n17806), .B(n17807), .Z(n17782) );
  ANDN U20063 ( .B(n17808), .A(n17809), .Z(n17806) );
  XOR U20064 ( .A(n17807), .B(n17810), .Z(n17808) );
  IV U20065 ( .A(n17780), .Z(n17805) );
  XOR U20066 ( .A(n17778), .B(n17811), .Z(n17780) );
  XOR U20067 ( .A(n17812), .B(n17813), .Z(n17811) );
  ANDN U20068 ( .B(n17814), .A(n17815), .Z(n17812) );
  XOR U20069 ( .A(n17816), .B(n17813), .Z(n17814) );
  IV U20070 ( .A(n17781), .Z(n17778) );
  XOR U20071 ( .A(n17817), .B(n17818), .Z(n17781) );
  ANDN U20072 ( .B(n17819), .A(n17820), .Z(n17817) );
  XOR U20073 ( .A(n17818), .B(n17821), .Z(n17819) );
  XOR U20074 ( .A(n17822), .B(n17823), .Z(n17794) );
  XNOR U20075 ( .A(n17789), .B(n17824), .Z(n17823) );
  IV U20076 ( .A(n17792), .Z(n17824) );
  XOR U20077 ( .A(n17825), .B(n17826), .Z(n17792) );
  ANDN U20078 ( .B(n17827), .A(n17828), .Z(n17825) );
  XOR U20079 ( .A(n17826), .B(n17829), .Z(n17827) );
  XNOR U20080 ( .A(n17830), .B(n17831), .Z(n17789) );
  ANDN U20081 ( .B(n17832), .A(n17833), .Z(n17830) );
  XOR U20082 ( .A(n17831), .B(n17834), .Z(n17832) );
  IV U20083 ( .A(n17788), .Z(n17822) );
  XOR U20084 ( .A(n17786), .B(n17835), .Z(n17788) );
  XOR U20085 ( .A(n17836), .B(n17837), .Z(n17835) );
  ANDN U20086 ( .B(n17838), .A(n17839), .Z(n17836) );
  XOR U20087 ( .A(n17840), .B(n17837), .Z(n17838) );
  IV U20088 ( .A(n17790), .Z(n17786) );
  XOR U20089 ( .A(n17841), .B(n17842), .Z(n17790) );
  ANDN U20090 ( .B(n17843), .A(n17844), .Z(n17841) );
  XOR U20091 ( .A(n17845), .B(n17842), .Z(n17843) );
  IV U20092 ( .A(n17800), .Z(n17804) );
  XOR U20093 ( .A(n17800), .B(n17755), .Z(n17802) );
  XOR U20094 ( .A(n17846), .B(n17847), .Z(n17755) );
  AND U20095 ( .A(n262), .B(n17848), .Z(n17846) );
  XOR U20096 ( .A(n17849), .B(n17847), .Z(n17848) );
  NANDN U20097 ( .A(n17757), .B(n17759), .Z(n17800) );
  XOR U20098 ( .A(n17850), .B(n17851), .Z(n17759) );
  AND U20099 ( .A(n262), .B(n17852), .Z(n17850) );
  XOR U20100 ( .A(n17851), .B(n17853), .Z(n17852) );
  XNOR U20101 ( .A(n17854), .B(n17855), .Z(n262) );
  AND U20102 ( .A(n17856), .B(n17857), .Z(n17854) );
  XOR U20103 ( .A(n17855), .B(n17770), .Z(n17857) );
  XNOR U20104 ( .A(n17858), .B(n17859), .Z(n17770) );
  ANDN U20105 ( .B(n17860), .A(n17861), .Z(n17858) );
  XOR U20106 ( .A(n17859), .B(n17862), .Z(n17860) );
  XNOR U20107 ( .A(n17855), .B(n17772), .Z(n17856) );
  XOR U20108 ( .A(n17863), .B(n17864), .Z(n17772) );
  AND U20109 ( .A(n266), .B(n17865), .Z(n17863) );
  XOR U20110 ( .A(n17866), .B(n17864), .Z(n17865) );
  XNOR U20111 ( .A(n17867), .B(n17868), .Z(n17855) );
  AND U20112 ( .A(n17869), .B(n17870), .Z(n17867) );
  XNOR U20113 ( .A(n17868), .B(n17797), .Z(n17870) );
  XOR U20114 ( .A(n17861), .B(n17862), .Z(n17797) );
  XNOR U20115 ( .A(n17871), .B(n17872), .Z(n17862) );
  ANDN U20116 ( .B(n17873), .A(n17874), .Z(n17871) );
  XOR U20117 ( .A(n17875), .B(n17876), .Z(n17873) );
  XOR U20118 ( .A(n17877), .B(n17878), .Z(n17861) );
  XNOR U20119 ( .A(n17879), .B(n17880), .Z(n17878) );
  ANDN U20120 ( .B(n17881), .A(n17882), .Z(n17879) );
  XNOR U20121 ( .A(n17883), .B(n17884), .Z(n17881) );
  IV U20122 ( .A(n17859), .Z(n17877) );
  XOR U20123 ( .A(n17885), .B(n17886), .Z(n17859) );
  ANDN U20124 ( .B(n17887), .A(n17888), .Z(n17885) );
  XOR U20125 ( .A(n17886), .B(n17889), .Z(n17887) );
  XOR U20126 ( .A(n17868), .B(n17799), .Z(n17869) );
  XOR U20127 ( .A(n17890), .B(n17891), .Z(n17799) );
  AND U20128 ( .A(n266), .B(n17892), .Z(n17890) );
  XOR U20129 ( .A(n17893), .B(n17891), .Z(n17892) );
  XNOR U20130 ( .A(n17894), .B(n17895), .Z(n17868) );
  NAND U20131 ( .A(n17896), .B(n17897), .Z(n17895) );
  XOR U20132 ( .A(n17898), .B(n17847), .Z(n17897) );
  XOR U20133 ( .A(n17888), .B(n17889), .Z(n17847) );
  XOR U20134 ( .A(n17899), .B(n17876), .Z(n17889) );
  XOR U20135 ( .A(n17900), .B(n17901), .Z(n17876) );
  ANDN U20136 ( .B(n17902), .A(n17903), .Z(n17900) );
  XOR U20137 ( .A(n17901), .B(n17904), .Z(n17902) );
  IV U20138 ( .A(n17874), .Z(n17899) );
  XOR U20139 ( .A(n17872), .B(n17905), .Z(n17874) );
  XOR U20140 ( .A(n17906), .B(n17907), .Z(n17905) );
  ANDN U20141 ( .B(n17908), .A(n17909), .Z(n17906) );
  XOR U20142 ( .A(n17910), .B(n17907), .Z(n17908) );
  IV U20143 ( .A(n17875), .Z(n17872) );
  XOR U20144 ( .A(n17911), .B(n17912), .Z(n17875) );
  ANDN U20145 ( .B(n17913), .A(n17914), .Z(n17911) );
  XOR U20146 ( .A(n17912), .B(n17915), .Z(n17913) );
  XOR U20147 ( .A(n17916), .B(n17917), .Z(n17888) );
  XNOR U20148 ( .A(n17883), .B(n17918), .Z(n17917) );
  IV U20149 ( .A(n17886), .Z(n17918) );
  XOR U20150 ( .A(n17919), .B(n17920), .Z(n17886) );
  ANDN U20151 ( .B(n17921), .A(n17922), .Z(n17919) );
  XOR U20152 ( .A(n17920), .B(n17923), .Z(n17921) );
  XNOR U20153 ( .A(n17924), .B(n17925), .Z(n17883) );
  ANDN U20154 ( .B(n17926), .A(n17927), .Z(n17924) );
  XOR U20155 ( .A(n17925), .B(n17928), .Z(n17926) );
  IV U20156 ( .A(n17882), .Z(n17916) );
  XOR U20157 ( .A(n17880), .B(n17929), .Z(n17882) );
  XOR U20158 ( .A(n17930), .B(n17931), .Z(n17929) );
  ANDN U20159 ( .B(n17932), .A(n17933), .Z(n17930) );
  XOR U20160 ( .A(n17934), .B(n17931), .Z(n17932) );
  IV U20161 ( .A(n17884), .Z(n17880) );
  XOR U20162 ( .A(n17935), .B(n17936), .Z(n17884) );
  ANDN U20163 ( .B(n17937), .A(n17938), .Z(n17935) );
  XOR U20164 ( .A(n17939), .B(n17936), .Z(n17937) );
  IV U20165 ( .A(n17894), .Z(n17898) );
  XOR U20166 ( .A(n17894), .B(n17849), .Z(n17896) );
  XOR U20167 ( .A(n17940), .B(n17941), .Z(n17849) );
  AND U20168 ( .A(n266), .B(n17942), .Z(n17940) );
  XOR U20169 ( .A(n17943), .B(n17941), .Z(n17942) );
  NANDN U20170 ( .A(n17851), .B(n17853), .Z(n17894) );
  XOR U20171 ( .A(n17944), .B(n17945), .Z(n17853) );
  AND U20172 ( .A(n266), .B(n17946), .Z(n17944) );
  XOR U20173 ( .A(n17945), .B(n17947), .Z(n17946) );
  XNOR U20174 ( .A(n17948), .B(n17949), .Z(n266) );
  AND U20175 ( .A(n17950), .B(n17951), .Z(n17948) );
  XOR U20176 ( .A(n17949), .B(n17864), .Z(n17951) );
  XNOR U20177 ( .A(n17952), .B(n17953), .Z(n17864) );
  ANDN U20178 ( .B(n17954), .A(n17955), .Z(n17952) );
  XOR U20179 ( .A(n17953), .B(n17956), .Z(n17954) );
  XNOR U20180 ( .A(n17949), .B(n17866), .Z(n17950) );
  XOR U20181 ( .A(n17957), .B(n17958), .Z(n17866) );
  AND U20182 ( .A(n270), .B(n17959), .Z(n17957) );
  XOR U20183 ( .A(n17960), .B(n17958), .Z(n17959) );
  XNOR U20184 ( .A(n17961), .B(n17962), .Z(n17949) );
  AND U20185 ( .A(n17963), .B(n17964), .Z(n17961) );
  XNOR U20186 ( .A(n17962), .B(n17891), .Z(n17964) );
  XOR U20187 ( .A(n17955), .B(n17956), .Z(n17891) );
  XNOR U20188 ( .A(n17965), .B(n17966), .Z(n17956) );
  ANDN U20189 ( .B(n17967), .A(n17968), .Z(n17965) );
  XOR U20190 ( .A(n17969), .B(n17970), .Z(n17967) );
  XOR U20191 ( .A(n17971), .B(n17972), .Z(n17955) );
  XNOR U20192 ( .A(n17973), .B(n17974), .Z(n17972) );
  ANDN U20193 ( .B(n17975), .A(n17976), .Z(n17973) );
  XNOR U20194 ( .A(n17977), .B(n17978), .Z(n17975) );
  IV U20195 ( .A(n17953), .Z(n17971) );
  XOR U20196 ( .A(n17979), .B(n17980), .Z(n17953) );
  ANDN U20197 ( .B(n17981), .A(n17982), .Z(n17979) );
  XOR U20198 ( .A(n17980), .B(n17983), .Z(n17981) );
  XOR U20199 ( .A(n17962), .B(n17893), .Z(n17963) );
  XOR U20200 ( .A(n17984), .B(n17985), .Z(n17893) );
  AND U20201 ( .A(n270), .B(n17986), .Z(n17984) );
  XOR U20202 ( .A(n17987), .B(n17985), .Z(n17986) );
  XNOR U20203 ( .A(n17988), .B(n17989), .Z(n17962) );
  NAND U20204 ( .A(n17990), .B(n17991), .Z(n17989) );
  XOR U20205 ( .A(n17992), .B(n17941), .Z(n17991) );
  XOR U20206 ( .A(n17982), .B(n17983), .Z(n17941) );
  XOR U20207 ( .A(n17993), .B(n17970), .Z(n17983) );
  XOR U20208 ( .A(n17994), .B(n17995), .Z(n17970) );
  ANDN U20209 ( .B(n17996), .A(n17997), .Z(n17994) );
  XOR U20210 ( .A(n17995), .B(n17998), .Z(n17996) );
  IV U20211 ( .A(n17968), .Z(n17993) );
  XOR U20212 ( .A(n17966), .B(n17999), .Z(n17968) );
  XOR U20213 ( .A(n18000), .B(n18001), .Z(n17999) );
  ANDN U20214 ( .B(n18002), .A(n18003), .Z(n18000) );
  XOR U20215 ( .A(n18004), .B(n18001), .Z(n18002) );
  IV U20216 ( .A(n17969), .Z(n17966) );
  XOR U20217 ( .A(n18005), .B(n18006), .Z(n17969) );
  ANDN U20218 ( .B(n18007), .A(n18008), .Z(n18005) );
  XOR U20219 ( .A(n18006), .B(n18009), .Z(n18007) );
  XOR U20220 ( .A(n18010), .B(n18011), .Z(n17982) );
  XNOR U20221 ( .A(n17977), .B(n18012), .Z(n18011) );
  IV U20222 ( .A(n17980), .Z(n18012) );
  XOR U20223 ( .A(n18013), .B(n18014), .Z(n17980) );
  ANDN U20224 ( .B(n18015), .A(n18016), .Z(n18013) );
  XOR U20225 ( .A(n18014), .B(n18017), .Z(n18015) );
  XNOR U20226 ( .A(n18018), .B(n18019), .Z(n17977) );
  ANDN U20227 ( .B(n18020), .A(n18021), .Z(n18018) );
  XOR U20228 ( .A(n18019), .B(n18022), .Z(n18020) );
  IV U20229 ( .A(n17976), .Z(n18010) );
  XOR U20230 ( .A(n17974), .B(n18023), .Z(n17976) );
  XOR U20231 ( .A(n18024), .B(n18025), .Z(n18023) );
  ANDN U20232 ( .B(n18026), .A(n18027), .Z(n18024) );
  XOR U20233 ( .A(n18028), .B(n18025), .Z(n18026) );
  IV U20234 ( .A(n17978), .Z(n17974) );
  XOR U20235 ( .A(n18029), .B(n18030), .Z(n17978) );
  ANDN U20236 ( .B(n18031), .A(n18032), .Z(n18029) );
  XOR U20237 ( .A(n18033), .B(n18030), .Z(n18031) );
  IV U20238 ( .A(n17988), .Z(n17992) );
  XOR U20239 ( .A(n17988), .B(n17943), .Z(n17990) );
  XOR U20240 ( .A(n18034), .B(n18035), .Z(n17943) );
  AND U20241 ( .A(n270), .B(n18036), .Z(n18034) );
  XOR U20242 ( .A(n18037), .B(n18035), .Z(n18036) );
  NANDN U20243 ( .A(n17945), .B(n17947), .Z(n17988) );
  XOR U20244 ( .A(n18038), .B(n18039), .Z(n17947) );
  AND U20245 ( .A(n270), .B(n18040), .Z(n18038) );
  XOR U20246 ( .A(n18039), .B(n18041), .Z(n18040) );
  XNOR U20247 ( .A(n18042), .B(n18043), .Z(n270) );
  AND U20248 ( .A(n18044), .B(n18045), .Z(n18042) );
  XOR U20249 ( .A(n18043), .B(n17958), .Z(n18045) );
  XNOR U20250 ( .A(n18046), .B(n18047), .Z(n17958) );
  ANDN U20251 ( .B(n18048), .A(n18049), .Z(n18046) );
  XOR U20252 ( .A(n18047), .B(n18050), .Z(n18048) );
  XNOR U20253 ( .A(n18043), .B(n17960), .Z(n18044) );
  XOR U20254 ( .A(n18051), .B(n18052), .Z(n17960) );
  AND U20255 ( .A(n274), .B(n18053), .Z(n18051) );
  XOR U20256 ( .A(n18054), .B(n18052), .Z(n18053) );
  XNOR U20257 ( .A(n18055), .B(n18056), .Z(n18043) );
  AND U20258 ( .A(n18057), .B(n18058), .Z(n18055) );
  XNOR U20259 ( .A(n18056), .B(n17985), .Z(n18058) );
  XOR U20260 ( .A(n18049), .B(n18050), .Z(n17985) );
  XNOR U20261 ( .A(n18059), .B(n18060), .Z(n18050) );
  ANDN U20262 ( .B(n18061), .A(n18062), .Z(n18059) );
  XOR U20263 ( .A(n18063), .B(n18064), .Z(n18061) );
  XOR U20264 ( .A(n18065), .B(n18066), .Z(n18049) );
  XNOR U20265 ( .A(n18067), .B(n18068), .Z(n18066) );
  ANDN U20266 ( .B(n18069), .A(n18070), .Z(n18067) );
  XNOR U20267 ( .A(n18071), .B(n18072), .Z(n18069) );
  IV U20268 ( .A(n18047), .Z(n18065) );
  XOR U20269 ( .A(n18073), .B(n18074), .Z(n18047) );
  ANDN U20270 ( .B(n18075), .A(n18076), .Z(n18073) );
  XOR U20271 ( .A(n18074), .B(n18077), .Z(n18075) );
  XOR U20272 ( .A(n18056), .B(n17987), .Z(n18057) );
  XOR U20273 ( .A(n18078), .B(n18079), .Z(n17987) );
  AND U20274 ( .A(n274), .B(n18080), .Z(n18078) );
  XOR U20275 ( .A(n18081), .B(n18079), .Z(n18080) );
  XNOR U20276 ( .A(n18082), .B(n18083), .Z(n18056) );
  NAND U20277 ( .A(n18084), .B(n18085), .Z(n18083) );
  XOR U20278 ( .A(n18086), .B(n18035), .Z(n18085) );
  XOR U20279 ( .A(n18076), .B(n18077), .Z(n18035) );
  XOR U20280 ( .A(n18087), .B(n18064), .Z(n18077) );
  XOR U20281 ( .A(n18088), .B(n18089), .Z(n18064) );
  ANDN U20282 ( .B(n18090), .A(n18091), .Z(n18088) );
  XOR U20283 ( .A(n18089), .B(n18092), .Z(n18090) );
  IV U20284 ( .A(n18062), .Z(n18087) );
  XOR U20285 ( .A(n18060), .B(n18093), .Z(n18062) );
  XOR U20286 ( .A(n18094), .B(n18095), .Z(n18093) );
  ANDN U20287 ( .B(n18096), .A(n18097), .Z(n18094) );
  XOR U20288 ( .A(n18098), .B(n18095), .Z(n18096) );
  IV U20289 ( .A(n18063), .Z(n18060) );
  XOR U20290 ( .A(n18099), .B(n18100), .Z(n18063) );
  ANDN U20291 ( .B(n18101), .A(n18102), .Z(n18099) );
  XOR U20292 ( .A(n18100), .B(n18103), .Z(n18101) );
  XOR U20293 ( .A(n18104), .B(n18105), .Z(n18076) );
  XNOR U20294 ( .A(n18071), .B(n18106), .Z(n18105) );
  IV U20295 ( .A(n18074), .Z(n18106) );
  XOR U20296 ( .A(n18107), .B(n18108), .Z(n18074) );
  ANDN U20297 ( .B(n18109), .A(n18110), .Z(n18107) );
  XOR U20298 ( .A(n18108), .B(n18111), .Z(n18109) );
  XNOR U20299 ( .A(n18112), .B(n18113), .Z(n18071) );
  ANDN U20300 ( .B(n18114), .A(n18115), .Z(n18112) );
  XOR U20301 ( .A(n18113), .B(n18116), .Z(n18114) );
  IV U20302 ( .A(n18070), .Z(n18104) );
  XOR U20303 ( .A(n18068), .B(n18117), .Z(n18070) );
  XOR U20304 ( .A(n18118), .B(n18119), .Z(n18117) );
  ANDN U20305 ( .B(n18120), .A(n18121), .Z(n18118) );
  XOR U20306 ( .A(n18122), .B(n18119), .Z(n18120) );
  IV U20307 ( .A(n18072), .Z(n18068) );
  XOR U20308 ( .A(n18123), .B(n18124), .Z(n18072) );
  ANDN U20309 ( .B(n18125), .A(n18126), .Z(n18123) );
  XOR U20310 ( .A(n18127), .B(n18124), .Z(n18125) );
  IV U20311 ( .A(n18082), .Z(n18086) );
  XOR U20312 ( .A(n18082), .B(n18037), .Z(n18084) );
  XOR U20313 ( .A(n18128), .B(n18129), .Z(n18037) );
  AND U20314 ( .A(n274), .B(n18130), .Z(n18128) );
  XOR U20315 ( .A(n18131), .B(n18129), .Z(n18130) );
  NANDN U20316 ( .A(n18039), .B(n18041), .Z(n18082) );
  XOR U20317 ( .A(n18132), .B(n18133), .Z(n18041) );
  AND U20318 ( .A(n274), .B(n18134), .Z(n18132) );
  XOR U20319 ( .A(n18133), .B(n18135), .Z(n18134) );
  XNOR U20320 ( .A(n18136), .B(n18137), .Z(n274) );
  AND U20321 ( .A(n18138), .B(n18139), .Z(n18136) );
  XOR U20322 ( .A(n18137), .B(n18052), .Z(n18139) );
  XNOR U20323 ( .A(n18140), .B(n18141), .Z(n18052) );
  ANDN U20324 ( .B(n18142), .A(n18143), .Z(n18140) );
  XOR U20325 ( .A(n18141), .B(n18144), .Z(n18142) );
  XNOR U20326 ( .A(n18137), .B(n18054), .Z(n18138) );
  XOR U20327 ( .A(n18145), .B(n18146), .Z(n18054) );
  AND U20328 ( .A(n278), .B(n18147), .Z(n18145) );
  XOR U20329 ( .A(n18148), .B(n18146), .Z(n18147) );
  XNOR U20330 ( .A(n18149), .B(n18150), .Z(n18137) );
  AND U20331 ( .A(n18151), .B(n18152), .Z(n18149) );
  XNOR U20332 ( .A(n18150), .B(n18079), .Z(n18152) );
  XOR U20333 ( .A(n18143), .B(n18144), .Z(n18079) );
  XNOR U20334 ( .A(n18153), .B(n18154), .Z(n18144) );
  ANDN U20335 ( .B(n18155), .A(n18156), .Z(n18153) );
  XOR U20336 ( .A(n18157), .B(n18158), .Z(n18155) );
  XOR U20337 ( .A(n18159), .B(n18160), .Z(n18143) );
  XNOR U20338 ( .A(n18161), .B(n18162), .Z(n18160) );
  ANDN U20339 ( .B(n18163), .A(n18164), .Z(n18161) );
  XNOR U20340 ( .A(n18165), .B(n18166), .Z(n18163) );
  IV U20341 ( .A(n18141), .Z(n18159) );
  XOR U20342 ( .A(n18167), .B(n18168), .Z(n18141) );
  ANDN U20343 ( .B(n18169), .A(n18170), .Z(n18167) );
  XOR U20344 ( .A(n18168), .B(n18171), .Z(n18169) );
  XOR U20345 ( .A(n18150), .B(n18081), .Z(n18151) );
  XOR U20346 ( .A(n18172), .B(n18173), .Z(n18081) );
  AND U20347 ( .A(n278), .B(n18174), .Z(n18172) );
  XOR U20348 ( .A(n18175), .B(n18173), .Z(n18174) );
  XNOR U20349 ( .A(n18176), .B(n18177), .Z(n18150) );
  NAND U20350 ( .A(n18178), .B(n18179), .Z(n18177) );
  XOR U20351 ( .A(n18180), .B(n18129), .Z(n18179) );
  XOR U20352 ( .A(n18170), .B(n18171), .Z(n18129) );
  XOR U20353 ( .A(n18181), .B(n18158), .Z(n18171) );
  XOR U20354 ( .A(n18182), .B(n18183), .Z(n18158) );
  ANDN U20355 ( .B(n18184), .A(n18185), .Z(n18182) );
  XOR U20356 ( .A(n18183), .B(n18186), .Z(n18184) );
  IV U20357 ( .A(n18156), .Z(n18181) );
  XOR U20358 ( .A(n18154), .B(n18187), .Z(n18156) );
  XOR U20359 ( .A(n18188), .B(n18189), .Z(n18187) );
  ANDN U20360 ( .B(n18190), .A(n18191), .Z(n18188) );
  XOR U20361 ( .A(n18192), .B(n18189), .Z(n18190) );
  IV U20362 ( .A(n18157), .Z(n18154) );
  XOR U20363 ( .A(n18193), .B(n18194), .Z(n18157) );
  ANDN U20364 ( .B(n18195), .A(n18196), .Z(n18193) );
  XOR U20365 ( .A(n18194), .B(n18197), .Z(n18195) );
  XOR U20366 ( .A(n18198), .B(n18199), .Z(n18170) );
  XNOR U20367 ( .A(n18165), .B(n18200), .Z(n18199) );
  IV U20368 ( .A(n18168), .Z(n18200) );
  XOR U20369 ( .A(n18201), .B(n18202), .Z(n18168) );
  ANDN U20370 ( .B(n18203), .A(n18204), .Z(n18201) );
  XOR U20371 ( .A(n18202), .B(n18205), .Z(n18203) );
  XNOR U20372 ( .A(n18206), .B(n18207), .Z(n18165) );
  ANDN U20373 ( .B(n18208), .A(n18209), .Z(n18206) );
  XOR U20374 ( .A(n18207), .B(n18210), .Z(n18208) );
  IV U20375 ( .A(n18164), .Z(n18198) );
  XOR U20376 ( .A(n18162), .B(n18211), .Z(n18164) );
  XOR U20377 ( .A(n18212), .B(n18213), .Z(n18211) );
  ANDN U20378 ( .B(n18214), .A(n18215), .Z(n18212) );
  XOR U20379 ( .A(n18216), .B(n18213), .Z(n18214) );
  IV U20380 ( .A(n18166), .Z(n18162) );
  XOR U20381 ( .A(n18217), .B(n18218), .Z(n18166) );
  ANDN U20382 ( .B(n18219), .A(n18220), .Z(n18217) );
  XOR U20383 ( .A(n18221), .B(n18218), .Z(n18219) );
  IV U20384 ( .A(n18176), .Z(n18180) );
  XOR U20385 ( .A(n18176), .B(n18131), .Z(n18178) );
  XOR U20386 ( .A(n18222), .B(n18223), .Z(n18131) );
  AND U20387 ( .A(n278), .B(n18224), .Z(n18222) );
  XOR U20388 ( .A(n18225), .B(n18223), .Z(n18224) );
  NANDN U20389 ( .A(n18133), .B(n18135), .Z(n18176) );
  XOR U20390 ( .A(n18226), .B(n18227), .Z(n18135) );
  AND U20391 ( .A(n278), .B(n18228), .Z(n18226) );
  XOR U20392 ( .A(n18227), .B(n18229), .Z(n18228) );
  XNOR U20393 ( .A(n18230), .B(n18231), .Z(n278) );
  AND U20394 ( .A(n18232), .B(n18233), .Z(n18230) );
  XOR U20395 ( .A(n18231), .B(n18146), .Z(n18233) );
  XNOR U20396 ( .A(n18234), .B(n18235), .Z(n18146) );
  ANDN U20397 ( .B(n18236), .A(n18237), .Z(n18234) );
  XOR U20398 ( .A(n18235), .B(n18238), .Z(n18236) );
  XNOR U20399 ( .A(n18231), .B(n18148), .Z(n18232) );
  XOR U20400 ( .A(n18239), .B(n18240), .Z(n18148) );
  AND U20401 ( .A(n282), .B(n18241), .Z(n18239) );
  XOR U20402 ( .A(n18242), .B(n18240), .Z(n18241) );
  XNOR U20403 ( .A(n18243), .B(n18244), .Z(n18231) );
  AND U20404 ( .A(n18245), .B(n18246), .Z(n18243) );
  XNOR U20405 ( .A(n18244), .B(n18173), .Z(n18246) );
  XOR U20406 ( .A(n18237), .B(n18238), .Z(n18173) );
  XNOR U20407 ( .A(n18247), .B(n18248), .Z(n18238) );
  ANDN U20408 ( .B(n18249), .A(n18250), .Z(n18247) );
  XOR U20409 ( .A(n18251), .B(n18252), .Z(n18249) );
  XOR U20410 ( .A(n18253), .B(n18254), .Z(n18237) );
  XNOR U20411 ( .A(n18255), .B(n18256), .Z(n18254) );
  ANDN U20412 ( .B(n18257), .A(n18258), .Z(n18255) );
  XNOR U20413 ( .A(n18259), .B(n18260), .Z(n18257) );
  IV U20414 ( .A(n18235), .Z(n18253) );
  XOR U20415 ( .A(n18261), .B(n18262), .Z(n18235) );
  ANDN U20416 ( .B(n18263), .A(n18264), .Z(n18261) );
  XOR U20417 ( .A(n18262), .B(n18265), .Z(n18263) );
  XOR U20418 ( .A(n18244), .B(n18175), .Z(n18245) );
  XOR U20419 ( .A(n18266), .B(n18267), .Z(n18175) );
  AND U20420 ( .A(n282), .B(n18268), .Z(n18266) );
  XOR U20421 ( .A(n18269), .B(n18267), .Z(n18268) );
  XNOR U20422 ( .A(n18270), .B(n18271), .Z(n18244) );
  NAND U20423 ( .A(n18272), .B(n18273), .Z(n18271) );
  XOR U20424 ( .A(n18274), .B(n18223), .Z(n18273) );
  XOR U20425 ( .A(n18264), .B(n18265), .Z(n18223) );
  XOR U20426 ( .A(n18275), .B(n18252), .Z(n18265) );
  XOR U20427 ( .A(n18276), .B(n18277), .Z(n18252) );
  ANDN U20428 ( .B(n18278), .A(n18279), .Z(n18276) );
  XOR U20429 ( .A(n18277), .B(n18280), .Z(n18278) );
  IV U20430 ( .A(n18250), .Z(n18275) );
  XOR U20431 ( .A(n18248), .B(n18281), .Z(n18250) );
  XOR U20432 ( .A(n18282), .B(n18283), .Z(n18281) );
  ANDN U20433 ( .B(n18284), .A(n18285), .Z(n18282) );
  XOR U20434 ( .A(n18286), .B(n18283), .Z(n18284) );
  IV U20435 ( .A(n18251), .Z(n18248) );
  XOR U20436 ( .A(n18287), .B(n18288), .Z(n18251) );
  ANDN U20437 ( .B(n18289), .A(n18290), .Z(n18287) );
  XOR U20438 ( .A(n18288), .B(n18291), .Z(n18289) );
  XOR U20439 ( .A(n18292), .B(n18293), .Z(n18264) );
  XNOR U20440 ( .A(n18259), .B(n18294), .Z(n18293) );
  IV U20441 ( .A(n18262), .Z(n18294) );
  XOR U20442 ( .A(n18295), .B(n18296), .Z(n18262) );
  ANDN U20443 ( .B(n18297), .A(n18298), .Z(n18295) );
  XOR U20444 ( .A(n18296), .B(n18299), .Z(n18297) );
  XNOR U20445 ( .A(n18300), .B(n18301), .Z(n18259) );
  ANDN U20446 ( .B(n18302), .A(n18303), .Z(n18300) );
  XOR U20447 ( .A(n18301), .B(n18304), .Z(n18302) );
  IV U20448 ( .A(n18258), .Z(n18292) );
  XOR U20449 ( .A(n18256), .B(n18305), .Z(n18258) );
  XOR U20450 ( .A(n18306), .B(n18307), .Z(n18305) );
  ANDN U20451 ( .B(n18308), .A(n18309), .Z(n18306) );
  XOR U20452 ( .A(n18310), .B(n18307), .Z(n18308) );
  IV U20453 ( .A(n18260), .Z(n18256) );
  XOR U20454 ( .A(n18311), .B(n18312), .Z(n18260) );
  ANDN U20455 ( .B(n18313), .A(n18314), .Z(n18311) );
  XOR U20456 ( .A(n18315), .B(n18312), .Z(n18313) );
  IV U20457 ( .A(n18270), .Z(n18274) );
  XOR U20458 ( .A(n18270), .B(n18225), .Z(n18272) );
  XOR U20459 ( .A(n18316), .B(n18317), .Z(n18225) );
  AND U20460 ( .A(n282), .B(n18318), .Z(n18316) );
  XOR U20461 ( .A(n18319), .B(n18317), .Z(n18318) );
  NANDN U20462 ( .A(n18227), .B(n18229), .Z(n18270) );
  XOR U20463 ( .A(n18320), .B(n18321), .Z(n18229) );
  AND U20464 ( .A(n282), .B(n18322), .Z(n18320) );
  XOR U20465 ( .A(n18321), .B(n18323), .Z(n18322) );
  XNOR U20466 ( .A(n18324), .B(n18325), .Z(n282) );
  AND U20467 ( .A(n18326), .B(n18327), .Z(n18324) );
  XOR U20468 ( .A(n18325), .B(n18240), .Z(n18327) );
  XNOR U20469 ( .A(n18328), .B(n18329), .Z(n18240) );
  ANDN U20470 ( .B(n18330), .A(n18331), .Z(n18328) );
  XOR U20471 ( .A(n18329), .B(n18332), .Z(n18330) );
  XNOR U20472 ( .A(n18325), .B(n18242), .Z(n18326) );
  XOR U20473 ( .A(n18333), .B(n18334), .Z(n18242) );
  AND U20474 ( .A(n286), .B(n18335), .Z(n18333) );
  XOR U20475 ( .A(n18336), .B(n18334), .Z(n18335) );
  XNOR U20476 ( .A(n18337), .B(n18338), .Z(n18325) );
  AND U20477 ( .A(n18339), .B(n18340), .Z(n18337) );
  XNOR U20478 ( .A(n18338), .B(n18267), .Z(n18340) );
  XOR U20479 ( .A(n18331), .B(n18332), .Z(n18267) );
  XNOR U20480 ( .A(n18341), .B(n18342), .Z(n18332) );
  ANDN U20481 ( .B(n18343), .A(n18344), .Z(n18341) );
  XOR U20482 ( .A(n18345), .B(n18346), .Z(n18343) );
  XOR U20483 ( .A(n18347), .B(n18348), .Z(n18331) );
  XNOR U20484 ( .A(n18349), .B(n18350), .Z(n18348) );
  ANDN U20485 ( .B(n18351), .A(n18352), .Z(n18349) );
  XNOR U20486 ( .A(n18353), .B(n18354), .Z(n18351) );
  IV U20487 ( .A(n18329), .Z(n18347) );
  XOR U20488 ( .A(n18355), .B(n18356), .Z(n18329) );
  ANDN U20489 ( .B(n18357), .A(n18358), .Z(n18355) );
  XOR U20490 ( .A(n18356), .B(n18359), .Z(n18357) );
  XOR U20491 ( .A(n18338), .B(n18269), .Z(n18339) );
  XOR U20492 ( .A(n18360), .B(n18361), .Z(n18269) );
  AND U20493 ( .A(n286), .B(n18362), .Z(n18360) );
  XOR U20494 ( .A(n18363), .B(n18361), .Z(n18362) );
  XNOR U20495 ( .A(n18364), .B(n18365), .Z(n18338) );
  NAND U20496 ( .A(n18366), .B(n18367), .Z(n18365) );
  XOR U20497 ( .A(n18368), .B(n18317), .Z(n18367) );
  XOR U20498 ( .A(n18358), .B(n18359), .Z(n18317) );
  XOR U20499 ( .A(n18369), .B(n18346), .Z(n18359) );
  XOR U20500 ( .A(n18370), .B(n18371), .Z(n18346) );
  ANDN U20501 ( .B(n18372), .A(n18373), .Z(n18370) );
  XOR U20502 ( .A(n18371), .B(n18374), .Z(n18372) );
  IV U20503 ( .A(n18344), .Z(n18369) );
  XOR U20504 ( .A(n18342), .B(n18375), .Z(n18344) );
  XOR U20505 ( .A(n18376), .B(n18377), .Z(n18375) );
  ANDN U20506 ( .B(n18378), .A(n18379), .Z(n18376) );
  XOR U20507 ( .A(n18380), .B(n18377), .Z(n18378) );
  IV U20508 ( .A(n18345), .Z(n18342) );
  XOR U20509 ( .A(n18381), .B(n18382), .Z(n18345) );
  ANDN U20510 ( .B(n18383), .A(n18384), .Z(n18381) );
  XOR U20511 ( .A(n18382), .B(n18385), .Z(n18383) );
  XOR U20512 ( .A(n18386), .B(n18387), .Z(n18358) );
  XNOR U20513 ( .A(n18353), .B(n18388), .Z(n18387) );
  IV U20514 ( .A(n18356), .Z(n18388) );
  XOR U20515 ( .A(n18389), .B(n18390), .Z(n18356) );
  ANDN U20516 ( .B(n18391), .A(n18392), .Z(n18389) );
  XOR U20517 ( .A(n18390), .B(n18393), .Z(n18391) );
  XNOR U20518 ( .A(n18394), .B(n18395), .Z(n18353) );
  ANDN U20519 ( .B(n18396), .A(n18397), .Z(n18394) );
  XOR U20520 ( .A(n18395), .B(n18398), .Z(n18396) );
  IV U20521 ( .A(n18352), .Z(n18386) );
  XOR U20522 ( .A(n18350), .B(n18399), .Z(n18352) );
  XOR U20523 ( .A(n18400), .B(n18401), .Z(n18399) );
  ANDN U20524 ( .B(n18402), .A(n18403), .Z(n18400) );
  XOR U20525 ( .A(n18404), .B(n18401), .Z(n18402) );
  IV U20526 ( .A(n18354), .Z(n18350) );
  XOR U20527 ( .A(n18405), .B(n18406), .Z(n18354) );
  ANDN U20528 ( .B(n18407), .A(n18408), .Z(n18405) );
  XOR U20529 ( .A(n18409), .B(n18406), .Z(n18407) );
  IV U20530 ( .A(n18364), .Z(n18368) );
  XOR U20531 ( .A(n18364), .B(n18319), .Z(n18366) );
  XOR U20532 ( .A(n18410), .B(n18411), .Z(n18319) );
  AND U20533 ( .A(n286), .B(n18412), .Z(n18410) );
  XOR U20534 ( .A(n18413), .B(n18411), .Z(n18412) );
  NANDN U20535 ( .A(n18321), .B(n18323), .Z(n18364) );
  XOR U20536 ( .A(n18414), .B(n18415), .Z(n18323) );
  AND U20537 ( .A(n286), .B(n18416), .Z(n18414) );
  XOR U20538 ( .A(n18415), .B(n18417), .Z(n18416) );
  XNOR U20539 ( .A(n18418), .B(n18419), .Z(n286) );
  AND U20540 ( .A(n18420), .B(n18421), .Z(n18418) );
  XOR U20541 ( .A(n18419), .B(n18334), .Z(n18421) );
  XNOR U20542 ( .A(n18422), .B(n18423), .Z(n18334) );
  ANDN U20543 ( .B(n18424), .A(n18425), .Z(n18422) );
  XOR U20544 ( .A(n18423), .B(n18426), .Z(n18424) );
  XNOR U20545 ( .A(n18419), .B(n18336), .Z(n18420) );
  XOR U20546 ( .A(n18427), .B(n18428), .Z(n18336) );
  AND U20547 ( .A(n290), .B(n18429), .Z(n18427) );
  XOR U20548 ( .A(n18430), .B(n18428), .Z(n18429) );
  XNOR U20549 ( .A(n18431), .B(n18432), .Z(n18419) );
  AND U20550 ( .A(n18433), .B(n18434), .Z(n18431) );
  XNOR U20551 ( .A(n18432), .B(n18361), .Z(n18434) );
  XOR U20552 ( .A(n18425), .B(n18426), .Z(n18361) );
  XNOR U20553 ( .A(n18435), .B(n18436), .Z(n18426) );
  ANDN U20554 ( .B(n18437), .A(n18438), .Z(n18435) );
  XOR U20555 ( .A(n18439), .B(n18440), .Z(n18437) );
  XOR U20556 ( .A(n18441), .B(n18442), .Z(n18425) );
  XNOR U20557 ( .A(n18443), .B(n18444), .Z(n18442) );
  ANDN U20558 ( .B(n18445), .A(n18446), .Z(n18443) );
  XNOR U20559 ( .A(n18447), .B(n18448), .Z(n18445) );
  IV U20560 ( .A(n18423), .Z(n18441) );
  XOR U20561 ( .A(n18449), .B(n18450), .Z(n18423) );
  ANDN U20562 ( .B(n18451), .A(n18452), .Z(n18449) );
  XOR U20563 ( .A(n18450), .B(n18453), .Z(n18451) );
  XOR U20564 ( .A(n18432), .B(n18363), .Z(n18433) );
  XOR U20565 ( .A(n18454), .B(n18455), .Z(n18363) );
  AND U20566 ( .A(n290), .B(n18456), .Z(n18454) );
  XOR U20567 ( .A(n18457), .B(n18455), .Z(n18456) );
  XNOR U20568 ( .A(n18458), .B(n18459), .Z(n18432) );
  NAND U20569 ( .A(n18460), .B(n18461), .Z(n18459) );
  XOR U20570 ( .A(n18462), .B(n18411), .Z(n18461) );
  XOR U20571 ( .A(n18452), .B(n18453), .Z(n18411) );
  XOR U20572 ( .A(n18463), .B(n18440), .Z(n18453) );
  XOR U20573 ( .A(n18464), .B(n18465), .Z(n18440) );
  ANDN U20574 ( .B(n18466), .A(n18467), .Z(n18464) );
  XOR U20575 ( .A(n18465), .B(n18468), .Z(n18466) );
  IV U20576 ( .A(n18438), .Z(n18463) );
  XOR U20577 ( .A(n18436), .B(n18469), .Z(n18438) );
  XOR U20578 ( .A(n18470), .B(n18471), .Z(n18469) );
  ANDN U20579 ( .B(n18472), .A(n18473), .Z(n18470) );
  XOR U20580 ( .A(n18474), .B(n18471), .Z(n18472) );
  IV U20581 ( .A(n18439), .Z(n18436) );
  XOR U20582 ( .A(n18475), .B(n18476), .Z(n18439) );
  ANDN U20583 ( .B(n18477), .A(n18478), .Z(n18475) );
  XOR U20584 ( .A(n18476), .B(n18479), .Z(n18477) );
  XOR U20585 ( .A(n18480), .B(n18481), .Z(n18452) );
  XNOR U20586 ( .A(n18447), .B(n18482), .Z(n18481) );
  IV U20587 ( .A(n18450), .Z(n18482) );
  XOR U20588 ( .A(n18483), .B(n18484), .Z(n18450) );
  ANDN U20589 ( .B(n18485), .A(n18486), .Z(n18483) );
  XOR U20590 ( .A(n18484), .B(n18487), .Z(n18485) );
  XNOR U20591 ( .A(n18488), .B(n18489), .Z(n18447) );
  ANDN U20592 ( .B(n18490), .A(n18491), .Z(n18488) );
  XOR U20593 ( .A(n18489), .B(n18492), .Z(n18490) );
  IV U20594 ( .A(n18446), .Z(n18480) );
  XOR U20595 ( .A(n18444), .B(n18493), .Z(n18446) );
  XOR U20596 ( .A(n18494), .B(n18495), .Z(n18493) );
  ANDN U20597 ( .B(n18496), .A(n18497), .Z(n18494) );
  XOR U20598 ( .A(n18498), .B(n18495), .Z(n18496) );
  IV U20599 ( .A(n18448), .Z(n18444) );
  XOR U20600 ( .A(n18499), .B(n18500), .Z(n18448) );
  ANDN U20601 ( .B(n18501), .A(n18502), .Z(n18499) );
  XOR U20602 ( .A(n18503), .B(n18500), .Z(n18501) );
  IV U20603 ( .A(n18458), .Z(n18462) );
  XOR U20604 ( .A(n18458), .B(n18413), .Z(n18460) );
  XOR U20605 ( .A(n18504), .B(n18505), .Z(n18413) );
  AND U20606 ( .A(n290), .B(n18506), .Z(n18504) );
  XOR U20607 ( .A(n18507), .B(n18505), .Z(n18506) );
  NANDN U20608 ( .A(n18415), .B(n18417), .Z(n18458) );
  XOR U20609 ( .A(n18508), .B(n18509), .Z(n18417) );
  AND U20610 ( .A(n290), .B(n18510), .Z(n18508) );
  XOR U20611 ( .A(n18509), .B(n18511), .Z(n18510) );
  XNOR U20612 ( .A(n18512), .B(n18513), .Z(n290) );
  AND U20613 ( .A(n18514), .B(n18515), .Z(n18512) );
  XOR U20614 ( .A(n18513), .B(n18428), .Z(n18515) );
  XNOR U20615 ( .A(n18516), .B(n18517), .Z(n18428) );
  ANDN U20616 ( .B(n18518), .A(n18519), .Z(n18516) );
  XOR U20617 ( .A(n18517), .B(n18520), .Z(n18518) );
  XNOR U20618 ( .A(n18513), .B(n18430), .Z(n18514) );
  XOR U20619 ( .A(n18521), .B(n18522), .Z(n18430) );
  AND U20620 ( .A(n294), .B(n18523), .Z(n18521) );
  XOR U20621 ( .A(n18524), .B(n18522), .Z(n18523) );
  XNOR U20622 ( .A(n18525), .B(n18526), .Z(n18513) );
  AND U20623 ( .A(n18527), .B(n18528), .Z(n18525) );
  XNOR U20624 ( .A(n18526), .B(n18455), .Z(n18528) );
  XOR U20625 ( .A(n18519), .B(n18520), .Z(n18455) );
  XNOR U20626 ( .A(n18529), .B(n18530), .Z(n18520) );
  ANDN U20627 ( .B(n18531), .A(n18532), .Z(n18529) );
  XOR U20628 ( .A(n18533), .B(n18534), .Z(n18531) );
  XOR U20629 ( .A(n18535), .B(n18536), .Z(n18519) );
  XNOR U20630 ( .A(n18537), .B(n18538), .Z(n18536) );
  ANDN U20631 ( .B(n18539), .A(n18540), .Z(n18537) );
  XNOR U20632 ( .A(n18541), .B(n18542), .Z(n18539) );
  IV U20633 ( .A(n18517), .Z(n18535) );
  XOR U20634 ( .A(n18543), .B(n18544), .Z(n18517) );
  ANDN U20635 ( .B(n18545), .A(n18546), .Z(n18543) );
  XOR U20636 ( .A(n18544), .B(n18547), .Z(n18545) );
  XOR U20637 ( .A(n18526), .B(n18457), .Z(n18527) );
  XOR U20638 ( .A(n18548), .B(n18549), .Z(n18457) );
  AND U20639 ( .A(n294), .B(n18550), .Z(n18548) );
  XOR U20640 ( .A(n18551), .B(n18549), .Z(n18550) );
  XNOR U20641 ( .A(n18552), .B(n18553), .Z(n18526) );
  NAND U20642 ( .A(n18554), .B(n18555), .Z(n18553) );
  XOR U20643 ( .A(n18556), .B(n18505), .Z(n18555) );
  XOR U20644 ( .A(n18546), .B(n18547), .Z(n18505) );
  XOR U20645 ( .A(n18557), .B(n18534), .Z(n18547) );
  XOR U20646 ( .A(n18558), .B(n18559), .Z(n18534) );
  ANDN U20647 ( .B(n18560), .A(n18561), .Z(n18558) );
  XOR U20648 ( .A(n18559), .B(n18562), .Z(n18560) );
  IV U20649 ( .A(n18532), .Z(n18557) );
  XOR U20650 ( .A(n18530), .B(n18563), .Z(n18532) );
  XOR U20651 ( .A(n18564), .B(n18565), .Z(n18563) );
  ANDN U20652 ( .B(n18566), .A(n18567), .Z(n18564) );
  XOR U20653 ( .A(n18568), .B(n18565), .Z(n18566) );
  IV U20654 ( .A(n18533), .Z(n18530) );
  XOR U20655 ( .A(n18569), .B(n18570), .Z(n18533) );
  ANDN U20656 ( .B(n18571), .A(n18572), .Z(n18569) );
  XOR U20657 ( .A(n18570), .B(n18573), .Z(n18571) );
  XOR U20658 ( .A(n18574), .B(n18575), .Z(n18546) );
  XNOR U20659 ( .A(n18541), .B(n18576), .Z(n18575) );
  IV U20660 ( .A(n18544), .Z(n18576) );
  XOR U20661 ( .A(n18577), .B(n18578), .Z(n18544) );
  ANDN U20662 ( .B(n18579), .A(n18580), .Z(n18577) );
  XOR U20663 ( .A(n18578), .B(n18581), .Z(n18579) );
  XNOR U20664 ( .A(n18582), .B(n18583), .Z(n18541) );
  ANDN U20665 ( .B(n18584), .A(n18585), .Z(n18582) );
  XOR U20666 ( .A(n18583), .B(n18586), .Z(n18584) );
  IV U20667 ( .A(n18540), .Z(n18574) );
  XOR U20668 ( .A(n18538), .B(n18587), .Z(n18540) );
  XOR U20669 ( .A(n18588), .B(n18589), .Z(n18587) );
  ANDN U20670 ( .B(n18590), .A(n18591), .Z(n18588) );
  XOR U20671 ( .A(n18592), .B(n18589), .Z(n18590) );
  IV U20672 ( .A(n18542), .Z(n18538) );
  XOR U20673 ( .A(n18593), .B(n18594), .Z(n18542) );
  ANDN U20674 ( .B(n18595), .A(n18596), .Z(n18593) );
  XOR U20675 ( .A(n18597), .B(n18594), .Z(n18595) );
  IV U20676 ( .A(n18552), .Z(n18556) );
  XOR U20677 ( .A(n18552), .B(n18507), .Z(n18554) );
  XOR U20678 ( .A(n18598), .B(n18599), .Z(n18507) );
  AND U20679 ( .A(n294), .B(n18600), .Z(n18598) );
  XOR U20680 ( .A(n18601), .B(n18599), .Z(n18600) );
  NANDN U20681 ( .A(n18509), .B(n18511), .Z(n18552) );
  XOR U20682 ( .A(n18602), .B(n18603), .Z(n18511) );
  AND U20683 ( .A(n294), .B(n18604), .Z(n18602) );
  XOR U20684 ( .A(n18603), .B(n18605), .Z(n18604) );
  XNOR U20685 ( .A(n18606), .B(n18607), .Z(n294) );
  AND U20686 ( .A(n18608), .B(n18609), .Z(n18606) );
  XOR U20687 ( .A(n18607), .B(n18522), .Z(n18609) );
  XNOR U20688 ( .A(n18610), .B(n18611), .Z(n18522) );
  ANDN U20689 ( .B(n18612), .A(n18613), .Z(n18610) );
  XOR U20690 ( .A(n18611), .B(n18614), .Z(n18612) );
  XNOR U20691 ( .A(n18607), .B(n18524), .Z(n18608) );
  XOR U20692 ( .A(n18615), .B(n18616), .Z(n18524) );
  AND U20693 ( .A(n298), .B(n18617), .Z(n18615) );
  XOR U20694 ( .A(n18618), .B(n18616), .Z(n18617) );
  XNOR U20695 ( .A(n18619), .B(n18620), .Z(n18607) );
  AND U20696 ( .A(n18621), .B(n18622), .Z(n18619) );
  XNOR U20697 ( .A(n18620), .B(n18549), .Z(n18622) );
  XOR U20698 ( .A(n18613), .B(n18614), .Z(n18549) );
  XNOR U20699 ( .A(n18623), .B(n18624), .Z(n18614) );
  ANDN U20700 ( .B(n18625), .A(n18626), .Z(n18623) );
  XOR U20701 ( .A(n18627), .B(n18628), .Z(n18625) );
  XOR U20702 ( .A(n18629), .B(n18630), .Z(n18613) );
  XNOR U20703 ( .A(n18631), .B(n18632), .Z(n18630) );
  ANDN U20704 ( .B(n18633), .A(n18634), .Z(n18631) );
  XNOR U20705 ( .A(n18635), .B(n18636), .Z(n18633) );
  IV U20706 ( .A(n18611), .Z(n18629) );
  XOR U20707 ( .A(n18637), .B(n18638), .Z(n18611) );
  ANDN U20708 ( .B(n18639), .A(n18640), .Z(n18637) );
  XOR U20709 ( .A(n18638), .B(n18641), .Z(n18639) );
  XOR U20710 ( .A(n18620), .B(n18551), .Z(n18621) );
  XOR U20711 ( .A(n18642), .B(n18643), .Z(n18551) );
  AND U20712 ( .A(n298), .B(n18644), .Z(n18642) );
  XOR U20713 ( .A(n18645), .B(n18643), .Z(n18644) );
  XNOR U20714 ( .A(n18646), .B(n18647), .Z(n18620) );
  NAND U20715 ( .A(n18648), .B(n18649), .Z(n18647) );
  XOR U20716 ( .A(n18650), .B(n18599), .Z(n18649) );
  XOR U20717 ( .A(n18640), .B(n18641), .Z(n18599) );
  XOR U20718 ( .A(n18651), .B(n18628), .Z(n18641) );
  XOR U20719 ( .A(n18652), .B(n18653), .Z(n18628) );
  ANDN U20720 ( .B(n18654), .A(n18655), .Z(n18652) );
  XOR U20721 ( .A(n18653), .B(n18656), .Z(n18654) );
  IV U20722 ( .A(n18626), .Z(n18651) );
  XOR U20723 ( .A(n18624), .B(n18657), .Z(n18626) );
  XOR U20724 ( .A(n18658), .B(n18659), .Z(n18657) );
  ANDN U20725 ( .B(n18660), .A(n18661), .Z(n18658) );
  XOR U20726 ( .A(n18662), .B(n18659), .Z(n18660) );
  IV U20727 ( .A(n18627), .Z(n18624) );
  XOR U20728 ( .A(n18663), .B(n18664), .Z(n18627) );
  ANDN U20729 ( .B(n18665), .A(n18666), .Z(n18663) );
  XOR U20730 ( .A(n18664), .B(n18667), .Z(n18665) );
  XOR U20731 ( .A(n18668), .B(n18669), .Z(n18640) );
  XNOR U20732 ( .A(n18635), .B(n18670), .Z(n18669) );
  IV U20733 ( .A(n18638), .Z(n18670) );
  XOR U20734 ( .A(n18671), .B(n18672), .Z(n18638) );
  ANDN U20735 ( .B(n18673), .A(n18674), .Z(n18671) );
  XOR U20736 ( .A(n18672), .B(n18675), .Z(n18673) );
  XNOR U20737 ( .A(n18676), .B(n18677), .Z(n18635) );
  ANDN U20738 ( .B(n18678), .A(n18679), .Z(n18676) );
  XOR U20739 ( .A(n18677), .B(n18680), .Z(n18678) );
  IV U20740 ( .A(n18634), .Z(n18668) );
  XOR U20741 ( .A(n18632), .B(n18681), .Z(n18634) );
  XOR U20742 ( .A(n18682), .B(n18683), .Z(n18681) );
  ANDN U20743 ( .B(n18684), .A(n18685), .Z(n18682) );
  XOR U20744 ( .A(n18686), .B(n18683), .Z(n18684) );
  IV U20745 ( .A(n18636), .Z(n18632) );
  XOR U20746 ( .A(n18687), .B(n18688), .Z(n18636) );
  ANDN U20747 ( .B(n18689), .A(n18690), .Z(n18687) );
  XOR U20748 ( .A(n18691), .B(n18688), .Z(n18689) );
  IV U20749 ( .A(n18646), .Z(n18650) );
  XOR U20750 ( .A(n18646), .B(n18601), .Z(n18648) );
  XOR U20751 ( .A(n18692), .B(n18693), .Z(n18601) );
  AND U20752 ( .A(n298), .B(n18694), .Z(n18692) );
  XOR U20753 ( .A(n18695), .B(n18693), .Z(n18694) );
  NANDN U20754 ( .A(n18603), .B(n18605), .Z(n18646) );
  XOR U20755 ( .A(n18696), .B(n18697), .Z(n18605) );
  AND U20756 ( .A(n298), .B(n18698), .Z(n18696) );
  XOR U20757 ( .A(n18697), .B(n18699), .Z(n18698) );
  XNOR U20758 ( .A(n18700), .B(n18701), .Z(n298) );
  AND U20759 ( .A(n18702), .B(n18703), .Z(n18700) );
  XOR U20760 ( .A(n18701), .B(n18616), .Z(n18703) );
  XNOR U20761 ( .A(n18704), .B(n18705), .Z(n18616) );
  ANDN U20762 ( .B(n18706), .A(n18707), .Z(n18704) );
  XOR U20763 ( .A(n18705), .B(n18708), .Z(n18706) );
  XNOR U20764 ( .A(n18701), .B(n18618), .Z(n18702) );
  XOR U20765 ( .A(n18709), .B(n18710), .Z(n18618) );
  AND U20766 ( .A(n302), .B(n18711), .Z(n18709) );
  XOR U20767 ( .A(n18712), .B(n18710), .Z(n18711) );
  XNOR U20768 ( .A(n18713), .B(n18714), .Z(n18701) );
  AND U20769 ( .A(n18715), .B(n18716), .Z(n18713) );
  XNOR U20770 ( .A(n18714), .B(n18643), .Z(n18716) );
  XOR U20771 ( .A(n18707), .B(n18708), .Z(n18643) );
  XNOR U20772 ( .A(n18717), .B(n18718), .Z(n18708) );
  ANDN U20773 ( .B(n18719), .A(n18720), .Z(n18717) );
  XOR U20774 ( .A(n18721), .B(n18722), .Z(n18719) );
  XOR U20775 ( .A(n18723), .B(n18724), .Z(n18707) );
  XNOR U20776 ( .A(n18725), .B(n18726), .Z(n18724) );
  ANDN U20777 ( .B(n18727), .A(n18728), .Z(n18725) );
  XNOR U20778 ( .A(n18729), .B(n18730), .Z(n18727) );
  IV U20779 ( .A(n18705), .Z(n18723) );
  XOR U20780 ( .A(n18731), .B(n18732), .Z(n18705) );
  ANDN U20781 ( .B(n18733), .A(n18734), .Z(n18731) );
  XOR U20782 ( .A(n18732), .B(n18735), .Z(n18733) );
  XOR U20783 ( .A(n18714), .B(n18645), .Z(n18715) );
  XOR U20784 ( .A(n18736), .B(n18737), .Z(n18645) );
  AND U20785 ( .A(n302), .B(n18738), .Z(n18736) );
  XOR U20786 ( .A(n18739), .B(n18737), .Z(n18738) );
  XNOR U20787 ( .A(n18740), .B(n18741), .Z(n18714) );
  NAND U20788 ( .A(n18742), .B(n18743), .Z(n18741) );
  XOR U20789 ( .A(n18744), .B(n18693), .Z(n18743) );
  XOR U20790 ( .A(n18734), .B(n18735), .Z(n18693) );
  XOR U20791 ( .A(n18745), .B(n18722), .Z(n18735) );
  XOR U20792 ( .A(n18746), .B(n18747), .Z(n18722) );
  ANDN U20793 ( .B(n18748), .A(n18749), .Z(n18746) );
  XOR U20794 ( .A(n18747), .B(n18750), .Z(n18748) );
  IV U20795 ( .A(n18720), .Z(n18745) );
  XOR U20796 ( .A(n18718), .B(n18751), .Z(n18720) );
  XOR U20797 ( .A(n18752), .B(n18753), .Z(n18751) );
  ANDN U20798 ( .B(n18754), .A(n18755), .Z(n18752) );
  XOR U20799 ( .A(n18756), .B(n18753), .Z(n18754) );
  IV U20800 ( .A(n18721), .Z(n18718) );
  XOR U20801 ( .A(n18757), .B(n18758), .Z(n18721) );
  ANDN U20802 ( .B(n18759), .A(n18760), .Z(n18757) );
  XOR U20803 ( .A(n18758), .B(n18761), .Z(n18759) );
  XOR U20804 ( .A(n18762), .B(n18763), .Z(n18734) );
  XNOR U20805 ( .A(n18729), .B(n18764), .Z(n18763) );
  IV U20806 ( .A(n18732), .Z(n18764) );
  XOR U20807 ( .A(n18765), .B(n18766), .Z(n18732) );
  ANDN U20808 ( .B(n18767), .A(n18768), .Z(n18765) );
  XOR U20809 ( .A(n18766), .B(n18769), .Z(n18767) );
  XNOR U20810 ( .A(n18770), .B(n18771), .Z(n18729) );
  ANDN U20811 ( .B(n18772), .A(n18773), .Z(n18770) );
  XOR U20812 ( .A(n18771), .B(n18774), .Z(n18772) );
  IV U20813 ( .A(n18728), .Z(n18762) );
  XOR U20814 ( .A(n18726), .B(n18775), .Z(n18728) );
  XOR U20815 ( .A(n18776), .B(n18777), .Z(n18775) );
  ANDN U20816 ( .B(n18778), .A(n18779), .Z(n18776) );
  XOR U20817 ( .A(n18780), .B(n18777), .Z(n18778) );
  IV U20818 ( .A(n18730), .Z(n18726) );
  XOR U20819 ( .A(n18781), .B(n18782), .Z(n18730) );
  ANDN U20820 ( .B(n18783), .A(n18784), .Z(n18781) );
  XOR U20821 ( .A(n18785), .B(n18782), .Z(n18783) );
  IV U20822 ( .A(n18740), .Z(n18744) );
  XOR U20823 ( .A(n18740), .B(n18695), .Z(n18742) );
  XOR U20824 ( .A(n18786), .B(n18787), .Z(n18695) );
  AND U20825 ( .A(n302), .B(n18788), .Z(n18786) );
  XOR U20826 ( .A(n18789), .B(n18787), .Z(n18788) );
  NANDN U20827 ( .A(n18697), .B(n18699), .Z(n18740) );
  XOR U20828 ( .A(n18790), .B(n18791), .Z(n18699) );
  AND U20829 ( .A(n302), .B(n18792), .Z(n18790) );
  XOR U20830 ( .A(n18791), .B(n18793), .Z(n18792) );
  XNOR U20831 ( .A(n18794), .B(n18795), .Z(n302) );
  AND U20832 ( .A(n18796), .B(n18797), .Z(n18794) );
  XOR U20833 ( .A(n18795), .B(n18710), .Z(n18797) );
  XNOR U20834 ( .A(n18798), .B(n18799), .Z(n18710) );
  ANDN U20835 ( .B(n18800), .A(n18801), .Z(n18798) );
  XOR U20836 ( .A(n18799), .B(n18802), .Z(n18800) );
  XNOR U20837 ( .A(n18795), .B(n18712), .Z(n18796) );
  XOR U20838 ( .A(n18803), .B(n18804), .Z(n18712) );
  AND U20839 ( .A(n306), .B(n18805), .Z(n18803) );
  XOR U20840 ( .A(n18806), .B(n18804), .Z(n18805) );
  XNOR U20841 ( .A(n18807), .B(n18808), .Z(n18795) );
  AND U20842 ( .A(n18809), .B(n18810), .Z(n18807) );
  XNOR U20843 ( .A(n18808), .B(n18737), .Z(n18810) );
  XOR U20844 ( .A(n18801), .B(n18802), .Z(n18737) );
  XNOR U20845 ( .A(n18811), .B(n18812), .Z(n18802) );
  ANDN U20846 ( .B(n18813), .A(n18814), .Z(n18811) );
  XOR U20847 ( .A(n18815), .B(n18816), .Z(n18813) );
  XOR U20848 ( .A(n18817), .B(n18818), .Z(n18801) );
  XNOR U20849 ( .A(n18819), .B(n18820), .Z(n18818) );
  ANDN U20850 ( .B(n18821), .A(n18822), .Z(n18819) );
  XNOR U20851 ( .A(n18823), .B(n18824), .Z(n18821) );
  IV U20852 ( .A(n18799), .Z(n18817) );
  XOR U20853 ( .A(n18825), .B(n18826), .Z(n18799) );
  ANDN U20854 ( .B(n18827), .A(n18828), .Z(n18825) );
  XOR U20855 ( .A(n18826), .B(n18829), .Z(n18827) );
  XOR U20856 ( .A(n18808), .B(n18739), .Z(n18809) );
  XOR U20857 ( .A(n18830), .B(n18831), .Z(n18739) );
  AND U20858 ( .A(n306), .B(n18832), .Z(n18830) );
  XOR U20859 ( .A(n18833), .B(n18831), .Z(n18832) );
  XNOR U20860 ( .A(n18834), .B(n18835), .Z(n18808) );
  NAND U20861 ( .A(n18836), .B(n18837), .Z(n18835) );
  XOR U20862 ( .A(n18838), .B(n18787), .Z(n18837) );
  XOR U20863 ( .A(n18828), .B(n18829), .Z(n18787) );
  XOR U20864 ( .A(n18839), .B(n18816), .Z(n18829) );
  XOR U20865 ( .A(n18840), .B(n18841), .Z(n18816) );
  ANDN U20866 ( .B(n18842), .A(n18843), .Z(n18840) );
  XOR U20867 ( .A(n18841), .B(n18844), .Z(n18842) );
  IV U20868 ( .A(n18814), .Z(n18839) );
  XOR U20869 ( .A(n18812), .B(n18845), .Z(n18814) );
  XOR U20870 ( .A(n18846), .B(n18847), .Z(n18845) );
  ANDN U20871 ( .B(n18848), .A(n18849), .Z(n18846) );
  XOR U20872 ( .A(n18850), .B(n18847), .Z(n18848) );
  IV U20873 ( .A(n18815), .Z(n18812) );
  XOR U20874 ( .A(n18851), .B(n18852), .Z(n18815) );
  ANDN U20875 ( .B(n18853), .A(n18854), .Z(n18851) );
  XOR U20876 ( .A(n18852), .B(n18855), .Z(n18853) );
  XOR U20877 ( .A(n18856), .B(n18857), .Z(n18828) );
  XNOR U20878 ( .A(n18823), .B(n18858), .Z(n18857) );
  IV U20879 ( .A(n18826), .Z(n18858) );
  XOR U20880 ( .A(n18859), .B(n18860), .Z(n18826) );
  ANDN U20881 ( .B(n18861), .A(n18862), .Z(n18859) );
  XOR U20882 ( .A(n18860), .B(n18863), .Z(n18861) );
  XNOR U20883 ( .A(n18864), .B(n18865), .Z(n18823) );
  ANDN U20884 ( .B(n18866), .A(n18867), .Z(n18864) );
  XOR U20885 ( .A(n18865), .B(n18868), .Z(n18866) );
  IV U20886 ( .A(n18822), .Z(n18856) );
  XOR U20887 ( .A(n18820), .B(n18869), .Z(n18822) );
  XOR U20888 ( .A(n18870), .B(n18871), .Z(n18869) );
  ANDN U20889 ( .B(n18872), .A(n18873), .Z(n18870) );
  XOR U20890 ( .A(n18874), .B(n18871), .Z(n18872) );
  IV U20891 ( .A(n18824), .Z(n18820) );
  XOR U20892 ( .A(n18875), .B(n18876), .Z(n18824) );
  ANDN U20893 ( .B(n18877), .A(n18878), .Z(n18875) );
  XOR U20894 ( .A(n18879), .B(n18876), .Z(n18877) );
  IV U20895 ( .A(n18834), .Z(n18838) );
  XOR U20896 ( .A(n18834), .B(n18789), .Z(n18836) );
  XOR U20897 ( .A(n18880), .B(n18881), .Z(n18789) );
  AND U20898 ( .A(n306), .B(n18882), .Z(n18880) );
  XOR U20899 ( .A(n18883), .B(n18881), .Z(n18882) );
  NANDN U20900 ( .A(n18791), .B(n18793), .Z(n18834) );
  XOR U20901 ( .A(n18884), .B(n18885), .Z(n18793) );
  AND U20902 ( .A(n306), .B(n18886), .Z(n18884) );
  XOR U20903 ( .A(n18885), .B(n18887), .Z(n18886) );
  XNOR U20904 ( .A(n18888), .B(n18889), .Z(n306) );
  AND U20905 ( .A(n18890), .B(n18891), .Z(n18888) );
  XOR U20906 ( .A(n18889), .B(n18804), .Z(n18891) );
  XNOR U20907 ( .A(n18892), .B(n18893), .Z(n18804) );
  ANDN U20908 ( .B(n18894), .A(n18895), .Z(n18892) );
  XOR U20909 ( .A(n18893), .B(n18896), .Z(n18894) );
  XNOR U20910 ( .A(n18889), .B(n18806), .Z(n18890) );
  XOR U20911 ( .A(n18897), .B(n18898), .Z(n18806) );
  AND U20912 ( .A(n310), .B(n18899), .Z(n18897) );
  XOR U20913 ( .A(n18900), .B(n18898), .Z(n18899) );
  XNOR U20914 ( .A(n18901), .B(n18902), .Z(n18889) );
  AND U20915 ( .A(n18903), .B(n18904), .Z(n18901) );
  XNOR U20916 ( .A(n18902), .B(n18831), .Z(n18904) );
  XOR U20917 ( .A(n18895), .B(n18896), .Z(n18831) );
  XNOR U20918 ( .A(n18905), .B(n18906), .Z(n18896) );
  ANDN U20919 ( .B(n18907), .A(n18908), .Z(n18905) );
  XOR U20920 ( .A(n18909), .B(n18910), .Z(n18907) );
  XOR U20921 ( .A(n18911), .B(n18912), .Z(n18895) );
  XNOR U20922 ( .A(n18913), .B(n18914), .Z(n18912) );
  ANDN U20923 ( .B(n18915), .A(n18916), .Z(n18913) );
  XNOR U20924 ( .A(n18917), .B(n18918), .Z(n18915) );
  IV U20925 ( .A(n18893), .Z(n18911) );
  XOR U20926 ( .A(n18919), .B(n18920), .Z(n18893) );
  ANDN U20927 ( .B(n18921), .A(n18922), .Z(n18919) );
  XOR U20928 ( .A(n18920), .B(n18923), .Z(n18921) );
  XOR U20929 ( .A(n18902), .B(n18833), .Z(n18903) );
  XOR U20930 ( .A(n18924), .B(n18925), .Z(n18833) );
  AND U20931 ( .A(n310), .B(n18926), .Z(n18924) );
  XOR U20932 ( .A(n18927), .B(n18925), .Z(n18926) );
  XNOR U20933 ( .A(n18928), .B(n18929), .Z(n18902) );
  NAND U20934 ( .A(n18930), .B(n18931), .Z(n18929) );
  XOR U20935 ( .A(n18932), .B(n18881), .Z(n18931) );
  XOR U20936 ( .A(n18922), .B(n18923), .Z(n18881) );
  XOR U20937 ( .A(n18933), .B(n18910), .Z(n18923) );
  XOR U20938 ( .A(n18934), .B(n18935), .Z(n18910) );
  ANDN U20939 ( .B(n18936), .A(n18937), .Z(n18934) );
  XOR U20940 ( .A(n18935), .B(n18938), .Z(n18936) );
  IV U20941 ( .A(n18908), .Z(n18933) );
  XOR U20942 ( .A(n18906), .B(n18939), .Z(n18908) );
  XOR U20943 ( .A(n18940), .B(n18941), .Z(n18939) );
  ANDN U20944 ( .B(n18942), .A(n18943), .Z(n18940) );
  XOR U20945 ( .A(n18944), .B(n18941), .Z(n18942) );
  IV U20946 ( .A(n18909), .Z(n18906) );
  XOR U20947 ( .A(n18945), .B(n18946), .Z(n18909) );
  ANDN U20948 ( .B(n18947), .A(n18948), .Z(n18945) );
  XOR U20949 ( .A(n18946), .B(n18949), .Z(n18947) );
  XOR U20950 ( .A(n18950), .B(n18951), .Z(n18922) );
  XNOR U20951 ( .A(n18917), .B(n18952), .Z(n18951) );
  IV U20952 ( .A(n18920), .Z(n18952) );
  XOR U20953 ( .A(n18953), .B(n18954), .Z(n18920) );
  ANDN U20954 ( .B(n18955), .A(n18956), .Z(n18953) );
  XOR U20955 ( .A(n18954), .B(n18957), .Z(n18955) );
  XNOR U20956 ( .A(n18958), .B(n18959), .Z(n18917) );
  ANDN U20957 ( .B(n18960), .A(n18961), .Z(n18958) );
  XOR U20958 ( .A(n18959), .B(n18962), .Z(n18960) );
  IV U20959 ( .A(n18916), .Z(n18950) );
  XOR U20960 ( .A(n18914), .B(n18963), .Z(n18916) );
  XOR U20961 ( .A(n18964), .B(n18965), .Z(n18963) );
  ANDN U20962 ( .B(n18966), .A(n18967), .Z(n18964) );
  XOR U20963 ( .A(n18968), .B(n18965), .Z(n18966) );
  IV U20964 ( .A(n18918), .Z(n18914) );
  XOR U20965 ( .A(n18969), .B(n18970), .Z(n18918) );
  ANDN U20966 ( .B(n18971), .A(n18972), .Z(n18969) );
  XOR U20967 ( .A(n18973), .B(n18970), .Z(n18971) );
  IV U20968 ( .A(n18928), .Z(n18932) );
  XOR U20969 ( .A(n18928), .B(n18883), .Z(n18930) );
  XOR U20970 ( .A(n18974), .B(n18975), .Z(n18883) );
  AND U20971 ( .A(n310), .B(n18976), .Z(n18974) );
  XOR U20972 ( .A(n18977), .B(n18975), .Z(n18976) );
  NANDN U20973 ( .A(n18885), .B(n18887), .Z(n18928) );
  XOR U20974 ( .A(n18978), .B(n18979), .Z(n18887) );
  AND U20975 ( .A(n310), .B(n18980), .Z(n18978) );
  XOR U20976 ( .A(n18979), .B(n18981), .Z(n18980) );
  XNOR U20977 ( .A(n18982), .B(n18983), .Z(n310) );
  AND U20978 ( .A(n18984), .B(n18985), .Z(n18982) );
  XOR U20979 ( .A(n18983), .B(n18898), .Z(n18985) );
  XNOR U20980 ( .A(n18986), .B(n18987), .Z(n18898) );
  ANDN U20981 ( .B(n18988), .A(n18989), .Z(n18986) );
  XOR U20982 ( .A(n18987), .B(n18990), .Z(n18988) );
  XNOR U20983 ( .A(n18983), .B(n18900), .Z(n18984) );
  XOR U20984 ( .A(n18991), .B(n18992), .Z(n18900) );
  AND U20985 ( .A(n314), .B(n18993), .Z(n18991) );
  XOR U20986 ( .A(n18994), .B(n18992), .Z(n18993) );
  XNOR U20987 ( .A(n18995), .B(n18996), .Z(n18983) );
  AND U20988 ( .A(n18997), .B(n18998), .Z(n18995) );
  XNOR U20989 ( .A(n18996), .B(n18925), .Z(n18998) );
  XOR U20990 ( .A(n18989), .B(n18990), .Z(n18925) );
  XNOR U20991 ( .A(n18999), .B(n19000), .Z(n18990) );
  ANDN U20992 ( .B(n19001), .A(n19002), .Z(n18999) );
  XOR U20993 ( .A(n19003), .B(n19004), .Z(n19001) );
  XOR U20994 ( .A(n19005), .B(n19006), .Z(n18989) );
  XNOR U20995 ( .A(n19007), .B(n19008), .Z(n19006) );
  ANDN U20996 ( .B(n19009), .A(n19010), .Z(n19007) );
  XNOR U20997 ( .A(n19011), .B(n19012), .Z(n19009) );
  IV U20998 ( .A(n18987), .Z(n19005) );
  XOR U20999 ( .A(n19013), .B(n19014), .Z(n18987) );
  ANDN U21000 ( .B(n19015), .A(n19016), .Z(n19013) );
  XOR U21001 ( .A(n19014), .B(n19017), .Z(n19015) );
  XOR U21002 ( .A(n18996), .B(n18927), .Z(n18997) );
  XOR U21003 ( .A(n19018), .B(n19019), .Z(n18927) );
  AND U21004 ( .A(n314), .B(n19020), .Z(n19018) );
  XOR U21005 ( .A(n19021), .B(n19019), .Z(n19020) );
  XNOR U21006 ( .A(n19022), .B(n19023), .Z(n18996) );
  NAND U21007 ( .A(n19024), .B(n19025), .Z(n19023) );
  XOR U21008 ( .A(n19026), .B(n18975), .Z(n19025) );
  XOR U21009 ( .A(n19016), .B(n19017), .Z(n18975) );
  XOR U21010 ( .A(n19027), .B(n19004), .Z(n19017) );
  XOR U21011 ( .A(n19028), .B(n19029), .Z(n19004) );
  ANDN U21012 ( .B(n19030), .A(n19031), .Z(n19028) );
  XOR U21013 ( .A(n19029), .B(n19032), .Z(n19030) );
  IV U21014 ( .A(n19002), .Z(n19027) );
  XOR U21015 ( .A(n19000), .B(n19033), .Z(n19002) );
  XOR U21016 ( .A(n19034), .B(n19035), .Z(n19033) );
  ANDN U21017 ( .B(n19036), .A(n19037), .Z(n19034) );
  XOR U21018 ( .A(n19038), .B(n19035), .Z(n19036) );
  IV U21019 ( .A(n19003), .Z(n19000) );
  XOR U21020 ( .A(n19039), .B(n19040), .Z(n19003) );
  ANDN U21021 ( .B(n19041), .A(n19042), .Z(n19039) );
  XOR U21022 ( .A(n19040), .B(n19043), .Z(n19041) );
  XOR U21023 ( .A(n19044), .B(n19045), .Z(n19016) );
  XNOR U21024 ( .A(n19011), .B(n19046), .Z(n19045) );
  IV U21025 ( .A(n19014), .Z(n19046) );
  XOR U21026 ( .A(n19047), .B(n19048), .Z(n19014) );
  ANDN U21027 ( .B(n19049), .A(n19050), .Z(n19047) );
  XOR U21028 ( .A(n19048), .B(n19051), .Z(n19049) );
  XNOR U21029 ( .A(n19052), .B(n19053), .Z(n19011) );
  ANDN U21030 ( .B(n19054), .A(n19055), .Z(n19052) );
  XOR U21031 ( .A(n19053), .B(n19056), .Z(n19054) );
  IV U21032 ( .A(n19010), .Z(n19044) );
  XOR U21033 ( .A(n19008), .B(n19057), .Z(n19010) );
  XOR U21034 ( .A(n19058), .B(n19059), .Z(n19057) );
  ANDN U21035 ( .B(n19060), .A(n19061), .Z(n19058) );
  XOR U21036 ( .A(n19062), .B(n19059), .Z(n19060) );
  IV U21037 ( .A(n19012), .Z(n19008) );
  XOR U21038 ( .A(n19063), .B(n19064), .Z(n19012) );
  ANDN U21039 ( .B(n19065), .A(n19066), .Z(n19063) );
  XOR U21040 ( .A(n19067), .B(n19064), .Z(n19065) );
  IV U21041 ( .A(n19022), .Z(n19026) );
  XOR U21042 ( .A(n19022), .B(n18977), .Z(n19024) );
  XOR U21043 ( .A(n19068), .B(n19069), .Z(n18977) );
  AND U21044 ( .A(n314), .B(n19070), .Z(n19068) );
  XOR U21045 ( .A(n19071), .B(n19069), .Z(n19070) );
  NANDN U21046 ( .A(n18979), .B(n18981), .Z(n19022) );
  XOR U21047 ( .A(n19072), .B(n19073), .Z(n18981) );
  AND U21048 ( .A(n314), .B(n19074), .Z(n19072) );
  XOR U21049 ( .A(n19073), .B(n19075), .Z(n19074) );
  XNOR U21050 ( .A(n19076), .B(n19077), .Z(n314) );
  AND U21051 ( .A(n19078), .B(n19079), .Z(n19076) );
  XOR U21052 ( .A(n19077), .B(n18992), .Z(n19079) );
  XNOR U21053 ( .A(n19080), .B(n19081), .Z(n18992) );
  ANDN U21054 ( .B(n19082), .A(n19083), .Z(n19080) );
  XOR U21055 ( .A(n19081), .B(n19084), .Z(n19082) );
  XNOR U21056 ( .A(n19077), .B(n18994), .Z(n19078) );
  XOR U21057 ( .A(n19085), .B(n19086), .Z(n18994) );
  AND U21058 ( .A(n318), .B(n19087), .Z(n19085) );
  XOR U21059 ( .A(n19088), .B(n19086), .Z(n19087) );
  XNOR U21060 ( .A(n19089), .B(n19090), .Z(n19077) );
  AND U21061 ( .A(n19091), .B(n19092), .Z(n19089) );
  XNOR U21062 ( .A(n19090), .B(n19019), .Z(n19092) );
  XOR U21063 ( .A(n19083), .B(n19084), .Z(n19019) );
  XNOR U21064 ( .A(n19093), .B(n19094), .Z(n19084) );
  ANDN U21065 ( .B(n19095), .A(n19096), .Z(n19093) );
  XOR U21066 ( .A(n19097), .B(n19098), .Z(n19095) );
  XOR U21067 ( .A(n19099), .B(n19100), .Z(n19083) );
  XNOR U21068 ( .A(n19101), .B(n19102), .Z(n19100) );
  ANDN U21069 ( .B(n19103), .A(n19104), .Z(n19101) );
  XNOR U21070 ( .A(n19105), .B(n19106), .Z(n19103) );
  IV U21071 ( .A(n19081), .Z(n19099) );
  XOR U21072 ( .A(n19107), .B(n19108), .Z(n19081) );
  ANDN U21073 ( .B(n19109), .A(n19110), .Z(n19107) );
  XOR U21074 ( .A(n19108), .B(n19111), .Z(n19109) );
  XOR U21075 ( .A(n19090), .B(n19021), .Z(n19091) );
  XOR U21076 ( .A(n19112), .B(n19113), .Z(n19021) );
  AND U21077 ( .A(n318), .B(n19114), .Z(n19112) );
  XOR U21078 ( .A(n19115), .B(n19113), .Z(n19114) );
  XNOR U21079 ( .A(n19116), .B(n19117), .Z(n19090) );
  NAND U21080 ( .A(n19118), .B(n19119), .Z(n19117) );
  XOR U21081 ( .A(n19120), .B(n19069), .Z(n19119) );
  XOR U21082 ( .A(n19110), .B(n19111), .Z(n19069) );
  XOR U21083 ( .A(n19121), .B(n19098), .Z(n19111) );
  XOR U21084 ( .A(n19122), .B(n19123), .Z(n19098) );
  ANDN U21085 ( .B(n19124), .A(n19125), .Z(n19122) );
  XOR U21086 ( .A(n19123), .B(n19126), .Z(n19124) );
  IV U21087 ( .A(n19096), .Z(n19121) );
  XOR U21088 ( .A(n19094), .B(n19127), .Z(n19096) );
  XOR U21089 ( .A(n19128), .B(n19129), .Z(n19127) );
  ANDN U21090 ( .B(n19130), .A(n19131), .Z(n19128) );
  XOR U21091 ( .A(n19132), .B(n19129), .Z(n19130) );
  IV U21092 ( .A(n19097), .Z(n19094) );
  XOR U21093 ( .A(n19133), .B(n19134), .Z(n19097) );
  ANDN U21094 ( .B(n19135), .A(n19136), .Z(n19133) );
  XOR U21095 ( .A(n19134), .B(n19137), .Z(n19135) );
  XOR U21096 ( .A(n19138), .B(n19139), .Z(n19110) );
  XNOR U21097 ( .A(n19105), .B(n19140), .Z(n19139) );
  IV U21098 ( .A(n19108), .Z(n19140) );
  XOR U21099 ( .A(n19141), .B(n19142), .Z(n19108) );
  ANDN U21100 ( .B(n19143), .A(n19144), .Z(n19141) );
  XOR U21101 ( .A(n19142), .B(n19145), .Z(n19143) );
  XNOR U21102 ( .A(n19146), .B(n19147), .Z(n19105) );
  ANDN U21103 ( .B(n19148), .A(n19149), .Z(n19146) );
  XOR U21104 ( .A(n19147), .B(n19150), .Z(n19148) );
  IV U21105 ( .A(n19104), .Z(n19138) );
  XOR U21106 ( .A(n19102), .B(n19151), .Z(n19104) );
  XOR U21107 ( .A(n19152), .B(n19153), .Z(n19151) );
  ANDN U21108 ( .B(n19154), .A(n19155), .Z(n19152) );
  XOR U21109 ( .A(n19156), .B(n19153), .Z(n19154) );
  IV U21110 ( .A(n19106), .Z(n19102) );
  XOR U21111 ( .A(n19157), .B(n19158), .Z(n19106) );
  ANDN U21112 ( .B(n19159), .A(n19160), .Z(n19157) );
  XOR U21113 ( .A(n19161), .B(n19158), .Z(n19159) );
  IV U21114 ( .A(n19116), .Z(n19120) );
  XOR U21115 ( .A(n19116), .B(n19071), .Z(n19118) );
  XOR U21116 ( .A(n19162), .B(n19163), .Z(n19071) );
  AND U21117 ( .A(n318), .B(n19164), .Z(n19162) );
  XOR U21118 ( .A(n19165), .B(n19163), .Z(n19164) );
  NANDN U21119 ( .A(n19073), .B(n19075), .Z(n19116) );
  XOR U21120 ( .A(n19166), .B(n19167), .Z(n19075) );
  AND U21121 ( .A(n318), .B(n19168), .Z(n19166) );
  XOR U21122 ( .A(n19167), .B(n19169), .Z(n19168) );
  XNOR U21123 ( .A(n19170), .B(n19171), .Z(n318) );
  AND U21124 ( .A(n19172), .B(n19173), .Z(n19170) );
  XOR U21125 ( .A(n19171), .B(n19086), .Z(n19173) );
  XNOR U21126 ( .A(n19174), .B(n19175), .Z(n19086) );
  ANDN U21127 ( .B(n19176), .A(n19177), .Z(n19174) );
  XOR U21128 ( .A(n19175), .B(n19178), .Z(n19176) );
  XNOR U21129 ( .A(n19171), .B(n19088), .Z(n19172) );
  XOR U21130 ( .A(n19179), .B(n19180), .Z(n19088) );
  AND U21131 ( .A(n322), .B(n19181), .Z(n19179) );
  XOR U21132 ( .A(n19182), .B(n19180), .Z(n19181) );
  XNOR U21133 ( .A(n19183), .B(n19184), .Z(n19171) );
  AND U21134 ( .A(n19185), .B(n19186), .Z(n19183) );
  XNOR U21135 ( .A(n19184), .B(n19113), .Z(n19186) );
  XOR U21136 ( .A(n19177), .B(n19178), .Z(n19113) );
  XNOR U21137 ( .A(n19187), .B(n19188), .Z(n19178) );
  ANDN U21138 ( .B(n19189), .A(n19190), .Z(n19187) );
  XOR U21139 ( .A(n19191), .B(n19192), .Z(n19189) );
  XOR U21140 ( .A(n19193), .B(n19194), .Z(n19177) );
  XNOR U21141 ( .A(n19195), .B(n19196), .Z(n19194) );
  ANDN U21142 ( .B(n19197), .A(n19198), .Z(n19195) );
  XNOR U21143 ( .A(n19199), .B(n19200), .Z(n19197) );
  IV U21144 ( .A(n19175), .Z(n19193) );
  XOR U21145 ( .A(n19201), .B(n19202), .Z(n19175) );
  ANDN U21146 ( .B(n19203), .A(n19204), .Z(n19201) );
  XOR U21147 ( .A(n19202), .B(n19205), .Z(n19203) );
  XOR U21148 ( .A(n19184), .B(n19115), .Z(n19185) );
  XOR U21149 ( .A(n19206), .B(n19207), .Z(n19115) );
  AND U21150 ( .A(n322), .B(n19208), .Z(n19206) );
  XOR U21151 ( .A(n19209), .B(n19207), .Z(n19208) );
  XNOR U21152 ( .A(n19210), .B(n19211), .Z(n19184) );
  NAND U21153 ( .A(n19212), .B(n19213), .Z(n19211) );
  XOR U21154 ( .A(n19214), .B(n19163), .Z(n19213) );
  XOR U21155 ( .A(n19204), .B(n19205), .Z(n19163) );
  XOR U21156 ( .A(n19215), .B(n19192), .Z(n19205) );
  XOR U21157 ( .A(n19216), .B(n19217), .Z(n19192) );
  ANDN U21158 ( .B(n19218), .A(n19219), .Z(n19216) );
  XOR U21159 ( .A(n19217), .B(n19220), .Z(n19218) );
  IV U21160 ( .A(n19190), .Z(n19215) );
  XOR U21161 ( .A(n19188), .B(n19221), .Z(n19190) );
  XOR U21162 ( .A(n19222), .B(n19223), .Z(n19221) );
  ANDN U21163 ( .B(n19224), .A(n19225), .Z(n19222) );
  XOR U21164 ( .A(n19226), .B(n19223), .Z(n19224) );
  IV U21165 ( .A(n19191), .Z(n19188) );
  XOR U21166 ( .A(n19227), .B(n19228), .Z(n19191) );
  ANDN U21167 ( .B(n19229), .A(n19230), .Z(n19227) );
  XOR U21168 ( .A(n19228), .B(n19231), .Z(n19229) );
  XOR U21169 ( .A(n19232), .B(n19233), .Z(n19204) );
  XNOR U21170 ( .A(n19199), .B(n19234), .Z(n19233) );
  IV U21171 ( .A(n19202), .Z(n19234) );
  XOR U21172 ( .A(n19235), .B(n19236), .Z(n19202) );
  ANDN U21173 ( .B(n19237), .A(n19238), .Z(n19235) );
  XOR U21174 ( .A(n19236), .B(n19239), .Z(n19237) );
  XNOR U21175 ( .A(n19240), .B(n19241), .Z(n19199) );
  ANDN U21176 ( .B(n19242), .A(n19243), .Z(n19240) );
  XOR U21177 ( .A(n19241), .B(n19244), .Z(n19242) );
  IV U21178 ( .A(n19198), .Z(n19232) );
  XOR U21179 ( .A(n19196), .B(n19245), .Z(n19198) );
  XOR U21180 ( .A(n19246), .B(n19247), .Z(n19245) );
  ANDN U21181 ( .B(n19248), .A(n19249), .Z(n19246) );
  XOR U21182 ( .A(n19250), .B(n19247), .Z(n19248) );
  IV U21183 ( .A(n19200), .Z(n19196) );
  XOR U21184 ( .A(n19251), .B(n19252), .Z(n19200) );
  ANDN U21185 ( .B(n19253), .A(n19254), .Z(n19251) );
  XOR U21186 ( .A(n19255), .B(n19252), .Z(n19253) );
  IV U21187 ( .A(n19210), .Z(n19214) );
  XOR U21188 ( .A(n19210), .B(n19165), .Z(n19212) );
  XOR U21189 ( .A(n19256), .B(n19257), .Z(n19165) );
  AND U21190 ( .A(n322), .B(n19258), .Z(n19256) );
  XOR U21191 ( .A(n19259), .B(n19257), .Z(n19258) );
  NANDN U21192 ( .A(n19167), .B(n19169), .Z(n19210) );
  XOR U21193 ( .A(n19260), .B(n19261), .Z(n19169) );
  AND U21194 ( .A(n322), .B(n19262), .Z(n19260) );
  XOR U21195 ( .A(n19261), .B(n19263), .Z(n19262) );
  XNOR U21196 ( .A(n19264), .B(n19265), .Z(n322) );
  AND U21197 ( .A(n19266), .B(n19267), .Z(n19264) );
  XOR U21198 ( .A(n19265), .B(n19180), .Z(n19267) );
  XNOR U21199 ( .A(n19268), .B(n19269), .Z(n19180) );
  ANDN U21200 ( .B(n19270), .A(n19271), .Z(n19268) );
  XOR U21201 ( .A(n19269), .B(n19272), .Z(n19270) );
  XNOR U21202 ( .A(n19265), .B(n19182), .Z(n19266) );
  XOR U21203 ( .A(n19273), .B(n19274), .Z(n19182) );
  AND U21204 ( .A(n326), .B(n19275), .Z(n19273) );
  XOR U21205 ( .A(n19276), .B(n19274), .Z(n19275) );
  XNOR U21206 ( .A(n19277), .B(n19278), .Z(n19265) );
  AND U21207 ( .A(n19279), .B(n19280), .Z(n19277) );
  XNOR U21208 ( .A(n19278), .B(n19207), .Z(n19280) );
  XOR U21209 ( .A(n19271), .B(n19272), .Z(n19207) );
  XNOR U21210 ( .A(n19281), .B(n19282), .Z(n19272) );
  ANDN U21211 ( .B(n19283), .A(n19284), .Z(n19281) );
  XOR U21212 ( .A(n19285), .B(n19286), .Z(n19283) );
  XOR U21213 ( .A(n19287), .B(n19288), .Z(n19271) );
  XNOR U21214 ( .A(n19289), .B(n19290), .Z(n19288) );
  ANDN U21215 ( .B(n19291), .A(n19292), .Z(n19289) );
  XNOR U21216 ( .A(n19293), .B(n19294), .Z(n19291) );
  IV U21217 ( .A(n19269), .Z(n19287) );
  XOR U21218 ( .A(n19295), .B(n19296), .Z(n19269) );
  ANDN U21219 ( .B(n19297), .A(n19298), .Z(n19295) );
  XOR U21220 ( .A(n19296), .B(n19299), .Z(n19297) );
  XOR U21221 ( .A(n19278), .B(n19209), .Z(n19279) );
  XOR U21222 ( .A(n19300), .B(n19301), .Z(n19209) );
  AND U21223 ( .A(n326), .B(n19302), .Z(n19300) );
  XOR U21224 ( .A(n19303), .B(n19301), .Z(n19302) );
  XNOR U21225 ( .A(n19304), .B(n19305), .Z(n19278) );
  NAND U21226 ( .A(n19306), .B(n19307), .Z(n19305) );
  XOR U21227 ( .A(n19308), .B(n19257), .Z(n19307) );
  XOR U21228 ( .A(n19298), .B(n19299), .Z(n19257) );
  XOR U21229 ( .A(n19309), .B(n19286), .Z(n19299) );
  XOR U21230 ( .A(n19310), .B(n19311), .Z(n19286) );
  ANDN U21231 ( .B(n19312), .A(n19313), .Z(n19310) );
  XOR U21232 ( .A(n19311), .B(n19314), .Z(n19312) );
  IV U21233 ( .A(n19284), .Z(n19309) );
  XOR U21234 ( .A(n19282), .B(n19315), .Z(n19284) );
  XOR U21235 ( .A(n19316), .B(n19317), .Z(n19315) );
  ANDN U21236 ( .B(n19318), .A(n19319), .Z(n19316) );
  XOR U21237 ( .A(n19320), .B(n19317), .Z(n19318) );
  IV U21238 ( .A(n19285), .Z(n19282) );
  XOR U21239 ( .A(n19321), .B(n19322), .Z(n19285) );
  ANDN U21240 ( .B(n19323), .A(n19324), .Z(n19321) );
  XOR U21241 ( .A(n19322), .B(n19325), .Z(n19323) );
  XOR U21242 ( .A(n19326), .B(n19327), .Z(n19298) );
  XNOR U21243 ( .A(n19293), .B(n19328), .Z(n19327) );
  IV U21244 ( .A(n19296), .Z(n19328) );
  XOR U21245 ( .A(n19329), .B(n19330), .Z(n19296) );
  ANDN U21246 ( .B(n19331), .A(n19332), .Z(n19329) );
  XOR U21247 ( .A(n19330), .B(n19333), .Z(n19331) );
  XNOR U21248 ( .A(n19334), .B(n19335), .Z(n19293) );
  ANDN U21249 ( .B(n19336), .A(n19337), .Z(n19334) );
  XOR U21250 ( .A(n19335), .B(n19338), .Z(n19336) );
  IV U21251 ( .A(n19292), .Z(n19326) );
  XOR U21252 ( .A(n19290), .B(n19339), .Z(n19292) );
  XOR U21253 ( .A(n19340), .B(n19341), .Z(n19339) );
  ANDN U21254 ( .B(n19342), .A(n19343), .Z(n19340) );
  XOR U21255 ( .A(n19344), .B(n19341), .Z(n19342) );
  IV U21256 ( .A(n19294), .Z(n19290) );
  XOR U21257 ( .A(n19345), .B(n19346), .Z(n19294) );
  ANDN U21258 ( .B(n19347), .A(n19348), .Z(n19345) );
  XOR U21259 ( .A(n19349), .B(n19346), .Z(n19347) );
  IV U21260 ( .A(n19304), .Z(n19308) );
  XOR U21261 ( .A(n19304), .B(n19259), .Z(n19306) );
  XOR U21262 ( .A(n19350), .B(n19351), .Z(n19259) );
  AND U21263 ( .A(n326), .B(n19352), .Z(n19350) );
  XOR U21264 ( .A(n19353), .B(n19351), .Z(n19352) );
  NANDN U21265 ( .A(n19261), .B(n19263), .Z(n19304) );
  XOR U21266 ( .A(n19354), .B(n19355), .Z(n19263) );
  AND U21267 ( .A(n326), .B(n19356), .Z(n19354) );
  XOR U21268 ( .A(n19355), .B(n19357), .Z(n19356) );
  XNOR U21269 ( .A(n19358), .B(n19359), .Z(n326) );
  AND U21270 ( .A(n19360), .B(n19361), .Z(n19358) );
  XOR U21271 ( .A(n19359), .B(n19274), .Z(n19361) );
  XNOR U21272 ( .A(n19362), .B(n19363), .Z(n19274) );
  ANDN U21273 ( .B(n19364), .A(n19365), .Z(n19362) );
  XOR U21274 ( .A(n19363), .B(n19366), .Z(n19364) );
  XNOR U21275 ( .A(n19359), .B(n19276), .Z(n19360) );
  XOR U21276 ( .A(n19367), .B(n19368), .Z(n19276) );
  AND U21277 ( .A(n330), .B(n19369), .Z(n19367) );
  XOR U21278 ( .A(n19370), .B(n19368), .Z(n19369) );
  XNOR U21279 ( .A(n19371), .B(n19372), .Z(n19359) );
  AND U21280 ( .A(n19373), .B(n19374), .Z(n19371) );
  XNOR U21281 ( .A(n19372), .B(n19301), .Z(n19374) );
  XOR U21282 ( .A(n19365), .B(n19366), .Z(n19301) );
  XNOR U21283 ( .A(n19375), .B(n19376), .Z(n19366) );
  ANDN U21284 ( .B(n19377), .A(n19378), .Z(n19375) );
  XOR U21285 ( .A(n19379), .B(n19380), .Z(n19377) );
  XOR U21286 ( .A(n19381), .B(n19382), .Z(n19365) );
  XNOR U21287 ( .A(n19383), .B(n19384), .Z(n19382) );
  ANDN U21288 ( .B(n19385), .A(n19386), .Z(n19383) );
  XNOR U21289 ( .A(n19387), .B(n19388), .Z(n19385) );
  IV U21290 ( .A(n19363), .Z(n19381) );
  XOR U21291 ( .A(n19389), .B(n19390), .Z(n19363) );
  ANDN U21292 ( .B(n19391), .A(n19392), .Z(n19389) );
  XOR U21293 ( .A(n19390), .B(n19393), .Z(n19391) );
  XOR U21294 ( .A(n19372), .B(n19303), .Z(n19373) );
  XOR U21295 ( .A(n19394), .B(n19395), .Z(n19303) );
  AND U21296 ( .A(n330), .B(n19396), .Z(n19394) );
  XOR U21297 ( .A(n19397), .B(n19395), .Z(n19396) );
  XNOR U21298 ( .A(n19398), .B(n19399), .Z(n19372) );
  NAND U21299 ( .A(n19400), .B(n19401), .Z(n19399) );
  XOR U21300 ( .A(n19402), .B(n19351), .Z(n19401) );
  XOR U21301 ( .A(n19392), .B(n19393), .Z(n19351) );
  XOR U21302 ( .A(n19403), .B(n19380), .Z(n19393) );
  XOR U21303 ( .A(n19404), .B(n19405), .Z(n19380) );
  ANDN U21304 ( .B(n19406), .A(n19407), .Z(n19404) );
  XOR U21305 ( .A(n19405), .B(n19408), .Z(n19406) );
  IV U21306 ( .A(n19378), .Z(n19403) );
  XOR U21307 ( .A(n19376), .B(n19409), .Z(n19378) );
  XOR U21308 ( .A(n19410), .B(n19411), .Z(n19409) );
  ANDN U21309 ( .B(n19412), .A(n19413), .Z(n19410) );
  XOR U21310 ( .A(n19414), .B(n19411), .Z(n19412) );
  IV U21311 ( .A(n19379), .Z(n19376) );
  XOR U21312 ( .A(n19415), .B(n19416), .Z(n19379) );
  ANDN U21313 ( .B(n19417), .A(n19418), .Z(n19415) );
  XOR U21314 ( .A(n19416), .B(n19419), .Z(n19417) );
  XOR U21315 ( .A(n19420), .B(n19421), .Z(n19392) );
  XNOR U21316 ( .A(n19387), .B(n19422), .Z(n19421) );
  IV U21317 ( .A(n19390), .Z(n19422) );
  XOR U21318 ( .A(n19423), .B(n19424), .Z(n19390) );
  ANDN U21319 ( .B(n19425), .A(n19426), .Z(n19423) );
  XOR U21320 ( .A(n19424), .B(n19427), .Z(n19425) );
  XNOR U21321 ( .A(n19428), .B(n19429), .Z(n19387) );
  ANDN U21322 ( .B(n19430), .A(n19431), .Z(n19428) );
  XOR U21323 ( .A(n19429), .B(n19432), .Z(n19430) );
  IV U21324 ( .A(n19386), .Z(n19420) );
  XOR U21325 ( .A(n19384), .B(n19433), .Z(n19386) );
  XOR U21326 ( .A(n19434), .B(n19435), .Z(n19433) );
  ANDN U21327 ( .B(n19436), .A(n19437), .Z(n19434) );
  XOR U21328 ( .A(n19438), .B(n19435), .Z(n19436) );
  IV U21329 ( .A(n19388), .Z(n19384) );
  XOR U21330 ( .A(n19439), .B(n19440), .Z(n19388) );
  ANDN U21331 ( .B(n19441), .A(n19442), .Z(n19439) );
  XOR U21332 ( .A(n19443), .B(n19440), .Z(n19441) );
  IV U21333 ( .A(n19398), .Z(n19402) );
  XOR U21334 ( .A(n19398), .B(n19353), .Z(n19400) );
  XOR U21335 ( .A(n19444), .B(n19445), .Z(n19353) );
  AND U21336 ( .A(n330), .B(n19446), .Z(n19444) );
  XOR U21337 ( .A(n19447), .B(n19445), .Z(n19446) );
  NANDN U21338 ( .A(n19355), .B(n19357), .Z(n19398) );
  XOR U21339 ( .A(n19448), .B(n19449), .Z(n19357) );
  AND U21340 ( .A(n330), .B(n19450), .Z(n19448) );
  XOR U21341 ( .A(n19449), .B(n19451), .Z(n19450) );
  XNOR U21342 ( .A(n19452), .B(n19453), .Z(n330) );
  AND U21343 ( .A(n19454), .B(n19455), .Z(n19452) );
  XOR U21344 ( .A(n19453), .B(n19368), .Z(n19455) );
  XNOR U21345 ( .A(n19456), .B(n19457), .Z(n19368) );
  ANDN U21346 ( .B(n19458), .A(n19459), .Z(n19456) );
  XOR U21347 ( .A(n19457), .B(n19460), .Z(n19458) );
  XNOR U21348 ( .A(n19453), .B(n19370), .Z(n19454) );
  XOR U21349 ( .A(n19461), .B(n19462), .Z(n19370) );
  AND U21350 ( .A(n334), .B(n19463), .Z(n19461) );
  XOR U21351 ( .A(n19464), .B(n19462), .Z(n19463) );
  XNOR U21352 ( .A(n19465), .B(n19466), .Z(n19453) );
  AND U21353 ( .A(n19467), .B(n19468), .Z(n19465) );
  XNOR U21354 ( .A(n19466), .B(n19395), .Z(n19468) );
  XOR U21355 ( .A(n19459), .B(n19460), .Z(n19395) );
  XNOR U21356 ( .A(n19469), .B(n19470), .Z(n19460) );
  ANDN U21357 ( .B(n19471), .A(n19472), .Z(n19469) );
  XOR U21358 ( .A(n19473), .B(n19474), .Z(n19471) );
  XOR U21359 ( .A(n19475), .B(n19476), .Z(n19459) );
  XNOR U21360 ( .A(n19477), .B(n19478), .Z(n19476) );
  ANDN U21361 ( .B(n19479), .A(n19480), .Z(n19477) );
  XNOR U21362 ( .A(n19481), .B(n19482), .Z(n19479) );
  IV U21363 ( .A(n19457), .Z(n19475) );
  XOR U21364 ( .A(n19483), .B(n19484), .Z(n19457) );
  ANDN U21365 ( .B(n19485), .A(n19486), .Z(n19483) );
  XOR U21366 ( .A(n19484), .B(n19487), .Z(n19485) );
  XOR U21367 ( .A(n19466), .B(n19397), .Z(n19467) );
  XOR U21368 ( .A(n19488), .B(n19489), .Z(n19397) );
  AND U21369 ( .A(n334), .B(n19490), .Z(n19488) );
  XOR U21370 ( .A(n19491), .B(n19489), .Z(n19490) );
  XNOR U21371 ( .A(n19492), .B(n19493), .Z(n19466) );
  NAND U21372 ( .A(n19494), .B(n19495), .Z(n19493) );
  XOR U21373 ( .A(n19496), .B(n19445), .Z(n19495) );
  XOR U21374 ( .A(n19486), .B(n19487), .Z(n19445) );
  XOR U21375 ( .A(n19497), .B(n19474), .Z(n19487) );
  XOR U21376 ( .A(n19498), .B(n19499), .Z(n19474) );
  ANDN U21377 ( .B(n19500), .A(n19501), .Z(n19498) );
  XOR U21378 ( .A(n19499), .B(n19502), .Z(n19500) );
  IV U21379 ( .A(n19472), .Z(n19497) );
  XOR U21380 ( .A(n19470), .B(n19503), .Z(n19472) );
  XOR U21381 ( .A(n19504), .B(n19505), .Z(n19503) );
  ANDN U21382 ( .B(n19506), .A(n19507), .Z(n19504) );
  XOR U21383 ( .A(n19508), .B(n19505), .Z(n19506) );
  IV U21384 ( .A(n19473), .Z(n19470) );
  XOR U21385 ( .A(n19509), .B(n19510), .Z(n19473) );
  ANDN U21386 ( .B(n19511), .A(n19512), .Z(n19509) );
  XOR U21387 ( .A(n19510), .B(n19513), .Z(n19511) );
  XOR U21388 ( .A(n19514), .B(n19515), .Z(n19486) );
  XNOR U21389 ( .A(n19481), .B(n19516), .Z(n19515) );
  IV U21390 ( .A(n19484), .Z(n19516) );
  XOR U21391 ( .A(n19517), .B(n19518), .Z(n19484) );
  ANDN U21392 ( .B(n19519), .A(n19520), .Z(n19517) );
  XOR U21393 ( .A(n19518), .B(n19521), .Z(n19519) );
  XNOR U21394 ( .A(n19522), .B(n19523), .Z(n19481) );
  ANDN U21395 ( .B(n19524), .A(n19525), .Z(n19522) );
  XOR U21396 ( .A(n19523), .B(n19526), .Z(n19524) );
  IV U21397 ( .A(n19480), .Z(n19514) );
  XOR U21398 ( .A(n19478), .B(n19527), .Z(n19480) );
  XOR U21399 ( .A(n19528), .B(n19529), .Z(n19527) );
  ANDN U21400 ( .B(n19530), .A(n19531), .Z(n19528) );
  XOR U21401 ( .A(n19532), .B(n19529), .Z(n19530) );
  IV U21402 ( .A(n19482), .Z(n19478) );
  XOR U21403 ( .A(n19533), .B(n19534), .Z(n19482) );
  ANDN U21404 ( .B(n19535), .A(n19536), .Z(n19533) );
  XOR U21405 ( .A(n19537), .B(n19534), .Z(n19535) );
  IV U21406 ( .A(n19492), .Z(n19496) );
  XOR U21407 ( .A(n19492), .B(n19447), .Z(n19494) );
  XOR U21408 ( .A(n19538), .B(n19539), .Z(n19447) );
  AND U21409 ( .A(n334), .B(n19540), .Z(n19538) );
  XOR U21410 ( .A(n19541), .B(n19539), .Z(n19540) );
  NANDN U21411 ( .A(n19449), .B(n19451), .Z(n19492) );
  XOR U21412 ( .A(n19542), .B(n19543), .Z(n19451) );
  AND U21413 ( .A(n334), .B(n19544), .Z(n19542) );
  XOR U21414 ( .A(n19543), .B(n19545), .Z(n19544) );
  XNOR U21415 ( .A(n19546), .B(n19547), .Z(n334) );
  AND U21416 ( .A(n19548), .B(n19549), .Z(n19546) );
  XOR U21417 ( .A(n19547), .B(n19462), .Z(n19549) );
  XNOR U21418 ( .A(n19550), .B(n19551), .Z(n19462) );
  ANDN U21419 ( .B(n19552), .A(n19553), .Z(n19550) );
  XOR U21420 ( .A(n19551), .B(n19554), .Z(n19552) );
  XNOR U21421 ( .A(n19547), .B(n19464), .Z(n19548) );
  XOR U21422 ( .A(n19555), .B(n19556), .Z(n19464) );
  AND U21423 ( .A(n338), .B(n19557), .Z(n19555) );
  XOR U21424 ( .A(n19558), .B(n19556), .Z(n19557) );
  XNOR U21425 ( .A(n19559), .B(n19560), .Z(n19547) );
  AND U21426 ( .A(n19561), .B(n19562), .Z(n19559) );
  XNOR U21427 ( .A(n19560), .B(n19489), .Z(n19562) );
  XOR U21428 ( .A(n19553), .B(n19554), .Z(n19489) );
  XNOR U21429 ( .A(n19563), .B(n19564), .Z(n19554) );
  ANDN U21430 ( .B(n19565), .A(n19566), .Z(n19563) );
  XOR U21431 ( .A(n19567), .B(n19568), .Z(n19565) );
  XOR U21432 ( .A(n19569), .B(n19570), .Z(n19553) );
  XNOR U21433 ( .A(n19571), .B(n19572), .Z(n19570) );
  ANDN U21434 ( .B(n19573), .A(n19574), .Z(n19571) );
  XNOR U21435 ( .A(n19575), .B(n19576), .Z(n19573) );
  IV U21436 ( .A(n19551), .Z(n19569) );
  XOR U21437 ( .A(n19577), .B(n19578), .Z(n19551) );
  ANDN U21438 ( .B(n19579), .A(n19580), .Z(n19577) );
  XOR U21439 ( .A(n19578), .B(n19581), .Z(n19579) );
  XOR U21440 ( .A(n19560), .B(n19491), .Z(n19561) );
  XOR U21441 ( .A(n19582), .B(n19583), .Z(n19491) );
  AND U21442 ( .A(n338), .B(n19584), .Z(n19582) );
  XOR U21443 ( .A(n19585), .B(n19583), .Z(n19584) );
  XNOR U21444 ( .A(n19586), .B(n19587), .Z(n19560) );
  NAND U21445 ( .A(n19588), .B(n19589), .Z(n19587) );
  XOR U21446 ( .A(n19590), .B(n19539), .Z(n19589) );
  XOR U21447 ( .A(n19580), .B(n19581), .Z(n19539) );
  XOR U21448 ( .A(n19591), .B(n19568), .Z(n19581) );
  XOR U21449 ( .A(n19592), .B(n19593), .Z(n19568) );
  ANDN U21450 ( .B(n19594), .A(n19595), .Z(n19592) );
  XOR U21451 ( .A(n19593), .B(n19596), .Z(n19594) );
  IV U21452 ( .A(n19566), .Z(n19591) );
  XOR U21453 ( .A(n19564), .B(n19597), .Z(n19566) );
  XOR U21454 ( .A(n19598), .B(n19599), .Z(n19597) );
  ANDN U21455 ( .B(n19600), .A(n19601), .Z(n19598) );
  XOR U21456 ( .A(n19602), .B(n19599), .Z(n19600) );
  IV U21457 ( .A(n19567), .Z(n19564) );
  XOR U21458 ( .A(n19603), .B(n19604), .Z(n19567) );
  ANDN U21459 ( .B(n19605), .A(n19606), .Z(n19603) );
  XOR U21460 ( .A(n19604), .B(n19607), .Z(n19605) );
  XOR U21461 ( .A(n19608), .B(n19609), .Z(n19580) );
  XNOR U21462 ( .A(n19575), .B(n19610), .Z(n19609) );
  IV U21463 ( .A(n19578), .Z(n19610) );
  XOR U21464 ( .A(n19611), .B(n19612), .Z(n19578) );
  ANDN U21465 ( .B(n19613), .A(n19614), .Z(n19611) );
  XOR U21466 ( .A(n19612), .B(n19615), .Z(n19613) );
  XNOR U21467 ( .A(n19616), .B(n19617), .Z(n19575) );
  ANDN U21468 ( .B(n19618), .A(n19619), .Z(n19616) );
  XOR U21469 ( .A(n19617), .B(n19620), .Z(n19618) );
  IV U21470 ( .A(n19574), .Z(n19608) );
  XOR U21471 ( .A(n19572), .B(n19621), .Z(n19574) );
  XOR U21472 ( .A(n19622), .B(n19623), .Z(n19621) );
  ANDN U21473 ( .B(n19624), .A(n19625), .Z(n19622) );
  XOR U21474 ( .A(n19626), .B(n19623), .Z(n19624) );
  IV U21475 ( .A(n19576), .Z(n19572) );
  XOR U21476 ( .A(n19627), .B(n19628), .Z(n19576) );
  ANDN U21477 ( .B(n19629), .A(n19630), .Z(n19627) );
  XOR U21478 ( .A(n19631), .B(n19628), .Z(n19629) );
  IV U21479 ( .A(n19586), .Z(n19590) );
  XOR U21480 ( .A(n19586), .B(n19541), .Z(n19588) );
  XOR U21481 ( .A(n19632), .B(n19633), .Z(n19541) );
  AND U21482 ( .A(n338), .B(n19634), .Z(n19632) );
  XOR U21483 ( .A(n19635), .B(n19633), .Z(n19634) );
  NANDN U21484 ( .A(n19543), .B(n19545), .Z(n19586) );
  XOR U21485 ( .A(n19636), .B(n19637), .Z(n19545) );
  AND U21486 ( .A(n338), .B(n19638), .Z(n19636) );
  XOR U21487 ( .A(n19637), .B(n19639), .Z(n19638) );
  XNOR U21488 ( .A(n19640), .B(n19641), .Z(n338) );
  AND U21489 ( .A(n19642), .B(n19643), .Z(n19640) );
  XOR U21490 ( .A(n19641), .B(n19556), .Z(n19643) );
  XNOR U21491 ( .A(n19644), .B(n19645), .Z(n19556) );
  ANDN U21492 ( .B(n19646), .A(n19647), .Z(n19644) );
  XOR U21493 ( .A(n19645), .B(n19648), .Z(n19646) );
  XNOR U21494 ( .A(n19641), .B(n19558), .Z(n19642) );
  XOR U21495 ( .A(n19649), .B(n19650), .Z(n19558) );
  AND U21496 ( .A(n342), .B(n19651), .Z(n19649) );
  XOR U21497 ( .A(n19652), .B(n19650), .Z(n19651) );
  XNOR U21498 ( .A(n19653), .B(n19654), .Z(n19641) );
  AND U21499 ( .A(n19655), .B(n19656), .Z(n19653) );
  XNOR U21500 ( .A(n19654), .B(n19583), .Z(n19656) );
  XOR U21501 ( .A(n19647), .B(n19648), .Z(n19583) );
  XNOR U21502 ( .A(n19657), .B(n19658), .Z(n19648) );
  ANDN U21503 ( .B(n19659), .A(n19660), .Z(n19657) );
  XOR U21504 ( .A(n19661), .B(n19662), .Z(n19659) );
  XOR U21505 ( .A(n19663), .B(n19664), .Z(n19647) );
  XNOR U21506 ( .A(n19665), .B(n19666), .Z(n19664) );
  ANDN U21507 ( .B(n19667), .A(n19668), .Z(n19665) );
  XNOR U21508 ( .A(n19669), .B(n19670), .Z(n19667) );
  IV U21509 ( .A(n19645), .Z(n19663) );
  XOR U21510 ( .A(n19671), .B(n19672), .Z(n19645) );
  ANDN U21511 ( .B(n19673), .A(n19674), .Z(n19671) );
  XOR U21512 ( .A(n19672), .B(n19675), .Z(n19673) );
  XOR U21513 ( .A(n19654), .B(n19585), .Z(n19655) );
  XOR U21514 ( .A(n19676), .B(n19677), .Z(n19585) );
  AND U21515 ( .A(n342), .B(n19678), .Z(n19676) );
  XOR U21516 ( .A(n19679), .B(n19677), .Z(n19678) );
  XNOR U21517 ( .A(n19680), .B(n19681), .Z(n19654) );
  NAND U21518 ( .A(n19682), .B(n19683), .Z(n19681) );
  XOR U21519 ( .A(n19684), .B(n19633), .Z(n19683) );
  XOR U21520 ( .A(n19674), .B(n19675), .Z(n19633) );
  XOR U21521 ( .A(n19685), .B(n19662), .Z(n19675) );
  XOR U21522 ( .A(n19686), .B(n19687), .Z(n19662) );
  ANDN U21523 ( .B(n19688), .A(n19689), .Z(n19686) );
  XOR U21524 ( .A(n19687), .B(n19690), .Z(n19688) );
  IV U21525 ( .A(n19660), .Z(n19685) );
  XOR U21526 ( .A(n19658), .B(n19691), .Z(n19660) );
  XOR U21527 ( .A(n19692), .B(n19693), .Z(n19691) );
  ANDN U21528 ( .B(n19694), .A(n19695), .Z(n19692) );
  XOR U21529 ( .A(n19696), .B(n19693), .Z(n19694) );
  IV U21530 ( .A(n19661), .Z(n19658) );
  XOR U21531 ( .A(n19697), .B(n19698), .Z(n19661) );
  ANDN U21532 ( .B(n19699), .A(n19700), .Z(n19697) );
  XOR U21533 ( .A(n19698), .B(n19701), .Z(n19699) );
  XOR U21534 ( .A(n19702), .B(n19703), .Z(n19674) );
  XNOR U21535 ( .A(n19669), .B(n19704), .Z(n19703) );
  IV U21536 ( .A(n19672), .Z(n19704) );
  XOR U21537 ( .A(n19705), .B(n19706), .Z(n19672) );
  ANDN U21538 ( .B(n19707), .A(n19708), .Z(n19705) );
  XOR U21539 ( .A(n19706), .B(n19709), .Z(n19707) );
  XNOR U21540 ( .A(n19710), .B(n19711), .Z(n19669) );
  ANDN U21541 ( .B(n19712), .A(n19713), .Z(n19710) );
  XOR U21542 ( .A(n19711), .B(n19714), .Z(n19712) );
  IV U21543 ( .A(n19668), .Z(n19702) );
  XOR U21544 ( .A(n19666), .B(n19715), .Z(n19668) );
  XOR U21545 ( .A(n19716), .B(n19717), .Z(n19715) );
  ANDN U21546 ( .B(n19718), .A(n19719), .Z(n19716) );
  XOR U21547 ( .A(n19720), .B(n19717), .Z(n19718) );
  IV U21548 ( .A(n19670), .Z(n19666) );
  XOR U21549 ( .A(n19721), .B(n19722), .Z(n19670) );
  ANDN U21550 ( .B(n19723), .A(n19724), .Z(n19721) );
  XOR U21551 ( .A(n19725), .B(n19722), .Z(n19723) );
  IV U21552 ( .A(n19680), .Z(n19684) );
  XOR U21553 ( .A(n19680), .B(n19635), .Z(n19682) );
  XOR U21554 ( .A(n19726), .B(n19727), .Z(n19635) );
  AND U21555 ( .A(n342), .B(n19728), .Z(n19726) );
  XOR U21556 ( .A(n19729), .B(n19727), .Z(n19728) );
  NANDN U21557 ( .A(n19637), .B(n19639), .Z(n19680) );
  XOR U21558 ( .A(n19730), .B(n19731), .Z(n19639) );
  AND U21559 ( .A(n342), .B(n19732), .Z(n19730) );
  XOR U21560 ( .A(n19731), .B(n19733), .Z(n19732) );
  XNOR U21561 ( .A(n19734), .B(n19735), .Z(n342) );
  AND U21562 ( .A(n19736), .B(n19737), .Z(n19734) );
  XOR U21563 ( .A(n19735), .B(n19650), .Z(n19737) );
  XNOR U21564 ( .A(n19738), .B(n19739), .Z(n19650) );
  ANDN U21565 ( .B(n19740), .A(n19741), .Z(n19738) );
  XOR U21566 ( .A(n19739), .B(n19742), .Z(n19740) );
  XNOR U21567 ( .A(n19735), .B(n19652), .Z(n19736) );
  XOR U21568 ( .A(n19743), .B(n19744), .Z(n19652) );
  AND U21569 ( .A(n346), .B(n19745), .Z(n19743) );
  XOR U21570 ( .A(n19746), .B(n19744), .Z(n19745) );
  XNOR U21571 ( .A(n19747), .B(n19748), .Z(n19735) );
  AND U21572 ( .A(n19749), .B(n19750), .Z(n19747) );
  XNOR U21573 ( .A(n19748), .B(n19677), .Z(n19750) );
  XOR U21574 ( .A(n19741), .B(n19742), .Z(n19677) );
  XNOR U21575 ( .A(n19751), .B(n19752), .Z(n19742) );
  ANDN U21576 ( .B(n19753), .A(n19754), .Z(n19751) );
  XOR U21577 ( .A(n19755), .B(n19756), .Z(n19753) );
  XOR U21578 ( .A(n19757), .B(n19758), .Z(n19741) );
  XNOR U21579 ( .A(n19759), .B(n19760), .Z(n19758) );
  ANDN U21580 ( .B(n19761), .A(n19762), .Z(n19759) );
  XNOR U21581 ( .A(n19763), .B(n19764), .Z(n19761) );
  IV U21582 ( .A(n19739), .Z(n19757) );
  XOR U21583 ( .A(n19765), .B(n19766), .Z(n19739) );
  ANDN U21584 ( .B(n19767), .A(n19768), .Z(n19765) );
  XOR U21585 ( .A(n19766), .B(n19769), .Z(n19767) );
  XOR U21586 ( .A(n19748), .B(n19679), .Z(n19749) );
  XOR U21587 ( .A(n19770), .B(n19771), .Z(n19679) );
  AND U21588 ( .A(n346), .B(n19772), .Z(n19770) );
  XOR U21589 ( .A(n19773), .B(n19771), .Z(n19772) );
  XNOR U21590 ( .A(n19774), .B(n19775), .Z(n19748) );
  NAND U21591 ( .A(n19776), .B(n19777), .Z(n19775) );
  XOR U21592 ( .A(n19778), .B(n19727), .Z(n19777) );
  XOR U21593 ( .A(n19768), .B(n19769), .Z(n19727) );
  XOR U21594 ( .A(n19779), .B(n19756), .Z(n19769) );
  XOR U21595 ( .A(n19780), .B(n19781), .Z(n19756) );
  ANDN U21596 ( .B(n19782), .A(n19783), .Z(n19780) );
  XOR U21597 ( .A(n19781), .B(n19784), .Z(n19782) );
  IV U21598 ( .A(n19754), .Z(n19779) );
  XOR U21599 ( .A(n19752), .B(n19785), .Z(n19754) );
  XOR U21600 ( .A(n19786), .B(n19787), .Z(n19785) );
  ANDN U21601 ( .B(n19788), .A(n19789), .Z(n19786) );
  XOR U21602 ( .A(n19790), .B(n19787), .Z(n19788) );
  IV U21603 ( .A(n19755), .Z(n19752) );
  XOR U21604 ( .A(n19791), .B(n19792), .Z(n19755) );
  ANDN U21605 ( .B(n19793), .A(n19794), .Z(n19791) );
  XOR U21606 ( .A(n19792), .B(n19795), .Z(n19793) );
  XOR U21607 ( .A(n19796), .B(n19797), .Z(n19768) );
  XNOR U21608 ( .A(n19763), .B(n19798), .Z(n19797) );
  IV U21609 ( .A(n19766), .Z(n19798) );
  XOR U21610 ( .A(n19799), .B(n19800), .Z(n19766) );
  ANDN U21611 ( .B(n19801), .A(n19802), .Z(n19799) );
  XOR U21612 ( .A(n19800), .B(n19803), .Z(n19801) );
  XNOR U21613 ( .A(n19804), .B(n19805), .Z(n19763) );
  ANDN U21614 ( .B(n19806), .A(n19807), .Z(n19804) );
  XOR U21615 ( .A(n19805), .B(n19808), .Z(n19806) );
  IV U21616 ( .A(n19762), .Z(n19796) );
  XOR U21617 ( .A(n19760), .B(n19809), .Z(n19762) );
  XOR U21618 ( .A(n19810), .B(n19811), .Z(n19809) );
  ANDN U21619 ( .B(n19812), .A(n19813), .Z(n19810) );
  XOR U21620 ( .A(n19814), .B(n19811), .Z(n19812) );
  IV U21621 ( .A(n19764), .Z(n19760) );
  XOR U21622 ( .A(n19815), .B(n19816), .Z(n19764) );
  ANDN U21623 ( .B(n19817), .A(n19818), .Z(n19815) );
  XOR U21624 ( .A(n19819), .B(n19816), .Z(n19817) );
  IV U21625 ( .A(n19774), .Z(n19778) );
  XOR U21626 ( .A(n19774), .B(n19729), .Z(n19776) );
  XOR U21627 ( .A(n19820), .B(n19821), .Z(n19729) );
  AND U21628 ( .A(n346), .B(n19822), .Z(n19820) );
  XOR U21629 ( .A(n19823), .B(n19821), .Z(n19822) );
  NANDN U21630 ( .A(n19731), .B(n19733), .Z(n19774) );
  XOR U21631 ( .A(n19824), .B(n19825), .Z(n19733) );
  AND U21632 ( .A(n346), .B(n19826), .Z(n19824) );
  XOR U21633 ( .A(n19825), .B(n19827), .Z(n19826) );
  XNOR U21634 ( .A(n19828), .B(n19829), .Z(n346) );
  AND U21635 ( .A(n19830), .B(n19831), .Z(n19828) );
  XOR U21636 ( .A(n19829), .B(n19744), .Z(n19831) );
  XNOR U21637 ( .A(n19832), .B(n19833), .Z(n19744) );
  ANDN U21638 ( .B(n19834), .A(n19835), .Z(n19832) );
  XOR U21639 ( .A(n19833), .B(n19836), .Z(n19834) );
  XNOR U21640 ( .A(n19829), .B(n19746), .Z(n19830) );
  XOR U21641 ( .A(n19837), .B(n19838), .Z(n19746) );
  AND U21642 ( .A(n350), .B(n19839), .Z(n19837) );
  XOR U21643 ( .A(n19840), .B(n19838), .Z(n19839) );
  XNOR U21644 ( .A(n19841), .B(n19842), .Z(n19829) );
  AND U21645 ( .A(n19843), .B(n19844), .Z(n19841) );
  XNOR U21646 ( .A(n19842), .B(n19771), .Z(n19844) );
  XOR U21647 ( .A(n19835), .B(n19836), .Z(n19771) );
  XNOR U21648 ( .A(n19845), .B(n19846), .Z(n19836) );
  ANDN U21649 ( .B(n19847), .A(n19848), .Z(n19845) );
  XOR U21650 ( .A(n19849), .B(n19850), .Z(n19847) );
  XOR U21651 ( .A(n19851), .B(n19852), .Z(n19835) );
  XNOR U21652 ( .A(n19853), .B(n19854), .Z(n19852) );
  ANDN U21653 ( .B(n19855), .A(n19856), .Z(n19853) );
  XNOR U21654 ( .A(n19857), .B(n19858), .Z(n19855) );
  IV U21655 ( .A(n19833), .Z(n19851) );
  XOR U21656 ( .A(n19859), .B(n19860), .Z(n19833) );
  ANDN U21657 ( .B(n19861), .A(n19862), .Z(n19859) );
  XOR U21658 ( .A(n19860), .B(n19863), .Z(n19861) );
  XOR U21659 ( .A(n19842), .B(n19773), .Z(n19843) );
  XOR U21660 ( .A(n19864), .B(n19865), .Z(n19773) );
  AND U21661 ( .A(n350), .B(n19866), .Z(n19864) );
  XOR U21662 ( .A(n19867), .B(n19865), .Z(n19866) );
  XNOR U21663 ( .A(n19868), .B(n19869), .Z(n19842) );
  NAND U21664 ( .A(n19870), .B(n19871), .Z(n19869) );
  XOR U21665 ( .A(n19872), .B(n19821), .Z(n19871) );
  XOR U21666 ( .A(n19862), .B(n19863), .Z(n19821) );
  XOR U21667 ( .A(n19873), .B(n19850), .Z(n19863) );
  XOR U21668 ( .A(n19874), .B(n19875), .Z(n19850) );
  ANDN U21669 ( .B(n19876), .A(n19877), .Z(n19874) );
  XOR U21670 ( .A(n19875), .B(n19878), .Z(n19876) );
  IV U21671 ( .A(n19848), .Z(n19873) );
  XOR U21672 ( .A(n19846), .B(n19879), .Z(n19848) );
  XOR U21673 ( .A(n19880), .B(n19881), .Z(n19879) );
  ANDN U21674 ( .B(n19882), .A(n19883), .Z(n19880) );
  XOR U21675 ( .A(n19884), .B(n19881), .Z(n19882) );
  IV U21676 ( .A(n19849), .Z(n19846) );
  XOR U21677 ( .A(n19885), .B(n19886), .Z(n19849) );
  ANDN U21678 ( .B(n19887), .A(n19888), .Z(n19885) );
  XOR U21679 ( .A(n19886), .B(n19889), .Z(n19887) );
  XOR U21680 ( .A(n19890), .B(n19891), .Z(n19862) );
  XNOR U21681 ( .A(n19857), .B(n19892), .Z(n19891) );
  IV U21682 ( .A(n19860), .Z(n19892) );
  XOR U21683 ( .A(n19893), .B(n19894), .Z(n19860) );
  ANDN U21684 ( .B(n19895), .A(n19896), .Z(n19893) );
  XOR U21685 ( .A(n19894), .B(n19897), .Z(n19895) );
  XNOR U21686 ( .A(n19898), .B(n19899), .Z(n19857) );
  ANDN U21687 ( .B(n19900), .A(n19901), .Z(n19898) );
  XOR U21688 ( .A(n19899), .B(n19902), .Z(n19900) );
  IV U21689 ( .A(n19856), .Z(n19890) );
  XOR U21690 ( .A(n19854), .B(n19903), .Z(n19856) );
  XOR U21691 ( .A(n19904), .B(n19905), .Z(n19903) );
  ANDN U21692 ( .B(n19906), .A(n19907), .Z(n19904) );
  XOR U21693 ( .A(n19908), .B(n19905), .Z(n19906) );
  IV U21694 ( .A(n19858), .Z(n19854) );
  XOR U21695 ( .A(n19909), .B(n19910), .Z(n19858) );
  ANDN U21696 ( .B(n19911), .A(n19912), .Z(n19909) );
  XOR U21697 ( .A(n19913), .B(n19910), .Z(n19911) );
  IV U21698 ( .A(n19868), .Z(n19872) );
  XOR U21699 ( .A(n19868), .B(n19823), .Z(n19870) );
  XOR U21700 ( .A(n19914), .B(n19915), .Z(n19823) );
  AND U21701 ( .A(n350), .B(n19916), .Z(n19914) );
  XOR U21702 ( .A(n19917), .B(n19915), .Z(n19916) );
  NANDN U21703 ( .A(n19825), .B(n19827), .Z(n19868) );
  XOR U21704 ( .A(n19918), .B(n19919), .Z(n19827) );
  AND U21705 ( .A(n350), .B(n19920), .Z(n19918) );
  XOR U21706 ( .A(n19919), .B(n19921), .Z(n19920) );
  XNOR U21707 ( .A(n19922), .B(n19923), .Z(n350) );
  AND U21708 ( .A(n19924), .B(n19925), .Z(n19922) );
  XOR U21709 ( .A(n19923), .B(n19838), .Z(n19925) );
  XNOR U21710 ( .A(n19926), .B(n19927), .Z(n19838) );
  ANDN U21711 ( .B(n19928), .A(n19929), .Z(n19926) );
  XOR U21712 ( .A(n19927), .B(n19930), .Z(n19928) );
  XNOR U21713 ( .A(n19923), .B(n19840), .Z(n19924) );
  XOR U21714 ( .A(n19931), .B(n19932), .Z(n19840) );
  AND U21715 ( .A(n354), .B(n19933), .Z(n19931) );
  XOR U21716 ( .A(n19934), .B(n19932), .Z(n19933) );
  XNOR U21717 ( .A(n19935), .B(n19936), .Z(n19923) );
  AND U21718 ( .A(n19937), .B(n19938), .Z(n19935) );
  XNOR U21719 ( .A(n19936), .B(n19865), .Z(n19938) );
  XOR U21720 ( .A(n19929), .B(n19930), .Z(n19865) );
  XNOR U21721 ( .A(n19939), .B(n19940), .Z(n19930) );
  ANDN U21722 ( .B(n19941), .A(n19942), .Z(n19939) );
  XOR U21723 ( .A(n19943), .B(n19944), .Z(n19941) );
  XOR U21724 ( .A(n19945), .B(n19946), .Z(n19929) );
  XNOR U21725 ( .A(n19947), .B(n19948), .Z(n19946) );
  ANDN U21726 ( .B(n19949), .A(n19950), .Z(n19947) );
  XNOR U21727 ( .A(n19951), .B(n19952), .Z(n19949) );
  IV U21728 ( .A(n19927), .Z(n19945) );
  XOR U21729 ( .A(n19953), .B(n19954), .Z(n19927) );
  ANDN U21730 ( .B(n19955), .A(n19956), .Z(n19953) );
  XOR U21731 ( .A(n19954), .B(n19957), .Z(n19955) );
  XOR U21732 ( .A(n19936), .B(n19867), .Z(n19937) );
  XOR U21733 ( .A(n19958), .B(n19959), .Z(n19867) );
  AND U21734 ( .A(n354), .B(n19960), .Z(n19958) );
  XOR U21735 ( .A(n19961), .B(n19959), .Z(n19960) );
  XNOR U21736 ( .A(n19962), .B(n19963), .Z(n19936) );
  NAND U21737 ( .A(n19964), .B(n19965), .Z(n19963) );
  XOR U21738 ( .A(n19966), .B(n19915), .Z(n19965) );
  XOR U21739 ( .A(n19956), .B(n19957), .Z(n19915) );
  XOR U21740 ( .A(n19967), .B(n19944), .Z(n19957) );
  XOR U21741 ( .A(n19968), .B(n19969), .Z(n19944) );
  ANDN U21742 ( .B(n19970), .A(n19971), .Z(n19968) );
  XOR U21743 ( .A(n19969), .B(n19972), .Z(n19970) );
  IV U21744 ( .A(n19942), .Z(n19967) );
  XOR U21745 ( .A(n19940), .B(n19973), .Z(n19942) );
  XOR U21746 ( .A(n19974), .B(n19975), .Z(n19973) );
  ANDN U21747 ( .B(n19976), .A(n19977), .Z(n19974) );
  XOR U21748 ( .A(n19978), .B(n19975), .Z(n19976) );
  IV U21749 ( .A(n19943), .Z(n19940) );
  XOR U21750 ( .A(n19979), .B(n19980), .Z(n19943) );
  ANDN U21751 ( .B(n19981), .A(n19982), .Z(n19979) );
  XOR U21752 ( .A(n19980), .B(n19983), .Z(n19981) );
  XOR U21753 ( .A(n19984), .B(n19985), .Z(n19956) );
  XNOR U21754 ( .A(n19951), .B(n19986), .Z(n19985) );
  IV U21755 ( .A(n19954), .Z(n19986) );
  XOR U21756 ( .A(n19987), .B(n19988), .Z(n19954) );
  ANDN U21757 ( .B(n19989), .A(n19990), .Z(n19987) );
  XOR U21758 ( .A(n19988), .B(n19991), .Z(n19989) );
  XNOR U21759 ( .A(n19992), .B(n19993), .Z(n19951) );
  ANDN U21760 ( .B(n19994), .A(n19995), .Z(n19992) );
  XOR U21761 ( .A(n19993), .B(n19996), .Z(n19994) );
  IV U21762 ( .A(n19950), .Z(n19984) );
  XOR U21763 ( .A(n19948), .B(n19997), .Z(n19950) );
  XOR U21764 ( .A(n19998), .B(n19999), .Z(n19997) );
  ANDN U21765 ( .B(n20000), .A(n20001), .Z(n19998) );
  XOR U21766 ( .A(n20002), .B(n19999), .Z(n20000) );
  IV U21767 ( .A(n19952), .Z(n19948) );
  XOR U21768 ( .A(n20003), .B(n20004), .Z(n19952) );
  ANDN U21769 ( .B(n20005), .A(n20006), .Z(n20003) );
  XOR U21770 ( .A(n20007), .B(n20004), .Z(n20005) );
  IV U21771 ( .A(n19962), .Z(n19966) );
  XOR U21772 ( .A(n19962), .B(n19917), .Z(n19964) );
  XOR U21773 ( .A(n20008), .B(n20009), .Z(n19917) );
  AND U21774 ( .A(n354), .B(n20010), .Z(n20008) );
  XOR U21775 ( .A(n20011), .B(n20009), .Z(n20010) );
  NANDN U21776 ( .A(n19919), .B(n19921), .Z(n19962) );
  XOR U21777 ( .A(n20012), .B(n20013), .Z(n19921) );
  AND U21778 ( .A(n354), .B(n20014), .Z(n20012) );
  XOR U21779 ( .A(n20013), .B(n20015), .Z(n20014) );
  XNOR U21780 ( .A(n20016), .B(n20017), .Z(n354) );
  AND U21781 ( .A(n20018), .B(n20019), .Z(n20016) );
  XOR U21782 ( .A(n20017), .B(n19932), .Z(n20019) );
  XNOR U21783 ( .A(n20020), .B(n20021), .Z(n19932) );
  ANDN U21784 ( .B(n20022), .A(n20023), .Z(n20020) );
  XOR U21785 ( .A(n20021), .B(n20024), .Z(n20022) );
  XNOR U21786 ( .A(n20017), .B(n19934), .Z(n20018) );
  XOR U21787 ( .A(n20025), .B(n20026), .Z(n19934) );
  AND U21788 ( .A(n358), .B(n20027), .Z(n20025) );
  XOR U21789 ( .A(n20028), .B(n20026), .Z(n20027) );
  XNOR U21790 ( .A(n20029), .B(n20030), .Z(n20017) );
  AND U21791 ( .A(n20031), .B(n20032), .Z(n20029) );
  XNOR U21792 ( .A(n20030), .B(n19959), .Z(n20032) );
  XOR U21793 ( .A(n20023), .B(n20024), .Z(n19959) );
  XNOR U21794 ( .A(n20033), .B(n20034), .Z(n20024) );
  ANDN U21795 ( .B(n20035), .A(n20036), .Z(n20033) );
  XOR U21796 ( .A(n20037), .B(n20038), .Z(n20035) );
  XOR U21797 ( .A(n20039), .B(n20040), .Z(n20023) );
  XNOR U21798 ( .A(n20041), .B(n20042), .Z(n20040) );
  ANDN U21799 ( .B(n20043), .A(n20044), .Z(n20041) );
  XNOR U21800 ( .A(n20045), .B(n20046), .Z(n20043) );
  IV U21801 ( .A(n20021), .Z(n20039) );
  XOR U21802 ( .A(n20047), .B(n20048), .Z(n20021) );
  ANDN U21803 ( .B(n20049), .A(n20050), .Z(n20047) );
  XOR U21804 ( .A(n20048), .B(n20051), .Z(n20049) );
  XOR U21805 ( .A(n20030), .B(n19961), .Z(n20031) );
  XOR U21806 ( .A(n20052), .B(n20053), .Z(n19961) );
  AND U21807 ( .A(n358), .B(n20054), .Z(n20052) );
  XOR U21808 ( .A(n20055), .B(n20053), .Z(n20054) );
  XNOR U21809 ( .A(n20056), .B(n20057), .Z(n20030) );
  NAND U21810 ( .A(n20058), .B(n20059), .Z(n20057) );
  XOR U21811 ( .A(n20060), .B(n20009), .Z(n20059) );
  XOR U21812 ( .A(n20050), .B(n20051), .Z(n20009) );
  XOR U21813 ( .A(n20061), .B(n20038), .Z(n20051) );
  XOR U21814 ( .A(n20062), .B(n20063), .Z(n20038) );
  ANDN U21815 ( .B(n20064), .A(n20065), .Z(n20062) );
  XOR U21816 ( .A(n20063), .B(n20066), .Z(n20064) );
  IV U21817 ( .A(n20036), .Z(n20061) );
  XOR U21818 ( .A(n20034), .B(n20067), .Z(n20036) );
  XOR U21819 ( .A(n20068), .B(n20069), .Z(n20067) );
  ANDN U21820 ( .B(n20070), .A(n20071), .Z(n20068) );
  XOR U21821 ( .A(n20072), .B(n20069), .Z(n20070) );
  IV U21822 ( .A(n20037), .Z(n20034) );
  XOR U21823 ( .A(n20073), .B(n20074), .Z(n20037) );
  ANDN U21824 ( .B(n20075), .A(n20076), .Z(n20073) );
  XOR U21825 ( .A(n20074), .B(n20077), .Z(n20075) );
  XOR U21826 ( .A(n20078), .B(n20079), .Z(n20050) );
  XNOR U21827 ( .A(n20045), .B(n20080), .Z(n20079) );
  IV U21828 ( .A(n20048), .Z(n20080) );
  XOR U21829 ( .A(n20081), .B(n20082), .Z(n20048) );
  ANDN U21830 ( .B(n20083), .A(n20084), .Z(n20081) );
  XOR U21831 ( .A(n20082), .B(n20085), .Z(n20083) );
  XNOR U21832 ( .A(n20086), .B(n20087), .Z(n20045) );
  ANDN U21833 ( .B(n20088), .A(n20089), .Z(n20086) );
  XOR U21834 ( .A(n20087), .B(n20090), .Z(n20088) );
  IV U21835 ( .A(n20044), .Z(n20078) );
  XOR U21836 ( .A(n20042), .B(n20091), .Z(n20044) );
  XOR U21837 ( .A(n20092), .B(n20093), .Z(n20091) );
  ANDN U21838 ( .B(n20094), .A(n20095), .Z(n20092) );
  XOR U21839 ( .A(n20096), .B(n20093), .Z(n20094) );
  IV U21840 ( .A(n20046), .Z(n20042) );
  XOR U21841 ( .A(n20097), .B(n20098), .Z(n20046) );
  ANDN U21842 ( .B(n20099), .A(n20100), .Z(n20097) );
  XOR U21843 ( .A(n20101), .B(n20098), .Z(n20099) );
  IV U21844 ( .A(n20056), .Z(n20060) );
  XOR U21845 ( .A(n20056), .B(n20011), .Z(n20058) );
  XOR U21846 ( .A(n20102), .B(n20103), .Z(n20011) );
  AND U21847 ( .A(n358), .B(n20104), .Z(n20102) );
  XOR U21848 ( .A(n20105), .B(n20103), .Z(n20104) );
  NANDN U21849 ( .A(n20013), .B(n20015), .Z(n20056) );
  XOR U21850 ( .A(n20106), .B(n20107), .Z(n20015) );
  AND U21851 ( .A(n358), .B(n20108), .Z(n20106) );
  XOR U21852 ( .A(n20107), .B(n20109), .Z(n20108) );
  XNOR U21853 ( .A(n20110), .B(n20111), .Z(n358) );
  AND U21854 ( .A(n20112), .B(n20113), .Z(n20110) );
  XOR U21855 ( .A(n20111), .B(n20026), .Z(n20113) );
  XNOR U21856 ( .A(n20114), .B(n20115), .Z(n20026) );
  ANDN U21857 ( .B(n20116), .A(n20117), .Z(n20114) );
  XOR U21858 ( .A(n20115), .B(n20118), .Z(n20116) );
  XNOR U21859 ( .A(n20111), .B(n20028), .Z(n20112) );
  XOR U21860 ( .A(n20119), .B(n20120), .Z(n20028) );
  AND U21861 ( .A(n362), .B(n20121), .Z(n20119) );
  XOR U21862 ( .A(n20122), .B(n20120), .Z(n20121) );
  XNOR U21863 ( .A(n20123), .B(n20124), .Z(n20111) );
  AND U21864 ( .A(n20125), .B(n20126), .Z(n20123) );
  XNOR U21865 ( .A(n20124), .B(n20053), .Z(n20126) );
  XOR U21866 ( .A(n20117), .B(n20118), .Z(n20053) );
  XNOR U21867 ( .A(n20127), .B(n20128), .Z(n20118) );
  ANDN U21868 ( .B(n20129), .A(n20130), .Z(n20127) );
  XOR U21869 ( .A(n20131), .B(n20132), .Z(n20129) );
  XOR U21870 ( .A(n20133), .B(n20134), .Z(n20117) );
  XNOR U21871 ( .A(n20135), .B(n20136), .Z(n20134) );
  ANDN U21872 ( .B(n20137), .A(n20138), .Z(n20135) );
  XNOR U21873 ( .A(n20139), .B(n20140), .Z(n20137) );
  IV U21874 ( .A(n20115), .Z(n20133) );
  XOR U21875 ( .A(n20141), .B(n20142), .Z(n20115) );
  ANDN U21876 ( .B(n20143), .A(n20144), .Z(n20141) );
  XOR U21877 ( .A(n20142), .B(n20145), .Z(n20143) );
  XOR U21878 ( .A(n20124), .B(n20055), .Z(n20125) );
  XOR U21879 ( .A(n20146), .B(n20147), .Z(n20055) );
  AND U21880 ( .A(n362), .B(n20148), .Z(n20146) );
  XOR U21881 ( .A(n20149), .B(n20147), .Z(n20148) );
  XNOR U21882 ( .A(n20150), .B(n20151), .Z(n20124) );
  NAND U21883 ( .A(n20152), .B(n20153), .Z(n20151) );
  XOR U21884 ( .A(n20154), .B(n20103), .Z(n20153) );
  XOR U21885 ( .A(n20144), .B(n20145), .Z(n20103) );
  XOR U21886 ( .A(n20155), .B(n20132), .Z(n20145) );
  XOR U21887 ( .A(n20156), .B(n20157), .Z(n20132) );
  ANDN U21888 ( .B(n20158), .A(n20159), .Z(n20156) );
  XOR U21889 ( .A(n20157), .B(n20160), .Z(n20158) );
  IV U21890 ( .A(n20130), .Z(n20155) );
  XOR U21891 ( .A(n20128), .B(n20161), .Z(n20130) );
  XOR U21892 ( .A(n20162), .B(n20163), .Z(n20161) );
  ANDN U21893 ( .B(n20164), .A(n20165), .Z(n20162) );
  XOR U21894 ( .A(n20166), .B(n20163), .Z(n20164) );
  IV U21895 ( .A(n20131), .Z(n20128) );
  XOR U21896 ( .A(n20167), .B(n20168), .Z(n20131) );
  ANDN U21897 ( .B(n20169), .A(n20170), .Z(n20167) );
  XOR U21898 ( .A(n20168), .B(n20171), .Z(n20169) );
  XOR U21899 ( .A(n20172), .B(n20173), .Z(n20144) );
  XNOR U21900 ( .A(n20139), .B(n20174), .Z(n20173) );
  IV U21901 ( .A(n20142), .Z(n20174) );
  XOR U21902 ( .A(n20175), .B(n20176), .Z(n20142) );
  ANDN U21903 ( .B(n20177), .A(n20178), .Z(n20175) );
  XOR U21904 ( .A(n20176), .B(n20179), .Z(n20177) );
  XNOR U21905 ( .A(n20180), .B(n20181), .Z(n20139) );
  ANDN U21906 ( .B(n20182), .A(n20183), .Z(n20180) );
  XOR U21907 ( .A(n20181), .B(n20184), .Z(n20182) );
  IV U21908 ( .A(n20138), .Z(n20172) );
  XOR U21909 ( .A(n20136), .B(n20185), .Z(n20138) );
  XOR U21910 ( .A(n20186), .B(n20187), .Z(n20185) );
  ANDN U21911 ( .B(n20188), .A(n20189), .Z(n20186) );
  XOR U21912 ( .A(n20190), .B(n20187), .Z(n20188) );
  IV U21913 ( .A(n20140), .Z(n20136) );
  XOR U21914 ( .A(n20191), .B(n20192), .Z(n20140) );
  ANDN U21915 ( .B(n20193), .A(n20194), .Z(n20191) );
  XOR U21916 ( .A(n20195), .B(n20192), .Z(n20193) );
  IV U21917 ( .A(n20150), .Z(n20154) );
  XOR U21918 ( .A(n20150), .B(n20105), .Z(n20152) );
  XOR U21919 ( .A(n20196), .B(n20197), .Z(n20105) );
  AND U21920 ( .A(n362), .B(n20198), .Z(n20196) );
  XOR U21921 ( .A(n20199), .B(n20197), .Z(n20198) );
  NANDN U21922 ( .A(n20107), .B(n20109), .Z(n20150) );
  XOR U21923 ( .A(n20200), .B(n20201), .Z(n20109) );
  AND U21924 ( .A(n362), .B(n20202), .Z(n20200) );
  XOR U21925 ( .A(n20201), .B(n20203), .Z(n20202) );
  XNOR U21926 ( .A(n20204), .B(n20205), .Z(n362) );
  AND U21927 ( .A(n20206), .B(n20207), .Z(n20204) );
  XOR U21928 ( .A(n20205), .B(n20120), .Z(n20207) );
  XNOR U21929 ( .A(n20208), .B(n20209), .Z(n20120) );
  ANDN U21930 ( .B(n20210), .A(n20211), .Z(n20208) );
  XOR U21931 ( .A(n20209), .B(n20212), .Z(n20210) );
  XNOR U21932 ( .A(n20205), .B(n20122), .Z(n20206) );
  XOR U21933 ( .A(n20213), .B(n20214), .Z(n20122) );
  AND U21934 ( .A(n366), .B(n20215), .Z(n20213) );
  XOR U21935 ( .A(n20216), .B(n20214), .Z(n20215) );
  XNOR U21936 ( .A(n20217), .B(n20218), .Z(n20205) );
  AND U21937 ( .A(n20219), .B(n20220), .Z(n20217) );
  XNOR U21938 ( .A(n20218), .B(n20147), .Z(n20220) );
  XOR U21939 ( .A(n20211), .B(n20212), .Z(n20147) );
  XNOR U21940 ( .A(n20221), .B(n20222), .Z(n20212) );
  ANDN U21941 ( .B(n20223), .A(n20224), .Z(n20221) );
  XOR U21942 ( .A(n20225), .B(n20226), .Z(n20223) );
  XOR U21943 ( .A(n20227), .B(n20228), .Z(n20211) );
  XNOR U21944 ( .A(n20229), .B(n20230), .Z(n20228) );
  ANDN U21945 ( .B(n20231), .A(n20232), .Z(n20229) );
  XNOR U21946 ( .A(n20233), .B(n20234), .Z(n20231) );
  IV U21947 ( .A(n20209), .Z(n20227) );
  XOR U21948 ( .A(n20235), .B(n20236), .Z(n20209) );
  ANDN U21949 ( .B(n20237), .A(n20238), .Z(n20235) );
  XOR U21950 ( .A(n20236), .B(n20239), .Z(n20237) );
  XOR U21951 ( .A(n20218), .B(n20149), .Z(n20219) );
  XOR U21952 ( .A(n20240), .B(n20241), .Z(n20149) );
  AND U21953 ( .A(n366), .B(n20242), .Z(n20240) );
  XOR U21954 ( .A(n20243), .B(n20241), .Z(n20242) );
  XNOR U21955 ( .A(n20244), .B(n20245), .Z(n20218) );
  NAND U21956 ( .A(n20246), .B(n20247), .Z(n20245) );
  XOR U21957 ( .A(n20248), .B(n20197), .Z(n20247) );
  XOR U21958 ( .A(n20238), .B(n20239), .Z(n20197) );
  XOR U21959 ( .A(n20249), .B(n20226), .Z(n20239) );
  XOR U21960 ( .A(n20250), .B(n20251), .Z(n20226) );
  ANDN U21961 ( .B(n20252), .A(n20253), .Z(n20250) );
  XOR U21962 ( .A(n20251), .B(n20254), .Z(n20252) );
  IV U21963 ( .A(n20224), .Z(n20249) );
  XOR U21964 ( .A(n20222), .B(n20255), .Z(n20224) );
  XOR U21965 ( .A(n20256), .B(n20257), .Z(n20255) );
  ANDN U21966 ( .B(n20258), .A(n20259), .Z(n20256) );
  XOR U21967 ( .A(n20260), .B(n20257), .Z(n20258) );
  IV U21968 ( .A(n20225), .Z(n20222) );
  XOR U21969 ( .A(n20261), .B(n20262), .Z(n20225) );
  ANDN U21970 ( .B(n20263), .A(n20264), .Z(n20261) );
  XOR U21971 ( .A(n20262), .B(n20265), .Z(n20263) );
  XOR U21972 ( .A(n20266), .B(n20267), .Z(n20238) );
  XNOR U21973 ( .A(n20233), .B(n20268), .Z(n20267) );
  IV U21974 ( .A(n20236), .Z(n20268) );
  XOR U21975 ( .A(n20269), .B(n20270), .Z(n20236) );
  ANDN U21976 ( .B(n20271), .A(n20272), .Z(n20269) );
  XOR U21977 ( .A(n20270), .B(n20273), .Z(n20271) );
  XNOR U21978 ( .A(n20274), .B(n20275), .Z(n20233) );
  ANDN U21979 ( .B(n20276), .A(n20277), .Z(n20274) );
  XOR U21980 ( .A(n20275), .B(n20278), .Z(n20276) );
  IV U21981 ( .A(n20232), .Z(n20266) );
  XOR U21982 ( .A(n20230), .B(n20279), .Z(n20232) );
  XOR U21983 ( .A(n20280), .B(n20281), .Z(n20279) );
  ANDN U21984 ( .B(n20282), .A(n20283), .Z(n20280) );
  XOR U21985 ( .A(n20284), .B(n20281), .Z(n20282) );
  IV U21986 ( .A(n20234), .Z(n20230) );
  XOR U21987 ( .A(n20285), .B(n20286), .Z(n20234) );
  ANDN U21988 ( .B(n20287), .A(n20288), .Z(n20285) );
  XOR U21989 ( .A(n20289), .B(n20286), .Z(n20287) );
  IV U21990 ( .A(n20244), .Z(n20248) );
  XOR U21991 ( .A(n20244), .B(n20199), .Z(n20246) );
  XOR U21992 ( .A(n20290), .B(n20291), .Z(n20199) );
  AND U21993 ( .A(n366), .B(n20292), .Z(n20290) );
  XOR U21994 ( .A(n20293), .B(n20291), .Z(n20292) );
  NANDN U21995 ( .A(n20201), .B(n20203), .Z(n20244) );
  XOR U21996 ( .A(n20294), .B(n20295), .Z(n20203) );
  AND U21997 ( .A(n366), .B(n20296), .Z(n20294) );
  XOR U21998 ( .A(n20295), .B(n20297), .Z(n20296) );
  XNOR U21999 ( .A(n20298), .B(n20299), .Z(n366) );
  AND U22000 ( .A(n20300), .B(n20301), .Z(n20298) );
  XOR U22001 ( .A(n20299), .B(n20214), .Z(n20301) );
  XNOR U22002 ( .A(n20302), .B(n20303), .Z(n20214) );
  ANDN U22003 ( .B(n20304), .A(n20305), .Z(n20302) );
  XOR U22004 ( .A(n20303), .B(n20306), .Z(n20304) );
  XNOR U22005 ( .A(n20299), .B(n20216), .Z(n20300) );
  XOR U22006 ( .A(n20307), .B(n20308), .Z(n20216) );
  AND U22007 ( .A(n370), .B(n20309), .Z(n20307) );
  XOR U22008 ( .A(n20310), .B(n20308), .Z(n20309) );
  XNOR U22009 ( .A(n20311), .B(n20312), .Z(n20299) );
  AND U22010 ( .A(n20313), .B(n20314), .Z(n20311) );
  XNOR U22011 ( .A(n20312), .B(n20241), .Z(n20314) );
  XOR U22012 ( .A(n20305), .B(n20306), .Z(n20241) );
  XNOR U22013 ( .A(n20315), .B(n20316), .Z(n20306) );
  ANDN U22014 ( .B(n20317), .A(n20318), .Z(n20315) );
  XOR U22015 ( .A(n20319), .B(n20320), .Z(n20317) );
  XOR U22016 ( .A(n20321), .B(n20322), .Z(n20305) );
  XNOR U22017 ( .A(n20323), .B(n20324), .Z(n20322) );
  ANDN U22018 ( .B(n20325), .A(n20326), .Z(n20323) );
  XNOR U22019 ( .A(n20327), .B(n20328), .Z(n20325) );
  IV U22020 ( .A(n20303), .Z(n20321) );
  XOR U22021 ( .A(n20329), .B(n20330), .Z(n20303) );
  ANDN U22022 ( .B(n20331), .A(n20332), .Z(n20329) );
  XOR U22023 ( .A(n20330), .B(n20333), .Z(n20331) );
  XOR U22024 ( .A(n20312), .B(n20243), .Z(n20313) );
  XOR U22025 ( .A(n20334), .B(n20335), .Z(n20243) );
  AND U22026 ( .A(n370), .B(n20336), .Z(n20334) );
  XOR U22027 ( .A(n20337), .B(n20335), .Z(n20336) );
  XNOR U22028 ( .A(n20338), .B(n20339), .Z(n20312) );
  NAND U22029 ( .A(n20340), .B(n20341), .Z(n20339) );
  XOR U22030 ( .A(n20342), .B(n20291), .Z(n20341) );
  XOR U22031 ( .A(n20332), .B(n20333), .Z(n20291) );
  XOR U22032 ( .A(n20343), .B(n20320), .Z(n20333) );
  XOR U22033 ( .A(n20344), .B(n20345), .Z(n20320) );
  ANDN U22034 ( .B(n20346), .A(n20347), .Z(n20344) );
  XOR U22035 ( .A(n20345), .B(n20348), .Z(n20346) );
  IV U22036 ( .A(n20318), .Z(n20343) );
  XOR U22037 ( .A(n20316), .B(n20349), .Z(n20318) );
  XOR U22038 ( .A(n20350), .B(n20351), .Z(n20349) );
  ANDN U22039 ( .B(n20352), .A(n20353), .Z(n20350) );
  XOR U22040 ( .A(n20354), .B(n20351), .Z(n20352) );
  IV U22041 ( .A(n20319), .Z(n20316) );
  XOR U22042 ( .A(n20355), .B(n20356), .Z(n20319) );
  ANDN U22043 ( .B(n20357), .A(n20358), .Z(n20355) );
  XOR U22044 ( .A(n20356), .B(n20359), .Z(n20357) );
  XOR U22045 ( .A(n20360), .B(n20361), .Z(n20332) );
  XNOR U22046 ( .A(n20327), .B(n20362), .Z(n20361) );
  IV U22047 ( .A(n20330), .Z(n20362) );
  XOR U22048 ( .A(n20363), .B(n20364), .Z(n20330) );
  ANDN U22049 ( .B(n20365), .A(n20366), .Z(n20363) );
  XOR U22050 ( .A(n20364), .B(n20367), .Z(n20365) );
  XNOR U22051 ( .A(n20368), .B(n20369), .Z(n20327) );
  ANDN U22052 ( .B(n20370), .A(n20371), .Z(n20368) );
  XOR U22053 ( .A(n20369), .B(n20372), .Z(n20370) );
  IV U22054 ( .A(n20326), .Z(n20360) );
  XOR U22055 ( .A(n20324), .B(n20373), .Z(n20326) );
  XOR U22056 ( .A(n20374), .B(n20375), .Z(n20373) );
  ANDN U22057 ( .B(n20376), .A(n20377), .Z(n20374) );
  XOR U22058 ( .A(n20378), .B(n20375), .Z(n20376) );
  IV U22059 ( .A(n20328), .Z(n20324) );
  XOR U22060 ( .A(n20379), .B(n20380), .Z(n20328) );
  ANDN U22061 ( .B(n20381), .A(n20382), .Z(n20379) );
  XOR U22062 ( .A(n20383), .B(n20380), .Z(n20381) );
  IV U22063 ( .A(n20338), .Z(n20342) );
  XOR U22064 ( .A(n20338), .B(n20293), .Z(n20340) );
  XOR U22065 ( .A(n20384), .B(n20385), .Z(n20293) );
  AND U22066 ( .A(n370), .B(n20386), .Z(n20384) );
  XOR U22067 ( .A(n20387), .B(n20385), .Z(n20386) );
  NANDN U22068 ( .A(n20295), .B(n20297), .Z(n20338) );
  XOR U22069 ( .A(n20388), .B(n20389), .Z(n20297) );
  AND U22070 ( .A(n370), .B(n20390), .Z(n20388) );
  XOR U22071 ( .A(n20389), .B(n20391), .Z(n20390) );
  XNOR U22072 ( .A(n20392), .B(n20393), .Z(n370) );
  AND U22073 ( .A(n20394), .B(n20395), .Z(n20392) );
  XOR U22074 ( .A(n20393), .B(n20308), .Z(n20395) );
  XNOR U22075 ( .A(n20396), .B(n20397), .Z(n20308) );
  ANDN U22076 ( .B(n20398), .A(n20399), .Z(n20396) );
  XOR U22077 ( .A(n20397), .B(n20400), .Z(n20398) );
  XNOR U22078 ( .A(n20393), .B(n20310), .Z(n20394) );
  XOR U22079 ( .A(n20401), .B(n20402), .Z(n20310) );
  AND U22080 ( .A(n374), .B(n20403), .Z(n20401) );
  XOR U22081 ( .A(n20404), .B(n20402), .Z(n20403) );
  XNOR U22082 ( .A(n20405), .B(n20406), .Z(n20393) );
  AND U22083 ( .A(n20407), .B(n20408), .Z(n20405) );
  XNOR U22084 ( .A(n20406), .B(n20335), .Z(n20408) );
  XOR U22085 ( .A(n20399), .B(n20400), .Z(n20335) );
  XNOR U22086 ( .A(n20409), .B(n20410), .Z(n20400) );
  ANDN U22087 ( .B(n20411), .A(n20412), .Z(n20409) );
  XOR U22088 ( .A(n20413), .B(n20414), .Z(n20411) );
  XOR U22089 ( .A(n20415), .B(n20416), .Z(n20399) );
  XNOR U22090 ( .A(n20417), .B(n20418), .Z(n20416) );
  ANDN U22091 ( .B(n20419), .A(n20420), .Z(n20417) );
  XNOR U22092 ( .A(n20421), .B(n20422), .Z(n20419) );
  IV U22093 ( .A(n20397), .Z(n20415) );
  XOR U22094 ( .A(n20423), .B(n20424), .Z(n20397) );
  ANDN U22095 ( .B(n20425), .A(n20426), .Z(n20423) );
  XOR U22096 ( .A(n20424), .B(n20427), .Z(n20425) );
  XOR U22097 ( .A(n20406), .B(n20337), .Z(n20407) );
  XOR U22098 ( .A(n20428), .B(n20429), .Z(n20337) );
  AND U22099 ( .A(n374), .B(n20430), .Z(n20428) );
  XOR U22100 ( .A(n20431), .B(n20429), .Z(n20430) );
  XNOR U22101 ( .A(n20432), .B(n20433), .Z(n20406) );
  NAND U22102 ( .A(n20434), .B(n20435), .Z(n20433) );
  XOR U22103 ( .A(n20436), .B(n20385), .Z(n20435) );
  XOR U22104 ( .A(n20426), .B(n20427), .Z(n20385) );
  XOR U22105 ( .A(n20437), .B(n20414), .Z(n20427) );
  XOR U22106 ( .A(n20438), .B(n20439), .Z(n20414) );
  ANDN U22107 ( .B(n20440), .A(n20441), .Z(n20438) );
  XOR U22108 ( .A(n20439), .B(n20442), .Z(n20440) );
  IV U22109 ( .A(n20412), .Z(n20437) );
  XOR U22110 ( .A(n20410), .B(n20443), .Z(n20412) );
  XOR U22111 ( .A(n20444), .B(n20445), .Z(n20443) );
  ANDN U22112 ( .B(n20446), .A(n20447), .Z(n20444) );
  XOR U22113 ( .A(n20448), .B(n20445), .Z(n20446) );
  IV U22114 ( .A(n20413), .Z(n20410) );
  XOR U22115 ( .A(n20449), .B(n20450), .Z(n20413) );
  ANDN U22116 ( .B(n20451), .A(n20452), .Z(n20449) );
  XOR U22117 ( .A(n20450), .B(n20453), .Z(n20451) );
  XOR U22118 ( .A(n20454), .B(n20455), .Z(n20426) );
  XNOR U22119 ( .A(n20421), .B(n20456), .Z(n20455) );
  IV U22120 ( .A(n20424), .Z(n20456) );
  XOR U22121 ( .A(n20457), .B(n20458), .Z(n20424) );
  ANDN U22122 ( .B(n20459), .A(n20460), .Z(n20457) );
  XOR U22123 ( .A(n20458), .B(n20461), .Z(n20459) );
  XNOR U22124 ( .A(n20462), .B(n20463), .Z(n20421) );
  ANDN U22125 ( .B(n20464), .A(n20465), .Z(n20462) );
  XOR U22126 ( .A(n20463), .B(n20466), .Z(n20464) );
  IV U22127 ( .A(n20420), .Z(n20454) );
  XOR U22128 ( .A(n20418), .B(n20467), .Z(n20420) );
  XOR U22129 ( .A(n20468), .B(n20469), .Z(n20467) );
  ANDN U22130 ( .B(n20470), .A(n20471), .Z(n20468) );
  XOR U22131 ( .A(n20472), .B(n20469), .Z(n20470) );
  IV U22132 ( .A(n20422), .Z(n20418) );
  XOR U22133 ( .A(n20473), .B(n20474), .Z(n20422) );
  ANDN U22134 ( .B(n20475), .A(n20476), .Z(n20473) );
  XOR U22135 ( .A(n20477), .B(n20474), .Z(n20475) );
  IV U22136 ( .A(n20432), .Z(n20436) );
  XOR U22137 ( .A(n20432), .B(n20387), .Z(n20434) );
  XOR U22138 ( .A(n20478), .B(n20479), .Z(n20387) );
  AND U22139 ( .A(n374), .B(n20480), .Z(n20478) );
  XOR U22140 ( .A(n20481), .B(n20479), .Z(n20480) );
  NANDN U22141 ( .A(n20389), .B(n20391), .Z(n20432) );
  XOR U22142 ( .A(n20482), .B(n20483), .Z(n20391) );
  AND U22143 ( .A(n374), .B(n20484), .Z(n20482) );
  XOR U22144 ( .A(n20483), .B(n20485), .Z(n20484) );
  XNOR U22145 ( .A(n20486), .B(n20487), .Z(n374) );
  AND U22146 ( .A(n20488), .B(n20489), .Z(n20486) );
  XOR U22147 ( .A(n20487), .B(n20402), .Z(n20489) );
  XNOR U22148 ( .A(n20490), .B(n20491), .Z(n20402) );
  ANDN U22149 ( .B(n20492), .A(n20493), .Z(n20490) );
  XOR U22150 ( .A(n20491), .B(n20494), .Z(n20492) );
  XNOR U22151 ( .A(n20487), .B(n20404), .Z(n20488) );
  XOR U22152 ( .A(n20495), .B(n20496), .Z(n20404) );
  AND U22153 ( .A(n378), .B(n20497), .Z(n20495) );
  XOR U22154 ( .A(n20498), .B(n20496), .Z(n20497) );
  XNOR U22155 ( .A(n20499), .B(n20500), .Z(n20487) );
  AND U22156 ( .A(n20501), .B(n20502), .Z(n20499) );
  XNOR U22157 ( .A(n20500), .B(n20429), .Z(n20502) );
  XOR U22158 ( .A(n20493), .B(n20494), .Z(n20429) );
  XNOR U22159 ( .A(n20503), .B(n20504), .Z(n20494) );
  ANDN U22160 ( .B(n20505), .A(n20506), .Z(n20503) );
  XOR U22161 ( .A(n20507), .B(n20508), .Z(n20505) );
  XOR U22162 ( .A(n20509), .B(n20510), .Z(n20493) );
  XNOR U22163 ( .A(n20511), .B(n20512), .Z(n20510) );
  ANDN U22164 ( .B(n20513), .A(n20514), .Z(n20511) );
  XNOR U22165 ( .A(n20515), .B(n20516), .Z(n20513) );
  IV U22166 ( .A(n20491), .Z(n20509) );
  XOR U22167 ( .A(n20517), .B(n20518), .Z(n20491) );
  ANDN U22168 ( .B(n20519), .A(n20520), .Z(n20517) );
  XOR U22169 ( .A(n20518), .B(n20521), .Z(n20519) );
  XOR U22170 ( .A(n20500), .B(n20431), .Z(n20501) );
  XOR U22171 ( .A(n20522), .B(n20523), .Z(n20431) );
  AND U22172 ( .A(n378), .B(n20524), .Z(n20522) );
  XOR U22173 ( .A(n20525), .B(n20523), .Z(n20524) );
  XNOR U22174 ( .A(n20526), .B(n20527), .Z(n20500) );
  NAND U22175 ( .A(n20528), .B(n20529), .Z(n20527) );
  XOR U22176 ( .A(n20530), .B(n20479), .Z(n20529) );
  XOR U22177 ( .A(n20520), .B(n20521), .Z(n20479) );
  XOR U22178 ( .A(n20531), .B(n20508), .Z(n20521) );
  XOR U22179 ( .A(n20532), .B(n20533), .Z(n20508) );
  ANDN U22180 ( .B(n20534), .A(n20535), .Z(n20532) );
  XOR U22181 ( .A(n20533), .B(n20536), .Z(n20534) );
  IV U22182 ( .A(n20506), .Z(n20531) );
  XOR U22183 ( .A(n20504), .B(n20537), .Z(n20506) );
  XOR U22184 ( .A(n20538), .B(n20539), .Z(n20537) );
  ANDN U22185 ( .B(n20540), .A(n20541), .Z(n20538) );
  XOR U22186 ( .A(n20542), .B(n20539), .Z(n20540) );
  IV U22187 ( .A(n20507), .Z(n20504) );
  XOR U22188 ( .A(n20543), .B(n20544), .Z(n20507) );
  ANDN U22189 ( .B(n20545), .A(n20546), .Z(n20543) );
  XOR U22190 ( .A(n20544), .B(n20547), .Z(n20545) );
  XOR U22191 ( .A(n20548), .B(n20549), .Z(n20520) );
  XNOR U22192 ( .A(n20515), .B(n20550), .Z(n20549) );
  IV U22193 ( .A(n20518), .Z(n20550) );
  XOR U22194 ( .A(n20551), .B(n20552), .Z(n20518) );
  ANDN U22195 ( .B(n20553), .A(n20554), .Z(n20551) );
  XOR U22196 ( .A(n20552), .B(n20555), .Z(n20553) );
  XNOR U22197 ( .A(n20556), .B(n20557), .Z(n20515) );
  ANDN U22198 ( .B(n20558), .A(n20559), .Z(n20556) );
  XOR U22199 ( .A(n20557), .B(n20560), .Z(n20558) );
  IV U22200 ( .A(n20514), .Z(n20548) );
  XOR U22201 ( .A(n20512), .B(n20561), .Z(n20514) );
  XOR U22202 ( .A(n20562), .B(n20563), .Z(n20561) );
  ANDN U22203 ( .B(n20564), .A(n20565), .Z(n20562) );
  XOR U22204 ( .A(n20566), .B(n20563), .Z(n20564) );
  IV U22205 ( .A(n20516), .Z(n20512) );
  XOR U22206 ( .A(n20567), .B(n20568), .Z(n20516) );
  ANDN U22207 ( .B(n20569), .A(n20570), .Z(n20567) );
  XOR U22208 ( .A(n20571), .B(n20568), .Z(n20569) );
  IV U22209 ( .A(n20526), .Z(n20530) );
  XOR U22210 ( .A(n20526), .B(n20481), .Z(n20528) );
  XOR U22211 ( .A(n20572), .B(n20573), .Z(n20481) );
  AND U22212 ( .A(n378), .B(n20574), .Z(n20572) );
  XOR U22213 ( .A(n20575), .B(n20573), .Z(n20574) );
  NANDN U22214 ( .A(n20483), .B(n20485), .Z(n20526) );
  XOR U22215 ( .A(n20576), .B(n20577), .Z(n20485) );
  AND U22216 ( .A(n378), .B(n20578), .Z(n20576) );
  XOR U22217 ( .A(n20577), .B(n20579), .Z(n20578) );
  XNOR U22218 ( .A(n20580), .B(n20581), .Z(n378) );
  AND U22219 ( .A(n20582), .B(n20583), .Z(n20580) );
  XOR U22220 ( .A(n20581), .B(n20496), .Z(n20583) );
  XNOR U22221 ( .A(n20584), .B(n20585), .Z(n20496) );
  ANDN U22222 ( .B(n20586), .A(n20587), .Z(n20584) );
  XOR U22223 ( .A(n20585), .B(n20588), .Z(n20586) );
  XNOR U22224 ( .A(n20581), .B(n20498), .Z(n20582) );
  XOR U22225 ( .A(n20589), .B(n20590), .Z(n20498) );
  AND U22226 ( .A(n382), .B(n20591), .Z(n20589) );
  XOR U22227 ( .A(n20592), .B(n20590), .Z(n20591) );
  XNOR U22228 ( .A(n20593), .B(n20594), .Z(n20581) );
  AND U22229 ( .A(n20595), .B(n20596), .Z(n20593) );
  XNOR U22230 ( .A(n20594), .B(n20523), .Z(n20596) );
  XOR U22231 ( .A(n20587), .B(n20588), .Z(n20523) );
  XNOR U22232 ( .A(n20597), .B(n20598), .Z(n20588) );
  ANDN U22233 ( .B(n20599), .A(n20600), .Z(n20597) );
  XOR U22234 ( .A(n20601), .B(n20602), .Z(n20599) );
  XOR U22235 ( .A(n20603), .B(n20604), .Z(n20587) );
  XNOR U22236 ( .A(n20605), .B(n20606), .Z(n20604) );
  ANDN U22237 ( .B(n20607), .A(n20608), .Z(n20605) );
  XNOR U22238 ( .A(n20609), .B(n20610), .Z(n20607) );
  IV U22239 ( .A(n20585), .Z(n20603) );
  XOR U22240 ( .A(n20611), .B(n20612), .Z(n20585) );
  ANDN U22241 ( .B(n20613), .A(n20614), .Z(n20611) );
  XOR U22242 ( .A(n20612), .B(n20615), .Z(n20613) );
  XOR U22243 ( .A(n20594), .B(n20525), .Z(n20595) );
  XOR U22244 ( .A(n20616), .B(n20617), .Z(n20525) );
  AND U22245 ( .A(n382), .B(n20618), .Z(n20616) );
  XOR U22246 ( .A(n20619), .B(n20617), .Z(n20618) );
  XNOR U22247 ( .A(n20620), .B(n20621), .Z(n20594) );
  NAND U22248 ( .A(n20622), .B(n20623), .Z(n20621) );
  XOR U22249 ( .A(n20624), .B(n20573), .Z(n20623) );
  XOR U22250 ( .A(n20614), .B(n20615), .Z(n20573) );
  XOR U22251 ( .A(n20625), .B(n20602), .Z(n20615) );
  XOR U22252 ( .A(n20626), .B(n20627), .Z(n20602) );
  ANDN U22253 ( .B(n20628), .A(n20629), .Z(n20626) );
  XOR U22254 ( .A(n20627), .B(n20630), .Z(n20628) );
  IV U22255 ( .A(n20600), .Z(n20625) );
  XOR U22256 ( .A(n20598), .B(n20631), .Z(n20600) );
  XOR U22257 ( .A(n20632), .B(n20633), .Z(n20631) );
  ANDN U22258 ( .B(n20634), .A(n20635), .Z(n20632) );
  XOR U22259 ( .A(n20636), .B(n20633), .Z(n20634) );
  IV U22260 ( .A(n20601), .Z(n20598) );
  XOR U22261 ( .A(n20637), .B(n20638), .Z(n20601) );
  ANDN U22262 ( .B(n20639), .A(n20640), .Z(n20637) );
  XOR U22263 ( .A(n20638), .B(n20641), .Z(n20639) );
  XOR U22264 ( .A(n20642), .B(n20643), .Z(n20614) );
  XNOR U22265 ( .A(n20609), .B(n20644), .Z(n20643) );
  IV U22266 ( .A(n20612), .Z(n20644) );
  XOR U22267 ( .A(n20645), .B(n20646), .Z(n20612) );
  ANDN U22268 ( .B(n20647), .A(n20648), .Z(n20645) );
  XOR U22269 ( .A(n20646), .B(n20649), .Z(n20647) );
  XNOR U22270 ( .A(n20650), .B(n20651), .Z(n20609) );
  ANDN U22271 ( .B(n20652), .A(n20653), .Z(n20650) );
  XOR U22272 ( .A(n20651), .B(n20654), .Z(n20652) );
  IV U22273 ( .A(n20608), .Z(n20642) );
  XOR U22274 ( .A(n20606), .B(n20655), .Z(n20608) );
  XOR U22275 ( .A(n20656), .B(n20657), .Z(n20655) );
  ANDN U22276 ( .B(n20658), .A(n20659), .Z(n20656) );
  XOR U22277 ( .A(n20660), .B(n20657), .Z(n20658) );
  IV U22278 ( .A(n20610), .Z(n20606) );
  XOR U22279 ( .A(n20661), .B(n20662), .Z(n20610) );
  ANDN U22280 ( .B(n20663), .A(n20664), .Z(n20661) );
  XOR U22281 ( .A(n20665), .B(n20662), .Z(n20663) );
  IV U22282 ( .A(n20620), .Z(n20624) );
  XOR U22283 ( .A(n20620), .B(n20575), .Z(n20622) );
  XOR U22284 ( .A(n20666), .B(n20667), .Z(n20575) );
  AND U22285 ( .A(n382), .B(n20668), .Z(n20666) );
  XOR U22286 ( .A(n20669), .B(n20667), .Z(n20668) );
  NANDN U22287 ( .A(n20577), .B(n20579), .Z(n20620) );
  XOR U22288 ( .A(n20670), .B(n20671), .Z(n20579) );
  AND U22289 ( .A(n382), .B(n20672), .Z(n20670) );
  XOR U22290 ( .A(n20671), .B(n20673), .Z(n20672) );
  XNOR U22291 ( .A(n20674), .B(n20675), .Z(n382) );
  AND U22292 ( .A(n20676), .B(n20677), .Z(n20674) );
  XOR U22293 ( .A(n20675), .B(n20590), .Z(n20677) );
  XNOR U22294 ( .A(n20678), .B(n20679), .Z(n20590) );
  ANDN U22295 ( .B(n20680), .A(n20681), .Z(n20678) );
  XOR U22296 ( .A(n20679), .B(n20682), .Z(n20680) );
  XNOR U22297 ( .A(n20675), .B(n20592), .Z(n20676) );
  XOR U22298 ( .A(n20683), .B(n20684), .Z(n20592) );
  AND U22299 ( .A(n386), .B(n20685), .Z(n20683) );
  XOR U22300 ( .A(n20686), .B(n20684), .Z(n20685) );
  XNOR U22301 ( .A(n20687), .B(n20688), .Z(n20675) );
  AND U22302 ( .A(n20689), .B(n20690), .Z(n20687) );
  XNOR U22303 ( .A(n20688), .B(n20617), .Z(n20690) );
  XOR U22304 ( .A(n20681), .B(n20682), .Z(n20617) );
  XNOR U22305 ( .A(n20691), .B(n20692), .Z(n20682) );
  ANDN U22306 ( .B(n20693), .A(n20694), .Z(n20691) );
  XOR U22307 ( .A(n20695), .B(n20696), .Z(n20693) );
  XOR U22308 ( .A(n20697), .B(n20698), .Z(n20681) );
  XNOR U22309 ( .A(n20699), .B(n20700), .Z(n20698) );
  ANDN U22310 ( .B(n20701), .A(n20702), .Z(n20699) );
  XNOR U22311 ( .A(n20703), .B(n20704), .Z(n20701) );
  IV U22312 ( .A(n20679), .Z(n20697) );
  XOR U22313 ( .A(n20705), .B(n20706), .Z(n20679) );
  ANDN U22314 ( .B(n20707), .A(n20708), .Z(n20705) );
  XOR U22315 ( .A(n20706), .B(n20709), .Z(n20707) );
  XOR U22316 ( .A(n20688), .B(n20619), .Z(n20689) );
  XOR U22317 ( .A(n20710), .B(n20711), .Z(n20619) );
  AND U22318 ( .A(n386), .B(n20712), .Z(n20710) );
  XOR U22319 ( .A(n20713), .B(n20711), .Z(n20712) );
  XNOR U22320 ( .A(n20714), .B(n20715), .Z(n20688) );
  NAND U22321 ( .A(n20716), .B(n20717), .Z(n20715) );
  XOR U22322 ( .A(n20718), .B(n20667), .Z(n20717) );
  XOR U22323 ( .A(n20708), .B(n20709), .Z(n20667) );
  XOR U22324 ( .A(n20719), .B(n20696), .Z(n20709) );
  XOR U22325 ( .A(n20720), .B(n20721), .Z(n20696) );
  ANDN U22326 ( .B(n20722), .A(n20723), .Z(n20720) );
  XOR U22327 ( .A(n20721), .B(n20724), .Z(n20722) );
  IV U22328 ( .A(n20694), .Z(n20719) );
  XOR U22329 ( .A(n20692), .B(n20725), .Z(n20694) );
  XOR U22330 ( .A(n20726), .B(n20727), .Z(n20725) );
  ANDN U22331 ( .B(n20728), .A(n20729), .Z(n20726) );
  XOR U22332 ( .A(n20730), .B(n20727), .Z(n20728) );
  IV U22333 ( .A(n20695), .Z(n20692) );
  XOR U22334 ( .A(n20731), .B(n20732), .Z(n20695) );
  ANDN U22335 ( .B(n20733), .A(n20734), .Z(n20731) );
  XOR U22336 ( .A(n20732), .B(n20735), .Z(n20733) );
  XOR U22337 ( .A(n20736), .B(n20737), .Z(n20708) );
  XNOR U22338 ( .A(n20703), .B(n20738), .Z(n20737) );
  IV U22339 ( .A(n20706), .Z(n20738) );
  XOR U22340 ( .A(n20739), .B(n20740), .Z(n20706) );
  ANDN U22341 ( .B(n20741), .A(n20742), .Z(n20739) );
  XOR U22342 ( .A(n20740), .B(n20743), .Z(n20741) );
  XNOR U22343 ( .A(n20744), .B(n20745), .Z(n20703) );
  ANDN U22344 ( .B(n20746), .A(n20747), .Z(n20744) );
  XOR U22345 ( .A(n20745), .B(n20748), .Z(n20746) );
  IV U22346 ( .A(n20702), .Z(n20736) );
  XOR U22347 ( .A(n20700), .B(n20749), .Z(n20702) );
  XOR U22348 ( .A(n20750), .B(n20751), .Z(n20749) );
  ANDN U22349 ( .B(n20752), .A(n20753), .Z(n20750) );
  XOR U22350 ( .A(n20754), .B(n20751), .Z(n20752) );
  IV U22351 ( .A(n20704), .Z(n20700) );
  XOR U22352 ( .A(n20755), .B(n20756), .Z(n20704) );
  ANDN U22353 ( .B(n20757), .A(n20758), .Z(n20755) );
  XOR U22354 ( .A(n20759), .B(n20756), .Z(n20757) );
  IV U22355 ( .A(n20714), .Z(n20718) );
  XOR U22356 ( .A(n20714), .B(n20669), .Z(n20716) );
  XOR U22357 ( .A(n20760), .B(n20761), .Z(n20669) );
  AND U22358 ( .A(n386), .B(n20762), .Z(n20760) );
  XOR U22359 ( .A(n20763), .B(n20761), .Z(n20762) );
  NANDN U22360 ( .A(n20671), .B(n20673), .Z(n20714) );
  XOR U22361 ( .A(n20764), .B(n20765), .Z(n20673) );
  AND U22362 ( .A(n386), .B(n20766), .Z(n20764) );
  XOR U22363 ( .A(n20765), .B(n20767), .Z(n20766) );
  XNOR U22364 ( .A(n20768), .B(n20769), .Z(n386) );
  AND U22365 ( .A(n20770), .B(n20771), .Z(n20768) );
  XOR U22366 ( .A(n20769), .B(n20684), .Z(n20771) );
  XNOR U22367 ( .A(n20772), .B(n20773), .Z(n20684) );
  ANDN U22368 ( .B(n20774), .A(n20775), .Z(n20772) );
  XOR U22369 ( .A(n20773), .B(n20776), .Z(n20774) );
  XNOR U22370 ( .A(n20769), .B(n20686), .Z(n20770) );
  XOR U22371 ( .A(n20777), .B(n20778), .Z(n20686) );
  AND U22372 ( .A(n390), .B(n20779), .Z(n20777) );
  XOR U22373 ( .A(n20780), .B(n20778), .Z(n20779) );
  XNOR U22374 ( .A(n20781), .B(n20782), .Z(n20769) );
  AND U22375 ( .A(n20783), .B(n20784), .Z(n20781) );
  XNOR U22376 ( .A(n20782), .B(n20711), .Z(n20784) );
  XOR U22377 ( .A(n20775), .B(n20776), .Z(n20711) );
  XNOR U22378 ( .A(n20785), .B(n20786), .Z(n20776) );
  ANDN U22379 ( .B(n20787), .A(n20788), .Z(n20785) );
  XOR U22380 ( .A(n20789), .B(n20790), .Z(n20787) );
  XOR U22381 ( .A(n20791), .B(n20792), .Z(n20775) );
  XNOR U22382 ( .A(n20793), .B(n20794), .Z(n20792) );
  ANDN U22383 ( .B(n20795), .A(n20796), .Z(n20793) );
  XNOR U22384 ( .A(n20797), .B(n20798), .Z(n20795) );
  IV U22385 ( .A(n20773), .Z(n20791) );
  XOR U22386 ( .A(n20799), .B(n20800), .Z(n20773) );
  ANDN U22387 ( .B(n20801), .A(n20802), .Z(n20799) );
  XOR U22388 ( .A(n20800), .B(n20803), .Z(n20801) );
  XOR U22389 ( .A(n20782), .B(n20713), .Z(n20783) );
  XOR U22390 ( .A(n20804), .B(n20805), .Z(n20713) );
  AND U22391 ( .A(n390), .B(n20806), .Z(n20804) );
  XOR U22392 ( .A(n20807), .B(n20805), .Z(n20806) );
  XNOR U22393 ( .A(n20808), .B(n20809), .Z(n20782) );
  NAND U22394 ( .A(n20810), .B(n20811), .Z(n20809) );
  XOR U22395 ( .A(n20812), .B(n20761), .Z(n20811) );
  XOR U22396 ( .A(n20802), .B(n20803), .Z(n20761) );
  XOR U22397 ( .A(n20813), .B(n20790), .Z(n20803) );
  XOR U22398 ( .A(n20814), .B(n20815), .Z(n20790) );
  ANDN U22399 ( .B(n20816), .A(n20817), .Z(n20814) );
  XOR U22400 ( .A(n20815), .B(n20818), .Z(n20816) );
  IV U22401 ( .A(n20788), .Z(n20813) );
  XOR U22402 ( .A(n20786), .B(n20819), .Z(n20788) );
  XOR U22403 ( .A(n20820), .B(n20821), .Z(n20819) );
  ANDN U22404 ( .B(n20822), .A(n20823), .Z(n20820) );
  XOR U22405 ( .A(n20824), .B(n20821), .Z(n20822) );
  IV U22406 ( .A(n20789), .Z(n20786) );
  XOR U22407 ( .A(n20825), .B(n20826), .Z(n20789) );
  ANDN U22408 ( .B(n20827), .A(n20828), .Z(n20825) );
  XOR U22409 ( .A(n20826), .B(n20829), .Z(n20827) );
  XOR U22410 ( .A(n20830), .B(n20831), .Z(n20802) );
  XNOR U22411 ( .A(n20797), .B(n20832), .Z(n20831) );
  IV U22412 ( .A(n20800), .Z(n20832) );
  XOR U22413 ( .A(n20833), .B(n20834), .Z(n20800) );
  ANDN U22414 ( .B(n20835), .A(n20836), .Z(n20833) );
  XOR U22415 ( .A(n20834), .B(n20837), .Z(n20835) );
  XNOR U22416 ( .A(n20838), .B(n20839), .Z(n20797) );
  ANDN U22417 ( .B(n20840), .A(n20841), .Z(n20838) );
  XOR U22418 ( .A(n20839), .B(n20842), .Z(n20840) );
  IV U22419 ( .A(n20796), .Z(n20830) );
  XOR U22420 ( .A(n20794), .B(n20843), .Z(n20796) );
  XOR U22421 ( .A(n20844), .B(n20845), .Z(n20843) );
  ANDN U22422 ( .B(n20846), .A(n20847), .Z(n20844) );
  XOR U22423 ( .A(n20848), .B(n20845), .Z(n20846) );
  IV U22424 ( .A(n20798), .Z(n20794) );
  XOR U22425 ( .A(n20849), .B(n20850), .Z(n20798) );
  ANDN U22426 ( .B(n20851), .A(n20852), .Z(n20849) );
  XOR U22427 ( .A(n20853), .B(n20850), .Z(n20851) );
  IV U22428 ( .A(n20808), .Z(n20812) );
  XOR U22429 ( .A(n20808), .B(n20763), .Z(n20810) );
  XOR U22430 ( .A(n20854), .B(n20855), .Z(n20763) );
  AND U22431 ( .A(n390), .B(n20856), .Z(n20854) );
  XOR U22432 ( .A(n20857), .B(n20855), .Z(n20856) );
  NANDN U22433 ( .A(n20765), .B(n20767), .Z(n20808) );
  XOR U22434 ( .A(n20858), .B(n20859), .Z(n20767) );
  AND U22435 ( .A(n390), .B(n20860), .Z(n20858) );
  XOR U22436 ( .A(n20859), .B(n20861), .Z(n20860) );
  XNOR U22437 ( .A(n20862), .B(n20863), .Z(n390) );
  AND U22438 ( .A(n20864), .B(n20865), .Z(n20862) );
  XOR U22439 ( .A(n20863), .B(n20778), .Z(n20865) );
  XNOR U22440 ( .A(n20866), .B(n20867), .Z(n20778) );
  ANDN U22441 ( .B(n20868), .A(n20869), .Z(n20866) );
  XOR U22442 ( .A(n20867), .B(n20870), .Z(n20868) );
  XNOR U22443 ( .A(n20863), .B(n20780), .Z(n20864) );
  XOR U22444 ( .A(n20871), .B(n20872), .Z(n20780) );
  AND U22445 ( .A(n394), .B(n20873), .Z(n20871) );
  XOR U22446 ( .A(n20874), .B(n20872), .Z(n20873) );
  XNOR U22447 ( .A(n20875), .B(n20876), .Z(n20863) );
  AND U22448 ( .A(n20877), .B(n20878), .Z(n20875) );
  XNOR U22449 ( .A(n20876), .B(n20805), .Z(n20878) );
  XOR U22450 ( .A(n20869), .B(n20870), .Z(n20805) );
  XNOR U22451 ( .A(n20879), .B(n20880), .Z(n20870) );
  ANDN U22452 ( .B(n20881), .A(n20882), .Z(n20879) );
  XOR U22453 ( .A(n20883), .B(n20884), .Z(n20881) );
  XOR U22454 ( .A(n20885), .B(n20886), .Z(n20869) );
  XNOR U22455 ( .A(n20887), .B(n20888), .Z(n20886) );
  ANDN U22456 ( .B(n20889), .A(n20890), .Z(n20887) );
  XNOR U22457 ( .A(n20891), .B(n20892), .Z(n20889) );
  IV U22458 ( .A(n20867), .Z(n20885) );
  XOR U22459 ( .A(n20893), .B(n20894), .Z(n20867) );
  ANDN U22460 ( .B(n20895), .A(n20896), .Z(n20893) );
  XOR U22461 ( .A(n20894), .B(n20897), .Z(n20895) );
  XOR U22462 ( .A(n20876), .B(n20807), .Z(n20877) );
  XOR U22463 ( .A(n20898), .B(n20899), .Z(n20807) );
  AND U22464 ( .A(n394), .B(n20900), .Z(n20898) );
  XOR U22465 ( .A(n20901), .B(n20899), .Z(n20900) );
  XNOR U22466 ( .A(n20902), .B(n20903), .Z(n20876) );
  NAND U22467 ( .A(n20904), .B(n20905), .Z(n20903) );
  XOR U22468 ( .A(n20906), .B(n20855), .Z(n20905) );
  XOR U22469 ( .A(n20896), .B(n20897), .Z(n20855) );
  XOR U22470 ( .A(n20907), .B(n20884), .Z(n20897) );
  XOR U22471 ( .A(n20908), .B(n20909), .Z(n20884) );
  ANDN U22472 ( .B(n20910), .A(n20911), .Z(n20908) );
  XOR U22473 ( .A(n20909), .B(n20912), .Z(n20910) );
  IV U22474 ( .A(n20882), .Z(n20907) );
  XOR U22475 ( .A(n20880), .B(n20913), .Z(n20882) );
  XOR U22476 ( .A(n20914), .B(n20915), .Z(n20913) );
  ANDN U22477 ( .B(n20916), .A(n20917), .Z(n20914) );
  XOR U22478 ( .A(n20918), .B(n20915), .Z(n20916) );
  IV U22479 ( .A(n20883), .Z(n20880) );
  XOR U22480 ( .A(n20919), .B(n20920), .Z(n20883) );
  ANDN U22481 ( .B(n20921), .A(n20922), .Z(n20919) );
  XOR U22482 ( .A(n20920), .B(n20923), .Z(n20921) );
  XOR U22483 ( .A(n20924), .B(n20925), .Z(n20896) );
  XNOR U22484 ( .A(n20891), .B(n20926), .Z(n20925) );
  IV U22485 ( .A(n20894), .Z(n20926) );
  XOR U22486 ( .A(n20927), .B(n20928), .Z(n20894) );
  ANDN U22487 ( .B(n20929), .A(n20930), .Z(n20927) );
  XOR U22488 ( .A(n20928), .B(n20931), .Z(n20929) );
  XNOR U22489 ( .A(n20932), .B(n20933), .Z(n20891) );
  ANDN U22490 ( .B(n20934), .A(n20935), .Z(n20932) );
  XOR U22491 ( .A(n20933), .B(n20936), .Z(n20934) );
  IV U22492 ( .A(n20890), .Z(n20924) );
  XOR U22493 ( .A(n20888), .B(n20937), .Z(n20890) );
  XOR U22494 ( .A(n20938), .B(n20939), .Z(n20937) );
  ANDN U22495 ( .B(n20940), .A(n20941), .Z(n20938) );
  XOR U22496 ( .A(n20942), .B(n20939), .Z(n20940) );
  IV U22497 ( .A(n20892), .Z(n20888) );
  XOR U22498 ( .A(n20943), .B(n20944), .Z(n20892) );
  ANDN U22499 ( .B(n20945), .A(n20946), .Z(n20943) );
  XOR U22500 ( .A(n20947), .B(n20944), .Z(n20945) );
  IV U22501 ( .A(n20902), .Z(n20906) );
  XOR U22502 ( .A(n20902), .B(n20857), .Z(n20904) );
  XOR U22503 ( .A(n20948), .B(n20949), .Z(n20857) );
  AND U22504 ( .A(n394), .B(n20950), .Z(n20948) );
  XOR U22505 ( .A(n20951), .B(n20949), .Z(n20950) );
  NANDN U22506 ( .A(n20859), .B(n20861), .Z(n20902) );
  XOR U22507 ( .A(n20952), .B(n20953), .Z(n20861) );
  AND U22508 ( .A(n394), .B(n20954), .Z(n20952) );
  XOR U22509 ( .A(n20953), .B(n20955), .Z(n20954) );
  XNOR U22510 ( .A(n20956), .B(n20957), .Z(n394) );
  AND U22511 ( .A(n20958), .B(n20959), .Z(n20956) );
  XOR U22512 ( .A(n20957), .B(n20872), .Z(n20959) );
  XNOR U22513 ( .A(n20960), .B(n20961), .Z(n20872) );
  ANDN U22514 ( .B(n20962), .A(n20963), .Z(n20960) );
  XOR U22515 ( .A(n20961), .B(n20964), .Z(n20962) );
  XNOR U22516 ( .A(n20957), .B(n20874), .Z(n20958) );
  XOR U22517 ( .A(n20965), .B(n20966), .Z(n20874) );
  AND U22518 ( .A(n398), .B(n20967), .Z(n20965) );
  XOR U22519 ( .A(n20968), .B(n20966), .Z(n20967) );
  XNOR U22520 ( .A(n20969), .B(n20970), .Z(n20957) );
  AND U22521 ( .A(n20971), .B(n20972), .Z(n20969) );
  XNOR U22522 ( .A(n20970), .B(n20899), .Z(n20972) );
  XOR U22523 ( .A(n20963), .B(n20964), .Z(n20899) );
  XNOR U22524 ( .A(n20973), .B(n20974), .Z(n20964) );
  ANDN U22525 ( .B(n20975), .A(n20976), .Z(n20973) );
  XOR U22526 ( .A(n20977), .B(n20978), .Z(n20975) );
  XOR U22527 ( .A(n20979), .B(n20980), .Z(n20963) );
  XNOR U22528 ( .A(n20981), .B(n20982), .Z(n20980) );
  ANDN U22529 ( .B(n20983), .A(n20984), .Z(n20981) );
  XNOR U22530 ( .A(n20985), .B(n20986), .Z(n20983) );
  IV U22531 ( .A(n20961), .Z(n20979) );
  XOR U22532 ( .A(n20987), .B(n20988), .Z(n20961) );
  ANDN U22533 ( .B(n20989), .A(n20990), .Z(n20987) );
  XOR U22534 ( .A(n20988), .B(n20991), .Z(n20989) );
  XOR U22535 ( .A(n20970), .B(n20901), .Z(n20971) );
  XOR U22536 ( .A(n20992), .B(n20993), .Z(n20901) );
  AND U22537 ( .A(n398), .B(n20994), .Z(n20992) );
  XOR U22538 ( .A(n20995), .B(n20993), .Z(n20994) );
  XNOR U22539 ( .A(n20996), .B(n20997), .Z(n20970) );
  NAND U22540 ( .A(n20998), .B(n20999), .Z(n20997) );
  XOR U22541 ( .A(n21000), .B(n20949), .Z(n20999) );
  XOR U22542 ( .A(n20990), .B(n20991), .Z(n20949) );
  XOR U22543 ( .A(n21001), .B(n20978), .Z(n20991) );
  XOR U22544 ( .A(n21002), .B(n21003), .Z(n20978) );
  ANDN U22545 ( .B(n21004), .A(n21005), .Z(n21002) );
  XOR U22546 ( .A(n21003), .B(n21006), .Z(n21004) );
  IV U22547 ( .A(n20976), .Z(n21001) );
  XOR U22548 ( .A(n20974), .B(n21007), .Z(n20976) );
  XOR U22549 ( .A(n21008), .B(n21009), .Z(n21007) );
  ANDN U22550 ( .B(n21010), .A(n21011), .Z(n21008) );
  XOR U22551 ( .A(n21012), .B(n21009), .Z(n21010) );
  IV U22552 ( .A(n20977), .Z(n20974) );
  XOR U22553 ( .A(n21013), .B(n21014), .Z(n20977) );
  ANDN U22554 ( .B(n21015), .A(n21016), .Z(n21013) );
  XOR U22555 ( .A(n21014), .B(n21017), .Z(n21015) );
  XOR U22556 ( .A(n21018), .B(n21019), .Z(n20990) );
  XNOR U22557 ( .A(n20985), .B(n21020), .Z(n21019) );
  IV U22558 ( .A(n20988), .Z(n21020) );
  XOR U22559 ( .A(n21021), .B(n21022), .Z(n20988) );
  ANDN U22560 ( .B(n21023), .A(n21024), .Z(n21021) );
  XOR U22561 ( .A(n21022), .B(n21025), .Z(n21023) );
  XNOR U22562 ( .A(n21026), .B(n21027), .Z(n20985) );
  ANDN U22563 ( .B(n21028), .A(n21029), .Z(n21026) );
  XOR U22564 ( .A(n21027), .B(n21030), .Z(n21028) );
  IV U22565 ( .A(n20984), .Z(n21018) );
  XOR U22566 ( .A(n20982), .B(n21031), .Z(n20984) );
  XOR U22567 ( .A(n21032), .B(n21033), .Z(n21031) );
  ANDN U22568 ( .B(n21034), .A(n21035), .Z(n21032) );
  XOR U22569 ( .A(n21036), .B(n21033), .Z(n21034) );
  IV U22570 ( .A(n20986), .Z(n20982) );
  XOR U22571 ( .A(n21037), .B(n21038), .Z(n20986) );
  ANDN U22572 ( .B(n21039), .A(n21040), .Z(n21037) );
  XOR U22573 ( .A(n21041), .B(n21038), .Z(n21039) );
  IV U22574 ( .A(n20996), .Z(n21000) );
  XOR U22575 ( .A(n20996), .B(n20951), .Z(n20998) );
  XOR U22576 ( .A(n21042), .B(n21043), .Z(n20951) );
  AND U22577 ( .A(n398), .B(n21044), .Z(n21042) );
  XOR U22578 ( .A(n21045), .B(n21043), .Z(n21044) );
  NANDN U22579 ( .A(n20953), .B(n20955), .Z(n20996) );
  XOR U22580 ( .A(n21046), .B(n21047), .Z(n20955) );
  AND U22581 ( .A(n398), .B(n21048), .Z(n21046) );
  XOR U22582 ( .A(n21047), .B(n21049), .Z(n21048) );
  XNOR U22583 ( .A(n21050), .B(n21051), .Z(n398) );
  AND U22584 ( .A(n21052), .B(n21053), .Z(n21050) );
  XOR U22585 ( .A(n21051), .B(n20966), .Z(n21053) );
  XNOR U22586 ( .A(n21054), .B(n21055), .Z(n20966) );
  ANDN U22587 ( .B(n21056), .A(n21057), .Z(n21054) );
  XOR U22588 ( .A(n21055), .B(n21058), .Z(n21056) );
  XNOR U22589 ( .A(n21051), .B(n20968), .Z(n21052) );
  XOR U22590 ( .A(n21059), .B(n21060), .Z(n20968) );
  AND U22591 ( .A(n402), .B(n21061), .Z(n21059) );
  XOR U22592 ( .A(n21062), .B(n21060), .Z(n21061) );
  XNOR U22593 ( .A(n21063), .B(n21064), .Z(n21051) );
  AND U22594 ( .A(n21065), .B(n21066), .Z(n21063) );
  XNOR U22595 ( .A(n21064), .B(n20993), .Z(n21066) );
  XOR U22596 ( .A(n21057), .B(n21058), .Z(n20993) );
  XNOR U22597 ( .A(n21067), .B(n21068), .Z(n21058) );
  ANDN U22598 ( .B(n21069), .A(n21070), .Z(n21067) );
  XOR U22599 ( .A(n21071), .B(n21072), .Z(n21069) );
  XOR U22600 ( .A(n21073), .B(n21074), .Z(n21057) );
  XNOR U22601 ( .A(n21075), .B(n21076), .Z(n21074) );
  ANDN U22602 ( .B(n21077), .A(n21078), .Z(n21075) );
  XNOR U22603 ( .A(n21079), .B(n21080), .Z(n21077) );
  IV U22604 ( .A(n21055), .Z(n21073) );
  XOR U22605 ( .A(n21081), .B(n21082), .Z(n21055) );
  ANDN U22606 ( .B(n21083), .A(n21084), .Z(n21081) );
  XOR U22607 ( .A(n21082), .B(n21085), .Z(n21083) );
  XOR U22608 ( .A(n21064), .B(n20995), .Z(n21065) );
  XOR U22609 ( .A(n21086), .B(n21087), .Z(n20995) );
  AND U22610 ( .A(n402), .B(n21088), .Z(n21086) );
  XOR U22611 ( .A(n21089), .B(n21087), .Z(n21088) );
  XNOR U22612 ( .A(n21090), .B(n21091), .Z(n21064) );
  NAND U22613 ( .A(n21092), .B(n21093), .Z(n21091) );
  XOR U22614 ( .A(n21094), .B(n21043), .Z(n21093) );
  XOR U22615 ( .A(n21084), .B(n21085), .Z(n21043) );
  XOR U22616 ( .A(n21095), .B(n21072), .Z(n21085) );
  XOR U22617 ( .A(n21096), .B(n21097), .Z(n21072) );
  ANDN U22618 ( .B(n21098), .A(n21099), .Z(n21096) );
  XOR U22619 ( .A(n21097), .B(n21100), .Z(n21098) );
  IV U22620 ( .A(n21070), .Z(n21095) );
  XOR U22621 ( .A(n21068), .B(n21101), .Z(n21070) );
  XOR U22622 ( .A(n21102), .B(n21103), .Z(n21101) );
  ANDN U22623 ( .B(n21104), .A(n21105), .Z(n21102) );
  XOR U22624 ( .A(n21106), .B(n21103), .Z(n21104) );
  IV U22625 ( .A(n21071), .Z(n21068) );
  XOR U22626 ( .A(n21107), .B(n21108), .Z(n21071) );
  ANDN U22627 ( .B(n21109), .A(n21110), .Z(n21107) );
  XOR U22628 ( .A(n21108), .B(n21111), .Z(n21109) );
  XOR U22629 ( .A(n21112), .B(n21113), .Z(n21084) );
  XNOR U22630 ( .A(n21079), .B(n21114), .Z(n21113) );
  IV U22631 ( .A(n21082), .Z(n21114) );
  XOR U22632 ( .A(n21115), .B(n21116), .Z(n21082) );
  ANDN U22633 ( .B(n21117), .A(n21118), .Z(n21115) );
  XOR U22634 ( .A(n21116), .B(n21119), .Z(n21117) );
  XNOR U22635 ( .A(n21120), .B(n21121), .Z(n21079) );
  ANDN U22636 ( .B(n21122), .A(n21123), .Z(n21120) );
  XOR U22637 ( .A(n21121), .B(n21124), .Z(n21122) );
  IV U22638 ( .A(n21078), .Z(n21112) );
  XOR U22639 ( .A(n21076), .B(n21125), .Z(n21078) );
  XOR U22640 ( .A(n21126), .B(n21127), .Z(n21125) );
  ANDN U22641 ( .B(n21128), .A(n21129), .Z(n21126) );
  XOR U22642 ( .A(n21130), .B(n21127), .Z(n21128) );
  IV U22643 ( .A(n21080), .Z(n21076) );
  XOR U22644 ( .A(n21131), .B(n21132), .Z(n21080) );
  ANDN U22645 ( .B(n21133), .A(n21134), .Z(n21131) );
  XOR U22646 ( .A(n21135), .B(n21132), .Z(n21133) );
  IV U22647 ( .A(n21090), .Z(n21094) );
  XOR U22648 ( .A(n21090), .B(n21045), .Z(n21092) );
  XOR U22649 ( .A(n21136), .B(n21137), .Z(n21045) );
  AND U22650 ( .A(n402), .B(n21138), .Z(n21136) );
  XOR U22651 ( .A(n21139), .B(n21137), .Z(n21138) );
  NANDN U22652 ( .A(n21047), .B(n21049), .Z(n21090) );
  XOR U22653 ( .A(n21140), .B(n21141), .Z(n21049) );
  AND U22654 ( .A(n402), .B(n21142), .Z(n21140) );
  XOR U22655 ( .A(n21141), .B(n21143), .Z(n21142) );
  XNOR U22656 ( .A(n21144), .B(n21145), .Z(n402) );
  AND U22657 ( .A(n21146), .B(n21147), .Z(n21144) );
  XOR U22658 ( .A(n21145), .B(n21060), .Z(n21147) );
  XNOR U22659 ( .A(n21148), .B(n21149), .Z(n21060) );
  ANDN U22660 ( .B(n21150), .A(n21151), .Z(n21148) );
  XOR U22661 ( .A(n21149), .B(n21152), .Z(n21150) );
  XNOR U22662 ( .A(n21145), .B(n21062), .Z(n21146) );
  XOR U22663 ( .A(n21153), .B(n21154), .Z(n21062) );
  AND U22664 ( .A(n406), .B(n21155), .Z(n21153) );
  XOR U22665 ( .A(n21156), .B(n21154), .Z(n21155) );
  XNOR U22666 ( .A(n21157), .B(n21158), .Z(n21145) );
  AND U22667 ( .A(n21159), .B(n21160), .Z(n21157) );
  XNOR U22668 ( .A(n21158), .B(n21087), .Z(n21160) );
  XOR U22669 ( .A(n21151), .B(n21152), .Z(n21087) );
  XNOR U22670 ( .A(n21161), .B(n21162), .Z(n21152) );
  ANDN U22671 ( .B(n21163), .A(n21164), .Z(n21161) );
  XOR U22672 ( .A(n21165), .B(n21166), .Z(n21163) );
  XOR U22673 ( .A(n21167), .B(n21168), .Z(n21151) );
  XNOR U22674 ( .A(n21169), .B(n21170), .Z(n21168) );
  ANDN U22675 ( .B(n21171), .A(n21172), .Z(n21169) );
  XNOR U22676 ( .A(n21173), .B(n21174), .Z(n21171) );
  IV U22677 ( .A(n21149), .Z(n21167) );
  XOR U22678 ( .A(n21175), .B(n21176), .Z(n21149) );
  ANDN U22679 ( .B(n21177), .A(n21178), .Z(n21175) );
  XOR U22680 ( .A(n21176), .B(n21179), .Z(n21177) );
  XOR U22681 ( .A(n21158), .B(n21089), .Z(n21159) );
  XOR U22682 ( .A(n21180), .B(n21181), .Z(n21089) );
  AND U22683 ( .A(n406), .B(n21182), .Z(n21180) );
  XOR U22684 ( .A(n21183), .B(n21181), .Z(n21182) );
  XNOR U22685 ( .A(n21184), .B(n21185), .Z(n21158) );
  NAND U22686 ( .A(n21186), .B(n21187), .Z(n21185) );
  XOR U22687 ( .A(n21188), .B(n21137), .Z(n21187) );
  XOR U22688 ( .A(n21178), .B(n21179), .Z(n21137) );
  XOR U22689 ( .A(n21189), .B(n21166), .Z(n21179) );
  XOR U22690 ( .A(n21190), .B(n21191), .Z(n21166) );
  ANDN U22691 ( .B(n21192), .A(n21193), .Z(n21190) );
  XOR U22692 ( .A(n21191), .B(n21194), .Z(n21192) );
  IV U22693 ( .A(n21164), .Z(n21189) );
  XOR U22694 ( .A(n21162), .B(n21195), .Z(n21164) );
  XOR U22695 ( .A(n21196), .B(n21197), .Z(n21195) );
  ANDN U22696 ( .B(n21198), .A(n21199), .Z(n21196) );
  XOR U22697 ( .A(n21200), .B(n21197), .Z(n21198) );
  IV U22698 ( .A(n21165), .Z(n21162) );
  XOR U22699 ( .A(n21201), .B(n21202), .Z(n21165) );
  ANDN U22700 ( .B(n21203), .A(n21204), .Z(n21201) );
  XOR U22701 ( .A(n21202), .B(n21205), .Z(n21203) );
  XOR U22702 ( .A(n21206), .B(n21207), .Z(n21178) );
  XNOR U22703 ( .A(n21173), .B(n21208), .Z(n21207) );
  IV U22704 ( .A(n21176), .Z(n21208) );
  XOR U22705 ( .A(n21209), .B(n21210), .Z(n21176) );
  ANDN U22706 ( .B(n21211), .A(n21212), .Z(n21209) );
  XOR U22707 ( .A(n21210), .B(n21213), .Z(n21211) );
  XNOR U22708 ( .A(n21214), .B(n21215), .Z(n21173) );
  ANDN U22709 ( .B(n21216), .A(n21217), .Z(n21214) );
  XOR U22710 ( .A(n21215), .B(n21218), .Z(n21216) );
  IV U22711 ( .A(n21172), .Z(n21206) );
  XOR U22712 ( .A(n21170), .B(n21219), .Z(n21172) );
  XOR U22713 ( .A(n21220), .B(n21221), .Z(n21219) );
  ANDN U22714 ( .B(n21222), .A(n21223), .Z(n21220) );
  XOR U22715 ( .A(n21224), .B(n21221), .Z(n21222) );
  IV U22716 ( .A(n21174), .Z(n21170) );
  XOR U22717 ( .A(n21225), .B(n21226), .Z(n21174) );
  ANDN U22718 ( .B(n21227), .A(n21228), .Z(n21225) );
  XOR U22719 ( .A(n21229), .B(n21226), .Z(n21227) );
  IV U22720 ( .A(n21184), .Z(n21188) );
  XOR U22721 ( .A(n21184), .B(n21139), .Z(n21186) );
  XOR U22722 ( .A(n21230), .B(n21231), .Z(n21139) );
  AND U22723 ( .A(n406), .B(n21232), .Z(n21230) );
  XOR U22724 ( .A(n21233), .B(n21231), .Z(n21232) );
  NANDN U22725 ( .A(n21141), .B(n21143), .Z(n21184) );
  XOR U22726 ( .A(n21234), .B(n21235), .Z(n21143) );
  AND U22727 ( .A(n406), .B(n21236), .Z(n21234) );
  XOR U22728 ( .A(n21235), .B(n21237), .Z(n21236) );
  XNOR U22729 ( .A(n21238), .B(n21239), .Z(n406) );
  AND U22730 ( .A(n21240), .B(n21241), .Z(n21238) );
  XOR U22731 ( .A(n21239), .B(n21154), .Z(n21241) );
  XNOR U22732 ( .A(n21242), .B(n21243), .Z(n21154) );
  ANDN U22733 ( .B(n21244), .A(n21245), .Z(n21242) );
  XOR U22734 ( .A(n21243), .B(n21246), .Z(n21244) );
  XNOR U22735 ( .A(n21239), .B(n21156), .Z(n21240) );
  XOR U22736 ( .A(n21247), .B(n21248), .Z(n21156) );
  AND U22737 ( .A(n410), .B(n21249), .Z(n21247) );
  XOR U22738 ( .A(n21250), .B(n21248), .Z(n21249) );
  XNOR U22739 ( .A(n21251), .B(n21252), .Z(n21239) );
  AND U22740 ( .A(n21253), .B(n21254), .Z(n21251) );
  XNOR U22741 ( .A(n21252), .B(n21181), .Z(n21254) );
  XOR U22742 ( .A(n21245), .B(n21246), .Z(n21181) );
  XNOR U22743 ( .A(n21255), .B(n21256), .Z(n21246) );
  ANDN U22744 ( .B(n21257), .A(n21258), .Z(n21255) );
  XOR U22745 ( .A(n21259), .B(n21260), .Z(n21257) );
  XOR U22746 ( .A(n21261), .B(n21262), .Z(n21245) );
  XNOR U22747 ( .A(n21263), .B(n21264), .Z(n21262) );
  ANDN U22748 ( .B(n21265), .A(n21266), .Z(n21263) );
  XNOR U22749 ( .A(n21267), .B(n21268), .Z(n21265) );
  IV U22750 ( .A(n21243), .Z(n21261) );
  XOR U22751 ( .A(n21269), .B(n21270), .Z(n21243) );
  ANDN U22752 ( .B(n21271), .A(n21272), .Z(n21269) );
  XOR U22753 ( .A(n21270), .B(n21273), .Z(n21271) );
  XOR U22754 ( .A(n21252), .B(n21183), .Z(n21253) );
  XOR U22755 ( .A(n21274), .B(n21275), .Z(n21183) );
  AND U22756 ( .A(n410), .B(n21276), .Z(n21274) );
  XOR U22757 ( .A(n21277), .B(n21275), .Z(n21276) );
  XNOR U22758 ( .A(n21278), .B(n21279), .Z(n21252) );
  NAND U22759 ( .A(n21280), .B(n21281), .Z(n21279) );
  XOR U22760 ( .A(n21282), .B(n21231), .Z(n21281) );
  XOR U22761 ( .A(n21272), .B(n21273), .Z(n21231) );
  XOR U22762 ( .A(n21283), .B(n21260), .Z(n21273) );
  XOR U22763 ( .A(n21284), .B(n21285), .Z(n21260) );
  ANDN U22764 ( .B(n21286), .A(n21287), .Z(n21284) );
  XOR U22765 ( .A(n21285), .B(n21288), .Z(n21286) );
  IV U22766 ( .A(n21258), .Z(n21283) );
  XOR U22767 ( .A(n21256), .B(n21289), .Z(n21258) );
  XOR U22768 ( .A(n21290), .B(n21291), .Z(n21289) );
  ANDN U22769 ( .B(n21292), .A(n21293), .Z(n21290) );
  XOR U22770 ( .A(n21294), .B(n21291), .Z(n21292) );
  IV U22771 ( .A(n21259), .Z(n21256) );
  XOR U22772 ( .A(n21295), .B(n21296), .Z(n21259) );
  ANDN U22773 ( .B(n21297), .A(n21298), .Z(n21295) );
  XOR U22774 ( .A(n21296), .B(n21299), .Z(n21297) );
  XOR U22775 ( .A(n21300), .B(n21301), .Z(n21272) );
  XNOR U22776 ( .A(n21267), .B(n21302), .Z(n21301) );
  IV U22777 ( .A(n21270), .Z(n21302) );
  XOR U22778 ( .A(n21303), .B(n21304), .Z(n21270) );
  ANDN U22779 ( .B(n21305), .A(n21306), .Z(n21303) );
  XOR U22780 ( .A(n21304), .B(n21307), .Z(n21305) );
  XNOR U22781 ( .A(n21308), .B(n21309), .Z(n21267) );
  ANDN U22782 ( .B(n21310), .A(n21311), .Z(n21308) );
  XOR U22783 ( .A(n21309), .B(n21312), .Z(n21310) );
  IV U22784 ( .A(n21266), .Z(n21300) );
  XOR U22785 ( .A(n21264), .B(n21313), .Z(n21266) );
  XOR U22786 ( .A(n21314), .B(n21315), .Z(n21313) );
  ANDN U22787 ( .B(n21316), .A(n21317), .Z(n21314) );
  XOR U22788 ( .A(n21318), .B(n21315), .Z(n21316) );
  IV U22789 ( .A(n21268), .Z(n21264) );
  XOR U22790 ( .A(n21319), .B(n21320), .Z(n21268) );
  ANDN U22791 ( .B(n21321), .A(n21322), .Z(n21319) );
  XOR U22792 ( .A(n21323), .B(n21320), .Z(n21321) );
  IV U22793 ( .A(n21278), .Z(n21282) );
  XOR U22794 ( .A(n21278), .B(n21233), .Z(n21280) );
  XOR U22795 ( .A(n21324), .B(n21325), .Z(n21233) );
  AND U22796 ( .A(n410), .B(n21326), .Z(n21324) );
  XOR U22797 ( .A(n21327), .B(n21325), .Z(n21326) );
  NANDN U22798 ( .A(n21235), .B(n21237), .Z(n21278) );
  XOR U22799 ( .A(n21328), .B(n21329), .Z(n21237) );
  AND U22800 ( .A(n410), .B(n21330), .Z(n21328) );
  XOR U22801 ( .A(n21329), .B(n21331), .Z(n21330) );
  XNOR U22802 ( .A(n21332), .B(n21333), .Z(n410) );
  AND U22803 ( .A(n21334), .B(n21335), .Z(n21332) );
  XOR U22804 ( .A(n21333), .B(n21248), .Z(n21335) );
  XNOR U22805 ( .A(n21336), .B(n21337), .Z(n21248) );
  ANDN U22806 ( .B(n21338), .A(n21339), .Z(n21336) );
  XOR U22807 ( .A(n21337), .B(n21340), .Z(n21338) );
  XNOR U22808 ( .A(n21333), .B(n21250), .Z(n21334) );
  XOR U22809 ( .A(n21341), .B(n21342), .Z(n21250) );
  AND U22810 ( .A(n414), .B(n21343), .Z(n21341) );
  XOR U22811 ( .A(n21344), .B(n21342), .Z(n21343) );
  XNOR U22812 ( .A(n21345), .B(n21346), .Z(n21333) );
  AND U22813 ( .A(n21347), .B(n21348), .Z(n21345) );
  XNOR U22814 ( .A(n21346), .B(n21275), .Z(n21348) );
  XOR U22815 ( .A(n21339), .B(n21340), .Z(n21275) );
  XNOR U22816 ( .A(n21349), .B(n21350), .Z(n21340) );
  ANDN U22817 ( .B(n21351), .A(n21352), .Z(n21349) );
  XOR U22818 ( .A(n21353), .B(n21354), .Z(n21351) );
  XOR U22819 ( .A(n21355), .B(n21356), .Z(n21339) );
  XNOR U22820 ( .A(n21357), .B(n21358), .Z(n21356) );
  ANDN U22821 ( .B(n21359), .A(n21360), .Z(n21357) );
  XNOR U22822 ( .A(n21361), .B(n21362), .Z(n21359) );
  IV U22823 ( .A(n21337), .Z(n21355) );
  XOR U22824 ( .A(n21363), .B(n21364), .Z(n21337) );
  ANDN U22825 ( .B(n21365), .A(n21366), .Z(n21363) );
  XOR U22826 ( .A(n21364), .B(n21367), .Z(n21365) );
  XOR U22827 ( .A(n21346), .B(n21277), .Z(n21347) );
  XOR U22828 ( .A(n21368), .B(n21369), .Z(n21277) );
  AND U22829 ( .A(n414), .B(n21370), .Z(n21368) );
  XOR U22830 ( .A(n21371), .B(n21369), .Z(n21370) );
  XNOR U22831 ( .A(n21372), .B(n21373), .Z(n21346) );
  NAND U22832 ( .A(n21374), .B(n21375), .Z(n21373) );
  XOR U22833 ( .A(n21376), .B(n21325), .Z(n21375) );
  XOR U22834 ( .A(n21366), .B(n21367), .Z(n21325) );
  XOR U22835 ( .A(n21377), .B(n21354), .Z(n21367) );
  XOR U22836 ( .A(n21378), .B(n21379), .Z(n21354) );
  ANDN U22837 ( .B(n21380), .A(n21381), .Z(n21378) );
  XOR U22838 ( .A(n21379), .B(n21382), .Z(n21380) );
  IV U22839 ( .A(n21352), .Z(n21377) );
  XOR U22840 ( .A(n21350), .B(n21383), .Z(n21352) );
  XOR U22841 ( .A(n21384), .B(n21385), .Z(n21383) );
  ANDN U22842 ( .B(n21386), .A(n21387), .Z(n21384) );
  XOR U22843 ( .A(n21388), .B(n21385), .Z(n21386) );
  IV U22844 ( .A(n21353), .Z(n21350) );
  XOR U22845 ( .A(n21389), .B(n21390), .Z(n21353) );
  ANDN U22846 ( .B(n21391), .A(n21392), .Z(n21389) );
  XOR U22847 ( .A(n21390), .B(n21393), .Z(n21391) );
  XOR U22848 ( .A(n21394), .B(n21395), .Z(n21366) );
  XNOR U22849 ( .A(n21361), .B(n21396), .Z(n21395) );
  IV U22850 ( .A(n21364), .Z(n21396) );
  XOR U22851 ( .A(n21397), .B(n21398), .Z(n21364) );
  ANDN U22852 ( .B(n21399), .A(n21400), .Z(n21397) );
  XOR U22853 ( .A(n21398), .B(n21401), .Z(n21399) );
  XNOR U22854 ( .A(n21402), .B(n21403), .Z(n21361) );
  ANDN U22855 ( .B(n21404), .A(n21405), .Z(n21402) );
  XOR U22856 ( .A(n21403), .B(n21406), .Z(n21404) );
  IV U22857 ( .A(n21360), .Z(n21394) );
  XOR U22858 ( .A(n21358), .B(n21407), .Z(n21360) );
  XOR U22859 ( .A(n21408), .B(n21409), .Z(n21407) );
  ANDN U22860 ( .B(n21410), .A(n21411), .Z(n21408) );
  XOR U22861 ( .A(n21412), .B(n21409), .Z(n21410) );
  IV U22862 ( .A(n21362), .Z(n21358) );
  XOR U22863 ( .A(n21413), .B(n21414), .Z(n21362) );
  ANDN U22864 ( .B(n21415), .A(n21416), .Z(n21413) );
  XOR U22865 ( .A(n21417), .B(n21414), .Z(n21415) );
  IV U22866 ( .A(n21372), .Z(n21376) );
  XOR U22867 ( .A(n21372), .B(n21327), .Z(n21374) );
  XOR U22868 ( .A(n21418), .B(n21419), .Z(n21327) );
  AND U22869 ( .A(n414), .B(n21420), .Z(n21418) );
  XOR U22870 ( .A(n21421), .B(n21419), .Z(n21420) );
  NANDN U22871 ( .A(n21329), .B(n21331), .Z(n21372) );
  XOR U22872 ( .A(n21422), .B(n21423), .Z(n21331) );
  AND U22873 ( .A(n414), .B(n21424), .Z(n21422) );
  XOR U22874 ( .A(n21423), .B(n21425), .Z(n21424) );
  XNOR U22875 ( .A(n21426), .B(n21427), .Z(n414) );
  AND U22876 ( .A(n21428), .B(n21429), .Z(n21426) );
  XOR U22877 ( .A(n21427), .B(n21342), .Z(n21429) );
  XNOR U22878 ( .A(n21430), .B(n21431), .Z(n21342) );
  ANDN U22879 ( .B(n21432), .A(n21433), .Z(n21430) );
  XOR U22880 ( .A(n21431), .B(n21434), .Z(n21432) );
  XNOR U22881 ( .A(n21427), .B(n21344), .Z(n21428) );
  XOR U22882 ( .A(n21435), .B(n21436), .Z(n21344) );
  AND U22883 ( .A(n418), .B(n21437), .Z(n21435) );
  XOR U22884 ( .A(n21438), .B(n21436), .Z(n21437) );
  XNOR U22885 ( .A(n21439), .B(n21440), .Z(n21427) );
  AND U22886 ( .A(n21441), .B(n21442), .Z(n21439) );
  XNOR U22887 ( .A(n21440), .B(n21369), .Z(n21442) );
  XOR U22888 ( .A(n21433), .B(n21434), .Z(n21369) );
  XNOR U22889 ( .A(n21443), .B(n21444), .Z(n21434) );
  ANDN U22890 ( .B(n21445), .A(n21446), .Z(n21443) );
  XOR U22891 ( .A(n21447), .B(n21448), .Z(n21445) );
  XOR U22892 ( .A(n21449), .B(n21450), .Z(n21433) );
  XNOR U22893 ( .A(n21451), .B(n21452), .Z(n21450) );
  ANDN U22894 ( .B(n21453), .A(n21454), .Z(n21451) );
  XNOR U22895 ( .A(n21455), .B(n21456), .Z(n21453) );
  IV U22896 ( .A(n21431), .Z(n21449) );
  XOR U22897 ( .A(n21457), .B(n21458), .Z(n21431) );
  ANDN U22898 ( .B(n21459), .A(n21460), .Z(n21457) );
  XOR U22899 ( .A(n21458), .B(n21461), .Z(n21459) );
  XOR U22900 ( .A(n21440), .B(n21371), .Z(n21441) );
  XOR U22901 ( .A(n21462), .B(n21463), .Z(n21371) );
  AND U22902 ( .A(n418), .B(n21464), .Z(n21462) );
  XOR U22903 ( .A(n21465), .B(n21463), .Z(n21464) );
  XNOR U22904 ( .A(n21466), .B(n21467), .Z(n21440) );
  NAND U22905 ( .A(n21468), .B(n21469), .Z(n21467) );
  XOR U22906 ( .A(n21470), .B(n21419), .Z(n21469) );
  XOR U22907 ( .A(n21460), .B(n21461), .Z(n21419) );
  XOR U22908 ( .A(n21471), .B(n21448), .Z(n21461) );
  XOR U22909 ( .A(n21472), .B(n21473), .Z(n21448) );
  ANDN U22910 ( .B(n21474), .A(n21475), .Z(n21472) );
  XOR U22911 ( .A(n21473), .B(n21476), .Z(n21474) );
  IV U22912 ( .A(n21446), .Z(n21471) );
  XOR U22913 ( .A(n21444), .B(n21477), .Z(n21446) );
  XOR U22914 ( .A(n21478), .B(n21479), .Z(n21477) );
  ANDN U22915 ( .B(n21480), .A(n21481), .Z(n21478) );
  XOR U22916 ( .A(n21482), .B(n21479), .Z(n21480) );
  IV U22917 ( .A(n21447), .Z(n21444) );
  XOR U22918 ( .A(n21483), .B(n21484), .Z(n21447) );
  ANDN U22919 ( .B(n21485), .A(n21486), .Z(n21483) );
  XOR U22920 ( .A(n21484), .B(n21487), .Z(n21485) );
  XOR U22921 ( .A(n21488), .B(n21489), .Z(n21460) );
  XNOR U22922 ( .A(n21455), .B(n21490), .Z(n21489) );
  IV U22923 ( .A(n21458), .Z(n21490) );
  XOR U22924 ( .A(n21491), .B(n21492), .Z(n21458) );
  ANDN U22925 ( .B(n21493), .A(n21494), .Z(n21491) );
  XOR U22926 ( .A(n21492), .B(n21495), .Z(n21493) );
  XNOR U22927 ( .A(n21496), .B(n21497), .Z(n21455) );
  ANDN U22928 ( .B(n21498), .A(n21499), .Z(n21496) );
  XOR U22929 ( .A(n21497), .B(n21500), .Z(n21498) );
  IV U22930 ( .A(n21454), .Z(n21488) );
  XOR U22931 ( .A(n21452), .B(n21501), .Z(n21454) );
  XOR U22932 ( .A(n21502), .B(n21503), .Z(n21501) );
  ANDN U22933 ( .B(n21504), .A(n21505), .Z(n21502) );
  XOR U22934 ( .A(n21506), .B(n21503), .Z(n21504) );
  IV U22935 ( .A(n21456), .Z(n21452) );
  XOR U22936 ( .A(n21507), .B(n21508), .Z(n21456) );
  ANDN U22937 ( .B(n21509), .A(n21510), .Z(n21507) );
  XOR U22938 ( .A(n21511), .B(n21508), .Z(n21509) );
  IV U22939 ( .A(n21466), .Z(n21470) );
  XOR U22940 ( .A(n21466), .B(n21421), .Z(n21468) );
  XOR U22941 ( .A(n21512), .B(n21513), .Z(n21421) );
  AND U22942 ( .A(n418), .B(n21514), .Z(n21512) );
  XOR U22943 ( .A(n21515), .B(n21513), .Z(n21514) );
  NANDN U22944 ( .A(n21423), .B(n21425), .Z(n21466) );
  XOR U22945 ( .A(n21516), .B(n21517), .Z(n21425) );
  AND U22946 ( .A(n418), .B(n21518), .Z(n21516) );
  XOR U22947 ( .A(n21517), .B(n21519), .Z(n21518) );
  XNOR U22948 ( .A(n21520), .B(n21521), .Z(n418) );
  AND U22949 ( .A(n21522), .B(n21523), .Z(n21520) );
  XOR U22950 ( .A(n21521), .B(n21436), .Z(n21523) );
  XNOR U22951 ( .A(n21524), .B(n21525), .Z(n21436) );
  ANDN U22952 ( .B(n21526), .A(n21527), .Z(n21524) );
  XOR U22953 ( .A(n21525), .B(n21528), .Z(n21526) );
  XNOR U22954 ( .A(n21521), .B(n21438), .Z(n21522) );
  XOR U22955 ( .A(n21529), .B(n21530), .Z(n21438) );
  AND U22956 ( .A(n422), .B(n21531), .Z(n21529) );
  XOR U22957 ( .A(n21532), .B(n21530), .Z(n21531) );
  XNOR U22958 ( .A(n21533), .B(n21534), .Z(n21521) );
  AND U22959 ( .A(n21535), .B(n21536), .Z(n21533) );
  XNOR U22960 ( .A(n21534), .B(n21463), .Z(n21536) );
  XOR U22961 ( .A(n21527), .B(n21528), .Z(n21463) );
  XNOR U22962 ( .A(n21537), .B(n21538), .Z(n21528) );
  ANDN U22963 ( .B(n21539), .A(n21540), .Z(n21537) );
  XOR U22964 ( .A(n21541), .B(n21542), .Z(n21539) );
  XOR U22965 ( .A(n21543), .B(n21544), .Z(n21527) );
  XNOR U22966 ( .A(n21545), .B(n21546), .Z(n21544) );
  ANDN U22967 ( .B(n21547), .A(n21548), .Z(n21545) );
  XNOR U22968 ( .A(n21549), .B(n21550), .Z(n21547) );
  IV U22969 ( .A(n21525), .Z(n21543) );
  XOR U22970 ( .A(n21551), .B(n21552), .Z(n21525) );
  ANDN U22971 ( .B(n21553), .A(n21554), .Z(n21551) );
  XOR U22972 ( .A(n21552), .B(n21555), .Z(n21553) );
  XOR U22973 ( .A(n21534), .B(n21465), .Z(n21535) );
  XOR U22974 ( .A(n21556), .B(n21557), .Z(n21465) );
  AND U22975 ( .A(n422), .B(n21558), .Z(n21556) );
  XOR U22976 ( .A(n21559), .B(n21557), .Z(n21558) );
  XNOR U22977 ( .A(n21560), .B(n21561), .Z(n21534) );
  NAND U22978 ( .A(n21562), .B(n21563), .Z(n21561) );
  XOR U22979 ( .A(n21564), .B(n21513), .Z(n21563) );
  XOR U22980 ( .A(n21554), .B(n21555), .Z(n21513) );
  XOR U22981 ( .A(n21565), .B(n21542), .Z(n21555) );
  XOR U22982 ( .A(n21566), .B(n21567), .Z(n21542) );
  ANDN U22983 ( .B(n21568), .A(n21569), .Z(n21566) );
  XOR U22984 ( .A(n21567), .B(n21570), .Z(n21568) );
  IV U22985 ( .A(n21540), .Z(n21565) );
  XOR U22986 ( .A(n21538), .B(n21571), .Z(n21540) );
  XOR U22987 ( .A(n21572), .B(n21573), .Z(n21571) );
  ANDN U22988 ( .B(n21574), .A(n21575), .Z(n21572) );
  XOR U22989 ( .A(n21576), .B(n21573), .Z(n21574) );
  IV U22990 ( .A(n21541), .Z(n21538) );
  XOR U22991 ( .A(n21577), .B(n21578), .Z(n21541) );
  ANDN U22992 ( .B(n21579), .A(n21580), .Z(n21577) );
  XOR U22993 ( .A(n21578), .B(n21581), .Z(n21579) );
  XOR U22994 ( .A(n21582), .B(n21583), .Z(n21554) );
  XNOR U22995 ( .A(n21549), .B(n21584), .Z(n21583) );
  IV U22996 ( .A(n21552), .Z(n21584) );
  XOR U22997 ( .A(n21585), .B(n21586), .Z(n21552) );
  ANDN U22998 ( .B(n21587), .A(n21588), .Z(n21585) );
  XOR U22999 ( .A(n21586), .B(n21589), .Z(n21587) );
  XNOR U23000 ( .A(n21590), .B(n21591), .Z(n21549) );
  ANDN U23001 ( .B(n21592), .A(n21593), .Z(n21590) );
  XOR U23002 ( .A(n21591), .B(n21594), .Z(n21592) );
  IV U23003 ( .A(n21548), .Z(n21582) );
  XOR U23004 ( .A(n21546), .B(n21595), .Z(n21548) );
  XOR U23005 ( .A(n21596), .B(n21597), .Z(n21595) );
  ANDN U23006 ( .B(n21598), .A(n21599), .Z(n21596) );
  XOR U23007 ( .A(n21600), .B(n21597), .Z(n21598) );
  IV U23008 ( .A(n21550), .Z(n21546) );
  XOR U23009 ( .A(n21601), .B(n21602), .Z(n21550) );
  ANDN U23010 ( .B(n21603), .A(n21604), .Z(n21601) );
  XOR U23011 ( .A(n21605), .B(n21602), .Z(n21603) );
  IV U23012 ( .A(n21560), .Z(n21564) );
  XOR U23013 ( .A(n21560), .B(n21515), .Z(n21562) );
  XOR U23014 ( .A(n21606), .B(n21607), .Z(n21515) );
  AND U23015 ( .A(n422), .B(n21608), .Z(n21606) );
  XOR U23016 ( .A(n21609), .B(n21607), .Z(n21608) );
  NANDN U23017 ( .A(n21517), .B(n21519), .Z(n21560) );
  XOR U23018 ( .A(n21610), .B(n21611), .Z(n21519) );
  AND U23019 ( .A(n422), .B(n21612), .Z(n21610) );
  XOR U23020 ( .A(n21611), .B(n21613), .Z(n21612) );
  XNOR U23021 ( .A(n21614), .B(n21615), .Z(n422) );
  AND U23022 ( .A(n21616), .B(n21617), .Z(n21614) );
  XOR U23023 ( .A(n21615), .B(n21530), .Z(n21617) );
  XNOR U23024 ( .A(n21618), .B(n21619), .Z(n21530) );
  ANDN U23025 ( .B(n21620), .A(n21621), .Z(n21618) );
  XOR U23026 ( .A(n21619), .B(n21622), .Z(n21620) );
  XNOR U23027 ( .A(n21615), .B(n21532), .Z(n21616) );
  XOR U23028 ( .A(n21623), .B(n21624), .Z(n21532) );
  AND U23029 ( .A(n426), .B(n21625), .Z(n21623) );
  XOR U23030 ( .A(n21626), .B(n21624), .Z(n21625) );
  XNOR U23031 ( .A(n21627), .B(n21628), .Z(n21615) );
  AND U23032 ( .A(n21629), .B(n21630), .Z(n21627) );
  XNOR U23033 ( .A(n21628), .B(n21557), .Z(n21630) );
  XOR U23034 ( .A(n21621), .B(n21622), .Z(n21557) );
  XNOR U23035 ( .A(n21631), .B(n21632), .Z(n21622) );
  ANDN U23036 ( .B(n21633), .A(n21634), .Z(n21631) );
  XOR U23037 ( .A(n21635), .B(n21636), .Z(n21633) );
  XOR U23038 ( .A(n21637), .B(n21638), .Z(n21621) );
  XNOR U23039 ( .A(n21639), .B(n21640), .Z(n21638) );
  ANDN U23040 ( .B(n21641), .A(n21642), .Z(n21639) );
  XNOR U23041 ( .A(n21643), .B(n21644), .Z(n21641) );
  IV U23042 ( .A(n21619), .Z(n21637) );
  XOR U23043 ( .A(n21645), .B(n21646), .Z(n21619) );
  ANDN U23044 ( .B(n21647), .A(n21648), .Z(n21645) );
  XOR U23045 ( .A(n21646), .B(n21649), .Z(n21647) );
  XOR U23046 ( .A(n21628), .B(n21559), .Z(n21629) );
  XOR U23047 ( .A(n21650), .B(n21651), .Z(n21559) );
  AND U23048 ( .A(n426), .B(n21652), .Z(n21650) );
  XOR U23049 ( .A(n21653), .B(n21651), .Z(n21652) );
  XNOR U23050 ( .A(n21654), .B(n21655), .Z(n21628) );
  NAND U23051 ( .A(n21656), .B(n21657), .Z(n21655) );
  XOR U23052 ( .A(n21658), .B(n21607), .Z(n21657) );
  XOR U23053 ( .A(n21648), .B(n21649), .Z(n21607) );
  XOR U23054 ( .A(n21659), .B(n21636), .Z(n21649) );
  XOR U23055 ( .A(n21660), .B(n21661), .Z(n21636) );
  ANDN U23056 ( .B(n21662), .A(n21663), .Z(n21660) );
  XOR U23057 ( .A(n21661), .B(n21664), .Z(n21662) );
  IV U23058 ( .A(n21634), .Z(n21659) );
  XOR U23059 ( .A(n21632), .B(n21665), .Z(n21634) );
  XOR U23060 ( .A(n21666), .B(n21667), .Z(n21665) );
  ANDN U23061 ( .B(n21668), .A(n21669), .Z(n21666) );
  XOR U23062 ( .A(n21670), .B(n21667), .Z(n21668) );
  IV U23063 ( .A(n21635), .Z(n21632) );
  XOR U23064 ( .A(n21671), .B(n21672), .Z(n21635) );
  ANDN U23065 ( .B(n21673), .A(n21674), .Z(n21671) );
  XOR U23066 ( .A(n21672), .B(n21675), .Z(n21673) );
  XOR U23067 ( .A(n21676), .B(n21677), .Z(n21648) );
  XNOR U23068 ( .A(n21643), .B(n21678), .Z(n21677) );
  IV U23069 ( .A(n21646), .Z(n21678) );
  XOR U23070 ( .A(n21679), .B(n21680), .Z(n21646) );
  ANDN U23071 ( .B(n21681), .A(n21682), .Z(n21679) );
  XOR U23072 ( .A(n21680), .B(n21683), .Z(n21681) );
  XNOR U23073 ( .A(n21684), .B(n21685), .Z(n21643) );
  ANDN U23074 ( .B(n21686), .A(n21687), .Z(n21684) );
  XOR U23075 ( .A(n21685), .B(n21688), .Z(n21686) );
  IV U23076 ( .A(n21642), .Z(n21676) );
  XOR U23077 ( .A(n21640), .B(n21689), .Z(n21642) );
  XOR U23078 ( .A(n21690), .B(n21691), .Z(n21689) );
  ANDN U23079 ( .B(n21692), .A(n21693), .Z(n21690) );
  XOR U23080 ( .A(n21694), .B(n21691), .Z(n21692) );
  IV U23081 ( .A(n21644), .Z(n21640) );
  XOR U23082 ( .A(n21695), .B(n21696), .Z(n21644) );
  ANDN U23083 ( .B(n21697), .A(n21698), .Z(n21695) );
  XOR U23084 ( .A(n21699), .B(n21696), .Z(n21697) );
  IV U23085 ( .A(n21654), .Z(n21658) );
  XOR U23086 ( .A(n21654), .B(n21609), .Z(n21656) );
  XOR U23087 ( .A(n21700), .B(n21701), .Z(n21609) );
  AND U23088 ( .A(n426), .B(n21702), .Z(n21700) );
  XOR U23089 ( .A(n21703), .B(n21701), .Z(n21702) );
  NANDN U23090 ( .A(n21611), .B(n21613), .Z(n21654) );
  XOR U23091 ( .A(n21704), .B(n21705), .Z(n21613) );
  AND U23092 ( .A(n426), .B(n21706), .Z(n21704) );
  XOR U23093 ( .A(n21705), .B(n21707), .Z(n21706) );
  XNOR U23094 ( .A(n21708), .B(n21709), .Z(n426) );
  AND U23095 ( .A(n21710), .B(n21711), .Z(n21708) );
  XOR U23096 ( .A(n21709), .B(n21624), .Z(n21711) );
  XNOR U23097 ( .A(n21712), .B(n21713), .Z(n21624) );
  ANDN U23098 ( .B(n21714), .A(n21715), .Z(n21712) );
  XOR U23099 ( .A(n21713), .B(n21716), .Z(n21714) );
  XNOR U23100 ( .A(n21709), .B(n21626), .Z(n21710) );
  XOR U23101 ( .A(n21717), .B(n21718), .Z(n21626) );
  AND U23102 ( .A(n430), .B(n21719), .Z(n21717) );
  XOR U23103 ( .A(n21720), .B(n21718), .Z(n21719) );
  XNOR U23104 ( .A(n21721), .B(n21722), .Z(n21709) );
  AND U23105 ( .A(n21723), .B(n21724), .Z(n21721) );
  XNOR U23106 ( .A(n21722), .B(n21651), .Z(n21724) );
  XOR U23107 ( .A(n21715), .B(n21716), .Z(n21651) );
  XNOR U23108 ( .A(n21725), .B(n21726), .Z(n21716) );
  ANDN U23109 ( .B(n21727), .A(n21728), .Z(n21725) );
  XOR U23110 ( .A(n21729), .B(n21730), .Z(n21727) );
  XOR U23111 ( .A(n21731), .B(n21732), .Z(n21715) );
  XNOR U23112 ( .A(n21733), .B(n21734), .Z(n21732) );
  ANDN U23113 ( .B(n21735), .A(n21736), .Z(n21733) );
  XNOR U23114 ( .A(n21737), .B(n21738), .Z(n21735) );
  IV U23115 ( .A(n21713), .Z(n21731) );
  XOR U23116 ( .A(n21739), .B(n21740), .Z(n21713) );
  ANDN U23117 ( .B(n21741), .A(n21742), .Z(n21739) );
  XOR U23118 ( .A(n21740), .B(n21743), .Z(n21741) );
  XOR U23119 ( .A(n21722), .B(n21653), .Z(n21723) );
  XOR U23120 ( .A(n21744), .B(n21745), .Z(n21653) );
  AND U23121 ( .A(n430), .B(n21746), .Z(n21744) );
  XOR U23122 ( .A(n21747), .B(n21745), .Z(n21746) );
  XNOR U23123 ( .A(n21748), .B(n21749), .Z(n21722) );
  NAND U23124 ( .A(n21750), .B(n21751), .Z(n21749) );
  XOR U23125 ( .A(n21752), .B(n21701), .Z(n21751) );
  XOR U23126 ( .A(n21742), .B(n21743), .Z(n21701) );
  XOR U23127 ( .A(n21753), .B(n21730), .Z(n21743) );
  XOR U23128 ( .A(n21754), .B(n21755), .Z(n21730) );
  ANDN U23129 ( .B(n21756), .A(n21757), .Z(n21754) );
  XOR U23130 ( .A(n21755), .B(n21758), .Z(n21756) );
  IV U23131 ( .A(n21728), .Z(n21753) );
  XOR U23132 ( .A(n21726), .B(n21759), .Z(n21728) );
  XOR U23133 ( .A(n21760), .B(n21761), .Z(n21759) );
  ANDN U23134 ( .B(n21762), .A(n21763), .Z(n21760) );
  XOR U23135 ( .A(n21764), .B(n21761), .Z(n21762) );
  IV U23136 ( .A(n21729), .Z(n21726) );
  XOR U23137 ( .A(n21765), .B(n21766), .Z(n21729) );
  ANDN U23138 ( .B(n21767), .A(n21768), .Z(n21765) );
  XOR U23139 ( .A(n21766), .B(n21769), .Z(n21767) );
  XOR U23140 ( .A(n21770), .B(n21771), .Z(n21742) );
  XNOR U23141 ( .A(n21737), .B(n21772), .Z(n21771) );
  IV U23142 ( .A(n21740), .Z(n21772) );
  XOR U23143 ( .A(n21773), .B(n21774), .Z(n21740) );
  ANDN U23144 ( .B(n21775), .A(n21776), .Z(n21773) );
  XOR U23145 ( .A(n21774), .B(n21777), .Z(n21775) );
  XNOR U23146 ( .A(n21778), .B(n21779), .Z(n21737) );
  ANDN U23147 ( .B(n21780), .A(n21781), .Z(n21778) );
  XOR U23148 ( .A(n21779), .B(n21782), .Z(n21780) );
  IV U23149 ( .A(n21736), .Z(n21770) );
  XOR U23150 ( .A(n21734), .B(n21783), .Z(n21736) );
  XOR U23151 ( .A(n21784), .B(n21785), .Z(n21783) );
  ANDN U23152 ( .B(n21786), .A(n21787), .Z(n21784) );
  XOR U23153 ( .A(n21788), .B(n21785), .Z(n21786) );
  IV U23154 ( .A(n21738), .Z(n21734) );
  XOR U23155 ( .A(n21789), .B(n21790), .Z(n21738) );
  ANDN U23156 ( .B(n21791), .A(n21792), .Z(n21789) );
  XOR U23157 ( .A(n21793), .B(n21790), .Z(n21791) );
  IV U23158 ( .A(n21748), .Z(n21752) );
  XOR U23159 ( .A(n21748), .B(n21703), .Z(n21750) );
  XOR U23160 ( .A(n21794), .B(n21795), .Z(n21703) );
  AND U23161 ( .A(n430), .B(n21796), .Z(n21794) );
  XOR U23162 ( .A(n21797), .B(n21795), .Z(n21796) );
  NANDN U23163 ( .A(n21705), .B(n21707), .Z(n21748) );
  XOR U23164 ( .A(n21798), .B(n21799), .Z(n21707) );
  AND U23165 ( .A(n430), .B(n21800), .Z(n21798) );
  XOR U23166 ( .A(n21799), .B(n21801), .Z(n21800) );
  XNOR U23167 ( .A(n21802), .B(n21803), .Z(n430) );
  AND U23168 ( .A(n21804), .B(n21805), .Z(n21802) );
  XOR U23169 ( .A(n21803), .B(n21718), .Z(n21805) );
  XNOR U23170 ( .A(n21806), .B(n21807), .Z(n21718) );
  ANDN U23171 ( .B(n21808), .A(n21809), .Z(n21806) );
  XOR U23172 ( .A(n21807), .B(n21810), .Z(n21808) );
  XNOR U23173 ( .A(n21803), .B(n21720), .Z(n21804) );
  XOR U23174 ( .A(n21811), .B(n21812), .Z(n21720) );
  AND U23175 ( .A(n434), .B(n21813), .Z(n21811) );
  XOR U23176 ( .A(n21814), .B(n21812), .Z(n21813) );
  XNOR U23177 ( .A(n21815), .B(n21816), .Z(n21803) );
  AND U23178 ( .A(n21817), .B(n21818), .Z(n21815) );
  XNOR U23179 ( .A(n21816), .B(n21745), .Z(n21818) );
  XOR U23180 ( .A(n21809), .B(n21810), .Z(n21745) );
  XNOR U23181 ( .A(n21819), .B(n21820), .Z(n21810) );
  ANDN U23182 ( .B(n21821), .A(n21822), .Z(n21819) );
  XOR U23183 ( .A(n21823), .B(n21824), .Z(n21821) );
  XOR U23184 ( .A(n21825), .B(n21826), .Z(n21809) );
  XNOR U23185 ( .A(n21827), .B(n21828), .Z(n21826) );
  ANDN U23186 ( .B(n21829), .A(n21830), .Z(n21827) );
  XNOR U23187 ( .A(n21831), .B(n21832), .Z(n21829) );
  IV U23188 ( .A(n21807), .Z(n21825) );
  XOR U23189 ( .A(n21833), .B(n21834), .Z(n21807) );
  ANDN U23190 ( .B(n21835), .A(n21836), .Z(n21833) );
  XOR U23191 ( .A(n21834), .B(n21837), .Z(n21835) );
  XOR U23192 ( .A(n21816), .B(n21747), .Z(n21817) );
  XOR U23193 ( .A(n21838), .B(n21839), .Z(n21747) );
  AND U23194 ( .A(n434), .B(n21840), .Z(n21838) );
  XOR U23195 ( .A(n21841), .B(n21839), .Z(n21840) );
  XNOR U23196 ( .A(n21842), .B(n21843), .Z(n21816) );
  NAND U23197 ( .A(n21844), .B(n21845), .Z(n21843) );
  XOR U23198 ( .A(n21846), .B(n21795), .Z(n21845) );
  XOR U23199 ( .A(n21836), .B(n21837), .Z(n21795) );
  XOR U23200 ( .A(n21847), .B(n21824), .Z(n21837) );
  XOR U23201 ( .A(n21848), .B(n21849), .Z(n21824) );
  ANDN U23202 ( .B(n21850), .A(n21851), .Z(n21848) );
  XOR U23203 ( .A(n21849), .B(n21852), .Z(n21850) );
  IV U23204 ( .A(n21822), .Z(n21847) );
  XOR U23205 ( .A(n21820), .B(n21853), .Z(n21822) );
  XOR U23206 ( .A(n21854), .B(n21855), .Z(n21853) );
  ANDN U23207 ( .B(n21856), .A(n21857), .Z(n21854) );
  XOR U23208 ( .A(n21858), .B(n21855), .Z(n21856) );
  IV U23209 ( .A(n21823), .Z(n21820) );
  XOR U23210 ( .A(n21859), .B(n21860), .Z(n21823) );
  ANDN U23211 ( .B(n21861), .A(n21862), .Z(n21859) );
  XOR U23212 ( .A(n21860), .B(n21863), .Z(n21861) );
  XOR U23213 ( .A(n21864), .B(n21865), .Z(n21836) );
  XNOR U23214 ( .A(n21831), .B(n21866), .Z(n21865) );
  IV U23215 ( .A(n21834), .Z(n21866) );
  XOR U23216 ( .A(n21867), .B(n21868), .Z(n21834) );
  ANDN U23217 ( .B(n21869), .A(n21870), .Z(n21867) );
  XOR U23218 ( .A(n21868), .B(n21871), .Z(n21869) );
  XNOR U23219 ( .A(n21872), .B(n21873), .Z(n21831) );
  ANDN U23220 ( .B(n21874), .A(n21875), .Z(n21872) );
  XOR U23221 ( .A(n21873), .B(n21876), .Z(n21874) );
  IV U23222 ( .A(n21830), .Z(n21864) );
  XOR U23223 ( .A(n21828), .B(n21877), .Z(n21830) );
  XOR U23224 ( .A(n21878), .B(n21879), .Z(n21877) );
  ANDN U23225 ( .B(n21880), .A(n21881), .Z(n21878) );
  XOR U23226 ( .A(n21882), .B(n21879), .Z(n21880) );
  IV U23227 ( .A(n21832), .Z(n21828) );
  XOR U23228 ( .A(n21883), .B(n21884), .Z(n21832) );
  ANDN U23229 ( .B(n21885), .A(n21886), .Z(n21883) );
  XOR U23230 ( .A(n21887), .B(n21884), .Z(n21885) );
  IV U23231 ( .A(n21842), .Z(n21846) );
  XOR U23232 ( .A(n21842), .B(n21797), .Z(n21844) );
  XOR U23233 ( .A(n21888), .B(n21889), .Z(n21797) );
  AND U23234 ( .A(n434), .B(n21890), .Z(n21888) );
  XOR U23235 ( .A(n21891), .B(n21889), .Z(n21890) );
  NANDN U23236 ( .A(n21799), .B(n21801), .Z(n21842) );
  XOR U23237 ( .A(n21892), .B(n21893), .Z(n21801) );
  AND U23238 ( .A(n434), .B(n21894), .Z(n21892) );
  XOR U23239 ( .A(n21893), .B(n21895), .Z(n21894) );
  XNOR U23240 ( .A(n21896), .B(n21897), .Z(n434) );
  AND U23241 ( .A(n21898), .B(n21899), .Z(n21896) );
  XOR U23242 ( .A(n21897), .B(n21812), .Z(n21899) );
  XNOR U23243 ( .A(n21900), .B(n21901), .Z(n21812) );
  ANDN U23244 ( .B(n21902), .A(n21903), .Z(n21900) );
  XOR U23245 ( .A(n21901), .B(n21904), .Z(n21902) );
  XNOR U23246 ( .A(n21897), .B(n21814), .Z(n21898) );
  XOR U23247 ( .A(n21905), .B(n21906), .Z(n21814) );
  AND U23248 ( .A(n438), .B(n21907), .Z(n21905) );
  XOR U23249 ( .A(n21908), .B(n21906), .Z(n21907) );
  XNOR U23250 ( .A(n21909), .B(n21910), .Z(n21897) );
  AND U23251 ( .A(n21911), .B(n21912), .Z(n21909) );
  XNOR U23252 ( .A(n21910), .B(n21839), .Z(n21912) );
  XOR U23253 ( .A(n21903), .B(n21904), .Z(n21839) );
  XNOR U23254 ( .A(n21913), .B(n21914), .Z(n21904) );
  ANDN U23255 ( .B(n21915), .A(n21916), .Z(n21913) );
  XOR U23256 ( .A(n21917), .B(n21918), .Z(n21915) );
  XOR U23257 ( .A(n21919), .B(n21920), .Z(n21903) );
  XNOR U23258 ( .A(n21921), .B(n21922), .Z(n21920) );
  ANDN U23259 ( .B(n21923), .A(n21924), .Z(n21921) );
  XNOR U23260 ( .A(n21925), .B(n21926), .Z(n21923) );
  IV U23261 ( .A(n21901), .Z(n21919) );
  XOR U23262 ( .A(n21927), .B(n21928), .Z(n21901) );
  ANDN U23263 ( .B(n21929), .A(n21930), .Z(n21927) );
  XOR U23264 ( .A(n21928), .B(n21931), .Z(n21929) );
  XOR U23265 ( .A(n21910), .B(n21841), .Z(n21911) );
  XOR U23266 ( .A(n21932), .B(n21933), .Z(n21841) );
  AND U23267 ( .A(n438), .B(n21934), .Z(n21932) );
  XOR U23268 ( .A(n21935), .B(n21933), .Z(n21934) );
  XNOR U23269 ( .A(n21936), .B(n21937), .Z(n21910) );
  NAND U23270 ( .A(n21938), .B(n21939), .Z(n21937) );
  XOR U23271 ( .A(n21940), .B(n21889), .Z(n21939) );
  XOR U23272 ( .A(n21930), .B(n21931), .Z(n21889) );
  XOR U23273 ( .A(n21941), .B(n21918), .Z(n21931) );
  XOR U23274 ( .A(n21942), .B(n21943), .Z(n21918) );
  ANDN U23275 ( .B(n21944), .A(n21945), .Z(n21942) );
  XOR U23276 ( .A(n21943), .B(n21946), .Z(n21944) );
  IV U23277 ( .A(n21916), .Z(n21941) );
  XOR U23278 ( .A(n21914), .B(n21947), .Z(n21916) );
  XOR U23279 ( .A(n21948), .B(n21949), .Z(n21947) );
  ANDN U23280 ( .B(n21950), .A(n21951), .Z(n21948) );
  XOR U23281 ( .A(n21952), .B(n21949), .Z(n21950) );
  IV U23282 ( .A(n21917), .Z(n21914) );
  XOR U23283 ( .A(n21953), .B(n21954), .Z(n21917) );
  ANDN U23284 ( .B(n21955), .A(n21956), .Z(n21953) );
  XOR U23285 ( .A(n21954), .B(n21957), .Z(n21955) );
  XOR U23286 ( .A(n21958), .B(n21959), .Z(n21930) );
  XNOR U23287 ( .A(n21925), .B(n21960), .Z(n21959) );
  IV U23288 ( .A(n21928), .Z(n21960) );
  XOR U23289 ( .A(n21961), .B(n21962), .Z(n21928) );
  ANDN U23290 ( .B(n21963), .A(n21964), .Z(n21961) );
  XOR U23291 ( .A(n21962), .B(n21965), .Z(n21963) );
  XNOR U23292 ( .A(n21966), .B(n21967), .Z(n21925) );
  ANDN U23293 ( .B(n21968), .A(n21969), .Z(n21966) );
  XOR U23294 ( .A(n21967), .B(n21970), .Z(n21968) );
  IV U23295 ( .A(n21924), .Z(n21958) );
  XOR U23296 ( .A(n21922), .B(n21971), .Z(n21924) );
  XOR U23297 ( .A(n21972), .B(n21973), .Z(n21971) );
  ANDN U23298 ( .B(n21974), .A(n21975), .Z(n21972) );
  XOR U23299 ( .A(n21976), .B(n21973), .Z(n21974) );
  IV U23300 ( .A(n21926), .Z(n21922) );
  XOR U23301 ( .A(n21977), .B(n21978), .Z(n21926) );
  ANDN U23302 ( .B(n21979), .A(n21980), .Z(n21977) );
  XOR U23303 ( .A(n21981), .B(n21978), .Z(n21979) );
  IV U23304 ( .A(n21936), .Z(n21940) );
  XOR U23305 ( .A(n21936), .B(n21891), .Z(n21938) );
  XOR U23306 ( .A(n21982), .B(n21983), .Z(n21891) );
  AND U23307 ( .A(n438), .B(n21984), .Z(n21982) );
  XOR U23308 ( .A(n21985), .B(n21983), .Z(n21984) );
  NANDN U23309 ( .A(n21893), .B(n21895), .Z(n21936) );
  XOR U23310 ( .A(n21986), .B(n21987), .Z(n21895) );
  AND U23311 ( .A(n438), .B(n21988), .Z(n21986) );
  XOR U23312 ( .A(n21987), .B(n21989), .Z(n21988) );
  XNOR U23313 ( .A(n21990), .B(n21991), .Z(n438) );
  AND U23314 ( .A(n21992), .B(n21993), .Z(n21990) );
  XOR U23315 ( .A(n21991), .B(n21906), .Z(n21993) );
  XNOR U23316 ( .A(n21994), .B(n21995), .Z(n21906) );
  ANDN U23317 ( .B(n21996), .A(n21997), .Z(n21994) );
  XOR U23318 ( .A(n21995), .B(n21998), .Z(n21996) );
  XNOR U23319 ( .A(n21991), .B(n21908), .Z(n21992) );
  XOR U23320 ( .A(n21999), .B(n22000), .Z(n21908) );
  AND U23321 ( .A(n442), .B(n22001), .Z(n21999) );
  XOR U23322 ( .A(n22002), .B(n22000), .Z(n22001) );
  XNOR U23323 ( .A(n22003), .B(n22004), .Z(n21991) );
  AND U23324 ( .A(n22005), .B(n22006), .Z(n22003) );
  XNOR U23325 ( .A(n22004), .B(n21933), .Z(n22006) );
  XOR U23326 ( .A(n21997), .B(n21998), .Z(n21933) );
  XNOR U23327 ( .A(n22007), .B(n22008), .Z(n21998) );
  ANDN U23328 ( .B(n22009), .A(n22010), .Z(n22007) );
  XOR U23329 ( .A(n22011), .B(n22012), .Z(n22009) );
  XOR U23330 ( .A(n22013), .B(n22014), .Z(n21997) );
  XNOR U23331 ( .A(n22015), .B(n22016), .Z(n22014) );
  ANDN U23332 ( .B(n22017), .A(n22018), .Z(n22015) );
  XNOR U23333 ( .A(n22019), .B(n22020), .Z(n22017) );
  IV U23334 ( .A(n21995), .Z(n22013) );
  XOR U23335 ( .A(n22021), .B(n22022), .Z(n21995) );
  ANDN U23336 ( .B(n22023), .A(n22024), .Z(n22021) );
  XOR U23337 ( .A(n22022), .B(n22025), .Z(n22023) );
  XOR U23338 ( .A(n22004), .B(n21935), .Z(n22005) );
  XOR U23339 ( .A(n22026), .B(n22027), .Z(n21935) );
  AND U23340 ( .A(n442), .B(n22028), .Z(n22026) );
  XOR U23341 ( .A(n22029), .B(n22027), .Z(n22028) );
  XNOR U23342 ( .A(n22030), .B(n22031), .Z(n22004) );
  NAND U23343 ( .A(n22032), .B(n22033), .Z(n22031) );
  XOR U23344 ( .A(n22034), .B(n21983), .Z(n22033) );
  XOR U23345 ( .A(n22024), .B(n22025), .Z(n21983) );
  XOR U23346 ( .A(n22035), .B(n22012), .Z(n22025) );
  XOR U23347 ( .A(n22036), .B(n22037), .Z(n22012) );
  ANDN U23348 ( .B(n22038), .A(n22039), .Z(n22036) );
  XOR U23349 ( .A(n22037), .B(n22040), .Z(n22038) );
  IV U23350 ( .A(n22010), .Z(n22035) );
  XOR U23351 ( .A(n22008), .B(n22041), .Z(n22010) );
  XOR U23352 ( .A(n22042), .B(n22043), .Z(n22041) );
  ANDN U23353 ( .B(n22044), .A(n22045), .Z(n22042) );
  XOR U23354 ( .A(n22046), .B(n22043), .Z(n22044) );
  IV U23355 ( .A(n22011), .Z(n22008) );
  XOR U23356 ( .A(n22047), .B(n22048), .Z(n22011) );
  ANDN U23357 ( .B(n22049), .A(n22050), .Z(n22047) );
  XOR U23358 ( .A(n22048), .B(n22051), .Z(n22049) );
  XOR U23359 ( .A(n22052), .B(n22053), .Z(n22024) );
  XNOR U23360 ( .A(n22019), .B(n22054), .Z(n22053) );
  IV U23361 ( .A(n22022), .Z(n22054) );
  XOR U23362 ( .A(n22055), .B(n22056), .Z(n22022) );
  ANDN U23363 ( .B(n22057), .A(n22058), .Z(n22055) );
  XOR U23364 ( .A(n22056), .B(n22059), .Z(n22057) );
  XNOR U23365 ( .A(n22060), .B(n22061), .Z(n22019) );
  ANDN U23366 ( .B(n22062), .A(n22063), .Z(n22060) );
  XOR U23367 ( .A(n22061), .B(n22064), .Z(n22062) );
  IV U23368 ( .A(n22018), .Z(n22052) );
  XOR U23369 ( .A(n22016), .B(n22065), .Z(n22018) );
  XOR U23370 ( .A(n22066), .B(n22067), .Z(n22065) );
  ANDN U23371 ( .B(n22068), .A(n22069), .Z(n22066) );
  XOR U23372 ( .A(n22070), .B(n22067), .Z(n22068) );
  IV U23373 ( .A(n22020), .Z(n22016) );
  XOR U23374 ( .A(n22071), .B(n22072), .Z(n22020) );
  ANDN U23375 ( .B(n22073), .A(n22074), .Z(n22071) );
  XOR U23376 ( .A(n22075), .B(n22072), .Z(n22073) );
  IV U23377 ( .A(n22030), .Z(n22034) );
  XOR U23378 ( .A(n22030), .B(n21985), .Z(n22032) );
  XOR U23379 ( .A(n22076), .B(n22077), .Z(n21985) );
  AND U23380 ( .A(n442), .B(n22078), .Z(n22076) );
  XOR U23381 ( .A(n22079), .B(n22077), .Z(n22078) );
  NANDN U23382 ( .A(n21987), .B(n21989), .Z(n22030) );
  XOR U23383 ( .A(n22080), .B(n22081), .Z(n21989) );
  AND U23384 ( .A(n442), .B(n22082), .Z(n22080) );
  XOR U23385 ( .A(n22081), .B(n22083), .Z(n22082) );
  XNOR U23386 ( .A(n22084), .B(n22085), .Z(n442) );
  AND U23387 ( .A(n22086), .B(n22087), .Z(n22084) );
  XOR U23388 ( .A(n22085), .B(n22000), .Z(n22087) );
  XNOR U23389 ( .A(n22088), .B(n22089), .Z(n22000) );
  ANDN U23390 ( .B(n22090), .A(n22091), .Z(n22088) );
  XOR U23391 ( .A(n22089), .B(n22092), .Z(n22090) );
  XNOR U23392 ( .A(n22085), .B(n22002), .Z(n22086) );
  XOR U23393 ( .A(n22093), .B(n22094), .Z(n22002) );
  AND U23394 ( .A(n446), .B(n22095), .Z(n22093) );
  XOR U23395 ( .A(n22096), .B(n22094), .Z(n22095) );
  XNOR U23396 ( .A(n22097), .B(n22098), .Z(n22085) );
  AND U23397 ( .A(n22099), .B(n22100), .Z(n22097) );
  XNOR U23398 ( .A(n22098), .B(n22027), .Z(n22100) );
  XOR U23399 ( .A(n22091), .B(n22092), .Z(n22027) );
  XNOR U23400 ( .A(n22101), .B(n22102), .Z(n22092) );
  ANDN U23401 ( .B(n22103), .A(n22104), .Z(n22101) );
  XOR U23402 ( .A(n22105), .B(n22106), .Z(n22103) );
  XOR U23403 ( .A(n22107), .B(n22108), .Z(n22091) );
  XNOR U23404 ( .A(n22109), .B(n22110), .Z(n22108) );
  ANDN U23405 ( .B(n22111), .A(n22112), .Z(n22109) );
  XNOR U23406 ( .A(n22113), .B(n22114), .Z(n22111) );
  IV U23407 ( .A(n22089), .Z(n22107) );
  XOR U23408 ( .A(n22115), .B(n22116), .Z(n22089) );
  ANDN U23409 ( .B(n22117), .A(n22118), .Z(n22115) );
  XOR U23410 ( .A(n22116), .B(n22119), .Z(n22117) );
  XOR U23411 ( .A(n22098), .B(n22029), .Z(n22099) );
  XOR U23412 ( .A(n22120), .B(n22121), .Z(n22029) );
  AND U23413 ( .A(n446), .B(n22122), .Z(n22120) );
  XOR U23414 ( .A(n22123), .B(n22121), .Z(n22122) );
  XNOR U23415 ( .A(n22124), .B(n22125), .Z(n22098) );
  NAND U23416 ( .A(n22126), .B(n22127), .Z(n22125) );
  XOR U23417 ( .A(n22128), .B(n22077), .Z(n22127) );
  XOR U23418 ( .A(n22118), .B(n22119), .Z(n22077) );
  XOR U23419 ( .A(n22129), .B(n22106), .Z(n22119) );
  XOR U23420 ( .A(n22130), .B(n22131), .Z(n22106) );
  ANDN U23421 ( .B(n22132), .A(n22133), .Z(n22130) );
  XOR U23422 ( .A(n22131), .B(n22134), .Z(n22132) );
  IV U23423 ( .A(n22104), .Z(n22129) );
  XOR U23424 ( .A(n22102), .B(n22135), .Z(n22104) );
  XOR U23425 ( .A(n22136), .B(n22137), .Z(n22135) );
  ANDN U23426 ( .B(n22138), .A(n22139), .Z(n22136) );
  XOR U23427 ( .A(n22140), .B(n22137), .Z(n22138) );
  IV U23428 ( .A(n22105), .Z(n22102) );
  XOR U23429 ( .A(n22141), .B(n22142), .Z(n22105) );
  ANDN U23430 ( .B(n22143), .A(n22144), .Z(n22141) );
  XOR U23431 ( .A(n22142), .B(n22145), .Z(n22143) );
  XOR U23432 ( .A(n22146), .B(n22147), .Z(n22118) );
  XNOR U23433 ( .A(n22113), .B(n22148), .Z(n22147) );
  IV U23434 ( .A(n22116), .Z(n22148) );
  XOR U23435 ( .A(n22149), .B(n22150), .Z(n22116) );
  ANDN U23436 ( .B(n22151), .A(n22152), .Z(n22149) );
  XOR U23437 ( .A(n22150), .B(n22153), .Z(n22151) );
  XNOR U23438 ( .A(n22154), .B(n22155), .Z(n22113) );
  ANDN U23439 ( .B(n22156), .A(n22157), .Z(n22154) );
  XOR U23440 ( .A(n22155), .B(n22158), .Z(n22156) );
  IV U23441 ( .A(n22112), .Z(n22146) );
  XOR U23442 ( .A(n22110), .B(n22159), .Z(n22112) );
  XOR U23443 ( .A(n22160), .B(n22161), .Z(n22159) );
  ANDN U23444 ( .B(n22162), .A(n22163), .Z(n22160) );
  XOR U23445 ( .A(n22164), .B(n22161), .Z(n22162) );
  IV U23446 ( .A(n22114), .Z(n22110) );
  XOR U23447 ( .A(n22165), .B(n22166), .Z(n22114) );
  ANDN U23448 ( .B(n22167), .A(n22168), .Z(n22165) );
  XOR U23449 ( .A(n22169), .B(n22166), .Z(n22167) );
  IV U23450 ( .A(n22124), .Z(n22128) );
  XOR U23451 ( .A(n22124), .B(n22079), .Z(n22126) );
  XOR U23452 ( .A(n22170), .B(n22171), .Z(n22079) );
  AND U23453 ( .A(n446), .B(n22172), .Z(n22170) );
  XOR U23454 ( .A(n22173), .B(n22171), .Z(n22172) );
  NANDN U23455 ( .A(n22081), .B(n22083), .Z(n22124) );
  XOR U23456 ( .A(n22174), .B(n22175), .Z(n22083) );
  AND U23457 ( .A(n446), .B(n22176), .Z(n22174) );
  XOR U23458 ( .A(n22175), .B(n22177), .Z(n22176) );
  XNOR U23459 ( .A(n22178), .B(n22179), .Z(n446) );
  AND U23460 ( .A(n22180), .B(n22181), .Z(n22178) );
  XOR U23461 ( .A(n22179), .B(n22094), .Z(n22181) );
  XNOR U23462 ( .A(n22182), .B(n22183), .Z(n22094) );
  ANDN U23463 ( .B(n22184), .A(n22185), .Z(n22182) );
  XOR U23464 ( .A(n22183), .B(n22186), .Z(n22184) );
  XNOR U23465 ( .A(n22179), .B(n22096), .Z(n22180) );
  XOR U23466 ( .A(n22187), .B(n22188), .Z(n22096) );
  AND U23467 ( .A(n450), .B(n22189), .Z(n22187) );
  XOR U23468 ( .A(n22190), .B(n22188), .Z(n22189) );
  XNOR U23469 ( .A(n22191), .B(n22192), .Z(n22179) );
  AND U23470 ( .A(n22193), .B(n22194), .Z(n22191) );
  XNOR U23471 ( .A(n22192), .B(n22121), .Z(n22194) );
  XOR U23472 ( .A(n22185), .B(n22186), .Z(n22121) );
  XNOR U23473 ( .A(n22195), .B(n22196), .Z(n22186) );
  ANDN U23474 ( .B(n22197), .A(n22198), .Z(n22195) );
  XOR U23475 ( .A(n22199), .B(n22200), .Z(n22197) );
  XOR U23476 ( .A(n22201), .B(n22202), .Z(n22185) );
  XNOR U23477 ( .A(n22203), .B(n22204), .Z(n22202) );
  ANDN U23478 ( .B(n22205), .A(n22206), .Z(n22203) );
  XNOR U23479 ( .A(n22207), .B(n22208), .Z(n22205) );
  IV U23480 ( .A(n22183), .Z(n22201) );
  XOR U23481 ( .A(n22209), .B(n22210), .Z(n22183) );
  ANDN U23482 ( .B(n22211), .A(n22212), .Z(n22209) );
  XOR U23483 ( .A(n22210), .B(n22213), .Z(n22211) );
  XOR U23484 ( .A(n22192), .B(n22123), .Z(n22193) );
  XOR U23485 ( .A(n22214), .B(n22215), .Z(n22123) );
  AND U23486 ( .A(n450), .B(n22216), .Z(n22214) );
  XOR U23487 ( .A(n22217), .B(n22215), .Z(n22216) );
  XNOR U23488 ( .A(n22218), .B(n22219), .Z(n22192) );
  NAND U23489 ( .A(n22220), .B(n22221), .Z(n22219) );
  XOR U23490 ( .A(n22222), .B(n22171), .Z(n22221) );
  XOR U23491 ( .A(n22212), .B(n22213), .Z(n22171) );
  XOR U23492 ( .A(n22223), .B(n22200), .Z(n22213) );
  XOR U23493 ( .A(n22224), .B(n22225), .Z(n22200) );
  ANDN U23494 ( .B(n22226), .A(n22227), .Z(n22224) );
  XOR U23495 ( .A(n22225), .B(n22228), .Z(n22226) );
  IV U23496 ( .A(n22198), .Z(n22223) );
  XOR U23497 ( .A(n22196), .B(n22229), .Z(n22198) );
  XOR U23498 ( .A(n22230), .B(n22231), .Z(n22229) );
  ANDN U23499 ( .B(n22232), .A(n22233), .Z(n22230) );
  XOR U23500 ( .A(n22234), .B(n22231), .Z(n22232) );
  IV U23501 ( .A(n22199), .Z(n22196) );
  XOR U23502 ( .A(n22235), .B(n22236), .Z(n22199) );
  ANDN U23503 ( .B(n22237), .A(n22238), .Z(n22235) );
  XOR U23504 ( .A(n22236), .B(n22239), .Z(n22237) );
  XOR U23505 ( .A(n22240), .B(n22241), .Z(n22212) );
  XNOR U23506 ( .A(n22207), .B(n22242), .Z(n22241) );
  IV U23507 ( .A(n22210), .Z(n22242) );
  XOR U23508 ( .A(n22243), .B(n22244), .Z(n22210) );
  ANDN U23509 ( .B(n22245), .A(n22246), .Z(n22243) );
  XOR U23510 ( .A(n22244), .B(n22247), .Z(n22245) );
  XNOR U23511 ( .A(n22248), .B(n22249), .Z(n22207) );
  ANDN U23512 ( .B(n22250), .A(n22251), .Z(n22248) );
  XOR U23513 ( .A(n22249), .B(n22252), .Z(n22250) );
  IV U23514 ( .A(n22206), .Z(n22240) );
  XOR U23515 ( .A(n22204), .B(n22253), .Z(n22206) );
  XOR U23516 ( .A(n22254), .B(n22255), .Z(n22253) );
  ANDN U23517 ( .B(n22256), .A(n22257), .Z(n22254) );
  XOR U23518 ( .A(n22258), .B(n22255), .Z(n22256) );
  IV U23519 ( .A(n22208), .Z(n22204) );
  XOR U23520 ( .A(n22259), .B(n22260), .Z(n22208) );
  ANDN U23521 ( .B(n22261), .A(n22262), .Z(n22259) );
  XOR U23522 ( .A(n22263), .B(n22260), .Z(n22261) );
  IV U23523 ( .A(n22218), .Z(n22222) );
  XOR U23524 ( .A(n22218), .B(n22173), .Z(n22220) );
  XOR U23525 ( .A(n22264), .B(n22265), .Z(n22173) );
  AND U23526 ( .A(n450), .B(n22266), .Z(n22264) );
  XOR U23527 ( .A(n22267), .B(n22265), .Z(n22266) );
  NANDN U23528 ( .A(n22175), .B(n22177), .Z(n22218) );
  XOR U23529 ( .A(n22268), .B(n22269), .Z(n22177) );
  AND U23530 ( .A(n450), .B(n22270), .Z(n22268) );
  XOR U23531 ( .A(n22269), .B(n22271), .Z(n22270) );
  XNOR U23532 ( .A(n22272), .B(n22273), .Z(n450) );
  AND U23533 ( .A(n22274), .B(n22275), .Z(n22272) );
  XOR U23534 ( .A(n22273), .B(n22188), .Z(n22275) );
  XNOR U23535 ( .A(n22276), .B(n22277), .Z(n22188) );
  ANDN U23536 ( .B(n22278), .A(n22279), .Z(n22276) );
  XOR U23537 ( .A(n22277), .B(n22280), .Z(n22278) );
  XNOR U23538 ( .A(n22273), .B(n22190), .Z(n22274) );
  XOR U23539 ( .A(n22281), .B(n22282), .Z(n22190) );
  AND U23540 ( .A(n454), .B(n22283), .Z(n22281) );
  XOR U23541 ( .A(n22284), .B(n22282), .Z(n22283) );
  XNOR U23542 ( .A(n22285), .B(n22286), .Z(n22273) );
  AND U23543 ( .A(n22287), .B(n22288), .Z(n22285) );
  XNOR U23544 ( .A(n22286), .B(n22215), .Z(n22288) );
  XOR U23545 ( .A(n22279), .B(n22280), .Z(n22215) );
  XNOR U23546 ( .A(n22289), .B(n22290), .Z(n22280) );
  ANDN U23547 ( .B(n22291), .A(n22292), .Z(n22289) );
  XOR U23548 ( .A(n22293), .B(n22294), .Z(n22291) );
  XOR U23549 ( .A(n22295), .B(n22296), .Z(n22279) );
  XNOR U23550 ( .A(n22297), .B(n22298), .Z(n22296) );
  ANDN U23551 ( .B(n22299), .A(n22300), .Z(n22297) );
  XNOR U23552 ( .A(n22301), .B(n22302), .Z(n22299) );
  IV U23553 ( .A(n22277), .Z(n22295) );
  XOR U23554 ( .A(n22303), .B(n22304), .Z(n22277) );
  ANDN U23555 ( .B(n22305), .A(n22306), .Z(n22303) );
  XOR U23556 ( .A(n22304), .B(n22307), .Z(n22305) );
  XOR U23557 ( .A(n22286), .B(n22217), .Z(n22287) );
  XOR U23558 ( .A(n22308), .B(n22309), .Z(n22217) );
  AND U23559 ( .A(n454), .B(n22310), .Z(n22308) );
  XOR U23560 ( .A(n22311), .B(n22309), .Z(n22310) );
  XNOR U23561 ( .A(n22312), .B(n22313), .Z(n22286) );
  NAND U23562 ( .A(n22314), .B(n22315), .Z(n22313) );
  XOR U23563 ( .A(n22316), .B(n22265), .Z(n22315) );
  XOR U23564 ( .A(n22306), .B(n22307), .Z(n22265) );
  XOR U23565 ( .A(n22317), .B(n22294), .Z(n22307) );
  XOR U23566 ( .A(n22318), .B(n22319), .Z(n22294) );
  ANDN U23567 ( .B(n22320), .A(n22321), .Z(n22318) );
  XOR U23568 ( .A(n22319), .B(n22322), .Z(n22320) );
  IV U23569 ( .A(n22292), .Z(n22317) );
  XOR U23570 ( .A(n22290), .B(n22323), .Z(n22292) );
  XOR U23571 ( .A(n22324), .B(n22325), .Z(n22323) );
  ANDN U23572 ( .B(n22326), .A(n22327), .Z(n22324) );
  XOR U23573 ( .A(n22328), .B(n22325), .Z(n22326) );
  IV U23574 ( .A(n22293), .Z(n22290) );
  XOR U23575 ( .A(n22329), .B(n22330), .Z(n22293) );
  ANDN U23576 ( .B(n22331), .A(n22332), .Z(n22329) );
  XOR U23577 ( .A(n22330), .B(n22333), .Z(n22331) );
  XOR U23578 ( .A(n22334), .B(n22335), .Z(n22306) );
  XNOR U23579 ( .A(n22301), .B(n22336), .Z(n22335) );
  IV U23580 ( .A(n22304), .Z(n22336) );
  XOR U23581 ( .A(n22337), .B(n22338), .Z(n22304) );
  ANDN U23582 ( .B(n22339), .A(n22340), .Z(n22337) );
  XOR U23583 ( .A(n22338), .B(n22341), .Z(n22339) );
  XNOR U23584 ( .A(n22342), .B(n22343), .Z(n22301) );
  ANDN U23585 ( .B(n22344), .A(n22345), .Z(n22342) );
  XOR U23586 ( .A(n22343), .B(n22346), .Z(n22344) );
  IV U23587 ( .A(n22300), .Z(n22334) );
  XOR U23588 ( .A(n22298), .B(n22347), .Z(n22300) );
  XOR U23589 ( .A(n22348), .B(n22349), .Z(n22347) );
  ANDN U23590 ( .B(n22350), .A(n22351), .Z(n22348) );
  XOR U23591 ( .A(n22352), .B(n22349), .Z(n22350) );
  IV U23592 ( .A(n22302), .Z(n22298) );
  XOR U23593 ( .A(n22353), .B(n22354), .Z(n22302) );
  ANDN U23594 ( .B(n22355), .A(n22356), .Z(n22353) );
  XOR U23595 ( .A(n22357), .B(n22354), .Z(n22355) );
  IV U23596 ( .A(n22312), .Z(n22316) );
  XOR U23597 ( .A(n22312), .B(n22267), .Z(n22314) );
  XOR U23598 ( .A(n22358), .B(n22359), .Z(n22267) );
  AND U23599 ( .A(n454), .B(n22360), .Z(n22358) );
  XOR U23600 ( .A(n22361), .B(n22359), .Z(n22360) );
  NANDN U23601 ( .A(n22269), .B(n22271), .Z(n22312) );
  XOR U23602 ( .A(n22362), .B(n22363), .Z(n22271) );
  AND U23603 ( .A(n454), .B(n22364), .Z(n22362) );
  XOR U23604 ( .A(n22363), .B(n22365), .Z(n22364) );
  XNOR U23605 ( .A(n22366), .B(n22367), .Z(n454) );
  AND U23606 ( .A(n22368), .B(n22369), .Z(n22366) );
  XOR U23607 ( .A(n22367), .B(n22282), .Z(n22369) );
  XNOR U23608 ( .A(n22370), .B(n22371), .Z(n22282) );
  ANDN U23609 ( .B(n22372), .A(n22373), .Z(n22370) );
  XOR U23610 ( .A(n22371), .B(n22374), .Z(n22372) );
  XNOR U23611 ( .A(n22367), .B(n22284), .Z(n22368) );
  XOR U23612 ( .A(n22375), .B(n22376), .Z(n22284) );
  AND U23613 ( .A(n458), .B(n22377), .Z(n22375) );
  XOR U23614 ( .A(n22378), .B(n22376), .Z(n22377) );
  XNOR U23615 ( .A(n22379), .B(n22380), .Z(n22367) );
  AND U23616 ( .A(n22381), .B(n22382), .Z(n22379) );
  XNOR U23617 ( .A(n22380), .B(n22309), .Z(n22382) );
  XOR U23618 ( .A(n22373), .B(n22374), .Z(n22309) );
  XNOR U23619 ( .A(n22383), .B(n22384), .Z(n22374) );
  ANDN U23620 ( .B(n22385), .A(n22386), .Z(n22383) );
  XOR U23621 ( .A(n22387), .B(n22388), .Z(n22385) );
  XOR U23622 ( .A(n22389), .B(n22390), .Z(n22373) );
  XNOR U23623 ( .A(n22391), .B(n22392), .Z(n22390) );
  ANDN U23624 ( .B(n22393), .A(n22394), .Z(n22391) );
  XNOR U23625 ( .A(n22395), .B(n22396), .Z(n22393) );
  IV U23626 ( .A(n22371), .Z(n22389) );
  XOR U23627 ( .A(n22397), .B(n22398), .Z(n22371) );
  ANDN U23628 ( .B(n22399), .A(n22400), .Z(n22397) );
  XOR U23629 ( .A(n22398), .B(n22401), .Z(n22399) );
  XOR U23630 ( .A(n22380), .B(n22311), .Z(n22381) );
  XOR U23631 ( .A(n22402), .B(n22403), .Z(n22311) );
  AND U23632 ( .A(n458), .B(n22404), .Z(n22402) );
  XOR U23633 ( .A(n22405), .B(n22403), .Z(n22404) );
  XNOR U23634 ( .A(n22406), .B(n22407), .Z(n22380) );
  NAND U23635 ( .A(n22408), .B(n22409), .Z(n22407) );
  XOR U23636 ( .A(n22410), .B(n22359), .Z(n22409) );
  XOR U23637 ( .A(n22400), .B(n22401), .Z(n22359) );
  XOR U23638 ( .A(n22411), .B(n22388), .Z(n22401) );
  XOR U23639 ( .A(n22412), .B(n22413), .Z(n22388) );
  ANDN U23640 ( .B(n22414), .A(n22415), .Z(n22412) );
  XOR U23641 ( .A(n22413), .B(n22416), .Z(n22414) );
  IV U23642 ( .A(n22386), .Z(n22411) );
  XOR U23643 ( .A(n22384), .B(n22417), .Z(n22386) );
  XOR U23644 ( .A(n22418), .B(n22419), .Z(n22417) );
  ANDN U23645 ( .B(n22420), .A(n22421), .Z(n22418) );
  XOR U23646 ( .A(n22422), .B(n22419), .Z(n22420) );
  IV U23647 ( .A(n22387), .Z(n22384) );
  XOR U23648 ( .A(n22423), .B(n22424), .Z(n22387) );
  ANDN U23649 ( .B(n22425), .A(n22426), .Z(n22423) );
  XOR U23650 ( .A(n22424), .B(n22427), .Z(n22425) );
  XOR U23651 ( .A(n22428), .B(n22429), .Z(n22400) );
  XNOR U23652 ( .A(n22395), .B(n22430), .Z(n22429) );
  IV U23653 ( .A(n22398), .Z(n22430) );
  XOR U23654 ( .A(n22431), .B(n22432), .Z(n22398) );
  ANDN U23655 ( .B(n22433), .A(n22434), .Z(n22431) );
  XOR U23656 ( .A(n22432), .B(n22435), .Z(n22433) );
  XNOR U23657 ( .A(n22436), .B(n22437), .Z(n22395) );
  ANDN U23658 ( .B(n22438), .A(n22439), .Z(n22436) );
  XOR U23659 ( .A(n22437), .B(n22440), .Z(n22438) );
  IV U23660 ( .A(n22394), .Z(n22428) );
  XOR U23661 ( .A(n22392), .B(n22441), .Z(n22394) );
  XOR U23662 ( .A(n22442), .B(n22443), .Z(n22441) );
  ANDN U23663 ( .B(n22444), .A(n22445), .Z(n22442) );
  XOR U23664 ( .A(n22446), .B(n22443), .Z(n22444) );
  IV U23665 ( .A(n22396), .Z(n22392) );
  XOR U23666 ( .A(n22447), .B(n22448), .Z(n22396) );
  ANDN U23667 ( .B(n22449), .A(n22450), .Z(n22447) );
  XOR U23668 ( .A(n22451), .B(n22448), .Z(n22449) );
  IV U23669 ( .A(n22406), .Z(n22410) );
  XOR U23670 ( .A(n22406), .B(n22361), .Z(n22408) );
  XOR U23671 ( .A(n22452), .B(n22453), .Z(n22361) );
  AND U23672 ( .A(n458), .B(n22454), .Z(n22452) );
  XOR U23673 ( .A(n22455), .B(n22453), .Z(n22454) );
  NANDN U23674 ( .A(n22363), .B(n22365), .Z(n22406) );
  XOR U23675 ( .A(n22456), .B(n22457), .Z(n22365) );
  AND U23676 ( .A(n458), .B(n22458), .Z(n22456) );
  XOR U23677 ( .A(n22457), .B(n22459), .Z(n22458) );
  XNOR U23678 ( .A(n22460), .B(n22461), .Z(n458) );
  AND U23679 ( .A(n22462), .B(n22463), .Z(n22460) );
  XOR U23680 ( .A(n22461), .B(n22376), .Z(n22463) );
  XNOR U23681 ( .A(n22464), .B(n22465), .Z(n22376) );
  ANDN U23682 ( .B(n22466), .A(n22467), .Z(n22464) );
  XOR U23683 ( .A(n22465), .B(n22468), .Z(n22466) );
  XNOR U23684 ( .A(n22461), .B(n22378), .Z(n22462) );
  XOR U23685 ( .A(n22469), .B(n22470), .Z(n22378) );
  AND U23686 ( .A(n462), .B(n22471), .Z(n22469) );
  XOR U23687 ( .A(n22472), .B(n22470), .Z(n22471) );
  XNOR U23688 ( .A(n22473), .B(n22474), .Z(n22461) );
  AND U23689 ( .A(n22475), .B(n22476), .Z(n22473) );
  XNOR U23690 ( .A(n22474), .B(n22403), .Z(n22476) );
  XOR U23691 ( .A(n22467), .B(n22468), .Z(n22403) );
  XNOR U23692 ( .A(n22477), .B(n22478), .Z(n22468) );
  ANDN U23693 ( .B(n22479), .A(n22480), .Z(n22477) );
  XOR U23694 ( .A(n22481), .B(n22482), .Z(n22479) );
  XOR U23695 ( .A(n22483), .B(n22484), .Z(n22467) );
  XNOR U23696 ( .A(n22485), .B(n22486), .Z(n22484) );
  ANDN U23697 ( .B(n22487), .A(n22488), .Z(n22485) );
  XNOR U23698 ( .A(n22489), .B(n22490), .Z(n22487) );
  IV U23699 ( .A(n22465), .Z(n22483) );
  XOR U23700 ( .A(n22491), .B(n22492), .Z(n22465) );
  ANDN U23701 ( .B(n22493), .A(n22494), .Z(n22491) );
  XOR U23702 ( .A(n22492), .B(n22495), .Z(n22493) );
  XOR U23703 ( .A(n22474), .B(n22405), .Z(n22475) );
  XOR U23704 ( .A(n22496), .B(n22497), .Z(n22405) );
  AND U23705 ( .A(n462), .B(n22498), .Z(n22496) );
  XOR U23706 ( .A(n22499), .B(n22497), .Z(n22498) );
  XNOR U23707 ( .A(n22500), .B(n22501), .Z(n22474) );
  NAND U23708 ( .A(n22502), .B(n22503), .Z(n22501) );
  XOR U23709 ( .A(n22504), .B(n22453), .Z(n22503) );
  XOR U23710 ( .A(n22494), .B(n22495), .Z(n22453) );
  XOR U23711 ( .A(n22505), .B(n22482), .Z(n22495) );
  XOR U23712 ( .A(n22506), .B(n22507), .Z(n22482) );
  ANDN U23713 ( .B(n22508), .A(n22509), .Z(n22506) );
  XOR U23714 ( .A(n22507), .B(n22510), .Z(n22508) );
  IV U23715 ( .A(n22480), .Z(n22505) );
  XOR U23716 ( .A(n22478), .B(n22511), .Z(n22480) );
  XOR U23717 ( .A(n22512), .B(n22513), .Z(n22511) );
  ANDN U23718 ( .B(n22514), .A(n22515), .Z(n22512) );
  XOR U23719 ( .A(n22516), .B(n22513), .Z(n22514) );
  IV U23720 ( .A(n22481), .Z(n22478) );
  XOR U23721 ( .A(n22517), .B(n22518), .Z(n22481) );
  ANDN U23722 ( .B(n22519), .A(n22520), .Z(n22517) );
  XOR U23723 ( .A(n22518), .B(n22521), .Z(n22519) );
  XOR U23724 ( .A(n22522), .B(n22523), .Z(n22494) );
  XNOR U23725 ( .A(n22489), .B(n22524), .Z(n22523) );
  IV U23726 ( .A(n22492), .Z(n22524) );
  XOR U23727 ( .A(n22525), .B(n22526), .Z(n22492) );
  ANDN U23728 ( .B(n22527), .A(n22528), .Z(n22525) );
  XOR U23729 ( .A(n22526), .B(n22529), .Z(n22527) );
  XNOR U23730 ( .A(n22530), .B(n22531), .Z(n22489) );
  ANDN U23731 ( .B(n22532), .A(n22533), .Z(n22530) );
  XOR U23732 ( .A(n22531), .B(n22534), .Z(n22532) );
  IV U23733 ( .A(n22488), .Z(n22522) );
  XOR U23734 ( .A(n22486), .B(n22535), .Z(n22488) );
  XOR U23735 ( .A(n22536), .B(n22537), .Z(n22535) );
  ANDN U23736 ( .B(n22538), .A(n22539), .Z(n22536) );
  XOR U23737 ( .A(n22540), .B(n22537), .Z(n22538) );
  IV U23738 ( .A(n22490), .Z(n22486) );
  XOR U23739 ( .A(n22541), .B(n22542), .Z(n22490) );
  ANDN U23740 ( .B(n22543), .A(n22544), .Z(n22541) );
  XOR U23741 ( .A(n22545), .B(n22542), .Z(n22543) );
  IV U23742 ( .A(n22500), .Z(n22504) );
  XOR U23743 ( .A(n22500), .B(n22455), .Z(n22502) );
  XOR U23744 ( .A(n22546), .B(n22547), .Z(n22455) );
  AND U23745 ( .A(n462), .B(n22548), .Z(n22546) );
  XOR U23746 ( .A(n22549), .B(n22547), .Z(n22548) );
  NANDN U23747 ( .A(n22457), .B(n22459), .Z(n22500) );
  XOR U23748 ( .A(n22550), .B(n22551), .Z(n22459) );
  AND U23749 ( .A(n462), .B(n22552), .Z(n22550) );
  XOR U23750 ( .A(n22551), .B(n22553), .Z(n22552) );
  XNOR U23751 ( .A(n22554), .B(n22555), .Z(n462) );
  AND U23752 ( .A(n22556), .B(n22557), .Z(n22554) );
  XOR U23753 ( .A(n22555), .B(n22470), .Z(n22557) );
  XNOR U23754 ( .A(n22558), .B(n22559), .Z(n22470) );
  ANDN U23755 ( .B(n22560), .A(n22561), .Z(n22558) );
  XOR U23756 ( .A(n22559), .B(n22562), .Z(n22560) );
  XNOR U23757 ( .A(n22555), .B(n22472), .Z(n22556) );
  XOR U23758 ( .A(n22563), .B(n22564), .Z(n22472) );
  AND U23759 ( .A(n466), .B(n22565), .Z(n22563) );
  XOR U23760 ( .A(n22566), .B(n22564), .Z(n22565) );
  XNOR U23761 ( .A(n22567), .B(n22568), .Z(n22555) );
  AND U23762 ( .A(n22569), .B(n22570), .Z(n22567) );
  XNOR U23763 ( .A(n22568), .B(n22497), .Z(n22570) );
  XOR U23764 ( .A(n22561), .B(n22562), .Z(n22497) );
  XNOR U23765 ( .A(n22571), .B(n22572), .Z(n22562) );
  ANDN U23766 ( .B(n22573), .A(n22574), .Z(n22571) );
  XOR U23767 ( .A(n22575), .B(n22576), .Z(n22573) );
  XOR U23768 ( .A(n22577), .B(n22578), .Z(n22561) );
  XNOR U23769 ( .A(n22579), .B(n22580), .Z(n22578) );
  ANDN U23770 ( .B(n22581), .A(n22582), .Z(n22579) );
  XNOR U23771 ( .A(n22583), .B(n22584), .Z(n22581) );
  IV U23772 ( .A(n22559), .Z(n22577) );
  XOR U23773 ( .A(n22585), .B(n22586), .Z(n22559) );
  ANDN U23774 ( .B(n22587), .A(n22588), .Z(n22585) );
  XOR U23775 ( .A(n22586), .B(n22589), .Z(n22587) );
  XOR U23776 ( .A(n22568), .B(n22499), .Z(n22569) );
  XOR U23777 ( .A(n22590), .B(n22591), .Z(n22499) );
  AND U23778 ( .A(n466), .B(n22592), .Z(n22590) );
  XOR U23779 ( .A(n22593), .B(n22591), .Z(n22592) );
  XNOR U23780 ( .A(n22594), .B(n22595), .Z(n22568) );
  NAND U23781 ( .A(n22596), .B(n22597), .Z(n22595) );
  XOR U23782 ( .A(n22598), .B(n22547), .Z(n22597) );
  XOR U23783 ( .A(n22588), .B(n22589), .Z(n22547) );
  XOR U23784 ( .A(n22599), .B(n22576), .Z(n22589) );
  XOR U23785 ( .A(n22600), .B(n22601), .Z(n22576) );
  ANDN U23786 ( .B(n22602), .A(n22603), .Z(n22600) );
  XOR U23787 ( .A(n22601), .B(n22604), .Z(n22602) );
  IV U23788 ( .A(n22574), .Z(n22599) );
  XOR U23789 ( .A(n22572), .B(n22605), .Z(n22574) );
  XOR U23790 ( .A(n22606), .B(n22607), .Z(n22605) );
  ANDN U23791 ( .B(n22608), .A(n22609), .Z(n22606) );
  XOR U23792 ( .A(n22610), .B(n22607), .Z(n22608) );
  IV U23793 ( .A(n22575), .Z(n22572) );
  XOR U23794 ( .A(n22611), .B(n22612), .Z(n22575) );
  ANDN U23795 ( .B(n22613), .A(n22614), .Z(n22611) );
  XOR U23796 ( .A(n22612), .B(n22615), .Z(n22613) );
  XOR U23797 ( .A(n22616), .B(n22617), .Z(n22588) );
  XNOR U23798 ( .A(n22583), .B(n22618), .Z(n22617) );
  IV U23799 ( .A(n22586), .Z(n22618) );
  XOR U23800 ( .A(n22619), .B(n22620), .Z(n22586) );
  ANDN U23801 ( .B(n22621), .A(n22622), .Z(n22619) );
  XOR U23802 ( .A(n22620), .B(n22623), .Z(n22621) );
  XNOR U23803 ( .A(n22624), .B(n22625), .Z(n22583) );
  ANDN U23804 ( .B(n22626), .A(n22627), .Z(n22624) );
  XOR U23805 ( .A(n22625), .B(n22628), .Z(n22626) );
  IV U23806 ( .A(n22582), .Z(n22616) );
  XOR U23807 ( .A(n22580), .B(n22629), .Z(n22582) );
  XOR U23808 ( .A(n22630), .B(n22631), .Z(n22629) );
  ANDN U23809 ( .B(n22632), .A(n22633), .Z(n22630) );
  XOR U23810 ( .A(n22634), .B(n22631), .Z(n22632) );
  IV U23811 ( .A(n22584), .Z(n22580) );
  XOR U23812 ( .A(n22635), .B(n22636), .Z(n22584) );
  ANDN U23813 ( .B(n22637), .A(n22638), .Z(n22635) );
  XOR U23814 ( .A(n22639), .B(n22636), .Z(n22637) );
  IV U23815 ( .A(n22594), .Z(n22598) );
  XOR U23816 ( .A(n22594), .B(n22549), .Z(n22596) );
  XOR U23817 ( .A(n22640), .B(n22641), .Z(n22549) );
  AND U23818 ( .A(n466), .B(n22642), .Z(n22640) );
  XOR U23819 ( .A(n22643), .B(n22641), .Z(n22642) );
  NANDN U23820 ( .A(n22551), .B(n22553), .Z(n22594) );
  XOR U23821 ( .A(n22644), .B(n22645), .Z(n22553) );
  AND U23822 ( .A(n466), .B(n22646), .Z(n22644) );
  XOR U23823 ( .A(n22645), .B(n22647), .Z(n22646) );
  XNOR U23824 ( .A(n22648), .B(n22649), .Z(n466) );
  AND U23825 ( .A(n22650), .B(n22651), .Z(n22648) );
  XOR U23826 ( .A(n22649), .B(n22564), .Z(n22651) );
  XNOR U23827 ( .A(n22652), .B(n22653), .Z(n22564) );
  ANDN U23828 ( .B(n22654), .A(n22655), .Z(n22652) );
  XOR U23829 ( .A(n22653), .B(n22656), .Z(n22654) );
  XNOR U23830 ( .A(n22649), .B(n22566), .Z(n22650) );
  XOR U23831 ( .A(n22657), .B(n22658), .Z(n22566) );
  AND U23832 ( .A(n470), .B(n22659), .Z(n22657) );
  XOR U23833 ( .A(n22660), .B(n22658), .Z(n22659) );
  XNOR U23834 ( .A(n22661), .B(n22662), .Z(n22649) );
  AND U23835 ( .A(n22663), .B(n22664), .Z(n22661) );
  XNOR U23836 ( .A(n22662), .B(n22591), .Z(n22664) );
  XOR U23837 ( .A(n22655), .B(n22656), .Z(n22591) );
  XNOR U23838 ( .A(n22665), .B(n22666), .Z(n22656) );
  ANDN U23839 ( .B(n22667), .A(n22668), .Z(n22665) );
  XOR U23840 ( .A(n22669), .B(n22670), .Z(n22667) );
  XOR U23841 ( .A(n22671), .B(n22672), .Z(n22655) );
  XNOR U23842 ( .A(n22673), .B(n22674), .Z(n22672) );
  ANDN U23843 ( .B(n22675), .A(n22676), .Z(n22673) );
  XNOR U23844 ( .A(n22677), .B(n22678), .Z(n22675) );
  IV U23845 ( .A(n22653), .Z(n22671) );
  XOR U23846 ( .A(n22679), .B(n22680), .Z(n22653) );
  ANDN U23847 ( .B(n22681), .A(n22682), .Z(n22679) );
  XOR U23848 ( .A(n22680), .B(n22683), .Z(n22681) );
  XOR U23849 ( .A(n22662), .B(n22593), .Z(n22663) );
  XOR U23850 ( .A(n22684), .B(n22685), .Z(n22593) );
  AND U23851 ( .A(n470), .B(n22686), .Z(n22684) );
  XOR U23852 ( .A(n22687), .B(n22685), .Z(n22686) );
  XNOR U23853 ( .A(n22688), .B(n22689), .Z(n22662) );
  NAND U23854 ( .A(n22690), .B(n22691), .Z(n22689) );
  XOR U23855 ( .A(n22692), .B(n22641), .Z(n22691) );
  XOR U23856 ( .A(n22682), .B(n22683), .Z(n22641) );
  XOR U23857 ( .A(n22693), .B(n22670), .Z(n22683) );
  XOR U23858 ( .A(n22694), .B(n22695), .Z(n22670) );
  ANDN U23859 ( .B(n22696), .A(n22697), .Z(n22694) );
  XOR U23860 ( .A(n22695), .B(n22698), .Z(n22696) );
  IV U23861 ( .A(n22668), .Z(n22693) );
  XOR U23862 ( .A(n22666), .B(n22699), .Z(n22668) );
  XOR U23863 ( .A(n22700), .B(n22701), .Z(n22699) );
  ANDN U23864 ( .B(n22702), .A(n22703), .Z(n22700) );
  XOR U23865 ( .A(n22704), .B(n22701), .Z(n22702) );
  IV U23866 ( .A(n22669), .Z(n22666) );
  XOR U23867 ( .A(n22705), .B(n22706), .Z(n22669) );
  ANDN U23868 ( .B(n22707), .A(n22708), .Z(n22705) );
  XOR U23869 ( .A(n22706), .B(n22709), .Z(n22707) );
  XOR U23870 ( .A(n22710), .B(n22711), .Z(n22682) );
  XNOR U23871 ( .A(n22677), .B(n22712), .Z(n22711) );
  IV U23872 ( .A(n22680), .Z(n22712) );
  XOR U23873 ( .A(n22713), .B(n22714), .Z(n22680) );
  ANDN U23874 ( .B(n22715), .A(n22716), .Z(n22713) );
  XOR U23875 ( .A(n22714), .B(n22717), .Z(n22715) );
  XNOR U23876 ( .A(n22718), .B(n22719), .Z(n22677) );
  ANDN U23877 ( .B(n22720), .A(n22721), .Z(n22718) );
  XOR U23878 ( .A(n22719), .B(n22722), .Z(n22720) );
  IV U23879 ( .A(n22676), .Z(n22710) );
  XOR U23880 ( .A(n22674), .B(n22723), .Z(n22676) );
  XOR U23881 ( .A(n22724), .B(n22725), .Z(n22723) );
  ANDN U23882 ( .B(n22726), .A(n22727), .Z(n22724) );
  XOR U23883 ( .A(n22728), .B(n22725), .Z(n22726) );
  IV U23884 ( .A(n22678), .Z(n22674) );
  XOR U23885 ( .A(n22729), .B(n22730), .Z(n22678) );
  ANDN U23886 ( .B(n22731), .A(n22732), .Z(n22729) );
  XOR U23887 ( .A(n22733), .B(n22730), .Z(n22731) );
  IV U23888 ( .A(n22688), .Z(n22692) );
  XOR U23889 ( .A(n22688), .B(n22643), .Z(n22690) );
  XOR U23890 ( .A(n22734), .B(n22735), .Z(n22643) );
  AND U23891 ( .A(n470), .B(n22736), .Z(n22734) );
  XOR U23892 ( .A(n22737), .B(n22735), .Z(n22736) );
  NANDN U23893 ( .A(n22645), .B(n22647), .Z(n22688) );
  XOR U23894 ( .A(n22738), .B(n22739), .Z(n22647) );
  AND U23895 ( .A(n470), .B(n22740), .Z(n22738) );
  XOR U23896 ( .A(n22739), .B(n22741), .Z(n22740) );
  XNOR U23897 ( .A(n22742), .B(n22743), .Z(n470) );
  AND U23898 ( .A(n22744), .B(n22745), .Z(n22742) );
  XOR U23899 ( .A(n22743), .B(n22658), .Z(n22745) );
  XNOR U23900 ( .A(n22746), .B(n22747), .Z(n22658) );
  ANDN U23901 ( .B(n22748), .A(n22749), .Z(n22746) );
  XOR U23902 ( .A(n22747), .B(n22750), .Z(n22748) );
  XNOR U23903 ( .A(n22743), .B(n22660), .Z(n22744) );
  XOR U23904 ( .A(n22751), .B(n22752), .Z(n22660) );
  AND U23905 ( .A(n474), .B(n22753), .Z(n22751) );
  XOR U23906 ( .A(n22754), .B(n22752), .Z(n22753) );
  XNOR U23907 ( .A(n22755), .B(n22756), .Z(n22743) );
  AND U23908 ( .A(n22757), .B(n22758), .Z(n22755) );
  XNOR U23909 ( .A(n22756), .B(n22685), .Z(n22758) );
  XOR U23910 ( .A(n22749), .B(n22750), .Z(n22685) );
  XNOR U23911 ( .A(n22759), .B(n22760), .Z(n22750) );
  ANDN U23912 ( .B(n22761), .A(n22762), .Z(n22759) );
  XOR U23913 ( .A(n22763), .B(n22764), .Z(n22761) );
  XOR U23914 ( .A(n22765), .B(n22766), .Z(n22749) );
  XNOR U23915 ( .A(n22767), .B(n22768), .Z(n22766) );
  ANDN U23916 ( .B(n22769), .A(n22770), .Z(n22767) );
  XNOR U23917 ( .A(n22771), .B(n22772), .Z(n22769) );
  IV U23918 ( .A(n22747), .Z(n22765) );
  XOR U23919 ( .A(n22773), .B(n22774), .Z(n22747) );
  ANDN U23920 ( .B(n22775), .A(n22776), .Z(n22773) );
  XOR U23921 ( .A(n22774), .B(n22777), .Z(n22775) );
  XOR U23922 ( .A(n22756), .B(n22687), .Z(n22757) );
  XOR U23923 ( .A(n22778), .B(n22779), .Z(n22687) );
  AND U23924 ( .A(n474), .B(n22780), .Z(n22778) );
  XOR U23925 ( .A(n22781), .B(n22779), .Z(n22780) );
  XNOR U23926 ( .A(n22782), .B(n22783), .Z(n22756) );
  NAND U23927 ( .A(n22784), .B(n22785), .Z(n22783) );
  XOR U23928 ( .A(n22786), .B(n22735), .Z(n22785) );
  XOR U23929 ( .A(n22776), .B(n22777), .Z(n22735) );
  XOR U23930 ( .A(n22787), .B(n22764), .Z(n22777) );
  XOR U23931 ( .A(n22788), .B(n22789), .Z(n22764) );
  ANDN U23932 ( .B(n22790), .A(n22791), .Z(n22788) );
  XOR U23933 ( .A(n22789), .B(n22792), .Z(n22790) );
  IV U23934 ( .A(n22762), .Z(n22787) );
  XOR U23935 ( .A(n22760), .B(n22793), .Z(n22762) );
  XOR U23936 ( .A(n22794), .B(n22795), .Z(n22793) );
  ANDN U23937 ( .B(n22796), .A(n22797), .Z(n22794) );
  XOR U23938 ( .A(n22798), .B(n22795), .Z(n22796) );
  IV U23939 ( .A(n22763), .Z(n22760) );
  XOR U23940 ( .A(n22799), .B(n22800), .Z(n22763) );
  ANDN U23941 ( .B(n22801), .A(n22802), .Z(n22799) );
  XOR U23942 ( .A(n22800), .B(n22803), .Z(n22801) );
  XOR U23943 ( .A(n22804), .B(n22805), .Z(n22776) );
  XNOR U23944 ( .A(n22771), .B(n22806), .Z(n22805) );
  IV U23945 ( .A(n22774), .Z(n22806) );
  XOR U23946 ( .A(n22807), .B(n22808), .Z(n22774) );
  ANDN U23947 ( .B(n22809), .A(n22810), .Z(n22807) );
  XOR U23948 ( .A(n22808), .B(n22811), .Z(n22809) );
  XNOR U23949 ( .A(n22812), .B(n22813), .Z(n22771) );
  ANDN U23950 ( .B(n22814), .A(n22815), .Z(n22812) );
  XOR U23951 ( .A(n22813), .B(n22816), .Z(n22814) );
  IV U23952 ( .A(n22770), .Z(n22804) );
  XOR U23953 ( .A(n22768), .B(n22817), .Z(n22770) );
  XOR U23954 ( .A(n22818), .B(n22819), .Z(n22817) );
  ANDN U23955 ( .B(n22820), .A(n22821), .Z(n22818) );
  XOR U23956 ( .A(n22822), .B(n22819), .Z(n22820) );
  IV U23957 ( .A(n22772), .Z(n22768) );
  XOR U23958 ( .A(n22823), .B(n22824), .Z(n22772) );
  ANDN U23959 ( .B(n22825), .A(n22826), .Z(n22823) );
  XOR U23960 ( .A(n22827), .B(n22824), .Z(n22825) );
  IV U23961 ( .A(n22782), .Z(n22786) );
  XOR U23962 ( .A(n22782), .B(n22737), .Z(n22784) );
  XOR U23963 ( .A(n22828), .B(n22829), .Z(n22737) );
  AND U23964 ( .A(n474), .B(n22830), .Z(n22828) );
  XOR U23965 ( .A(n22831), .B(n22829), .Z(n22830) );
  NANDN U23966 ( .A(n22739), .B(n22741), .Z(n22782) );
  XOR U23967 ( .A(n22832), .B(n22833), .Z(n22741) );
  AND U23968 ( .A(n474), .B(n22834), .Z(n22832) );
  XOR U23969 ( .A(n22833), .B(n22835), .Z(n22834) );
  XNOR U23970 ( .A(n22836), .B(n22837), .Z(n474) );
  AND U23971 ( .A(n22838), .B(n22839), .Z(n22836) );
  XOR U23972 ( .A(n22837), .B(n22752), .Z(n22839) );
  XNOR U23973 ( .A(n22840), .B(n22841), .Z(n22752) );
  ANDN U23974 ( .B(n22842), .A(n22843), .Z(n22840) );
  XOR U23975 ( .A(n22841), .B(n22844), .Z(n22842) );
  XNOR U23976 ( .A(n22837), .B(n22754), .Z(n22838) );
  XOR U23977 ( .A(n22845), .B(n22846), .Z(n22754) );
  AND U23978 ( .A(n478), .B(n22847), .Z(n22845) );
  XOR U23979 ( .A(n22848), .B(n22846), .Z(n22847) );
  XNOR U23980 ( .A(n22849), .B(n22850), .Z(n22837) );
  AND U23981 ( .A(n22851), .B(n22852), .Z(n22849) );
  XNOR U23982 ( .A(n22850), .B(n22779), .Z(n22852) );
  XOR U23983 ( .A(n22843), .B(n22844), .Z(n22779) );
  XNOR U23984 ( .A(n22853), .B(n22854), .Z(n22844) );
  ANDN U23985 ( .B(n22855), .A(n22856), .Z(n22853) );
  XOR U23986 ( .A(n22857), .B(n22858), .Z(n22855) );
  XOR U23987 ( .A(n22859), .B(n22860), .Z(n22843) );
  XNOR U23988 ( .A(n22861), .B(n22862), .Z(n22860) );
  ANDN U23989 ( .B(n22863), .A(n22864), .Z(n22861) );
  XNOR U23990 ( .A(n22865), .B(n22866), .Z(n22863) );
  IV U23991 ( .A(n22841), .Z(n22859) );
  XOR U23992 ( .A(n22867), .B(n22868), .Z(n22841) );
  ANDN U23993 ( .B(n22869), .A(n22870), .Z(n22867) );
  XOR U23994 ( .A(n22868), .B(n22871), .Z(n22869) );
  XOR U23995 ( .A(n22850), .B(n22781), .Z(n22851) );
  XOR U23996 ( .A(n22872), .B(n22873), .Z(n22781) );
  AND U23997 ( .A(n478), .B(n22874), .Z(n22872) );
  XOR U23998 ( .A(n22875), .B(n22873), .Z(n22874) );
  XNOR U23999 ( .A(n22876), .B(n22877), .Z(n22850) );
  NAND U24000 ( .A(n22878), .B(n22879), .Z(n22877) );
  XOR U24001 ( .A(n22880), .B(n22829), .Z(n22879) );
  XOR U24002 ( .A(n22870), .B(n22871), .Z(n22829) );
  XOR U24003 ( .A(n22881), .B(n22858), .Z(n22871) );
  XOR U24004 ( .A(n22882), .B(n22883), .Z(n22858) );
  ANDN U24005 ( .B(n22884), .A(n22885), .Z(n22882) );
  XOR U24006 ( .A(n22883), .B(n22886), .Z(n22884) );
  IV U24007 ( .A(n22856), .Z(n22881) );
  XOR U24008 ( .A(n22854), .B(n22887), .Z(n22856) );
  XOR U24009 ( .A(n22888), .B(n22889), .Z(n22887) );
  ANDN U24010 ( .B(n22890), .A(n22891), .Z(n22888) );
  XOR U24011 ( .A(n22892), .B(n22889), .Z(n22890) );
  IV U24012 ( .A(n22857), .Z(n22854) );
  XOR U24013 ( .A(n22893), .B(n22894), .Z(n22857) );
  ANDN U24014 ( .B(n22895), .A(n22896), .Z(n22893) );
  XOR U24015 ( .A(n22894), .B(n22897), .Z(n22895) );
  XOR U24016 ( .A(n22898), .B(n22899), .Z(n22870) );
  XNOR U24017 ( .A(n22865), .B(n22900), .Z(n22899) );
  IV U24018 ( .A(n22868), .Z(n22900) );
  XOR U24019 ( .A(n22901), .B(n22902), .Z(n22868) );
  ANDN U24020 ( .B(n22903), .A(n22904), .Z(n22901) );
  XOR U24021 ( .A(n22902), .B(n22905), .Z(n22903) );
  XNOR U24022 ( .A(n22906), .B(n22907), .Z(n22865) );
  ANDN U24023 ( .B(n22908), .A(n22909), .Z(n22906) );
  XOR U24024 ( .A(n22907), .B(n22910), .Z(n22908) );
  IV U24025 ( .A(n22864), .Z(n22898) );
  XOR U24026 ( .A(n22862), .B(n22911), .Z(n22864) );
  XOR U24027 ( .A(n22912), .B(n22913), .Z(n22911) );
  ANDN U24028 ( .B(n22914), .A(n22915), .Z(n22912) );
  XOR U24029 ( .A(n22916), .B(n22913), .Z(n22914) );
  IV U24030 ( .A(n22866), .Z(n22862) );
  XOR U24031 ( .A(n22917), .B(n22918), .Z(n22866) );
  ANDN U24032 ( .B(n22919), .A(n22920), .Z(n22917) );
  XOR U24033 ( .A(n22921), .B(n22918), .Z(n22919) );
  IV U24034 ( .A(n22876), .Z(n22880) );
  XOR U24035 ( .A(n22876), .B(n22831), .Z(n22878) );
  XOR U24036 ( .A(n22922), .B(n22923), .Z(n22831) );
  AND U24037 ( .A(n478), .B(n22924), .Z(n22922) );
  XOR U24038 ( .A(n22925), .B(n22923), .Z(n22924) );
  NANDN U24039 ( .A(n22833), .B(n22835), .Z(n22876) );
  XOR U24040 ( .A(n22926), .B(n22927), .Z(n22835) );
  AND U24041 ( .A(n478), .B(n22928), .Z(n22926) );
  XOR U24042 ( .A(n22927), .B(n22929), .Z(n22928) );
  XNOR U24043 ( .A(n22930), .B(n22931), .Z(n478) );
  AND U24044 ( .A(n22932), .B(n22933), .Z(n22930) );
  XOR U24045 ( .A(n22931), .B(n22846), .Z(n22933) );
  XNOR U24046 ( .A(n22934), .B(n22935), .Z(n22846) );
  ANDN U24047 ( .B(n22936), .A(n22937), .Z(n22934) );
  XOR U24048 ( .A(n22935), .B(n22938), .Z(n22936) );
  XNOR U24049 ( .A(n22931), .B(n22848), .Z(n22932) );
  XOR U24050 ( .A(n22939), .B(n22940), .Z(n22848) );
  AND U24051 ( .A(n482), .B(n22941), .Z(n22939) );
  XOR U24052 ( .A(n22942), .B(n22940), .Z(n22941) );
  XNOR U24053 ( .A(n22943), .B(n22944), .Z(n22931) );
  AND U24054 ( .A(n22945), .B(n22946), .Z(n22943) );
  XNOR U24055 ( .A(n22944), .B(n22873), .Z(n22946) );
  XOR U24056 ( .A(n22937), .B(n22938), .Z(n22873) );
  XNOR U24057 ( .A(n22947), .B(n22948), .Z(n22938) );
  ANDN U24058 ( .B(n22949), .A(n22950), .Z(n22947) );
  XOR U24059 ( .A(n22951), .B(n22952), .Z(n22949) );
  XOR U24060 ( .A(n22953), .B(n22954), .Z(n22937) );
  XNOR U24061 ( .A(n22955), .B(n22956), .Z(n22954) );
  ANDN U24062 ( .B(n22957), .A(n22958), .Z(n22955) );
  XNOR U24063 ( .A(n22959), .B(n22960), .Z(n22957) );
  IV U24064 ( .A(n22935), .Z(n22953) );
  XOR U24065 ( .A(n22961), .B(n22962), .Z(n22935) );
  ANDN U24066 ( .B(n22963), .A(n22964), .Z(n22961) );
  XOR U24067 ( .A(n22962), .B(n22965), .Z(n22963) );
  XOR U24068 ( .A(n22944), .B(n22875), .Z(n22945) );
  XOR U24069 ( .A(n22966), .B(n22967), .Z(n22875) );
  AND U24070 ( .A(n482), .B(n22968), .Z(n22966) );
  XOR U24071 ( .A(n22969), .B(n22967), .Z(n22968) );
  XNOR U24072 ( .A(n22970), .B(n22971), .Z(n22944) );
  NAND U24073 ( .A(n22972), .B(n22973), .Z(n22971) );
  XOR U24074 ( .A(n22974), .B(n22923), .Z(n22973) );
  XOR U24075 ( .A(n22964), .B(n22965), .Z(n22923) );
  XOR U24076 ( .A(n22975), .B(n22952), .Z(n22965) );
  XOR U24077 ( .A(n22976), .B(n22977), .Z(n22952) );
  ANDN U24078 ( .B(n22978), .A(n22979), .Z(n22976) );
  XOR U24079 ( .A(n22977), .B(n22980), .Z(n22978) );
  IV U24080 ( .A(n22950), .Z(n22975) );
  XOR U24081 ( .A(n22948), .B(n22981), .Z(n22950) );
  XOR U24082 ( .A(n22982), .B(n22983), .Z(n22981) );
  ANDN U24083 ( .B(n22984), .A(n22985), .Z(n22982) );
  XOR U24084 ( .A(n22986), .B(n22983), .Z(n22984) );
  IV U24085 ( .A(n22951), .Z(n22948) );
  XOR U24086 ( .A(n22987), .B(n22988), .Z(n22951) );
  ANDN U24087 ( .B(n22989), .A(n22990), .Z(n22987) );
  XOR U24088 ( .A(n22988), .B(n22991), .Z(n22989) );
  XOR U24089 ( .A(n22992), .B(n22993), .Z(n22964) );
  XNOR U24090 ( .A(n22959), .B(n22994), .Z(n22993) );
  IV U24091 ( .A(n22962), .Z(n22994) );
  XOR U24092 ( .A(n22995), .B(n22996), .Z(n22962) );
  ANDN U24093 ( .B(n22997), .A(n22998), .Z(n22995) );
  XOR U24094 ( .A(n22996), .B(n22999), .Z(n22997) );
  XNOR U24095 ( .A(n23000), .B(n23001), .Z(n22959) );
  ANDN U24096 ( .B(n23002), .A(n23003), .Z(n23000) );
  XOR U24097 ( .A(n23001), .B(n23004), .Z(n23002) );
  IV U24098 ( .A(n22958), .Z(n22992) );
  XOR U24099 ( .A(n22956), .B(n23005), .Z(n22958) );
  XOR U24100 ( .A(n23006), .B(n23007), .Z(n23005) );
  ANDN U24101 ( .B(n23008), .A(n23009), .Z(n23006) );
  XOR U24102 ( .A(n23010), .B(n23007), .Z(n23008) );
  IV U24103 ( .A(n22960), .Z(n22956) );
  XOR U24104 ( .A(n23011), .B(n23012), .Z(n22960) );
  ANDN U24105 ( .B(n23013), .A(n23014), .Z(n23011) );
  XOR U24106 ( .A(n23015), .B(n23012), .Z(n23013) );
  IV U24107 ( .A(n22970), .Z(n22974) );
  XOR U24108 ( .A(n22970), .B(n22925), .Z(n22972) );
  XOR U24109 ( .A(n23016), .B(n23017), .Z(n22925) );
  AND U24110 ( .A(n482), .B(n23018), .Z(n23016) );
  XOR U24111 ( .A(n23019), .B(n23017), .Z(n23018) );
  NANDN U24112 ( .A(n22927), .B(n22929), .Z(n22970) );
  XOR U24113 ( .A(n23020), .B(n23021), .Z(n22929) );
  AND U24114 ( .A(n482), .B(n23022), .Z(n23020) );
  XOR U24115 ( .A(n23021), .B(n23023), .Z(n23022) );
  XNOR U24116 ( .A(n23024), .B(n23025), .Z(n482) );
  AND U24117 ( .A(n23026), .B(n23027), .Z(n23024) );
  XOR U24118 ( .A(n23025), .B(n22940), .Z(n23027) );
  XNOR U24119 ( .A(n23028), .B(n23029), .Z(n22940) );
  ANDN U24120 ( .B(n23030), .A(n23031), .Z(n23028) );
  XOR U24121 ( .A(n23029), .B(n23032), .Z(n23030) );
  XNOR U24122 ( .A(n23025), .B(n22942), .Z(n23026) );
  XOR U24123 ( .A(n23033), .B(n23034), .Z(n22942) );
  AND U24124 ( .A(n486), .B(n23035), .Z(n23033) );
  XOR U24125 ( .A(n23036), .B(n23034), .Z(n23035) );
  XNOR U24126 ( .A(n23037), .B(n23038), .Z(n23025) );
  AND U24127 ( .A(n23039), .B(n23040), .Z(n23037) );
  XNOR U24128 ( .A(n23038), .B(n22967), .Z(n23040) );
  XOR U24129 ( .A(n23031), .B(n23032), .Z(n22967) );
  XNOR U24130 ( .A(n23041), .B(n23042), .Z(n23032) );
  ANDN U24131 ( .B(n23043), .A(n23044), .Z(n23041) );
  XOR U24132 ( .A(n23045), .B(n23046), .Z(n23043) );
  XOR U24133 ( .A(n23047), .B(n23048), .Z(n23031) );
  XNOR U24134 ( .A(n23049), .B(n23050), .Z(n23048) );
  ANDN U24135 ( .B(n23051), .A(n23052), .Z(n23049) );
  XNOR U24136 ( .A(n23053), .B(n23054), .Z(n23051) );
  IV U24137 ( .A(n23029), .Z(n23047) );
  XOR U24138 ( .A(n23055), .B(n23056), .Z(n23029) );
  ANDN U24139 ( .B(n23057), .A(n23058), .Z(n23055) );
  XOR U24140 ( .A(n23056), .B(n23059), .Z(n23057) );
  XOR U24141 ( .A(n23038), .B(n22969), .Z(n23039) );
  XOR U24142 ( .A(n23060), .B(n23061), .Z(n22969) );
  AND U24143 ( .A(n486), .B(n23062), .Z(n23060) );
  XOR U24144 ( .A(n23063), .B(n23061), .Z(n23062) );
  XNOR U24145 ( .A(n23064), .B(n23065), .Z(n23038) );
  NAND U24146 ( .A(n23066), .B(n23067), .Z(n23065) );
  XOR U24147 ( .A(n23068), .B(n23017), .Z(n23067) );
  XOR U24148 ( .A(n23058), .B(n23059), .Z(n23017) );
  XOR U24149 ( .A(n23069), .B(n23046), .Z(n23059) );
  XOR U24150 ( .A(n23070), .B(n23071), .Z(n23046) );
  ANDN U24151 ( .B(n23072), .A(n23073), .Z(n23070) );
  XOR U24152 ( .A(n23071), .B(n23074), .Z(n23072) );
  IV U24153 ( .A(n23044), .Z(n23069) );
  XOR U24154 ( .A(n23042), .B(n23075), .Z(n23044) );
  XOR U24155 ( .A(n23076), .B(n23077), .Z(n23075) );
  ANDN U24156 ( .B(n23078), .A(n23079), .Z(n23076) );
  XOR U24157 ( .A(n23080), .B(n23077), .Z(n23078) );
  IV U24158 ( .A(n23045), .Z(n23042) );
  XOR U24159 ( .A(n23081), .B(n23082), .Z(n23045) );
  ANDN U24160 ( .B(n23083), .A(n23084), .Z(n23081) );
  XOR U24161 ( .A(n23082), .B(n23085), .Z(n23083) );
  XOR U24162 ( .A(n23086), .B(n23087), .Z(n23058) );
  XNOR U24163 ( .A(n23053), .B(n23088), .Z(n23087) );
  IV U24164 ( .A(n23056), .Z(n23088) );
  XOR U24165 ( .A(n23089), .B(n23090), .Z(n23056) );
  ANDN U24166 ( .B(n23091), .A(n23092), .Z(n23089) );
  XOR U24167 ( .A(n23090), .B(n23093), .Z(n23091) );
  XNOR U24168 ( .A(n23094), .B(n23095), .Z(n23053) );
  ANDN U24169 ( .B(n23096), .A(n23097), .Z(n23094) );
  XOR U24170 ( .A(n23095), .B(n23098), .Z(n23096) );
  IV U24171 ( .A(n23052), .Z(n23086) );
  XOR U24172 ( .A(n23050), .B(n23099), .Z(n23052) );
  XOR U24173 ( .A(n23100), .B(n23101), .Z(n23099) );
  ANDN U24174 ( .B(n23102), .A(n23103), .Z(n23100) );
  XOR U24175 ( .A(n23104), .B(n23101), .Z(n23102) );
  IV U24176 ( .A(n23054), .Z(n23050) );
  XOR U24177 ( .A(n23105), .B(n23106), .Z(n23054) );
  ANDN U24178 ( .B(n23107), .A(n23108), .Z(n23105) );
  XOR U24179 ( .A(n23109), .B(n23106), .Z(n23107) );
  IV U24180 ( .A(n23064), .Z(n23068) );
  XOR U24181 ( .A(n23064), .B(n23019), .Z(n23066) );
  XOR U24182 ( .A(n23110), .B(n23111), .Z(n23019) );
  AND U24183 ( .A(n486), .B(n23112), .Z(n23110) );
  XOR U24184 ( .A(n23113), .B(n23111), .Z(n23112) );
  NANDN U24185 ( .A(n23021), .B(n23023), .Z(n23064) );
  XOR U24186 ( .A(n23114), .B(n23115), .Z(n23023) );
  AND U24187 ( .A(n486), .B(n23116), .Z(n23114) );
  XOR U24188 ( .A(n23115), .B(n23117), .Z(n23116) );
  XNOR U24189 ( .A(n23118), .B(n23119), .Z(n486) );
  AND U24190 ( .A(n23120), .B(n23121), .Z(n23118) );
  XOR U24191 ( .A(n23119), .B(n23034), .Z(n23121) );
  XNOR U24192 ( .A(n23122), .B(n23123), .Z(n23034) );
  ANDN U24193 ( .B(n23124), .A(n23125), .Z(n23122) );
  XOR U24194 ( .A(n23123), .B(n23126), .Z(n23124) );
  XNOR U24195 ( .A(n23119), .B(n23036), .Z(n23120) );
  XOR U24196 ( .A(n23127), .B(n23128), .Z(n23036) );
  AND U24197 ( .A(n490), .B(n23129), .Z(n23127) );
  XOR U24198 ( .A(n23130), .B(n23128), .Z(n23129) );
  XNOR U24199 ( .A(n23131), .B(n23132), .Z(n23119) );
  AND U24200 ( .A(n23133), .B(n23134), .Z(n23131) );
  XNOR U24201 ( .A(n23132), .B(n23061), .Z(n23134) );
  XOR U24202 ( .A(n23125), .B(n23126), .Z(n23061) );
  XNOR U24203 ( .A(n23135), .B(n23136), .Z(n23126) );
  ANDN U24204 ( .B(n23137), .A(n23138), .Z(n23135) );
  XOR U24205 ( .A(n23139), .B(n23140), .Z(n23137) );
  XOR U24206 ( .A(n23141), .B(n23142), .Z(n23125) );
  XNOR U24207 ( .A(n23143), .B(n23144), .Z(n23142) );
  ANDN U24208 ( .B(n23145), .A(n23146), .Z(n23143) );
  XNOR U24209 ( .A(n23147), .B(n23148), .Z(n23145) );
  IV U24210 ( .A(n23123), .Z(n23141) );
  XOR U24211 ( .A(n23149), .B(n23150), .Z(n23123) );
  ANDN U24212 ( .B(n23151), .A(n23152), .Z(n23149) );
  XOR U24213 ( .A(n23150), .B(n23153), .Z(n23151) );
  XOR U24214 ( .A(n23132), .B(n23063), .Z(n23133) );
  XOR U24215 ( .A(n23154), .B(n23155), .Z(n23063) );
  AND U24216 ( .A(n490), .B(n23156), .Z(n23154) );
  XOR U24217 ( .A(n23157), .B(n23155), .Z(n23156) );
  XNOR U24218 ( .A(n23158), .B(n23159), .Z(n23132) );
  NAND U24219 ( .A(n23160), .B(n23161), .Z(n23159) );
  XOR U24220 ( .A(n23162), .B(n23111), .Z(n23161) );
  XOR U24221 ( .A(n23152), .B(n23153), .Z(n23111) );
  XOR U24222 ( .A(n23163), .B(n23140), .Z(n23153) );
  XOR U24223 ( .A(n23164), .B(n23165), .Z(n23140) );
  ANDN U24224 ( .B(n23166), .A(n23167), .Z(n23164) );
  XOR U24225 ( .A(n23165), .B(n23168), .Z(n23166) );
  IV U24226 ( .A(n23138), .Z(n23163) );
  XOR U24227 ( .A(n23136), .B(n23169), .Z(n23138) );
  XOR U24228 ( .A(n23170), .B(n23171), .Z(n23169) );
  ANDN U24229 ( .B(n23172), .A(n23173), .Z(n23170) );
  XOR U24230 ( .A(n23174), .B(n23171), .Z(n23172) );
  IV U24231 ( .A(n23139), .Z(n23136) );
  XOR U24232 ( .A(n23175), .B(n23176), .Z(n23139) );
  ANDN U24233 ( .B(n23177), .A(n23178), .Z(n23175) );
  XOR U24234 ( .A(n23176), .B(n23179), .Z(n23177) );
  XOR U24235 ( .A(n23180), .B(n23181), .Z(n23152) );
  XNOR U24236 ( .A(n23147), .B(n23182), .Z(n23181) );
  IV U24237 ( .A(n23150), .Z(n23182) );
  XOR U24238 ( .A(n23183), .B(n23184), .Z(n23150) );
  ANDN U24239 ( .B(n23185), .A(n23186), .Z(n23183) );
  XOR U24240 ( .A(n23184), .B(n23187), .Z(n23185) );
  XNOR U24241 ( .A(n23188), .B(n23189), .Z(n23147) );
  ANDN U24242 ( .B(n23190), .A(n23191), .Z(n23188) );
  XOR U24243 ( .A(n23189), .B(n23192), .Z(n23190) );
  IV U24244 ( .A(n23146), .Z(n23180) );
  XOR U24245 ( .A(n23144), .B(n23193), .Z(n23146) );
  XOR U24246 ( .A(n23194), .B(n23195), .Z(n23193) );
  ANDN U24247 ( .B(n23196), .A(n23197), .Z(n23194) );
  XOR U24248 ( .A(n23198), .B(n23195), .Z(n23196) );
  IV U24249 ( .A(n23148), .Z(n23144) );
  XOR U24250 ( .A(n23199), .B(n23200), .Z(n23148) );
  ANDN U24251 ( .B(n23201), .A(n23202), .Z(n23199) );
  XOR U24252 ( .A(n23203), .B(n23200), .Z(n23201) );
  IV U24253 ( .A(n23158), .Z(n23162) );
  XOR U24254 ( .A(n23158), .B(n23113), .Z(n23160) );
  XOR U24255 ( .A(n23204), .B(n23205), .Z(n23113) );
  AND U24256 ( .A(n490), .B(n23206), .Z(n23204) );
  XOR U24257 ( .A(n23207), .B(n23205), .Z(n23206) );
  NANDN U24258 ( .A(n23115), .B(n23117), .Z(n23158) );
  XOR U24259 ( .A(n23208), .B(n23209), .Z(n23117) );
  AND U24260 ( .A(n490), .B(n23210), .Z(n23208) );
  XOR U24261 ( .A(n23209), .B(n23211), .Z(n23210) );
  XNOR U24262 ( .A(n23212), .B(n23213), .Z(n490) );
  AND U24263 ( .A(n23214), .B(n23215), .Z(n23212) );
  XOR U24264 ( .A(n23213), .B(n23128), .Z(n23215) );
  XNOR U24265 ( .A(n23216), .B(n23217), .Z(n23128) );
  ANDN U24266 ( .B(n23218), .A(n23219), .Z(n23216) );
  XOR U24267 ( .A(n23217), .B(n23220), .Z(n23218) );
  XNOR U24268 ( .A(n23213), .B(n23130), .Z(n23214) );
  XOR U24269 ( .A(n23221), .B(n23222), .Z(n23130) );
  AND U24270 ( .A(n494), .B(n23223), .Z(n23221) );
  XOR U24271 ( .A(n23224), .B(n23222), .Z(n23223) );
  XNOR U24272 ( .A(n23225), .B(n23226), .Z(n23213) );
  AND U24273 ( .A(n23227), .B(n23228), .Z(n23225) );
  XNOR U24274 ( .A(n23226), .B(n23155), .Z(n23228) );
  XOR U24275 ( .A(n23219), .B(n23220), .Z(n23155) );
  XNOR U24276 ( .A(n23229), .B(n23230), .Z(n23220) );
  ANDN U24277 ( .B(n23231), .A(n23232), .Z(n23229) );
  XOR U24278 ( .A(n23233), .B(n23234), .Z(n23231) );
  XOR U24279 ( .A(n23235), .B(n23236), .Z(n23219) );
  XNOR U24280 ( .A(n23237), .B(n23238), .Z(n23236) );
  ANDN U24281 ( .B(n23239), .A(n23240), .Z(n23237) );
  XNOR U24282 ( .A(n23241), .B(n23242), .Z(n23239) );
  IV U24283 ( .A(n23217), .Z(n23235) );
  XOR U24284 ( .A(n23243), .B(n23244), .Z(n23217) );
  ANDN U24285 ( .B(n23245), .A(n23246), .Z(n23243) );
  XOR U24286 ( .A(n23244), .B(n23247), .Z(n23245) );
  XOR U24287 ( .A(n23226), .B(n23157), .Z(n23227) );
  XOR U24288 ( .A(n23248), .B(n23249), .Z(n23157) );
  AND U24289 ( .A(n494), .B(n23250), .Z(n23248) );
  XOR U24290 ( .A(n23251), .B(n23249), .Z(n23250) );
  XNOR U24291 ( .A(n23252), .B(n23253), .Z(n23226) );
  NAND U24292 ( .A(n23254), .B(n23255), .Z(n23253) );
  XOR U24293 ( .A(n23256), .B(n23205), .Z(n23255) );
  XOR U24294 ( .A(n23246), .B(n23247), .Z(n23205) );
  XOR U24295 ( .A(n23257), .B(n23234), .Z(n23247) );
  XOR U24296 ( .A(n23258), .B(n23259), .Z(n23234) );
  ANDN U24297 ( .B(n23260), .A(n23261), .Z(n23258) );
  XOR U24298 ( .A(n23259), .B(n23262), .Z(n23260) );
  IV U24299 ( .A(n23232), .Z(n23257) );
  XOR U24300 ( .A(n23230), .B(n23263), .Z(n23232) );
  XOR U24301 ( .A(n23264), .B(n23265), .Z(n23263) );
  ANDN U24302 ( .B(n23266), .A(n23267), .Z(n23264) );
  XOR U24303 ( .A(n23268), .B(n23265), .Z(n23266) );
  IV U24304 ( .A(n23233), .Z(n23230) );
  XOR U24305 ( .A(n23269), .B(n23270), .Z(n23233) );
  ANDN U24306 ( .B(n23271), .A(n23272), .Z(n23269) );
  XOR U24307 ( .A(n23270), .B(n23273), .Z(n23271) );
  XOR U24308 ( .A(n23274), .B(n23275), .Z(n23246) );
  XNOR U24309 ( .A(n23241), .B(n23276), .Z(n23275) );
  IV U24310 ( .A(n23244), .Z(n23276) );
  XOR U24311 ( .A(n23277), .B(n23278), .Z(n23244) );
  ANDN U24312 ( .B(n23279), .A(n23280), .Z(n23277) );
  XOR U24313 ( .A(n23278), .B(n23281), .Z(n23279) );
  XNOR U24314 ( .A(n23282), .B(n23283), .Z(n23241) );
  ANDN U24315 ( .B(n23284), .A(n23285), .Z(n23282) );
  XOR U24316 ( .A(n23283), .B(n23286), .Z(n23284) );
  IV U24317 ( .A(n23240), .Z(n23274) );
  XOR U24318 ( .A(n23238), .B(n23287), .Z(n23240) );
  XOR U24319 ( .A(n23288), .B(n23289), .Z(n23287) );
  ANDN U24320 ( .B(n23290), .A(n23291), .Z(n23288) );
  XOR U24321 ( .A(n23292), .B(n23289), .Z(n23290) );
  IV U24322 ( .A(n23242), .Z(n23238) );
  XOR U24323 ( .A(n23293), .B(n23294), .Z(n23242) );
  ANDN U24324 ( .B(n23295), .A(n23296), .Z(n23293) );
  XOR U24325 ( .A(n23297), .B(n23294), .Z(n23295) );
  IV U24326 ( .A(n23252), .Z(n23256) );
  XOR U24327 ( .A(n23252), .B(n23207), .Z(n23254) );
  XOR U24328 ( .A(n23298), .B(n23299), .Z(n23207) );
  AND U24329 ( .A(n494), .B(n23300), .Z(n23298) );
  XOR U24330 ( .A(n23301), .B(n23299), .Z(n23300) );
  NANDN U24331 ( .A(n23209), .B(n23211), .Z(n23252) );
  XOR U24332 ( .A(n23302), .B(n23303), .Z(n23211) );
  AND U24333 ( .A(n494), .B(n23304), .Z(n23302) );
  XOR U24334 ( .A(n23303), .B(n23305), .Z(n23304) );
  XNOR U24335 ( .A(n23306), .B(n23307), .Z(n494) );
  AND U24336 ( .A(n23308), .B(n23309), .Z(n23306) );
  XOR U24337 ( .A(n23307), .B(n23222), .Z(n23309) );
  XNOR U24338 ( .A(n23310), .B(n23311), .Z(n23222) );
  ANDN U24339 ( .B(n23312), .A(n23313), .Z(n23310) );
  XOR U24340 ( .A(n23311), .B(n23314), .Z(n23312) );
  XNOR U24341 ( .A(n23307), .B(n23224), .Z(n23308) );
  XOR U24342 ( .A(n23315), .B(n23316), .Z(n23224) );
  AND U24343 ( .A(n498), .B(n23317), .Z(n23315) );
  XOR U24344 ( .A(n23318), .B(n23316), .Z(n23317) );
  XNOR U24345 ( .A(n23319), .B(n23320), .Z(n23307) );
  AND U24346 ( .A(n23321), .B(n23322), .Z(n23319) );
  XNOR U24347 ( .A(n23320), .B(n23249), .Z(n23322) );
  XOR U24348 ( .A(n23313), .B(n23314), .Z(n23249) );
  XNOR U24349 ( .A(n23323), .B(n23324), .Z(n23314) );
  ANDN U24350 ( .B(n23325), .A(n23326), .Z(n23323) );
  XOR U24351 ( .A(n23327), .B(n23328), .Z(n23325) );
  XOR U24352 ( .A(n23329), .B(n23330), .Z(n23313) );
  XNOR U24353 ( .A(n23331), .B(n23332), .Z(n23330) );
  ANDN U24354 ( .B(n23333), .A(n23334), .Z(n23331) );
  XNOR U24355 ( .A(n23335), .B(n23336), .Z(n23333) );
  IV U24356 ( .A(n23311), .Z(n23329) );
  XOR U24357 ( .A(n23337), .B(n23338), .Z(n23311) );
  ANDN U24358 ( .B(n23339), .A(n23340), .Z(n23337) );
  XOR U24359 ( .A(n23338), .B(n23341), .Z(n23339) );
  XOR U24360 ( .A(n23320), .B(n23251), .Z(n23321) );
  XOR U24361 ( .A(n23342), .B(n23343), .Z(n23251) );
  AND U24362 ( .A(n498), .B(n23344), .Z(n23342) );
  XOR U24363 ( .A(n23345), .B(n23343), .Z(n23344) );
  XNOR U24364 ( .A(n23346), .B(n23347), .Z(n23320) );
  NAND U24365 ( .A(n23348), .B(n23349), .Z(n23347) );
  XOR U24366 ( .A(n23350), .B(n23299), .Z(n23349) );
  XOR U24367 ( .A(n23340), .B(n23341), .Z(n23299) );
  XOR U24368 ( .A(n23351), .B(n23328), .Z(n23341) );
  XOR U24369 ( .A(n23352), .B(n23353), .Z(n23328) );
  ANDN U24370 ( .B(n23354), .A(n23355), .Z(n23352) );
  XOR U24371 ( .A(n23353), .B(n23356), .Z(n23354) );
  IV U24372 ( .A(n23326), .Z(n23351) );
  XOR U24373 ( .A(n23324), .B(n23357), .Z(n23326) );
  XOR U24374 ( .A(n23358), .B(n23359), .Z(n23357) );
  ANDN U24375 ( .B(n23360), .A(n23361), .Z(n23358) );
  XOR U24376 ( .A(n23362), .B(n23359), .Z(n23360) );
  IV U24377 ( .A(n23327), .Z(n23324) );
  XOR U24378 ( .A(n23363), .B(n23364), .Z(n23327) );
  ANDN U24379 ( .B(n23365), .A(n23366), .Z(n23363) );
  XOR U24380 ( .A(n23364), .B(n23367), .Z(n23365) );
  XOR U24381 ( .A(n23368), .B(n23369), .Z(n23340) );
  XNOR U24382 ( .A(n23335), .B(n23370), .Z(n23369) );
  IV U24383 ( .A(n23338), .Z(n23370) );
  XOR U24384 ( .A(n23371), .B(n23372), .Z(n23338) );
  ANDN U24385 ( .B(n23373), .A(n23374), .Z(n23371) );
  XOR U24386 ( .A(n23372), .B(n23375), .Z(n23373) );
  XNOR U24387 ( .A(n23376), .B(n23377), .Z(n23335) );
  ANDN U24388 ( .B(n23378), .A(n23379), .Z(n23376) );
  XOR U24389 ( .A(n23377), .B(n23380), .Z(n23378) );
  IV U24390 ( .A(n23334), .Z(n23368) );
  XOR U24391 ( .A(n23332), .B(n23381), .Z(n23334) );
  XOR U24392 ( .A(n23382), .B(n23383), .Z(n23381) );
  ANDN U24393 ( .B(n23384), .A(n23385), .Z(n23382) );
  XOR U24394 ( .A(n23386), .B(n23383), .Z(n23384) );
  IV U24395 ( .A(n23336), .Z(n23332) );
  XOR U24396 ( .A(n23387), .B(n23388), .Z(n23336) );
  ANDN U24397 ( .B(n23389), .A(n23390), .Z(n23387) );
  XOR U24398 ( .A(n23391), .B(n23388), .Z(n23389) );
  IV U24399 ( .A(n23346), .Z(n23350) );
  XOR U24400 ( .A(n23346), .B(n23301), .Z(n23348) );
  XOR U24401 ( .A(n23392), .B(n23393), .Z(n23301) );
  AND U24402 ( .A(n498), .B(n23394), .Z(n23392) );
  XOR U24403 ( .A(n23395), .B(n23393), .Z(n23394) );
  NANDN U24404 ( .A(n23303), .B(n23305), .Z(n23346) );
  XOR U24405 ( .A(n23396), .B(n23397), .Z(n23305) );
  AND U24406 ( .A(n498), .B(n23398), .Z(n23396) );
  XOR U24407 ( .A(n23397), .B(n23399), .Z(n23398) );
  XNOR U24408 ( .A(n23400), .B(n23401), .Z(n498) );
  AND U24409 ( .A(n23402), .B(n23403), .Z(n23400) );
  XOR U24410 ( .A(n23401), .B(n23316), .Z(n23403) );
  XNOR U24411 ( .A(n23404), .B(n23405), .Z(n23316) );
  ANDN U24412 ( .B(n23406), .A(n23407), .Z(n23404) );
  XOR U24413 ( .A(n23405), .B(n23408), .Z(n23406) );
  XNOR U24414 ( .A(n23401), .B(n23318), .Z(n23402) );
  XOR U24415 ( .A(n23409), .B(n23410), .Z(n23318) );
  AND U24416 ( .A(n502), .B(n23411), .Z(n23409) );
  XOR U24417 ( .A(n23412), .B(n23410), .Z(n23411) );
  XNOR U24418 ( .A(n23413), .B(n23414), .Z(n23401) );
  AND U24419 ( .A(n23415), .B(n23416), .Z(n23413) );
  XNOR U24420 ( .A(n23414), .B(n23343), .Z(n23416) );
  XOR U24421 ( .A(n23407), .B(n23408), .Z(n23343) );
  XNOR U24422 ( .A(n23417), .B(n23418), .Z(n23408) );
  ANDN U24423 ( .B(n23419), .A(n23420), .Z(n23417) );
  XOR U24424 ( .A(n23421), .B(n23422), .Z(n23419) );
  XOR U24425 ( .A(n23423), .B(n23424), .Z(n23407) );
  XNOR U24426 ( .A(n23425), .B(n23426), .Z(n23424) );
  ANDN U24427 ( .B(n23427), .A(n23428), .Z(n23425) );
  XNOR U24428 ( .A(n23429), .B(n23430), .Z(n23427) );
  IV U24429 ( .A(n23405), .Z(n23423) );
  XOR U24430 ( .A(n23431), .B(n23432), .Z(n23405) );
  ANDN U24431 ( .B(n23433), .A(n23434), .Z(n23431) );
  XOR U24432 ( .A(n23432), .B(n23435), .Z(n23433) );
  XOR U24433 ( .A(n23414), .B(n23345), .Z(n23415) );
  XOR U24434 ( .A(n23436), .B(n23437), .Z(n23345) );
  AND U24435 ( .A(n502), .B(n23438), .Z(n23436) );
  XOR U24436 ( .A(n23439), .B(n23437), .Z(n23438) );
  XNOR U24437 ( .A(n23440), .B(n23441), .Z(n23414) );
  NAND U24438 ( .A(n23442), .B(n23443), .Z(n23441) );
  XOR U24439 ( .A(n23444), .B(n23393), .Z(n23443) );
  XOR U24440 ( .A(n23434), .B(n23435), .Z(n23393) );
  XOR U24441 ( .A(n23445), .B(n23422), .Z(n23435) );
  XOR U24442 ( .A(n23446), .B(n23447), .Z(n23422) );
  ANDN U24443 ( .B(n23448), .A(n23449), .Z(n23446) );
  XOR U24444 ( .A(n23447), .B(n23450), .Z(n23448) );
  IV U24445 ( .A(n23420), .Z(n23445) );
  XOR U24446 ( .A(n23418), .B(n23451), .Z(n23420) );
  XOR U24447 ( .A(n23452), .B(n23453), .Z(n23451) );
  ANDN U24448 ( .B(n23454), .A(n23455), .Z(n23452) );
  XOR U24449 ( .A(n23456), .B(n23453), .Z(n23454) );
  IV U24450 ( .A(n23421), .Z(n23418) );
  XOR U24451 ( .A(n23457), .B(n23458), .Z(n23421) );
  ANDN U24452 ( .B(n23459), .A(n23460), .Z(n23457) );
  XOR U24453 ( .A(n23458), .B(n23461), .Z(n23459) );
  XOR U24454 ( .A(n23462), .B(n23463), .Z(n23434) );
  XNOR U24455 ( .A(n23429), .B(n23464), .Z(n23463) );
  IV U24456 ( .A(n23432), .Z(n23464) );
  XOR U24457 ( .A(n23465), .B(n23466), .Z(n23432) );
  ANDN U24458 ( .B(n23467), .A(n23468), .Z(n23465) );
  XOR U24459 ( .A(n23466), .B(n23469), .Z(n23467) );
  XNOR U24460 ( .A(n23470), .B(n23471), .Z(n23429) );
  ANDN U24461 ( .B(n23472), .A(n23473), .Z(n23470) );
  XOR U24462 ( .A(n23471), .B(n23474), .Z(n23472) );
  IV U24463 ( .A(n23428), .Z(n23462) );
  XOR U24464 ( .A(n23426), .B(n23475), .Z(n23428) );
  XOR U24465 ( .A(n23476), .B(n23477), .Z(n23475) );
  ANDN U24466 ( .B(n23478), .A(n23479), .Z(n23476) );
  XOR U24467 ( .A(n23480), .B(n23477), .Z(n23478) );
  IV U24468 ( .A(n23430), .Z(n23426) );
  XOR U24469 ( .A(n23481), .B(n23482), .Z(n23430) );
  ANDN U24470 ( .B(n23483), .A(n23484), .Z(n23481) );
  XOR U24471 ( .A(n23485), .B(n23482), .Z(n23483) );
  IV U24472 ( .A(n23440), .Z(n23444) );
  XOR U24473 ( .A(n23440), .B(n23395), .Z(n23442) );
  XOR U24474 ( .A(n23486), .B(n23487), .Z(n23395) );
  AND U24475 ( .A(n502), .B(n23488), .Z(n23486) );
  XOR U24476 ( .A(n23489), .B(n23487), .Z(n23488) );
  NANDN U24477 ( .A(n23397), .B(n23399), .Z(n23440) );
  XOR U24478 ( .A(n23490), .B(n23491), .Z(n23399) );
  AND U24479 ( .A(n502), .B(n23492), .Z(n23490) );
  XOR U24480 ( .A(n23491), .B(n23493), .Z(n23492) );
  XNOR U24481 ( .A(n23494), .B(n23495), .Z(n502) );
  AND U24482 ( .A(n23496), .B(n23497), .Z(n23494) );
  XOR U24483 ( .A(n23495), .B(n23410), .Z(n23497) );
  XNOR U24484 ( .A(n23498), .B(n23499), .Z(n23410) );
  ANDN U24485 ( .B(n23500), .A(n23501), .Z(n23498) );
  XOR U24486 ( .A(n23499), .B(n23502), .Z(n23500) );
  XNOR U24487 ( .A(n23495), .B(n23412), .Z(n23496) );
  XOR U24488 ( .A(n23503), .B(n23504), .Z(n23412) );
  AND U24489 ( .A(n506), .B(n23505), .Z(n23503) );
  XOR U24490 ( .A(n23506), .B(n23504), .Z(n23505) );
  XNOR U24491 ( .A(n23507), .B(n23508), .Z(n23495) );
  AND U24492 ( .A(n23509), .B(n23510), .Z(n23507) );
  XNOR U24493 ( .A(n23508), .B(n23437), .Z(n23510) );
  XOR U24494 ( .A(n23501), .B(n23502), .Z(n23437) );
  XNOR U24495 ( .A(n23511), .B(n23512), .Z(n23502) );
  ANDN U24496 ( .B(n23513), .A(n23514), .Z(n23511) );
  XOR U24497 ( .A(n23515), .B(n23516), .Z(n23513) );
  XOR U24498 ( .A(n23517), .B(n23518), .Z(n23501) );
  XNOR U24499 ( .A(n23519), .B(n23520), .Z(n23518) );
  ANDN U24500 ( .B(n23521), .A(n23522), .Z(n23519) );
  XNOR U24501 ( .A(n23523), .B(n23524), .Z(n23521) );
  IV U24502 ( .A(n23499), .Z(n23517) );
  XOR U24503 ( .A(n23525), .B(n23526), .Z(n23499) );
  ANDN U24504 ( .B(n23527), .A(n23528), .Z(n23525) );
  XOR U24505 ( .A(n23526), .B(n23529), .Z(n23527) );
  XOR U24506 ( .A(n23508), .B(n23439), .Z(n23509) );
  XOR U24507 ( .A(n23530), .B(n23531), .Z(n23439) );
  AND U24508 ( .A(n506), .B(n23532), .Z(n23530) );
  XOR U24509 ( .A(n23533), .B(n23531), .Z(n23532) );
  XNOR U24510 ( .A(n23534), .B(n23535), .Z(n23508) );
  NAND U24511 ( .A(n23536), .B(n23537), .Z(n23535) );
  XOR U24512 ( .A(n23538), .B(n23487), .Z(n23537) );
  XOR U24513 ( .A(n23528), .B(n23529), .Z(n23487) );
  XOR U24514 ( .A(n23539), .B(n23516), .Z(n23529) );
  XOR U24515 ( .A(n23540), .B(n23541), .Z(n23516) );
  ANDN U24516 ( .B(n23542), .A(n23543), .Z(n23540) );
  XOR U24517 ( .A(n23541), .B(n23544), .Z(n23542) );
  IV U24518 ( .A(n23514), .Z(n23539) );
  XOR U24519 ( .A(n23512), .B(n23545), .Z(n23514) );
  XOR U24520 ( .A(n23546), .B(n23547), .Z(n23545) );
  ANDN U24521 ( .B(n23548), .A(n23549), .Z(n23546) );
  XOR U24522 ( .A(n23550), .B(n23547), .Z(n23548) );
  IV U24523 ( .A(n23515), .Z(n23512) );
  XOR U24524 ( .A(n23551), .B(n23552), .Z(n23515) );
  ANDN U24525 ( .B(n23553), .A(n23554), .Z(n23551) );
  XOR U24526 ( .A(n23552), .B(n23555), .Z(n23553) );
  XOR U24527 ( .A(n23556), .B(n23557), .Z(n23528) );
  XNOR U24528 ( .A(n23523), .B(n23558), .Z(n23557) );
  IV U24529 ( .A(n23526), .Z(n23558) );
  XOR U24530 ( .A(n23559), .B(n23560), .Z(n23526) );
  ANDN U24531 ( .B(n23561), .A(n23562), .Z(n23559) );
  XOR U24532 ( .A(n23560), .B(n23563), .Z(n23561) );
  XNOR U24533 ( .A(n23564), .B(n23565), .Z(n23523) );
  ANDN U24534 ( .B(n23566), .A(n23567), .Z(n23564) );
  XOR U24535 ( .A(n23565), .B(n23568), .Z(n23566) );
  IV U24536 ( .A(n23522), .Z(n23556) );
  XOR U24537 ( .A(n23520), .B(n23569), .Z(n23522) );
  XOR U24538 ( .A(n23570), .B(n23571), .Z(n23569) );
  ANDN U24539 ( .B(n23572), .A(n23573), .Z(n23570) );
  XOR U24540 ( .A(n23574), .B(n23571), .Z(n23572) );
  IV U24541 ( .A(n23524), .Z(n23520) );
  XOR U24542 ( .A(n23575), .B(n23576), .Z(n23524) );
  ANDN U24543 ( .B(n23577), .A(n23578), .Z(n23575) );
  XOR U24544 ( .A(n23579), .B(n23576), .Z(n23577) );
  IV U24545 ( .A(n23534), .Z(n23538) );
  XOR U24546 ( .A(n23534), .B(n23489), .Z(n23536) );
  XOR U24547 ( .A(n23580), .B(n23581), .Z(n23489) );
  AND U24548 ( .A(n506), .B(n23582), .Z(n23580) );
  XOR U24549 ( .A(n23583), .B(n23581), .Z(n23582) );
  NANDN U24550 ( .A(n23491), .B(n23493), .Z(n23534) );
  XOR U24551 ( .A(n23584), .B(n23585), .Z(n23493) );
  AND U24552 ( .A(n506), .B(n23586), .Z(n23584) );
  XOR U24553 ( .A(n23585), .B(n23587), .Z(n23586) );
  XNOR U24554 ( .A(n23588), .B(n23589), .Z(n506) );
  AND U24555 ( .A(n23590), .B(n23591), .Z(n23588) );
  XOR U24556 ( .A(n23589), .B(n23504), .Z(n23591) );
  XNOR U24557 ( .A(n23592), .B(n23593), .Z(n23504) );
  ANDN U24558 ( .B(n23594), .A(n23595), .Z(n23592) );
  XOR U24559 ( .A(n23593), .B(n23596), .Z(n23594) );
  XNOR U24560 ( .A(n23589), .B(n23506), .Z(n23590) );
  XOR U24561 ( .A(n23597), .B(n23598), .Z(n23506) );
  AND U24562 ( .A(n510), .B(n23599), .Z(n23597) );
  XOR U24563 ( .A(n23600), .B(n23598), .Z(n23599) );
  XNOR U24564 ( .A(n23601), .B(n23602), .Z(n23589) );
  AND U24565 ( .A(n23603), .B(n23604), .Z(n23601) );
  XNOR U24566 ( .A(n23602), .B(n23531), .Z(n23604) );
  XOR U24567 ( .A(n23595), .B(n23596), .Z(n23531) );
  XNOR U24568 ( .A(n23605), .B(n23606), .Z(n23596) );
  ANDN U24569 ( .B(n23607), .A(n23608), .Z(n23605) );
  XOR U24570 ( .A(n23609), .B(n23610), .Z(n23607) );
  XOR U24571 ( .A(n23611), .B(n23612), .Z(n23595) );
  XNOR U24572 ( .A(n23613), .B(n23614), .Z(n23612) );
  ANDN U24573 ( .B(n23615), .A(n23616), .Z(n23613) );
  XNOR U24574 ( .A(n23617), .B(n23618), .Z(n23615) );
  IV U24575 ( .A(n23593), .Z(n23611) );
  XOR U24576 ( .A(n23619), .B(n23620), .Z(n23593) );
  ANDN U24577 ( .B(n23621), .A(n23622), .Z(n23619) );
  XOR U24578 ( .A(n23620), .B(n23623), .Z(n23621) );
  XOR U24579 ( .A(n23602), .B(n23533), .Z(n23603) );
  XOR U24580 ( .A(n23624), .B(n23625), .Z(n23533) );
  AND U24581 ( .A(n510), .B(n23626), .Z(n23624) );
  XOR U24582 ( .A(n23627), .B(n23625), .Z(n23626) );
  XNOR U24583 ( .A(n23628), .B(n23629), .Z(n23602) );
  NAND U24584 ( .A(n23630), .B(n23631), .Z(n23629) );
  XOR U24585 ( .A(n23632), .B(n23581), .Z(n23631) );
  XOR U24586 ( .A(n23622), .B(n23623), .Z(n23581) );
  XOR U24587 ( .A(n23633), .B(n23610), .Z(n23623) );
  XOR U24588 ( .A(n23634), .B(n23635), .Z(n23610) );
  ANDN U24589 ( .B(n23636), .A(n23637), .Z(n23634) );
  XOR U24590 ( .A(n23635), .B(n23638), .Z(n23636) );
  IV U24591 ( .A(n23608), .Z(n23633) );
  XOR U24592 ( .A(n23606), .B(n23639), .Z(n23608) );
  XOR U24593 ( .A(n23640), .B(n23641), .Z(n23639) );
  ANDN U24594 ( .B(n23642), .A(n23643), .Z(n23640) );
  XOR U24595 ( .A(n23644), .B(n23641), .Z(n23642) );
  IV U24596 ( .A(n23609), .Z(n23606) );
  XOR U24597 ( .A(n23645), .B(n23646), .Z(n23609) );
  ANDN U24598 ( .B(n23647), .A(n23648), .Z(n23645) );
  XOR U24599 ( .A(n23646), .B(n23649), .Z(n23647) );
  XOR U24600 ( .A(n23650), .B(n23651), .Z(n23622) );
  XNOR U24601 ( .A(n23617), .B(n23652), .Z(n23651) );
  IV U24602 ( .A(n23620), .Z(n23652) );
  XOR U24603 ( .A(n23653), .B(n23654), .Z(n23620) );
  ANDN U24604 ( .B(n23655), .A(n23656), .Z(n23653) );
  XOR U24605 ( .A(n23654), .B(n23657), .Z(n23655) );
  XNOR U24606 ( .A(n23658), .B(n23659), .Z(n23617) );
  ANDN U24607 ( .B(n23660), .A(n23661), .Z(n23658) );
  XOR U24608 ( .A(n23659), .B(n23662), .Z(n23660) );
  IV U24609 ( .A(n23616), .Z(n23650) );
  XOR U24610 ( .A(n23614), .B(n23663), .Z(n23616) );
  XOR U24611 ( .A(n23664), .B(n23665), .Z(n23663) );
  ANDN U24612 ( .B(n23666), .A(n23667), .Z(n23664) );
  XOR U24613 ( .A(n23668), .B(n23665), .Z(n23666) );
  IV U24614 ( .A(n23618), .Z(n23614) );
  XOR U24615 ( .A(n23669), .B(n23670), .Z(n23618) );
  ANDN U24616 ( .B(n23671), .A(n23672), .Z(n23669) );
  XOR U24617 ( .A(n23673), .B(n23670), .Z(n23671) );
  IV U24618 ( .A(n23628), .Z(n23632) );
  XOR U24619 ( .A(n23628), .B(n23583), .Z(n23630) );
  XOR U24620 ( .A(n23674), .B(n23675), .Z(n23583) );
  AND U24621 ( .A(n510), .B(n23676), .Z(n23674) );
  XOR U24622 ( .A(n23677), .B(n23675), .Z(n23676) );
  NANDN U24623 ( .A(n23585), .B(n23587), .Z(n23628) );
  XOR U24624 ( .A(n23678), .B(n23679), .Z(n23587) );
  AND U24625 ( .A(n510), .B(n23680), .Z(n23678) );
  XOR U24626 ( .A(n23679), .B(n23681), .Z(n23680) );
  XNOR U24627 ( .A(n23682), .B(n23683), .Z(n510) );
  AND U24628 ( .A(n23684), .B(n23685), .Z(n23682) );
  XOR U24629 ( .A(n23683), .B(n23598), .Z(n23685) );
  XNOR U24630 ( .A(n23686), .B(n23687), .Z(n23598) );
  ANDN U24631 ( .B(n23688), .A(n23689), .Z(n23686) );
  XOR U24632 ( .A(n23687), .B(n23690), .Z(n23688) );
  XNOR U24633 ( .A(n23683), .B(n23600), .Z(n23684) );
  XOR U24634 ( .A(n23691), .B(n23692), .Z(n23600) );
  AND U24635 ( .A(n514), .B(n23693), .Z(n23691) );
  XOR U24636 ( .A(n23694), .B(n23692), .Z(n23693) );
  XNOR U24637 ( .A(n23695), .B(n23696), .Z(n23683) );
  AND U24638 ( .A(n23697), .B(n23698), .Z(n23695) );
  XNOR U24639 ( .A(n23696), .B(n23625), .Z(n23698) );
  XOR U24640 ( .A(n23689), .B(n23690), .Z(n23625) );
  XNOR U24641 ( .A(n23699), .B(n23700), .Z(n23690) );
  ANDN U24642 ( .B(n23701), .A(n23702), .Z(n23699) );
  XOR U24643 ( .A(n23703), .B(n23704), .Z(n23701) );
  XOR U24644 ( .A(n23705), .B(n23706), .Z(n23689) );
  XNOR U24645 ( .A(n23707), .B(n23708), .Z(n23706) );
  ANDN U24646 ( .B(n23709), .A(n23710), .Z(n23707) );
  XNOR U24647 ( .A(n23711), .B(n23712), .Z(n23709) );
  IV U24648 ( .A(n23687), .Z(n23705) );
  XOR U24649 ( .A(n23713), .B(n23714), .Z(n23687) );
  ANDN U24650 ( .B(n23715), .A(n23716), .Z(n23713) );
  XOR U24651 ( .A(n23714), .B(n23717), .Z(n23715) );
  XOR U24652 ( .A(n23696), .B(n23627), .Z(n23697) );
  XOR U24653 ( .A(n23718), .B(n23719), .Z(n23627) );
  AND U24654 ( .A(n514), .B(n23720), .Z(n23718) );
  XOR U24655 ( .A(n23721), .B(n23719), .Z(n23720) );
  XNOR U24656 ( .A(n23722), .B(n23723), .Z(n23696) );
  NAND U24657 ( .A(n23724), .B(n23725), .Z(n23723) );
  XOR U24658 ( .A(n23726), .B(n23675), .Z(n23725) );
  XOR U24659 ( .A(n23716), .B(n23717), .Z(n23675) );
  XOR U24660 ( .A(n23727), .B(n23704), .Z(n23717) );
  XOR U24661 ( .A(n23728), .B(n23729), .Z(n23704) );
  ANDN U24662 ( .B(n23730), .A(n23731), .Z(n23728) );
  XOR U24663 ( .A(n23729), .B(n23732), .Z(n23730) );
  IV U24664 ( .A(n23702), .Z(n23727) );
  XOR U24665 ( .A(n23700), .B(n23733), .Z(n23702) );
  XOR U24666 ( .A(n23734), .B(n23735), .Z(n23733) );
  ANDN U24667 ( .B(n23736), .A(n23737), .Z(n23734) );
  XOR U24668 ( .A(n23738), .B(n23735), .Z(n23736) );
  IV U24669 ( .A(n23703), .Z(n23700) );
  XOR U24670 ( .A(n23739), .B(n23740), .Z(n23703) );
  ANDN U24671 ( .B(n23741), .A(n23742), .Z(n23739) );
  XOR U24672 ( .A(n23740), .B(n23743), .Z(n23741) );
  XOR U24673 ( .A(n23744), .B(n23745), .Z(n23716) );
  XNOR U24674 ( .A(n23711), .B(n23746), .Z(n23745) );
  IV U24675 ( .A(n23714), .Z(n23746) );
  XOR U24676 ( .A(n23747), .B(n23748), .Z(n23714) );
  ANDN U24677 ( .B(n23749), .A(n23750), .Z(n23747) );
  XOR U24678 ( .A(n23748), .B(n23751), .Z(n23749) );
  XNOR U24679 ( .A(n23752), .B(n23753), .Z(n23711) );
  ANDN U24680 ( .B(n23754), .A(n23755), .Z(n23752) );
  XOR U24681 ( .A(n23753), .B(n23756), .Z(n23754) );
  IV U24682 ( .A(n23710), .Z(n23744) );
  XOR U24683 ( .A(n23708), .B(n23757), .Z(n23710) );
  XOR U24684 ( .A(n23758), .B(n23759), .Z(n23757) );
  ANDN U24685 ( .B(n23760), .A(n23761), .Z(n23758) );
  XOR U24686 ( .A(n23762), .B(n23759), .Z(n23760) );
  IV U24687 ( .A(n23712), .Z(n23708) );
  XOR U24688 ( .A(n23763), .B(n23764), .Z(n23712) );
  ANDN U24689 ( .B(n23765), .A(n23766), .Z(n23763) );
  XOR U24690 ( .A(n23767), .B(n23764), .Z(n23765) );
  IV U24691 ( .A(n23722), .Z(n23726) );
  XOR U24692 ( .A(n23722), .B(n23677), .Z(n23724) );
  XOR U24693 ( .A(n23768), .B(n23769), .Z(n23677) );
  AND U24694 ( .A(n514), .B(n23770), .Z(n23768) );
  XOR U24695 ( .A(n23771), .B(n23769), .Z(n23770) );
  NANDN U24696 ( .A(n23679), .B(n23681), .Z(n23722) );
  XOR U24697 ( .A(n23772), .B(n23773), .Z(n23681) );
  AND U24698 ( .A(n514), .B(n23774), .Z(n23772) );
  XOR U24699 ( .A(n23773), .B(n23775), .Z(n23774) );
  XNOR U24700 ( .A(n23776), .B(n23777), .Z(n514) );
  AND U24701 ( .A(n23778), .B(n23779), .Z(n23776) );
  XOR U24702 ( .A(n23777), .B(n23692), .Z(n23779) );
  XNOR U24703 ( .A(n23780), .B(n23781), .Z(n23692) );
  ANDN U24704 ( .B(n23782), .A(n23783), .Z(n23780) );
  XOR U24705 ( .A(n23781), .B(n23784), .Z(n23782) );
  XNOR U24706 ( .A(n23777), .B(n23694), .Z(n23778) );
  XOR U24707 ( .A(n23785), .B(n23786), .Z(n23694) );
  AND U24708 ( .A(n518), .B(n23787), .Z(n23785) );
  XOR U24709 ( .A(n23788), .B(n23786), .Z(n23787) );
  XNOR U24710 ( .A(n23789), .B(n23790), .Z(n23777) );
  AND U24711 ( .A(n23791), .B(n23792), .Z(n23789) );
  XNOR U24712 ( .A(n23790), .B(n23719), .Z(n23792) );
  XOR U24713 ( .A(n23783), .B(n23784), .Z(n23719) );
  XNOR U24714 ( .A(n23793), .B(n23794), .Z(n23784) );
  ANDN U24715 ( .B(n23795), .A(n23796), .Z(n23793) );
  XOR U24716 ( .A(n23797), .B(n23798), .Z(n23795) );
  XOR U24717 ( .A(n23799), .B(n23800), .Z(n23783) );
  XNOR U24718 ( .A(n23801), .B(n23802), .Z(n23800) );
  ANDN U24719 ( .B(n23803), .A(n23804), .Z(n23801) );
  XNOR U24720 ( .A(n23805), .B(n23806), .Z(n23803) );
  IV U24721 ( .A(n23781), .Z(n23799) );
  XOR U24722 ( .A(n23807), .B(n23808), .Z(n23781) );
  ANDN U24723 ( .B(n23809), .A(n23810), .Z(n23807) );
  XOR U24724 ( .A(n23808), .B(n23811), .Z(n23809) );
  XOR U24725 ( .A(n23790), .B(n23721), .Z(n23791) );
  XOR U24726 ( .A(n23812), .B(n23813), .Z(n23721) );
  AND U24727 ( .A(n518), .B(n23814), .Z(n23812) );
  XOR U24728 ( .A(n23815), .B(n23813), .Z(n23814) );
  XNOR U24729 ( .A(n23816), .B(n23817), .Z(n23790) );
  NAND U24730 ( .A(n23818), .B(n23819), .Z(n23817) );
  XOR U24731 ( .A(n23820), .B(n23769), .Z(n23819) );
  XOR U24732 ( .A(n23810), .B(n23811), .Z(n23769) );
  XOR U24733 ( .A(n23821), .B(n23798), .Z(n23811) );
  XOR U24734 ( .A(n23822), .B(n23823), .Z(n23798) );
  ANDN U24735 ( .B(n23824), .A(n23825), .Z(n23822) );
  XOR U24736 ( .A(n23823), .B(n23826), .Z(n23824) );
  IV U24737 ( .A(n23796), .Z(n23821) );
  XOR U24738 ( .A(n23794), .B(n23827), .Z(n23796) );
  XOR U24739 ( .A(n23828), .B(n23829), .Z(n23827) );
  ANDN U24740 ( .B(n23830), .A(n23831), .Z(n23828) );
  XOR U24741 ( .A(n23832), .B(n23829), .Z(n23830) );
  IV U24742 ( .A(n23797), .Z(n23794) );
  XOR U24743 ( .A(n23833), .B(n23834), .Z(n23797) );
  ANDN U24744 ( .B(n23835), .A(n23836), .Z(n23833) );
  XOR U24745 ( .A(n23834), .B(n23837), .Z(n23835) );
  XOR U24746 ( .A(n23838), .B(n23839), .Z(n23810) );
  XNOR U24747 ( .A(n23805), .B(n23840), .Z(n23839) );
  IV U24748 ( .A(n23808), .Z(n23840) );
  XOR U24749 ( .A(n23841), .B(n23842), .Z(n23808) );
  ANDN U24750 ( .B(n23843), .A(n23844), .Z(n23841) );
  XOR U24751 ( .A(n23842), .B(n23845), .Z(n23843) );
  XNOR U24752 ( .A(n23846), .B(n23847), .Z(n23805) );
  ANDN U24753 ( .B(n23848), .A(n23849), .Z(n23846) );
  XOR U24754 ( .A(n23847), .B(n23850), .Z(n23848) );
  IV U24755 ( .A(n23804), .Z(n23838) );
  XOR U24756 ( .A(n23802), .B(n23851), .Z(n23804) );
  XOR U24757 ( .A(n23852), .B(n23853), .Z(n23851) );
  ANDN U24758 ( .B(n23854), .A(n23855), .Z(n23852) );
  XOR U24759 ( .A(n23856), .B(n23853), .Z(n23854) );
  IV U24760 ( .A(n23806), .Z(n23802) );
  XOR U24761 ( .A(n23857), .B(n23858), .Z(n23806) );
  ANDN U24762 ( .B(n23859), .A(n23860), .Z(n23857) );
  XOR U24763 ( .A(n23861), .B(n23858), .Z(n23859) );
  IV U24764 ( .A(n23816), .Z(n23820) );
  XOR U24765 ( .A(n23816), .B(n23771), .Z(n23818) );
  XOR U24766 ( .A(n23862), .B(n23863), .Z(n23771) );
  AND U24767 ( .A(n518), .B(n23864), .Z(n23862) );
  XOR U24768 ( .A(n23865), .B(n23863), .Z(n23864) );
  NANDN U24769 ( .A(n23773), .B(n23775), .Z(n23816) );
  XOR U24770 ( .A(n23866), .B(n23867), .Z(n23775) );
  AND U24771 ( .A(n518), .B(n23868), .Z(n23866) );
  XOR U24772 ( .A(n23867), .B(n23869), .Z(n23868) );
  XNOR U24773 ( .A(n23870), .B(n23871), .Z(n518) );
  AND U24774 ( .A(n23872), .B(n23873), .Z(n23870) );
  XOR U24775 ( .A(n23871), .B(n23786), .Z(n23873) );
  XNOR U24776 ( .A(n23874), .B(n23875), .Z(n23786) );
  ANDN U24777 ( .B(n23876), .A(n23877), .Z(n23874) );
  XOR U24778 ( .A(n23875), .B(n23878), .Z(n23876) );
  XNOR U24779 ( .A(n23871), .B(n23788), .Z(n23872) );
  XOR U24780 ( .A(n23879), .B(n23880), .Z(n23788) );
  AND U24781 ( .A(n522), .B(n23881), .Z(n23879) );
  XOR U24782 ( .A(n23882), .B(n23880), .Z(n23881) );
  XNOR U24783 ( .A(n23883), .B(n23884), .Z(n23871) );
  AND U24784 ( .A(n23885), .B(n23886), .Z(n23883) );
  XNOR U24785 ( .A(n23884), .B(n23813), .Z(n23886) );
  XOR U24786 ( .A(n23877), .B(n23878), .Z(n23813) );
  XNOR U24787 ( .A(n23887), .B(n23888), .Z(n23878) );
  ANDN U24788 ( .B(n23889), .A(n23890), .Z(n23887) );
  XOR U24789 ( .A(n23891), .B(n23892), .Z(n23889) );
  XOR U24790 ( .A(n23893), .B(n23894), .Z(n23877) );
  XNOR U24791 ( .A(n23895), .B(n23896), .Z(n23894) );
  ANDN U24792 ( .B(n23897), .A(n23898), .Z(n23895) );
  XNOR U24793 ( .A(n23899), .B(n23900), .Z(n23897) );
  IV U24794 ( .A(n23875), .Z(n23893) );
  XOR U24795 ( .A(n23901), .B(n23902), .Z(n23875) );
  ANDN U24796 ( .B(n23903), .A(n23904), .Z(n23901) );
  XOR U24797 ( .A(n23902), .B(n23905), .Z(n23903) );
  XOR U24798 ( .A(n23884), .B(n23815), .Z(n23885) );
  XOR U24799 ( .A(n23906), .B(n23907), .Z(n23815) );
  AND U24800 ( .A(n522), .B(n23908), .Z(n23906) );
  XOR U24801 ( .A(n23909), .B(n23907), .Z(n23908) );
  XNOR U24802 ( .A(n23910), .B(n23911), .Z(n23884) );
  NAND U24803 ( .A(n23912), .B(n23913), .Z(n23911) );
  XOR U24804 ( .A(n23914), .B(n23863), .Z(n23913) );
  XOR U24805 ( .A(n23904), .B(n23905), .Z(n23863) );
  XOR U24806 ( .A(n23915), .B(n23892), .Z(n23905) );
  XOR U24807 ( .A(n23916), .B(n23917), .Z(n23892) );
  ANDN U24808 ( .B(n23918), .A(n23919), .Z(n23916) );
  XOR U24809 ( .A(n23917), .B(n23920), .Z(n23918) );
  IV U24810 ( .A(n23890), .Z(n23915) );
  XOR U24811 ( .A(n23888), .B(n23921), .Z(n23890) );
  XOR U24812 ( .A(n23922), .B(n23923), .Z(n23921) );
  ANDN U24813 ( .B(n23924), .A(n23925), .Z(n23922) );
  XOR U24814 ( .A(n23926), .B(n23923), .Z(n23924) );
  IV U24815 ( .A(n23891), .Z(n23888) );
  XOR U24816 ( .A(n23927), .B(n23928), .Z(n23891) );
  ANDN U24817 ( .B(n23929), .A(n23930), .Z(n23927) );
  XOR U24818 ( .A(n23928), .B(n23931), .Z(n23929) );
  XOR U24819 ( .A(n23932), .B(n23933), .Z(n23904) );
  XNOR U24820 ( .A(n23899), .B(n23934), .Z(n23933) );
  IV U24821 ( .A(n23902), .Z(n23934) );
  XOR U24822 ( .A(n23935), .B(n23936), .Z(n23902) );
  ANDN U24823 ( .B(n23937), .A(n23938), .Z(n23935) );
  XOR U24824 ( .A(n23936), .B(n23939), .Z(n23937) );
  XNOR U24825 ( .A(n23940), .B(n23941), .Z(n23899) );
  ANDN U24826 ( .B(n23942), .A(n23943), .Z(n23940) );
  XOR U24827 ( .A(n23941), .B(n23944), .Z(n23942) );
  IV U24828 ( .A(n23898), .Z(n23932) );
  XOR U24829 ( .A(n23896), .B(n23945), .Z(n23898) );
  XOR U24830 ( .A(n23946), .B(n23947), .Z(n23945) );
  ANDN U24831 ( .B(n23948), .A(n23949), .Z(n23946) );
  XOR U24832 ( .A(n23950), .B(n23947), .Z(n23948) );
  IV U24833 ( .A(n23900), .Z(n23896) );
  XOR U24834 ( .A(n23951), .B(n23952), .Z(n23900) );
  ANDN U24835 ( .B(n23953), .A(n23954), .Z(n23951) );
  XOR U24836 ( .A(n23955), .B(n23952), .Z(n23953) );
  IV U24837 ( .A(n23910), .Z(n23914) );
  XOR U24838 ( .A(n23910), .B(n23865), .Z(n23912) );
  XOR U24839 ( .A(n23956), .B(n23957), .Z(n23865) );
  AND U24840 ( .A(n522), .B(n23958), .Z(n23956) );
  XOR U24841 ( .A(n23959), .B(n23957), .Z(n23958) );
  NANDN U24842 ( .A(n23867), .B(n23869), .Z(n23910) );
  XOR U24843 ( .A(n23960), .B(n23961), .Z(n23869) );
  AND U24844 ( .A(n522), .B(n23962), .Z(n23960) );
  XOR U24845 ( .A(n23961), .B(n23963), .Z(n23962) );
  XNOR U24846 ( .A(n23964), .B(n23965), .Z(n522) );
  AND U24847 ( .A(n23966), .B(n23967), .Z(n23964) );
  XOR U24848 ( .A(n23965), .B(n23880), .Z(n23967) );
  XNOR U24849 ( .A(n23968), .B(n23969), .Z(n23880) );
  ANDN U24850 ( .B(n23970), .A(n23971), .Z(n23968) );
  XOR U24851 ( .A(n23969), .B(n23972), .Z(n23970) );
  XNOR U24852 ( .A(n23965), .B(n23882), .Z(n23966) );
  XOR U24853 ( .A(n23973), .B(n23974), .Z(n23882) );
  AND U24854 ( .A(n526), .B(n23975), .Z(n23973) );
  XOR U24855 ( .A(n23976), .B(n23974), .Z(n23975) );
  XNOR U24856 ( .A(n23977), .B(n23978), .Z(n23965) );
  AND U24857 ( .A(n23979), .B(n23980), .Z(n23977) );
  XNOR U24858 ( .A(n23978), .B(n23907), .Z(n23980) );
  XOR U24859 ( .A(n23971), .B(n23972), .Z(n23907) );
  XNOR U24860 ( .A(n23981), .B(n23982), .Z(n23972) );
  ANDN U24861 ( .B(n23983), .A(n23984), .Z(n23981) );
  XOR U24862 ( .A(n23985), .B(n23986), .Z(n23983) );
  XOR U24863 ( .A(n23987), .B(n23988), .Z(n23971) );
  XNOR U24864 ( .A(n23989), .B(n23990), .Z(n23988) );
  ANDN U24865 ( .B(n23991), .A(n23992), .Z(n23989) );
  XNOR U24866 ( .A(n23993), .B(n23994), .Z(n23991) );
  IV U24867 ( .A(n23969), .Z(n23987) );
  XOR U24868 ( .A(n23995), .B(n23996), .Z(n23969) );
  ANDN U24869 ( .B(n23997), .A(n23998), .Z(n23995) );
  XOR U24870 ( .A(n23996), .B(n23999), .Z(n23997) );
  XOR U24871 ( .A(n23978), .B(n23909), .Z(n23979) );
  XOR U24872 ( .A(n24000), .B(n24001), .Z(n23909) );
  AND U24873 ( .A(n526), .B(n24002), .Z(n24000) );
  XOR U24874 ( .A(n24003), .B(n24001), .Z(n24002) );
  XNOR U24875 ( .A(n24004), .B(n24005), .Z(n23978) );
  NAND U24876 ( .A(n24006), .B(n24007), .Z(n24005) );
  XOR U24877 ( .A(n24008), .B(n23957), .Z(n24007) );
  XOR U24878 ( .A(n23998), .B(n23999), .Z(n23957) );
  XOR U24879 ( .A(n24009), .B(n23986), .Z(n23999) );
  XOR U24880 ( .A(n24010), .B(n24011), .Z(n23986) );
  ANDN U24881 ( .B(n24012), .A(n24013), .Z(n24010) );
  XOR U24882 ( .A(n24011), .B(n24014), .Z(n24012) );
  IV U24883 ( .A(n23984), .Z(n24009) );
  XOR U24884 ( .A(n23982), .B(n24015), .Z(n23984) );
  XOR U24885 ( .A(n24016), .B(n24017), .Z(n24015) );
  ANDN U24886 ( .B(n24018), .A(n24019), .Z(n24016) );
  XOR U24887 ( .A(n24020), .B(n24017), .Z(n24018) );
  IV U24888 ( .A(n23985), .Z(n23982) );
  XOR U24889 ( .A(n24021), .B(n24022), .Z(n23985) );
  ANDN U24890 ( .B(n24023), .A(n24024), .Z(n24021) );
  XOR U24891 ( .A(n24022), .B(n24025), .Z(n24023) );
  XOR U24892 ( .A(n24026), .B(n24027), .Z(n23998) );
  XNOR U24893 ( .A(n23993), .B(n24028), .Z(n24027) );
  IV U24894 ( .A(n23996), .Z(n24028) );
  XOR U24895 ( .A(n24029), .B(n24030), .Z(n23996) );
  ANDN U24896 ( .B(n24031), .A(n24032), .Z(n24029) );
  XOR U24897 ( .A(n24030), .B(n24033), .Z(n24031) );
  XNOR U24898 ( .A(n24034), .B(n24035), .Z(n23993) );
  ANDN U24899 ( .B(n24036), .A(n24037), .Z(n24034) );
  XOR U24900 ( .A(n24035), .B(n24038), .Z(n24036) );
  IV U24901 ( .A(n23992), .Z(n24026) );
  XOR U24902 ( .A(n23990), .B(n24039), .Z(n23992) );
  XOR U24903 ( .A(n24040), .B(n24041), .Z(n24039) );
  ANDN U24904 ( .B(n24042), .A(n24043), .Z(n24040) );
  XOR U24905 ( .A(n24044), .B(n24041), .Z(n24042) );
  IV U24906 ( .A(n23994), .Z(n23990) );
  XOR U24907 ( .A(n24045), .B(n24046), .Z(n23994) );
  ANDN U24908 ( .B(n24047), .A(n24048), .Z(n24045) );
  XOR U24909 ( .A(n24049), .B(n24046), .Z(n24047) );
  IV U24910 ( .A(n24004), .Z(n24008) );
  XOR U24911 ( .A(n24004), .B(n23959), .Z(n24006) );
  XOR U24912 ( .A(n24050), .B(n24051), .Z(n23959) );
  AND U24913 ( .A(n526), .B(n24052), .Z(n24050) );
  XOR U24914 ( .A(n24053), .B(n24051), .Z(n24052) );
  NANDN U24915 ( .A(n23961), .B(n23963), .Z(n24004) );
  XOR U24916 ( .A(n24054), .B(n24055), .Z(n23963) );
  AND U24917 ( .A(n526), .B(n24056), .Z(n24054) );
  XOR U24918 ( .A(n24055), .B(n24057), .Z(n24056) );
  XNOR U24919 ( .A(n24058), .B(n24059), .Z(n526) );
  AND U24920 ( .A(n24060), .B(n24061), .Z(n24058) );
  XOR U24921 ( .A(n24059), .B(n23974), .Z(n24061) );
  XNOR U24922 ( .A(n24062), .B(n24063), .Z(n23974) );
  ANDN U24923 ( .B(n24064), .A(n24065), .Z(n24062) );
  XOR U24924 ( .A(n24063), .B(n24066), .Z(n24064) );
  XNOR U24925 ( .A(n24059), .B(n23976), .Z(n24060) );
  XOR U24926 ( .A(n24067), .B(n24068), .Z(n23976) );
  AND U24927 ( .A(n530), .B(n24069), .Z(n24067) );
  XOR U24928 ( .A(n24070), .B(n24068), .Z(n24069) );
  XNOR U24929 ( .A(n24071), .B(n24072), .Z(n24059) );
  AND U24930 ( .A(n24073), .B(n24074), .Z(n24071) );
  XNOR U24931 ( .A(n24072), .B(n24001), .Z(n24074) );
  XOR U24932 ( .A(n24065), .B(n24066), .Z(n24001) );
  XNOR U24933 ( .A(n24075), .B(n24076), .Z(n24066) );
  ANDN U24934 ( .B(n24077), .A(n24078), .Z(n24075) );
  XOR U24935 ( .A(n24079), .B(n24080), .Z(n24077) );
  XOR U24936 ( .A(n24081), .B(n24082), .Z(n24065) );
  XNOR U24937 ( .A(n24083), .B(n24084), .Z(n24082) );
  ANDN U24938 ( .B(n24085), .A(n24086), .Z(n24083) );
  XNOR U24939 ( .A(n24087), .B(n24088), .Z(n24085) );
  IV U24940 ( .A(n24063), .Z(n24081) );
  XOR U24941 ( .A(n24089), .B(n24090), .Z(n24063) );
  ANDN U24942 ( .B(n24091), .A(n24092), .Z(n24089) );
  XOR U24943 ( .A(n24090), .B(n24093), .Z(n24091) );
  XOR U24944 ( .A(n24072), .B(n24003), .Z(n24073) );
  XOR U24945 ( .A(n24094), .B(n24095), .Z(n24003) );
  AND U24946 ( .A(n530), .B(n24096), .Z(n24094) );
  XOR U24947 ( .A(n24097), .B(n24095), .Z(n24096) );
  XNOR U24948 ( .A(n24098), .B(n24099), .Z(n24072) );
  NAND U24949 ( .A(n24100), .B(n24101), .Z(n24099) );
  XOR U24950 ( .A(n24102), .B(n24051), .Z(n24101) );
  XOR U24951 ( .A(n24092), .B(n24093), .Z(n24051) );
  XOR U24952 ( .A(n24103), .B(n24080), .Z(n24093) );
  XOR U24953 ( .A(n24104), .B(n24105), .Z(n24080) );
  ANDN U24954 ( .B(n24106), .A(n24107), .Z(n24104) );
  XOR U24955 ( .A(n24105), .B(n24108), .Z(n24106) );
  IV U24956 ( .A(n24078), .Z(n24103) );
  XOR U24957 ( .A(n24076), .B(n24109), .Z(n24078) );
  XOR U24958 ( .A(n24110), .B(n24111), .Z(n24109) );
  ANDN U24959 ( .B(n24112), .A(n24113), .Z(n24110) );
  XOR U24960 ( .A(n24114), .B(n24111), .Z(n24112) );
  IV U24961 ( .A(n24079), .Z(n24076) );
  XOR U24962 ( .A(n24115), .B(n24116), .Z(n24079) );
  ANDN U24963 ( .B(n24117), .A(n24118), .Z(n24115) );
  XOR U24964 ( .A(n24116), .B(n24119), .Z(n24117) );
  XOR U24965 ( .A(n24120), .B(n24121), .Z(n24092) );
  XNOR U24966 ( .A(n24087), .B(n24122), .Z(n24121) );
  IV U24967 ( .A(n24090), .Z(n24122) );
  XOR U24968 ( .A(n24123), .B(n24124), .Z(n24090) );
  ANDN U24969 ( .B(n24125), .A(n24126), .Z(n24123) );
  XOR U24970 ( .A(n24124), .B(n24127), .Z(n24125) );
  XNOR U24971 ( .A(n24128), .B(n24129), .Z(n24087) );
  ANDN U24972 ( .B(n24130), .A(n24131), .Z(n24128) );
  XOR U24973 ( .A(n24129), .B(n24132), .Z(n24130) );
  IV U24974 ( .A(n24086), .Z(n24120) );
  XOR U24975 ( .A(n24084), .B(n24133), .Z(n24086) );
  XOR U24976 ( .A(n24134), .B(n24135), .Z(n24133) );
  ANDN U24977 ( .B(n24136), .A(n24137), .Z(n24134) );
  XOR U24978 ( .A(n24138), .B(n24135), .Z(n24136) );
  IV U24979 ( .A(n24088), .Z(n24084) );
  XOR U24980 ( .A(n24139), .B(n24140), .Z(n24088) );
  ANDN U24981 ( .B(n24141), .A(n24142), .Z(n24139) );
  XOR U24982 ( .A(n24143), .B(n24140), .Z(n24141) );
  IV U24983 ( .A(n24098), .Z(n24102) );
  XOR U24984 ( .A(n24098), .B(n24053), .Z(n24100) );
  XOR U24985 ( .A(n24144), .B(n24145), .Z(n24053) );
  AND U24986 ( .A(n530), .B(n24146), .Z(n24144) );
  XOR U24987 ( .A(n24147), .B(n24145), .Z(n24146) );
  NANDN U24988 ( .A(n24055), .B(n24057), .Z(n24098) );
  XOR U24989 ( .A(n24148), .B(n24149), .Z(n24057) );
  AND U24990 ( .A(n530), .B(n24150), .Z(n24148) );
  XOR U24991 ( .A(n24149), .B(n24151), .Z(n24150) );
  XNOR U24992 ( .A(n24152), .B(n24153), .Z(n530) );
  AND U24993 ( .A(n24154), .B(n24155), .Z(n24152) );
  XOR U24994 ( .A(n24153), .B(n24068), .Z(n24155) );
  XNOR U24995 ( .A(n24156), .B(n24157), .Z(n24068) );
  ANDN U24996 ( .B(n24158), .A(n24159), .Z(n24156) );
  XOR U24997 ( .A(n24157), .B(n24160), .Z(n24158) );
  XNOR U24998 ( .A(n24153), .B(n24070), .Z(n24154) );
  XOR U24999 ( .A(n24161), .B(n24162), .Z(n24070) );
  AND U25000 ( .A(n534), .B(n24163), .Z(n24161) );
  XOR U25001 ( .A(n24164), .B(n24162), .Z(n24163) );
  XNOR U25002 ( .A(n24165), .B(n24166), .Z(n24153) );
  AND U25003 ( .A(n24167), .B(n24168), .Z(n24165) );
  XNOR U25004 ( .A(n24166), .B(n24095), .Z(n24168) );
  XOR U25005 ( .A(n24159), .B(n24160), .Z(n24095) );
  XNOR U25006 ( .A(n24169), .B(n24170), .Z(n24160) );
  ANDN U25007 ( .B(n24171), .A(n24172), .Z(n24169) );
  XOR U25008 ( .A(n24173), .B(n24174), .Z(n24171) );
  XOR U25009 ( .A(n24175), .B(n24176), .Z(n24159) );
  XNOR U25010 ( .A(n24177), .B(n24178), .Z(n24176) );
  ANDN U25011 ( .B(n24179), .A(n24180), .Z(n24177) );
  XNOR U25012 ( .A(n24181), .B(n24182), .Z(n24179) );
  IV U25013 ( .A(n24157), .Z(n24175) );
  XOR U25014 ( .A(n24183), .B(n24184), .Z(n24157) );
  ANDN U25015 ( .B(n24185), .A(n24186), .Z(n24183) );
  XOR U25016 ( .A(n24184), .B(n24187), .Z(n24185) );
  XOR U25017 ( .A(n24166), .B(n24097), .Z(n24167) );
  XOR U25018 ( .A(n24188), .B(n24189), .Z(n24097) );
  AND U25019 ( .A(n534), .B(n24190), .Z(n24188) );
  XOR U25020 ( .A(n24191), .B(n24189), .Z(n24190) );
  XNOR U25021 ( .A(n24192), .B(n24193), .Z(n24166) );
  NAND U25022 ( .A(n24194), .B(n24195), .Z(n24193) );
  XOR U25023 ( .A(n24196), .B(n24145), .Z(n24195) );
  XOR U25024 ( .A(n24186), .B(n24187), .Z(n24145) );
  XOR U25025 ( .A(n24197), .B(n24174), .Z(n24187) );
  XOR U25026 ( .A(n24198), .B(n24199), .Z(n24174) );
  ANDN U25027 ( .B(n24200), .A(n24201), .Z(n24198) );
  XOR U25028 ( .A(n24199), .B(n24202), .Z(n24200) );
  IV U25029 ( .A(n24172), .Z(n24197) );
  XOR U25030 ( .A(n24170), .B(n24203), .Z(n24172) );
  XOR U25031 ( .A(n24204), .B(n24205), .Z(n24203) );
  ANDN U25032 ( .B(n24206), .A(n24207), .Z(n24204) );
  XOR U25033 ( .A(n24208), .B(n24205), .Z(n24206) );
  IV U25034 ( .A(n24173), .Z(n24170) );
  XOR U25035 ( .A(n24209), .B(n24210), .Z(n24173) );
  ANDN U25036 ( .B(n24211), .A(n24212), .Z(n24209) );
  XOR U25037 ( .A(n24210), .B(n24213), .Z(n24211) );
  XOR U25038 ( .A(n24214), .B(n24215), .Z(n24186) );
  XNOR U25039 ( .A(n24181), .B(n24216), .Z(n24215) );
  IV U25040 ( .A(n24184), .Z(n24216) );
  XOR U25041 ( .A(n24217), .B(n24218), .Z(n24184) );
  ANDN U25042 ( .B(n24219), .A(n24220), .Z(n24217) );
  XOR U25043 ( .A(n24218), .B(n24221), .Z(n24219) );
  XNOR U25044 ( .A(n24222), .B(n24223), .Z(n24181) );
  ANDN U25045 ( .B(n24224), .A(n24225), .Z(n24222) );
  XOR U25046 ( .A(n24223), .B(n24226), .Z(n24224) );
  IV U25047 ( .A(n24180), .Z(n24214) );
  XOR U25048 ( .A(n24178), .B(n24227), .Z(n24180) );
  XOR U25049 ( .A(n24228), .B(n24229), .Z(n24227) );
  ANDN U25050 ( .B(n24230), .A(n24231), .Z(n24228) );
  XOR U25051 ( .A(n24232), .B(n24229), .Z(n24230) );
  IV U25052 ( .A(n24182), .Z(n24178) );
  XOR U25053 ( .A(n24233), .B(n24234), .Z(n24182) );
  ANDN U25054 ( .B(n24235), .A(n24236), .Z(n24233) );
  XOR U25055 ( .A(n24237), .B(n24234), .Z(n24235) );
  IV U25056 ( .A(n24192), .Z(n24196) );
  XOR U25057 ( .A(n24192), .B(n24147), .Z(n24194) );
  XOR U25058 ( .A(n24238), .B(n24239), .Z(n24147) );
  AND U25059 ( .A(n534), .B(n24240), .Z(n24238) );
  XOR U25060 ( .A(n24241), .B(n24239), .Z(n24240) );
  NANDN U25061 ( .A(n24149), .B(n24151), .Z(n24192) );
  XOR U25062 ( .A(n24242), .B(n24243), .Z(n24151) );
  AND U25063 ( .A(n534), .B(n24244), .Z(n24242) );
  XOR U25064 ( .A(n24243), .B(n24245), .Z(n24244) );
  XNOR U25065 ( .A(n24246), .B(n24247), .Z(n534) );
  AND U25066 ( .A(n24248), .B(n24249), .Z(n24246) );
  XOR U25067 ( .A(n24247), .B(n24162), .Z(n24249) );
  XNOR U25068 ( .A(n24250), .B(n24251), .Z(n24162) );
  ANDN U25069 ( .B(n24252), .A(n24253), .Z(n24250) );
  XOR U25070 ( .A(n24251), .B(n24254), .Z(n24252) );
  XNOR U25071 ( .A(n24247), .B(n24164), .Z(n24248) );
  XOR U25072 ( .A(n24255), .B(n24256), .Z(n24164) );
  AND U25073 ( .A(n538), .B(n24257), .Z(n24255) );
  XOR U25074 ( .A(n24258), .B(n24256), .Z(n24257) );
  XNOR U25075 ( .A(n24259), .B(n24260), .Z(n24247) );
  AND U25076 ( .A(n24261), .B(n24262), .Z(n24259) );
  XNOR U25077 ( .A(n24260), .B(n24189), .Z(n24262) );
  XOR U25078 ( .A(n24253), .B(n24254), .Z(n24189) );
  XNOR U25079 ( .A(n24263), .B(n24264), .Z(n24254) );
  ANDN U25080 ( .B(n24265), .A(n24266), .Z(n24263) );
  XOR U25081 ( .A(n24267), .B(n24268), .Z(n24265) );
  XOR U25082 ( .A(n24269), .B(n24270), .Z(n24253) );
  XNOR U25083 ( .A(n24271), .B(n24272), .Z(n24270) );
  ANDN U25084 ( .B(n24273), .A(n24274), .Z(n24271) );
  XNOR U25085 ( .A(n24275), .B(n24276), .Z(n24273) );
  IV U25086 ( .A(n24251), .Z(n24269) );
  XOR U25087 ( .A(n24277), .B(n24278), .Z(n24251) );
  ANDN U25088 ( .B(n24279), .A(n24280), .Z(n24277) );
  XOR U25089 ( .A(n24278), .B(n24281), .Z(n24279) );
  XOR U25090 ( .A(n24260), .B(n24191), .Z(n24261) );
  XOR U25091 ( .A(n24282), .B(n24283), .Z(n24191) );
  AND U25092 ( .A(n538), .B(n24284), .Z(n24282) );
  XOR U25093 ( .A(n24285), .B(n24283), .Z(n24284) );
  XNOR U25094 ( .A(n24286), .B(n24287), .Z(n24260) );
  NAND U25095 ( .A(n24288), .B(n24289), .Z(n24287) );
  XOR U25096 ( .A(n24290), .B(n24239), .Z(n24289) );
  XOR U25097 ( .A(n24280), .B(n24281), .Z(n24239) );
  XOR U25098 ( .A(n24291), .B(n24268), .Z(n24281) );
  XOR U25099 ( .A(n24292), .B(n24293), .Z(n24268) );
  ANDN U25100 ( .B(n24294), .A(n24295), .Z(n24292) );
  XOR U25101 ( .A(n24293), .B(n24296), .Z(n24294) );
  IV U25102 ( .A(n24266), .Z(n24291) );
  XOR U25103 ( .A(n24264), .B(n24297), .Z(n24266) );
  XOR U25104 ( .A(n24298), .B(n24299), .Z(n24297) );
  ANDN U25105 ( .B(n24300), .A(n24301), .Z(n24298) );
  XOR U25106 ( .A(n24302), .B(n24299), .Z(n24300) );
  IV U25107 ( .A(n24267), .Z(n24264) );
  XOR U25108 ( .A(n24303), .B(n24304), .Z(n24267) );
  ANDN U25109 ( .B(n24305), .A(n24306), .Z(n24303) );
  XOR U25110 ( .A(n24304), .B(n24307), .Z(n24305) );
  XOR U25111 ( .A(n24308), .B(n24309), .Z(n24280) );
  XNOR U25112 ( .A(n24275), .B(n24310), .Z(n24309) );
  IV U25113 ( .A(n24278), .Z(n24310) );
  XOR U25114 ( .A(n24311), .B(n24312), .Z(n24278) );
  ANDN U25115 ( .B(n24313), .A(n24314), .Z(n24311) );
  XOR U25116 ( .A(n24312), .B(n24315), .Z(n24313) );
  XNOR U25117 ( .A(n24316), .B(n24317), .Z(n24275) );
  ANDN U25118 ( .B(n24318), .A(n24319), .Z(n24316) );
  XOR U25119 ( .A(n24317), .B(n24320), .Z(n24318) );
  IV U25120 ( .A(n24274), .Z(n24308) );
  XOR U25121 ( .A(n24272), .B(n24321), .Z(n24274) );
  XOR U25122 ( .A(n24322), .B(n24323), .Z(n24321) );
  ANDN U25123 ( .B(n24324), .A(n24325), .Z(n24322) );
  XOR U25124 ( .A(n24326), .B(n24323), .Z(n24324) );
  IV U25125 ( .A(n24276), .Z(n24272) );
  XOR U25126 ( .A(n24327), .B(n24328), .Z(n24276) );
  ANDN U25127 ( .B(n24329), .A(n24330), .Z(n24327) );
  XOR U25128 ( .A(n24331), .B(n24328), .Z(n24329) );
  IV U25129 ( .A(n24286), .Z(n24290) );
  XOR U25130 ( .A(n24286), .B(n24241), .Z(n24288) );
  XOR U25131 ( .A(n24332), .B(n24333), .Z(n24241) );
  AND U25132 ( .A(n538), .B(n24334), .Z(n24332) );
  XOR U25133 ( .A(n24335), .B(n24333), .Z(n24334) );
  NANDN U25134 ( .A(n24243), .B(n24245), .Z(n24286) );
  XOR U25135 ( .A(n24336), .B(n24337), .Z(n24245) );
  AND U25136 ( .A(n538), .B(n24338), .Z(n24336) );
  XOR U25137 ( .A(n24337), .B(n24339), .Z(n24338) );
  XNOR U25138 ( .A(n24340), .B(n24341), .Z(n538) );
  AND U25139 ( .A(n24342), .B(n24343), .Z(n24340) );
  XOR U25140 ( .A(n24341), .B(n24256), .Z(n24343) );
  XNOR U25141 ( .A(n24344), .B(n24345), .Z(n24256) );
  ANDN U25142 ( .B(n24346), .A(n24347), .Z(n24344) );
  XOR U25143 ( .A(n24345), .B(n24348), .Z(n24346) );
  XNOR U25144 ( .A(n24341), .B(n24258), .Z(n24342) );
  XOR U25145 ( .A(n24349), .B(n24350), .Z(n24258) );
  AND U25146 ( .A(n542), .B(n24351), .Z(n24349) );
  XOR U25147 ( .A(n24352), .B(n24350), .Z(n24351) );
  XNOR U25148 ( .A(n24353), .B(n24354), .Z(n24341) );
  AND U25149 ( .A(n24355), .B(n24356), .Z(n24353) );
  XNOR U25150 ( .A(n24354), .B(n24283), .Z(n24356) );
  XOR U25151 ( .A(n24347), .B(n24348), .Z(n24283) );
  XNOR U25152 ( .A(n24357), .B(n24358), .Z(n24348) );
  ANDN U25153 ( .B(n24359), .A(n24360), .Z(n24357) );
  XOR U25154 ( .A(n24361), .B(n24362), .Z(n24359) );
  XOR U25155 ( .A(n24363), .B(n24364), .Z(n24347) );
  XNOR U25156 ( .A(n24365), .B(n24366), .Z(n24364) );
  ANDN U25157 ( .B(n24367), .A(n24368), .Z(n24365) );
  XNOR U25158 ( .A(n24369), .B(n24370), .Z(n24367) );
  IV U25159 ( .A(n24345), .Z(n24363) );
  XOR U25160 ( .A(n24371), .B(n24372), .Z(n24345) );
  ANDN U25161 ( .B(n24373), .A(n24374), .Z(n24371) );
  XOR U25162 ( .A(n24372), .B(n24375), .Z(n24373) );
  XOR U25163 ( .A(n24354), .B(n24285), .Z(n24355) );
  XOR U25164 ( .A(n24376), .B(n24377), .Z(n24285) );
  AND U25165 ( .A(n542), .B(n24378), .Z(n24376) );
  XOR U25166 ( .A(n24379), .B(n24377), .Z(n24378) );
  XNOR U25167 ( .A(n24380), .B(n24381), .Z(n24354) );
  NAND U25168 ( .A(n24382), .B(n24383), .Z(n24381) );
  XOR U25169 ( .A(n24384), .B(n24333), .Z(n24383) );
  XOR U25170 ( .A(n24374), .B(n24375), .Z(n24333) );
  XOR U25171 ( .A(n24385), .B(n24362), .Z(n24375) );
  XOR U25172 ( .A(n24386), .B(n24387), .Z(n24362) );
  ANDN U25173 ( .B(n24388), .A(n24389), .Z(n24386) );
  XOR U25174 ( .A(n24387), .B(n24390), .Z(n24388) );
  IV U25175 ( .A(n24360), .Z(n24385) );
  XOR U25176 ( .A(n24358), .B(n24391), .Z(n24360) );
  XOR U25177 ( .A(n24392), .B(n24393), .Z(n24391) );
  ANDN U25178 ( .B(n24394), .A(n24395), .Z(n24392) );
  XOR U25179 ( .A(n24396), .B(n24393), .Z(n24394) );
  IV U25180 ( .A(n24361), .Z(n24358) );
  XOR U25181 ( .A(n24397), .B(n24398), .Z(n24361) );
  ANDN U25182 ( .B(n24399), .A(n24400), .Z(n24397) );
  XOR U25183 ( .A(n24398), .B(n24401), .Z(n24399) );
  XOR U25184 ( .A(n24402), .B(n24403), .Z(n24374) );
  XNOR U25185 ( .A(n24369), .B(n24404), .Z(n24403) );
  IV U25186 ( .A(n24372), .Z(n24404) );
  XOR U25187 ( .A(n24405), .B(n24406), .Z(n24372) );
  ANDN U25188 ( .B(n24407), .A(n24408), .Z(n24405) );
  XOR U25189 ( .A(n24406), .B(n24409), .Z(n24407) );
  XNOR U25190 ( .A(n24410), .B(n24411), .Z(n24369) );
  ANDN U25191 ( .B(n24412), .A(n24413), .Z(n24410) );
  XOR U25192 ( .A(n24411), .B(n24414), .Z(n24412) );
  IV U25193 ( .A(n24368), .Z(n24402) );
  XOR U25194 ( .A(n24366), .B(n24415), .Z(n24368) );
  XOR U25195 ( .A(n24416), .B(n24417), .Z(n24415) );
  ANDN U25196 ( .B(n24418), .A(n24419), .Z(n24416) );
  XOR U25197 ( .A(n24420), .B(n24417), .Z(n24418) );
  IV U25198 ( .A(n24370), .Z(n24366) );
  XOR U25199 ( .A(n24421), .B(n24422), .Z(n24370) );
  ANDN U25200 ( .B(n24423), .A(n24424), .Z(n24421) );
  XOR U25201 ( .A(n24425), .B(n24422), .Z(n24423) );
  IV U25202 ( .A(n24380), .Z(n24384) );
  XOR U25203 ( .A(n24380), .B(n24335), .Z(n24382) );
  XOR U25204 ( .A(n24426), .B(n24427), .Z(n24335) );
  AND U25205 ( .A(n542), .B(n24428), .Z(n24426) );
  XOR U25206 ( .A(n24429), .B(n24427), .Z(n24428) );
  NANDN U25207 ( .A(n24337), .B(n24339), .Z(n24380) );
  XOR U25208 ( .A(n24430), .B(n24431), .Z(n24339) );
  AND U25209 ( .A(n542), .B(n24432), .Z(n24430) );
  XOR U25210 ( .A(n24431), .B(n24433), .Z(n24432) );
  XNOR U25211 ( .A(n24434), .B(n24435), .Z(n542) );
  AND U25212 ( .A(n24436), .B(n24437), .Z(n24434) );
  XOR U25213 ( .A(n24435), .B(n24350), .Z(n24437) );
  XNOR U25214 ( .A(n24438), .B(n24439), .Z(n24350) );
  ANDN U25215 ( .B(n24440), .A(n24441), .Z(n24438) );
  XOR U25216 ( .A(n24439), .B(n24442), .Z(n24440) );
  XNOR U25217 ( .A(n24435), .B(n24352), .Z(n24436) );
  XOR U25218 ( .A(n24443), .B(n24444), .Z(n24352) );
  AND U25219 ( .A(n546), .B(n24445), .Z(n24443) );
  XOR U25220 ( .A(n24446), .B(n24444), .Z(n24445) );
  XNOR U25221 ( .A(n24447), .B(n24448), .Z(n24435) );
  AND U25222 ( .A(n24449), .B(n24450), .Z(n24447) );
  XNOR U25223 ( .A(n24448), .B(n24377), .Z(n24450) );
  XOR U25224 ( .A(n24441), .B(n24442), .Z(n24377) );
  XNOR U25225 ( .A(n24451), .B(n24452), .Z(n24442) );
  ANDN U25226 ( .B(n24453), .A(n24454), .Z(n24451) );
  XOR U25227 ( .A(n24455), .B(n24456), .Z(n24453) );
  XOR U25228 ( .A(n24457), .B(n24458), .Z(n24441) );
  XNOR U25229 ( .A(n24459), .B(n24460), .Z(n24458) );
  ANDN U25230 ( .B(n24461), .A(n24462), .Z(n24459) );
  XNOR U25231 ( .A(n24463), .B(n24464), .Z(n24461) );
  IV U25232 ( .A(n24439), .Z(n24457) );
  XOR U25233 ( .A(n24465), .B(n24466), .Z(n24439) );
  ANDN U25234 ( .B(n24467), .A(n24468), .Z(n24465) );
  XOR U25235 ( .A(n24466), .B(n24469), .Z(n24467) );
  XOR U25236 ( .A(n24448), .B(n24379), .Z(n24449) );
  XOR U25237 ( .A(n24470), .B(n24471), .Z(n24379) );
  AND U25238 ( .A(n546), .B(n24472), .Z(n24470) );
  XOR U25239 ( .A(n24473), .B(n24471), .Z(n24472) );
  XNOR U25240 ( .A(n24474), .B(n24475), .Z(n24448) );
  NAND U25241 ( .A(n24476), .B(n24477), .Z(n24475) );
  XOR U25242 ( .A(n24478), .B(n24427), .Z(n24477) );
  XOR U25243 ( .A(n24468), .B(n24469), .Z(n24427) );
  XOR U25244 ( .A(n24479), .B(n24456), .Z(n24469) );
  XOR U25245 ( .A(n24480), .B(n24481), .Z(n24456) );
  ANDN U25246 ( .B(n24482), .A(n24483), .Z(n24480) );
  XOR U25247 ( .A(n24481), .B(n24484), .Z(n24482) );
  IV U25248 ( .A(n24454), .Z(n24479) );
  XOR U25249 ( .A(n24452), .B(n24485), .Z(n24454) );
  XOR U25250 ( .A(n24486), .B(n24487), .Z(n24485) );
  ANDN U25251 ( .B(n24488), .A(n24489), .Z(n24486) );
  XOR U25252 ( .A(n24490), .B(n24487), .Z(n24488) );
  IV U25253 ( .A(n24455), .Z(n24452) );
  XOR U25254 ( .A(n24491), .B(n24492), .Z(n24455) );
  ANDN U25255 ( .B(n24493), .A(n24494), .Z(n24491) );
  XOR U25256 ( .A(n24492), .B(n24495), .Z(n24493) );
  XOR U25257 ( .A(n24496), .B(n24497), .Z(n24468) );
  XNOR U25258 ( .A(n24463), .B(n24498), .Z(n24497) );
  IV U25259 ( .A(n24466), .Z(n24498) );
  XOR U25260 ( .A(n24499), .B(n24500), .Z(n24466) );
  ANDN U25261 ( .B(n24501), .A(n24502), .Z(n24499) );
  XOR U25262 ( .A(n24500), .B(n24503), .Z(n24501) );
  XNOR U25263 ( .A(n24504), .B(n24505), .Z(n24463) );
  ANDN U25264 ( .B(n24506), .A(n24507), .Z(n24504) );
  XOR U25265 ( .A(n24505), .B(n24508), .Z(n24506) );
  IV U25266 ( .A(n24462), .Z(n24496) );
  XOR U25267 ( .A(n24460), .B(n24509), .Z(n24462) );
  XOR U25268 ( .A(n24510), .B(n24511), .Z(n24509) );
  ANDN U25269 ( .B(n24512), .A(n24513), .Z(n24510) );
  XOR U25270 ( .A(n24514), .B(n24511), .Z(n24512) );
  IV U25271 ( .A(n24464), .Z(n24460) );
  XOR U25272 ( .A(n24515), .B(n24516), .Z(n24464) );
  ANDN U25273 ( .B(n24517), .A(n24518), .Z(n24515) );
  XOR U25274 ( .A(n24519), .B(n24516), .Z(n24517) );
  IV U25275 ( .A(n24474), .Z(n24478) );
  XOR U25276 ( .A(n24474), .B(n24429), .Z(n24476) );
  XOR U25277 ( .A(n24520), .B(n24521), .Z(n24429) );
  AND U25278 ( .A(n546), .B(n24522), .Z(n24520) );
  XOR U25279 ( .A(n24523), .B(n24521), .Z(n24522) );
  NANDN U25280 ( .A(n24431), .B(n24433), .Z(n24474) );
  XOR U25281 ( .A(n24524), .B(n24525), .Z(n24433) );
  AND U25282 ( .A(n546), .B(n24526), .Z(n24524) );
  XOR U25283 ( .A(n24525), .B(n24527), .Z(n24526) );
  XNOR U25284 ( .A(n24528), .B(n24529), .Z(n546) );
  AND U25285 ( .A(n24530), .B(n24531), .Z(n24528) );
  XOR U25286 ( .A(n24529), .B(n24444), .Z(n24531) );
  XNOR U25287 ( .A(n24532), .B(n24533), .Z(n24444) );
  ANDN U25288 ( .B(n24534), .A(n24535), .Z(n24532) );
  XOR U25289 ( .A(n24533), .B(n24536), .Z(n24534) );
  XNOR U25290 ( .A(n24529), .B(n24446), .Z(n24530) );
  XOR U25291 ( .A(n24537), .B(n24538), .Z(n24446) );
  AND U25292 ( .A(n550), .B(n24539), .Z(n24537) );
  XOR U25293 ( .A(n24540), .B(n24538), .Z(n24539) );
  XNOR U25294 ( .A(n24541), .B(n24542), .Z(n24529) );
  AND U25295 ( .A(n24543), .B(n24544), .Z(n24541) );
  XNOR U25296 ( .A(n24542), .B(n24471), .Z(n24544) );
  XOR U25297 ( .A(n24535), .B(n24536), .Z(n24471) );
  XNOR U25298 ( .A(n24545), .B(n24546), .Z(n24536) );
  ANDN U25299 ( .B(n24547), .A(n24548), .Z(n24545) );
  XOR U25300 ( .A(n24549), .B(n24550), .Z(n24547) );
  XOR U25301 ( .A(n24551), .B(n24552), .Z(n24535) );
  XNOR U25302 ( .A(n24553), .B(n24554), .Z(n24552) );
  ANDN U25303 ( .B(n24555), .A(n24556), .Z(n24553) );
  XNOR U25304 ( .A(n24557), .B(n24558), .Z(n24555) );
  IV U25305 ( .A(n24533), .Z(n24551) );
  XOR U25306 ( .A(n24559), .B(n24560), .Z(n24533) );
  ANDN U25307 ( .B(n24561), .A(n24562), .Z(n24559) );
  XOR U25308 ( .A(n24560), .B(n24563), .Z(n24561) );
  XOR U25309 ( .A(n24542), .B(n24473), .Z(n24543) );
  XOR U25310 ( .A(n24564), .B(n24565), .Z(n24473) );
  AND U25311 ( .A(n550), .B(n24566), .Z(n24564) );
  XOR U25312 ( .A(n24567), .B(n24565), .Z(n24566) );
  XNOR U25313 ( .A(n24568), .B(n24569), .Z(n24542) );
  NAND U25314 ( .A(n24570), .B(n24571), .Z(n24569) );
  XOR U25315 ( .A(n24572), .B(n24521), .Z(n24571) );
  XOR U25316 ( .A(n24562), .B(n24563), .Z(n24521) );
  XOR U25317 ( .A(n24573), .B(n24550), .Z(n24563) );
  XOR U25318 ( .A(n24574), .B(n24575), .Z(n24550) );
  ANDN U25319 ( .B(n24576), .A(n24577), .Z(n24574) );
  XOR U25320 ( .A(n24575), .B(n24578), .Z(n24576) );
  IV U25321 ( .A(n24548), .Z(n24573) );
  XOR U25322 ( .A(n24546), .B(n24579), .Z(n24548) );
  XOR U25323 ( .A(n24580), .B(n24581), .Z(n24579) );
  ANDN U25324 ( .B(n24582), .A(n24583), .Z(n24580) );
  XOR U25325 ( .A(n24584), .B(n24581), .Z(n24582) );
  IV U25326 ( .A(n24549), .Z(n24546) );
  XOR U25327 ( .A(n24585), .B(n24586), .Z(n24549) );
  ANDN U25328 ( .B(n24587), .A(n24588), .Z(n24585) );
  XOR U25329 ( .A(n24586), .B(n24589), .Z(n24587) );
  XOR U25330 ( .A(n24590), .B(n24591), .Z(n24562) );
  XNOR U25331 ( .A(n24557), .B(n24592), .Z(n24591) );
  IV U25332 ( .A(n24560), .Z(n24592) );
  XOR U25333 ( .A(n24593), .B(n24594), .Z(n24560) );
  ANDN U25334 ( .B(n24595), .A(n24596), .Z(n24593) );
  XOR U25335 ( .A(n24594), .B(n24597), .Z(n24595) );
  XNOR U25336 ( .A(n24598), .B(n24599), .Z(n24557) );
  ANDN U25337 ( .B(n24600), .A(n24601), .Z(n24598) );
  XOR U25338 ( .A(n24599), .B(n24602), .Z(n24600) );
  IV U25339 ( .A(n24556), .Z(n24590) );
  XOR U25340 ( .A(n24554), .B(n24603), .Z(n24556) );
  XOR U25341 ( .A(n24604), .B(n24605), .Z(n24603) );
  ANDN U25342 ( .B(n24606), .A(n24607), .Z(n24604) );
  XOR U25343 ( .A(n24608), .B(n24605), .Z(n24606) );
  IV U25344 ( .A(n24558), .Z(n24554) );
  XOR U25345 ( .A(n24609), .B(n24610), .Z(n24558) );
  ANDN U25346 ( .B(n24611), .A(n24612), .Z(n24609) );
  XOR U25347 ( .A(n24613), .B(n24610), .Z(n24611) );
  IV U25348 ( .A(n24568), .Z(n24572) );
  XOR U25349 ( .A(n24568), .B(n24523), .Z(n24570) );
  XOR U25350 ( .A(n24614), .B(n24615), .Z(n24523) );
  AND U25351 ( .A(n550), .B(n24616), .Z(n24614) );
  XOR U25352 ( .A(n24617), .B(n24615), .Z(n24616) );
  NANDN U25353 ( .A(n24525), .B(n24527), .Z(n24568) );
  XOR U25354 ( .A(n24618), .B(n24619), .Z(n24527) );
  AND U25355 ( .A(n550), .B(n24620), .Z(n24618) );
  XOR U25356 ( .A(n24619), .B(n24621), .Z(n24620) );
  XNOR U25357 ( .A(n24622), .B(n24623), .Z(n550) );
  AND U25358 ( .A(n24624), .B(n24625), .Z(n24622) );
  XOR U25359 ( .A(n24623), .B(n24538), .Z(n24625) );
  XNOR U25360 ( .A(n24626), .B(n24627), .Z(n24538) );
  ANDN U25361 ( .B(n24628), .A(n24629), .Z(n24626) );
  XOR U25362 ( .A(n24627), .B(n24630), .Z(n24628) );
  XNOR U25363 ( .A(n24623), .B(n24540), .Z(n24624) );
  XOR U25364 ( .A(n24631), .B(n24632), .Z(n24540) );
  AND U25365 ( .A(n554), .B(n24633), .Z(n24631) );
  XOR U25366 ( .A(n24634), .B(n24632), .Z(n24633) );
  XNOR U25367 ( .A(n24635), .B(n24636), .Z(n24623) );
  AND U25368 ( .A(n24637), .B(n24638), .Z(n24635) );
  XNOR U25369 ( .A(n24636), .B(n24565), .Z(n24638) );
  XOR U25370 ( .A(n24629), .B(n24630), .Z(n24565) );
  XNOR U25371 ( .A(n24639), .B(n24640), .Z(n24630) );
  ANDN U25372 ( .B(n24641), .A(n24642), .Z(n24639) );
  XOR U25373 ( .A(n24643), .B(n24644), .Z(n24641) );
  XOR U25374 ( .A(n24645), .B(n24646), .Z(n24629) );
  XNOR U25375 ( .A(n24647), .B(n24648), .Z(n24646) );
  ANDN U25376 ( .B(n24649), .A(n24650), .Z(n24647) );
  XNOR U25377 ( .A(n24651), .B(n24652), .Z(n24649) );
  IV U25378 ( .A(n24627), .Z(n24645) );
  XOR U25379 ( .A(n24653), .B(n24654), .Z(n24627) );
  ANDN U25380 ( .B(n24655), .A(n24656), .Z(n24653) );
  XOR U25381 ( .A(n24654), .B(n24657), .Z(n24655) );
  XOR U25382 ( .A(n24636), .B(n24567), .Z(n24637) );
  XOR U25383 ( .A(n24658), .B(n24659), .Z(n24567) );
  AND U25384 ( .A(n554), .B(n24660), .Z(n24658) );
  XOR U25385 ( .A(n24661), .B(n24659), .Z(n24660) );
  XNOR U25386 ( .A(n24662), .B(n24663), .Z(n24636) );
  NAND U25387 ( .A(n24664), .B(n24665), .Z(n24663) );
  XOR U25388 ( .A(n24666), .B(n24615), .Z(n24665) );
  XOR U25389 ( .A(n24656), .B(n24657), .Z(n24615) );
  XOR U25390 ( .A(n24667), .B(n24644), .Z(n24657) );
  XOR U25391 ( .A(n24668), .B(n24669), .Z(n24644) );
  ANDN U25392 ( .B(n24670), .A(n24671), .Z(n24668) );
  XOR U25393 ( .A(n24669), .B(n24672), .Z(n24670) );
  IV U25394 ( .A(n24642), .Z(n24667) );
  XOR U25395 ( .A(n24640), .B(n24673), .Z(n24642) );
  XOR U25396 ( .A(n24674), .B(n24675), .Z(n24673) );
  ANDN U25397 ( .B(n24676), .A(n24677), .Z(n24674) );
  XOR U25398 ( .A(n24678), .B(n24675), .Z(n24676) );
  IV U25399 ( .A(n24643), .Z(n24640) );
  XOR U25400 ( .A(n24679), .B(n24680), .Z(n24643) );
  ANDN U25401 ( .B(n24681), .A(n24682), .Z(n24679) );
  XOR U25402 ( .A(n24680), .B(n24683), .Z(n24681) );
  XOR U25403 ( .A(n24684), .B(n24685), .Z(n24656) );
  XNOR U25404 ( .A(n24651), .B(n24686), .Z(n24685) );
  IV U25405 ( .A(n24654), .Z(n24686) );
  XOR U25406 ( .A(n24687), .B(n24688), .Z(n24654) );
  ANDN U25407 ( .B(n24689), .A(n24690), .Z(n24687) );
  XOR U25408 ( .A(n24688), .B(n24691), .Z(n24689) );
  XNOR U25409 ( .A(n24692), .B(n24693), .Z(n24651) );
  ANDN U25410 ( .B(n24694), .A(n24695), .Z(n24692) );
  XOR U25411 ( .A(n24693), .B(n24696), .Z(n24694) );
  IV U25412 ( .A(n24650), .Z(n24684) );
  XOR U25413 ( .A(n24648), .B(n24697), .Z(n24650) );
  XOR U25414 ( .A(n24698), .B(n24699), .Z(n24697) );
  ANDN U25415 ( .B(n24700), .A(n24701), .Z(n24698) );
  XOR U25416 ( .A(n24702), .B(n24699), .Z(n24700) );
  IV U25417 ( .A(n24652), .Z(n24648) );
  XOR U25418 ( .A(n24703), .B(n24704), .Z(n24652) );
  ANDN U25419 ( .B(n24705), .A(n24706), .Z(n24703) );
  XOR U25420 ( .A(n24707), .B(n24704), .Z(n24705) );
  IV U25421 ( .A(n24662), .Z(n24666) );
  XOR U25422 ( .A(n24662), .B(n24617), .Z(n24664) );
  XOR U25423 ( .A(n24708), .B(n24709), .Z(n24617) );
  AND U25424 ( .A(n554), .B(n24710), .Z(n24708) );
  XOR U25425 ( .A(n24711), .B(n24709), .Z(n24710) );
  NANDN U25426 ( .A(n24619), .B(n24621), .Z(n24662) );
  XOR U25427 ( .A(n24712), .B(n24713), .Z(n24621) );
  AND U25428 ( .A(n554), .B(n24714), .Z(n24712) );
  XOR U25429 ( .A(n24713), .B(n24715), .Z(n24714) );
  XNOR U25430 ( .A(n24716), .B(n24717), .Z(n554) );
  AND U25431 ( .A(n24718), .B(n24719), .Z(n24716) );
  XOR U25432 ( .A(n24717), .B(n24632), .Z(n24719) );
  XNOR U25433 ( .A(n24720), .B(n24721), .Z(n24632) );
  ANDN U25434 ( .B(n24722), .A(n24723), .Z(n24720) );
  XOR U25435 ( .A(n24721), .B(n24724), .Z(n24722) );
  XNOR U25436 ( .A(n24717), .B(n24634), .Z(n24718) );
  XOR U25437 ( .A(n24725), .B(n24726), .Z(n24634) );
  AND U25438 ( .A(n558), .B(n24727), .Z(n24725) );
  XOR U25439 ( .A(n24728), .B(n24726), .Z(n24727) );
  XNOR U25440 ( .A(n24729), .B(n24730), .Z(n24717) );
  AND U25441 ( .A(n24731), .B(n24732), .Z(n24729) );
  XNOR U25442 ( .A(n24730), .B(n24659), .Z(n24732) );
  XOR U25443 ( .A(n24723), .B(n24724), .Z(n24659) );
  XNOR U25444 ( .A(n24733), .B(n24734), .Z(n24724) );
  ANDN U25445 ( .B(n24735), .A(n24736), .Z(n24733) );
  XOR U25446 ( .A(n24737), .B(n24738), .Z(n24735) );
  XOR U25447 ( .A(n24739), .B(n24740), .Z(n24723) );
  XNOR U25448 ( .A(n24741), .B(n24742), .Z(n24740) );
  ANDN U25449 ( .B(n24743), .A(n24744), .Z(n24741) );
  XNOR U25450 ( .A(n24745), .B(n24746), .Z(n24743) );
  IV U25451 ( .A(n24721), .Z(n24739) );
  XOR U25452 ( .A(n24747), .B(n24748), .Z(n24721) );
  ANDN U25453 ( .B(n24749), .A(n24750), .Z(n24747) );
  XOR U25454 ( .A(n24748), .B(n24751), .Z(n24749) );
  XOR U25455 ( .A(n24730), .B(n24661), .Z(n24731) );
  XOR U25456 ( .A(n24752), .B(n24753), .Z(n24661) );
  AND U25457 ( .A(n558), .B(n24754), .Z(n24752) );
  XOR U25458 ( .A(n24755), .B(n24753), .Z(n24754) );
  XNOR U25459 ( .A(n24756), .B(n24757), .Z(n24730) );
  NAND U25460 ( .A(n24758), .B(n24759), .Z(n24757) );
  XOR U25461 ( .A(n24760), .B(n24709), .Z(n24759) );
  XOR U25462 ( .A(n24750), .B(n24751), .Z(n24709) );
  XOR U25463 ( .A(n24761), .B(n24738), .Z(n24751) );
  XOR U25464 ( .A(n24762), .B(n24763), .Z(n24738) );
  ANDN U25465 ( .B(n24764), .A(n24765), .Z(n24762) );
  XOR U25466 ( .A(n24763), .B(n24766), .Z(n24764) );
  IV U25467 ( .A(n24736), .Z(n24761) );
  XOR U25468 ( .A(n24734), .B(n24767), .Z(n24736) );
  XOR U25469 ( .A(n24768), .B(n24769), .Z(n24767) );
  ANDN U25470 ( .B(n24770), .A(n24771), .Z(n24768) );
  XOR U25471 ( .A(n24772), .B(n24769), .Z(n24770) );
  IV U25472 ( .A(n24737), .Z(n24734) );
  XOR U25473 ( .A(n24773), .B(n24774), .Z(n24737) );
  ANDN U25474 ( .B(n24775), .A(n24776), .Z(n24773) );
  XOR U25475 ( .A(n24774), .B(n24777), .Z(n24775) );
  XOR U25476 ( .A(n24778), .B(n24779), .Z(n24750) );
  XNOR U25477 ( .A(n24745), .B(n24780), .Z(n24779) );
  IV U25478 ( .A(n24748), .Z(n24780) );
  XOR U25479 ( .A(n24781), .B(n24782), .Z(n24748) );
  ANDN U25480 ( .B(n24783), .A(n24784), .Z(n24781) );
  XOR U25481 ( .A(n24782), .B(n24785), .Z(n24783) );
  XNOR U25482 ( .A(n24786), .B(n24787), .Z(n24745) );
  ANDN U25483 ( .B(n24788), .A(n24789), .Z(n24786) );
  XOR U25484 ( .A(n24787), .B(n24790), .Z(n24788) );
  IV U25485 ( .A(n24744), .Z(n24778) );
  XOR U25486 ( .A(n24742), .B(n24791), .Z(n24744) );
  XOR U25487 ( .A(n24792), .B(n24793), .Z(n24791) );
  ANDN U25488 ( .B(n24794), .A(n24795), .Z(n24792) );
  XOR U25489 ( .A(n24796), .B(n24793), .Z(n24794) );
  IV U25490 ( .A(n24746), .Z(n24742) );
  XOR U25491 ( .A(n24797), .B(n24798), .Z(n24746) );
  ANDN U25492 ( .B(n24799), .A(n24800), .Z(n24797) );
  XOR U25493 ( .A(n24801), .B(n24798), .Z(n24799) );
  IV U25494 ( .A(n24756), .Z(n24760) );
  XOR U25495 ( .A(n24756), .B(n24711), .Z(n24758) );
  XOR U25496 ( .A(n24802), .B(n24803), .Z(n24711) );
  AND U25497 ( .A(n558), .B(n24804), .Z(n24802) );
  XOR U25498 ( .A(n24805), .B(n24803), .Z(n24804) );
  NANDN U25499 ( .A(n24713), .B(n24715), .Z(n24756) );
  XOR U25500 ( .A(n24806), .B(n24807), .Z(n24715) );
  AND U25501 ( .A(n558), .B(n24808), .Z(n24806) );
  XOR U25502 ( .A(n24807), .B(n24809), .Z(n24808) );
  XNOR U25503 ( .A(n24810), .B(n24811), .Z(n558) );
  AND U25504 ( .A(n24812), .B(n24813), .Z(n24810) );
  XOR U25505 ( .A(n24811), .B(n24726), .Z(n24813) );
  XNOR U25506 ( .A(n24814), .B(n24815), .Z(n24726) );
  ANDN U25507 ( .B(n24816), .A(n24817), .Z(n24814) );
  XOR U25508 ( .A(n24815), .B(n24818), .Z(n24816) );
  XNOR U25509 ( .A(n24811), .B(n24728), .Z(n24812) );
  XOR U25510 ( .A(n24819), .B(n24820), .Z(n24728) );
  AND U25511 ( .A(n562), .B(n24821), .Z(n24819) );
  XOR U25512 ( .A(n24822), .B(n24820), .Z(n24821) );
  XNOR U25513 ( .A(n24823), .B(n24824), .Z(n24811) );
  AND U25514 ( .A(n24825), .B(n24826), .Z(n24823) );
  XNOR U25515 ( .A(n24824), .B(n24753), .Z(n24826) );
  XOR U25516 ( .A(n24817), .B(n24818), .Z(n24753) );
  XNOR U25517 ( .A(n24827), .B(n24828), .Z(n24818) );
  ANDN U25518 ( .B(n24829), .A(n24830), .Z(n24827) );
  XOR U25519 ( .A(n24831), .B(n24832), .Z(n24829) );
  XOR U25520 ( .A(n24833), .B(n24834), .Z(n24817) );
  XNOR U25521 ( .A(n24835), .B(n24836), .Z(n24834) );
  ANDN U25522 ( .B(n24837), .A(n24838), .Z(n24835) );
  XNOR U25523 ( .A(n24839), .B(n24840), .Z(n24837) );
  IV U25524 ( .A(n24815), .Z(n24833) );
  XOR U25525 ( .A(n24841), .B(n24842), .Z(n24815) );
  ANDN U25526 ( .B(n24843), .A(n24844), .Z(n24841) );
  XOR U25527 ( .A(n24842), .B(n24845), .Z(n24843) );
  XOR U25528 ( .A(n24824), .B(n24755), .Z(n24825) );
  XOR U25529 ( .A(n24846), .B(n24847), .Z(n24755) );
  AND U25530 ( .A(n562), .B(n24848), .Z(n24846) );
  XOR U25531 ( .A(n24849), .B(n24847), .Z(n24848) );
  XNOR U25532 ( .A(n24850), .B(n24851), .Z(n24824) );
  NAND U25533 ( .A(n24852), .B(n24853), .Z(n24851) );
  XOR U25534 ( .A(n24854), .B(n24803), .Z(n24853) );
  XOR U25535 ( .A(n24844), .B(n24845), .Z(n24803) );
  XOR U25536 ( .A(n24855), .B(n24832), .Z(n24845) );
  XOR U25537 ( .A(n24856), .B(n24857), .Z(n24832) );
  ANDN U25538 ( .B(n24858), .A(n24859), .Z(n24856) );
  XOR U25539 ( .A(n24857), .B(n24860), .Z(n24858) );
  IV U25540 ( .A(n24830), .Z(n24855) );
  XOR U25541 ( .A(n24828), .B(n24861), .Z(n24830) );
  XOR U25542 ( .A(n24862), .B(n24863), .Z(n24861) );
  ANDN U25543 ( .B(n24864), .A(n24865), .Z(n24862) );
  XOR U25544 ( .A(n24866), .B(n24863), .Z(n24864) );
  IV U25545 ( .A(n24831), .Z(n24828) );
  XOR U25546 ( .A(n24867), .B(n24868), .Z(n24831) );
  ANDN U25547 ( .B(n24869), .A(n24870), .Z(n24867) );
  XOR U25548 ( .A(n24868), .B(n24871), .Z(n24869) );
  XOR U25549 ( .A(n24872), .B(n24873), .Z(n24844) );
  XNOR U25550 ( .A(n24839), .B(n24874), .Z(n24873) );
  IV U25551 ( .A(n24842), .Z(n24874) );
  XOR U25552 ( .A(n24875), .B(n24876), .Z(n24842) );
  ANDN U25553 ( .B(n24877), .A(n24878), .Z(n24875) );
  XOR U25554 ( .A(n24876), .B(n24879), .Z(n24877) );
  XNOR U25555 ( .A(n24880), .B(n24881), .Z(n24839) );
  ANDN U25556 ( .B(n24882), .A(n24883), .Z(n24880) );
  XOR U25557 ( .A(n24881), .B(n24884), .Z(n24882) );
  IV U25558 ( .A(n24838), .Z(n24872) );
  XOR U25559 ( .A(n24836), .B(n24885), .Z(n24838) );
  XOR U25560 ( .A(n24886), .B(n24887), .Z(n24885) );
  ANDN U25561 ( .B(n24888), .A(n24889), .Z(n24886) );
  XOR U25562 ( .A(n24890), .B(n24887), .Z(n24888) );
  IV U25563 ( .A(n24840), .Z(n24836) );
  XOR U25564 ( .A(n24891), .B(n24892), .Z(n24840) );
  ANDN U25565 ( .B(n24893), .A(n24894), .Z(n24891) );
  XOR U25566 ( .A(n24895), .B(n24892), .Z(n24893) );
  IV U25567 ( .A(n24850), .Z(n24854) );
  XOR U25568 ( .A(n24850), .B(n24805), .Z(n24852) );
  XOR U25569 ( .A(n24896), .B(n24897), .Z(n24805) );
  AND U25570 ( .A(n562), .B(n24898), .Z(n24896) );
  XOR U25571 ( .A(n24899), .B(n24897), .Z(n24898) );
  NANDN U25572 ( .A(n24807), .B(n24809), .Z(n24850) );
  XOR U25573 ( .A(n24900), .B(n24901), .Z(n24809) );
  AND U25574 ( .A(n562), .B(n24902), .Z(n24900) );
  XOR U25575 ( .A(n24901), .B(n24903), .Z(n24902) );
  XNOR U25576 ( .A(n24904), .B(n24905), .Z(n562) );
  AND U25577 ( .A(n24906), .B(n24907), .Z(n24904) );
  XOR U25578 ( .A(n24905), .B(n24820), .Z(n24907) );
  XNOR U25579 ( .A(n24908), .B(n24909), .Z(n24820) );
  ANDN U25580 ( .B(n24910), .A(n24911), .Z(n24908) );
  XOR U25581 ( .A(n24909), .B(n24912), .Z(n24910) );
  XNOR U25582 ( .A(n24905), .B(n24822), .Z(n24906) );
  XOR U25583 ( .A(n24913), .B(n24914), .Z(n24822) );
  AND U25584 ( .A(n566), .B(n24915), .Z(n24913) );
  XOR U25585 ( .A(n24916), .B(n24914), .Z(n24915) );
  XNOR U25586 ( .A(n24917), .B(n24918), .Z(n24905) );
  AND U25587 ( .A(n24919), .B(n24920), .Z(n24917) );
  XNOR U25588 ( .A(n24918), .B(n24847), .Z(n24920) );
  XOR U25589 ( .A(n24911), .B(n24912), .Z(n24847) );
  XNOR U25590 ( .A(n24921), .B(n24922), .Z(n24912) );
  ANDN U25591 ( .B(n24923), .A(n24924), .Z(n24921) );
  XOR U25592 ( .A(n24925), .B(n24926), .Z(n24923) );
  XOR U25593 ( .A(n24927), .B(n24928), .Z(n24911) );
  XNOR U25594 ( .A(n24929), .B(n24930), .Z(n24928) );
  ANDN U25595 ( .B(n24931), .A(n24932), .Z(n24929) );
  XNOR U25596 ( .A(n24933), .B(n24934), .Z(n24931) );
  IV U25597 ( .A(n24909), .Z(n24927) );
  XOR U25598 ( .A(n24935), .B(n24936), .Z(n24909) );
  ANDN U25599 ( .B(n24937), .A(n24938), .Z(n24935) );
  XOR U25600 ( .A(n24936), .B(n24939), .Z(n24937) );
  XOR U25601 ( .A(n24918), .B(n24849), .Z(n24919) );
  XOR U25602 ( .A(n24940), .B(n24941), .Z(n24849) );
  AND U25603 ( .A(n566), .B(n24942), .Z(n24940) );
  XOR U25604 ( .A(n24943), .B(n24941), .Z(n24942) );
  XNOR U25605 ( .A(n24944), .B(n24945), .Z(n24918) );
  NAND U25606 ( .A(n24946), .B(n24947), .Z(n24945) );
  XOR U25607 ( .A(n24948), .B(n24897), .Z(n24947) );
  XOR U25608 ( .A(n24938), .B(n24939), .Z(n24897) );
  XOR U25609 ( .A(n24949), .B(n24926), .Z(n24939) );
  XOR U25610 ( .A(n24950), .B(n24951), .Z(n24926) );
  ANDN U25611 ( .B(n24952), .A(n24953), .Z(n24950) );
  XOR U25612 ( .A(n24951), .B(n24954), .Z(n24952) );
  IV U25613 ( .A(n24924), .Z(n24949) );
  XOR U25614 ( .A(n24922), .B(n24955), .Z(n24924) );
  XOR U25615 ( .A(n24956), .B(n24957), .Z(n24955) );
  ANDN U25616 ( .B(n24958), .A(n24959), .Z(n24956) );
  XOR U25617 ( .A(n24960), .B(n24957), .Z(n24958) );
  IV U25618 ( .A(n24925), .Z(n24922) );
  XOR U25619 ( .A(n24961), .B(n24962), .Z(n24925) );
  ANDN U25620 ( .B(n24963), .A(n24964), .Z(n24961) );
  XOR U25621 ( .A(n24962), .B(n24965), .Z(n24963) );
  XOR U25622 ( .A(n24966), .B(n24967), .Z(n24938) );
  XNOR U25623 ( .A(n24933), .B(n24968), .Z(n24967) );
  IV U25624 ( .A(n24936), .Z(n24968) );
  XOR U25625 ( .A(n24969), .B(n24970), .Z(n24936) );
  ANDN U25626 ( .B(n24971), .A(n24972), .Z(n24969) );
  XOR U25627 ( .A(n24970), .B(n24973), .Z(n24971) );
  XNOR U25628 ( .A(n24974), .B(n24975), .Z(n24933) );
  ANDN U25629 ( .B(n24976), .A(n24977), .Z(n24974) );
  XOR U25630 ( .A(n24975), .B(n24978), .Z(n24976) );
  IV U25631 ( .A(n24932), .Z(n24966) );
  XOR U25632 ( .A(n24930), .B(n24979), .Z(n24932) );
  XOR U25633 ( .A(n24980), .B(n24981), .Z(n24979) );
  ANDN U25634 ( .B(n24982), .A(n24983), .Z(n24980) );
  XOR U25635 ( .A(n24984), .B(n24981), .Z(n24982) );
  IV U25636 ( .A(n24934), .Z(n24930) );
  XOR U25637 ( .A(n24985), .B(n24986), .Z(n24934) );
  ANDN U25638 ( .B(n24987), .A(n24988), .Z(n24985) );
  XOR U25639 ( .A(n24989), .B(n24986), .Z(n24987) );
  IV U25640 ( .A(n24944), .Z(n24948) );
  XOR U25641 ( .A(n24944), .B(n24899), .Z(n24946) );
  XOR U25642 ( .A(n24990), .B(n24991), .Z(n24899) );
  AND U25643 ( .A(n566), .B(n24992), .Z(n24990) );
  XOR U25644 ( .A(n24993), .B(n24991), .Z(n24992) );
  NANDN U25645 ( .A(n24901), .B(n24903), .Z(n24944) );
  XOR U25646 ( .A(n24994), .B(n24995), .Z(n24903) );
  AND U25647 ( .A(n566), .B(n24996), .Z(n24994) );
  XOR U25648 ( .A(n24995), .B(n24997), .Z(n24996) );
  XNOR U25649 ( .A(n24998), .B(n24999), .Z(n566) );
  AND U25650 ( .A(n25000), .B(n25001), .Z(n24998) );
  XOR U25651 ( .A(n24999), .B(n24914), .Z(n25001) );
  XNOR U25652 ( .A(n25002), .B(n25003), .Z(n24914) );
  ANDN U25653 ( .B(n25004), .A(n25005), .Z(n25002) );
  XOR U25654 ( .A(n25003), .B(n25006), .Z(n25004) );
  XNOR U25655 ( .A(n24999), .B(n24916), .Z(n25000) );
  XOR U25656 ( .A(n25007), .B(n25008), .Z(n24916) );
  AND U25657 ( .A(n570), .B(n25009), .Z(n25007) );
  XOR U25658 ( .A(n25010), .B(n25008), .Z(n25009) );
  XNOR U25659 ( .A(n25011), .B(n25012), .Z(n24999) );
  AND U25660 ( .A(n25013), .B(n25014), .Z(n25011) );
  XNOR U25661 ( .A(n25012), .B(n24941), .Z(n25014) );
  XOR U25662 ( .A(n25005), .B(n25006), .Z(n24941) );
  XNOR U25663 ( .A(n25015), .B(n25016), .Z(n25006) );
  ANDN U25664 ( .B(n25017), .A(n25018), .Z(n25015) );
  XOR U25665 ( .A(n25019), .B(n25020), .Z(n25017) );
  XOR U25666 ( .A(n25021), .B(n25022), .Z(n25005) );
  XNOR U25667 ( .A(n25023), .B(n25024), .Z(n25022) );
  ANDN U25668 ( .B(n25025), .A(n25026), .Z(n25023) );
  XNOR U25669 ( .A(n25027), .B(n25028), .Z(n25025) );
  IV U25670 ( .A(n25003), .Z(n25021) );
  XOR U25671 ( .A(n25029), .B(n25030), .Z(n25003) );
  ANDN U25672 ( .B(n25031), .A(n25032), .Z(n25029) );
  XOR U25673 ( .A(n25030), .B(n25033), .Z(n25031) );
  XOR U25674 ( .A(n25012), .B(n24943), .Z(n25013) );
  XOR U25675 ( .A(n25034), .B(n25035), .Z(n24943) );
  AND U25676 ( .A(n570), .B(n25036), .Z(n25034) );
  XOR U25677 ( .A(n25037), .B(n25035), .Z(n25036) );
  XNOR U25678 ( .A(n25038), .B(n25039), .Z(n25012) );
  NAND U25679 ( .A(n25040), .B(n25041), .Z(n25039) );
  XOR U25680 ( .A(n25042), .B(n24991), .Z(n25041) );
  XOR U25681 ( .A(n25032), .B(n25033), .Z(n24991) );
  XOR U25682 ( .A(n25043), .B(n25020), .Z(n25033) );
  XOR U25683 ( .A(n25044), .B(n25045), .Z(n25020) );
  ANDN U25684 ( .B(n25046), .A(n25047), .Z(n25044) );
  XOR U25685 ( .A(n25045), .B(n25048), .Z(n25046) );
  IV U25686 ( .A(n25018), .Z(n25043) );
  XOR U25687 ( .A(n25016), .B(n25049), .Z(n25018) );
  XOR U25688 ( .A(n25050), .B(n25051), .Z(n25049) );
  ANDN U25689 ( .B(n25052), .A(n25053), .Z(n25050) );
  XOR U25690 ( .A(n25054), .B(n25051), .Z(n25052) );
  IV U25691 ( .A(n25019), .Z(n25016) );
  XOR U25692 ( .A(n25055), .B(n25056), .Z(n25019) );
  ANDN U25693 ( .B(n25057), .A(n25058), .Z(n25055) );
  XOR U25694 ( .A(n25056), .B(n25059), .Z(n25057) );
  XOR U25695 ( .A(n25060), .B(n25061), .Z(n25032) );
  XNOR U25696 ( .A(n25027), .B(n25062), .Z(n25061) );
  IV U25697 ( .A(n25030), .Z(n25062) );
  XOR U25698 ( .A(n25063), .B(n25064), .Z(n25030) );
  ANDN U25699 ( .B(n25065), .A(n25066), .Z(n25063) );
  XOR U25700 ( .A(n25064), .B(n25067), .Z(n25065) );
  XNOR U25701 ( .A(n25068), .B(n25069), .Z(n25027) );
  ANDN U25702 ( .B(n25070), .A(n25071), .Z(n25068) );
  XOR U25703 ( .A(n25069), .B(n25072), .Z(n25070) );
  IV U25704 ( .A(n25026), .Z(n25060) );
  XOR U25705 ( .A(n25024), .B(n25073), .Z(n25026) );
  XOR U25706 ( .A(n25074), .B(n25075), .Z(n25073) );
  ANDN U25707 ( .B(n25076), .A(n25077), .Z(n25074) );
  XOR U25708 ( .A(n25078), .B(n25075), .Z(n25076) );
  IV U25709 ( .A(n25028), .Z(n25024) );
  XOR U25710 ( .A(n25079), .B(n25080), .Z(n25028) );
  ANDN U25711 ( .B(n25081), .A(n25082), .Z(n25079) );
  XOR U25712 ( .A(n25083), .B(n25080), .Z(n25081) );
  IV U25713 ( .A(n25038), .Z(n25042) );
  XOR U25714 ( .A(n25038), .B(n24993), .Z(n25040) );
  XOR U25715 ( .A(n25084), .B(n25085), .Z(n24993) );
  AND U25716 ( .A(n570), .B(n25086), .Z(n25084) );
  XOR U25717 ( .A(n25087), .B(n25085), .Z(n25086) );
  NANDN U25718 ( .A(n24995), .B(n24997), .Z(n25038) );
  XOR U25719 ( .A(n25088), .B(n25089), .Z(n24997) );
  AND U25720 ( .A(n570), .B(n25090), .Z(n25088) );
  XOR U25721 ( .A(n25089), .B(n25091), .Z(n25090) );
  XNOR U25722 ( .A(n25092), .B(n25093), .Z(n570) );
  AND U25723 ( .A(n25094), .B(n25095), .Z(n25092) );
  XOR U25724 ( .A(n25093), .B(n25008), .Z(n25095) );
  XNOR U25725 ( .A(n25096), .B(n25097), .Z(n25008) );
  ANDN U25726 ( .B(n25098), .A(n25099), .Z(n25096) );
  XOR U25727 ( .A(n25097), .B(n25100), .Z(n25098) );
  XNOR U25728 ( .A(n25093), .B(n25010), .Z(n25094) );
  XOR U25729 ( .A(n25101), .B(n25102), .Z(n25010) );
  AND U25730 ( .A(n574), .B(n25103), .Z(n25101) );
  XOR U25731 ( .A(n25104), .B(n25102), .Z(n25103) );
  XNOR U25732 ( .A(n25105), .B(n25106), .Z(n25093) );
  AND U25733 ( .A(n25107), .B(n25108), .Z(n25105) );
  XNOR U25734 ( .A(n25106), .B(n25035), .Z(n25108) );
  XOR U25735 ( .A(n25099), .B(n25100), .Z(n25035) );
  XNOR U25736 ( .A(n25109), .B(n25110), .Z(n25100) );
  ANDN U25737 ( .B(n25111), .A(n25112), .Z(n25109) );
  XOR U25738 ( .A(n25113), .B(n25114), .Z(n25111) );
  XOR U25739 ( .A(n25115), .B(n25116), .Z(n25099) );
  XNOR U25740 ( .A(n25117), .B(n25118), .Z(n25116) );
  ANDN U25741 ( .B(n25119), .A(n25120), .Z(n25117) );
  XNOR U25742 ( .A(n25121), .B(n25122), .Z(n25119) );
  IV U25743 ( .A(n25097), .Z(n25115) );
  XOR U25744 ( .A(n25123), .B(n25124), .Z(n25097) );
  ANDN U25745 ( .B(n25125), .A(n25126), .Z(n25123) );
  XOR U25746 ( .A(n25124), .B(n25127), .Z(n25125) );
  XOR U25747 ( .A(n25106), .B(n25037), .Z(n25107) );
  XOR U25748 ( .A(n25128), .B(n25129), .Z(n25037) );
  AND U25749 ( .A(n574), .B(n25130), .Z(n25128) );
  XOR U25750 ( .A(n25131), .B(n25129), .Z(n25130) );
  XNOR U25751 ( .A(n25132), .B(n25133), .Z(n25106) );
  NAND U25752 ( .A(n25134), .B(n25135), .Z(n25133) );
  XOR U25753 ( .A(n25136), .B(n25085), .Z(n25135) );
  XOR U25754 ( .A(n25126), .B(n25127), .Z(n25085) );
  XOR U25755 ( .A(n25137), .B(n25114), .Z(n25127) );
  XOR U25756 ( .A(n25138), .B(n25139), .Z(n25114) );
  ANDN U25757 ( .B(n25140), .A(n25141), .Z(n25138) );
  XOR U25758 ( .A(n25139), .B(n25142), .Z(n25140) );
  IV U25759 ( .A(n25112), .Z(n25137) );
  XOR U25760 ( .A(n25110), .B(n25143), .Z(n25112) );
  XOR U25761 ( .A(n25144), .B(n25145), .Z(n25143) );
  ANDN U25762 ( .B(n25146), .A(n25147), .Z(n25144) );
  XOR U25763 ( .A(n25148), .B(n25145), .Z(n25146) );
  IV U25764 ( .A(n25113), .Z(n25110) );
  XOR U25765 ( .A(n25149), .B(n25150), .Z(n25113) );
  ANDN U25766 ( .B(n25151), .A(n25152), .Z(n25149) );
  XOR U25767 ( .A(n25150), .B(n25153), .Z(n25151) );
  XOR U25768 ( .A(n25154), .B(n25155), .Z(n25126) );
  XNOR U25769 ( .A(n25121), .B(n25156), .Z(n25155) );
  IV U25770 ( .A(n25124), .Z(n25156) );
  XOR U25771 ( .A(n25157), .B(n25158), .Z(n25124) );
  ANDN U25772 ( .B(n25159), .A(n25160), .Z(n25157) );
  XOR U25773 ( .A(n25158), .B(n25161), .Z(n25159) );
  XNOR U25774 ( .A(n25162), .B(n25163), .Z(n25121) );
  ANDN U25775 ( .B(n25164), .A(n25165), .Z(n25162) );
  XOR U25776 ( .A(n25163), .B(n25166), .Z(n25164) );
  IV U25777 ( .A(n25120), .Z(n25154) );
  XOR U25778 ( .A(n25118), .B(n25167), .Z(n25120) );
  XOR U25779 ( .A(n25168), .B(n25169), .Z(n25167) );
  ANDN U25780 ( .B(n25170), .A(n25171), .Z(n25168) );
  XOR U25781 ( .A(n25172), .B(n25169), .Z(n25170) );
  IV U25782 ( .A(n25122), .Z(n25118) );
  XOR U25783 ( .A(n25173), .B(n25174), .Z(n25122) );
  ANDN U25784 ( .B(n25175), .A(n25176), .Z(n25173) );
  XOR U25785 ( .A(n25177), .B(n25174), .Z(n25175) );
  IV U25786 ( .A(n25132), .Z(n25136) );
  XOR U25787 ( .A(n25132), .B(n25087), .Z(n25134) );
  XOR U25788 ( .A(n25178), .B(n25179), .Z(n25087) );
  AND U25789 ( .A(n574), .B(n25180), .Z(n25178) );
  XOR U25790 ( .A(n25181), .B(n25179), .Z(n25180) );
  NANDN U25791 ( .A(n25089), .B(n25091), .Z(n25132) );
  XOR U25792 ( .A(n25182), .B(n25183), .Z(n25091) );
  AND U25793 ( .A(n574), .B(n25184), .Z(n25182) );
  XOR U25794 ( .A(n25183), .B(n25185), .Z(n25184) );
  XNOR U25795 ( .A(n25186), .B(n25187), .Z(n574) );
  AND U25796 ( .A(n25188), .B(n25189), .Z(n25186) );
  XOR U25797 ( .A(n25187), .B(n25102), .Z(n25189) );
  XNOR U25798 ( .A(n25190), .B(n25191), .Z(n25102) );
  ANDN U25799 ( .B(n25192), .A(n25193), .Z(n25190) );
  XOR U25800 ( .A(n25191), .B(n25194), .Z(n25192) );
  XNOR U25801 ( .A(n25187), .B(n25104), .Z(n25188) );
  XOR U25802 ( .A(n25195), .B(n25196), .Z(n25104) );
  AND U25803 ( .A(n578), .B(n25197), .Z(n25195) );
  XOR U25804 ( .A(n25198), .B(n25196), .Z(n25197) );
  XNOR U25805 ( .A(n25199), .B(n25200), .Z(n25187) );
  AND U25806 ( .A(n25201), .B(n25202), .Z(n25199) );
  XNOR U25807 ( .A(n25200), .B(n25129), .Z(n25202) );
  XOR U25808 ( .A(n25193), .B(n25194), .Z(n25129) );
  XNOR U25809 ( .A(n25203), .B(n25204), .Z(n25194) );
  ANDN U25810 ( .B(n25205), .A(n25206), .Z(n25203) );
  XOR U25811 ( .A(n25207), .B(n25208), .Z(n25205) );
  XOR U25812 ( .A(n25209), .B(n25210), .Z(n25193) );
  XNOR U25813 ( .A(n25211), .B(n25212), .Z(n25210) );
  ANDN U25814 ( .B(n25213), .A(n25214), .Z(n25211) );
  XNOR U25815 ( .A(n25215), .B(n25216), .Z(n25213) );
  IV U25816 ( .A(n25191), .Z(n25209) );
  XOR U25817 ( .A(n25217), .B(n25218), .Z(n25191) );
  ANDN U25818 ( .B(n25219), .A(n25220), .Z(n25217) );
  XOR U25819 ( .A(n25218), .B(n25221), .Z(n25219) );
  XOR U25820 ( .A(n25200), .B(n25131), .Z(n25201) );
  XOR U25821 ( .A(n25222), .B(n25223), .Z(n25131) );
  AND U25822 ( .A(n578), .B(n25224), .Z(n25222) );
  XOR U25823 ( .A(n25225), .B(n25223), .Z(n25224) );
  XNOR U25824 ( .A(n25226), .B(n25227), .Z(n25200) );
  NAND U25825 ( .A(n25228), .B(n25229), .Z(n25227) );
  XOR U25826 ( .A(n25230), .B(n25179), .Z(n25229) );
  XOR U25827 ( .A(n25220), .B(n25221), .Z(n25179) );
  XOR U25828 ( .A(n25231), .B(n25208), .Z(n25221) );
  XOR U25829 ( .A(n25232), .B(n25233), .Z(n25208) );
  ANDN U25830 ( .B(n25234), .A(n25235), .Z(n25232) );
  XOR U25831 ( .A(n25233), .B(n25236), .Z(n25234) );
  IV U25832 ( .A(n25206), .Z(n25231) );
  XOR U25833 ( .A(n25204), .B(n25237), .Z(n25206) );
  XOR U25834 ( .A(n25238), .B(n25239), .Z(n25237) );
  ANDN U25835 ( .B(n25240), .A(n25241), .Z(n25238) );
  XOR U25836 ( .A(n25242), .B(n25239), .Z(n25240) );
  IV U25837 ( .A(n25207), .Z(n25204) );
  XOR U25838 ( .A(n25243), .B(n25244), .Z(n25207) );
  ANDN U25839 ( .B(n25245), .A(n25246), .Z(n25243) );
  XOR U25840 ( .A(n25244), .B(n25247), .Z(n25245) );
  XOR U25841 ( .A(n25248), .B(n25249), .Z(n25220) );
  XNOR U25842 ( .A(n25215), .B(n25250), .Z(n25249) );
  IV U25843 ( .A(n25218), .Z(n25250) );
  XOR U25844 ( .A(n25251), .B(n25252), .Z(n25218) );
  ANDN U25845 ( .B(n25253), .A(n25254), .Z(n25251) );
  XOR U25846 ( .A(n25252), .B(n25255), .Z(n25253) );
  XNOR U25847 ( .A(n25256), .B(n25257), .Z(n25215) );
  ANDN U25848 ( .B(n25258), .A(n25259), .Z(n25256) );
  XOR U25849 ( .A(n25257), .B(n25260), .Z(n25258) );
  IV U25850 ( .A(n25214), .Z(n25248) );
  XOR U25851 ( .A(n25212), .B(n25261), .Z(n25214) );
  XOR U25852 ( .A(n25262), .B(n25263), .Z(n25261) );
  ANDN U25853 ( .B(n25264), .A(n25265), .Z(n25262) );
  XOR U25854 ( .A(n25266), .B(n25263), .Z(n25264) );
  IV U25855 ( .A(n25216), .Z(n25212) );
  XOR U25856 ( .A(n25267), .B(n25268), .Z(n25216) );
  ANDN U25857 ( .B(n25269), .A(n25270), .Z(n25267) );
  XOR U25858 ( .A(n25271), .B(n25268), .Z(n25269) );
  IV U25859 ( .A(n25226), .Z(n25230) );
  XOR U25860 ( .A(n25226), .B(n25181), .Z(n25228) );
  XOR U25861 ( .A(n25272), .B(n25273), .Z(n25181) );
  AND U25862 ( .A(n578), .B(n25274), .Z(n25272) );
  XOR U25863 ( .A(n25275), .B(n25273), .Z(n25274) );
  NANDN U25864 ( .A(n25183), .B(n25185), .Z(n25226) );
  XOR U25865 ( .A(n25276), .B(n25277), .Z(n25185) );
  AND U25866 ( .A(n578), .B(n25278), .Z(n25276) );
  XOR U25867 ( .A(n25277), .B(n25279), .Z(n25278) );
  XNOR U25868 ( .A(n25280), .B(n25281), .Z(n578) );
  AND U25869 ( .A(n25282), .B(n25283), .Z(n25280) );
  XOR U25870 ( .A(n25281), .B(n25196), .Z(n25283) );
  XNOR U25871 ( .A(n25284), .B(n25285), .Z(n25196) );
  ANDN U25872 ( .B(n25286), .A(n25287), .Z(n25284) );
  XOR U25873 ( .A(n25285), .B(n25288), .Z(n25286) );
  XNOR U25874 ( .A(n25281), .B(n25198), .Z(n25282) );
  XOR U25875 ( .A(n25289), .B(n25290), .Z(n25198) );
  AND U25876 ( .A(n582), .B(n25291), .Z(n25289) );
  XOR U25877 ( .A(n25292), .B(n25290), .Z(n25291) );
  XNOR U25878 ( .A(n25293), .B(n25294), .Z(n25281) );
  AND U25879 ( .A(n25295), .B(n25296), .Z(n25293) );
  XNOR U25880 ( .A(n25294), .B(n25223), .Z(n25296) );
  XOR U25881 ( .A(n25287), .B(n25288), .Z(n25223) );
  XNOR U25882 ( .A(n25297), .B(n25298), .Z(n25288) );
  ANDN U25883 ( .B(n25299), .A(n25300), .Z(n25297) );
  XOR U25884 ( .A(n25301), .B(n25302), .Z(n25299) );
  XOR U25885 ( .A(n25303), .B(n25304), .Z(n25287) );
  XNOR U25886 ( .A(n25305), .B(n25306), .Z(n25304) );
  ANDN U25887 ( .B(n25307), .A(n25308), .Z(n25305) );
  XNOR U25888 ( .A(n25309), .B(n25310), .Z(n25307) );
  IV U25889 ( .A(n25285), .Z(n25303) );
  XOR U25890 ( .A(n25311), .B(n25312), .Z(n25285) );
  ANDN U25891 ( .B(n25313), .A(n25314), .Z(n25311) );
  XOR U25892 ( .A(n25312), .B(n25315), .Z(n25313) );
  XOR U25893 ( .A(n25294), .B(n25225), .Z(n25295) );
  XOR U25894 ( .A(n25316), .B(n25317), .Z(n25225) );
  AND U25895 ( .A(n582), .B(n25318), .Z(n25316) );
  XOR U25896 ( .A(n25319), .B(n25317), .Z(n25318) );
  XNOR U25897 ( .A(n25320), .B(n25321), .Z(n25294) );
  NAND U25898 ( .A(n25322), .B(n25323), .Z(n25321) );
  XOR U25899 ( .A(n25324), .B(n25273), .Z(n25323) );
  XOR U25900 ( .A(n25314), .B(n25315), .Z(n25273) );
  XOR U25901 ( .A(n25325), .B(n25302), .Z(n25315) );
  XOR U25902 ( .A(n25326), .B(n25327), .Z(n25302) );
  ANDN U25903 ( .B(n25328), .A(n25329), .Z(n25326) );
  XOR U25904 ( .A(n25327), .B(n25330), .Z(n25328) );
  IV U25905 ( .A(n25300), .Z(n25325) );
  XOR U25906 ( .A(n25298), .B(n25331), .Z(n25300) );
  XOR U25907 ( .A(n25332), .B(n25333), .Z(n25331) );
  ANDN U25908 ( .B(n25334), .A(n25335), .Z(n25332) );
  XOR U25909 ( .A(n25336), .B(n25333), .Z(n25334) );
  IV U25910 ( .A(n25301), .Z(n25298) );
  XOR U25911 ( .A(n25337), .B(n25338), .Z(n25301) );
  ANDN U25912 ( .B(n25339), .A(n25340), .Z(n25337) );
  XOR U25913 ( .A(n25338), .B(n25341), .Z(n25339) );
  XOR U25914 ( .A(n25342), .B(n25343), .Z(n25314) );
  XNOR U25915 ( .A(n25309), .B(n25344), .Z(n25343) );
  IV U25916 ( .A(n25312), .Z(n25344) );
  XOR U25917 ( .A(n25345), .B(n25346), .Z(n25312) );
  ANDN U25918 ( .B(n25347), .A(n25348), .Z(n25345) );
  XOR U25919 ( .A(n25346), .B(n25349), .Z(n25347) );
  XNOR U25920 ( .A(n25350), .B(n25351), .Z(n25309) );
  ANDN U25921 ( .B(n25352), .A(n25353), .Z(n25350) );
  XOR U25922 ( .A(n25351), .B(n25354), .Z(n25352) );
  IV U25923 ( .A(n25308), .Z(n25342) );
  XOR U25924 ( .A(n25306), .B(n25355), .Z(n25308) );
  XOR U25925 ( .A(n25356), .B(n25357), .Z(n25355) );
  ANDN U25926 ( .B(n25358), .A(n25359), .Z(n25356) );
  XOR U25927 ( .A(n25360), .B(n25357), .Z(n25358) );
  IV U25928 ( .A(n25310), .Z(n25306) );
  XOR U25929 ( .A(n25361), .B(n25362), .Z(n25310) );
  ANDN U25930 ( .B(n25363), .A(n25364), .Z(n25361) );
  XOR U25931 ( .A(n25365), .B(n25362), .Z(n25363) );
  IV U25932 ( .A(n25320), .Z(n25324) );
  XOR U25933 ( .A(n25320), .B(n25275), .Z(n25322) );
  XOR U25934 ( .A(n25366), .B(n25367), .Z(n25275) );
  AND U25935 ( .A(n582), .B(n25368), .Z(n25366) );
  XOR U25936 ( .A(n25369), .B(n25367), .Z(n25368) );
  NANDN U25937 ( .A(n25277), .B(n25279), .Z(n25320) );
  XOR U25938 ( .A(n25370), .B(n25371), .Z(n25279) );
  AND U25939 ( .A(n582), .B(n25372), .Z(n25370) );
  XOR U25940 ( .A(n25371), .B(n25373), .Z(n25372) );
  XNOR U25941 ( .A(n25374), .B(n25375), .Z(n582) );
  AND U25942 ( .A(n25376), .B(n25377), .Z(n25374) );
  XOR U25943 ( .A(n25375), .B(n25290), .Z(n25377) );
  XNOR U25944 ( .A(n25378), .B(n25379), .Z(n25290) );
  ANDN U25945 ( .B(n25380), .A(n25381), .Z(n25378) );
  XOR U25946 ( .A(n25379), .B(n25382), .Z(n25380) );
  XNOR U25947 ( .A(n25375), .B(n25292), .Z(n25376) );
  XOR U25948 ( .A(n25383), .B(n25384), .Z(n25292) );
  AND U25949 ( .A(n586), .B(n25385), .Z(n25383) );
  XOR U25950 ( .A(n25386), .B(n25384), .Z(n25385) );
  XNOR U25951 ( .A(n25387), .B(n25388), .Z(n25375) );
  AND U25952 ( .A(n25389), .B(n25390), .Z(n25387) );
  XNOR U25953 ( .A(n25388), .B(n25317), .Z(n25390) );
  XOR U25954 ( .A(n25381), .B(n25382), .Z(n25317) );
  XNOR U25955 ( .A(n25391), .B(n25392), .Z(n25382) );
  ANDN U25956 ( .B(n25393), .A(n25394), .Z(n25391) );
  XOR U25957 ( .A(n25395), .B(n25396), .Z(n25393) );
  XOR U25958 ( .A(n25397), .B(n25398), .Z(n25381) );
  XNOR U25959 ( .A(n25399), .B(n25400), .Z(n25398) );
  ANDN U25960 ( .B(n25401), .A(n25402), .Z(n25399) );
  XNOR U25961 ( .A(n25403), .B(n25404), .Z(n25401) );
  IV U25962 ( .A(n25379), .Z(n25397) );
  XOR U25963 ( .A(n25405), .B(n25406), .Z(n25379) );
  ANDN U25964 ( .B(n25407), .A(n25408), .Z(n25405) );
  XOR U25965 ( .A(n25406), .B(n25409), .Z(n25407) );
  XOR U25966 ( .A(n25388), .B(n25319), .Z(n25389) );
  XOR U25967 ( .A(n25410), .B(n25411), .Z(n25319) );
  AND U25968 ( .A(n586), .B(n25412), .Z(n25410) );
  XOR U25969 ( .A(n25413), .B(n25411), .Z(n25412) );
  XNOR U25970 ( .A(n25414), .B(n25415), .Z(n25388) );
  NAND U25971 ( .A(n25416), .B(n25417), .Z(n25415) );
  XOR U25972 ( .A(n25418), .B(n25367), .Z(n25417) );
  XOR U25973 ( .A(n25408), .B(n25409), .Z(n25367) );
  XOR U25974 ( .A(n25419), .B(n25396), .Z(n25409) );
  XOR U25975 ( .A(n25420), .B(n25421), .Z(n25396) );
  ANDN U25976 ( .B(n25422), .A(n25423), .Z(n25420) );
  XOR U25977 ( .A(n25421), .B(n25424), .Z(n25422) );
  IV U25978 ( .A(n25394), .Z(n25419) );
  XOR U25979 ( .A(n25392), .B(n25425), .Z(n25394) );
  XOR U25980 ( .A(n25426), .B(n25427), .Z(n25425) );
  ANDN U25981 ( .B(n25428), .A(n25429), .Z(n25426) );
  XOR U25982 ( .A(n25430), .B(n25427), .Z(n25428) );
  IV U25983 ( .A(n25395), .Z(n25392) );
  XOR U25984 ( .A(n25431), .B(n25432), .Z(n25395) );
  ANDN U25985 ( .B(n25433), .A(n25434), .Z(n25431) );
  XOR U25986 ( .A(n25432), .B(n25435), .Z(n25433) );
  XOR U25987 ( .A(n25436), .B(n25437), .Z(n25408) );
  XNOR U25988 ( .A(n25403), .B(n25438), .Z(n25437) );
  IV U25989 ( .A(n25406), .Z(n25438) );
  XOR U25990 ( .A(n25439), .B(n25440), .Z(n25406) );
  ANDN U25991 ( .B(n25441), .A(n25442), .Z(n25439) );
  XOR U25992 ( .A(n25440), .B(n25443), .Z(n25441) );
  XNOR U25993 ( .A(n25444), .B(n25445), .Z(n25403) );
  ANDN U25994 ( .B(n25446), .A(n25447), .Z(n25444) );
  XOR U25995 ( .A(n25445), .B(n25448), .Z(n25446) );
  IV U25996 ( .A(n25402), .Z(n25436) );
  XOR U25997 ( .A(n25400), .B(n25449), .Z(n25402) );
  XOR U25998 ( .A(n25450), .B(n25451), .Z(n25449) );
  ANDN U25999 ( .B(n25452), .A(n25453), .Z(n25450) );
  XOR U26000 ( .A(n25454), .B(n25451), .Z(n25452) );
  IV U26001 ( .A(n25404), .Z(n25400) );
  XOR U26002 ( .A(n25455), .B(n25456), .Z(n25404) );
  ANDN U26003 ( .B(n25457), .A(n25458), .Z(n25455) );
  XOR U26004 ( .A(n25459), .B(n25456), .Z(n25457) );
  IV U26005 ( .A(n25414), .Z(n25418) );
  XOR U26006 ( .A(n25414), .B(n25369), .Z(n25416) );
  XOR U26007 ( .A(n25460), .B(n25461), .Z(n25369) );
  AND U26008 ( .A(n586), .B(n25462), .Z(n25460) );
  XOR U26009 ( .A(n25463), .B(n25461), .Z(n25462) );
  NANDN U26010 ( .A(n25371), .B(n25373), .Z(n25414) );
  XOR U26011 ( .A(n25464), .B(n25465), .Z(n25373) );
  AND U26012 ( .A(n586), .B(n25466), .Z(n25464) );
  XOR U26013 ( .A(n25465), .B(n25467), .Z(n25466) );
  XNOR U26014 ( .A(n25468), .B(n25469), .Z(n586) );
  AND U26015 ( .A(n25470), .B(n25471), .Z(n25468) );
  XOR U26016 ( .A(n25469), .B(n25384), .Z(n25471) );
  XNOR U26017 ( .A(n25472), .B(n25473), .Z(n25384) );
  ANDN U26018 ( .B(n25474), .A(n25475), .Z(n25472) );
  XOR U26019 ( .A(n25473), .B(n25476), .Z(n25474) );
  XNOR U26020 ( .A(n25469), .B(n25386), .Z(n25470) );
  XOR U26021 ( .A(n25477), .B(n25478), .Z(n25386) );
  AND U26022 ( .A(n590), .B(n25479), .Z(n25477) );
  XOR U26023 ( .A(n25480), .B(n25478), .Z(n25479) );
  XNOR U26024 ( .A(n25481), .B(n25482), .Z(n25469) );
  AND U26025 ( .A(n25483), .B(n25484), .Z(n25481) );
  XNOR U26026 ( .A(n25482), .B(n25411), .Z(n25484) );
  XOR U26027 ( .A(n25475), .B(n25476), .Z(n25411) );
  XNOR U26028 ( .A(n25485), .B(n25486), .Z(n25476) );
  ANDN U26029 ( .B(n25487), .A(n25488), .Z(n25485) );
  XOR U26030 ( .A(n25489), .B(n25490), .Z(n25487) );
  XOR U26031 ( .A(n25491), .B(n25492), .Z(n25475) );
  XNOR U26032 ( .A(n25493), .B(n25494), .Z(n25492) );
  ANDN U26033 ( .B(n25495), .A(n25496), .Z(n25493) );
  XNOR U26034 ( .A(n25497), .B(n25498), .Z(n25495) );
  IV U26035 ( .A(n25473), .Z(n25491) );
  XOR U26036 ( .A(n25499), .B(n25500), .Z(n25473) );
  ANDN U26037 ( .B(n25501), .A(n25502), .Z(n25499) );
  XOR U26038 ( .A(n25500), .B(n25503), .Z(n25501) );
  XOR U26039 ( .A(n25482), .B(n25413), .Z(n25483) );
  XOR U26040 ( .A(n25504), .B(n25505), .Z(n25413) );
  AND U26041 ( .A(n590), .B(n25506), .Z(n25504) );
  XOR U26042 ( .A(n25507), .B(n25505), .Z(n25506) );
  XNOR U26043 ( .A(n25508), .B(n25509), .Z(n25482) );
  NAND U26044 ( .A(n25510), .B(n25511), .Z(n25509) );
  XOR U26045 ( .A(n25512), .B(n25461), .Z(n25511) );
  XOR U26046 ( .A(n25502), .B(n25503), .Z(n25461) );
  XOR U26047 ( .A(n25513), .B(n25490), .Z(n25503) );
  XOR U26048 ( .A(n25514), .B(n25515), .Z(n25490) );
  ANDN U26049 ( .B(n25516), .A(n25517), .Z(n25514) );
  XOR U26050 ( .A(n25515), .B(n25518), .Z(n25516) );
  IV U26051 ( .A(n25488), .Z(n25513) );
  XOR U26052 ( .A(n25486), .B(n25519), .Z(n25488) );
  XOR U26053 ( .A(n25520), .B(n25521), .Z(n25519) );
  ANDN U26054 ( .B(n25522), .A(n25523), .Z(n25520) );
  XOR U26055 ( .A(n25524), .B(n25521), .Z(n25522) );
  IV U26056 ( .A(n25489), .Z(n25486) );
  XOR U26057 ( .A(n25525), .B(n25526), .Z(n25489) );
  ANDN U26058 ( .B(n25527), .A(n25528), .Z(n25525) );
  XOR U26059 ( .A(n25526), .B(n25529), .Z(n25527) );
  XOR U26060 ( .A(n25530), .B(n25531), .Z(n25502) );
  XNOR U26061 ( .A(n25497), .B(n25532), .Z(n25531) );
  IV U26062 ( .A(n25500), .Z(n25532) );
  XOR U26063 ( .A(n25533), .B(n25534), .Z(n25500) );
  ANDN U26064 ( .B(n25535), .A(n25536), .Z(n25533) );
  XOR U26065 ( .A(n25534), .B(n25537), .Z(n25535) );
  XNOR U26066 ( .A(n25538), .B(n25539), .Z(n25497) );
  ANDN U26067 ( .B(n25540), .A(n25541), .Z(n25538) );
  XOR U26068 ( .A(n25539), .B(n25542), .Z(n25540) );
  IV U26069 ( .A(n25496), .Z(n25530) );
  XOR U26070 ( .A(n25494), .B(n25543), .Z(n25496) );
  XOR U26071 ( .A(n25544), .B(n25545), .Z(n25543) );
  ANDN U26072 ( .B(n25546), .A(n25547), .Z(n25544) );
  XOR U26073 ( .A(n25548), .B(n25545), .Z(n25546) );
  IV U26074 ( .A(n25498), .Z(n25494) );
  XOR U26075 ( .A(n25549), .B(n25550), .Z(n25498) );
  ANDN U26076 ( .B(n25551), .A(n25552), .Z(n25549) );
  XOR U26077 ( .A(n25553), .B(n25550), .Z(n25551) );
  IV U26078 ( .A(n25508), .Z(n25512) );
  XOR U26079 ( .A(n25508), .B(n25463), .Z(n25510) );
  XOR U26080 ( .A(n25554), .B(n25555), .Z(n25463) );
  AND U26081 ( .A(n590), .B(n25556), .Z(n25554) );
  XOR U26082 ( .A(n25557), .B(n25555), .Z(n25556) );
  NANDN U26083 ( .A(n25465), .B(n25467), .Z(n25508) );
  XOR U26084 ( .A(n25558), .B(n25559), .Z(n25467) );
  AND U26085 ( .A(n590), .B(n25560), .Z(n25558) );
  XOR U26086 ( .A(n25559), .B(n25561), .Z(n25560) );
  XNOR U26087 ( .A(n25562), .B(n25563), .Z(n590) );
  AND U26088 ( .A(n25564), .B(n25565), .Z(n25562) );
  XOR U26089 ( .A(n25563), .B(n25478), .Z(n25565) );
  XNOR U26090 ( .A(n25566), .B(n25567), .Z(n25478) );
  ANDN U26091 ( .B(n25568), .A(n25569), .Z(n25566) );
  XOR U26092 ( .A(n25567), .B(n25570), .Z(n25568) );
  XNOR U26093 ( .A(n25563), .B(n25480), .Z(n25564) );
  XOR U26094 ( .A(n25571), .B(n25572), .Z(n25480) );
  AND U26095 ( .A(n594), .B(n25573), .Z(n25571) );
  XOR U26096 ( .A(n25574), .B(n25572), .Z(n25573) );
  XNOR U26097 ( .A(n25575), .B(n25576), .Z(n25563) );
  AND U26098 ( .A(n25577), .B(n25578), .Z(n25575) );
  XNOR U26099 ( .A(n25576), .B(n25505), .Z(n25578) );
  XOR U26100 ( .A(n25569), .B(n25570), .Z(n25505) );
  XNOR U26101 ( .A(n25579), .B(n25580), .Z(n25570) );
  ANDN U26102 ( .B(n25581), .A(n25582), .Z(n25579) );
  XOR U26103 ( .A(n25583), .B(n25584), .Z(n25581) );
  XOR U26104 ( .A(n25585), .B(n25586), .Z(n25569) );
  XNOR U26105 ( .A(n25587), .B(n25588), .Z(n25586) );
  ANDN U26106 ( .B(n25589), .A(n25590), .Z(n25587) );
  XNOR U26107 ( .A(n25591), .B(n25592), .Z(n25589) );
  IV U26108 ( .A(n25567), .Z(n25585) );
  XOR U26109 ( .A(n25593), .B(n25594), .Z(n25567) );
  ANDN U26110 ( .B(n25595), .A(n25596), .Z(n25593) );
  XOR U26111 ( .A(n25594), .B(n25597), .Z(n25595) );
  XOR U26112 ( .A(n25576), .B(n25507), .Z(n25577) );
  XOR U26113 ( .A(n25598), .B(n25599), .Z(n25507) );
  AND U26114 ( .A(n594), .B(n25600), .Z(n25598) );
  XOR U26115 ( .A(n25601), .B(n25599), .Z(n25600) );
  XNOR U26116 ( .A(n25602), .B(n25603), .Z(n25576) );
  NAND U26117 ( .A(n25604), .B(n25605), .Z(n25603) );
  XOR U26118 ( .A(n25606), .B(n25555), .Z(n25605) );
  XOR U26119 ( .A(n25596), .B(n25597), .Z(n25555) );
  XOR U26120 ( .A(n25607), .B(n25584), .Z(n25597) );
  XOR U26121 ( .A(n25608), .B(n25609), .Z(n25584) );
  ANDN U26122 ( .B(n25610), .A(n25611), .Z(n25608) );
  XOR U26123 ( .A(n25609), .B(n25612), .Z(n25610) );
  IV U26124 ( .A(n25582), .Z(n25607) );
  XOR U26125 ( .A(n25580), .B(n25613), .Z(n25582) );
  XOR U26126 ( .A(n25614), .B(n25615), .Z(n25613) );
  ANDN U26127 ( .B(n25616), .A(n25617), .Z(n25614) );
  XOR U26128 ( .A(n25618), .B(n25615), .Z(n25616) );
  IV U26129 ( .A(n25583), .Z(n25580) );
  XOR U26130 ( .A(n25619), .B(n25620), .Z(n25583) );
  ANDN U26131 ( .B(n25621), .A(n25622), .Z(n25619) );
  XOR U26132 ( .A(n25620), .B(n25623), .Z(n25621) );
  XOR U26133 ( .A(n25624), .B(n25625), .Z(n25596) );
  XNOR U26134 ( .A(n25591), .B(n25626), .Z(n25625) );
  IV U26135 ( .A(n25594), .Z(n25626) );
  XOR U26136 ( .A(n25627), .B(n25628), .Z(n25594) );
  ANDN U26137 ( .B(n25629), .A(n25630), .Z(n25627) );
  XOR U26138 ( .A(n25628), .B(n25631), .Z(n25629) );
  XNOR U26139 ( .A(n25632), .B(n25633), .Z(n25591) );
  ANDN U26140 ( .B(n25634), .A(n25635), .Z(n25632) );
  XOR U26141 ( .A(n25633), .B(n25636), .Z(n25634) );
  IV U26142 ( .A(n25590), .Z(n25624) );
  XOR U26143 ( .A(n25588), .B(n25637), .Z(n25590) );
  XOR U26144 ( .A(n25638), .B(n25639), .Z(n25637) );
  ANDN U26145 ( .B(n25640), .A(n25641), .Z(n25638) );
  XOR U26146 ( .A(n25642), .B(n25639), .Z(n25640) );
  IV U26147 ( .A(n25592), .Z(n25588) );
  XOR U26148 ( .A(n25643), .B(n25644), .Z(n25592) );
  ANDN U26149 ( .B(n25645), .A(n25646), .Z(n25643) );
  XOR U26150 ( .A(n25647), .B(n25644), .Z(n25645) );
  IV U26151 ( .A(n25602), .Z(n25606) );
  XOR U26152 ( .A(n25602), .B(n25557), .Z(n25604) );
  XOR U26153 ( .A(n25648), .B(n25649), .Z(n25557) );
  AND U26154 ( .A(n594), .B(n25650), .Z(n25648) );
  XOR U26155 ( .A(n25651), .B(n25649), .Z(n25650) );
  NANDN U26156 ( .A(n25559), .B(n25561), .Z(n25602) );
  XOR U26157 ( .A(n25652), .B(n25653), .Z(n25561) );
  AND U26158 ( .A(n594), .B(n25654), .Z(n25652) );
  XOR U26159 ( .A(n25653), .B(n25655), .Z(n25654) );
  XNOR U26160 ( .A(n25656), .B(n25657), .Z(n594) );
  AND U26161 ( .A(n25658), .B(n25659), .Z(n25656) );
  XOR U26162 ( .A(n25657), .B(n25572), .Z(n25659) );
  XNOR U26163 ( .A(n25660), .B(n25661), .Z(n25572) );
  ANDN U26164 ( .B(n25662), .A(n25663), .Z(n25660) );
  XOR U26165 ( .A(n25661), .B(n25664), .Z(n25662) );
  XNOR U26166 ( .A(n25657), .B(n25574), .Z(n25658) );
  XOR U26167 ( .A(n25665), .B(n25666), .Z(n25574) );
  AND U26168 ( .A(n598), .B(n25667), .Z(n25665) );
  XOR U26169 ( .A(n25668), .B(n25666), .Z(n25667) );
  XNOR U26170 ( .A(n25669), .B(n25670), .Z(n25657) );
  AND U26171 ( .A(n25671), .B(n25672), .Z(n25669) );
  XNOR U26172 ( .A(n25670), .B(n25599), .Z(n25672) );
  XOR U26173 ( .A(n25663), .B(n25664), .Z(n25599) );
  XNOR U26174 ( .A(n25673), .B(n25674), .Z(n25664) );
  ANDN U26175 ( .B(n25675), .A(n25676), .Z(n25673) );
  XOR U26176 ( .A(n25677), .B(n25678), .Z(n25675) );
  XOR U26177 ( .A(n25679), .B(n25680), .Z(n25663) );
  XNOR U26178 ( .A(n25681), .B(n25682), .Z(n25680) );
  ANDN U26179 ( .B(n25683), .A(n25684), .Z(n25681) );
  XNOR U26180 ( .A(n25685), .B(n25686), .Z(n25683) );
  IV U26181 ( .A(n25661), .Z(n25679) );
  XOR U26182 ( .A(n25687), .B(n25688), .Z(n25661) );
  ANDN U26183 ( .B(n25689), .A(n25690), .Z(n25687) );
  XOR U26184 ( .A(n25688), .B(n25691), .Z(n25689) );
  XOR U26185 ( .A(n25670), .B(n25601), .Z(n25671) );
  XOR U26186 ( .A(n25692), .B(n25693), .Z(n25601) );
  AND U26187 ( .A(n598), .B(n25694), .Z(n25692) );
  XOR U26188 ( .A(n25695), .B(n25693), .Z(n25694) );
  XNOR U26189 ( .A(n25696), .B(n25697), .Z(n25670) );
  NAND U26190 ( .A(n25698), .B(n25699), .Z(n25697) );
  XOR U26191 ( .A(n25700), .B(n25649), .Z(n25699) );
  XOR U26192 ( .A(n25690), .B(n25691), .Z(n25649) );
  XOR U26193 ( .A(n25701), .B(n25678), .Z(n25691) );
  XOR U26194 ( .A(n25702), .B(n25703), .Z(n25678) );
  ANDN U26195 ( .B(n25704), .A(n25705), .Z(n25702) );
  XOR U26196 ( .A(n25703), .B(n25706), .Z(n25704) );
  IV U26197 ( .A(n25676), .Z(n25701) );
  XOR U26198 ( .A(n25674), .B(n25707), .Z(n25676) );
  XOR U26199 ( .A(n25708), .B(n25709), .Z(n25707) );
  ANDN U26200 ( .B(n25710), .A(n25711), .Z(n25708) );
  XOR U26201 ( .A(n25712), .B(n25709), .Z(n25710) );
  IV U26202 ( .A(n25677), .Z(n25674) );
  XOR U26203 ( .A(n25713), .B(n25714), .Z(n25677) );
  ANDN U26204 ( .B(n25715), .A(n25716), .Z(n25713) );
  XOR U26205 ( .A(n25714), .B(n25717), .Z(n25715) );
  XOR U26206 ( .A(n25718), .B(n25719), .Z(n25690) );
  XNOR U26207 ( .A(n25685), .B(n25720), .Z(n25719) );
  IV U26208 ( .A(n25688), .Z(n25720) );
  XOR U26209 ( .A(n25721), .B(n25722), .Z(n25688) );
  ANDN U26210 ( .B(n25723), .A(n25724), .Z(n25721) );
  XOR U26211 ( .A(n25722), .B(n25725), .Z(n25723) );
  XNOR U26212 ( .A(n25726), .B(n25727), .Z(n25685) );
  ANDN U26213 ( .B(n25728), .A(n25729), .Z(n25726) );
  XOR U26214 ( .A(n25727), .B(n25730), .Z(n25728) );
  IV U26215 ( .A(n25684), .Z(n25718) );
  XOR U26216 ( .A(n25682), .B(n25731), .Z(n25684) );
  XOR U26217 ( .A(n25732), .B(n25733), .Z(n25731) );
  ANDN U26218 ( .B(n25734), .A(n25735), .Z(n25732) );
  XOR U26219 ( .A(n25736), .B(n25733), .Z(n25734) );
  IV U26220 ( .A(n25686), .Z(n25682) );
  XOR U26221 ( .A(n25737), .B(n25738), .Z(n25686) );
  ANDN U26222 ( .B(n25739), .A(n25740), .Z(n25737) );
  XOR U26223 ( .A(n25741), .B(n25738), .Z(n25739) );
  IV U26224 ( .A(n25696), .Z(n25700) );
  XOR U26225 ( .A(n25696), .B(n25651), .Z(n25698) );
  XOR U26226 ( .A(n25742), .B(n25743), .Z(n25651) );
  AND U26227 ( .A(n598), .B(n25744), .Z(n25742) );
  XOR U26228 ( .A(n25745), .B(n25743), .Z(n25744) );
  NANDN U26229 ( .A(n25653), .B(n25655), .Z(n25696) );
  XOR U26230 ( .A(n25746), .B(n25747), .Z(n25655) );
  AND U26231 ( .A(n598), .B(n25748), .Z(n25746) );
  XOR U26232 ( .A(n25747), .B(n25749), .Z(n25748) );
  XNOR U26233 ( .A(n25750), .B(n25751), .Z(n598) );
  AND U26234 ( .A(n25752), .B(n25753), .Z(n25750) );
  XOR U26235 ( .A(n25751), .B(n25666), .Z(n25753) );
  XNOR U26236 ( .A(n25754), .B(n25755), .Z(n25666) );
  ANDN U26237 ( .B(n25756), .A(n25757), .Z(n25754) );
  XOR U26238 ( .A(n25755), .B(n25758), .Z(n25756) );
  XNOR U26239 ( .A(n25751), .B(n25668), .Z(n25752) );
  XOR U26240 ( .A(n25759), .B(n25760), .Z(n25668) );
  AND U26241 ( .A(n602), .B(n25761), .Z(n25759) );
  XOR U26242 ( .A(n25762), .B(n25760), .Z(n25761) );
  XNOR U26243 ( .A(n25763), .B(n25764), .Z(n25751) );
  AND U26244 ( .A(n25765), .B(n25766), .Z(n25763) );
  XNOR U26245 ( .A(n25764), .B(n25693), .Z(n25766) );
  XOR U26246 ( .A(n25757), .B(n25758), .Z(n25693) );
  XNOR U26247 ( .A(n25767), .B(n25768), .Z(n25758) );
  ANDN U26248 ( .B(n25769), .A(n25770), .Z(n25767) );
  XOR U26249 ( .A(n25771), .B(n25772), .Z(n25769) );
  XOR U26250 ( .A(n25773), .B(n25774), .Z(n25757) );
  XNOR U26251 ( .A(n25775), .B(n25776), .Z(n25774) );
  ANDN U26252 ( .B(n25777), .A(n25778), .Z(n25775) );
  XNOR U26253 ( .A(n25779), .B(n25780), .Z(n25777) );
  IV U26254 ( .A(n25755), .Z(n25773) );
  XOR U26255 ( .A(n25781), .B(n25782), .Z(n25755) );
  ANDN U26256 ( .B(n25783), .A(n25784), .Z(n25781) );
  XOR U26257 ( .A(n25782), .B(n25785), .Z(n25783) );
  XOR U26258 ( .A(n25764), .B(n25695), .Z(n25765) );
  XOR U26259 ( .A(n25786), .B(n25787), .Z(n25695) );
  AND U26260 ( .A(n602), .B(n25788), .Z(n25786) );
  XOR U26261 ( .A(n25789), .B(n25787), .Z(n25788) );
  XNOR U26262 ( .A(n25790), .B(n25791), .Z(n25764) );
  NAND U26263 ( .A(n25792), .B(n25793), .Z(n25791) );
  XOR U26264 ( .A(n25794), .B(n25743), .Z(n25793) );
  XOR U26265 ( .A(n25784), .B(n25785), .Z(n25743) );
  XOR U26266 ( .A(n25795), .B(n25772), .Z(n25785) );
  XOR U26267 ( .A(n25796), .B(n25797), .Z(n25772) );
  ANDN U26268 ( .B(n25798), .A(n25799), .Z(n25796) );
  XOR U26269 ( .A(n25797), .B(n25800), .Z(n25798) );
  IV U26270 ( .A(n25770), .Z(n25795) );
  XOR U26271 ( .A(n25768), .B(n25801), .Z(n25770) );
  XOR U26272 ( .A(n25802), .B(n25803), .Z(n25801) );
  ANDN U26273 ( .B(n25804), .A(n25805), .Z(n25802) );
  XOR U26274 ( .A(n25806), .B(n25803), .Z(n25804) );
  IV U26275 ( .A(n25771), .Z(n25768) );
  XOR U26276 ( .A(n25807), .B(n25808), .Z(n25771) );
  ANDN U26277 ( .B(n25809), .A(n25810), .Z(n25807) );
  XOR U26278 ( .A(n25808), .B(n25811), .Z(n25809) );
  XOR U26279 ( .A(n25812), .B(n25813), .Z(n25784) );
  XNOR U26280 ( .A(n25779), .B(n25814), .Z(n25813) );
  IV U26281 ( .A(n25782), .Z(n25814) );
  XOR U26282 ( .A(n25815), .B(n25816), .Z(n25782) );
  ANDN U26283 ( .B(n25817), .A(n25818), .Z(n25815) );
  XOR U26284 ( .A(n25816), .B(n25819), .Z(n25817) );
  XNOR U26285 ( .A(n25820), .B(n25821), .Z(n25779) );
  ANDN U26286 ( .B(n25822), .A(n25823), .Z(n25820) );
  XOR U26287 ( .A(n25821), .B(n25824), .Z(n25822) );
  IV U26288 ( .A(n25778), .Z(n25812) );
  XOR U26289 ( .A(n25776), .B(n25825), .Z(n25778) );
  XOR U26290 ( .A(n25826), .B(n25827), .Z(n25825) );
  ANDN U26291 ( .B(n25828), .A(n25829), .Z(n25826) );
  XOR U26292 ( .A(n25830), .B(n25827), .Z(n25828) );
  IV U26293 ( .A(n25780), .Z(n25776) );
  XOR U26294 ( .A(n25831), .B(n25832), .Z(n25780) );
  ANDN U26295 ( .B(n25833), .A(n25834), .Z(n25831) );
  XOR U26296 ( .A(n25835), .B(n25832), .Z(n25833) );
  IV U26297 ( .A(n25790), .Z(n25794) );
  XOR U26298 ( .A(n25790), .B(n25745), .Z(n25792) );
  XOR U26299 ( .A(n25836), .B(n25837), .Z(n25745) );
  AND U26300 ( .A(n602), .B(n25838), .Z(n25836) );
  XOR U26301 ( .A(n25839), .B(n25837), .Z(n25838) );
  NANDN U26302 ( .A(n25747), .B(n25749), .Z(n25790) );
  XOR U26303 ( .A(n25840), .B(n25841), .Z(n25749) );
  AND U26304 ( .A(n602), .B(n25842), .Z(n25840) );
  XOR U26305 ( .A(n25841), .B(n25843), .Z(n25842) );
  XNOR U26306 ( .A(n25844), .B(n25845), .Z(n602) );
  AND U26307 ( .A(n25846), .B(n25847), .Z(n25844) );
  XOR U26308 ( .A(n25845), .B(n25760), .Z(n25847) );
  XNOR U26309 ( .A(n25848), .B(n25849), .Z(n25760) );
  ANDN U26310 ( .B(n25850), .A(n25851), .Z(n25848) );
  XOR U26311 ( .A(n25849), .B(n25852), .Z(n25850) );
  XNOR U26312 ( .A(n25845), .B(n25762), .Z(n25846) );
  XOR U26313 ( .A(n25853), .B(n25854), .Z(n25762) );
  AND U26314 ( .A(n606), .B(n25855), .Z(n25853) );
  XOR U26315 ( .A(n25856), .B(n25854), .Z(n25855) );
  XNOR U26316 ( .A(n25857), .B(n25858), .Z(n25845) );
  AND U26317 ( .A(n25859), .B(n25860), .Z(n25857) );
  XNOR U26318 ( .A(n25858), .B(n25787), .Z(n25860) );
  XOR U26319 ( .A(n25851), .B(n25852), .Z(n25787) );
  XNOR U26320 ( .A(n25861), .B(n25862), .Z(n25852) );
  ANDN U26321 ( .B(n25863), .A(n25864), .Z(n25861) );
  XOR U26322 ( .A(n25865), .B(n25866), .Z(n25863) );
  XOR U26323 ( .A(n25867), .B(n25868), .Z(n25851) );
  XNOR U26324 ( .A(n25869), .B(n25870), .Z(n25868) );
  ANDN U26325 ( .B(n25871), .A(n25872), .Z(n25869) );
  XNOR U26326 ( .A(n25873), .B(n25874), .Z(n25871) );
  IV U26327 ( .A(n25849), .Z(n25867) );
  XOR U26328 ( .A(n25875), .B(n25876), .Z(n25849) );
  ANDN U26329 ( .B(n25877), .A(n25878), .Z(n25875) );
  XOR U26330 ( .A(n25876), .B(n25879), .Z(n25877) );
  XOR U26331 ( .A(n25858), .B(n25789), .Z(n25859) );
  XOR U26332 ( .A(n25880), .B(n25881), .Z(n25789) );
  AND U26333 ( .A(n606), .B(n25882), .Z(n25880) );
  XOR U26334 ( .A(n25883), .B(n25881), .Z(n25882) );
  XNOR U26335 ( .A(n25884), .B(n25885), .Z(n25858) );
  NAND U26336 ( .A(n25886), .B(n25887), .Z(n25885) );
  XOR U26337 ( .A(n25888), .B(n25837), .Z(n25887) );
  XOR U26338 ( .A(n25878), .B(n25879), .Z(n25837) );
  XOR U26339 ( .A(n25889), .B(n25866), .Z(n25879) );
  XOR U26340 ( .A(n25890), .B(n25891), .Z(n25866) );
  ANDN U26341 ( .B(n25892), .A(n25893), .Z(n25890) );
  XOR U26342 ( .A(n25891), .B(n25894), .Z(n25892) );
  IV U26343 ( .A(n25864), .Z(n25889) );
  XOR U26344 ( .A(n25862), .B(n25895), .Z(n25864) );
  XOR U26345 ( .A(n25896), .B(n25897), .Z(n25895) );
  ANDN U26346 ( .B(n25898), .A(n25899), .Z(n25896) );
  XOR U26347 ( .A(n25900), .B(n25897), .Z(n25898) );
  IV U26348 ( .A(n25865), .Z(n25862) );
  XOR U26349 ( .A(n25901), .B(n25902), .Z(n25865) );
  ANDN U26350 ( .B(n25903), .A(n25904), .Z(n25901) );
  XOR U26351 ( .A(n25902), .B(n25905), .Z(n25903) );
  XOR U26352 ( .A(n25906), .B(n25907), .Z(n25878) );
  XNOR U26353 ( .A(n25873), .B(n25908), .Z(n25907) );
  IV U26354 ( .A(n25876), .Z(n25908) );
  XOR U26355 ( .A(n25909), .B(n25910), .Z(n25876) );
  ANDN U26356 ( .B(n25911), .A(n25912), .Z(n25909) );
  XOR U26357 ( .A(n25910), .B(n25913), .Z(n25911) );
  XNOR U26358 ( .A(n25914), .B(n25915), .Z(n25873) );
  ANDN U26359 ( .B(n25916), .A(n25917), .Z(n25914) );
  XOR U26360 ( .A(n25915), .B(n25918), .Z(n25916) );
  IV U26361 ( .A(n25872), .Z(n25906) );
  XOR U26362 ( .A(n25870), .B(n25919), .Z(n25872) );
  XOR U26363 ( .A(n25920), .B(n25921), .Z(n25919) );
  ANDN U26364 ( .B(n25922), .A(n25923), .Z(n25920) );
  XOR U26365 ( .A(n25924), .B(n25921), .Z(n25922) );
  IV U26366 ( .A(n25874), .Z(n25870) );
  XOR U26367 ( .A(n25925), .B(n25926), .Z(n25874) );
  ANDN U26368 ( .B(n25927), .A(n25928), .Z(n25925) );
  XOR U26369 ( .A(n25929), .B(n25926), .Z(n25927) );
  IV U26370 ( .A(n25884), .Z(n25888) );
  XOR U26371 ( .A(n25884), .B(n25839), .Z(n25886) );
  XOR U26372 ( .A(n25930), .B(n25931), .Z(n25839) );
  AND U26373 ( .A(n606), .B(n25932), .Z(n25930) );
  XOR U26374 ( .A(n25933), .B(n25931), .Z(n25932) );
  NANDN U26375 ( .A(n25841), .B(n25843), .Z(n25884) );
  XOR U26376 ( .A(n25934), .B(n25935), .Z(n25843) );
  AND U26377 ( .A(n606), .B(n25936), .Z(n25934) );
  XOR U26378 ( .A(n25935), .B(n25937), .Z(n25936) );
  XNOR U26379 ( .A(n25938), .B(n25939), .Z(n606) );
  AND U26380 ( .A(n25940), .B(n25941), .Z(n25938) );
  XOR U26381 ( .A(n25939), .B(n25854), .Z(n25941) );
  XNOR U26382 ( .A(n25942), .B(n25943), .Z(n25854) );
  ANDN U26383 ( .B(n25944), .A(n25945), .Z(n25942) );
  XOR U26384 ( .A(n25943), .B(n25946), .Z(n25944) );
  XNOR U26385 ( .A(n25939), .B(n25856), .Z(n25940) );
  XOR U26386 ( .A(n25947), .B(n25948), .Z(n25856) );
  AND U26387 ( .A(n610), .B(n25949), .Z(n25947) );
  XOR U26388 ( .A(n25950), .B(n25948), .Z(n25949) );
  XNOR U26389 ( .A(n25951), .B(n25952), .Z(n25939) );
  AND U26390 ( .A(n25953), .B(n25954), .Z(n25951) );
  XNOR U26391 ( .A(n25952), .B(n25881), .Z(n25954) );
  XOR U26392 ( .A(n25945), .B(n25946), .Z(n25881) );
  XNOR U26393 ( .A(n25955), .B(n25956), .Z(n25946) );
  ANDN U26394 ( .B(n25957), .A(n25958), .Z(n25955) );
  XOR U26395 ( .A(n25959), .B(n25960), .Z(n25957) );
  XOR U26396 ( .A(n25961), .B(n25962), .Z(n25945) );
  XNOR U26397 ( .A(n25963), .B(n25964), .Z(n25962) );
  ANDN U26398 ( .B(n25965), .A(n25966), .Z(n25963) );
  XNOR U26399 ( .A(n25967), .B(n25968), .Z(n25965) );
  IV U26400 ( .A(n25943), .Z(n25961) );
  XOR U26401 ( .A(n25969), .B(n25970), .Z(n25943) );
  ANDN U26402 ( .B(n25971), .A(n25972), .Z(n25969) );
  XOR U26403 ( .A(n25970), .B(n25973), .Z(n25971) );
  XOR U26404 ( .A(n25952), .B(n25883), .Z(n25953) );
  XOR U26405 ( .A(n25974), .B(n25975), .Z(n25883) );
  AND U26406 ( .A(n610), .B(n25976), .Z(n25974) );
  XOR U26407 ( .A(n25977), .B(n25975), .Z(n25976) );
  XNOR U26408 ( .A(n25978), .B(n25979), .Z(n25952) );
  NAND U26409 ( .A(n25980), .B(n25981), .Z(n25979) );
  XOR U26410 ( .A(n25982), .B(n25931), .Z(n25981) );
  XOR U26411 ( .A(n25972), .B(n25973), .Z(n25931) );
  XOR U26412 ( .A(n25983), .B(n25960), .Z(n25973) );
  XOR U26413 ( .A(n25984), .B(n25985), .Z(n25960) );
  ANDN U26414 ( .B(n25986), .A(n25987), .Z(n25984) );
  XOR U26415 ( .A(n25985), .B(n25988), .Z(n25986) );
  IV U26416 ( .A(n25958), .Z(n25983) );
  XOR U26417 ( .A(n25956), .B(n25989), .Z(n25958) );
  XOR U26418 ( .A(n25990), .B(n25991), .Z(n25989) );
  ANDN U26419 ( .B(n25992), .A(n25993), .Z(n25990) );
  XOR U26420 ( .A(n25994), .B(n25991), .Z(n25992) );
  IV U26421 ( .A(n25959), .Z(n25956) );
  XOR U26422 ( .A(n25995), .B(n25996), .Z(n25959) );
  ANDN U26423 ( .B(n25997), .A(n25998), .Z(n25995) );
  XOR U26424 ( .A(n25996), .B(n25999), .Z(n25997) );
  XOR U26425 ( .A(n26000), .B(n26001), .Z(n25972) );
  XNOR U26426 ( .A(n25967), .B(n26002), .Z(n26001) );
  IV U26427 ( .A(n25970), .Z(n26002) );
  XOR U26428 ( .A(n26003), .B(n26004), .Z(n25970) );
  ANDN U26429 ( .B(n26005), .A(n26006), .Z(n26003) );
  XOR U26430 ( .A(n26004), .B(n26007), .Z(n26005) );
  XNOR U26431 ( .A(n26008), .B(n26009), .Z(n25967) );
  ANDN U26432 ( .B(n26010), .A(n26011), .Z(n26008) );
  XOR U26433 ( .A(n26009), .B(n26012), .Z(n26010) );
  IV U26434 ( .A(n25966), .Z(n26000) );
  XOR U26435 ( .A(n25964), .B(n26013), .Z(n25966) );
  XOR U26436 ( .A(n26014), .B(n26015), .Z(n26013) );
  ANDN U26437 ( .B(n26016), .A(n26017), .Z(n26014) );
  XOR U26438 ( .A(n26018), .B(n26015), .Z(n26016) );
  IV U26439 ( .A(n25968), .Z(n25964) );
  XOR U26440 ( .A(n26019), .B(n26020), .Z(n25968) );
  ANDN U26441 ( .B(n26021), .A(n26022), .Z(n26019) );
  XOR U26442 ( .A(n26023), .B(n26020), .Z(n26021) );
  IV U26443 ( .A(n25978), .Z(n25982) );
  XOR U26444 ( .A(n25978), .B(n25933), .Z(n25980) );
  XOR U26445 ( .A(n26024), .B(n26025), .Z(n25933) );
  AND U26446 ( .A(n610), .B(n26026), .Z(n26024) );
  XOR U26447 ( .A(n26027), .B(n26025), .Z(n26026) );
  NANDN U26448 ( .A(n25935), .B(n25937), .Z(n25978) );
  XOR U26449 ( .A(n26028), .B(n26029), .Z(n25937) );
  AND U26450 ( .A(n610), .B(n26030), .Z(n26028) );
  XOR U26451 ( .A(n26029), .B(n26031), .Z(n26030) );
  XNOR U26452 ( .A(n26032), .B(n26033), .Z(n610) );
  AND U26453 ( .A(n26034), .B(n26035), .Z(n26032) );
  XOR U26454 ( .A(n26033), .B(n25948), .Z(n26035) );
  XNOR U26455 ( .A(n26036), .B(n26037), .Z(n25948) );
  ANDN U26456 ( .B(n26038), .A(n26039), .Z(n26036) );
  XOR U26457 ( .A(n26037), .B(n26040), .Z(n26038) );
  XNOR U26458 ( .A(n26033), .B(n25950), .Z(n26034) );
  XOR U26459 ( .A(n26041), .B(n26042), .Z(n25950) );
  AND U26460 ( .A(n614), .B(n26043), .Z(n26041) );
  XOR U26461 ( .A(n26044), .B(n26042), .Z(n26043) );
  XNOR U26462 ( .A(n26045), .B(n26046), .Z(n26033) );
  AND U26463 ( .A(n26047), .B(n26048), .Z(n26045) );
  XNOR U26464 ( .A(n26046), .B(n25975), .Z(n26048) );
  XOR U26465 ( .A(n26039), .B(n26040), .Z(n25975) );
  XNOR U26466 ( .A(n26049), .B(n26050), .Z(n26040) );
  ANDN U26467 ( .B(n26051), .A(n26052), .Z(n26049) );
  XOR U26468 ( .A(n26053), .B(n26054), .Z(n26051) );
  XOR U26469 ( .A(n26055), .B(n26056), .Z(n26039) );
  XNOR U26470 ( .A(n26057), .B(n26058), .Z(n26056) );
  ANDN U26471 ( .B(n26059), .A(n26060), .Z(n26057) );
  XNOR U26472 ( .A(n26061), .B(n26062), .Z(n26059) );
  IV U26473 ( .A(n26037), .Z(n26055) );
  XOR U26474 ( .A(n26063), .B(n26064), .Z(n26037) );
  ANDN U26475 ( .B(n26065), .A(n26066), .Z(n26063) );
  XOR U26476 ( .A(n26064), .B(n26067), .Z(n26065) );
  XOR U26477 ( .A(n26046), .B(n25977), .Z(n26047) );
  XOR U26478 ( .A(n26068), .B(n26069), .Z(n25977) );
  AND U26479 ( .A(n614), .B(n26070), .Z(n26068) );
  XOR U26480 ( .A(n26071), .B(n26069), .Z(n26070) );
  XNOR U26481 ( .A(n26072), .B(n26073), .Z(n26046) );
  NAND U26482 ( .A(n26074), .B(n26075), .Z(n26073) );
  XOR U26483 ( .A(n26076), .B(n26025), .Z(n26075) );
  XOR U26484 ( .A(n26066), .B(n26067), .Z(n26025) );
  XOR U26485 ( .A(n26077), .B(n26054), .Z(n26067) );
  XOR U26486 ( .A(n26078), .B(n26079), .Z(n26054) );
  ANDN U26487 ( .B(n26080), .A(n26081), .Z(n26078) );
  XOR U26488 ( .A(n26079), .B(n26082), .Z(n26080) );
  IV U26489 ( .A(n26052), .Z(n26077) );
  XOR U26490 ( .A(n26050), .B(n26083), .Z(n26052) );
  XOR U26491 ( .A(n26084), .B(n26085), .Z(n26083) );
  ANDN U26492 ( .B(n26086), .A(n26087), .Z(n26084) );
  XOR U26493 ( .A(n26088), .B(n26085), .Z(n26086) );
  IV U26494 ( .A(n26053), .Z(n26050) );
  XOR U26495 ( .A(n26089), .B(n26090), .Z(n26053) );
  ANDN U26496 ( .B(n26091), .A(n26092), .Z(n26089) );
  XOR U26497 ( .A(n26090), .B(n26093), .Z(n26091) );
  XOR U26498 ( .A(n26094), .B(n26095), .Z(n26066) );
  XNOR U26499 ( .A(n26061), .B(n26096), .Z(n26095) );
  IV U26500 ( .A(n26064), .Z(n26096) );
  XOR U26501 ( .A(n26097), .B(n26098), .Z(n26064) );
  ANDN U26502 ( .B(n26099), .A(n26100), .Z(n26097) );
  XOR U26503 ( .A(n26098), .B(n26101), .Z(n26099) );
  XNOR U26504 ( .A(n26102), .B(n26103), .Z(n26061) );
  ANDN U26505 ( .B(n26104), .A(n26105), .Z(n26102) );
  XOR U26506 ( .A(n26103), .B(n26106), .Z(n26104) );
  IV U26507 ( .A(n26060), .Z(n26094) );
  XOR U26508 ( .A(n26058), .B(n26107), .Z(n26060) );
  XOR U26509 ( .A(n26108), .B(n26109), .Z(n26107) );
  ANDN U26510 ( .B(n26110), .A(n26111), .Z(n26108) );
  XOR U26511 ( .A(n26112), .B(n26109), .Z(n26110) );
  IV U26512 ( .A(n26062), .Z(n26058) );
  XOR U26513 ( .A(n26113), .B(n26114), .Z(n26062) );
  ANDN U26514 ( .B(n26115), .A(n26116), .Z(n26113) );
  XOR U26515 ( .A(n26117), .B(n26114), .Z(n26115) );
  IV U26516 ( .A(n26072), .Z(n26076) );
  XOR U26517 ( .A(n26072), .B(n26027), .Z(n26074) );
  XOR U26518 ( .A(n26118), .B(n26119), .Z(n26027) );
  AND U26519 ( .A(n614), .B(n26120), .Z(n26118) );
  XOR U26520 ( .A(n26121), .B(n26119), .Z(n26120) );
  NANDN U26521 ( .A(n26029), .B(n26031), .Z(n26072) );
  XOR U26522 ( .A(n26122), .B(n26123), .Z(n26031) );
  AND U26523 ( .A(n614), .B(n26124), .Z(n26122) );
  XOR U26524 ( .A(n26123), .B(n26125), .Z(n26124) );
  XNOR U26525 ( .A(n26126), .B(n26127), .Z(n614) );
  AND U26526 ( .A(n26128), .B(n26129), .Z(n26126) );
  XOR U26527 ( .A(n26127), .B(n26042), .Z(n26129) );
  XNOR U26528 ( .A(n26130), .B(n26131), .Z(n26042) );
  ANDN U26529 ( .B(n26132), .A(n26133), .Z(n26130) );
  XOR U26530 ( .A(n26131), .B(n26134), .Z(n26132) );
  XNOR U26531 ( .A(n26127), .B(n26044), .Z(n26128) );
  XOR U26532 ( .A(n26135), .B(n26136), .Z(n26044) );
  AND U26533 ( .A(n618), .B(n26137), .Z(n26135) );
  XOR U26534 ( .A(n26138), .B(n26136), .Z(n26137) );
  XNOR U26535 ( .A(n26139), .B(n26140), .Z(n26127) );
  AND U26536 ( .A(n26141), .B(n26142), .Z(n26139) );
  XNOR U26537 ( .A(n26140), .B(n26069), .Z(n26142) );
  XOR U26538 ( .A(n26133), .B(n26134), .Z(n26069) );
  XNOR U26539 ( .A(n26143), .B(n26144), .Z(n26134) );
  ANDN U26540 ( .B(n26145), .A(n26146), .Z(n26143) );
  XOR U26541 ( .A(n26147), .B(n26148), .Z(n26145) );
  XOR U26542 ( .A(n26149), .B(n26150), .Z(n26133) );
  XNOR U26543 ( .A(n26151), .B(n26152), .Z(n26150) );
  ANDN U26544 ( .B(n26153), .A(n26154), .Z(n26151) );
  XNOR U26545 ( .A(n26155), .B(n26156), .Z(n26153) );
  IV U26546 ( .A(n26131), .Z(n26149) );
  XOR U26547 ( .A(n26157), .B(n26158), .Z(n26131) );
  ANDN U26548 ( .B(n26159), .A(n26160), .Z(n26157) );
  XOR U26549 ( .A(n26158), .B(n26161), .Z(n26159) );
  XOR U26550 ( .A(n26140), .B(n26071), .Z(n26141) );
  XOR U26551 ( .A(n26162), .B(n26163), .Z(n26071) );
  AND U26552 ( .A(n618), .B(n26164), .Z(n26162) );
  XOR U26553 ( .A(n26165), .B(n26163), .Z(n26164) );
  XNOR U26554 ( .A(n26166), .B(n26167), .Z(n26140) );
  NAND U26555 ( .A(n26168), .B(n26169), .Z(n26167) );
  XOR U26556 ( .A(n26170), .B(n26119), .Z(n26169) );
  XOR U26557 ( .A(n26160), .B(n26161), .Z(n26119) );
  XOR U26558 ( .A(n26171), .B(n26148), .Z(n26161) );
  XOR U26559 ( .A(n26172), .B(n26173), .Z(n26148) );
  ANDN U26560 ( .B(n26174), .A(n26175), .Z(n26172) );
  XOR U26561 ( .A(n26173), .B(n26176), .Z(n26174) );
  IV U26562 ( .A(n26146), .Z(n26171) );
  XOR U26563 ( .A(n26144), .B(n26177), .Z(n26146) );
  XOR U26564 ( .A(n26178), .B(n26179), .Z(n26177) );
  ANDN U26565 ( .B(n26180), .A(n26181), .Z(n26178) );
  XOR U26566 ( .A(n26182), .B(n26179), .Z(n26180) );
  IV U26567 ( .A(n26147), .Z(n26144) );
  XOR U26568 ( .A(n26183), .B(n26184), .Z(n26147) );
  ANDN U26569 ( .B(n26185), .A(n26186), .Z(n26183) );
  XOR U26570 ( .A(n26184), .B(n26187), .Z(n26185) );
  XOR U26571 ( .A(n26188), .B(n26189), .Z(n26160) );
  XNOR U26572 ( .A(n26155), .B(n26190), .Z(n26189) );
  IV U26573 ( .A(n26158), .Z(n26190) );
  XOR U26574 ( .A(n26191), .B(n26192), .Z(n26158) );
  ANDN U26575 ( .B(n26193), .A(n26194), .Z(n26191) );
  XOR U26576 ( .A(n26192), .B(n26195), .Z(n26193) );
  XNOR U26577 ( .A(n26196), .B(n26197), .Z(n26155) );
  ANDN U26578 ( .B(n26198), .A(n26199), .Z(n26196) );
  XOR U26579 ( .A(n26197), .B(n26200), .Z(n26198) );
  IV U26580 ( .A(n26154), .Z(n26188) );
  XOR U26581 ( .A(n26152), .B(n26201), .Z(n26154) );
  XOR U26582 ( .A(n26202), .B(n26203), .Z(n26201) );
  ANDN U26583 ( .B(n26204), .A(n26205), .Z(n26202) );
  XOR U26584 ( .A(n26206), .B(n26203), .Z(n26204) );
  IV U26585 ( .A(n26156), .Z(n26152) );
  XOR U26586 ( .A(n26207), .B(n26208), .Z(n26156) );
  ANDN U26587 ( .B(n26209), .A(n26210), .Z(n26207) );
  XOR U26588 ( .A(n26211), .B(n26208), .Z(n26209) );
  IV U26589 ( .A(n26166), .Z(n26170) );
  XOR U26590 ( .A(n26166), .B(n26121), .Z(n26168) );
  XOR U26591 ( .A(n26212), .B(n26213), .Z(n26121) );
  AND U26592 ( .A(n618), .B(n26214), .Z(n26212) );
  XOR U26593 ( .A(n26215), .B(n26213), .Z(n26214) );
  NANDN U26594 ( .A(n26123), .B(n26125), .Z(n26166) );
  XOR U26595 ( .A(n26216), .B(n26217), .Z(n26125) );
  AND U26596 ( .A(n618), .B(n26218), .Z(n26216) );
  XOR U26597 ( .A(n26217), .B(n26219), .Z(n26218) );
  XNOR U26598 ( .A(n26220), .B(n26221), .Z(n618) );
  AND U26599 ( .A(n26222), .B(n26223), .Z(n26220) );
  XOR U26600 ( .A(n26221), .B(n26136), .Z(n26223) );
  XNOR U26601 ( .A(n26224), .B(n26225), .Z(n26136) );
  ANDN U26602 ( .B(n26226), .A(n26227), .Z(n26224) );
  XOR U26603 ( .A(n26225), .B(n26228), .Z(n26226) );
  XNOR U26604 ( .A(n26221), .B(n26138), .Z(n26222) );
  XOR U26605 ( .A(n26229), .B(n26230), .Z(n26138) );
  AND U26606 ( .A(n622), .B(n26231), .Z(n26229) );
  XOR U26607 ( .A(n26232), .B(n26230), .Z(n26231) );
  XNOR U26608 ( .A(n26233), .B(n26234), .Z(n26221) );
  AND U26609 ( .A(n26235), .B(n26236), .Z(n26233) );
  XNOR U26610 ( .A(n26234), .B(n26163), .Z(n26236) );
  XOR U26611 ( .A(n26227), .B(n26228), .Z(n26163) );
  XNOR U26612 ( .A(n26237), .B(n26238), .Z(n26228) );
  ANDN U26613 ( .B(n26239), .A(n26240), .Z(n26237) );
  XOR U26614 ( .A(n26241), .B(n26242), .Z(n26239) );
  XOR U26615 ( .A(n26243), .B(n26244), .Z(n26227) );
  XNOR U26616 ( .A(n26245), .B(n26246), .Z(n26244) );
  ANDN U26617 ( .B(n26247), .A(n26248), .Z(n26245) );
  XNOR U26618 ( .A(n26249), .B(n26250), .Z(n26247) );
  IV U26619 ( .A(n26225), .Z(n26243) );
  XOR U26620 ( .A(n26251), .B(n26252), .Z(n26225) );
  ANDN U26621 ( .B(n26253), .A(n26254), .Z(n26251) );
  XOR U26622 ( .A(n26252), .B(n26255), .Z(n26253) );
  XOR U26623 ( .A(n26234), .B(n26165), .Z(n26235) );
  XOR U26624 ( .A(n26256), .B(n26257), .Z(n26165) );
  AND U26625 ( .A(n622), .B(n26258), .Z(n26256) );
  XOR U26626 ( .A(n26259), .B(n26257), .Z(n26258) );
  XNOR U26627 ( .A(n26260), .B(n26261), .Z(n26234) );
  NAND U26628 ( .A(n26262), .B(n26263), .Z(n26261) );
  XOR U26629 ( .A(n26264), .B(n26213), .Z(n26263) );
  XOR U26630 ( .A(n26254), .B(n26255), .Z(n26213) );
  XOR U26631 ( .A(n26265), .B(n26242), .Z(n26255) );
  XOR U26632 ( .A(n26266), .B(n26267), .Z(n26242) );
  ANDN U26633 ( .B(n26268), .A(n26269), .Z(n26266) );
  XOR U26634 ( .A(n26267), .B(n26270), .Z(n26268) );
  IV U26635 ( .A(n26240), .Z(n26265) );
  XOR U26636 ( .A(n26238), .B(n26271), .Z(n26240) );
  XOR U26637 ( .A(n26272), .B(n26273), .Z(n26271) );
  ANDN U26638 ( .B(n26274), .A(n26275), .Z(n26272) );
  XOR U26639 ( .A(n26276), .B(n26273), .Z(n26274) );
  IV U26640 ( .A(n26241), .Z(n26238) );
  XOR U26641 ( .A(n26277), .B(n26278), .Z(n26241) );
  ANDN U26642 ( .B(n26279), .A(n26280), .Z(n26277) );
  XOR U26643 ( .A(n26278), .B(n26281), .Z(n26279) );
  XOR U26644 ( .A(n26282), .B(n26283), .Z(n26254) );
  XNOR U26645 ( .A(n26249), .B(n26284), .Z(n26283) );
  IV U26646 ( .A(n26252), .Z(n26284) );
  XOR U26647 ( .A(n26285), .B(n26286), .Z(n26252) );
  ANDN U26648 ( .B(n26287), .A(n26288), .Z(n26285) );
  XOR U26649 ( .A(n26286), .B(n26289), .Z(n26287) );
  XNOR U26650 ( .A(n26290), .B(n26291), .Z(n26249) );
  ANDN U26651 ( .B(n26292), .A(n26293), .Z(n26290) );
  XOR U26652 ( .A(n26291), .B(n26294), .Z(n26292) );
  IV U26653 ( .A(n26248), .Z(n26282) );
  XOR U26654 ( .A(n26246), .B(n26295), .Z(n26248) );
  XOR U26655 ( .A(n26296), .B(n26297), .Z(n26295) );
  ANDN U26656 ( .B(n26298), .A(n26299), .Z(n26296) );
  XOR U26657 ( .A(n26300), .B(n26297), .Z(n26298) );
  IV U26658 ( .A(n26250), .Z(n26246) );
  XOR U26659 ( .A(n26301), .B(n26302), .Z(n26250) );
  ANDN U26660 ( .B(n26303), .A(n26304), .Z(n26301) );
  XOR U26661 ( .A(n26305), .B(n26302), .Z(n26303) );
  IV U26662 ( .A(n26260), .Z(n26264) );
  XOR U26663 ( .A(n26260), .B(n26215), .Z(n26262) );
  XOR U26664 ( .A(n26306), .B(n26307), .Z(n26215) );
  AND U26665 ( .A(n622), .B(n26308), .Z(n26306) );
  XOR U26666 ( .A(n26309), .B(n26307), .Z(n26308) );
  NANDN U26667 ( .A(n26217), .B(n26219), .Z(n26260) );
  XOR U26668 ( .A(n26310), .B(n26311), .Z(n26219) );
  AND U26669 ( .A(n622), .B(n26312), .Z(n26310) );
  XOR U26670 ( .A(n26311), .B(n26313), .Z(n26312) );
  XNOR U26671 ( .A(n26314), .B(n26315), .Z(n622) );
  AND U26672 ( .A(n26316), .B(n26317), .Z(n26314) );
  XOR U26673 ( .A(n26315), .B(n26230), .Z(n26317) );
  XNOR U26674 ( .A(n26318), .B(n26319), .Z(n26230) );
  ANDN U26675 ( .B(n26320), .A(n26321), .Z(n26318) );
  XOR U26676 ( .A(n26319), .B(n26322), .Z(n26320) );
  XNOR U26677 ( .A(n26315), .B(n26232), .Z(n26316) );
  XOR U26678 ( .A(n26323), .B(n26324), .Z(n26232) );
  AND U26679 ( .A(n626), .B(n26325), .Z(n26323) );
  XOR U26680 ( .A(n26326), .B(n26324), .Z(n26325) );
  XNOR U26681 ( .A(n26327), .B(n26328), .Z(n26315) );
  AND U26682 ( .A(n26329), .B(n26330), .Z(n26327) );
  XNOR U26683 ( .A(n26328), .B(n26257), .Z(n26330) );
  XOR U26684 ( .A(n26321), .B(n26322), .Z(n26257) );
  XNOR U26685 ( .A(n26331), .B(n26332), .Z(n26322) );
  ANDN U26686 ( .B(n26333), .A(n26334), .Z(n26331) );
  XOR U26687 ( .A(n26335), .B(n26336), .Z(n26333) );
  XOR U26688 ( .A(n26337), .B(n26338), .Z(n26321) );
  XNOR U26689 ( .A(n26339), .B(n26340), .Z(n26338) );
  ANDN U26690 ( .B(n26341), .A(n26342), .Z(n26339) );
  XNOR U26691 ( .A(n26343), .B(n26344), .Z(n26341) );
  IV U26692 ( .A(n26319), .Z(n26337) );
  XOR U26693 ( .A(n26345), .B(n26346), .Z(n26319) );
  ANDN U26694 ( .B(n26347), .A(n26348), .Z(n26345) );
  XOR U26695 ( .A(n26346), .B(n26349), .Z(n26347) );
  XOR U26696 ( .A(n26328), .B(n26259), .Z(n26329) );
  XOR U26697 ( .A(n26350), .B(n26351), .Z(n26259) );
  AND U26698 ( .A(n626), .B(n26352), .Z(n26350) );
  XOR U26699 ( .A(n26353), .B(n26351), .Z(n26352) );
  XNOR U26700 ( .A(n26354), .B(n26355), .Z(n26328) );
  NAND U26701 ( .A(n26356), .B(n26357), .Z(n26355) );
  XOR U26702 ( .A(n26358), .B(n26307), .Z(n26357) );
  XOR U26703 ( .A(n26348), .B(n26349), .Z(n26307) );
  XOR U26704 ( .A(n26359), .B(n26336), .Z(n26349) );
  XOR U26705 ( .A(n26360), .B(n26361), .Z(n26336) );
  ANDN U26706 ( .B(n26362), .A(n26363), .Z(n26360) );
  XOR U26707 ( .A(n26361), .B(n26364), .Z(n26362) );
  IV U26708 ( .A(n26334), .Z(n26359) );
  XOR U26709 ( .A(n26332), .B(n26365), .Z(n26334) );
  XOR U26710 ( .A(n26366), .B(n26367), .Z(n26365) );
  ANDN U26711 ( .B(n26368), .A(n26369), .Z(n26366) );
  XOR U26712 ( .A(n26370), .B(n26367), .Z(n26368) );
  IV U26713 ( .A(n26335), .Z(n26332) );
  XOR U26714 ( .A(n26371), .B(n26372), .Z(n26335) );
  ANDN U26715 ( .B(n26373), .A(n26374), .Z(n26371) );
  XOR U26716 ( .A(n26372), .B(n26375), .Z(n26373) );
  XOR U26717 ( .A(n26376), .B(n26377), .Z(n26348) );
  XNOR U26718 ( .A(n26343), .B(n26378), .Z(n26377) );
  IV U26719 ( .A(n26346), .Z(n26378) );
  XOR U26720 ( .A(n26379), .B(n26380), .Z(n26346) );
  ANDN U26721 ( .B(n26381), .A(n26382), .Z(n26379) );
  XOR U26722 ( .A(n26380), .B(n26383), .Z(n26381) );
  XNOR U26723 ( .A(n26384), .B(n26385), .Z(n26343) );
  ANDN U26724 ( .B(n26386), .A(n26387), .Z(n26384) );
  XOR U26725 ( .A(n26385), .B(n26388), .Z(n26386) );
  IV U26726 ( .A(n26342), .Z(n26376) );
  XOR U26727 ( .A(n26340), .B(n26389), .Z(n26342) );
  XOR U26728 ( .A(n26390), .B(n26391), .Z(n26389) );
  ANDN U26729 ( .B(n26392), .A(n26393), .Z(n26390) );
  XOR U26730 ( .A(n26394), .B(n26391), .Z(n26392) );
  IV U26731 ( .A(n26344), .Z(n26340) );
  XOR U26732 ( .A(n26395), .B(n26396), .Z(n26344) );
  ANDN U26733 ( .B(n26397), .A(n26398), .Z(n26395) );
  XOR U26734 ( .A(n26399), .B(n26396), .Z(n26397) );
  IV U26735 ( .A(n26354), .Z(n26358) );
  XOR U26736 ( .A(n26354), .B(n26309), .Z(n26356) );
  XOR U26737 ( .A(n26400), .B(n26401), .Z(n26309) );
  AND U26738 ( .A(n626), .B(n26402), .Z(n26400) );
  XOR U26739 ( .A(n26403), .B(n26401), .Z(n26402) );
  NANDN U26740 ( .A(n26311), .B(n26313), .Z(n26354) );
  XOR U26741 ( .A(n26404), .B(n26405), .Z(n26313) );
  AND U26742 ( .A(n626), .B(n26406), .Z(n26404) );
  XOR U26743 ( .A(n26405), .B(n26407), .Z(n26406) );
  XNOR U26744 ( .A(n26408), .B(n26409), .Z(n626) );
  AND U26745 ( .A(n26410), .B(n26411), .Z(n26408) );
  XOR U26746 ( .A(n26409), .B(n26324), .Z(n26411) );
  XNOR U26747 ( .A(n26412), .B(n26413), .Z(n26324) );
  ANDN U26748 ( .B(n26414), .A(n26415), .Z(n26412) );
  XOR U26749 ( .A(n26413), .B(n26416), .Z(n26414) );
  XNOR U26750 ( .A(n26409), .B(n26326), .Z(n26410) );
  XOR U26751 ( .A(n26417), .B(n26418), .Z(n26326) );
  AND U26752 ( .A(n630), .B(n26419), .Z(n26417) );
  XOR U26753 ( .A(n26420), .B(n26418), .Z(n26419) );
  XNOR U26754 ( .A(n26421), .B(n26422), .Z(n26409) );
  AND U26755 ( .A(n26423), .B(n26424), .Z(n26421) );
  XNOR U26756 ( .A(n26422), .B(n26351), .Z(n26424) );
  XOR U26757 ( .A(n26415), .B(n26416), .Z(n26351) );
  XNOR U26758 ( .A(n26425), .B(n26426), .Z(n26416) );
  ANDN U26759 ( .B(n26427), .A(n26428), .Z(n26425) );
  XOR U26760 ( .A(n26429), .B(n26430), .Z(n26427) );
  XOR U26761 ( .A(n26431), .B(n26432), .Z(n26415) );
  XNOR U26762 ( .A(n26433), .B(n26434), .Z(n26432) );
  ANDN U26763 ( .B(n26435), .A(n26436), .Z(n26433) );
  XNOR U26764 ( .A(n26437), .B(n26438), .Z(n26435) );
  IV U26765 ( .A(n26413), .Z(n26431) );
  XOR U26766 ( .A(n26439), .B(n26440), .Z(n26413) );
  ANDN U26767 ( .B(n26441), .A(n26442), .Z(n26439) );
  XOR U26768 ( .A(n26440), .B(n26443), .Z(n26441) );
  XOR U26769 ( .A(n26422), .B(n26353), .Z(n26423) );
  XOR U26770 ( .A(n26444), .B(n26445), .Z(n26353) );
  AND U26771 ( .A(n630), .B(n26446), .Z(n26444) );
  XOR U26772 ( .A(n26447), .B(n26445), .Z(n26446) );
  XNOR U26773 ( .A(n26448), .B(n26449), .Z(n26422) );
  NAND U26774 ( .A(n26450), .B(n26451), .Z(n26449) );
  XOR U26775 ( .A(n26452), .B(n26401), .Z(n26451) );
  XOR U26776 ( .A(n26442), .B(n26443), .Z(n26401) );
  XOR U26777 ( .A(n26453), .B(n26430), .Z(n26443) );
  XOR U26778 ( .A(n26454), .B(n26455), .Z(n26430) );
  ANDN U26779 ( .B(n26456), .A(n26457), .Z(n26454) );
  XOR U26780 ( .A(n26455), .B(n26458), .Z(n26456) );
  IV U26781 ( .A(n26428), .Z(n26453) );
  XOR U26782 ( .A(n26426), .B(n26459), .Z(n26428) );
  XOR U26783 ( .A(n26460), .B(n26461), .Z(n26459) );
  ANDN U26784 ( .B(n26462), .A(n26463), .Z(n26460) );
  XOR U26785 ( .A(n26464), .B(n26461), .Z(n26462) );
  IV U26786 ( .A(n26429), .Z(n26426) );
  XOR U26787 ( .A(n26465), .B(n26466), .Z(n26429) );
  ANDN U26788 ( .B(n26467), .A(n26468), .Z(n26465) );
  XOR U26789 ( .A(n26466), .B(n26469), .Z(n26467) );
  XOR U26790 ( .A(n26470), .B(n26471), .Z(n26442) );
  XNOR U26791 ( .A(n26437), .B(n26472), .Z(n26471) );
  IV U26792 ( .A(n26440), .Z(n26472) );
  XOR U26793 ( .A(n26473), .B(n26474), .Z(n26440) );
  ANDN U26794 ( .B(n26475), .A(n26476), .Z(n26473) );
  XOR U26795 ( .A(n26474), .B(n26477), .Z(n26475) );
  XNOR U26796 ( .A(n26478), .B(n26479), .Z(n26437) );
  ANDN U26797 ( .B(n26480), .A(n26481), .Z(n26478) );
  XOR U26798 ( .A(n26479), .B(n26482), .Z(n26480) );
  IV U26799 ( .A(n26436), .Z(n26470) );
  XOR U26800 ( .A(n26434), .B(n26483), .Z(n26436) );
  XOR U26801 ( .A(n26484), .B(n26485), .Z(n26483) );
  ANDN U26802 ( .B(n26486), .A(n26487), .Z(n26484) );
  XOR U26803 ( .A(n26488), .B(n26485), .Z(n26486) );
  IV U26804 ( .A(n26438), .Z(n26434) );
  XOR U26805 ( .A(n26489), .B(n26490), .Z(n26438) );
  ANDN U26806 ( .B(n26491), .A(n26492), .Z(n26489) );
  XOR U26807 ( .A(n26493), .B(n26490), .Z(n26491) );
  IV U26808 ( .A(n26448), .Z(n26452) );
  XOR U26809 ( .A(n26448), .B(n26403), .Z(n26450) );
  XOR U26810 ( .A(n26494), .B(n26495), .Z(n26403) );
  AND U26811 ( .A(n630), .B(n26496), .Z(n26494) );
  XOR U26812 ( .A(n26497), .B(n26495), .Z(n26496) );
  NANDN U26813 ( .A(n26405), .B(n26407), .Z(n26448) );
  XOR U26814 ( .A(n26498), .B(n26499), .Z(n26407) );
  AND U26815 ( .A(n630), .B(n26500), .Z(n26498) );
  XOR U26816 ( .A(n26499), .B(n26501), .Z(n26500) );
  XNOR U26817 ( .A(n26502), .B(n26503), .Z(n630) );
  AND U26818 ( .A(n26504), .B(n26505), .Z(n26502) );
  XOR U26819 ( .A(n26503), .B(n26418), .Z(n26505) );
  XNOR U26820 ( .A(n26506), .B(n26507), .Z(n26418) );
  ANDN U26821 ( .B(n26508), .A(n26509), .Z(n26506) );
  XOR U26822 ( .A(n26507), .B(n26510), .Z(n26508) );
  XNOR U26823 ( .A(n26503), .B(n26420), .Z(n26504) );
  XOR U26824 ( .A(n26511), .B(n26512), .Z(n26420) );
  AND U26825 ( .A(n634), .B(n26513), .Z(n26511) );
  XOR U26826 ( .A(n26514), .B(n26512), .Z(n26513) );
  XNOR U26827 ( .A(n26515), .B(n26516), .Z(n26503) );
  AND U26828 ( .A(n26517), .B(n26518), .Z(n26515) );
  XNOR U26829 ( .A(n26516), .B(n26445), .Z(n26518) );
  XOR U26830 ( .A(n26509), .B(n26510), .Z(n26445) );
  XNOR U26831 ( .A(n26519), .B(n26520), .Z(n26510) );
  ANDN U26832 ( .B(n26521), .A(n26522), .Z(n26519) );
  XOR U26833 ( .A(n26523), .B(n26524), .Z(n26521) );
  XOR U26834 ( .A(n26525), .B(n26526), .Z(n26509) );
  XNOR U26835 ( .A(n26527), .B(n26528), .Z(n26526) );
  ANDN U26836 ( .B(n26529), .A(n26530), .Z(n26527) );
  XNOR U26837 ( .A(n26531), .B(n26532), .Z(n26529) );
  IV U26838 ( .A(n26507), .Z(n26525) );
  XOR U26839 ( .A(n26533), .B(n26534), .Z(n26507) );
  ANDN U26840 ( .B(n26535), .A(n26536), .Z(n26533) );
  XOR U26841 ( .A(n26534), .B(n26537), .Z(n26535) );
  XOR U26842 ( .A(n26516), .B(n26447), .Z(n26517) );
  XOR U26843 ( .A(n26538), .B(n26539), .Z(n26447) );
  AND U26844 ( .A(n634), .B(n26540), .Z(n26538) );
  XOR U26845 ( .A(n26541), .B(n26539), .Z(n26540) );
  XNOR U26846 ( .A(n26542), .B(n26543), .Z(n26516) );
  NAND U26847 ( .A(n26544), .B(n26545), .Z(n26543) );
  XOR U26848 ( .A(n26546), .B(n26495), .Z(n26545) );
  XOR U26849 ( .A(n26536), .B(n26537), .Z(n26495) );
  XOR U26850 ( .A(n26547), .B(n26524), .Z(n26537) );
  XOR U26851 ( .A(n26548), .B(n26549), .Z(n26524) );
  ANDN U26852 ( .B(n26550), .A(n26551), .Z(n26548) );
  XOR U26853 ( .A(n26549), .B(n26552), .Z(n26550) );
  IV U26854 ( .A(n26522), .Z(n26547) );
  XOR U26855 ( .A(n26520), .B(n26553), .Z(n26522) );
  XOR U26856 ( .A(n26554), .B(n26555), .Z(n26553) );
  ANDN U26857 ( .B(n26556), .A(n26557), .Z(n26554) );
  XOR U26858 ( .A(n26558), .B(n26555), .Z(n26556) );
  IV U26859 ( .A(n26523), .Z(n26520) );
  XOR U26860 ( .A(n26559), .B(n26560), .Z(n26523) );
  ANDN U26861 ( .B(n26561), .A(n26562), .Z(n26559) );
  XOR U26862 ( .A(n26560), .B(n26563), .Z(n26561) );
  XOR U26863 ( .A(n26564), .B(n26565), .Z(n26536) );
  XNOR U26864 ( .A(n26531), .B(n26566), .Z(n26565) );
  IV U26865 ( .A(n26534), .Z(n26566) );
  XOR U26866 ( .A(n26567), .B(n26568), .Z(n26534) );
  ANDN U26867 ( .B(n26569), .A(n26570), .Z(n26567) );
  XOR U26868 ( .A(n26568), .B(n26571), .Z(n26569) );
  XNOR U26869 ( .A(n26572), .B(n26573), .Z(n26531) );
  ANDN U26870 ( .B(n26574), .A(n26575), .Z(n26572) );
  XOR U26871 ( .A(n26573), .B(n26576), .Z(n26574) );
  IV U26872 ( .A(n26530), .Z(n26564) );
  XOR U26873 ( .A(n26528), .B(n26577), .Z(n26530) );
  XOR U26874 ( .A(n26578), .B(n26579), .Z(n26577) );
  ANDN U26875 ( .B(n26580), .A(n26581), .Z(n26578) );
  XOR U26876 ( .A(n26582), .B(n26579), .Z(n26580) );
  IV U26877 ( .A(n26532), .Z(n26528) );
  XOR U26878 ( .A(n26583), .B(n26584), .Z(n26532) );
  ANDN U26879 ( .B(n26585), .A(n26586), .Z(n26583) );
  XOR U26880 ( .A(n26587), .B(n26584), .Z(n26585) );
  IV U26881 ( .A(n26542), .Z(n26546) );
  XOR U26882 ( .A(n26542), .B(n26497), .Z(n26544) );
  XOR U26883 ( .A(n26588), .B(n26589), .Z(n26497) );
  AND U26884 ( .A(n634), .B(n26590), .Z(n26588) );
  XOR U26885 ( .A(n26591), .B(n26589), .Z(n26590) );
  NANDN U26886 ( .A(n26499), .B(n26501), .Z(n26542) );
  XOR U26887 ( .A(n26592), .B(n26593), .Z(n26501) );
  AND U26888 ( .A(n634), .B(n26594), .Z(n26592) );
  XOR U26889 ( .A(n26593), .B(n26595), .Z(n26594) );
  XNOR U26890 ( .A(n26596), .B(n26597), .Z(n634) );
  AND U26891 ( .A(n26598), .B(n26599), .Z(n26596) );
  XOR U26892 ( .A(n26597), .B(n26512), .Z(n26599) );
  XNOR U26893 ( .A(n26600), .B(n26601), .Z(n26512) );
  ANDN U26894 ( .B(n26602), .A(n26603), .Z(n26600) );
  XOR U26895 ( .A(n26601), .B(n26604), .Z(n26602) );
  XNOR U26896 ( .A(n26597), .B(n26514), .Z(n26598) );
  XOR U26897 ( .A(n26605), .B(n26606), .Z(n26514) );
  AND U26898 ( .A(n638), .B(n26607), .Z(n26605) );
  XOR U26899 ( .A(n26608), .B(n26606), .Z(n26607) );
  XNOR U26900 ( .A(n26609), .B(n26610), .Z(n26597) );
  AND U26901 ( .A(n26611), .B(n26612), .Z(n26609) );
  XNOR U26902 ( .A(n26610), .B(n26539), .Z(n26612) );
  XOR U26903 ( .A(n26603), .B(n26604), .Z(n26539) );
  XNOR U26904 ( .A(n26613), .B(n26614), .Z(n26604) );
  ANDN U26905 ( .B(n26615), .A(n26616), .Z(n26613) );
  XOR U26906 ( .A(n26617), .B(n26618), .Z(n26615) );
  XOR U26907 ( .A(n26619), .B(n26620), .Z(n26603) );
  XNOR U26908 ( .A(n26621), .B(n26622), .Z(n26620) );
  ANDN U26909 ( .B(n26623), .A(n26624), .Z(n26621) );
  XNOR U26910 ( .A(n26625), .B(n26626), .Z(n26623) );
  IV U26911 ( .A(n26601), .Z(n26619) );
  XOR U26912 ( .A(n26627), .B(n26628), .Z(n26601) );
  ANDN U26913 ( .B(n26629), .A(n26630), .Z(n26627) );
  XOR U26914 ( .A(n26628), .B(n26631), .Z(n26629) );
  XOR U26915 ( .A(n26610), .B(n26541), .Z(n26611) );
  XOR U26916 ( .A(n26632), .B(n26633), .Z(n26541) );
  AND U26917 ( .A(n638), .B(n26634), .Z(n26632) );
  XOR U26918 ( .A(n26635), .B(n26633), .Z(n26634) );
  XNOR U26919 ( .A(n26636), .B(n26637), .Z(n26610) );
  NAND U26920 ( .A(n26638), .B(n26639), .Z(n26637) );
  XOR U26921 ( .A(n26640), .B(n26589), .Z(n26639) );
  XOR U26922 ( .A(n26630), .B(n26631), .Z(n26589) );
  XOR U26923 ( .A(n26641), .B(n26618), .Z(n26631) );
  XOR U26924 ( .A(n26642), .B(n26643), .Z(n26618) );
  ANDN U26925 ( .B(n26644), .A(n26645), .Z(n26642) );
  XOR U26926 ( .A(n26643), .B(n26646), .Z(n26644) );
  IV U26927 ( .A(n26616), .Z(n26641) );
  XOR U26928 ( .A(n26614), .B(n26647), .Z(n26616) );
  XOR U26929 ( .A(n26648), .B(n26649), .Z(n26647) );
  ANDN U26930 ( .B(n26650), .A(n26651), .Z(n26648) );
  XOR U26931 ( .A(n26652), .B(n26649), .Z(n26650) );
  IV U26932 ( .A(n26617), .Z(n26614) );
  XOR U26933 ( .A(n26653), .B(n26654), .Z(n26617) );
  ANDN U26934 ( .B(n26655), .A(n26656), .Z(n26653) );
  XOR U26935 ( .A(n26654), .B(n26657), .Z(n26655) );
  XOR U26936 ( .A(n26658), .B(n26659), .Z(n26630) );
  XNOR U26937 ( .A(n26625), .B(n26660), .Z(n26659) );
  IV U26938 ( .A(n26628), .Z(n26660) );
  XOR U26939 ( .A(n26661), .B(n26662), .Z(n26628) );
  ANDN U26940 ( .B(n26663), .A(n26664), .Z(n26661) );
  XOR U26941 ( .A(n26662), .B(n26665), .Z(n26663) );
  XNOR U26942 ( .A(n26666), .B(n26667), .Z(n26625) );
  ANDN U26943 ( .B(n26668), .A(n26669), .Z(n26666) );
  XOR U26944 ( .A(n26667), .B(n26670), .Z(n26668) );
  IV U26945 ( .A(n26624), .Z(n26658) );
  XOR U26946 ( .A(n26622), .B(n26671), .Z(n26624) );
  XOR U26947 ( .A(n26672), .B(n26673), .Z(n26671) );
  ANDN U26948 ( .B(n26674), .A(n26675), .Z(n26672) );
  XOR U26949 ( .A(n26676), .B(n26673), .Z(n26674) );
  IV U26950 ( .A(n26626), .Z(n26622) );
  XOR U26951 ( .A(n26677), .B(n26678), .Z(n26626) );
  ANDN U26952 ( .B(n26679), .A(n26680), .Z(n26677) );
  XOR U26953 ( .A(n26681), .B(n26678), .Z(n26679) );
  IV U26954 ( .A(n26636), .Z(n26640) );
  XOR U26955 ( .A(n26636), .B(n26591), .Z(n26638) );
  XOR U26956 ( .A(n26682), .B(n26683), .Z(n26591) );
  AND U26957 ( .A(n638), .B(n26684), .Z(n26682) );
  XOR U26958 ( .A(n26685), .B(n26683), .Z(n26684) );
  NANDN U26959 ( .A(n26593), .B(n26595), .Z(n26636) );
  XOR U26960 ( .A(n26686), .B(n26687), .Z(n26595) );
  AND U26961 ( .A(n638), .B(n26688), .Z(n26686) );
  XOR U26962 ( .A(n26687), .B(n26689), .Z(n26688) );
  XNOR U26963 ( .A(n26690), .B(n26691), .Z(n638) );
  AND U26964 ( .A(n26692), .B(n26693), .Z(n26690) );
  XOR U26965 ( .A(n26691), .B(n26606), .Z(n26693) );
  XNOR U26966 ( .A(n26694), .B(n26695), .Z(n26606) );
  ANDN U26967 ( .B(n26696), .A(n26697), .Z(n26694) );
  XOR U26968 ( .A(n26695), .B(n26698), .Z(n26696) );
  XNOR U26969 ( .A(n26691), .B(n26608), .Z(n26692) );
  XOR U26970 ( .A(n26699), .B(n26700), .Z(n26608) );
  AND U26971 ( .A(n642), .B(n26701), .Z(n26699) );
  XOR U26972 ( .A(n26702), .B(n26700), .Z(n26701) );
  XNOR U26973 ( .A(n26703), .B(n26704), .Z(n26691) );
  AND U26974 ( .A(n26705), .B(n26706), .Z(n26703) );
  XNOR U26975 ( .A(n26704), .B(n26633), .Z(n26706) );
  XOR U26976 ( .A(n26697), .B(n26698), .Z(n26633) );
  XNOR U26977 ( .A(n26707), .B(n26708), .Z(n26698) );
  ANDN U26978 ( .B(n26709), .A(n26710), .Z(n26707) );
  XOR U26979 ( .A(n26711), .B(n26712), .Z(n26709) );
  XOR U26980 ( .A(n26713), .B(n26714), .Z(n26697) );
  XNOR U26981 ( .A(n26715), .B(n26716), .Z(n26714) );
  ANDN U26982 ( .B(n26717), .A(n26718), .Z(n26715) );
  XNOR U26983 ( .A(n26719), .B(n26720), .Z(n26717) );
  IV U26984 ( .A(n26695), .Z(n26713) );
  XOR U26985 ( .A(n26721), .B(n26722), .Z(n26695) );
  ANDN U26986 ( .B(n26723), .A(n26724), .Z(n26721) );
  XOR U26987 ( .A(n26722), .B(n26725), .Z(n26723) );
  XOR U26988 ( .A(n26704), .B(n26635), .Z(n26705) );
  XOR U26989 ( .A(n26726), .B(n26727), .Z(n26635) );
  AND U26990 ( .A(n642), .B(n26728), .Z(n26726) );
  XOR U26991 ( .A(n26729), .B(n26727), .Z(n26728) );
  XNOR U26992 ( .A(n26730), .B(n26731), .Z(n26704) );
  NAND U26993 ( .A(n26732), .B(n26733), .Z(n26731) );
  XOR U26994 ( .A(n26734), .B(n26683), .Z(n26733) );
  XOR U26995 ( .A(n26724), .B(n26725), .Z(n26683) );
  XOR U26996 ( .A(n26735), .B(n26712), .Z(n26725) );
  XOR U26997 ( .A(n26736), .B(n26737), .Z(n26712) );
  ANDN U26998 ( .B(n26738), .A(n26739), .Z(n26736) );
  XOR U26999 ( .A(n26737), .B(n26740), .Z(n26738) );
  IV U27000 ( .A(n26710), .Z(n26735) );
  XOR U27001 ( .A(n26708), .B(n26741), .Z(n26710) );
  XOR U27002 ( .A(n26742), .B(n26743), .Z(n26741) );
  ANDN U27003 ( .B(n26744), .A(n26745), .Z(n26742) );
  XOR U27004 ( .A(n26746), .B(n26743), .Z(n26744) );
  IV U27005 ( .A(n26711), .Z(n26708) );
  XOR U27006 ( .A(n26747), .B(n26748), .Z(n26711) );
  ANDN U27007 ( .B(n26749), .A(n26750), .Z(n26747) );
  XOR U27008 ( .A(n26748), .B(n26751), .Z(n26749) );
  XOR U27009 ( .A(n26752), .B(n26753), .Z(n26724) );
  XNOR U27010 ( .A(n26719), .B(n26754), .Z(n26753) );
  IV U27011 ( .A(n26722), .Z(n26754) );
  XOR U27012 ( .A(n26755), .B(n26756), .Z(n26722) );
  ANDN U27013 ( .B(n26757), .A(n26758), .Z(n26755) );
  XOR U27014 ( .A(n26756), .B(n26759), .Z(n26757) );
  XNOR U27015 ( .A(n26760), .B(n26761), .Z(n26719) );
  ANDN U27016 ( .B(n26762), .A(n26763), .Z(n26760) );
  XOR U27017 ( .A(n26761), .B(n26764), .Z(n26762) );
  IV U27018 ( .A(n26718), .Z(n26752) );
  XOR U27019 ( .A(n26716), .B(n26765), .Z(n26718) );
  XOR U27020 ( .A(n26766), .B(n26767), .Z(n26765) );
  ANDN U27021 ( .B(n26768), .A(n26769), .Z(n26766) );
  XOR U27022 ( .A(n26770), .B(n26767), .Z(n26768) );
  IV U27023 ( .A(n26720), .Z(n26716) );
  XOR U27024 ( .A(n26771), .B(n26772), .Z(n26720) );
  ANDN U27025 ( .B(n26773), .A(n26774), .Z(n26771) );
  XOR U27026 ( .A(n26775), .B(n26772), .Z(n26773) );
  IV U27027 ( .A(n26730), .Z(n26734) );
  XOR U27028 ( .A(n26730), .B(n26685), .Z(n26732) );
  XOR U27029 ( .A(n26776), .B(n26777), .Z(n26685) );
  AND U27030 ( .A(n642), .B(n26778), .Z(n26776) );
  XOR U27031 ( .A(n26779), .B(n26777), .Z(n26778) );
  NANDN U27032 ( .A(n26687), .B(n26689), .Z(n26730) );
  XOR U27033 ( .A(n26780), .B(n26781), .Z(n26689) );
  AND U27034 ( .A(n642), .B(n26782), .Z(n26780) );
  XOR U27035 ( .A(n26781), .B(n26783), .Z(n26782) );
  XNOR U27036 ( .A(n26784), .B(n26785), .Z(n642) );
  AND U27037 ( .A(n26786), .B(n26787), .Z(n26784) );
  XOR U27038 ( .A(n26785), .B(n26700), .Z(n26787) );
  XNOR U27039 ( .A(n26788), .B(n26789), .Z(n26700) );
  ANDN U27040 ( .B(n26790), .A(n26791), .Z(n26788) );
  XOR U27041 ( .A(n26789), .B(n26792), .Z(n26790) );
  XNOR U27042 ( .A(n26785), .B(n26702), .Z(n26786) );
  XOR U27043 ( .A(n26793), .B(n26794), .Z(n26702) );
  AND U27044 ( .A(n646), .B(n26795), .Z(n26793) );
  XOR U27045 ( .A(n26796), .B(n26794), .Z(n26795) );
  XNOR U27046 ( .A(n26797), .B(n26798), .Z(n26785) );
  AND U27047 ( .A(n26799), .B(n26800), .Z(n26797) );
  XNOR U27048 ( .A(n26798), .B(n26727), .Z(n26800) );
  XOR U27049 ( .A(n26791), .B(n26792), .Z(n26727) );
  XNOR U27050 ( .A(n26801), .B(n26802), .Z(n26792) );
  ANDN U27051 ( .B(n26803), .A(n26804), .Z(n26801) );
  XOR U27052 ( .A(n26805), .B(n26806), .Z(n26803) );
  XOR U27053 ( .A(n26807), .B(n26808), .Z(n26791) );
  XNOR U27054 ( .A(n26809), .B(n26810), .Z(n26808) );
  ANDN U27055 ( .B(n26811), .A(n26812), .Z(n26809) );
  XNOR U27056 ( .A(n26813), .B(n26814), .Z(n26811) );
  IV U27057 ( .A(n26789), .Z(n26807) );
  XOR U27058 ( .A(n26815), .B(n26816), .Z(n26789) );
  ANDN U27059 ( .B(n26817), .A(n26818), .Z(n26815) );
  XOR U27060 ( .A(n26816), .B(n26819), .Z(n26817) );
  XOR U27061 ( .A(n26798), .B(n26729), .Z(n26799) );
  XOR U27062 ( .A(n26820), .B(n26821), .Z(n26729) );
  AND U27063 ( .A(n646), .B(n26822), .Z(n26820) );
  XOR U27064 ( .A(n26823), .B(n26821), .Z(n26822) );
  XNOR U27065 ( .A(n26824), .B(n26825), .Z(n26798) );
  NAND U27066 ( .A(n26826), .B(n26827), .Z(n26825) );
  XOR U27067 ( .A(n26828), .B(n26777), .Z(n26827) );
  XOR U27068 ( .A(n26818), .B(n26819), .Z(n26777) );
  XOR U27069 ( .A(n26829), .B(n26806), .Z(n26819) );
  XOR U27070 ( .A(n26830), .B(n26831), .Z(n26806) );
  ANDN U27071 ( .B(n26832), .A(n26833), .Z(n26830) );
  XOR U27072 ( .A(n26831), .B(n26834), .Z(n26832) );
  IV U27073 ( .A(n26804), .Z(n26829) );
  XOR U27074 ( .A(n26802), .B(n26835), .Z(n26804) );
  XOR U27075 ( .A(n26836), .B(n26837), .Z(n26835) );
  ANDN U27076 ( .B(n26838), .A(n26839), .Z(n26836) );
  XOR U27077 ( .A(n26840), .B(n26837), .Z(n26838) );
  IV U27078 ( .A(n26805), .Z(n26802) );
  XOR U27079 ( .A(n26841), .B(n26842), .Z(n26805) );
  ANDN U27080 ( .B(n26843), .A(n26844), .Z(n26841) );
  XOR U27081 ( .A(n26842), .B(n26845), .Z(n26843) );
  XOR U27082 ( .A(n26846), .B(n26847), .Z(n26818) );
  XNOR U27083 ( .A(n26813), .B(n26848), .Z(n26847) );
  IV U27084 ( .A(n26816), .Z(n26848) );
  XOR U27085 ( .A(n26849), .B(n26850), .Z(n26816) );
  ANDN U27086 ( .B(n26851), .A(n26852), .Z(n26849) );
  XOR U27087 ( .A(n26850), .B(n26853), .Z(n26851) );
  XNOR U27088 ( .A(n26854), .B(n26855), .Z(n26813) );
  ANDN U27089 ( .B(n26856), .A(n26857), .Z(n26854) );
  XOR U27090 ( .A(n26855), .B(n26858), .Z(n26856) );
  IV U27091 ( .A(n26812), .Z(n26846) );
  XOR U27092 ( .A(n26810), .B(n26859), .Z(n26812) );
  XOR U27093 ( .A(n26860), .B(n26861), .Z(n26859) );
  ANDN U27094 ( .B(n26862), .A(n26863), .Z(n26860) );
  XOR U27095 ( .A(n26864), .B(n26861), .Z(n26862) );
  IV U27096 ( .A(n26814), .Z(n26810) );
  XOR U27097 ( .A(n26865), .B(n26866), .Z(n26814) );
  ANDN U27098 ( .B(n26867), .A(n26868), .Z(n26865) );
  XOR U27099 ( .A(n26869), .B(n26866), .Z(n26867) );
  IV U27100 ( .A(n26824), .Z(n26828) );
  XOR U27101 ( .A(n26824), .B(n26779), .Z(n26826) );
  XOR U27102 ( .A(n26870), .B(n26871), .Z(n26779) );
  AND U27103 ( .A(n646), .B(n26872), .Z(n26870) );
  XOR U27104 ( .A(n26873), .B(n26871), .Z(n26872) );
  NANDN U27105 ( .A(n26781), .B(n26783), .Z(n26824) );
  XOR U27106 ( .A(n26874), .B(n26875), .Z(n26783) );
  AND U27107 ( .A(n646), .B(n26876), .Z(n26874) );
  XOR U27108 ( .A(n26875), .B(n26877), .Z(n26876) );
  XNOR U27109 ( .A(n26878), .B(n26879), .Z(n646) );
  AND U27110 ( .A(n26880), .B(n26881), .Z(n26878) );
  XOR U27111 ( .A(n26879), .B(n26794), .Z(n26881) );
  XNOR U27112 ( .A(n26882), .B(n26883), .Z(n26794) );
  ANDN U27113 ( .B(n26884), .A(n26885), .Z(n26882) );
  XOR U27114 ( .A(n26883), .B(n26886), .Z(n26884) );
  XNOR U27115 ( .A(n26879), .B(n26796), .Z(n26880) );
  XOR U27116 ( .A(n26887), .B(n26888), .Z(n26796) );
  AND U27117 ( .A(n650), .B(n26889), .Z(n26887) );
  XOR U27118 ( .A(n26890), .B(n26888), .Z(n26889) );
  XNOR U27119 ( .A(n26891), .B(n26892), .Z(n26879) );
  AND U27120 ( .A(n26893), .B(n26894), .Z(n26891) );
  XNOR U27121 ( .A(n26892), .B(n26821), .Z(n26894) );
  XOR U27122 ( .A(n26885), .B(n26886), .Z(n26821) );
  XNOR U27123 ( .A(n26895), .B(n26896), .Z(n26886) );
  ANDN U27124 ( .B(n26897), .A(n26898), .Z(n26895) );
  XOR U27125 ( .A(n26899), .B(n26900), .Z(n26897) );
  XOR U27126 ( .A(n26901), .B(n26902), .Z(n26885) );
  XNOR U27127 ( .A(n26903), .B(n26904), .Z(n26902) );
  ANDN U27128 ( .B(n26905), .A(n26906), .Z(n26903) );
  XNOR U27129 ( .A(n26907), .B(n26908), .Z(n26905) );
  IV U27130 ( .A(n26883), .Z(n26901) );
  XOR U27131 ( .A(n26909), .B(n26910), .Z(n26883) );
  ANDN U27132 ( .B(n26911), .A(n26912), .Z(n26909) );
  XOR U27133 ( .A(n26910), .B(n26913), .Z(n26911) );
  XOR U27134 ( .A(n26892), .B(n26823), .Z(n26893) );
  XOR U27135 ( .A(n26914), .B(n26915), .Z(n26823) );
  AND U27136 ( .A(n650), .B(n26916), .Z(n26914) );
  XOR U27137 ( .A(n26917), .B(n26915), .Z(n26916) );
  XNOR U27138 ( .A(n26918), .B(n26919), .Z(n26892) );
  NAND U27139 ( .A(n26920), .B(n26921), .Z(n26919) );
  XOR U27140 ( .A(n26922), .B(n26871), .Z(n26921) );
  XOR U27141 ( .A(n26912), .B(n26913), .Z(n26871) );
  XOR U27142 ( .A(n26923), .B(n26900), .Z(n26913) );
  XOR U27143 ( .A(n26924), .B(n26925), .Z(n26900) );
  ANDN U27144 ( .B(n26926), .A(n26927), .Z(n26924) );
  XOR U27145 ( .A(n26925), .B(n26928), .Z(n26926) );
  IV U27146 ( .A(n26898), .Z(n26923) );
  XOR U27147 ( .A(n26896), .B(n26929), .Z(n26898) );
  XOR U27148 ( .A(n26930), .B(n26931), .Z(n26929) );
  ANDN U27149 ( .B(n26932), .A(n26933), .Z(n26930) );
  XOR U27150 ( .A(n26934), .B(n26931), .Z(n26932) );
  IV U27151 ( .A(n26899), .Z(n26896) );
  XOR U27152 ( .A(n26935), .B(n26936), .Z(n26899) );
  ANDN U27153 ( .B(n26937), .A(n26938), .Z(n26935) );
  XOR U27154 ( .A(n26936), .B(n26939), .Z(n26937) );
  XOR U27155 ( .A(n26940), .B(n26941), .Z(n26912) );
  XNOR U27156 ( .A(n26907), .B(n26942), .Z(n26941) );
  IV U27157 ( .A(n26910), .Z(n26942) );
  XOR U27158 ( .A(n26943), .B(n26944), .Z(n26910) );
  ANDN U27159 ( .B(n26945), .A(n26946), .Z(n26943) );
  XOR U27160 ( .A(n26944), .B(n26947), .Z(n26945) );
  XNOR U27161 ( .A(n26948), .B(n26949), .Z(n26907) );
  ANDN U27162 ( .B(n26950), .A(n26951), .Z(n26948) );
  XOR U27163 ( .A(n26949), .B(n26952), .Z(n26950) );
  IV U27164 ( .A(n26906), .Z(n26940) );
  XOR U27165 ( .A(n26904), .B(n26953), .Z(n26906) );
  XOR U27166 ( .A(n26954), .B(n26955), .Z(n26953) );
  ANDN U27167 ( .B(n26956), .A(n26957), .Z(n26954) );
  XOR U27168 ( .A(n26958), .B(n26955), .Z(n26956) );
  IV U27169 ( .A(n26908), .Z(n26904) );
  XOR U27170 ( .A(n26959), .B(n26960), .Z(n26908) );
  ANDN U27171 ( .B(n26961), .A(n26962), .Z(n26959) );
  XOR U27172 ( .A(n26963), .B(n26960), .Z(n26961) );
  IV U27173 ( .A(n26918), .Z(n26922) );
  XOR U27174 ( .A(n26918), .B(n26873), .Z(n26920) );
  XOR U27175 ( .A(n26964), .B(n26965), .Z(n26873) );
  AND U27176 ( .A(n650), .B(n26966), .Z(n26964) );
  XOR U27177 ( .A(n26967), .B(n26965), .Z(n26966) );
  NANDN U27178 ( .A(n26875), .B(n26877), .Z(n26918) );
  XOR U27179 ( .A(n26968), .B(n26969), .Z(n26877) );
  AND U27180 ( .A(n650), .B(n26970), .Z(n26968) );
  XOR U27181 ( .A(n26969), .B(n26971), .Z(n26970) );
  XNOR U27182 ( .A(n26972), .B(n26973), .Z(n650) );
  AND U27183 ( .A(n26974), .B(n26975), .Z(n26972) );
  XOR U27184 ( .A(n26973), .B(n26888), .Z(n26975) );
  XNOR U27185 ( .A(n26976), .B(n26977), .Z(n26888) );
  ANDN U27186 ( .B(n26978), .A(n26979), .Z(n26976) );
  XOR U27187 ( .A(n26977), .B(n26980), .Z(n26978) );
  XNOR U27188 ( .A(n26973), .B(n26890), .Z(n26974) );
  XOR U27189 ( .A(n26981), .B(n26982), .Z(n26890) );
  AND U27190 ( .A(n654), .B(n26983), .Z(n26981) );
  XOR U27191 ( .A(n26984), .B(n26982), .Z(n26983) );
  XNOR U27192 ( .A(n26985), .B(n26986), .Z(n26973) );
  AND U27193 ( .A(n26987), .B(n26988), .Z(n26985) );
  XNOR U27194 ( .A(n26986), .B(n26915), .Z(n26988) );
  XOR U27195 ( .A(n26979), .B(n26980), .Z(n26915) );
  XNOR U27196 ( .A(n26989), .B(n26990), .Z(n26980) );
  ANDN U27197 ( .B(n26991), .A(n26992), .Z(n26989) );
  XOR U27198 ( .A(n26993), .B(n26994), .Z(n26991) );
  XOR U27199 ( .A(n26995), .B(n26996), .Z(n26979) );
  XNOR U27200 ( .A(n26997), .B(n26998), .Z(n26996) );
  ANDN U27201 ( .B(n26999), .A(n27000), .Z(n26997) );
  XNOR U27202 ( .A(n27001), .B(n27002), .Z(n26999) );
  IV U27203 ( .A(n26977), .Z(n26995) );
  XOR U27204 ( .A(n27003), .B(n27004), .Z(n26977) );
  ANDN U27205 ( .B(n27005), .A(n27006), .Z(n27003) );
  XOR U27206 ( .A(n27004), .B(n27007), .Z(n27005) );
  XOR U27207 ( .A(n26986), .B(n26917), .Z(n26987) );
  XOR U27208 ( .A(n27008), .B(n27009), .Z(n26917) );
  AND U27209 ( .A(n654), .B(n27010), .Z(n27008) );
  XOR U27210 ( .A(n27011), .B(n27009), .Z(n27010) );
  XNOR U27211 ( .A(n27012), .B(n27013), .Z(n26986) );
  NAND U27212 ( .A(n27014), .B(n27015), .Z(n27013) );
  XOR U27213 ( .A(n27016), .B(n26965), .Z(n27015) );
  XOR U27214 ( .A(n27006), .B(n27007), .Z(n26965) );
  XOR U27215 ( .A(n27017), .B(n26994), .Z(n27007) );
  XOR U27216 ( .A(n27018), .B(n27019), .Z(n26994) );
  ANDN U27217 ( .B(n27020), .A(n27021), .Z(n27018) );
  XOR U27218 ( .A(n27019), .B(n27022), .Z(n27020) );
  IV U27219 ( .A(n26992), .Z(n27017) );
  XOR U27220 ( .A(n26990), .B(n27023), .Z(n26992) );
  XOR U27221 ( .A(n27024), .B(n27025), .Z(n27023) );
  ANDN U27222 ( .B(n27026), .A(n27027), .Z(n27024) );
  XOR U27223 ( .A(n27028), .B(n27025), .Z(n27026) );
  IV U27224 ( .A(n26993), .Z(n26990) );
  XOR U27225 ( .A(n27029), .B(n27030), .Z(n26993) );
  ANDN U27226 ( .B(n27031), .A(n27032), .Z(n27029) );
  XOR U27227 ( .A(n27030), .B(n27033), .Z(n27031) );
  XOR U27228 ( .A(n27034), .B(n27035), .Z(n27006) );
  XNOR U27229 ( .A(n27001), .B(n27036), .Z(n27035) );
  IV U27230 ( .A(n27004), .Z(n27036) );
  XOR U27231 ( .A(n27037), .B(n27038), .Z(n27004) );
  ANDN U27232 ( .B(n27039), .A(n27040), .Z(n27037) );
  XOR U27233 ( .A(n27038), .B(n27041), .Z(n27039) );
  XNOR U27234 ( .A(n27042), .B(n27043), .Z(n27001) );
  ANDN U27235 ( .B(n27044), .A(n27045), .Z(n27042) );
  XOR U27236 ( .A(n27043), .B(n27046), .Z(n27044) );
  IV U27237 ( .A(n27000), .Z(n27034) );
  XOR U27238 ( .A(n26998), .B(n27047), .Z(n27000) );
  XOR U27239 ( .A(n27048), .B(n27049), .Z(n27047) );
  ANDN U27240 ( .B(n27050), .A(n27051), .Z(n27048) );
  XOR U27241 ( .A(n27052), .B(n27049), .Z(n27050) );
  IV U27242 ( .A(n27002), .Z(n26998) );
  XOR U27243 ( .A(n27053), .B(n27054), .Z(n27002) );
  ANDN U27244 ( .B(n27055), .A(n27056), .Z(n27053) );
  XOR U27245 ( .A(n27057), .B(n27054), .Z(n27055) );
  IV U27246 ( .A(n27012), .Z(n27016) );
  XOR U27247 ( .A(n27012), .B(n26967), .Z(n27014) );
  XOR U27248 ( .A(n27058), .B(n27059), .Z(n26967) );
  AND U27249 ( .A(n654), .B(n27060), .Z(n27058) );
  XOR U27250 ( .A(n27061), .B(n27059), .Z(n27060) );
  NANDN U27251 ( .A(n26969), .B(n26971), .Z(n27012) );
  XOR U27252 ( .A(n27062), .B(n27063), .Z(n26971) );
  AND U27253 ( .A(n654), .B(n27064), .Z(n27062) );
  XOR U27254 ( .A(n27063), .B(n27065), .Z(n27064) );
  XNOR U27255 ( .A(n27066), .B(n27067), .Z(n654) );
  AND U27256 ( .A(n27068), .B(n27069), .Z(n27066) );
  XOR U27257 ( .A(n27067), .B(n26982), .Z(n27069) );
  XNOR U27258 ( .A(n27070), .B(n27071), .Z(n26982) );
  ANDN U27259 ( .B(n27072), .A(n27073), .Z(n27070) );
  XOR U27260 ( .A(n27071), .B(n27074), .Z(n27072) );
  XNOR U27261 ( .A(n27067), .B(n26984), .Z(n27068) );
  XOR U27262 ( .A(n27075), .B(n27076), .Z(n26984) );
  AND U27263 ( .A(n658), .B(n27077), .Z(n27075) );
  XOR U27264 ( .A(n27078), .B(n27076), .Z(n27077) );
  XNOR U27265 ( .A(n27079), .B(n27080), .Z(n27067) );
  AND U27266 ( .A(n27081), .B(n27082), .Z(n27079) );
  XNOR U27267 ( .A(n27080), .B(n27009), .Z(n27082) );
  XOR U27268 ( .A(n27073), .B(n27074), .Z(n27009) );
  XNOR U27269 ( .A(n27083), .B(n27084), .Z(n27074) );
  ANDN U27270 ( .B(n27085), .A(n27086), .Z(n27083) );
  XOR U27271 ( .A(n27087), .B(n27088), .Z(n27085) );
  XOR U27272 ( .A(n27089), .B(n27090), .Z(n27073) );
  XNOR U27273 ( .A(n27091), .B(n27092), .Z(n27090) );
  ANDN U27274 ( .B(n27093), .A(n27094), .Z(n27091) );
  XNOR U27275 ( .A(n27095), .B(n27096), .Z(n27093) );
  IV U27276 ( .A(n27071), .Z(n27089) );
  XOR U27277 ( .A(n27097), .B(n27098), .Z(n27071) );
  ANDN U27278 ( .B(n27099), .A(n27100), .Z(n27097) );
  XOR U27279 ( .A(n27098), .B(n27101), .Z(n27099) );
  XOR U27280 ( .A(n27080), .B(n27011), .Z(n27081) );
  XOR U27281 ( .A(n27102), .B(n27103), .Z(n27011) );
  AND U27282 ( .A(n658), .B(n27104), .Z(n27102) );
  XOR U27283 ( .A(n27105), .B(n27103), .Z(n27104) );
  XNOR U27284 ( .A(n27106), .B(n27107), .Z(n27080) );
  NAND U27285 ( .A(n27108), .B(n27109), .Z(n27107) );
  XOR U27286 ( .A(n27110), .B(n27059), .Z(n27109) );
  XOR U27287 ( .A(n27100), .B(n27101), .Z(n27059) );
  XOR U27288 ( .A(n27111), .B(n27088), .Z(n27101) );
  XOR U27289 ( .A(n27112), .B(n27113), .Z(n27088) );
  ANDN U27290 ( .B(n27114), .A(n27115), .Z(n27112) );
  XOR U27291 ( .A(n27113), .B(n27116), .Z(n27114) );
  IV U27292 ( .A(n27086), .Z(n27111) );
  XOR U27293 ( .A(n27084), .B(n27117), .Z(n27086) );
  XOR U27294 ( .A(n27118), .B(n27119), .Z(n27117) );
  ANDN U27295 ( .B(n27120), .A(n27121), .Z(n27118) );
  XOR U27296 ( .A(n27122), .B(n27119), .Z(n27120) );
  IV U27297 ( .A(n27087), .Z(n27084) );
  XOR U27298 ( .A(n27123), .B(n27124), .Z(n27087) );
  ANDN U27299 ( .B(n27125), .A(n27126), .Z(n27123) );
  XOR U27300 ( .A(n27124), .B(n27127), .Z(n27125) );
  XOR U27301 ( .A(n27128), .B(n27129), .Z(n27100) );
  XNOR U27302 ( .A(n27095), .B(n27130), .Z(n27129) );
  IV U27303 ( .A(n27098), .Z(n27130) );
  XOR U27304 ( .A(n27131), .B(n27132), .Z(n27098) );
  ANDN U27305 ( .B(n27133), .A(n27134), .Z(n27131) );
  XOR U27306 ( .A(n27132), .B(n27135), .Z(n27133) );
  XNOR U27307 ( .A(n27136), .B(n27137), .Z(n27095) );
  ANDN U27308 ( .B(n27138), .A(n27139), .Z(n27136) );
  XOR U27309 ( .A(n27137), .B(n27140), .Z(n27138) );
  IV U27310 ( .A(n27094), .Z(n27128) );
  XOR U27311 ( .A(n27092), .B(n27141), .Z(n27094) );
  XOR U27312 ( .A(n27142), .B(n27143), .Z(n27141) );
  ANDN U27313 ( .B(n27144), .A(n27145), .Z(n27142) );
  XOR U27314 ( .A(n27146), .B(n27143), .Z(n27144) );
  IV U27315 ( .A(n27096), .Z(n27092) );
  XOR U27316 ( .A(n27147), .B(n27148), .Z(n27096) );
  ANDN U27317 ( .B(n27149), .A(n27150), .Z(n27147) );
  XOR U27318 ( .A(n27151), .B(n27148), .Z(n27149) );
  IV U27319 ( .A(n27106), .Z(n27110) );
  XOR U27320 ( .A(n27106), .B(n27061), .Z(n27108) );
  XOR U27321 ( .A(n27152), .B(n27153), .Z(n27061) );
  AND U27322 ( .A(n658), .B(n27154), .Z(n27152) );
  XOR U27323 ( .A(n27155), .B(n27153), .Z(n27154) );
  NANDN U27324 ( .A(n27063), .B(n27065), .Z(n27106) );
  XOR U27325 ( .A(n27156), .B(n27157), .Z(n27065) );
  AND U27326 ( .A(n658), .B(n27158), .Z(n27156) );
  XOR U27327 ( .A(n27157), .B(n27159), .Z(n27158) );
  XNOR U27328 ( .A(n27160), .B(n27161), .Z(n658) );
  AND U27329 ( .A(n27162), .B(n27163), .Z(n27160) );
  XOR U27330 ( .A(n27161), .B(n27076), .Z(n27163) );
  XNOR U27331 ( .A(n27164), .B(n27165), .Z(n27076) );
  ANDN U27332 ( .B(n27166), .A(n27167), .Z(n27164) );
  XOR U27333 ( .A(n27165), .B(n27168), .Z(n27166) );
  XNOR U27334 ( .A(n27161), .B(n27078), .Z(n27162) );
  XOR U27335 ( .A(n27169), .B(n27170), .Z(n27078) );
  AND U27336 ( .A(n662), .B(n27171), .Z(n27169) );
  XOR U27337 ( .A(n27172), .B(n27170), .Z(n27171) );
  XNOR U27338 ( .A(n27173), .B(n27174), .Z(n27161) );
  AND U27339 ( .A(n27175), .B(n27176), .Z(n27173) );
  XNOR U27340 ( .A(n27174), .B(n27103), .Z(n27176) );
  XOR U27341 ( .A(n27167), .B(n27168), .Z(n27103) );
  XNOR U27342 ( .A(n27177), .B(n27178), .Z(n27168) );
  ANDN U27343 ( .B(n27179), .A(n27180), .Z(n27177) );
  XOR U27344 ( .A(n27181), .B(n27182), .Z(n27179) );
  XOR U27345 ( .A(n27183), .B(n27184), .Z(n27167) );
  XNOR U27346 ( .A(n27185), .B(n27186), .Z(n27184) );
  ANDN U27347 ( .B(n27187), .A(n27188), .Z(n27185) );
  XNOR U27348 ( .A(n27189), .B(n27190), .Z(n27187) );
  IV U27349 ( .A(n27165), .Z(n27183) );
  XOR U27350 ( .A(n27191), .B(n27192), .Z(n27165) );
  ANDN U27351 ( .B(n27193), .A(n27194), .Z(n27191) );
  XOR U27352 ( .A(n27192), .B(n27195), .Z(n27193) );
  XOR U27353 ( .A(n27174), .B(n27105), .Z(n27175) );
  XOR U27354 ( .A(n27196), .B(n27197), .Z(n27105) );
  AND U27355 ( .A(n662), .B(n27198), .Z(n27196) );
  XOR U27356 ( .A(n27199), .B(n27197), .Z(n27198) );
  XNOR U27357 ( .A(n27200), .B(n27201), .Z(n27174) );
  NAND U27358 ( .A(n27202), .B(n27203), .Z(n27201) );
  XOR U27359 ( .A(n27204), .B(n27153), .Z(n27203) );
  XOR U27360 ( .A(n27194), .B(n27195), .Z(n27153) );
  XOR U27361 ( .A(n27205), .B(n27182), .Z(n27195) );
  XOR U27362 ( .A(n27206), .B(n27207), .Z(n27182) );
  ANDN U27363 ( .B(n27208), .A(n27209), .Z(n27206) );
  XOR U27364 ( .A(n27207), .B(n27210), .Z(n27208) );
  IV U27365 ( .A(n27180), .Z(n27205) );
  XOR U27366 ( .A(n27178), .B(n27211), .Z(n27180) );
  XOR U27367 ( .A(n27212), .B(n27213), .Z(n27211) );
  ANDN U27368 ( .B(n27214), .A(n27215), .Z(n27212) );
  XOR U27369 ( .A(n27216), .B(n27213), .Z(n27214) );
  IV U27370 ( .A(n27181), .Z(n27178) );
  XOR U27371 ( .A(n27217), .B(n27218), .Z(n27181) );
  ANDN U27372 ( .B(n27219), .A(n27220), .Z(n27217) );
  XOR U27373 ( .A(n27218), .B(n27221), .Z(n27219) );
  XOR U27374 ( .A(n27222), .B(n27223), .Z(n27194) );
  XNOR U27375 ( .A(n27189), .B(n27224), .Z(n27223) );
  IV U27376 ( .A(n27192), .Z(n27224) );
  XOR U27377 ( .A(n27225), .B(n27226), .Z(n27192) );
  ANDN U27378 ( .B(n27227), .A(n27228), .Z(n27225) );
  XOR U27379 ( .A(n27226), .B(n27229), .Z(n27227) );
  XNOR U27380 ( .A(n27230), .B(n27231), .Z(n27189) );
  ANDN U27381 ( .B(n27232), .A(n27233), .Z(n27230) );
  XOR U27382 ( .A(n27231), .B(n27234), .Z(n27232) );
  IV U27383 ( .A(n27188), .Z(n27222) );
  XOR U27384 ( .A(n27186), .B(n27235), .Z(n27188) );
  XOR U27385 ( .A(n27236), .B(n27237), .Z(n27235) );
  ANDN U27386 ( .B(n27238), .A(n27239), .Z(n27236) );
  XOR U27387 ( .A(n27240), .B(n27237), .Z(n27238) );
  IV U27388 ( .A(n27190), .Z(n27186) );
  XOR U27389 ( .A(n27241), .B(n27242), .Z(n27190) );
  ANDN U27390 ( .B(n27243), .A(n27244), .Z(n27241) );
  XOR U27391 ( .A(n27245), .B(n27242), .Z(n27243) );
  IV U27392 ( .A(n27200), .Z(n27204) );
  XOR U27393 ( .A(n27200), .B(n27155), .Z(n27202) );
  XOR U27394 ( .A(n27246), .B(n27247), .Z(n27155) );
  AND U27395 ( .A(n662), .B(n27248), .Z(n27246) );
  XOR U27396 ( .A(n27249), .B(n27247), .Z(n27248) );
  NANDN U27397 ( .A(n27157), .B(n27159), .Z(n27200) );
  XOR U27398 ( .A(n27250), .B(n27251), .Z(n27159) );
  AND U27399 ( .A(n662), .B(n27252), .Z(n27250) );
  XOR U27400 ( .A(n27251), .B(n27253), .Z(n27252) );
  XNOR U27401 ( .A(n27254), .B(n27255), .Z(n662) );
  AND U27402 ( .A(n27256), .B(n27257), .Z(n27254) );
  XOR U27403 ( .A(n27255), .B(n27170), .Z(n27257) );
  XNOR U27404 ( .A(n27258), .B(n27259), .Z(n27170) );
  ANDN U27405 ( .B(n27260), .A(n27261), .Z(n27258) );
  XOR U27406 ( .A(n27259), .B(n27262), .Z(n27260) );
  XNOR U27407 ( .A(n27255), .B(n27172), .Z(n27256) );
  XOR U27408 ( .A(n27263), .B(n27264), .Z(n27172) );
  AND U27409 ( .A(n666), .B(n27265), .Z(n27263) );
  XOR U27410 ( .A(n27266), .B(n27264), .Z(n27265) );
  XNOR U27411 ( .A(n27267), .B(n27268), .Z(n27255) );
  AND U27412 ( .A(n27269), .B(n27270), .Z(n27267) );
  XNOR U27413 ( .A(n27268), .B(n27197), .Z(n27270) );
  XOR U27414 ( .A(n27261), .B(n27262), .Z(n27197) );
  XNOR U27415 ( .A(n27271), .B(n27272), .Z(n27262) );
  ANDN U27416 ( .B(n27273), .A(n27274), .Z(n27271) );
  XOR U27417 ( .A(n27275), .B(n27276), .Z(n27273) );
  XOR U27418 ( .A(n27277), .B(n27278), .Z(n27261) );
  XNOR U27419 ( .A(n27279), .B(n27280), .Z(n27278) );
  ANDN U27420 ( .B(n27281), .A(n27282), .Z(n27279) );
  XNOR U27421 ( .A(n27283), .B(n27284), .Z(n27281) );
  IV U27422 ( .A(n27259), .Z(n27277) );
  XOR U27423 ( .A(n27285), .B(n27286), .Z(n27259) );
  ANDN U27424 ( .B(n27287), .A(n27288), .Z(n27285) );
  XOR U27425 ( .A(n27286), .B(n27289), .Z(n27287) );
  XOR U27426 ( .A(n27268), .B(n27199), .Z(n27269) );
  XOR U27427 ( .A(n27290), .B(n27291), .Z(n27199) );
  AND U27428 ( .A(n666), .B(n27292), .Z(n27290) );
  XOR U27429 ( .A(n27293), .B(n27291), .Z(n27292) );
  XNOR U27430 ( .A(n27294), .B(n27295), .Z(n27268) );
  NAND U27431 ( .A(n27296), .B(n27297), .Z(n27295) );
  XOR U27432 ( .A(n27298), .B(n27247), .Z(n27297) );
  XOR U27433 ( .A(n27288), .B(n27289), .Z(n27247) );
  XOR U27434 ( .A(n27299), .B(n27276), .Z(n27289) );
  XOR U27435 ( .A(n27300), .B(n27301), .Z(n27276) );
  ANDN U27436 ( .B(n27302), .A(n27303), .Z(n27300) );
  XOR U27437 ( .A(n27301), .B(n27304), .Z(n27302) );
  IV U27438 ( .A(n27274), .Z(n27299) );
  XOR U27439 ( .A(n27272), .B(n27305), .Z(n27274) );
  XOR U27440 ( .A(n27306), .B(n27307), .Z(n27305) );
  ANDN U27441 ( .B(n27308), .A(n27309), .Z(n27306) );
  XOR U27442 ( .A(n27310), .B(n27307), .Z(n27308) );
  IV U27443 ( .A(n27275), .Z(n27272) );
  XOR U27444 ( .A(n27311), .B(n27312), .Z(n27275) );
  ANDN U27445 ( .B(n27313), .A(n27314), .Z(n27311) );
  XOR U27446 ( .A(n27312), .B(n27315), .Z(n27313) );
  XOR U27447 ( .A(n27316), .B(n27317), .Z(n27288) );
  XNOR U27448 ( .A(n27283), .B(n27318), .Z(n27317) );
  IV U27449 ( .A(n27286), .Z(n27318) );
  XOR U27450 ( .A(n27319), .B(n27320), .Z(n27286) );
  ANDN U27451 ( .B(n27321), .A(n27322), .Z(n27319) );
  XOR U27452 ( .A(n27320), .B(n27323), .Z(n27321) );
  XNOR U27453 ( .A(n27324), .B(n27325), .Z(n27283) );
  ANDN U27454 ( .B(n27326), .A(n27327), .Z(n27324) );
  XOR U27455 ( .A(n27325), .B(n27328), .Z(n27326) );
  IV U27456 ( .A(n27282), .Z(n27316) );
  XOR U27457 ( .A(n27280), .B(n27329), .Z(n27282) );
  XOR U27458 ( .A(n27330), .B(n27331), .Z(n27329) );
  ANDN U27459 ( .B(n27332), .A(n27333), .Z(n27330) );
  XOR U27460 ( .A(n27334), .B(n27331), .Z(n27332) );
  IV U27461 ( .A(n27284), .Z(n27280) );
  XOR U27462 ( .A(n27335), .B(n27336), .Z(n27284) );
  ANDN U27463 ( .B(n27337), .A(n27338), .Z(n27335) );
  XOR U27464 ( .A(n27339), .B(n27336), .Z(n27337) );
  IV U27465 ( .A(n27294), .Z(n27298) );
  XOR U27466 ( .A(n27294), .B(n27249), .Z(n27296) );
  XOR U27467 ( .A(n27340), .B(n27341), .Z(n27249) );
  AND U27468 ( .A(n666), .B(n27342), .Z(n27340) );
  XOR U27469 ( .A(n27343), .B(n27341), .Z(n27342) );
  NANDN U27470 ( .A(n27251), .B(n27253), .Z(n27294) );
  XOR U27471 ( .A(n27344), .B(n27345), .Z(n27253) );
  AND U27472 ( .A(n666), .B(n27346), .Z(n27344) );
  XOR U27473 ( .A(n27345), .B(n27347), .Z(n27346) );
  XNOR U27474 ( .A(n27348), .B(n27349), .Z(n666) );
  AND U27475 ( .A(n27350), .B(n27351), .Z(n27348) );
  XOR U27476 ( .A(n27349), .B(n27264), .Z(n27351) );
  XNOR U27477 ( .A(n27352), .B(n27353), .Z(n27264) );
  ANDN U27478 ( .B(n27354), .A(n27355), .Z(n27352) );
  XOR U27479 ( .A(n27353), .B(n27356), .Z(n27354) );
  XNOR U27480 ( .A(n27349), .B(n27266), .Z(n27350) );
  XOR U27481 ( .A(n27357), .B(n27358), .Z(n27266) );
  AND U27482 ( .A(n670), .B(n27359), .Z(n27357) );
  XOR U27483 ( .A(n27360), .B(n27358), .Z(n27359) );
  XNOR U27484 ( .A(n27361), .B(n27362), .Z(n27349) );
  AND U27485 ( .A(n27363), .B(n27364), .Z(n27361) );
  XNOR U27486 ( .A(n27362), .B(n27291), .Z(n27364) );
  XOR U27487 ( .A(n27355), .B(n27356), .Z(n27291) );
  XNOR U27488 ( .A(n27365), .B(n27366), .Z(n27356) );
  ANDN U27489 ( .B(n27367), .A(n27368), .Z(n27365) );
  XOR U27490 ( .A(n27369), .B(n27370), .Z(n27367) );
  XOR U27491 ( .A(n27371), .B(n27372), .Z(n27355) );
  XNOR U27492 ( .A(n27373), .B(n27374), .Z(n27372) );
  ANDN U27493 ( .B(n27375), .A(n27376), .Z(n27373) );
  XNOR U27494 ( .A(n27377), .B(n27378), .Z(n27375) );
  IV U27495 ( .A(n27353), .Z(n27371) );
  XOR U27496 ( .A(n27379), .B(n27380), .Z(n27353) );
  ANDN U27497 ( .B(n27381), .A(n27382), .Z(n27379) );
  XOR U27498 ( .A(n27380), .B(n27383), .Z(n27381) );
  XOR U27499 ( .A(n27362), .B(n27293), .Z(n27363) );
  XOR U27500 ( .A(n27384), .B(n27385), .Z(n27293) );
  AND U27501 ( .A(n670), .B(n27386), .Z(n27384) );
  XOR U27502 ( .A(n27387), .B(n27385), .Z(n27386) );
  XNOR U27503 ( .A(n27388), .B(n27389), .Z(n27362) );
  NAND U27504 ( .A(n27390), .B(n27391), .Z(n27389) );
  XOR U27505 ( .A(n27392), .B(n27341), .Z(n27391) );
  XOR U27506 ( .A(n27382), .B(n27383), .Z(n27341) );
  XOR U27507 ( .A(n27393), .B(n27370), .Z(n27383) );
  XOR U27508 ( .A(n27394), .B(n27395), .Z(n27370) );
  ANDN U27509 ( .B(n27396), .A(n27397), .Z(n27394) );
  XOR U27510 ( .A(n27395), .B(n27398), .Z(n27396) );
  IV U27511 ( .A(n27368), .Z(n27393) );
  XOR U27512 ( .A(n27366), .B(n27399), .Z(n27368) );
  XOR U27513 ( .A(n27400), .B(n27401), .Z(n27399) );
  ANDN U27514 ( .B(n27402), .A(n27403), .Z(n27400) );
  XOR U27515 ( .A(n27404), .B(n27401), .Z(n27402) );
  IV U27516 ( .A(n27369), .Z(n27366) );
  XOR U27517 ( .A(n27405), .B(n27406), .Z(n27369) );
  ANDN U27518 ( .B(n27407), .A(n27408), .Z(n27405) );
  XOR U27519 ( .A(n27406), .B(n27409), .Z(n27407) );
  XOR U27520 ( .A(n27410), .B(n27411), .Z(n27382) );
  XNOR U27521 ( .A(n27377), .B(n27412), .Z(n27411) );
  IV U27522 ( .A(n27380), .Z(n27412) );
  XOR U27523 ( .A(n27413), .B(n27414), .Z(n27380) );
  ANDN U27524 ( .B(n27415), .A(n27416), .Z(n27413) );
  XOR U27525 ( .A(n27414), .B(n27417), .Z(n27415) );
  XNOR U27526 ( .A(n27418), .B(n27419), .Z(n27377) );
  ANDN U27527 ( .B(n27420), .A(n27421), .Z(n27418) );
  XOR U27528 ( .A(n27419), .B(n27422), .Z(n27420) );
  IV U27529 ( .A(n27376), .Z(n27410) );
  XOR U27530 ( .A(n27374), .B(n27423), .Z(n27376) );
  XOR U27531 ( .A(n27424), .B(n27425), .Z(n27423) );
  ANDN U27532 ( .B(n27426), .A(n27427), .Z(n27424) );
  XOR U27533 ( .A(n27428), .B(n27425), .Z(n27426) );
  IV U27534 ( .A(n27378), .Z(n27374) );
  XOR U27535 ( .A(n27429), .B(n27430), .Z(n27378) );
  ANDN U27536 ( .B(n27431), .A(n27432), .Z(n27429) );
  XOR U27537 ( .A(n27433), .B(n27430), .Z(n27431) );
  IV U27538 ( .A(n27388), .Z(n27392) );
  XOR U27539 ( .A(n27388), .B(n27343), .Z(n27390) );
  XOR U27540 ( .A(n27434), .B(n27435), .Z(n27343) );
  AND U27541 ( .A(n670), .B(n27436), .Z(n27434) );
  XOR U27542 ( .A(n27437), .B(n27435), .Z(n27436) );
  NANDN U27543 ( .A(n27345), .B(n27347), .Z(n27388) );
  XOR U27544 ( .A(n27438), .B(n27439), .Z(n27347) );
  AND U27545 ( .A(n670), .B(n27440), .Z(n27438) );
  XOR U27546 ( .A(n27439), .B(n27441), .Z(n27440) );
  XNOR U27547 ( .A(n27442), .B(n27443), .Z(n670) );
  AND U27548 ( .A(n27444), .B(n27445), .Z(n27442) );
  XOR U27549 ( .A(n27443), .B(n27358), .Z(n27445) );
  XNOR U27550 ( .A(n27446), .B(n27447), .Z(n27358) );
  ANDN U27551 ( .B(n27448), .A(n27449), .Z(n27446) );
  XOR U27552 ( .A(n27447), .B(n27450), .Z(n27448) );
  XNOR U27553 ( .A(n27443), .B(n27360), .Z(n27444) );
  XOR U27554 ( .A(n27451), .B(n27452), .Z(n27360) );
  AND U27555 ( .A(n674), .B(n27453), .Z(n27451) );
  XOR U27556 ( .A(n27454), .B(n27452), .Z(n27453) );
  XNOR U27557 ( .A(n27455), .B(n27456), .Z(n27443) );
  AND U27558 ( .A(n27457), .B(n27458), .Z(n27455) );
  XNOR U27559 ( .A(n27456), .B(n27385), .Z(n27458) );
  XOR U27560 ( .A(n27449), .B(n27450), .Z(n27385) );
  XNOR U27561 ( .A(n27459), .B(n27460), .Z(n27450) );
  ANDN U27562 ( .B(n27461), .A(n27462), .Z(n27459) );
  XOR U27563 ( .A(n27463), .B(n27464), .Z(n27461) );
  XOR U27564 ( .A(n27465), .B(n27466), .Z(n27449) );
  XNOR U27565 ( .A(n27467), .B(n27468), .Z(n27466) );
  ANDN U27566 ( .B(n27469), .A(n27470), .Z(n27467) );
  XNOR U27567 ( .A(n27471), .B(n27472), .Z(n27469) );
  IV U27568 ( .A(n27447), .Z(n27465) );
  XOR U27569 ( .A(n27473), .B(n27474), .Z(n27447) );
  ANDN U27570 ( .B(n27475), .A(n27476), .Z(n27473) );
  XOR U27571 ( .A(n27474), .B(n27477), .Z(n27475) );
  XOR U27572 ( .A(n27456), .B(n27387), .Z(n27457) );
  XOR U27573 ( .A(n27478), .B(n27479), .Z(n27387) );
  AND U27574 ( .A(n674), .B(n27480), .Z(n27478) );
  XOR U27575 ( .A(n27481), .B(n27479), .Z(n27480) );
  XNOR U27576 ( .A(n27482), .B(n27483), .Z(n27456) );
  NAND U27577 ( .A(n27484), .B(n27485), .Z(n27483) );
  XOR U27578 ( .A(n27486), .B(n27435), .Z(n27485) );
  XOR U27579 ( .A(n27476), .B(n27477), .Z(n27435) );
  XOR U27580 ( .A(n27487), .B(n27464), .Z(n27477) );
  XOR U27581 ( .A(n27488), .B(n27489), .Z(n27464) );
  ANDN U27582 ( .B(n27490), .A(n27491), .Z(n27488) );
  XOR U27583 ( .A(n27489), .B(n27492), .Z(n27490) );
  IV U27584 ( .A(n27462), .Z(n27487) );
  XOR U27585 ( .A(n27460), .B(n27493), .Z(n27462) );
  XOR U27586 ( .A(n27494), .B(n27495), .Z(n27493) );
  ANDN U27587 ( .B(n27496), .A(n27497), .Z(n27494) );
  XOR U27588 ( .A(n27498), .B(n27495), .Z(n27496) );
  IV U27589 ( .A(n27463), .Z(n27460) );
  XOR U27590 ( .A(n27499), .B(n27500), .Z(n27463) );
  ANDN U27591 ( .B(n27501), .A(n27502), .Z(n27499) );
  XOR U27592 ( .A(n27500), .B(n27503), .Z(n27501) );
  XOR U27593 ( .A(n27504), .B(n27505), .Z(n27476) );
  XNOR U27594 ( .A(n27471), .B(n27506), .Z(n27505) );
  IV U27595 ( .A(n27474), .Z(n27506) );
  XOR U27596 ( .A(n27507), .B(n27508), .Z(n27474) );
  ANDN U27597 ( .B(n27509), .A(n27510), .Z(n27507) );
  XOR U27598 ( .A(n27508), .B(n27511), .Z(n27509) );
  XNOR U27599 ( .A(n27512), .B(n27513), .Z(n27471) );
  ANDN U27600 ( .B(n27514), .A(n27515), .Z(n27512) );
  XOR U27601 ( .A(n27513), .B(n27516), .Z(n27514) );
  IV U27602 ( .A(n27470), .Z(n27504) );
  XOR U27603 ( .A(n27468), .B(n27517), .Z(n27470) );
  XOR U27604 ( .A(n27518), .B(n27519), .Z(n27517) );
  ANDN U27605 ( .B(n27520), .A(n27521), .Z(n27518) );
  XOR U27606 ( .A(n27522), .B(n27519), .Z(n27520) );
  IV U27607 ( .A(n27472), .Z(n27468) );
  XOR U27608 ( .A(n27523), .B(n27524), .Z(n27472) );
  ANDN U27609 ( .B(n27525), .A(n27526), .Z(n27523) );
  XOR U27610 ( .A(n27527), .B(n27524), .Z(n27525) );
  IV U27611 ( .A(n27482), .Z(n27486) );
  XOR U27612 ( .A(n27482), .B(n27437), .Z(n27484) );
  XOR U27613 ( .A(n27528), .B(n27529), .Z(n27437) );
  AND U27614 ( .A(n674), .B(n27530), .Z(n27528) );
  XOR U27615 ( .A(n27531), .B(n27529), .Z(n27530) );
  NANDN U27616 ( .A(n27439), .B(n27441), .Z(n27482) );
  XOR U27617 ( .A(n27532), .B(n27533), .Z(n27441) );
  AND U27618 ( .A(n674), .B(n27534), .Z(n27532) );
  XOR U27619 ( .A(n27533), .B(n27535), .Z(n27534) );
  XNOR U27620 ( .A(n27536), .B(n27537), .Z(n674) );
  AND U27621 ( .A(n27538), .B(n27539), .Z(n27536) );
  XOR U27622 ( .A(n27537), .B(n27452), .Z(n27539) );
  XNOR U27623 ( .A(n27540), .B(n27541), .Z(n27452) );
  ANDN U27624 ( .B(n27542), .A(n27543), .Z(n27540) );
  XOR U27625 ( .A(n27541), .B(n27544), .Z(n27542) );
  XNOR U27626 ( .A(n27537), .B(n27454), .Z(n27538) );
  XOR U27627 ( .A(n27545), .B(n27546), .Z(n27454) );
  AND U27628 ( .A(n678), .B(n27547), .Z(n27545) );
  XOR U27629 ( .A(n27548), .B(n27546), .Z(n27547) );
  XNOR U27630 ( .A(n27549), .B(n27550), .Z(n27537) );
  AND U27631 ( .A(n27551), .B(n27552), .Z(n27549) );
  XNOR U27632 ( .A(n27550), .B(n27479), .Z(n27552) );
  XOR U27633 ( .A(n27543), .B(n27544), .Z(n27479) );
  XNOR U27634 ( .A(n27553), .B(n27554), .Z(n27544) );
  ANDN U27635 ( .B(n27555), .A(n27556), .Z(n27553) );
  XOR U27636 ( .A(n27557), .B(n27558), .Z(n27555) );
  XOR U27637 ( .A(n27559), .B(n27560), .Z(n27543) );
  XNOR U27638 ( .A(n27561), .B(n27562), .Z(n27560) );
  ANDN U27639 ( .B(n27563), .A(n27564), .Z(n27561) );
  XNOR U27640 ( .A(n27565), .B(n27566), .Z(n27563) );
  IV U27641 ( .A(n27541), .Z(n27559) );
  XOR U27642 ( .A(n27567), .B(n27568), .Z(n27541) );
  ANDN U27643 ( .B(n27569), .A(n27570), .Z(n27567) );
  XOR U27644 ( .A(n27568), .B(n27571), .Z(n27569) );
  XOR U27645 ( .A(n27550), .B(n27481), .Z(n27551) );
  XOR U27646 ( .A(n27572), .B(n27573), .Z(n27481) );
  AND U27647 ( .A(n678), .B(n27574), .Z(n27572) );
  XOR U27648 ( .A(n27575), .B(n27573), .Z(n27574) );
  XNOR U27649 ( .A(n27576), .B(n27577), .Z(n27550) );
  NAND U27650 ( .A(n27578), .B(n27579), .Z(n27577) );
  XOR U27651 ( .A(n27580), .B(n27529), .Z(n27579) );
  XOR U27652 ( .A(n27570), .B(n27571), .Z(n27529) );
  XOR U27653 ( .A(n27581), .B(n27558), .Z(n27571) );
  XOR U27654 ( .A(n27582), .B(n27583), .Z(n27558) );
  ANDN U27655 ( .B(n27584), .A(n27585), .Z(n27582) );
  XOR U27656 ( .A(n27583), .B(n27586), .Z(n27584) );
  IV U27657 ( .A(n27556), .Z(n27581) );
  XOR U27658 ( .A(n27554), .B(n27587), .Z(n27556) );
  XOR U27659 ( .A(n27588), .B(n27589), .Z(n27587) );
  ANDN U27660 ( .B(n27590), .A(n27591), .Z(n27588) );
  XOR U27661 ( .A(n27592), .B(n27589), .Z(n27590) );
  IV U27662 ( .A(n27557), .Z(n27554) );
  XOR U27663 ( .A(n27593), .B(n27594), .Z(n27557) );
  ANDN U27664 ( .B(n27595), .A(n27596), .Z(n27593) );
  XOR U27665 ( .A(n27594), .B(n27597), .Z(n27595) );
  XOR U27666 ( .A(n27598), .B(n27599), .Z(n27570) );
  XNOR U27667 ( .A(n27565), .B(n27600), .Z(n27599) );
  IV U27668 ( .A(n27568), .Z(n27600) );
  XOR U27669 ( .A(n27601), .B(n27602), .Z(n27568) );
  ANDN U27670 ( .B(n27603), .A(n27604), .Z(n27601) );
  XOR U27671 ( .A(n27602), .B(n27605), .Z(n27603) );
  XNOR U27672 ( .A(n27606), .B(n27607), .Z(n27565) );
  ANDN U27673 ( .B(n27608), .A(n27609), .Z(n27606) );
  XOR U27674 ( .A(n27607), .B(n27610), .Z(n27608) );
  IV U27675 ( .A(n27564), .Z(n27598) );
  XOR U27676 ( .A(n27562), .B(n27611), .Z(n27564) );
  XOR U27677 ( .A(n27612), .B(n27613), .Z(n27611) );
  ANDN U27678 ( .B(n27614), .A(n27615), .Z(n27612) );
  XOR U27679 ( .A(n27616), .B(n27613), .Z(n27614) );
  IV U27680 ( .A(n27566), .Z(n27562) );
  XOR U27681 ( .A(n27617), .B(n27618), .Z(n27566) );
  ANDN U27682 ( .B(n27619), .A(n27620), .Z(n27617) );
  XOR U27683 ( .A(n27621), .B(n27618), .Z(n27619) );
  IV U27684 ( .A(n27576), .Z(n27580) );
  XOR U27685 ( .A(n27576), .B(n27531), .Z(n27578) );
  XOR U27686 ( .A(n27622), .B(n27623), .Z(n27531) );
  AND U27687 ( .A(n678), .B(n27624), .Z(n27622) );
  XOR U27688 ( .A(n27625), .B(n27623), .Z(n27624) );
  NANDN U27689 ( .A(n27533), .B(n27535), .Z(n27576) );
  XOR U27690 ( .A(n27626), .B(n27627), .Z(n27535) );
  AND U27691 ( .A(n678), .B(n27628), .Z(n27626) );
  XOR U27692 ( .A(n27627), .B(n27629), .Z(n27628) );
  XNOR U27693 ( .A(n27630), .B(n27631), .Z(n678) );
  AND U27694 ( .A(n27632), .B(n27633), .Z(n27630) );
  XOR U27695 ( .A(n27631), .B(n27546), .Z(n27633) );
  XNOR U27696 ( .A(n27634), .B(n27635), .Z(n27546) );
  ANDN U27697 ( .B(n27636), .A(n27637), .Z(n27634) );
  XOR U27698 ( .A(n27635), .B(n27638), .Z(n27636) );
  XNOR U27699 ( .A(n27631), .B(n27548), .Z(n27632) );
  XOR U27700 ( .A(n27639), .B(n27640), .Z(n27548) );
  AND U27701 ( .A(n682), .B(n27641), .Z(n27639) );
  XOR U27702 ( .A(n27642), .B(n27640), .Z(n27641) );
  XNOR U27703 ( .A(n27643), .B(n27644), .Z(n27631) );
  AND U27704 ( .A(n27645), .B(n27646), .Z(n27643) );
  XNOR U27705 ( .A(n27644), .B(n27573), .Z(n27646) );
  XOR U27706 ( .A(n27637), .B(n27638), .Z(n27573) );
  XNOR U27707 ( .A(n27647), .B(n27648), .Z(n27638) );
  ANDN U27708 ( .B(n27649), .A(n27650), .Z(n27647) );
  XOR U27709 ( .A(n27651), .B(n27652), .Z(n27649) );
  XOR U27710 ( .A(n27653), .B(n27654), .Z(n27637) );
  XNOR U27711 ( .A(n27655), .B(n27656), .Z(n27654) );
  ANDN U27712 ( .B(n27657), .A(n27658), .Z(n27655) );
  XNOR U27713 ( .A(n27659), .B(n27660), .Z(n27657) );
  IV U27714 ( .A(n27635), .Z(n27653) );
  XOR U27715 ( .A(n27661), .B(n27662), .Z(n27635) );
  ANDN U27716 ( .B(n27663), .A(n27664), .Z(n27661) );
  XOR U27717 ( .A(n27662), .B(n27665), .Z(n27663) );
  XOR U27718 ( .A(n27644), .B(n27575), .Z(n27645) );
  XOR U27719 ( .A(n27666), .B(n27667), .Z(n27575) );
  AND U27720 ( .A(n682), .B(n27668), .Z(n27666) );
  XOR U27721 ( .A(n27669), .B(n27667), .Z(n27668) );
  XNOR U27722 ( .A(n27670), .B(n27671), .Z(n27644) );
  NAND U27723 ( .A(n27672), .B(n27673), .Z(n27671) );
  XOR U27724 ( .A(n27674), .B(n27623), .Z(n27673) );
  XOR U27725 ( .A(n27664), .B(n27665), .Z(n27623) );
  XOR U27726 ( .A(n27675), .B(n27652), .Z(n27665) );
  XOR U27727 ( .A(n27676), .B(n27677), .Z(n27652) );
  ANDN U27728 ( .B(n27678), .A(n27679), .Z(n27676) );
  XOR U27729 ( .A(n27677), .B(n27680), .Z(n27678) );
  IV U27730 ( .A(n27650), .Z(n27675) );
  XOR U27731 ( .A(n27648), .B(n27681), .Z(n27650) );
  XOR U27732 ( .A(n27682), .B(n27683), .Z(n27681) );
  ANDN U27733 ( .B(n27684), .A(n27685), .Z(n27682) );
  XOR U27734 ( .A(n27686), .B(n27683), .Z(n27684) );
  IV U27735 ( .A(n27651), .Z(n27648) );
  XOR U27736 ( .A(n27687), .B(n27688), .Z(n27651) );
  ANDN U27737 ( .B(n27689), .A(n27690), .Z(n27687) );
  XOR U27738 ( .A(n27688), .B(n27691), .Z(n27689) );
  XOR U27739 ( .A(n27692), .B(n27693), .Z(n27664) );
  XNOR U27740 ( .A(n27659), .B(n27694), .Z(n27693) );
  IV U27741 ( .A(n27662), .Z(n27694) );
  XOR U27742 ( .A(n27695), .B(n27696), .Z(n27662) );
  ANDN U27743 ( .B(n27697), .A(n27698), .Z(n27695) );
  XOR U27744 ( .A(n27696), .B(n27699), .Z(n27697) );
  XNOR U27745 ( .A(n27700), .B(n27701), .Z(n27659) );
  ANDN U27746 ( .B(n27702), .A(n27703), .Z(n27700) );
  XOR U27747 ( .A(n27701), .B(n27704), .Z(n27702) );
  IV U27748 ( .A(n27658), .Z(n27692) );
  XOR U27749 ( .A(n27656), .B(n27705), .Z(n27658) );
  XOR U27750 ( .A(n27706), .B(n27707), .Z(n27705) );
  ANDN U27751 ( .B(n27708), .A(n27709), .Z(n27706) );
  XOR U27752 ( .A(n27710), .B(n27707), .Z(n27708) );
  IV U27753 ( .A(n27660), .Z(n27656) );
  XOR U27754 ( .A(n27711), .B(n27712), .Z(n27660) );
  ANDN U27755 ( .B(n27713), .A(n27714), .Z(n27711) );
  XOR U27756 ( .A(n27715), .B(n27712), .Z(n27713) );
  IV U27757 ( .A(n27670), .Z(n27674) );
  XOR U27758 ( .A(n27670), .B(n27625), .Z(n27672) );
  XOR U27759 ( .A(n27716), .B(n27717), .Z(n27625) );
  AND U27760 ( .A(n682), .B(n27718), .Z(n27716) );
  XOR U27761 ( .A(n27719), .B(n27717), .Z(n27718) );
  NANDN U27762 ( .A(n27627), .B(n27629), .Z(n27670) );
  XOR U27763 ( .A(n27720), .B(n27721), .Z(n27629) );
  AND U27764 ( .A(n682), .B(n27722), .Z(n27720) );
  XOR U27765 ( .A(n27721), .B(n27723), .Z(n27722) );
  XNOR U27766 ( .A(n27724), .B(n27725), .Z(n682) );
  AND U27767 ( .A(n27726), .B(n27727), .Z(n27724) );
  XOR U27768 ( .A(n27725), .B(n27640), .Z(n27727) );
  XNOR U27769 ( .A(n27728), .B(n27729), .Z(n27640) );
  ANDN U27770 ( .B(n27730), .A(n27731), .Z(n27728) );
  XOR U27771 ( .A(n27729), .B(n27732), .Z(n27730) );
  XNOR U27772 ( .A(n27725), .B(n27642), .Z(n27726) );
  XOR U27773 ( .A(n27733), .B(n27734), .Z(n27642) );
  AND U27774 ( .A(n686), .B(n27735), .Z(n27733) );
  XOR U27775 ( .A(n27736), .B(n27734), .Z(n27735) );
  XNOR U27776 ( .A(n27737), .B(n27738), .Z(n27725) );
  AND U27777 ( .A(n27739), .B(n27740), .Z(n27737) );
  XNOR U27778 ( .A(n27738), .B(n27667), .Z(n27740) );
  XOR U27779 ( .A(n27731), .B(n27732), .Z(n27667) );
  XNOR U27780 ( .A(n27741), .B(n27742), .Z(n27732) );
  ANDN U27781 ( .B(n27743), .A(n27744), .Z(n27741) );
  XOR U27782 ( .A(n27745), .B(n27746), .Z(n27743) );
  XOR U27783 ( .A(n27747), .B(n27748), .Z(n27731) );
  XNOR U27784 ( .A(n27749), .B(n27750), .Z(n27748) );
  ANDN U27785 ( .B(n27751), .A(n27752), .Z(n27749) );
  XNOR U27786 ( .A(n27753), .B(n27754), .Z(n27751) );
  IV U27787 ( .A(n27729), .Z(n27747) );
  XOR U27788 ( .A(n27755), .B(n27756), .Z(n27729) );
  ANDN U27789 ( .B(n27757), .A(n27758), .Z(n27755) );
  XOR U27790 ( .A(n27756), .B(n27759), .Z(n27757) );
  XOR U27791 ( .A(n27738), .B(n27669), .Z(n27739) );
  XOR U27792 ( .A(n27760), .B(n27761), .Z(n27669) );
  AND U27793 ( .A(n686), .B(n27762), .Z(n27760) );
  XOR U27794 ( .A(n27763), .B(n27761), .Z(n27762) );
  XNOR U27795 ( .A(n27764), .B(n27765), .Z(n27738) );
  NAND U27796 ( .A(n27766), .B(n27767), .Z(n27765) );
  XOR U27797 ( .A(n27768), .B(n27717), .Z(n27767) );
  XOR U27798 ( .A(n27758), .B(n27759), .Z(n27717) );
  XOR U27799 ( .A(n27769), .B(n27746), .Z(n27759) );
  XOR U27800 ( .A(n27770), .B(n27771), .Z(n27746) );
  ANDN U27801 ( .B(n27772), .A(n27773), .Z(n27770) );
  XOR U27802 ( .A(n27771), .B(n27774), .Z(n27772) );
  IV U27803 ( .A(n27744), .Z(n27769) );
  XOR U27804 ( .A(n27742), .B(n27775), .Z(n27744) );
  XOR U27805 ( .A(n27776), .B(n27777), .Z(n27775) );
  ANDN U27806 ( .B(n27778), .A(n27779), .Z(n27776) );
  XOR U27807 ( .A(n27780), .B(n27777), .Z(n27778) );
  IV U27808 ( .A(n27745), .Z(n27742) );
  XOR U27809 ( .A(n27781), .B(n27782), .Z(n27745) );
  ANDN U27810 ( .B(n27783), .A(n27784), .Z(n27781) );
  XOR U27811 ( .A(n27782), .B(n27785), .Z(n27783) );
  XOR U27812 ( .A(n27786), .B(n27787), .Z(n27758) );
  XNOR U27813 ( .A(n27753), .B(n27788), .Z(n27787) );
  IV U27814 ( .A(n27756), .Z(n27788) );
  XOR U27815 ( .A(n27789), .B(n27790), .Z(n27756) );
  ANDN U27816 ( .B(n27791), .A(n27792), .Z(n27789) );
  XOR U27817 ( .A(n27790), .B(n27793), .Z(n27791) );
  XNOR U27818 ( .A(n27794), .B(n27795), .Z(n27753) );
  ANDN U27819 ( .B(n27796), .A(n27797), .Z(n27794) );
  XOR U27820 ( .A(n27795), .B(n27798), .Z(n27796) );
  IV U27821 ( .A(n27752), .Z(n27786) );
  XOR U27822 ( .A(n27750), .B(n27799), .Z(n27752) );
  XOR U27823 ( .A(n27800), .B(n27801), .Z(n27799) );
  ANDN U27824 ( .B(n27802), .A(n27803), .Z(n27800) );
  XOR U27825 ( .A(n27804), .B(n27801), .Z(n27802) );
  IV U27826 ( .A(n27754), .Z(n27750) );
  XOR U27827 ( .A(n27805), .B(n27806), .Z(n27754) );
  ANDN U27828 ( .B(n27807), .A(n27808), .Z(n27805) );
  XOR U27829 ( .A(n27809), .B(n27806), .Z(n27807) );
  IV U27830 ( .A(n27764), .Z(n27768) );
  XOR U27831 ( .A(n27764), .B(n27719), .Z(n27766) );
  XOR U27832 ( .A(n27810), .B(n27811), .Z(n27719) );
  AND U27833 ( .A(n686), .B(n27812), .Z(n27810) );
  XOR U27834 ( .A(n27813), .B(n27811), .Z(n27812) );
  NANDN U27835 ( .A(n27721), .B(n27723), .Z(n27764) );
  XOR U27836 ( .A(n27814), .B(n27815), .Z(n27723) );
  AND U27837 ( .A(n686), .B(n27816), .Z(n27814) );
  XOR U27838 ( .A(n27815), .B(n27817), .Z(n27816) );
  XNOR U27839 ( .A(n27818), .B(n27819), .Z(n686) );
  AND U27840 ( .A(n27820), .B(n27821), .Z(n27818) );
  XOR U27841 ( .A(n27819), .B(n27734), .Z(n27821) );
  XNOR U27842 ( .A(n27822), .B(n27823), .Z(n27734) );
  ANDN U27843 ( .B(n27824), .A(n27825), .Z(n27822) );
  XOR U27844 ( .A(n27823), .B(n27826), .Z(n27824) );
  XNOR U27845 ( .A(n27819), .B(n27736), .Z(n27820) );
  XOR U27846 ( .A(n27827), .B(n27828), .Z(n27736) );
  AND U27847 ( .A(n690), .B(n27829), .Z(n27827) );
  XOR U27848 ( .A(n27830), .B(n27828), .Z(n27829) );
  XNOR U27849 ( .A(n27831), .B(n27832), .Z(n27819) );
  AND U27850 ( .A(n27833), .B(n27834), .Z(n27831) );
  XNOR U27851 ( .A(n27832), .B(n27761), .Z(n27834) );
  XOR U27852 ( .A(n27825), .B(n27826), .Z(n27761) );
  XNOR U27853 ( .A(n27835), .B(n27836), .Z(n27826) );
  ANDN U27854 ( .B(n27837), .A(n27838), .Z(n27835) );
  XOR U27855 ( .A(n27839), .B(n27840), .Z(n27837) );
  XOR U27856 ( .A(n27841), .B(n27842), .Z(n27825) );
  XNOR U27857 ( .A(n27843), .B(n27844), .Z(n27842) );
  ANDN U27858 ( .B(n27845), .A(n27846), .Z(n27843) );
  XNOR U27859 ( .A(n27847), .B(n27848), .Z(n27845) );
  IV U27860 ( .A(n27823), .Z(n27841) );
  XOR U27861 ( .A(n27849), .B(n27850), .Z(n27823) );
  ANDN U27862 ( .B(n27851), .A(n27852), .Z(n27849) );
  XOR U27863 ( .A(n27850), .B(n27853), .Z(n27851) );
  XOR U27864 ( .A(n27832), .B(n27763), .Z(n27833) );
  XOR U27865 ( .A(n27854), .B(n27855), .Z(n27763) );
  AND U27866 ( .A(n690), .B(n27856), .Z(n27854) );
  XOR U27867 ( .A(n27857), .B(n27855), .Z(n27856) );
  XNOR U27868 ( .A(n27858), .B(n27859), .Z(n27832) );
  NAND U27869 ( .A(n27860), .B(n27861), .Z(n27859) );
  XOR U27870 ( .A(n27862), .B(n27811), .Z(n27861) );
  XOR U27871 ( .A(n27852), .B(n27853), .Z(n27811) );
  XOR U27872 ( .A(n27863), .B(n27840), .Z(n27853) );
  XOR U27873 ( .A(n27864), .B(n27865), .Z(n27840) );
  ANDN U27874 ( .B(n27866), .A(n27867), .Z(n27864) );
  XOR U27875 ( .A(n27865), .B(n27868), .Z(n27866) );
  IV U27876 ( .A(n27838), .Z(n27863) );
  XOR U27877 ( .A(n27836), .B(n27869), .Z(n27838) );
  XOR U27878 ( .A(n27870), .B(n27871), .Z(n27869) );
  ANDN U27879 ( .B(n27872), .A(n27873), .Z(n27870) );
  XOR U27880 ( .A(n27874), .B(n27871), .Z(n27872) );
  IV U27881 ( .A(n27839), .Z(n27836) );
  XOR U27882 ( .A(n27875), .B(n27876), .Z(n27839) );
  ANDN U27883 ( .B(n27877), .A(n27878), .Z(n27875) );
  XOR U27884 ( .A(n27876), .B(n27879), .Z(n27877) );
  XOR U27885 ( .A(n27880), .B(n27881), .Z(n27852) );
  XNOR U27886 ( .A(n27847), .B(n27882), .Z(n27881) );
  IV U27887 ( .A(n27850), .Z(n27882) );
  XOR U27888 ( .A(n27883), .B(n27884), .Z(n27850) );
  ANDN U27889 ( .B(n27885), .A(n27886), .Z(n27883) );
  XOR U27890 ( .A(n27884), .B(n27887), .Z(n27885) );
  XNOR U27891 ( .A(n27888), .B(n27889), .Z(n27847) );
  ANDN U27892 ( .B(n27890), .A(n27891), .Z(n27888) );
  XOR U27893 ( .A(n27889), .B(n27892), .Z(n27890) );
  IV U27894 ( .A(n27846), .Z(n27880) );
  XOR U27895 ( .A(n27844), .B(n27893), .Z(n27846) );
  XOR U27896 ( .A(n27894), .B(n27895), .Z(n27893) );
  ANDN U27897 ( .B(n27896), .A(n27897), .Z(n27894) );
  XOR U27898 ( .A(n27898), .B(n27895), .Z(n27896) );
  IV U27899 ( .A(n27848), .Z(n27844) );
  XOR U27900 ( .A(n27899), .B(n27900), .Z(n27848) );
  ANDN U27901 ( .B(n27901), .A(n27902), .Z(n27899) );
  XOR U27902 ( .A(n27903), .B(n27900), .Z(n27901) );
  IV U27903 ( .A(n27858), .Z(n27862) );
  XOR U27904 ( .A(n27858), .B(n27813), .Z(n27860) );
  XOR U27905 ( .A(n27904), .B(n27905), .Z(n27813) );
  AND U27906 ( .A(n690), .B(n27906), .Z(n27904) );
  XOR U27907 ( .A(n27907), .B(n27905), .Z(n27906) );
  NANDN U27908 ( .A(n27815), .B(n27817), .Z(n27858) );
  XOR U27909 ( .A(n27908), .B(n27909), .Z(n27817) );
  AND U27910 ( .A(n690), .B(n27910), .Z(n27908) );
  XOR U27911 ( .A(n27909), .B(n27911), .Z(n27910) );
  XNOR U27912 ( .A(n27912), .B(n27913), .Z(n690) );
  AND U27913 ( .A(n27914), .B(n27915), .Z(n27912) );
  XOR U27914 ( .A(n27913), .B(n27828), .Z(n27915) );
  XNOR U27915 ( .A(n27916), .B(n27917), .Z(n27828) );
  ANDN U27916 ( .B(n27918), .A(n27919), .Z(n27916) );
  XOR U27917 ( .A(n27917), .B(n27920), .Z(n27918) );
  XNOR U27918 ( .A(n27913), .B(n27830), .Z(n27914) );
  XOR U27919 ( .A(n27921), .B(n27922), .Z(n27830) );
  AND U27920 ( .A(n694), .B(n27923), .Z(n27921) );
  XOR U27921 ( .A(n27924), .B(n27922), .Z(n27923) );
  XNOR U27922 ( .A(n27925), .B(n27926), .Z(n27913) );
  AND U27923 ( .A(n27927), .B(n27928), .Z(n27925) );
  XNOR U27924 ( .A(n27926), .B(n27855), .Z(n27928) );
  XOR U27925 ( .A(n27919), .B(n27920), .Z(n27855) );
  XNOR U27926 ( .A(n27929), .B(n27930), .Z(n27920) );
  ANDN U27927 ( .B(n27931), .A(n27932), .Z(n27929) );
  XOR U27928 ( .A(n27933), .B(n27934), .Z(n27931) );
  XOR U27929 ( .A(n27935), .B(n27936), .Z(n27919) );
  XNOR U27930 ( .A(n27937), .B(n27938), .Z(n27936) );
  ANDN U27931 ( .B(n27939), .A(n27940), .Z(n27937) );
  XNOR U27932 ( .A(n27941), .B(n27942), .Z(n27939) );
  IV U27933 ( .A(n27917), .Z(n27935) );
  XOR U27934 ( .A(n27943), .B(n27944), .Z(n27917) );
  ANDN U27935 ( .B(n27945), .A(n27946), .Z(n27943) );
  XOR U27936 ( .A(n27944), .B(n27947), .Z(n27945) );
  XOR U27937 ( .A(n27926), .B(n27857), .Z(n27927) );
  XOR U27938 ( .A(n27948), .B(n27949), .Z(n27857) );
  AND U27939 ( .A(n694), .B(n27950), .Z(n27948) );
  XOR U27940 ( .A(n27951), .B(n27949), .Z(n27950) );
  XNOR U27941 ( .A(n27952), .B(n27953), .Z(n27926) );
  NAND U27942 ( .A(n27954), .B(n27955), .Z(n27953) );
  XOR U27943 ( .A(n27956), .B(n27905), .Z(n27955) );
  XOR U27944 ( .A(n27946), .B(n27947), .Z(n27905) );
  XOR U27945 ( .A(n27957), .B(n27934), .Z(n27947) );
  XOR U27946 ( .A(n27958), .B(n27959), .Z(n27934) );
  ANDN U27947 ( .B(n27960), .A(n27961), .Z(n27958) );
  XOR U27948 ( .A(n27959), .B(n27962), .Z(n27960) );
  IV U27949 ( .A(n27932), .Z(n27957) );
  XOR U27950 ( .A(n27930), .B(n27963), .Z(n27932) );
  XOR U27951 ( .A(n27964), .B(n27965), .Z(n27963) );
  ANDN U27952 ( .B(n27966), .A(n27967), .Z(n27964) );
  XOR U27953 ( .A(n27968), .B(n27965), .Z(n27966) );
  IV U27954 ( .A(n27933), .Z(n27930) );
  XOR U27955 ( .A(n27969), .B(n27970), .Z(n27933) );
  ANDN U27956 ( .B(n27971), .A(n27972), .Z(n27969) );
  XOR U27957 ( .A(n27970), .B(n27973), .Z(n27971) );
  XOR U27958 ( .A(n27974), .B(n27975), .Z(n27946) );
  XNOR U27959 ( .A(n27941), .B(n27976), .Z(n27975) );
  IV U27960 ( .A(n27944), .Z(n27976) );
  XOR U27961 ( .A(n27977), .B(n27978), .Z(n27944) );
  ANDN U27962 ( .B(n27979), .A(n27980), .Z(n27977) );
  XOR U27963 ( .A(n27978), .B(n27981), .Z(n27979) );
  XNOR U27964 ( .A(n27982), .B(n27983), .Z(n27941) );
  ANDN U27965 ( .B(n27984), .A(n27985), .Z(n27982) );
  XOR U27966 ( .A(n27983), .B(n27986), .Z(n27984) );
  IV U27967 ( .A(n27940), .Z(n27974) );
  XOR U27968 ( .A(n27938), .B(n27987), .Z(n27940) );
  XOR U27969 ( .A(n27988), .B(n27989), .Z(n27987) );
  ANDN U27970 ( .B(n27990), .A(n27991), .Z(n27988) );
  XOR U27971 ( .A(n27992), .B(n27989), .Z(n27990) );
  IV U27972 ( .A(n27942), .Z(n27938) );
  XOR U27973 ( .A(n27993), .B(n27994), .Z(n27942) );
  ANDN U27974 ( .B(n27995), .A(n27996), .Z(n27993) );
  XOR U27975 ( .A(n27997), .B(n27994), .Z(n27995) );
  IV U27976 ( .A(n27952), .Z(n27956) );
  XOR U27977 ( .A(n27952), .B(n27907), .Z(n27954) );
  XOR U27978 ( .A(n27998), .B(n27999), .Z(n27907) );
  AND U27979 ( .A(n694), .B(n28000), .Z(n27998) );
  XOR U27980 ( .A(n28001), .B(n27999), .Z(n28000) );
  NANDN U27981 ( .A(n27909), .B(n27911), .Z(n27952) );
  XOR U27982 ( .A(n28002), .B(n28003), .Z(n27911) );
  AND U27983 ( .A(n694), .B(n28004), .Z(n28002) );
  XOR U27984 ( .A(n28003), .B(n28005), .Z(n28004) );
  XNOR U27985 ( .A(n28006), .B(n28007), .Z(n694) );
  AND U27986 ( .A(n28008), .B(n28009), .Z(n28006) );
  XOR U27987 ( .A(n28007), .B(n27922), .Z(n28009) );
  XNOR U27988 ( .A(n28010), .B(n28011), .Z(n27922) );
  ANDN U27989 ( .B(n28012), .A(n28013), .Z(n28010) );
  XOR U27990 ( .A(n28011), .B(n28014), .Z(n28012) );
  XNOR U27991 ( .A(n28007), .B(n27924), .Z(n28008) );
  XOR U27992 ( .A(n28015), .B(n28016), .Z(n27924) );
  AND U27993 ( .A(n698), .B(n28017), .Z(n28015) );
  XOR U27994 ( .A(n28018), .B(n28016), .Z(n28017) );
  XNOR U27995 ( .A(n28019), .B(n28020), .Z(n28007) );
  AND U27996 ( .A(n28021), .B(n28022), .Z(n28019) );
  XNOR U27997 ( .A(n28020), .B(n27949), .Z(n28022) );
  XOR U27998 ( .A(n28013), .B(n28014), .Z(n27949) );
  XNOR U27999 ( .A(n28023), .B(n28024), .Z(n28014) );
  ANDN U28000 ( .B(n28025), .A(n28026), .Z(n28023) );
  XOR U28001 ( .A(n28027), .B(n28028), .Z(n28025) );
  XOR U28002 ( .A(n28029), .B(n28030), .Z(n28013) );
  XNOR U28003 ( .A(n28031), .B(n28032), .Z(n28030) );
  ANDN U28004 ( .B(n28033), .A(n28034), .Z(n28031) );
  XNOR U28005 ( .A(n28035), .B(n28036), .Z(n28033) );
  IV U28006 ( .A(n28011), .Z(n28029) );
  XOR U28007 ( .A(n28037), .B(n28038), .Z(n28011) );
  ANDN U28008 ( .B(n28039), .A(n28040), .Z(n28037) );
  XOR U28009 ( .A(n28038), .B(n28041), .Z(n28039) );
  XOR U28010 ( .A(n28020), .B(n27951), .Z(n28021) );
  XOR U28011 ( .A(n28042), .B(n28043), .Z(n27951) );
  AND U28012 ( .A(n698), .B(n28044), .Z(n28042) );
  XOR U28013 ( .A(n28045), .B(n28043), .Z(n28044) );
  XNOR U28014 ( .A(n28046), .B(n28047), .Z(n28020) );
  NAND U28015 ( .A(n28048), .B(n28049), .Z(n28047) );
  XOR U28016 ( .A(n28050), .B(n27999), .Z(n28049) );
  XOR U28017 ( .A(n28040), .B(n28041), .Z(n27999) );
  XOR U28018 ( .A(n28051), .B(n28028), .Z(n28041) );
  XOR U28019 ( .A(n28052), .B(n28053), .Z(n28028) );
  ANDN U28020 ( .B(n28054), .A(n28055), .Z(n28052) );
  XOR U28021 ( .A(n28053), .B(n28056), .Z(n28054) );
  IV U28022 ( .A(n28026), .Z(n28051) );
  XOR U28023 ( .A(n28024), .B(n28057), .Z(n28026) );
  XOR U28024 ( .A(n28058), .B(n28059), .Z(n28057) );
  ANDN U28025 ( .B(n28060), .A(n28061), .Z(n28058) );
  XOR U28026 ( .A(n28062), .B(n28059), .Z(n28060) );
  IV U28027 ( .A(n28027), .Z(n28024) );
  XOR U28028 ( .A(n28063), .B(n28064), .Z(n28027) );
  ANDN U28029 ( .B(n28065), .A(n28066), .Z(n28063) );
  XOR U28030 ( .A(n28064), .B(n28067), .Z(n28065) );
  XOR U28031 ( .A(n28068), .B(n28069), .Z(n28040) );
  XNOR U28032 ( .A(n28035), .B(n28070), .Z(n28069) );
  IV U28033 ( .A(n28038), .Z(n28070) );
  XOR U28034 ( .A(n28071), .B(n28072), .Z(n28038) );
  ANDN U28035 ( .B(n28073), .A(n28074), .Z(n28071) );
  XOR U28036 ( .A(n28072), .B(n28075), .Z(n28073) );
  XNOR U28037 ( .A(n28076), .B(n28077), .Z(n28035) );
  ANDN U28038 ( .B(n28078), .A(n28079), .Z(n28076) );
  XOR U28039 ( .A(n28077), .B(n28080), .Z(n28078) );
  IV U28040 ( .A(n28034), .Z(n28068) );
  XOR U28041 ( .A(n28032), .B(n28081), .Z(n28034) );
  XOR U28042 ( .A(n28082), .B(n28083), .Z(n28081) );
  ANDN U28043 ( .B(n28084), .A(n28085), .Z(n28082) );
  XOR U28044 ( .A(n28086), .B(n28083), .Z(n28084) );
  IV U28045 ( .A(n28036), .Z(n28032) );
  XOR U28046 ( .A(n28087), .B(n28088), .Z(n28036) );
  ANDN U28047 ( .B(n28089), .A(n28090), .Z(n28087) );
  XOR U28048 ( .A(n28091), .B(n28088), .Z(n28089) );
  IV U28049 ( .A(n28046), .Z(n28050) );
  XOR U28050 ( .A(n28046), .B(n28001), .Z(n28048) );
  XOR U28051 ( .A(n28092), .B(n28093), .Z(n28001) );
  AND U28052 ( .A(n698), .B(n28094), .Z(n28092) );
  XOR U28053 ( .A(n28095), .B(n28093), .Z(n28094) );
  NANDN U28054 ( .A(n28003), .B(n28005), .Z(n28046) );
  XOR U28055 ( .A(n28096), .B(n28097), .Z(n28005) );
  AND U28056 ( .A(n698), .B(n28098), .Z(n28096) );
  XOR U28057 ( .A(n28097), .B(n28099), .Z(n28098) );
  XNOR U28058 ( .A(n28100), .B(n28101), .Z(n698) );
  AND U28059 ( .A(n28102), .B(n28103), .Z(n28100) );
  XOR U28060 ( .A(n28101), .B(n28016), .Z(n28103) );
  XNOR U28061 ( .A(n28104), .B(n28105), .Z(n28016) );
  ANDN U28062 ( .B(n28106), .A(n28107), .Z(n28104) );
  XOR U28063 ( .A(n28105), .B(n28108), .Z(n28106) );
  XNOR U28064 ( .A(n28101), .B(n28018), .Z(n28102) );
  XOR U28065 ( .A(n28109), .B(n28110), .Z(n28018) );
  AND U28066 ( .A(n702), .B(n28111), .Z(n28109) );
  XOR U28067 ( .A(n28112), .B(n28110), .Z(n28111) );
  XNOR U28068 ( .A(n28113), .B(n28114), .Z(n28101) );
  AND U28069 ( .A(n28115), .B(n28116), .Z(n28113) );
  XNOR U28070 ( .A(n28114), .B(n28043), .Z(n28116) );
  XOR U28071 ( .A(n28107), .B(n28108), .Z(n28043) );
  XNOR U28072 ( .A(n28117), .B(n28118), .Z(n28108) );
  ANDN U28073 ( .B(n28119), .A(n28120), .Z(n28117) );
  XOR U28074 ( .A(n28121), .B(n28122), .Z(n28119) );
  XOR U28075 ( .A(n28123), .B(n28124), .Z(n28107) );
  XNOR U28076 ( .A(n28125), .B(n28126), .Z(n28124) );
  ANDN U28077 ( .B(n28127), .A(n28128), .Z(n28125) );
  XNOR U28078 ( .A(n28129), .B(n28130), .Z(n28127) );
  IV U28079 ( .A(n28105), .Z(n28123) );
  XOR U28080 ( .A(n28131), .B(n28132), .Z(n28105) );
  ANDN U28081 ( .B(n28133), .A(n28134), .Z(n28131) );
  XOR U28082 ( .A(n28132), .B(n28135), .Z(n28133) );
  XOR U28083 ( .A(n28114), .B(n28045), .Z(n28115) );
  XOR U28084 ( .A(n28136), .B(n28137), .Z(n28045) );
  AND U28085 ( .A(n702), .B(n28138), .Z(n28136) );
  XOR U28086 ( .A(n28139), .B(n28137), .Z(n28138) );
  XNOR U28087 ( .A(n28140), .B(n28141), .Z(n28114) );
  NAND U28088 ( .A(n28142), .B(n28143), .Z(n28141) );
  XOR U28089 ( .A(n28144), .B(n28093), .Z(n28143) );
  XOR U28090 ( .A(n28134), .B(n28135), .Z(n28093) );
  XOR U28091 ( .A(n28145), .B(n28122), .Z(n28135) );
  XOR U28092 ( .A(n28146), .B(n28147), .Z(n28122) );
  ANDN U28093 ( .B(n28148), .A(n28149), .Z(n28146) );
  XOR U28094 ( .A(n28147), .B(n28150), .Z(n28148) );
  IV U28095 ( .A(n28120), .Z(n28145) );
  XOR U28096 ( .A(n28118), .B(n28151), .Z(n28120) );
  XOR U28097 ( .A(n28152), .B(n28153), .Z(n28151) );
  ANDN U28098 ( .B(n28154), .A(n28155), .Z(n28152) );
  XOR U28099 ( .A(n28156), .B(n28153), .Z(n28154) );
  IV U28100 ( .A(n28121), .Z(n28118) );
  XOR U28101 ( .A(n28157), .B(n28158), .Z(n28121) );
  ANDN U28102 ( .B(n28159), .A(n28160), .Z(n28157) );
  XOR U28103 ( .A(n28158), .B(n28161), .Z(n28159) );
  XOR U28104 ( .A(n28162), .B(n28163), .Z(n28134) );
  XNOR U28105 ( .A(n28129), .B(n28164), .Z(n28163) );
  IV U28106 ( .A(n28132), .Z(n28164) );
  XOR U28107 ( .A(n28165), .B(n28166), .Z(n28132) );
  ANDN U28108 ( .B(n28167), .A(n28168), .Z(n28165) );
  XOR U28109 ( .A(n28166), .B(n28169), .Z(n28167) );
  XNOR U28110 ( .A(n28170), .B(n28171), .Z(n28129) );
  ANDN U28111 ( .B(n28172), .A(n28173), .Z(n28170) );
  XOR U28112 ( .A(n28171), .B(n28174), .Z(n28172) );
  IV U28113 ( .A(n28128), .Z(n28162) );
  XOR U28114 ( .A(n28126), .B(n28175), .Z(n28128) );
  XOR U28115 ( .A(n28176), .B(n28177), .Z(n28175) );
  ANDN U28116 ( .B(n28178), .A(n28179), .Z(n28176) );
  XOR U28117 ( .A(n28180), .B(n28177), .Z(n28178) );
  IV U28118 ( .A(n28130), .Z(n28126) );
  XOR U28119 ( .A(n28181), .B(n28182), .Z(n28130) );
  ANDN U28120 ( .B(n28183), .A(n28184), .Z(n28181) );
  XOR U28121 ( .A(n28185), .B(n28182), .Z(n28183) );
  IV U28122 ( .A(n28140), .Z(n28144) );
  XOR U28123 ( .A(n28140), .B(n28095), .Z(n28142) );
  XOR U28124 ( .A(n28186), .B(n28187), .Z(n28095) );
  AND U28125 ( .A(n702), .B(n28188), .Z(n28186) );
  XOR U28126 ( .A(n28189), .B(n28187), .Z(n28188) );
  NANDN U28127 ( .A(n28097), .B(n28099), .Z(n28140) );
  XOR U28128 ( .A(n28190), .B(n28191), .Z(n28099) );
  AND U28129 ( .A(n702), .B(n28192), .Z(n28190) );
  XOR U28130 ( .A(n28191), .B(n28193), .Z(n28192) );
  XNOR U28131 ( .A(n28194), .B(n28195), .Z(n702) );
  AND U28132 ( .A(n28196), .B(n28197), .Z(n28194) );
  XOR U28133 ( .A(n28195), .B(n28110), .Z(n28197) );
  XNOR U28134 ( .A(n28198), .B(n28199), .Z(n28110) );
  ANDN U28135 ( .B(n28200), .A(n28201), .Z(n28198) );
  XOR U28136 ( .A(n28199), .B(n28202), .Z(n28200) );
  XNOR U28137 ( .A(n28195), .B(n28112), .Z(n28196) );
  XOR U28138 ( .A(n28203), .B(n28204), .Z(n28112) );
  AND U28139 ( .A(n706), .B(n28205), .Z(n28203) );
  XOR U28140 ( .A(n28206), .B(n28204), .Z(n28205) );
  XNOR U28141 ( .A(n28207), .B(n28208), .Z(n28195) );
  AND U28142 ( .A(n28209), .B(n28210), .Z(n28207) );
  XNOR U28143 ( .A(n28208), .B(n28137), .Z(n28210) );
  XOR U28144 ( .A(n28201), .B(n28202), .Z(n28137) );
  XNOR U28145 ( .A(n28211), .B(n28212), .Z(n28202) );
  ANDN U28146 ( .B(n28213), .A(n28214), .Z(n28211) );
  XOR U28147 ( .A(n28215), .B(n28216), .Z(n28213) );
  XOR U28148 ( .A(n28217), .B(n28218), .Z(n28201) );
  XNOR U28149 ( .A(n28219), .B(n28220), .Z(n28218) );
  ANDN U28150 ( .B(n28221), .A(n28222), .Z(n28219) );
  XNOR U28151 ( .A(n28223), .B(n28224), .Z(n28221) );
  IV U28152 ( .A(n28199), .Z(n28217) );
  XOR U28153 ( .A(n28225), .B(n28226), .Z(n28199) );
  ANDN U28154 ( .B(n28227), .A(n28228), .Z(n28225) );
  XOR U28155 ( .A(n28226), .B(n28229), .Z(n28227) );
  XOR U28156 ( .A(n28208), .B(n28139), .Z(n28209) );
  XOR U28157 ( .A(n28230), .B(n28231), .Z(n28139) );
  AND U28158 ( .A(n706), .B(n28232), .Z(n28230) );
  XOR U28159 ( .A(n28233), .B(n28231), .Z(n28232) );
  XNOR U28160 ( .A(n28234), .B(n28235), .Z(n28208) );
  NAND U28161 ( .A(n28236), .B(n28237), .Z(n28235) );
  XOR U28162 ( .A(n28238), .B(n28187), .Z(n28237) );
  XOR U28163 ( .A(n28228), .B(n28229), .Z(n28187) );
  XOR U28164 ( .A(n28239), .B(n28216), .Z(n28229) );
  XOR U28165 ( .A(n28240), .B(n28241), .Z(n28216) );
  ANDN U28166 ( .B(n28242), .A(n28243), .Z(n28240) );
  XOR U28167 ( .A(n28241), .B(n28244), .Z(n28242) );
  IV U28168 ( .A(n28214), .Z(n28239) );
  XOR U28169 ( .A(n28212), .B(n28245), .Z(n28214) );
  XOR U28170 ( .A(n28246), .B(n28247), .Z(n28245) );
  ANDN U28171 ( .B(n28248), .A(n28249), .Z(n28246) );
  XOR U28172 ( .A(n28250), .B(n28247), .Z(n28248) );
  IV U28173 ( .A(n28215), .Z(n28212) );
  XOR U28174 ( .A(n28251), .B(n28252), .Z(n28215) );
  ANDN U28175 ( .B(n28253), .A(n28254), .Z(n28251) );
  XOR U28176 ( .A(n28252), .B(n28255), .Z(n28253) );
  XOR U28177 ( .A(n28256), .B(n28257), .Z(n28228) );
  XNOR U28178 ( .A(n28223), .B(n28258), .Z(n28257) );
  IV U28179 ( .A(n28226), .Z(n28258) );
  XOR U28180 ( .A(n28259), .B(n28260), .Z(n28226) );
  ANDN U28181 ( .B(n28261), .A(n28262), .Z(n28259) );
  XOR U28182 ( .A(n28260), .B(n28263), .Z(n28261) );
  XNOR U28183 ( .A(n28264), .B(n28265), .Z(n28223) );
  ANDN U28184 ( .B(n28266), .A(n28267), .Z(n28264) );
  XOR U28185 ( .A(n28265), .B(n28268), .Z(n28266) );
  IV U28186 ( .A(n28222), .Z(n28256) );
  XOR U28187 ( .A(n28220), .B(n28269), .Z(n28222) );
  XOR U28188 ( .A(n28270), .B(n28271), .Z(n28269) );
  ANDN U28189 ( .B(n28272), .A(n28273), .Z(n28270) );
  XOR U28190 ( .A(n28274), .B(n28271), .Z(n28272) );
  IV U28191 ( .A(n28224), .Z(n28220) );
  XOR U28192 ( .A(n28275), .B(n28276), .Z(n28224) );
  ANDN U28193 ( .B(n28277), .A(n28278), .Z(n28275) );
  XOR U28194 ( .A(n28279), .B(n28276), .Z(n28277) );
  IV U28195 ( .A(n28234), .Z(n28238) );
  XOR U28196 ( .A(n28234), .B(n28189), .Z(n28236) );
  XOR U28197 ( .A(n28280), .B(n28281), .Z(n28189) );
  AND U28198 ( .A(n706), .B(n28282), .Z(n28280) );
  XOR U28199 ( .A(n28283), .B(n28281), .Z(n28282) );
  NANDN U28200 ( .A(n28191), .B(n28193), .Z(n28234) );
  XOR U28201 ( .A(n28284), .B(n28285), .Z(n28193) );
  AND U28202 ( .A(n706), .B(n28286), .Z(n28284) );
  XOR U28203 ( .A(n28285), .B(n28287), .Z(n28286) );
  XNOR U28204 ( .A(n28288), .B(n28289), .Z(n706) );
  AND U28205 ( .A(n28290), .B(n28291), .Z(n28288) );
  XOR U28206 ( .A(n28289), .B(n28204), .Z(n28291) );
  XNOR U28207 ( .A(n28292), .B(n28293), .Z(n28204) );
  ANDN U28208 ( .B(n28294), .A(n28295), .Z(n28292) );
  XOR U28209 ( .A(n28293), .B(n28296), .Z(n28294) );
  XNOR U28210 ( .A(n28289), .B(n28206), .Z(n28290) );
  XOR U28211 ( .A(n28297), .B(n28298), .Z(n28206) );
  AND U28212 ( .A(n710), .B(n28299), .Z(n28297) );
  XOR U28213 ( .A(n28300), .B(n28298), .Z(n28299) );
  XNOR U28214 ( .A(n28301), .B(n28302), .Z(n28289) );
  AND U28215 ( .A(n28303), .B(n28304), .Z(n28301) );
  XNOR U28216 ( .A(n28302), .B(n28231), .Z(n28304) );
  XOR U28217 ( .A(n28295), .B(n28296), .Z(n28231) );
  XNOR U28218 ( .A(n28305), .B(n28306), .Z(n28296) );
  ANDN U28219 ( .B(n28307), .A(n28308), .Z(n28305) );
  XOR U28220 ( .A(n28309), .B(n28310), .Z(n28307) );
  XOR U28221 ( .A(n28311), .B(n28312), .Z(n28295) );
  XNOR U28222 ( .A(n28313), .B(n28314), .Z(n28312) );
  ANDN U28223 ( .B(n28315), .A(n28316), .Z(n28313) );
  XNOR U28224 ( .A(n28317), .B(n28318), .Z(n28315) );
  IV U28225 ( .A(n28293), .Z(n28311) );
  XOR U28226 ( .A(n28319), .B(n28320), .Z(n28293) );
  ANDN U28227 ( .B(n28321), .A(n28322), .Z(n28319) );
  XOR U28228 ( .A(n28320), .B(n28323), .Z(n28321) );
  XOR U28229 ( .A(n28302), .B(n28233), .Z(n28303) );
  XOR U28230 ( .A(n28324), .B(n28325), .Z(n28233) );
  AND U28231 ( .A(n710), .B(n28326), .Z(n28324) );
  XOR U28232 ( .A(n28327), .B(n28325), .Z(n28326) );
  XNOR U28233 ( .A(n28328), .B(n28329), .Z(n28302) );
  NAND U28234 ( .A(n28330), .B(n28331), .Z(n28329) );
  XOR U28235 ( .A(n28332), .B(n28281), .Z(n28331) );
  XOR U28236 ( .A(n28322), .B(n28323), .Z(n28281) );
  XOR U28237 ( .A(n28333), .B(n28310), .Z(n28323) );
  XOR U28238 ( .A(n28334), .B(n28335), .Z(n28310) );
  ANDN U28239 ( .B(n28336), .A(n28337), .Z(n28334) );
  XOR U28240 ( .A(n28335), .B(n28338), .Z(n28336) );
  IV U28241 ( .A(n28308), .Z(n28333) );
  XOR U28242 ( .A(n28306), .B(n28339), .Z(n28308) );
  XOR U28243 ( .A(n28340), .B(n28341), .Z(n28339) );
  ANDN U28244 ( .B(n28342), .A(n28343), .Z(n28340) );
  XOR U28245 ( .A(n28344), .B(n28341), .Z(n28342) );
  IV U28246 ( .A(n28309), .Z(n28306) );
  XOR U28247 ( .A(n28345), .B(n28346), .Z(n28309) );
  ANDN U28248 ( .B(n28347), .A(n28348), .Z(n28345) );
  XOR U28249 ( .A(n28346), .B(n28349), .Z(n28347) );
  XOR U28250 ( .A(n28350), .B(n28351), .Z(n28322) );
  XNOR U28251 ( .A(n28317), .B(n28352), .Z(n28351) );
  IV U28252 ( .A(n28320), .Z(n28352) );
  XOR U28253 ( .A(n28353), .B(n28354), .Z(n28320) );
  ANDN U28254 ( .B(n28355), .A(n28356), .Z(n28353) );
  XOR U28255 ( .A(n28354), .B(n28357), .Z(n28355) );
  XNOR U28256 ( .A(n28358), .B(n28359), .Z(n28317) );
  ANDN U28257 ( .B(n28360), .A(n28361), .Z(n28358) );
  XOR U28258 ( .A(n28359), .B(n28362), .Z(n28360) );
  IV U28259 ( .A(n28316), .Z(n28350) );
  XOR U28260 ( .A(n28314), .B(n28363), .Z(n28316) );
  XOR U28261 ( .A(n28364), .B(n28365), .Z(n28363) );
  ANDN U28262 ( .B(n28366), .A(n28367), .Z(n28364) );
  XOR U28263 ( .A(n28368), .B(n28365), .Z(n28366) );
  IV U28264 ( .A(n28318), .Z(n28314) );
  XOR U28265 ( .A(n28369), .B(n28370), .Z(n28318) );
  ANDN U28266 ( .B(n28371), .A(n28372), .Z(n28369) );
  XOR U28267 ( .A(n28373), .B(n28370), .Z(n28371) );
  IV U28268 ( .A(n28328), .Z(n28332) );
  XOR U28269 ( .A(n28328), .B(n28283), .Z(n28330) );
  XOR U28270 ( .A(n28374), .B(n28375), .Z(n28283) );
  AND U28271 ( .A(n710), .B(n28376), .Z(n28374) );
  XOR U28272 ( .A(n28377), .B(n28375), .Z(n28376) );
  NANDN U28273 ( .A(n28285), .B(n28287), .Z(n28328) );
  XOR U28274 ( .A(n28378), .B(n28379), .Z(n28287) );
  AND U28275 ( .A(n710), .B(n28380), .Z(n28378) );
  XOR U28276 ( .A(n28379), .B(n28381), .Z(n28380) );
  XNOR U28277 ( .A(n28382), .B(n28383), .Z(n710) );
  AND U28278 ( .A(n28384), .B(n28385), .Z(n28382) );
  XOR U28279 ( .A(n28383), .B(n28298), .Z(n28385) );
  XNOR U28280 ( .A(n28386), .B(n28387), .Z(n28298) );
  ANDN U28281 ( .B(n28388), .A(n28389), .Z(n28386) );
  XOR U28282 ( .A(n28387), .B(n28390), .Z(n28388) );
  XNOR U28283 ( .A(n28383), .B(n28300), .Z(n28384) );
  XOR U28284 ( .A(n28391), .B(n28392), .Z(n28300) );
  AND U28285 ( .A(n714), .B(n28393), .Z(n28391) );
  XOR U28286 ( .A(n28394), .B(n28392), .Z(n28393) );
  XNOR U28287 ( .A(n28395), .B(n28396), .Z(n28383) );
  AND U28288 ( .A(n28397), .B(n28398), .Z(n28395) );
  XNOR U28289 ( .A(n28396), .B(n28325), .Z(n28398) );
  XOR U28290 ( .A(n28389), .B(n28390), .Z(n28325) );
  XNOR U28291 ( .A(n28399), .B(n28400), .Z(n28390) );
  ANDN U28292 ( .B(n28401), .A(n28402), .Z(n28399) );
  XOR U28293 ( .A(n28403), .B(n28404), .Z(n28401) );
  XOR U28294 ( .A(n28405), .B(n28406), .Z(n28389) );
  XNOR U28295 ( .A(n28407), .B(n28408), .Z(n28406) );
  ANDN U28296 ( .B(n28409), .A(n28410), .Z(n28407) );
  XNOR U28297 ( .A(n28411), .B(n28412), .Z(n28409) );
  IV U28298 ( .A(n28387), .Z(n28405) );
  XOR U28299 ( .A(n28413), .B(n28414), .Z(n28387) );
  ANDN U28300 ( .B(n28415), .A(n28416), .Z(n28413) );
  XOR U28301 ( .A(n28414), .B(n28417), .Z(n28415) );
  XOR U28302 ( .A(n28396), .B(n28327), .Z(n28397) );
  XOR U28303 ( .A(n28418), .B(n28419), .Z(n28327) );
  AND U28304 ( .A(n714), .B(n28420), .Z(n28418) );
  XOR U28305 ( .A(n28421), .B(n28419), .Z(n28420) );
  XNOR U28306 ( .A(n28422), .B(n28423), .Z(n28396) );
  NAND U28307 ( .A(n28424), .B(n28425), .Z(n28423) );
  XOR U28308 ( .A(n28426), .B(n28375), .Z(n28425) );
  XOR U28309 ( .A(n28416), .B(n28417), .Z(n28375) );
  XOR U28310 ( .A(n28427), .B(n28404), .Z(n28417) );
  XOR U28311 ( .A(n28428), .B(n28429), .Z(n28404) );
  ANDN U28312 ( .B(n28430), .A(n28431), .Z(n28428) );
  XOR U28313 ( .A(n28429), .B(n28432), .Z(n28430) );
  IV U28314 ( .A(n28402), .Z(n28427) );
  XOR U28315 ( .A(n28400), .B(n28433), .Z(n28402) );
  XOR U28316 ( .A(n28434), .B(n28435), .Z(n28433) );
  ANDN U28317 ( .B(n28436), .A(n28437), .Z(n28434) );
  XOR U28318 ( .A(n28438), .B(n28435), .Z(n28436) );
  IV U28319 ( .A(n28403), .Z(n28400) );
  XOR U28320 ( .A(n28439), .B(n28440), .Z(n28403) );
  ANDN U28321 ( .B(n28441), .A(n28442), .Z(n28439) );
  XOR U28322 ( .A(n28440), .B(n28443), .Z(n28441) );
  XOR U28323 ( .A(n28444), .B(n28445), .Z(n28416) );
  XNOR U28324 ( .A(n28411), .B(n28446), .Z(n28445) );
  IV U28325 ( .A(n28414), .Z(n28446) );
  XOR U28326 ( .A(n28447), .B(n28448), .Z(n28414) );
  ANDN U28327 ( .B(n28449), .A(n28450), .Z(n28447) );
  XOR U28328 ( .A(n28448), .B(n28451), .Z(n28449) );
  XNOR U28329 ( .A(n28452), .B(n28453), .Z(n28411) );
  ANDN U28330 ( .B(n28454), .A(n28455), .Z(n28452) );
  XOR U28331 ( .A(n28453), .B(n28456), .Z(n28454) );
  IV U28332 ( .A(n28410), .Z(n28444) );
  XOR U28333 ( .A(n28408), .B(n28457), .Z(n28410) );
  XOR U28334 ( .A(n28458), .B(n28459), .Z(n28457) );
  ANDN U28335 ( .B(n28460), .A(n28461), .Z(n28458) );
  XOR U28336 ( .A(n28462), .B(n28459), .Z(n28460) );
  IV U28337 ( .A(n28412), .Z(n28408) );
  XOR U28338 ( .A(n28463), .B(n28464), .Z(n28412) );
  ANDN U28339 ( .B(n28465), .A(n28466), .Z(n28463) );
  XOR U28340 ( .A(n28467), .B(n28464), .Z(n28465) );
  IV U28341 ( .A(n28422), .Z(n28426) );
  XOR U28342 ( .A(n28422), .B(n28377), .Z(n28424) );
  XOR U28343 ( .A(n28468), .B(n28469), .Z(n28377) );
  AND U28344 ( .A(n714), .B(n28470), .Z(n28468) );
  XOR U28345 ( .A(n28471), .B(n28469), .Z(n28470) );
  NANDN U28346 ( .A(n28379), .B(n28381), .Z(n28422) );
  XOR U28347 ( .A(n28472), .B(n28473), .Z(n28381) );
  AND U28348 ( .A(n714), .B(n28474), .Z(n28472) );
  XOR U28349 ( .A(n28473), .B(n28475), .Z(n28474) );
  XNOR U28350 ( .A(n28476), .B(n28477), .Z(n714) );
  AND U28351 ( .A(n28478), .B(n28479), .Z(n28476) );
  XOR U28352 ( .A(n28477), .B(n28392), .Z(n28479) );
  XNOR U28353 ( .A(n28480), .B(n28481), .Z(n28392) );
  ANDN U28354 ( .B(n28482), .A(n28483), .Z(n28480) );
  XOR U28355 ( .A(n28481), .B(n28484), .Z(n28482) );
  XNOR U28356 ( .A(n28477), .B(n28394), .Z(n28478) );
  XOR U28357 ( .A(n28485), .B(n28486), .Z(n28394) );
  AND U28358 ( .A(n718), .B(n28487), .Z(n28485) );
  XOR U28359 ( .A(n28488), .B(n28486), .Z(n28487) );
  XNOR U28360 ( .A(n28489), .B(n28490), .Z(n28477) );
  AND U28361 ( .A(n28491), .B(n28492), .Z(n28489) );
  XNOR U28362 ( .A(n28490), .B(n28419), .Z(n28492) );
  XOR U28363 ( .A(n28483), .B(n28484), .Z(n28419) );
  XNOR U28364 ( .A(n28493), .B(n28494), .Z(n28484) );
  ANDN U28365 ( .B(n28495), .A(n28496), .Z(n28493) );
  XOR U28366 ( .A(n28497), .B(n28498), .Z(n28495) );
  XOR U28367 ( .A(n28499), .B(n28500), .Z(n28483) );
  XNOR U28368 ( .A(n28501), .B(n28502), .Z(n28500) );
  ANDN U28369 ( .B(n28503), .A(n28504), .Z(n28501) );
  XNOR U28370 ( .A(n28505), .B(n28506), .Z(n28503) );
  IV U28371 ( .A(n28481), .Z(n28499) );
  XOR U28372 ( .A(n28507), .B(n28508), .Z(n28481) );
  ANDN U28373 ( .B(n28509), .A(n28510), .Z(n28507) );
  XOR U28374 ( .A(n28508), .B(n28511), .Z(n28509) );
  XOR U28375 ( .A(n28490), .B(n28421), .Z(n28491) );
  XOR U28376 ( .A(n28512), .B(n28513), .Z(n28421) );
  AND U28377 ( .A(n718), .B(n28514), .Z(n28512) );
  XOR U28378 ( .A(n28515), .B(n28513), .Z(n28514) );
  XNOR U28379 ( .A(n28516), .B(n28517), .Z(n28490) );
  NAND U28380 ( .A(n28518), .B(n28519), .Z(n28517) );
  XOR U28381 ( .A(n28520), .B(n28469), .Z(n28519) );
  XOR U28382 ( .A(n28510), .B(n28511), .Z(n28469) );
  XOR U28383 ( .A(n28521), .B(n28498), .Z(n28511) );
  XOR U28384 ( .A(n28522), .B(n28523), .Z(n28498) );
  ANDN U28385 ( .B(n28524), .A(n28525), .Z(n28522) );
  XOR U28386 ( .A(n28523), .B(n28526), .Z(n28524) );
  IV U28387 ( .A(n28496), .Z(n28521) );
  XOR U28388 ( .A(n28494), .B(n28527), .Z(n28496) );
  XOR U28389 ( .A(n28528), .B(n28529), .Z(n28527) );
  ANDN U28390 ( .B(n28530), .A(n28531), .Z(n28528) );
  XOR U28391 ( .A(n28532), .B(n28529), .Z(n28530) );
  IV U28392 ( .A(n28497), .Z(n28494) );
  XOR U28393 ( .A(n28533), .B(n28534), .Z(n28497) );
  ANDN U28394 ( .B(n28535), .A(n28536), .Z(n28533) );
  XOR U28395 ( .A(n28534), .B(n28537), .Z(n28535) );
  XOR U28396 ( .A(n28538), .B(n28539), .Z(n28510) );
  XNOR U28397 ( .A(n28505), .B(n28540), .Z(n28539) );
  IV U28398 ( .A(n28508), .Z(n28540) );
  XOR U28399 ( .A(n28541), .B(n28542), .Z(n28508) );
  ANDN U28400 ( .B(n28543), .A(n28544), .Z(n28541) );
  XOR U28401 ( .A(n28542), .B(n28545), .Z(n28543) );
  XNOR U28402 ( .A(n28546), .B(n28547), .Z(n28505) );
  ANDN U28403 ( .B(n28548), .A(n28549), .Z(n28546) );
  XOR U28404 ( .A(n28547), .B(n28550), .Z(n28548) );
  IV U28405 ( .A(n28504), .Z(n28538) );
  XOR U28406 ( .A(n28502), .B(n28551), .Z(n28504) );
  XOR U28407 ( .A(n28552), .B(n28553), .Z(n28551) );
  ANDN U28408 ( .B(n28554), .A(n28555), .Z(n28552) );
  XOR U28409 ( .A(n28556), .B(n28553), .Z(n28554) );
  IV U28410 ( .A(n28506), .Z(n28502) );
  XOR U28411 ( .A(n28557), .B(n28558), .Z(n28506) );
  ANDN U28412 ( .B(n28559), .A(n28560), .Z(n28557) );
  XOR U28413 ( .A(n28561), .B(n28558), .Z(n28559) );
  IV U28414 ( .A(n28516), .Z(n28520) );
  XOR U28415 ( .A(n28516), .B(n28471), .Z(n28518) );
  XOR U28416 ( .A(n28562), .B(n28563), .Z(n28471) );
  AND U28417 ( .A(n718), .B(n28564), .Z(n28562) );
  XOR U28418 ( .A(n28565), .B(n28563), .Z(n28564) );
  NANDN U28419 ( .A(n28473), .B(n28475), .Z(n28516) );
  XOR U28420 ( .A(n28566), .B(n28567), .Z(n28475) );
  AND U28421 ( .A(n718), .B(n28568), .Z(n28566) );
  XOR U28422 ( .A(n28567), .B(n28569), .Z(n28568) );
  XNOR U28423 ( .A(n28570), .B(n28571), .Z(n718) );
  AND U28424 ( .A(n28572), .B(n28573), .Z(n28570) );
  XOR U28425 ( .A(n28571), .B(n28486), .Z(n28573) );
  XNOR U28426 ( .A(n28574), .B(n28575), .Z(n28486) );
  ANDN U28427 ( .B(n28576), .A(n28577), .Z(n28574) );
  XOR U28428 ( .A(n28575), .B(n28578), .Z(n28576) );
  XNOR U28429 ( .A(n28571), .B(n28488), .Z(n28572) );
  XOR U28430 ( .A(n28579), .B(n28580), .Z(n28488) );
  AND U28431 ( .A(n722), .B(n28581), .Z(n28579) );
  XOR U28432 ( .A(n28582), .B(n28580), .Z(n28581) );
  XNOR U28433 ( .A(n28583), .B(n28584), .Z(n28571) );
  AND U28434 ( .A(n28585), .B(n28586), .Z(n28583) );
  XNOR U28435 ( .A(n28584), .B(n28513), .Z(n28586) );
  XOR U28436 ( .A(n28577), .B(n28578), .Z(n28513) );
  XNOR U28437 ( .A(n28587), .B(n28588), .Z(n28578) );
  ANDN U28438 ( .B(n28589), .A(n28590), .Z(n28587) );
  XOR U28439 ( .A(n28591), .B(n28592), .Z(n28589) );
  XOR U28440 ( .A(n28593), .B(n28594), .Z(n28577) );
  XNOR U28441 ( .A(n28595), .B(n28596), .Z(n28594) );
  ANDN U28442 ( .B(n28597), .A(n28598), .Z(n28595) );
  XNOR U28443 ( .A(n28599), .B(n28600), .Z(n28597) );
  IV U28444 ( .A(n28575), .Z(n28593) );
  XOR U28445 ( .A(n28601), .B(n28602), .Z(n28575) );
  ANDN U28446 ( .B(n28603), .A(n28604), .Z(n28601) );
  XOR U28447 ( .A(n28602), .B(n28605), .Z(n28603) );
  XOR U28448 ( .A(n28584), .B(n28515), .Z(n28585) );
  XOR U28449 ( .A(n28606), .B(n28607), .Z(n28515) );
  AND U28450 ( .A(n722), .B(n28608), .Z(n28606) );
  XOR U28451 ( .A(n28609), .B(n28607), .Z(n28608) );
  XNOR U28452 ( .A(n28610), .B(n28611), .Z(n28584) );
  NAND U28453 ( .A(n28612), .B(n28613), .Z(n28611) );
  XOR U28454 ( .A(n28614), .B(n28563), .Z(n28613) );
  XOR U28455 ( .A(n28604), .B(n28605), .Z(n28563) );
  XOR U28456 ( .A(n28615), .B(n28592), .Z(n28605) );
  XOR U28457 ( .A(n28616), .B(n28617), .Z(n28592) );
  ANDN U28458 ( .B(n28618), .A(n28619), .Z(n28616) );
  XOR U28459 ( .A(n28617), .B(n28620), .Z(n28618) );
  IV U28460 ( .A(n28590), .Z(n28615) );
  XOR U28461 ( .A(n28588), .B(n28621), .Z(n28590) );
  XOR U28462 ( .A(n28622), .B(n28623), .Z(n28621) );
  ANDN U28463 ( .B(n28624), .A(n28625), .Z(n28622) );
  XOR U28464 ( .A(n28626), .B(n28623), .Z(n28624) );
  IV U28465 ( .A(n28591), .Z(n28588) );
  XOR U28466 ( .A(n28627), .B(n28628), .Z(n28591) );
  ANDN U28467 ( .B(n28629), .A(n28630), .Z(n28627) );
  XOR U28468 ( .A(n28628), .B(n28631), .Z(n28629) );
  XOR U28469 ( .A(n28632), .B(n28633), .Z(n28604) );
  XNOR U28470 ( .A(n28599), .B(n28634), .Z(n28633) );
  IV U28471 ( .A(n28602), .Z(n28634) );
  XOR U28472 ( .A(n28635), .B(n28636), .Z(n28602) );
  ANDN U28473 ( .B(n28637), .A(n28638), .Z(n28635) );
  XOR U28474 ( .A(n28636), .B(n28639), .Z(n28637) );
  XNOR U28475 ( .A(n28640), .B(n28641), .Z(n28599) );
  ANDN U28476 ( .B(n28642), .A(n28643), .Z(n28640) );
  XOR U28477 ( .A(n28641), .B(n28644), .Z(n28642) );
  IV U28478 ( .A(n28598), .Z(n28632) );
  XOR U28479 ( .A(n28596), .B(n28645), .Z(n28598) );
  XOR U28480 ( .A(n28646), .B(n28647), .Z(n28645) );
  ANDN U28481 ( .B(n28648), .A(n28649), .Z(n28646) );
  XOR U28482 ( .A(n28650), .B(n28647), .Z(n28648) );
  IV U28483 ( .A(n28600), .Z(n28596) );
  XOR U28484 ( .A(n28651), .B(n28652), .Z(n28600) );
  ANDN U28485 ( .B(n28653), .A(n28654), .Z(n28651) );
  XOR U28486 ( .A(n28655), .B(n28652), .Z(n28653) );
  IV U28487 ( .A(n28610), .Z(n28614) );
  XOR U28488 ( .A(n28610), .B(n28565), .Z(n28612) );
  XOR U28489 ( .A(n28656), .B(n28657), .Z(n28565) );
  AND U28490 ( .A(n722), .B(n28658), .Z(n28656) );
  XOR U28491 ( .A(n28659), .B(n28657), .Z(n28658) );
  NANDN U28492 ( .A(n28567), .B(n28569), .Z(n28610) );
  XOR U28493 ( .A(n28660), .B(n28661), .Z(n28569) );
  AND U28494 ( .A(n722), .B(n28662), .Z(n28660) );
  XOR U28495 ( .A(n28661), .B(n28663), .Z(n28662) );
  XNOR U28496 ( .A(n28664), .B(n28665), .Z(n722) );
  AND U28497 ( .A(n28666), .B(n28667), .Z(n28664) );
  XOR U28498 ( .A(n28665), .B(n28580), .Z(n28667) );
  XNOR U28499 ( .A(n28668), .B(n28669), .Z(n28580) );
  ANDN U28500 ( .B(n28670), .A(n28671), .Z(n28668) );
  XOR U28501 ( .A(n28669), .B(n28672), .Z(n28670) );
  XNOR U28502 ( .A(n28665), .B(n28582), .Z(n28666) );
  XOR U28503 ( .A(n28673), .B(n28674), .Z(n28582) );
  AND U28504 ( .A(n726), .B(n28675), .Z(n28673) );
  XOR U28505 ( .A(n28676), .B(n28674), .Z(n28675) );
  XNOR U28506 ( .A(n28677), .B(n28678), .Z(n28665) );
  AND U28507 ( .A(n28679), .B(n28680), .Z(n28677) );
  XNOR U28508 ( .A(n28678), .B(n28607), .Z(n28680) );
  XOR U28509 ( .A(n28671), .B(n28672), .Z(n28607) );
  XNOR U28510 ( .A(n28681), .B(n28682), .Z(n28672) );
  ANDN U28511 ( .B(n28683), .A(n28684), .Z(n28681) );
  XOR U28512 ( .A(n28685), .B(n28686), .Z(n28683) );
  XOR U28513 ( .A(n28687), .B(n28688), .Z(n28671) );
  XNOR U28514 ( .A(n28689), .B(n28690), .Z(n28688) );
  ANDN U28515 ( .B(n28691), .A(n28692), .Z(n28689) );
  XNOR U28516 ( .A(n28693), .B(n28694), .Z(n28691) );
  IV U28517 ( .A(n28669), .Z(n28687) );
  XOR U28518 ( .A(n28695), .B(n28696), .Z(n28669) );
  ANDN U28519 ( .B(n28697), .A(n28698), .Z(n28695) );
  XOR U28520 ( .A(n28696), .B(n28699), .Z(n28697) );
  XOR U28521 ( .A(n28678), .B(n28609), .Z(n28679) );
  XOR U28522 ( .A(n28700), .B(n28701), .Z(n28609) );
  AND U28523 ( .A(n726), .B(n28702), .Z(n28700) );
  XOR U28524 ( .A(n28703), .B(n28701), .Z(n28702) );
  XNOR U28525 ( .A(n28704), .B(n28705), .Z(n28678) );
  NAND U28526 ( .A(n28706), .B(n28707), .Z(n28705) );
  XOR U28527 ( .A(n28708), .B(n28657), .Z(n28707) );
  XOR U28528 ( .A(n28698), .B(n28699), .Z(n28657) );
  XOR U28529 ( .A(n28709), .B(n28686), .Z(n28699) );
  XOR U28530 ( .A(n28710), .B(n28711), .Z(n28686) );
  ANDN U28531 ( .B(n28712), .A(n28713), .Z(n28710) );
  XOR U28532 ( .A(n28711), .B(n28714), .Z(n28712) );
  IV U28533 ( .A(n28684), .Z(n28709) );
  XOR U28534 ( .A(n28682), .B(n28715), .Z(n28684) );
  XOR U28535 ( .A(n28716), .B(n28717), .Z(n28715) );
  ANDN U28536 ( .B(n28718), .A(n28719), .Z(n28716) );
  XOR U28537 ( .A(n28720), .B(n28717), .Z(n28718) );
  IV U28538 ( .A(n28685), .Z(n28682) );
  XOR U28539 ( .A(n28721), .B(n28722), .Z(n28685) );
  ANDN U28540 ( .B(n28723), .A(n28724), .Z(n28721) );
  XOR U28541 ( .A(n28722), .B(n28725), .Z(n28723) );
  XOR U28542 ( .A(n28726), .B(n28727), .Z(n28698) );
  XNOR U28543 ( .A(n28693), .B(n28728), .Z(n28727) );
  IV U28544 ( .A(n28696), .Z(n28728) );
  XOR U28545 ( .A(n28729), .B(n28730), .Z(n28696) );
  ANDN U28546 ( .B(n28731), .A(n28732), .Z(n28729) );
  XOR U28547 ( .A(n28730), .B(n28733), .Z(n28731) );
  XNOR U28548 ( .A(n28734), .B(n28735), .Z(n28693) );
  ANDN U28549 ( .B(n28736), .A(n28737), .Z(n28734) );
  XOR U28550 ( .A(n28735), .B(n28738), .Z(n28736) );
  IV U28551 ( .A(n28692), .Z(n28726) );
  XOR U28552 ( .A(n28690), .B(n28739), .Z(n28692) );
  XOR U28553 ( .A(n28740), .B(n28741), .Z(n28739) );
  ANDN U28554 ( .B(n28742), .A(n28743), .Z(n28740) );
  XOR U28555 ( .A(n28744), .B(n28741), .Z(n28742) );
  IV U28556 ( .A(n28694), .Z(n28690) );
  XOR U28557 ( .A(n28745), .B(n28746), .Z(n28694) );
  ANDN U28558 ( .B(n28747), .A(n28748), .Z(n28745) );
  XOR U28559 ( .A(n28749), .B(n28746), .Z(n28747) );
  IV U28560 ( .A(n28704), .Z(n28708) );
  XOR U28561 ( .A(n28704), .B(n28659), .Z(n28706) );
  XOR U28562 ( .A(n28750), .B(n28751), .Z(n28659) );
  AND U28563 ( .A(n726), .B(n28752), .Z(n28750) );
  XOR U28564 ( .A(n28753), .B(n28751), .Z(n28752) );
  NANDN U28565 ( .A(n28661), .B(n28663), .Z(n28704) );
  XOR U28566 ( .A(n28754), .B(n28755), .Z(n28663) );
  AND U28567 ( .A(n726), .B(n28756), .Z(n28754) );
  XOR U28568 ( .A(n28755), .B(n28757), .Z(n28756) );
  XNOR U28569 ( .A(n28758), .B(n28759), .Z(n726) );
  AND U28570 ( .A(n28760), .B(n28761), .Z(n28758) );
  XOR U28571 ( .A(n28759), .B(n28674), .Z(n28761) );
  XNOR U28572 ( .A(n28762), .B(n28763), .Z(n28674) );
  ANDN U28573 ( .B(n28764), .A(n28765), .Z(n28762) );
  XOR U28574 ( .A(n28763), .B(n28766), .Z(n28764) );
  XNOR U28575 ( .A(n28759), .B(n28676), .Z(n28760) );
  XOR U28576 ( .A(n28767), .B(n28768), .Z(n28676) );
  AND U28577 ( .A(n730), .B(n28769), .Z(n28767) );
  XOR U28578 ( .A(n28770), .B(n28768), .Z(n28769) );
  XNOR U28579 ( .A(n28771), .B(n28772), .Z(n28759) );
  AND U28580 ( .A(n28773), .B(n28774), .Z(n28771) );
  XNOR U28581 ( .A(n28772), .B(n28701), .Z(n28774) );
  XOR U28582 ( .A(n28765), .B(n28766), .Z(n28701) );
  XNOR U28583 ( .A(n28775), .B(n28776), .Z(n28766) );
  ANDN U28584 ( .B(n28777), .A(n28778), .Z(n28775) );
  XOR U28585 ( .A(n28779), .B(n28780), .Z(n28777) );
  XOR U28586 ( .A(n28781), .B(n28782), .Z(n28765) );
  XNOR U28587 ( .A(n28783), .B(n28784), .Z(n28782) );
  ANDN U28588 ( .B(n28785), .A(n28786), .Z(n28783) );
  XNOR U28589 ( .A(n28787), .B(n28788), .Z(n28785) );
  IV U28590 ( .A(n28763), .Z(n28781) );
  XOR U28591 ( .A(n28789), .B(n28790), .Z(n28763) );
  ANDN U28592 ( .B(n28791), .A(n28792), .Z(n28789) );
  XOR U28593 ( .A(n28790), .B(n28793), .Z(n28791) );
  XOR U28594 ( .A(n28772), .B(n28703), .Z(n28773) );
  XOR U28595 ( .A(n28794), .B(n28795), .Z(n28703) );
  AND U28596 ( .A(n730), .B(n28796), .Z(n28794) );
  XOR U28597 ( .A(n28797), .B(n28795), .Z(n28796) );
  XNOR U28598 ( .A(n28798), .B(n28799), .Z(n28772) );
  NAND U28599 ( .A(n28800), .B(n28801), .Z(n28799) );
  XOR U28600 ( .A(n28802), .B(n28751), .Z(n28801) );
  XOR U28601 ( .A(n28792), .B(n28793), .Z(n28751) );
  XOR U28602 ( .A(n28803), .B(n28780), .Z(n28793) );
  XOR U28603 ( .A(n28804), .B(n28805), .Z(n28780) );
  ANDN U28604 ( .B(n28806), .A(n28807), .Z(n28804) );
  XOR U28605 ( .A(n28805), .B(n28808), .Z(n28806) );
  IV U28606 ( .A(n28778), .Z(n28803) );
  XOR U28607 ( .A(n28776), .B(n28809), .Z(n28778) );
  XOR U28608 ( .A(n28810), .B(n28811), .Z(n28809) );
  ANDN U28609 ( .B(n28812), .A(n28813), .Z(n28810) );
  XOR U28610 ( .A(n28814), .B(n28811), .Z(n28812) );
  IV U28611 ( .A(n28779), .Z(n28776) );
  XOR U28612 ( .A(n28815), .B(n28816), .Z(n28779) );
  ANDN U28613 ( .B(n28817), .A(n28818), .Z(n28815) );
  XOR U28614 ( .A(n28816), .B(n28819), .Z(n28817) );
  XOR U28615 ( .A(n28820), .B(n28821), .Z(n28792) );
  XNOR U28616 ( .A(n28787), .B(n28822), .Z(n28821) );
  IV U28617 ( .A(n28790), .Z(n28822) );
  XOR U28618 ( .A(n28823), .B(n28824), .Z(n28790) );
  ANDN U28619 ( .B(n28825), .A(n28826), .Z(n28823) );
  XOR U28620 ( .A(n28824), .B(n28827), .Z(n28825) );
  XNOR U28621 ( .A(n28828), .B(n28829), .Z(n28787) );
  ANDN U28622 ( .B(n28830), .A(n28831), .Z(n28828) );
  XOR U28623 ( .A(n28829), .B(n28832), .Z(n28830) );
  IV U28624 ( .A(n28786), .Z(n28820) );
  XOR U28625 ( .A(n28784), .B(n28833), .Z(n28786) );
  XOR U28626 ( .A(n28834), .B(n28835), .Z(n28833) );
  ANDN U28627 ( .B(n28836), .A(n28837), .Z(n28834) );
  XOR U28628 ( .A(n28838), .B(n28835), .Z(n28836) );
  IV U28629 ( .A(n28788), .Z(n28784) );
  XOR U28630 ( .A(n28839), .B(n28840), .Z(n28788) );
  ANDN U28631 ( .B(n28841), .A(n28842), .Z(n28839) );
  XOR U28632 ( .A(n28843), .B(n28840), .Z(n28841) );
  IV U28633 ( .A(n28798), .Z(n28802) );
  XOR U28634 ( .A(n28798), .B(n28753), .Z(n28800) );
  XOR U28635 ( .A(n28844), .B(n28845), .Z(n28753) );
  AND U28636 ( .A(n730), .B(n28846), .Z(n28844) );
  XOR U28637 ( .A(n28847), .B(n28845), .Z(n28846) );
  NANDN U28638 ( .A(n28755), .B(n28757), .Z(n28798) );
  XOR U28639 ( .A(n28848), .B(n28849), .Z(n28757) );
  AND U28640 ( .A(n730), .B(n28850), .Z(n28848) );
  XOR U28641 ( .A(n28849), .B(n28851), .Z(n28850) );
  XNOR U28642 ( .A(n28852), .B(n28853), .Z(n730) );
  AND U28643 ( .A(n28854), .B(n28855), .Z(n28852) );
  XOR U28644 ( .A(n28853), .B(n28768), .Z(n28855) );
  XNOR U28645 ( .A(n28856), .B(n28857), .Z(n28768) );
  ANDN U28646 ( .B(n28858), .A(n28859), .Z(n28856) );
  XOR U28647 ( .A(n28857), .B(n28860), .Z(n28858) );
  XNOR U28648 ( .A(n28853), .B(n28770), .Z(n28854) );
  XOR U28649 ( .A(n28861), .B(n28862), .Z(n28770) );
  AND U28650 ( .A(n734), .B(n28863), .Z(n28861) );
  XOR U28651 ( .A(n28864), .B(n28862), .Z(n28863) );
  XNOR U28652 ( .A(n28865), .B(n28866), .Z(n28853) );
  AND U28653 ( .A(n28867), .B(n28868), .Z(n28865) );
  XNOR U28654 ( .A(n28866), .B(n28795), .Z(n28868) );
  XOR U28655 ( .A(n28859), .B(n28860), .Z(n28795) );
  XNOR U28656 ( .A(n28869), .B(n28870), .Z(n28860) );
  ANDN U28657 ( .B(n28871), .A(n28872), .Z(n28869) );
  XOR U28658 ( .A(n28873), .B(n28874), .Z(n28871) );
  XOR U28659 ( .A(n28875), .B(n28876), .Z(n28859) );
  XNOR U28660 ( .A(n28877), .B(n28878), .Z(n28876) );
  ANDN U28661 ( .B(n28879), .A(n28880), .Z(n28877) );
  XNOR U28662 ( .A(n28881), .B(n28882), .Z(n28879) );
  IV U28663 ( .A(n28857), .Z(n28875) );
  XOR U28664 ( .A(n28883), .B(n28884), .Z(n28857) );
  ANDN U28665 ( .B(n28885), .A(n28886), .Z(n28883) );
  XOR U28666 ( .A(n28884), .B(n28887), .Z(n28885) );
  XOR U28667 ( .A(n28866), .B(n28797), .Z(n28867) );
  XOR U28668 ( .A(n28888), .B(n28889), .Z(n28797) );
  AND U28669 ( .A(n734), .B(n28890), .Z(n28888) );
  XOR U28670 ( .A(n28891), .B(n28889), .Z(n28890) );
  XNOR U28671 ( .A(n28892), .B(n28893), .Z(n28866) );
  NAND U28672 ( .A(n28894), .B(n28895), .Z(n28893) );
  XOR U28673 ( .A(n28896), .B(n28845), .Z(n28895) );
  XOR U28674 ( .A(n28886), .B(n28887), .Z(n28845) );
  XOR U28675 ( .A(n28897), .B(n28874), .Z(n28887) );
  XOR U28676 ( .A(n28898), .B(n28899), .Z(n28874) );
  ANDN U28677 ( .B(n28900), .A(n28901), .Z(n28898) );
  XOR U28678 ( .A(n28899), .B(n28902), .Z(n28900) );
  IV U28679 ( .A(n28872), .Z(n28897) );
  XOR U28680 ( .A(n28870), .B(n28903), .Z(n28872) );
  XOR U28681 ( .A(n28904), .B(n28905), .Z(n28903) );
  ANDN U28682 ( .B(n28906), .A(n28907), .Z(n28904) );
  XOR U28683 ( .A(n28908), .B(n28905), .Z(n28906) );
  IV U28684 ( .A(n28873), .Z(n28870) );
  XOR U28685 ( .A(n28909), .B(n28910), .Z(n28873) );
  ANDN U28686 ( .B(n28911), .A(n28912), .Z(n28909) );
  XOR U28687 ( .A(n28910), .B(n28913), .Z(n28911) );
  XOR U28688 ( .A(n28914), .B(n28915), .Z(n28886) );
  XNOR U28689 ( .A(n28881), .B(n28916), .Z(n28915) );
  IV U28690 ( .A(n28884), .Z(n28916) );
  XOR U28691 ( .A(n28917), .B(n28918), .Z(n28884) );
  ANDN U28692 ( .B(n28919), .A(n28920), .Z(n28917) );
  XOR U28693 ( .A(n28918), .B(n28921), .Z(n28919) );
  XNOR U28694 ( .A(n28922), .B(n28923), .Z(n28881) );
  ANDN U28695 ( .B(n28924), .A(n28925), .Z(n28922) );
  XOR U28696 ( .A(n28923), .B(n28926), .Z(n28924) );
  IV U28697 ( .A(n28880), .Z(n28914) );
  XOR U28698 ( .A(n28878), .B(n28927), .Z(n28880) );
  XOR U28699 ( .A(n28928), .B(n28929), .Z(n28927) );
  ANDN U28700 ( .B(n28930), .A(n28931), .Z(n28928) );
  XOR U28701 ( .A(n28932), .B(n28929), .Z(n28930) );
  IV U28702 ( .A(n28882), .Z(n28878) );
  XOR U28703 ( .A(n28933), .B(n28934), .Z(n28882) );
  ANDN U28704 ( .B(n28935), .A(n28936), .Z(n28933) );
  XOR U28705 ( .A(n28937), .B(n28934), .Z(n28935) );
  IV U28706 ( .A(n28892), .Z(n28896) );
  XOR U28707 ( .A(n28892), .B(n28847), .Z(n28894) );
  XOR U28708 ( .A(n28938), .B(n28939), .Z(n28847) );
  AND U28709 ( .A(n734), .B(n28940), .Z(n28938) );
  XOR U28710 ( .A(n28941), .B(n28939), .Z(n28940) );
  NANDN U28711 ( .A(n28849), .B(n28851), .Z(n28892) );
  XOR U28712 ( .A(n28942), .B(n28943), .Z(n28851) );
  AND U28713 ( .A(n734), .B(n28944), .Z(n28942) );
  XOR U28714 ( .A(n28943), .B(n28945), .Z(n28944) );
  XNOR U28715 ( .A(n28946), .B(n28947), .Z(n734) );
  AND U28716 ( .A(n28948), .B(n28949), .Z(n28946) );
  XOR U28717 ( .A(n28947), .B(n28862), .Z(n28949) );
  XNOR U28718 ( .A(n28950), .B(n28951), .Z(n28862) );
  ANDN U28719 ( .B(n28952), .A(n28953), .Z(n28950) );
  XOR U28720 ( .A(n28951), .B(n28954), .Z(n28952) );
  XNOR U28721 ( .A(n28947), .B(n28864), .Z(n28948) );
  XOR U28722 ( .A(n28955), .B(n28956), .Z(n28864) );
  AND U28723 ( .A(n738), .B(n28957), .Z(n28955) );
  XOR U28724 ( .A(n28958), .B(n28956), .Z(n28957) );
  XNOR U28725 ( .A(n28959), .B(n28960), .Z(n28947) );
  AND U28726 ( .A(n28961), .B(n28962), .Z(n28959) );
  XNOR U28727 ( .A(n28960), .B(n28889), .Z(n28962) );
  XOR U28728 ( .A(n28953), .B(n28954), .Z(n28889) );
  XNOR U28729 ( .A(n28963), .B(n28964), .Z(n28954) );
  ANDN U28730 ( .B(n28965), .A(n28966), .Z(n28963) );
  XOR U28731 ( .A(n28967), .B(n28968), .Z(n28965) );
  XOR U28732 ( .A(n28969), .B(n28970), .Z(n28953) );
  XNOR U28733 ( .A(n28971), .B(n28972), .Z(n28970) );
  ANDN U28734 ( .B(n28973), .A(n28974), .Z(n28971) );
  XNOR U28735 ( .A(n28975), .B(n28976), .Z(n28973) );
  IV U28736 ( .A(n28951), .Z(n28969) );
  XOR U28737 ( .A(n28977), .B(n28978), .Z(n28951) );
  ANDN U28738 ( .B(n28979), .A(n28980), .Z(n28977) );
  XOR U28739 ( .A(n28978), .B(n28981), .Z(n28979) );
  XOR U28740 ( .A(n28960), .B(n28891), .Z(n28961) );
  XOR U28741 ( .A(n28982), .B(n28983), .Z(n28891) );
  AND U28742 ( .A(n738), .B(n28984), .Z(n28982) );
  XOR U28743 ( .A(n28985), .B(n28983), .Z(n28984) );
  XNOR U28744 ( .A(n28986), .B(n28987), .Z(n28960) );
  NAND U28745 ( .A(n28988), .B(n28989), .Z(n28987) );
  XOR U28746 ( .A(n28990), .B(n28939), .Z(n28989) );
  XOR U28747 ( .A(n28980), .B(n28981), .Z(n28939) );
  XOR U28748 ( .A(n28991), .B(n28968), .Z(n28981) );
  XOR U28749 ( .A(n28992), .B(n28993), .Z(n28968) );
  ANDN U28750 ( .B(n28994), .A(n28995), .Z(n28992) );
  XOR U28751 ( .A(n28993), .B(n28996), .Z(n28994) );
  IV U28752 ( .A(n28966), .Z(n28991) );
  XOR U28753 ( .A(n28964), .B(n28997), .Z(n28966) );
  XOR U28754 ( .A(n28998), .B(n28999), .Z(n28997) );
  ANDN U28755 ( .B(n29000), .A(n29001), .Z(n28998) );
  XOR U28756 ( .A(n29002), .B(n28999), .Z(n29000) );
  IV U28757 ( .A(n28967), .Z(n28964) );
  XOR U28758 ( .A(n29003), .B(n29004), .Z(n28967) );
  ANDN U28759 ( .B(n29005), .A(n29006), .Z(n29003) );
  XOR U28760 ( .A(n29004), .B(n29007), .Z(n29005) );
  XOR U28761 ( .A(n29008), .B(n29009), .Z(n28980) );
  XNOR U28762 ( .A(n28975), .B(n29010), .Z(n29009) );
  IV U28763 ( .A(n28978), .Z(n29010) );
  XOR U28764 ( .A(n29011), .B(n29012), .Z(n28978) );
  ANDN U28765 ( .B(n29013), .A(n29014), .Z(n29011) );
  XOR U28766 ( .A(n29012), .B(n29015), .Z(n29013) );
  XNOR U28767 ( .A(n29016), .B(n29017), .Z(n28975) );
  ANDN U28768 ( .B(n29018), .A(n29019), .Z(n29016) );
  XOR U28769 ( .A(n29017), .B(n29020), .Z(n29018) );
  IV U28770 ( .A(n28974), .Z(n29008) );
  XOR U28771 ( .A(n28972), .B(n29021), .Z(n28974) );
  XOR U28772 ( .A(n29022), .B(n29023), .Z(n29021) );
  ANDN U28773 ( .B(n29024), .A(n29025), .Z(n29022) );
  XOR U28774 ( .A(n29026), .B(n29023), .Z(n29024) );
  IV U28775 ( .A(n28976), .Z(n28972) );
  XOR U28776 ( .A(n29027), .B(n29028), .Z(n28976) );
  ANDN U28777 ( .B(n29029), .A(n29030), .Z(n29027) );
  XOR U28778 ( .A(n29031), .B(n29028), .Z(n29029) );
  IV U28779 ( .A(n28986), .Z(n28990) );
  XOR U28780 ( .A(n28986), .B(n28941), .Z(n28988) );
  XOR U28781 ( .A(n29032), .B(n29033), .Z(n28941) );
  AND U28782 ( .A(n738), .B(n29034), .Z(n29032) );
  XOR U28783 ( .A(n29035), .B(n29033), .Z(n29034) );
  NANDN U28784 ( .A(n28943), .B(n28945), .Z(n28986) );
  XOR U28785 ( .A(n29036), .B(n29037), .Z(n28945) );
  AND U28786 ( .A(n738), .B(n29038), .Z(n29036) );
  XOR U28787 ( .A(n29037), .B(n29039), .Z(n29038) );
  XNOR U28788 ( .A(n29040), .B(n29041), .Z(n738) );
  AND U28789 ( .A(n29042), .B(n29043), .Z(n29040) );
  XOR U28790 ( .A(n29041), .B(n28956), .Z(n29043) );
  XNOR U28791 ( .A(n29044), .B(n29045), .Z(n28956) );
  ANDN U28792 ( .B(n29046), .A(n29047), .Z(n29044) );
  XOR U28793 ( .A(n29045), .B(n29048), .Z(n29046) );
  XNOR U28794 ( .A(n29041), .B(n28958), .Z(n29042) );
  XOR U28795 ( .A(n29049), .B(n29050), .Z(n28958) );
  AND U28796 ( .A(n742), .B(n29051), .Z(n29049) );
  XOR U28797 ( .A(n29052), .B(n29050), .Z(n29051) );
  XNOR U28798 ( .A(n29053), .B(n29054), .Z(n29041) );
  AND U28799 ( .A(n29055), .B(n29056), .Z(n29053) );
  XNOR U28800 ( .A(n29054), .B(n28983), .Z(n29056) );
  XOR U28801 ( .A(n29047), .B(n29048), .Z(n28983) );
  XNOR U28802 ( .A(n29057), .B(n29058), .Z(n29048) );
  ANDN U28803 ( .B(n29059), .A(n29060), .Z(n29057) );
  XOR U28804 ( .A(n29061), .B(n29062), .Z(n29059) );
  XOR U28805 ( .A(n29063), .B(n29064), .Z(n29047) );
  XNOR U28806 ( .A(n29065), .B(n29066), .Z(n29064) );
  ANDN U28807 ( .B(n29067), .A(n29068), .Z(n29065) );
  XNOR U28808 ( .A(n29069), .B(n29070), .Z(n29067) );
  IV U28809 ( .A(n29045), .Z(n29063) );
  XOR U28810 ( .A(n29071), .B(n29072), .Z(n29045) );
  ANDN U28811 ( .B(n29073), .A(n29074), .Z(n29071) );
  XOR U28812 ( .A(n29072), .B(n29075), .Z(n29073) );
  XOR U28813 ( .A(n29054), .B(n28985), .Z(n29055) );
  XOR U28814 ( .A(n29076), .B(n29077), .Z(n28985) );
  AND U28815 ( .A(n742), .B(n29078), .Z(n29076) );
  XOR U28816 ( .A(n29079), .B(n29077), .Z(n29078) );
  XNOR U28817 ( .A(n29080), .B(n29081), .Z(n29054) );
  NAND U28818 ( .A(n29082), .B(n29083), .Z(n29081) );
  XOR U28819 ( .A(n29084), .B(n29033), .Z(n29083) );
  XOR U28820 ( .A(n29074), .B(n29075), .Z(n29033) );
  XOR U28821 ( .A(n29085), .B(n29062), .Z(n29075) );
  XOR U28822 ( .A(n29086), .B(n29087), .Z(n29062) );
  ANDN U28823 ( .B(n29088), .A(n29089), .Z(n29086) );
  XOR U28824 ( .A(n29087), .B(n29090), .Z(n29088) );
  IV U28825 ( .A(n29060), .Z(n29085) );
  XOR U28826 ( .A(n29058), .B(n29091), .Z(n29060) );
  XOR U28827 ( .A(n29092), .B(n29093), .Z(n29091) );
  ANDN U28828 ( .B(n29094), .A(n29095), .Z(n29092) );
  XOR U28829 ( .A(n29096), .B(n29093), .Z(n29094) );
  IV U28830 ( .A(n29061), .Z(n29058) );
  XOR U28831 ( .A(n29097), .B(n29098), .Z(n29061) );
  ANDN U28832 ( .B(n29099), .A(n29100), .Z(n29097) );
  XOR U28833 ( .A(n29098), .B(n29101), .Z(n29099) );
  XOR U28834 ( .A(n29102), .B(n29103), .Z(n29074) );
  XNOR U28835 ( .A(n29069), .B(n29104), .Z(n29103) );
  IV U28836 ( .A(n29072), .Z(n29104) );
  XOR U28837 ( .A(n29105), .B(n29106), .Z(n29072) );
  ANDN U28838 ( .B(n29107), .A(n29108), .Z(n29105) );
  XOR U28839 ( .A(n29106), .B(n29109), .Z(n29107) );
  XNOR U28840 ( .A(n29110), .B(n29111), .Z(n29069) );
  ANDN U28841 ( .B(n29112), .A(n29113), .Z(n29110) );
  XOR U28842 ( .A(n29111), .B(n29114), .Z(n29112) );
  IV U28843 ( .A(n29068), .Z(n29102) );
  XOR U28844 ( .A(n29066), .B(n29115), .Z(n29068) );
  XOR U28845 ( .A(n29116), .B(n29117), .Z(n29115) );
  ANDN U28846 ( .B(n29118), .A(n29119), .Z(n29116) );
  XOR U28847 ( .A(n29120), .B(n29117), .Z(n29118) );
  IV U28848 ( .A(n29070), .Z(n29066) );
  XOR U28849 ( .A(n29121), .B(n29122), .Z(n29070) );
  ANDN U28850 ( .B(n29123), .A(n29124), .Z(n29121) );
  XOR U28851 ( .A(n29125), .B(n29122), .Z(n29123) );
  IV U28852 ( .A(n29080), .Z(n29084) );
  XOR U28853 ( .A(n29080), .B(n29035), .Z(n29082) );
  XOR U28854 ( .A(n29126), .B(n29127), .Z(n29035) );
  AND U28855 ( .A(n742), .B(n29128), .Z(n29126) );
  XOR U28856 ( .A(n29129), .B(n29127), .Z(n29128) );
  NANDN U28857 ( .A(n29037), .B(n29039), .Z(n29080) );
  XOR U28858 ( .A(n29130), .B(n29131), .Z(n29039) );
  AND U28859 ( .A(n742), .B(n29132), .Z(n29130) );
  XOR U28860 ( .A(n29131), .B(n29133), .Z(n29132) );
  XNOR U28861 ( .A(n29134), .B(n29135), .Z(n742) );
  AND U28862 ( .A(n29136), .B(n29137), .Z(n29134) );
  XOR U28863 ( .A(n29135), .B(n29050), .Z(n29137) );
  XNOR U28864 ( .A(n29138), .B(n29139), .Z(n29050) );
  ANDN U28865 ( .B(n29140), .A(n29141), .Z(n29138) );
  XOR U28866 ( .A(n29139), .B(n29142), .Z(n29140) );
  XNOR U28867 ( .A(n29135), .B(n29052), .Z(n29136) );
  XOR U28868 ( .A(n29143), .B(n29144), .Z(n29052) );
  AND U28869 ( .A(n746), .B(n29145), .Z(n29143) );
  XOR U28870 ( .A(n29146), .B(n29144), .Z(n29145) );
  XNOR U28871 ( .A(n29147), .B(n29148), .Z(n29135) );
  AND U28872 ( .A(n29149), .B(n29150), .Z(n29147) );
  XNOR U28873 ( .A(n29148), .B(n29077), .Z(n29150) );
  XOR U28874 ( .A(n29141), .B(n29142), .Z(n29077) );
  XNOR U28875 ( .A(n29151), .B(n29152), .Z(n29142) );
  ANDN U28876 ( .B(n29153), .A(n29154), .Z(n29151) );
  XOR U28877 ( .A(n29155), .B(n29156), .Z(n29153) );
  XOR U28878 ( .A(n29157), .B(n29158), .Z(n29141) );
  XNOR U28879 ( .A(n29159), .B(n29160), .Z(n29158) );
  ANDN U28880 ( .B(n29161), .A(n29162), .Z(n29159) );
  XNOR U28881 ( .A(n29163), .B(n29164), .Z(n29161) );
  IV U28882 ( .A(n29139), .Z(n29157) );
  XOR U28883 ( .A(n29165), .B(n29166), .Z(n29139) );
  ANDN U28884 ( .B(n29167), .A(n29168), .Z(n29165) );
  XOR U28885 ( .A(n29166), .B(n29169), .Z(n29167) );
  XOR U28886 ( .A(n29148), .B(n29079), .Z(n29149) );
  XOR U28887 ( .A(n29170), .B(n29171), .Z(n29079) );
  AND U28888 ( .A(n746), .B(n29172), .Z(n29170) );
  XOR U28889 ( .A(n29173), .B(n29171), .Z(n29172) );
  XNOR U28890 ( .A(n29174), .B(n29175), .Z(n29148) );
  NAND U28891 ( .A(n29176), .B(n29177), .Z(n29175) );
  XOR U28892 ( .A(n29178), .B(n29127), .Z(n29177) );
  XOR U28893 ( .A(n29168), .B(n29169), .Z(n29127) );
  XOR U28894 ( .A(n29179), .B(n29156), .Z(n29169) );
  XOR U28895 ( .A(n29180), .B(n29181), .Z(n29156) );
  ANDN U28896 ( .B(n29182), .A(n29183), .Z(n29180) );
  XOR U28897 ( .A(n29181), .B(n29184), .Z(n29182) );
  IV U28898 ( .A(n29154), .Z(n29179) );
  XOR U28899 ( .A(n29152), .B(n29185), .Z(n29154) );
  XOR U28900 ( .A(n29186), .B(n29187), .Z(n29185) );
  ANDN U28901 ( .B(n29188), .A(n29189), .Z(n29186) );
  XOR U28902 ( .A(n29190), .B(n29187), .Z(n29188) );
  IV U28903 ( .A(n29155), .Z(n29152) );
  XOR U28904 ( .A(n29191), .B(n29192), .Z(n29155) );
  ANDN U28905 ( .B(n29193), .A(n29194), .Z(n29191) );
  XOR U28906 ( .A(n29192), .B(n29195), .Z(n29193) );
  XOR U28907 ( .A(n29196), .B(n29197), .Z(n29168) );
  XNOR U28908 ( .A(n29163), .B(n29198), .Z(n29197) );
  IV U28909 ( .A(n29166), .Z(n29198) );
  XOR U28910 ( .A(n29199), .B(n29200), .Z(n29166) );
  ANDN U28911 ( .B(n29201), .A(n29202), .Z(n29199) );
  XOR U28912 ( .A(n29200), .B(n29203), .Z(n29201) );
  XNOR U28913 ( .A(n29204), .B(n29205), .Z(n29163) );
  ANDN U28914 ( .B(n29206), .A(n29207), .Z(n29204) );
  XOR U28915 ( .A(n29205), .B(n29208), .Z(n29206) );
  IV U28916 ( .A(n29162), .Z(n29196) );
  XOR U28917 ( .A(n29160), .B(n29209), .Z(n29162) );
  XOR U28918 ( .A(n29210), .B(n29211), .Z(n29209) );
  ANDN U28919 ( .B(n29212), .A(n29213), .Z(n29210) );
  XOR U28920 ( .A(n29214), .B(n29211), .Z(n29212) );
  IV U28921 ( .A(n29164), .Z(n29160) );
  XOR U28922 ( .A(n29215), .B(n29216), .Z(n29164) );
  ANDN U28923 ( .B(n29217), .A(n29218), .Z(n29215) );
  XOR U28924 ( .A(n29219), .B(n29216), .Z(n29217) );
  IV U28925 ( .A(n29174), .Z(n29178) );
  XOR U28926 ( .A(n29174), .B(n29129), .Z(n29176) );
  XOR U28927 ( .A(n29220), .B(n29221), .Z(n29129) );
  AND U28928 ( .A(n746), .B(n29222), .Z(n29220) );
  XOR U28929 ( .A(n29223), .B(n29221), .Z(n29222) );
  NANDN U28930 ( .A(n29131), .B(n29133), .Z(n29174) );
  XOR U28931 ( .A(n29224), .B(n29225), .Z(n29133) );
  AND U28932 ( .A(n746), .B(n29226), .Z(n29224) );
  XOR U28933 ( .A(n29225), .B(n29227), .Z(n29226) );
  XNOR U28934 ( .A(n29228), .B(n29229), .Z(n746) );
  AND U28935 ( .A(n29230), .B(n29231), .Z(n29228) );
  XOR U28936 ( .A(n29229), .B(n29144), .Z(n29231) );
  XNOR U28937 ( .A(n29232), .B(n29233), .Z(n29144) );
  ANDN U28938 ( .B(n29234), .A(n29235), .Z(n29232) );
  XOR U28939 ( .A(n29233), .B(n29236), .Z(n29234) );
  XNOR U28940 ( .A(n29229), .B(n29146), .Z(n29230) );
  XOR U28941 ( .A(n29237), .B(n29238), .Z(n29146) );
  AND U28942 ( .A(n750), .B(n29239), .Z(n29237) );
  XOR U28943 ( .A(n29240), .B(n29238), .Z(n29239) );
  XNOR U28944 ( .A(n29241), .B(n29242), .Z(n29229) );
  AND U28945 ( .A(n29243), .B(n29244), .Z(n29241) );
  XNOR U28946 ( .A(n29242), .B(n29171), .Z(n29244) );
  XOR U28947 ( .A(n29235), .B(n29236), .Z(n29171) );
  XNOR U28948 ( .A(n29245), .B(n29246), .Z(n29236) );
  ANDN U28949 ( .B(n29247), .A(n29248), .Z(n29245) );
  XOR U28950 ( .A(n29249), .B(n29250), .Z(n29247) );
  XOR U28951 ( .A(n29251), .B(n29252), .Z(n29235) );
  XNOR U28952 ( .A(n29253), .B(n29254), .Z(n29252) );
  ANDN U28953 ( .B(n29255), .A(n29256), .Z(n29253) );
  XNOR U28954 ( .A(n29257), .B(n29258), .Z(n29255) );
  IV U28955 ( .A(n29233), .Z(n29251) );
  XOR U28956 ( .A(n29259), .B(n29260), .Z(n29233) );
  ANDN U28957 ( .B(n29261), .A(n29262), .Z(n29259) );
  XOR U28958 ( .A(n29260), .B(n29263), .Z(n29261) );
  XOR U28959 ( .A(n29242), .B(n29173), .Z(n29243) );
  XOR U28960 ( .A(n29264), .B(n29265), .Z(n29173) );
  AND U28961 ( .A(n750), .B(n29266), .Z(n29264) );
  XOR U28962 ( .A(n29267), .B(n29265), .Z(n29266) );
  XNOR U28963 ( .A(n29268), .B(n29269), .Z(n29242) );
  NAND U28964 ( .A(n29270), .B(n29271), .Z(n29269) );
  XOR U28965 ( .A(n29272), .B(n29221), .Z(n29271) );
  XOR U28966 ( .A(n29262), .B(n29263), .Z(n29221) );
  XOR U28967 ( .A(n29273), .B(n29250), .Z(n29263) );
  XOR U28968 ( .A(n29274), .B(n29275), .Z(n29250) );
  ANDN U28969 ( .B(n29276), .A(n29277), .Z(n29274) );
  XOR U28970 ( .A(n29275), .B(n29278), .Z(n29276) );
  IV U28971 ( .A(n29248), .Z(n29273) );
  XOR U28972 ( .A(n29246), .B(n29279), .Z(n29248) );
  XOR U28973 ( .A(n29280), .B(n29281), .Z(n29279) );
  ANDN U28974 ( .B(n29282), .A(n29283), .Z(n29280) );
  XOR U28975 ( .A(n29284), .B(n29281), .Z(n29282) );
  IV U28976 ( .A(n29249), .Z(n29246) );
  XOR U28977 ( .A(n29285), .B(n29286), .Z(n29249) );
  ANDN U28978 ( .B(n29287), .A(n29288), .Z(n29285) );
  XOR U28979 ( .A(n29286), .B(n29289), .Z(n29287) );
  XOR U28980 ( .A(n29290), .B(n29291), .Z(n29262) );
  XNOR U28981 ( .A(n29257), .B(n29292), .Z(n29291) );
  IV U28982 ( .A(n29260), .Z(n29292) );
  XOR U28983 ( .A(n29293), .B(n29294), .Z(n29260) );
  ANDN U28984 ( .B(n29295), .A(n29296), .Z(n29293) );
  XOR U28985 ( .A(n29294), .B(n29297), .Z(n29295) );
  XNOR U28986 ( .A(n29298), .B(n29299), .Z(n29257) );
  ANDN U28987 ( .B(n29300), .A(n29301), .Z(n29298) );
  XOR U28988 ( .A(n29299), .B(n29302), .Z(n29300) );
  IV U28989 ( .A(n29256), .Z(n29290) );
  XOR U28990 ( .A(n29254), .B(n29303), .Z(n29256) );
  XOR U28991 ( .A(n29304), .B(n29305), .Z(n29303) );
  ANDN U28992 ( .B(n29306), .A(n29307), .Z(n29304) );
  XOR U28993 ( .A(n29308), .B(n29305), .Z(n29306) );
  IV U28994 ( .A(n29258), .Z(n29254) );
  XOR U28995 ( .A(n29309), .B(n29310), .Z(n29258) );
  ANDN U28996 ( .B(n29311), .A(n29312), .Z(n29309) );
  XOR U28997 ( .A(n29313), .B(n29310), .Z(n29311) );
  IV U28998 ( .A(n29268), .Z(n29272) );
  XOR U28999 ( .A(n29268), .B(n29223), .Z(n29270) );
  XOR U29000 ( .A(n29314), .B(n29315), .Z(n29223) );
  AND U29001 ( .A(n750), .B(n29316), .Z(n29314) );
  XOR U29002 ( .A(n29317), .B(n29315), .Z(n29316) );
  NANDN U29003 ( .A(n29225), .B(n29227), .Z(n29268) );
  XOR U29004 ( .A(n29318), .B(n29319), .Z(n29227) );
  AND U29005 ( .A(n750), .B(n29320), .Z(n29318) );
  XOR U29006 ( .A(n29319), .B(n29321), .Z(n29320) );
  XNOR U29007 ( .A(n29322), .B(n29323), .Z(n750) );
  AND U29008 ( .A(n29324), .B(n29325), .Z(n29322) );
  XOR U29009 ( .A(n29323), .B(n29238), .Z(n29325) );
  XNOR U29010 ( .A(n29326), .B(n29327), .Z(n29238) );
  ANDN U29011 ( .B(n29328), .A(n29329), .Z(n29326) );
  XOR U29012 ( .A(n29327), .B(n29330), .Z(n29328) );
  XNOR U29013 ( .A(n29323), .B(n29240), .Z(n29324) );
  XOR U29014 ( .A(n29331), .B(n29332), .Z(n29240) );
  AND U29015 ( .A(n754), .B(n29333), .Z(n29331) );
  XOR U29016 ( .A(n29334), .B(n29332), .Z(n29333) );
  XNOR U29017 ( .A(n29335), .B(n29336), .Z(n29323) );
  AND U29018 ( .A(n29337), .B(n29338), .Z(n29335) );
  XNOR U29019 ( .A(n29336), .B(n29265), .Z(n29338) );
  XOR U29020 ( .A(n29329), .B(n29330), .Z(n29265) );
  XNOR U29021 ( .A(n29339), .B(n29340), .Z(n29330) );
  ANDN U29022 ( .B(n29341), .A(n29342), .Z(n29339) );
  XOR U29023 ( .A(n29343), .B(n29344), .Z(n29341) );
  XOR U29024 ( .A(n29345), .B(n29346), .Z(n29329) );
  XNOR U29025 ( .A(n29347), .B(n29348), .Z(n29346) );
  ANDN U29026 ( .B(n29349), .A(n29350), .Z(n29347) );
  XNOR U29027 ( .A(n29351), .B(n29352), .Z(n29349) );
  IV U29028 ( .A(n29327), .Z(n29345) );
  XOR U29029 ( .A(n29353), .B(n29354), .Z(n29327) );
  ANDN U29030 ( .B(n29355), .A(n29356), .Z(n29353) );
  XOR U29031 ( .A(n29354), .B(n29357), .Z(n29355) );
  XOR U29032 ( .A(n29336), .B(n29267), .Z(n29337) );
  XOR U29033 ( .A(n29358), .B(n29359), .Z(n29267) );
  AND U29034 ( .A(n754), .B(n29360), .Z(n29358) );
  XOR U29035 ( .A(n29361), .B(n29359), .Z(n29360) );
  XNOR U29036 ( .A(n29362), .B(n29363), .Z(n29336) );
  NAND U29037 ( .A(n29364), .B(n29365), .Z(n29363) );
  XOR U29038 ( .A(n29366), .B(n29315), .Z(n29365) );
  XOR U29039 ( .A(n29356), .B(n29357), .Z(n29315) );
  XOR U29040 ( .A(n29367), .B(n29344), .Z(n29357) );
  XOR U29041 ( .A(n29368), .B(n29369), .Z(n29344) );
  ANDN U29042 ( .B(n29370), .A(n29371), .Z(n29368) );
  XOR U29043 ( .A(n29369), .B(n29372), .Z(n29370) );
  IV U29044 ( .A(n29342), .Z(n29367) );
  XOR U29045 ( .A(n29340), .B(n29373), .Z(n29342) );
  XOR U29046 ( .A(n29374), .B(n29375), .Z(n29373) );
  ANDN U29047 ( .B(n29376), .A(n29377), .Z(n29374) );
  XOR U29048 ( .A(n29378), .B(n29375), .Z(n29376) );
  IV U29049 ( .A(n29343), .Z(n29340) );
  XOR U29050 ( .A(n29379), .B(n29380), .Z(n29343) );
  ANDN U29051 ( .B(n29381), .A(n29382), .Z(n29379) );
  XOR U29052 ( .A(n29380), .B(n29383), .Z(n29381) );
  XOR U29053 ( .A(n29384), .B(n29385), .Z(n29356) );
  XNOR U29054 ( .A(n29351), .B(n29386), .Z(n29385) );
  IV U29055 ( .A(n29354), .Z(n29386) );
  XOR U29056 ( .A(n29387), .B(n29388), .Z(n29354) );
  ANDN U29057 ( .B(n29389), .A(n29390), .Z(n29387) );
  XOR U29058 ( .A(n29388), .B(n29391), .Z(n29389) );
  XNOR U29059 ( .A(n29392), .B(n29393), .Z(n29351) );
  ANDN U29060 ( .B(n29394), .A(n29395), .Z(n29392) );
  XOR U29061 ( .A(n29393), .B(n29396), .Z(n29394) );
  IV U29062 ( .A(n29350), .Z(n29384) );
  XOR U29063 ( .A(n29348), .B(n29397), .Z(n29350) );
  XOR U29064 ( .A(n29398), .B(n29399), .Z(n29397) );
  ANDN U29065 ( .B(n29400), .A(n29401), .Z(n29398) );
  XOR U29066 ( .A(n29402), .B(n29399), .Z(n29400) );
  IV U29067 ( .A(n29352), .Z(n29348) );
  XOR U29068 ( .A(n29403), .B(n29404), .Z(n29352) );
  ANDN U29069 ( .B(n29405), .A(n29406), .Z(n29403) );
  XOR U29070 ( .A(n29407), .B(n29404), .Z(n29405) );
  IV U29071 ( .A(n29362), .Z(n29366) );
  XOR U29072 ( .A(n29362), .B(n29317), .Z(n29364) );
  XOR U29073 ( .A(n29408), .B(n29409), .Z(n29317) );
  AND U29074 ( .A(n754), .B(n29410), .Z(n29408) );
  XOR U29075 ( .A(n29411), .B(n29409), .Z(n29410) );
  NANDN U29076 ( .A(n29319), .B(n29321), .Z(n29362) );
  XOR U29077 ( .A(n29412), .B(n29413), .Z(n29321) );
  AND U29078 ( .A(n754), .B(n29414), .Z(n29412) );
  XOR U29079 ( .A(n29413), .B(n29415), .Z(n29414) );
  XNOR U29080 ( .A(n29416), .B(n29417), .Z(n754) );
  AND U29081 ( .A(n29418), .B(n29419), .Z(n29416) );
  XOR U29082 ( .A(n29417), .B(n29332), .Z(n29419) );
  XNOR U29083 ( .A(n29420), .B(n29421), .Z(n29332) );
  ANDN U29084 ( .B(n29422), .A(n29423), .Z(n29420) );
  XOR U29085 ( .A(n29421), .B(n29424), .Z(n29422) );
  XNOR U29086 ( .A(n29417), .B(n29334), .Z(n29418) );
  XOR U29087 ( .A(n29425), .B(n29426), .Z(n29334) );
  AND U29088 ( .A(n758), .B(n29427), .Z(n29425) );
  XOR U29089 ( .A(n29428), .B(n29426), .Z(n29427) );
  XNOR U29090 ( .A(n29429), .B(n29430), .Z(n29417) );
  AND U29091 ( .A(n29431), .B(n29432), .Z(n29429) );
  XNOR U29092 ( .A(n29430), .B(n29359), .Z(n29432) );
  XOR U29093 ( .A(n29423), .B(n29424), .Z(n29359) );
  XNOR U29094 ( .A(n29433), .B(n29434), .Z(n29424) );
  ANDN U29095 ( .B(n29435), .A(n29436), .Z(n29433) );
  XOR U29096 ( .A(n29437), .B(n29438), .Z(n29435) );
  XOR U29097 ( .A(n29439), .B(n29440), .Z(n29423) );
  XNOR U29098 ( .A(n29441), .B(n29442), .Z(n29440) );
  ANDN U29099 ( .B(n29443), .A(n29444), .Z(n29441) );
  XNOR U29100 ( .A(n29445), .B(n29446), .Z(n29443) );
  IV U29101 ( .A(n29421), .Z(n29439) );
  XOR U29102 ( .A(n29447), .B(n29448), .Z(n29421) );
  ANDN U29103 ( .B(n29449), .A(n29450), .Z(n29447) );
  XOR U29104 ( .A(n29448), .B(n29451), .Z(n29449) );
  XOR U29105 ( .A(n29430), .B(n29361), .Z(n29431) );
  XOR U29106 ( .A(n29452), .B(n29453), .Z(n29361) );
  AND U29107 ( .A(n758), .B(n29454), .Z(n29452) );
  XOR U29108 ( .A(n29455), .B(n29453), .Z(n29454) );
  XNOR U29109 ( .A(n29456), .B(n29457), .Z(n29430) );
  NAND U29110 ( .A(n29458), .B(n29459), .Z(n29457) );
  XOR U29111 ( .A(n29460), .B(n29409), .Z(n29459) );
  XOR U29112 ( .A(n29450), .B(n29451), .Z(n29409) );
  XOR U29113 ( .A(n29461), .B(n29438), .Z(n29451) );
  XOR U29114 ( .A(n29462), .B(n29463), .Z(n29438) );
  ANDN U29115 ( .B(n29464), .A(n29465), .Z(n29462) );
  XOR U29116 ( .A(n29463), .B(n29466), .Z(n29464) );
  IV U29117 ( .A(n29436), .Z(n29461) );
  XOR U29118 ( .A(n29434), .B(n29467), .Z(n29436) );
  XOR U29119 ( .A(n29468), .B(n29469), .Z(n29467) );
  ANDN U29120 ( .B(n29470), .A(n29471), .Z(n29468) );
  XOR U29121 ( .A(n29472), .B(n29469), .Z(n29470) );
  IV U29122 ( .A(n29437), .Z(n29434) );
  XOR U29123 ( .A(n29473), .B(n29474), .Z(n29437) );
  ANDN U29124 ( .B(n29475), .A(n29476), .Z(n29473) );
  XOR U29125 ( .A(n29474), .B(n29477), .Z(n29475) );
  XOR U29126 ( .A(n29478), .B(n29479), .Z(n29450) );
  XNOR U29127 ( .A(n29445), .B(n29480), .Z(n29479) );
  IV U29128 ( .A(n29448), .Z(n29480) );
  XOR U29129 ( .A(n29481), .B(n29482), .Z(n29448) );
  ANDN U29130 ( .B(n29483), .A(n29484), .Z(n29481) );
  XOR U29131 ( .A(n29482), .B(n29485), .Z(n29483) );
  XNOR U29132 ( .A(n29486), .B(n29487), .Z(n29445) );
  ANDN U29133 ( .B(n29488), .A(n29489), .Z(n29486) );
  XOR U29134 ( .A(n29487), .B(n29490), .Z(n29488) );
  IV U29135 ( .A(n29444), .Z(n29478) );
  XOR U29136 ( .A(n29442), .B(n29491), .Z(n29444) );
  XOR U29137 ( .A(n29492), .B(n29493), .Z(n29491) );
  ANDN U29138 ( .B(n29494), .A(n29495), .Z(n29492) );
  XOR U29139 ( .A(n29496), .B(n29493), .Z(n29494) );
  IV U29140 ( .A(n29446), .Z(n29442) );
  XOR U29141 ( .A(n29497), .B(n29498), .Z(n29446) );
  ANDN U29142 ( .B(n29499), .A(n29500), .Z(n29497) );
  XOR U29143 ( .A(n29501), .B(n29498), .Z(n29499) );
  IV U29144 ( .A(n29456), .Z(n29460) );
  XOR U29145 ( .A(n29456), .B(n29411), .Z(n29458) );
  XOR U29146 ( .A(n29502), .B(n29503), .Z(n29411) );
  AND U29147 ( .A(n758), .B(n29504), .Z(n29502) );
  XOR U29148 ( .A(n29505), .B(n29503), .Z(n29504) );
  NANDN U29149 ( .A(n29413), .B(n29415), .Z(n29456) );
  XOR U29150 ( .A(n29506), .B(n29507), .Z(n29415) );
  AND U29151 ( .A(n758), .B(n29508), .Z(n29506) );
  XOR U29152 ( .A(n29507), .B(n29509), .Z(n29508) );
  XNOR U29153 ( .A(n29510), .B(n29511), .Z(n758) );
  AND U29154 ( .A(n29512), .B(n29513), .Z(n29510) );
  XOR U29155 ( .A(n29511), .B(n29426), .Z(n29513) );
  XNOR U29156 ( .A(n29514), .B(n29515), .Z(n29426) );
  ANDN U29157 ( .B(n29516), .A(n29517), .Z(n29514) );
  XOR U29158 ( .A(n29515), .B(n29518), .Z(n29516) );
  XNOR U29159 ( .A(n29511), .B(n29428), .Z(n29512) );
  XOR U29160 ( .A(n29519), .B(n29520), .Z(n29428) );
  AND U29161 ( .A(n762), .B(n29521), .Z(n29519) );
  XOR U29162 ( .A(n29522), .B(n29520), .Z(n29521) );
  XNOR U29163 ( .A(n29523), .B(n29524), .Z(n29511) );
  AND U29164 ( .A(n29525), .B(n29526), .Z(n29523) );
  XNOR U29165 ( .A(n29524), .B(n29453), .Z(n29526) );
  XOR U29166 ( .A(n29517), .B(n29518), .Z(n29453) );
  XNOR U29167 ( .A(n29527), .B(n29528), .Z(n29518) );
  ANDN U29168 ( .B(n29529), .A(n29530), .Z(n29527) );
  XOR U29169 ( .A(n29531), .B(n29532), .Z(n29529) );
  XOR U29170 ( .A(n29533), .B(n29534), .Z(n29517) );
  XNOR U29171 ( .A(n29535), .B(n29536), .Z(n29534) );
  ANDN U29172 ( .B(n29537), .A(n29538), .Z(n29535) );
  XNOR U29173 ( .A(n29539), .B(n29540), .Z(n29537) );
  IV U29174 ( .A(n29515), .Z(n29533) );
  XOR U29175 ( .A(n29541), .B(n29542), .Z(n29515) );
  ANDN U29176 ( .B(n29543), .A(n29544), .Z(n29541) );
  XOR U29177 ( .A(n29542), .B(n29545), .Z(n29543) );
  XOR U29178 ( .A(n29524), .B(n29455), .Z(n29525) );
  XOR U29179 ( .A(n29546), .B(n29547), .Z(n29455) );
  AND U29180 ( .A(n762), .B(n29548), .Z(n29546) );
  XOR U29181 ( .A(n29549), .B(n29547), .Z(n29548) );
  XNOR U29182 ( .A(n29550), .B(n29551), .Z(n29524) );
  NAND U29183 ( .A(n29552), .B(n29553), .Z(n29551) );
  XOR U29184 ( .A(n29554), .B(n29503), .Z(n29553) );
  XOR U29185 ( .A(n29544), .B(n29545), .Z(n29503) );
  XOR U29186 ( .A(n29555), .B(n29532), .Z(n29545) );
  XOR U29187 ( .A(n29556), .B(n29557), .Z(n29532) );
  ANDN U29188 ( .B(n29558), .A(n29559), .Z(n29556) );
  XOR U29189 ( .A(n29557), .B(n29560), .Z(n29558) );
  IV U29190 ( .A(n29530), .Z(n29555) );
  XOR U29191 ( .A(n29528), .B(n29561), .Z(n29530) );
  XOR U29192 ( .A(n29562), .B(n29563), .Z(n29561) );
  ANDN U29193 ( .B(n29564), .A(n29565), .Z(n29562) );
  XOR U29194 ( .A(n29566), .B(n29563), .Z(n29564) );
  IV U29195 ( .A(n29531), .Z(n29528) );
  XOR U29196 ( .A(n29567), .B(n29568), .Z(n29531) );
  ANDN U29197 ( .B(n29569), .A(n29570), .Z(n29567) );
  XOR U29198 ( .A(n29568), .B(n29571), .Z(n29569) );
  XOR U29199 ( .A(n29572), .B(n29573), .Z(n29544) );
  XNOR U29200 ( .A(n29539), .B(n29574), .Z(n29573) );
  IV U29201 ( .A(n29542), .Z(n29574) );
  XOR U29202 ( .A(n29575), .B(n29576), .Z(n29542) );
  ANDN U29203 ( .B(n29577), .A(n29578), .Z(n29575) );
  XOR U29204 ( .A(n29576), .B(n29579), .Z(n29577) );
  XNOR U29205 ( .A(n29580), .B(n29581), .Z(n29539) );
  ANDN U29206 ( .B(n29582), .A(n29583), .Z(n29580) );
  XOR U29207 ( .A(n29581), .B(n29584), .Z(n29582) );
  IV U29208 ( .A(n29538), .Z(n29572) );
  XOR U29209 ( .A(n29536), .B(n29585), .Z(n29538) );
  XOR U29210 ( .A(n29586), .B(n29587), .Z(n29585) );
  ANDN U29211 ( .B(n29588), .A(n29589), .Z(n29586) );
  XOR U29212 ( .A(n29590), .B(n29587), .Z(n29588) );
  IV U29213 ( .A(n29540), .Z(n29536) );
  XOR U29214 ( .A(n29591), .B(n29592), .Z(n29540) );
  ANDN U29215 ( .B(n29593), .A(n29594), .Z(n29591) );
  XOR U29216 ( .A(n29595), .B(n29592), .Z(n29593) );
  IV U29217 ( .A(n29550), .Z(n29554) );
  XOR U29218 ( .A(n29550), .B(n29505), .Z(n29552) );
  XOR U29219 ( .A(n29596), .B(n29597), .Z(n29505) );
  AND U29220 ( .A(n762), .B(n29598), .Z(n29596) );
  XOR U29221 ( .A(n29599), .B(n29597), .Z(n29598) );
  NANDN U29222 ( .A(n29507), .B(n29509), .Z(n29550) );
  XOR U29223 ( .A(n29600), .B(n29601), .Z(n29509) );
  AND U29224 ( .A(n762), .B(n29602), .Z(n29600) );
  XOR U29225 ( .A(n29601), .B(n29603), .Z(n29602) );
  XNOR U29226 ( .A(n29604), .B(n29605), .Z(n762) );
  AND U29227 ( .A(n29606), .B(n29607), .Z(n29604) );
  XOR U29228 ( .A(n29605), .B(n29520), .Z(n29607) );
  XNOR U29229 ( .A(n29608), .B(n29609), .Z(n29520) );
  ANDN U29230 ( .B(n29610), .A(n29611), .Z(n29608) );
  XOR U29231 ( .A(n29609), .B(n29612), .Z(n29610) );
  XNOR U29232 ( .A(n29605), .B(n29522), .Z(n29606) );
  XOR U29233 ( .A(n29613), .B(n29614), .Z(n29522) );
  AND U29234 ( .A(n766), .B(n29615), .Z(n29613) );
  XOR U29235 ( .A(n29616), .B(n29614), .Z(n29615) );
  XNOR U29236 ( .A(n29617), .B(n29618), .Z(n29605) );
  AND U29237 ( .A(n29619), .B(n29620), .Z(n29617) );
  XNOR U29238 ( .A(n29618), .B(n29547), .Z(n29620) );
  XOR U29239 ( .A(n29611), .B(n29612), .Z(n29547) );
  XNOR U29240 ( .A(n29621), .B(n29622), .Z(n29612) );
  ANDN U29241 ( .B(n29623), .A(n29624), .Z(n29621) );
  XOR U29242 ( .A(n29625), .B(n29626), .Z(n29623) );
  XOR U29243 ( .A(n29627), .B(n29628), .Z(n29611) );
  XNOR U29244 ( .A(n29629), .B(n29630), .Z(n29628) );
  ANDN U29245 ( .B(n29631), .A(n29632), .Z(n29629) );
  XNOR U29246 ( .A(n29633), .B(n29634), .Z(n29631) );
  IV U29247 ( .A(n29609), .Z(n29627) );
  XOR U29248 ( .A(n29635), .B(n29636), .Z(n29609) );
  ANDN U29249 ( .B(n29637), .A(n29638), .Z(n29635) );
  XOR U29250 ( .A(n29636), .B(n29639), .Z(n29637) );
  XOR U29251 ( .A(n29618), .B(n29549), .Z(n29619) );
  XOR U29252 ( .A(n29640), .B(n29641), .Z(n29549) );
  AND U29253 ( .A(n766), .B(n29642), .Z(n29640) );
  XOR U29254 ( .A(n29643), .B(n29641), .Z(n29642) );
  XNOR U29255 ( .A(n29644), .B(n29645), .Z(n29618) );
  NAND U29256 ( .A(n29646), .B(n29647), .Z(n29645) );
  XOR U29257 ( .A(n29648), .B(n29597), .Z(n29647) );
  XOR U29258 ( .A(n29638), .B(n29639), .Z(n29597) );
  XOR U29259 ( .A(n29649), .B(n29626), .Z(n29639) );
  XOR U29260 ( .A(n29650), .B(n29651), .Z(n29626) );
  ANDN U29261 ( .B(n29652), .A(n29653), .Z(n29650) );
  XOR U29262 ( .A(n29651), .B(n29654), .Z(n29652) );
  IV U29263 ( .A(n29624), .Z(n29649) );
  XOR U29264 ( .A(n29622), .B(n29655), .Z(n29624) );
  XOR U29265 ( .A(n29656), .B(n29657), .Z(n29655) );
  ANDN U29266 ( .B(n29658), .A(n29659), .Z(n29656) );
  XOR U29267 ( .A(n29660), .B(n29657), .Z(n29658) );
  IV U29268 ( .A(n29625), .Z(n29622) );
  XOR U29269 ( .A(n29661), .B(n29662), .Z(n29625) );
  ANDN U29270 ( .B(n29663), .A(n29664), .Z(n29661) );
  XOR U29271 ( .A(n29662), .B(n29665), .Z(n29663) );
  XOR U29272 ( .A(n29666), .B(n29667), .Z(n29638) );
  XNOR U29273 ( .A(n29633), .B(n29668), .Z(n29667) );
  IV U29274 ( .A(n29636), .Z(n29668) );
  XOR U29275 ( .A(n29669), .B(n29670), .Z(n29636) );
  ANDN U29276 ( .B(n29671), .A(n29672), .Z(n29669) );
  XOR U29277 ( .A(n29670), .B(n29673), .Z(n29671) );
  XNOR U29278 ( .A(n29674), .B(n29675), .Z(n29633) );
  ANDN U29279 ( .B(n29676), .A(n29677), .Z(n29674) );
  XOR U29280 ( .A(n29675), .B(n29678), .Z(n29676) );
  IV U29281 ( .A(n29632), .Z(n29666) );
  XOR U29282 ( .A(n29630), .B(n29679), .Z(n29632) );
  XOR U29283 ( .A(n29680), .B(n29681), .Z(n29679) );
  ANDN U29284 ( .B(n29682), .A(n29683), .Z(n29680) );
  XOR U29285 ( .A(n29684), .B(n29681), .Z(n29682) );
  IV U29286 ( .A(n29634), .Z(n29630) );
  XOR U29287 ( .A(n29685), .B(n29686), .Z(n29634) );
  ANDN U29288 ( .B(n29687), .A(n29688), .Z(n29685) );
  XOR U29289 ( .A(n29689), .B(n29686), .Z(n29687) );
  IV U29290 ( .A(n29644), .Z(n29648) );
  XOR U29291 ( .A(n29644), .B(n29599), .Z(n29646) );
  XOR U29292 ( .A(n29690), .B(n29691), .Z(n29599) );
  AND U29293 ( .A(n766), .B(n29692), .Z(n29690) );
  XOR U29294 ( .A(n29693), .B(n29691), .Z(n29692) );
  NANDN U29295 ( .A(n29601), .B(n29603), .Z(n29644) );
  XOR U29296 ( .A(n29694), .B(n29695), .Z(n29603) );
  AND U29297 ( .A(n766), .B(n29696), .Z(n29694) );
  XOR U29298 ( .A(n29695), .B(n29697), .Z(n29696) );
  XNOR U29299 ( .A(n29698), .B(n29699), .Z(n766) );
  AND U29300 ( .A(n29700), .B(n29701), .Z(n29698) );
  XOR U29301 ( .A(n29699), .B(n29614), .Z(n29701) );
  XNOR U29302 ( .A(n29702), .B(n29703), .Z(n29614) );
  ANDN U29303 ( .B(n29704), .A(n29705), .Z(n29702) );
  XOR U29304 ( .A(n29703), .B(n29706), .Z(n29704) );
  XNOR U29305 ( .A(n29699), .B(n29616), .Z(n29700) );
  XOR U29306 ( .A(n29707), .B(n29708), .Z(n29616) );
  AND U29307 ( .A(n770), .B(n29709), .Z(n29707) );
  XOR U29308 ( .A(n29710), .B(n29708), .Z(n29709) );
  XNOR U29309 ( .A(n29711), .B(n29712), .Z(n29699) );
  AND U29310 ( .A(n29713), .B(n29714), .Z(n29711) );
  XNOR U29311 ( .A(n29712), .B(n29641), .Z(n29714) );
  XOR U29312 ( .A(n29705), .B(n29706), .Z(n29641) );
  XNOR U29313 ( .A(n29715), .B(n29716), .Z(n29706) );
  ANDN U29314 ( .B(n29717), .A(n29718), .Z(n29715) );
  XOR U29315 ( .A(n29719), .B(n29720), .Z(n29717) );
  XOR U29316 ( .A(n29721), .B(n29722), .Z(n29705) );
  XNOR U29317 ( .A(n29723), .B(n29724), .Z(n29722) );
  ANDN U29318 ( .B(n29725), .A(n29726), .Z(n29723) );
  XNOR U29319 ( .A(n29727), .B(n29728), .Z(n29725) );
  IV U29320 ( .A(n29703), .Z(n29721) );
  XOR U29321 ( .A(n29729), .B(n29730), .Z(n29703) );
  ANDN U29322 ( .B(n29731), .A(n29732), .Z(n29729) );
  XOR U29323 ( .A(n29730), .B(n29733), .Z(n29731) );
  XOR U29324 ( .A(n29712), .B(n29643), .Z(n29713) );
  XOR U29325 ( .A(n29734), .B(n29735), .Z(n29643) );
  AND U29326 ( .A(n770), .B(n29736), .Z(n29734) );
  XOR U29327 ( .A(n29737), .B(n29735), .Z(n29736) );
  XNOR U29328 ( .A(n29738), .B(n29739), .Z(n29712) );
  NAND U29329 ( .A(n29740), .B(n29741), .Z(n29739) );
  XOR U29330 ( .A(n29742), .B(n29691), .Z(n29741) );
  XOR U29331 ( .A(n29732), .B(n29733), .Z(n29691) );
  XOR U29332 ( .A(n29743), .B(n29720), .Z(n29733) );
  XOR U29333 ( .A(n29744), .B(n29745), .Z(n29720) );
  ANDN U29334 ( .B(n29746), .A(n29747), .Z(n29744) );
  XOR U29335 ( .A(n29745), .B(n29748), .Z(n29746) );
  IV U29336 ( .A(n29718), .Z(n29743) );
  XOR U29337 ( .A(n29716), .B(n29749), .Z(n29718) );
  XOR U29338 ( .A(n29750), .B(n29751), .Z(n29749) );
  ANDN U29339 ( .B(n29752), .A(n29753), .Z(n29750) );
  XOR U29340 ( .A(n29754), .B(n29751), .Z(n29752) );
  IV U29341 ( .A(n29719), .Z(n29716) );
  XOR U29342 ( .A(n29755), .B(n29756), .Z(n29719) );
  ANDN U29343 ( .B(n29757), .A(n29758), .Z(n29755) );
  XOR U29344 ( .A(n29756), .B(n29759), .Z(n29757) );
  XOR U29345 ( .A(n29760), .B(n29761), .Z(n29732) );
  XNOR U29346 ( .A(n29727), .B(n29762), .Z(n29761) );
  IV U29347 ( .A(n29730), .Z(n29762) );
  XOR U29348 ( .A(n29763), .B(n29764), .Z(n29730) );
  ANDN U29349 ( .B(n29765), .A(n29766), .Z(n29763) );
  XOR U29350 ( .A(n29764), .B(n29767), .Z(n29765) );
  XNOR U29351 ( .A(n29768), .B(n29769), .Z(n29727) );
  ANDN U29352 ( .B(n29770), .A(n29771), .Z(n29768) );
  XOR U29353 ( .A(n29769), .B(n29772), .Z(n29770) );
  IV U29354 ( .A(n29726), .Z(n29760) );
  XOR U29355 ( .A(n29724), .B(n29773), .Z(n29726) );
  XOR U29356 ( .A(n29774), .B(n29775), .Z(n29773) );
  ANDN U29357 ( .B(n29776), .A(n29777), .Z(n29774) );
  XOR U29358 ( .A(n29778), .B(n29775), .Z(n29776) );
  IV U29359 ( .A(n29728), .Z(n29724) );
  XOR U29360 ( .A(n29779), .B(n29780), .Z(n29728) );
  ANDN U29361 ( .B(n29781), .A(n29782), .Z(n29779) );
  XOR U29362 ( .A(n29783), .B(n29780), .Z(n29781) );
  IV U29363 ( .A(n29738), .Z(n29742) );
  XOR U29364 ( .A(n29738), .B(n29693), .Z(n29740) );
  XOR U29365 ( .A(n29784), .B(n29785), .Z(n29693) );
  AND U29366 ( .A(n770), .B(n29786), .Z(n29784) );
  XOR U29367 ( .A(n29787), .B(n29785), .Z(n29786) );
  NANDN U29368 ( .A(n29695), .B(n29697), .Z(n29738) );
  XOR U29369 ( .A(n29788), .B(n29789), .Z(n29697) );
  AND U29370 ( .A(n770), .B(n29790), .Z(n29788) );
  XOR U29371 ( .A(n29789), .B(n29791), .Z(n29790) );
  XNOR U29372 ( .A(n29792), .B(n29793), .Z(n770) );
  AND U29373 ( .A(n29794), .B(n29795), .Z(n29792) );
  XOR U29374 ( .A(n29793), .B(n29708), .Z(n29795) );
  XNOR U29375 ( .A(n29796), .B(n29797), .Z(n29708) );
  ANDN U29376 ( .B(n29798), .A(n29799), .Z(n29796) );
  XOR U29377 ( .A(n29797), .B(n29800), .Z(n29798) );
  XNOR U29378 ( .A(n29793), .B(n29710), .Z(n29794) );
  XOR U29379 ( .A(n29801), .B(n29802), .Z(n29710) );
  AND U29380 ( .A(n774), .B(n29803), .Z(n29801) );
  XOR U29381 ( .A(n29804), .B(n29802), .Z(n29803) );
  XNOR U29382 ( .A(n29805), .B(n29806), .Z(n29793) );
  AND U29383 ( .A(n29807), .B(n29808), .Z(n29805) );
  XNOR U29384 ( .A(n29806), .B(n29735), .Z(n29808) );
  XOR U29385 ( .A(n29799), .B(n29800), .Z(n29735) );
  XNOR U29386 ( .A(n29809), .B(n29810), .Z(n29800) );
  ANDN U29387 ( .B(n29811), .A(n29812), .Z(n29809) );
  XOR U29388 ( .A(n29813), .B(n29814), .Z(n29811) );
  XOR U29389 ( .A(n29815), .B(n29816), .Z(n29799) );
  XNOR U29390 ( .A(n29817), .B(n29818), .Z(n29816) );
  ANDN U29391 ( .B(n29819), .A(n29820), .Z(n29817) );
  XNOR U29392 ( .A(n29821), .B(n29822), .Z(n29819) );
  IV U29393 ( .A(n29797), .Z(n29815) );
  XOR U29394 ( .A(n29823), .B(n29824), .Z(n29797) );
  ANDN U29395 ( .B(n29825), .A(n29826), .Z(n29823) );
  XOR U29396 ( .A(n29824), .B(n29827), .Z(n29825) );
  XOR U29397 ( .A(n29806), .B(n29737), .Z(n29807) );
  XOR U29398 ( .A(n29828), .B(n29829), .Z(n29737) );
  AND U29399 ( .A(n774), .B(n29830), .Z(n29828) );
  XOR U29400 ( .A(n29831), .B(n29829), .Z(n29830) );
  XNOR U29401 ( .A(n29832), .B(n29833), .Z(n29806) );
  NAND U29402 ( .A(n29834), .B(n29835), .Z(n29833) );
  XOR U29403 ( .A(n29836), .B(n29785), .Z(n29835) );
  XOR U29404 ( .A(n29826), .B(n29827), .Z(n29785) );
  XOR U29405 ( .A(n29837), .B(n29814), .Z(n29827) );
  XOR U29406 ( .A(n29838), .B(n29839), .Z(n29814) );
  ANDN U29407 ( .B(n29840), .A(n29841), .Z(n29838) );
  XOR U29408 ( .A(n29839), .B(n29842), .Z(n29840) );
  IV U29409 ( .A(n29812), .Z(n29837) );
  XOR U29410 ( .A(n29810), .B(n29843), .Z(n29812) );
  XOR U29411 ( .A(n29844), .B(n29845), .Z(n29843) );
  ANDN U29412 ( .B(n29846), .A(n29847), .Z(n29844) );
  XOR U29413 ( .A(n29848), .B(n29845), .Z(n29846) );
  IV U29414 ( .A(n29813), .Z(n29810) );
  XOR U29415 ( .A(n29849), .B(n29850), .Z(n29813) );
  ANDN U29416 ( .B(n29851), .A(n29852), .Z(n29849) );
  XOR U29417 ( .A(n29850), .B(n29853), .Z(n29851) );
  XOR U29418 ( .A(n29854), .B(n29855), .Z(n29826) );
  XNOR U29419 ( .A(n29821), .B(n29856), .Z(n29855) );
  IV U29420 ( .A(n29824), .Z(n29856) );
  XOR U29421 ( .A(n29857), .B(n29858), .Z(n29824) );
  ANDN U29422 ( .B(n29859), .A(n29860), .Z(n29857) );
  XOR U29423 ( .A(n29858), .B(n29861), .Z(n29859) );
  XNOR U29424 ( .A(n29862), .B(n29863), .Z(n29821) );
  ANDN U29425 ( .B(n29864), .A(n29865), .Z(n29862) );
  XOR U29426 ( .A(n29863), .B(n29866), .Z(n29864) );
  IV U29427 ( .A(n29820), .Z(n29854) );
  XOR U29428 ( .A(n29818), .B(n29867), .Z(n29820) );
  XOR U29429 ( .A(n29868), .B(n29869), .Z(n29867) );
  ANDN U29430 ( .B(n29870), .A(n29871), .Z(n29868) );
  XOR U29431 ( .A(n29872), .B(n29869), .Z(n29870) );
  IV U29432 ( .A(n29822), .Z(n29818) );
  XOR U29433 ( .A(n29873), .B(n29874), .Z(n29822) );
  ANDN U29434 ( .B(n29875), .A(n29876), .Z(n29873) );
  XOR U29435 ( .A(n29877), .B(n29874), .Z(n29875) );
  IV U29436 ( .A(n29832), .Z(n29836) );
  XOR U29437 ( .A(n29832), .B(n29787), .Z(n29834) );
  XOR U29438 ( .A(n29878), .B(n29879), .Z(n29787) );
  AND U29439 ( .A(n774), .B(n29880), .Z(n29878) );
  XOR U29440 ( .A(n29881), .B(n29879), .Z(n29880) );
  NANDN U29441 ( .A(n29789), .B(n29791), .Z(n29832) );
  XOR U29442 ( .A(n29882), .B(n29883), .Z(n29791) );
  AND U29443 ( .A(n774), .B(n29884), .Z(n29882) );
  XOR U29444 ( .A(n29883), .B(n29885), .Z(n29884) );
  XNOR U29445 ( .A(n29886), .B(n29887), .Z(n774) );
  AND U29446 ( .A(n29888), .B(n29889), .Z(n29886) );
  XOR U29447 ( .A(n29887), .B(n29802), .Z(n29889) );
  XNOR U29448 ( .A(n29890), .B(n29891), .Z(n29802) );
  ANDN U29449 ( .B(n29892), .A(n29893), .Z(n29890) );
  XOR U29450 ( .A(n29891), .B(n29894), .Z(n29892) );
  XNOR U29451 ( .A(n29887), .B(n29804), .Z(n29888) );
  XOR U29452 ( .A(n29895), .B(n29896), .Z(n29804) );
  AND U29453 ( .A(n778), .B(n29897), .Z(n29895) );
  XOR U29454 ( .A(n29898), .B(n29896), .Z(n29897) );
  XNOR U29455 ( .A(n29899), .B(n29900), .Z(n29887) );
  AND U29456 ( .A(n29901), .B(n29902), .Z(n29899) );
  XNOR U29457 ( .A(n29900), .B(n29829), .Z(n29902) );
  XOR U29458 ( .A(n29893), .B(n29894), .Z(n29829) );
  XNOR U29459 ( .A(n29903), .B(n29904), .Z(n29894) );
  ANDN U29460 ( .B(n29905), .A(n29906), .Z(n29903) );
  XOR U29461 ( .A(n29907), .B(n29908), .Z(n29905) );
  XOR U29462 ( .A(n29909), .B(n29910), .Z(n29893) );
  XNOR U29463 ( .A(n29911), .B(n29912), .Z(n29910) );
  ANDN U29464 ( .B(n29913), .A(n29914), .Z(n29911) );
  XNOR U29465 ( .A(n29915), .B(n29916), .Z(n29913) );
  IV U29466 ( .A(n29891), .Z(n29909) );
  XOR U29467 ( .A(n29917), .B(n29918), .Z(n29891) );
  ANDN U29468 ( .B(n29919), .A(n29920), .Z(n29917) );
  XOR U29469 ( .A(n29918), .B(n29921), .Z(n29919) );
  XOR U29470 ( .A(n29900), .B(n29831), .Z(n29901) );
  XOR U29471 ( .A(n29922), .B(n29923), .Z(n29831) );
  AND U29472 ( .A(n778), .B(n29924), .Z(n29922) );
  XOR U29473 ( .A(n29925), .B(n29923), .Z(n29924) );
  XNOR U29474 ( .A(n29926), .B(n29927), .Z(n29900) );
  NAND U29475 ( .A(n29928), .B(n29929), .Z(n29927) );
  XOR U29476 ( .A(n29930), .B(n29879), .Z(n29929) );
  XOR U29477 ( .A(n29920), .B(n29921), .Z(n29879) );
  XOR U29478 ( .A(n29931), .B(n29908), .Z(n29921) );
  XOR U29479 ( .A(n29932), .B(n29933), .Z(n29908) );
  ANDN U29480 ( .B(n29934), .A(n29935), .Z(n29932) );
  XOR U29481 ( .A(n29933), .B(n29936), .Z(n29934) );
  IV U29482 ( .A(n29906), .Z(n29931) );
  XOR U29483 ( .A(n29904), .B(n29937), .Z(n29906) );
  XOR U29484 ( .A(n29938), .B(n29939), .Z(n29937) );
  ANDN U29485 ( .B(n29940), .A(n29941), .Z(n29938) );
  XOR U29486 ( .A(n29942), .B(n29939), .Z(n29940) );
  IV U29487 ( .A(n29907), .Z(n29904) );
  XOR U29488 ( .A(n29943), .B(n29944), .Z(n29907) );
  ANDN U29489 ( .B(n29945), .A(n29946), .Z(n29943) );
  XOR U29490 ( .A(n29944), .B(n29947), .Z(n29945) );
  XOR U29491 ( .A(n29948), .B(n29949), .Z(n29920) );
  XNOR U29492 ( .A(n29915), .B(n29950), .Z(n29949) );
  IV U29493 ( .A(n29918), .Z(n29950) );
  XOR U29494 ( .A(n29951), .B(n29952), .Z(n29918) );
  ANDN U29495 ( .B(n29953), .A(n29954), .Z(n29951) );
  XOR U29496 ( .A(n29952), .B(n29955), .Z(n29953) );
  XNOR U29497 ( .A(n29956), .B(n29957), .Z(n29915) );
  ANDN U29498 ( .B(n29958), .A(n29959), .Z(n29956) );
  XOR U29499 ( .A(n29957), .B(n29960), .Z(n29958) );
  IV U29500 ( .A(n29914), .Z(n29948) );
  XOR U29501 ( .A(n29912), .B(n29961), .Z(n29914) );
  XOR U29502 ( .A(n29962), .B(n29963), .Z(n29961) );
  ANDN U29503 ( .B(n29964), .A(n29965), .Z(n29962) );
  XOR U29504 ( .A(n29966), .B(n29963), .Z(n29964) );
  IV U29505 ( .A(n29916), .Z(n29912) );
  XOR U29506 ( .A(n29967), .B(n29968), .Z(n29916) );
  ANDN U29507 ( .B(n29969), .A(n29970), .Z(n29967) );
  XOR U29508 ( .A(n29971), .B(n29968), .Z(n29969) );
  IV U29509 ( .A(n29926), .Z(n29930) );
  XOR U29510 ( .A(n29926), .B(n29881), .Z(n29928) );
  XOR U29511 ( .A(n29972), .B(n29973), .Z(n29881) );
  AND U29512 ( .A(n778), .B(n29974), .Z(n29972) );
  XOR U29513 ( .A(n29975), .B(n29973), .Z(n29974) );
  NANDN U29514 ( .A(n29883), .B(n29885), .Z(n29926) );
  XOR U29515 ( .A(n29976), .B(n29977), .Z(n29885) );
  AND U29516 ( .A(n778), .B(n29978), .Z(n29976) );
  XOR U29517 ( .A(n29977), .B(n29979), .Z(n29978) );
  XNOR U29518 ( .A(n29980), .B(n29981), .Z(n778) );
  AND U29519 ( .A(n29982), .B(n29983), .Z(n29980) );
  XOR U29520 ( .A(n29981), .B(n29896), .Z(n29983) );
  XNOR U29521 ( .A(n29984), .B(n29985), .Z(n29896) );
  ANDN U29522 ( .B(n29986), .A(n29987), .Z(n29984) );
  XOR U29523 ( .A(n29985), .B(n29988), .Z(n29986) );
  XNOR U29524 ( .A(n29981), .B(n29898), .Z(n29982) );
  XOR U29525 ( .A(n29989), .B(n29990), .Z(n29898) );
  AND U29526 ( .A(n782), .B(n29991), .Z(n29989) );
  XOR U29527 ( .A(n29992), .B(n29990), .Z(n29991) );
  XNOR U29528 ( .A(n29993), .B(n29994), .Z(n29981) );
  AND U29529 ( .A(n29995), .B(n29996), .Z(n29993) );
  XNOR U29530 ( .A(n29994), .B(n29923), .Z(n29996) );
  XOR U29531 ( .A(n29987), .B(n29988), .Z(n29923) );
  XNOR U29532 ( .A(n29997), .B(n29998), .Z(n29988) );
  ANDN U29533 ( .B(n29999), .A(n30000), .Z(n29997) );
  XOR U29534 ( .A(n30001), .B(n30002), .Z(n29999) );
  XOR U29535 ( .A(n30003), .B(n30004), .Z(n29987) );
  XNOR U29536 ( .A(n30005), .B(n30006), .Z(n30004) );
  ANDN U29537 ( .B(n30007), .A(n30008), .Z(n30005) );
  XNOR U29538 ( .A(n30009), .B(n30010), .Z(n30007) );
  IV U29539 ( .A(n29985), .Z(n30003) );
  XOR U29540 ( .A(n30011), .B(n30012), .Z(n29985) );
  ANDN U29541 ( .B(n30013), .A(n30014), .Z(n30011) );
  XOR U29542 ( .A(n30012), .B(n30015), .Z(n30013) );
  XOR U29543 ( .A(n29994), .B(n29925), .Z(n29995) );
  XOR U29544 ( .A(n30016), .B(n30017), .Z(n29925) );
  AND U29545 ( .A(n782), .B(n30018), .Z(n30016) );
  XOR U29546 ( .A(n30019), .B(n30017), .Z(n30018) );
  XNOR U29547 ( .A(n30020), .B(n30021), .Z(n29994) );
  NAND U29548 ( .A(n30022), .B(n30023), .Z(n30021) );
  XOR U29549 ( .A(n30024), .B(n29973), .Z(n30023) );
  XOR U29550 ( .A(n30014), .B(n30015), .Z(n29973) );
  XOR U29551 ( .A(n30025), .B(n30002), .Z(n30015) );
  XOR U29552 ( .A(n30026), .B(n30027), .Z(n30002) );
  ANDN U29553 ( .B(n30028), .A(n30029), .Z(n30026) );
  XOR U29554 ( .A(n30027), .B(n30030), .Z(n30028) );
  IV U29555 ( .A(n30000), .Z(n30025) );
  XOR U29556 ( .A(n29998), .B(n30031), .Z(n30000) );
  XOR U29557 ( .A(n30032), .B(n30033), .Z(n30031) );
  ANDN U29558 ( .B(n30034), .A(n30035), .Z(n30032) );
  XOR U29559 ( .A(n30036), .B(n30033), .Z(n30034) );
  IV U29560 ( .A(n30001), .Z(n29998) );
  XOR U29561 ( .A(n30037), .B(n30038), .Z(n30001) );
  ANDN U29562 ( .B(n30039), .A(n30040), .Z(n30037) );
  XOR U29563 ( .A(n30038), .B(n30041), .Z(n30039) );
  XOR U29564 ( .A(n30042), .B(n30043), .Z(n30014) );
  XNOR U29565 ( .A(n30009), .B(n30044), .Z(n30043) );
  IV U29566 ( .A(n30012), .Z(n30044) );
  XOR U29567 ( .A(n30045), .B(n30046), .Z(n30012) );
  ANDN U29568 ( .B(n30047), .A(n30048), .Z(n30045) );
  XOR U29569 ( .A(n30046), .B(n30049), .Z(n30047) );
  XNOR U29570 ( .A(n30050), .B(n30051), .Z(n30009) );
  ANDN U29571 ( .B(n30052), .A(n30053), .Z(n30050) );
  XOR U29572 ( .A(n30051), .B(n30054), .Z(n30052) );
  IV U29573 ( .A(n30008), .Z(n30042) );
  XOR U29574 ( .A(n30006), .B(n30055), .Z(n30008) );
  XOR U29575 ( .A(n30056), .B(n30057), .Z(n30055) );
  ANDN U29576 ( .B(n30058), .A(n30059), .Z(n30056) );
  XOR U29577 ( .A(n30060), .B(n30057), .Z(n30058) );
  IV U29578 ( .A(n30010), .Z(n30006) );
  XOR U29579 ( .A(n30061), .B(n30062), .Z(n30010) );
  ANDN U29580 ( .B(n30063), .A(n30064), .Z(n30061) );
  XOR U29581 ( .A(n30065), .B(n30062), .Z(n30063) );
  IV U29582 ( .A(n30020), .Z(n30024) );
  XOR U29583 ( .A(n30020), .B(n29975), .Z(n30022) );
  XOR U29584 ( .A(n30066), .B(n30067), .Z(n29975) );
  AND U29585 ( .A(n782), .B(n30068), .Z(n30066) );
  XOR U29586 ( .A(n30069), .B(n30067), .Z(n30068) );
  NANDN U29587 ( .A(n29977), .B(n29979), .Z(n30020) );
  XOR U29588 ( .A(n30070), .B(n30071), .Z(n29979) );
  AND U29589 ( .A(n782), .B(n30072), .Z(n30070) );
  XOR U29590 ( .A(n30071), .B(n30073), .Z(n30072) );
  XNOR U29591 ( .A(n30074), .B(n30075), .Z(n782) );
  AND U29592 ( .A(n30076), .B(n30077), .Z(n30074) );
  XOR U29593 ( .A(n30075), .B(n29990), .Z(n30077) );
  XNOR U29594 ( .A(n30078), .B(n30079), .Z(n29990) );
  ANDN U29595 ( .B(n30080), .A(n30081), .Z(n30078) );
  XOR U29596 ( .A(n30079), .B(n30082), .Z(n30080) );
  XNOR U29597 ( .A(n30075), .B(n29992), .Z(n30076) );
  XOR U29598 ( .A(n30083), .B(n30084), .Z(n29992) );
  AND U29599 ( .A(n786), .B(n30085), .Z(n30083) );
  XOR U29600 ( .A(n30086), .B(n30084), .Z(n30085) );
  XNOR U29601 ( .A(n30087), .B(n30088), .Z(n30075) );
  AND U29602 ( .A(n30089), .B(n30090), .Z(n30087) );
  XNOR U29603 ( .A(n30088), .B(n30017), .Z(n30090) );
  XOR U29604 ( .A(n30081), .B(n30082), .Z(n30017) );
  XNOR U29605 ( .A(n30091), .B(n30092), .Z(n30082) );
  ANDN U29606 ( .B(n30093), .A(n30094), .Z(n30091) );
  XOR U29607 ( .A(n30095), .B(n30096), .Z(n30093) );
  XOR U29608 ( .A(n30097), .B(n30098), .Z(n30081) );
  XNOR U29609 ( .A(n30099), .B(n30100), .Z(n30098) );
  ANDN U29610 ( .B(n30101), .A(n30102), .Z(n30099) );
  XNOR U29611 ( .A(n30103), .B(n30104), .Z(n30101) );
  IV U29612 ( .A(n30079), .Z(n30097) );
  XOR U29613 ( .A(n30105), .B(n30106), .Z(n30079) );
  ANDN U29614 ( .B(n30107), .A(n30108), .Z(n30105) );
  XOR U29615 ( .A(n30106), .B(n30109), .Z(n30107) );
  XOR U29616 ( .A(n30088), .B(n30019), .Z(n30089) );
  XOR U29617 ( .A(n30110), .B(n30111), .Z(n30019) );
  AND U29618 ( .A(n786), .B(n30112), .Z(n30110) );
  XOR U29619 ( .A(n30113), .B(n30111), .Z(n30112) );
  XNOR U29620 ( .A(n30114), .B(n30115), .Z(n30088) );
  NAND U29621 ( .A(n30116), .B(n30117), .Z(n30115) );
  XOR U29622 ( .A(n30118), .B(n30067), .Z(n30117) );
  XOR U29623 ( .A(n30108), .B(n30109), .Z(n30067) );
  XOR U29624 ( .A(n30119), .B(n30096), .Z(n30109) );
  XOR U29625 ( .A(n30120), .B(n30121), .Z(n30096) );
  ANDN U29626 ( .B(n30122), .A(n30123), .Z(n30120) );
  XOR U29627 ( .A(n30121), .B(n30124), .Z(n30122) );
  IV U29628 ( .A(n30094), .Z(n30119) );
  XOR U29629 ( .A(n30092), .B(n30125), .Z(n30094) );
  XOR U29630 ( .A(n30126), .B(n30127), .Z(n30125) );
  ANDN U29631 ( .B(n30128), .A(n30129), .Z(n30126) );
  XOR U29632 ( .A(n30130), .B(n30127), .Z(n30128) );
  IV U29633 ( .A(n30095), .Z(n30092) );
  XOR U29634 ( .A(n30131), .B(n30132), .Z(n30095) );
  ANDN U29635 ( .B(n30133), .A(n30134), .Z(n30131) );
  XOR U29636 ( .A(n30132), .B(n30135), .Z(n30133) );
  XOR U29637 ( .A(n30136), .B(n30137), .Z(n30108) );
  XNOR U29638 ( .A(n30103), .B(n30138), .Z(n30137) );
  IV U29639 ( .A(n30106), .Z(n30138) );
  XOR U29640 ( .A(n30139), .B(n30140), .Z(n30106) );
  ANDN U29641 ( .B(n30141), .A(n30142), .Z(n30139) );
  XOR U29642 ( .A(n30140), .B(n30143), .Z(n30141) );
  XNOR U29643 ( .A(n30144), .B(n30145), .Z(n30103) );
  ANDN U29644 ( .B(n30146), .A(n30147), .Z(n30144) );
  XOR U29645 ( .A(n30145), .B(n30148), .Z(n30146) );
  IV U29646 ( .A(n30102), .Z(n30136) );
  XOR U29647 ( .A(n30100), .B(n30149), .Z(n30102) );
  XOR U29648 ( .A(n30150), .B(n30151), .Z(n30149) );
  ANDN U29649 ( .B(n30152), .A(n30153), .Z(n30150) );
  XOR U29650 ( .A(n30154), .B(n30151), .Z(n30152) );
  IV U29651 ( .A(n30104), .Z(n30100) );
  XOR U29652 ( .A(n30155), .B(n30156), .Z(n30104) );
  ANDN U29653 ( .B(n30157), .A(n30158), .Z(n30155) );
  XOR U29654 ( .A(n30159), .B(n30156), .Z(n30157) );
  IV U29655 ( .A(n30114), .Z(n30118) );
  XOR U29656 ( .A(n30114), .B(n30069), .Z(n30116) );
  XOR U29657 ( .A(n30160), .B(n30161), .Z(n30069) );
  AND U29658 ( .A(n786), .B(n30162), .Z(n30160) );
  XOR U29659 ( .A(n30163), .B(n30161), .Z(n30162) );
  NANDN U29660 ( .A(n30071), .B(n30073), .Z(n30114) );
  XOR U29661 ( .A(n30164), .B(n30165), .Z(n30073) );
  AND U29662 ( .A(n786), .B(n30166), .Z(n30164) );
  XOR U29663 ( .A(n30165), .B(n30167), .Z(n30166) );
  XNOR U29664 ( .A(n30168), .B(n30169), .Z(n786) );
  AND U29665 ( .A(n30170), .B(n30171), .Z(n30168) );
  XOR U29666 ( .A(n30169), .B(n30084), .Z(n30171) );
  XNOR U29667 ( .A(n30172), .B(n30173), .Z(n30084) );
  ANDN U29668 ( .B(n30174), .A(n30175), .Z(n30172) );
  XOR U29669 ( .A(n30173), .B(n30176), .Z(n30174) );
  XNOR U29670 ( .A(n30169), .B(n30086), .Z(n30170) );
  XOR U29671 ( .A(n30177), .B(n30178), .Z(n30086) );
  AND U29672 ( .A(n790), .B(n30179), .Z(n30177) );
  XOR U29673 ( .A(n30180), .B(n30178), .Z(n30179) );
  XNOR U29674 ( .A(n30181), .B(n30182), .Z(n30169) );
  AND U29675 ( .A(n30183), .B(n30184), .Z(n30181) );
  XNOR U29676 ( .A(n30182), .B(n30111), .Z(n30184) );
  XOR U29677 ( .A(n30175), .B(n30176), .Z(n30111) );
  XNOR U29678 ( .A(n30185), .B(n30186), .Z(n30176) );
  ANDN U29679 ( .B(n30187), .A(n30188), .Z(n30185) );
  XOR U29680 ( .A(n30189), .B(n30190), .Z(n30187) );
  XOR U29681 ( .A(n30191), .B(n30192), .Z(n30175) );
  XNOR U29682 ( .A(n30193), .B(n30194), .Z(n30192) );
  ANDN U29683 ( .B(n30195), .A(n30196), .Z(n30193) );
  XNOR U29684 ( .A(n30197), .B(n30198), .Z(n30195) );
  IV U29685 ( .A(n30173), .Z(n30191) );
  XOR U29686 ( .A(n30199), .B(n30200), .Z(n30173) );
  ANDN U29687 ( .B(n30201), .A(n30202), .Z(n30199) );
  XOR U29688 ( .A(n30200), .B(n30203), .Z(n30201) );
  XOR U29689 ( .A(n30182), .B(n30113), .Z(n30183) );
  XOR U29690 ( .A(n30204), .B(n30205), .Z(n30113) );
  AND U29691 ( .A(n790), .B(n30206), .Z(n30204) );
  XOR U29692 ( .A(n30207), .B(n30205), .Z(n30206) );
  XNOR U29693 ( .A(n30208), .B(n30209), .Z(n30182) );
  NAND U29694 ( .A(n30210), .B(n30211), .Z(n30209) );
  XOR U29695 ( .A(n30212), .B(n30161), .Z(n30211) );
  XOR U29696 ( .A(n30202), .B(n30203), .Z(n30161) );
  XOR U29697 ( .A(n30213), .B(n30190), .Z(n30203) );
  XOR U29698 ( .A(n30214), .B(n30215), .Z(n30190) );
  ANDN U29699 ( .B(n30216), .A(n30217), .Z(n30214) );
  XOR U29700 ( .A(n30215), .B(n30218), .Z(n30216) );
  IV U29701 ( .A(n30188), .Z(n30213) );
  XOR U29702 ( .A(n30186), .B(n30219), .Z(n30188) );
  XOR U29703 ( .A(n30220), .B(n30221), .Z(n30219) );
  ANDN U29704 ( .B(n30222), .A(n30223), .Z(n30220) );
  XOR U29705 ( .A(n30224), .B(n30221), .Z(n30222) );
  IV U29706 ( .A(n30189), .Z(n30186) );
  XOR U29707 ( .A(n30225), .B(n30226), .Z(n30189) );
  ANDN U29708 ( .B(n30227), .A(n30228), .Z(n30225) );
  XOR U29709 ( .A(n30226), .B(n30229), .Z(n30227) );
  XOR U29710 ( .A(n30230), .B(n30231), .Z(n30202) );
  XNOR U29711 ( .A(n30197), .B(n30232), .Z(n30231) );
  IV U29712 ( .A(n30200), .Z(n30232) );
  XOR U29713 ( .A(n30233), .B(n30234), .Z(n30200) );
  ANDN U29714 ( .B(n30235), .A(n30236), .Z(n30233) );
  XOR U29715 ( .A(n30234), .B(n30237), .Z(n30235) );
  XNOR U29716 ( .A(n30238), .B(n30239), .Z(n30197) );
  ANDN U29717 ( .B(n30240), .A(n30241), .Z(n30238) );
  XOR U29718 ( .A(n30239), .B(n30242), .Z(n30240) );
  IV U29719 ( .A(n30196), .Z(n30230) );
  XOR U29720 ( .A(n30194), .B(n30243), .Z(n30196) );
  XOR U29721 ( .A(n30244), .B(n30245), .Z(n30243) );
  ANDN U29722 ( .B(n30246), .A(n30247), .Z(n30244) );
  XOR U29723 ( .A(n30248), .B(n30245), .Z(n30246) );
  IV U29724 ( .A(n30198), .Z(n30194) );
  XOR U29725 ( .A(n30249), .B(n30250), .Z(n30198) );
  ANDN U29726 ( .B(n30251), .A(n30252), .Z(n30249) );
  XOR U29727 ( .A(n30253), .B(n30250), .Z(n30251) );
  IV U29728 ( .A(n30208), .Z(n30212) );
  XOR U29729 ( .A(n30208), .B(n30163), .Z(n30210) );
  XOR U29730 ( .A(n30254), .B(n30255), .Z(n30163) );
  AND U29731 ( .A(n790), .B(n30256), .Z(n30254) );
  XOR U29732 ( .A(n30257), .B(n30255), .Z(n30256) );
  NANDN U29733 ( .A(n30165), .B(n30167), .Z(n30208) );
  XOR U29734 ( .A(n30258), .B(n30259), .Z(n30167) );
  AND U29735 ( .A(n790), .B(n30260), .Z(n30258) );
  XOR U29736 ( .A(n30259), .B(n30261), .Z(n30260) );
  XNOR U29737 ( .A(n30262), .B(n30263), .Z(n790) );
  AND U29738 ( .A(n30264), .B(n30265), .Z(n30262) );
  XOR U29739 ( .A(n30263), .B(n30178), .Z(n30265) );
  XNOR U29740 ( .A(n30266), .B(n30267), .Z(n30178) );
  ANDN U29741 ( .B(n30268), .A(n30269), .Z(n30266) );
  XOR U29742 ( .A(n30267), .B(n30270), .Z(n30268) );
  XNOR U29743 ( .A(n30263), .B(n30180), .Z(n30264) );
  XOR U29744 ( .A(n30271), .B(n30272), .Z(n30180) );
  AND U29745 ( .A(n794), .B(n30273), .Z(n30271) );
  XOR U29746 ( .A(n30274), .B(n30272), .Z(n30273) );
  XNOR U29747 ( .A(n30275), .B(n30276), .Z(n30263) );
  AND U29748 ( .A(n30277), .B(n30278), .Z(n30275) );
  XNOR U29749 ( .A(n30276), .B(n30205), .Z(n30278) );
  XOR U29750 ( .A(n30269), .B(n30270), .Z(n30205) );
  XNOR U29751 ( .A(n30279), .B(n30280), .Z(n30270) );
  ANDN U29752 ( .B(n30281), .A(n30282), .Z(n30279) );
  XOR U29753 ( .A(n30283), .B(n30284), .Z(n30281) );
  XOR U29754 ( .A(n30285), .B(n30286), .Z(n30269) );
  XNOR U29755 ( .A(n30287), .B(n30288), .Z(n30286) );
  ANDN U29756 ( .B(n30289), .A(n30290), .Z(n30287) );
  XNOR U29757 ( .A(n30291), .B(n30292), .Z(n30289) );
  IV U29758 ( .A(n30267), .Z(n30285) );
  XOR U29759 ( .A(n30293), .B(n30294), .Z(n30267) );
  ANDN U29760 ( .B(n30295), .A(n30296), .Z(n30293) );
  XOR U29761 ( .A(n30294), .B(n30297), .Z(n30295) );
  XOR U29762 ( .A(n30276), .B(n30207), .Z(n30277) );
  XOR U29763 ( .A(n30298), .B(n30299), .Z(n30207) );
  AND U29764 ( .A(n794), .B(n30300), .Z(n30298) );
  XOR U29765 ( .A(n30301), .B(n30299), .Z(n30300) );
  XNOR U29766 ( .A(n30302), .B(n30303), .Z(n30276) );
  NAND U29767 ( .A(n30304), .B(n30305), .Z(n30303) );
  XOR U29768 ( .A(n30306), .B(n30255), .Z(n30305) );
  XOR U29769 ( .A(n30296), .B(n30297), .Z(n30255) );
  XOR U29770 ( .A(n30307), .B(n30284), .Z(n30297) );
  XOR U29771 ( .A(n30308), .B(n30309), .Z(n30284) );
  ANDN U29772 ( .B(n30310), .A(n30311), .Z(n30308) );
  XOR U29773 ( .A(n30309), .B(n30312), .Z(n30310) );
  IV U29774 ( .A(n30282), .Z(n30307) );
  XOR U29775 ( .A(n30280), .B(n30313), .Z(n30282) );
  XOR U29776 ( .A(n30314), .B(n30315), .Z(n30313) );
  ANDN U29777 ( .B(n30316), .A(n30317), .Z(n30314) );
  XOR U29778 ( .A(n30318), .B(n30315), .Z(n30316) );
  IV U29779 ( .A(n30283), .Z(n30280) );
  XOR U29780 ( .A(n30319), .B(n30320), .Z(n30283) );
  ANDN U29781 ( .B(n30321), .A(n30322), .Z(n30319) );
  XOR U29782 ( .A(n30320), .B(n30323), .Z(n30321) );
  XOR U29783 ( .A(n30324), .B(n30325), .Z(n30296) );
  XNOR U29784 ( .A(n30291), .B(n30326), .Z(n30325) );
  IV U29785 ( .A(n30294), .Z(n30326) );
  XOR U29786 ( .A(n30327), .B(n30328), .Z(n30294) );
  ANDN U29787 ( .B(n30329), .A(n30330), .Z(n30327) );
  XOR U29788 ( .A(n30328), .B(n30331), .Z(n30329) );
  XNOR U29789 ( .A(n30332), .B(n30333), .Z(n30291) );
  ANDN U29790 ( .B(n30334), .A(n30335), .Z(n30332) );
  XOR U29791 ( .A(n30333), .B(n30336), .Z(n30334) );
  IV U29792 ( .A(n30290), .Z(n30324) );
  XOR U29793 ( .A(n30288), .B(n30337), .Z(n30290) );
  XOR U29794 ( .A(n30338), .B(n30339), .Z(n30337) );
  ANDN U29795 ( .B(n30340), .A(n30341), .Z(n30338) );
  XOR U29796 ( .A(n30342), .B(n30339), .Z(n30340) );
  IV U29797 ( .A(n30292), .Z(n30288) );
  XOR U29798 ( .A(n30343), .B(n30344), .Z(n30292) );
  ANDN U29799 ( .B(n30345), .A(n30346), .Z(n30343) );
  XOR U29800 ( .A(n30347), .B(n30344), .Z(n30345) );
  IV U29801 ( .A(n30302), .Z(n30306) );
  XOR U29802 ( .A(n30302), .B(n30257), .Z(n30304) );
  XOR U29803 ( .A(n30348), .B(n30349), .Z(n30257) );
  AND U29804 ( .A(n794), .B(n30350), .Z(n30348) );
  XOR U29805 ( .A(n30351), .B(n30349), .Z(n30350) );
  NANDN U29806 ( .A(n30259), .B(n30261), .Z(n30302) );
  XOR U29807 ( .A(n30352), .B(n30353), .Z(n30261) );
  AND U29808 ( .A(n794), .B(n30354), .Z(n30352) );
  XOR U29809 ( .A(n30353), .B(n30355), .Z(n30354) );
  XNOR U29810 ( .A(n30356), .B(n30357), .Z(n794) );
  AND U29811 ( .A(n30358), .B(n30359), .Z(n30356) );
  XOR U29812 ( .A(n30357), .B(n30272), .Z(n30359) );
  XNOR U29813 ( .A(n30360), .B(n30361), .Z(n30272) );
  ANDN U29814 ( .B(n30362), .A(n30363), .Z(n30360) );
  XOR U29815 ( .A(n30361), .B(n30364), .Z(n30362) );
  XNOR U29816 ( .A(n30357), .B(n30274), .Z(n30358) );
  XOR U29817 ( .A(n30365), .B(n30366), .Z(n30274) );
  AND U29818 ( .A(n798), .B(n30367), .Z(n30365) );
  XOR U29819 ( .A(n30368), .B(n30366), .Z(n30367) );
  XNOR U29820 ( .A(n30369), .B(n30370), .Z(n30357) );
  AND U29821 ( .A(n30371), .B(n30372), .Z(n30369) );
  XNOR U29822 ( .A(n30370), .B(n30299), .Z(n30372) );
  XOR U29823 ( .A(n30363), .B(n30364), .Z(n30299) );
  XNOR U29824 ( .A(n30373), .B(n30374), .Z(n30364) );
  ANDN U29825 ( .B(n30375), .A(n30376), .Z(n30373) );
  XOR U29826 ( .A(n30377), .B(n30378), .Z(n30375) );
  XOR U29827 ( .A(n30379), .B(n30380), .Z(n30363) );
  XNOR U29828 ( .A(n30381), .B(n30382), .Z(n30380) );
  ANDN U29829 ( .B(n30383), .A(n30384), .Z(n30381) );
  XNOR U29830 ( .A(n30385), .B(n30386), .Z(n30383) );
  IV U29831 ( .A(n30361), .Z(n30379) );
  XOR U29832 ( .A(n30387), .B(n30388), .Z(n30361) );
  ANDN U29833 ( .B(n30389), .A(n30390), .Z(n30387) );
  XOR U29834 ( .A(n30388), .B(n30391), .Z(n30389) );
  XOR U29835 ( .A(n30370), .B(n30301), .Z(n30371) );
  XOR U29836 ( .A(n30392), .B(n30393), .Z(n30301) );
  AND U29837 ( .A(n798), .B(n30394), .Z(n30392) );
  XOR U29838 ( .A(n30395), .B(n30393), .Z(n30394) );
  XNOR U29839 ( .A(n30396), .B(n30397), .Z(n30370) );
  NAND U29840 ( .A(n30398), .B(n30399), .Z(n30397) );
  XOR U29841 ( .A(n30400), .B(n30349), .Z(n30399) );
  XOR U29842 ( .A(n30390), .B(n30391), .Z(n30349) );
  XOR U29843 ( .A(n30401), .B(n30378), .Z(n30391) );
  XOR U29844 ( .A(n30402), .B(n30403), .Z(n30378) );
  ANDN U29845 ( .B(n30404), .A(n30405), .Z(n30402) );
  XOR U29846 ( .A(n30403), .B(n30406), .Z(n30404) );
  IV U29847 ( .A(n30376), .Z(n30401) );
  XOR U29848 ( .A(n30374), .B(n30407), .Z(n30376) );
  XOR U29849 ( .A(n30408), .B(n30409), .Z(n30407) );
  ANDN U29850 ( .B(n30410), .A(n30411), .Z(n30408) );
  XOR U29851 ( .A(n30412), .B(n30409), .Z(n30410) );
  IV U29852 ( .A(n30377), .Z(n30374) );
  XOR U29853 ( .A(n30413), .B(n30414), .Z(n30377) );
  ANDN U29854 ( .B(n30415), .A(n30416), .Z(n30413) );
  XOR U29855 ( .A(n30414), .B(n30417), .Z(n30415) );
  XOR U29856 ( .A(n30418), .B(n30419), .Z(n30390) );
  XNOR U29857 ( .A(n30385), .B(n30420), .Z(n30419) );
  IV U29858 ( .A(n30388), .Z(n30420) );
  XOR U29859 ( .A(n30421), .B(n30422), .Z(n30388) );
  ANDN U29860 ( .B(n30423), .A(n30424), .Z(n30421) );
  XOR U29861 ( .A(n30422), .B(n30425), .Z(n30423) );
  XNOR U29862 ( .A(n30426), .B(n30427), .Z(n30385) );
  ANDN U29863 ( .B(n30428), .A(n30429), .Z(n30426) );
  XOR U29864 ( .A(n30427), .B(n30430), .Z(n30428) );
  IV U29865 ( .A(n30384), .Z(n30418) );
  XOR U29866 ( .A(n30382), .B(n30431), .Z(n30384) );
  XOR U29867 ( .A(n30432), .B(n30433), .Z(n30431) );
  ANDN U29868 ( .B(n30434), .A(n30435), .Z(n30432) );
  XOR U29869 ( .A(n30436), .B(n30433), .Z(n30434) );
  IV U29870 ( .A(n30386), .Z(n30382) );
  XOR U29871 ( .A(n30437), .B(n30438), .Z(n30386) );
  ANDN U29872 ( .B(n30439), .A(n30440), .Z(n30437) );
  XOR U29873 ( .A(n30441), .B(n30438), .Z(n30439) );
  IV U29874 ( .A(n30396), .Z(n30400) );
  XOR U29875 ( .A(n30396), .B(n30351), .Z(n30398) );
  XOR U29876 ( .A(n30442), .B(n30443), .Z(n30351) );
  AND U29877 ( .A(n798), .B(n30444), .Z(n30442) );
  XOR U29878 ( .A(n30445), .B(n30443), .Z(n30444) );
  NANDN U29879 ( .A(n30353), .B(n30355), .Z(n30396) );
  XOR U29880 ( .A(n30446), .B(n30447), .Z(n30355) );
  AND U29881 ( .A(n798), .B(n30448), .Z(n30446) );
  XOR U29882 ( .A(n30447), .B(n30449), .Z(n30448) );
  XNOR U29883 ( .A(n30450), .B(n30451), .Z(n798) );
  AND U29884 ( .A(n30452), .B(n30453), .Z(n30450) );
  XOR U29885 ( .A(n30451), .B(n30366), .Z(n30453) );
  XNOR U29886 ( .A(n30454), .B(n30455), .Z(n30366) );
  ANDN U29887 ( .B(n30456), .A(n30457), .Z(n30454) );
  XOR U29888 ( .A(n30455), .B(n30458), .Z(n30456) );
  XNOR U29889 ( .A(n30451), .B(n30368), .Z(n30452) );
  XOR U29890 ( .A(n30459), .B(n30460), .Z(n30368) );
  AND U29891 ( .A(n802), .B(n30461), .Z(n30459) );
  XOR U29892 ( .A(n30462), .B(n30460), .Z(n30461) );
  XNOR U29893 ( .A(n30463), .B(n30464), .Z(n30451) );
  AND U29894 ( .A(n30465), .B(n30466), .Z(n30463) );
  XNOR U29895 ( .A(n30464), .B(n30393), .Z(n30466) );
  XOR U29896 ( .A(n30457), .B(n30458), .Z(n30393) );
  XNOR U29897 ( .A(n30467), .B(n30468), .Z(n30458) );
  ANDN U29898 ( .B(n30469), .A(n30470), .Z(n30467) );
  XOR U29899 ( .A(n30471), .B(n30472), .Z(n30469) );
  XOR U29900 ( .A(n30473), .B(n30474), .Z(n30457) );
  XNOR U29901 ( .A(n30475), .B(n30476), .Z(n30474) );
  ANDN U29902 ( .B(n30477), .A(n30478), .Z(n30475) );
  XNOR U29903 ( .A(n30479), .B(n30480), .Z(n30477) );
  IV U29904 ( .A(n30455), .Z(n30473) );
  XOR U29905 ( .A(n30481), .B(n30482), .Z(n30455) );
  ANDN U29906 ( .B(n30483), .A(n30484), .Z(n30481) );
  XOR U29907 ( .A(n30482), .B(n30485), .Z(n30483) );
  XOR U29908 ( .A(n30464), .B(n30395), .Z(n30465) );
  XOR U29909 ( .A(n30486), .B(n30487), .Z(n30395) );
  AND U29910 ( .A(n802), .B(n30488), .Z(n30486) );
  XOR U29911 ( .A(n30489), .B(n30487), .Z(n30488) );
  XNOR U29912 ( .A(n30490), .B(n30491), .Z(n30464) );
  NAND U29913 ( .A(n30492), .B(n30493), .Z(n30491) );
  XOR U29914 ( .A(n30494), .B(n30443), .Z(n30493) );
  XOR U29915 ( .A(n30484), .B(n30485), .Z(n30443) );
  XOR U29916 ( .A(n30495), .B(n30472), .Z(n30485) );
  XOR U29917 ( .A(n30496), .B(n30497), .Z(n30472) );
  ANDN U29918 ( .B(n30498), .A(n30499), .Z(n30496) );
  XOR U29919 ( .A(n30497), .B(n30500), .Z(n30498) );
  IV U29920 ( .A(n30470), .Z(n30495) );
  XOR U29921 ( .A(n30468), .B(n30501), .Z(n30470) );
  XOR U29922 ( .A(n30502), .B(n30503), .Z(n30501) );
  ANDN U29923 ( .B(n30504), .A(n30505), .Z(n30502) );
  XOR U29924 ( .A(n30506), .B(n30503), .Z(n30504) );
  IV U29925 ( .A(n30471), .Z(n30468) );
  XOR U29926 ( .A(n30507), .B(n30508), .Z(n30471) );
  ANDN U29927 ( .B(n30509), .A(n30510), .Z(n30507) );
  XOR U29928 ( .A(n30508), .B(n30511), .Z(n30509) );
  XOR U29929 ( .A(n30512), .B(n30513), .Z(n30484) );
  XNOR U29930 ( .A(n30479), .B(n30514), .Z(n30513) );
  IV U29931 ( .A(n30482), .Z(n30514) );
  XOR U29932 ( .A(n30515), .B(n30516), .Z(n30482) );
  ANDN U29933 ( .B(n30517), .A(n30518), .Z(n30515) );
  XOR U29934 ( .A(n30516), .B(n30519), .Z(n30517) );
  XNOR U29935 ( .A(n30520), .B(n30521), .Z(n30479) );
  ANDN U29936 ( .B(n30522), .A(n30523), .Z(n30520) );
  XOR U29937 ( .A(n30521), .B(n30524), .Z(n30522) );
  IV U29938 ( .A(n30478), .Z(n30512) );
  XOR U29939 ( .A(n30476), .B(n30525), .Z(n30478) );
  XOR U29940 ( .A(n30526), .B(n30527), .Z(n30525) );
  ANDN U29941 ( .B(n30528), .A(n30529), .Z(n30526) );
  XOR U29942 ( .A(n30530), .B(n30527), .Z(n30528) );
  IV U29943 ( .A(n30480), .Z(n30476) );
  XOR U29944 ( .A(n30531), .B(n30532), .Z(n30480) );
  ANDN U29945 ( .B(n30533), .A(n30534), .Z(n30531) );
  XOR U29946 ( .A(n30535), .B(n30532), .Z(n30533) );
  IV U29947 ( .A(n30490), .Z(n30494) );
  XOR U29948 ( .A(n30490), .B(n30445), .Z(n30492) );
  XOR U29949 ( .A(n30536), .B(n30537), .Z(n30445) );
  AND U29950 ( .A(n802), .B(n30538), .Z(n30536) );
  XOR U29951 ( .A(n30539), .B(n30537), .Z(n30538) );
  NANDN U29952 ( .A(n30447), .B(n30449), .Z(n30490) );
  XOR U29953 ( .A(n30540), .B(n30541), .Z(n30449) );
  AND U29954 ( .A(n802), .B(n30542), .Z(n30540) );
  XOR U29955 ( .A(n30541), .B(n30543), .Z(n30542) );
  XNOR U29956 ( .A(n30544), .B(n30545), .Z(n802) );
  AND U29957 ( .A(n30546), .B(n30547), .Z(n30544) );
  XOR U29958 ( .A(n30545), .B(n30460), .Z(n30547) );
  XNOR U29959 ( .A(n30548), .B(n30549), .Z(n30460) );
  ANDN U29960 ( .B(n30550), .A(n30551), .Z(n30548) );
  XOR U29961 ( .A(n30549), .B(n30552), .Z(n30550) );
  XNOR U29962 ( .A(n30545), .B(n30462), .Z(n30546) );
  XOR U29963 ( .A(n30553), .B(n30554), .Z(n30462) );
  AND U29964 ( .A(n806), .B(n30555), .Z(n30553) );
  XOR U29965 ( .A(n30556), .B(n30554), .Z(n30555) );
  XNOR U29966 ( .A(n30557), .B(n30558), .Z(n30545) );
  AND U29967 ( .A(n30559), .B(n30560), .Z(n30557) );
  XNOR U29968 ( .A(n30558), .B(n30487), .Z(n30560) );
  XOR U29969 ( .A(n30551), .B(n30552), .Z(n30487) );
  XNOR U29970 ( .A(n30561), .B(n30562), .Z(n30552) );
  ANDN U29971 ( .B(n30563), .A(n30564), .Z(n30561) );
  XOR U29972 ( .A(n30565), .B(n30566), .Z(n30563) );
  XOR U29973 ( .A(n30567), .B(n30568), .Z(n30551) );
  XNOR U29974 ( .A(n30569), .B(n30570), .Z(n30568) );
  ANDN U29975 ( .B(n30571), .A(n30572), .Z(n30569) );
  XNOR U29976 ( .A(n30573), .B(n30574), .Z(n30571) );
  IV U29977 ( .A(n30549), .Z(n30567) );
  XOR U29978 ( .A(n30575), .B(n30576), .Z(n30549) );
  ANDN U29979 ( .B(n30577), .A(n30578), .Z(n30575) );
  XOR U29980 ( .A(n30576), .B(n30579), .Z(n30577) );
  XOR U29981 ( .A(n30558), .B(n30489), .Z(n30559) );
  XOR U29982 ( .A(n30580), .B(n30581), .Z(n30489) );
  AND U29983 ( .A(n806), .B(n30582), .Z(n30580) );
  XOR U29984 ( .A(n30583), .B(n30581), .Z(n30582) );
  XNOR U29985 ( .A(n30584), .B(n30585), .Z(n30558) );
  NAND U29986 ( .A(n30586), .B(n30587), .Z(n30585) );
  XOR U29987 ( .A(n30588), .B(n30537), .Z(n30587) );
  XOR U29988 ( .A(n30578), .B(n30579), .Z(n30537) );
  XOR U29989 ( .A(n30589), .B(n30566), .Z(n30579) );
  XOR U29990 ( .A(n30590), .B(n30591), .Z(n30566) );
  ANDN U29991 ( .B(n30592), .A(n30593), .Z(n30590) );
  XOR U29992 ( .A(n30591), .B(n30594), .Z(n30592) );
  IV U29993 ( .A(n30564), .Z(n30589) );
  XOR U29994 ( .A(n30562), .B(n30595), .Z(n30564) );
  XOR U29995 ( .A(n30596), .B(n30597), .Z(n30595) );
  ANDN U29996 ( .B(n30598), .A(n30599), .Z(n30596) );
  XOR U29997 ( .A(n30600), .B(n30597), .Z(n30598) );
  IV U29998 ( .A(n30565), .Z(n30562) );
  XOR U29999 ( .A(n30601), .B(n30602), .Z(n30565) );
  ANDN U30000 ( .B(n30603), .A(n30604), .Z(n30601) );
  XOR U30001 ( .A(n30602), .B(n30605), .Z(n30603) );
  XOR U30002 ( .A(n30606), .B(n30607), .Z(n30578) );
  XNOR U30003 ( .A(n30573), .B(n30608), .Z(n30607) );
  IV U30004 ( .A(n30576), .Z(n30608) );
  XOR U30005 ( .A(n30609), .B(n30610), .Z(n30576) );
  ANDN U30006 ( .B(n30611), .A(n30612), .Z(n30609) );
  XOR U30007 ( .A(n30610), .B(n30613), .Z(n30611) );
  XNOR U30008 ( .A(n30614), .B(n30615), .Z(n30573) );
  ANDN U30009 ( .B(n30616), .A(n30617), .Z(n30614) );
  XOR U30010 ( .A(n30615), .B(n30618), .Z(n30616) );
  IV U30011 ( .A(n30572), .Z(n30606) );
  XOR U30012 ( .A(n30570), .B(n30619), .Z(n30572) );
  XOR U30013 ( .A(n30620), .B(n30621), .Z(n30619) );
  ANDN U30014 ( .B(n30622), .A(n30623), .Z(n30620) );
  XOR U30015 ( .A(n30624), .B(n30621), .Z(n30622) );
  IV U30016 ( .A(n30574), .Z(n30570) );
  XOR U30017 ( .A(n30625), .B(n30626), .Z(n30574) );
  ANDN U30018 ( .B(n30627), .A(n30628), .Z(n30625) );
  XOR U30019 ( .A(n30629), .B(n30626), .Z(n30627) );
  IV U30020 ( .A(n30584), .Z(n30588) );
  XOR U30021 ( .A(n30584), .B(n30539), .Z(n30586) );
  XOR U30022 ( .A(n30630), .B(n30631), .Z(n30539) );
  AND U30023 ( .A(n806), .B(n30632), .Z(n30630) );
  XOR U30024 ( .A(n30633), .B(n30631), .Z(n30632) );
  NANDN U30025 ( .A(n30541), .B(n30543), .Z(n30584) );
  XOR U30026 ( .A(n30634), .B(n30635), .Z(n30543) );
  AND U30027 ( .A(n806), .B(n30636), .Z(n30634) );
  XOR U30028 ( .A(n30635), .B(n30637), .Z(n30636) );
  XNOR U30029 ( .A(n30638), .B(n30639), .Z(n806) );
  AND U30030 ( .A(n30640), .B(n30641), .Z(n30638) );
  XOR U30031 ( .A(n30639), .B(n30554), .Z(n30641) );
  XNOR U30032 ( .A(n30642), .B(n30643), .Z(n30554) );
  ANDN U30033 ( .B(n30644), .A(n30645), .Z(n30642) );
  XOR U30034 ( .A(n30643), .B(n30646), .Z(n30644) );
  XNOR U30035 ( .A(n30639), .B(n30556), .Z(n30640) );
  XOR U30036 ( .A(n30647), .B(n30648), .Z(n30556) );
  AND U30037 ( .A(n810), .B(n30649), .Z(n30647) );
  XOR U30038 ( .A(n30650), .B(n30648), .Z(n30649) );
  XNOR U30039 ( .A(n30651), .B(n30652), .Z(n30639) );
  AND U30040 ( .A(n30653), .B(n30654), .Z(n30651) );
  XNOR U30041 ( .A(n30652), .B(n30581), .Z(n30654) );
  XOR U30042 ( .A(n30645), .B(n30646), .Z(n30581) );
  XNOR U30043 ( .A(n30655), .B(n30656), .Z(n30646) );
  ANDN U30044 ( .B(n30657), .A(n30658), .Z(n30655) );
  XOR U30045 ( .A(n30659), .B(n30660), .Z(n30657) );
  XOR U30046 ( .A(n30661), .B(n30662), .Z(n30645) );
  XNOR U30047 ( .A(n30663), .B(n30664), .Z(n30662) );
  ANDN U30048 ( .B(n30665), .A(n30666), .Z(n30663) );
  XNOR U30049 ( .A(n30667), .B(n30668), .Z(n30665) );
  IV U30050 ( .A(n30643), .Z(n30661) );
  XOR U30051 ( .A(n30669), .B(n30670), .Z(n30643) );
  ANDN U30052 ( .B(n30671), .A(n30672), .Z(n30669) );
  XOR U30053 ( .A(n30670), .B(n30673), .Z(n30671) );
  XOR U30054 ( .A(n30652), .B(n30583), .Z(n30653) );
  XOR U30055 ( .A(n30674), .B(n30675), .Z(n30583) );
  AND U30056 ( .A(n810), .B(n30676), .Z(n30674) );
  XOR U30057 ( .A(n30677), .B(n30675), .Z(n30676) );
  XNOR U30058 ( .A(n30678), .B(n30679), .Z(n30652) );
  NAND U30059 ( .A(n30680), .B(n30681), .Z(n30679) );
  XOR U30060 ( .A(n30682), .B(n30631), .Z(n30681) );
  XOR U30061 ( .A(n30672), .B(n30673), .Z(n30631) );
  XOR U30062 ( .A(n30683), .B(n30660), .Z(n30673) );
  XOR U30063 ( .A(n30684), .B(n30685), .Z(n30660) );
  ANDN U30064 ( .B(n30686), .A(n30687), .Z(n30684) );
  XOR U30065 ( .A(n30685), .B(n30688), .Z(n30686) );
  IV U30066 ( .A(n30658), .Z(n30683) );
  XOR U30067 ( .A(n30656), .B(n30689), .Z(n30658) );
  XOR U30068 ( .A(n30690), .B(n30691), .Z(n30689) );
  ANDN U30069 ( .B(n30692), .A(n30693), .Z(n30690) );
  XOR U30070 ( .A(n30694), .B(n30691), .Z(n30692) );
  IV U30071 ( .A(n30659), .Z(n30656) );
  XOR U30072 ( .A(n30695), .B(n30696), .Z(n30659) );
  ANDN U30073 ( .B(n30697), .A(n30698), .Z(n30695) );
  XOR U30074 ( .A(n30696), .B(n30699), .Z(n30697) );
  XOR U30075 ( .A(n30700), .B(n30701), .Z(n30672) );
  XNOR U30076 ( .A(n30667), .B(n30702), .Z(n30701) );
  IV U30077 ( .A(n30670), .Z(n30702) );
  XOR U30078 ( .A(n30703), .B(n30704), .Z(n30670) );
  ANDN U30079 ( .B(n30705), .A(n30706), .Z(n30703) );
  XOR U30080 ( .A(n30704), .B(n30707), .Z(n30705) );
  XNOR U30081 ( .A(n30708), .B(n30709), .Z(n30667) );
  ANDN U30082 ( .B(n30710), .A(n30711), .Z(n30708) );
  XOR U30083 ( .A(n30709), .B(n30712), .Z(n30710) );
  IV U30084 ( .A(n30666), .Z(n30700) );
  XOR U30085 ( .A(n30664), .B(n30713), .Z(n30666) );
  XOR U30086 ( .A(n30714), .B(n30715), .Z(n30713) );
  ANDN U30087 ( .B(n30716), .A(n30717), .Z(n30714) );
  XOR U30088 ( .A(n30718), .B(n30715), .Z(n30716) );
  IV U30089 ( .A(n30668), .Z(n30664) );
  XOR U30090 ( .A(n30719), .B(n30720), .Z(n30668) );
  ANDN U30091 ( .B(n30721), .A(n30722), .Z(n30719) );
  XOR U30092 ( .A(n30723), .B(n30720), .Z(n30721) );
  IV U30093 ( .A(n30678), .Z(n30682) );
  XOR U30094 ( .A(n30678), .B(n30633), .Z(n30680) );
  XOR U30095 ( .A(n30724), .B(n30725), .Z(n30633) );
  AND U30096 ( .A(n810), .B(n30726), .Z(n30724) );
  XOR U30097 ( .A(n30727), .B(n30725), .Z(n30726) );
  NANDN U30098 ( .A(n30635), .B(n30637), .Z(n30678) );
  XOR U30099 ( .A(n30728), .B(n30729), .Z(n30637) );
  AND U30100 ( .A(n810), .B(n30730), .Z(n30728) );
  XOR U30101 ( .A(n30729), .B(n30731), .Z(n30730) );
  XNOR U30102 ( .A(n30732), .B(n30733), .Z(n810) );
  AND U30103 ( .A(n30734), .B(n30735), .Z(n30732) );
  XOR U30104 ( .A(n30733), .B(n30648), .Z(n30735) );
  XNOR U30105 ( .A(n30736), .B(n30737), .Z(n30648) );
  ANDN U30106 ( .B(n30738), .A(n30739), .Z(n30736) );
  XOR U30107 ( .A(n30737), .B(n30740), .Z(n30738) );
  XNOR U30108 ( .A(n30733), .B(n30650), .Z(n30734) );
  XOR U30109 ( .A(n30741), .B(n30742), .Z(n30650) );
  AND U30110 ( .A(n814), .B(n30743), .Z(n30741) );
  XOR U30111 ( .A(n30744), .B(n30742), .Z(n30743) );
  XNOR U30112 ( .A(n30745), .B(n30746), .Z(n30733) );
  AND U30113 ( .A(n30747), .B(n30748), .Z(n30745) );
  XNOR U30114 ( .A(n30746), .B(n30675), .Z(n30748) );
  XOR U30115 ( .A(n30739), .B(n30740), .Z(n30675) );
  XNOR U30116 ( .A(n30749), .B(n30750), .Z(n30740) );
  ANDN U30117 ( .B(n30751), .A(n30752), .Z(n30749) );
  XOR U30118 ( .A(n30753), .B(n30754), .Z(n30751) );
  XOR U30119 ( .A(n30755), .B(n30756), .Z(n30739) );
  XNOR U30120 ( .A(n30757), .B(n30758), .Z(n30756) );
  ANDN U30121 ( .B(n30759), .A(n30760), .Z(n30757) );
  XNOR U30122 ( .A(n30761), .B(n30762), .Z(n30759) );
  IV U30123 ( .A(n30737), .Z(n30755) );
  XOR U30124 ( .A(n30763), .B(n30764), .Z(n30737) );
  ANDN U30125 ( .B(n30765), .A(n30766), .Z(n30763) );
  XOR U30126 ( .A(n30764), .B(n30767), .Z(n30765) );
  XOR U30127 ( .A(n30746), .B(n30677), .Z(n30747) );
  XOR U30128 ( .A(n30768), .B(n30769), .Z(n30677) );
  AND U30129 ( .A(n814), .B(n30770), .Z(n30768) );
  XOR U30130 ( .A(n30771), .B(n30769), .Z(n30770) );
  XNOR U30131 ( .A(n30772), .B(n30773), .Z(n30746) );
  NAND U30132 ( .A(n30774), .B(n30775), .Z(n30773) );
  XOR U30133 ( .A(n30776), .B(n30725), .Z(n30775) );
  XOR U30134 ( .A(n30766), .B(n30767), .Z(n30725) );
  XOR U30135 ( .A(n30777), .B(n30754), .Z(n30767) );
  XOR U30136 ( .A(n30778), .B(n30779), .Z(n30754) );
  ANDN U30137 ( .B(n30780), .A(n30781), .Z(n30778) );
  XOR U30138 ( .A(n30779), .B(n30782), .Z(n30780) );
  IV U30139 ( .A(n30752), .Z(n30777) );
  XOR U30140 ( .A(n30750), .B(n30783), .Z(n30752) );
  XOR U30141 ( .A(n30784), .B(n30785), .Z(n30783) );
  ANDN U30142 ( .B(n30786), .A(n30787), .Z(n30784) );
  XOR U30143 ( .A(n30788), .B(n30785), .Z(n30786) );
  IV U30144 ( .A(n30753), .Z(n30750) );
  XOR U30145 ( .A(n30789), .B(n30790), .Z(n30753) );
  ANDN U30146 ( .B(n30791), .A(n30792), .Z(n30789) );
  XOR U30147 ( .A(n30790), .B(n30793), .Z(n30791) );
  XOR U30148 ( .A(n30794), .B(n30795), .Z(n30766) );
  XNOR U30149 ( .A(n30761), .B(n30796), .Z(n30795) );
  IV U30150 ( .A(n30764), .Z(n30796) );
  XOR U30151 ( .A(n30797), .B(n30798), .Z(n30764) );
  ANDN U30152 ( .B(n30799), .A(n30800), .Z(n30797) );
  XOR U30153 ( .A(n30798), .B(n30801), .Z(n30799) );
  XNOR U30154 ( .A(n30802), .B(n30803), .Z(n30761) );
  ANDN U30155 ( .B(n30804), .A(n30805), .Z(n30802) );
  XOR U30156 ( .A(n30803), .B(n30806), .Z(n30804) );
  IV U30157 ( .A(n30760), .Z(n30794) );
  XOR U30158 ( .A(n30758), .B(n30807), .Z(n30760) );
  XOR U30159 ( .A(n30808), .B(n30809), .Z(n30807) );
  ANDN U30160 ( .B(n30810), .A(n30811), .Z(n30808) );
  XOR U30161 ( .A(n30812), .B(n30809), .Z(n30810) );
  IV U30162 ( .A(n30762), .Z(n30758) );
  XOR U30163 ( .A(n30813), .B(n30814), .Z(n30762) );
  ANDN U30164 ( .B(n30815), .A(n30816), .Z(n30813) );
  XOR U30165 ( .A(n30817), .B(n30814), .Z(n30815) );
  IV U30166 ( .A(n30772), .Z(n30776) );
  XOR U30167 ( .A(n30772), .B(n30727), .Z(n30774) );
  XOR U30168 ( .A(n30818), .B(n30819), .Z(n30727) );
  AND U30169 ( .A(n814), .B(n30820), .Z(n30818) );
  XOR U30170 ( .A(n30821), .B(n30819), .Z(n30820) );
  NANDN U30171 ( .A(n30729), .B(n30731), .Z(n30772) );
  XOR U30172 ( .A(n30822), .B(n30823), .Z(n30731) );
  AND U30173 ( .A(n814), .B(n30824), .Z(n30822) );
  XOR U30174 ( .A(n30823), .B(n30825), .Z(n30824) );
  XNOR U30175 ( .A(n30826), .B(n30827), .Z(n814) );
  AND U30176 ( .A(n30828), .B(n30829), .Z(n30826) );
  XOR U30177 ( .A(n30827), .B(n30742), .Z(n30829) );
  XNOR U30178 ( .A(n30830), .B(n30831), .Z(n30742) );
  ANDN U30179 ( .B(n30832), .A(n30833), .Z(n30830) );
  XOR U30180 ( .A(n30831), .B(n30834), .Z(n30832) );
  XNOR U30181 ( .A(n30827), .B(n30744), .Z(n30828) );
  XOR U30182 ( .A(n30835), .B(n30836), .Z(n30744) );
  AND U30183 ( .A(n818), .B(n30837), .Z(n30835) );
  XOR U30184 ( .A(n30838), .B(n30836), .Z(n30837) );
  XNOR U30185 ( .A(n30839), .B(n30840), .Z(n30827) );
  AND U30186 ( .A(n30841), .B(n30842), .Z(n30839) );
  XNOR U30187 ( .A(n30840), .B(n30769), .Z(n30842) );
  XOR U30188 ( .A(n30833), .B(n30834), .Z(n30769) );
  XNOR U30189 ( .A(n30843), .B(n30844), .Z(n30834) );
  ANDN U30190 ( .B(n30845), .A(n30846), .Z(n30843) );
  XOR U30191 ( .A(n30847), .B(n30848), .Z(n30845) );
  XOR U30192 ( .A(n30849), .B(n30850), .Z(n30833) );
  XNOR U30193 ( .A(n30851), .B(n30852), .Z(n30850) );
  ANDN U30194 ( .B(n30853), .A(n30854), .Z(n30851) );
  XNOR U30195 ( .A(n30855), .B(n30856), .Z(n30853) );
  IV U30196 ( .A(n30831), .Z(n30849) );
  XOR U30197 ( .A(n30857), .B(n30858), .Z(n30831) );
  ANDN U30198 ( .B(n30859), .A(n30860), .Z(n30857) );
  XOR U30199 ( .A(n30858), .B(n30861), .Z(n30859) );
  XOR U30200 ( .A(n30840), .B(n30771), .Z(n30841) );
  XOR U30201 ( .A(n30862), .B(n30863), .Z(n30771) );
  AND U30202 ( .A(n818), .B(n30864), .Z(n30862) );
  XOR U30203 ( .A(n30865), .B(n30863), .Z(n30864) );
  XNOR U30204 ( .A(n30866), .B(n30867), .Z(n30840) );
  NAND U30205 ( .A(n30868), .B(n30869), .Z(n30867) );
  XOR U30206 ( .A(n30870), .B(n30819), .Z(n30869) );
  XOR U30207 ( .A(n30860), .B(n30861), .Z(n30819) );
  XOR U30208 ( .A(n30871), .B(n30848), .Z(n30861) );
  XOR U30209 ( .A(n30872), .B(n30873), .Z(n30848) );
  ANDN U30210 ( .B(n30874), .A(n30875), .Z(n30872) );
  XOR U30211 ( .A(n30873), .B(n30876), .Z(n30874) );
  IV U30212 ( .A(n30846), .Z(n30871) );
  XOR U30213 ( .A(n30844), .B(n30877), .Z(n30846) );
  XOR U30214 ( .A(n30878), .B(n30879), .Z(n30877) );
  ANDN U30215 ( .B(n30880), .A(n30881), .Z(n30878) );
  XOR U30216 ( .A(n30882), .B(n30879), .Z(n30880) );
  IV U30217 ( .A(n30847), .Z(n30844) );
  XOR U30218 ( .A(n30883), .B(n30884), .Z(n30847) );
  ANDN U30219 ( .B(n30885), .A(n30886), .Z(n30883) );
  XOR U30220 ( .A(n30884), .B(n30887), .Z(n30885) );
  XOR U30221 ( .A(n30888), .B(n30889), .Z(n30860) );
  XNOR U30222 ( .A(n30855), .B(n30890), .Z(n30889) );
  IV U30223 ( .A(n30858), .Z(n30890) );
  XOR U30224 ( .A(n30891), .B(n30892), .Z(n30858) );
  ANDN U30225 ( .B(n30893), .A(n30894), .Z(n30891) );
  XOR U30226 ( .A(n30892), .B(n30895), .Z(n30893) );
  XNOR U30227 ( .A(n30896), .B(n30897), .Z(n30855) );
  ANDN U30228 ( .B(n30898), .A(n30899), .Z(n30896) );
  XOR U30229 ( .A(n30897), .B(n30900), .Z(n30898) );
  IV U30230 ( .A(n30854), .Z(n30888) );
  XOR U30231 ( .A(n30852), .B(n30901), .Z(n30854) );
  XOR U30232 ( .A(n30902), .B(n30903), .Z(n30901) );
  ANDN U30233 ( .B(n30904), .A(n30905), .Z(n30902) );
  XOR U30234 ( .A(n30906), .B(n30903), .Z(n30904) );
  IV U30235 ( .A(n30856), .Z(n30852) );
  XOR U30236 ( .A(n30907), .B(n30908), .Z(n30856) );
  ANDN U30237 ( .B(n30909), .A(n30910), .Z(n30907) );
  XOR U30238 ( .A(n30911), .B(n30908), .Z(n30909) );
  IV U30239 ( .A(n30866), .Z(n30870) );
  XOR U30240 ( .A(n30866), .B(n30821), .Z(n30868) );
  XOR U30241 ( .A(n30912), .B(n30913), .Z(n30821) );
  AND U30242 ( .A(n818), .B(n30914), .Z(n30912) );
  XOR U30243 ( .A(n30915), .B(n30913), .Z(n30914) );
  NANDN U30244 ( .A(n30823), .B(n30825), .Z(n30866) );
  XOR U30245 ( .A(n30916), .B(n30917), .Z(n30825) );
  AND U30246 ( .A(n818), .B(n30918), .Z(n30916) );
  XOR U30247 ( .A(n30917), .B(n30919), .Z(n30918) );
  XNOR U30248 ( .A(n30920), .B(n30921), .Z(n818) );
  AND U30249 ( .A(n30922), .B(n30923), .Z(n30920) );
  XOR U30250 ( .A(n30921), .B(n30836), .Z(n30923) );
  XNOR U30251 ( .A(n30924), .B(n30925), .Z(n30836) );
  ANDN U30252 ( .B(n30926), .A(n30927), .Z(n30924) );
  XOR U30253 ( .A(n30925), .B(n30928), .Z(n30926) );
  XNOR U30254 ( .A(n30921), .B(n30838), .Z(n30922) );
  XOR U30255 ( .A(n30929), .B(n30930), .Z(n30838) );
  AND U30256 ( .A(n822), .B(n30931), .Z(n30929) );
  XOR U30257 ( .A(n30932), .B(n30930), .Z(n30931) );
  XNOR U30258 ( .A(n30933), .B(n30934), .Z(n30921) );
  AND U30259 ( .A(n30935), .B(n30936), .Z(n30933) );
  XNOR U30260 ( .A(n30934), .B(n30863), .Z(n30936) );
  XOR U30261 ( .A(n30927), .B(n30928), .Z(n30863) );
  XNOR U30262 ( .A(n30937), .B(n30938), .Z(n30928) );
  ANDN U30263 ( .B(n30939), .A(n30940), .Z(n30937) );
  XOR U30264 ( .A(n30941), .B(n30942), .Z(n30939) );
  XOR U30265 ( .A(n30943), .B(n30944), .Z(n30927) );
  XNOR U30266 ( .A(n30945), .B(n30946), .Z(n30944) );
  ANDN U30267 ( .B(n30947), .A(n30948), .Z(n30945) );
  XNOR U30268 ( .A(n30949), .B(n30950), .Z(n30947) );
  IV U30269 ( .A(n30925), .Z(n30943) );
  XOR U30270 ( .A(n30951), .B(n30952), .Z(n30925) );
  ANDN U30271 ( .B(n30953), .A(n30954), .Z(n30951) );
  XOR U30272 ( .A(n30952), .B(n30955), .Z(n30953) );
  XOR U30273 ( .A(n30934), .B(n30865), .Z(n30935) );
  XOR U30274 ( .A(n30956), .B(n30957), .Z(n30865) );
  AND U30275 ( .A(n822), .B(n30958), .Z(n30956) );
  XOR U30276 ( .A(n30959), .B(n30957), .Z(n30958) );
  XNOR U30277 ( .A(n30960), .B(n30961), .Z(n30934) );
  NAND U30278 ( .A(n30962), .B(n30963), .Z(n30961) );
  XOR U30279 ( .A(n30964), .B(n30913), .Z(n30963) );
  XOR U30280 ( .A(n30954), .B(n30955), .Z(n30913) );
  XOR U30281 ( .A(n30965), .B(n30942), .Z(n30955) );
  XOR U30282 ( .A(n30966), .B(n30967), .Z(n30942) );
  ANDN U30283 ( .B(n30968), .A(n30969), .Z(n30966) );
  XOR U30284 ( .A(n30967), .B(n30970), .Z(n30968) );
  IV U30285 ( .A(n30940), .Z(n30965) );
  XOR U30286 ( .A(n30938), .B(n30971), .Z(n30940) );
  XOR U30287 ( .A(n30972), .B(n30973), .Z(n30971) );
  ANDN U30288 ( .B(n30974), .A(n30975), .Z(n30972) );
  XOR U30289 ( .A(n30976), .B(n30973), .Z(n30974) );
  IV U30290 ( .A(n30941), .Z(n30938) );
  XOR U30291 ( .A(n30977), .B(n30978), .Z(n30941) );
  ANDN U30292 ( .B(n30979), .A(n30980), .Z(n30977) );
  XOR U30293 ( .A(n30978), .B(n30981), .Z(n30979) );
  XOR U30294 ( .A(n30982), .B(n30983), .Z(n30954) );
  XNOR U30295 ( .A(n30949), .B(n30984), .Z(n30983) );
  IV U30296 ( .A(n30952), .Z(n30984) );
  XOR U30297 ( .A(n30985), .B(n30986), .Z(n30952) );
  ANDN U30298 ( .B(n30987), .A(n30988), .Z(n30985) );
  XOR U30299 ( .A(n30986), .B(n30989), .Z(n30987) );
  XNOR U30300 ( .A(n30990), .B(n30991), .Z(n30949) );
  ANDN U30301 ( .B(n30992), .A(n30993), .Z(n30990) );
  XOR U30302 ( .A(n30991), .B(n30994), .Z(n30992) );
  IV U30303 ( .A(n30948), .Z(n30982) );
  XOR U30304 ( .A(n30946), .B(n30995), .Z(n30948) );
  XOR U30305 ( .A(n30996), .B(n30997), .Z(n30995) );
  ANDN U30306 ( .B(n30998), .A(n30999), .Z(n30996) );
  XOR U30307 ( .A(n31000), .B(n30997), .Z(n30998) );
  IV U30308 ( .A(n30950), .Z(n30946) );
  XOR U30309 ( .A(n31001), .B(n31002), .Z(n30950) );
  ANDN U30310 ( .B(n31003), .A(n31004), .Z(n31001) );
  XOR U30311 ( .A(n31005), .B(n31002), .Z(n31003) );
  IV U30312 ( .A(n30960), .Z(n30964) );
  XOR U30313 ( .A(n30960), .B(n30915), .Z(n30962) );
  XOR U30314 ( .A(n31006), .B(n31007), .Z(n30915) );
  AND U30315 ( .A(n822), .B(n31008), .Z(n31006) );
  XOR U30316 ( .A(n31009), .B(n31007), .Z(n31008) );
  NANDN U30317 ( .A(n30917), .B(n30919), .Z(n30960) );
  XOR U30318 ( .A(n31010), .B(n31011), .Z(n30919) );
  AND U30319 ( .A(n822), .B(n31012), .Z(n31010) );
  XOR U30320 ( .A(n31011), .B(n31013), .Z(n31012) );
  XNOR U30321 ( .A(n31014), .B(n31015), .Z(n822) );
  AND U30322 ( .A(n31016), .B(n31017), .Z(n31014) );
  XOR U30323 ( .A(n31015), .B(n30930), .Z(n31017) );
  XNOR U30324 ( .A(n31018), .B(n31019), .Z(n30930) );
  ANDN U30325 ( .B(n31020), .A(n31021), .Z(n31018) );
  XOR U30326 ( .A(n31019), .B(n31022), .Z(n31020) );
  XNOR U30327 ( .A(n31015), .B(n30932), .Z(n31016) );
  XOR U30328 ( .A(n31023), .B(n31024), .Z(n30932) );
  AND U30329 ( .A(n826), .B(n31025), .Z(n31023) );
  XOR U30330 ( .A(n31026), .B(n31024), .Z(n31025) );
  XNOR U30331 ( .A(n31027), .B(n31028), .Z(n31015) );
  AND U30332 ( .A(n31029), .B(n31030), .Z(n31027) );
  XNOR U30333 ( .A(n31028), .B(n30957), .Z(n31030) );
  XOR U30334 ( .A(n31021), .B(n31022), .Z(n30957) );
  XNOR U30335 ( .A(n31031), .B(n31032), .Z(n31022) );
  ANDN U30336 ( .B(n31033), .A(n31034), .Z(n31031) );
  XOR U30337 ( .A(n31035), .B(n31036), .Z(n31033) );
  XOR U30338 ( .A(n31037), .B(n31038), .Z(n31021) );
  XNOR U30339 ( .A(n31039), .B(n31040), .Z(n31038) );
  ANDN U30340 ( .B(n31041), .A(n31042), .Z(n31039) );
  XNOR U30341 ( .A(n31043), .B(n31044), .Z(n31041) );
  IV U30342 ( .A(n31019), .Z(n31037) );
  XOR U30343 ( .A(n31045), .B(n31046), .Z(n31019) );
  ANDN U30344 ( .B(n31047), .A(n31048), .Z(n31045) );
  XOR U30345 ( .A(n31046), .B(n31049), .Z(n31047) );
  XOR U30346 ( .A(n31028), .B(n30959), .Z(n31029) );
  XOR U30347 ( .A(n31050), .B(n31051), .Z(n30959) );
  AND U30348 ( .A(n826), .B(n31052), .Z(n31050) );
  XOR U30349 ( .A(n31053), .B(n31051), .Z(n31052) );
  XNOR U30350 ( .A(n31054), .B(n31055), .Z(n31028) );
  NAND U30351 ( .A(n31056), .B(n31057), .Z(n31055) );
  XOR U30352 ( .A(n31058), .B(n31007), .Z(n31057) );
  XOR U30353 ( .A(n31048), .B(n31049), .Z(n31007) );
  XOR U30354 ( .A(n31059), .B(n31036), .Z(n31049) );
  XOR U30355 ( .A(n31060), .B(n31061), .Z(n31036) );
  ANDN U30356 ( .B(n31062), .A(n31063), .Z(n31060) );
  XOR U30357 ( .A(n31061), .B(n31064), .Z(n31062) );
  IV U30358 ( .A(n31034), .Z(n31059) );
  XOR U30359 ( .A(n31032), .B(n31065), .Z(n31034) );
  XOR U30360 ( .A(n31066), .B(n31067), .Z(n31065) );
  ANDN U30361 ( .B(n31068), .A(n31069), .Z(n31066) );
  XOR U30362 ( .A(n31070), .B(n31067), .Z(n31068) );
  IV U30363 ( .A(n31035), .Z(n31032) );
  XOR U30364 ( .A(n31071), .B(n31072), .Z(n31035) );
  ANDN U30365 ( .B(n31073), .A(n31074), .Z(n31071) );
  XOR U30366 ( .A(n31072), .B(n31075), .Z(n31073) );
  XOR U30367 ( .A(n31076), .B(n31077), .Z(n31048) );
  XNOR U30368 ( .A(n31043), .B(n31078), .Z(n31077) );
  IV U30369 ( .A(n31046), .Z(n31078) );
  XOR U30370 ( .A(n31079), .B(n31080), .Z(n31046) );
  ANDN U30371 ( .B(n31081), .A(n31082), .Z(n31079) );
  XOR U30372 ( .A(n31080), .B(n31083), .Z(n31081) );
  XNOR U30373 ( .A(n31084), .B(n31085), .Z(n31043) );
  ANDN U30374 ( .B(n31086), .A(n31087), .Z(n31084) );
  XOR U30375 ( .A(n31085), .B(n31088), .Z(n31086) );
  IV U30376 ( .A(n31042), .Z(n31076) );
  XOR U30377 ( .A(n31040), .B(n31089), .Z(n31042) );
  XOR U30378 ( .A(n31090), .B(n31091), .Z(n31089) );
  ANDN U30379 ( .B(n31092), .A(n31093), .Z(n31090) );
  XOR U30380 ( .A(n31094), .B(n31091), .Z(n31092) );
  IV U30381 ( .A(n31044), .Z(n31040) );
  XOR U30382 ( .A(n31095), .B(n31096), .Z(n31044) );
  ANDN U30383 ( .B(n31097), .A(n31098), .Z(n31095) );
  XOR U30384 ( .A(n31099), .B(n31096), .Z(n31097) );
  IV U30385 ( .A(n31054), .Z(n31058) );
  XOR U30386 ( .A(n31054), .B(n31009), .Z(n31056) );
  XOR U30387 ( .A(n31100), .B(n31101), .Z(n31009) );
  AND U30388 ( .A(n826), .B(n31102), .Z(n31100) );
  XOR U30389 ( .A(n31103), .B(n31101), .Z(n31102) );
  NANDN U30390 ( .A(n31011), .B(n31013), .Z(n31054) );
  XOR U30391 ( .A(n31104), .B(n31105), .Z(n31013) );
  AND U30392 ( .A(n826), .B(n31106), .Z(n31104) );
  XOR U30393 ( .A(n31105), .B(n31107), .Z(n31106) );
  XNOR U30394 ( .A(n31108), .B(n31109), .Z(n826) );
  AND U30395 ( .A(n31110), .B(n31111), .Z(n31108) );
  XOR U30396 ( .A(n31109), .B(n31024), .Z(n31111) );
  XNOR U30397 ( .A(n31112), .B(n31113), .Z(n31024) );
  ANDN U30398 ( .B(n31114), .A(n31115), .Z(n31112) );
  XOR U30399 ( .A(n31113), .B(n31116), .Z(n31114) );
  XNOR U30400 ( .A(n31109), .B(n31026), .Z(n31110) );
  XOR U30401 ( .A(n31117), .B(n31118), .Z(n31026) );
  AND U30402 ( .A(n830), .B(n31119), .Z(n31117) );
  XOR U30403 ( .A(n31120), .B(n31118), .Z(n31119) );
  XNOR U30404 ( .A(n31121), .B(n31122), .Z(n31109) );
  AND U30405 ( .A(n31123), .B(n31124), .Z(n31121) );
  XNOR U30406 ( .A(n31122), .B(n31051), .Z(n31124) );
  XOR U30407 ( .A(n31115), .B(n31116), .Z(n31051) );
  XNOR U30408 ( .A(n31125), .B(n31126), .Z(n31116) );
  ANDN U30409 ( .B(n31127), .A(n31128), .Z(n31125) );
  XOR U30410 ( .A(n31129), .B(n31130), .Z(n31127) );
  XOR U30411 ( .A(n31131), .B(n31132), .Z(n31115) );
  XNOR U30412 ( .A(n31133), .B(n31134), .Z(n31132) );
  ANDN U30413 ( .B(n31135), .A(n31136), .Z(n31133) );
  XNOR U30414 ( .A(n31137), .B(n31138), .Z(n31135) );
  IV U30415 ( .A(n31113), .Z(n31131) );
  XOR U30416 ( .A(n31139), .B(n31140), .Z(n31113) );
  ANDN U30417 ( .B(n31141), .A(n31142), .Z(n31139) );
  XOR U30418 ( .A(n31140), .B(n31143), .Z(n31141) );
  XOR U30419 ( .A(n31122), .B(n31053), .Z(n31123) );
  XOR U30420 ( .A(n31144), .B(n31145), .Z(n31053) );
  AND U30421 ( .A(n830), .B(n31146), .Z(n31144) );
  XOR U30422 ( .A(n31147), .B(n31145), .Z(n31146) );
  XNOR U30423 ( .A(n31148), .B(n31149), .Z(n31122) );
  NAND U30424 ( .A(n31150), .B(n31151), .Z(n31149) );
  XOR U30425 ( .A(n31152), .B(n31101), .Z(n31151) );
  XOR U30426 ( .A(n31142), .B(n31143), .Z(n31101) );
  XOR U30427 ( .A(n31153), .B(n31130), .Z(n31143) );
  XOR U30428 ( .A(n31154), .B(n31155), .Z(n31130) );
  ANDN U30429 ( .B(n31156), .A(n31157), .Z(n31154) );
  XOR U30430 ( .A(n31155), .B(n31158), .Z(n31156) );
  IV U30431 ( .A(n31128), .Z(n31153) );
  XOR U30432 ( .A(n31126), .B(n31159), .Z(n31128) );
  XOR U30433 ( .A(n31160), .B(n31161), .Z(n31159) );
  ANDN U30434 ( .B(n31162), .A(n31163), .Z(n31160) );
  XOR U30435 ( .A(n31164), .B(n31161), .Z(n31162) );
  IV U30436 ( .A(n31129), .Z(n31126) );
  XOR U30437 ( .A(n31165), .B(n31166), .Z(n31129) );
  ANDN U30438 ( .B(n31167), .A(n31168), .Z(n31165) );
  XOR U30439 ( .A(n31166), .B(n31169), .Z(n31167) );
  XOR U30440 ( .A(n31170), .B(n31171), .Z(n31142) );
  XNOR U30441 ( .A(n31137), .B(n31172), .Z(n31171) );
  IV U30442 ( .A(n31140), .Z(n31172) );
  XOR U30443 ( .A(n31173), .B(n31174), .Z(n31140) );
  ANDN U30444 ( .B(n31175), .A(n31176), .Z(n31173) );
  XOR U30445 ( .A(n31174), .B(n31177), .Z(n31175) );
  XNOR U30446 ( .A(n31178), .B(n31179), .Z(n31137) );
  ANDN U30447 ( .B(n31180), .A(n31181), .Z(n31178) );
  XOR U30448 ( .A(n31179), .B(n31182), .Z(n31180) );
  IV U30449 ( .A(n31136), .Z(n31170) );
  XOR U30450 ( .A(n31134), .B(n31183), .Z(n31136) );
  XOR U30451 ( .A(n31184), .B(n31185), .Z(n31183) );
  ANDN U30452 ( .B(n31186), .A(n31187), .Z(n31184) );
  XOR U30453 ( .A(n31188), .B(n31185), .Z(n31186) );
  IV U30454 ( .A(n31138), .Z(n31134) );
  XOR U30455 ( .A(n31189), .B(n31190), .Z(n31138) );
  ANDN U30456 ( .B(n31191), .A(n31192), .Z(n31189) );
  XOR U30457 ( .A(n31193), .B(n31190), .Z(n31191) );
  IV U30458 ( .A(n31148), .Z(n31152) );
  XOR U30459 ( .A(n31148), .B(n31103), .Z(n31150) );
  XOR U30460 ( .A(n31194), .B(n31195), .Z(n31103) );
  AND U30461 ( .A(n830), .B(n31196), .Z(n31194) );
  XOR U30462 ( .A(n31197), .B(n31195), .Z(n31196) );
  NANDN U30463 ( .A(n31105), .B(n31107), .Z(n31148) );
  XOR U30464 ( .A(n31198), .B(n31199), .Z(n31107) );
  AND U30465 ( .A(n830), .B(n31200), .Z(n31198) );
  XOR U30466 ( .A(n31199), .B(n31201), .Z(n31200) );
  XNOR U30467 ( .A(n31202), .B(n31203), .Z(n830) );
  AND U30468 ( .A(n31204), .B(n31205), .Z(n31202) );
  XOR U30469 ( .A(n31203), .B(n31118), .Z(n31205) );
  XNOR U30470 ( .A(n31206), .B(n31207), .Z(n31118) );
  ANDN U30471 ( .B(n31208), .A(n31209), .Z(n31206) );
  XOR U30472 ( .A(n31207), .B(n31210), .Z(n31208) );
  XNOR U30473 ( .A(n31203), .B(n31120), .Z(n31204) );
  XOR U30474 ( .A(n31211), .B(n31212), .Z(n31120) );
  AND U30475 ( .A(n834), .B(n31213), .Z(n31211) );
  XOR U30476 ( .A(n31214), .B(n31212), .Z(n31213) );
  XNOR U30477 ( .A(n31215), .B(n31216), .Z(n31203) );
  AND U30478 ( .A(n31217), .B(n31218), .Z(n31215) );
  XNOR U30479 ( .A(n31216), .B(n31145), .Z(n31218) );
  XOR U30480 ( .A(n31209), .B(n31210), .Z(n31145) );
  XNOR U30481 ( .A(n31219), .B(n31220), .Z(n31210) );
  ANDN U30482 ( .B(n31221), .A(n31222), .Z(n31219) );
  XOR U30483 ( .A(n31223), .B(n31224), .Z(n31221) );
  XOR U30484 ( .A(n31225), .B(n31226), .Z(n31209) );
  XNOR U30485 ( .A(n31227), .B(n31228), .Z(n31226) );
  ANDN U30486 ( .B(n31229), .A(n31230), .Z(n31227) );
  XNOR U30487 ( .A(n31231), .B(n31232), .Z(n31229) );
  IV U30488 ( .A(n31207), .Z(n31225) );
  XOR U30489 ( .A(n31233), .B(n31234), .Z(n31207) );
  ANDN U30490 ( .B(n31235), .A(n31236), .Z(n31233) );
  XOR U30491 ( .A(n31234), .B(n31237), .Z(n31235) );
  XOR U30492 ( .A(n31216), .B(n31147), .Z(n31217) );
  XOR U30493 ( .A(n31238), .B(n31239), .Z(n31147) );
  AND U30494 ( .A(n834), .B(n31240), .Z(n31238) );
  XOR U30495 ( .A(n31241), .B(n31239), .Z(n31240) );
  XNOR U30496 ( .A(n31242), .B(n31243), .Z(n31216) );
  NAND U30497 ( .A(n31244), .B(n31245), .Z(n31243) );
  XOR U30498 ( .A(n31246), .B(n31195), .Z(n31245) );
  XOR U30499 ( .A(n31236), .B(n31237), .Z(n31195) );
  XOR U30500 ( .A(n31247), .B(n31224), .Z(n31237) );
  XOR U30501 ( .A(n31248), .B(n31249), .Z(n31224) );
  ANDN U30502 ( .B(n31250), .A(n31251), .Z(n31248) );
  XOR U30503 ( .A(n31249), .B(n31252), .Z(n31250) );
  IV U30504 ( .A(n31222), .Z(n31247) );
  XOR U30505 ( .A(n31220), .B(n31253), .Z(n31222) );
  XOR U30506 ( .A(n31254), .B(n31255), .Z(n31253) );
  ANDN U30507 ( .B(n31256), .A(n31257), .Z(n31254) );
  XOR U30508 ( .A(n31258), .B(n31255), .Z(n31256) );
  IV U30509 ( .A(n31223), .Z(n31220) );
  XOR U30510 ( .A(n31259), .B(n31260), .Z(n31223) );
  ANDN U30511 ( .B(n31261), .A(n31262), .Z(n31259) );
  XOR U30512 ( .A(n31260), .B(n31263), .Z(n31261) );
  XOR U30513 ( .A(n31264), .B(n31265), .Z(n31236) );
  XNOR U30514 ( .A(n31231), .B(n31266), .Z(n31265) );
  IV U30515 ( .A(n31234), .Z(n31266) );
  XOR U30516 ( .A(n31267), .B(n31268), .Z(n31234) );
  ANDN U30517 ( .B(n31269), .A(n31270), .Z(n31267) );
  XOR U30518 ( .A(n31268), .B(n31271), .Z(n31269) );
  XNOR U30519 ( .A(n31272), .B(n31273), .Z(n31231) );
  ANDN U30520 ( .B(n31274), .A(n31275), .Z(n31272) );
  XOR U30521 ( .A(n31273), .B(n31276), .Z(n31274) );
  IV U30522 ( .A(n31230), .Z(n31264) );
  XOR U30523 ( .A(n31228), .B(n31277), .Z(n31230) );
  XOR U30524 ( .A(n31278), .B(n31279), .Z(n31277) );
  ANDN U30525 ( .B(n31280), .A(n31281), .Z(n31278) );
  XOR U30526 ( .A(n31282), .B(n31279), .Z(n31280) );
  IV U30527 ( .A(n31232), .Z(n31228) );
  XOR U30528 ( .A(n31283), .B(n31284), .Z(n31232) );
  ANDN U30529 ( .B(n31285), .A(n31286), .Z(n31283) );
  XOR U30530 ( .A(n31287), .B(n31284), .Z(n31285) );
  IV U30531 ( .A(n31242), .Z(n31246) );
  XOR U30532 ( .A(n31242), .B(n31197), .Z(n31244) );
  XOR U30533 ( .A(n31288), .B(n31289), .Z(n31197) );
  AND U30534 ( .A(n834), .B(n31290), .Z(n31288) );
  XOR U30535 ( .A(n31291), .B(n31289), .Z(n31290) );
  NANDN U30536 ( .A(n31199), .B(n31201), .Z(n31242) );
  XOR U30537 ( .A(n31292), .B(n31293), .Z(n31201) );
  AND U30538 ( .A(n834), .B(n31294), .Z(n31292) );
  XOR U30539 ( .A(n31293), .B(n31295), .Z(n31294) );
  XNOR U30540 ( .A(n31296), .B(n31297), .Z(n834) );
  AND U30541 ( .A(n31298), .B(n31299), .Z(n31296) );
  XOR U30542 ( .A(n31297), .B(n31212), .Z(n31299) );
  XNOR U30543 ( .A(n31300), .B(n31301), .Z(n31212) );
  ANDN U30544 ( .B(n31302), .A(n31303), .Z(n31300) );
  XOR U30545 ( .A(n31301), .B(n31304), .Z(n31302) );
  XNOR U30546 ( .A(n31297), .B(n31214), .Z(n31298) );
  XOR U30547 ( .A(n31305), .B(n31306), .Z(n31214) );
  AND U30548 ( .A(n838), .B(n31307), .Z(n31305) );
  XOR U30549 ( .A(n31308), .B(n31306), .Z(n31307) );
  XNOR U30550 ( .A(n31309), .B(n31310), .Z(n31297) );
  AND U30551 ( .A(n31311), .B(n31312), .Z(n31309) );
  XNOR U30552 ( .A(n31310), .B(n31239), .Z(n31312) );
  XOR U30553 ( .A(n31303), .B(n31304), .Z(n31239) );
  XNOR U30554 ( .A(n31313), .B(n31314), .Z(n31304) );
  ANDN U30555 ( .B(n31315), .A(n31316), .Z(n31313) );
  XOR U30556 ( .A(n31317), .B(n31318), .Z(n31315) );
  XOR U30557 ( .A(n31319), .B(n31320), .Z(n31303) );
  XNOR U30558 ( .A(n31321), .B(n31322), .Z(n31320) );
  ANDN U30559 ( .B(n31323), .A(n31324), .Z(n31321) );
  XNOR U30560 ( .A(n31325), .B(n31326), .Z(n31323) );
  IV U30561 ( .A(n31301), .Z(n31319) );
  XOR U30562 ( .A(n31327), .B(n31328), .Z(n31301) );
  ANDN U30563 ( .B(n31329), .A(n31330), .Z(n31327) );
  XOR U30564 ( .A(n31328), .B(n31331), .Z(n31329) );
  XOR U30565 ( .A(n31310), .B(n31241), .Z(n31311) );
  XOR U30566 ( .A(n31332), .B(n31333), .Z(n31241) );
  AND U30567 ( .A(n838), .B(n31334), .Z(n31332) );
  XOR U30568 ( .A(n31335), .B(n31333), .Z(n31334) );
  XNOR U30569 ( .A(n31336), .B(n31337), .Z(n31310) );
  NAND U30570 ( .A(n31338), .B(n31339), .Z(n31337) );
  XOR U30571 ( .A(n31340), .B(n31289), .Z(n31339) );
  XOR U30572 ( .A(n31330), .B(n31331), .Z(n31289) );
  XOR U30573 ( .A(n31341), .B(n31318), .Z(n31331) );
  XOR U30574 ( .A(n31342), .B(n31343), .Z(n31318) );
  ANDN U30575 ( .B(n31344), .A(n31345), .Z(n31342) );
  XOR U30576 ( .A(n31343), .B(n31346), .Z(n31344) );
  IV U30577 ( .A(n31316), .Z(n31341) );
  XOR U30578 ( .A(n31314), .B(n31347), .Z(n31316) );
  XOR U30579 ( .A(n31348), .B(n31349), .Z(n31347) );
  ANDN U30580 ( .B(n31350), .A(n31351), .Z(n31348) );
  XOR U30581 ( .A(n31352), .B(n31349), .Z(n31350) );
  IV U30582 ( .A(n31317), .Z(n31314) );
  XOR U30583 ( .A(n31353), .B(n31354), .Z(n31317) );
  ANDN U30584 ( .B(n31355), .A(n31356), .Z(n31353) );
  XOR U30585 ( .A(n31354), .B(n31357), .Z(n31355) );
  XOR U30586 ( .A(n31358), .B(n31359), .Z(n31330) );
  XNOR U30587 ( .A(n31325), .B(n31360), .Z(n31359) );
  IV U30588 ( .A(n31328), .Z(n31360) );
  XOR U30589 ( .A(n31361), .B(n31362), .Z(n31328) );
  ANDN U30590 ( .B(n31363), .A(n31364), .Z(n31361) );
  XOR U30591 ( .A(n31362), .B(n31365), .Z(n31363) );
  XNOR U30592 ( .A(n31366), .B(n31367), .Z(n31325) );
  ANDN U30593 ( .B(n31368), .A(n31369), .Z(n31366) );
  XOR U30594 ( .A(n31367), .B(n31370), .Z(n31368) );
  IV U30595 ( .A(n31324), .Z(n31358) );
  XOR U30596 ( .A(n31322), .B(n31371), .Z(n31324) );
  XOR U30597 ( .A(n31372), .B(n31373), .Z(n31371) );
  ANDN U30598 ( .B(n31374), .A(n31375), .Z(n31372) );
  XOR U30599 ( .A(n31376), .B(n31373), .Z(n31374) );
  IV U30600 ( .A(n31326), .Z(n31322) );
  XOR U30601 ( .A(n31377), .B(n31378), .Z(n31326) );
  ANDN U30602 ( .B(n31379), .A(n31380), .Z(n31377) );
  XOR U30603 ( .A(n31381), .B(n31378), .Z(n31379) );
  IV U30604 ( .A(n31336), .Z(n31340) );
  XOR U30605 ( .A(n31336), .B(n31291), .Z(n31338) );
  XOR U30606 ( .A(n31382), .B(n31383), .Z(n31291) );
  AND U30607 ( .A(n838), .B(n31384), .Z(n31382) );
  XOR U30608 ( .A(n31385), .B(n31383), .Z(n31384) );
  NANDN U30609 ( .A(n31293), .B(n31295), .Z(n31336) );
  XOR U30610 ( .A(n31386), .B(n31387), .Z(n31295) );
  AND U30611 ( .A(n838), .B(n31388), .Z(n31386) );
  XOR U30612 ( .A(n31387), .B(n31389), .Z(n31388) );
  XNOR U30613 ( .A(n31390), .B(n31391), .Z(n838) );
  AND U30614 ( .A(n31392), .B(n31393), .Z(n31390) );
  XOR U30615 ( .A(n31391), .B(n31306), .Z(n31393) );
  XNOR U30616 ( .A(n31394), .B(n31395), .Z(n31306) );
  ANDN U30617 ( .B(n31396), .A(n31397), .Z(n31394) );
  XOR U30618 ( .A(n31395), .B(n31398), .Z(n31396) );
  XNOR U30619 ( .A(n31391), .B(n31308), .Z(n31392) );
  XOR U30620 ( .A(n31399), .B(n31400), .Z(n31308) );
  AND U30621 ( .A(n842), .B(n31401), .Z(n31399) );
  XOR U30622 ( .A(n31402), .B(n31400), .Z(n31401) );
  XNOR U30623 ( .A(n31403), .B(n31404), .Z(n31391) );
  AND U30624 ( .A(n31405), .B(n31406), .Z(n31403) );
  XNOR U30625 ( .A(n31404), .B(n31333), .Z(n31406) );
  XOR U30626 ( .A(n31397), .B(n31398), .Z(n31333) );
  XNOR U30627 ( .A(n31407), .B(n31408), .Z(n31398) );
  ANDN U30628 ( .B(n31409), .A(n31410), .Z(n31407) );
  XOR U30629 ( .A(n31411), .B(n31412), .Z(n31409) );
  XOR U30630 ( .A(n31413), .B(n31414), .Z(n31397) );
  XNOR U30631 ( .A(n31415), .B(n31416), .Z(n31414) );
  ANDN U30632 ( .B(n31417), .A(n31418), .Z(n31415) );
  XNOR U30633 ( .A(n31419), .B(n31420), .Z(n31417) );
  IV U30634 ( .A(n31395), .Z(n31413) );
  XOR U30635 ( .A(n31421), .B(n31422), .Z(n31395) );
  ANDN U30636 ( .B(n31423), .A(n31424), .Z(n31421) );
  XOR U30637 ( .A(n31422), .B(n31425), .Z(n31423) );
  XOR U30638 ( .A(n31404), .B(n31335), .Z(n31405) );
  XOR U30639 ( .A(n31426), .B(n31427), .Z(n31335) );
  AND U30640 ( .A(n842), .B(n31428), .Z(n31426) );
  XOR U30641 ( .A(n31429), .B(n31427), .Z(n31428) );
  XNOR U30642 ( .A(n31430), .B(n31431), .Z(n31404) );
  NAND U30643 ( .A(n31432), .B(n31433), .Z(n31431) );
  XOR U30644 ( .A(n31434), .B(n31383), .Z(n31433) );
  XOR U30645 ( .A(n31424), .B(n31425), .Z(n31383) );
  XOR U30646 ( .A(n31435), .B(n31412), .Z(n31425) );
  XOR U30647 ( .A(n31436), .B(n31437), .Z(n31412) );
  ANDN U30648 ( .B(n31438), .A(n31439), .Z(n31436) );
  XOR U30649 ( .A(n31437), .B(n31440), .Z(n31438) );
  IV U30650 ( .A(n31410), .Z(n31435) );
  XOR U30651 ( .A(n31408), .B(n31441), .Z(n31410) );
  XOR U30652 ( .A(n31442), .B(n31443), .Z(n31441) );
  ANDN U30653 ( .B(n31444), .A(n31445), .Z(n31442) );
  XOR U30654 ( .A(n31446), .B(n31443), .Z(n31444) );
  IV U30655 ( .A(n31411), .Z(n31408) );
  XOR U30656 ( .A(n31447), .B(n31448), .Z(n31411) );
  ANDN U30657 ( .B(n31449), .A(n31450), .Z(n31447) );
  XOR U30658 ( .A(n31448), .B(n31451), .Z(n31449) );
  XOR U30659 ( .A(n31452), .B(n31453), .Z(n31424) );
  XNOR U30660 ( .A(n31419), .B(n31454), .Z(n31453) );
  IV U30661 ( .A(n31422), .Z(n31454) );
  XOR U30662 ( .A(n31455), .B(n31456), .Z(n31422) );
  ANDN U30663 ( .B(n31457), .A(n31458), .Z(n31455) );
  XOR U30664 ( .A(n31456), .B(n31459), .Z(n31457) );
  XNOR U30665 ( .A(n31460), .B(n31461), .Z(n31419) );
  ANDN U30666 ( .B(n31462), .A(n31463), .Z(n31460) );
  XOR U30667 ( .A(n31461), .B(n31464), .Z(n31462) );
  IV U30668 ( .A(n31418), .Z(n31452) );
  XOR U30669 ( .A(n31416), .B(n31465), .Z(n31418) );
  XOR U30670 ( .A(n31466), .B(n31467), .Z(n31465) );
  ANDN U30671 ( .B(n31468), .A(n31469), .Z(n31466) );
  XOR U30672 ( .A(n31470), .B(n31467), .Z(n31468) );
  IV U30673 ( .A(n31420), .Z(n31416) );
  XOR U30674 ( .A(n31471), .B(n31472), .Z(n31420) );
  ANDN U30675 ( .B(n31473), .A(n31474), .Z(n31471) );
  XOR U30676 ( .A(n31475), .B(n31472), .Z(n31473) );
  IV U30677 ( .A(n31430), .Z(n31434) );
  XOR U30678 ( .A(n31430), .B(n31385), .Z(n31432) );
  XOR U30679 ( .A(n31476), .B(n31477), .Z(n31385) );
  AND U30680 ( .A(n842), .B(n31478), .Z(n31476) );
  XOR U30681 ( .A(n31479), .B(n31477), .Z(n31478) );
  NANDN U30682 ( .A(n31387), .B(n31389), .Z(n31430) );
  XOR U30683 ( .A(n31480), .B(n31481), .Z(n31389) );
  AND U30684 ( .A(n842), .B(n31482), .Z(n31480) );
  XOR U30685 ( .A(n31481), .B(n31483), .Z(n31482) );
  XNOR U30686 ( .A(n31484), .B(n31485), .Z(n842) );
  AND U30687 ( .A(n31486), .B(n31487), .Z(n31484) );
  XOR U30688 ( .A(n31485), .B(n31400), .Z(n31487) );
  XNOR U30689 ( .A(n31488), .B(n31489), .Z(n31400) );
  ANDN U30690 ( .B(n31490), .A(n31491), .Z(n31488) );
  XOR U30691 ( .A(n31489), .B(n31492), .Z(n31490) );
  XNOR U30692 ( .A(n31485), .B(n31402), .Z(n31486) );
  XOR U30693 ( .A(n31493), .B(n31494), .Z(n31402) );
  AND U30694 ( .A(n846), .B(n31495), .Z(n31493) );
  XOR U30695 ( .A(n31496), .B(n31494), .Z(n31495) );
  XNOR U30696 ( .A(n31497), .B(n31498), .Z(n31485) );
  AND U30697 ( .A(n31499), .B(n31500), .Z(n31497) );
  XNOR U30698 ( .A(n31498), .B(n31427), .Z(n31500) );
  XOR U30699 ( .A(n31491), .B(n31492), .Z(n31427) );
  XNOR U30700 ( .A(n31501), .B(n31502), .Z(n31492) );
  ANDN U30701 ( .B(n31503), .A(n31504), .Z(n31501) );
  XOR U30702 ( .A(n31505), .B(n31506), .Z(n31503) );
  XOR U30703 ( .A(n31507), .B(n31508), .Z(n31491) );
  XNOR U30704 ( .A(n31509), .B(n31510), .Z(n31508) );
  ANDN U30705 ( .B(n31511), .A(n31512), .Z(n31509) );
  XNOR U30706 ( .A(n31513), .B(n31514), .Z(n31511) );
  IV U30707 ( .A(n31489), .Z(n31507) );
  XOR U30708 ( .A(n31515), .B(n31516), .Z(n31489) );
  ANDN U30709 ( .B(n31517), .A(n31518), .Z(n31515) );
  XOR U30710 ( .A(n31516), .B(n31519), .Z(n31517) );
  XOR U30711 ( .A(n31498), .B(n31429), .Z(n31499) );
  XOR U30712 ( .A(n31520), .B(n31521), .Z(n31429) );
  AND U30713 ( .A(n846), .B(n31522), .Z(n31520) );
  XOR U30714 ( .A(n31523), .B(n31521), .Z(n31522) );
  XNOR U30715 ( .A(n31524), .B(n31525), .Z(n31498) );
  NAND U30716 ( .A(n31526), .B(n31527), .Z(n31525) );
  XOR U30717 ( .A(n31528), .B(n31477), .Z(n31527) );
  XOR U30718 ( .A(n31518), .B(n31519), .Z(n31477) );
  XOR U30719 ( .A(n31529), .B(n31506), .Z(n31519) );
  XOR U30720 ( .A(n31530), .B(n31531), .Z(n31506) );
  ANDN U30721 ( .B(n31532), .A(n31533), .Z(n31530) );
  XOR U30722 ( .A(n31531), .B(n31534), .Z(n31532) );
  IV U30723 ( .A(n31504), .Z(n31529) );
  XOR U30724 ( .A(n31502), .B(n31535), .Z(n31504) );
  XOR U30725 ( .A(n31536), .B(n31537), .Z(n31535) );
  ANDN U30726 ( .B(n31538), .A(n31539), .Z(n31536) );
  XOR U30727 ( .A(n31540), .B(n31537), .Z(n31538) );
  IV U30728 ( .A(n31505), .Z(n31502) );
  XOR U30729 ( .A(n31541), .B(n31542), .Z(n31505) );
  ANDN U30730 ( .B(n31543), .A(n31544), .Z(n31541) );
  XOR U30731 ( .A(n31542), .B(n31545), .Z(n31543) );
  XOR U30732 ( .A(n31546), .B(n31547), .Z(n31518) );
  XNOR U30733 ( .A(n31513), .B(n31548), .Z(n31547) );
  IV U30734 ( .A(n31516), .Z(n31548) );
  XOR U30735 ( .A(n31549), .B(n31550), .Z(n31516) );
  ANDN U30736 ( .B(n31551), .A(n31552), .Z(n31549) );
  XOR U30737 ( .A(n31550), .B(n31553), .Z(n31551) );
  XNOR U30738 ( .A(n31554), .B(n31555), .Z(n31513) );
  ANDN U30739 ( .B(n31556), .A(n31557), .Z(n31554) );
  XOR U30740 ( .A(n31555), .B(n31558), .Z(n31556) );
  IV U30741 ( .A(n31512), .Z(n31546) );
  XOR U30742 ( .A(n31510), .B(n31559), .Z(n31512) );
  XOR U30743 ( .A(n31560), .B(n31561), .Z(n31559) );
  ANDN U30744 ( .B(n31562), .A(n31563), .Z(n31560) );
  XOR U30745 ( .A(n31564), .B(n31561), .Z(n31562) );
  IV U30746 ( .A(n31514), .Z(n31510) );
  XOR U30747 ( .A(n31565), .B(n31566), .Z(n31514) );
  ANDN U30748 ( .B(n31567), .A(n31568), .Z(n31565) );
  XOR U30749 ( .A(n31569), .B(n31566), .Z(n31567) );
  IV U30750 ( .A(n31524), .Z(n31528) );
  XOR U30751 ( .A(n31524), .B(n31479), .Z(n31526) );
  XOR U30752 ( .A(n31570), .B(n31571), .Z(n31479) );
  AND U30753 ( .A(n846), .B(n31572), .Z(n31570) );
  XOR U30754 ( .A(n31573), .B(n31571), .Z(n31572) );
  NANDN U30755 ( .A(n31481), .B(n31483), .Z(n31524) );
  XOR U30756 ( .A(n31574), .B(n31575), .Z(n31483) );
  AND U30757 ( .A(n846), .B(n31576), .Z(n31574) );
  XOR U30758 ( .A(n31575), .B(n31577), .Z(n31576) );
  XNOR U30759 ( .A(n31578), .B(n31579), .Z(n846) );
  AND U30760 ( .A(n31580), .B(n31581), .Z(n31578) );
  XOR U30761 ( .A(n31579), .B(n31494), .Z(n31581) );
  XNOR U30762 ( .A(n31582), .B(n31583), .Z(n31494) );
  ANDN U30763 ( .B(n31584), .A(n31585), .Z(n31582) );
  XOR U30764 ( .A(n31583), .B(n31586), .Z(n31584) );
  XNOR U30765 ( .A(n31579), .B(n31496), .Z(n31580) );
  XOR U30766 ( .A(n31587), .B(n31588), .Z(n31496) );
  AND U30767 ( .A(n850), .B(n31589), .Z(n31587) );
  XOR U30768 ( .A(n31590), .B(n31588), .Z(n31589) );
  XNOR U30769 ( .A(n31591), .B(n31592), .Z(n31579) );
  AND U30770 ( .A(n31593), .B(n31594), .Z(n31591) );
  XNOR U30771 ( .A(n31592), .B(n31521), .Z(n31594) );
  XOR U30772 ( .A(n31585), .B(n31586), .Z(n31521) );
  XNOR U30773 ( .A(n31595), .B(n31596), .Z(n31586) );
  ANDN U30774 ( .B(n31597), .A(n31598), .Z(n31595) );
  XOR U30775 ( .A(n31599), .B(n31600), .Z(n31597) );
  XOR U30776 ( .A(n31601), .B(n31602), .Z(n31585) );
  XNOR U30777 ( .A(n31603), .B(n31604), .Z(n31602) );
  ANDN U30778 ( .B(n31605), .A(n31606), .Z(n31603) );
  XNOR U30779 ( .A(n31607), .B(n31608), .Z(n31605) );
  IV U30780 ( .A(n31583), .Z(n31601) );
  XOR U30781 ( .A(n31609), .B(n31610), .Z(n31583) );
  ANDN U30782 ( .B(n31611), .A(n31612), .Z(n31609) );
  XOR U30783 ( .A(n31610), .B(n31613), .Z(n31611) );
  XOR U30784 ( .A(n31592), .B(n31523), .Z(n31593) );
  XOR U30785 ( .A(n31614), .B(n31615), .Z(n31523) );
  AND U30786 ( .A(n850), .B(n31616), .Z(n31614) );
  XOR U30787 ( .A(n31617), .B(n31615), .Z(n31616) );
  XNOR U30788 ( .A(n31618), .B(n31619), .Z(n31592) );
  NAND U30789 ( .A(n31620), .B(n31621), .Z(n31619) );
  XOR U30790 ( .A(n31622), .B(n31571), .Z(n31621) );
  XOR U30791 ( .A(n31612), .B(n31613), .Z(n31571) );
  XOR U30792 ( .A(n31623), .B(n31600), .Z(n31613) );
  XOR U30793 ( .A(n31624), .B(n31625), .Z(n31600) );
  ANDN U30794 ( .B(n31626), .A(n31627), .Z(n31624) );
  XOR U30795 ( .A(n31625), .B(n31628), .Z(n31626) );
  IV U30796 ( .A(n31598), .Z(n31623) );
  XOR U30797 ( .A(n31596), .B(n31629), .Z(n31598) );
  XOR U30798 ( .A(n31630), .B(n31631), .Z(n31629) );
  ANDN U30799 ( .B(n31632), .A(n31633), .Z(n31630) );
  XOR U30800 ( .A(n31634), .B(n31631), .Z(n31632) );
  IV U30801 ( .A(n31599), .Z(n31596) );
  XOR U30802 ( .A(n31635), .B(n31636), .Z(n31599) );
  ANDN U30803 ( .B(n31637), .A(n31638), .Z(n31635) );
  XOR U30804 ( .A(n31636), .B(n31639), .Z(n31637) );
  XOR U30805 ( .A(n31640), .B(n31641), .Z(n31612) );
  XNOR U30806 ( .A(n31607), .B(n31642), .Z(n31641) );
  IV U30807 ( .A(n31610), .Z(n31642) );
  XOR U30808 ( .A(n31643), .B(n31644), .Z(n31610) );
  ANDN U30809 ( .B(n31645), .A(n31646), .Z(n31643) );
  XOR U30810 ( .A(n31644), .B(n31647), .Z(n31645) );
  XNOR U30811 ( .A(n31648), .B(n31649), .Z(n31607) );
  ANDN U30812 ( .B(n31650), .A(n31651), .Z(n31648) );
  XOR U30813 ( .A(n31649), .B(n31652), .Z(n31650) );
  IV U30814 ( .A(n31606), .Z(n31640) );
  XOR U30815 ( .A(n31604), .B(n31653), .Z(n31606) );
  XOR U30816 ( .A(n31654), .B(n31655), .Z(n31653) );
  ANDN U30817 ( .B(n31656), .A(n31657), .Z(n31654) );
  XOR U30818 ( .A(n31658), .B(n31655), .Z(n31656) );
  IV U30819 ( .A(n31608), .Z(n31604) );
  XOR U30820 ( .A(n31659), .B(n31660), .Z(n31608) );
  ANDN U30821 ( .B(n31661), .A(n31662), .Z(n31659) );
  XOR U30822 ( .A(n31663), .B(n31660), .Z(n31661) );
  IV U30823 ( .A(n31618), .Z(n31622) );
  XOR U30824 ( .A(n31618), .B(n31573), .Z(n31620) );
  XOR U30825 ( .A(n31664), .B(n31665), .Z(n31573) );
  AND U30826 ( .A(n850), .B(n31666), .Z(n31664) );
  XOR U30827 ( .A(n31667), .B(n31665), .Z(n31666) );
  NANDN U30828 ( .A(n31575), .B(n31577), .Z(n31618) );
  XOR U30829 ( .A(n31668), .B(n31669), .Z(n31577) );
  AND U30830 ( .A(n850), .B(n31670), .Z(n31668) );
  XOR U30831 ( .A(n31669), .B(n31671), .Z(n31670) );
  XNOR U30832 ( .A(n31672), .B(n31673), .Z(n850) );
  AND U30833 ( .A(n31674), .B(n31675), .Z(n31672) );
  XOR U30834 ( .A(n31673), .B(n31588), .Z(n31675) );
  XNOR U30835 ( .A(n31676), .B(n31677), .Z(n31588) );
  ANDN U30836 ( .B(n31678), .A(n31679), .Z(n31676) );
  XOR U30837 ( .A(n31677), .B(n31680), .Z(n31678) );
  XNOR U30838 ( .A(n31673), .B(n31590), .Z(n31674) );
  XOR U30839 ( .A(n31681), .B(n31682), .Z(n31590) );
  AND U30840 ( .A(n854), .B(n31683), .Z(n31681) );
  XOR U30841 ( .A(n31684), .B(n31682), .Z(n31683) );
  XNOR U30842 ( .A(n31685), .B(n31686), .Z(n31673) );
  AND U30843 ( .A(n31687), .B(n31688), .Z(n31685) );
  XNOR U30844 ( .A(n31686), .B(n31615), .Z(n31688) );
  XOR U30845 ( .A(n31679), .B(n31680), .Z(n31615) );
  XNOR U30846 ( .A(n31689), .B(n31690), .Z(n31680) );
  ANDN U30847 ( .B(n31691), .A(n31692), .Z(n31689) );
  XOR U30848 ( .A(n31693), .B(n31694), .Z(n31691) );
  XOR U30849 ( .A(n31695), .B(n31696), .Z(n31679) );
  XNOR U30850 ( .A(n31697), .B(n31698), .Z(n31696) );
  ANDN U30851 ( .B(n31699), .A(n31700), .Z(n31697) );
  XNOR U30852 ( .A(n31701), .B(n31702), .Z(n31699) );
  IV U30853 ( .A(n31677), .Z(n31695) );
  XOR U30854 ( .A(n31703), .B(n31704), .Z(n31677) );
  ANDN U30855 ( .B(n31705), .A(n31706), .Z(n31703) );
  XOR U30856 ( .A(n31704), .B(n31707), .Z(n31705) );
  XOR U30857 ( .A(n31686), .B(n31617), .Z(n31687) );
  XOR U30858 ( .A(n31708), .B(n31709), .Z(n31617) );
  AND U30859 ( .A(n854), .B(n31710), .Z(n31708) );
  XOR U30860 ( .A(n31711), .B(n31709), .Z(n31710) );
  XNOR U30861 ( .A(n31712), .B(n31713), .Z(n31686) );
  NAND U30862 ( .A(n31714), .B(n31715), .Z(n31713) );
  XOR U30863 ( .A(n31716), .B(n31665), .Z(n31715) );
  XOR U30864 ( .A(n31706), .B(n31707), .Z(n31665) );
  XOR U30865 ( .A(n31717), .B(n31694), .Z(n31707) );
  XOR U30866 ( .A(n31718), .B(n31719), .Z(n31694) );
  ANDN U30867 ( .B(n31720), .A(n31721), .Z(n31718) );
  XOR U30868 ( .A(n31719), .B(n31722), .Z(n31720) );
  IV U30869 ( .A(n31692), .Z(n31717) );
  XOR U30870 ( .A(n31690), .B(n31723), .Z(n31692) );
  XOR U30871 ( .A(n31724), .B(n31725), .Z(n31723) );
  ANDN U30872 ( .B(n31726), .A(n31727), .Z(n31724) );
  XOR U30873 ( .A(n31728), .B(n31725), .Z(n31726) );
  IV U30874 ( .A(n31693), .Z(n31690) );
  XOR U30875 ( .A(n31729), .B(n31730), .Z(n31693) );
  ANDN U30876 ( .B(n31731), .A(n31732), .Z(n31729) );
  XOR U30877 ( .A(n31730), .B(n31733), .Z(n31731) );
  XOR U30878 ( .A(n31734), .B(n31735), .Z(n31706) );
  XNOR U30879 ( .A(n31701), .B(n31736), .Z(n31735) );
  IV U30880 ( .A(n31704), .Z(n31736) );
  XOR U30881 ( .A(n31737), .B(n31738), .Z(n31704) );
  ANDN U30882 ( .B(n31739), .A(n31740), .Z(n31737) );
  XOR U30883 ( .A(n31738), .B(n31741), .Z(n31739) );
  XNOR U30884 ( .A(n31742), .B(n31743), .Z(n31701) );
  ANDN U30885 ( .B(n31744), .A(n31745), .Z(n31742) );
  XOR U30886 ( .A(n31743), .B(n31746), .Z(n31744) );
  IV U30887 ( .A(n31700), .Z(n31734) );
  XOR U30888 ( .A(n31698), .B(n31747), .Z(n31700) );
  XOR U30889 ( .A(n31748), .B(n31749), .Z(n31747) );
  ANDN U30890 ( .B(n31750), .A(n31751), .Z(n31748) );
  XOR U30891 ( .A(n31752), .B(n31749), .Z(n31750) );
  IV U30892 ( .A(n31702), .Z(n31698) );
  XOR U30893 ( .A(n31753), .B(n31754), .Z(n31702) );
  ANDN U30894 ( .B(n31755), .A(n31756), .Z(n31753) );
  XOR U30895 ( .A(n31757), .B(n31754), .Z(n31755) );
  IV U30896 ( .A(n31712), .Z(n31716) );
  XOR U30897 ( .A(n31712), .B(n31667), .Z(n31714) );
  XOR U30898 ( .A(n31758), .B(n31759), .Z(n31667) );
  AND U30899 ( .A(n854), .B(n31760), .Z(n31758) );
  XOR U30900 ( .A(n31761), .B(n31759), .Z(n31760) );
  NANDN U30901 ( .A(n31669), .B(n31671), .Z(n31712) );
  XOR U30902 ( .A(n31762), .B(n31763), .Z(n31671) );
  AND U30903 ( .A(n854), .B(n31764), .Z(n31762) );
  XOR U30904 ( .A(n31763), .B(n31765), .Z(n31764) );
  XNOR U30905 ( .A(n31766), .B(n31767), .Z(n854) );
  AND U30906 ( .A(n31768), .B(n31769), .Z(n31766) );
  XOR U30907 ( .A(n31767), .B(n31682), .Z(n31769) );
  XNOR U30908 ( .A(n31770), .B(n31771), .Z(n31682) );
  ANDN U30909 ( .B(n31772), .A(n31773), .Z(n31770) );
  XOR U30910 ( .A(n31771), .B(n31774), .Z(n31772) );
  XNOR U30911 ( .A(n31767), .B(n31684), .Z(n31768) );
  XOR U30912 ( .A(n31775), .B(n31776), .Z(n31684) );
  AND U30913 ( .A(n858), .B(n31777), .Z(n31775) );
  XOR U30914 ( .A(n31778), .B(n31776), .Z(n31777) );
  XNOR U30915 ( .A(n31779), .B(n31780), .Z(n31767) );
  AND U30916 ( .A(n31781), .B(n31782), .Z(n31779) );
  XNOR U30917 ( .A(n31780), .B(n31709), .Z(n31782) );
  XOR U30918 ( .A(n31773), .B(n31774), .Z(n31709) );
  XNOR U30919 ( .A(n31783), .B(n31784), .Z(n31774) );
  ANDN U30920 ( .B(n31785), .A(n31786), .Z(n31783) );
  XOR U30921 ( .A(n31787), .B(n31788), .Z(n31785) );
  XOR U30922 ( .A(n31789), .B(n31790), .Z(n31773) );
  XNOR U30923 ( .A(n31791), .B(n31792), .Z(n31790) );
  ANDN U30924 ( .B(n31793), .A(n31794), .Z(n31791) );
  XNOR U30925 ( .A(n31795), .B(n31796), .Z(n31793) );
  IV U30926 ( .A(n31771), .Z(n31789) );
  XOR U30927 ( .A(n31797), .B(n31798), .Z(n31771) );
  ANDN U30928 ( .B(n31799), .A(n31800), .Z(n31797) );
  XOR U30929 ( .A(n31798), .B(n31801), .Z(n31799) );
  XOR U30930 ( .A(n31780), .B(n31711), .Z(n31781) );
  XOR U30931 ( .A(n31802), .B(n31803), .Z(n31711) );
  AND U30932 ( .A(n858), .B(n31804), .Z(n31802) );
  XOR U30933 ( .A(n31805), .B(n31803), .Z(n31804) );
  XNOR U30934 ( .A(n31806), .B(n31807), .Z(n31780) );
  NAND U30935 ( .A(n31808), .B(n31809), .Z(n31807) );
  XOR U30936 ( .A(n31810), .B(n31759), .Z(n31809) );
  XOR U30937 ( .A(n31800), .B(n31801), .Z(n31759) );
  XOR U30938 ( .A(n31811), .B(n31788), .Z(n31801) );
  XOR U30939 ( .A(n31812), .B(n31813), .Z(n31788) );
  ANDN U30940 ( .B(n31814), .A(n31815), .Z(n31812) );
  XOR U30941 ( .A(n31813), .B(n31816), .Z(n31814) );
  IV U30942 ( .A(n31786), .Z(n31811) );
  XOR U30943 ( .A(n31784), .B(n31817), .Z(n31786) );
  XOR U30944 ( .A(n31818), .B(n31819), .Z(n31817) );
  ANDN U30945 ( .B(n31820), .A(n31821), .Z(n31818) );
  XOR U30946 ( .A(n31822), .B(n31819), .Z(n31820) );
  IV U30947 ( .A(n31787), .Z(n31784) );
  XOR U30948 ( .A(n31823), .B(n31824), .Z(n31787) );
  ANDN U30949 ( .B(n31825), .A(n31826), .Z(n31823) );
  XOR U30950 ( .A(n31824), .B(n31827), .Z(n31825) );
  XOR U30951 ( .A(n31828), .B(n31829), .Z(n31800) );
  XNOR U30952 ( .A(n31795), .B(n31830), .Z(n31829) );
  IV U30953 ( .A(n31798), .Z(n31830) );
  XOR U30954 ( .A(n31831), .B(n31832), .Z(n31798) );
  ANDN U30955 ( .B(n31833), .A(n31834), .Z(n31831) );
  XOR U30956 ( .A(n31832), .B(n31835), .Z(n31833) );
  XNOR U30957 ( .A(n31836), .B(n31837), .Z(n31795) );
  ANDN U30958 ( .B(n31838), .A(n31839), .Z(n31836) );
  XOR U30959 ( .A(n31837), .B(n31840), .Z(n31838) );
  IV U30960 ( .A(n31794), .Z(n31828) );
  XOR U30961 ( .A(n31792), .B(n31841), .Z(n31794) );
  XOR U30962 ( .A(n31842), .B(n31843), .Z(n31841) );
  ANDN U30963 ( .B(n31844), .A(n31845), .Z(n31842) );
  XOR U30964 ( .A(n31846), .B(n31843), .Z(n31844) );
  IV U30965 ( .A(n31796), .Z(n31792) );
  XOR U30966 ( .A(n31847), .B(n31848), .Z(n31796) );
  ANDN U30967 ( .B(n31849), .A(n31850), .Z(n31847) );
  XOR U30968 ( .A(n31851), .B(n31848), .Z(n31849) );
  IV U30969 ( .A(n31806), .Z(n31810) );
  XOR U30970 ( .A(n31806), .B(n31761), .Z(n31808) );
  XOR U30971 ( .A(n31852), .B(n31853), .Z(n31761) );
  AND U30972 ( .A(n858), .B(n31854), .Z(n31852) );
  XOR U30973 ( .A(n31855), .B(n31853), .Z(n31854) );
  NANDN U30974 ( .A(n31763), .B(n31765), .Z(n31806) );
  XOR U30975 ( .A(n31856), .B(n31857), .Z(n31765) );
  AND U30976 ( .A(n858), .B(n31858), .Z(n31856) );
  XOR U30977 ( .A(n31857), .B(n31859), .Z(n31858) );
  XNOR U30978 ( .A(n31860), .B(n31861), .Z(n858) );
  AND U30979 ( .A(n31862), .B(n31863), .Z(n31860) );
  XOR U30980 ( .A(n31861), .B(n31776), .Z(n31863) );
  XNOR U30981 ( .A(n31864), .B(n31865), .Z(n31776) );
  ANDN U30982 ( .B(n31866), .A(n31867), .Z(n31864) );
  XOR U30983 ( .A(n31865), .B(n31868), .Z(n31866) );
  XNOR U30984 ( .A(n31861), .B(n31778), .Z(n31862) );
  XOR U30985 ( .A(n31869), .B(n31870), .Z(n31778) );
  AND U30986 ( .A(n862), .B(n31871), .Z(n31869) );
  XOR U30987 ( .A(n31872), .B(n31870), .Z(n31871) );
  XNOR U30988 ( .A(n31873), .B(n31874), .Z(n31861) );
  AND U30989 ( .A(n31875), .B(n31876), .Z(n31873) );
  XNOR U30990 ( .A(n31874), .B(n31803), .Z(n31876) );
  XOR U30991 ( .A(n31867), .B(n31868), .Z(n31803) );
  XNOR U30992 ( .A(n31877), .B(n31878), .Z(n31868) );
  ANDN U30993 ( .B(n31879), .A(n31880), .Z(n31877) );
  XOR U30994 ( .A(n31881), .B(n31882), .Z(n31879) );
  XOR U30995 ( .A(n31883), .B(n31884), .Z(n31867) );
  XNOR U30996 ( .A(n31885), .B(n31886), .Z(n31884) );
  ANDN U30997 ( .B(n31887), .A(n31888), .Z(n31885) );
  XNOR U30998 ( .A(n31889), .B(n31890), .Z(n31887) );
  IV U30999 ( .A(n31865), .Z(n31883) );
  XOR U31000 ( .A(n31891), .B(n31892), .Z(n31865) );
  ANDN U31001 ( .B(n31893), .A(n31894), .Z(n31891) );
  XOR U31002 ( .A(n31892), .B(n31895), .Z(n31893) );
  XOR U31003 ( .A(n31874), .B(n31805), .Z(n31875) );
  XOR U31004 ( .A(n31896), .B(n31897), .Z(n31805) );
  AND U31005 ( .A(n862), .B(n31898), .Z(n31896) );
  XOR U31006 ( .A(n31899), .B(n31897), .Z(n31898) );
  XNOR U31007 ( .A(n31900), .B(n31901), .Z(n31874) );
  NAND U31008 ( .A(n31902), .B(n31903), .Z(n31901) );
  XOR U31009 ( .A(n31904), .B(n31853), .Z(n31903) );
  XOR U31010 ( .A(n31894), .B(n31895), .Z(n31853) );
  XOR U31011 ( .A(n31905), .B(n31882), .Z(n31895) );
  XOR U31012 ( .A(n31906), .B(n31907), .Z(n31882) );
  ANDN U31013 ( .B(n31908), .A(n31909), .Z(n31906) );
  XOR U31014 ( .A(n31907), .B(n31910), .Z(n31908) );
  IV U31015 ( .A(n31880), .Z(n31905) );
  XOR U31016 ( .A(n31878), .B(n31911), .Z(n31880) );
  XOR U31017 ( .A(n31912), .B(n31913), .Z(n31911) );
  ANDN U31018 ( .B(n31914), .A(n31915), .Z(n31912) );
  XOR U31019 ( .A(n31916), .B(n31913), .Z(n31914) );
  IV U31020 ( .A(n31881), .Z(n31878) );
  XOR U31021 ( .A(n31917), .B(n31918), .Z(n31881) );
  ANDN U31022 ( .B(n31919), .A(n31920), .Z(n31917) );
  XOR U31023 ( .A(n31918), .B(n31921), .Z(n31919) );
  XOR U31024 ( .A(n31922), .B(n31923), .Z(n31894) );
  XNOR U31025 ( .A(n31889), .B(n31924), .Z(n31923) );
  IV U31026 ( .A(n31892), .Z(n31924) );
  XOR U31027 ( .A(n31925), .B(n31926), .Z(n31892) );
  ANDN U31028 ( .B(n31927), .A(n31928), .Z(n31925) );
  XOR U31029 ( .A(n31926), .B(n31929), .Z(n31927) );
  XNOR U31030 ( .A(n31930), .B(n31931), .Z(n31889) );
  ANDN U31031 ( .B(n31932), .A(n31933), .Z(n31930) );
  XOR U31032 ( .A(n31931), .B(n31934), .Z(n31932) );
  IV U31033 ( .A(n31888), .Z(n31922) );
  XOR U31034 ( .A(n31886), .B(n31935), .Z(n31888) );
  XOR U31035 ( .A(n31936), .B(n31937), .Z(n31935) );
  ANDN U31036 ( .B(n31938), .A(n31939), .Z(n31936) );
  XOR U31037 ( .A(n31940), .B(n31937), .Z(n31938) );
  IV U31038 ( .A(n31890), .Z(n31886) );
  XOR U31039 ( .A(n31941), .B(n31942), .Z(n31890) );
  ANDN U31040 ( .B(n31943), .A(n31944), .Z(n31941) );
  XOR U31041 ( .A(n31945), .B(n31942), .Z(n31943) );
  IV U31042 ( .A(n31900), .Z(n31904) );
  XOR U31043 ( .A(n31900), .B(n31855), .Z(n31902) );
  XOR U31044 ( .A(n31946), .B(n31947), .Z(n31855) );
  AND U31045 ( .A(n862), .B(n31948), .Z(n31946) );
  XOR U31046 ( .A(n31949), .B(n31947), .Z(n31948) );
  NANDN U31047 ( .A(n31857), .B(n31859), .Z(n31900) );
  XOR U31048 ( .A(n31950), .B(n31951), .Z(n31859) );
  AND U31049 ( .A(n862), .B(n31952), .Z(n31950) );
  XOR U31050 ( .A(n31951), .B(n31953), .Z(n31952) );
  XNOR U31051 ( .A(n31954), .B(n31955), .Z(n862) );
  AND U31052 ( .A(n31956), .B(n31957), .Z(n31954) );
  XOR U31053 ( .A(n31955), .B(n31870), .Z(n31957) );
  XNOR U31054 ( .A(n31958), .B(n31959), .Z(n31870) );
  ANDN U31055 ( .B(n31960), .A(n31961), .Z(n31958) );
  XOR U31056 ( .A(n31959), .B(n31962), .Z(n31960) );
  XNOR U31057 ( .A(n31955), .B(n31872), .Z(n31956) );
  XOR U31058 ( .A(n31963), .B(n31964), .Z(n31872) );
  AND U31059 ( .A(n866), .B(n31965), .Z(n31963) );
  XOR U31060 ( .A(n31966), .B(n31964), .Z(n31965) );
  XNOR U31061 ( .A(n31967), .B(n31968), .Z(n31955) );
  AND U31062 ( .A(n31969), .B(n31970), .Z(n31967) );
  XNOR U31063 ( .A(n31968), .B(n31897), .Z(n31970) );
  XOR U31064 ( .A(n31961), .B(n31962), .Z(n31897) );
  XNOR U31065 ( .A(n31971), .B(n31972), .Z(n31962) );
  ANDN U31066 ( .B(n31973), .A(n31974), .Z(n31971) );
  XOR U31067 ( .A(n31975), .B(n31976), .Z(n31973) );
  XOR U31068 ( .A(n31977), .B(n31978), .Z(n31961) );
  XNOR U31069 ( .A(n31979), .B(n31980), .Z(n31978) );
  ANDN U31070 ( .B(n31981), .A(n31982), .Z(n31979) );
  XNOR U31071 ( .A(n31983), .B(n31984), .Z(n31981) );
  IV U31072 ( .A(n31959), .Z(n31977) );
  XOR U31073 ( .A(n31985), .B(n31986), .Z(n31959) );
  ANDN U31074 ( .B(n31987), .A(n31988), .Z(n31985) );
  XOR U31075 ( .A(n31986), .B(n31989), .Z(n31987) );
  XOR U31076 ( .A(n31968), .B(n31899), .Z(n31969) );
  XOR U31077 ( .A(n31990), .B(n31991), .Z(n31899) );
  AND U31078 ( .A(n866), .B(n31992), .Z(n31990) );
  XOR U31079 ( .A(n31993), .B(n31991), .Z(n31992) );
  XNOR U31080 ( .A(n31994), .B(n31995), .Z(n31968) );
  NAND U31081 ( .A(n31996), .B(n31997), .Z(n31995) );
  XOR U31082 ( .A(n31998), .B(n31947), .Z(n31997) );
  XOR U31083 ( .A(n31988), .B(n31989), .Z(n31947) );
  XOR U31084 ( .A(n31999), .B(n31976), .Z(n31989) );
  XOR U31085 ( .A(n32000), .B(n32001), .Z(n31976) );
  ANDN U31086 ( .B(n32002), .A(n32003), .Z(n32000) );
  XOR U31087 ( .A(n32001), .B(n32004), .Z(n32002) );
  IV U31088 ( .A(n31974), .Z(n31999) );
  XOR U31089 ( .A(n31972), .B(n32005), .Z(n31974) );
  XOR U31090 ( .A(n32006), .B(n32007), .Z(n32005) );
  ANDN U31091 ( .B(n32008), .A(n32009), .Z(n32006) );
  XOR U31092 ( .A(n32010), .B(n32007), .Z(n32008) );
  IV U31093 ( .A(n31975), .Z(n31972) );
  XOR U31094 ( .A(n32011), .B(n32012), .Z(n31975) );
  ANDN U31095 ( .B(n32013), .A(n32014), .Z(n32011) );
  XOR U31096 ( .A(n32012), .B(n32015), .Z(n32013) );
  XOR U31097 ( .A(n32016), .B(n32017), .Z(n31988) );
  XNOR U31098 ( .A(n31983), .B(n32018), .Z(n32017) );
  IV U31099 ( .A(n31986), .Z(n32018) );
  XOR U31100 ( .A(n32019), .B(n32020), .Z(n31986) );
  ANDN U31101 ( .B(n32021), .A(n32022), .Z(n32019) );
  XOR U31102 ( .A(n32020), .B(n32023), .Z(n32021) );
  XNOR U31103 ( .A(n32024), .B(n32025), .Z(n31983) );
  ANDN U31104 ( .B(n32026), .A(n32027), .Z(n32024) );
  XOR U31105 ( .A(n32025), .B(n32028), .Z(n32026) );
  IV U31106 ( .A(n31982), .Z(n32016) );
  XOR U31107 ( .A(n31980), .B(n32029), .Z(n31982) );
  XOR U31108 ( .A(n32030), .B(n32031), .Z(n32029) );
  ANDN U31109 ( .B(n32032), .A(n32033), .Z(n32030) );
  XOR U31110 ( .A(n32034), .B(n32031), .Z(n32032) );
  IV U31111 ( .A(n31984), .Z(n31980) );
  XOR U31112 ( .A(n32035), .B(n32036), .Z(n31984) );
  ANDN U31113 ( .B(n32037), .A(n32038), .Z(n32035) );
  XOR U31114 ( .A(n32039), .B(n32036), .Z(n32037) );
  IV U31115 ( .A(n31994), .Z(n31998) );
  XOR U31116 ( .A(n31994), .B(n31949), .Z(n31996) );
  XOR U31117 ( .A(n32040), .B(n32041), .Z(n31949) );
  AND U31118 ( .A(n866), .B(n32042), .Z(n32040) );
  XOR U31119 ( .A(n32043), .B(n32041), .Z(n32042) );
  NANDN U31120 ( .A(n31951), .B(n31953), .Z(n31994) );
  XOR U31121 ( .A(n32044), .B(n32045), .Z(n31953) );
  AND U31122 ( .A(n866), .B(n32046), .Z(n32044) );
  XOR U31123 ( .A(n32045), .B(n32047), .Z(n32046) );
  XNOR U31124 ( .A(n32048), .B(n32049), .Z(n866) );
  AND U31125 ( .A(n32050), .B(n32051), .Z(n32048) );
  XOR U31126 ( .A(n32049), .B(n31964), .Z(n32051) );
  XNOR U31127 ( .A(n32052), .B(n32053), .Z(n31964) );
  ANDN U31128 ( .B(n32054), .A(n32055), .Z(n32052) );
  XOR U31129 ( .A(n32053), .B(n32056), .Z(n32054) );
  XNOR U31130 ( .A(n32049), .B(n31966), .Z(n32050) );
  XOR U31131 ( .A(n32057), .B(n32058), .Z(n31966) );
  AND U31132 ( .A(n870), .B(n32059), .Z(n32057) );
  XOR U31133 ( .A(n32060), .B(n32058), .Z(n32059) );
  XNOR U31134 ( .A(n32061), .B(n32062), .Z(n32049) );
  AND U31135 ( .A(n32063), .B(n32064), .Z(n32061) );
  XNOR U31136 ( .A(n32062), .B(n31991), .Z(n32064) );
  XOR U31137 ( .A(n32055), .B(n32056), .Z(n31991) );
  XNOR U31138 ( .A(n32065), .B(n32066), .Z(n32056) );
  ANDN U31139 ( .B(n32067), .A(n32068), .Z(n32065) );
  XOR U31140 ( .A(n32069), .B(n32070), .Z(n32067) );
  XOR U31141 ( .A(n32071), .B(n32072), .Z(n32055) );
  XNOR U31142 ( .A(n32073), .B(n32074), .Z(n32072) );
  ANDN U31143 ( .B(n32075), .A(n32076), .Z(n32073) );
  XNOR U31144 ( .A(n32077), .B(n32078), .Z(n32075) );
  IV U31145 ( .A(n32053), .Z(n32071) );
  XOR U31146 ( .A(n32079), .B(n32080), .Z(n32053) );
  ANDN U31147 ( .B(n32081), .A(n32082), .Z(n32079) );
  XOR U31148 ( .A(n32080), .B(n32083), .Z(n32081) );
  XOR U31149 ( .A(n32062), .B(n31993), .Z(n32063) );
  XOR U31150 ( .A(n32084), .B(n32085), .Z(n31993) );
  AND U31151 ( .A(n870), .B(n32086), .Z(n32084) );
  XOR U31152 ( .A(n32087), .B(n32085), .Z(n32086) );
  XNOR U31153 ( .A(n32088), .B(n32089), .Z(n32062) );
  NAND U31154 ( .A(n32090), .B(n32091), .Z(n32089) );
  XOR U31155 ( .A(n32092), .B(n32041), .Z(n32091) );
  XOR U31156 ( .A(n32082), .B(n32083), .Z(n32041) );
  XOR U31157 ( .A(n32093), .B(n32070), .Z(n32083) );
  XOR U31158 ( .A(n32094), .B(n32095), .Z(n32070) );
  ANDN U31159 ( .B(n32096), .A(n32097), .Z(n32094) );
  XOR U31160 ( .A(n32095), .B(n32098), .Z(n32096) );
  IV U31161 ( .A(n32068), .Z(n32093) );
  XOR U31162 ( .A(n32066), .B(n32099), .Z(n32068) );
  XOR U31163 ( .A(n32100), .B(n32101), .Z(n32099) );
  ANDN U31164 ( .B(n32102), .A(n32103), .Z(n32100) );
  XOR U31165 ( .A(n32104), .B(n32101), .Z(n32102) );
  IV U31166 ( .A(n32069), .Z(n32066) );
  XOR U31167 ( .A(n32105), .B(n32106), .Z(n32069) );
  ANDN U31168 ( .B(n32107), .A(n32108), .Z(n32105) );
  XOR U31169 ( .A(n32106), .B(n32109), .Z(n32107) );
  XOR U31170 ( .A(n32110), .B(n32111), .Z(n32082) );
  XNOR U31171 ( .A(n32077), .B(n32112), .Z(n32111) );
  IV U31172 ( .A(n32080), .Z(n32112) );
  XOR U31173 ( .A(n32113), .B(n32114), .Z(n32080) );
  ANDN U31174 ( .B(n32115), .A(n32116), .Z(n32113) );
  XOR U31175 ( .A(n32114), .B(n32117), .Z(n32115) );
  XNOR U31176 ( .A(n32118), .B(n32119), .Z(n32077) );
  ANDN U31177 ( .B(n32120), .A(n32121), .Z(n32118) );
  XOR U31178 ( .A(n32119), .B(n32122), .Z(n32120) );
  IV U31179 ( .A(n32076), .Z(n32110) );
  XOR U31180 ( .A(n32074), .B(n32123), .Z(n32076) );
  XOR U31181 ( .A(n32124), .B(n32125), .Z(n32123) );
  ANDN U31182 ( .B(n32126), .A(n32127), .Z(n32124) );
  XOR U31183 ( .A(n32128), .B(n32125), .Z(n32126) );
  IV U31184 ( .A(n32078), .Z(n32074) );
  XOR U31185 ( .A(n32129), .B(n32130), .Z(n32078) );
  ANDN U31186 ( .B(n32131), .A(n32132), .Z(n32129) );
  XOR U31187 ( .A(n32133), .B(n32130), .Z(n32131) );
  IV U31188 ( .A(n32088), .Z(n32092) );
  XOR U31189 ( .A(n32088), .B(n32043), .Z(n32090) );
  XOR U31190 ( .A(n32134), .B(n32135), .Z(n32043) );
  AND U31191 ( .A(n870), .B(n32136), .Z(n32134) );
  XOR U31192 ( .A(n32137), .B(n32135), .Z(n32136) );
  NANDN U31193 ( .A(n32045), .B(n32047), .Z(n32088) );
  XOR U31194 ( .A(n32138), .B(n32139), .Z(n32047) );
  AND U31195 ( .A(n870), .B(n32140), .Z(n32138) );
  XOR U31196 ( .A(n32139), .B(n32141), .Z(n32140) );
  XNOR U31197 ( .A(n32142), .B(n32143), .Z(n870) );
  AND U31198 ( .A(n32144), .B(n32145), .Z(n32142) );
  XOR U31199 ( .A(n32143), .B(n32058), .Z(n32145) );
  XNOR U31200 ( .A(n32146), .B(n32147), .Z(n32058) );
  ANDN U31201 ( .B(n32148), .A(n32149), .Z(n32146) );
  XOR U31202 ( .A(n32147), .B(n32150), .Z(n32148) );
  XNOR U31203 ( .A(n32143), .B(n32060), .Z(n32144) );
  XOR U31204 ( .A(n32151), .B(n32152), .Z(n32060) );
  AND U31205 ( .A(n874), .B(n32153), .Z(n32151) );
  XOR U31206 ( .A(n32154), .B(n32152), .Z(n32153) );
  XNOR U31207 ( .A(n32155), .B(n32156), .Z(n32143) );
  AND U31208 ( .A(n32157), .B(n32158), .Z(n32155) );
  XNOR U31209 ( .A(n32156), .B(n32085), .Z(n32158) );
  XOR U31210 ( .A(n32149), .B(n32150), .Z(n32085) );
  XNOR U31211 ( .A(n32159), .B(n32160), .Z(n32150) );
  ANDN U31212 ( .B(n32161), .A(n32162), .Z(n32159) );
  XOR U31213 ( .A(n32163), .B(n32164), .Z(n32161) );
  XOR U31214 ( .A(n32165), .B(n32166), .Z(n32149) );
  XNOR U31215 ( .A(n32167), .B(n32168), .Z(n32166) );
  ANDN U31216 ( .B(n32169), .A(n32170), .Z(n32167) );
  XNOR U31217 ( .A(n32171), .B(n32172), .Z(n32169) );
  IV U31218 ( .A(n32147), .Z(n32165) );
  XOR U31219 ( .A(n32173), .B(n32174), .Z(n32147) );
  ANDN U31220 ( .B(n32175), .A(n32176), .Z(n32173) );
  XOR U31221 ( .A(n32174), .B(n32177), .Z(n32175) );
  XOR U31222 ( .A(n32156), .B(n32087), .Z(n32157) );
  XOR U31223 ( .A(n32178), .B(n32179), .Z(n32087) );
  AND U31224 ( .A(n874), .B(n32180), .Z(n32178) );
  XOR U31225 ( .A(n32181), .B(n32179), .Z(n32180) );
  XNOR U31226 ( .A(n32182), .B(n32183), .Z(n32156) );
  NAND U31227 ( .A(n32184), .B(n32185), .Z(n32183) );
  XOR U31228 ( .A(n32186), .B(n32135), .Z(n32185) );
  XOR U31229 ( .A(n32176), .B(n32177), .Z(n32135) );
  XOR U31230 ( .A(n32187), .B(n32164), .Z(n32177) );
  XOR U31231 ( .A(n32188), .B(n32189), .Z(n32164) );
  ANDN U31232 ( .B(n32190), .A(n32191), .Z(n32188) );
  XOR U31233 ( .A(n32189), .B(n32192), .Z(n32190) );
  IV U31234 ( .A(n32162), .Z(n32187) );
  XOR U31235 ( .A(n32160), .B(n32193), .Z(n32162) );
  XOR U31236 ( .A(n32194), .B(n32195), .Z(n32193) );
  ANDN U31237 ( .B(n32196), .A(n32197), .Z(n32194) );
  XOR U31238 ( .A(n32198), .B(n32195), .Z(n32196) );
  IV U31239 ( .A(n32163), .Z(n32160) );
  XOR U31240 ( .A(n32199), .B(n32200), .Z(n32163) );
  ANDN U31241 ( .B(n32201), .A(n32202), .Z(n32199) );
  XOR U31242 ( .A(n32200), .B(n32203), .Z(n32201) );
  XOR U31243 ( .A(n32204), .B(n32205), .Z(n32176) );
  XNOR U31244 ( .A(n32171), .B(n32206), .Z(n32205) );
  IV U31245 ( .A(n32174), .Z(n32206) );
  XOR U31246 ( .A(n32207), .B(n32208), .Z(n32174) );
  ANDN U31247 ( .B(n32209), .A(n32210), .Z(n32207) );
  XOR U31248 ( .A(n32208), .B(n32211), .Z(n32209) );
  XNOR U31249 ( .A(n32212), .B(n32213), .Z(n32171) );
  ANDN U31250 ( .B(n32214), .A(n32215), .Z(n32212) );
  XOR U31251 ( .A(n32213), .B(n32216), .Z(n32214) );
  IV U31252 ( .A(n32170), .Z(n32204) );
  XOR U31253 ( .A(n32168), .B(n32217), .Z(n32170) );
  XOR U31254 ( .A(n32218), .B(n32219), .Z(n32217) );
  ANDN U31255 ( .B(n32220), .A(n32221), .Z(n32218) );
  XOR U31256 ( .A(n32222), .B(n32219), .Z(n32220) );
  IV U31257 ( .A(n32172), .Z(n32168) );
  XOR U31258 ( .A(n32223), .B(n32224), .Z(n32172) );
  ANDN U31259 ( .B(n32225), .A(n32226), .Z(n32223) );
  XOR U31260 ( .A(n32227), .B(n32224), .Z(n32225) );
  IV U31261 ( .A(n32182), .Z(n32186) );
  XOR U31262 ( .A(n32182), .B(n32137), .Z(n32184) );
  XOR U31263 ( .A(n32228), .B(n32229), .Z(n32137) );
  AND U31264 ( .A(n874), .B(n32230), .Z(n32228) );
  XOR U31265 ( .A(n32231), .B(n32229), .Z(n32230) );
  NANDN U31266 ( .A(n32139), .B(n32141), .Z(n32182) );
  XOR U31267 ( .A(n32232), .B(n32233), .Z(n32141) );
  AND U31268 ( .A(n874), .B(n32234), .Z(n32232) );
  XOR U31269 ( .A(n32233), .B(n32235), .Z(n32234) );
  XNOR U31270 ( .A(n32236), .B(n32237), .Z(n874) );
  AND U31271 ( .A(n32238), .B(n32239), .Z(n32236) );
  XOR U31272 ( .A(n32237), .B(n32152), .Z(n32239) );
  XNOR U31273 ( .A(n32240), .B(n32241), .Z(n32152) );
  ANDN U31274 ( .B(n32242), .A(n32243), .Z(n32240) );
  XOR U31275 ( .A(n32241), .B(n32244), .Z(n32242) );
  XNOR U31276 ( .A(n32237), .B(n32154), .Z(n32238) );
  XOR U31277 ( .A(n32245), .B(n32246), .Z(n32154) );
  AND U31278 ( .A(n878), .B(n32247), .Z(n32245) );
  XOR U31279 ( .A(n32248), .B(n32246), .Z(n32247) );
  XNOR U31280 ( .A(n32249), .B(n32250), .Z(n32237) );
  AND U31281 ( .A(n32251), .B(n32252), .Z(n32249) );
  XNOR U31282 ( .A(n32250), .B(n32179), .Z(n32252) );
  XOR U31283 ( .A(n32243), .B(n32244), .Z(n32179) );
  XNOR U31284 ( .A(n32253), .B(n32254), .Z(n32244) );
  ANDN U31285 ( .B(n32255), .A(n32256), .Z(n32253) );
  XOR U31286 ( .A(n32257), .B(n32258), .Z(n32255) );
  XOR U31287 ( .A(n32259), .B(n32260), .Z(n32243) );
  XNOR U31288 ( .A(n32261), .B(n32262), .Z(n32260) );
  ANDN U31289 ( .B(n32263), .A(n32264), .Z(n32261) );
  XNOR U31290 ( .A(n32265), .B(n32266), .Z(n32263) );
  IV U31291 ( .A(n32241), .Z(n32259) );
  XOR U31292 ( .A(n32267), .B(n32268), .Z(n32241) );
  ANDN U31293 ( .B(n32269), .A(n32270), .Z(n32267) );
  XOR U31294 ( .A(n32268), .B(n32271), .Z(n32269) );
  XOR U31295 ( .A(n32250), .B(n32181), .Z(n32251) );
  XOR U31296 ( .A(n32272), .B(n32273), .Z(n32181) );
  AND U31297 ( .A(n878), .B(n32274), .Z(n32272) );
  XOR U31298 ( .A(n32275), .B(n32273), .Z(n32274) );
  XNOR U31299 ( .A(n32276), .B(n32277), .Z(n32250) );
  NAND U31300 ( .A(n32278), .B(n32279), .Z(n32277) );
  XOR U31301 ( .A(n32280), .B(n32229), .Z(n32279) );
  XOR U31302 ( .A(n32270), .B(n32271), .Z(n32229) );
  XOR U31303 ( .A(n32281), .B(n32258), .Z(n32271) );
  XOR U31304 ( .A(n32282), .B(n32283), .Z(n32258) );
  ANDN U31305 ( .B(n32284), .A(n32285), .Z(n32282) );
  XOR U31306 ( .A(n32283), .B(n32286), .Z(n32284) );
  IV U31307 ( .A(n32256), .Z(n32281) );
  XOR U31308 ( .A(n32254), .B(n32287), .Z(n32256) );
  XOR U31309 ( .A(n32288), .B(n32289), .Z(n32287) );
  ANDN U31310 ( .B(n32290), .A(n32291), .Z(n32288) );
  XOR U31311 ( .A(n32292), .B(n32289), .Z(n32290) );
  IV U31312 ( .A(n32257), .Z(n32254) );
  XOR U31313 ( .A(n32293), .B(n32294), .Z(n32257) );
  ANDN U31314 ( .B(n32295), .A(n32296), .Z(n32293) );
  XOR U31315 ( .A(n32294), .B(n32297), .Z(n32295) );
  XOR U31316 ( .A(n32298), .B(n32299), .Z(n32270) );
  XNOR U31317 ( .A(n32265), .B(n32300), .Z(n32299) );
  IV U31318 ( .A(n32268), .Z(n32300) );
  XOR U31319 ( .A(n32301), .B(n32302), .Z(n32268) );
  ANDN U31320 ( .B(n32303), .A(n32304), .Z(n32301) );
  XOR U31321 ( .A(n32302), .B(n32305), .Z(n32303) );
  XNOR U31322 ( .A(n32306), .B(n32307), .Z(n32265) );
  ANDN U31323 ( .B(n32308), .A(n32309), .Z(n32306) );
  XOR U31324 ( .A(n32307), .B(n32310), .Z(n32308) );
  IV U31325 ( .A(n32264), .Z(n32298) );
  XOR U31326 ( .A(n32262), .B(n32311), .Z(n32264) );
  XOR U31327 ( .A(n32312), .B(n32313), .Z(n32311) );
  ANDN U31328 ( .B(n32314), .A(n32315), .Z(n32312) );
  XOR U31329 ( .A(n32316), .B(n32313), .Z(n32314) );
  IV U31330 ( .A(n32266), .Z(n32262) );
  XOR U31331 ( .A(n32317), .B(n32318), .Z(n32266) );
  ANDN U31332 ( .B(n32319), .A(n32320), .Z(n32317) );
  XOR U31333 ( .A(n32321), .B(n32318), .Z(n32319) );
  IV U31334 ( .A(n32276), .Z(n32280) );
  XOR U31335 ( .A(n32276), .B(n32231), .Z(n32278) );
  XOR U31336 ( .A(n32322), .B(n32323), .Z(n32231) );
  AND U31337 ( .A(n878), .B(n32324), .Z(n32322) );
  XOR U31338 ( .A(n32325), .B(n32323), .Z(n32324) );
  NANDN U31339 ( .A(n32233), .B(n32235), .Z(n32276) );
  XOR U31340 ( .A(n32326), .B(n32327), .Z(n32235) );
  AND U31341 ( .A(n878), .B(n32328), .Z(n32326) );
  XOR U31342 ( .A(n32327), .B(n32329), .Z(n32328) );
  XNOR U31343 ( .A(n32330), .B(n32331), .Z(n878) );
  AND U31344 ( .A(n32332), .B(n32333), .Z(n32330) );
  XOR U31345 ( .A(n32331), .B(n32246), .Z(n32333) );
  XNOR U31346 ( .A(n32334), .B(n32335), .Z(n32246) );
  ANDN U31347 ( .B(n32336), .A(n32337), .Z(n32334) );
  XOR U31348 ( .A(n32335), .B(n32338), .Z(n32336) );
  XNOR U31349 ( .A(n32331), .B(n32248), .Z(n32332) );
  XOR U31350 ( .A(n32339), .B(n32340), .Z(n32248) );
  AND U31351 ( .A(n882), .B(n32341), .Z(n32339) );
  XOR U31352 ( .A(n32342), .B(n32340), .Z(n32341) );
  XNOR U31353 ( .A(n32343), .B(n32344), .Z(n32331) );
  AND U31354 ( .A(n32345), .B(n32346), .Z(n32343) );
  XNOR U31355 ( .A(n32344), .B(n32273), .Z(n32346) );
  XOR U31356 ( .A(n32337), .B(n32338), .Z(n32273) );
  XNOR U31357 ( .A(n32347), .B(n32348), .Z(n32338) );
  ANDN U31358 ( .B(n32349), .A(n32350), .Z(n32347) );
  XOR U31359 ( .A(n32351), .B(n32352), .Z(n32349) );
  XOR U31360 ( .A(n32353), .B(n32354), .Z(n32337) );
  XNOR U31361 ( .A(n32355), .B(n32356), .Z(n32354) );
  ANDN U31362 ( .B(n32357), .A(n32358), .Z(n32355) );
  XNOR U31363 ( .A(n32359), .B(n32360), .Z(n32357) );
  IV U31364 ( .A(n32335), .Z(n32353) );
  XOR U31365 ( .A(n32361), .B(n32362), .Z(n32335) );
  ANDN U31366 ( .B(n32363), .A(n32364), .Z(n32361) );
  XOR U31367 ( .A(n32362), .B(n32365), .Z(n32363) );
  XOR U31368 ( .A(n32344), .B(n32275), .Z(n32345) );
  XOR U31369 ( .A(n32366), .B(n32367), .Z(n32275) );
  AND U31370 ( .A(n882), .B(n32368), .Z(n32366) );
  XOR U31371 ( .A(n32369), .B(n32367), .Z(n32368) );
  XNOR U31372 ( .A(n32370), .B(n32371), .Z(n32344) );
  NAND U31373 ( .A(n32372), .B(n32373), .Z(n32371) );
  XOR U31374 ( .A(n32374), .B(n32323), .Z(n32373) );
  XOR U31375 ( .A(n32364), .B(n32365), .Z(n32323) );
  XOR U31376 ( .A(n32375), .B(n32352), .Z(n32365) );
  XOR U31377 ( .A(n32376), .B(n32377), .Z(n32352) );
  ANDN U31378 ( .B(n32378), .A(n32379), .Z(n32376) );
  XOR U31379 ( .A(n32377), .B(n32380), .Z(n32378) );
  IV U31380 ( .A(n32350), .Z(n32375) );
  XOR U31381 ( .A(n32348), .B(n32381), .Z(n32350) );
  XOR U31382 ( .A(n32382), .B(n32383), .Z(n32381) );
  ANDN U31383 ( .B(n32384), .A(n32385), .Z(n32382) );
  XOR U31384 ( .A(n32386), .B(n32383), .Z(n32384) );
  IV U31385 ( .A(n32351), .Z(n32348) );
  XOR U31386 ( .A(n32387), .B(n32388), .Z(n32351) );
  ANDN U31387 ( .B(n32389), .A(n32390), .Z(n32387) );
  XOR U31388 ( .A(n32388), .B(n32391), .Z(n32389) );
  XOR U31389 ( .A(n32392), .B(n32393), .Z(n32364) );
  XNOR U31390 ( .A(n32359), .B(n32394), .Z(n32393) );
  IV U31391 ( .A(n32362), .Z(n32394) );
  XOR U31392 ( .A(n32395), .B(n32396), .Z(n32362) );
  ANDN U31393 ( .B(n32397), .A(n32398), .Z(n32395) );
  XOR U31394 ( .A(n32396), .B(n32399), .Z(n32397) );
  XNOR U31395 ( .A(n32400), .B(n32401), .Z(n32359) );
  ANDN U31396 ( .B(n32402), .A(n32403), .Z(n32400) );
  XOR U31397 ( .A(n32401), .B(n32404), .Z(n32402) );
  IV U31398 ( .A(n32358), .Z(n32392) );
  XOR U31399 ( .A(n32356), .B(n32405), .Z(n32358) );
  XOR U31400 ( .A(n32406), .B(n32407), .Z(n32405) );
  ANDN U31401 ( .B(n32408), .A(n32409), .Z(n32406) );
  XOR U31402 ( .A(n32410), .B(n32407), .Z(n32408) );
  IV U31403 ( .A(n32360), .Z(n32356) );
  XOR U31404 ( .A(n32411), .B(n32412), .Z(n32360) );
  ANDN U31405 ( .B(n32413), .A(n32414), .Z(n32411) );
  XOR U31406 ( .A(n32415), .B(n32412), .Z(n32413) );
  IV U31407 ( .A(n32370), .Z(n32374) );
  XOR U31408 ( .A(n32370), .B(n32325), .Z(n32372) );
  XOR U31409 ( .A(n32416), .B(n32417), .Z(n32325) );
  AND U31410 ( .A(n882), .B(n32418), .Z(n32416) );
  XOR U31411 ( .A(n32419), .B(n32417), .Z(n32418) );
  NANDN U31412 ( .A(n32327), .B(n32329), .Z(n32370) );
  XOR U31413 ( .A(n32420), .B(n32421), .Z(n32329) );
  AND U31414 ( .A(n882), .B(n32422), .Z(n32420) );
  XOR U31415 ( .A(n32421), .B(n32423), .Z(n32422) );
  XNOR U31416 ( .A(n32424), .B(n32425), .Z(n882) );
  AND U31417 ( .A(n32426), .B(n32427), .Z(n32424) );
  XOR U31418 ( .A(n32425), .B(n32340), .Z(n32427) );
  XNOR U31419 ( .A(n32428), .B(n32429), .Z(n32340) );
  ANDN U31420 ( .B(n32430), .A(n32431), .Z(n32428) );
  XOR U31421 ( .A(n32429), .B(n32432), .Z(n32430) );
  XNOR U31422 ( .A(n32425), .B(n32342), .Z(n32426) );
  XOR U31423 ( .A(n32433), .B(n32434), .Z(n32342) );
  AND U31424 ( .A(n886), .B(n32435), .Z(n32433) );
  XOR U31425 ( .A(n32436), .B(n32434), .Z(n32435) );
  XNOR U31426 ( .A(n32437), .B(n32438), .Z(n32425) );
  AND U31427 ( .A(n32439), .B(n32440), .Z(n32437) );
  XNOR U31428 ( .A(n32438), .B(n32367), .Z(n32440) );
  XOR U31429 ( .A(n32431), .B(n32432), .Z(n32367) );
  XNOR U31430 ( .A(n32441), .B(n32442), .Z(n32432) );
  ANDN U31431 ( .B(n32443), .A(n32444), .Z(n32441) );
  XOR U31432 ( .A(n32445), .B(n32446), .Z(n32443) );
  XOR U31433 ( .A(n32447), .B(n32448), .Z(n32431) );
  XNOR U31434 ( .A(n32449), .B(n32450), .Z(n32448) );
  ANDN U31435 ( .B(n32451), .A(n32452), .Z(n32449) );
  XNOR U31436 ( .A(n32453), .B(n32454), .Z(n32451) );
  IV U31437 ( .A(n32429), .Z(n32447) );
  XOR U31438 ( .A(n32455), .B(n32456), .Z(n32429) );
  ANDN U31439 ( .B(n32457), .A(n32458), .Z(n32455) );
  XOR U31440 ( .A(n32456), .B(n32459), .Z(n32457) );
  XOR U31441 ( .A(n32438), .B(n32369), .Z(n32439) );
  XOR U31442 ( .A(n32460), .B(n32461), .Z(n32369) );
  AND U31443 ( .A(n886), .B(n32462), .Z(n32460) );
  XOR U31444 ( .A(n32463), .B(n32461), .Z(n32462) );
  XNOR U31445 ( .A(n32464), .B(n32465), .Z(n32438) );
  NAND U31446 ( .A(n32466), .B(n32467), .Z(n32465) );
  XOR U31447 ( .A(n32468), .B(n32417), .Z(n32467) );
  XOR U31448 ( .A(n32458), .B(n32459), .Z(n32417) );
  XOR U31449 ( .A(n32469), .B(n32446), .Z(n32459) );
  XOR U31450 ( .A(n32470), .B(n32471), .Z(n32446) );
  ANDN U31451 ( .B(n32472), .A(n32473), .Z(n32470) );
  XOR U31452 ( .A(n32471), .B(n32474), .Z(n32472) );
  IV U31453 ( .A(n32444), .Z(n32469) );
  XOR U31454 ( .A(n32442), .B(n32475), .Z(n32444) );
  XOR U31455 ( .A(n32476), .B(n32477), .Z(n32475) );
  ANDN U31456 ( .B(n32478), .A(n32479), .Z(n32476) );
  XOR U31457 ( .A(n32480), .B(n32477), .Z(n32478) );
  IV U31458 ( .A(n32445), .Z(n32442) );
  XOR U31459 ( .A(n32481), .B(n32482), .Z(n32445) );
  ANDN U31460 ( .B(n32483), .A(n32484), .Z(n32481) );
  XOR U31461 ( .A(n32482), .B(n32485), .Z(n32483) );
  XOR U31462 ( .A(n32486), .B(n32487), .Z(n32458) );
  XNOR U31463 ( .A(n32453), .B(n32488), .Z(n32487) );
  IV U31464 ( .A(n32456), .Z(n32488) );
  XOR U31465 ( .A(n32489), .B(n32490), .Z(n32456) );
  ANDN U31466 ( .B(n32491), .A(n32492), .Z(n32489) );
  XOR U31467 ( .A(n32490), .B(n32493), .Z(n32491) );
  XNOR U31468 ( .A(n32494), .B(n32495), .Z(n32453) );
  ANDN U31469 ( .B(n32496), .A(n32497), .Z(n32494) );
  XOR U31470 ( .A(n32495), .B(n32498), .Z(n32496) );
  IV U31471 ( .A(n32452), .Z(n32486) );
  XOR U31472 ( .A(n32450), .B(n32499), .Z(n32452) );
  XOR U31473 ( .A(n32500), .B(n32501), .Z(n32499) );
  ANDN U31474 ( .B(n32502), .A(n32503), .Z(n32500) );
  XOR U31475 ( .A(n32504), .B(n32501), .Z(n32502) );
  IV U31476 ( .A(n32454), .Z(n32450) );
  XOR U31477 ( .A(n32505), .B(n32506), .Z(n32454) );
  ANDN U31478 ( .B(n32507), .A(n32508), .Z(n32505) );
  XOR U31479 ( .A(n32509), .B(n32506), .Z(n32507) );
  IV U31480 ( .A(n32464), .Z(n32468) );
  XOR U31481 ( .A(n32464), .B(n32419), .Z(n32466) );
  XOR U31482 ( .A(n32510), .B(n32511), .Z(n32419) );
  AND U31483 ( .A(n886), .B(n32512), .Z(n32510) );
  XOR U31484 ( .A(n32513), .B(n32511), .Z(n32512) );
  NANDN U31485 ( .A(n32421), .B(n32423), .Z(n32464) );
  XOR U31486 ( .A(n32514), .B(n32515), .Z(n32423) );
  AND U31487 ( .A(n886), .B(n32516), .Z(n32514) );
  XOR U31488 ( .A(n32515), .B(n32517), .Z(n32516) );
  XNOR U31489 ( .A(n32518), .B(n32519), .Z(n886) );
  AND U31490 ( .A(n32520), .B(n32521), .Z(n32518) );
  XOR U31491 ( .A(n32519), .B(n32434), .Z(n32521) );
  XNOR U31492 ( .A(n32522), .B(n32523), .Z(n32434) );
  ANDN U31493 ( .B(n32524), .A(n32525), .Z(n32522) );
  XOR U31494 ( .A(n32523), .B(n32526), .Z(n32524) );
  XNOR U31495 ( .A(n32519), .B(n32436), .Z(n32520) );
  XOR U31496 ( .A(n32527), .B(n32528), .Z(n32436) );
  AND U31497 ( .A(n890), .B(n32529), .Z(n32527) );
  XOR U31498 ( .A(n32530), .B(n32528), .Z(n32529) );
  XNOR U31499 ( .A(n32531), .B(n32532), .Z(n32519) );
  AND U31500 ( .A(n32533), .B(n32534), .Z(n32531) );
  XNOR U31501 ( .A(n32532), .B(n32461), .Z(n32534) );
  XOR U31502 ( .A(n32525), .B(n32526), .Z(n32461) );
  XNOR U31503 ( .A(n32535), .B(n32536), .Z(n32526) );
  ANDN U31504 ( .B(n32537), .A(n32538), .Z(n32535) );
  XOR U31505 ( .A(n32539), .B(n32540), .Z(n32537) );
  XOR U31506 ( .A(n32541), .B(n32542), .Z(n32525) );
  XNOR U31507 ( .A(n32543), .B(n32544), .Z(n32542) );
  ANDN U31508 ( .B(n32545), .A(n32546), .Z(n32543) );
  XNOR U31509 ( .A(n32547), .B(n32548), .Z(n32545) );
  IV U31510 ( .A(n32523), .Z(n32541) );
  XOR U31511 ( .A(n32549), .B(n32550), .Z(n32523) );
  ANDN U31512 ( .B(n32551), .A(n32552), .Z(n32549) );
  XOR U31513 ( .A(n32550), .B(n32553), .Z(n32551) );
  XOR U31514 ( .A(n32532), .B(n32463), .Z(n32533) );
  XOR U31515 ( .A(n32554), .B(n32555), .Z(n32463) );
  AND U31516 ( .A(n890), .B(n32556), .Z(n32554) );
  XOR U31517 ( .A(n32557), .B(n32555), .Z(n32556) );
  XNOR U31518 ( .A(n32558), .B(n32559), .Z(n32532) );
  NAND U31519 ( .A(n32560), .B(n32561), .Z(n32559) );
  XOR U31520 ( .A(n32562), .B(n32511), .Z(n32561) );
  XOR U31521 ( .A(n32552), .B(n32553), .Z(n32511) );
  XOR U31522 ( .A(n32563), .B(n32540), .Z(n32553) );
  XOR U31523 ( .A(n32564), .B(n32565), .Z(n32540) );
  ANDN U31524 ( .B(n32566), .A(n32567), .Z(n32564) );
  XOR U31525 ( .A(n32565), .B(n32568), .Z(n32566) );
  IV U31526 ( .A(n32538), .Z(n32563) );
  XOR U31527 ( .A(n32536), .B(n32569), .Z(n32538) );
  XOR U31528 ( .A(n32570), .B(n32571), .Z(n32569) );
  ANDN U31529 ( .B(n32572), .A(n32573), .Z(n32570) );
  XOR U31530 ( .A(n32574), .B(n32571), .Z(n32572) );
  IV U31531 ( .A(n32539), .Z(n32536) );
  XOR U31532 ( .A(n32575), .B(n32576), .Z(n32539) );
  ANDN U31533 ( .B(n32577), .A(n32578), .Z(n32575) );
  XOR U31534 ( .A(n32576), .B(n32579), .Z(n32577) );
  XOR U31535 ( .A(n32580), .B(n32581), .Z(n32552) );
  XNOR U31536 ( .A(n32547), .B(n32582), .Z(n32581) );
  IV U31537 ( .A(n32550), .Z(n32582) );
  XOR U31538 ( .A(n32583), .B(n32584), .Z(n32550) );
  ANDN U31539 ( .B(n32585), .A(n32586), .Z(n32583) );
  XOR U31540 ( .A(n32584), .B(n32587), .Z(n32585) );
  XNOR U31541 ( .A(n32588), .B(n32589), .Z(n32547) );
  ANDN U31542 ( .B(n32590), .A(n32591), .Z(n32588) );
  XOR U31543 ( .A(n32589), .B(n32592), .Z(n32590) );
  IV U31544 ( .A(n32546), .Z(n32580) );
  XOR U31545 ( .A(n32544), .B(n32593), .Z(n32546) );
  XOR U31546 ( .A(n32594), .B(n32595), .Z(n32593) );
  ANDN U31547 ( .B(n32596), .A(n32597), .Z(n32594) );
  XOR U31548 ( .A(n32598), .B(n32595), .Z(n32596) );
  IV U31549 ( .A(n32548), .Z(n32544) );
  XOR U31550 ( .A(n32599), .B(n32600), .Z(n32548) );
  ANDN U31551 ( .B(n32601), .A(n32602), .Z(n32599) );
  XOR U31552 ( .A(n32603), .B(n32600), .Z(n32601) );
  IV U31553 ( .A(n32558), .Z(n32562) );
  XOR U31554 ( .A(n32558), .B(n32513), .Z(n32560) );
  XOR U31555 ( .A(n32604), .B(n32605), .Z(n32513) );
  AND U31556 ( .A(n890), .B(n32606), .Z(n32604) );
  XOR U31557 ( .A(n32607), .B(n32605), .Z(n32606) );
  NANDN U31558 ( .A(n32515), .B(n32517), .Z(n32558) );
  XOR U31559 ( .A(n32608), .B(n32609), .Z(n32517) );
  AND U31560 ( .A(n890), .B(n32610), .Z(n32608) );
  XOR U31561 ( .A(n32609), .B(n32611), .Z(n32610) );
  XNOR U31562 ( .A(n32612), .B(n32613), .Z(n890) );
  AND U31563 ( .A(n32614), .B(n32615), .Z(n32612) );
  XOR U31564 ( .A(n32613), .B(n32528), .Z(n32615) );
  XNOR U31565 ( .A(n32616), .B(n32617), .Z(n32528) );
  ANDN U31566 ( .B(n32618), .A(n32619), .Z(n32616) );
  XOR U31567 ( .A(n32617), .B(n32620), .Z(n32618) );
  XNOR U31568 ( .A(n32613), .B(n32530), .Z(n32614) );
  XOR U31569 ( .A(n32621), .B(n32622), .Z(n32530) );
  AND U31570 ( .A(n894), .B(n32623), .Z(n32621) );
  XOR U31571 ( .A(n32624), .B(n32622), .Z(n32623) );
  XNOR U31572 ( .A(n32625), .B(n32626), .Z(n32613) );
  AND U31573 ( .A(n32627), .B(n32628), .Z(n32625) );
  XNOR U31574 ( .A(n32626), .B(n32555), .Z(n32628) );
  XOR U31575 ( .A(n32619), .B(n32620), .Z(n32555) );
  XNOR U31576 ( .A(n32629), .B(n32630), .Z(n32620) );
  ANDN U31577 ( .B(n32631), .A(n32632), .Z(n32629) );
  XOR U31578 ( .A(n32633), .B(n32634), .Z(n32631) );
  XOR U31579 ( .A(n32635), .B(n32636), .Z(n32619) );
  XNOR U31580 ( .A(n32637), .B(n32638), .Z(n32636) );
  ANDN U31581 ( .B(n32639), .A(n32640), .Z(n32637) );
  XNOR U31582 ( .A(n32641), .B(n32642), .Z(n32639) );
  IV U31583 ( .A(n32617), .Z(n32635) );
  XOR U31584 ( .A(n32643), .B(n32644), .Z(n32617) );
  ANDN U31585 ( .B(n32645), .A(n32646), .Z(n32643) );
  XOR U31586 ( .A(n32644), .B(n32647), .Z(n32645) );
  XOR U31587 ( .A(n32626), .B(n32557), .Z(n32627) );
  XOR U31588 ( .A(n32648), .B(n32649), .Z(n32557) );
  AND U31589 ( .A(n894), .B(n32650), .Z(n32648) );
  XOR U31590 ( .A(n32651), .B(n32649), .Z(n32650) );
  XNOR U31591 ( .A(n32652), .B(n32653), .Z(n32626) );
  NAND U31592 ( .A(n32654), .B(n32655), .Z(n32653) );
  XOR U31593 ( .A(n32656), .B(n32605), .Z(n32655) );
  XOR U31594 ( .A(n32646), .B(n32647), .Z(n32605) );
  XOR U31595 ( .A(n32657), .B(n32634), .Z(n32647) );
  XOR U31596 ( .A(n32658), .B(n32659), .Z(n32634) );
  ANDN U31597 ( .B(n32660), .A(n32661), .Z(n32658) );
  XOR U31598 ( .A(n32659), .B(n32662), .Z(n32660) );
  IV U31599 ( .A(n32632), .Z(n32657) );
  XOR U31600 ( .A(n32630), .B(n32663), .Z(n32632) );
  XOR U31601 ( .A(n32664), .B(n32665), .Z(n32663) );
  ANDN U31602 ( .B(n32666), .A(n32667), .Z(n32664) );
  XOR U31603 ( .A(n32668), .B(n32665), .Z(n32666) );
  IV U31604 ( .A(n32633), .Z(n32630) );
  XOR U31605 ( .A(n32669), .B(n32670), .Z(n32633) );
  ANDN U31606 ( .B(n32671), .A(n32672), .Z(n32669) );
  XOR U31607 ( .A(n32670), .B(n32673), .Z(n32671) );
  XOR U31608 ( .A(n32674), .B(n32675), .Z(n32646) );
  XNOR U31609 ( .A(n32641), .B(n32676), .Z(n32675) );
  IV U31610 ( .A(n32644), .Z(n32676) );
  XOR U31611 ( .A(n32677), .B(n32678), .Z(n32644) );
  ANDN U31612 ( .B(n32679), .A(n32680), .Z(n32677) );
  XOR U31613 ( .A(n32678), .B(n32681), .Z(n32679) );
  XNOR U31614 ( .A(n32682), .B(n32683), .Z(n32641) );
  ANDN U31615 ( .B(n32684), .A(n32685), .Z(n32682) );
  XOR U31616 ( .A(n32683), .B(n32686), .Z(n32684) );
  IV U31617 ( .A(n32640), .Z(n32674) );
  XOR U31618 ( .A(n32638), .B(n32687), .Z(n32640) );
  XOR U31619 ( .A(n32688), .B(n32689), .Z(n32687) );
  ANDN U31620 ( .B(n32690), .A(n32691), .Z(n32688) );
  XOR U31621 ( .A(n32692), .B(n32689), .Z(n32690) );
  IV U31622 ( .A(n32642), .Z(n32638) );
  XOR U31623 ( .A(n32693), .B(n32694), .Z(n32642) );
  ANDN U31624 ( .B(n32695), .A(n32696), .Z(n32693) );
  XOR U31625 ( .A(n32697), .B(n32694), .Z(n32695) );
  IV U31626 ( .A(n32652), .Z(n32656) );
  XOR U31627 ( .A(n32652), .B(n32607), .Z(n32654) );
  XOR U31628 ( .A(n32698), .B(n32699), .Z(n32607) );
  AND U31629 ( .A(n894), .B(n32700), .Z(n32698) );
  XOR U31630 ( .A(n32701), .B(n32699), .Z(n32700) );
  NANDN U31631 ( .A(n32609), .B(n32611), .Z(n32652) );
  XOR U31632 ( .A(n32702), .B(n32703), .Z(n32611) );
  AND U31633 ( .A(n894), .B(n32704), .Z(n32702) );
  XOR U31634 ( .A(n32703), .B(n32705), .Z(n32704) );
  XNOR U31635 ( .A(n32706), .B(n32707), .Z(n894) );
  AND U31636 ( .A(n32708), .B(n32709), .Z(n32706) );
  XOR U31637 ( .A(n32707), .B(n32622), .Z(n32709) );
  XNOR U31638 ( .A(n32710), .B(n32711), .Z(n32622) );
  ANDN U31639 ( .B(n32712), .A(n32713), .Z(n32710) );
  XOR U31640 ( .A(n32711), .B(n32714), .Z(n32712) );
  XNOR U31641 ( .A(n32707), .B(n32624), .Z(n32708) );
  XOR U31642 ( .A(n32715), .B(n32716), .Z(n32624) );
  AND U31643 ( .A(n898), .B(n32717), .Z(n32715) );
  XOR U31644 ( .A(n32718), .B(n32716), .Z(n32717) );
  XNOR U31645 ( .A(n32719), .B(n32720), .Z(n32707) );
  AND U31646 ( .A(n32721), .B(n32722), .Z(n32719) );
  XNOR U31647 ( .A(n32720), .B(n32649), .Z(n32722) );
  XOR U31648 ( .A(n32713), .B(n32714), .Z(n32649) );
  XNOR U31649 ( .A(n32723), .B(n32724), .Z(n32714) );
  ANDN U31650 ( .B(n32725), .A(n32726), .Z(n32723) );
  XOR U31651 ( .A(n32727), .B(n32728), .Z(n32725) );
  XOR U31652 ( .A(n32729), .B(n32730), .Z(n32713) );
  XNOR U31653 ( .A(n32731), .B(n32732), .Z(n32730) );
  ANDN U31654 ( .B(n32733), .A(n32734), .Z(n32731) );
  XNOR U31655 ( .A(n32735), .B(n32736), .Z(n32733) );
  IV U31656 ( .A(n32711), .Z(n32729) );
  XOR U31657 ( .A(n32737), .B(n32738), .Z(n32711) );
  ANDN U31658 ( .B(n32739), .A(n32740), .Z(n32737) );
  XOR U31659 ( .A(n32738), .B(n32741), .Z(n32739) );
  XOR U31660 ( .A(n32720), .B(n32651), .Z(n32721) );
  XOR U31661 ( .A(n32742), .B(n32743), .Z(n32651) );
  AND U31662 ( .A(n898), .B(n32744), .Z(n32742) );
  XOR U31663 ( .A(n32745), .B(n32743), .Z(n32744) );
  XNOR U31664 ( .A(n32746), .B(n32747), .Z(n32720) );
  NAND U31665 ( .A(n32748), .B(n32749), .Z(n32747) );
  XOR U31666 ( .A(n32750), .B(n32699), .Z(n32749) );
  XOR U31667 ( .A(n32740), .B(n32741), .Z(n32699) );
  XOR U31668 ( .A(n32751), .B(n32728), .Z(n32741) );
  XOR U31669 ( .A(n32752), .B(n32753), .Z(n32728) );
  ANDN U31670 ( .B(n32754), .A(n32755), .Z(n32752) );
  XOR U31671 ( .A(n32753), .B(n32756), .Z(n32754) );
  IV U31672 ( .A(n32726), .Z(n32751) );
  XOR U31673 ( .A(n32724), .B(n32757), .Z(n32726) );
  XOR U31674 ( .A(n32758), .B(n32759), .Z(n32757) );
  ANDN U31675 ( .B(n32760), .A(n32761), .Z(n32758) );
  XOR U31676 ( .A(n32762), .B(n32759), .Z(n32760) );
  IV U31677 ( .A(n32727), .Z(n32724) );
  XOR U31678 ( .A(n32763), .B(n32764), .Z(n32727) );
  ANDN U31679 ( .B(n32765), .A(n32766), .Z(n32763) );
  XOR U31680 ( .A(n32764), .B(n32767), .Z(n32765) );
  XOR U31681 ( .A(n32768), .B(n32769), .Z(n32740) );
  XNOR U31682 ( .A(n32735), .B(n32770), .Z(n32769) );
  IV U31683 ( .A(n32738), .Z(n32770) );
  XOR U31684 ( .A(n32771), .B(n32772), .Z(n32738) );
  ANDN U31685 ( .B(n32773), .A(n32774), .Z(n32771) );
  XOR U31686 ( .A(n32772), .B(n32775), .Z(n32773) );
  XNOR U31687 ( .A(n32776), .B(n32777), .Z(n32735) );
  ANDN U31688 ( .B(n32778), .A(n32779), .Z(n32776) );
  XOR U31689 ( .A(n32777), .B(n32780), .Z(n32778) );
  IV U31690 ( .A(n32734), .Z(n32768) );
  XOR U31691 ( .A(n32732), .B(n32781), .Z(n32734) );
  XOR U31692 ( .A(n32782), .B(n32783), .Z(n32781) );
  ANDN U31693 ( .B(n32784), .A(n32785), .Z(n32782) );
  XOR U31694 ( .A(n32786), .B(n32783), .Z(n32784) );
  IV U31695 ( .A(n32736), .Z(n32732) );
  XOR U31696 ( .A(n32787), .B(n32788), .Z(n32736) );
  ANDN U31697 ( .B(n32789), .A(n32790), .Z(n32787) );
  XOR U31698 ( .A(n32791), .B(n32788), .Z(n32789) );
  IV U31699 ( .A(n32746), .Z(n32750) );
  XOR U31700 ( .A(n32746), .B(n32701), .Z(n32748) );
  XOR U31701 ( .A(n32792), .B(n32793), .Z(n32701) );
  AND U31702 ( .A(n898), .B(n32794), .Z(n32792) );
  XOR U31703 ( .A(n32795), .B(n32793), .Z(n32794) );
  NANDN U31704 ( .A(n32703), .B(n32705), .Z(n32746) );
  XOR U31705 ( .A(n32796), .B(n32797), .Z(n32705) );
  AND U31706 ( .A(n898), .B(n32798), .Z(n32796) );
  XOR U31707 ( .A(n32797), .B(n32799), .Z(n32798) );
  XNOR U31708 ( .A(n32800), .B(n32801), .Z(n898) );
  AND U31709 ( .A(n32802), .B(n32803), .Z(n32800) );
  XOR U31710 ( .A(n32801), .B(n32716), .Z(n32803) );
  XNOR U31711 ( .A(n32804), .B(n32805), .Z(n32716) );
  ANDN U31712 ( .B(n32806), .A(n32807), .Z(n32804) );
  XOR U31713 ( .A(n32805), .B(n32808), .Z(n32806) );
  XNOR U31714 ( .A(n32801), .B(n32718), .Z(n32802) );
  XOR U31715 ( .A(n32809), .B(n32810), .Z(n32718) );
  AND U31716 ( .A(n902), .B(n32811), .Z(n32809) );
  XOR U31717 ( .A(n32812), .B(n32810), .Z(n32811) );
  XNOR U31718 ( .A(n32813), .B(n32814), .Z(n32801) );
  AND U31719 ( .A(n32815), .B(n32816), .Z(n32813) );
  XNOR U31720 ( .A(n32814), .B(n32743), .Z(n32816) );
  XOR U31721 ( .A(n32807), .B(n32808), .Z(n32743) );
  XNOR U31722 ( .A(n32817), .B(n32818), .Z(n32808) );
  ANDN U31723 ( .B(n32819), .A(n32820), .Z(n32817) );
  XOR U31724 ( .A(n32821), .B(n32822), .Z(n32819) );
  XOR U31725 ( .A(n32823), .B(n32824), .Z(n32807) );
  XNOR U31726 ( .A(n32825), .B(n32826), .Z(n32824) );
  ANDN U31727 ( .B(n32827), .A(n32828), .Z(n32825) );
  XNOR U31728 ( .A(n32829), .B(n32830), .Z(n32827) );
  IV U31729 ( .A(n32805), .Z(n32823) );
  XOR U31730 ( .A(n32831), .B(n32832), .Z(n32805) );
  ANDN U31731 ( .B(n32833), .A(n32834), .Z(n32831) );
  XOR U31732 ( .A(n32832), .B(n32835), .Z(n32833) );
  XOR U31733 ( .A(n32814), .B(n32745), .Z(n32815) );
  XOR U31734 ( .A(n32836), .B(n32837), .Z(n32745) );
  AND U31735 ( .A(n902), .B(n32838), .Z(n32836) );
  XOR U31736 ( .A(n32839), .B(n32837), .Z(n32838) );
  XNOR U31737 ( .A(n32840), .B(n32841), .Z(n32814) );
  NAND U31738 ( .A(n32842), .B(n32843), .Z(n32841) );
  XOR U31739 ( .A(n32844), .B(n32793), .Z(n32843) );
  XOR U31740 ( .A(n32834), .B(n32835), .Z(n32793) );
  XOR U31741 ( .A(n32845), .B(n32822), .Z(n32835) );
  XOR U31742 ( .A(n32846), .B(n32847), .Z(n32822) );
  ANDN U31743 ( .B(n32848), .A(n32849), .Z(n32846) );
  XOR U31744 ( .A(n32847), .B(n32850), .Z(n32848) );
  IV U31745 ( .A(n32820), .Z(n32845) );
  XOR U31746 ( .A(n32818), .B(n32851), .Z(n32820) );
  XOR U31747 ( .A(n32852), .B(n32853), .Z(n32851) );
  ANDN U31748 ( .B(n32854), .A(n32855), .Z(n32852) );
  XOR U31749 ( .A(n32856), .B(n32853), .Z(n32854) );
  IV U31750 ( .A(n32821), .Z(n32818) );
  XOR U31751 ( .A(n32857), .B(n32858), .Z(n32821) );
  ANDN U31752 ( .B(n32859), .A(n32860), .Z(n32857) );
  XOR U31753 ( .A(n32858), .B(n32861), .Z(n32859) );
  XOR U31754 ( .A(n32862), .B(n32863), .Z(n32834) );
  XNOR U31755 ( .A(n32829), .B(n32864), .Z(n32863) );
  IV U31756 ( .A(n32832), .Z(n32864) );
  XOR U31757 ( .A(n32865), .B(n32866), .Z(n32832) );
  ANDN U31758 ( .B(n32867), .A(n32868), .Z(n32865) );
  XOR U31759 ( .A(n32866), .B(n32869), .Z(n32867) );
  XNOR U31760 ( .A(n32870), .B(n32871), .Z(n32829) );
  ANDN U31761 ( .B(n32872), .A(n32873), .Z(n32870) );
  XOR U31762 ( .A(n32871), .B(n32874), .Z(n32872) );
  IV U31763 ( .A(n32828), .Z(n32862) );
  XOR U31764 ( .A(n32826), .B(n32875), .Z(n32828) );
  XOR U31765 ( .A(n32876), .B(n32877), .Z(n32875) );
  ANDN U31766 ( .B(n32878), .A(n32879), .Z(n32876) );
  XOR U31767 ( .A(n32880), .B(n32877), .Z(n32878) );
  IV U31768 ( .A(n32830), .Z(n32826) );
  XOR U31769 ( .A(n32881), .B(n32882), .Z(n32830) );
  ANDN U31770 ( .B(n32883), .A(n32884), .Z(n32881) );
  XOR U31771 ( .A(n32885), .B(n32882), .Z(n32883) );
  IV U31772 ( .A(n32840), .Z(n32844) );
  XOR U31773 ( .A(n32840), .B(n32795), .Z(n32842) );
  XOR U31774 ( .A(n32886), .B(n32887), .Z(n32795) );
  AND U31775 ( .A(n902), .B(n32888), .Z(n32886) );
  XOR U31776 ( .A(n32889), .B(n32887), .Z(n32888) );
  NANDN U31777 ( .A(n32797), .B(n32799), .Z(n32840) );
  XOR U31778 ( .A(n32890), .B(n32891), .Z(n32799) );
  AND U31779 ( .A(n902), .B(n32892), .Z(n32890) );
  XOR U31780 ( .A(n32891), .B(n32893), .Z(n32892) );
  XNOR U31781 ( .A(n32894), .B(n32895), .Z(n902) );
  AND U31782 ( .A(n32896), .B(n32897), .Z(n32894) );
  XOR U31783 ( .A(n32895), .B(n32810), .Z(n32897) );
  XNOR U31784 ( .A(n32898), .B(n32899), .Z(n32810) );
  ANDN U31785 ( .B(n32900), .A(n32901), .Z(n32898) );
  XOR U31786 ( .A(n32899), .B(n32902), .Z(n32900) );
  XNOR U31787 ( .A(n32895), .B(n32812), .Z(n32896) );
  XOR U31788 ( .A(n32903), .B(n32904), .Z(n32812) );
  AND U31789 ( .A(n906), .B(n32905), .Z(n32903) );
  XOR U31790 ( .A(n32906), .B(n32904), .Z(n32905) );
  XNOR U31791 ( .A(n32907), .B(n32908), .Z(n32895) );
  AND U31792 ( .A(n32909), .B(n32910), .Z(n32907) );
  XNOR U31793 ( .A(n32908), .B(n32837), .Z(n32910) );
  XOR U31794 ( .A(n32901), .B(n32902), .Z(n32837) );
  XNOR U31795 ( .A(n32911), .B(n32912), .Z(n32902) );
  ANDN U31796 ( .B(n32913), .A(n32914), .Z(n32911) );
  XOR U31797 ( .A(n32915), .B(n32916), .Z(n32913) );
  XOR U31798 ( .A(n32917), .B(n32918), .Z(n32901) );
  XNOR U31799 ( .A(n32919), .B(n32920), .Z(n32918) );
  ANDN U31800 ( .B(n32921), .A(n32922), .Z(n32919) );
  XNOR U31801 ( .A(n32923), .B(n32924), .Z(n32921) );
  IV U31802 ( .A(n32899), .Z(n32917) );
  XOR U31803 ( .A(n32925), .B(n32926), .Z(n32899) );
  ANDN U31804 ( .B(n32927), .A(n32928), .Z(n32925) );
  XOR U31805 ( .A(n32926), .B(n32929), .Z(n32927) );
  XOR U31806 ( .A(n32908), .B(n32839), .Z(n32909) );
  XOR U31807 ( .A(n32930), .B(n32931), .Z(n32839) );
  AND U31808 ( .A(n906), .B(n32932), .Z(n32930) );
  XOR U31809 ( .A(n32933), .B(n32931), .Z(n32932) );
  XNOR U31810 ( .A(n32934), .B(n32935), .Z(n32908) );
  NAND U31811 ( .A(n32936), .B(n32937), .Z(n32935) );
  XOR U31812 ( .A(n32938), .B(n32887), .Z(n32937) );
  XOR U31813 ( .A(n32928), .B(n32929), .Z(n32887) );
  XOR U31814 ( .A(n32939), .B(n32916), .Z(n32929) );
  XOR U31815 ( .A(n32940), .B(n32941), .Z(n32916) );
  ANDN U31816 ( .B(n32942), .A(n32943), .Z(n32940) );
  XOR U31817 ( .A(n32941), .B(n32944), .Z(n32942) );
  IV U31818 ( .A(n32914), .Z(n32939) );
  XOR U31819 ( .A(n32912), .B(n32945), .Z(n32914) );
  XOR U31820 ( .A(n32946), .B(n32947), .Z(n32945) );
  ANDN U31821 ( .B(n32948), .A(n32949), .Z(n32946) );
  XOR U31822 ( .A(n32950), .B(n32947), .Z(n32948) );
  IV U31823 ( .A(n32915), .Z(n32912) );
  XOR U31824 ( .A(n32951), .B(n32952), .Z(n32915) );
  ANDN U31825 ( .B(n32953), .A(n32954), .Z(n32951) );
  XOR U31826 ( .A(n32952), .B(n32955), .Z(n32953) );
  XOR U31827 ( .A(n32956), .B(n32957), .Z(n32928) );
  XNOR U31828 ( .A(n32923), .B(n32958), .Z(n32957) );
  IV U31829 ( .A(n32926), .Z(n32958) );
  XOR U31830 ( .A(n32959), .B(n32960), .Z(n32926) );
  ANDN U31831 ( .B(n32961), .A(n32962), .Z(n32959) );
  XOR U31832 ( .A(n32960), .B(n32963), .Z(n32961) );
  XNOR U31833 ( .A(n32964), .B(n32965), .Z(n32923) );
  ANDN U31834 ( .B(n32966), .A(n32967), .Z(n32964) );
  XOR U31835 ( .A(n32965), .B(n32968), .Z(n32966) );
  IV U31836 ( .A(n32922), .Z(n32956) );
  XOR U31837 ( .A(n32920), .B(n32969), .Z(n32922) );
  XOR U31838 ( .A(n32970), .B(n32971), .Z(n32969) );
  ANDN U31839 ( .B(n32972), .A(n32973), .Z(n32970) );
  XOR U31840 ( .A(n32974), .B(n32971), .Z(n32972) );
  IV U31841 ( .A(n32924), .Z(n32920) );
  XOR U31842 ( .A(n32975), .B(n32976), .Z(n32924) );
  ANDN U31843 ( .B(n32977), .A(n32978), .Z(n32975) );
  XOR U31844 ( .A(n32979), .B(n32976), .Z(n32977) );
  IV U31845 ( .A(n32934), .Z(n32938) );
  XOR U31846 ( .A(n32934), .B(n32889), .Z(n32936) );
  XOR U31847 ( .A(n32980), .B(n32981), .Z(n32889) );
  AND U31848 ( .A(n906), .B(n32982), .Z(n32980) );
  XOR U31849 ( .A(n32983), .B(n32981), .Z(n32982) );
  NANDN U31850 ( .A(n32891), .B(n32893), .Z(n32934) );
  XOR U31851 ( .A(n32984), .B(n32985), .Z(n32893) );
  AND U31852 ( .A(n906), .B(n32986), .Z(n32984) );
  XOR U31853 ( .A(n32985), .B(n32987), .Z(n32986) );
  XNOR U31854 ( .A(n32988), .B(n32989), .Z(n906) );
  AND U31855 ( .A(n32990), .B(n32991), .Z(n32988) );
  XOR U31856 ( .A(n32989), .B(n32904), .Z(n32991) );
  XNOR U31857 ( .A(n32992), .B(n32993), .Z(n32904) );
  ANDN U31858 ( .B(n32994), .A(n32995), .Z(n32992) );
  XOR U31859 ( .A(n32993), .B(n32996), .Z(n32994) );
  XNOR U31860 ( .A(n32989), .B(n32906), .Z(n32990) );
  XOR U31861 ( .A(n32997), .B(n32998), .Z(n32906) );
  AND U31862 ( .A(n910), .B(n32999), .Z(n32997) );
  XOR U31863 ( .A(n33000), .B(n32998), .Z(n32999) );
  XNOR U31864 ( .A(n33001), .B(n33002), .Z(n32989) );
  AND U31865 ( .A(n33003), .B(n33004), .Z(n33001) );
  XNOR U31866 ( .A(n33002), .B(n32931), .Z(n33004) );
  XOR U31867 ( .A(n32995), .B(n32996), .Z(n32931) );
  XNOR U31868 ( .A(n33005), .B(n33006), .Z(n32996) );
  ANDN U31869 ( .B(n33007), .A(n33008), .Z(n33005) );
  XOR U31870 ( .A(n33009), .B(n33010), .Z(n33007) );
  XOR U31871 ( .A(n33011), .B(n33012), .Z(n32995) );
  XNOR U31872 ( .A(n33013), .B(n33014), .Z(n33012) );
  ANDN U31873 ( .B(n33015), .A(n33016), .Z(n33013) );
  XNOR U31874 ( .A(n33017), .B(n33018), .Z(n33015) );
  IV U31875 ( .A(n32993), .Z(n33011) );
  XOR U31876 ( .A(n33019), .B(n33020), .Z(n32993) );
  ANDN U31877 ( .B(n33021), .A(n33022), .Z(n33019) );
  XOR U31878 ( .A(n33020), .B(n33023), .Z(n33021) );
  XOR U31879 ( .A(n33002), .B(n32933), .Z(n33003) );
  XOR U31880 ( .A(n33024), .B(n33025), .Z(n32933) );
  AND U31881 ( .A(n910), .B(n33026), .Z(n33024) );
  XOR U31882 ( .A(n33027), .B(n33025), .Z(n33026) );
  XNOR U31883 ( .A(n33028), .B(n33029), .Z(n33002) );
  NAND U31884 ( .A(n33030), .B(n33031), .Z(n33029) );
  XOR U31885 ( .A(n33032), .B(n32981), .Z(n33031) );
  XOR U31886 ( .A(n33022), .B(n33023), .Z(n32981) );
  XOR U31887 ( .A(n33033), .B(n33010), .Z(n33023) );
  XOR U31888 ( .A(n33034), .B(n33035), .Z(n33010) );
  ANDN U31889 ( .B(n33036), .A(n33037), .Z(n33034) );
  XOR U31890 ( .A(n33035), .B(n33038), .Z(n33036) );
  IV U31891 ( .A(n33008), .Z(n33033) );
  XOR U31892 ( .A(n33006), .B(n33039), .Z(n33008) );
  XOR U31893 ( .A(n33040), .B(n33041), .Z(n33039) );
  ANDN U31894 ( .B(n33042), .A(n33043), .Z(n33040) );
  XOR U31895 ( .A(n33044), .B(n33041), .Z(n33042) );
  IV U31896 ( .A(n33009), .Z(n33006) );
  XOR U31897 ( .A(n33045), .B(n33046), .Z(n33009) );
  ANDN U31898 ( .B(n33047), .A(n33048), .Z(n33045) );
  XOR U31899 ( .A(n33046), .B(n33049), .Z(n33047) );
  XOR U31900 ( .A(n33050), .B(n33051), .Z(n33022) );
  XNOR U31901 ( .A(n33017), .B(n33052), .Z(n33051) );
  IV U31902 ( .A(n33020), .Z(n33052) );
  XOR U31903 ( .A(n33053), .B(n33054), .Z(n33020) );
  ANDN U31904 ( .B(n33055), .A(n33056), .Z(n33053) );
  XOR U31905 ( .A(n33054), .B(n33057), .Z(n33055) );
  XNOR U31906 ( .A(n33058), .B(n33059), .Z(n33017) );
  ANDN U31907 ( .B(n33060), .A(n33061), .Z(n33058) );
  XOR U31908 ( .A(n33059), .B(n33062), .Z(n33060) );
  IV U31909 ( .A(n33016), .Z(n33050) );
  XOR U31910 ( .A(n33014), .B(n33063), .Z(n33016) );
  XOR U31911 ( .A(n33064), .B(n33065), .Z(n33063) );
  ANDN U31912 ( .B(n33066), .A(n33067), .Z(n33064) );
  XOR U31913 ( .A(n33068), .B(n33065), .Z(n33066) );
  IV U31914 ( .A(n33018), .Z(n33014) );
  XOR U31915 ( .A(n33069), .B(n33070), .Z(n33018) );
  ANDN U31916 ( .B(n33071), .A(n33072), .Z(n33069) );
  XOR U31917 ( .A(n33073), .B(n33070), .Z(n33071) );
  IV U31918 ( .A(n33028), .Z(n33032) );
  XOR U31919 ( .A(n33028), .B(n32983), .Z(n33030) );
  XOR U31920 ( .A(n33074), .B(n33075), .Z(n32983) );
  AND U31921 ( .A(n910), .B(n33076), .Z(n33074) );
  XOR U31922 ( .A(n33077), .B(n33075), .Z(n33076) );
  NANDN U31923 ( .A(n32985), .B(n32987), .Z(n33028) );
  XOR U31924 ( .A(n33078), .B(n33079), .Z(n32987) );
  AND U31925 ( .A(n910), .B(n33080), .Z(n33078) );
  XOR U31926 ( .A(n33079), .B(n33081), .Z(n33080) );
  XNOR U31927 ( .A(n33082), .B(n33083), .Z(n910) );
  AND U31928 ( .A(n33084), .B(n33085), .Z(n33082) );
  XOR U31929 ( .A(n33083), .B(n32998), .Z(n33085) );
  XNOR U31930 ( .A(n33086), .B(n33087), .Z(n32998) );
  ANDN U31931 ( .B(n33088), .A(n33089), .Z(n33086) );
  XOR U31932 ( .A(n33087), .B(n33090), .Z(n33088) );
  XNOR U31933 ( .A(n33083), .B(n33000), .Z(n33084) );
  XOR U31934 ( .A(n33091), .B(n33092), .Z(n33000) );
  AND U31935 ( .A(n914), .B(n33093), .Z(n33091) );
  XOR U31936 ( .A(n33094), .B(n33092), .Z(n33093) );
  XNOR U31937 ( .A(n33095), .B(n33096), .Z(n33083) );
  AND U31938 ( .A(n33097), .B(n33098), .Z(n33095) );
  XNOR U31939 ( .A(n33096), .B(n33025), .Z(n33098) );
  XOR U31940 ( .A(n33089), .B(n33090), .Z(n33025) );
  XNOR U31941 ( .A(n33099), .B(n33100), .Z(n33090) );
  ANDN U31942 ( .B(n33101), .A(n33102), .Z(n33099) );
  XOR U31943 ( .A(n33103), .B(n33104), .Z(n33101) );
  XOR U31944 ( .A(n33105), .B(n33106), .Z(n33089) );
  XNOR U31945 ( .A(n33107), .B(n33108), .Z(n33106) );
  ANDN U31946 ( .B(n33109), .A(n33110), .Z(n33107) );
  XNOR U31947 ( .A(n33111), .B(n33112), .Z(n33109) );
  IV U31948 ( .A(n33087), .Z(n33105) );
  XOR U31949 ( .A(n33113), .B(n33114), .Z(n33087) );
  ANDN U31950 ( .B(n33115), .A(n33116), .Z(n33113) );
  XOR U31951 ( .A(n33114), .B(n33117), .Z(n33115) );
  XOR U31952 ( .A(n33096), .B(n33027), .Z(n33097) );
  XOR U31953 ( .A(n33118), .B(n33119), .Z(n33027) );
  AND U31954 ( .A(n914), .B(n33120), .Z(n33118) );
  XOR U31955 ( .A(n33121), .B(n33119), .Z(n33120) );
  XNOR U31956 ( .A(n33122), .B(n33123), .Z(n33096) );
  NAND U31957 ( .A(n33124), .B(n33125), .Z(n33123) );
  XOR U31958 ( .A(n33126), .B(n33075), .Z(n33125) );
  XOR U31959 ( .A(n33116), .B(n33117), .Z(n33075) );
  XOR U31960 ( .A(n33127), .B(n33104), .Z(n33117) );
  XOR U31961 ( .A(n33128), .B(n33129), .Z(n33104) );
  ANDN U31962 ( .B(n33130), .A(n33131), .Z(n33128) );
  XOR U31963 ( .A(n33129), .B(n33132), .Z(n33130) );
  IV U31964 ( .A(n33102), .Z(n33127) );
  XOR U31965 ( .A(n33100), .B(n33133), .Z(n33102) );
  XOR U31966 ( .A(n33134), .B(n33135), .Z(n33133) );
  ANDN U31967 ( .B(n33136), .A(n33137), .Z(n33134) );
  XOR U31968 ( .A(n33138), .B(n33135), .Z(n33136) );
  IV U31969 ( .A(n33103), .Z(n33100) );
  XOR U31970 ( .A(n33139), .B(n33140), .Z(n33103) );
  ANDN U31971 ( .B(n33141), .A(n33142), .Z(n33139) );
  XOR U31972 ( .A(n33140), .B(n33143), .Z(n33141) );
  XOR U31973 ( .A(n33144), .B(n33145), .Z(n33116) );
  XNOR U31974 ( .A(n33111), .B(n33146), .Z(n33145) );
  IV U31975 ( .A(n33114), .Z(n33146) );
  XOR U31976 ( .A(n33147), .B(n33148), .Z(n33114) );
  ANDN U31977 ( .B(n33149), .A(n33150), .Z(n33147) );
  XOR U31978 ( .A(n33148), .B(n33151), .Z(n33149) );
  XNOR U31979 ( .A(n33152), .B(n33153), .Z(n33111) );
  ANDN U31980 ( .B(n33154), .A(n33155), .Z(n33152) );
  XOR U31981 ( .A(n33153), .B(n33156), .Z(n33154) );
  IV U31982 ( .A(n33110), .Z(n33144) );
  XOR U31983 ( .A(n33108), .B(n33157), .Z(n33110) );
  XOR U31984 ( .A(n33158), .B(n33159), .Z(n33157) );
  ANDN U31985 ( .B(n33160), .A(n33161), .Z(n33158) );
  XOR U31986 ( .A(n33162), .B(n33159), .Z(n33160) );
  IV U31987 ( .A(n33112), .Z(n33108) );
  XOR U31988 ( .A(n33163), .B(n33164), .Z(n33112) );
  ANDN U31989 ( .B(n33165), .A(n33166), .Z(n33163) );
  XOR U31990 ( .A(n33167), .B(n33164), .Z(n33165) );
  IV U31991 ( .A(n33122), .Z(n33126) );
  XOR U31992 ( .A(n33122), .B(n33077), .Z(n33124) );
  XOR U31993 ( .A(n33168), .B(n33169), .Z(n33077) );
  AND U31994 ( .A(n914), .B(n33170), .Z(n33168) );
  XOR U31995 ( .A(n33171), .B(n33169), .Z(n33170) );
  NANDN U31996 ( .A(n33079), .B(n33081), .Z(n33122) );
  XOR U31997 ( .A(n33172), .B(n33173), .Z(n33081) );
  AND U31998 ( .A(n914), .B(n33174), .Z(n33172) );
  XOR U31999 ( .A(n33173), .B(n33175), .Z(n33174) );
  XNOR U32000 ( .A(n33176), .B(n33177), .Z(n914) );
  AND U32001 ( .A(n33178), .B(n33179), .Z(n33176) );
  XOR U32002 ( .A(n33177), .B(n33092), .Z(n33179) );
  XNOR U32003 ( .A(n33180), .B(n33181), .Z(n33092) );
  ANDN U32004 ( .B(n33182), .A(n33183), .Z(n33180) );
  XOR U32005 ( .A(n33181), .B(n33184), .Z(n33182) );
  XNOR U32006 ( .A(n33177), .B(n33094), .Z(n33178) );
  XOR U32007 ( .A(n33185), .B(n33186), .Z(n33094) );
  AND U32008 ( .A(n918), .B(n33187), .Z(n33185) );
  XOR U32009 ( .A(n33188), .B(n33186), .Z(n33187) );
  XNOR U32010 ( .A(n33189), .B(n33190), .Z(n33177) );
  AND U32011 ( .A(n33191), .B(n33192), .Z(n33189) );
  XNOR U32012 ( .A(n33190), .B(n33119), .Z(n33192) );
  XOR U32013 ( .A(n33183), .B(n33184), .Z(n33119) );
  XNOR U32014 ( .A(n33193), .B(n33194), .Z(n33184) );
  ANDN U32015 ( .B(n33195), .A(n33196), .Z(n33193) );
  XOR U32016 ( .A(n33197), .B(n33198), .Z(n33195) );
  XOR U32017 ( .A(n33199), .B(n33200), .Z(n33183) );
  XNOR U32018 ( .A(n33201), .B(n33202), .Z(n33200) );
  ANDN U32019 ( .B(n33203), .A(n33204), .Z(n33201) );
  XNOR U32020 ( .A(n33205), .B(n33206), .Z(n33203) );
  IV U32021 ( .A(n33181), .Z(n33199) );
  XOR U32022 ( .A(n33207), .B(n33208), .Z(n33181) );
  ANDN U32023 ( .B(n33209), .A(n33210), .Z(n33207) );
  XOR U32024 ( .A(n33208), .B(n33211), .Z(n33209) );
  XOR U32025 ( .A(n33190), .B(n33121), .Z(n33191) );
  XOR U32026 ( .A(n33212), .B(n33213), .Z(n33121) );
  AND U32027 ( .A(n918), .B(n33214), .Z(n33212) );
  XOR U32028 ( .A(n33215), .B(n33213), .Z(n33214) );
  XNOR U32029 ( .A(n33216), .B(n33217), .Z(n33190) );
  NAND U32030 ( .A(n33218), .B(n33219), .Z(n33217) );
  XOR U32031 ( .A(n33220), .B(n33169), .Z(n33219) );
  XOR U32032 ( .A(n33210), .B(n33211), .Z(n33169) );
  XOR U32033 ( .A(n33221), .B(n33198), .Z(n33211) );
  XOR U32034 ( .A(n33222), .B(n33223), .Z(n33198) );
  ANDN U32035 ( .B(n33224), .A(n33225), .Z(n33222) );
  XOR U32036 ( .A(n33223), .B(n33226), .Z(n33224) );
  IV U32037 ( .A(n33196), .Z(n33221) );
  XOR U32038 ( .A(n33194), .B(n33227), .Z(n33196) );
  XOR U32039 ( .A(n33228), .B(n33229), .Z(n33227) );
  ANDN U32040 ( .B(n33230), .A(n33231), .Z(n33228) );
  XOR U32041 ( .A(n33232), .B(n33229), .Z(n33230) );
  IV U32042 ( .A(n33197), .Z(n33194) );
  XOR U32043 ( .A(n33233), .B(n33234), .Z(n33197) );
  ANDN U32044 ( .B(n33235), .A(n33236), .Z(n33233) );
  XOR U32045 ( .A(n33234), .B(n33237), .Z(n33235) );
  XOR U32046 ( .A(n33238), .B(n33239), .Z(n33210) );
  XNOR U32047 ( .A(n33205), .B(n33240), .Z(n33239) );
  IV U32048 ( .A(n33208), .Z(n33240) );
  XOR U32049 ( .A(n33241), .B(n33242), .Z(n33208) );
  ANDN U32050 ( .B(n33243), .A(n33244), .Z(n33241) );
  XOR U32051 ( .A(n33242), .B(n33245), .Z(n33243) );
  XNOR U32052 ( .A(n33246), .B(n33247), .Z(n33205) );
  ANDN U32053 ( .B(n33248), .A(n33249), .Z(n33246) );
  XOR U32054 ( .A(n33247), .B(n33250), .Z(n33248) );
  IV U32055 ( .A(n33204), .Z(n33238) );
  XOR U32056 ( .A(n33202), .B(n33251), .Z(n33204) );
  XOR U32057 ( .A(n33252), .B(n33253), .Z(n33251) );
  ANDN U32058 ( .B(n33254), .A(n33255), .Z(n33252) );
  XOR U32059 ( .A(n33256), .B(n33253), .Z(n33254) );
  IV U32060 ( .A(n33206), .Z(n33202) );
  XOR U32061 ( .A(n33257), .B(n33258), .Z(n33206) );
  ANDN U32062 ( .B(n33259), .A(n33260), .Z(n33257) );
  XOR U32063 ( .A(n33261), .B(n33258), .Z(n33259) );
  IV U32064 ( .A(n33216), .Z(n33220) );
  XOR U32065 ( .A(n33216), .B(n33171), .Z(n33218) );
  XOR U32066 ( .A(n33262), .B(n33263), .Z(n33171) );
  AND U32067 ( .A(n918), .B(n33264), .Z(n33262) );
  XOR U32068 ( .A(n33265), .B(n33263), .Z(n33264) );
  NANDN U32069 ( .A(n33173), .B(n33175), .Z(n33216) );
  XOR U32070 ( .A(n33266), .B(n33267), .Z(n33175) );
  AND U32071 ( .A(n918), .B(n33268), .Z(n33266) );
  XOR U32072 ( .A(n33267), .B(n33269), .Z(n33268) );
  XNOR U32073 ( .A(n33270), .B(n33271), .Z(n918) );
  AND U32074 ( .A(n33272), .B(n33273), .Z(n33270) );
  XOR U32075 ( .A(n33271), .B(n33186), .Z(n33273) );
  XNOR U32076 ( .A(n33274), .B(n33275), .Z(n33186) );
  ANDN U32077 ( .B(n33276), .A(n33277), .Z(n33274) );
  XOR U32078 ( .A(n33275), .B(n33278), .Z(n33276) );
  XNOR U32079 ( .A(n33271), .B(n33188), .Z(n33272) );
  XOR U32080 ( .A(n33279), .B(n33280), .Z(n33188) );
  AND U32081 ( .A(n922), .B(n33281), .Z(n33279) );
  XOR U32082 ( .A(n33282), .B(n33280), .Z(n33281) );
  XNOR U32083 ( .A(n33283), .B(n33284), .Z(n33271) );
  AND U32084 ( .A(n33285), .B(n33286), .Z(n33283) );
  XNOR U32085 ( .A(n33284), .B(n33213), .Z(n33286) );
  XOR U32086 ( .A(n33277), .B(n33278), .Z(n33213) );
  XNOR U32087 ( .A(n33287), .B(n33288), .Z(n33278) );
  ANDN U32088 ( .B(n33289), .A(n33290), .Z(n33287) );
  XOR U32089 ( .A(n33291), .B(n33292), .Z(n33289) );
  XOR U32090 ( .A(n33293), .B(n33294), .Z(n33277) );
  XNOR U32091 ( .A(n33295), .B(n33296), .Z(n33294) );
  ANDN U32092 ( .B(n33297), .A(n33298), .Z(n33295) );
  XNOR U32093 ( .A(n33299), .B(n33300), .Z(n33297) );
  IV U32094 ( .A(n33275), .Z(n33293) );
  XOR U32095 ( .A(n33301), .B(n33302), .Z(n33275) );
  ANDN U32096 ( .B(n33303), .A(n33304), .Z(n33301) );
  XOR U32097 ( .A(n33302), .B(n33305), .Z(n33303) );
  XOR U32098 ( .A(n33284), .B(n33215), .Z(n33285) );
  XOR U32099 ( .A(n33306), .B(n33307), .Z(n33215) );
  AND U32100 ( .A(n922), .B(n33308), .Z(n33306) );
  XOR U32101 ( .A(n33309), .B(n33307), .Z(n33308) );
  XNOR U32102 ( .A(n33310), .B(n33311), .Z(n33284) );
  NAND U32103 ( .A(n33312), .B(n33313), .Z(n33311) );
  XOR U32104 ( .A(n33314), .B(n33263), .Z(n33313) );
  XOR U32105 ( .A(n33304), .B(n33305), .Z(n33263) );
  XOR U32106 ( .A(n33315), .B(n33292), .Z(n33305) );
  XOR U32107 ( .A(n33316), .B(n33317), .Z(n33292) );
  ANDN U32108 ( .B(n33318), .A(n33319), .Z(n33316) );
  XOR U32109 ( .A(n33317), .B(n33320), .Z(n33318) );
  IV U32110 ( .A(n33290), .Z(n33315) );
  XOR U32111 ( .A(n33288), .B(n33321), .Z(n33290) );
  XOR U32112 ( .A(n33322), .B(n33323), .Z(n33321) );
  ANDN U32113 ( .B(n33324), .A(n33325), .Z(n33322) );
  XOR U32114 ( .A(n33326), .B(n33323), .Z(n33324) );
  IV U32115 ( .A(n33291), .Z(n33288) );
  XOR U32116 ( .A(n33327), .B(n33328), .Z(n33291) );
  ANDN U32117 ( .B(n33329), .A(n33330), .Z(n33327) );
  XOR U32118 ( .A(n33328), .B(n33331), .Z(n33329) );
  XOR U32119 ( .A(n33332), .B(n33333), .Z(n33304) );
  XNOR U32120 ( .A(n33299), .B(n33334), .Z(n33333) );
  IV U32121 ( .A(n33302), .Z(n33334) );
  XOR U32122 ( .A(n33335), .B(n33336), .Z(n33302) );
  ANDN U32123 ( .B(n33337), .A(n33338), .Z(n33335) );
  XOR U32124 ( .A(n33336), .B(n33339), .Z(n33337) );
  XNOR U32125 ( .A(n33340), .B(n33341), .Z(n33299) );
  ANDN U32126 ( .B(n33342), .A(n33343), .Z(n33340) );
  XOR U32127 ( .A(n33341), .B(n33344), .Z(n33342) );
  IV U32128 ( .A(n33298), .Z(n33332) );
  XOR U32129 ( .A(n33296), .B(n33345), .Z(n33298) );
  XOR U32130 ( .A(n33346), .B(n33347), .Z(n33345) );
  ANDN U32131 ( .B(n33348), .A(n33349), .Z(n33346) );
  XOR U32132 ( .A(n33350), .B(n33347), .Z(n33348) );
  IV U32133 ( .A(n33300), .Z(n33296) );
  XOR U32134 ( .A(n33351), .B(n33352), .Z(n33300) );
  ANDN U32135 ( .B(n33353), .A(n33354), .Z(n33351) );
  XOR U32136 ( .A(n33355), .B(n33352), .Z(n33353) );
  IV U32137 ( .A(n33310), .Z(n33314) );
  XOR U32138 ( .A(n33310), .B(n33265), .Z(n33312) );
  XOR U32139 ( .A(n33356), .B(n33357), .Z(n33265) );
  AND U32140 ( .A(n922), .B(n33358), .Z(n33356) );
  XOR U32141 ( .A(n33359), .B(n33357), .Z(n33358) );
  NANDN U32142 ( .A(n33267), .B(n33269), .Z(n33310) );
  XOR U32143 ( .A(n33360), .B(n33361), .Z(n33269) );
  AND U32144 ( .A(n922), .B(n33362), .Z(n33360) );
  XOR U32145 ( .A(n33361), .B(n33363), .Z(n33362) );
  XNOR U32146 ( .A(n33364), .B(n33365), .Z(n922) );
  AND U32147 ( .A(n33366), .B(n33367), .Z(n33364) );
  XOR U32148 ( .A(n33365), .B(n33280), .Z(n33367) );
  XNOR U32149 ( .A(n33368), .B(n33369), .Z(n33280) );
  ANDN U32150 ( .B(n33370), .A(n33371), .Z(n33368) );
  XOR U32151 ( .A(n33369), .B(n33372), .Z(n33370) );
  XNOR U32152 ( .A(n33365), .B(n33282), .Z(n33366) );
  XOR U32153 ( .A(n33373), .B(n33374), .Z(n33282) );
  AND U32154 ( .A(n926), .B(n33375), .Z(n33373) );
  XOR U32155 ( .A(n33376), .B(n33374), .Z(n33375) );
  XNOR U32156 ( .A(n33377), .B(n33378), .Z(n33365) );
  AND U32157 ( .A(n33379), .B(n33380), .Z(n33377) );
  XNOR U32158 ( .A(n33378), .B(n33307), .Z(n33380) );
  XOR U32159 ( .A(n33371), .B(n33372), .Z(n33307) );
  XNOR U32160 ( .A(n33381), .B(n33382), .Z(n33372) );
  ANDN U32161 ( .B(n33383), .A(n33384), .Z(n33381) );
  XOR U32162 ( .A(n33385), .B(n33386), .Z(n33383) );
  XOR U32163 ( .A(n33387), .B(n33388), .Z(n33371) );
  XNOR U32164 ( .A(n33389), .B(n33390), .Z(n33388) );
  ANDN U32165 ( .B(n33391), .A(n33392), .Z(n33389) );
  XNOR U32166 ( .A(n33393), .B(n33394), .Z(n33391) );
  IV U32167 ( .A(n33369), .Z(n33387) );
  XOR U32168 ( .A(n33395), .B(n33396), .Z(n33369) );
  ANDN U32169 ( .B(n33397), .A(n33398), .Z(n33395) );
  XOR U32170 ( .A(n33396), .B(n33399), .Z(n33397) );
  XOR U32171 ( .A(n33378), .B(n33309), .Z(n33379) );
  XOR U32172 ( .A(n33400), .B(n33401), .Z(n33309) );
  AND U32173 ( .A(n926), .B(n33402), .Z(n33400) );
  XOR U32174 ( .A(n33403), .B(n33401), .Z(n33402) );
  XNOR U32175 ( .A(n33404), .B(n33405), .Z(n33378) );
  NAND U32176 ( .A(n33406), .B(n33407), .Z(n33405) );
  XOR U32177 ( .A(n33408), .B(n33357), .Z(n33407) );
  XOR U32178 ( .A(n33398), .B(n33399), .Z(n33357) );
  XOR U32179 ( .A(n33409), .B(n33386), .Z(n33399) );
  XOR U32180 ( .A(n33410), .B(n33411), .Z(n33386) );
  ANDN U32181 ( .B(n33412), .A(n33413), .Z(n33410) );
  XOR U32182 ( .A(n33411), .B(n33414), .Z(n33412) );
  IV U32183 ( .A(n33384), .Z(n33409) );
  XOR U32184 ( .A(n33382), .B(n33415), .Z(n33384) );
  XOR U32185 ( .A(n33416), .B(n33417), .Z(n33415) );
  ANDN U32186 ( .B(n33418), .A(n33419), .Z(n33416) );
  XOR U32187 ( .A(n33420), .B(n33417), .Z(n33418) );
  IV U32188 ( .A(n33385), .Z(n33382) );
  XOR U32189 ( .A(n33421), .B(n33422), .Z(n33385) );
  ANDN U32190 ( .B(n33423), .A(n33424), .Z(n33421) );
  XOR U32191 ( .A(n33422), .B(n33425), .Z(n33423) );
  XOR U32192 ( .A(n33426), .B(n33427), .Z(n33398) );
  XNOR U32193 ( .A(n33393), .B(n33428), .Z(n33427) );
  IV U32194 ( .A(n33396), .Z(n33428) );
  XOR U32195 ( .A(n33429), .B(n33430), .Z(n33396) );
  ANDN U32196 ( .B(n33431), .A(n33432), .Z(n33429) );
  XOR U32197 ( .A(n33430), .B(n33433), .Z(n33431) );
  XNOR U32198 ( .A(n33434), .B(n33435), .Z(n33393) );
  ANDN U32199 ( .B(n33436), .A(n33437), .Z(n33434) );
  XOR U32200 ( .A(n33435), .B(n33438), .Z(n33436) );
  IV U32201 ( .A(n33392), .Z(n33426) );
  XOR U32202 ( .A(n33390), .B(n33439), .Z(n33392) );
  XOR U32203 ( .A(n33440), .B(n33441), .Z(n33439) );
  ANDN U32204 ( .B(n33442), .A(n33443), .Z(n33440) );
  XOR U32205 ( .A(n33444), .B(n33441), .Z(n33442) );
  IV U32206 ( .A(n33394), .Z(n33390) );
  XOR U32207 ( .A(n33445), .B(n33446), .Z(n33394) );
  ANDN U32208 ( .B(n33447), .A(n33448), .Z(n33445) );
  XOR U32209 ( .A(n33449), .B(n33446), .Z(n33447) );
  IV U32210 ( .A(n33404), .Z(n33408) );
  XOR U32211 ( .A(n33404), .B(n33359), .Z(n33406) );
  XOR U32212 ( .A(n33450), .B(n33451), .Z(n33359) );
  AND U32213 ( .A(n926), .B(n33452), .Z(n33450) );
  XOR U32214 ( .A(n33453), .B(n33451), .Z(n33452) );
  NANDN U32215 ( .A(n33361), .B(n33363), .Z(n33404) );
  XOR U32216 ( .A(n33454), .B(n33455), .Z(n33363) );
  AND U32217 ( .A(n926), .B(n33456), .Z(n33454) );
  XOR U32218 ( .A(n33455), .B(n33457), .Z(n33456) );
  XNOR U32219 ( .A(n33458), .B(n33459), .Z(n926) );
  AND U32220 ( .A(n33460), .B(n33461), .Z(n33458) );
  XOR U32221 ( .A(n33459), .B(n33374), .Z(n33461) );
  XNOR U32222 ( .A(n33462), .B(n33463), .Z(n33374) );
  ANDN U32223 ( .B(n33464), .A(n33465), .Z(n33462) );
  XOR U32224 ( .A(n33463), .B(n33466), .Z(n33464) );
  XNOR U32225 ( .A(n33459), .B(n33376), .Z(n33460) );
  XOR U32226 ( .A(n33467), .B(n33468), .Z(n33376) );
  AND U32227 ( .A(n930), .B(n33469), .Z(n33467) );
  XOR U32228 ( .A(n33470), .B(n33468), .Z(n33469) );
  XNOR U32229 ( .A(n33471), .B(n33472), .Z(n33459) );
  AND U32230 ( .A(n33473), .B(n33474), .Z(n33471) );
  XNOR U32231 ( .A(n33472), .B(n33401), .Z(n33474) );
  XOR U32232 ( .A(n33465), .B(n33466), .Z(n33401) );
  XNOR U32233 ( .A(n33475), .B(n33476), .Z(n33466) );
  ANDN U32234 ( .B(n33477), .A(n33478), .Z(n33475) );
  XOR U32235 ( .A(n33479), .B(n33480), .Z(n33477) );
  XOR U32236 ( .A(n33481), .B(n33482), .Z(n33465) );
  XNOR U32237 ( .A(n33483), .B(n33484), .Z(n33482) );
  ANDN U32238 ( .B(n33485), .A(n33486), .Z(n33483) );
  XNOR U32239 ( .A(n33487), .B(n33488), .Z(n33485) );
  IV U32240 ( .A(n33463), .Z(n33481) );
  XOR U32241 ( .A(n33489), .B(n33490), .Z(n33463) );
  ANDN U32242 ( .B(n33491), .A(n33492), .Z(n33489) );
  XOR U32243 ( .A(n33490), .B(n33493), .Z(n33491) );
  XOR U32244 ( .A(n33472), .B(n33403), .Z(n33473) );
  XOR U32245 ( .A(n33494), .B(n33495), .Z(n33403) );
  AND U32246 ( .A(n930), .B(n33496), .Z(n33494) );
  XOR U32247 ( .A(n33497), .B(n33495), .Z(n33496) );
  XNOR U32248 ( .A(n33498), .B(n33499), .Z(n33472) );
  NAND U32249 ( .A(n33500), .B(n33501), .Z(n33499) );
  XOR U32250 ( .A(n33502), .B(n33451), .Z(n33501) );
  XOR U32251 ( .A(n33492), .B(n33493), .Z(n33451) );
  XOR U32252 ( .A(n33503), .B(n33480), .Z(n33493) );
  XOR U32253 ( .A(n33504), .B(n33505), .Z(n33480) );
  ANDN U32254 ( .B(n33506), .A(n33507), .Z(n33504) );
  XOR U32255 ( .A(n33505), .B(n33508), .Z(n33506) );
  IV U32256 ( .A(n33478), .Z(n33503) );
  XOR U32257 ( .A(n33476), .B(n33509), .Z(n33478) );
  XOR U32258 ( .A(n33510), .B(n33511), .Z(n33509) );
  ANDN U32259 ( .B(n33512), .A(n33513), .Z(n33510) );
  XOR U32260 ( .A(n33514), .B(n33511), .Z(n33512) );
  IV U32261 ( .A(n33479), .Z(n33476) );
  XOR U32262 ( .A(n33515), .B(n33516), .Z(n33479) );
  ANDN U32263 ( .B(n33517), .A(n33518), .Z(n33515) );
  XOR U32264 ( .A(n33516), .B(n33519), .Z(n33517) );
  XOR U32265 ( .A(n33520), .B(n33521), .Z(n33492) );
  XNOR U32266 ( .A(n33487), .B(n33522), .Z(n33521) );
  IV U32267 ( .A(n33490), .Z(n33522) );
  XOR U32268 ( .A(n33523), .B(n33524), .Z(n33490) );
  ANDN U32269 ( .B(n33525), .A(n33526), .Z(n33523) );
  XOR U32270 ( .A(n33524), .B(n33527), .Z(n33525) );
  XNOR U32271 ( .A(n33528), .B(n33529), .Z(n33487) );
  ANDN U32272 ( .B(n33530), .A(n33531), .Z(n33528) );
  XOR U32273 ( .A(n33529), .B(n33532), .Z(n33530) );
  IV U32274 ( .A(n33486), .Z(n33520) );
  XOR U32275 ( .A(n33484), .B(n33533), .Z(n33486) );
  XOR U32276 ( .A(n33534), .B(n33535), .Z(n33533) );
  ANDN U32277 ( .B(n33536), .A(n33537), .Z(n33534) );
  XOR U32278 ( .A(n33538), .B(n33535), .Z(n33536) );
  IV U32279 ( .A(n33488), .Z(n33484) );
  XOR U32280 ( .A(n33539), .B(n33540), .Z(n33488) );
  ANDN U32281 ( .B(n33541), .A(n33542), .Z(n33539) );
  XOR U32282 ( .A(n33543), .B(n33540), .Z(n33541) );
  IV U32283 ( .A(n33498), .Z(n33502) );
  XOR U32284 ( .A(n33498), .B(n33453), .Z(n33500) );
  XOR U32285 ( .A(n33544), .B(n33545), .Z(n33453) );
  AND U32286 ( .A(n930), .B(n33546), .Z(n33544) );
  XOR U32287 ( .A(n33547), .B(n33545), .Z(n33546) );
  NANDN U32288 ( .A(n33455), .B(n33457), .Z(n33498) );
  XOR U32289 ( .A(n33548), .B(n33549), .Z(n33457) );
  AND U32290 ( .A(n930), .B(n33550), .Z(n33548) );
  XOR U32291 ( .A(n33549), .B(n33551), .Z(n33550) );
  XNOR U32292 ( .A(n33552), .B(n33553), .Z(n930) );
  AND U32293 ( .A(n33554), .B(n33555), .Z(n33552) );
  XOR U32294 ( .A(n33553), .B(n33468), .Z(n33555) );
  XNOR U32295 ( .A(n33556), .B(n33557), .Z(n33468) );
  ANDN U32296 ( .B(n33558), .A(n33559), .Z(n33556) );
  XOR U32297 ( .A(n33557), .B(n33560), .Z(n33558) );
  XNOR U32298 ( .A(n33553), .B(n33470), .Z(n33554) );
  XOR U32299 ( .A(n33561), .B(n33562), .Z(n33470) );
  AND U32300 ( .A(n934), .B(n33563), .Z(n33561) );
  XOR U32301 ( .A(n33564), .B(n33562), .Z(n33563) );
  XNOR U32302 ( .A(n33565), .B(n33566), .Z(n33553) );
  AND U32303 ( .A(n33567), .B(n33568), .Z(n33565) );
  XNOR U32304 ( .A(n33566), .B(n33495), .Z(n33568) );
  XOR U32305 ( .A(n33559), .B(n33560), .Z(n33495) );
  XNOR U32306 ( .A(n33569), .B(n33570), .Z(n33560) );
  ANDN U32307 ( .B(n33571), .A(n33572), .Z(n33569) );
  XOR U32308 ( .A(n33573), .B(n33574), .Z(n33571) );
  XOR U32309 ( .A(n33575), .B(n33576), .Z(n33559) );
  XNOR U32310 ( .A(n33577), .B(n33578), .Z(n33576) );
  ANDN U32311 ( .B(n33579), .A(n33580), .Z(n33577) );
  XNOR U32312 ( .A(n33581), .B(n33582), .Z(n33579) );
  IV U32313 ( .A(n33557), .Z(n33575) );
  XOR U32314 ( .A(n33583), .B(n33584), .Z(n33557) );
  ANDN U32315 ( .B(n33585), .A(n33586), .Z(n33583) );
  XOR U32316 ( .A(n33584), .B(n33587), .Z(n33585) );
  XOR U32317 ( .A(n33566), .B(n33497), .Z(n33567) );
  XOR U32318 ( .A(n33588), .B(n33589), .Z(n33497) );
  AND U32319 ( .A(n934), .B(n33590), .Z(n33588) );
  XOR U32320 ( .A(n33591), .B(n33589), .Z(n33590) );
  XNOR U32321 ( .A(n33592), .B(n33593), .Z(n33566) );
  NAND U32322 ( .A(n33594), .B(n33595), .Z(n33593) );
  XOR U32323 ( .A(n33596), .B(n33545), .Z(n33595) );
  XOR U32324 ( .A(n33586), .B(n33587), .Z(n33545) );
  XOR U32325 ( .A(n33597), .B(n33574), .Z(n33587) );
  XOR U32326 ( .A(n33598), .B(n33599), .Z(n33574) );
  ANDN U32327 ( .B(n33600), .A(n33601), .Z(n33598) );
  XOR U32328 ( .A(n33599), .B(n33602), .Z(n33600) );
  IV U32329 ( .A(n33572), .Z(n33597) );
  XOR U32330 ( .A(n33570), .B(n33603), .Z(n33572) );
  XOR U32331 ( .A(n33604), .B(n33605), .Z(n33603) );
  ANDN U32332 ( .B(n33606), .A(n33607), .Z(n33604) );
  XOR U32333 ( .A(n33608), .B(n33605), .Z(n33606) );
  IV U32334 ( .A(n33573), .Z(n33570) );
  XOR U32335 ( .A(n33609), .B(n33610), .Z(n33573) );
  ANDN U32336 ( .B(n33611), .A(n33612), .Z(n33609) );
  XOR U32337 ( .A(n33610), .B(n33613), .Z(n33611) );
  XOR U32338 ( .A(n33614), .B(n33615), .Z(n33586) );
  XNOR U32339 ( .A(n33581), .B(n33616), .Z(n33615) );
  IV U32340 ( .A(n33584), .Z(n33616) );
  XOR U32341 ( .A(n33617), .B(n33618), .Z(n33584) );
  ANDN U32342 ( .B(n33619), .A(n33620), .Z(n33617) );
  XOR U32343 ( .A(n33618), .B(n33621), .Z(n33619) );
  XNOR U32344 ( .A(n33622), .B(n33623), .Z(n33581) );
  ANDN U32345 ( .B(n33624), .A(n33625), .Z(n33622) );
  XOR U32346 ( .A(n33623), .B(n33626), .Z(n33624) );
  IV U32347 ( .A(n33580), .Z(n33614) );
  XOR U32348 ( .A(n33578), .B(n33627), .Z(n33580) );
  XOR U32349 ( .A(n33628), .B(n33629), .Z(n33627) );
  ANDN U32350 ( .B(n33630), .A(n33631), .Z(n33628) );
  XOR U32351 ( .A(n33632), .B(n33629), .Z(n33630) );
  IV U32352 ( .A(n33582), .Z(n33578) );
  XOR U32353 ( .A(n33633), .B(n33634), .Z(n33582) );
  ANDN U32354 ( .B(n33635), .A(n33636), .Z(n33633) );
  XOR U32355 ( .A(n33637), .B(n33634), .Z(n33635) );
  IV U32356 ( .A(n33592), .Z(n33596) );
  XOR U32357 ( .A(n33592), .B(n33547), .Z(n33594) );
  XOR U32358 ( .A(n33638), .B(n33639), .Z(n33547) );
  AND U32359 ( .A(n934), .B(n33640), .Z(n33638) );
  XOR U32360 ( .A(n33641), .B(n33639), .Z(n33640) );
  NANDN U32361 ( .A(n33549), .B(n33551), .Z(n33592) );
  XOR U32362 ( .A(n33642), .B(n33643), .Z(n33551) );
  AND U32363 ( .A(n934), .B(n33644), .Z(n33642) );
  XOR U32364 ( .A(n33643), .B(n33645), .Z(n33644) );
  XNOR U32365 ( .A(n33646), .B(n33647), .Z(n934) );
  AND U32366 ( .A(n33648), .B(n33649), .Z(n33646) );
  XOR U32367 ( .A(n33647), .B(n33562), .Z(n33649) );
  XNOR U32368 ( .A(n33650), .B(n33651), .Z(n33562) );
  ANDN U32369 ( .B(n33652), .A(n33653), .Z(n33650) );
  XOR U32370 ( .A(n33651), .B(n33654), .Z(n33652) );
  XNOR U32371 ( .A(n33647), .B(n33564), .Z(n33648) );
  XOR U32372 ( .A(n33655), .B(n33656), .Z(n33564) );
  AND U32373 ( .A(n938), .B(n33657), .Z(n33655) );
  XOR U32374 ( .A(n33658), .B(n33656), .Z(n33657) );
  XNOR U32375 ( .A(n33659), .B(n33660), .Z(n33647) );
  AND U32376 ( .A(n33661), .B(n33662), .Z(n33659) );
  XNOR U32377 ( .A(n33660), .B(n33589), .Z(n33662) );
  XOR U32378 ( .A(n33653), .B(n33654), .Z(n33589) );
  XNOR U32379 ( .A(n33663), .B(n33664), .Z(n33654) );
  ANDN U32380 ( .B(n33665), .A(n33666), .Z(n33663) );
  XOR U32381 ( .A(n33667), .B(n33668), .Z(n33665) );
  XOR U32382 ( .A(n33669), .B(n33670), .Z(n33653) );
  XNOR U32383 ( .A(n33671), .B(n33672), .Z(n33670) );
  ANDN U32384 ( .B(n33673), .A(n33674), .Z(n33671) );
  XNOR U32385 ( .A(n33675), .B(n33676), .Z(n33673) );
  IV U32386 ( .A(n33651), .Z(n33669) );
  XOR U32387 ( .A(n33677), .B(n33678), .Z(n33651) );
  ANDN U32388 ( .B(n33679), .A(n33680), .Z(n33677) );
  XOR U32389 ( .A(n33678), .B(n33681), .Z(n33679) );
  XOR U32390 ( .A(n33660), .B(n33591), .Z(n33661) );
  XOR U32391 ( .A(n33682), .B(n33683), .Z(n33591) );
  AND U32392 ( .A(n938), .B(n33684), .Z(n33682) );
  XOR U32393 ( .A(n33685), .B(n33683), .Z(n33684) );
  XNOR U32394 ( .A(n33686), .B(n33687), .Z(n33660) );
  NAND U32395 ( .A(n33688), .B(n33689), .Z(n33687) );
  XOR U32396 ( .A(n33690), .B(n33639), .Z(n33689) );
  XOR U32397 ( .A(n33680), .B(n33681), .Z(n33639) );
  XOR U32398 ( .A(n33691), .B(n33668), .Z(n33681) );
  XOR U32399 ( .A(n33692), .B(n33693), .Z(n33668) );
  ANDN U32400 ( .B(n33694), .A(n33695), .Z(n33692) );
  XOR U32401 ( .A(n33693), .B(n33696), .Z(n33694) );
  IV U32402 ( .A(n33666), .Z(n33691) );
  XOR U32403 ( .A(n33664), .B(n33697), .Z(n33666) );
  XOR U32404 ( .A(n33698), .B(n33699), .Z(n33697) );
  ANDN U32405 ( .B(n33700), .A(n33701), .Z(n33698) );
  XOR U32406 ( .A(n33702), .B(n33699), .Z(n33700) );
  IV U32407 ( .A(n33667), .Z(n33664) );
  XOR U32408 ( .A(n33703), .B(n33704), .Z(n33667) );
  ANDN U32409 ( .B(n33705), .A(n33706), .Z(n33703) );
  XOR U32410 ( .A(n33704), .B(n33707), .Z(n33705) );
  XOR U32411 ( .A(n33708), .B(n33709), .Z(n33680) );
  XNOR U32412 ( .A(n33675), .B(n33710), .Z(n33709) );
  IV U32413 ( .A(n33678), .Z(n33710) );
  XOR U32414 ( .A(n33711), .B(n33712), .Z(n33678) );
  ANDN U32415 ( .B(n33713), .A(n33714), .Z(n33711) );
  XOR U32416 ( .A(n33712), .B(n33715), .Z(n33713) );
  XNOR U32417 ( .A(n33716), .B(n33717), .Z(n33675) );
  ANDN U32418 ( .B(n33718), .A(n33719), .Z(n33716) );
  XOR U32419 ( .A(n33717), .B(n33720), .Z(n33718) );
  IV U32420 ( .A(n33674), .Z(n33708) );
  XOR U32421 ( .A(n33672), .B(n33721), .Z(n33674) );
  XOR U32422 ( .A(n33722), .B(n33723), .Z(n33721) );
  ANDN U32423 ( .B(n33724), .A(n33725), .Z(n33722) );
  XOR U32424 ( .A(n33726), .B(n33723), .Z(n33724) );
  IV U32425 ( .A(n33676), .Z(n33672) );
  XOR U32426 ( .A(n33727), .B(n33728), .Z(n33676) );
  ANDN U32427 ( .B(n33729), .A(n33730), .Z(n33727) );
  XOR U32428 ( .A(n33731), .B(n33728), .Z(n33729) );
  IV U32429 ( .A(n33686), .Z(n33690) );
  XOR U32430 ( .A(n33686), .B(n33641), .Z(n33688) );
  XOR U32431 ( .A(n33732), .B(n33733), .Z(n33641) );
  AND U32432 ( .A(n938), .B(n33734), .Z(n33732) );
  XOR U32433 ( .A(n33735), .B(n33733), .Z(n33734) );
  NANDN U32434 ( .A(n33643), .B(n33645), .Z(n33686) );
  XOR U32435 ( .A(n33736), .B(n33737), .Z(n33645) );
  AND U32436 ( .A(n938), .B(n33738), .Z(n33736) );
  XOR U32437 ( .A(n33737), .B(n33739), .Z(n33738) );
  XNOR U32438 ( .A(n33740), .B(n33741), .Z(n938) );
  AND U32439 ( .A(n33742), .B(n33743), .Z(n33740) );
  XOR U32440 ( .A(n33741), .B(n33656), .Z(n33743) );
  XNOR U32441 ( .A(n33744), .B(n33745), .Z(n33656) );
  ANDN U32442 ( .B(n33746), .A(n33747), .Z(n33744) );
  XOR U32443 ( .A(n33745), .B(n33748), .Z(n33746) );
  XNOR U32444 ( .A(n33741), .B(n33658), .Z(n33742) );
  XOR U32445 ( .A(n33749), .B(n33750), .Z(n33658) );
  AND U32446 ( .A(n942), .B(n33751), .Z(n33749) );
  XOR U32447 ( .A(n33752), .B(n33750), .Z(n33751) );
  XNOR U32448 ( .A(n33753), .B(n33754), .Z(n33741) );
  AND U32449 ( .A(n33755), .B(n33756), .Z(n33753) );
  XNOR U32450 ( .A(n33754), .B(n33683), .Z(n33756) );
  XOR U32451 ( .A(n33747), .B(n33748), .Z(n33683) );
  XNOR U32452 ( .A(n33757), .B(n33758), .Z(n33748) );
  ANDN U32453 ( .B(n33759), .A(n33760), .Z(n33757) );
  XOR U32454 ( .A(n33761), .B(n33762), .Z(n33759) );
  XOR U32455 ( .A(n33763), .B(n33764), .Z(n33747) );
  XNOR U32456 ( .A(n33765), .B(n33766), .Z(n33764) );
  ANDN U32457 ( .B(n33767), .A(n33768), .Z(n33765) );
  XNOR U32458 ( .A(n33769), .B(n33770), .Z(n33767) );
  IV U32459 ( .A(n33745), .Z(n33763) );
  XOR U32460 ( .A(n33771), .B(n33772), .Z(n33745) );
  ANDN U32461 ( .B(n33773), .A(n33774), .Z(n33771) );
  XOR U32462 ( .A(n33772), .B(n33775), .Z(n33773) );
  XOR U32463 ( .A(n33754), .B(n33685), .Z(n33755) );
  XOR U32464 ( .A(n33776), .B(n33777), .Z(n33685) );
  AND U32465 ( .A(n942), .B(n33778), .Z(n33776) );
  XOR U32466 ( .A(n33779), .B(n33777), .Z(n33778) );
  XNOR U32467 ( .A(n33780), .B(n33781), .Z(n33754) );
  NAND U32468 ( .A(n33782), .B(n33783), .Z(n33781) );
  XOR U32469 ( .A(n33784), .B(n33733), .Z(n33783) );
  XOR U32470 ( .A(n33774), .B(n33775), .Z(n33733) );
  XOR U32471 ( .A(n33785), .B(n33762), .Z(n33775) );
  XOR U32472 ( .A(n33786), .B(n33787), .Z(n33762) );
  ANDN U32473 ( .B(n33788), .A(n33789), .Z(n33786) );
  XOR U32474 ( .A(n33787), .B(n33790), .Z(n33788) );
  IV U32475 ( .A(n33760), .Z(n33785) );
  XOR U32476 ( .A(n33758), .B(n33791), .Z(n33760) );
  XOR U32477 ( .A(n33792), .B(n33793), .Z(n33791) );
  ANDN U32478 ( .B(n33794), .A(n33795), .Z(n33792) );
  XOR U32479 ( .A(n33796), .B(n33793), .Z(n33794) );
  IV U32480 ( .A(n33761), .Z(n33758) );
  XOR U32481 ( .A(n33797), .B(n33798), .Z(n33761) );
  ANDN U32482 ( .B(n33799), .A(n33800), .Z(n33797) );
  XOR U32483 ( .A(n33798), .B(n33801), .Z(n33799) );
  XOR U32484 ( .A(n33802), .B(n33803), .Z(n33774) );
  XNOR U32485 ( .A(n33769), .B(n33804), .Z(n33803) );
  IV U32486 ( .A(n33772), .Z(n33804) );
  XOR U32487 ( .A(n33805), .B(n33806), .Z(n33772) );
  ANDN U32488 ( .B(n33807), .A(n33808), .Z(n33805) );
  XOR U32489 ( .A(n33806), .B(n33809), .Z(n33807) );
  XNOR U32490 ( .A(n33810), .B(n33811), .Z(n33769) );
  ANDN U32491 ( .B(n33812), .A(n33813), .Z(n33810) );
  XOR U32492 ( .A(n33811), .B(n33814), .Z(n33812) );
  IV U32493 ( .A(n33768), .Z(n33802) );
  XOR U32494 ( .A(n33766), .B(n33815), .Z(n33768) );
  XOR U32495 ( .A(n33816), .B(n33817), .Z(n33815) );
  ANDN U32496 ( .B(n33818), .A(n33819), .Z(n33816) );
  XOR U32497 ( .A(n33820), .B(n33817), .Z(n33818) );
  IV U32498 ( .A(n33770), .Z(n33766) );
  XOR U32499 ( .A(n33821), .B(n33822), .Z(n33770) );
  ANDN U32500 ( .B(n33823), .A(n33824), .Z(n33821) );
  XOR U32501 ( .A(n33825), .B(n33822), .Z(n33823) );
  IV U32502 ( .A(n33780), .Z(n33784) );
  XOR U32503 ( .A(n33780), .B(n33735), .Z(n33782) );
  XOR U32504 ( .A(n33826), .B(n33827), .Z(n33735) );
  AND U32505 ( .A(n942), .B(n33828), .Z(n33826) );
  XOR U32506 ( .A(n33829), .B(n33827), .Z(n33828) );
  NANDN U32507 ( .A(n33737), .B(n33739), .Z(n33780) );
  XOR U32508 ( .A(n33830), .B(n33831), .Z(n33739) );
  AND U32509 ( .A(n942), .B(n33832), .Z(n33830) );
  XOR U32510 ( .A(n33831), .B(n33833), .Z(n33832) );
  XNOR U32511 ( .A(n33834), .B(n33835), .Z(n942) );
  AND U32512 ( .A(n33836), .B(n33837), .Z(n33834) );
  XOR U32513 ( .A(n33835), .B(n33750), .Z(n33837) );
  XNOR U32514 ( .A(n33838), .B(n33839), .Z(n33750) );
  ANDN U32515 ( .B(n33840), .A(n33841), .Z(n33838) );
  XOR U32516 ( .A(n33839), .B(n33842), .Z(n33840) );
  XNOR U32517 ( .A(n33835), .B(n33752), .Z(n33836) );
  XOR U32518 ( .A(n33843), .B(n33844), .Z(n33752) );
  AND U32519 ( .A(n946), .B(n33845), .Z(n33843) );
  XOR U32520 ( .A(n33846), .B(n33844), .Z(n33845) );
  XNOR U32521 ( .A(n33847), .B(n33848), .Z(n33835) );
  AND U32522 ( .A(n33849), .B(n33850), .Z(n33847) );
  XNOR U32523 ( .A(n33848), .B(n33777), .Z(n33850) );
  XOR U32524 ( .A(n33841), .B(n33842), .Z(n33777) );
  XNOR U32525 ( .A(n33851), .B(n33852), .Z(n33842) );
  ANDN U32526 ( .B(n33853), .A(n33854), .Z(n33851) );
  XOR U32527 ( .A(n33855), .B(n33856), .Z(n33853) );
  XOR U32528 ( .A(n33857), .B(n33858), .Z(n33841) );
  XNOR U32529 ( .A(n33859), .B(n33860), .Z(n33858) );
  ANDN U32530 ( .B(n33861), .A(n33862), .Z(n33859) );
  XNOR U32531 ( .A(n33863), .B(n33864), .Z(n33861) );
  IV U32532 ( .A(n33839), .Z(n33857) );
  XOR U32533 ( .A(n33865), .B(n33866), .Z(n33839) );
  ANDN U32534 ( .B(n33867), .A(n33868), .Z(n33865) );
  XOR U32535 ( .A(n33866), .B(n33869), .Z(n33867) );
  XOR U32536 ( .A(n33848), .B(n33779), .Z(n33849) );
  XOR U32537 ( .A(n33870), .B(n33871), .Z(n33779) );
  AND U32538 ( .A(n946), .B(n33872), .Z(n33870) );
  XOR U32539 ( .A(n33873), .B(n33871), .Z(n33872) );
  XNOR U32540 ( .A(n33874), .B(n33875), .Z(n33848) );
  NAND U32541 ( .A(n33876), .B(n33877), .Z(n33875) );
  XOR U32542 ( .A(n33878), .B(n33827), .Z(n33877) );
  XOR U32543 ( .A(n33868), .B(n33869), .Z(n33827) );
  XOR U32544 ( .A(n33879), .B(n33856), .Z(n33869) );
  XOR U32545 ( .A(n33880), .B(n33881), .Z(n33856) );
  ANDN U32546 ( .B(n33882), .A(n33883), .Z(n33880) );
  XOR U32547 ( .A(n33881), .B(n33884), .Z(n33882) );
  IV U32548 ( .A(n33854), .Z(n33879) );
  XOR U32549 ( .A(n33852), .B(n33885), .Z(n33854) );
  XOR U32550 ( .A(n33886), .B(n33887), .Z(n33885) );
  ANDN U32551 ( .B(n33888), .A(n33889), .Z(n33886) );
  XOR U32552 ( .A(n33890), .B(n33887), .Z(n33888) );
  IV U32553 ( .A(n33855), .Z(n33852) );
  XOR U32554 ( .A(n33891), .B(n33892), .Z(n33855) );
  ANDN U32555 ( .B(n33893), .A(n33894), .Z(n33891) );
  XOR U32556 ( .A(n33892), .B(n33895), .Z(n33893) );
  XOR U32557 ( .A(n33896), .B(n33897), .Z(n33868) );
  XNOR U32558 ( .A(n33863), .B(n33898), .Z(n33897) );
  IV U32559 ( .A(n33866), .Z(n33898) );
  XOR U32560 ( .A(n33899), .B(n33900), .Z(n33866) );
  ANDN U32561 ( .B(n33901), .A(n33902), .Z(n33899) );
  XOR U32562 ( .A(n33900), .B(n33903), .Z(n33901) );
  XNOR U32563 ( .A(n33904), .B(n33905), .Z(n33863) );
  ANDN U32564 ( .B(n33906), .A(n33907), .Z(n33904) );
  XOR U32565 ( .A(n33905), .B(n33908), .Z(n33906) );
  IV U32566 ( .A(n33862), .Z(n33896) );
  XOR U32567 ( .A(n33860), .B(n33909), .Z(n33862) );
  XOR U32568 ( .A(n33910), .B(n33911), .Z(n33909) );
  ANDN U32569 ( .B(n33912), .A(n33913), .Z(n33910) );
  XOR U32570 ( .A(n33914), .B(n33911), .Z(n33912) );
  IV U32571 ( .A(n33864), .Z(n33860) );
  XOR U32572 ( .A(n33915), .B(n33916), .Z(n33864) );
  ANDN U32573 ( .B(n33917), .A(n33918), .Z(n33915) );
  XOR U32574 ( .A(n33919), .B(n33916), .Z(n33917) );
  IV U32575 ( .A(n33874), .Z(n33878) );
  XOR U32576 ( .A(n33874), .B(n33829), .Z(n33876) );
  XOR U32577 ( .A(n33920), .B(n33921), .Z(n33829) );
  AND U32578 ( .A(n946), .B(n33922), .Z(n33920) );
  XOR U32579 ( .A(n33923), .B(n33921), .Z(n33922) );
  NANDN U32580 ( .A(n33831), .B(n33833), .Z(n33874) );
  XOR U32581 ( .A(n33924), .B(n33925), .Z(n33833) );
  AND U32582 ( .A(n946), .B(n33926), .Z(n33924) );
  XOR U32583 ( .A(n33925), .B(n33927), .Z(n33926) );
  XNOR U32584 ( .A(n33928), .B(n33929), .Z(n946) );
  AND U32585 ( .A(n33930), .B(n33931), .Z(n33928) );
  XOR U32586 ( .A(n33929), .B(n33844), .Z(n33931) );
  XNOR U32587 ( .A(n33932), .B(n33933), .Z(n33844) );
  ANDN U32588 ( .B(n33934), .A(n33935), .Z(n33932) );
  XOR U32589 ( .A(n33933), .B(n33936), .Z(n33934) );
  XNOR U32590 ( .A(n33929), .B(n33846), .Z(n33930) );
  XOR U32591 ( .A(n33937), .B(n33938), .Z(n33846) );
  AND U32592 ( .A(n950), .B(n33939), .Z(n33937) );
  XOR U32593 ( .A(n33940), .B(n33938), .Z(n33939) );
  XNOR U32594 ( .A(n33941), .B(n33942), .Z(n33929) );
  AND U32595 ( .A(n33943), .B(n33944), .Z(n33941) );
  XNOR U32596 ( .A(n33942), .B(n33871), .Z(n33944) );
  XOR U32597 ( .A(n33935), .B(n33936), .Z(n33871) );
  XNOR U32598 ( .A(n33945), .B(n33946), .Z(n33936) );
  ANDN U32599 ( .B(n33947), .A(n33948), .Z(n33945) );
  XOR U32600 ( .A(n33949), .B(n33950), .Z(n33947) );
  XOR U32601 ( .A(n33951), .B(n33952), .Z(n33935) );
  XNOR U32602 ( .A(n33953), .B(n33954), .Z(n33952) );
  ANDN U32603 ( .B(n33955), .A(n33956), .Z(n33953) );
  XNOR U32604 ( .A(n33957), .B(n33958), .Z(n33955) );
  IV U32605 ( .A(n33933), .Z(n33951) );
  XOR U32606 ( .A(n33959), .B(n33960), .Z(n33933) );
  ANDN U32607 ( .B(n33961), .A(n33962), .Z(n33959) );
  XOR U32608 ( .A(n33960), .B(n33963), .Z(n33961) );
  XOR U32609 ( .A(n33942), .B(n33873), .Z(n33943) );
  XOR U32610 ( .A(n33964), .B(n33965), .Z(n33873) );
  AND U32611 ( .A(n950), .B(n33966), .Z(n33964) );
  XOR U32612 ( .A(n33967), .B(n33965), .Z(n33966) );
  XNOR U32613 ( .A(n33968), .B(n33969), .Z(n33942) );
  NAND U32614 ( .A(n33970), .B(n33971), .Z(n33969) );
  XOR U32615 ( .A(n33972), .B(n33921), .Z(n33971) );
  XOR U32616 ( .A(n33962), .B(n33963), .Z(n33921) );
  XOR U32617 ( .A(n33973), .B(n33950), .Z(n33963) );
  XOR U32618 ( .A(n33974), .B(n33975), .Z(n33950) );
  ANDN U32619 ( .B(n33976), .A(n33977), .Z(n33974) );
  XOR U32620 ( .A(n33975), .B(n33978), .Z(n33976) );
  IV U32621 ( .A(n33948), .Z(n33973) );
  XOR U32622 ( .A(n33946), .B(n33979), .Z(n33948) );
  XOR U32623 ( .A(n33980), .B(n33981), .Z(n33979) );
  ANDN U32624 ( .B(n33982), .A(n33983), .Z(n33980) );
  XOR U32625 ( .A(n33984), .B(n33981), .Z(n33982) );
  IV U32626 ( .A(n33949), .Z(n33946) );
  XOR U32627 ( .A(n33985), .B(n33986), .Z(n33949) );
  ANDN U32628 ( .B(n33987), .A(n33988), .Z(n33985) );
  XOR U32629 ( .A(n33986), .B(n33989), .Z(n33987) );
  XOR U32630 ( .A(n33990), .B(n33991), .Z(n33962) );
  XNOR U32631 ( .A(n33957), .B(n33992), .Z(n33991) );
  IV U32632 ( .A(n33960), .Z(n33992) );
  XOR U32633 ( .A(n33993), .B(n33994), .Z(n33960) );
  ANDN U32634 ( .B(n33995), .A(n33996), .Z(n33993) );
  XOR U32635 ( .A(n33994), .B(n33997), .Z(n33995) );
  XNOR U32636 ( .A(n33998), .B(n33999), .Z(n33957) );
  ANDN U32637 ( .B(n34000), .A(n34001), .Z(n33998) );
  XOR U32638 ( .A(n33999), .B(n34002), .Z(n34000) );
  IV U32639 ( .A(n33956), .Z(n33990) );
  XOR U32640 ( .A(n33954), .B(n34003), .Z(n33956) );
  XOR U32641 ( .A(n34004), .B(n34005), .Z(n34003) );
  ANDN U32642 ( .B(n34006), .A(n34007), .Z(n34004) );
  XOR U32643 ( .A(n34008), .B(n34005), .Z(n34006) );
  IV U32644 ( .A(n33958), .Z(n33954) );
  XOR U32645 ( .A(n34009), .B(n34010), .Z(n33958) );
  ANDN U32646 ( .B(n34011), .A(n34012), .Z(n34009) );
  XOR U32647 ( .A(n34013), .B(n34010), .Z(n34011) );
  IV U32648 ( .A(n33968), .Z(n33972) );
  XOR U32649 ( .A(n33968), .B(n33923), .Z(n33970) );
  XOR U32650 ( .A(n34014), .B(n34015), .Z(n33923) );
  AND U32651 ( .A(n950), .B(n34016), .Z(n34014) );
  XOR U32652 ( .A(n34017), .B(n34015), .Z(n34016) );
  NANDN U32653 ( .A(n33925), .B(n33927), .Z(n33968) );
  XOR U32654 ( .A(n34018), .B(n34019), .Z(n33927) );
  AND U32655 ( .A(n950), .B(n34020), .Z(n34018) );
  XOR U32656 ( .A(n34019), .B(n34021), .Z(n34020) );
  XNOR U32657 ( .A(n34022), .B(n34023), .Z(n950) );
  AND U32658 ( .A(n34024), .B(n34025), .Z(n34022) );
  XOR U32659 ( .A(n34023), .B(n33938), .Z(n34025) );
  XNOR U32660 ( .A(n34026), .B(n34027), .Z(n33938) );
  ANDN U32661 ( .B(n34028), .A(n34029), .Z(n34026) );
  XOR U32662 ( .A(n34027), .B(n34030), .Z(n34028) );
  XNOR U32663 ( .A(n34023), .B(n33940), .Z(n34024) );
  XOR U32664 ( .A(n34031), .B(n34032), .Z(n33940) );
  AND U32665 ( .A(n954), .B(n34033), .Z(n34031) );
  XOR U32666 ( .A(n34034), .B(n34032), .Z(n34033) );
  XNOR U32667 ( .A(n34035), .B(n34036), .Z(n34023) );
  AND U32668 ( .A(n34037), .B(n34038), .Z(n34035) );
  XNOR U32669 ( .A(n34036), .B(n33965), .Z(n34038) );
  XOR U32670 ( .A(n34029), .B(n34030), .Z(n33965) );
  XNOR U32671 ( .A(n34039), .B(n34040), .Z(n34030) );
  ANDN U32672 ( .B(n34041), .A(n34042), .Z(n34039) );
  XOR U32673 ( .A(n34043), .B(n34044), .Z(n34041) );
  XOR U32674 ( .A(n34045), .B(n34046), .Z(n34029) );
  XNOR U32675 ( .A(n34047), .B(n34048), .Z(n34046) );
  ANDN U32676 ( .B(n34049), .A(n34050), .Z(n34047) );
  XNOR U32677 ( .A(n34051), .B(n34052), .Z(n34049) );
  IV U32678 ( .A(n34027), .Z(n34045) );
  XOR U32679 ( .A(n34053), .B(n34054), .Z(n34027) );
  ANDN U32680 ( .B(n34055), .A(n34056), .Z(n34053) );
  XOR U32681 ( .A(n34054), .B(n34057), .Z(n34055) );
  XOR U32682 ( .A(n34036), .B(n33967), .Z(n34037) );
  XOR U32683 ( .A(n34058), .B(n34059), .Z(n33967) );
  AND U32684 ( .A(n954), .B(n34060), .Z(n34058) );
  XOR U32685 ( .A(n34061), .B(n34059), .Z(n34060) );
  XNOR U32686 ( .A(n34062), .B(n34063), .Z(n34036) );
  NAND U32687 ( .A(n34064), .B(n34065), .Z(n34063) );
  XOR U32688 ( .A(n34066), .B(n34015), .Z(n34065) );
  XOR U32689 ( .A(n34056), .B(n34057), .Z(n34015) );
  XOR U32690 ( .A(n34067), .B(n34044), .Z(n34057) );
  XOR U32691 ( .A(n34068), .B(n34069), .Z(n34044) );
  ANDN U32692 ( .B(n34070), .A(n34071), .Z(n34068) );
  XOR U32693 ( .A(n34069), .B(n34072), .Z(n34070) );
  IV U32694 ( .A(n34042), .Z(n34067) );
  XOR U32695 ( .A(n34040), .B(n34073), .Z(n34042) );
  XOR U32696 ( .A(n34074), .B(n34075), .Z(n34073) );
  ANDN U32697 ( .B(n34076), .A(n34077), .Z(n34074) );
  XOR U32698 ( .A(n34078), .B(n34075), .Z(n34076) );
  IV U32699 ( .A(n34043), .Z(n34040) );
  XOR U32700 ( .A(n34079), .B(n34080), .Z(n34043) );
  ANDN U32701 ( .B(n34081), .A(n34082), .Z(n34079) );
  XOR U32702 ( .A(n34080), .B(n34083), .Z(n34081) );
  XOR U32703 ( .A(n34084), .B(n34085), .Z(n34056) );
  XNOR U32704 ( .A(n34051), .B(n34086), .Z(n34085) );
  IV U32705 ( .A(n34054), .Z(n34086) );
  XOR U32706 ( .A(n34087), .B(n34088), .Z(n34054) );
  ANDN U32707 ( .B(n34089), .A(n34090), .Z(n34087) );
  XOR U32708 ( .A(n34088), .B(n34091), .Z(n34089) );
  XNOR U32709 ( .A(n34092), .B(n34093), .Z(n34051) );
  ANDN U32710 ( .B(n34094), .A(n34095), .Z(n34092) );
  XOR U32711 ( .A(n34093), .B(n34096), .Z(n34094) );
  IV U32712 ( .A(n34050), .Z(n34084) );
  XOR U32713 ( .A(n34048), .B(n34097), .Z(n34050) );
  XOR U32714 ( .A(n34098), .B(n34099), .Z(n34097) );
  ANDN U32715 ( .B(n34100), .A(n34101), .Z(n34098) );
  XOR U32716 ( .A(n34102), .B(n34099), .Z(n34100) );
  IV U32717 ( .A(n34052), .Z(n34048) );
  XOR U32718 ( .A(n34103), .B(n34104), .Z(n34052) );
  ANDN U32719 ( .B(n34105), .A(n34106), .Z(n34103) );
  XOR U32720 ( .A(n34107), .B(n34104), .Z(n34105) );
  IV U32721 ( .A(n34062), .Z(n34066) );
  XOR U32722 ( .A(n34062), .B(n34017), .Z(n34064) );
  XOR U32723 ( .A(n34108), .B(n34109), .Z(n34017) );
  AND U32724 ( .A(n954), .B(n34110), .Z(n34108) );
  XOR U32725 ( .A(n34111), .B(n34109), .Z(n34110) );
  NANDN U32726 ( .A(n34019), .B(n34021), .Z(n34062) );
  XOR U32727 ( .A(n34112), .B(n34113), .Z(n34021) );
  AND U32728 ( .A(n954), .B(n34114), .Z(n34112) );
  XOR U32729 ( .A(n34113), .B(n34115), .Z(n34114) );
  XNOR U32730 ( .A(n34116), .B(n34117), .Z(n954) );
  AND U32731 ( .A(n34118), .B(n34119), .Z(n34116) );
  XOR U32732 ( .A(n34117), .B(n34032), .Z(n34119) );
  XNOR U32733 ( .A(n34120), .B(n34121), .Z(n34032) );
  ANDN U32734 ( .B(n34122), .A(n34123), .Z(n34120) );
  XOR U32735 ( .A(n34121), .B(n34124), .Z(n34122) );
  XNOR U32736 ( .A(n34117), .B(n34034), .Z(n34118) );
  XOR U32737 ( .A(n34125), .B(n34126), .Z(n34034) );
  AND U32738 ( .A(n958), .B(n34127), .Z(n34125) );
  XOR U32739 ( .A(n34128), .B(n34126), .Z(n34127) );
  XNOR U32740 ( .A(n34129), .B(n34130), .Z(n34117) );
  AND U32741 ( .A(n34131), .B(n34132), .Z(n34129) );
  XNOR U32742 ( .A(n34130), .B(n34059), .Z(n34132) );
  XOR U32743 ( .A(n34123), .B(n34124), .Z(n34059) );
  XNOR U32744 ( .A(n34133), .B(n34134), .Z(n34124) );
  ANDN U32745 ( .B(n34135), .A(n34136), .Z(n34133) );
  XOR U32746 ( .A(n34137), .B(n34138), .Z(n34135) );
  XOR U32747 ( .A(n34139), .B(n34140), .Z(n34123) );
  XNOR U32748 ( .A(n34141), .B(n34142), .Z(n34140) );
  ANDN U32749 ( .B(n34143), .A(n34144), .Z(n34141) );
  XNOR U32750 ( .A(n34145), .B(n34146), .Z(n34143) );
  IV U32751 ( .A(n34121), .Z(n34139) );
  XOR U32752 ( .A(n34147), .B(n34148), .Z(n34121) );
  ANDN U32753 ( .B(n34149), .A(n34150), .Z(n34147) );
  XOR U32754 ( .A(n34148), .B(n34151), .Z(n34149) );
  XOR U32755 ( .A(n34130), .B(n34061), .Z(n34131) );
  XOR U32756 ( .A(n34152), .B(n34153), .Z(n34061) );
  AND U32757 ( .A(n958), .B(n34154), .Z(n34152) );
  XOR U32758 ( .A(n34155), .B(n34153), .Z(n34154) );
  XNOR U32759 ( .A(n34156), .B(n34157), .Z(n34130) );
  NAND U32760 ( .A(n34158), .B(n34159), .Z(n34157) );
  XOR U32761 ( .A(n34160), .B(n34109), .Z(n34159) );
  XOR U32762 ( .A(n34150), .B(n34151), .Z(n34109) );
  XOR U32763 ( .A(n34161), .B(n34138), .Z(n34151) );
  XOR U32764 ( .A(n34162), .B(n34163), .Z(n34138) );
  ANDN U32765 ( .B(n34164), .A(n34165), .Z(n34162) );
  XOR U32766 ( .A(n34163), .B(n34166), .Z(n34164) );
  IV U32767 ( .A(n34136), .Z(n34161) );
  XOR U32768 ( .A(n34134), .B(n34167), .Z(n34136) );
  XOR U32769 ( .A(n34168), .B(n34169), .Z(n34167) );
  ANDN U32770 ( .B(n34170), .A(n34171), .Z(n34168) );
  XOR U32771 ( .A(n34172), .B(n34169), .Z(n34170) );
  IV U32772 ( .A(n34137), .Z(n34134) );
  XOR U32773 ( .A(n34173), .B(n34174), .Z(n34137) );
  ANDN U32774 ( .B(n34175), .A(n34176), .Z(n34173) );
  XOR U32775 ( .A(n34174), .B(n34177), .Z(n34175) );
  XOR U32776 ( .A(n34178), .B(n34179), .Z(n34150) );
  XNOR U32777 ( .A(n34145), .B(n34180), .Z(n34179) );
  IV U32778 ( .A(n34148), .Z(n34180) );
  XOR U32779 ( .A(n34181), .B(n34182), .Z(n34148) );
  ANDN U32780 ( .B(n34183), .A(n34184), .Z(n34181) );
  XOR U32781 ( .A(n34182), .B(n34185), .Z(n34183) );
  XNOR U32782 ( .A(n34186), .B(n34187), .Z(n34145) );
  ANDN U32783 ( .B(n34188), .A(n34189), .Z(n34186) );
  XOR U32784 ( .A(n34187), .B(n34190), .Z(n34188) );
  IV U32785 ( .A(n34144), .Z(n34178) );
  XOR U32786 ( .A(n34142), .B(n34191), .Z(n34144) );
  XOR U32787 ( .A(n34192), .B(n34193), .Z(n34191) );
  ANDN U32788 ( .B(n34194), .A(n34195), .Z(n34192) );
  XOR U32789 ( .A(n34196), .B(n34193), .Z(n34194) );
  IV U32790 ( .A(n34146), .Z(n34142) );
  XOR U32791 ( .A(n34197), .B(n34198), .Z(n34146) );
  ANDN U32792 ( .B(n34199), .A(n34200), .Z(n34197) );
  XOR U32793 ( .A(n34201), .B(n34198), .Z(n34199) );
  IV U32794 ( .A(n34156), .Z(n34160) );
  XOR U32795 ( .A(n34156), .B(n34111), .Z(n34158) );
  XOR U32796 ( .A(n34202), .B(n34203), .Z(n34111) );
  AND U32797 ( .A(n958), .B(n34204), .Z(n34202) );
  XOR U32798 ( .A(n34205), .B(n34203), .Z(n34204) );
  NANDN U32799 ( .A(n34113), .B(n34115), .Z(n34156) );
  XOR U32800 ( .A(n34206), .B(n34207), .Z(n34115) );
  AND U32801 ( .A(n958), .B(n34208), .Z(n34206) );
  XOR U32802 ( .A(n34207), .B(n34209), .Z(n34208) );
  XNOR U32803 ( .A(n34210), .B(n34211), .Z(n958) );
  AND U32804 ( .A(n34212), .B(n34213), .Z(n34210) );
  XOR U32805 ( .A(n34211), .B(n34126), .Z(n34213) );
  XNOR U32806 ( .A(n34214), .B(n34215), .Z(n34126) );
  ANDN U32807 ( .B(n34216), .A(n34217), .Z(n34214) );
  XOR U32808 ( .A(n34215), .B(n34218), .Z(n34216) );
  XNOR U32809 ( .A(n34211), .B(n34128), .Z(n34212) );
  XOR U32810 ( .A(n34219), .B(n34220), .Z(n34128) );
  AND U32811 ( .A(n962), .B(n34221), .Z(n34219) );
  XOR U32812 ( .A(n34222), .B(n34220), .Z(n34221) );
  XNOR U32813 ( .A(n34223), .B(n34224), .Z(n34211) );
  AND U32814 ( .A(n34225), .B(n34226), .Z(n34223) );
  XNOR U32815 ( .A(n34224), .B(n34153), .Z(n34226) );
  XOR U32816 ( .A(n34217), .B(n34218), .Z(n34153) );
  XNOR U32817 ( .A(n34227), .B(n34228), .Z(n34218) );
  ANDN U32818 ( .B(n34229), .A(n34230), .Z(n34227) );
  XOR U32819 ( .A(n34231), .B(n34232), .Z(n34229) );
  XOR U32820 ( .A(n34233), .B(n34234), .Z(n34217) );
  XNOR U32821 ( .A(n34235), .B(n34236), .Z(n34234) );
  ANDN U32822 ( .B(n34237), .A(n34238), .Z(n34235) );
  XNOR U32823 ( .A(n34239), .B(n34240), .Z(n34237) );
  IV U32824 ( .A(n34215), .Z(n34233) );
  XOR U32825 ( .A(n34241), .B(n34242), .Z(n34215) );
  ANDN U32826 ( .B(n34243), .A(n34244), .Z(n34241) );
  XOR U32827 ( .A(n34242), .B(n34245), .Z(n34243) );
  XOR U32828 ( .A(n34224), .B(n34155), .Z(n34225) );
  XOR U32829 ( .A(n34246), .B(n34247), .Z(n34155) );
  AND U32830 ( .A(n962), .B(n34248), .Z(n34246) );
  XOR U32831 ( .A(n34249), .B(n34247), .Z(n34248) );
  XNOR U32832 ( .A(n34250), .B(n34251), .Z(n34224) );
  NAND U32833 ( .A(n34252), .B(n34253), .Z(n34251) );
  XOR U32834 ( .A(n34254), .B(n34203), .Z(n34253) );
  XOR U32835 ( .A(n34244), .B(n34245), .Z(n34203) );
  XOR U32836 ( .A(n34255), .B(n34232), .Z(n34245) );
  XOR U32837 ( .A(n34256), .B(n34257), .Z(n34232) );
  ANDN U32838 ( .B(n34258), .A(n34259), .Z(n34256) );
  XOR U32839 ( .A(n34257), .B(n34260), .Z(n34258) );
  IV U32840 ( .A(n34230), .Z(n34255) );
  XOR U32841 ( .A(n34228), .B(n34261), .Z(n34230) );
  XOR U32842 ( .A(n34262), .B(n34263), .Z(n34261) );
  ANDN U32843 ( .B(n34264), .A(n34265), .Z(n34262) );
  XOR U32844 ( .A(n34266), .B(n34263), .Z(n34264) );
  IV U32845 ( .A(n34231), .Z(n34228) );
  XOR U32846 ( .A(n34267), .B(n34268), .Z(n34231) );
  ANDN U32847 ( .B(n34269), .A(n34270), .Z(n34267) );
  XOR U32848 ( .A(n34268), .B(n34271), .Z(n34269) );
  XOR U32849 ( .A(n34272), .B(n34273), .Z(n34244) );
  XNOR U32850 ( .A(n34239), .B(n34274), .Z(n34273) );
  IV U32851 ( .A(n34242), .Z(n34274) );
  XOR U32852 ( .A(n34275), .B(n34276), .Z(n34242) );
  ANDN U32853 ( .B(n34277), .A(n34278), .Z(n34275) );
  XOR U32854 ( .A(n34276), .B(n34279), .Z(n34277) );
  XNOR U32855 ( .A(n34280), .B(n34281), .Z(n34239) );
  ANDN U32856 ( .B(n34282), .A(n34283), .Z(n34280) );
  XOR U32857 ( .A(n34281), .B(n34284), .Z(n34282) );
  IV U32858 ( .A(n34238), .Z(n34272) );
  XOR U32859 ( .A(n34236), .B(n34285), .Z(n34238) );
  XOR U32860 ( .A(n34286), .B(n34287), .Z(n34285) );
  ANDN U32861 ( .B(n34288), .A(n34289), .Z(n34286) );
  XOR U32862 ( .A(n34290), .B(n34287), .Z(n34288) );
  IV U32863 ( .A(n34240), .Z(n34236) );
  XOR U32864 ( .A(n34291), .B(n34292), .Z(n34240) );
  ANDN U32865 ( .B(n34293), .A(n34294), .Z(n34291) );
  XOR U32866 ( .A(n34295), .B(n34292), .Z(n34293) );
  IV U32867 ( .A(n34250), .Z(n34254) );
  XOR U32868 ( .A(n34250), .B(n34205), .Z(n34252) );
  XOR U32869 ( .A(n34296), .B(n34297), .Z(n34205) );
  AND U32870 ( .A(n962), .B(n34298), .Z(n34296) );
  XOR U32871 ( .A(n34299), .B(n34297), .Z(n34298) );
  NANDN U32872 ( .A(n34207), .B(n34209), .Z(n34250) );
  XOR U32873 ( .A(n34300), .B(n34301), .Z(n34209) );
  AND U32874 ( .A(n962), .B(n34302), .Z(n34300) );
  XOR U32875 ( .A(n34301), .B(n34303), .Z(n34302) );
  XNOR U32876 ( .A(n34304), .B(n34305), .Z(n962) );
  AND U32877 ( .A(n34306), .B(n34307), .Z(n34304) );
  XOR U32878 ( .A(n34305), .B(n34220), .Z(n34307) );
  XNOR U32879 ( .A(n34308), .B(n34309), .Z(n34220) );
  ANDN U32880 ( .B(n34310), .A(n34311), .Z(n34308) );
  XOR U32881 ( .A(n34309), .B(n34312), .Z(n34310) );
  XNOR U32882 ( .A(n34305), .B(n34222), .Z(n34306) );
  XOR U32883 ( .A(n34313), .B(n34314), .Z(n34222) );
  AND U32884 ( .A(n966), .B(n34315), .Z(n34313) );
  XOR U32885 ( .A(n34316), .B(n34314), .Z(n34315) );
  XNOR U32886 ( .A(n34317), .B(n34318), .Z(n34305) );
  AND U32887 ( .A(n34319), .B(n34320), .Z(n34317) );
  XNOR U32888 ( .A(n34318), .B(n34247), .Z(n34320) );
  XOR U32889 ( .A(n34311), .B(n34312), .Z(n34247) );
  XNOR U32890 ( .A(n34321), .B(n34322), .Z(n34312) );
  ANDN U32891 ( .B(n34323), .A(n34324), .Z(n34321) );
  XOR U32892 ( .A(n34325), .B(n34326), .Z(n34323) );
  XOR U32893 ( .A(n34327), .B(n34328), .Z(n34311) );
  XNOR U32894 ( .A(n34329), .B(n34330), .Z(n34328) );
  ANDN U32895 ( .B(n34331), .A(n34332), .Z(n34329) );
  XNOR U32896 ( .A(n34333), .B(n34334), .Z(n34331) );
  IV U32897 ( .A(n34309), .Z(n34327) );
  XOR U32898 ( .A(n34335), .B(n34336), .Z(n34309) );
  ANDN U32899 ( .B(n34337), .A(n34338), .Z(n34335) );
  XOR U32900 ( .A(n34336), .B(n34339), .Z(n34337) );
  XOR U32901 ( .A(n34318), .B(n34249), .Z(n34319) );
  XOR U32902 ( .A(n34340), .B(n34341), .Z(n34249) );
  AND U32903 ( .A(n966), .B(n34342), .Z(n34340) );
  XOR U32904 ( .A(n34343), .B(n34341), .Z(n34342) );
  XNOR U32905 ( .A(n34344), .B(n34345), .Z(n34318) );
  NAND U32906 ( .A(n34346), .B(n34347), .Z(n34345) );
  XOR U32907 ( .A(n34348), .B(n34297), .Z(n34347) );
  XOR U32908 ( .A(n34338), .B(n34339), .Z(n34297) );
  XOR U32909 ( .A(n34349), .B(n34326), .Z(n34339) );
  XOR U32910 ( .A(n34350), .B(n34351), .Z(n34326) );
  ANDN U32911 ( .B(n34352), .A(n34353), .Z(n34350) );
  XOR U32912 ( .A(n34351), .B(n34354), .Z(n34352) );
  IV U32913 ( .A(n34324), .Z(n34349) );
  XOR U32914 ( .A(n34322), .B(n34355), .Z(n34324) );
  XOR U32915 ( .A(n34356), .B(n34357), .Z(n34355) );
  ANDN U32916 ( .B(n34358), .A(n34359), .Z(n34356) );
  XOR U32917 ( .A(n34360), .B(n34357), .Z(n34358) );
  IV U32918 ( .A(n34325), .Z(n34322) );
  XOR U32919 ( .A(n34361), .B(n34362), .Z(n34325) );
  ANDN U32920 ( .B(n34363), .A(n34364), .Z(n34361) );
  XOR U32921 ( .A(n34362), .B(n34365), .Z(n34363) );
  XOR U32922 ( .A(n34366), .B(n34367), .Z(n34338) );
  XNOR U32923 ( .A(n34333), .B(n34368), .Z(n34367) );
  IV U32924 ( .A(n34336), .Z(n34368) );
  XOR U32925 ( .A(n34369), .B(n34370), .Z(n34336) );
  ANDN U32926 ( .B(n34371), .A(n34372), .Z(n34369) );
  XOR U32927 ( .A(n34370), .B(n34373), .Z(n34371) );
  XNOR U32928 ( .A(n34374), .B(n34375), .Z(n34333) );
  ANDN U32929 ( .B(n34376), .A(n34377), .Z(n34374) );
  XOR U32930 ( .A(n34375), .B(n34378), .Z(n34376) );
  IV U32931 ( .A(n34332), .Z(n34366) );
  XOR U32932 ( .A(n34330), .B(n34379), .Z(n34332) );
  XOR U32933 ( .A(n34380), .B(n34381), .Z(n34379) );
  ANDN U32934 ( .B(n34382), .A(n34383), .Z(n34380) );
  XOR U32935 ( .A(n34384), .B(n34381), .Z(n34382) );
  IV U32936 ( .A(n34334), .Z(n34330) );
  XOR U32937 ( .A(n34385), .B(n34386), .Z(n34334) );
  ANDN U32938 ( .B(n34387), .A(n34388), .Z(n34385) );
  XOR U32939 ( .A(n34389), .B(n34386), .Z(n34387) );
  IV U32940 ( .A(n34344), .Z(n34348) );
  XOR U32941 ( .A(n34344), .B(n34299), .Z(n34346) );
  XOR U32942 ( .A(n34390), .B(n34391), .Z(n34299) );
  AND U32943 ( .A(n966), .B(n34392), .Z(n34390) );
  XOR U32944 ( .A(n34393), .B(n34391), .Z(n34392) );
  NANDN U32945 ( .A(n34301), .B(n34303), .Z(n34344) );
  XOR U32946 ( .A(n34394), .B(n34395), .Z(n34303) );
  AND U32947 ( .A(n966), .B(n34396), .Z(n34394) );
  XOR U32948 ( .A(n34395), .B(n34397), .Z(n34396) );
  XNOR U32949 ( .A(n34398), .B(n34399), .Z(n966) );
  AND U32950 ( .A(n34400), .B(n34401), .Z(n34398) );
  XOR U32951 ( .A(n34399), .B(n34314), .Z(n34401) );
  XNOR U32952 ( .A(n34402), .B(n34403), .Z(n34314) );
  ANDN U32953 ( .B(n34404), .A(n34405), .Z(n34402) );
  XOR U32954 ( .A(n34403), .B(n34406), .Z(n34404) );
  XNOR U32955 ( .A(n34399), .B(n34316), .Z(n34400) );
  XOR U32956 ( .A(n34407), .B(n34408), .Z(n34316) );
  AND U32957 ( .A(n970), .B(n34409), .Z(n34407) );
  XOR U32958 ( .A(n34410), .B(n34408), .Z(n34409) );
  XNOR U32959 ( .A(n34411), .B(n34412), .Z(n34399) );
  AND U32960 ( .A(n34413), .B(n34414), .Z(n34411) );
  XNOR U32961 ( .A(n34412), .B(n34341), .Z(n34414) );
  XOR U32962 ( .A(n34405), .B(n34406), .Z(n34341) );
  XNOR U32963 ( .A(n34415), .B(n34416), .Z(n34406) );
  ANDN U32964 ( .B(n34417), .A(n34418), .Z(n34415) );
  XOR U32965 ( .A(n34419), .B(n34420), .Z(n34417) );
  XOR U32966 ( .A(n34421), .B(n34422), .Z(n34405) );
  XNOR U32967 ( .A(n34423), .B(n34424), .Z(n34422) );
  ANDN U32968 ( .B(n34425), .A(n34426), .Z(n34423) );
  XNOR U32969 ( .A(n34427), .B(n34428), .Z(n34425) );
  IV U32970 ( .A(n34403), .Z(n34421) );
  XOR U32971 ( .A(n34429), .B(n34430), .Z(n34403) );
  ANDN U32972 ( .B(n34431), .A(n34432), .Z(n34429) );
  XOR U32973 ( .A(n34430), .B(n34433), .Z(n34431) );
  XOR U32974 ( .A(n34412), .B(n34343), .Z(n34413) );
  XOR U32975 ( .A(n34434), .B(n34435), .Z(n34343) );
  AND U32976 ( .A(n970), .B(n34436), .Z(n34434) );
  XOR U32977 ( .A(n34437), .B(n34435), .Z(n34436) );
  XNOR U32978 ( .A(n34438), .B(n34439), .Z(n34412) );
  NAND U32979 ( .A(n34440), .B(n34441), .Z(n34439) );
  XOR U32980 ( .A(n34442), .B(n34391), .Z(n34441) );
  XOR U32981 ( .A(n34432), .B(n34433), .Z(n34391) );
  XOR U32982 ( .A(n34443), .B(n34420), .Z(n34433) );
  XOR U32983 ( .A(n34444), .B(n34445), .Z(n34420) );
  ANDN U32984 ( .B(n34446), .A(n34447), .Z(n34444) );
  XOR U32985 ( .A(n34445), .B(n34448), .Z(n34446) );
  IV U32986 ( .A(n34418), .Z(n34443) );
  XOR U32987 ( .A(n34416), .B(n34449), .Z(n34418) );
  XOR U32988 ( .A(n34450), .B(n34451), .Z(n34449) );
  ANDN U32989 ( .B(n34452), .A(n34453), .Z(n34450) );
  XOR U32990 ( .A(n34454), .B(n34451), .Z(n34452) );
  IV U32991 ( .A(n34419), .Z(n34416) );
  XOR U32992 ( .A(n34455), .B(n34456), .Z(n34419) );
  ANDN U32993 ( .B(n34457), .A(n34458), .Z(n34455) );
  XOR U32994 ( .A(n34456), .B(n34459), .Z(n34457) );
  XOR U32995 ( .A(n34460), .B(n34461), .Z(n34432) );
  XNOR U32996 ( .A(n34427), .B(n34462), .Z(n34461) );
  IV U32997 ( .A(n34430), .Z(n34462) );
  XOR U32998 ( .A(n34463), .B(n34464), .Z(n34430) );
  ANDN U32999 ( .B(n34465), .A(n34466), .Z(n34463) );
  XOR U33000 ( .A(n34464), .B(n34467), .Z(n34465) );
  XNOR U33001 ( .A(n34468), .B(n34469), .Z(n34427) );
  ANDN U33002 ( .B(n34470), .A(n34471), .Z(n34468) );
  XOR U33003 ( .A(n34469), .B(n34472), .Z(n34470) );
  IV U33004 ( .A(n34426), .Z(n34460) );
  XOR U33005 ( .A(n34424), .B(n34473), .Z(n34426) );
  XOR U33006 ( .A(n34474), .B(n34475), .Z(n34473) );
  ANDN U33007 ( .B(n34476), .A(n34477), .Z(n34474) );
  XOR U33008 ( .A(n34478), .B(n34475), .Z(n34476) );
  IV U33009 ( .A(n34428), .Z(n34424) );
  XOR U33010 ( .A(n34479), .B(n34480), .Z(n34428) );
  ANDN U33011 ( .B(n34481), .A(n34482), .Z(n34479) );
  XOR U33012 ( .A(n34483), .B(n34480), .Z(n34481) );
  IV U33013 ( .A(n34438), .Z(n34442) );
  XOR U33014 ( .A(n34438), .B(n34393), .Z(n34440) );
  XOR U33015 ( .A(n34484), .B(n34485), .Z(n34393) );
  AND U33016 ( .A(n970), .B(n34486), .Z(n34484) );
  XOR U33017 ( .A(n34487), .B(n34485), .Z(n34486) );
  NANDN U33018 ( .A(n34395), .B(n34397), .Z(n34438) );
  XOR U33019 ( .A(n34488), .B(n34489), .Z(n34397) );
  AND U33020 ( .A(n970), .B(n34490), .Z(n34488) );
  XOR U33021 ( .A(n34489), .B(n34491), .Z(n34490) );
  XNOR U33022 ( .A(n34492), .B(n34493), .Z(n970) );
  AND U33023 ( .A(n34494), .B(n34495), .Z(n34492) );
  XOR U33024 ( .A(n34493), .B(n34408), .Z(n34495) );
  XNOR U33025 ( .A(n34496), .B(n34497), .Z(n34408) );
  ANDN U33026 ( .B(n34498), .A(n34499), .Z(n34496) );
  XOR U33027 ( .A(n34497), .B(n34500), .Z(n34498) );
  XNOR U33028 ( .A(n34493), .B(n34410), .Z(n34494) );
  XOR U33029 ( .A(n34501), .B(n34502), .Z(n34410) );
  AND U33030 ( .A(n974), .B(n34503), .Z(n34501) );
  XOR U33031 ( .A(n34504), .B(n34502), .Z(n34503) );
  XNOR U33032 ( .A(n34505), .B(n34506), .Z(n34493) );
  AND U33033 ( .A(n34507), .B(n34508), .Z(n34505) );
  XNOR U33034 ( .A(n34506), .B(n34435), .Z(n34508) );
  XOR U33035 ( .A(n34499), .B(n34500), .Z(n34435) );
  XNOR U33036 ( .A(n34509), .B(n34510), .Z(n34500) );
  ANDN U33037 ( .B(n34511), .A(n34512), .Z(n34509) );
  XOR U33038 ( .A(n34513), .B(n34514), .Z(n34511) );
  XOR U33039 ( .A(n34515), .B(n34516), .Z(n34499) );
  XNOR U33040 ( .A(n34517), .B(n34518), .Z(n34516) );
  ANDN U33041 ( .B(n34519), .A(n34520), .Z(n34517) );
  XNOR U33042 ( .A(n34521), .B(n34522), .Z(n34519) );
  IV U33043 ( .A(n34497), .Z(n34515) );
  XOR U33044 ( .A(n34523), .B(n34524), .Z(n34497) );
  ANDN U33045 ( .B(n34525), .A(n34526), .Z(n34523) );
  XOR U33046 ( .A(n34524), .B(n34527), .Z(n34525) );
  XOR U33047 ( .A(n34506), .B(n34437), .Z(n34507) );
  XOR U33048 ( .A(n34528), .B(n34529), .Z(n34437) );
  AND U33049 ( .A(n974), .B(n34530), .Z(n34528) );
  XOR U33050 ( .A(n34531), .B(n34529), .Z(n34530) );
  XNOR U33051 ( .A(n34532), .B(n34533), .Z(n34506) );
  NAND U33052 ( .A(n34534), .B(n34535), .Z(n34533) );
  XOR U33053 ( .A(n34536), .B(n34485), .Z(n34535) );
  XOR U33054 ( .A(n34526), .B(n34527), .Z(n34485) );
  XOR U33055 ( .A(n34537), .B(n34514), .Z(n34527) );
  XOR U33056 ( .A(n34538), .B(n34539), .Z(n34514) );
  ANDN U33057 ( .B(n34540), .A(n34541), .Z(n34538) );
  XOR U33058 ( .A(n34539), .B(n34542), .Z(n34540) );
  IV U33059 ( .A(n34512), .Z(n34537) );
  XOR U33060 ( .A(n34510), .B(n34543), .Z(n34512) );
  XOR U33061 ( .A(n34544), .B(n34545), .Z(n34543) );
  ANDN U33062 ( .B(n34546), .A(n34547), .Z(n34544) );
  XOR U33063 ( .A(n34548), .B(n34545), .Z(n34546) );
  IV U33064 ( .A(n34513), .Z(n34510) );
  XOR U33065 ( .A(n34549), .B(n34550), .Z(n34513) );
  ANDN U33066 ( .B(n34551), .A(n34552), .Z(n34549) );
  XOR U33067 ( .A(n34550), .B(n34553), .Z(n34551) );
  XOR U33068 ( .A(n34554), .B(n34555), .Z(n34526) );
  XNOR U33069 ( .A(n34521), .B(n34556), .Z(n34555) );
  IV U33070 ( .A(n34524), .Z(n34556) );
  XOR U33071 ( .A(n34557), .B(n34558), .Z(n34524) );
  ANDN U33072 ( .B(n34559), .A(n34560), .Z(n34557) );
  XOR U33073 ( .A(n34558), .B(n34561), .Z(n34559) );
  XNOR U33074 ( .A(n34562), .B(n34563), .Z(n34521) );
  ANDN U33075 ( .B(n34564), .A(n34565), .Z(n34562) );
  XOR U33076 ( .A(n34563), .B(n34566), .Z(n34564) );
  IV U33077 ( .A(n34520), .Z(n34554) );
  XOR U33078 ( .A(n34518), .B(n34567), .Z(n34520) );
  XOR U33079 ( .A(n34568), .B(n34569), .Z(n34567) );
  ANDN U33080 ( .B(n34570), .A(n34571), .Z(n34568) );
  XOR U33081 ( .A(n34572), .B(n34569), .Z(n34570) );
  IV U33082 ( .A(n34522), .Z(n34518) );
  XOR U33083 ( .A(n34573), .B(n34574), .Z(n34522) );
  ANDN U33084 ( .B(n34575), .A(n34576), .Z(n34573) );
  XOR U33085 ( .A(n34577), .B(n34574), .Z(n34575) );
  IV U33086 ( .A(n34532), .Z(n34536) );
  XOR U33087 ( .A(n34532), .B(n34487), .Z(n34534) );
  XOR U33088 ( .A(n34578), .B(n34579), .Z(n34487) );
  AND U33089 ( .A(n974), .B(n34580), .Z(n34578) );
  XOR U33090 ( .A(n34581), .B(n34579), .Z(n34580) );
  NANDN U33091 ( .A(n34489), .B(n34491), .Z(n34532) );
  XOR U33092 ( .A(n34582), .B(n34583), .Z(n34491) );
  AND U33093 ( .A(n974), .B(n34584), .Z(n34582) );
  XOR U33094 ( .A(n34583), .B(n34585), .Z(n34584) );
  XNOR U33095 ( .A(n34586), .B(n34587), .Z(n974) );
  AND U33096 ( .A(n34588), .B(n34589), .Z(n34586) );
  XOR U33097 ( .A(n34587), .B(n34502), .Z(n34589) );
  XNOR U33098 ( .A(n34590), .B(n34591), .Z(n34502) );
  ANDN U33099 ( .B(n34592), .A(n34593), .Z(n34590) );
  XOR U33100 ( .A(n34591), .B(n34594), .Z(n34592) );
  XNOR U33101 ( .A(n34587), .B(n34504), .Z(n34588) );
  XOR U33102 ( .A(n34595), .B(n34596), .Z(n34504) );
  AND U33103 ( .A(n978), .B(n34597), .Z(n34595) );
  XOR U33104 ( .A(n34598), .B(n34596), .Z(n34597) );
  XNOR U33105 ( .A(n34599), .B(n34600), .Z(n34587) );
  AND U33106 ( .A(n34601), .B(n34602), .Z(n34599) );
  XNOR U33107 ( .A(n34600), .B(n34529), .Z(n34602) );
  XOR U33108 ( .A(n34593), .B(n34594), .Z(n34529) );
  XNOR U33109 ( .A(n34603), .B(n34604), .Z(n34594) );
  ANDN U33110 ( .B(n34605), .A(n34606), .Z(n34603) );
  XOR U33111 ( .A(n34607), .B(n34608), .Z(n34605) );
  XOR U33112 ( .A(n34609), .B(n34610), .Z(n34593) );
  XNOR U33113 ( .A(n34611), .B(n34612), .Z(n34610) );
  ANDN U33114 ( .B(n34613), .A(n34614), .Z(n34611) );
  XNOR U33115 ( .A(n34615), .B(n34616), .Z(n34613) );
  IV U33116 ( .A(n34591), .Z(n34609) );
  XOR U33117 ( .A(n34617), .B(n34618), .Z(n34591) );
  ANDN U33118 ( .B(n34619), .A(n34620), .Z(n34617) );
  XOR U33119 ( .A(n34618), .B(n34621), .Z(n34619) );
  XOR U33120 ( .A(n34600), .B(n34531), .Z(n34601) );
  XOR U33121 ( .A(n34622), .B(n34623), .Z(n34531) );
  AND U33122 ( .A(n978), .B(n34624), .Z(n34622) );
  XOR U33123 ( .A(n34625), .B(n34623), .Z(n34624) );
  XNOR U33124 ( .A(n34626), .B(n34627), .Z(n34600) );
  NAND U33125 ( .A(n34628), .B(n34629), .Z(n34627) );
  XOR U33126 ( .A(n34630), .B(n34579), .Z(n34629) );
  XOR U33127 ( .A(n34620), .B(n34621), .Z(n34579) );
  XOR U33128 ( .A(n34631), .B(n34608), .Z(n34621) );
  XOR U33129 ( .A(n34632), .B(n34633), .Z(n34608) );
  ANDN U33130 ( .B(n34634), .A(n34635), .Z(n34632) );
  XOR U33131 ( .A(n34633), .B(n34636), .Z(n34634) );
  IV U33132 ( .A(n34606), .Z(n34631) );
  XOR U33133 ( .A(n34604), .B(n34637), .Z(n34606) );
  XOR U33134 ( .A(n34638), .B(n34639), .Z(n34637) );
  ANDN U33135 ( .B(n34640), .A(n34641), .Z(n34638) );
  XOR U33136 ( .A(n34642), .B(n34639), .Z(n34640) );
  IV U33137 ( .A(n34607), .Z(n34604) );
  XOR U33138 ( .A(n34643), .B(n34644), .Z(n34607) );
  ANDN U33139 ( .B(n34645), .A(n34646), .Z(n34643) );
  XOR U33140 ( .A(n34644), .B(n34647), .Z(n34645) );
  XOR U33141 ( .A(n34648), .B(n34649), .Z(n34620) );
  XNOR U33142 ( .A(n34615), .B(n34650), .Z(n34649) );
  IV U33143 ( .A(n34618), .Z(n34650) );
  XOR U33144 ( .A(n34651), .B(n34652), .Z(n34618) );
  ANDN U33145 ( .B(n34653), .A(n34654), .Z(n34651) );
  XOR U33146 ( .A(n34652), .B(n34655), .Z(n34653) );
  XNOR U33147 ( .A(n34656), .B(n34657), .Z(n34615) );
  ANDN U33148 ( .B(n34658), .A(n34659), .Z(n34656) );
  XOR U33149 ( .A(n34657), .B(n34660), .Z(n34658) );
  IV U33150 ( .A(n34614), .Z(n34648) );
  XOR U33151 ( .A(n34612), .B(n34661), .Z(n34614) );
  XOR U33152 ( .A(n34662), .B(n34663), .Z(n34661) );
  ANDN U33153 ( .B(n34664), .A(n34665), .Z(n34662) );
  XOR U33154 ( .A(n34666), .B(n34663), .Z(n34664) );
  IV U33155 ( .A(n34616), .Z(n34612) );
  XOR U33156 ( .A(n34667), .B(n34668), .Z(n34616) );
  ANDN U33157 ( .B(n34669), .A(n34670), .Z(n34667) );
  XOR U33158 ( .A(n34671), .B(n34668), .Z(n34669) );
  IV U33159 ( .A(n34626), .Z(n34630) );
  XOR U33160 ( .A(n34626), .B(n34581), .Z(n34628) );
  XOR U33161 ( .A(n34672), .B(n34673), .Z(n34581) );
  AND U33162 ( .A(n978), .B(n34674), .Z(n34672) );
  XOR U33163 ( .A(n34675), .B(n34673), .Z(n34674) );
  NANDN U33164 ( .A(n34583), .B(n34585), .Z(n34626) );
  XOR U33165 ( .A(n34676), .B(n34677), .Z(n34585) );
  AND U33166 ( .A(n978), .B(n34678), .Z(n34676) );
  XOR U33167 ( .A(n34677), .B(n34679), .Z(n34678) );
  XNOR U33168 ( .A(n34680), .B(n34681), .Z(n978) );
  AND U33169 ( .A(n34682), .B(n34683), .Z(n34680) );
  XOR U33170 ( .A(n34681), .B(n34596), .Z(n34683) );
  XNOR U33171 ( .A(n34684), .B(n34685), .Z(n34596) );
  ANDN U33172 ( .B(n34686), .A(n34687), .Z(n34684) );
  XOR U33173 ( .A(n34685), .B(n34688), .Z(n34686) );
  XNOR U33174 ( .A(n34681), .B(n34598), .Z(n34682) );
  XOR U33175 ( .A(n34689), .B(n34690), .Z(n34598) );
  AND U33176 ( .A(n982), .B(n34691), .Z(n34689) );
  XOR U33177 ( .A(n34692), .B(n34690), .Z(n34691) );
  XNOR U33178 ( .A(n34693), .B(n34694), .Z(n34681) );
  AND U33179 ( .A(n34695), .B(n34696), .Z(n34693) );
  XNOR U33180 ( .A(n34694), .B(n34623), .Z(n34696) );
  XOR U33181 ( .A(n34687), .B(n34688), .Z(n34623) );
  XNOR U33182 ( .A(n34697), .B(n34698), .Z(n34688) );
  ANDN U33183 ( .B(n34699), .A(n34700), .Z(n34697) );
  XOR U33184 ( .A(n34701), .B(n34702), .Z(n34699) );
  XOR U33185 ( .A(n34703), .B(n34704), .Z(n34687) );
  XNOR U33186 ( .A(n34705), .B(n34706), .Z(n34704) );
  ANDN U33187 ( .B(n34707), .A(n34708), .Z(n34705) );
  XNOR U33188 ( .A(n34709), .B(n34710), .Z(n34707) );
  IV U33189 ( .A(n34685), .Z(n34703) );
  XOR U33190 ( .A(n34711), .B(n34712), .Z(n34685) );
  ANDN U33191 ( .B(n34713), .A(n34714), .Z(n34711) );
  XOR U33192 ( .A(n34712), .B(n34715), .Z(n34713) );
  XOR U33193 ( .A(n34694), .B(n34625), .Z(n34695) );
  XOR U33194 ( .A(n34716), .B(n34717), .Z(n34625) );
  AND U33195 ( .A(n982), .B(n34718), .Z(n34716) );
  XOR U33196 ( .A(n34719), .B(n34717), .Z(n34718) );
  XNOR U33197 ( .A(n34720), .B(n34721), .Z(n34694) );
  NAND U33198 ( .A(n34722), .B(n34723), .Z(n34721) );
  XOR U33199 ( .A(n34724), .B(n34673), .Z(n34723) );
  XOR U33200 ( .A(n34714), .B(n34715), .Z(n34673) );
  XOR U33201 ( .A(n34725), .B(n34702), .Z(n34715) );
  XOR U33202 ( .A(n34726), .B(n34727), .Z(n34702) );
  ANDN U33203 ( .B(n34728), .A(n34729), .Z(n34726) );
  XOR U33204 ( .A(n34727), .B(n34730), .Z(n34728) );
  IV U33205 ( .A(n34700), .Z(n34725) );
  XOR U33206 ( .A(n34698), .B(n34731), .Z(n34700) );
  XOR U33207 ( .A(n34732), .B(n34733), .Z(n34731) );
  ANDN U33208 ( .B(n34734), .A(n34735), .Z(n34732) );
  XOR U33209 ( .A(n34736), .B(n34733), .Z(n34734) );
  IV U33210 ( .A(n34701), .Z(n34698) );
  XOR U33211 ( .A(n34737), .B(n34738), .Z(n34701) );
  ANDN U33212 ( .B(n34739), .A(n34740), .Z(n34737) );
  XOR U33213 ( .A(n34738), .B(n34741), .Z(n34739) );
  XOR U33214 ( .A(n34742), .B(n34743), .Z(n34714) );
  XNOR U33215 ( .A(n34709), .B(n34744), .Z(n34743) );
  IV U33216 ( .A(n34712), .Z(n34744) );
  XOR U33217 ( .A(n34745), .B(n34746), .Z(n34712) );
  ANDN U33218 ( .B(n34747), .A(n34748), .Z(n34745) );
  XOR U33219 ( .A(n34746), .B(n34749), .Z(n34747) );
  XNOR U33220 ( .A(n34750), .B(n34751), .Z(n34709) );
  ANDN U33221 ( .B(n34752), .A(n34753), .Z(n34750) );
  XOR U33222 ( .A(n34751), .B(n34754), .Z(n34752) );
  IV U33223 ( .A(n34708), .Z(n34742) );
  XOR U33224 ( .A(n34706), .B(n34755), .Z(n34708) );
  XOR U33225 ( .A(n34756), .B(n34757), .Z(n34755) );
  ANDN U33226 ( .B(n34758), .A(n34759), .Z(n34756) );
  XOR U33227 ( .A(n34760), .B(n34757), .Z(n34758) );
  IV U33228 ( .A(n34710), .Z(n34706) );
  XOR U33229 ( .A(n34761), .B(n34762), .Z(n34710) );
  ANDN U33230 ( .B(n34763), .A(n34764), .Z(n34761) );
  XOR U33231 ( .A(n34765), .B(n34762), .Z(n34763) );
  IV U33232 ( .A(n34720), .Z(n34724) );
  XOR U33233 ( .A(n34720), .B(n34675), .Z(n34722) );
  XOR U33234 ( .A(n34766), .B(n34767), .Z(n34675) );
  AND U33235 ( .A(n982), .B(n34768), .Z(n34766) );
  XOR U33236 ( .A(n34769), .B(n34767), .Z(n34768) );
  NANDN U33237 ( .A(n34677), .B(n34679), .Z(n34720) );
  XOR U33238 ( .A(n34770), .B(n34771), .Z(n34679) );
  AND U33239 ( .A(n982), .B(n34772), .Z(n34770) );
  XOR U33240 ( .A(n34771), .B(n34773), .Z(n34772) );
  XNOR U33241 ( .A(n34774), .B(n34775), .Z(n982) );
  AND U33242 ( .A(n34776), .B(n34777), .Z(n34774) );
  XOR U33243 ( .A(n34775), .B(n34690), .Z(n34777) );
  XNOR U33244 ( .A(n34778), .B(n34779), .Z(n34690) );
  ANDN U33245 ( .B(n34780), .A(n34781), .Z(n34778) );
  XOR U33246 ( .A(n34779), .B(n34782), .Z(n34780) );
  XNOR U33247 ( .A(n34775), .B(n34692), .Z(n34776) );
  XOR U33248 ( .A(n34783), .B(n34784), .Z(n34692) );
  AND U33249 ( .A(n986), .B(n34785), .Z(n34783) );
  XOR U33250 ( .A(n34786), .B(n34784), .Z(n34785) );
  XNOR U33251 ( .A(n34787), .B(n34788), .Z(n34775) );
  AND U33252 ( .A(n34789), .B(n34790), .Z(n34787) );
  XNOR U33253 ( .A(n34788), .B(n34717), .Z(n34790) );
  XOR U33254 ( .A(n34781), .B(n34782), .Z(n34717) );
  XNOR U33255 ( .A(n34791), .B(n34792), .Z(n34782) );
  ANDN U33256 ( .B(n34793), .A(n34794), .Z(n34791) );
  XOR U33257 ( .A(n34795), .B(n34796), .Z(n34793) );
  XOR U33258 ( .A(n34797), .B(n34798), .Z(n34781) );
  XNOR U33259 ( .A(n34799), .B(n34800), .Z(n34798) );
  ANDN U33260 ( .B(n34801), .A(n34802), .Z(n34799) );
  XNOR U33261 ( .A(n34803), .B(n34804), .Z(n34801) );
  IV U33262 ( .A(n34779), .Z(n34797) );
  XOR U33263 ( .A(n34805), .B(n34806), .Z(n34779) );
  ANDN U33264 ( .B(n34807), .A(n34808), .Z(n34805) );
  XOR U33265 ( .A(n34806), .B(n34809), .Z(n34807) );
  XOR U33266 ( .A(n34788), .B(n34719), .Z(n34789) );
  XOR U33267 ( .A(n34810), .B(n34811), .Z(n34719) );
  AND U33268 ( .A(n986), .B(n34812), .Z(n34810) );
  XOR U33269 ( .A(n34813), .B(n34811), .Z(n34812) );
  XNOR U33270 ( .A(n34814), .B(n34815), .Z(n34788) );
  NAND U33271 ( .A(n34816), .B(n34817), .Z(n34815) );
  XOR U33272 ( .A(n34818), .B(n34767), .Z(n34817) );
  XOR U33273 ( .A(n34808), .B(n34809), .Z(n34767) );
  XOR U33274 ( .A(n34819), .B(n34796), .Z(n34809) );
  XOR U33275 ( .A(n34820), .B(n34821), .Z(n34796) );
  ANDN U33276 ( .B(n34822), .A(n34823), .Z(n34820) );
  XOR U33277 ( .A(n34821), .B(n34824), .Z(n34822) );
  IV U33278 ( .A(n34794), .Z(n34819) );
  XOR U33279 ( .A(n34792), .B(n34825), .Z(n34794) );
  XOR U33280 ( .A(n34826), .B(n34827), .Z(n34825) );
  ANDN U33281 ( .B(n34828), .A(n34829), .Z(n34826) );
  XOR U33282 ( .A(n34830), .B(n34827), .Z(n34828) );
  IV U33283 ( .A(n34795), .Z(n34792) );
  XOR U33284 ( .A(n34831), .B(n34832), .Z(n34795) );
  ANDN U33285 ( .B(n34833), .A(n34834), .Z(n34831) );
  XOR U33286 ( .A(n34832), .B(n34835), .Z(n34833) );
  XOR U33287 ( .A(n34836), .B(n34837), .Z(n34808) );
  XNOR U33288 ( .A(n34803), .B(n34838), .Z(n34837) );
  IV U33289 ( .A(n34806), .Z(n34838) );
  XOR U33290 ( .A(n34839), .B(n34840), .Z(n34806) );
  ANDN U33291 ( .B(n34841), .A(n34842), .Z(n34839) );
  XOR U33292 ( .A(n34840), .B(n34843), .Z(n34841) );
  XNOR U33293 ( .A(n34844), .B(n34845), .Z(n34803) );
  ANDN U33294 ( .B(n34846), .A(n34847), .Z(n34844) );
  XOR U33295 ( .A(n34845), .B(n34848), .Z(n34846) );
  IV U33296 ( .A(n34802), .Z(n34836) );
  XOR U33297 ( .A(n34800), .B(n34849), .Z(n34802) );
  XOR U33298 ( .A(n34850), .B(n34851), .Z(n34849) );
  ANDN U33299 ( .B(n34852), .A(n34853), .Z(n34850) );
  XOR U33300 ( .A(n34854), .B(n34851), .Z(n34852) );
  IV U33301 ( .A(n34804), .Z(n34800) );
  XOR U33302 ( .A(n34855), .B(n34856), .Z(n34804) );
  ANDN U33303 ( .B(n34857), .A(n34858), .Z(n34855) );
  XOR U33304 ( .A(n34859), .B(n34856), .Z(n34857) );
  IV U33305 ( .A(n34814), .Z(n34818) );
  XOR U33306 ( .A(n34814), .B(n34769), .Z(n34816) );
  XOR U33307 ( .A(n34860), .B(n34861), .Z(n34769) );
  AND U33308 ( .A(n986), .B(n34862), .Z(n34860) );
  XOR U33309 ( .A(n34863), .B(n34861), .Z(n34862) );
  NANDN U33310 ( .A(n34771), .B(n34773), .Z(n34814) );
  XOR U33311 ( .A(n34864), .B(n34865), .Z(n34773) );
  AND U33312 ( .A(n986), .B(n34866), .Z(n34864) );
  XOR U33313 ( .A(n34865), .B(n34867), .Z(n34866) );
  XNOR U33314 ( .A(n34868), .B(n34869), .Z(n986) );
  AND U33315 ( .A(n34870), .B(n34871), .Z(n34868) );
  XOR U33316 ( .A(n34869), .B(n34784), .Z(n34871) );
  XNOR U33317 ( .A(n34872), .B(n34873), .Z(n34784) );
  ANDN U33318 ( .B(n34874), .A(n34875), .Z(n34872) );
  XOR U33319 ( .A(n34873), .B(n34876), .Z(n34874) );
  XNOR U33320 ( .A(n34869), .B(n34786), .Z(n34870) );
  XOR U33321 ( .A(n34877), .B(n34878), .Z(n34786) );
  AND U33322 ( .A(n990), .B(n34879), .Z(n34877) );
  XOR U33323 ( .A(n34880), .B(n34878), .Z(n34879) );
  XNOR U33324 ( .A(n34881), .B(n34882), .Z(n34869) );
  AND U33325 ( .A(n34883), .B(n34884), .Z(n34881) );
  XNOR U33326 ( .A(n34882), .B(n34811), .Z(n34884) );
  XOR U33327 ( .A(n34875), .B(n34876), .Z(n34811) );
  XNOR U33328 ( .A(n34885), .B(n34886), .Z(n34876) );
  ANDN U33329 ( .B(n34887), .A(n34888), .Z(n34885) );
  XOR U33330 ( .A(n34889), .B(n34890), .Z(n34887) );
  XOR U33331 ( .A(n34891), .B(n34892), .Z(n34875) );
  XNOR U33332 ( .A(n34893), .B(n34894), .Z(n34892) );
  ANDN U33333 ( .B(n34895), .A(n34896), .Z(n34893) );
  XNOR U33334 ( .A(n34897), .B(n34898), .Z(n34895) );
  IV U33335 ( .A(n34873), .Z(n34891) );
  XOR U33336 ( .A(n34899), .B(n34900), .Z(n34873) );
  ANDN U33337 ( .B(n34901), .A(n34902), .Z(n34899) );
  XOR U33338 ( .A(n34900), .B(n34903), .Z(n34901) );
  XOR U33339 ( .A(n34882), .B(n34813), .Z(n34883) );
  XOR U33340 ( .A(n34904), .B(n34905), .Z(n34813) );
  AND U33341 ( .A(n990), .B(n34906), .Z(n34904) );
  XOR U33342 ( .A(n34907), .B(n34905), .Z(n34906) );
  XNOR U33343 ( .A(n34908), .B(n34909), .Z(n34882) );
  NAND U33344 ( .A(n34910), .B(n34911), .Z(n34909) );
  XOR U33345 ( .A(n34912), .B(n34861), .Z(n34911) );
  XOR U33346 ( .A(n34902), .B(n34903), .Z(n34861) );
  XOR U33347 ( .A(n34913), .B(n34890), .Z(n34903) );
  XOR U33348 ( .A(n34914), .B(n34915), .Z(n34890) );
  ANDN U33349 ( .B(n34916), .A(n34917), .Z(n34914) );
  XOR U33350 ( .A(n34915), .B(n34918), .Z(n34916) );
  IV U33351 ( .A(n34888), .Z(n34913) );
  XOR U33352 ( .A(n34886), .B(n34919), .Z(n34888) );
  XOR U33353 ( .A(n34920), .B(n34921), .Z(n34919) );
  ANDN U33354 ( .B(n34922), .A(n34923), .Z(n34920) );
  XOR U33355 ( .A(n34924), .B(n34921), .Z(n34922) );
  IV U33356 ( .A(n34889), .Z(n34886) );
  XOR U33357 ( .A(n34925), .B(n34926), .Z(n34889) );
  ANDN U33358 ( .B(n34927), .A(n34928), .Z(n34925) );
  XOR U33359 ( .A(n34926), .B(n34929), .Z(n34927) );
  XOR U33360 ( .A(n34930), .B(n34931), .Z(n34902) );
  XNOR U33361 ( .A(n34897), .B(n34932), .Z(n34931) );
  IV U33362 ( .A(n34900), .Z(n34932) );
  XOR U33363 ( .A(n34933), .B(n34934), .Z(n34900) );
  ANDN U33364 ( .B(n34935), .A(n34936), .Z(n34933) );
  XOR U33365 ( .A(n34934), .B(n34937), .Z(n34935) );
  XNOR U33366 ( .A(n34938), .B(n34939), .Z(n34897) );
  ANDN U33367 ( .B(n34940), .A(n34941), .Z(n34938) );
  XOR U33368 ( .A(n34939), .B(n34942), .Z(n34940) );
  IV U33369 ( .A(n34896), .Z(n34930) );
  XOR U33370 ( .A(n34894), .B(n34943), .Z(n34896) );
  XOR U33371 ( .A(n34944), .B(n34945), .Z(n34943) );
  ANDN U33372 ( .B(n34946), .A(n34947), .Z(n34944) );
  XOR U33373 ( .A(n34948), .B(n34945), .Z(n34946) );
  IV U33374 ( .A(n34898), .Z(n34894) );
  XOR U33375 ( .A(n34949), .B(n34950), .Z(n34898) );
  ANDN U33376 ( .B(n34951), .A(n34952), .Z(n34949) );
  XOR U33377 ( .A(n34953), .B(n34950), .Z(n34951) );
  IV U33378 ( .A(n34908), .Z(n34912) );
  XOR U33379 ( .A(n34908), .B(n34863), .Z(n34910) );
  XOR U33380 ( .A(n34954), .B(n34955), .Z(n34863) );
  AND U33381 ( .A(n990), .B(n34956), .Z(n34954) );
  XOR U33382 ( .A(n34957), .B(n34955), .Z(n34956) );
  NANDN U33383 ( .A(n34865), .B(n34867), .Z(n34908) );
  XOR U33384 ( .A(n34958), .B(n34959), .Z(n34867) );
  AND U33385 ( .A(n990), .B(n34960), .Z(n34958) );
  XOR U33386 ( .A(n34959), .B(n34961), .Z(n34960) );
  XNOR U33387 ( .A(n34962), .B(n34963), .Z(n990) );
  AND U33388 ( .A(n34964), .B(n34965), .Z(n34962) );
  XOR U33389 ( .A(n34963), .B(n34878), .Z(n34965) );
  XNOR U33390 ( .A(n34966), .B(n34967), .Z(n34878) );
  ANDN U33391 ( .B(n34968), .A(n34969), .Z(n34966) );
  XOR U33392 ( .A(n34967), .B(n34970), .Z(n34968) );
  XNOR U33393 ( .A(n34963), .B(n34880), .Z(n34964) );
  XOR U33394 ( .A(n34971), .B(n34972), .Z(n34880) );
  AND U33395 ( .A(n994), .B(n34973), .Z(n34971) );
  XOR U33396 ( .A(n34974), .B(n34972), .Z(n34973) );
  XNOR U33397 ( .A(n34975), .B(n34976), .Z(n34963) );
  AND U33398 ( .A(n34977), .B(n34978), .Z(n34975) );
  XNOR U33399 ( .A(n34976), .B(n34905), .Z(n34978) );
  XOR U33400 ( .A(n34969), .B(n34970), .Z(n34905) );
  XNOR U33401 ( .A(n34979), .B(n34980), .Z(n34970) );
  ANDN U33402 ( .B(n34981), .A(n34982), .Z(n34979) );
  XOR U33403 ( .A(n34983), .B(n34984), .Z(n34981) );
  XOR U33404 ( .A(n34985), .B(n34986), .Z(n34969) );
  XNOR U33405 ( .A(n34987), .B(n34988), .Z(n34986) );
  ANDN U33406 ( .B(n34989), .A(n34990), .Z(n34987) );
  XNOR U33407 ( .A(n34991), .B(n34992), .Z(n34989) );
  IV U33408 ( .A(n34967), .Z(n34985) );
  XOR U33409 ( .A(n34993), .B(n34994), .Z(n34967) );
  ANDN U33410 ( .B(n34995), .A(n34996), .Z(n34993) );
  XOR U33411 ( .A(n34994), .B(n34997), .Z(n34995) );
  XOR U33412 ( .A(n34976), .B(n34907), .Z(n34977) );
  XOR U33413 ( .A(n34998), .B(n34999), .Z(n34907) );
  AND U33414 ( .A(n994), .B(n35000), .Z(n34998) );
  XOR U33415 ( .A(n35001), .B(n34999), .Z(n35000) );
  XNOR U33416 ( .A(n35002), .B(n35003), .Z(n34976) );
  NAND U33417 ( .A(n35004), .B(n35005), .Z(n35003) );
  XOR U33418 ( .A(n35006), .B(n34955), .Z(n35005) );
  XOR U33419 ( .A(n34996), .B(n34997), .Z(n34955) );
  XOR U33420 ( .A(n35007), .B(n34984), .Z(n34997) );
  XOR U33421 ( .A(n35008), .B(n35009), .Z(n34984) );
  ANDN U33422 ( .B(n35010), .A(n35011), .Z(n35008) );
  XOR U33423 ( .A(n35009), .B(n35012), .Z(n35010) );
  IV U33424 ( .A(n34982), .Z(n35007) );
  XOR U33425 ( .A(n34980), .B(n35013), .Z(n34982) );
  XOR U33426 ( .A(n35014), .B(n35015), .Z(n35013) );
  ANDN U33427 ( .B(n35016), .A(n35017), .Z(n35014) );
  XOR U33428 ( .A(n35018), .B(n35015), .Z(n35016) );
  IV U33429 ( .A(n34983), .Z(n34980) );
  XOR U33430 ( .A(n35019), .B(n35020), .Z(n34983) );
  ANDN U33431 ( .B(n35021), .A(n35022), .Z(n35019) );
  XOR U33432 ( .A(n35020), .B(n35023), .Z(n35021) );
  XOR U33433 ( .A(n35024), .B(n35025), .Z(n34996) );
  XNOR U33434 ( .A(n34991), .B(n35026), .Z(n35025) );
  IV U33435 ( .A(n34994), .Z(n35026) );
  XOR U33436 ( .A(n35027), .B(n35028), .Z(n34994) );
  ANDN U33437 ( .B(n35029), .A(n35030), .Z(n35027) );
  XOR U33438 ( .A(n35028), .B(n35031), .Z(n35029) );
  XNOR U33439 ( .A(n35032), .B(n35033), .Z(n34991) );
  ANDN U33440 ( .B(n35034), .A(n35035), .Z(n35032) );
  XOR U33441 ( .A(n35033), .B(n35036), .Z(n35034) );
  IV U33442 ( .A(n34990), .Z(n35024) );
  XOR U33443 ( .A(n34988), .B(n35037), .Z(n34990) );
  XOR U33444 ( .A(n35038), .B(n35039), .Z(n35037) );
  ANDN U33445 ( .B(n35040), .A(n35041), .Z(n35038) );
  XOR U33446 ( .A(n35042), .B(n35039), .Z(n35040) );
  IV U33447 ( .A(n34992), .Z(n34988) );
  XOR U33448 ( .A(n35043), .B(n35044), .Z(n34992) );
  ANDN U33449 ( .B(n35045), .A(n35046), .Z(n35043) );
  XOR U33450 ( .A(n35047), .B(n35044), .Z(n35045) );
  IV U33451 ( .A(n35002), .Z(n35006) );
  XOR U33452 ( .A(n35002), .B(n34957), .Z(n35004) );
  XOR U33453 ( .A(n35048), .B(n35049), .Z(n34957) );
  AND U33454 ( .A(n994), .B(n35050), .Z(n35048) );
  XOR U33455 ( .A(n35051), .B(n35049), .Z(n35050) );
  NANDN U33456 ( .A(n34959), .B(n34961), .Z(n35002) );
  XOR U33457 ( .A(n35052), .B(n35053), .Z(n34961) );
  AND U33458 ( .A(n994), .B(n35054), .Z(n35052) );
  XOR U33459 ( .A(n35053), .B(n35055), .Z(n35054) );
  XNOR U33460 ( .A(n35056), .B(n35057), .Z(n994) );
  AND U33461 ( .A(n35058), .B(n35059), .Z(n35056) );
  XOR U33462 ( .A(n35057), .B(n34972), .Z(n35059) );
  XNOR U33463 ( .A(n35060), .B(n35061), .Z(n34972) );
  ANDN U33464 ( .B(n35062), .A(n35063), .Z(n35060) );
  XOR U33465 ( .A(n35061), .B(n35064), .Z(n35062) );
  XNOR U33466 ( .A(n35057), .B(n34974), .Z(n35058) );
  XOR U33467 ( .A(n35065), .B(n35066), .Z(n34974) );
  AND U33468 ( .A(n998), .B(n35067), .Z(n35065) );
  XOR U33469 ( .A(n35068), .B(n35066), .Z(n35067) );
  XNOR U33470 ( .A(n35069), .B(n35070), .Z(n35057) );
  AND U33471 ( .A(n35071), .B(n35072), .Z(n35069) );
  XNOR U33472 ( .A(n35070), .B(n34999), .Z(n35072) );
  XOR U33473 ( .A(n35063), .B(n35064), .Z(n34999) );
  XNOR U33474 ( .A(n35073), .B(n35074), .Z(n35064) );
  ANDN U33475 ( .B(n35075), .A(n35076), .Z(n35073) );
  XOR U33476 ( .A(n35077), .B(n35078), .Z(n35075) );
  XOR U33477 ( .A(n35079), .B(n35080), .Z(n35063) );
  XNOR U33478 ( .A(n35081), .B(n35082), .Z(n35080) );
  ANDN U33479 ( .B(n35083), .A(n35084), .Z(n35081) );
  XNOR U33480 ( .A(n35085), .B(n35086), .Z(n35083) );
  IV U33481 ( .A(n35061), .Z(n35079) );
  XOR U33482 ( .A(n35087), .B(n35088), .Z(n35061) );
  ANDN U33483 ( .B(n35089), .A(n35090), .Z(n35087) );
  XOR U33484 ( .A(n35088), .B(n35091), .Z(n35089) );
  XOR U33485 ( .A(n35070), .B(n35001), .Z(n35071) );
  XOR U33486 ( .A(n35092), .B(n35093), .Z(n35001) );
  AND U33487 ( .A(n998), .B(n35094), .Z(n35092) );
  XOR U33488 ( .A(n35095), .B(n35093), .Z(n35094) );
  XNOR U33489 ( .A(n35096), .B(n35097), .Z(n35070) );
  NAND U33490 ( .A(n35098), .B(n35099), .Z(n35097) );
  XOR U33491 ( .A(n35100), .B(n35049), .Z(n35099) );
  XOR U33492 ( .A(n35090), .B(n35091), .Z(n35049) );
  XOR U33493 ( .A(n35101), .B(n35078), .Z(n35091) );
  XOR U33494 ( .A(n35102), .B(n35103), .Z(n35078) );
  ANDN U33495 ( .B(n35104), .A(n35105), .Z(n35102) );
  XOR U33496 ( .A(n35103), .B(n35106), .Z(n35104) );
  IV U33497 ( .A(n35076), .Z(n35101) );
  XOR U33498 ( .A(n35074), .B(n35107), .Z(n35076) );
  XOR U33499 ( .A(n35108), .B(n35109), .Z(n35107) );
  ANDN U33500 ( .B(n35110), .A(n35111), .Z(n35108) );
  XOR U33501 ( .A(n35112), .B(n35109), .Z(n35110) );
  IV U33502 ( .A(n35077), .Z(n35074) );
  XOR U33503 ( .A(n35113), .B(n35114), .Z(n35077) );
  ANDN U33504 ( .B(n35115), .A(n35116), .Z(n35113) );
  XOR U33505 ( .A(n35114), .B(n35117), .Z(n35115) );
  XOR U33506 ( .A(n35118), .B(n35119), .Z(n35090) );
  XNOR U33507 ( .A(n35085), .B(n35120), .Z(n35119) );
  IV U33508 ( .A(n35088), .Z(n35120) );
  XOR U33509 ( .A(n35121), .B(n35122), .Z(n35088) );
  ANDN U33510 ( .B(n35123), .A(n35124), .Z(n35121) );
  XOR U33511 ( .A(n35122), .B(n35125), .Z(n35123) );
  XNOR U33512 ( .A(n35126), .B(n35127), .Z(n35085) );
  ANDN U33513 ( .B(n35128), .A(n35129), .Z(n35126) );
  XOR U33514 ( .A(n35127), .B(n35130), .Z(n35128) );
  IV U33515 ( .A(n35084), .Z(n35118) );
  XOR U33516 ( .A(n35082), .B(n35131), .Z(n35084) );
  XOR U33517 ( .A(n35132), .B(n35133), .Z(n35131) );
  ANDN U33518 ( .B(n35134), .A(n35135), .Z(n35132) );
  XOR U33519 ( .A(n35136), .B(n35133), .Z(n35134) );
  IV U33520 ( .A(n35086), .Z(n35082) );
  XOR U33521 ( .A(n35137), .B(n35138), .Z(n35086) );
  ANDN U33522 ( .B(n35139), .A(n35140), .Z(n35137) );
  XOR U33523 ( .A(n35141), .B(n35138), .Z(n35139) );
  IV U33524 ( .A(n35096), .Z(n35100) );
  XOR U33525 ( .A(n35096), .B(n35051), .Z(n35098) );
  XOR U33526 ( .A(n35142), .B(n35143), .Z(n35051) );
  AND U33527 ( .A(n998), .B(n35144), .Z(n35142) );
  XOR U33528 ( .A(n35145), .B(n35143), .Z(n35144) );
  NANDN U33529 ( .A(n35053), .B(n35055), .Z(n35096) );
  XOR U33530 ( .A(n35146), .B(n35147), .Z(n35055) );
  AND U33531 ( .A(n998), .B(n35148), .Z(n35146) );
  XOR U33532 ( .A(n35147), .B(n35149), .Z(n35148) );
  XNOR U33533 ( .A(n35150), .B(n35151), .Z(n998) );
  AND U33534 ( .A(n35152), .B(n35153), .Z(n35150) );
  XOR U33535 ( .A(n35151), .B(n35066), .Z(n35153) );
  XNOR U33536 ( .A(n35154), .B(n35155), .Z(n35066) );
  ANDN U33537 ( .B(n35156), .A(n35157), .Z(n35154) );
  XOR U33538 ( .A(n35155), .B(n35158), .Z(n35156) );
  XNOR U33539 ( .A(n35151), .B(n35068), .Z(n35152) );
  XOR U33540 ( .A(n35159), .B(n35160), .Z(n35068) );
  AND U33541 ( .A(n1002), .B(n35161), .Z(n35159) );
  XOR U33542 ( .A(n35162), .B(n35160), .Z(n35161) );
  XNOR U33543 ( .A(n35163), .B(n35164), .Z(n35151) );
  AND U33544 ( .A(n35165), .B(n35166), .Z(n35163) );
  XNOR U33545 ( .A(n35164), .B(n35093), .Z(n35166) );
  XOR U33546 ( .A(n35157), .B(n35158), .Z(n35093) );
  XNOR U33547 ( .A(n35167), .B(n35168), .Z(n35158) );
  ANDN U33548 ( .B(n35169), .A(n35170), .Z(n35167) );
  XOR U33549 ( .A(n35171), .B(n35172), .Z(n35169) );
  XOR U33550 ( .A(n35173), .B(n35174), .Z(n35157) );
  XNOR U33551 ( .A(n35175), .B(n35176), .Z(n35174) );
  ANDN U33552 ( .B(n35177), .A(n35178), .Z(n35175) );
  XNOR U33553 ( .A(n35179), .B(n35180), .Z(n35177) );
  IV U33554 ( .A(n35155), .Z(n35173) );
  XOR U33555 ( .A(n35181), .B(n35182), .Z(n35155) );
  ANDN U33556 ( .B(n35183), .A(n35184), .Z(n35181) );
  XOR U33557 ( .A(n35182), .B(n35185), .Z(n35183) );
  XOR U33558 ( .A(n35164), .B(n35095), .Z(n35165) );
  XOR U33559 ( .A(n35186), .B(n35187), .Z(n35095) );
  AND U33560 ( .A(n1002), .B(n35188), .Z(n35186) );
  XOR U33561 ( .A(n35189), .B(n35187), .Z(n35188) );
  XNOR U33562 ( .A(n35190), .B(n35191), .Z(n35164) );
  NAND U33563 ( .A(n35192), .B(n35193), .Z(n35191) );
  XOR U33564 ( .A(n35194), .B(n35143), .Z(n35193) );
  XOR U33565 ( .A(n35184), .B(n35185), .Z(n35143) );
  XOR U33566 ( .A(n35195), .B(n35172), .Z(n35185) );
  XOR U33567 ( .A(n35196), .B(n35197), .Z(n35172) );
  ANDN U33568 ( .B(n35198), .A(n35199), .Z(n35196) );
  XOR U33569 ( .A(n35197), .B(n35200), .Z(n35198) );
  IV U33570 ( .A(n35170), .Z(n35195) );
  XOR U33571 ( .A(n35168), .B(n35201), .Z(n35170) );
  XOR U33572 ( .A(n35202), .B(n35203), .Z(n35201) );
  ANDN U33573 ( .B(n35204), .A(n35205), .Z(n35202) );
  XOR U33574 ( .A(n35206), .B(n35203), .Z(n35204) );
  IV U33575 ( .A(n35171), .Z(n35168) );
  XOR U33576 ( .A(n35207), .B(n35208), .Z(n35171) );
  ANDN U33577 ( .B(n35209), .A(n35210), .Z(n35207) );
  XOR U33578 ( .A(n35208), .B(n35211), .Z(n35209) );
  XOR U33579 ( .A(n35212), .B(n35213), .Z(n35184) );
  XNOR U33580 ( .A(n35179), .B(n35214), .Z(n35213) );
  IV U33581 ( .A(n35182), .Z(n35214) );
  XOR U33582 ( .A(n35215), .B(n35216), .Z(n35182) );
  ANDN U33583 ( .B(n35217), .A(n35218), .Z(n35215) );
  XOR U33584 ( .A(n35216), .B(n35219), .Z(n35217) );
  XNOR U33585 ( .A(n35220), .B(n35221), .Z(n35179) );
  ANDN U33586 ( .B(n35222), .A(n35223), .Z(n35220) );
  XOR U33587 ( .A(n35221), .B(n35224), .Z(n35222) );
  IV U33588 ( .A(n35178), .Z(n35212) );
  XOR U33589 ( .A(n35176), .B(n35225), .Z(n35178) );
  XOR U33590 ( .A(n35226), .B(n35227), .Z(n35225) );
  ANDN U33591 ( .B(n35228), .A(n35229), .Z(n35226) );
  XOR U33592 ( .A(n35230), .B(n35227), .Z(n35228) );
  IV U33593 ( .A(n35180), .Z(n35176) );
  XOR U33594 ( .A(n35231), .B(n35232), .Z(n35180) );
  ANDN U33595 ( .B(n35233), .A(n35234), .Z(n35231) );
  XOR U33596 ( .A(n35235), .B(n35232), .Z(n35233) );
  IV U33597 ( .A(n35190), .Z(n35194) );
  XOR U33598 ( .A(n35190), .B(n35145), .Z(n35192) );
  XOR U33599 ( .A(n35236), .B(n35237), .Z(n35145) );
  AND U33600 ( .A(n1002), .B(n35238), .Z(n35236) );
  XOR U33601 ( .A(n35239), .B(n35237), .Z(n35238) );
  NANDN U33602 ( .A(n35147), .B(n35149), .Z(n35190) );
  XOR U33603 ( .A(n35240), .B(n35241), .Z(n35149) );
  AND U33604 ( .A(n1002), .B(n35242), .Z(n35240) );
  XOR U33605 ( .A(n35241), .B(n35243), .Z(n35242) );
  XNOR U33606 ( .A(n35244), .B(n35245), .Z(n1002) );
  AND U33607 ( .A(n35246), .B(n35247), .Z(n35244) );
  XOR U33608 ( .A(n35245), .B(n35160), .Z(n35247) );
  XNOR U33609 ( .A(n35248), .B(n35249), .Z(n35160) );
  ANDN U33610 ( .B(n35250), .A(n35251), .Z(n35248) );
  XOR U33611 ( .A(n35249), .B(n35252), .Z(n35250) );
  XNOR U33612 ( .A(n35245), .B(n35162), .Z(n35246) );
  XOR U33613 ( .A(n35253), .B(n35254), .Z(n35162) );
  AND U33614 ( .A(n1006), .B(n35255), .Z(n35253) );
  XOR U33615 ( .A(n35256), .B(n35254), .Z(n35255) );
  XNOR U33616 ( .A(n35257), .B(n35258), .Z(n35245) );
  AND U33617 ( .A(n35259), .B(n35260), .Z(n35257) );
  XNOR U33618 ( .A(n35258), .B(n35187), .Z(n35260) );
  XOR U33619 ( .A(n35251), .B(n35252), .Z(n35187) );
  XNOR U33620 ( .A(n35261), .B(n35262), .Z(n35252) );
  ANDN U33621 ( .B(n35263), .A(n35264), .Z(n35261) );
  XOR U33622 ( .A(n35265), .B(n35266), .Z(n35263) );
  XOR U33623 ( .A(n35267), .B(n35268), .Z(n35251) );
  XNOR U33624 ( .A(n35269), .B(n35270), .Z(n35268) );
  ANDN U33625 ( .B(n35271), .A(n35272), .Z(n35269) );
  XNOR U33626 ( .A(n35273), .B(n35274), .Z(n35271) );
  IV U33627 ( .A(n35249), .Z(n35267) );
  XOR U33628 ( .A(n35275), .B(n35276), .Z(n35249) );
  ANDN U33629 ( .B(n35277), .A(n35278), .Z(n35275) );
  XOR U33630 ( .A(n35276), .B(n35279), .Z(n35277) );
  XOR U33631 ( .A(n35258), .B(n35189), .Z(n35259) );
  XOR U33632 ( .A(n35280), .B(n35281), .Z(n35189) );
  AND U33633 ( .A(n1006), .B(n35282), .Z(n35280) );
  XOR U33634 ( .A(n35283), .B(n35281), .Z(n35282) );
  XNOR U33635 ( .A(n35284), .B(n35285), .Z(n35258) );
  NAND U33636 ( .A(n35286), .B(n35287), .Z(n35285) );
  XOR U33637 ( .A(n35288), .B(n35237), .Z(n35287) );
  XOR U33638 ( .A(n35278), .B(n35279), .Z(n35237) );
  XOR U33639 ( .A(n35289), .B(n35266), .Z(n35279) );
  XOR U33640 ( .A(n35290), .B(n35291), .Z(n35266) );
  ANDN U33641 ( .B(n35292), .A(n35293), .Z(n35290) );
  XOR U33642 ( .A(n35291), .B(n35294), .Z(n35292) );
  IV U33643 ( .A(n35264), .Z(n35289) );
  XOR U33644 ( .A(n35262), .B(n35295), .Z(n35264) );
  XOR U33645 ( .A(n35296), .B(n35297), .Z(n35295) );
  ANDN U33646 ( .B(n35298), .A(n35299), .Z(n35296) );
  XOR U33647 ( .A(n35300), .B(n35297), .Z(n35298) );
  IV U33648 ( .A(n35265), .Z(n35262) );
  XOR U33649 ( .A(n35301), .B(n35302), .Z(n35265) );
  ANDN U33650 ( .B(n35303), .A(n35304), .Z(n35301) );
  XOR U33651 ( .A(n35302), .B(n35305), .Z(n35303) );
  XOR U33652 ( .A(n35306), .B(n35307), .Z(n35278) );
  XNOR U33653 ( .A(n35273), .B(n35308), .Z(n35307) );
  IV U33654 ( .A(n35276), .Z(n35308) );
  XOR U33655 ( .A(n35309), .B(n35310), .Z(n35276) );
  ANDN U33656 ( .B(n35311), .A(n35312), .Z(n35309) );
  XOR U33657 ( .A(n35310), .B(n35313), .Z(n35311) );
  XNOR U33658 ( .A(n35314), .B(n35315), .Z(n35273) );
  ANDN U33659 ( .B(n35316), .A(n35317), .Z(n35314) );
  XOR U33660 ( .A(n35315), .B(n35318), .Z(n35316) );
  IV U33661 ( .A(n35272), .Z(n35306) );
  XOR U33662 ( .A(n35270), .B(n35319), .Z(n35272) );
  XOR U33663 ( .A(n35320), .B(n35321), .Z(n35319) );
  ANDN U33664 ( .B(n35322), .A(n35323), .Z(n35320) );
  XOR U33665 ( .A(n35324), .B(n35321), .Z(n35322) );
  IV U33666 ( .A(n35274), .Z(n35270) );
  XOR U33667 ( .A(n35325), .B(n35326), .Z(n35274) );
  ANDN U33668 ( .B(n35327), .A(n35328), .Z(n35325) );
  XOR U33669 ( .A(n35329), .B(n35326), .Z(n35327) );
  IV U33670 ( .A(n35284), .Z(n35288) );
  XOR U33671 ( .A(n35284), .B(n35239), .Z(n35286) );
  XOR U33672 ( .A(n35330), .B(n35331), .Z(n35239) );
  AND U33673 ( .A(n1006), .B(n35332), .Z(n35330) );
  XOR U33674 ( .A(n35333), .B(n35331), .Z(n35332) );
  NANDN U33675 ( .A(n35241), .B(n35243), .Z(n35284) );
  XOR U33676 ( .A(n35334), .B(n35335), .Z(n35243) );
  AND U33677 ( .A(n1006), .B(n35336), .Z(n35334) );
  XOR U33678 ( .A(n35335), .B(n35337), .Z(n35336) );
  XNOR U33679 ( .A(n35338), .B(n35339), .Z(n1006) );
  AND U33680 ( .A(n35340), .B(n35341), .Z(n35338) );
  XOR U33681 ( .A(n35339), .B(n35254), .Z(n35341) );
  XNOR U33682 ( .A(n35342), .B(n35343), .Z(n35254) );
  ANDN U33683 ( .B(n35344), .A(n35345), .Z(n35342) );
  XOR U33684 ( .A(n35343), .B(n35346), .Z(n35344) );
  XNOR U33685 ( .A(n35339), .B(n35256), .Z(n35340) );
  XOR U33686 ( .A(n35347), .B(n35348), .Z(n35256) );
  AND U33687 ( .A(n1010), .B(n35349), .Z(n35347) );
  XOR U33688 ( .A(n35350), .B(n35348), .Z(n35349) );
  XNOR U33689 ( .A(n35351), .B(n35352), .Z(n35339) );
  AND U33690 ( .A(n35353), .B(n35354), .Z(n35351) );
  XNOR U33691 ( .A(n35352), .B(n35281), .Z(n35354) );
  XOR U33692 ( .A(n35345), .B(n35346), .Z(n35281) );
  XNOR U33693 ( .A(n35355), .B(n35356), .Z(n35346) );
  ANDN U33694 ( .B(n35357), .A(n35358), .Z(n35355) );
  XOR U33695 ( .A(n35359), .B(n35360), .Z(n35357) );
  XOR U33696 ( .A(n35361), .B(n35362), .Z(n35345) );
  XNOR U33697 ( .A(n35363), .B(n35364), .Z(n35362) );
  ANDN U33698 ( .B(n35365), .A(n35366), .Z(n35363) );
  XNOR U33699 ( .A(n35367), .B(n35368), .Z(n35365) );
  IV U33700 ( .A(n35343), .Z(n35361) );
  XOR U33701 ( .A(n35369), .B(n35370), .Z(n35343) );
  ANDN U33702 ( .B(n35371), .A(n35372), .Z(n35369) );
  XOR U33703 ( .A(n35370), .B(n35373), .Z(n35371) );
  XOR U33704 ( .A(n35352), .B(n35283), .Z(n35353) );
  XOR U33705 ( .A(n35374), .B(n35375), .Z(n35283) );
  AND U33706 ( .A(n1010), .B(n35376), .Z(n35374) );
  XOR U33707 ( .A(n35377), .B(n35375), .Z(n35376) );
  XNOR U33708 ( .A(n35378), .B(n35379), .Z(n35352) );
  NAND U33709 ( .A(n35380), .B(n35381), .Z(n35379) );
  XOR U33710 ( .A(n35382), .B(n35331), .Z(n35381) );
  XOR U33711 ( .A(n35372), .B(n35373), .Z(n35331) );
  XOR U33712 ( .A(n35383), .B(n35360), .Z(n35373) );
  XOR U33713 ( .A(n35384), .B(n35385), .Z(n35360) );
  ANDN U33714 ( .B(n35386), .A(n35387), .Z(n35384) );
  XOR U33715 ( .A(n35385), .B(n35388), .Z(n35386) );
  IV U33716 ( .A(n35358), .Z(n35383) );
  XOR U33717 ( .A(n35356), .B(n35389), .Z(n35358) );
  XOR U33718 ( .A(n35390), .B(n35391), .Z(n35389) );
  ANDN U33719 ( .B(n35392), .A(n35393), .Z(n35390) );
  XOR U33720 ( .A(n35394), .B(n35391), .Z(n35392) );
  IV U33721 ( .A(n35359), .Z(n35356) );
  XOR U33722 ( .A(n35395), .B(n35396), .Z(n35359) );
  ANDN U33723 ( .B(n35397), .A(n35398), .Z(n35395) );
  XOR U33724 ( .A(n35396), .B(n35399), .Z(n35397) );
  XOR U33725 ( .A(n35400), .B(n35401), .Z(n35372) );
  XNOR U33726 ( .A(n35367), .B(n35402), .Z(n35401) );
  IV U33727 ( .A(n35370), .Z(n35402) );
  XOR U33728 ( .A(n35403), .B(n35404), .Z(n35370) );
  ANDN U33729 ( .B(n35405), .A(n35406), .Z(n35403) );
  XOR U33730 ( .A(n35404), .B(n35407), .Z(n35405) );
  XNOR U33731 ( .A(n35408), .B(n35409), .Z(n35367) );
  ANDN U33732 ( .B(n35410), .A(n35411), .Z(n35408) );
  XOR U33733 ( .A(n35409), .B(n35412), .Z(n35410) );
  IV U33734 ( .A(n35366), .Z(n35400) );
  XOR U33735 ( .A(n35364), .B(n35413), .Z(n35366) );
  XOR U33736 ( .A(n35414), .B(n35415), .Z(n35413) );
  ANDN U33737 ( .B(n35416), .A(n35417), .Z(n35414) );
  XOR U33738 ( .A(n35418), .B(n35415), .Z(n35416) );
  IV U33739 ( .A(n35368), .Z(n35364) );
  XOR U33740 ( .A(n35419), .B(n35420), .Z(n35368) );
  ANDN U33741 ( .B(n35421), .A(n35422), .Z(n35419) );
  XOR U33742 ( .A(n35423), .B(n35420), .Z(n35421) );
  IV U33743 ( .A(n35378), .Z(n35382) );
  XOR U33744 ( .A(n35378), .B(n35333), .Z(n35380) );
  XOR U33745 ( .A(n35424), .B(n35425), .Z(n35333) );
  AND U33746 ( .A(n1010), .B(n35426), .Z(n35424) );
  XOR U33747 ( .A(n35427), .B(n35425), .Z(n35426) );
  NANDN U33748 ( .A(n35335), .B(n35337), .Z(n35378) );
  XOR U33749 ( .A(n35428), .B(n35429), .Z(n35337) );
  AND U33750 ( .A(n1010), .B(n35430), .Z(n35428) );
  XOR U33751 ( .A(n35429), .B(n35431), .Z(n35430) );
  XNOR U33752 ( .A(n35432), .B(n35433), .Z(n1010) );
  AND U33753 ( .A(n35434), .B(n35435), .Z(n35432) );
  XOR U33754 ( .A(n35433), .B(n35348), .Z(n35435) );
  XNOR U33755 ( .A(n35436), .B(n35437), .Z(n35348) );
  ANDN U33756 ( .B(n35438), .A(n35439), .Z(n35436) );
  XOR U33757 ( .A(n35437), .B(n35440), .Z(n35438) );
  XNOR U33758 ( .A(n35433), .B(n35350), .Z(n35434) );
  XOR U33759 ( .A(n35441), .B(n35442), .Z(n35350) );
  AND U33760 ( .A(n1014), .B(n35443), .Z(n35441) );
  XOR U33761 ( .A(n35444), .B(n35442), .Z(n35443) );
  XNOR U33762 ( .A(n35445), .B(n35446), .Z(n35433) );
  AND U33763 ( .A(n35447), .B(n35448), .Z(n35445) );
  XNOR U33764 ( .A(n35446), .B(n35375), .Z(n35448) );
  XOR U33765 ( .A(n35439), .B(n35440), .Z(n35375) );
  XNOR U33766 ( .A(n35449), .B(n35450), .Z(n35440) );
  ANDN U33767 ( .B(n35451), .A(n35452), .Z(n35449) );
  XOR U33768 ( .A(n35453), .B(n35454), .Z(n35451) );
  XOR U33769 ( .A(n35455), .B(n35456), .Z(n35439) );
  XNOR U33770 ( .A(n35457), .B(n35458), .Z(n35456) );
  ANDN U33771 ( .B(n35459), .A(n35460), .Z(n35457) );
  XNOR U33772 ( .A(n35461), .B(n35462), .Z(n35459) );
  IV U33773 ( .A(n35437), .Z(n35455) );
  XOR U33774 ( .A(n35463), .B(n35464), .Z(n35437) );
  ANDN U33775 ( .B(n35465), .A(n35466), .Z(n35463) );
  XOR U33776 ( .A(n35464), .B(n35467), .Z(n35465) );
  XOR U33777 ( .A(n35446), .B(n35377), .Z(n35447) );
  XOR U33778 ( .A(n35468), .B(n35469), .Z(n35377) );
  AND U33779 ( .A(n1014), .B(n35470), .Z(n35468) );
  XOR U33780 ( .A(n35471), .B(n35469), .Z(n35470) );
  XNOR U33781 ( .A(n35472), .B(n35473), .Z(n35446) );
  NAND U33782 ( .A(n35474), .B(n35475), .Z(n35473) );
  XOR U33783 ( .A(n35476), .B(n35425), .Z(n35475) );
  XOR U33784 ( .A(n35466), .B(n35467), .Z(n35425) );
  XOR U33785 ( .A(n35477), .B(n35454), .Z(n35467) );
  XOR U33786 ( .A(n35478), .B(n35479), .Z(n35454) );
  ANDN U33787 ( .B(n35480), .A(n35481), .Z(n35478) );
  XOR U33788 ( .A(n35479), .B(n35482), .Z(n35480) );
  IV U33789 ( .A(n35452), .Z(n35477) );
  XOR U33790 ( .A(n35450), .B(n35483), .Z(n35452) );
  XOR U33791 ( .A(n35484), .B(n35485), .Z(n35483) );
  ANDN U33792 ( .B(n35486), .A(n35487), .Z(n35484) );
  XOR U33793 ( .A(n35488), .B(n35485), .Z(n35486) );
  IV U33794 ( .A(n35453), .Z(n35450) );
  XOR U33795 ( .A(n35489), .B(n35490), .Z(n35453) );
  ANDN U33796 ( .B(n35491), .A(n35492), .Z(n35489) );
  XOR U33797 ( .A(n35490), .B(n35493), .Z(n35491) );
  XOR U33798 ( .A(n35494), .B(n35495), .Z(n35466) );
  XNOR U33799 ( .A(n35461), .B(n35496), .Z(n35495) );
  IV U33800 ( .A(n35464), .Z(n35496) );
  XOR U33801 ( .A(n35497), .B(n35498), .Z(n35464) );
  ANDN U33802 ( .B(n35499), .A(n35500), .Z(n35497) );
  XOR U33803 ( .A(n35498), .B(n35501), .Z(n35499) );
  XNOR U33804 ( .A(n35502), .B(n35503), .Z(n35461) );
  ANDN U33805 ( .B(n35504), .A(n35505), .Z(n35502) );
  XOR U33806 ( .A(n35503), .B(n35506), .Z(n35504) );
  IV U33807 ( .A(n35460), .Z(n35494) );
  XOR U33808 ( .A(n35458), .B(n35507), .Z(n35460) );
  XOR U33809 ( .A(n35508), .B(n35509), .Z(n35507) );
  ANDN U33810 ( .B(n35510), .A(n35511), .Z(n35508) );
  XOR U33811 ( .A(n35512), .B(n35509), .Z(n35510) );
  IV U33812 ( .A(n35462), .Z(n35458) );
  XOR U33813 ( .A(n35513), .B(n35514), .Z(n35462) );
  ANDN U33814 ( .B(n35515), .A(n35516), .Z(n35513) );
  XOR U33815 ( .A(n35517), .B(n35514), .Z(n35515) );
  IV U33816 ( .A(n35472), .Z(n35476) );
  XOR U33817 ( .A(n35472), .B(n35427), .Z(n35474) );
  XOR U33818 ( .A(n35518), .B(n35519), .Z(n35427) );
  AND U33819 ( .A(n1014), .B(n35520), .Z(n35518) );
  XOR U33820 ( .A(n35521), .B(n35519), .Z(n35520) );
  NANDN U33821 ( .A(n35429), .B(n35431), .Z(n35472) );
  XOR U33822 ( .A(n35522), .B(n35523), .Z(n35431) );
  AND U33823 ( .A(n1014), .B(n35524), .Z(n35522) );
  XOR U33824 ( .A(n35523), .B(n35525), .Z(n35524) );
  XNOR U33825 ( .A(n35526), .B(n35527), .Z(n1014) );
  AND U33826 ( .A(n35528), .B(n35529), .Z(n35526) );
  XOR U33827 ( .A(n35527), .B(n35442), .Z(n35529) );
  XNOR U33828 ( .A(n35530), .B(n35531), .Z(n35442) );
  ANDN U33829 ( .B(n35532), .A(n35533), .Z(n35530) );
  XOR U33830 ( .A(n35531), .B(n35534), .Z(n35532) );
  XNOR U33831 ( .A(n35527), .B(n35444), .Z(n35528) );
  XOR U33832 ( .A(n35535), .B(n35536), .Z(n35444) );
  AND U33833 ( .A(n1018), .B(n35537), .Z(n35535) );
  XOR U33834 ( .A(n35538), .B(n35536), .Z(n35537) );
  XNOR U33835 ( .A(n35539), .B(n35540), .Z(n35527) );
  AND U33836 ( .A(n35541), .B(n35542), .Z(n35539) );
  XNOR U33837 ( .A(n35540), .B(n35469), .Z(n35542) );
  XOR U33838 ( .A(n35533), .B(n35534), .Z(n35469) );
  XNOR U33839 ( .A(n35543), .B(n35544), .Z(n35534) );
  ANDN U33840 ( .B(n35545), .A(n35546), .Z(n35543) );
  XOR U33841 ( .A(n35547), .B(n35548), .Z(n35545) );
  XOR U33842 ( .A(n35549), .B(n35550), .Z(n35533) );
  XNOR U33843 ( .A(n35551), .B(n35552), .Z(n35550) );
  ANDN U33844 ( .B(n35553), .A(n35554), .Z(n35551) );
  XNOR U33845 ( .A(n35555), .B(n35556), .Z(n35553) );
  IV U33846 ( .A(n35531), .Z(n35549) );
  XOR U33847 ( .A(n35557), .B(n35558), .Z(n35531) );
  ANDN U33848 ( .B(n35559), .A(n35560), .Z(n35557) );
  XOR U33849 ( .A(n35558), .B(n35561), .Z(n35559) );
  XOR U33850 ( .A(n35540), .B(n35471), .Z(n35541) );
  XOR U33851 ( .A(n35562), .B(n35563), .Z(n35471) );
  AND U33852 ( .A(n1018), .B(n35564), .Z(n35562) );
  XNOR U33853 ( .A(n35565), .B(n35563), .Z(n35564) );
  XNOR U33854 ( .A(n35566), .B(n35567), .Z(n35540) );
  NAND U33855 ( .A(n35568), .B(n35569), .Z(n35567) );
  XOR U33856 ( .A(n35570), .B(n35519), .Z(n35569) );
  XOR U33857 ( .A(n35560), .B(n35561), .Z(n35519) );
  XOR U33858 ( .A(n35571), .B(n35548), .Z(n35561) );
  XOR U33859 ( .A(n35572), .B(n35573), .Z(n35548) );
  ANDN U33860 ( .B(n35574), .A(n35575), .Z(n35572) );
  XOR U33861 ( .A(n35573), .B(n35576), .Z(n35574) );
  IV U33862 ( .A(n35546), .Z(n35571) );
  XOR U33863 ( .A(n35544), .B(n35577), .Z(n35546) );
  XOR U33864 ( .A(n35578), .B(n35579), .Z(n35577) );
  ANDN U33865 ( .B(n35580), .A(n35581), .Z(n35578) );
  XOR U33866 ( .A(n35582), .B(n35579), .Z(n35580) );
  IV U33867 ( .A(n35547), .Z(n35544) );
  XOR U33868 ( .A(n35583), .B(n35584), .Z(n35547) );
  ANDN U33869 ( .B(n35585), .A(n35586), .Z(n35583) );
  XOR U33870 ( .A(n35584), .B(n35587), .Z(n35585) );
  XOR U33871 ( .A(n35588), .B(n35589), .Z(n35560) );
  XNOR U33872 ( .A(n35555), .B(n35590), .Z(n35589) );
  IV U33873 ( .A(n35558), .Z(n35590) );
  XOR U33874 ( .A(n35591), .B(n35592), .Z(n35558) );
  ANDN U33875 ( .B(n35593), .A(n35594), .Z(n35591) );
  XOR U33876 ( .A(n35592), .B(n35595), .Z(n35593) );
  XNOR U33877 ( .A(n35596), .B(n35597), .Z(n35555) );
  ANDN U33878 ( .B(n35598), .A(n35599), .Z(n35596) );
  XOR U33879 ( .A(n35597), .B(n35600), .Z(n35598) );
  IV U33880 ( .A(n35554), .Z(n35588) );
  XOR U33881 ( .A(n35552), .B(n35601), .Z(n35554) );
  XOR U33882 ( .A(n35602), .B(n35603), .Z(n35601) );
  ANDN U33883 ( .B(n35604), .A(n35605), .Z(n35602) );
  XOR U33884 ( .A(n35606), .B(n35603), .Z(n35604) );
  IV U33885 ( .A(n35556), .Z(n35552) );
  XOR U33886 ( .A(n35607), .B(n35608), .Z(n35556) );
  ANDN U33887 ( .B(n35609), .A(n35610), .Z(n35607) );
  XOR U33888 ( .A(n35611), .B(n35608), .Z(n35609) );
  IV U33889 ( .A(n35566), .Z(n35570) );
  XOR U33890 ( .A(n35566), .B(n35521), .Z(n35568) );
  XOR U33891 ( .A(n35612), .B(n35613), .Z(n35521) );
  AND U33892 ( .A(n1018), .B(n35614), .Z(n35612) );
  XNOR U33893 ( .A(n35615), .B(n35613), .Z(n35614) );
  NANDN U33894 ( .A(n35523), .B(n35525), .Z(n35566) );
  XOR U33895 ( .A(n35616), .B(n35617), .Z(n35525) );
  AND U33896 ( .A(n1018), .B(n35618), .Z(n35616) );
  XOR U33897 ( .A(n35617), .B(n35619), .Z(n35618) );
  XNOR U33898 ( .A(n35620), .B(n35621), .Z(n1018) );
  AND U33899 ( .A(n35622), .B(n35623), .Z(n35620) );
  XOR U33900 ( .A(n35621), .B(n35536), .Z(n35623) );
  XNOR U33901 ( .A(n35624), .B(n35625), .Z(n35536) );
  ANDN U33902 ( .B(n35626), .A(n35627), .Z(n35624) );
  XOR U33903 ( .A(n35625), .B(n35628), .Z(n35626) );
  XNOR U33904 ( .A(n35621), .B(n35538), .Z(n35622) );
  XNOR U33905 ( .A(n35629), .B(n35630), .Z(n35538) );
  ANDN U33906 ( .B(n35631), .A(n35632), .Z(n35629) );
  XOR U33907 ( .A(n35630), .B(n35633), .Z(n35631) );
  XNOR U33908 ( .A(n35634), .B(n35635), .Z(n35621) );
  AND U33909 ( .A(n35636), .B(n35637), .Z(n35634) );
  XNOR U33910 ( .A(n35635), .B(n35563), .Z(n35637) );
  XOR U33911 ( .A(n35627), .B(n35628), .Z(n35563) );
  XNOR U33912 ( .A(n35638), .B(n35639), .Z(n35628) );
  ANDN U33913 ( .B(n35640), .A(n35641), .Z(n35638) );
  XOR U33914 ( .A(n35642), .B(n35643), .Z(n35640) );
  XOR U33915 ( .A(n35644), .B(n35645), .Z(n35627) );
  XNOR U33916 ( .A(n35646), .B(n35647), .Z(n35645) );
  ANDN U33917 ( .B(n35648), .A(n35649), .Z(n35646) );
  XNOR U33918 ( .A(n35650), .B(n35651), .Z(n35648) );
  IV U33919 ( .A(n35625), .Z(n35644) );
  XOR U33920 ( .A(n35652), .B(n35653), .Z(n35625) );
  ANDN U33921 ( .B(n35654), .A(n35655), .Z(n35652) );
  XOR U33922 ( .A(n35653), .B(n35656), .Z(n35654) );
  XNOR U33923 ( .A(n35635), .B(n35565), .Z(n35636) );
  XOR U33924 ( .A(n35657), .B(n35633), .Z(n35565) );
  XNOR U33925 ( .A(n35658), .B(n35659), .Z(n35633) );
  ANDN U33926 ( .B(n35660), .A(n35661), .Z(n35658) );
  XOR U33927 ( .A(n35662), .B(n35663), .Z(n35660) );
  IV U33928 ( .A(n35632), .Z(n35657) );
  XOR U33929 ( .A(n35664), .B(n35665), .Z(n35632) );
  XNOR U33930 ( .A(n35666), .B(n35667), .Z(n35665) );
  ANDN U33931 ( .B(n35668), .A(n35669), .Z(n35666) );
  XNOR U33932 ( .A(n35670), .B(n35671), .Z(n35668) );
  IV U33933 ( .A(n35630), .Z(n35664) );
  XOR U33934 ( .A(n35672), .B(n35673), .Z(n35630) );
  ANDN U33935 ( .B(n35674), .A(n35675), .Z(n35672) );
  XOR U33936 ( .A(n35673), .B(n35676), .Z(n35674) );
  XNOR U33937 ( .A(n35677), .B(n35678), .Z(n35635) );
  NAND U33938 ( .A(n35679), .B(n35680), .Z(n35678) );
  XOR U33939 ( .A(n35681), .B(n35613), .Z(n35680) );
  XOR U33940 ( .A(n35655), .B(n35656), .Z(n35613) );
  XOR U33941 ( .A(n35682), .B(n35643), .Z(n35656) );
  XOR U33942 ( .A(n35683), .B(n35684), .Z(n35643) );
  ANDN U33943 ( .B(n35685), .A(n35686), .Z(n35683) );
  XOR U33944 ( .A(n35684), .B(n35687), .Z(n35685) );
  IV U33945 ( .A(n35641), .Z(n35682) );
  XOR U33946 ( .A(n35639), .B(n35688), .Z(n35641) );
  XOR U33947 ( .A(n35689), .B(n35690), .Z(n35688) );
  ANDN U33948 ( .B(n35691), .A(n35692), .Z(n35689) );
  XOR U33949 ( .A(n35693), .B(n35690), .Z(n35691) );
  IV U33950 ( .A(n35642), .Z(n35639) );
  XOR U33951 ( .A(n35694), .B(n35695), .Z(n35642) );
  ANDN U33952 ( .B(n35696), .A(n35697), .Z(n35694) );
  XOR U33953 ( .A(n35695), .B(n35698), .Z(n35696) );
  XOR U33954 ( .A(n35699), .B(n35700), .Z(n35655) );
  XNOR U33955 ( .A(n35650), .B(n35701), .Z(n35700) );
  IV U33956 ( .A(n35653), .Z(n35701) );
  XOR U33957 ( .A(n35702), .B(n35703), .Z(n35653) );
  ANDN U33958 ( .B(n35704), .A(n35705), .Z(n35702) );
  XOR U33959 ( .A(n35703), .B(n35706), .Z(n35704) );
  XNOR U33960 ( .A(n35707), .B(n35708), .Z(n35650) );
  ANDN U33961 ( .B(n35709), .A(n35710), .Z(n35707) );
  XOR U33962 ( .A(n35708), .B(n35711), .Z(n35709) );
  IV U33963 ( .A(n35649), .Z(n35699) );
  XOR U33964 ( .A(n35647), .B(n35712), .Z(n35649) );
  XOR U33965 ( .A(n35713), .B(n35714), .Z(n35712) );
  ANDN U33966 ( .B(n35715), .A(n35716), .Z(n35713) );
  XOR U33967 ( .A(n35717), .B(n35714), .Z(n35715) );
  IV U33968 ( .A(n35651), .Z(n35647) );
  XOR U33969 ( .A(n35718), .B(n35719), .Z(n35651) );
  ANDN U33970 ( .B(n35720), .A(n35721), .Z(n35718) );
  XOR U33971 ( .A(n35722), .B(n35719), .Z(n35720) );
  IV U33972 ( .A(n35677), .Z(n35681) );
  XNOR U33973 ( .A(n35677), .B(n35615), .Z(n35679) );
  XOR U33974 ( .A(n35723), .B(n35676), .Z(n35615) );
  XOR U33975 ( .A(n35724), .B(n35663), .Z(n35676) );
  XOR U33976 ( .A(n35725), .B(n35726), .Z(n35663) );
  ANDN U33977 ( .B(n35727), .A(n35728), .Z(n35725) );
  XOR U33978 ( .A(n35726), .B(n35729), .Z(n35727) );
  IV U33979 ( .A(n35661), .Z(n35724) );
  XOR U33980 ( .A(n35659), .B(n35730), .Z(n35661) );
  XOR U33981 ( .A(n35731), .B(n35732), .Z(n35730) );
  ANDN U33982 ( .B(n35733), .A(n35734), .Z(n35731) );
  XOR U33983 ( .A(n35735), .B(n35732), .Z(n35733) );
  IV U33984 ( .A(n35662), .Z(n35659) );
  XOR U33985 ( .A(n35736), .B(n35737), .Z(n35662) );
  ANDN U33986 ( .B(n35738), .A(n35739), .Z(n35736) );
  XOR U33987 ( .A(n35737), .B(n35740), .Z(n35738) );
  IV U33988 ( .A(n35675), .Z(n35723) );
  XOR U33989 ( .A(n35741), .B(n35742), .Z(n35675) );
  XNOR U33990 ( .A(n35670), .B(n35743), .Z(n35742) );
  IV U33991 ( .A(n35673), .Z(n35743) );
  XNOR U33992 ( .A(n35744), .B(n35745), .Z(n35673) );
  ANDN U33993 ( .B(n35746), .A(n35747), .Z(n35744) );
  XNOR U33994 ( .A(n35745), .B(n35748), .Z(n35746) );
  XNOR U33995 ( .A(n35749), .B(n35750), .Z(n35670) );
  ANDN U33996 ( .B(n35751), .A(n35752), .Z(n35749) );
  XOR U33997 ( .A(n35750), .B(n35753), .Z(n35751) );
  IV U33998 ( .A(n35669), .Z(n35741) );
  XOR U33999 ( .A(n35667), .B(n35754), .Z(n35669) );
  XOR U34000 ( .A(n35755), .B(n35756), .Z(n35754) );
  ANDN U34001 ( .B(n35757), .A(n35758), .Z(n35755) );
  XOR U34002 ( .A(n35759), .B(n35756), .Z(n35757) );
  IV U34003 ( .A(n35671), .Z(n35667) );
  XOR U34004 ( .A(n35760), .B(n35761), .Z(n35671) );
  ANDN U34005 ( .B(n35762), .A(n35763), .Z(n35760) );
  XOR U34006 ( .A(n35764), .B(n35761), .Z(n35762) );
  NANDN U34007 ( .A(n35617), .B(n35619), .Z(n35677) );
  XOR U34008 ( .A(n35765), .B(n35748), .Z(n35619) );
  XOR U34009 ( .A(n35766), .B(n35740), .Z(n35748) );
  XOR U34010 ( .A(n35767), .B(n35729), .Z(n35740) );
  XNOR U34011 ( .A(q[14]), .B(DB[14]), .Z(n35729) );
  IV U34012 ( .A(n35728), .Z(n35767) );
  XNOR U34013 ( .A(n35726), .B(n35768), .Z(n35728) );
  XNOR U34014 ( .A(q[13]), .B(DB[13]), .Z(n35768) );
  XNOR U34015 ( .A(q[12]), .B(DB[12]), .Z(n35726) );
  IV U34016 ( .A(n35739), .Z(n35766) );
  XOR U34017 ( .A(n35769), .B(n35770), .Z(n35739) );
  XNOR U34018 ( .A(n35735), .B(n35737), .Z(n35770) );
  XNOR U34019 ( .A(q[8]), .B(DB[8]), .Z(n35737) );
  XNOR U34020 ( .A(q[11]), .B(DB[11]), .Z(n35735) );
  IV U34021 ( .A(n35734), .Z(n35769) );
  XNOR U34022 ( .A(n35732), .B(n35771), .Z(n35734) );
  XNOR U34023 ( .A(q[10]), .B(DB[10]), .Z(n35771) );
  XNOR U34024 ( .A(q[9]), .B(DB[9]), .Z(n35732) );
  IV U34025 ( .A(n35747), .Z(n35765) );
  XOR U34026 ( .A(n35772), .B(n35773), .Z(n35747) );
  XOR U34027 ( .A(n35745), .B(n35764), .Z(n35773) );
  XOR U34028 ( .A(n35774), .B(n35753), .Z(n35764) );
  XNOR U34029 ( .A(q[7]), .B(DB[7]), .Z(n35753) );
  IV U34030 ( .A(n35752), .Z(n35774) );
  XNOR U34031 ( .A(n35750), .B(n35775), .Z(n35752) );
  XNOR U34032 ( .A(q[6]), .B(DB[6]), .Z(n35775) );
  XNOR U34033 ( .A(q[5]), .B(DB[5]), .Z(n35750) );
  XOR U34034 ( .A(q[0]), .B(DB[0]), .Z(n35745) );
  IV U34035 ( .A(n35763), .Z(n35772) );
  XOR U34036 ( .A(n35776), .B(n35777), .Z(n35763) );
  XNOR U34037 ( .A(n35759), .B(n35761), .Z(n35777) );
  XNOR U34038 ( .A(q[1]), .B(DB[1]), .Z(n35761) );
  XNOR U34039 ( .A(q[4]), .B(DB[4]), .Z(n35759) );
  IV U34040 ( .A(n35758), .Z(n35776) );
  XNOR U34041 ( .A(n35756), .B(n35778), .Z(n35758) );
  XNOR U34042 ( .A(q[3]), .B(DB[3]), .Z(n35778) );
  XNOR U34043 ( .A(q[2]), .B(DB[2]), .Z(n35756) );
  XOR U34044 ( .A(n35779), .B(n35706), .Z(n35617) );
  XOR U34045 ( .A(n35780), .B(n35698), .Z(n35706) );
  XOR U34046 ( .A(n35781), .B(n35687), .Z(n35698) );
  XNOR U34047 ( .A(q[14]), .B(DB[29]), .Z(n35687) );
  IV U34048 ( .A(n35686), .Z(n35781) );
  XNOR U34049 ( .A(n35684), .B(n35782), .Z(n35686) );
  XNOR U34050 ( .A(q[13]), .B(DB[28]), .Z(n35782) );
  XNOR U34051 ( .A(q[12]), .B(DB[27]), .Z(n35684) );
  IV U34052 ( .A(n35697), .Z(n35780) );
  XOR U34053 ( .A(n35783), .B(n35784), .Z(n35697) );
  XNOR U34054 ( .A(n35693), .B(n35695), .Z(n35784) );
  XNOR U34055 ( .A(q[8]), .B(DB[23]), .Z(n35695) );
  XNOR U34056 ( .A(q[11]), .B(DB[26]), .Z(n35693) );
  IV U34057 ( .A(n35692), .Z(n35783) );
  XNOR U34058 ( .A(n35690), .B(n35785), .Z(n35692) );
  XNOR U34059 ( .A(q[10]), .B(DB[25]), .Z(n35785) );
  XNOR U34060 ( .A(q[9]), .B(DB[24]), .Z(n35690) );
  IV U34061 ( .A(n35705), .Z(n35779) );
  XOR U34062 ( .A(n35786), .B(n35787), .Z(n35705) );
  XNOR U34063 ( .A(n35722), .B(n35703), .Z(n35787) );
  XNOR U34064 ( .A(q[0]), .B(DB[15]), .Z(n35703) );
  XOR U34065 ( .A(n35788), .B(n35711), .Z(n35722) );
  XNOR U34066 ( .A(q[7]), .B(DB[22]), .Z(n35711) );
  IV U34067 ( .A(n35710), .Z(n35788) );
  XNOR U34068 ( .A(n35708), .B(n35789), .Z(n35710) );
  XNOR U34069 ( .A(q[6]), .B(DB[21]), .Z(n35789) );
  XNOR U34070 ( .A(q[5]), .B(DB[20]), .Z(n35708) );
  IV U34071 ( .A(n35721), .Z(n35786) );
  XOR U34072 ( .A(n35790), .B(n35791), .Z(n35721) );
  XNOR U34073 ( .A(n35717), .B(n35719), .Z(n35791) );
  XNOR U34074 ( .A(q[1]), .B(DB[16]), .Z(n35719) );
  XNOR U34075 ( .A(q[4]), .B(DB[19]), .Z(n35717) );
  IV U34076 ( .A(n35716), .Z(n35790) );
  XNOR U34077 ( .A(n35714), .B(n35792), .Z(n35716) );
  XNOR U34078 ( .A(q[3]), .B(DB[18]), .Z(n35792) );
  XNOR U34079 ( .A(q[2]), .B(DB[17]), .Z(n35714) );
  XOR U34080 ( .A(n35793), .B(n35595), .Z(n35523) );
  XOR U34081 ( .A(n35794), .B(n35587), .Z(n35595) );
  XOR U34082 ( .A(n35795), .B(n35576), .Z(n35587) );
  XNOR U34083 ( .A(q[14]), .B(DB[44]), .Z(n35576) );
  IV U34084 ( .A(n35575), .Z(n35795) );
  XNOR U34085 ( .A(n35573), .B(n35796), .Z(n35575) );
  XNOR U34086 ( .A(q[13]), .B(DB[43]), .Z(n35796) );
  XNOR U34087 ( .A(q[12]), .B(DB[42]), .Z(n35573) );
  IV U34088 ( .A(n35586), .Z(n35794) );
  XOR U34089 ( .A(n35797), .B(n35798), .Z(n35586) );
  XNOR U34090 ( .A(n35582), .B(n35584), .Z(n35798) );
  XNOR U34091 ( .A(q[8]), .B(DB[38]), .Z(n35584) );
  XNOR U34092 ( .A(q[11]), .B(DB[41]), .Z(n35582) );
  IV U34093 ( .A(n35581), .Z(n35797) );
  XNOR U34094 ( .A(n35579), .B(n35799), .Z(n35581) );
  XNOR U34095 ( .A(q[10]), .B(DB[40]), .Z(n35799) );
  XNOR U34096 ( .A(q[9]), .B(DB[39]), .Z(n35579) );
  IV U34097 ( .A(n35594), .Z(n35793) );
  XOR U34098 ( .A(n35800), .B(n35801), .Z(n35594) );
  XNOR U34099 ( .A(n35611), .B(n35592), .Z(n35801) );
  XNOR U34100 ( .A(q[0]), .B(DB[30]), .Z(n35592) );
  XOR U34101 ( .A(n35802), .B(n35600), .Z(n35611) );
  XNOR U34102 ( .A(q[7]), .B(DB[37]), .Z(n35600) );
  IV U34103 ( .A(n35599), .Z(n35802) );
  XNOR U34104 ( .A(n35597), .B(n35803), .Z(n35599) );
  XNOR U34105 ( .A(q[6]), .B(DB[36]), .Z(n35803) );
  XNOR U34106 ( .A(q[5]), .B(DB[35]), .Z(n35597) );
  IV U34107 ( .A(n35610), .Z(n35800) );
  XOR U34108 ( .A(n35804), .B(n35805), .Z(n35610) );
  XNOR U34109 ( .A(n35606), .B(n35608), .Z(n35805) );
  XNOR U34110 ( .A(q[1]), .B(DB[31]), .Z(n35608) );
  XNOR U34111 ( .A(q[4]), .B(DB[34]), .Z(n35606) );
  IV U34112 ( .A(n35605), .Z(n35804) );
  XNOR U34113 ( .A(n35603), .B(n35806), .Z(n35605) );
  XNOR U34114 ( .A(q[3]), .B(DB[33]), .Z(n35806) );
  XNOR U34115 ( .A(q[2]), .B(DB[32]), .Z(n35603) );
  XOR U34116 ( .A(n35807), .B(n35501), .Z(n35429) );
  XOR U34117 ( .A(n35808), .B(n35493), .Z(n35501) );
  XOR U34118 ( .A(n35809), .B(n35482), .Z(n35493) );
  XNOR U34119 ( .A(q[14]), .B(DB[59]), .Z(n35482) );
  IV U34120 ( .A(n35481), .Z(n35809) );
  XNOR U34121 ( .A(n35479), .B(n35810), .Z(n35481) );
  XNOR U34122 ( .A(q[13]), .B(DB[58]), .Z(n35810) );
  XNOR U34123 ( .A(q[12]), .B(DB[57]), .Z(n35479) );
  IV U34124 ( .A(n35492), .Z(n35808) );
  XOR U34125 ( .A(n35811), .B(n35812), .Z(n35492) );
  XNOR U34126 ( .A(n35488), .B(n35490), .Z(n35812) );
  XNOR U34127 ( .A(q[8]), .B(DB[53]), .Z(n35490) );
  XNOR U34128 ( .A(q[11]), .B(DB[56]), .Z(n35488) );
  IV U34129 ( .A(n35487), .Z(n35811) );
  XNOR U34130 ( .A(n35485), .B(n35813), .Z(n35487) );
  XNOR U34131 ( .A(q[10]), .B(DB[55]), .Z(n35813) );
  XNOR U34132 ( .A(q[9]), .B(DB[54]), .Z(n35485) );
  IV U34133 ( .A(n35500), .Z(n35807) );
  XOR U34134 ( .A(n35814), .B(n35815), .Z(n35500) );
  XNOR U34135 ( .A(n35517), .B(n35498), .Z(n35815) );
  XNOR U34136 ( .A(q[0]), .B(DB[45]), .Z(n35498) );
  XOR U34137 ( .A(n35816), .B(n35506), .Z(n35517) );
  XNOR U34138 ( .A(q[7]), .B(DB[52]), .Z(n35506) );
  IV U34139 ( .A(n35505), .Z(n35816) );
  XNOR U34140 ( .A(n35503), .B(n35817), .Z(n35505) );
  XNOR U34141 ( .A(q[6]), .B(DB[51]), .Z(n35817) );
  XNOR U34142 ( .A(q[5]), .B(DB[50]), .Z(n35503) );
  IV U34143 ( .A(n35516), .Z(n35814) );
  XOR U34144 ( .A(n35818), .B(n35819), .Z(n35516) );
  XNOR U34145 ( .A(n35512), .B(n35514), .Z(n35819) );
  XNOR U34146 ( .A(q[1]), .B(DB[46]), .Z(n35514) );
  XNOR U34147 ( .A(q[4]), .B(DB[49]), .Z(n35512) );
  IV U34148 ( .A(n35511), .Z(n35818) );
  XNOR U34149 ( .A(n35509), .B(n35820), .Z(n35511) );
  XNOR U34150 ( .A(q[3]), .B(DB[48]), .Z(n35820) );
  XNOR U34151 ( .A(q[2]), .B(DB[47]), .Z(n35509) );
  XOR U34152 ( .A(n35821), .B(n35407), .Z(n35335) );
  XOR U34153 ( .A(n35822), .B(n35399), .Z(n35407) );
  XOR U34154 ( .A(n35823), .B(n35388), .Z(n35399) );
  XNOR U34155 ( .A(q[14]), .B(DB[74]), .Z(n35388) );
  IV U34156 ( .A(n35387), .Z(n35823) );
  XNOR U34157 ( .A(n35385), .B(n35824), .Z(n35387) );
  XNOR U34158 ( .A(q[13]), .B(DB[73]), .Z(n35824) );
  XNOR U34159 ( .A(q[12]), .B(DB[72]), .Z(n35385) );
  IV U34160 ( .A(n35398), .Z(n35822) );
  XOR U34161 ( .A(n35825), .B(n35826), .Z(n35398) );
  XNOR U34162 ( .A(n35394), .B(n35396), .Z(n35826) );
  XNOR U34163 ( .A(q[8]), .B(DB[68]), .Z(n35396) );
  XNOR U34164 ( .A(q[11]), .B(DB[71]), .Z(n35394) );
  IV U34165 ( .A(n35393), .Z(n35825) );
  XNOR U34166 ( .A(n35391), .B(n35827), .Z(n35393) );
  XNOR U34167 ( .A(q[10]), .B(DB[70]), .Z(n35827) );
  XNOR U34168 ( .A(q[9]), .B(DB[69]), .Z(n35391) );
  IV U34169 ( .A(n35406), .Z(n35821) );
  XOR U34170 ( .A(n35828), .B(n35829), .Z(n35406) );
  XNOR U34171 ( .A(n35423), .B(n35404), .Z(n35829) );
  XNOR U34172 ( .A(q[0]), .B(DB[60]), .Z(n35404) );
  XOR U34173 ( .A(n35830), .B(n35412), .Z(n35423) );
  XNOR U34174 ( .A(q[7]), .B(DB[67]), .Z(n35412) );
  IV U34175 ( .A(n35411), .Z(n35830) );
  XNOR U34176 ( .A(n35409), .B(n35831), .Z(n35411) );
  XNOR U34177 ( .A(q[6]), .B(DB[66]), .Z(n35831) );
  XNOR U34178 ( .A(q[5]), .B(DB[65]), .Z(n35409) );
  IV U34179 ( .A(n35422), .Z(n35828) );
  XOR U34180 ( .A(n35832), .B(n35833), .Z(n35422) );
  XNOR U34181 ( .A(n35418), .B(n35420), .Z(n35833) );
  XNOR U34182 ( .A(q[1]), .B(DB[61]), .Z(n35420) );
  XNOR U34183 ( .A(q[4]), .B(DB[64]), .Z(n35418) );
  IV U34184 ( .A(n35417), .Z(n35832) );
  XNOR U34185 ( .A(n35415), .B(n35834), .Z(n35417) );
  XNOR U34186 ( .A(q[3]), .B(DB[63]), .Z(n35834) );
  XNOR U34187 ( .A(q[2]), .B(DB[62]), .Z(n35415) );
  XOR U34188 ( .A(n35835), .B(n35313), .Z(n35241) );
  XOR U34189 ( .A(n35836), .B(n35305), .Z(n35313) );
  XOR U34190 ( .A(n35837), .B(n35294), .Z(n35305) );
  XNOR U34191 ( .A(q[14]), .B(DB[89]), .Z(n35294) );
  IV U34192 ( .A(n35293), .Z(n35837) );
  XNOR U34193 ( .A(n35291), .B(n35838), .Z(n35293) );
  XNOR U34194 ( .A(q[13]), .B(DB[88]), .Z(n35838) );
  XNOR U34195 ( .A(q[12]), .B(DB[87]), .Z(n35291) );
  IV U34196 ( .A(n35304), .Z(n35836) );
  XOR U34197 ( .A(n35839), .B(n35840), .Z(n35304) );
  XNOR U34198 ( .A(n35300), .B(n35302), .Z(n35840) );
  XNOR U34199 ( .A(q[8]), .B(DB[83]), .Z(n35302) );
  XNOR U34200 ( .A(q[11]), .B(DB[86]), .Z(n35300) );
  IV U34201 ( .A(n35299), .Z(n35839) );
  XNOR U34202 ( .A(n35297), .B(n35841), .Z(n35299) );
  XNOR U34203 ( .A(q[10]), .B(DB[85]), .Z(n35841) );
  XNOR U34204 ( .A(q[9]), .B(DB[84]), .Z(n35297) );
  IV U34205 ( .A(n35312), .Z(n35835) );
  XOR U34206 ( .A(n35842), .B(n35843), .Z(n35312) );
  XNOR U34207 ( .A(n35329), .B(n35310), .Z(n35843) );
  XNOR U34208 ( .A(q[0]), .B(DB[75]), .Z(n35310) );
  XOR U34209 ( .A(n35844), .B(n35318), .Z(n35329) );
  XNOR U34210 ( .A(q[7]), .B(DB[82]), .Z(n35318) );
  IV U34211 ( .A(n35317), .Z(n35844) );
  XNOR U34212 ( .A(n35315), .B(n35845), .Z(n35317) );
  XNOR U34213 ( .A(q[6]), .B(DB[81]), .Z(n35845) );
  XNOR U34214 ( .A(q[5]), .B(DB[80]), .Z(n35315) );
  IV U34215 ( .A(n35328), .Z(n35842) );
  XOR U34216 ( .A(n35846), .B(n35847), .Z(n35328) );
  XNOR U34217 ( .A(n35324), .B(n35326), .Z(n35847) );
  XNOR U34218 ( .A(q[1]), .B(DB[76]), .Z(n35326) );
  XNOR U34219 ( .A(q[4]), .B(DB[79]), .Z(n35324) );
  IV U34220 ( .A(n35323), .Z(n35846) );
  XNOR U34221 ( .A(n35321), .B(n35848), .Z(n35323) );
  XNOR U34222 ( .A(q[3]), .B(DB[78]), .Z(n35848) );
  XNOR U34223 ( .A(q[2]), .B(DB[77]), .Z(n35321) );
  XOR U34224 ( .A(n35849), .B(n35219), .Z(n35147) );
  XOR U34225 ( .A(n35850), .B(n35211), .Z(n35219) );
  XOR U34226 ( .A(n35851), .B(n35200), .Z(n35211) );
  XNOR U34227 ( .A(q[14]), .B(DB[104]), .Z(n35200) );
  IV U34228 ( .A(n35199), .Z(n35851) );
  XNOR U34229 ( .A(n35197), .B(n35852), .Z(n35199) );
  XNOR U34230 ( .A(q[13]), .B(DB[103]), .Z(n35852) );
  XNOR U34231 ( .A(q[12]), .B(DB[102]), .Z(n35197) );
  IV U34232 ( .A(n35210), .Z(n35850) );
  XOR U34233 ( .A(n35853), .B(n35854), .Z(n35210) );
  XNOR U34234 ( .A(n35206), .B(n35208), .Z(n35854) );
  XNOR U34235 ( .A(q[8]), .B(DB[98]), .Z(n35208) );
  XNOR U34236 ( .A(q[11]), .B(DB[101]), .Z(n35206) );
  IV U34237 ( .A(n35205), .Z(n35853) );
  XNOR U34238 ( .A(n35203), .B(n35855), .Z(n35205) );
  XNOR U34239 ( .A(q[10]), .B(DB[100]), .Z(n35855) );
  XNOR U34240 ( .A(q[9]), .B(DB[99]), .Z(n35203) );
  IV U34241 ( .A(n35218), .Z(n35849) );
  XOR U34242 ( .A(n35856), .B(n35857), .Z(n35218) );
  XNOR U34243 ( .A(n35235), .B(n35216), .Z(n35857) );
  XNOR U34244 ( .A(q[0]), .B(DB[90]), .Z(n35216) );
  XOR U34245 ( .A(n35858), .B(n35224), .Z(n35235) );
  XNOR U34246 ( .A(q[7]), .B(DB[97]), .Z(n35224) );
  IV U34247 ( .A(n35223), .Z(n35858) );
  XNOR U34248 ( .A(n35221), .B(n35859), .Z(n35223) );
  XNOR U34249 ( .A(q[6]), .B(DB[96]), .Z(n35859) );
  XNOR U34250 ( .A(q[5]), .B(DB[95]), .Z(n35221) );
  IV U34251 ( .A(n35234), .Z(n35856) );
  XOR U34252 ( .A(n35860), .B(n35861), .Z(n35234) );
  XNOR U34253 ( .A(n35230), .B(n35232), .Z(n35861) );
  XNOR U34254 ( .A(q[1]), .B(DB[91]), .Z(n35232) );
  XNOR U34255 ( .A(q[4]), .B(DB[94]), .Z(n35230) );
  IV U34256 ( .A(n35229), .Z(n35860) );
  XNOR U34257 ( .A(n35227), .B(n35862), .Z(n35229) );
  XNOR U34258 ( .A(q[3]), .B(DB[93]), .Z(n35862) );
  XNOR U34259 ( .A(q[2]), .B(DB[92]), .Z(n35227) );
  XOR U34260 ( .A(n35863), .B(n35125), .Z(n35053) );
  XOR U34261 ( .A(n35864), .B(n35117), .Z(n35125) );
  XOR U34262 ( .A(n35865), .B(n35106), .Z(n35117) );
  XNOR U34263 ( .A(q[14]), .B(DB[119]), .Z(n35106) );
  IV U34264 ( .A(n35105), .Z(n35865) );
  XNOR U34265 ( .A(n35103), .B(n35866), .Z(n35105) );
  XNOR U34266 ( .A(q[13]), .B(DB[118]), .Z(n35866) );
  XNOR U34267 ( .A(q[12]), .B(DB[117]), .Z(n35103) );
  IV U34268 ( .A(n35116), .Z(n35864) );
  XOR U34269 ( .A(n35867), .B(n35868), .Z(n35116) );
  XNOR U34270 ( .A(n35112), .B(n35114), .Z(n35868) );
  XNOR U34271 ( .A(q[8]), .B(DB[113]), .Z(n35114) );
  XNOR U34272 ( .A(q[11]), .B(DB[116]), .Z(n35112) );
  IV U34273 ( .A(n35111), .Z(n35867) );
  XNOR U34274 ( .A(n35109), .B(n35869), .Z(n35111) );
  XNOR U34275 ( .A(q[10]), .B(DB[115]), .Z(n35869) );
  XNOR U34276 ( .A(q[9]), .B(DB[114]), .Z(n35109) );
  IV U34277 ( .A(n35124), .Z(n35863) );
  XOR U34278 ( .A(n35870), .B(n35871), .Z(n35124) );
  XNOR U34279 ( .A(n35141), .B(n35122), .Z(n35871) );
  XNOR U34280 ( .A(q[0]), .B(DB[105]), .Z(n35122) );
  XOR U34281 ( .A(n35872), .B(n35130), .Z(n35141) );
  XNOR U34282 ( .A(q[7]), .B(DB[112]), .Z(n35130) );
  IV U34283 ( .A(n35129), .Z(n35872) );
  XNOR U34284 ( .A(n35127), .B(n35873), .Z(n35129) );
  XNOR U34285 ( .A(q[6]), .B(DB[111]), .Z(n35873) );
  XNOR U34286 ( .A(q[5]), .B(DB[110]), .Z(n35127) );
  IV U34287 ( .A(n35140), .Z(n35870) );
  XOR U34288 ( .A(n35874), .B(n35875), .Z(n35140) );
  XNOR U34289 ( .A(n35136), .B(n35138), .Z(n35875) );
  XNOR U34290 ( .A(q[1]), .B(DB[106]), .Z(n35138) );
  XNOR U34291 ( .A(q[4]), .B(DB[109]), .Z(n35136) );
  IV U34292 ( .A(n35135), .Z(n35874) );
  XNOR U34293 ( .A(n35133), .B(n35876), .Z(n35135) );
  XNOR U34294 ( .A(q[3]), .B(DB[108]), .Z(n35876) );
  XNOR U34295 ( .A(q[2]), .B(DB[107]), .Z(n35133) );
  XOR U34296 ( .A(n35877), .B(n35031), .Z(n34959) );
  XOR U34297 ( .A(n35878), .B(n35023), .Z(n35031) );
  XOR U34298 ( .A(n35879), .B(n35012), .Z(n35023) );
  XNOR U34299 ( .A(q[14]), .B(DB[134]), .Z(n35012) );
  IV U34300 ( .A(n35011), .Z(n35879) );
  XNOR U34301 ( .A(n35009), .B(n35880), .Z(n35011) );
  XNOR U34302 ( .A(q[13]), .B(DB[133]), .Z(n35880) );
  XNOR U34303 ( .A(q[12]), .B(DB[132]), .Z(n35009) );
  IV U34304 ( .A(n35022), .Z(n35878) );
  XOR U34305 ( .A(n35881), .B(n35882), .Z(n35022) );
  XNOR U34306 ( .A(n35018), .B(n35020), .Z(n35882) );
  XNOR U34307 ( .A(q[8]), .B(DB[128]), .Z(n35020) );
  XNOR U34308 ( .A(q[11]), .B(DB[131]), .Z(n35018) );
  IV U34309 ( .A(n35017), .Z(n35881) );
  XNOR U34310 ( .A(n35015), .B(n35883), .Z(n35017) );
  XNOR U34311 ( .A(q[10]), .B(DB[130]), .Z(n35883) );
  XNOR U34312 ( .A(q[9]), .B(DB[129]), .Z(n35015) );
  IV U34313 ( .A(n35030), .Z(n35877) );
  XOR U34314 ( .A(n35884), .B(n35885), .Z(n35030) );
  XNOR U34315 ( .A(n35047), .B(n35028), .Z(n35885) );
  XNOR U34316 ( .A(q[0]), .B(DB[120]), .Z(n35028) );
  XOR U34317 ( .A(n35886), .B(n35036), .Z(n35047) );
  XNOR U34318 ( .A(q[7]), .B(DB[127]), .Z(n35036) );
  IV U34319 ( .A(n35035), .Z(n35886) );
  XNOR U34320 ( .A(n35033), .B(n35887), .Z(n35035) );
  XNOR U34321 ( .A(q[6]), .B(DB[126]), .Z(n35887) );
  XNOR U34322 ( .A(q[5]), .B(DB[125]), .Z(n35033) );
  IV U34323 ( .A(n35046), .Z(n35884) );
  XOR U34324 ( .A(n35888), .B(n35889), .Z(n35046) );
  XNOR U34325 ( .A(n35042), .B(n35044), .Z(n35889) );
  XNOR U34326 ( .A(q[1]), .B(DB[121]), .Z(n35044) );
  XNOR U34327 ( .A(q[4]), .B(DB[124]), .Z(n35042) );
  IV U34328 ( .A(n35041), .Z(n35888) );
  XNOR U34329 ( .A(n35039), .B(n35890), .Z(n35041) );
  XNOR U34330 ( .A(q[3]), .B(DB[123]), .Z(n35890) );
  XNOR U34331 ( .A(q[2]), .B(DB[122]), .Z(n35039) );
  XOR U34332 ( .A(n35891), .B(n34937), .Z(n34865) );
  XOR U34333 ( .A(n35892), .B(n34929), .Z(n34937) );
  XOR U34334 ( .A(n35893), .B(n34918), .Z(n34929) );
  XNOR U34335 ( .A(q[14]), .B(DB[149]), .Z(n34918) );
  IV U34336 ( .A(n34917), .Z(n35893) );
  XNOR U34337 ( .A(n34915), .B(n35894), .Z(n34917) );
  XNOR U34338 ( .A(q[13]), .B(DB[148]), .Z(n35894) );
  XNOR U34339 ( .A(q[12]), .B(DB[147]), .Z(n34915) );
  IV U34340 ( .A(n34928), .Z(n35892) );
  XOR U34341 ( .A(n35895), .B(n35896), .Z(n34928) );
  XNOR U34342 ( .A(n34924), .B(n34926), .Z(n35896) );
  XNOR U34343 ( .A(q[8]), .B(DB[143]), .Z(n34926) );
  XNOR U34344 ( .A(q[11]), .B(DB[146]), .Z(n34924) );
  IV U34345 ( .A(n34923), .Z(n35895) );
  XNOR U34346 ( .A(n34921), .B(n35897), .Z(n34923) );
  XNOR U34347 ( .A(q[10]), .B(DB[145]), .Z(n35897) );
  XNOR U34348 ( .A(q[9]), .B(DB[144]), .Z(n34921) );
  IV U34349 ( .A(n34936), .Z(n35891) );
  XOR U34350 ( .A(n35898), .B(n35899), .Z(n34936) );
  XNOR U34351 ( .A(n34953), .B(n34934), .Z(n35899) );
  XNOR U34352 ( .A(q[0]), .B(DB[135]), .Z(n34934) );
  XOR U34353 ( .A(n35900), .B(n34942), .Z(n34953) );
  XNOR U34354 ( .A(q[7]), .B(DB[142]), .Z(n34942) );
  IV U34355 ( .A(n34941), .Z(n35900) );
  XNOR U34356 ( .A(n34939), .B(n35901), .Z(n34941) );
  XNOR U34357 ( .A(q[6]), .B(DB[141]), .Z(n35901) );
  XNOR U34358 ( .A(q[5]), .B(DB[140]), .Z(n34939) );
  IV U34359 ( .A(n34952), .Z(n35898) );
  XOR U34360 ( .A(n35902), .B(n35903), .Z(n34952) );
  XNOR U34361 ( .A(n34948), .B(n34950), .Z(n35903) );
  XNOR U34362 ( .A(q[1]), .B(DB[136]), .Z(n34950) );
  XNOR U34363 ( .A(q[4]), .B(DB[139]), .Z(n34948) );
  IV U34364 ( .A(n34947), .Z(n35902) );
  XNOR U34365 ( .A(n34945), .B(n35904), .Z(n34947) );
  XNOR U34366 ( .A(q[3]), .B(DB[138]), .Z(n35904) );
  XNOR U34367 ( .A(q[2]), .B(DB[137]), .Z(n34945) );
  XOR U34368 ( .A(n35905), .B(n34843), .Z(n34771) );
  XOR U34369 ( .A(n35906), .B(n34835), .Z(n34843) );
  XOR U34370 ( .A(n35907), .B(n34824), .Z(n34835) );
  XNOR U34371 ( .A(q[14]), .B(DB[164]), .Z(n34824) );
  IV U34372 ( .A(n34823), .Z(n35907) );
  XNOR U34373 ( .A(n34821), .B(n35908), .Z(n34823) );
  XNOR U34374 ( .A(q[13]), .B(DB[163]), .Z(n35908) );
  XNOR U34375 ( .A(q[12]), .B(DB[162]), .Z(n34821) );
  IV U34376 ( .A(n34834), .Z(n35906) );
  XOR U34377 ( .A(n35909), .B(n35910), .Z(n34834) );
  XNOR U34378 ( .A(n34830), .B(n34832), .Z(n35910) );
  XNOR U34379 ( .A(q[8]), .B(DB[158]), .Z(n34832) );
  XNOR U34380 ( .A(q[11]), .B(DB[161]), .Z(n34830) );
  IV U34381 ( .A(n34829), .Z(n35909) );
  XNOR U34382 ( .A(n34827), .B(n35911), .Z(n34829) );
  XNOR U34383 ( .A(q[10]), .B(DB[160]), .Z(n35911) );
  XNOR U34384 ( .A(q[9]), .B(DB[159]), .Z(n34827) );
  IV U34385 ( .A(n34842), .Z(n35905) );
  XOR U34386 ( .A(n35912), .B(n35913), .Z(n34842) );
  XNOR U34387 ( .A(n34859), .B(n34840), .Z(n35913) );
  XNOR U34388 ( .A(q[0]), .B(DB[150]), .Z(n34840) );
  XOR U34389 ( .A(n35914), .B(n34848), .Z(n34859) );
  XNOR U34390 ( .A(q[7]), .B(DB[157]), .Z(n34848) );
  IV U34391 ( .A(n34847), .Z(n35914) );
  XNOR U34392 ( .A(n34845), .B(n35915), .Z(n34847) );
  XNOR U34393 ( .A(q[6]), .B(DB[156]), .Z(n35915) );
  XNOR U34394 ( .A(q[5]), .B(DB[155]), .Z(n34845) );
  IV U34395 ( .A(n34858), .Z(n35912) );
  XOR U34396 ( .A(n35916), .B(n35917), .Z(n34858) );
  XNOR U34397 ( .A(n34854), .B(n34856), .Z(n35917) );
  XNOR U34398 ( .A(q[1]), .B(DB[151]), .Z(n34856) );
  XNOR U34399 ( .A(q[4]), .B(DB[154]), .Z(n34854) );
  IV U34400 ( .A(n34853), .Z(n35916) );
  XNOR U34401 ( .A(n34851), .B(n35918), .Z(n34853) );
  XNOR U34402 ( .A(q[3]), .B(DB[153]), .Z(n35918) );
  XNOR U34403 ( .A(q[2]), .B(DB[152]), .Z(n34851) );
  XOR U34404 ( .A(n35919), .B(n34749), .Z(n34677) );
  XOR U34405 ( .A(n35920), .B(n34741), .Z(n34749) );
  XOR U34406 ( .A(n35921), .B(n34730), .Z(n34741) );
  XNOR U34407 ( .A(q[14]), .B(DB[179]), .Z(n34730) );
  IV U34408 ( .A(n34729), .Z(n35921) );
  XNOR U34409 ( .A(n34727), .B(n35922), .Z(n34729) );
  XNOR U34410 ( .A(q[13]), .B(DB[178]), .Z(n35922) );
  XNOR U34411 ( .A(q[12]), .B(DB[177]), .Z(n34727) );
  IV U34412 ( .A(n34740), .Z(n35920) );
  XOR U34413 ( .A(n35923), .B(n35924), .Z(n34740) );
  XNOR U34414 ( .A(n34736), .B(n34738), .Z(n35924) );
  XNOR U34415 ( .A(q[8]), .B(DB[173]), .Z(n34738) );
  XNOR U34416 ( .A(q[11]), .B(DB[176]), .Z(n34736) );
  IV U34417 ( .A(n34735), .Z(n35923) );
  XNOR U34418 ( .A(n34733), .B(n35925), .Z(n34735) );
  XNOR U34419 ( .A(q[10]), .B(DB[175]), .Z(n35925) );
  XNOR U34420 ( .A(q[9]), .B(DB[174]), .Z(n34733) );
  IV U34421 ( .A(n34748), .Z(n35919) );
  XOR U34422 ( .A(n35926), .B(n35927), .Z(n34748) );
  XNOR U34423 ( .A(n34765), .B(n34746), .Z(n35927) );
  XNOR U34424 ( .A(q[0]), .B(DB[165]), .Z(n34746) );
  XOR U34425 ( .A(n35928), .B(n34754), .Z(n34765) );
  XNOR U34426 ( .A(q[7]), .B(DB[172]), .Z(n34754) );
  IV U34427 ( .A(n34753), .Z(n35928) );
  XNOR U34428 ( .A(n34751), .B(n35929), .Z(n34753) );
  XNOR U34429 ( .A(q[6]), .B(DB[171]), .Z(n35929) );
  XNOR U34430 ( .A(q[5]), .B(DB[170]), .Z(n34751) );
  IV U34431 ( .A(n34764), .Z(n35926) );
  XOR U34432 ( .A(n35930), .B(n35931), .Z(n34764) );
  XNOR U34433 ( .A(n34760), .B(n34762), .Z(n35931) );
  XNOR U34434 ( .A(q[1]), .B(DB[166]), .Z(n34762) );
  XNOR U34435 ( .A(q[4]), .B(DB[169]), .Z(n34760) );
  IV U34436 ( .A(n34759), .Z(n35930) );
  XNOR U34437 ( .A(n34757), .B(n35932), .Z(n34759) );
  XNOR U34438 ( .A(q[3]), .B(DB[168]), .Z(n35932) );
  XNOR U34439 ( .A(q[2]), .B(DB[167]), .Z(n34757) );
  XOR U34440 ( .A(n35933), .B(n34655), .Z(n34583) );
  XOR U34441 ( .A(n35934), .B(n34647), .Z(n34655) );
  XOR U34442 ( .A(n35935), .B(n34636), .Z(n34647) );
  XNOR U34443 ( .A(q[14]), .B(DB[194]), .Z(n34636) );
  IV U34444 ( .A(n34635), .Z(n35935) );
  XNOR U34445 ( .A(n34633), .B(n35936), .Z(n34635) );
  XNOR U34446 ( .A(q[13]), .B(DB[193]), .Z(n35936) );
  XNOR U34447 ( .A(q[12]), .B(DB[192]), .Z(n34633) );
  IV U34448 ( .A(n34646), .Z(n35934) );
  XOR U34449 ( .A(n35937), .B(n35938), .Z(n34646) );
  XNOR U34450 ( .A(n34642), .B(n34644), .Z(n35938) );
  XNOR U34451 ( .A(q[8]), .B(DB[188]), .Z(n34644) );
  XNOR U34452 ( .A(q[11]), .B(DB[191]), .Z(n34642) );
  IV U34453 ( .A(n34641), .Z(n35937) );
  XNOR U34454 ( .A(n34639), .B(n35939), .Z(n34641) );
  XNOR U34455 ( .A(q[10]), .B(DB[190]), .Z(n35939) );
  XNOR U34456 ( .A(q[9]), .B(DB[189]), .Z(n34639) );
  IV U34457 ( .A(n34654), .Z(n35933) );
  XOR U34458 ( .A(n35940), .B(n35941), .Z(n34654) );
  XNOR U34459 ( .A(n34671), .B(n34652), .Z(n35941) );
  XNOR U34460 ( .A(q[0]), .B(DB[180]), .Z(n34652) );
  XOR U34461 ( .A(n35942), .B(n34660), .Z(n34671) );
  XNOR U34462 ( .A(q[7]), .B(DB[187]), .Z(n34660) );
  IV U34463 ( .A(n34659), .Z(n35942) );
  XNOR U34464 ( .A(n34657), .B(n35943), .Z(n34659) );
  XNOR U34465 ( .A(q[6]), .B(DB[186]), .Z(n35943) );
  XNOR U34466 ( .A(q[5]), .B(DB[185]), .Z(n34657) );
  IV U34467 ( .A(n34670), .Z(n35940) );
  XOR U34468 ( .A(n35944), .B(n35945), .Z(n34670) );
  XNOR U34469 ( .A(n34666), .B(n34668), .Z(n35945) );
  XNOR U34470 ( .A(q[1]), .B(DB[181]), .Z(n34668) );
  XNOR U34471 ( .A(q[4]), .B(DB[184]), .Z(n34666) );
  IV U34472 ( .A(n34665), .Z(n35944) );
  XNOR U34473 ( .A(n34663), .B(n35946), .Z(n34665) );
  XNOR U34474 ( .A(q[3]), .B(DB[183]), .Z(n35946) );
  XNOR U34475 ( .A(q[2]), .B(DB[182]), .Z(n34663) );
  XOR U34476 ( .A(n35947), .B(n34561), .Z(n34489) );
  XOR U34477 ( .A(n35948), .B(n34553), .Z(n34561) );
  XOR U34478 ( .A(n35949), .B(n34542), .Z(n34553) );
  XNOR U34479 ( .A(q[14]), .B(DB[209]), .Z(n34542) );
  IV U34480 ( .A(n34541), .Z(n35949) );
  XNOR U34481 ( .A(n34539), .B(n35950), .Z(n34541) );
  XNOR U34482 ( .A(q[13]), .B(DB[208]), .Z(n35950) );
  XNOR U34483 ( .A(q[12]), .B(DB[207]), .Z(n34539) );
  IV U34484 ( .A(n34552), .Z(n35948) );
  XOR U34485 ( .A(n35951), .B(n35952), .Z(n34552) );
  XNOR U34486 ( .A(n34548), .B(n34550), .Z(n35952) );
  XNOR U34487 ( .A(q[8]), .B(DB[203]), .Z(n34550) );
  XNOR U34488 ( .A(q[11]), .B(DB[206]), .Z(n34548) );
  IV U34489 ( .A(n34547), .Z(n35951) );
  XNOR U34490 ( .A(n34545), .B(n35953), .Z(n34547) );
  XNOR U34491 ( .A(q[10]), .B(DB[205]), .Z(n35953) );
  XNOR U34492 ( .A(q[9]), .B(DB[204]), .Z(n34545) );
  IV U34493 ( .A(n34560), .Z(n35947) );
  XOR U34494 ( .A(n35954), .B(n35955), .Z(n34560) );
  XNOR U34495 ( .A(n34577), .B(n34558), .Z(n35955) );
  XNOR U34496 ( .A(q[0]), .B(DB[195]), .Z(n34558) );
  XOR U34497 ( .A(n35956), .B(n34566), .Z(n34577) );
  XNOR U34498 ( .A(q[7]), .B(DB[202]), .Z(n34566) );
  IV U34499 ( .A(n34565), .Z(n35956) );
  XNOR U34500 ( .A(n34563), .B(n35957), .Z(n34565) );
  XNOR U34501 ( .A(q[6]), .B(DB[201]), .Z(n35957) );
  XNOR U34502 ( .A(q[5]), .B(DB[200]), .Z(n34563) );
  IV U34503 ( .A(n34576), .Z(n35954) );
  XOR U34504 ( .A(n35958), .B(n35959), .Z(n34576) );
  XNOR U34505 ( .A(n34572), .B(n34574), .Z(n35959) );
  XNOR U34506 ( .A(q[1]), .B(DB[196]), .Z(n34574) );
  XNOR U34507 ( .A(q[4]), .B(DB[199]), .Z(n34572) );
  IV U34508 ( .A(n34571), .Z(n35958) );
  XNOR U34509 ( .A(n34569), .B(n35960), .Z(n34571) );
  XNOR U34510 ( .A(q[3]), .B(DB[198]), .Z(n35960) );
  XNOR U34511 ( .A(q[2]), .B(DB[197]), .Z(n34569) );
  XOR U34512 ( .A(n35961), .B(n34467), .Z(n34395) );
  XOR U34513 ( .A(n35962), .B(n34459), .Z(n34467) );
  XOR U34514 ( .A(n35963), .B(n34448), .Z(n34459) );
  XNOR U34515 ( .A(q[14]), .B(DB[224]), .Z(n34448) );
  IV U34516 ( .A(n34447), .Z(n35963) );
  XNOR U34517 ( .A(n34445), .B(n35964), .Z(n34447) );
  XNOR U34518 ( .A(q[13]), .B(DB[223]), .Z(n35964) );
  XNOR U34519 ( .A(q[12]), .B(DB[222]), .Z(n34445) );
  IV U34520 ( .A(n34458), .Z(n35962) );
  XOR U34521 ( .A(n35965), .B(n35966), .Z(n34458) );
  XNOR U34522 ( .A(n34454), .B(n34456), .Z(n35966) );
  XNOR U34523 ( .A(q[8]), .B(DB[218]), .Z(n34456) );
  XNOR U34524 ( .A(q[11]), .B(DB[221]), .Z(n34454) );
  IV U34525 ( .A(n34453), .Z(n35965) );
  XNOR U34526 ( .A(n34451), .B(n35967), .Z(n34453) );
  XNOR U34527 ( .A(q[10]), .B(DB[220]), .Z(n35967) );
  XNOR U34528 ( .A(q[9]), .B(DB[219]), .Z(n34451) );
  IV U34529 ( .A(n34466), .Z(n35961) );
  XOR U34530 ( .A(n35968), .B(n35969), .Z(n34466) );
  XNOR U34531 ( .A(n34483), .B(n34464), .Z(n35969) );
  XNOR U34532 ( .A(q[0]), .B(DB[210]), .Z(n34464) );
  XOR U34533 ( .A(n35970), .B(n34472), .Z(n34483) );
  XNOR U34534 ( .A(q[7]), .B(DB[217]), .Z(n34472) );
  IV U34535 ( .A(n34471), .Z(n35970) );
  XNOR U34536 ( .A(n34469), .B(n35971), .Z(n34471) );
  XNOR U34537 ( .A(q[6]), .B(DB[216]), .Z(n35971) );
  XNOR U34538 ( .A(q[5]), .B(DB[215]), .Z(n34469) );
  IV U34539 ( .A(n34482), .Z(n35968) );
  XOR U34540 ( .A(n35972), .B(n35973), .Z(n34482) );
  XNOR U34541 ( .A(n34478), .B(n34480), .Z(n35973) );
  XNOR U34542 ( .A(q[1]), .B(DB[211]), .Z(n34480) );
  XNOR U34543 ( .A(q[4]), .B(DB[214]), .Z(n34478) );
  IV U34544 ( .A(n34477), .Z(n35972) );
  XNOR U34545 ( .A(n34475), .B(n35974), .Z(n34477) );
  XNOR U34546 ( .A(q[3]), .B(DB[213]), .Z(n35974) );
  XNOR U34547 ( .A(q[2]), .B(DB[212]), .Z(n34475) );
  XOR U34548 ( .A(n35975), .B(n34373), .Z(n34301) );
  XOR U34549 ( .A(n35976), .B(n34365), .Z(n34373) );
  XOR U34550 ( .A(n35977), .B(n34354), .Z(n34365) );
  XNOR U34551 ( .A(q[14]), .B(DB[239]), .Z(n34354) );
  IV U34552 ( .A(n34353), .Z(n35977) );
  XNOR U34553 ( .A(n34351), .B(n35978), .Z(n34353) );
  XNOR U34554 ( .A(q[13]), .B(DB[238]), .Z(n35978) );
  XNOR U34555 ( .A(q[12]), .B(DB[237]), .Z(n34351) );
  IV U34556 ( .A(n34364), .Z(n35976) );
  XOR U34557 ( .A(n35979), .B(n35980), .Z(n34364) );
  XNOR U34558 ( .A(n34360), .B(n34362), .Z(n35980) );
  XNOR U34559 ( .A(q[8]), .B(DB[233]), .Z(n34362) );
  XNOR U34560 ( .A(q[11]), .B(DB[236]), .Z(n34360) );
  IV U34561 ( .A(n34359), .Z(n35979) );
  XNOR U34562 ( .A(n34357), .B(n35981), .Z(n34359) );
  XNOR U34563 ( .A(q[10]), .B(DB[235]), .Z(n35981) );
  XNOR U34564 ( .A(q[9]), .B(DB[234]), .Z(n34357) );
  IV U34565 ( .A(n34372), .Z(n35975) );
  XOR U34566 ( .A(n35982), .B(n35983), .Z(n34372) );
  XNOR U34567 ( .A(n34389), .B(n34370), .Z(n35983) );
  XNOR U34568 ( .A(q[0]), .B(DB[225]), .Z(n34370) );
  XOR U34569 ( .A(n35984), .B(n34378), .Z(n34389) );
  XNOR U34570 ( .A(q[7]), .B(DB[232]), .Z(n34378) );
  IV U34571 ( .A(n34377), .Z(n35984) );
  XNOR U34572 ( .A(n34375), .B(n35985), .Z(n34377) );
  XNOR U34573 ( .A(q[6]), .B(DB[231]), .Z(n35985) );
  XNOR U34574 ( .A(q[5]), .B(DB[230]), .Z(n34375) );
  IV U34575 ( .A(n34388), .Z(n35982) );
  XOR U34576 ( .A(n35986), .B(n35987), .Z(n34388) );
  XNOR U34577 ( .A(n34384), .B(n34386), .Z(n35987) );
  XNOR U34578 ( .A(q[1]), .B(DB[226]), .Z(n34386) );
  XNOR U34579 ( .A(q[4]), .B(DB[229]), .Z(n34384) );
  IV U34580 ( .A(n34383), .Z(n35986) );
  XNOR U34581 ( .A(n34381), .B(n35988), .Z(n34383) );
  XNOR U34582 ( .A(q[3]), .B(DB[228]), .Z(n35988) );
  XNOR U34583 ( .A(q[2]), .B(DB[227]), .Z(n34381) );
  XOR U34584 ( .A(n35989), .B(n34279), .Z(n34207) );
  XOR U34585 ( .A(n35990), .B(n34271), .Z(n34279) );
  XOR U34586 ( .A(n35991), .B(n34260), .Z(n34271) );
  XNOR U34587 ( .A(q[14]), .B(DB[254]), .Z(n34260) );
  IV U34588 ( .A(n34259), .Z(n35991) );
  XNOR U34589 ( .A(n34257), .B(n35992), .Z(n34259) );
  XNOR U34590 ( .A(q[13]), .B(DB[253]), .Z(n35992) );
  XNOR U34591 ( .A(q[12]), .B(DB[252]), .Z(n34257) );
  IV U34592 ( .A(n34270), .Z(n35990) );
  XOR U34593 ( .A(n35993), .B(n35994), .Z(n34270) );
  XNOR U34594 ( .A(n34266), .B(n34268), .Z(n35994) );
  XNOR U34595 ( .A(q[8]), .B(DB[248]), .Z(n34268) );
  XNOR U34596 ( .A(q[11]), .B(DB[251]), .Z(n34266) );
  IV U34597 ( .A(n34265), .Z(n35993) );
  XNOR U34598 ( .A(n34263), .B(n35995), .Z(n34265) );
  XNOR U34599 ( .A(q[10]), .B(DB[250]), .Z(n35995) );
  XNOR U34600 ( .A(q[9]), .B(DB[249]), .Z(n34263) );
  IV U34601 ( .A(n34278), .Z(n35989) );
  XOR U34602 ( .A(n35996), .B(n35997), .Z(n34278) );
  XNOR U34603 ( .A(n34295), .B(n34276), .Z(n35997) );
  XNOR U34604 ( .A(q[0]), .B(DB[240]), .Z(n34276) );
  XOR U34605 ( .A(n35998), .B(n34284), .Z(n34295) );
  XNOR U34606 ( .A(q[7]), .B(DB[247]), .Z(n34284) );
  IV U34607 ( .A(n34283), .Z(n35998) );
  XNOR U34608 ( .A(n34281), .B(n35999), .Z(n34283) );
  XNOR U34609 ( .A(q[6]), .B(DB[246]), .Z(n35999) );
  XNOR U34610 ( .A(q[5]), .B(DB[245]), .Z(n34281) );
  IV U34611 ( .A(n34294), .Z(n35996) );
  XOR U34612 ( .A(n36000), .B(n36001), .Z(n34294) );
  XNOR U34613 ( .A(n34290), .B(n34292), .Z(n36001) );
  XNOR U34614 ( .A(q[1]), .B(DB[241]), .Z(n34292) );
  XNOR U34615 ( .A(q[4]), .B(DB[244]), .Z(n34290) );
  IV U34616 ( .A(n34289), .Z(n36000) );
  XNOR U34617 ( .A(n34287), .B(n36002), .Z(n34289) );
  XNOR U34618 ( .A(q[3]), .B(DB[243]), .Z(n36002) );
  XNOR U34619 ( .A(q[2]), .B(DB[242]), .Z(n34287) );
  XOR U34620 ( .A(n36003), .B(n34185), .Z(n34113) );
  XOR U34621 ( .A(n36004), .B(n34177), .Z(n34185) );
  XOR U34622 ( .A(n36005), .B(n34166), .Z(n34177) );
  XNOR U34623 ( .A(q[14]), .B(DB[269]), .Z(n34166) );
  IV U34624 ( .A(n34165), .Z(n36005) );
  XNOR U34625 ( .A(n34163), .B(n36006), .Z(n34165) );
  XNOR U34626 ( .A(q[13]), .B(DB[268]), .Z(n36006) );
  XNOR U34627 ( .A(q[12]), .B(DB[267]), .Z(n34163) );
  IV U34628 ( .A(n34176), .Z(n36004) );
  XOR U34629 ( .A(n36007), .B(n36008), .Z(n34176) );
  XNOR U34630 ( .A(n34172), .B(n34174), .Z(n36008) );
  XNOR U34631 ( .A(q[8]), .B(DB[263]), .Z(n34174) );
  XNOR U34632 ( .A(q[11]), .B(DB[266]), .Z(n34172) );
  IV U34633 ( .A(n34171), .Z(n36007) );
  XNOR U34634 ( .A(n34169), .B(n36009), .Z(n34171) );
  XNOR U34635 ( .A(q[10]), .B(DB[265]), .Z(n36009) );
  XNOR U34636 ( .A(q[9]), .B(DB[264]), .Z(n34169) );
  IV U34637 ( .A(n34184), .Z(n36003) );
  XOR U34638 ( .A(n36010), .B(n36011), .Z(n34184) );
  XNOR U34639 ( .A(n34201), .B(n34182), .Z(n36011) );
  XNOR U34640 ( .A(q[0]), .B(DB[255]), .Z(n34182) );
  XOR U34641 ( .A(n36012), .B(n34190), .Z(n34201) );
  XNOR U34642 ( .A(q[7]), .B(DB[262]), .Z(n34190) );
  IV U34643 ( .A(n34189), .Z(n36012) );
  XNOR U34644 ( .A(n34187), .B(n36013), .Z(n34189) );
  XNOR U34645 ( .A(q[6]), .B(DB[261]), .Z(n36013) );
  XNOR U34646 ( .A(q[5]), .B(DB[260]), .Z(n34187) );
  IV U34647 ( .A(n34200), .Z(n36010) );
  XOR U34648 ( .A(n36014), .B(n36015), .Z(n34200) );
  XNOR U34649 ( .A(n34196), .B(n34198), .Z(n36015) );
  XNOR U34650 ( .A(q[1]), .B(DB[256]), .Z(n34198) );
  XNOR U34651 ( .A(q[4]), .B(DB[259]), .Z(n34196) );
  IV U34652 ( .A(n34195), .Z(n36014) );
  XNOR U34653 ( .A(n34193), .B(n36016), .Z(n34195) );
  XNOR U34654 ( .A(q[3]), .B(DB[258]), .Z(n36016) );
  XNOR U34655 ( .A(q[2]), .B(DB[257]), .Z(n34193) );
  XOR U34656 ( .A(n36017), .B(n34091), .Z(n34019) );
  XOR U34657 ( .A(n36018), .B(n34083), .Z(n34091) );
  XOR U34658 ( .A(n36019), .B(n34072), .Z(n34083) );
  XNOR U34659 ( .A(q[14]), .B(DB[284]), .Z(n34072) );
  IV U34660 ( .A(n34071), .Z(n36019) );
  XNOR U34661 ( .A(n34069), .B(n36020), .Z(n34071) );
  XNOR U34662 ( .A(q[13]), .B(DB[283]), .Z(n36020) );
  XNOR U34663 ( .A(q[12]), .B(DB[282]), .Z(n34069) );
  IV U34664 ( .A(n34082), .Z(n36018) );
  XOR U34665 ( .A(n36021), .B(n36022), .Z(n34082) );
  XNOR U34666 ( .A(n34078), .B(n34080), .Z(n36022) );
  XNOR U34667 ( .A(q[8]), .B(DB[278]), .Z(n34080) );
  XNOR U34668 ( .A(q[11]), .B(DB[281]), .Z(n34078) );
  IV U34669 ( .A(n34077), .Z(n36021) );
  XNOR U34670 ( .A(n34075), .B(n36023), .Z(n34077) );
  XNOR U34671 ( .A(q[10]), .B(DB[280]), .Z(n36023) );
  XNOR U34672 ( .A(q[9]), .B(DB[279]), .Z(n34075) );
  IV U34673 ( .A(n34090), .Z(n36017) );
  XOR U34674 ( .A(n36024), .B(n36025), .Z(n34090) );
  XNOR U34675 ( .A(n34107), .B(n34088), .Z(n36025) );
  XNOR U34676 ( .A(q[0]), .B(DB[270]), .Z(n34088) );
  XOR U34677 ( .A(n36026), .B(n34096), .Z(n34107) );
  XNOR U34678 ( .A(q[7]), .B(DB[277]), .Z(n34096) );
  IV U34679 ( .A(n34095), .Z(n36026) );
  XNOR U34680 ( .A(n34093), .B(n36027), .Z(n34095) );
  XNOR U34681 ( .A(q[6]), .B(DB[276]), .Z(n36027) );
  XNOR U34682 ( .A(q[5]), .B(DB[275]), .Z(n34093) );
  IV U34683 ( .A(n34106), .Z(n36024) );
  XOR U34684 ( .A(n36028), .B(n36029), .Z(n34106) );
  XNOR U34685 ( .A(n34102), .B(n34104), .Z(n36029) );
  XNOR U34686 ( .A(q[1]), .B(DB[271]), .Z(n34104) );
  XNOR U34687 ( .A(q[4]), .B(DB[274]), .Z(n34102) );
  IV U34688 ( .A(n34101), .Z(n36028) );
  XNOR U34689 ( .A(n34099), .B(n36030), .Z(n34101) );
  XNOR U34690 ( .A(q[3]), .B(DB[273]), .Z(n36030) );
  XNOR U34691 ( .A(q[2]), .B(DB[272]), .Z(n34099) );
  XOR U34692 ( .A(n36031), .B(n33997), .Z(n33925) );
  XOR U34693 ( .A(n36032), .B(n33989), .Z(n33997) );
  XOR U34694 ( .A(n36033), .B(n33978), .Z(n33989) );
  XNOR U34695 ( .A(q[14]), .B(DB[299]), .Z(n33978) );
  IV U34696 ( .A(n33977), .Z(n36033) );
  XNOR U34697 ( .A(n33975), .B(n36034), .Z(n33977) );
  XNOR U34698 ( .A(q[13]), .B(DB[298]), .Z(n36034) );
  XNOR U34699 ( .A(q[12]), .B(DB[297]), .Z(n33975) );
  IV U34700 ( .A(n33988), .Z(n36032) );
  XOR U34701 ( .A(n36035), .B(n36036), .Z(n33988) );
  XNOR U34702 ( .A(n33984), .B(n33986), .Z(n36036) );
  XNOR U34703 ( .A(q[8]), .B(DB[293]), .Z(n33986) );
  XNOR U34704 ( .A(q[11]), .B(DB[296]), .Z(n33984) );
  IV U34705 ( .A(n33983), .Z(n36035) );
  XNOR U34706 ( .A(n33981), .B(n36037), .Z(n33983) );
  XNOR U34707 ( .A(q[10]), .B(DB[295]), .Z(n36037) );
  XNOR U34708 ( .A(q[9]), .B(DB[294]), .Z(n33981) );
  IV U34709 ( .A(n33996), .Z(n36031) );
  XOR U34710 ( .A(n36038), .B(n36039), .Z(n33996) );
  XNOR U34711 ( .A(n34013), .B(n33994), .Z(n36039) );
  XNOR U34712 ( .A(q[0]), .B(DB[285]), .Z(n33994) );
  XOR U34713 ( .A(n36040), .B(n34002), .Z(n34013) );
  XNOR U34714 ( .A(q[7]), .B(DB[292]), .Z(n34002) );
  IV U34715 ( .A(n34001), .Z(n36040) );
  XNOR U34716 ( .A(n33999), .B(n36041), .Z(n34001) );
  XNOR U34717 ( .A(q[6]), .B(DB[291]), .Z(n36041) );
  XNOR U34718 ( .A(q[5]), .B(DB[290]), .Z(n33999) );
  IV U34719 ( .A(n34012), .Z(n36038) );
  XOR U34720 ( .A(n36042), .B(n36043), .Z(n34012) );
  XNOR U34721 ( .A(n34008), .B(n34010), .Z(n36043) );
  XNOR U34722 ( .A(q[1]), .B(DB[286]), .Z(n34010) );
  XNOR U34723 ( .A(q[4]), .B(DB[289]), .Z(n34008) );
  IV U34724 ( .A(n34007), .Z(n36042) );
  XNOR U34725 ( .A(n34005), .B(n36044), .Z(n34007) );
  XNOR U34726 ( .A(q[3]), .B(DB[288]), .Z(n36044) );
  XNOR U34727 ( .A(q[2]), .B(DB[287]), .Z(n34005) );
  XOR U34728 ( .A(n36045), .B(n33903), .Z(n33831) );
  XOR U34729 ( .A(n36046), .B(n33895), .Z(n33903) );
  XOR U34730 ( .A(n36047), .B(n33884), .Z(n33895) );
  XNOR U34731 ( .A(q[14]), .B(DB[314]), .Z(n33884) );
  IV U34732 ( .A(n33883), .Z(n36047) );
  XNOR U34733 ( .A(n33881), .B(n36048), .Z(n33883) );
  XNOR U34734 ( .A(q[13]), .B(DB[313]), .Z(n36048) );
  XNOR U34735 ( .A(q[12]), .B(DB[312]), .Z(n33881) );
  IV U34736 ( .A(n33894), .Z(n36046) );
  XOR U34737 ( .A(n36049), .B(n36050), .Z(n33894) );
  XNOR U34738 ( .A(n33890), .B(n33892), .Z(n36050) );
  XNOR U34739 ( .A(q[8]), .B(DB[308]), .Z(n33892) );
  XNOR U34740 ( .A(q[11]), .B(DB[311]), .Z(n33890) );
  IV U34741 ( .A(n33889), .Z(n36049) );
  XNOR U34742 ( .A(n33887), .B(n36051), .Z(n33889) );
  XNOR U34743 ( .A(q[10]), .B(DB[310]), .Z(n36051) );
  XNOR U34744 ( .A(q[9]), .B(DB[309]), .Z(n33887) );
  IV U34745 ( .A(n33902), .Z(n36045) );
  XOR U34746 ( .A(n36052), .B(n36053), .Z(n33902) );
  XNOR U34747 ( .A(n33919), .B(n33900), .Z(n36053) );
  XNOR U34748 ( .A(q[0]), .B(DB[300]), .Z(n33900) );
  XOR U34749 ( .A(n36054), .B(n33908), .Z(n33919) );
  XNOR U34750 ( .A(q[7]), .B(DB[307]), .Z(n33908) );
  IV U34751 ( .A(n33907), .Z(n36054) );
  XNOR U34752 ( .A(n33905), .B(n36055), .Z(n33907) );
  XNOR U34753 ( .A(q[6]), .B(DB[306]), .Z(n36055) );
  XNOR U34754 ( .A(q[5]), .B(DB[305]), .Z(n33905) );
  IV U34755 ( .A(n33918), .Z(n36052) );
  XOR U34756 ( .A(n36056), .B(n36057), .Z(n33918) );
  XNOR U34757 ( .A(n33914), .B(n33916), .Z(n36057) );
  XNOR U34758 ( .A(q[1]), .B(DB[301]), .Z(n33916) );
  XNOR U34759 ( .A(q[4]), .B(DB[304]), .Z(n33914) );
  IV U34760 ( .A(n33913), .Z(n36056) );
  XNOR U34761 ( .A(n33911), .B(n36058), .Z(n33913) );
  XNOR U34762 ( .A(q[3]), .B(DB[303]), .Z(n36058) );
  XNOR U34763 ( .A(q[2]), .B(DB[302]), .Z(n33911) );
  XOR U34764 ( .A(n36059), .B(n33809), .Z(n33737) );
  XOR U34765 ( .A(n36060), .B(n33801), .Z(n33809) );
  XOR U34766 ( .A(n36061), .B(n33790), .Z(n33801) );
  XNOR U34767 ( .A(q[14]), .B(DB[329]), .Z(n33790) );
  IV U34768 ( .A(n33789), .Z(n36061) );
  XNOR U34769 ( .A(n33787), .B(n36062), .Z(n33789) );
  XNOR U34770 ( .A(q[13]), .B(DB[328]), .Z(n36062) );
  XNOR U34771 ( .A(q[12]), .B(DB[327]), .Z(n33787) );
  IV U34772 ( .A(n33800), .Z(n36060) );
  XOR U34773 ( .A(n36063), .B(n36064), .Z(n33800) );
  XNOR U34774 ( .A(n33796), .B(n33798), .Z(n36064) );
  XNOR U34775 ( .A(q[8]), .B(DB[323]), .Z(n33798) );
  XNOR U34776 ( .A(q[11]), .B(DB[326]), .Z(n33796) );
  IV U34777 ( .A(n33795), .Z(n36063) );
  XNOR U34778 ( .A(n33793), .B(n36065), .Z(n33795) );
  XNOR U34779 ( .A(q[10]), .B(DB[325]), .Z(n36065) );
  XNOR U34780 ( .A(q[9]), .B(DB[324]), .Z(n33793) );
  IV U34781 ( .A(n33808), .Z(n36059) );
  XOR U34782 ( .A(n36066), .B(n36067), .Z(n33808) );
  XNOR U34783 ( .A(n33825), .B(n33806), .Z(n36067) );
  XNOR U34784 ( .A(q[0]), .B(DB[315]), .Z(n33806) );
  XOR U34785 ( .A(n36068), .B(n33814), .Z(n33825) );
  XNOR U34786 ( .A(q[7]), .B(DB[322]), .Z(n33814) );
  IV U34787 ( .A(n33813), .Z(n36068) );
  XNOR U34788 ( .A(n33811), .B(n36069), .Z(n33813) );
  XNOR U34789 ( .A(q[6]), .B(DB[321]), .Z(n36069) );
  XNOR U34790 ( .A(q[5]), .B(DB[320]), .Z(n33811) );
  IV U34791 ( .A(n33824), .Z(n36066) );
  XOR U34792 ( .A(n36070), .B(n36071), .Z(n33824) );
  XNOR U34793 ( .A(n33820), .B(n33822), .Z(n36071) );
  XNOR U34794 ( .A(q[1]), .B(DB[316]), .Z(n33822) );
  XNOR U34795 ( .A(q[4]), .B(DB[319]), .Z(n33820) );
  IV U34796 ( .A(n33819), .Z(n36070) );
  XNOR U34797 ( .A(n33817), .B(n36072), .Z(n33819) );
  XNOR U34798 ( .A(q[3]), .B(DB[318]), .Z(n36072) );
  XNOR U34799 ( .A(q[2]), .B(DB[317]), .Z(n33817) );
  XOR U34800 ( .A(n36073), .B(n33715), .Z(n33643) );
  XOR U34801 ( .A(n36074), .B(n33707), .Z(n33715) );
  XOR U34802 ( .A(n36075), .B(n33696), .Z(n33707) );
  XNOR U34803 ( .A(q[14]), .B(DB[344]), .Z(n33696) );
  IV U34804 ( .A(n33695), .Z(n36075) );
  XNOR U34805 ( .A(n33693), .B(n36076), .Z(n33695) );
  XNOR U34806 ( .A(q[13]), .B(DB[343]), .Z(n36076) );
  XNOR U34807 ( .A(q[12]), .B(DB[342]), .Z(n33693) );
  IV U34808 ( .A(n33706), .Z(n36074) );
  XOR U34809 ( .A(n36077), .B(n36078), .Z(n33706) );
  XNOR U34810 ( .A(n33702), .B(n33704), .Z(n36078) );
  XNOR U34811 ( .A(q[8]), .B(DB[338]), .Z(n33704) );
  XNOR U34812 ( .A(q[11]), .B(DB[341]), .Z(n33702) );
  IV U34813 ( .A(n33701), .Z(n36077) );
  XNOR U34814 ( .A(n33699), .B(n36079), .Z(n33701) );
  XNOR U34815 ( .A(q[10]), .B(DB[340]), .Z(n36079) );
  XNOR U34816 ( .A(q[9]), .B(DB[339]), .Z(n33699) );
  IV U34817 ( .A(n33714), .Z(n36073) );
  XOR U34818 ( .A(n36080), .B(n36081), .Z(n33714) );
  XNOR U34819 ( .A(n33731), .B(n33712), .Z(n36081) );
  XNOR U34820 ( .A(q[0]), .B(DB[330]), .Z(n33712) );
  XOR U34821 ( .A(n36082), .B(n33720), .Z(n33731) );
  XNOR U34822 ( .A(q[7]), .B(DB[337]), .Z(n33720) );
  IV U34823 ( .A(n33719), .Z(n36082) );
  XNOR U34824 ( .A(n33717), .B(n36083), .Z(n33719) );
  XNOR U34825 ( .A(q[6]), .B(DB[336]), .Z(n36083) );
  XNOR U34826 ( .A(q[5]), .B(DB[335]), .Z(n33717) );
  IV U34827 ( .A(n33730), .Z(n36080) );
  XOR U34828 ( .A(n36084), .B(n36085), .Z(n33730) );
  XNOR U34829 ( .A(n33726), .B(n33728), .Z(n36085) );
  XNOR U34830 ( .A(q[1]), .B(DB[331]), .Z(n33728) );
  XNOR U34831 ( .A(q[4]), .B(DB[334]), .Z(n33726) );
  IV U34832 ( .A(n33725), .Z(n36084) );
  XNOR U34833 ( .A(n33723), .B(n36086), .Z(n33725) );
  XNOR U34834 ( .A(q[3]), .B(DB[333]), .Z(n36086) );
  XNOR U34835 ( .A(q[2]), .B(DB[332]), .Z(n33723) );
  XOR U34836 ( .A(n36087), .B(n33621), .Z(n33549) );
  XOR U34837 ( .A(n36088), .B(n33613), .Z(n33621) );
  XOR U34838 ( .A(n36089), .B(n33602), .Z(n33613) );
  XNOR U34839 ( .A(q[14]), .B(DB[359]), .Z(n33602) );
  IV U34840 ( .A(n33601), .Z(n36089) );
  XNOR U34841 ( .A(n33599), .B(n36090), .Z(n33601) );
  XNOR U34842 ( .A(q[13]), .B(DB[358]), .Z(n36090) );
  XNOR U34843 ( .A(q[12]), .B(DB[357]), .Z(n33599) );
  IV U34844 ( .A(n33612), .Z(n36088) );
  XOR U34845 ( .A(n36091), .B(n36092), .Z(n33612) );
  XNOR U34846 ( .A(n33608), .B(n33610), .Z(n36092) );
  XNOR U34847 ( .A(q[8]), .B(DB[353]), .Z(n33610) );
  XNOR U34848 ( .A(q[11]), .B(DB[356]), .Z(n33608) );
  IV U34849 ( .A(n33607), .Z(n36091) );
  XNOR U34850 ( .A(n33605), .B(n36093), .Z(n33607) );
  XNOR U34851 ( .A(q[10]), .B(DB[355]), .Z(n36093) );
  XNOR U34852 ( .A(q[9]), .B(DB[354]), .Z(n33605) );
  IV U34853 ( .A(n33620), .Z(n36087) );
  XOR U34854 ( .A(n36094), .B(n36095), .Z(n33620) );
  XNOR U34855 ( .A(n33637), .B(n33618), .Z(n36095) );
  XNOR U34856 ( .A(q[0]), .B(DB[345]), .Z(n33618) );
  XOR U34857 ( .A(n36096), .B(n33626), .Z(n33637) );
  XNOR U34858 ( .A(q[7]), .B(DB[352]), .Z(n33626) );
  IV U34859 ( .A(n33625), .Z(n36096) );
  XNOR U34860 ( .A(n33623), .B(n36097), .Z(n33625) );
  XNOR U34861 ( .A(q[6]), .B(DB[351]), .Z(n36097) );
  XNOR U34862 ( .A(q[5]), .B(DB[350]), .Z(n33623) );
  IV U34863 ( .A(n33636), .Z(n36094) );
  XOR U34864 ( .A(n36098), .B(n36099), .Z(n33636) );
  XNOR U34865 ( .A(n33632), .B(n33634), .Z(n36099) );
  XNOR U34866 ( .A(q[1]), .B(DB[346]), .Z(n33634) );
  XNOR U34867 ( .A(q[4]), .B(DB[349]), .Z(n33632) );
  IV U34868 ( .A(n33631), .Z(n36098) );
  XNOR U34869 ( .A(n33629), .B(n36100), .Z(n33631) );
  XNOR U34870 ( .A(q[3]), .B(DB[348]), .Z(n36100) );
  XNOR U34871 ( .A(q[2]), .B(DB[347]), .Z(n33629) );
  XOR U34872 ( .A(n36101), .B(n33527), .Z(n33455) );
  XOR U34873 ( .A(n36102), .B(n33519), .Z(n33527) );
  XOR U34874 ( .A(n36103), .B(n33508), .Z(n33519) );
  XNOR U34875 ( .A(q[14]), .B(DB[374]), .Z(n33508) );
  IV U34876 ( .A(n33507), .Z(n36103) );
  XNOR U34877 ( .A(n33505), .B(n36104), .Z(n33507) );
  XNOR U34878 ( .A(q[13]), .B(DB[373]), .Z(n36104) );
  XNOR U34879 ( .A(q[12]), .B(DB[372]), .Z(n33505) );
  IV U34880 ( .A(n33518), .Z(n36102) );
  XOR U34881 ( .A(n36105), .B(n36106), .Z(n33518) );
  XNOR U34882 ( .A(n33514), .B(n33516), .Z(n36106) );
  XNOR U34883 ( .A(q[8]), .B(DB[368]), .Z(n33516) );
  XNOR U34884 ( .A(q[11]), .B(DB[371]), .Z(n33514) );
  IV U34885 ( .A(n33513), .Z(n36105) );
  XNOR U34886 ( .A(n33511), .B(n36107), .Z(n33513) );
  XNOR U34887 ( .A(q[10]), .B(DB[370]), .Z(n36107) );
  XNOR U34888 ( .A(q[9]), .B(DB[369]), .Z(n33511) );
  IV U34889 ( .A(n33526), .Z(n36101) );
  XOR U34890 ( .A(n36108), .B(n36109), .Z(n33526) );
  XNOR U34891 ( .A(n33543), .B(n33524), .Z(n36109) );
  XNOR U34892 ( .A(q[0]), .B(DB[360]), .Z(n33524) );
  XOR U34893 ( .A(n36110), .B(n33532), .Z(n33543) );
  XNOR U34894 ( .A(q[7]), .B(DB[367]), .Z(n33532) );
  IV U34895 ( .A(n33531), .Z(n36110) );
  XNOR U34896 ( .A(n33529), .B(n36111), .Z(n33531) );
  XNOR U34897 ( .A(q[6]), .B(DB[366]), .Z(n36111) );
  XNOR U34898 ( .A(q[5]), .B(DB[365]), .Z(n33529) );
  IV U34899 ( .A(n33542), .Z(n36108) );
  XOR U34900 ( .A(n36112), .B(n36113), .Z(n33542) );
  XNOR U34901 ( .A(n33538), .B(n33540), .Z(n36113) );
  XNOR U34902 ( .A(q[1]), .B(DB[361]), .Z(n33540) );
  XNOR U34903 ( .A(q[4]), .B(DB[364]), .Z(n33538) );
  IV U34904 ( .A(n33537), .Z(n36112) );
  XNOR U34905 ( .A(n33535), .B(n36114), .Z(n33537) );
  XNOR U34906 ( .A(q[3]), .B(DB[363]), .Z(n36114) );
  XNOR U34907 ( .A(q[2]), .B(DB[362]), .Z(n33535) );
  XOR U34908 ( .A(n36115), .B(n33433), .Z(n33361) );
  XOR U34909 ( .A(n36116), .B(n33425), .Z(n33433) );
  XOR U34910 ( .A(n36117), .B(n33414), .Z(n33425) );
  XNOR U34911 ( .A(q[14]), .B(DB[389]), .Z(n33414) );
  IV U34912 ( .A(n33413), .Z(n36117) );
  XNOR U34913 ( .A(n33411), .B(n36118), .Z(n33413) );
  XNOR U34914 ( .A(q[13]), .B(DB[388]), .Z(n36118) );
  XNOR U34915 ( .A(q[12]), .B(DB[387]), .Z(n33411) );
  IV U34916 ( .A(n33424), .Z(n36116) );
  XOR U34917 ( .A(n36119), .B(n36120), .Z(n33424) );
  XNOR U34918 ( .A(n33420), .B(n33422), .Z(n36120) );
  XNOR U34919 ( .A(q[8]), .B(DB[383]), .Z(n33422) );
  XNOR U34920 ( .A(q[11]), .B(DB[386]), .Z(n33420) );
  IV U34921 ( .A(n33419), .Z(n36119) );
  XNOR U34922 ( .A(n33417), .B(n36121), .Z(n33419) );
  XNOR U34923 ( .A(q[10]), .B(DB[385]), .Z(n36121) );
  XNOR U34924 ( .A(q[9]), .B(DB[384]), .Z(n33417) );
  IV U34925 ( .A(n33432), .Z(n36115) );
  XOR U34926 ( .A(n36122), .B(n36123), .Z(n33432) );
  XNOR U34927 ( .A(n33449), .B(n33430), .Z(n36123) );
  XNOR U34928 ( .A(q[0]), .B(DB[375]), .Z(n33430) );
  XOR U34929 ( .A(n36124), .B(n33438), .Z(n33449) );
  XNOR U34930 ( .A(q[7]), .B(DB[382]), .Z(n33438) );
  IV U34931 ( .A(n33437), .Z(n36124) );
  XNOR U34932 ( .A(n33435), .B(n36125), .Z(n33437) );
  XNOR U34933 ( .A(q[6]), .B(DB[381]), .Z(n36125) );
  XNOR U34934 ( .A(q[5]), .B(DB[380]), .Z(n33435) );
  IV U34935 ( .A(n33448), .Z(n36122) );
  XOR U34936 ( .A(n36126), .B(n36127), .Z(n33448) );
  XNOR U34937 ( .A(n33444), .B(n33446), .Z(n36127) );
  XNOR U34938 ( .A(q[1]), .B(DB[376]), .Z(n33446) );
  XNOR U34939 ( .A(q[4]), .B(DB[379]), .Z(n33444) );
  IV U34940 ( .A(n33443), .Z(n36126) );
  XNOR U34941 ( .A(n33441), .B(n36128), .Z(n33443) );
  XNOR U34942 ( .A(q[3]), .B(DB[378]), .Z(n36128) );
  XNOR U34943 ( .A(q[2]), .B(DB[377]), .Z(n33441) );
  XOR U34944 ( .A(n36129), .B(n33339), .Z(n33267) );
  XOR U34945 ( .A(n36130), .B(n33331), .Z(n33339) );
  XOR U34946 ( .A(n36131), .B(n33320), .Z(n33331) );
  XNOR U34947 ( .A(q[14]), .B(DB[404]), .Z(n33320) );
  IV U34948 ( .A(n33319), .Z(n36131) );
  XNOR U34949 ( .A(n33317), .B(n36132), .Z(n33319) );
  XNOR U34950 ( .A(q[13]), .B(DB[403]), .Z(n36132) );
  XNOR U34951 ( .A(q[12]), .B(DB[402]), .Z(n33317) );
  IV U34952 ( .A(n33330), .Z(n36130) );
  XOR U34953 ( .A(n36133), .B(n36134), .Z(n33330) );
  XNOR U34954 ( .A(n33326), .B(n33328), .Z(n36134) );
  XNOR U34955 ( .A(q[8]), .B(DB[398]), .Z(n33328) );
  XNOR U34956 ( .A(q[11]), .B(DB[401]), .Z(n33326) );
  IV U34957 ( .A(n33325), .Z(n36133) );
  XNOR U34958 ( .A(n33323), .B(n36135), .Z(n33325) );
  XNOR U34959 ( .A(q[10]), .B(DB[400]), .Z(n36135) );
  XNOR U34960 ( .A(q[9]), .B(DB[399]), .Z(n33323) );
  IV U34961 ( .A(n33338), .Z(n36129) );
  XOR U34962 ( .A(n36136), .B(n36137), .Z(n33338) );
  XNOR U34963 ( .A(n33355), .B(n33336), .Z(n36137) );
  XNOR U34964 ( .A(q[0]), .B(DB[390]), .Z(n33336) );
  XOR U34965 ( .A(n36138), .B(n33344), .Z(n33355) );
  XNOR U34966 ( .A(q[7]), .B(DB[397]), .Z(n33344) );
  IV U34967 ( .A(n33343), .Z(n36138) );
  XNOR U34968 ( .A(n33341), .B(n36139), .Z(n33343) );
  XNOR U34969 ( .A(q[6]), .B(DB[396]), .Z(n36139) );
  XNOR U34970 ( .A(q[5]), .B(DB[395]), .Z(n33341) );
  IV U34971 ( .A(n33354), .Z(n36136) );
  XOR U34972 ( .A(n36140), .B(n36141), .Z(n33354) );
  XNOR U34973 ( .A(n33350), .B(n33352), .Z(n36141) );
  XNOR U34974 ( .A(q[1]), .B(DB[391]), .Z(n33352) );
  XNOR U34975 ( .A(q[4]), .B(DB[394]), .Z(n33350) );
  IV U34976 ( .A(n33349), .Z(n36140) );
  XNOR U34977 ( .A(n33347), .B(n36142), .Z(n33349) );
  XNOR U34978 ( .A(q[3]), .B(DB[393]), .Z(n36142) );
  XNOR U34979 ( .A(q[2]), .B(DB[392]), .Z(n33347) );
  XOR U34980 ( .A(n36143), .B(n33245), .Z(n33173) );
  XOR U34981 ( .A(n36144), .B(n33237), .Z(n33245) );
  XOR U34982 ( .A(n36145), .B(n33226), .Z(n33237) );
  XNOR U34983 ( .A(q[14]), .B(DB[419]), .Z(n33226) );
  IV U34984 ( .A(n33225), .Z(n36145) );
  XNOR U34985 ( .A(n33223), .B(n36146), .Z(n33225) );
  XNOR U34986 ( .A(q[13]), .B(DB[418]), .Z(n36146) );
  XNOR U34987 ( .A(q[12]), .B(DB[417]), .Z(n33223) );
  IV U34988 ( .A(n33236), .Z(n36144) );
  XOR U34989 ( .A(n36147), .B(n36148), .Z(n33236) );
  XNOR U34990 ( .A(n33232), .B(n33234), .Z(n36148) );
  XNOR U34991 ( .A(q[8]), .B(DB[413]), .Z(n33234) );
  XNOR U34992 ( .A(q[11]), .B(DB[416]), .Z(n33232) );
  IV U34993 ( .A(n33231), .Z(n36147) );
  XNOR U34994 ( .A(n33229), .B(n36149), .Z(n33231) );
  XNOR U34995 ( .A(q[10]), .B(DB[415]), .Z(n36149) );
  XNOR U34996 ( .A(q[9]), .B(DB[414]), .Z(n33229) );
  IV U34997 ( .A(n33244), .Z(n36143) );
  XOR U34998 ( .A(n36150), .B(n36151), .Z(n33244) );
  XNOR U34999 ( .A(n33261), .B(n33242), .Z(n36151) );
  XNOR U35000 ( .A(q[0]), .B(DB[405]), .Z(n33242) );
  XOR U35001 ( .A(n36152), .B(n33250), .Z(n33261) );
  XNOR U35002 ( .A(q[7]), .B(DB[412]), .Z(n33250) );
  IV U35003 ( .A(n33249), .Z(n36152) );
  XNOR U35004 ( .A(n33247), .B(n36153), .Z(n33249) );
  XNOR U35005 ( .A(q[6]), .B(DB[411]), .Z(n36153) );
  XNOR U35006 ( .A(q[5]), .B(DB[410]), .Z(n33247) );
  IV U35007 ( .A(n33260), .Z(n36150) );
  XOR U35008 ( .A(n36154), .B(n36155), .Z(n33260) );
  XNOR U35009 ( .A(n33256), .B(n33258), .Z(n36155) );
  XNOR U35010 ( .A(q[1]), .B(DB[406]), .Z(n33258) );
  XNOR U35011 ( .A(q[4]), .B(DB[409]), .Z(n33256) );
  IV U35012 ( .A(n33255), .Z(n36154) );
  XNOR U35013 ( .A(n33253), .B(n36156), .Z(n33255) );
  XNOR U35014 ( .A(q[3]), .B(DB[408]), .Z(n36156) );
  XNOR U35015 ( .A(q[2]), .B(DB[407]), .Z(n33253) );
  XOR U35016 ( .A(n36157), .B(n33151), .Z(n33079) );
  XOR U35017 ( .A(n36158), .B(n33143), .Z(n33151) );
  XOR U35018 ( .A(n36159), .B(n33132), .Z(n33143) );
  XNOR U35019 ( .A(q[14]), .B(DB[434]), .Z(n33132) );
  IV U35020 ( .A(n33131), .Z(n36159) );
  XNOR U35021 ( .A(n33129), .B(n36160), .Z(n33131) );
  XNOR U35022 ( .A(q[13]), .B(DB[433]), .Z(n36160) );
  XNOR U35023 ( .A(q[12]), .B(DB[432]), .Z(n33129) );
  IV U35024 ( .A(n33142), .Z(n36158) );
  XOR U35025 ( .A(n36161), .B(n36162), .Z(n33142) );
  XNOR U35026 ( .A(n33138), .B(n33140), .Z(n36162) );
  XNOR U35027 ( .A(q[8]), .B(DB[428]), .Z(n33140) );
  XNOR U35028 ( .A(q[11]), .B(DB[431]), .Z(n33138) );
  IV U35029 ( .A(n33137), .Z(n36161) );
  XNOR U35030 ( .A(n33135), .B(n36163), .Z(n33137) );
  XNOR U35031 ( .A(q[10]), .B(DB[430]), .Z(n36163) );
  XNOR U35032 ( .A(q[9]), .B(DB[429]), .Z(n33135) );
  IV U35033 ( .A(n33150), .Z(n36157) );
  XOR U35034 ( .A(n36164), .B(n36165), .Z(n33150) );
  XNOR U35035 ( .A(n33167), .B(n33148), .Z(n36165) );
  XNOR U35036 ( .A(q[0]), .B(DB[420]), .Z(n33148) );
  XOR U35037 ( .A(n36166), .B(n33156), .Z(n33167) );
  XNOR U35038 ( .A(q[7]), .B(DB[427]), .Z(n33156) );
  IV U35039 ( .A(n33155), .Z(n36166) );
  XNOR U35040 ( .A(n33153), .B(n36167), .Z(n33155) );
  XNOR U35041 ( .A(q[6]), .B(DB[426]), .Z(n36167) );
  XNOR U35042 ( .A(q[5]), .B(DB[425]), .Z(n33153) );
  IV U35043 ( .A(n33166), .Z(n36164) );
  XOR U35044 ( .A(n36168), .B(n36169), .Z(n33166) );
  XNOR U35045 ( .A(n33162), .B(n33164), .Z(n36169) );
  XNOR U35046 ( .A(q[1]), .B(DB[421]), .Z(n33164) );
  XNOR U35047 ( .A(q[4]), .B(DB[424]), .Z(n33162) );
  IV U35048 ( .A(n33161), .Z(n36168) );
  XNOR U35049 ( .A(n33159), .B(n36170), .Z(n33161) );
  XNOR U35050 ( .A(q[3]), .B(DB[423]), .Z(n36170) );
  XNOR U35051 ( .A(q[2]), .B(DB[422]), .Z(n33159) );
  XOR U35052 ( .A(n36171), .B(n33057), .Z(n32985) );
  XOR U35053 ( .A(n36172), .B(n33049), .Z(n33057) );
  XOR U35054 ( .A(n36173), .B(n33038), .Z(n33049) );
  XNOR U35055 ( .A(q[14]), .B(DB[449]), .Z(n33038) );
  IV U35056 ( .A(n33037), .Z(n36173) );
  XNOR U35057 ( .A(n33035), .B(n36174), .Z(n33037) );
  XNOR U35058 ( .A(q[13]), .B(DB[448]), .Z(n36174) );
  XNOR U35059 ( .A(q[12]), .B(DB[447]), .Z(n33035) );
  IV U35060 ( .A(n33048), .Z(n36172) );
  XOR U35061 ( .A(n36175), .B(n36176), .Z(n33048) );
  XNOR U35062 ( .A(n33044), .B(n33046), .Z(n36176) );
  XNOR U35063 ( .A(q[8]), .B(DB[443]), .Z(n33046) );
  XNOR U35064 ( .A(q[11]), .B(DB[446]), .Z(n33044) );
  IV U35065 ( .A(n33043), .Z(n36175) );
  XNOR U35066 ( .A(n33041), .B(n36177), .Z(n33043) );
  XNOR U35067 ( .A(q[10]), .B(DB[445]), .Z(n36177) );
  XNOR U35068 ( .A(q[9]), .B(DB[444]), .Z(n33041) );
  IV U35069 ( .A(n33056), .Z(n36171) );
  XOR U35070 ( .A(n36178), .B(n36179), .Z(n33056) );
  XNOR U35071 ( .A(n33073), .B(n33054), .Z(n36179) );
  XNOR U35072 ( .A(q[0]), .B(DB[435]), .Z(n33054) );
  XOR U35073 ( .A(n36180), .B(n33062), .Z(n33073) );
  XNOR U35074 ( .A(q[7]), .B(DB[442]), .Z(n33062) );
  IV U35075 ( .A(n33061), .Z(n36180) );
  XNOR U35076 ( .A(n33059), .B(n36181), .Z(n33061) );
  XNOR U35077 ( .A(q[6]), .B(DB[441]), .Z(n36181) );
  XNOR U35078 ( .A(q[5]), .B(DB[440]), .Z(n33059) );
  IV U35079 ( .A(n33072), .Z(n36178) );
  XOR U35080 ( .A(n36182), .B(n36183), .Z(n33072) );
  XNOR U35081 ( .A(n33068), .B(n33070), .Z(n36183) );
  XNOR U35082 ( .A(q[1]), .B(DB[436]), .Z(n33070) );
  XNOR U35083 ( .A(q[4]), .B(DB[439]), .Z(n33068) );
  IV U35084 ( .A(n33067), .Z(n36182) );
  XNOR U35085 ( .A(n33065), .B(n36184), .Z(n33067) );
  XNOR U35086 ( .A(q[3]), .B(DB[438]), .Z(n36184) );
  XNOR U35087 ( .A(q[2]), .B(DB[437]), .Z(n33065) );
  XOR U35088 ( .A(n36185), .B(n32963), .Z(n32891) );
  XOR U35089 ( .A(n36186), .B(n32955), .Z(n32963) );
  XOR U35090 ( .A(n36187), .B(n32944), .Z(n32955) );
  XNOR U35091 ( .A(q[14]), .B(DB[464]), .Z(n32944) );
  IV U35092 ( .A(n32943), .Z(n36187) );
  XNOR U35093 ( .A(n32941), .B(n36188), .Z(n32943) );
  XNOR U35094 ( .A(q[13]), .B(DB[463]), .Z(n36188) );
  XNOR U35095 ( .A(q[12]), .B(DB[462]), .Z(n32941) );
  IV U35096 ( .A(n32954), .Z(n36186) );
  XOR U35097 ( .A(n36189), .B(n36190), .Z(n32954) );
  XNOR U35098 ( .A(n32950), .B(n32952), .Z(n36190) );
  XNOR U35099 ( .A(q[8]), .B(DB[458]), .Z(n32952) );
  XNOR U35100 ( .A(q[11]), .B(DB[461]), .Z(n32950) );
  IV U35101 ( .A(n32949), .Z(n36189) );
  XNOR U35102 ( .A(n32947), .B(n36191), .Z(n32949) );
  XNOR U35103 ( .A(q[10]), .B(DB[460]), .Z(n36191) );
  XNOR U35104 ( .A(q[9]), .B(DB[459]), .Z(n32947) );
  IV U35105 ( .A(n32962), .Z(n36185) );
  XOR U35106 ( .A(n36192), .B(n36193), .Z(n32962) );
  XNOR U35107 ( .A(n32979), .B(n32960), .Z(n36193) );
  XNOR U35108 ( .A(q[0]), .B(DB[450]), .Z(n32960) );
  XOR U35109 ( .A(n36194), .B(n32968), .Z(n32979) );
  XNOR U35110 ( .A(q[7]), .B(DB[457]), .Z(n32968) );
  IV U35111 ( .A(n32967), .Z(n36194) );
  XNOR U35112 ( .A(n32965), .B(n36195), .Z(n32967) );
  XNOR U35113 ( .A(q[6]), .B(DB[456]), .Z(n36195) );
  XNOR U35114 ( .A(q[5]), .B(DB[455]), .Z(n32965) );
  IV U35115 ( .A(n32978), .Z(n36192) );
  XOR U35116 ( .A(n36196), .B(n36197), .Z(n32978) );
  XNOR U35117 ( .A(n32974), .B(n32976), .Z(n36197) );
  XNOR U35118 ( .A(q[1]), .B(DB[451]), .Z(n32976) );
  XNOR U35119 ( .A(q[4]), .B(DB[454]), .Z(n32974) );
  IV U35120 ( .A(n32973), .Z(n36196) );
  XNOR U35121 ( .A(n32971), .B(n36198), .Z(n32973) );
  XNOR U35122 ( .A(q[3]), .B(DB[453]), .Z(n36198) );
  XNOR U35123 ( .A(q[2]), .B(DB[452]), .Z(n32971) );
  XOR U35124 ( .A(n36199), .B(n32869), .Z(n32797) );
  XOR U35125 ( .A(n36200), .B(n32861), .Z(n32869) );
  XOR U35126 ( .A(n36201), .B(n32850), .Z(n32861) );
  XNOR U35127 ( .A(q[14]), .B(DB[479]), .Z(n32850) );
  IV U35128 ( .A(n32849), .Z(n36201) );
  XNOR U35129 ( .A(n32847), .B(n36202), .Z(n32849) );
  XNOR U35130 ( .A(q[13]), .B(DB[478]), .Z(n36202) );
  XNOR U35131 ( .A(q[12]), .B(DB[477]), .Z(n32847) );
  IV U35132 ( .A(n32860), .Z(n36200) );
  XOR U35133 ( .A(n36203), .B(n36204), .Z(n32860) );
  XNOR U35134 ( .A(n32856), .B(n32858), .Z(n36204) );
  XNOR U35135 ( .A(q[8]), .B(DB[473]), .Z(n32858) );
  XNOR U35136 ( .A(q[11]), .B(DB[476]), .Z(n32856) );
  IV U35137 ( .A(n32855), .Z(n36203) );
  XNOR U35138 ( .A(n32853), .B(n36205), .Z(n32855) );
  XNOR U35139 ( .A(q[10]), .B(DB[475]), .Z(n36205) );
  XNOR U35140 ( .A(q[9]), .B(DB[474]), .Z(n32853) );
  IV U35141 ( .A(n32868), .Z(n36199) );
  XOR U35142 ( .A(n36206), .B(n36207), .Z(n32868) );
  XNOR U35143 ( .A(n32885), .B(n32866), .Z(n36207) );
  XNOR U35144 ( .A(q[0]), .B(DB[465]), .Z(n32866) );
  XOR U35145 ( .A(n36208), .B(n32874), .Z(n32885) );
  XNOR U35146 ( .A(q[7]), .B(DB[472]), .Z(n32874) );
  IV U35147 ( .A(n32873), .Z(n36208) );
  XNOR U35148 ( .A(n32871), .B(n36209), .Z(n32873) );
  XNOR U35149 ( .A(q[6]), .B(DB[471]), .Z(n36209) );
  XNOR U35150 ( .A(q[5]), .B(DB[470]), .Z(n32871) );
  IV U35151 ( .A(n32884), .Z(n36206) );
  XOR U35152 ( .A(n36210), .B(n36211), .Z(n32884) );
  XNOR U35153 ( .A(n32880), .B(n32882), .Z(n36211) );
  XNOR U35154 ( .A(q[1]), .B(DB[466]), .Z(n32882) );
  XNOR U35155 ( .A(q[4]), .B(DB[469]), .Z(n32880) );
  IV U35156 ( .A(n32879), .Z(n36210) );
  XNOR U35157 ( .A(n32877), .B(n36212), .Z(n32879) );
  XNOR U35158 ( .A(q[3]), .B(DB[468]), .Z(n36212) );
  XNOR U35159 ( .A(q[2]), .B(DB[467]), .Z(n32877) );
  XOR U35160 ( .A(n36213), .B(n32775), .Z(n32703) );
  XOR U35161 ( .A(n36214), .B(n32767), .Z(n32775) );
  XOR U35162 ( .A(n36215), .B(n32756), .Z(n32767) );
  XNOR U35163 ( .A(q[14]), .B(DB[494]), .Z(n32756) );
  IV U35164 ( .A(n32755), .Z(n36215) );
  XNOR U35165 ( .A(n32753), .B(n36216), .Z(n32755) );
  XNOR U35166 ( .A(q[13]), .B(DB[493]), .Z(n36216) );
  XNOR U35167 ( .A(q[12]), .B(DB[492]), .Z(n32753) );
  IV U35168 ( .A(n32766), .Z(n36214) );
  XOR U35169 ( .A(n36217), .B(n36218), .Z(n32766) );
  XNOR U35170 ( .A(n32762), .B(n32764), .Z(n36218) );
  XNOR U35171 ( .A(q[8]), .B(DB[488]), .Z(n32764) );
  XNOR U35172 ( .A(q[11]), .B(DB[491]), .Z(n32762) );
  IV U35173 ( .A(n32761), .Z(n36217) );
  XNOR U35174 ( .A(n32759), .B(n36219), .Z(n32761) );
  XNOR U35175 ( .A(q[10]), .B(DB[490]), .Z(n36219) );
  XNOR U35176 ( .A(q[9]), .B(DB[489]), .Z(n32759) );
  IV U35177 ( .A(n32774), .Z(n36213) );
  XOR U35178 ( .A(n36220), .B(n36221), .Z(n32774) );
  XNOR U35179 ( .A(n32791), .B(n32772), .Z(n36221) );
  XNOR U35180 ( .A(q[0]), .B(DB[480]), .Z(n32772) );
  XOR U35181 ( .A(n36222), .B(n32780), .Z(n32791) );
  XNOR U35182 ( .A(q[7]), .B(DB[487]), .Z(n32780) );
  IV U35183 ( .A(n32779), .Z(n36222) );
  XNOR U35184 ( .A(n32777), .B(n36223), .Z(n32779) );
  XNOR U35185 ( .A(q[6]), .B(DB[486]), .Z(n36223) );
  XNOR U35186 ( .A(q[5]), .B(DB[485]), .Z(n32777) );
  IV U35187 ( .A(n32790), .Z(n36220) );
  XOR U35188 ( .A(n36224), .B(n36225), .Z(n32790) );
  XNOR U35189 ( .A(n32786), .B(n32788), .Z(n36225) );
  XNOR U35190 ( .A(q[1]), .B(DB[481]), .Z(n32788) );
  XNOR U35191 ( .A(q[4]), .B(DB[484]), .Z(n32786) );
  IV U35192 ( .A(n32785), .Z(n36224) );
  XNOR U35193 ( .A(n32783), .B(n36226), .Z(n32785) );
  XNOR U35194 ( .A(q[3]), .B(DB[483]), .Z(n36226) );
  XNOR U35195 ( .A(q[2]), .B(DB[482]), .Z(n32783) );
  XOR U35196 ( .A(n36227), .B(n32681), .Z(n32609) );
  XOR U35197 ( .A(n36228), .B(n32673), .Z(n32681) );
  XOR U35198 ( .A(n36229), .B(n32662), .Z(n32673) );
  XNOR U35199 ( .A(q[14]), .B(DB[509]), .Z(n32662) );
  IV U35200 ( .A(n32661), .Z(n36229) );
  XNOR U35201 ( .A(n32659), .B(n36230), .Z(n32661) );
  XNOR U35202 ( .A(q[13]), .B(DB[508]), .Z(n36230) );
  XNOR U35203 ( .A(q[12]), .B(DB[507]), .Z(n32659) );
  IV U35204 ( .A(n32672), .Z(n36228) );
  XOR U35205 ( .A(n36231), .B(n36232), .Z(n32672) );
  XNOR U35206 ( .A(n32668), .B(n32670), .Z(n36232) );
  XNOR U35207 ( .A(q[8]), .B(DB[503]), .Z(n32670) );
  XNOR U35208 ( .A(q[11]), .B(DB[506]), .Z(n32668) );
  IV U35209 ( .A(n32667), .Z(n36231) );
  XNOR U35210 ( .A(n32665), .B(n36233), .Z(n32667) );
  XNOR U35211 ( .A(q[10]), .B(DB[505]), .Z(n36233) );
  XNOR U35212 ( .A(q[9]), .B(DB[504]), .Z(n32665) );
  IV U35213 ( .A(n32680), .Z(n36227) );
  XOR U35214 ( .A(n36234), .B(n36235), .Z(n32680) );
  XNOR U35215 ( .A(n32697), .B(n32678), .Z(n36235) );
  XNOR U35216 ( .A(q[0]), .B(DB[495]), .Z(n32678) );
  XOR U35217 ( .A(n36236), .B(n32686), .Z(n32697) );
  XNOR U35218 ( .A(q[7]), .B(DB[502]), .Z(n32686) );
  IV U35219 ( .A(n32685), .Z(n36236) );
  XNOR U35220 ( .A(n32683), .B(n36237), .Z(n32685) );
  XNOR U35221 ( .A(q[6]), .B(DB[501]), .Z(n36237) );
  XNOR U35222 ( .A(q[5]), .B(DB[500]), .Z(n32683) );
  IV U35223 ( .A(n32696), .Z(n36234) );
  XOR U35224 ( .A(n36238), .B(n36239), .Z(n32696) );
  XNOR U35225 ( .A(n32692), .B(n32694), .Z(n36239) );
  XNOR U35226 ( .A(q[1]), .B(DB[496]), .Z(n32694) );
  XNOR U35227 ( .A(q[4]), .B(DB[499]), .Z(n32692) );
  IV U35228 ( .A(n32691), .Z(n36238) );
  XNOR U35229 ( .A(n32689), .B(n36240), .Z(n32691) );
  XNOR U35230 ( .A(q[3]), .B(DB[498]), .Z(n36240) );
  XNOR U35231 ( .A(q[2]), .B(DB[497]), .Z(n32689) );
  XOR U35232 ( .A(n36241), .B(n32587), .Z(n32515) );
  XOR U35233 ( .A(n36242), .B(n32579), .Z(n32587) );
  XOR U35234 ( .A(n36243), .B(n32568), .Z(n32579) );
  XNOR U35235 ( .A(q[14]), .B(DB[524]), .Z(n32568) );
  IV U35236 ( .A(n32567), .Z(n36243) );
  XNOR U35237 ( .A(n32565), .B(n36244), .Z(n32567) );
  XNOR U35238 ( .A(q[13]), .B(DB[523]), .Z(n36244) );
  XNOR U35239 ( .A(q[12]), .B(DB[522]), .Z(n32565) );
  IV U35240 ( .A(n32578), .Z(n36242) );
  XOR U35241 ( .A(n36245), .B(n36246), .Z(n32578) );
  XNOR U35242 ( .A(n32574), .B(n32576), .Z(n36246) );
  XNOR U35243 ( .A(q[8]), .B(DB[518]), .Z(n32576) );
  XNOR U35244 ( .A(q[11]), .B(DB[521]), .Z(n32574) );
  IV U35245 ( .A(n32573), .Z(n36245) );
  XNOR U35246 ( .A(n32571), .B(n36247), .Z(n32573) );
  XNOR U35247 ( .A(q[10]), .B(DB[520]), .Z(n36247) );
  XNOR U35248 ( .A(q[9]), .B(DB[519]), .Z(n32571) );
  IV U35249 ( .A(n32586), .Z(n36241) );
  XOR U35250 ( .A(n36248), .B(n36249), .Z(n32586) );
  XNOR U35251 ( .A(n32603), .B(n32584), .Z(n36249) );
  XNOR U35252 ( .A(q[0]), .B(DB[510]), .Z(n32584) );
  XOR U35253 ( .A(n36250), .B(n32592), .Z(n32603) );
  XNOR U35254 ( .A(q[7]), .B(DB[517]), .Z(n32592) );
  IV U35255 ( .A(n32591), .Z(n36250) );
  XNOR U35256 ( .A(n32589), .B(n36251), .Z(n32591) );
  XNOR U35257 ( .A(q[6]), .B(DB[516]), .Z(n36251) );
  XNOR U35258 ( .A(q[5]), .B(DB[515]), .Z(n32589) );
  IV U35259 ( .A(n32602), .Z(n36248) );
  XOR U35260 ( .A(n36252), .B(n36253), .Z(n32602) );
  XNOR U35261 ( .A(n32598), .B(n32600), .Z(n36253) );
  XNOR U35262 ( .A(q[1]), .B(DB[511]), .Z(n32600) );
  XNOR U35263 ( .A(q[4]), .B(DB[514]), .Z(n32598) );
  IV U35264 ( .A(n32597), .Z(n36252) );
  XNOR U35265 ( .A(n32595), .B(n36254), .Z(n32597) );
  XNOR U35266 ( .A(q[3]), .B(DB[513]), .Z(n36254) );
  XNOR U35267 ( .A(q[2]), .B(DB[512]), .Z(n32595) );
  XOR U35268 ( .A(n36255), .B(n32493), .Z(n32421) );
  XOR U35269 ( .A(n36256), .B(n32485), .Z(n32493) );
  XOR U35270 ( .A(n36257), .B(n32474), .Z(n32485) );
  XNOR U35271 ( .A(q[14]), .B(DB[539]), .Z(n32474) );
  IV U35272 ( .A(n32473), .Z(n36257) );
  XNOR U35273 ( .A(n32471), .B(n36258), .Z(n32473) );
  XNOR U35274 ( .A(q[13]), .B(DB[538]), .Z(n36258) );
  XNOR U35275 ( .A(q[12]), .B(DB[537]), .Z(n32471) );
  IV U35276 ( .A(n32484), .Z(n36256) );
  XOR U35277 ( .A(n36259), .B(n36260), .Z(n32484) );
  XNOR U35278 ( .A(n32480), .B(n32482), .Z(n36260) );
  XNOR U35279 ( .A(q[8]), .B(DB[533]), .Z(n32482) );
  XNOR U35280 ( .A(q[11]), .B(DB[536]), .Z(n32480) );
  IV U35281 ( .A(n32479), .Z(n36259) );
  XNOR U35282 ( .A(n32477), .B(n36261), .Z(n32479) );
  XNOR U35283 ( .A(q[10]), .B(DB[535]), .Z(n36261) );
  XNOR U35284 ( .A(q[9]), .B(DB[534]), .Z(n32477) );
  IV U35285 ( .A(n32492), .Z(n36255) );
  XOR U35286 ( .A(n36262), .B(n36263), .Z(n32492) );
  XNOR U35287 ( .A(n32509), .B(n32490), .Z(n36263) );
  XNOR U35288 ( .A(q[0]), .B(DB[525]), .Z(n32490) );
  XOR U35289 ( .A(n36264), .B(n32498), .Z(n32509) );
  XNOR U35290 ( .A(q[7]), .B(DB[532]), .Z(n32498) );
  IV U35291 ( .A(n32497), .Z(n36264) );
  XNOR U35292 ( .A(n32495), .B(n36265), .Z(n32497) );
  XNOR U35293 ( .A(q[6]), .B(DB[531]), .Z(n36265) );
  XNOR U35294 ( .A(q[5]), .B(DB[530]), .Z(n32495) );
  IV U35295 ( .A(n32508), .Z(n36262) );
  XOR U35296 ( .A(n36266), .B(n36267), .Z(n32508) );
  XNOR U35297 ( .A(n32504), .B(n32506), .Z(n36267) );
  XNOR U35298 ( .A(q[1]), .B(DB[526]), .Z(n32506) );
  XNOR U35299 ( .A(q[4]), .B(DB[529]), .Z(n32504) );
  IV U35300 ( .A(n32503), .Z(n36266) );
  XNOR U35301 ( .A(n32501), .B(n36268), .Z(n32503) );
  XNOR U35302 ( .A(q[3]), .B(DB[528]), .Z(n36268) );
  XNOR U35303 ( .A(q[2]), .B(DB[527]), .Z(n32501) );
  XOR U35304 ( .A(n36269), .B(n32399), .Z(n32327) );
  XOR U35305 ( .A(n36270), .B(n32391), .Z(n32399) );
  XOR U35306 ( .A(n36271), .B(n32380), .Z(n32391) );
  XNOR U35307 ( .A(q[14]), .B(DB[554]), .Z(n32380) );
  IV U35308 ( .A(n32379), .Z(n36271) );
  XNOR U35309 ( .A(n32377), .B(n36272), .Z(n32379) );
  XNOR U35310 ( .A(q[13]), .B(DB[553]), .Z(n36272) );
  XNOR U35311 ( .A(q[12]), .B(DB[552]), .Z(n32377) );
  IV U35312 ( .A(n32390), .Z(n36270) );
  XOR U35313 ( .A(n36273), .B(n36274), .Z(n32390) );
  XNOR U35314 ( .A(n32386), .B(n32388), .Z(n36274) );
  XNOR U35315 ( .A(q[8]), .B(DB[548]), .Z(n32388) );
  XNOR U35316 ( .A(q[11]), .B(DB[551]), .Z(n32386) );
  IV U35317 ( .A(n32385), .Z(n36273) );
  XNOR U35318 ( .A(n32383), .B(n36275), .Z(n32385) );
  XNOR U35319 ( .A(q[10]), .B(DB[550]), .Z(n36275) );
  XNOR U35320 ( .A(q[9]), .B(DB[549]), .Z(n32383) );
  IV U35321 ( .A(n32398), .Z(n36269) );
  XOR U35322 ( .A(n36276), .B(n36277), .Z(n32398) );
  XNOR U35323 ( .A(n32415), .B(n32396), .Z(n36277) );
  XNOR U35324 ( .A(q[0]), .B(DB[540]), .Z(n32396) );
  XOR U35325 ( .A(n36278), .B(n32404), .Z(n32415) );
  XNOR U35326 ( .A(q[7]), .B(DB[547]), .Z(n32404) );
  IV U35327 ( .A(n32403), .Z(n36278) );
  XNOR U35328 ( .A(n32401), .B(n36279), .Z(n32403) );
  XNOR U35329 ( .A(q[6]), .B(DB[546]), .Z(n36279) );
  XNOR U35330 ( .A(q[5]), .B(DB[545]), .Z(n32401) );
  IV U35331 ( .A(n32414), .Z(n36276) );
  XOR U35332 ( .A(n36280), .B(n36281), .Z(n32414) );
  XNOR U35333 ( .A(n32410), .B(n32412), .Z(n36281) );
  XNOR U35334 ( .A(q[1]), .B(DB[541]), .Z(n32412) );
  XNOR U35335 ( .A(q[4]), .B(DB[544]), .Z(n32410) );
  IV U35336 ( .A(n32409), .Z(n36280) );
  XNOR U35337 ( .A(n32407), .B(n36282), .Z(n32409) );
  XNOR U35338 ( .A(q[3]), .B(DB[543]), .Z(n36282) );
  XNOR U35339 ( .A(q[2]), .B(DB[542]), .Z(n32407) );
  XOR U35340 ( .A(n36283), .B(n32305), .Z(n32233) );
  XOR U35341 ( .A(n36284), .B(n32297), .Z(n32305) );
  XOR U35342 ( .A(n36285), .B(n32286), .Z(n32297) );
  XNOR U35343 ( .A(q[14]), .B(DB[569]), .Z(n32286) );
  IV U35344 ( .A(n32285), .Z(n36285) );
  XNOR U35345 ( .A(n32283), .B(n36286), .Z(n32285) );
  XNOR U35346 ( .A(q[13]), .B(DB[568]), .Z(n36286) );
  XNOR U35347 ( .A(q[12]), .B(DB[567]), .Z(n32283) );
  IV U35348 ( .A(n32296), .Z(n36284) );
  XOR U35349 ( .A(n36287), .B(n36288), .Z(n32296) );
  XNOR U35350 ( .A(n32292), .B(n32294), .Z(n36288) );
  XNOR U35351 ( .A(q[8]), .B(DB[563]), .Z(n32294) );
  XNOR U35352 ( .A(q[11]), .B(DB[566]), .Z(n32292) );
  IV U35353 ( .A(n32291), .Z(n36287) );
  XNOR U35354 ( .A(n32289), .B(n36289), .Z(n32291) );
  XNOR U35355 ( .A(q[10]), .B(DB[565]), .Z(n36289) );
  XNOR U35356 ( .A(q[9]), .B(DB[564]), .Z(n32289) );
  IV U35357 ( .A(n32304), .Z(n36283) );
  XOR U35358 ( .A(n36290), .B(n36291), .Z(n32304) );
  XNOR U35359 ( .A(n32321), .B(n32302), .Z(n36291) );
  XNOR U35360 ( .A(q[0]), .B(DB[555]), .Z(n32302) );
  XOR U35361 ( .A(n36292), .B(n32310), .Z(n32321) );
  XNOR U35362 ( .A(q[7]), .B(DB[562]), .Z(n32310) );
  IV U35363 ( .A(n32309), .Z(n36292) );
  XNOR U35364 ( .A(n32307), .B(n36293), .Z(n32309) );
  XNOR U35365 ( .A(q[6]), .B(DB[561]), .Z(n36293) );
  XNOR U35366 ( .A(q[5]), .B(DB[560]), .Z(n32307) );
  IV U35367 ( .A(n32320), .Z(n36290) );
  XOR U35368 ( .A(n36294), .B(n36295), .Z(n32320) );
  XNOR U35369 ( .A(n32316), .B(n32318), .Z(n36295) );
  XNOR U35370 ( .A(q[1]), .B(DB[556]), .Z(n32318) );
  XNOR U35371 ( .A(q[4]), .B(DB[559]), .Z(n32316) );
  IV U35372 ( .A(n32315), .Z(n36294) );
  XNOR U35373 ( .A(n32313), .B(n36296), .Z(n32315) );
  XNOR U35374 ( .A(q[3]), .B(DB[558]), .Z(n36296) );
  XNOR U35375 ( .A(q[2]), .B(DB[557]), .Z(n32313) );
  XOR U35376 ( .A(n36297), .B(n32211), .Z(n32139) );
  XOR U35377 ( .A(n36298), .B(n32203), .Z(n32211) );
  XOR U35378 ( .A(n36299), .B(n32192), .Z(n32203) );
  XNOR U35379 ( .A(q[14]), .B(DB[584]), .Z(n32192) );
  IV U35380 ( .A(n32191), .Z(n36299) );
  XNOR U35381 ( .A(n32189), .B(n36300), .Z(n32191) );
  XNOR U35382 ( .A(q[13]), .B(DB[583]), .Z(n36300) );
  XNOR U35383 ( .A(q[12]), .B(DB[582]), .Z(n32189) );
  IV U35384 ( .A(n32202), .Z(n36298) );
  XOR U35385 ( .A(n36301), .B(n36302), .Z(n32202) );
  XNOR U35386 ( .A(n32198), .B(n32200), .Z(n36302) );
  XNOR U35387 ( .A(q[8]), .B(DB[578]), .Z(n32200) );
  XNOR U35388 ( .A(q[11]), .B(DB[581]), .Z(n32198) );
  IV U35389 ( .A(n32197), .Z(n36301) );
  XNOR U35390 ( .A(n32195), .B(n36303), .Z(n32197) );
  XNOR U35391 ( .A(q[10]), .B(DB[580]), .Z(n36303) );
  XNOR U35392 ( .A(q[9]), .B(DB[579]), .Z(n32195) );
  IV U35393 ( .A(n32210), .Z(n36297) );
  XOR U35394 ( .A(n36304), .B(n36305), .Z(n32210) );
  XNOR U35395 ( .A(n32227), .B(n32208), .Z(n36305) );
  XNOR U35396 ( .A(q[0]), .B(DB[570]), .Z(n32208) );
  XOR U35397 ( .A(n36306), .B(n32216), .Z(n32227) );
  XNOR U35398 ( .A(q[7]), .B(DB[577]), .Z(n32216) );
  IV U35399 ( .A(n32215), .Z(n36306) );
  XNOR U35400 ( .A(n32213), .B(n36307), .Z(n32215) );
  XNOR U35401 ( .A(q[6]), .B(DB[576]), .Z(n36307) );
  XNOR U35402 ( .A(q[5]), .B(DB[575]), .Z(n32213) );
  IV U35403 ( .A(n32226), .Z(n36304) );
  XOR U35404 ( .A(n36308), .B(n36309), .Z(n32226) );
  XNOR U35405 ( .A(n32222), .B(n32224), .Z(n36309) );
  XNOR U35406 ( .A(q[1]), .B(DB[571]), .Z(n32224) );
  XNOR U35407 ( .A(q[4]), .B(DB[574]), .Z(n32222) );
  IV U35408 ( .A(n32221), .Z(n36308) );
  XNOR U35409 ( .A(n32219), .B(n36310), .Z(n32221) );
  XNOR U35410 ( .A(q[3]), .B(DB[573]), .Z(n36310) );
  XNOR U35411 ( .A(q[2]), .B(DB[572]), .Z(n32219) );
  XOR U35412 ( .A(n36311), .B(n32117), .Z(n32045) );
  XOR U35413 ( .A(n36312), .B(n32109), .Z(n32117) );
  XOR U35414 ( .A(n36313), .B(n32098), .Z(n32109) );
  XNOR U35415 ( .A(q[14]), .B(DB[599]), .Z(n32098) );
  IV U35416 ( .A(n32097), .Z(n36313) );
  XNOR U35417 ( .A(n32095), .B(n36314), .Z(n32097) );
  XNOR U35418 ( .A(q[13]), .B(DB[598]), .Z(n36314) );
  XNOR U35419 ( .A(q[12]), .B(DB[597]), .Z(n32095) );
  IV U35420 ( .A(n32108), .Z(n36312) );
  XOR U35421 ( .A(n36315), .B(n36316), .Z(n32108) );
  XNOR U35422 ( .A(n32104), .B(n32106), .Z(n36316) );
  XNOR U35423 ( .A(q[8]), .B(DB[593]), .Z(n32106) );
  XNOR U35424 ( .A(q[11]), .B(DB[596]), .Z(n32104) );
  IV U35425 ( .A(n32103), .Z(n36315) );
  XNOR U35426 ( .A(n32101), .B(n36317), .Z(n32103) );
  XNOR U35427 ( .A(q[10]), .B(DB[595]), .Z(n36317) );
  XNOR U35428 ( .A(q[9]), .B(DB[594]), .Z(n32101) );
  IV U35429 ( .A(n32116), .Z(n36311) );
  XOR U35430 ( .A(n36318), .B(n36319), .Z(n32116) );
  XNOR U35431 ( .A(n32133), .B(n32114), .Z(n36319) );
  XNOR U35432 ( .A(q[0]), .B(DB[585]), .Z(n32114) );
  XOR U35433 ( .A(n36320), .B(n32122), .Z(n32133) );
  XNOR U35434 ( .A(q[7]), .B(DB[592]), .Z(n32122) );
  IV U35435 ( .A(n32121), .Z(n36320) );
  XNOR U35436 ( .A(n32119), .B(n36321), .Z(n32121) );
  XNOR U35437 ( .A(q[6]), .B(DB[591]), .Z(n36321) );
  XNOR U35438 ( .A(q[5]), .B(DB[590]), .Z(n32119) );
  IV U35439 ( .A(n32132), .Z(n36318) );
  XOR U35440 ( .A(n36322), .B(n36323), .Z(n32132) );
  XNOR U35441 ( .A(n32128), .B(n32130), .Z(n36323) );
  XNOR U35442 ( .A(q[1]), .B(DB[586]), .Z(n32130) );
  XNOR U35443 ( .A(q[4]), .B(DB[589]), .Z(n32128) );
  IV U35444 ( .A(n32127), .Z(n36322) );
  XNOR U35445 ( .A(n32125), .B(n36324), .Z(n32127) );
  XNOR U35446 ( .A(q[3]), .B(DB[588]), .Z(n36324) );
  XNOR U35447 ( .A(q[2]), .B(DB[587]), .Z(n32125) );
  XOR U35448 ( .A(n36325), .B(n32023), .Z(n31951) );
  XOR U35449 ( .A(n36326), .B(n32015), .Z(n32023) );
  XOR U35450 ( .A(n36327), .B(n32004), .Z(n32015) );
  XNOR U35451 ( .A(q[14]), .B(DB[614]), .Z(n32004) );
  IV U35452 ( .A(n32003), .Z(n36327) );
  XNOR U35453 ( .A(n32001), .B(n36328), .Z(n32003) );
  XNOR U35454 ( .A(q[13]), .B(DB[613]), .Z(n36328) );
  XNOR U35455 ( .A(q[12]), .B(DB[612]), .Z(n32001) );
  IV U35456 ( .A(n32014), .Z(n36326) );
  XOR U35457 ( .A(n36329), .B(n36330), .Z(n32014) );
  XNOR U35458 ( .A(n32010), .B(n32012), .Z(n36330) );
  XNOR U35459 ( .A(q[8]), .B(DB[608]), .Z(n32012) );
  XNOR U35460 ( .A(q[11]), .B(DB[611]), .Z(n32010) );
  IV U35461 ( .A(n32009), .Z(n36329) );
  XNOR U35462 ( .A(n32007), .B(n36331), .Z(n32009) );
  XNOR U35463 ( .A(q[10]), .B(DB[610]), .Z(n36331) );
  XNOR U35464 ( .A(q[9]), .B(DB[609]), .Z(n32007) );
  IV U35465 ( .A(n32022), .Z(n36325) );
  XOR U35466 ( .A(n36332), .B(n36333), .Z(n32022) );
  XNOR U35467 ( .A(n32039), .B(n32020), .Z(n36333) );
  XNOR U35468 ( .A(q[0]), .B(DB[600]), .Z(n32020) );
  XOR U35469 ( .A(n36334), .B(n32028), .Z(n32039) );
  XNOR U35470 ( .A(q[7]), .B(DB[607]), .Z(n32028) );
  IV U35471 ( .A(n32027), .Z(n36334) );
  XNOR U35472 ( .A(n32025), .B(n36335), .Z(n32027) );
  XNOR U35473 ( .A(q[6]), .B(DB[606]), .Z(n36335) );
  XNOR U35474 ( .A(q[5]), .B(DB[605]), .Z(n32025) );
  IV U35475 ( .A(n32038), .Z(n36332) );
  XOR U35476 ( .A(n36336), .B(n36337), .Z(n32038) );
  XNOR U35477 ( .A(n32034), .B(n32036), .Z(n36337) );
  XNOR U35478 ( .A(q[1]), .B(DB[601]), .Z(n32036) );
  XNOR U35479 ( .A(q[4]), .B(DB[604]), .Z(n32034) );
  IV U35480 ( .A(n32033), .Z(n36336) );
  XNOR U35481 ( .A(n32031), .B(n36338), .Z(n32033) );
  XNOR U35482 ( .A(q[3]), .B(DB[603]), .Z(n36338) );
  XNOR U35483 ( .A(q[2]), .B(DB[602]), .Z(n32031) );
  XOR U35484 ( .A(n36339), .B(n31929), .Z(n31857) );
  XOR U35485 ( .A(n36340), .B(n31921), .Z(n31929) );
  XOR U35486 ( .A(n36341), .B(n31910), .Z(n31921) );
  XNOR U35487 ( .A(q[14]), .B(DB[629]), .Z(n31910) );
  IV U35488 ( .A(n31909), .Z(n36341) );
  XNOR U35489 ( .A(n31907), .B(n36342), .Z(n31909) );
  XNOR U35490 ( .A(q[13]), .B(DB[628]), .Z(n36342) );
  XNOR U35491 ( .A(q[12]), .B(DB[627]), .Z(n31907) );
  IV U35492 ( .A(n31920), .Z(n36340) );
  XOR U35493 ( .A(n36343), .B(n36344), .Z(n31920) );
  XNOR U35494 ( .A(n31916), .B(n31918), .Z(n36344) );
  XNOR U35495 ( .A(q[8]), .B(DB[623]), .Z(n31918) );
  XNOR U35496 ( .A(q[11]), .B(DB[626]), .Z(n31916) );
  IV U35497 ( .A(n31915), .Z(n36343) );
  XNOR U35498 ( .A(n31913), .B(n36345), .Z(n31915) );
  XNOR U35499 ( .A(q[10]), .B(DB[625]), .Z(n36345) );
  XNOR U35500 ( .A(q[9]), .B(DB[624]), .Z(n31913) );
  IV U35501 ( .A(n31928), .Z(n36339) );
  XOR U35502 ( .A(n36346), .B(n36347), .Z(n31928) );
  XNOR U35503 ( .A(n31945), .B(n31926), .Z(n36347) );
  XNOR U35504 ( .A(q[0]), .B(DB[615]), .Z(n31926) );
  XOR U35505 ( .A(n36348), .B(n31934), .Z(n31945) );
  XNOR U35506 ( .A(q[7]), .B(DB[622]), .Z(n31934) );
  IV U35507 ( .A(n31933), .Z(n36348) );
  XNOR U35508 ( .A(n31931), .B(n36349), .Z(n31933) );
  XNOR U35509 ( .A(q[6]), .B(DB[621]), .Z(n36349) );
  XNOR U35510 ( .A(q[5]), .B(DB[620]), .Z(n31931) );
  IV U35511 ( .A(n31944), .Z(n36346) );
  XOR U35512 ( .A(n36350), .B(n36351), .Z(n31944) );
  XNOR U35513 ( .A(n31940), .B(n31942), .Z(n36351) );
  XNOR U35514 ( .A(q[1]), .B(DB[616]), .Z(n31942) );
  XNOR U35515 ( .A(q[4]), .B(DB[619]), .Z(n31940) );
  IV U35516 ( .A(n31939), .Z(n36350) );
  XNOR U35517 ( .A(n31937), .B(n36352), .Z(n31939) );
  XNOR U35518 ( .A(q[3]), .B(DB[618]), .Z(n36352) );
  XNOR U35519 ( .A(q[2]), .B(DB[617]), .Z(n31937) );
  XOR U35520 ( .A(n36353), .B(n31835), .Z(n31763) );
  XOR U35521 ( .A(n36354), .B(n31827), .Z(n31835) );
  XOR U35522 ( .A(n36355), .B(n31816), .Z(n31827) );
  XNOR U35523 ( .A(q[14]), .B(DB[644]), .Z(n31816) );
  IV U35524 ( .A(n31815), .Z(n36355) );
  XNOR U35525 ( .A(n31813), .B(n36356), .Z(n31815) );
  XNOR U35526 ( .A(q[13]), .B(DB[643]), .Z(n36356) );
  XNOR U35527 ( .A(q[12]), .B(DB[642]), .Z(n31813) );
  IV U35528 ( .A(n31826), .Z(n36354) );
  XOR U35529 ( .A(n36357), .B(n36358), .Z(n31826) );
  XNOR U35530 ( .A(n31822), .B(n31824), .Z(n36358) );
  XNOR U35531 ( .A(q[8]), .B(DB[638]), .Z(n31824) );
  XNOR U35532 ( .A(q[11]), .B(DB[641]), .Z(n31822) );
  IV U35533 ( .A(n31821), .Z(n36357) );
  XNOR U35534 ( .A(n31819), .B(n36359), .Z(n31821) );
  XNOR U35535 ( .A(q[10]), .B(DB[640]), .Z(n36359) );
  XNOR U35536 ( .A(q[9]), .B(DB[639]), .Z(n31819) );
  IV U35537 ( .A(n31834), .Z(n36353) );
  XOR U35538 ( .A(n36360), .B(n36361), .Z(n31834) );
  XNOR U35539 ( .A(n31851), .B(n31832), .Z(n36361) );
  XNOR U35540 ( .A(q[0]), .B(DB[630]), .Z(n31832) );
  XOR U35541 ( .A(n36362), .B(n31840), .Z(n31851) );
  XNOR U35542 ( .A(q[7]), .B(DB[637]), .Z(n31840) );
  IV U35543 ( .A(n31839), .Z(n36362) );
  XNOR U35544 ( .A(n31837), .B(n36363), .Z(n31839) );
  XNOR U35545 ( .A(q[6]), .B(DB[636]), .Z(n36363) );
  XNOR U35546 ( .A(q[5]), .B(DB[635]), .Z(n31837) );
  IV U35547 ( .A(n31850), .Z(n36360) );
  XOR U35548 ( .A(n36364), .B(n36365), .Z(n31850) );
  XNOR U35549 ( .A(n31846), .B(n31848), .Z(n36365) );
  XNOR U35550 ( .A(q[1]), .B(DB[631]), .Z(n31848) );
  XNOR U35551 ( .A(q[4]), .B(DB[634]), .Z(n31846) );
  IV U35552 ( .A(n31845), .Z(n36364) );
  XNOR U35553 ( .A(n31843), .B(n36366), .Z(n31845) );
  XNOR U35554 ( .A(q[3]), .B(DB[633]), .Z(n36366) );
  XNOR U35555 ( .A(q[2]), .B(DB[632]), .Z(n31843) );
  XOR U35556 ( .A(n36367), .B(n31741), .Z(n31669) );
  XOR U35557 ( .A(n36368), .B(n31733), .Z(n31741) );
  XOR U35558 ( .A(n36369), .B(n31722), .Z(n31733) );
  XNOR U35559 ( .A(q[14]), .B(DB[659]), .Z(n31722) );
  IV U35560 ( .A(n31721), .Z(n36369) );
  XNOR U35561 ( .A(n31719), .B(n36370), .Z(n31721) );
  XNOR U35562 ( .A(q[13]), .B(DB[658]), .Z(n36370) );
  XNOR U35563 ( .A(q[12]), .B(DB[657]), .Z(n31719) );
  IV U35564 ( .A(n31732), .Z(n36368) );
  XOR U35565 ( .A(n36371), .B(n36372), .Z(n31732) );
  XNOR U35566 ( .A(n31728), .B(n31730), .Z(n36372) );
  XNOR U35567 ( .A(q[8]), .B(DB[653]), .Z(n31730) );
  XNOR U35568 ( .A(q[11]), .B(DB[656]), .Z(n31728) );
  IV U35569 ( .A(n31727), .Z(n36371) );
  XNOR U35570 ( .A(n31725), .B(n36373), .Z(n31727) );
  XNOR U35571 ( .A(q[10]), .B(DB[655]), .Z(n36373) );
  XNOR U35572 ( .A(q[9]), .B(DB[654]), .Z(n31725) );
  IV U35573 ( .A(n31740), .Z(n36367) );
  XOR U35574 ( .A(n36374), .B(n36375), .Z(n31740) );
  XNOR U35575 ( .A(n31757), .B(n31738), .Z(n36375) );
  XNOR U35576 ( .A(q[0]), .B(DB[645]), .Z(n31738) );
  XOR U35577 ( .A(n36376), .B(n31746), .Z(n31757) );
  XNOR U35578 ( .A(q[7]), .B(DB[652]), .Z(n31746) );
  IV U35579 ( .A(n31745), .Z(n36376) );
  XNOR U35580 ( .A(n31743), .B(n36377), .Z(n31745) );
  XNOR U35581 ( .A(q[6]), .B(DB[651]), .Z(n36377) );
  XNOR U35582 ( .A(q[5]), .B(DB[650]), .Z(n31743) );
  IV U35583 ( .A(n31756), .Z(n36374) );
  XOR U35584 ( .A(n36378), .B(n36379), .Z(n31756) );
  XNOR U35585 ( .A(n31752), .B(n31754), .Z(n36379) );
  XNOR U35586 ( .A(q[1]), .B(DB[646]), .Z(n31754) );
  XNOR U35587 ( .A(q[4]), .B(DB[649]), .Z(n31752) );
  IV U35588 ( .A(n31751), .Z(n36378) );
  XNOR U35589 ( .A(n31749), .B(n36380), .Z(n31751) );
  XNOR U35590 ( .A(q[3]), .B(DB[648]), .Z(n36380) );
  XNOR U35591 ( .A(q[2]), .B(DB[647]), .Z(n31749) );
  XOR U35592 ( .A(n36381), .B(n31647), .Z(n31575) );
  XOR U35593 ( .A(n36382), .B(n31639), .Z(n31647) );
  XOR U35594 ( .A(n36383), .B(n31628), .Z(n31639) );
  XNOR U35595 ( .A(q[14]), .B(DB[674]), .Z(n31628) );
  IV U35596 ( .A(n31627), .Z(n36383) );
  XNOR U35597 ( .A(n31625), .B(n36384), .Z(n31627) );
  XNOR U35598 ( .A(q[13]), .B(DB[673]), .Z(n36384) );
  XNOR U35599 ( .A(q[12]), .B(DB[672]), .Z(n31625) );
  IV U35600 ( .A(n31638), .Z(n36382) );
  XOR U35601 ( .A(n36385), .B(n36386), .Z(n31638) );
  XNOR U35602 ( .A(n31634), .B(n31636), .Z(n36386) );
  XNOR U35603 ( .A(q[8]), .B(DB[668]), .Z(n31636) );
  XNOR U35604 ( .A(q[11]), .B(DB[671]), .Z(n31634) );
  IV U35605 ( .A(n31633), .Z(n36385) );
  XNOR U35606 ( .A(n31631), .B(n36387), .Z(n31633) );
  XNOR U35607 ( .A(q[10]), .B(DB[670]), .Z(n36387) );
  XNOR U35608 ( .A(q[9]), .B(DB[669]), .Z(n31631) );
  IV U35609 ( .A(n31646), .Z(n36381) );
  XOR U35610 ( .A(n36388), .B(n36389), .Z(n31646) );
  XNOR U35611 ( .A(n31663), .B(n31644), .Z(n36389) );
  XNOR U35612 ( .A(q[0]), .B(DB[660]), .Z(n31644) );
  XOR U35613 ( .A(n36390), .B(n31652), .Z(n31663) );
  XNOR U35614 ( .A(q[7]), .B(DB[667]), .Z(n31652) );
  IV U35615 ( .A(n31651), .Z(n36390) );
  XNOR U35616 ( .A(n31649), .B(n36391), .Z(n31651) );
  XNOR U35617 ( .A(q[6]), .B(DB[666]), .Z(n36391) );
  XNOR U35618 ( .A(q[5]), .B(DB[665]), .Z(n31649) );
  IV U35619 ( .A(n31662), .Z(n36388) );
  XOR U35620 ( .A(n36392), .B(n36393), .Z(n31662) );
  XNOR U35621 ( .A(n31658), .B(n31660), .Z(n36393) );
  XNOR U35622 ( .A(q[1]), .B(DB[661]), .Z(n31660) );
  XNOR U35623 ( .A(q[4]), .B(DB[664]), .Z(n31658) );
  IV U35624 ( .A(n31657), .Z(n36392) );
  XNOR U35625 ( .A(n31655), .B(n36394), .Z(n31657) );
  XNOR U35626 ( .A(q[3]), .B(DB[663]), .Z(n36394) );
  XNOR U35627 ( .A(q[2]), .B(DB[662]), .Z(n31655) );
  XOR U35628 ( .A(n36395), .B(n31553), .Z(n31481) );
  XOR U35629 ( .A(n36396), .B(n31545), .Z(n31553) );
  XOR U35630 ( .A(n36397), .B(n31534), .Z(n31545) );
  XNOR U35631 ( .A(q[14]), .B(DB[689]), .Z(n31534) );
  IV U35632 ( .A(n31533), .Z(n36397) );
  XNOR U35633 ( .A(n31531), .B(n36398), .Z(n31533) );
  XNOR U35634 ( .A(q[13]), .B(DB[688]), .Z(n36398) );
  XNOR U35635 ( .A(q[12]), .B(DB[687]), .Z(n31531) );
  IV U35636 ( .A(n31544), .Z(n36396) );
  XOR U35637 ( .A(n36399), .B(n36400), .Z(n31544) );
  XNOR U35638 ( .A(n31540), .B(n31542), .Z(n36400) );
  XNOR U35639 ( .A(q[8]), .B(DB[683]), .Z(n31542) );
  XNOR U35640 ( .A(q[11]), .B(DB[686]), .Z(n31540) );
  IV U35641 ( .A(n31539), .Z(n36399) );
  XNOR U35642 ( .A(n31537), .B(n36401), .Z(n31539) );
  XNOR U35643 ( .A(q[10]), .B(DB[685]), .Z(n36401) );
  XNOR U35644 ( .A(q[9]), .B(DB[684]), .Z(n31537) );
  IV U35645 ( .A(n31552), .Z(n36395) );
  XOR U35646 ( .A(n36402), .B(n36403), .Z(n31552) );
  XNOR U35647 ( .A(n31569), .B(n31550), .Z(n36403) );
  XNOR U35648 ( .A(q[0]), .B(DB[675]), .Z(n31550) );
  XOR U35649 ( .A(n36404), .B(n31558), .Z(n31569) );
  XNOR U35650 ( .A(q[7]), .B(DB[682]), .Z(n31558) );
  IV U35651 ( .A(n31557), .Z(n36404) );
  XNOR U35652 ( .A(n31555), .B(n36405), .Z(n31557) );
  XNOR U35653 ( .A(q[6]), .B(DB[681]), .Z(n36405) );
  XNOR U35654 ( .A(q[5]), .B(DB[680]), .Z(n31555) );
  IV U35655 ( .A(n31568), .Z(n36402) );
  XOR U35656 ( .A(n36406), .B(n36407), .Z(n31568) );
  XNOR U35657 ( .A(n31564), .B(n31566), .Z(n36407) );
  XNOR U35658 ( .A(q[1]), .B(DB[676]), .Z(n31566) );
  XNOR U35659 ( .A(q[4]), .B(DB[679]), .Z(n31564) );
  IV U35660 ( .A(n31563), .Z(n36406) );
  XNOR U35661 ( .A(n31561), .B(n36408), .Z(n31563) );
  XNOR U35662 ( .A(q[3]), .B(DB[678]), .Z(n36408) );
  XNOR U35663 ( .A(q[2]), .B(DB[677]), .Z(n31561) );
  XOR U35664 ( .A(n36409), .B(n31459), .Z(n31387) );
  XOR U35665 ( .A(n36410), .B(n31451), .Z(n31459) );
  XOR U35666 ( .A(n36411), .B(n31440), .Z(n31451) );
  XNOR U35667 ( .A(q[14]), .B(DB[704]), .Z(n31440) );
  IV U35668 ( .A(n31439), .Z(n36411) );
  XNOR U35669 ( .A(n31437), .B(n36412), .Z(n31439) );
  XNOR U35670 ( .A(q[13]), .B(DB[703]), .Z(n36412) );
  XNOR U35671 ( .A(q[12]), .B(DB[702]), .Z(n31437) );
  IV U35672 ( .A(n31450), .Z(n36410) );
  XOR U35673 ( .A(n36413), .B(n36414), .Z(n31450) );
  XNOR U35674 ( .A(n31446), .B(n31448), .Z(n36414) );
  XNOR U35675 ( .A(q[8]), .B(DB[698]), .Z(n31448) );
  XNOR U35676 ( .A(q[11]), .B(DB[701]), .Z(n31446) );
  IV U35677 ( .A(n31445), .Z(n36413) );
  XNOR U35678 ( .A(n31443), .B(n36415), .Z(n31445) );
  XNOR U35679 ( .A(q[10]), .B(DB[700]), .Z(n36415) );
  XNOR U35680 ( .A(q[9]), .B(DB[699]), .Z(n31443) );
  IV U35681 ( .A(n31458), .Z(n36409) );
  XOR U35682 ( .A(n36416), .B(n36417), .Z(n31458) );
  XNOR U35683 ( .A(n31475), .B(n31456), .Z(n36417) );
  XNOR U35684 ( .A(q[0]), .B(DB[690]), .Z(n31456) );
  XOR U35685 ( .A(n36418), .B(n31464), .Z(n31475) );
  XNOR U35686 ( .A(q[7]), .B(DB[697]), .Z(n31464) );
  IV U35687 ( .A(n31463), .Z(n36418) );
  XNOR U35688 ( .A(n31461), .B(n36419), .Z(n31463) );
  XNOR U35689 ( .A(q[6]), .B(DB[696]), .Z(n36419) );
  XNOR U35690 ( .A(q[5]), .B(DB[695]), .Z(n31461) );
  IV U35691 ( .A(n31474), .Z(n36416) );
  XOR U35692 ( .A(n36420), .B(n36421), .Z(n31474) );
  XNOR U35693 ( .A(n31470), .B(n31472), .Z(n36421) );
  XNOR U35694 ( .A(q[1]), .B(DB[691]), .Z(n31472) );
  XNOR U35695 ( .A(q[4]), .B(DB[694]), .Z(n31470) );
  IV U35696 ( .A(n31469), .Z(n36420) );
  XNOR U35697 ( .A(n31467), .B(n36422), .Z(n31469) );
  XNOR U35698 ( .A(q[3]), .B(DB[693]), .Z(n36422) );
  XNOR U35699 ( .A(q[2]), .B(DB[692]), .Z(n31467) );
  XOR U35700 ( .A(n36423), .B(n31365), .Z(n31293) );
  XOR U35701 ( .A(n36424), .B(n31357), .Z(n31365) );
  XOR U35702 ( .A(n36425), .B(n31346), .Z(n31357) );
  XNOR U35703 ( .A(q[14]), .B(DB[719]), .Z(n31346) );
  IV U35704 ( .A(n31345), .Z(n36425) );
  XNOR U35705 ( .A(n31343), .B(n36426), .Z(n31345) );
  XNOR U35706 ( .A(q[13]), .B(DB[718]), .Z(n36426) );
  XNOR U35707 ( .A(q[12]), .B(DB[717]), .Z(n31343) );
  IV U35708 ( .A(n31356), .Z(n36424) );
  XOR U35709 ( .A(n36427), .B(n36428), .Z(n31356) );
  XNOR U35710 ( .A(n31352), .B(n31354), .Z(n36428) );
  XNOR U35711 ( .A(q[8]), .B(DB[713]), .Z(n31354) );
  XNOR U35712 ( .A(q[11]), .B(DB[716]), .Z(n31352) );
  IV U35713 ( .A(n31351), .Z(n36427) );
  XNOR U35714 ( .A(n31349), .B(n36429), .Z(n31351) );
  XNOR U35715 ( .A(q[10]), .B(DB[715]), .Z(n36429) );
  XNOR U35716 ( .A(q[9]), .B(DB[714]), .Z(n31349) );
  IV U35717 ( .A(n31364), .Z(n36423) );
  XOR U35718 ( .A(n36430), .B(n36431), .Z(n31364) );
  XNOR U35719 ( .A(n31381), .B(n31362), .Z(n36431) );
  XNOR U35720 ( .A(q[0]), .B(DB[705]), .Z(n31362) );
  XOR U35721 ( .A(n36432), .B(n31370), .Z(n31381) );
  XNOR U35722 ( .A(q[7]), .B(DB[712]), .Z(n31370) );
  IV U35723 ( .A(n31369), .Z(n36432) );
  XNOR U35724 ( .A(n31367), .B(n36433), .Z(n31369) );
  XNOR U35725 ( .A(q[6]), .B(DB[711]), .Z(n36433) );
  XNOR U35726 ( .A(q[5]), .B(DB[710]), .Z(n31367) );
  IV U35727 ( .A(n31380), .Z(n36430) );
  XOR U35728 ( .A(n36434), .B(n36435), .Z(n31380) );
  XNOR U35729 ( .A(n31376), .B(n31378), .Z(n36435) );
  XNOR U35730 ( .A(q[1]), .B(DB[706]), .Z(n31378) );
  XNOR U35731 ( .A(q[4]), .B(DB[709]), .Z(n31376) );
  IV U35732 ( .A(n31375), .Z(n36434) );
  XNOR U35733 ( .A(n31373), .B(n36436), .Z(n31375) );
  XNOR U35734 ( .A(q[3]), .B(DB[708]), .Z(n36436) );
  XNOR U35735 ( .A(q[2]), .B(DB[707]), .Z(n31373) );
  XOR U35736 ( .A(n36437), .B(n31271), .Z(n31199) );
  XOR U35737 ( .A(n36438), .B(n31263), .Z(n31271) );
  XOR U35738 ( .A(n36439), .B(n31252), .Z(n31263) );
  XNOR U35739 ( .A(q[14]), .B(DB[734]), .Z(n31252) );
  IV U35740 ( .A(n31251), .Z(n36439) );
  XNOR U35741 ( .A(n31249), .B(n36440), .Z(n31251) );
  XNOR U35742 ( .A(q[13]), .B(DB[733]), .Z(n36440) );
  XNOR U35743 ( .A(q[12]), .B(DB[732]), .Z(n31249) );
  IV U35744 ( .A(n31262), .Z(n36438) );
  XOR U35745 ( .A(n36441), .B(n36442), .Z(n31262) );
  XNOR U35746 ( .A(n31258), .B(n31260), .Z(n36442) );
  XNOR U35747 ( .A(q[8]), .B(DB[728]), .Z(n31260) );
  XNOR U35748 ( .A(q[11]), .B(DB[731]), .Z(n31258) );
  IV U35749 ( .A(n31257), .Z(n36441) );
  XNOR U35750 ( .A(n31255), .B(n36443), .Z(n31257) );
  XNOR U35751 ( .A(q[10]), .B(DB[730]), .Z(n36443) );
  XNOR U35752 ( .A(q[9]), .B(DB[729]), .Z(n31255) );
  IV U35753 ( .A(n31270), .Z(n36437) );
  XOR U35754 ( .A(n36444), .B(n36445), .Z(n31270) );
  XNOR U35755 ( .A(n31287), .B(n31268), .Z(n36445) );
  XNOR U35756 ( .A(q[0]), .B(DB[720]), .Z(n31268) );
  XOR U35757 ( .A(n36446), .B(n31276), .Z(n31287) );
  XNOR U35758 ( .A(q[7]), .B(DB[727]), .Z(n31276) );
  IV U35759 ( .A(n31275), .Z(n36446) );
  XNOR U35760 ( .A(n31273), .B(n36447), .Z(n31275) );
  XNOR U35761 ( .A(q[6]), .B(DB[726]), .Z(n36447) );
  XNOR U35762 ( .A(q[5]), .B(DB[725]), .Z(n31273) );
  IV U35763 ( .A(n31286), .Z(n36444) );
  XOR U35764 ( .A(n36448), .B(n36449), .Z(n31286) );
  XNOR U35765 ( .A(n31282), .B(n31284), .Z(n36449) );
  XNOR U35766 ( .A(q[1]), .B(DB[721]), .Z(n31284) );
  XNOR U35767 ( .A(q[4]), .B(DB[724]), .Z(n31282) );
  IV U35768 ( .A(n31281), .Z(n36448) );
  XNOR U35769 ( .A(n31279), .B(n36450), .Z(n31281) );
  XNOR U35770 ( .A(q[3]), .B(DB[723]), .Z(n36450) );
  XNOR U35771 ( .A(q[2]), .B(DB[722]), .Z(n31279) );
  XOR U35772 ( .A(n36451), .B(n31177), .Z(n31105) );
  XOR U35773 ( .A(n36452), .B(n31169), .Z(n31177) );
  XOR U35774 ( .A(n36453), .B(n31158), .Z(n31169) );
  XNOR U35775 ( .A(q[14]), .B(DB[749]), .Z(n31158) );
  IV U35776 ( .A(n31157), .Z(n36453) );
  XNOR U35777 ( .A(n31155), .B(n36454), .Z(n31157) );
  XNOR U35778 ( .A(q[13]), .B(DB[748]), .Z(n36454) );
  XNOR U35779 ( .A(q[12]), .B(DB[747]), .Z(n31155) );
  IV U35780 ( .A(n31168), .Z(n36452) );
  XOR U35781 ( .A(n36455), .B(n36456), .Z(n31168) );
  XNOR U35782 ( .A(n31164), .B(n31166), .Z(n36456) );
  XNOR U35783 ( .A(q[8]), .B(DB[743]), .Z(n31166) );
  XNOR U35784 ( .A(q[11]), .B(DB[746]), .Z(n31164) );
  IV U35785 ( .A(n31163), .Z(n36455) );
  XNOR U35786 ( .A(n31161), .B(n36457), .Z(n31163) );
  XNOR U35787 ( .A(q[10]), .B(DB[745]), .Z(n36457) );
  XNOR U35788 ( .A(q[9]), .B(DB[744]), .Z(n31161) );
  IV U35789 ( .A(n31176), .Z(n36451) );
  XOR U35790 ( .A(n36458), .B(n36459), .Z(n31176) );
  XNOR U35791 ( .A(n31193), .B(n31174), .Z(n36459) );
  XNOR U35792 ( .A(q[0]), .B(DB[735]), .Z(n31174) );
  XOR U35793 ( .A(n36460), .B(n31182), .Z(n31193) );
  XNOR U35794 ( .A(q[7]), .B(DB[742]), .Z(n31182) );
  IV U35795 ( .A(n31181), .Z(n36460) );
  XNOR U35796 ( .A(n31179), .B(n36461), .Z(n31181) );
  XNOR U35797 ( .A(q[6]), .B(DB[741]), .Z(n36461) );
  XNOR U35798 ( .A(q[5]), .B(DB[740]), .Z(n31179) );
  IV U35799 ( .A(n31192), .Z(n36458) );
  XOR U35800 ( .A(n36462), .B(n36463), .Z(n31192) );
  XNOR U35801 ( .A(n31188), .B(n31190), .Z(n36463) );
  XNOR U35802 ( .A(q[1]), .B(DB[736]), .Z(n31190) );
  XNOR U35803 ( .A(q[4]), .B(DB[739]), .Z(n31188) );
  IV U35804 ( .A(n31187), .Z(n36462) );
  XNOR U35805 ( .A(n31185), .B(n36464), .Z(n31187) );
  XNOR U35806 ( .A(q[3]), .B(DB[738]), .Z(n36464) );
  XNOR U35807 ( .A(q[2]), .B(DB[737]), .Z(n31185) );
  XOR U35808 ( .A(n36465), .B(n31083), .Z(n31011) );
  XOR U35809 ( .A(n36466), .B(n31075), .Z(n31083) );
  XOR U35810 ( .A(n36467), .B(n31064), .Z(n31075) );
  XNOR U35811 ( .A(q[14]), .B(DB[764]), .Z(n31064) );
  IV U35812 ( .A(n31063), .Z(n36467) );
  XNOR U35813 ( .A(n31061), .B(n36468), .Z(n31063) );
  XNOR U35814 ( .A(q[13]), .B(DB[763]), .Z(n36468) );
  XNOR U35815 ( .A(q[12]), .B(DB[762]), .Z(n31061) );
  IV U35816 ( .A(n31074), .Z(n36466) );
  XOR U35817 ( .A(n36469), .B(n36470), .Z(n31074) );
  XNOR U35818 ( .A(n31070), .B(n31072), .Z(n36470) );
  XNOR U35819 ( .A(q[8]), .B(DB[758]), .Z(n31072) );
  XNOR U35820 ( .A(q[11]), .B(DB[761]), .Z(n31070) );
  IV U35821 ( .A(n31069), .Z(n36469) );
  XNOR U35822 ( .A(n31067), .B(n36471), .Z(n31069) );
  XNOR U35823 ( .A(q[10]), .B(DB[760]), .Z(n36471) );
  XNOR U35824 ( .A(q[9]), .B(DB[759]), .Z(n31067) );
  IV U35825 ( .A(n31082), .Z(n36465) );
  XOR U35826 ( .A(n36472), .B(n36473), .Z(n31082) );
  XNOR U35827 ( .A(n31099), .B(n31080), .Z(n36473) );
  XNOR U35828 ( .A(q[0]), .B(DB[750]), .Z(n31080) );
  XOR U35829 ( .A(n36474), .B(n31088), .Z(n31099) );
  XNOR U35830 ( .A(q[7]), .B(DB[757]), .Z(n31088) );
  IV U35831 ( .A(n31087), .Z(n36474) );
  XNOR U35832 ( .A(n31085), .B(n36475), .Z(n31087) );
  XNOR U35833 ( .A(q[6]), .B(DB[756]), .Z(n36475) );
  XNOR U35834 ( .A(q[5]), .B(DB[755]), .Z(n31085) );
  IV U35835 ( .A(n31098), .Z(n36472) );
  XOR U35836 ( .A(n36476), .B(n36477), .Z(n31098) );
  XNOR U35837 ( .A(n31094), .B(n31096), .Z(n36477) );
  XNOR U35838 ( .A(q[1]), .B(DB[751]), .Z(n31096) );
  XNOR U35839 ( .A(q[4]), .B(DB[754]), .Z(n31094) );
  IV U35840 ( .A(n31093), .Z(n36476) );
  XNOR U35841 ( .A(n31091), .B(n36478), .Z(n31093) );
  XNOR U35842 ( .A(q[3]), .B(DB[753]), .Z(n36478) );
  XNOR U35843 ( .A(q[2]), .B(DB[752]), .Z(n31091) );
  XOR U35844 ( .A(n36479), .B(n30989), .Z(n30917) );
  XOR U35845 ( .A(n36480), .B(n30981), .Z(n30989) );
  XOR U35846 ( .A(n36481), .B(n30970), .Z(n30981) );
  XNOR U35847 ( .A(q[14]), .B(DB[779]), .Z(n30970) );
  IV U35848 ( .A(n30969), .Z(n36481) );
  XNOR U35849 ( .A(n30967), .B(n36482), .Z(n30969) );
  XNOR U35850 ( .A(q[13]), .B(DB[778]), .Z(n36482) );
  XNOR U35851 ( .A(q[12]), .B(DB[777]), .Z(n30967) );
  IV U35852 ( .A(n30980), .Z(n36480) );
  XOR U35853 ( .A(n36483), .B(n36484), .Z(n30980) );
  XNOR U35854 ( .A(n30976), .B(n30978), .Z(n36484) );
  XNOR U35855 ( .A(q[8]), .B(DB[773]), .Z(n30978) );
  XNOR U35856 ( .A(q[11]), .B(DB[776]), .Z(n30976) );
  IV U35857 ( .A(n30975), .Z(n36483) );
  XNOR U35858 ( .A(n30973), .B(n36485), .Z(n30975) );
  XNOR U35859 ( .A(q[10]), .B(DB[775]), .Z(n36485) );
  XNOR U35860 ( .A(q[9]), .B(DB[774]), .Z(n30973) );
  IV U35861 ( .A(n30988), .Z(n36479) );
  XOR U35862 ( .A(n36486), .B(n36487), .Z(n30988) );
  XNOR U35863 ( .A(n31005), .B(n30986), .Z(n36487) );
  XNOR U35864 ( .A(q[0]), .B(DB[765]), .Z(n30986) );
  XOR U35865 ( .A(n36488), .B(n30994), .Z(n31005) );
  XNOR U35866 ( .A(q[7]), .B(DB[772]), .Z(n30994) );
  IV U35867 ( .A(n30993), .Z(n36488) );
  XNOR U35868 ( .A(n30991), .B(n36489), .Z(n30993) );
  XNOR U35869 ( .A(q[6]), .B(DB[771]), .Z(n36489) );
  XNOR U35870 ( .A(q[5]), .B(DB[770]), .Z(n30991) );
  IV U35871 ( .A(n31004), .Z(n36486) );
  XOR U35872 ( .A(n36490), .B(n36491), .Z(n31004) );
  XNOR U35873 ( .A(n31000), .B(n31002), .Z(n36491) );
  XNOR U35874 ( .A(q[1]), .B(DB[766]), .Z(n31002) );
  XNOR U35875 ( .A(q[4]), .B(DB[769]), .Z(n31000) );
  IV U35876 ( .A(n30999), .Z(n36490) );
  XNOR U35877 ( .A(n30997), .B(n36492), .Z(n30999) );
  XNOR U35878 ( .A(q[3]), .B(DB[768]), .Z(n36492) );
  XNOR U35879 ( .A(q[2]), .B(DB[767]), .Z(n30997) );
  XOR U35880 ( .A(n36493), .B(n30895), .Z(n30823) );
  XOR U35881 ( .A(n36494), .B(n30887), .Z(n30895) );
  XOR U35882 ( .A(n36495), .B(n30876), .Z(n30887) );
  XNOR U35883 ( .A(q[14]), .B(DB[794]), .Z(n30876) );
  IV U35884 ( .A(n30875), .Z(n36495) );
  XNOR U35885 ( .A(n30873), .B(n36496), .Z(n30875) );
  XNOR U35886 ( .A(q[13]), .B(DB[793]), .Z(n36496) );
  XNOR U35887 ( .A(q[12]), .B(DB[792]), .Z(n30873) );
  IV U35888 ( .A(n30886), .Z(n36494) );
  XOR U35889 ( .A(n36497), .B(n36498), .Z(n30886) );
  XNOR U35890 ( .A(n30882), .B(n30884), .Z(n36498) );
  XNOR U35891 ( .A(q[8]), .B(DB[788]), .Z(n30884) );
  XNOR U35892 ( .A(q[11]), .B(DB[791]), .Z(n30882) );
  IV U35893 ( .A(n30881), .Z(n36497) );
  XNOR U35894 ( .A(n30879), .B(n36499), .Z(n30881) );
  XNOR U35895 ( .A(q[10]), .B(DB[790]), .Z(n36499) );
  XNOR U35896 ( .A(q[9]), .B(DB[789]), .Z(n30879) );
  IV U35897 ( .A(n30894), .Z(n36493) );
  XOR U35898 ( .A(n36500), .B(n36501), .Z(n30894) );
  XNOR U35899 ( .A(n30911), .B(n30892), .Z(n36501) );
  XNOR U35900 ( .A(q[0]), .B(DB[780]), .Z(n30892) );
  XOR U35901 ( .A(n36502), .B(n30900), .Z(n30911) );
  XNOR U35902 ( .A(q[7]), .B(DB[787]), .Z(n30900) );
  IV U35903 ( .A(n30899), .Z(n36502) );
  XNOR U35904 ( .A(n30897), .B(n36503), .Z(n30899) );
  XNOR U35905 ( .A(q[6]), .B(DB[786]), .Z(n36503) );
  XNOR U35906 ( .A(q[5]), .B(DB[785]), .Z(n30897) );
  IV U35907 ( .A(n30910), .Z(n36500) );
  XOR U35908 ( .A(n36504), .B(n36505), .Z(n30910) );
  XNOR U35909 ( .A(n30906), .B(n30908), .Z(n36505) );
  XNOR U35910 ( .A(q[1]), .B(DB[781]), .Z(n30908) );
  XNOR U35911 ( .A(q[4]), .B(DB[784]), .Z(n30906) );
  IV U35912 ( .A(n30905), .Z(n36504) );
  XNOR U35913 ( .A(n30903), .B(n36506), .Z(n30905) );
  XNOR U35914 ( .A(q[3]), .B(DB[783]), .Z(n36506) );
  XNOR U35915 ( .A(q[2]), .B(DB[782]), .Z(n30903) );
  XOR U35916 ( .A(n36507), .B(n30801), .Z(n30729) );
  XOR U35917 ( .A(n36508), .B(n30793), .Z(n30801) );
  XOR U35918 ( .A(n36509), .B(n30782), .Z(n30793) );
  XNOR U35919 ( .A(q[14]), .B(DB[809]), .Z(n30782) );
  IV U35920 ( .A(n30781), .Z(n36509) );
  XNOR U35921 ( .A(n30779), .B(n36510), .Z(n30781) );
  XNOR U35922 ( .A(q[13]), .B(DB[808]), .Z(n36510) );
  XNOR U35923 ( .A(q[12]), .B(DB[807]), .Z(n30779) );
  IV U35924 ( .A(n30792), .Z(n36508) );
  XOR U35925 ( .A(n36511), .B(n36512), .Z(n30792) );
  XNOR U35926 ( .A(n30788), .B(n30790), .Z(n36512) );
  XNOR U35927 ( .A(q[8]), .B(DB[803]), .Z(n30790) );
  XNOR U35928 ( .A(q[11]), .B(DB[806]), .Z(n30788) );
  IV U35929 ( .A(n30787), .Z(n36511) );
  XNOR U35930 ( .A(n30785), .B(n36513), .Z(n30787) );
  XNOR U35931 ( .A(q[10]), .B(DB[805]), .Z(n36513) );
  XNOR U35932 ( .A(q[9]), .B(DB[804]), .Z(n30785) );
  IV U35933 ( .A(n30800), .Z(n36507) );
  XOR U35934 ( .A(n36514), .B(n36515), .Z(n30800) );
  XNOR U35935 ( .A(n30817), .B(n30798), .Z(n36515) );
  XNOR U35936 ( .A(q[0]), .B(DB[795]), .Z(n30798) );
  XOR U35937 ( .A(n36516), .B(n30806), .Z(n30817) );
  XNOR U35938 ( .A(q[7]), .B(DB[802]), .Z(n30806) );
  IV U35939 ( .A(n30805), .Z(n36516) );
  XNOR U35940 ( .A(n30803), .B(n36517), .Z(n30805) );
  XNOR U35941 ( .A(q[6]), .B(DB[801]), .Z(n36517) );
  XNOR U35942 ( .A(q[5]), .B(DB[800]), .Z(n30803) );
  IV U35943 ( .A(n30816), .Z(n36514) );
  XOR U35944 ( .A(n36518), .B(n36519), .Z(n30816) );
  XNOR U35945 ( .A(n30812), .B(n30814), .Z(n36519) );
  XNOR U35946 ( .A(q[1]), .B(DB[796]), .Z(n30814) );
  XNOR U35947 ( .A(q[4]), .B(DB[799]), .Z(n30812) );
  IV U35948 ( .A(n30811), .Z(n36518) );
  XNOR U35949 ( .A(n30809), .B(n36520), .Z(n30811) );
  XNOR U35950 ( .A(q[3]), .B(DB[798]), .Z(n36520) );
  XNOR U35951 ( .A(q[2]), .B(DB[797]), .Z(n30809) );
  XOR U35952 ( .A(n36521), .B(n30707), .Z(n30635) );
  XOR U35953 ( .A(n36522), .B(n30699), .Z(n30707) );
  XOR U35954 ( .A(n36523), .B(n30688), .Z(n30699) );
  XNOR U35955 ( .A(q[14]), .B(DB[824]), .Z(n30688) );
  IV U35956 ( .A(n30687), .Z(n36523) );
  XNOR U35957 ( .A(n30685), .B(n36524), .Z(n30687) );
  XNOR U35958 ( .A(q[13]), .B(DB[823]), .Z(n36524) );
  XNOR U35959 ( .A(q[12]), .B(DB[822]), .Z(n30685) );
  IV U35960 ( .A(n30698), .Z(n36522) );
  XOR U35961 ( .A(n36525), .B(n36526), .Z(n30698) );
  XNOR U35962 ( .A(n30694), .B(n30696), .Z(n36526) );
  XNOR U35963 ( .A(q[8]), .B(DB[818]), .Z(n30696) );
  XNOR U35964 ( .A(q[11]), .B(DB[821]), .Z(n30694) );
  IV U35965 ( .A(n30693), .Z(n36525) );
  XNOR U35966 ( .A(n30691), .B(n36527), .Z(n30693) );
  XNOR U35967 ( .A(q[10]), .B(DB[820]), .Z(n36527) );
  XNOR U35968 ( .A(q[9]), .B(DB[819]), .Z(n30691) );
  IV U35969 ( .A(n30706), .Z(n36521) );
  XOR U35970 ( .A(n36528), .B(n36529), .Z(n30706) );
  XNOR U35971 ( .A(n30723), .B(n30704), .Z(n36529) );
  XNOR U35972 ( .A(q[0]), .B(DB[810]), .Z(n30704) );
  XOR U35973 ( .A(n36530), .B(n30712), .Z(n30723) );
  XNOR U35974 ( .A(q[7]), .B(DB[817]), .Z(n30712) );
  IV U35975 ( .A(n30711), .Z(n36530) );
  XNOR U35976 ( .A(n30709), .B(n36531), .Z(n30711) );
  XNOR U35977 ( .A(q[6]), .B(DB[816]), .Z(n36531) );
  XNOR U35978 ( .A(q[5]), .B(DB[815]), .Z(n30709) );
  IV U35979 ( .A(n30722), .Z(n36528) );
  XOR U35980 ( .A(n36532), .B(n36533), .Z(n30722) );
  XNOR U35981 ( .A(n30718), .B(n30720), .Z(n36533) );
  XNOR U35982 ( .A(q[1]), .B(DB[811]), .Z(n30720) );
  XNOR U35983 ( .A(q[4]), .B(DB[814]), .Z(n30718) );
  IV U35984 ( .A(n30717), .Z(n36532) );
  XNOR U35985 ( .A(n30715), .B(n36534), .Z(n30717) );
  XNOR U35986 ( .A(q[3]), .B(DB[813]), .Z(n36534) );
  XNOR U35987 ( .A(q[2]), .B(DB[812]), .Z(n30715) );
  XOR U35988 ( .A(n36535), .B(n30613), .Z(n30541) );
  XOR U35989 ( .A(n36536), .B(n30605), .Z(n30613) );
  XOR U35990 ( .A(n36537), .B(n30594), .Z(n30605) );
  XNOR U35991 ( .A(q[14]), .B(DB[839]), .Z(n30594) );
  IV U35992 ( .A(n30593), .Z(n36537) );
  XNOR U35993 ( .A(n30591), .B(n36538), .Z(n30593) );
  XNOR U35994 ( .A(q[13]), .B(DB[838]), .Z(n36538) );
  XNOR U35995 ( .A(q[12]), .B(DB[837]), .Z(n30591) );
  IV U35996 ( .A(n30604), .Z(n36536) );
  XOR U35997 ( .A(n36539), .B(n36540), .Z(n30604) );
  XNOR U35998 ( .A(n30600), .B(n30602), .Z(n36540) );
  XNOR U35999 ( .A(q[8]), .B(DB[833]), .Z(n30602) );
  XNOR U36000 ( .A(q[11]), .B(DB[836]), .Z(n30600) );
  IV U36001 ( .A(n30599), .Z(n36539) );
  XNOR U36002 ( .A(n30597), .B(n36541), .Z(n30599) );
  XNOR U36003 ( .A(q[10]), .B(DB[835]), .Z(n36541) );
  XNOR U36004 ( .A(q[9]), .B(DB[834]), .Z(n30597) );
  IV U36005 ( .A(n30612), .Z(n36535) );
  XOR U36006 ( .A(n36542), .B(n36543), .Z(n30612) );
  XNOR U36007 ( .A(n30629), .B(n30610), .Z(n36543) );
  XNOR U36008 ( .A(q[0]), .B(DB[825]), .Z(n30610) );
  XOR U36009 ( .A(n36544), .B(n30618), .Z(n30629) );
  XNOR U36010 ( .A(q[7]), .B(DB[832]), .Z(n30618) );
  IV U36011 ( .A(n30617), .Z(n36544) );
  XNOR U36012 ( .A(n30615), .B(n36545), .Z(n30617) );
  XNOR U36013 ( .A(q[6]), .B(DB[831]), .Z(n36545) );
  XNOR U36014 ( .A(q[5]), .B(DB[830]), .Z(n30615) );
  IV U36015 ( .A(n30628), .Z(n36542) );
  XOR U36016 ( .A(n36546), .B(n36547), .Z(n30628) );
  XNOR U36017 ( .A(n30624), .B(n30626), .Z(n36547) );
  XNOR U36018 ( .A(q[1]), .B(DB[826]), .Z(n30626) );
  XNOR U36019 ( .A(q[4]), .B(DB[829]), .Z(n30624) );
  IV U36020 ( .A(n30623), .Z(n36546) );
  XNOR U36021 ( .A(n30621), .B(n36548), .Z(n30623) );
  XNOR U36022 ( .A(q[3]), .B(DB[828]), .Z(n36548) );
  XNOR U36023 ( .A(q[2]), .B(DB[827]), .Z(n30621) );
  XOR U36024 ( .A(n36549), .B(n30519), .Z(n30447) );
  XOR U36025 ( .A(n36550), .B(n30511), .Z(n30519) );
  XOR U36026 ( .A(n36551), .B(n30500), .Z(n30511) );
  XNOR U36027 ( .A(q[14]), .B(DB[854]), .Z(n30500) );
  IV U36028 ( .A(n30499), .Z(n36551) );
  XNOR U36029 ( .A(n30497), .B(n36552), .Z(n30499) );
  XNOR U36030 ( .A(q[13]), .B(DB[853]), .Z(n36552) );
  XNOR U36031 ( .A(q[12]), .B(DB[852]), .Z(n30497) );
  IV U36032 ( .A(n30510), .Z(n36550) );
  XOR U36033 ( .A(n36553), .B(n36554), .Z(n30510) );
  XNOR U36034 ( .A(n30506), .B(n30508), .Z(n36554) );
  XNOR U36035 ( .A(q[8]), .B(DB[848]), .Z(n30508) );
  XNOR U36036 ( .A(q[11]), .B(DB[851]), .Z(n30506) );
  IV U36037 ( .A(n30505), .Z(n36553) );
  XNOR U36038 ( .A(n30503), .B(n36555), .Z(n30505) );
  XNOR U36039 ( .A(q[10]), .B(DB[850]), .Z(n36555) );
  XNOR U36040 ( .A(q[9]), .B(DB[849]), .Z(n30503) );
  IV U36041 ( .A(n30518), .Z(n36549) );
  XOR U36042 ( .A(n36556), .B(n36557), .Z(n30518) );
  XNOR U36043 ( .A(n30535), .B(n30516), .Z(n36557) );
  XNOR U36044 ( .A(q[0]), .B(DB[840]), .Z(n30516) );
  XOR U36045 ( .A(n36558), .B(n30524), .Z(n30535) );
  XNOR U36046 ( .A(q[7]), .B(DB[847]), .Z(n30524) );
  IV U36047 ( .A(n30523), .Z(n36558) );
  XNOR U36048 ( .A(n30521), .B(n36559), .Z(n30523) );
  XNOR U36049 ( .A(q[6]), .B(DB[846]), .Z(n36559) );
  XNOR U36050 ( .A(q[5]), .B(DB[845]), .Z(n30521) );
  IV U36051 ( .A(n30534), .Z(n36556) );
  XOR U36052 ( .A(n36560), .B(n36561), .Z(n30534) );
  XNOR U36053 ( .A(n30530), .B(n30532), .Z(n36561) );
  XNOR U36054 ( .A(q[1]), .B(DB[841]), .Z(n30532) );
  XNOR U36055 ( .A(q[4]), .B(DB[844]), .Z(n30530) );
  IV U36056 ( .A(n30529), .Z(n36560) );
  XNOR U36057 ( .A(n30527), .B(n36562), .Z(n30529) );
  XNOR U36058 ( .A(q[3]), .B(DB[843]), .Z(n36562) );
  XNOR U36059 ( .A(q[2]), .B(DB[842]), .Z(n30527) );
  XOR U36060 ( .A(n36563), .B(n30425), .Z(n30353) );
  XOR U36061 ( .A(n36564), .B(n30417), .Z(n30425) );
  XOR U36062 ( .A(n36565), .B(n30406), .Z(n30417) );
  XNOR U36063 ( .A(q[14]), .B(DB[869]), .Z(n30406) );
  IV U36064 ( .A(n30405), .Z(n36565) );
  XNOR U36065 ( .A(n30403), .B(n36566), .Z(n30405) );
  XNOR U36066 ( .A(q[13]), .B(DB[868]), .Z(n36566) );
  XNOR U36067 ( .A(q[12]), .B(DB[867]), .Z(n30403) );
  IV U36068 ( .A(n30416), .Z(n36564) );
  XOR U36069 ( .A(n36567), .B(n36568), .Z(n30416) );
  XNOR U36070 ( .A(n30412), .B(n30414), .Z(n36568) );
  XNOR U36071 ( .A(q[8]), .B(DB[863]), .Z(n30414) );
  XNOR U36072 ( .A(q[11]), .B(DB[866]), .Z(n30412) );
  IV U36073 ( .A(n30411), .Z(n36567) );
  XNOR U36074 ( .A(n30409), .B(n36569), .Z(n30411) );
  XNOR U36075 ( .A(q[10]), .B(DB[865]), .Z(n36569) );
  XNOR U36076 ( .A(q[9]), .B(DB[864]), .Z(n30409) );
  IV U36077 ( .A(n30424), .Z(n36563) );
  XOR U36078 ( .A(n36570), .B(n36571), .Z(n30424) );
  XNOR U36079 ( .A(n30441), .B(n30422), .Z(n36571) );
  XNOR U36080 ( .A(q[0]), .B(DB[855]), .Z(n30422) );
  XOR U36081 ( .A(n36572), .B(n30430), .Z(n30441) );
  XNOR U36082 ( .A(q[7]), .B(DB[862]), .Z(n30430) );
  IV U36083 ( .A(n30429), .Z(n36572) );
  XNOR U36084 ( .A(n30427), .B(n36573), .Z(n30429) );
  XNOR U36085 ( .A(q[6]), .B(DB[861]), .Z(n36573) );
  XNOR U36086 ( .A(q[5]), .B(DB[860]), .Z(n30427) );
  IV U36087 ( .A(n30440), .Z(n36570) );
  XOR U36088 ( .A(n36574), .B(n36575), .Z(n30440) );
  XNOR U36089 ( .A(n30436), .B(n30438), .Z(n36575) );
  XNOR U36090 ( .A(q[1]), .B(DB[856]), .Z(n30438) );
  XNOR U36091 ( .A(q[4]), .B(DB[859]), .Z(n30436) );
  IV U36092 ( .A(n30435), .Z(n36574) );
  XNOR U36093 ( .A(n30433), .B(n36576), .Z(n30435) );
  XNOR U36094 ( .A(q[3]), .B(DB[858]), .Z(n36576) );
  XNOR U36095 ( .A(q[2]), .B(DB[857]), .Z(n30433) );
  XOR U36096 ( .A(n36577), .B(n30331), .Z(n30259) );
  XOR U36097 ( .A(n36578), .B(n30323), .Z(n30331) );
  XOR U36098 ( .A(n36579), .B(n30312), .Z(n30323) );
  XNOR U36099 ( .A(q[14]), .B(DB[884]), .Z(n30312) );
  IV U36100 ( .A(n30311), .Z(n36579) );
  XNOR U36101 ( .A(n30309), .B(n36580), .Z(n30311) );
  XNOR U36102 ( .A(q[13]), .B(DB[883]), .Z(n36580) );
  XNOR U36103 ( .A(q[12]), .B(DB[882]), .Z(n30309) );
  IV U36104 ( .A(n30322), .Z(n36578) );
  XOR U36105 ( .A(n36581), .B(n36582), .Z(n30322) );
  XNOR U36106 ( .A(n30318), .B(n30320), .Z(n36582) );
  XNOR U36107 ( .A(q[8]), .B(DB[878]), .Z(n30320) );
  XNOR U36108 ( .A(q[11]), .B(DB[881]), .Z(n30318) );
  IV U36109 ( .A(n30317), .Z(n36581) );
  XNOR U36110 ( .A(n30315), .B(n36583), .Z(n30317) );
  XNOR U36111 ( .A(q[10]), .B(DB[880]), .Z(n36583) );
  XNOR U36112 ( .A(q[9]), .B(DB[879]), .Z(n30315) );
  IV U36113 ( .A(n30330), .Z(n36577) );
  XOR U36114 ( .A(n36584), .B(n36585), .Z(n30330) );
  XNOR U36115 ( .A(n30347), .B(n30328), .Z(n36585) );
  XNOR U36116 ( .A(q[0]), .B(DB[870]), .Z(n30328) );
  XOR U36117 ( .A(n36586), .B(n30336), .Z(n30347) );
  XNOR U36118 ( .A(q[7]), .B(DB[877]), .Z(n30336) );
  IV U36119 ( .A(n30335), .Z(n36586) );
  XNOR U36120 ( .A(n30333), .B(n36587), .Z(n30335) );
  XNOR U36121 ( .A(q[6]), .B(DB[876]), .Z(n36587) );
  XNOR U36122 ( .A(q[5]), .B(DB[875]), .Z(n30333) );
  IV U36123 ( .A(n30346), .Z(n36584) );
  XOR U36124 ( .A(n36588), .B(n36589), .Z(n30346) );
  XNOR U36125 ( .A(n30342), .B(n30344), .Z(n36589) );
  XNOR U36126 ( .A(q[1]), .B(DB[871]), .Z(n30344) );
  XNOR U36127 ( .A(q[4]), .B(DB[874]), .Z(n30342) );
  IV U36128 ( .A(n30341), .Z(n36588) );
  XNOR U36129 ( .A(n30339), .B(n36590), .Z(n30341) );
  XNOR U36130 ( .A(q[3]), .B(DB[873]), .Z(n36590) );
  XNOR U36131 ( .A(q[2]), .B(DB[872]), .Z(n30339) );
  XOR U36132 ( .A(n36591), .B(n30237), .Z(n30165) );
  XOR U36133 ( .A(n36592), .B(n30229), .Z(n30237) );
  XOR U36134 ( .A(n36593), .B(n30218), .Z(n30229) );
  XNOR U36135 ( .A(q[14]), .B(DB[899]), .Z(n30218) );
  IV U36136 ( .A(n30217), .Z(n36593) );
  XNOR U36137 ( .A(n30215), .B(n36594), .Z(n30217) );
  XNOR U36138 ( .A(q[13]), .B(DB[898]), .Z(n36594) );
  XNOR U36139 ( .A(q[12]), .B(DB[897]), .Z(n30215) );
  IV U36140 ( .A(n30228), .Z(n36592) );
  XOR U36141 ( .A(n36595), .B(n36596), .Z(n30228) );
  XNOR U36142 ( .A(n30224), .B(n30226), .Z(n36596) );
  XNOR U36143 ( .A(q[8]), .B(DB[893]), .Z(n30226) );
  XNOR U36144 ( .A(q[11]), .B(DB[896]), .Z(n30224) );
  IV U36145 ( .A(n30223), .Z(n36595) );
  XNOR U36146 ( .A(n30221), .B(n36597), .Z(n30223) );
  XNOR U36147 ( .A(q[10]), .B(DB[895]), .Z(n36597) );
  XNOR U36148 ( .A(q[9]), .B(DB[894]), .Z(n30221) );
  IV U36149 ( .A(n30236), .Z(n36591) );
  XOR U36150 ( .A(n36598), .B(n36599), .Z(n30236) );
  XNOR U36151 ( .A(n30253), .B(n30234), .Z(n36599) );
  XNOR U36152 ( .A(q[0]), .B(DB[885]), .Z(n30234) );
  XOR U36153 ( .A(n36600), .B(n30242), .Z(n30253) );
  XNOR U36154 ( .A(q[7]), .B(DB[892]), .Z(n30242) );
  IV U36155 ( .A(n30241), .Z(n36600) );
  XNOR U36156 ( .A(n30239), .B(n36601), .Z(n30241) );
  XNOR U36157 ( .A(q[6]), .B(DB[891]), .Z(n36601) );
  XNOR U36158 ( .A(q[5]), .B(DB[890]), .Z(n30239) );
  IV U36159 ( .A(n30252), .Z(n36598) );
  XOR U36160 ( .A(n36602), .B(n36603), .Z(n30252) );
  XNOR U36161 ( .A(n30248), .B(n30250), .Z(n36603) );
  XNOR U36162 ( .A(q[1]), .B(DB[886]), .Z(n30250) );
  XNOR U36163 ( .A(q[4]), .B(DB[889]), .Z(n30248) );
  IV U36164 ( .A(n30247), .Z(n36602) );
  XNOR U36165 ( .A(n30245), .B(n36604), .Z(n30247) );
  XNOR U36166 ( .A(q[3]), .B(DB[888]), .Z(n36604) );
  XNOR U36167 ( .A(q[2]), .B(DB[887]), .Z(n30245) );
  XOR U36168 ( .A(n36605), .B(n30143), .Z(n30071) );
  XOR U36169 ( .A(n36606), .B(n30135), .Z(n30143) );
  XOR U36170 ( .A(n36607), .B(n30124), .Z(n30135) );
  XNOR U36171 ( .A(q[14]), .B(DB[914]), .Z(n30124) );
  IV U36172 ( .A(n30123), .Z(n36607) );
  XNOR U36173 ( .A(n30121), .B(n36608), .Z(n30123) );
  XNOR U36174 ( .A(q[13]), .B(DB[913]), .Z(n36608) );
  XNOR U36175 ( .A(q[12]), .B(DB[912]), .Z(n30121) );
  IV U36176 ( .A(n30134), .Z(n36606) );
  XOR U36177 ( .A(n36609), .B(n36610), .Z(n30134) );
  XNOR U36178 ( .A(n30130), .B(n30132), .Z(n36610) );
  XNOR U36179 ( .A(q[8]), .B(DB[908]), .Z(n30132) );
  XNOR U36180 ( .A(q[11]), .B(DB[911]), .Z(n30130) );
  IV U36181 ( .A(n30129), .Z(n36609) );
  XNOR U36182 ( .A(n30127), .B(n36611), .Z(n30129) );
  XNOR U36183 ( .A(q[10]), .B(DB[910]), .Z(n36611) );
  XNOR U36184 ( .A(q[9]), .B(DB[909]), .Z(n30127) );
  IV U36185 ( .A(n30142), .Z(n36605) );
  XOR U36186 ( .A(n36612), .B(n36613), .Z(n30142) );
  XNOR U36187 ( .A(n30159), .B(n30140), .Z(n36613) );
  XNOR U36188 ( .A(q[0]), .B(DB[900]), .Z(n30140) );
  XOR U36189 ( .A(n36614), .B(n30148), .Z(n30159) );
  XNOR U36190 ( .A(q[7]), .B(DB[907]), .Z(n30148) );
  IV U36191 ( .A(n30147), .Z(n36614) );
  XNOR U36192 ( .A(n30145), .B(n36615), .Z(n30147) );
  XNOR U36193 ( .A(q[6]), .B(DB[906]), .Z(n36615) );
  XNOR U36194 ( .A(q[5]), .B(DB[905]), .Z(n30145) );
  IV U36195 ( .A(n30158), .Z(n36612) );
  XOR U36196 ( .A(n36616), .B(n36617), .Z(n30158) );
  XNOR U36197 ( .A(n30154), .B(n30156), .Z(n36617) );
  XNOR U36198 ( .A(q[1]), .B(DB[901]), .Z(n30156) );
  XNOR U36199 ( .A(q[4]), .B(DB[904]), .Z(n30154) );
  IV U36200 ( .A(n30153), .Z(n36616) );
  XNOR U36201 ( .A(n30151), .B(n36618), .Z(n30153) );
  XNOR U36202 ( .A(q[3]), .B(DB[903]), .Z(n36618) );
  XNOR U36203 ( .A(q[2]), .B(DB[902]), .Z(n30151) );
  XOR U36204 ( .A(n36619), .B(n30049), .Z(n29977) );
  XOR U36205 ( .A(n36620), .B(n30041), .Z(n30049) );
  XOR U36206 ( .A(n36621), .B(n30030), .Z(n30041) );
  XNOR U36207 ( .A(q[14]), .B(DB[929]), .Z(n30030) );
  IV U36208 ( .A(n30029), .Z(n36621) );
  XNOR U36209 ( .A(n30027), .B(n36622), .Z(n30029) );
  XNOR U36210 ( .A(q[13]), .B(DB[928]), .Z(n36622) );
  XNOR U36211 ( .A(q[12]), .B(DB[927]), .Z(n30027) );
  IV U36212 ( .A(n30040), .Z(n36620) );
  XOR U36213 ( .A(n36623), .B(n36624), .Z(n30040) );
  XNOR U36214 ( .A(n30036), .B(n30038), .Z(n36624) );
  XNOR U36215 ( .A(q[8]), .B(DB[923]), .Z(n30038) );
  XNOR U36216 ( .A(q[11]), .B(DB[926]), .Z(n30036) );
  IV U36217 ( .A(n30035), .Z(n36623) );
  XNOR U36218 ( .A(n30033), .B(n36625), .Z(n30035) );
  XNOR U36219 ( .A(q[10]), .B(DB[925]), .Z(n36625) );
  XNOR U36220 ( .A(q[9]), .B(DB[924]), .Z(n30033) );
  IV U36221 ( .A(n30048), .Z(n36619) );
  XOR U36222 ( .A(n36626), .B(n36627), .Z(n30048) );
  XNOR U36223 ( .A(n30065), .B(n30046), .Z(n36627) );
  XNOR U36224 ( .A(q[0]), .B(DB[915]), .Z(n30046) );
  XOR U36225 ( .A(n36628), .B(n30054), .Z(n30065) );
  XNOR U36226 ( .A(q[7]), .B(DB[922]), .Z(n30054) );
  IV U36227 ( .A(n30053), .Z(n36628) );
  XNOR U36228 ( .A(n30051), .B(n36629), .Z(n30053) );
  XNOR U36229 ( .A(q[6]), .B(DB[921]), .Z(n36629) );
  XNOR U36230 ( .A(q[5]), .B(DB[920]), .Z(n30051) );
  IV U36231 ( .A(n30064), .Z(n36626) );
  XOR U36232 ( .A(n36630), .B(n36631), .Z(n30064) );
  XNOR U36233 ( .A(n30060), .B(n30062), .Z(n36631) );
  XNOR U36234 ( .A(q[1]), .B(DB[916]), .Z(n30062) );
  XNOR U36235 ( .A(q[4]), .B(DB[919]), .Z(n30060) );
  IV U36236 ( .A(n30059), .Z(n36630) );
  XNOR U36237 ( .A(n30057), .B(n36632), .Z(n30059) );
  XNOR U36238 ( .A(q[3]), .B(DB[918]), .Z(n36632) );
  XNOR U36239 ( .A(q[2]), .B(DB[917]), .Z(n30057) );
  XOR U36240 ( .A(n36633), .B(n29955), .Z(n29883) );
  XOR U36241 ( .A(n36634), .B(n29947), .Z(n29955) );
  XOR U36242 ( .A(n36635), .B(n29936), .Z(n29947) );
  XNOR U36243 ( .A(q[14]), .B(DB[944]), .Z(n29936) );
  IV U36244 ( .A(n29935), .Z(n36635) );
  XNOR U36245 ( .A(n29933), .B(n36636), .Z(n29935) );
  XNOR U36246 ( .A(q[13]), .B(DB[943]), .Z(n36636) );
  XNOR U36247 ( .A(q[12]), .B(DB[942]), .Z(n29933) );
  IV U36248 ( .A(n29946), .Z(n36634) );
  XOR U36249 ( .A(n36637), .B(n36638), .Z(n29946) );
  XNOR U36250 ( .A(n29942), .B(n29944), .Z(n36638) );
  XNOR U36251 ( .A(q[8]), .B(DB[938]), .Z(n29944) );
  XNOR U36252 ( .A(q[11]), .B(DB[941]), .Z(n29942) );
  IV U36253 ( .A(n29941), .Z(n36637) );
  XNOR U36254 ( .A(n29939), .B(n36639), .Z(n29941) );
  XNOR U36255 ( .A(q[10]), .B(DB[940]), .Z(n36639) );
  XNOR U36256 ( .A(q[9]), .B(DB[939]), .Z(n29939) );
  IV U36257 ( .A(n29954), .Z(n36633) );
  XOR U36258 ( .A(n36640), .B(n36641), .Z(n29954) );
  XNOR U36259 ( .A(n29971), .B(n29952), .Z(n36641) );
  XNOR U36260 ( .A(q[0]), .B(DB[930]), .Z(n29952) );
  XOR U36261 ( .A(n36642), .B(n29960), .Z(n29971) );
  XNOR U36262 ( .A(q[7]), .B(DB[937]), .Z(n29960) );
  IV U36263 ( .A(n29959), .Z(n36642) );
  XNOR U36264 ( .A(n29957), .B(n36643), .Z(n29959) );
  XNOR U36265 ( .A(q[6]), .B(DB[936]), .Z(n36643) );
  XNOR U36266 ( .A(q[5]), .B(DB[935]), .Z(n29957) );
  IV U36267 ( .A(n29970), .Z(n36640) );
  XOR U36268 ( .A(n36644), .B(n36645), .Z(n29970) );
  XNOR U36269 ( .A(n29966), .B(n29968), .Z(n36645) );
  XNOR U36270 ( .A(q[1]), .B(DB[931]), .Z(n29968) );
  XNOR U36271 ( .A(q[4]), .B(DB[934]), .Z(n29966) );
  IV U36272 ( .A(n29965), .Z(n36644) );
  XNOR U36273 ( .A(n29963), .B(n36646), .Z(n29965) );
  XNOR U36274 ( .A(q[3]), .B(DB[933]), .Z(n36646) );
  XNOR U36275 ( .A(q[2]), .B(DB[932]), .Z(n29963) );
  XOR U36276 ( .A(n36647), .B(n29861), .Z(n29789) );
  XOR U36277 ( .A(n36648), .B(n29853), .Z(n29861) );
  XOR U36278 ( .A(n36649), .B(n29842), .Z(n29853) );
  XNOR U36279 ( .A(q[14]), .B(DB[959]), .Z(n29842) );
  IV U36280 ( .A(n29841), .Z(n36649) );
  XNOR U36281 ( .A(n29839), .B(n36650), .Z(n29841) );
  XNOR U36282 ( .A(q[13]), .B(DB[958]), .Z(n36650) );
  XNOR U36283 ( .A(q[12]), .B(DB[957]), .Z(n29839) );
  IV U36284 ( .A(n29852), .Z(n36648) );
  XOR U36285 ( .A(n36651), .B(n36652), .Z(n29852) );
  XNOR U36286 ( .A(n29848), .B(n29850), .Z(n36652) );
  XNOR U36287 ( .A(q[8]), .B(DB[953]), .Z(n29850) );
  XNOR U36288 ( .A(q[11]), .B(DB[956]), .Z(n29848) );
  IV U36289 ( .A(n29847), .Z(n36651) );
  XNOR U36290 ( .A(n29845), .B(n36653), .Z(n29847) );
  XNOR U36291 ( .A(q[10]), .B(DB[955]), .Z(n36653) );
  XNOR U36292 ( .A(q[9]), .B(DB[954]), .Z(n29845) );
  IV U36293 ( .A(n29860), .Z(n36647) );
  XOR U36294 ( .A(n36654), .B(n36655), .Z(n29860) );
  XNOR U36295 ( .A(n29877), .B(n29858), .Z(n36655) );
  XNOR U36296 ( .A(q[0]), .B(DB[945]), .Z(n29858) );
  XOR U36297 ( .A(n36656), .B(n29866), .Z(n29877) );
  XNOR U36298 ( .A(q[7]), .B(DB[952]), .Z(n29866) );
  IV U36299 ( .A(n29865), .Z(n36656) );
  XNOR U36300 ( .A(n29863), .B(n36657), .Z(n29865) );
  XNOR U36301 ( .A(q[6]), .B(DB[951]), .Z(n36657) );
  XNOR U36302 ( .A(q[5]), .B(DB[950]), .Z(n29863) );
  IV U36303 ( .A(n29876), .Z(n36654) );
  XOR U36304 ( .A(n36658), .B(n36659), .Z(n29876) );
  XNOR U36305 ( .A(n29872), .B(n29874), .Z(n36659) );
  XNOR U36306 ( .A(q[1]), .B(DB[946]), .Z(n29874) );
  XNOR U36307 ( .A(q[4]), .B(DB[949]), .Z(n29872) );
  IV U36308 ( .A(n29871), .Z(n36658) );
  XNOR U36309 ( .A(n29869), .B(n36660), .Z(n29871) );
  XNOR U36310 ( .A(q[3]), .B(DB[948]), .Z(n36660) );
  XNOR U36311 ( .A(q[2]), .B(DB[947]), .Z(n29869) );
  XOR U36312 ( .A(n36661), .B(n29767), .Z(n29695) );
  XOR U36313 ( .A(n36662), .B(n29759), .Z(n29767) );
  XOR U36314 ( .A(n36663), .B(n29748), .Z(n29759) );
  XNOR U36315 ( .A(q[14]), .B(DB[974]), .Z(n29748) );
  IV U36316 ( .A(n29747), .Z(n36663) );
  XNOR U36317 ( .A(n29745), .B(n36664), .Z(n29747) );
  XNOR U36318 ( .A(q[13]), .B(DB[973]), .Z(n36664) );
  XNOR U36319 ( .A(q[12]), .B(DB[972]), .Z(n29745) );
  IV U36320 ( .A(n29758), .Z(n36662) );
  XOR U36321 ( .A(n36665), .B(n36666), .Z(n29758) );
  XNOR U36322 ( .A(n29754), .B(n29756), .Z(n36666) );
  XNOR U36323 ( .A(q[8]), .B(DB[968]), .Z(n29756) );
  XNOR U36324 ( .A(q[11]), .B(DB[971]), .Z(n29754) );
  IV U36325 ( .A(n29753), .Z(n36665) );
  XNOR U36326 ( .A(n29751), .B(n36667), .Z(n29753) );
  XNOR U36327 ( .A(q[10]), .B(DB[970]), .Z(n36667) );
  XNOR U36328 ( .A(q[9]), .B(DB[969]), .Z(n29751) );
  IV U36329 ( .A(n29766), .Z(n36661) );
  XOR U36330 ( .A(n36668), .B(n36669), .Z(n29766) );
  XNOR U36331 ( .A(n29783), .B(n29764), .Z(n36669) );
  XNOR U36332 ( .A(q[0]), .B(DB[960]), .Z(n29764) );
  XOR U36333 ( .A(n36670), .B(n29772), .Z(n29783) );
  XNOR U36334 ( .A(q[7]), .B(DB[967]), .Z(n29772) );
  IV U36335 ( .A(n29771), .Z(n36670) );
  XNOR U36336 ( .A(n29769), .B(n36671), .Z(n29771) );
  XNOR U36337 ( .A(q[6]), .B(DB[966]), .Z(n36671) );
  XNOR U36338 ( .A(q[5]), .B(DB[965]), .Z(n29769) );
  IV U36339 ( .A(n29782), .Z(n36668) );
  XOR U36340 ( .A(n36672), .B(n36673), .Z(n29782) );
  XNOR U36341 ( .A(n29778), .B(n29780), .Z(n36673) );
  XNOR U36342 ( .A(q[1]), .B(DB[961]), .Z(n29780) );
  XNOR U36343 ( .A(q[4]), .B(DB[964]), .Z(n29778) );
  IV U36344 ( .A(n29777), .Z(n36672) );
  XNOR U36345 ( .A(n29775), .B(n36674), .Z(n29777) );
  XNOR U36346 ( .A(q[3]), .B(DB[963]), .Z(n36674) );
  XNOR U36347 ( .A(q[2]), .B(DB[962]), .Z(n29775) );
  XOR U36348 ( .A(n36675), .B(n29673), .Z(n29601) );
  XOR U36349 ( .A(n36676), .B(n29665), .Z(n29673) );
  XOR U36350 ( .A(n36677), .B(n29654), .Z(n29665) );
  XNOR U36351 ( .A(q[14]), .B(DB[989]), .Z(n29654) );
  IV U36352 ( .A(n29653), .Z(n36677) );
  XNOR U36353 ( .A(n29651), .B(n36678), .Z(n29653) );
  XNOR U36354 ( .A(q[13]), .B(DB[988]), .Z(n36678) );
  XNOR U36355 ( .A(q[12]), .B(DB[987]), .Z(n29651) );
  IV U36356 ( .A(n29664), .Z(n36676) );
  XOR U36357 ( .A(n36679), .B(n36680), .Z(n29664) );
  XNOR U36358 ( .A(n29660), .B(n29662), .Z(n36680) );
  XNOR U36359 ( .A(q[8]), .B(DB[983]), .Z(n29662) );
  XNOR U36360 ( .A(q[11]), .B(DB[986]), .Z(n29660) );
  IV U36361 ( .A(n29659), .Z(n36679) );
  XNOR U36362 ( .A(n29657), .B(n36681), .Z(n29659) );
  XNOR U36363 ( .A(q[10]), .B(DB[985]), .Z(n36681) );
  XNOR U36364 ( .A(q[9]), .B(DB[984]), .Z(n29657) );
  IV U36365 ( .A(n29672), .Z(n36675) );
  XOR U36366 ( .A(n36682), .B(n36683), .Z(n29672) );
  XNOR U36367 ( .A(n29689), .B(n29670), .Z(n36683) );
  XNOR U36368 ( .A(q[0]), .B(DB[975]), .Z(n29670) );
  XOR U36369 ( .A(n36684), .B(n29678), .Z(n29689) );
  XNOR U36370 ( .A(q[7]), .B(DB[982]), .Z(n29678) );
  IV U36371 ( .A(n29677), .Z(n36684) );
  XNOR U36372 ( .A(n29675), .B(n36685), .Z(n29677) );
  XNOR U36373 ( .A(q[6]), .B(DB[981]), .Z(n36685) );
  XNOR U36374 ( .A(q[5]), .B(DB[980]), .Z(n29675) );
  IV U36375 ( .A(n29688), .Z(n36682) );
  XOR U36376 ( .A(n36686), .B(n36687), .Z(n29688) );
  XNOR U36377 ( .A(n29684), .B(n29686), .Z(n36687) );
  XNOR U36378 ( .A(q[1]), .B(DB[976]), .Z(n29686) );
  XNOR U36379 ( .A(q[4]), .B(DB[979]), .Z(n29684) );
  IV U36380 ( .A(n29683), .Z(n36686) );
  XNOR U36381 ( .A(n29681), .B(n36688), .Z(n29683) );
  XNOR U36382 ( .A(q[3]), .B(DB[978]), .Z(n36688) );
  XNOR U36383 ( .A(q[2]), .B(DB[977]), .Z(n29681) );
  XOR U36384 ( .A(n36689), .B(n29579), .Z(n29507) );
  XOR U36385 ( .A(n36690), .B(n29571), .Z(n29579) );
  XOR U36386 ( .A(n36691), .B(n29560), .Z(n29571) );
  XNOR U36387 ( .A(q[14]), .B(DB[1004]), .Z(n29560) );
  IV U36388 ( .A(n29559), .Z(n36691) );
  XNOR U36389 ( .A(n29557), .B(n36692), .Z(n29559) );
  XNOR U36390 ( .A(q[13]), .B(DB[1003]), .Z(n36692) );
  XNOR U36391 ( .A(q[12]), .B(DB[1002]), .Z(n29557) );
  IV U36392 ( .A(n29570), .Z(n36690) );
  XOR U36393 ( .A(n36693), .B(n36694), .Z(n29570) );
  XNOR U36394 ( .A(n29566), .B(n29568), .Z(n36694) );
  XNOR U36395 ( .A(q[8]), .B(DB[998]), .Z(n29568) );
  XNOR U36396 ( .A(q[11]), .B(DB[1001]), .Z(n29566) );
  IV U36397 ( .A(n29565), .Z(n36693) );
  XNOR U36398 ( .A(n29563), .B(n36695), .Z(n29565) );
  XNOR U36399 ( .A(q[10]), .B(DB[1000]), .Z(n36695) );
  XNOR U36400 ( .A(q[9]), .B(DB[999]), .Z(n29563) );
  IV U36401 ( .A(n29578), .Z(n36689) );
  XOR U36402 ( .A(n36696), .B(n36697), .Z(n29578) );
  XNOR U36403 ( .A(n29595), .B(n29576), .Z(n36697) );
  XNOR U36404 ( .A(q[0]), .B(DB[990]), .Z(n29576) );
  XOR U36405 ( .A(n36698), .B(n29584), .Z(n29595) );
  XNOR U36406 ( .A(q[7]), .B(DB[997]), .Z(n29584) );
  IV U36407 ( .A(n29583), .Z(n36698) );
  XNOR U36408 ( .A(n29581), .B(n36699), .Z(n29583) );
  XNOR U36409 ( .A(q[6]), .B(DB[996]), .Z(n36699) );
  XNOR U36410 ( .A(q[5]), .B(DB[995]), .Z(n29581) );
  IV U36411 ( .A(n29594), .Z(n36696) );
  XOR U36412 ( .A(n36700), .B(n36701), .Z(n29594) );
  XNOR U36413 ( .A(n29590), .B(n29592), .Z(n36701) );
  XNOR U36414 ( .A(q[1]), .B(DB[991]), .Z(n29592) );
  XNOR U36415 ( .A(q[4]), .B(DB[994]), .Z(n29590) );
  IV U36416 ( .A(n29589), .Z(n36700) );
  XNOR U36417 ( .A(n29587), .B(n36702), .Z(n29589) );
  XNOR U36418 ( .A(q[3]), .B(DB[993]), .Z(n36702) );
  XNOR U36419 ( .A(q[2]), .B(DB[992]), .Z(n29587) );
  XOR U36420 ( .A(n36703), .B(n29485), .Z(n29413) );
  XOR U36421 ( .A(n36704), .B(n29477), .Z(n29485) );
  XOR U36422 ( .A(n36705), .B(n29466), .Z(n29477) );
  XNOR U36423 ( .A(q[14]), .B(DB[1019]), .Z(n29466) );
  IV U36424 ( .A(n29465), .Z(n36705) );
  XNOR U36425 ( .A(n29463), .B(n36706), .Z(n29465) );
  XNOR U36426 ( .A(q[13]), .B(DB[1018]), .Z(n36706) );
  XNOR U36427 ( .A(q[12]), .B(DB[1017]), .Z(n29463) );
  IV U36428 ( .A(n29476), .Z(n36704) );
  XOR U36429 ( .A(n36707), .B(n36708), .Z(n29476) );
  XNOR U36430 ( .A(n29472), .B(n29474), .Z(n36708) );
  XNOR U36431 ( .A(q[8]), .B(DB[1013]), .Z(n29474) );
  XNOR U36432 ( .A(q[11]), .B(DB[1016]), .Z(n29472) );
  IV U36433 ( .A(n29471), .Z(n36707) );
  XNOR U36434 ( .A(n29469), .B(n36709), .Z(n29471) );
  XNOR U36435 ( .A(q[10]), .B(DB[1015]), .Z(n36709) );
  XNOR U36436 ( .A(q[9]), .B(DB[1014]), .Z(n29469) );
  IV U36437 ( .A(n29484), .Z(n36703) );
  XOR U36438 ( .A(n36710), .B(n36711), .Z(n29484) );
  XNOR U36439 ( .A(n29501), .B(n29482), .Z(n36711) );
  XNOR U36440 ( .A(q[0]), .B(DB[1005]), .Z(n29482) );
  XOR U36441 ( .A(n36712), .B(n29490), .Z(n29501) );
  XNOR U36442 ( .A(q[7]), .B(DB[1012]), .Z(n29490) );
  IV U36443 ( .A(n29489), .Z(n36712) );
  XNOR U36444 ( .A(n29487), .B(n36713), .Z(n29489) );
  XNOR U36445 ( .A(q[6]), .B(DB[1011]), .Z(n36713) );
  XNOR U36446 ( .A(q[5]), .B(DB[1010]), .Z(n29487) );
  IV U36447 ( .A(n29500), .Z(n36710) );
  XOR U36448 ( .A(n36714), .B(n36715), .Z(n29500) );
  XNOR U36449 ( .A(n29496), .B(n29498), .Z(n36715) );
  XNOR U36450 ( .A(q[1]), .B(DB[1006]), .Z(n29498) );
  XNOR U36451 ( .A(q[4]), .B(DB[1009]), .Z(n29496) );
  IV U36452 ( .A(n29495), .Z(n36714) );
  XNOR U36453 ( .A(n29493), .B(n36716), .Z(n29495) );
  XNOR U36454 ( .A(q[3]), .B(DB[1008]), .Z(n36716) );
  XNOR U36455 ( .A(q[2]), .B(DB[1007]), .Z(n29493) );
  XOR U36456 ( .A(n36717), .B(n29391), .Z(n29319) );
  XOR U36457 ( .A(n36718), .B(n29383), .Z(n29391) );
  XOR U36458 ( .A(n36719), .B(n29372), .Z(n29383) );
  XNOR U36459 ( .A(q[14]), .B(DB[1034]), .Z(n29372) );
  IV U36460 ( .A(n29371), .Z(n36719) );
  XNOR U36461 ( .A(n29369), .B(n36720), .Z(n29371) );
  XNOR U36462 ( .A(q[13]), .B(DB[1033]), .Z(n36720) );
  XNOR U36463 ( .A(q[12]), .B(DB[1032]), .Z(n29369) );
  IV U36464 ( .A(n29382), .Z(n36718) );
  XOR U36465 ( .A(n36721), .B(n36722), .Z(n29382) );
  XNOR U36466 ( .A(n29378), .B(n29380), .Z(n36722) );
  XNOR U36467 ( .A(q[8]), .B(DB[1028]), .Z(n29380) );
  XNOR U36468 ( .A(q[11]), .B(DB[1031]), .Z(n29378) );
  IV U36469 ( .A(n29377), .Z(n36721) );
  XNOR U36470 ( .A(n29375), .B(n36723), .Z(n29377) );
  XNOR U36471 ( .A(q[10]), .B(DB[1030]), .Z(n36723) );
  XNOR U36472 ( .A(q[9]), .B(DB[1029]), .Z(n29375) );
  IV U36473 ( .A(n29390), .Z(n36717) );
  XOR U36474 ( .A(n36724), .B(n36725), .Z(n29390) );
  XNOR U36475 ( .A(n29407), .B(n29388), .Z(n36725) );
  XNOR U36476 ( .A(q[0]), .B(DB[1020]), .Z(n29388) );
  XOR U36477 ( .A(n36726), .B(n29396), .Z(n29407) );
  XNOR U36478 ( .A(q[7]), .B(DB[1027]), .Z(n29396) );
  IV U36479 ( .A(n29395), .Z(n36726) );
  XNOR U36480 ( .A(n29393), .B(n36727), .Z(n29395) );
  XNOR U36481 ( .A(q[6]), .B(DB[1026]), .Z(n36727) );
  XNOR U36482 ( .A(q[5]), .B(DB[1025]), .Z(n29393) );
  IV U36483 ( .A(n29406), .Z(n36724) );
  XOR U36484 ( .A(n36728), .B(n36729), .Z(n29406) );
  XNOR U36485 ( .A(n29402), .B(n29404), .Z(n36729) );
  XNOR U36486 ( .A(q[1]), .B(DB[1021]), .Z(n29404) );
  XNOR U36487 ( .A(q[4]), .B(DB[1024]), .Z(n29402) );
  IV U36488 ( .A(n29401), .Z(n36728) );
  XNOR U36489 ( .A(n29399), .B(n36730), .Z(n29401) );
  XNOR U36490 ( .A(q[3]), .B(DB[1023]), .Z(n36730) );
  XNOR U36491 ( .A(q[2]), .B(DB[1022]), .Z(n29399) );
  XOR U36492 ( .A(n36731), .B(n29297), .Z(n29225) );
  XOR U36493 ( .A(n36732), .B(n29289), .Z(n29297) );
  XOR U36494 ( .A(n36733), .B(n29278), .Z(n29289) );
  XNOR U36495 ( .A(q[14]), .B(DB[1049]), .Z(n29278) );
  IV U36496 ( .A(n29277), .Z(n36733) );
  XNOR U36497 ( .A(n29275), .B(n36734), .Z(n29277) );
  XNOR U36498 ( .A(q[13]), .B(DB[1048]), .Z(n36734) );
  XNOR U36499 ( .A(q[12]), .B(DB[1047]), .Z(n29275) );
  IV U36500 ( .A(n29288), .Z(n36732) );
  XOR U36501 ( .A(n36735), .B(n36736), .Z(n29288) );
  XNOR U36502 ( .A(n29284), .B(n29286), .Z(n36736) );
  XNOR U36503 ( .A(q[8]), .B(DB[1043]), .Z(n29286) );
  XNOR U36504 ( .A(q[11]), .B(DB[1046]), .Z(n29284) );
  IV U36505 ( .A(n29283), .Z(n36735) );
  XNOR U36506 ( .A(n29281), .B(n36737), .Z(n29283) );
  XNOR U36507 ( .A(q[10]), .B(DB[1045]), .Z(n36737) );
  XNOR U36508 ( .A(q[9]), .B(DB[1044]), .Z(n29281) );
  IV U36509 ( .A(n29296), .Z(n36731) );
  XOR U36510 ( .A(n36738), .B(n36739), .Z(n29296) );
  XNOR U36511 ( .A(n29313), .B(n29294), .Z(n36739) );
  XNOR U36512 ( .A(q[0]), .B(DB[1035]), .Z(n29294) );
  XOR U36513 ( .A(n36740), .B(n29302), .Z(n29313) );
  XNOR U36514 ( .A(q[7]), .B(DB[1042]), .Z(n29302) );
  IV U36515 ( .A(n29301), .Z(n36740) );
  XNOR U36516 ( .A(n29299), .B(n36741), .Z(n29301) );
  XNOR U36517 ( .A(q[6]), .B(DB[1041]), .Z(n36741) );
  XNOR U36518 ( .A(q[5]), .B(DB[1040]), .Z(n29299) );
  IV U36519 ( .A(n29312), .Z(n36738) );
  XOR U36520 ( .A(n36742), .B(n36743), .Z(n29312) );
  XNOR U36521 ( .A(n29308), .B(n29310), .Z(n36743) );
  XNOR U36522 ( .A(q[1]), .B(DB[1036]), .Z(n29310) );
  XNOR U36523 ( .A(q[4]), .B(DB[1039]), .Z(n29308) );
  IV U36524 ( .A(n29307), .Z(n36742) );
  XNOR U36525 ( .A(n29305), .B(n36744), .Z(n29307) );
  XNOR U36526 ( .A(q[3]), .B(DB[1038]), .Z(n36744) );
  XNOR U36527 ( .A(q[2]), .B(DB[1037]), .Z(n29305) );
  XOR U36528 ( .A(n36745), .B(n29203), .Z(n29131) );
  XOR U36529 ( .A(n36746), .B(n29195), .Z(n29203) );
  XOR U36530 ( .A(n36747), .B(n29184), .Z(n29195) );
  XNOR U36531 ( .A(q[14]), .B(DB[1064]), .Z(n29184) );
  IV U36532 ( .A(n29183), .Z(n36747) );
  XNOR U36533 ( .A(n29181), .B(n36748), .Z(n29183) );
  XNOR U36534 ( .A(q[13]), .B(DB[1063]), .Z(n36748) );
  XNOR U36535 ( .A(q[12]), .B(DB[1062]), .Z(n29181) );
  IV U36536 ( .A(n29194), .Z(n36746) );
  XOR U36537 ( .A(n36749), .B(n36750), .Z(n29194) );
  XNOR U36538 ( .A(n29190), .B(n29192), .Z(n36750) );
  XNOR U36539 ( .A(q[8]), .B(DB[1058]), .Z(n29192) );
  XNOR U36540 ( .A(q[11]), .B(DB[1061]), .Z(n29190) );
  IV U36541 ( .A(n29189), .Z(n36749) );
  XNOR U36542 ( .A(n29187), .B(n36751), .Z(n29189) );
  XNOR U36543 ( .A(q[10]), .B(DB[1060]), .Z(n36751) );
  XNOR U36544 ( .A(q[9]), .B(DB[1059]), .Z(n29187) );
  IV U36545 ( .A(n29202), .Z(n36745) );
  XOR U36546 ( .A(n36752), .B(n36753), .Z(n29202) );
  XNOR U36547 ( .A(n29219), .B(n29200), .Z(n36753) );
  XNOR U36548 ( .A(q[0]), .B(DB[1050]), .Z(n29200) );
  XOR U36549 ( .A(n36754), .B(n29208), .Z(n29219) );
  XNOR U36550 ( .A(q[7]), .B(DB[1057]), .Z(n29208) );
  IV U36551 ( .A(n29207), .Z(n36754) );
  XNOR U36552 ( .A(n29205), .B(n36755), .Z(n29207) );
  XNOR U36553 ( .A(q[6]), .B(DB[1056]), .Z(n36755) );
  XNOR U36554 ( .A(q[5]), .B(DB[1055]), .Z(n29205) );
  IV U36555 ( .A(n29218), .Z(n36752) );
  XOR U36556 ( .A(n36756), .B(n36757), .Z(n29218) );
  XNOR U36557 ( .A(n29214), .B(n29216), .Z(n36757) );
  XNOR U36558 ( .A(q[1]), .B(DB[1051]), .Z(n29216) );
  XNOR U36559 ( .A(q[4]), .B(DB[1054]), .Z(n29214) );
  IV U36560 ( .A(n29213), .Z(n36756) );
  XNOR U36561 ( .A(n29211), .B(n36758), .Z(n29213) );
  XNOR U36562 ( .A(q[3]), .B(DB[1053]), .Z(n36758) );
  XNOR U36563 ( .A(q[2]), .B(DB[1052]), .Z(n29211) );
  XOR U36564 ( .A(n36759), .B(n29109), .Z(n29037) );
  XOR U36565 ( .A(n36760), .B(n29101), .Z(n29109) );
  XOR U36566 ( .A(n36761), .B(n29090), .Z(n29101) );
  XNOR U36567 ( .A(q[14]), .B(DB[1079]), .Z(n29090) );
  IV U36568 ( .A(n29089), .Z(n36761) );
  XNOR U36569 ( .A(n29087), .B(n36762), .Z(n29089) );
  XNOR U36570 ( .A(q[13]), .B(DB[1078]), .Z(n36762) );
  XNOR U36571 ( .A(q[12]), .B(DB[1077]), .Z(n29087) );
  IV U36572 ( .A(n29100), .Z(n36760) );
  XOR U36573 ( .A(n36763), .B(n36764), .Z(n29100) );
  XNOR U36574 ( .A(n29096), .B(n29098), .Z(n36764) );
  XNOR U36575 ( .A(q[8]), .B(DB[1073]), .Z(n29098) );
  XNOR U36576 ( .A(q[11]), .B(DB[1076]), .Z(n29096) );
  IV U36577 ( .A(n29095), .Z(n36763) );
  XNOR U36578 ( .A(n29093), .B(n36765), .Z(n29095) );
  XNOR U36579 ( .A(q[10]), .B(DB[1075]), .Z(n36765) );
  XNOR U36580 ( .A(q[9]), .B(DB[1074]), .Z(n29093) );
  IV U36581 ( .A(n29108), .Z(n36759) );
  XOR U36582 ( .A(n36766), .B(n36767), .Z(n29108) );
  XNOR U36583 ( .A(n29125), .B(n29106), .Z(n36767) );
  XNOR U36584 ( .A(q[0]), .B(DB[1065]), .Z(n29106) );
  XOR U36585 ( .A(n36768), .B(n29114), .Z(n29125) );
  XNOR U36586 ( .A(q[7]), .B(DB[1072]), .Z(n29114) );
  IV U36587 ( .A(n29113), .Z(n36768) );
  XNOR U36588 ( .A(n29111), .B(n36769), .Z(n29113) );
  XNOR U36589 ( .A(q[6]), .B(DB[1071]), .Z(n36769) );
  XNOR U36590 ( .A(q[5]), .B(DB[1070]), .Z(n29111) );
  IV U36591 ( .A(n29124), .Z(n36766) );
  XOR U36592 ( .A(n36770), .B(n36771), .Z(n29124) );
  XNOR U36593 ( .A(n29120), .B(n29122), .Z(n36771) );
  XNOR U36594 ( .A(q[1]), .B(DB[1066]), .Z(n29122) );
  XNOR U36595 ( .A(q[4]), .B(DB[1069]), .Z(n29120) );
  IV U36596 ( .A(n29119), .Z(n36770) );
  XNOR U36597 ( .A(n29117), .B(n36772), .Z(n29119) );
  XNOR U36598 ( .A(q[3]), .B(DB[1068]), .Z(n36772) );
  XNOR U36599 ( .A(q[2]), .B(DB[1067]), .Z(n29117) );
  XOR U36600 ( .A(n36773), .B(n29015), .Z(n28943) );
  XOR U36601 ( .A(n36774), .B(n29007), .Z(n29015) );
  XOR U36602 ( .A(n36775), .B(n28996), .Z(n29007) );
  XNOR U36603 ( .A(q[14]), .B(DB[1094]), .Z(n28996) );
  IV U36604 ( .A(n28995), .Z(n36775) );
  XNOR U36605 ( .A(n28993), .B(n36776), .Z(n28995) );
  XNOR U36606 ( .A(q[13]), .B(DB[1093]), .Z(n36776) );
  XNOR U36607 ( .A(q[12]), .B(DB[1092]), .Z(n28993) );
  IV U36608 ( .A(n29006), .Z(n36774) );
  XOR U36609 ( .A(n36777), .B(n36778), .Z(n29006) );
  XNOR U36610 ( .A(n29002), .B(n29004), .Z(n36778) );
  XNOR U36611 ( .A(q[8]), .B(DB[1088]), .Z(n29004) );
  XNOR U36612 ( .A(q[11]), .B(DB[1091]), .Z(n29002) );
  IV U36613 ( .A(n29001), .Z(n36777) );
  XNOR U36614 ( .A(n28999), .B(n36779), .Z(n29001) );
  XNOR U36615 ( .A(q[10]), .B(DB[1090]), .Z(n36779) );
  XNOR U36616 ( .A(q[9]), .B(DB[1089]), .Z(n28999) );
  IV U36617 ( .A(n29014), .Z(n36773) );
  XOR U36618 ( .A(n36780), .B(n36781), .Z(n29014) );
  XNOR U36619 ( .A(n29031), .B(n29012), .Z(n36781) );
  XNOR U36620 ( .A(q[0]), .B(DB[1080]), .Z(n29012) );
  XOR U36621 ( .A(n36782), .B(n29020), .Z(n29031) );
  XNOR U36622 ( .A(q[7]), .B(DB[1087]), .Z(n29020) );
  IV U36623 ( .A(n29019), .Z(n36782) );
  XNOR U36624 ( .A(n29017), .B(n36783), .Z(n29019) );
  XNOR U36625 ( .A(q[6]), .B(DB[1086]), .Z(n36783) );
  XNOR U36626 ( .A(q[5]), .B(DB[1085]), .Z(n29017) );
  IV U36627 ( .A(n29030), .Z(n36780) );
  XOR U36628 ( .A(n36784), .B(n36785), .Z(n29030) );
  XNOR U36629 ( .A(n29026), .B(n29028), .Z(n36785) );
  XNOR U36630 ( .A(q[1]), .B(DB[1081]), .Z(n29028) );
  XNOR U36631 ( .A(q[4]), .B(DB[1084]), .Z(n29026) );
  IV U36632 ( .A(n29025), .Z(n36784) );
  XNOR U36633 ( .A(n29023), .B(n36786), .Z(n29025) );
  XNOR U36634 ( .A(q[3]), .B(DB[1083]), .Z(n36786) );
  XNOR U36635 ( .A(q[2]), .B(DB[1082]), .Z(n29023) );
  XOR U36636 ( .A(n36787), .B(n28921), .Z(n28849) );
  XOR U36637 ( .A(n36788), .B(n28913), .Z(n28921) );
  XOR U36638 ( .A(n36789), .B(n28902), .Z(n28913) );
  XNOR U36639 ( .A(q[14]), .B(DB[1109]), .Z(n28902) );
  IV U36640 ( .A(n28901), .Z(n36789) );
  XNOR U36641 ( .A(n28899), .B(n36790), .Z(n28901) );
  XNOR U36642 ( .A(q[13]), .B(DB[1108]), .Z(n36790) );
  XNOR U36643 ( .A(q[12]), .B(DB[1107]), .Z(n28899) );
  IV U36644 ( .A(n28912), .Z(n36788) );
  XOR U36645 ( .A(n36791), .B(n36792), .Z(n28912) );
  XNOR U36646 ( .A(n28908), .B(n28910), .Z(n36792) );
  XNOR U36647 ( .A(q[8]), .B(DB[1103]), .Z(n28910) );
  XNOR U36648 ( .A(q[11]), .B(DB[1106]), .Z(n28908) );
  IV U36649 ( .A(n28907), .Z(n36791) );
  XNOR U36650 ( .A(n28905), .B(n36793), .Z(n28907) );
  XNOR U36651 ( .A(q[10]), .B(DB[1105]), .Z(n36793) );
  XNOR U36652 ( .A(q[9]), .B(DB[1104]), .Z(n28905) );
  IV U36653 ( .A(n28920), .Z(n36787) );
  XOR U36654 ( .A(n36794), .B(n36795), .Z(n28920) );
  XNOR U36655 ( .A(n28937), .B(n28918), .Z(n36795) );
  XNOR U36656 ( .A(q[0]), .B(DB[1095]), .Z(n28918) );
  XOR U36657 ( .A(n36796), .B(n28926), .Z(n28937) );
  XNOR U36658 ( .A(q[7]), .B(DB[1102]), .Z(n28926) );
  IV U36659 ( .A(n28925), .Z(n36796) );
  XNOR U36660 ( .A(n28923), .B(n36797), .Z(n28925) );
  XNOR U36661 ( .A(q[6]), .B(DB[1101]), .Z(n36797) );
  XNOR U36662 ( .A(q[5]), .B(DB[1100]), .Z(n28923) );
  IV U36663 ( .A(n28936), .Z(n36794) );
  XOR U36664 ( .A(n36798), .B(n36799), .Z(n28936) );
  XNOR U36665 ( .A(n28932), .B(n28934), .Z(n36799) );
  XNOR U36666 ( .A(q[1]), .B(DB[1096]), .Z(n28934) );
  XNOR U36667 ( .A(q[4]), .B(DB[1099]), .Z(n28932) );
  IV U36668 ( .A(n28931), .Z(n36798) );
  XNOR U36669 ( .A(n28929), .B(n36800), .Z(n28931) );
  XNOR U36670 ( .A(q[3]), .B(DB[1098]), .Z(n36800) );
  XNOR U36671 ( .A(q[2]), .B(DB[1097]), .Z(n28929) );
  XOR U36672 ( .A(n36801), .B(n28827), .Z(n28755) );
  XOR U36673 ( .A(n36802), .B(n28819), .Z(n28827) );
  XOR U36674 ( .A(n36803), .B(n28808), .Z(n28819) );
  XNOR U36675 ( .A(q[14]), .B(DB[1124]), .Z(n28808) );
  IV U36676 ( .A(n28807), .Z(n36803) );
  XNOR U36677 ( .A(n28805), .B(n36804), .Z(n28807) );
  XNOR U36678 ( .A(q[13]), .B(DB[1123]), .Z(n36804) );
  XNOR U36679 ( .A(q[12]), .B(DB[1122]), .Z(n28805) );
  IV U36680 ( .A(n28818), .Z(n36802) );
  XOR U36681 ( .A(n36805), .B(n36806), .Z(n28818) );
  XNOR U36682 ( .A(n28814), .B(n28816), .Z(n36806) );
  XNOR U36683 ( .A(q[8]), .B(DB[1118]), .Z(n28816) );
  XNOR U36684 ( .A(q[11]), .B(DB[1121]), .Z(n28814) );
  IV U36685 ( .A(n28813), .Z(n36805) );
  XNOR U36686 ( .A(n28811), .B(n36807), .Z(n28813) );
  XNOR U36687 ( .A(q[10]), .B(DB[1120]), .Z(n36807) );
  XNOR U36688 ( .A(q[9]), .B(DB[1119]), .Z(n28811) );
  IV U36689 ( .A(n28826), .Z(n36801) );
  XOR U36690 ( .A(n36808), .B(n36809), .Z(n28826) );
  XNOR U36691 ( .A(n28843), .B(n28824), .Z(n36809) );
  XNOR U36692 ( .A(q[0]), .B(DB[1110]), .Z(n28824) );
  XOR U36693 ( .A(n36810), .B(n28832), .Z(n28843) );
  XNOR U36694 ( .A(q[7]), .B(DB[1117]), .Z(n28832) );
  IV U36695 ( .A(n28831), .Z(n36810) );
  XNOR U36696 ( .A(n28829), .B(n36811), .Z(n28831) );
  XNOR U36697 ( .A(q[6]), .B(DB[1116]), .Z(n36811) );
  XNOR U36698 ( .A(q[5]), .B(DB[1115]), .Z(n28829) );
  IV U36699 ( .A(n28842), .Z(n36808) );
  XOR U36700 ( .A(n36812), .B(n36813), .Z(n28842) );
  XNOR U36701 ( .A(n28838), .B(n28840), .Z(n36813) );
  XNOR U36702 ( .A(q[1]), .B(DB[1111]), .Z(n28840) );
  XNOR U36703 ( .A(q[4]), .B(DB[1114]), .Z(n28838) );
  IV U36704 ( .A(n28837), .Z(n36812) );
  XNOR U36705 ( .A(n28835), .B(n36814), .Z(n28837) );
  XNOR U36706 ( .A(q[3]), .B(DB[1113]), .Z(n36814) );
  XNOR U36707 ( .A(q[2]), .B(DB[1112]), .Z(n28835) );
  XOR U36708 ( .A(n36815), .B(n28733), .Z(n28661) );
  XOR U36709 ( .A(n36816), .B(n28725), .Z(n28733) );
  XOR U36710 ( .A(n36817), .B(n28714), .Z(n28725) );
  XNOR U36711 ( .A(q[14]), .B(DB[1139]), .Z(n28714) );
  IV U36712 ( .A(n28713), .Z(n36817) );
  XNOR U36713 ( .A(n28711), .B(n36818), .Z(n28713) );
  XNOR U36714 ( .A(q[13]), .B(DB[1138]), .Z(n36818) );
  XNOR U36715 ( .A(q[12]), .B(DB[1137]), .Z(n28711) );
  IV U36716 ( .A(n28724), .Z(n36816) );
  XOR U36717 ( .A(n36819), .B(n36820), .Z(n28724) );
  XNOR U36718 ( .A(n28720), .B(n28722), .Z(n36820) );
  XNOR U36719 ( .A(q[8]), .B(DB[1133]), .Z(n28722) );
  XNOR U36720 ( .A(q[11]), .B(DB[1136]), .Z(n28720) );
  IV U36721 ( .A(n28719), .Z(n36819) );
  XNOR U36722 ( .A(n28717), .B(n36821), .Z(n28719) );
  XNOR U36723 ( .A(q[10]), .B(DB[1135]), .Z(n36821) );
  XNOR U36724 ( .A(q[9]), .B(DB[1134]), .Z(n28717) );
  IV U36725 ( .A(n28732), .Z(n36815) );
  XOR U36726 ( .A(n36822), .B(n36823), .Z(n28732) );
  XNOR U36727 ( .A(n28749), .B(n28730), .Z(n36823) );
  XNOR U36728 ( .A(q[0]), .B(DB[1125]), .Z(n28730) );
  XOR U36729 ( .A(n36824), .B(n28738), .Z(n28749) );
  XNOR U36730 ( .A(q[7]), .B(DB[1132]), .Z(n28738) );
  IV U36731 ( .A(n28737), .Z(n36824) );
  XNOR U36732 ( .A(n28735), .B(n36825), .Z(n28737) );
  XNOR U36733 ( .A(q[6]), .B(DB[1131]), .Z(n36825) );
  XNOR U36734 ( .A(q[5]), .B(DB[1130]), .Z(n28735) );
  IV U36735 ( .A(n28748), .Z(n36822) );
  XOR U36736 ( .A(n36826), .B(n36827), .Z(n28748) );
  XNOR U36737 ( .A(n28744), .B(n28746), .Z(n36827) );
  XNOR U36738 ( .A(q[1]), .B(DB[1126]), .Z(n28746) );
  XNOR U36739 ( .A(q[4]), .B(DB[1129]), .Z(n28744) );
  IV U36740 ( .A(n28743), .Z(n36826) );
  XNOR U36741 ( .A(n28741), .B(n36828), .Z(n28743) );
  XNOR U36742 ( .A(q[3]), .B(DB[1128]), .Z(n36828) );
  XNOR U36743 ( .A(q[2]), .B(DB[1127]), .Z(n28741) );
  XOR U36744 ( .A(n36829), .B(n28639), .Z(n28567) );
  XOR U36745 ( .A(n36830), .B(n28631), .Z(n28639) );
  XOR U36746 ( .A(n36831), .B(n28620), .Z(n28631) );
  XNOR U36747 ( .A(q[14]), .B(DB[1154]), .Z(n28620) );
  IV U36748 ( .A(n28619), .Z(n36831) );
  XNOR U36749 ( .A(n28617), .B(n36832), .Z(n28619) );
  XNOR U36750 ( .A(q[13]), .B(DB[1153]), .Z(n36832) );
  XNOR U36751 ( .A(q[12]), .B(DB[1152]), .Z(n28617) );
  IV U36752 ( .A(n28630), .Z(n36830) );
  XOR U36753 ( .A(n36833), .B(n36834), .Z(n28630) );
  XNOR U36754 ( .A(n28626), .B(n28628), .Z(n36834) );
  XNOR U36755 ( .A(q[8]), .B(DB[1148]), .Z(n28628) );
  XNOR U36756 ( .A(q[11]), .B(DB[1151]), .Z(n28626) );
  IV U36757 ( .A(n28625), .Z(n36833) );
  XNOR U36758 ( .A(n28623), .B(n36835), .Z(n28625) );
  XNOR U36759 ( .A(q[10]), .B(DB[1150]), .Z(n36835) );
  XNOR U36760 ( .A(q[9]), .B(DB[1149]), .Z(n28623) );
  IV U36761 ( .A(n28638), .Z(n36829) );
  XOR U36762 ( .A(n36836), .B(n36837), .Z(n28638) );
  XNOR U36763 ( .A(n28655), .B(n28636), .Z(n36837) );
  XNOR U36764 ( .A(q[0]), .B(DB[1140]), .Z(n28636) );
  XOR U36765 ( .A(n36838), .B(n28644), .Z(n28655) );
  XNOR U36766 ( .A(q[7]), .B(DB[1147]), .Z(n28644) );
  IV U36767 ( .A(n28643), .Z(n36838) );
  XNOR U36768 ( .A(n28641), .B(n36839), .Z(n28643) );
  XNOR U36769 ( .A(q[6]), .B(DB[1146]), .Z(n36839) );
  XNOR U36770 ( .A(q[5]), .B(DB[1145]), .Z(n28641) );
  IV U36771 ( .A(n28654), .Z(n36836) );
  XOR U36772 ( .A(n36840), .B(n36841), .Z(n28654) );
  XNOR U36773 ( .A(n28650), .B(n28652), .Z(n36841) );
  XNOR U36774 ( .A(q[1]), .B(DB[1141]), .Z(n28652) );
  XNOR U36775 ( .A(q[4]), .B(DB[1144]), .Z(n28650) );
  IV U36776 ( .A(n28649), .Z(n36840) );
  XNOR U36777 ( .A(n28647), .B(n36842), .Z(n28649) );
  XNOR U36778 ( .A(q[3]), .B(DB[1143]), .Z(n36842) );
  XNOR U36779 ( .A(q[2]), .B(DB[1142]), .Z(n28647) );
  XOR U36780 ( .A(n36843), .B(n28545), .Z(n28473) );
  XOR U36781 ( .A(n36844), .B(n28537), .Z(n28545) );
  XOR U36782 ( .A(n36845), .B(n28526), .Z(n28537) );
  XNOR U36783 ( .A(q[14]), .B(DB[1169]), .Z(n28526) );
  IV U36784 ( .A(n28525), .Z(n36845) );
  XNOR U36785 ( .A(n28523), .B(n36846), .Z(n28525) );
  XNOR U36786 ( .A(q[13]), .B(DB[1168]), .Z(n36846) );
  XNOR U36787 ( .A(q[12]), .B(DB[1167]), .Z(n28523) );
  IV U36788 ( .A(n28536), .Z(n36844) );
  XOR U36789 ( .A(n36847), .B(n36848), .Z(n28536) );
  XNOR U36790 ( .A(n28532), .B(n28534), .Z(n36848) );
  XNOR U36791 ( .A(q[8]), .B(DB[1163]), .Z(n28534) );
  XNOR U36792 ( .A(q[11]), .B(DB[1166]), .Z(n28532) );
  IV U36793 ( .A(n28531), .Z(n36847) );
  XNOR U36794 ( .A(n28529), .B(n36849), .Z(n28531) );
  XNOR U36795 ( .A(q[10]), .B(DB[1165]), .Z(n36849) );
  XNOR U36796 ( .A(q[9]), .B(DB[1164]), .Z(n28529) );
  IV U36797 ( .A(n28544), .Z(n36843) );
  XOR U36798 ( .A(n36850), .B(n36851), .Z(n28544) );
  XNOR U36799 ( .A(n28561), .B(n28542), .Z(n36851) );
  XNOR U36800 ( .A(q[0]), .B(DB[1155]), .Z(n28542) );
  XOR U36801 ( .A(n36852), .B(n28550), .Z(n28561) );
  XNOR U36802 ( .A(q[7]), .B(DB[1162]), .Z(n28550) );
  IV U36803 ( .A(n28549), .Z(n36852) );
  XNOR U36804 ( .A(n28547), .B(n36853), .Z(n28549) );
  XNOR U36805 ( .A(q[6]), .B(DB[1161]), .Z(n36853) );
  XNOR U36806 ( .A(q[5]), .B(DB[1160]), .Z(n28547) );
  IV U36807 ( .A(n28560), .Z(n36850) );
  XOR U36808 ( .A(n36854), .B(n36855), .Z(n28560) );
  XNOR U36809 ( .A(n28556), .B(n28558), .Z(n36855) );
  XNOR U36810 ( .A(q[1]), .B(DB[1156]), .Z(n28558) );
  XNOR U36811 ( .A(q[4]), .B(DB[1159]), .Z(n28556) );
  IV U36812 ( .A(n28555), .Z(n36854) );
  XNOR U36813 ( .A(n28553), .B(n36856), .Z(n28555) );
  XNOR U36814 ( .A(q[3]), .B(DB[1158]), .Z(n36856) );
  XNOR U36815 ( .A(q[2]), .B(DB[1157]), .Z(n28553) );
  XOR U36816 ( .A(n36857), .B(n28451), .Z(n28379) );
  XOR U36817 ( .A(n36858), .B(n28443), .Z(n28451) );
  XOR U36818 ( .A(n36859), .B(n28432), .Z(n28443) );
  XNOR U36819 ( .A(q[14]), .B(DB[1184]), .Z(n28432) );
  IV U36820 ( .A(n28431), .Z(n36859) );
  XNOR U36821 ( .A(n28429), .B(n36860), .Z(n28431) );
  XNOR U36822 ( .A(q[13]), .B(DB[1183]), .Z(n36860) );
  XNOR U36823 ( .A(q[12]), .B(DB[1182]), .Z(n28429) );
  IV U36824 ( .A(n28442), .Z(n36858) );
  XOR U36825 ( .A(n36861), .B(n36862), .Z(n28442) );
  XNOR U36826 ( .A(n28438), .B(n28440), .Z(n36862) );
  XNOR U36827 ( .A(q[8]), .B(DB[1178]), .Z(n28440) );
  XNOR U36828 ( .A(q[11]), .B(DB[1181]), .Z(n28438) );
  IV U36829 ( .A(n28437), .Z(n36861) );
  XNOR U36830 ( .A(n28435), .B(n36863), .Z(n28437) );
  XNOR U36831 ( .A(q[10]), .B(DB[1180]), .Z(n36863) );
  XNOR U36832 ( .A(q[9]), .B(DB[1179]), .Z(n28435) );
  IV U36833 ( .A(n28450), .Z(n36857) );
  XOR U36834 ( .A(n36864), .B(n36865), .Z(n28450) );
  XNOR U36835 ( .A(n28467), .B(n28448), .Z(n36865) );
  XNOR U36836 ( .A(q[0]), .B(DB[1170]), .Z(n28448) );
  XOR U36837 ( .A(n36866), .B(n28456), .Z(n28467) );
  XNOR U36838 ( .A(q[7]), .B(DB[1177]), .Z(n28456) );
  IV U36839 ( .A(n28455), .Z(n36866) );
  XNOR U36840 ( .A(n28453), .B(n36867), .Z(n28455) );
  XNOR U36841 ( .A(q[6]), .B(DB[1176]), .Z(n36867) );
  XNOR U36842 ( .A(q[5]), .B(DB[1175]), .Z(n28453) );
  IV U36843 ( .A(n28466), .Z(n36864) );
  XOR U36844 ( .A(n36868), .B(n36869), .Z(n28466) );
  XNOR U36845 ( .A(n28462), .B(n28464), .Z(n36869) );
  XNOR U36846 ( .A(q[1]), .B(DB[1171]), .Z(n28464) );
  XNOR U36847 ( .A(q[4]), .B(DB[1174]), .Z(n28462) );
  IV U36848 ( .A(n28461), .Z(n36868) );
  XNOR U36849 ( .A(n28459), .B(n36870), .Z(n28461) );
  XNOR U36850 ( .A(q[3]), .B(DB[1173]), .Z(n36870) );
  XNOR U36851 ( .A(q[2]), .B(DB[1172]), .Z(n28459) );
  XOR U36852 ( .A(n36871), .B(n28357), .Z(n28285) );
  XOR U36853 ( .A(n36872), .B(n28349), .Z(n28357) );
  XOR U36854 ( .A(n36873), .B(n28338), .Z(n28349) );
  XNOR U36855 ( .A(q[14]), .B(DB[1199]), .Z(n28338) );
  IV U36856 ( .A(n28337), .Z(n36873) );
  XNOR U36857 ( .A(n28335), .B(n36874), .Z(n28337) );
  XNOR U36858 ( .A(q[13]), .B(DB[1198]), .Z(n36874) );
  XNOR U36859 ( .A(q[12]), .B(DB[1197]), .Z(n28335) );
  IV U36860 ( .A(n28348), .Z(n36872) );
  XOR U36861 ( .A(n36875), .B(n36876), .Z(n28348) );
  XNOR U36862 ( .A(n28344), .B(n28346), .Z(n36876) );
  XNOR U36863 ( .A(q[8]), .B(DB[1193]), .Z(n28346) );
  XNOR U36864 ( .A(q[11]), .B(DB[1196]), .Z(n28344) );
  IV U36865 ( .A(n28343), .Z(n36875) );
  XNOR U36866 ( .A(n28341), .B(n36877), .Z(n28343) );
  XNOR U36867 ( .A(q[10]), .B(DB[1195]), .Z(n36877) );
  XNOR U36868 ( .A(q[9]), .B(DB[1194]), .Z(n28341) );
  IV U36869 ( .A(n28356), .Z(n36871) );
  XOR U36870 ( .A(n36878), .B(n36879), .Z(n28356) );
  XNOR U36871 ( .A(n28373), .B(n28354), .Z(n36879) );
  XNOR U36872 ( .A(q[0]), .B(DB[1185]), .Z(n28354) );
  XOR U36873 ( .A(n36880), .B(n28362), .Z(n28373) );
  XNOR U36874 ( .A(q[7]), .B(DB[1192]), .Z(n28362) );
  IV U36875 ( .A(n28361), .Z(n36880) );
  XNOR U36876 ( .A(n28359), .B(n36881), .Z(n28361) );
  XNOR U36877 ( .A(q[6]), .B(DB[1191]), .Z(n36881) );
  XNOR U36878 ( .A(q[5]), .B(DB[1190]), .Z(n28359) );
  IV U36879 ( .A(n28372), .Z(n36878) );
  XOR U36880 ( .A(n36882), .B(n36883), .Z(n28372) );
  XNOR U36881 ( .A(n28368), .B(n28370), .Z(n36883) );
  XNOR U36882 ( .A(q[1]), .B(DB[1186]), .Z(n28370) );
  XNOR U36883 ( .A(q[4]), .B(DB[1189]), .Z(n28368) );
  IV U36884 ( .A(n28367), .Z(n36882) );
  XNOR U36885 ( .A(n28365), .B(n36884), .Z(n28367) );
  XNOR U36886 ( .A(q[3]), .B(DB[1188]), .Z(n36884) );
  XNOR U36887 ( .A(q[2]), .B(DB[1187]), .Z(n28365) );
  XOR U36888 ( .A(n36885), .B(n28263), .Z(n28191) );
  XOR U36889 ( .A(n36886), .B(n28255), .Z(n28263) );
  XOR U36890 ( .A(n36887), .B(n28244), .Z(n28255) );
  XNOR U36891 ( .A(q[14]), .B(DB[1214]), .Z(n28244) );
  IV U36892 ( .A(n28243), .Z(n36887) );
  XNOR U36893 ( .A(n28241), .B(n36888), .Z(n28243) );
  XNOR U36894 ( .A(q[13]), .B(DB[1213]), .Z(n36888) );
  XNOR U36895 ( .A(q[12]), .B(DB[1212]), .Z(n28241) );
  IV U36896 ( .A(n28254), .Z(n36886) );
  XOR U36897 ( .A(n36889), .B(n36890), .Z(n28254) );
  XNOR U36898 ( .A(n28250), .B(n28252), .Z(n36890) );
  XNOR U36899 ( .A(q[8]), .B(DB[1208]), .Z(n28252) );
  XNOR U36900 ( .A(q[11]), .B(DB[1211]), .Z(n28250) );
  IV U36901 ( .A(n28249), .Z(n36889) );
  XNOR U36902 ( .A(n28247), .B(n36891), .Z(n28249) );
  XNOR U36903 ( .A(q[10]), .B(DB[1210]), .Z(n36891) );
  XNOR U36904 ( .A(q[9]), .B(DB[1209]), .Z(n28247) );
  IV U36905 ( .A(n28262), .Z(n36885) );
  XOR U36906 ( .A(n36892), .B(n36893), .Z(n28262) );
  XNOR U36907 ( .A(n28279), .B(n28260), .Z(n36893) );
  XNOR U36908 ( .A(q[0]), .B(DB[1200]), .Z(n28260) );
  XOR U36909 ( .A(n36894), .B(n28268), .Z(n28279) );
  XNOR U36910 ( .A(q[7]), .B(DB[1207]), .Z(n28268) );
  IV U36911 ( .A(n28267), .Z(n36894) );
  XNOR U36912 ( .A(n28265), .B(n36895), .Z(n28267) );
  XNOR U36913 ( .A(q[6]), .B(DB[1206]), .Z(n36895) );
  XNOR U36914 ( .A(q[5]), .B(DB[1205]), .Z(n28265) );
  IV U36915 ( .A(n28278), .Z(n36892) );
  XOR U36916 ( .A(n36896), .B(n36897), .Z(n28278) );
  XNOR U36917 ( .A(n28274), .B(n28276), .Z(n36897) );
  XNOR U36918 ( .A(q[1]), .B(DB[1201]), .Z(n28276) );
  XNOR U36919 ( .A(q[4]), .B(DB[1204]), .Z(n28274) );
  IV U36920 ( .A(n28273), .Z(n36896) );
  XNOR U36921 ( .A(n28271), .B(n36898), .Z(n28273) );
  XNOR U36922 ( .A(q[3]), .B(DB[1203]), .Z(n36898) );
  XNOR U36923 ( .A(q[2]), .B(DB[1202]), .Z(n28271) );
  XOR U36924 ( .A(n36899), .B(n28169), .Z(n28097) );
  XOR U36925 ( .A(n36900), .B(n28161), .Z(n28169) );
  XOR U36926 ( .A(n36901), .B(n28150), .Z(n28161) );
  XNOR U36927 ( .A(q[14]), .B(DB[1229]), .Z(n28150) );
  IV U36928 ( .A(n28149), .Z(n36901) );
  XNOR U36929 ( .A(n28147), .B(n36902), .Z(n28149) );
  XNOR U36930 ( .A(q[13]), .B(DB[1228]), .Z(n36902) );
  XNOR U36931 ( .A(q[12]), .B(DB[1227]), .Z(n28147) );
  IV U36932 ( .A(n28160), .Z(n36900) );
  XOR U36933 ( .A(n36903), .B(n36904), .Z(n28160) );
  XNOR U36934 ( .A(n28156), .B(n28158), .Z(n36904) );
  XNOR U36935 ( .A(q[8]), .B(DB[1223]), .Z(n28158) );
  XNOR U36936 ( .A(q[11]), .B(DB[1226]), .Z(n28156) );
  IV U36937 ( .A(n28155), .Z(n36903) );
  XNOR U36938 ( .A(n28153), .B(n36905), .Z(n28155) );
  XNOR U36939 ( .A(q[10]), .B(DB[1225]), .Z(n36905) );
  XNOR U36940 ( .A(q[9]), .B(DB[1224]), .Z(n28153) );
  IV U36941 ( .A(n28168), .Z(n36899) );
  XOR U36942 ( .A(n36906), .B(n36907), .Z(n28168) );
  XNOR U36943 ( .A(n28185), .B(n28166), .Z(n36907) );
  XNOR U36944 ( .A(q[0]), .B(DB[1215]), .Z(n28166) );
  XOR U36945 ( .A(n36908), .B(n28174), .Z(n28185) );
  XNOR U36946 ( .A(q[7]), .B(DB[1222]), .Z(n28174) );
  IV U36947 ( .A(n28173), .Z(n36908) );
  XNOR U36948 ( .A(n28171), .B(n36909), .Z(n28173) );
  XNOR U36949 ( .A(q[6]), .B(DB[1221]), .Z(n36909) );
  XNOR U36950 ( .A(q[5]), .B(DB[1220]), .Z(n28171) );
  IV U36951 ( .A(n28184), .Z(n36906) );
  XOR U36952 ( .A(n36910), .B(n36911), .Z(n28184) );
  XNOR U36953 ( .A(n28180), .B(n28182), .Z(n36911) );
  XNOR U36954 ( .A(q[1]), .B(DB[1216]), .Z(n28182) );
  XNOR U36955 ( .A(q[4]), .B(DB[1219]), .Z(n28180) );
  IV U36956 ( .A(n28179), .Z(n36910) );
  XNOR U36957 ( .A(n28177), .B(n36912), .Z(n28179) );
  XNOR U36958 ( .A(q[3]), .B(DB[1218]), .Z(n36912) );
  XNOR U36959 ( .A(q[2]), .B(DB[1217]), .Z(n28177) );
  XOR U36960 ( .A(n36913), .B(n28075), .Z(n28003) );
  XOR U36961 ( .A(n36914), .B(n28067), .Z(n28075) );
  XOR U36962 ( .A(n36915), .B(n28056), .Z(n28067) );
  XNOR U36963 ( .A(q[14]), .B(DB[1244]), .Z(n28056) );
  IV U36964 ( .A(n28055), .Z(n36915) );
  XNOR U36965 ( .A(n28053), .B(n36916), .Z(n28055) );
  XNOR U36966 ( .A(q[13]), .B(DB[1243]), .Z(n36916) );
  XNOR U36967 ( .A(q[12]), .B(DB[1242]), .Z(n28053) );
  IV U36968 ( .A(n28066), .Z(n36914) );
  XOR U36969 ( .A(n36917), .B(n36918), .Z(n28066) );
  XNOR U36970 ( .A(n28062), .B(n28064), .Z(n36918) );
  XNOR U36971 ( .A(q[8]), .B(DB[1238]), .Z(n28064) );
  XNOR U36972 ( .A(q[11]), .B(DB[1241]), .Z(n28062) );
  IV U36973 ( .A(n28061), .Z(n36917) );
  XNOR U36974 ( .A(n28059), .B(n36919), .Z(n28061) );
  XNOR U36975 ( .A(q[10]), .B(DB[1240]), .Z(n36919) );
  XNOR U36976 ( .A(q[9]), .B(DB[1239]), .Z(n28059) );
  IV U36977 ( .A(n28074), .Z(n36913) );
  XOR U36978 ( .A(n36920), .B(n36921), .Z(n28074) );
  XNOR U36979 ( .A(n28091), .B(n28072), .Z(n36921) );
  XNOR U36980 ( .A(q[0]), .B(DB[1230]), .Z(n28072) );
  XOR U36981 ( .A(n36922), .B(n28080), .Z(n28091) );
  XNOR U36982 ( .A(q[7]), .B(DB[1237]), .Z(n28080) );
  IV U36983 ( .A(n28079), .Z(n36922) );
  XNOR U36984 ( .A(n28077), .B(n36923), .Z(n28079) );
  XNOR U36985 ( .A(q[6]), .B(DB[1236]), .Z(n36923) );
  XNOR U36986 ( .A(q[5]), .B(DB[1235]), .Z(n28077) );
  IV U36987 ( .A(n28090), .Z(n36920) );
  XOR U36988 ( .A(n36924), .B(n36925), .Z(n28090) );
  XNOR U36989 ( .A(n28086), .B(n28088), .Z(n36925) );
  XNOR U36990 ( .A(q[1]), .B(DB[1231]), .Z(n28088) );
  XNOR U36991 ( .A(q[4]), .B(DB[1234]), .Z(n28086) );
  IV U36992 ( .A(n28085), .Z(n36924) );
  XNOR U36993 ( .A(n28083), .B(n36926), .Z(n28085) );
  XNOR U36994 ( .A(q[3]), .B(DB[1233]), .Z(n36926) );
  XNOR U36995 ( .A(q[2]), .B(DB[1232]), .Z(n28083) );
  XOR U36996 ( .A(n36927), .B(n27981), .Z(n27909) );
  XOR U36997 ( .A(n36928), .B(n27973), .Z(n27981) );
  XOR U36998 ( .A(n36929), .B(n27962), .Z(n27973) );
  XNOR U36999 ( .A(q[14]), .B(DB[1259]), .Z(n27962) );
  IV U37000 ( .A(n27961), .Z(n36929) );
  XNOR U37001 ( .A(n27959), .B(n36930), .Z(n27961) );
  XNOR U37002 ( .A(q[13]), .B(DB[1258]), .Z(n36930) );
  XNOR U37003 ( .A(q[12]), .B(DB[1257]), .Z(n27959) );
  IV U37004 ( .A(n27972), .Z(n36928) );
  XOR U37005 ( .A(n36931), .B(n36932), .Z(n27972) );
  XNOR U37006 ( .A(n27968), .B(n27970), .Z(n36932) );
  XNOR U37007 ( .A(q[8]), .B(DB[1253]), .Z(n27970) );
  XNOR U37008 ( .A(q[11]), .B(DB[1256]), .Z(n27968) );
  IV U37009 ( .A(n27967), .Z(n36931) );
  XNOR U37010 ( .A(n27965), .B(n36933), .Z(n27967) );
  XNOR U37011 ( .A(q[10]), .B(DB[1255]), .Z(n36933) );
  XNOR U37012 ( .A(q[9]), .B(DB[1254]), .Z(n27965) );
  IV U37013 ( .A(n27980), .Z(n36927) );
  XOR U37014 ( .A(n36934), .B(n36935), .Z(n27980) );
  XNOR U37015 ( .A(n27997), .B(n27978), .Z(n36935) );
  XNOR U37016 ( .A(q[0]), .B(DB[1245]), .Z(n27978) );
  XOR U37017 ( .A(n36936), .B(n27986), .Z(n27997) );
  XNOR U37018 ( .A(q[7]), .B(DB[1252]), .Z(n27986) );
  IV U37019 ( .A(n27985), .Z(n36936) );
  XNOR U37020 ( .A(n27983), .B(n36937), .Z(n27985) );
  XNOR U37021 ( .A(q[6]), .B(DB[1251]), .Z(n36937) );
  XNOR U37022 ( .A(q[5]), .B(DB[1250]), .Z(n27983) );
  IV U37023 ( .A(n27996), .Z(n36934) );
  XOR U37024 ( .A(n36938), .B(n36939), .Z(n27996) );
  XNOR U37025 ( .A(n27992), .B(n27994), .Z(n36939) );
  XNOR U37026 ( .A(q[1]), .B(DB[1246]), .Z(n27994) );
  XNOR U37027 ( .A(q[4]), .B(DB[1249]), .Z(n27992) );
  IV U37028 ( .A(n27991), .Z(n36938) );
  XNOR U37029 ( .A(n27989), .B(n36940), .Z(n27991) );
  XNOR U37030 ( .A(q[3]), .B(DB[1248]), .Z(n36940) );
  XNOR U37031 ( .A(q[2]), .B(DB[1247]), .Z(n27989) );
  XOR U37032 ( .A(n36941), .B(n27887), .Z(n27815) );
  XOR U37033 ( .A(n36942), .B(n27879), .Z(n27887) );
  XOR U37034 ( .A(n36943), .B(n27868), .Z(n27879) );
  XNOR U37035 ( .A(q[14]), .B(DB[1274]), .Z(n27868) );
  IV U37036 ( .A(n27867), .Z(n36943) );
  XNOR U37037 ( .A(n27865), .B(n36944), .Z(n27867) );
  XNOR U37038 ( .A(q[13]), .B(DB[1273]), .Z(n36944) );
  XNOR U37039 ( .A(q[12]), .B(DB[1272]), .Z(n27865) );
  IV U37040 ( .A(n27878), .Z(n36942) );
  XOR U37041 ( .A(n36945), .B(n36946), .Z(n27878) );
  XNOR U37042 ( .A(n27874), .B(n27876), .Z(n36946) );
  XNOR U37043 ( .A(q[8]), .B(DB[1268]), .Z(n27876) );
  XNOR U37044 ( .A(q[11]), .B(DB[1271]), .Z(n27874) );
  IV U37045 ( .A(n27873), .Z(n36945) );
  XNOR U37046 ( .A(n27871), .B(n36947), .Z(n27873) );
  XNOR U37047 ( .A(q[10]), .B(DB[1270]), .Z(n36947) );
  XNOR U37048 ( .A(q[9]), .B(DB[1269]), .Z(n27871) );
  IV U37049 ( .A(n27886), .Z(n36941) );
  XOR U37050 ( .A(n36948), .B(n36949), .Z(n27886) );
  XNOR U37051 ( .A(n27903), .B(n27884), .Z(n36949) );
  XNOR U37052 ( .A(q[0]), .B(DB[1260]), .Z(n27884) );
  XOR U37053 ( .A(n36950), .B(n27892), .Z(n27903) );
  XNOR U37054 ( .A(q[7]), .B(DB[1267]), .Z(n27892) );
  IV U37055 ( .A(n27891), .Z(n36950) );
  XNOR U37056 ( .A(n27889), .B(n36951), .Z(n27891) );
  XNOR U37057 ( .A(q[6]), .B(DB[1266]), .Z(n36951) );
  XNOR U37058 ( .A(q[5]), .B(DB[1265]), .Z(n27889) );
  IV U37059 ( .A(n27902), .Z(n36948) );
  XOR U37060 ( .A(n36952), .B(n36953), .Z(n27902) );
  XNOR U37061 ( .A(n27898), .B(n27900), .Z(n36953) );
  XNOR U37062 ( .A(q[1]), .B(DB[1261]), .Z(n27900) );
  XNOR U37063 ( .A(q[4]), .B(DB[1264]), .Z(n27898) );
  IV U37064 ( .A(n27897), .Z(n36952) );
  XNOR U37065 ( .A(n27895), .B(n36954), .Z(n27897) );
  XNOR U37066 ( .A(q[3]), .B(DB[1263]), .Z(n36954) );
  XNOR U37067 ( .A(q[2]), .B(DB[1262]), .Z(n27895) );
  XOR U37068 ( .A(n36955), .B(n27793), .Z(n27721) );
  XOR U37069 ( .A(n36956), .B(n27785), .Z(n27793) );
  XOR U37070 ( .A(n36957), .B(n27774), .Z(n27785) );
  XNOR U37071 ( .A(q[14]), .B(DB[1289]), .Z(n27774) );
  IV U37072 ( .A(n27773), .Z(n36957) );
  XNOR U37073 ( .A(n27771), .B(n36958), .Z(n27773) );
  XNOR U37074 ( .A(q[13]), .B(DB[1288]), .Z(n36958) );
  XNOR U37075 ( .A(q[12]), .B(DB[1287]), .Z(n27771) );
  IV U37076 ( .A(n27784), .Z(n36956) );
  XOR U37077 ( .A(n36959), .B(n36960), .Z(n27784) );
  XNOR U37078 ( .A(n27780), .B(n27782), .Z(n36960) );
  XNOR U37079 ( .A(q[8]), .B(DB[1283]), .Z(n27782) );
  XNOR U37080 ( .A(q[11]), .B(DB[1286]), .Z(n27780) );
  IV U37081 ( .A(n27779), .Z(n36959) );
  XNOR U37082 ( .A(n27777), .B(n36961), .Z(n27779) );
  XNOR U37083 ( .A(q[10]), .B(DB[1285]), .Z(n36961) );
  XNOR U37084 ( .A(q[9]), .B(DB[1284]), .Z(n27777) );
  IV U37085 ( .A(n27792), .Z(n36955) );
  XOR U37086 ( .A(n36962), .B(n36963), .Z(n27792) );
  XNOR U37087 ( .A(n27809), .B(n27790), .Z(n36963) );
  XNOR U37088 ( .A(q[0]), .B(DB[1275]), .Z(n27790) );
  XOR U37089 ( .A(n36964), .B(n27798), .Z(n27809) );
  XNOR U37090 ( .A(q[7]), .B(DB[1282]), .Z(n27798) );
  IV U37091 ( .A(n27797), .Z(n36964) );
  XNOR U37092 ( .A(n27795), .B(n36965), .Z(n27797) );
  XNOR U37093 ( .A(q[6]), .B(DB[1281]), .Z(n36965) );
  XNOR U37094 ( .A(q[5]), .B(DB[1280]), .Z(n27795) );
  IV U37095 ( .A(n27808), .Z(n36962) );
  XOR U37096 ( .A(n36966), .B(n36967), .Z(n27808) );
  XNOR U37097 ( .A(n27804), .B(n27806), .Z(n36967) );
  XNOR U37098 ( .A(q[1]), .B(DB[1276]), .Z(n27806) );
  XNOR U37099 ( .A(q[4]), .B(DB[1279]), .Z(n27804) );
  IV U37100 ( .A(n27803), .Z(n36966) );
  XNOR U37101 ( .A(n27801), .B(n36968), .Z(n27803) );
  XNOR U37102 ( .A(q[3]), .B(DB[1278]), .Z(n36968) );
  XNOR U37103 ( .A(q[2]), .B(DB[1277]), .Z(n27801) );
  XOR U37104 ( .A(n36969), .B(n27699), .Z(n27627) );
  XOR U37105 ( .A(n36970), .B(n27691), .Z(n27699) );
  XOR U37106 ( .A(n36971), .B(n27680), .Z(n27691) );
  XNOR U37107 ( .A(q[14]), .B(DB[1304]), .Z(n27680) );
  IV U37108 ( .A(n27679), .Z(n36971) );
  XNOR U37109 ( .A(n27677), .B(n36972), .Z(n27679) );
  XNOR U37110 ( .A(q[13]), .B(DB[1303]), .Z(n36972) );
  XNOR U37111 ( .A(q[12]), .B(DB[1302]), .Z(n27677) );
  IV U37112 ( .A(n27690), .Z(n36970) );
  XOR U37113 ( .A(n36973), .B(n36974), .Z(n27690) );
  XNOR U37114 ( .A(n27686), .B(n27688), .Z(n36974) );
  XNOR U37115 ( .A(q[8]), .B(DB[1298]), .Z(n27688) );
  XNOR U37116 ( .A(q[11]), .B(DB[1301]), .Z(n27686) );
  IV U37117 ( .A(n27685), .Z(n36973) );
  XNOR U37118 ( .A(n27683), .B(n36975), .Z(n27685) );
  XNOR U37119 ( .A(q[10]), .B(DB[1300]), .Z(n36975) );
  XNOR U37120 ( .A(q[9]), .B(DB[1299]), .Z(n27683) );
  IV U37121 ( .A(n27698), .Z(n36969) );
  XOR U37122 ( .A(n36976), .B(n36977), .Z(n27698) );
  XNOR U37123 ( .A(n27715), .B(n27696), .Z(n36977) );
  XNOR U37124 ( .A(q[0]), .B(DB[1290]), .Z(n27696) );
  XOR U37125 ( .A(n36978), .B(n27704), .Z(n27715) );
  XNOR U37126 ( .A(q[7]), .B(DB[1297]), .Z(n27704) );
  IV U37127 ( .A(n27703), .Z(n36978) );
  XNOR U37128 ( .A(n27701), .B(n36979), .Z(n27703) );
  XNOR U37129 ( .A(q[6]), .B(DB[1296]), .Z(n36979) );
  XNOR U37130 ( .A(q[5]), .B(DB[1295]), .Z(n27701) );
  IV U37131 ( .A(n27714), .Z(n36976) );
  XOR U37132 ( .A(n36980), .B(n36981), .Z(n27714) );
  XNOR U37133 ( .A(n27710), .B(n27712), .Z(n36981) );
  XNOR U37134 ( .A(q[1]), .B(DB[1291]), .Z(n27712) );
  XNOR U37135 ( .A(q[4]), .B(DB[1294]), .Z(n27710) );
  IV U37136 ( .A(n27709), .Z(n36980) );
  XNOR U37137 ( .A(n27707), .B(n36982), .Z(n27709) );
  XNOR U37138 ( .A(q[3]), .B(DB[1293]), .Z(n36982) );
  XNOR U37139 ( .A(q[2]), .B(DB[1292]), .Z(n27707) );
  XOR U37140 ( .A(n36983), .B(n27605), .Z(n27533) );
  XOR U37141 ( .A(n36984), .B(n27597), .Z(n27605) );
  XOR U37142 ( .A(n36985), .B(n27586), .Z(n27597) );
  XNOR U37143 ( .A(q[14]), .B(DB[1319]), .Z(n27586) );
  IV U37144 ( .A(n27585), .Z(n36985) );
  XNOR U37145 ( .A(n27583), .B(n36986), .Z(n27585) );
  XNOR U37146 ( .A(q[13]), .B(DB[1318]), .Z(n36986) );
  XNOR U37147 ( .A(q[12]), .B(DB[1317]), .Z(n27583) );
  IV U37148 ( .A(n27596), .Z(n36984) );
  XOR U37149 ( .A(n36987), .B(n36988), .Z(n27596) );
  XNOR U37150 ( .A(n27592), .B(n27594), .Z(n36988) );
  XNOR U37151 ( .A(q[8]), .B(DB[1313]), .Z(n27594) );
  XNOR U37152 ( .A(q[11]), .B(DB[1316]), .Z(n27592) );
  IV U37153 ( .A(n27591), .Z(n36987) );
  XNOR U37154 ( .A(n27589), .B(n36989), .Z(n27591) );
  XNOR U37155 ( .A(q[10]), .B(DB[1315]), .Z(n36989) );
  XNOR U37156 ( .A(q[9]), .B(DB[1314]), .Z(n27589) );
  IV U37157 ( .A(n27604), .Z(n36983) );
  XOR U37158 ( .A(n36990), .B(n36991), .Z(n27604) );
  XNOR U37159 ( .A(n27621), .B(n27602), .Z(n36991) );
  XNOR U37160 ( .A(q[0]), .B(DB[1305]), .Z(n27602) );
  XOR U37161 ( .A(n36992), .B(n27610), .Z(n27621) );
  XNOR U37162 ( .A(q[7]), .B(DB[1312]), .Z(n27610) );
  IV U37163 ( .A(n27609), .Z(n36992) );
  XNOR U37164 ( .A(n27607), .B(n36993), .Z(n27609) );
  XNOR U37165 ( .A(q[6]), .B(DB[1311]), .Z(n36993) );
  XNOR U37166 ( .A(q[5]), .B(DB[1310]), .Z(n27607) );
  IV U37167 ( .A(n27620), .Z(n36990) );
  XOR U37168 ( .A(n36994), .B(n36995), .Z(n27620) );
  XNOR U37169 ( .A(n27616), .B(n27618), .Z(n36995) );
  XNOR U37170 ( .A(q[1]), .B(DB[1306]), .Z(n27618) );
  XNOR U37171 ( .A(q[4]), .B(DB[1309]), .Z(n27616) );
  IV U37172 ( .A(n27615), .Z(n36994) );
  XNOR U37173 ( .A(n27613), .B(n36996), .Z(n27615) );
  XNOR U37174 ( .A(q[3]), .B(DB[1308]), .Z(n36996) );
  XNOR U37175 ( .A(q[2]), .B(DB[1307]), .Z(n27613) );
  XOR U37176 ( .A(n36997), .B(n27511), .Z(n27439) );
  XOR U37177 ( .A(n36998), .B(n27503), .Z(n27511) );
  XOR U37178 ( .A(n36999), .B(n27492), .Z(n27503) );
  XNOR U37179 ( .A(q[14]), .B(DB[1334]), .Z(n27492) );
  IV U37180 ( .A(n27491), .Z(n36999) );
  XNOR U37181 ( .A(n27489), .B(n37000), .Z(n27491) );
  XNOR U37182 ( .A(q[13]), .B(DB[1333]), .Z(n37000) );
  XNOR U37183 ( .A(q[12]), .B(DB[1332]), .Z(n27489) );
  IV U37184 ( .A(n27502), .Z(n36998) );
  XOR U37185 ( .A(n37001), .B(n37002), .Z(n27502) );
  XNOR U37186 ( .A(n27498), .B(n27500), .Z(n37002) );
  XNOR U37187 ( .A(q[8]), .B(DB[1328]), .Z(n27500) );
  XNOR U37188 ( .A(q[11]), .B(DB[1331]), .Z(n27498) );
  IV U37189 ( .A(n27497), .Z(n37001) );
  XNOR U37190 ( .A(n27495), .B(n37003), .Z(n27497) );
  XNOR U37191 ( .A(q[10]), .B(DB[1330]), .Z(n37003) );
  XNOR U37192 ( .A(q[9]), .B(DB[1329]), .Z(n27495) );
  IV U37193 ( .A(n27510), .Z(n36997) );
  XOR U37194 ( .A(n37004), .B(n37005), .Z(n27510) );
  XNOR U37195 ( .A(n27527), .B(n27508), .Z(n37005) );
  XNOR U37196 ( .A(q[0]), .B(DB[1320]), .Z(n27508) );
  XOR U37197 ( .A(n37006), .B(n27516), .Z(n27527) );
  XNOR U37198 ( .A(q[7]), .B(DB[1327]), .Z(n27516) );
  IV U37199 ( .A(n27515), .Z(n37006) );
  XNOR U37200 ( .A(n27513), .B(n37007), .Z(n27515) );
  XNOR U37201 ( .A(q[6]), .B(DB[1326]), .Z(n37007) );
  XNOR U37202 ( .A(q[5]), .B(DB[1325]), .Z(n27513) );
  IV U37203 ( .A(n27526), .Z(n37004) );
  XOR U37204 ( .A(n37008), .B(n37009), .Z(n27526) );
  XNOR U37205 ( .A(n27522), .B(n27524), .Z(n37009) );
  XNOR U37206 ( .A(q[1]), .B(DB[1321]), .Z(n27524) );
  XNOR U37207 ( .A(q[4]), .B(DB[1324]), .Z(n27522) );
  IV U37208 ( .A(n27521), .Z(n37008) );
  XNOR U37209 ( .A(n27519), .B(n37010), .Z(n27521) );
  XNOR U37210 ( .A(q[3]), .B(DB[1323]), .Z(n37010) );
  XNOR U37211 ( .A(q[2]), .B(DB[1322]), .Z(n27519) );
  XOR U37212 ( .A(n37011), .B(n27417), .Z(n27345) );
  XOR U37213 ( .A(n37012), .B(n27409), .Z(n27417) );
  XOR U37214 ( .A(n37013), .B(n27398), .Z(n27409) );
  XNOR U37215 ( .A(q[14]), .B(DB[1349]), .Z(n27398) );
  IV U37216 ( .A(n27397), .Z(n37013) );
  XNOR U37217 ( .A(n27395), .B(n37014), .Z(n27397) );
  XNOR U37218 ( .A(q[13]), .B(DB[1348]), .Z(n37014) );
  XNOR U37219 ( .A(q[12]), .B(DB[1347]), .Z(n27395) );
  IV U37220 ( .A(n27408), .Z(n37012) );
  XOR U37221 ( .A(n37015), .B(n37016), .Z(n27408) );
  XNOR U37222 ( .A(n27404), .B(n27406), .Z(n37016) );
  XNOR U37223 ( .A(q[8]), .B(DB[1343]), .Z(n27406) );
  XNOR U37224 ( .A(q[11]), .B(DB[1346]), .Z(n27404) );
  IV U37225 ( .A(n27403), .Z(n37015) );
  XNOR U37226 ( .A(n27401), .B(n37017), .Z(n27403) );
  XNOR U37227 ( .A(q[10]), .B(DB[1345]), .Z(n37017) );
  XNOR U37228 ( .A(q[9]), .B(DB[1344]), .Z(n27401) );
  IV U37229 ( .A(n27416), .Z(n37011) );
  XOR U37230 ( .A(n37018), .B(n37019), .Z(n27416) );
  XNOR U37231 ( .A(n27433), .B(n27414), .Z(n37019) );
  XNOR U37232 ( .A(q[0]), .B(DB[1335]), .Z(n27414) );
  XOR U37233 ( .A(n37020), .B(n27422), .Z(n27433) );
  XNOR U37234 ( .A(q[7]), .B(DB[1342]), .Z(n27422) );
  IV U37235 ( .A(n27421), .Z(n37020) );
  XNOR U37236 ( .A(n27419), .B(n37021), .Z(n27421) );
  XNOR U37237 ( .A(q[6]), .B(DB[1341]), .Z(n37021) );
  XNOR U37238 ( .A(q[5]), .B(DB[1340]), .Z(n27419) );
  IV U37239 ( .A(n27432), .Z(n37018) );
  XOR U37240 ( .A(n37022), .B(n37023), .Z(n27432) );
  XNOR U37241 ( .A(n27428), .B(n27430), .Z(n37023) );
  XNOR U37242 ( .A(q[1]), .B(DB[1336]), .Z(n27430) );
  XNOR U37243 ( .A(q[4]), .B(DB[1339]), .Z(n27428) );
  IV U37244 ( .A(n27427), .Z(n37022) );
  XNOR U37245 ( .A(n27425), .B(n37024), .Z(n27427) );
  XNOR U37246 ( .A(q[3]), .B(DB[1338]), .Z(n37024) );
  XNOR U37247 ( .A(q[2]), .B(DB[1337]), .Z(n27425) );
  XOR U37248 ( .A(n37025), .B(n27323), .Z(n27251) );
  XOR U37249 ( .A(n37026), .B(n27315), .Z(n27323) );
  XOR U37250 ( .A(n37027), .B(n27304), .Z(n27315) );
  XNOR U37251 ( .A(q[14]), .B(DB[1364]), .Z(n27304) );
  IV U37252 ( .A(n27303), .Z(n37027) );
  XNOR U37253 ( .A(n27301), .B(n37028), .Z(n27303) );
  XNOR U37254 ( .A(q[13]), .B(DB[1363]), .Z(n37028) );
  XNOR U37255 ( .A(q[12]), .B(DB[1362]), .Z(n27301) );
  IV U37256 ( .A(n27314), .Z(n37026) );
  XOR U37257 ( .A(n37029), .B(n37030), .Z(n27314) );
  XNOR U37258 ( .A(n27310), .B(n27312), .Z(n37030) );
  XNOR U37259 ( .A(q[8]), .B(DB[1358]), .Z(n27312) );
  XNOR U37260 ( .A(q[11]), .B(DB[1361]), .Z(n27310) );
  IV U37261 ( .A(n27309), .Z(n37029) );
  XNOR U37262 ( .A(n27307), .B(n37031), .Z(n27309) );
  XNOR U37263 ( .A(q[10]), .B(DB[1360]), .Z(n37031) );
  XNOR U37264 ( .A(q[9]), .B(DB[1359]), .Z(n27307) );
  IV U37265 ( .A(n27322), .Z(n37025) );
  XOR U37266 ( .A(n37032), .B(n37033), .Z(n27322) );
  XNOR U37267 ( .A(n27339), .B(n27320), .Z(n37033) );
  XNOR U37268 ( .A(q[0]), .B(DB[1350]), .Z(n27320) );
  XOR U37269 ( .A(n37034), .B(n27328), .Z(n27339) );
  XNOR U37270 ( .A(q[7]), .B(DB[1357]), .Z(n27328) );
  IV U37271 ( .A(n27327), .Z(n37034) );
  XNOR U37272 ( .A(n27325), .B(n37035), .Z(n27327) );
  XNOR U37273 ( .A(q[6]), .B(DB[1356]), .Z(n37035) );
  XNOR U37274 ( .A(q[5]), .B(DB[1355]), .Z(n27325) );
  IV U37275 ( .A(n27338), .Z(n37032) );
  XOR U37276 ( .A(n37036), .B(n37037), .Z(n27338) );
  XNOR U37277 ( .A(n27334), .B(n27336), .Z(n37037) );
  XNOR U37278 ( .A(q[1]), .B(DB[1351]), .Z(n27336) );
  XNOR U37279 ( .A(q[4]), .B(DB[1354]), .Z(n27334) );
  IV U37280 ( .A(n27333), .Z(n37036) );
  XNOR U37281 ( .A(n27331), .B(n37038), .Z(n27333) );
  XNOR U37282 ( .A(q[3]), .B(DB[1353]), .Z(n37038) );
  XNOR U37283 ( .A(q[2]), .B(DB[1352]), .Z(n27331) );
  XOR U37284 ( .A(n37039), .B(n27229), .Z(n27157) );
  XOR U37285 ( .A(n37040), .B(n27221), .Z(n27229) );
  XOR U37286 ( .A(n37041), .B(n27210), .Z(n27221) );
  XNOR U37287 ( .A(q[14]), .B(DB[1379]), .Z(n27210) );
  IV U37288 ( .A(n27209), .Z(n37041) );
  XNOR U37289 ( .A(n27207), .B(n37042), .Z(n27209) );
  XNOR U37290 ( .A(q[13]), .B(DB[1378]), .Z(n37042) );
  XNOR U37291 ( .A(q[12]), .B(DB[1377]), .Z(n27207) );
  IV U37292 ( .A(n27220), .Z(n37040) );
  XOR U37293 ( .A(n37043), .B(n37044), .Z(n27220) );
  XNOR U37294 ( .A(n27216), .B(n27218), .Z(n37044) );
  XNOR U37295 ( .A(q[8]), .B(DB[1373]), .Z(n27218) );
  XNOR U37296 ( .A(q[11]), .B(DB[1376]), .Z(n27216) );
  IV U37297 ( .A(n27215), .Z(n37043) );
  XNOR U37298 ( .A(n27213), .B(n37045), .Z(n27215) );
  XNOR U37299 ( .A(q[10]), .B(DB[1375]), .Z(n37045) );
  XNOR U37300 ( .A(q[9]), .B(DB[1374]), .Z(n27213) );
  IV U37301 ( .A(n27228), .Z(n37039) );
  XOR U37302 ( .A(n37046), .B(n37047), .Z(n27228) );
  XNOR U37303 ( .A(n27245), .B(n27226), .Z(n37047) );
  XNOR U37304 ( .A(q[0]), .B(DB[1365]), .Z(n27226) );
  XOR U37305 ( .A(n37048), .B(n27234), .Z(n27245) );
  XNOR U37306 ( .A(q[7]), .B(DB[1372]), .Z(n27234) );
  IV U37307 ( .A(n27233), .Z(n37048) );
  XNOR U37308 ( .A(n27231), .B(n37049), .Z(n27233) );
  XNOR U37309 ( .A(q[6]), .B(DB[1371]), .Z(n37049) );
  XNOR U37310 ( .A(q[5]), .B(DB[1370]), .Z(n27231) );
  IV U37311 ( .A(n27244), .Z(n37046) );
  XOR U37312 ( .A(n37050), .B(n37051), .Z(n27244) );
  XNOR U37313 ( .A(n27240), .B(n27242), .Z(n37051) );
  XNOR U37314 ( .A(q[1]), .B(DB[1366]), .Z(n27242) );
  XNOR U37315 ( .A(q[4]), .B(DB[1369]), .Z(n27240) );
  IV U37316 ( .A(n27239), .Z(n37050) );
  XNOR U37317 ( .A(n27237), .B(n37052), .Z(n27239) );
  XNOR U37318 ( .A(q[3]), .B(DB[1368]), .Z(n37052) );
  XNOR U37319 ( .A(q[2]), .B(DB[1367]), .Z(n27237) );
  XOR U37320 ( .A(n37053), .B(n27135), .Z(n27063) );
  XOR U37321 ( .A(n37054), .B(n27127), .Z(n27135) );
  XOR U37322 ( .A(n37055), .B(n27116), .Z(n27127) );
  XNOR U37323 ( .A(q[14]), .B(DB[1394]), .Z(n27116) );
  IV U37324 ( .A(n27115), .Z(n37055) );
  XNOR U37325 ( .A(n27113), .B(n37056), .Z(n27115) );
  XNOR U37326 ( .A(q[13]), .B(DB[1393]), .Z(n37056) );
  XNOR U37327 ( .A(q[12]), .B(DB[1392]), .Z(n27113) );
  IV U37328 ( .A(n27126), .Z(n37054) );
  XOR U37329 ( .A(n37057), .B(n37058), .Z(n27126) );
  XNOR U37330 ( .A(n27122), .B(n27124), .Z(n37058) );
  XNOR U37331 ( .A(q[8]), .B(DB[1388]), .Z(n27124) );
  XNOR U37332 ( .A(q[11]), .B(DB[1391]), .Z(n27122) );
  IV U37333 ( .A(n27121), .Z(n37057) );
  XNOR U37334 ( .A(n27119), .B(n37059), .Z(n27121) );
  XNOR U37335 ( .A(q[10]), .B(DB[1390]), .Z(n37059) );
  XNOR U37336 ( .A(q[9]), .B(DB[1389]), .Z(n27119) );
  IV U37337 ( .A(n27134), .Z(n37053) );
  XOR U37338 ( .A(n37060), .B(n37061), .Z(n27134) );
  XNOR U37339 ( .A(n27151), .B(n27132), .Z(n37061) );
  XNOR U37340 ( .A(q[0]), .B(DB[1380]), .Z(n27132) );
  XOR U37341 ( .A(n37062), .B(n27140), .Z(n27151) );
  XNOR U37342 ( .A(q[7]), .B(DB[1387]), .Z(n27140) );
  IV U37343 ( .A(n27139), .Z(n37062) );
  XNOR U37344 ( .A(n27137), .B(n37063), .Z(n27139) );
  XNOR U37345 ( .A(q[6]), .B(DB[1386]), .Z(n37063) );
  XNOR U37346 ( .A(q[5]), .B(DB[1385]), .Z(n27137) );
  IV U37347 ( .A(n27150), .Z(n37060) );
  XOR U37348 ( .A(n37064), .B(n37065), .Z(n27150) );
  XNOR U37349 ( .A(n27146), .B(n27148), .Z(n37065) );
  XNOR U37350 ( .A(q[1]), .B(DB[1381]), .Z(n27148) );
  XNOR U37351 ( .A(q[4]), .B(DB[1384]), .Z(n27146) );
  IV U37352 ( .A(n27145), .Z(n37064) );
  XNOR U37353 ( .A(n27143), .B(n37066), .Z(n27145) );
  XNOR U37354 ( .A(q[3]), .B(DB[1383]), .Z(n37066) );
  XNOR U37355 ( .A(q[2]), .B(DB[1382]), .Z(n27143) );
  XOR U37356 ( .A(n37067), .B(n27041), .Z(n26969) );
  XOR U37357 ( .A(n37068), .B(n27033), .Z(n27041) );
  XOR U37358 ( .A(n37069), .B(n27022), .Z(n27033) );
  XNOR U37359 ( .A(q[14]), .B(DB[1409]), .Z(n27022) );
  IV U37360 ( .A(n27021), .Z(n37069) );
  XNOR U37361 ( .A(n27019), .B(n37070), .Z(n27021) );
  XNOR U37362 ( .A(q[13]), .B(DB[1408]), .Z(n37070) );
  XNOR U37363 ( .A(q[12]), .B(DB[1407]), .Z(n27019) );
  IV U37364 ( .A(n27032), .Z(n37068) );
  XOR U37365 ( .A(n37071), .B(n37072), .Z(n27032) );
  XNOR U37366 ( .A(n27028), .B(n27030), .Z(n37072) );
  XNOR U37367 ( .A(q[8]), .B(DB[1403]), .Z(n27030) );
  XNOR U37368 ( .A(q[11]), .B(DB[1406]), .Z(n27028) );
  IV U37369 ( .A(n27027), .Z(n37071) );
  XNOR U37370 ( .A(n27025), .B(n37073), .Z(n27027) );
  XNOR U37371 ( .A(q[10]), .B(DB[1405]), .Z(n37073) );
  XNOR U37372 ( .A(q[9]), .B(DB[1404]), .Z(n27025) );
  IV U37373 ( .A(n27040), .Z(n37067) );
  XOR U37374 ( .A(n37074), .B(n37075), .Z(n27040) );
  XNOR U37375 ( .A(n27057), .B(n27038), .Z(n37075) );
  XNOR U37376 ( .A(q[0]), .B(DB[1395]), .Z(n27038) );
  XOR U37377 ( .A(n37076), .B(n27046), .Z(n27057) );
  XNOR U37378 ( .A(q[7]), .B(DB[1402]), .Z(n27046) );
  IV U37379 ( .A(n27045), .Z(n37076) );
  XNOR U37380 ( .A(n27043), .B(n37077), .Z(n27045) );
  XNOR U37381 ( .A(q[6]), .B(DB[1401]), .Z(n37077) );
  XNOR U37382 ( .A(q[5]), .B(DB[1400]), .Z(n27043) );
  IV U37383 ( .A(n27056), .Z(n37074) );
  XOR U37384 ( .A(n37078), .B(n37079), .Z(n27056) );
  XNOR U37385 ( .A(n27052), .B(n27054), .Z(n37079) );
  XNOR U37386 ( .A(q[1]), .B(DB[1396]), .Z(n27054) );
  XNOR U37387 ( .A(q[4]), .B(DB[1399]), .Z(n27052) );
  IV U37388 ( .A(n27051), .Z(n37078) );
  XNOR U37389 ( .A(n27049), .B(n37080), .Z(n27051) );
  XNOR U37390 ( .A(q[3]), .B(DB[1398]), .Z(n37080) );
  XNOR U37391 ( .A(q[2]), .B(DB[1397]), .Z(n27049) );
  XOR U37392 ( .A(n37081), .B(n26947), .Z(n26875) );
  XOR U37393 ( .A(n37082), .B(n26939), .Z(n26947) );
  XOR U37394 ( .A(n37083), .B(n26928), .Z(n26939) );
  XNOR U37395 ( .A(q[14]), .B(DB[1424]), .Z(n26928) );
  IV U37396 ( .A(n26927), .Z(n37083) );
  XNOR U37397 ( .A(n26925), .B(n37084), .Z(n26927) );
  XNOR U37398 ( .A(q[13]), .B(DB[1423]), .Z(n37084) );
  XNOR U37399 ( .A(q[12]), .B(DB[1422]), .Z(n26925) );
  IV U37400 ( .A(n26938), .Z(n37082) );
  XOR U37401 ( .A(n37085), .B(n37086), .Z(n26938) );
  XNOR U37402 ( .A(n26934), .B(n26936), .Z(n37086) );
  XNOR U37403 ( .A(q[8]), .B(DB[1418]), .Z(n26936) );
  XNOR U37404 ( .A(q[11]), .B(DB[1421]), .Z(n26934) );
  IV U37405 ( .A(n26933), .Z(n37085) );
  XNOR U37406 ( .A(n26931), .B(n37087), .Z(n26933) );
  XNOR U37407 ( .A(q[10]), .B(DB[1420]), .Z(n37087) );
  XNOR U37408 ( .A(q[9]), .B(DB[1419]), .Z(n26931) );
  IV U37409 ( .A(n26946), .Z(n37081) );
  XOR U37410 ( .A(n37088), .B(n37089), .Z(n26946) );
  XNOR U37411 ( .A(n26963), .B(n26944), .Z(n37089) );
  XNOR U37412 ( .A(q[0]), .B(DB[1410]), .Z(n26944) );
  XOR U37413 ( .A(n37090), .B(n26952), .Z(n26963) );
  XNOR U37414 ( .A(q[7]), .B(DB[1417]), .Z(n26952) );
  IV U37415 ( .A(n26951), .Z(n37090) );
  XNOR U37416 ( .A(n26949), .B(n37091), .Z(n26951) );
  XNOR U37417 ( .A(q[6]), .B(DB[1416]), .Z(n37091) );
  XNOR U37418 ( .A(q[5]), .B(DB[1415]), .Z(n26949) );
  IV U37419 ( .A(n26962), .Z(n37088) );
  XOR U37420 ( .A(n37092), .B(n37093), .Z(n26962) );
  XNOR U37421 ( .A(n26958), .B(n26960), .Z(n37093) );
  XNOR U37422 ( .A(q[1]), .B(DB[1411]), .Z(n26960) );
  XNOR U37423 ( .A(q[4]), .B(DB[1414]), .Z(n26958) );
  IV U37424 ( .A(n26957), .Z(n37092) );
  XNOR U37425 ( .A(n26955), .B(n37094), .Z(n26957) );
  XNOR U37426 ( .A(q[3]), .B(DB[1413]), .Z(n37094) );
  XNOR U37427 ( .A(q[2]), .B(DB[1412]), .Z(n26955) );
  XOR U37428 ( .A(n37095), .B(n26853), .Z(n26781) );
  XOR U37429 ( .A(n37096), .B(n26845), .Z(n26853) );
  XOR U37430 ( .A(n37097), .B(n26834), .Z(n26845) );
  XNOR U37431 ( .A(q[14]), .B(DB[1439]), .Z(n26834) );
  IV U37432 ( .A(n26833), .Z(n37097) );
  XNOR U37433 ( .A(n26831), .B(n37098), .Z(n26833) );
  XNOR U37434 ( .A(q[13]), .B(DB[1438]), .Z(n37098) );
  XNOR U37435 ( .A(q[12]), .B(DB[1437]), .Z(n26831) );
  IV U37436 ( .A(n26844), .Z(n37096) );
  XOR U37437 ( .A(n37099), .B(n37100), .Z(n26844) );
  XNOR U37438 ( .A(n26840), .B(n26842), .Z(n37100) );
  XNOR U37439 ( .A(q[8]), .B(DB[1433]), .Z(n26842) );
  XNOR U37440 ( .A(q[11]), .B(DB[1436]), .Z(n26840) );
  IV U37441 ( .A(n26839), .Z(n37099) );
  XNOR U37442 ( .A(n26837), .B(n37101), .Z(n26839) );
  XNOR U37443 ( .A(q[10]), .B(DB[1435]), .Z(n37101) );
  XNOR U37444 ( .A(q[9]), .B(DB[1434]), .Z(n26837) );
  IV U37445 ( .A(n26852), .Z(n37095) );
  XOR U37446 ( .A(n37102), .B(n37103), .Z(n26852) );
  XNOR U37447 ( .A(n26869), .B(n26850), .Z(n37103) );
  XNOR U37448 ( .A(q[0]), .B(DB[1425]), .Z(n26850) );
  XOR U37449 ( .A(n37104), .B(n26858), .Z(n26869) );
  XNOR U37450 ( .A(q[7]), .B(DB[1432]), .Z(n26858) );
  IV U37451 ( .A(n26857), .Z(n37104) );
  XNOR U37452 ( .A(n26855), .B(n37105), .Z(n26857) );
  XNOR U37453 ( .A(q[6]), .B(DB[1431]), .Z(n37105) );
  XNOR U37454 ( .A(q[5]), .B(DB[1430]), .Z(n26855) );
  IV U37455 ( .A(n26868), .Z(n37102) );
  XOR U37456 ( .A(n37106), .B(n37107), .Z(n26868) );
  XNOR U37457 ( .A(n26864), .B(n26866), .Z(n37107) );
  XNOR U37458 ( .A(q[1]), .B(DB[1426]), .Z(n26866) );
  XNOR U37459 ( .A(q[4]), .B(DB[1429]), .Z(n26864) );
  IV U37460 ( .A(n26863), .Z(n37106) );
  XNOR U37461 ( .A(n26861), .B(n37108), .Z(n26863) );
  XNOR U37462 ( .A(q[3]), .B(DB[1428]), .Z(n37108) );
  XNOR U37463 ( .A(q[2]), .B(DB[1427]), .Z(n26861) );
  XOR U37464 ( .A(n37109), .B(n26759), .Z(n26687) );
  XOR U37465 ( .A(n37110), .B(n26751), .Z(n26759) );
  XOR U37466 ( .A(n37111), .B(n26740), .Z(n26751) );
  XNOR U37467 ( .A(q[14]), .B(DB[1454]), .Z(n26740) );
  IV U37468 ( .A(n26739), .Z(n37111) );
  XNOR U37469 ( .A(n26737), .B(n37112), .Z(n26739) );
  XNOR U37470 ( .A(q[13]), .B(DB[1453]), .Z(n37112) );
  XNOR U37471 ( .A(q[12]), .B(DB[1452]), .Z(n26737) );
  IV U37472 ( .A(n26750), .Z(n37110) );
  XOR U37473 ( .A(n37113), .B(n37114), .Z(n26750) );
  XNOR U37474 ( .A(n26746), .B(n26748), .Z(n37114) );
  XNOR U37475 ( .A(q[8]), .B(DB[1448]), .Z(n26748) );
  XNOR U37476 ( .A(q[11]), .B(DB[1451]), .Z(n26746) );
  IV U37477 ( .A(n26745), .Z(n37113) );
  XNOR U37478 ( .A(n26743), .B(n37115), .Z(n26745) );
  XNOR U37479 ( .A(q[10]), .B(DB[1450]), .Z(n37115) );
  XNOR U37480 ( .A(q[9]), .B(DB[1449]), .Z(n26743) );
  IV U37481 ( .A(n26758), .Z(n37109) );
  XOR U37482 ( .A(n37116), .B(n37117), .Z(n26758) );
  XNOR U37483 ( .A(n26775), .B(n26756), .Z(n37117) );
  XNOR U37484 ( .A(q[0]), .B(DB[1440]), .Z(n26756) );
  XOR U37485 ( .A(n37118), .B(n26764), .Z(n26775) );
  XNOR U37486 ( .A(q[7]), .B(DB[1447]), .Z(n26764) );
  IV U37487 ( .A(n26763), .Z(n37118) );
  XNOR U37488 ( .A(n26761), .B(n37119), .Z(n26763) );
  XNOR U37489 ( .A(q[6]), .B(DB[1446]), .Z(n37119) );
  XNOR U37490 ( .A(q[5]), .B(DB[1445]), .Z(n26761) );
  IV U37491 ( .A(n26774), .Z(n37116) );
  XOR U37492 ( .A(n37120), .B(n37121), .Z(n26774) );
  XNOR U37493 ( .A(n26770), .B(n26772), .Z(n37121) );
  XNOR U37494 ( .A(q[1]), .B(DB[1441]), .Z(n26772) );
  XNOR U37495 ( .A(q[4]), .B(DB[1444]), .Z(n26770) );
  IV U37496 ( .A(n26769), .Z(n37120) );
  XNOR U37497 ( .A(n26767), .B(n37122), .Z(n26769) );
  XNOR U37498 ( .A(q[3]), .B(DB[1443]), .Z(n37122) );
  XNOR U37499 ( .A(q[2]), .B(DB[1442]), .Z(n26767) );
  XOR U37500 ( .A(n37123), .B(n26665), .Z(n26593) );
  XOR U37501 ( .A(n37124), .B(n26657), .Z(n26665) );
  XOR U37502 ( .A(n37125), .B(n26646), .Z(n26657) );
  XNOR U37503 ( .A(q[14]), .B(DB[1469]), .Z(n26646) );
  IV U37504 ( .A(n26645), .Z(n37125) );
  XNOR U37505 ( .A(n26643), .B(n37126), .Z(n26645) );
  XNOR U37506 ( .A(q[13]), .B(DB[1468]), .Z(n37126) );
  XNOR U37507 ( .A(q[12]), .B(DB[1467]), .Z(n26643) );
  IV U37508 ( .A(n26656), .Z(n37124) );
  XOR U37509 ( .A(n37127), .B(n37128), .Z(n26656) );
  XNOR U37510 ( .A(n26652), .B(n26654), .Z(n37128) );
  XNOR U37511 ( .A(q[8]), .B(DB[1463]), .Z(n26654) );
  XNOR U37512 ( .A(q[11]), .B(DB[1466]), .Z(n26652) );
  IV U37513 ( .A(n26651), .Z(n37127) );
  XNOR U37514 ( .A(n26649), .B(n37129), .Z(n26651) );
  XNOR U37515 ( .A(q[10]), .B(DB[1465]), .Z(n37129) );
  XNOR U37516 ( .A(q[9]), .B(DB[1464]), .Z(n26649) );
  IV U37517 ( .A(n26664), .Z(n37123) );
  XOR U37518 ( .A(n37130), .B(n37131), .Z(n26664) );
  XNOR U37519 ( .A(n26681), .B(n26662), .Z(n37131) );
  XNOR U37520 ( .A(q[0]), .B(DB[1455]), .Z(n26662) );
  XOR U37521 ( .A(n37132), .B(n26670), .Z(n26681) );
  XNOR U37522 ( .A(q[7]), .B(DB[1462]), .Z(n26670) );
  IV U37523 ( .A(n26669), .Z(n37132) );
  XNOR U37524 ( .A(n26667), .B(n37133), .Z(n26669) );
  XNOR U37525 ( .A(q[6]), .B(DB[1461]), .Z(n37133) );
  XNOR U37526 ( .A(q[5]), .B(DB[1460]), .Z(n26667) );
  IV U37527 ( .A(n26680), .Z(n37130) );
  XOR U37528 ( .A(n37134), .B(n37135), .Z(n26680) );
  XNOR U37529 ( .A(n26676), .B(n26678), .Z(n37135) );
  XNOR U37530 ( .A(q[1]), .B(DB[1456]), .Z(n26678) );
  XNOR U37531 ( .A(q[4]), .B(DB[1459]), .Z(n26676) );
  IV U37532 ( .A(n26675), .Z(n37134) );
  XNOR U37533 ( .A(n26673), .B(n37136), .Z(n26675) );
  XNOR U37534 ( .A(q[3]), .B(DB[1458]), .Z(n37136) );
  XNOR U37535 ( .A(q[2]), .B(DB[1457]), .Z(n26673) );
  XOR U37536 ( .A(n37137), .B(n26571), .Z(n26499) );
  XOR U37537 ( .A(n37138), .B(n26563), .Z(n26571) );
  XOR U37538 ( .A(n37139), .B(n26552), .Z(n26563) );
  XNOR U37539 ( .A(q[14]), .B(DB[1484]), .Z(n26552) );
  IV U37540 ( .A(n26551), .Z(n37139) );
  XNOR U37541 ( .A(n26549), .B(n37140), .Z(n26551) );
  XNOR U37542 ( .A(q[13]), .B(DB[1483]), .Z(n37140) );
  XNOR U37543 ( .A(q[12]), .B(DB[1482]), .Z(n26549) );
  IV U37544 ( .A(n26562), .Z(n37138) );
  XOR U37545 ( .A(n37141), .B(n37142), .Z(n26562) );
  XNOR U37546 ( .A(n26558), .B(n26560), .Z(n37142) );
  XNOR U37547 ( .A(q[8]), .B(DB[1478]), .Z(n26560) );
  XNOR U37548 ( .A(q[11]), .B(DB[1481]), .Z(n26558) );
  IV U37549 ( .A(n26557), .Z(n37141) );
  XNOR U37550 ( .A(n26555), .B(n37143), .Z(n26557) );
  XNOR U37551 ( .A(q[10]), .B(DB[1480]), .Z(n37143) );
  XNOR U37552 ( .A(q[9]), .B(DB[1479]), .Z(n26555) );
  IV U37553 ( .A(n26570), .Z(n37137) );
  XOR U37554 ( .A(n37144), .B(n37145), .Z(n26570) );
  XNOR U37555 ( .A(n26587), .B(n26568), .Z(n37145) );
  XNOR U37556 ( .A(q[0]), .B(DB[1470]), .Z(n26568) );
  XOR U37557 ( .A(n37146), .B(n26576), .Z(n26587) );
  XNOR U37558 ( .A(q[7]), .B(DB[1477]), .Z(n26576) );
  IV U37559 ( .A(n26575), .Z(n37146) );
  XNOR U37560 ( .A(n26573), .B(n37147), .Z(n26575) );
  XNOR U37561 ( .A(q[6]), .B(DB[1476]), .Z(n37147) );
  XNOR U37562 ( .A(q[5]), .B(DB[1475]), .Z(n26573) );
  IV U37563 ( .A(n26586), .Z(n37144) );
  XOR U37564 ( .A(n37148), .B(n37149), .Z(n26586) );
  XNOR U37565 ( .A(n26582), .B(n26584), .Z(n37149) );
  XNOR U37566 ( .A(q[1]), .B(DB[1471]), .Z(n26584) );
  XNOR U37567 ( .A(q[4]), .B(DB[1474]), .Z(n26582) );
  IV U37568 ( .A(n26581), .Z(n37148) );
  XNOR U37569 ( .A(n26579), .B(n37150), .Z(n26581) );
  XNOR U37570 ( .A(q[3]), .B(DB[1473]), .Z(n37150) );
  XNOR U37571 ( .A(q[2]), .B(DB[1472]), .Z(n26579) );
  XOR U37572 ( .A(n37151), .B(n26477), .Z(n26405) );
  XOR U37573 ( .A(n37152), .B(n26469), .Z(n26477) );
  XOR U37574 ( .A(n37153), .B(n26458), .Z(n26469) );
  XNOR U37575 ( .A(q[14]), .B(DB[1499]), .Z(n26458) );
  IV U37576 ( .A(n26457), .Z(n37153) );
  XNOR U37577 ( .A(n26455), .B(n37154), .Z(n26457) );
  XNOR U37578 ( .A(q[13]), .B(DB[1498]), .Z(n37154) );
  XNOR U37579 ( .A(q[12]), .B(DB[1497]), .Z(n26455) );
  IV U37580 ( .A(n26468), .Z(n37152) );
  XOR U37581 ( .A(n37155), .B(n37156), .Z(n26468) );
  XNOR U37582 ( .A(n26464), .B(n26466), .Z(n37156) );
  XNOR U37583 ( .A(q[8]), .B(DB[1493]), .Z(n26466) );
  XNOR U37584 ( .A(q[11]), .B(DB[1496]), .Z(n26464) );
  IV U37585 ( .A(n26463), .Z(n37155) );
  XNOR U37586 ( .A(n26461), .B(n37157), .Z(n26463) );
  XNOR U37587 ( .A(q[10]), .B(DB[1495]), .Z(n37157) );
  XNOR U37588 ( .A(q[9]), .B(DB[1494]), .Z(n26461) );
  IV U37589 ( .A(n26476), .Z(n37151) );
  XOR U37590 ( .A(n37158), .B(n37159), .Z(n26476) );
  XNOR U37591 ( .A(n26493), .B(n26474), .Z(n37159) );
  XNOR U37592 ( .A(q[0]), .B(DB[1485]), .Z(n26474) );
  XOR U37593 ( .A(n37160), .B(n26482), .Z(n26493) );
  XNOR U37594 ( .A(q[7]), .B(DB[1492]), .Z(n26482) );
  IV U37595 ( .A(n26481), .Z(n37160) );
  XNOR U37596 ( .A(n26479), .B(n37161), .Z(n26481) );
  XNOR U37597 ( .A(q[6]), .B(DB[1491]), .Z(n37161) );
  XNOR U37598 ( .A(q[5]), .B(DB[1490]), .Z(n26479) );
  IV U37599 ( .A(n26492), .Z(n37158) );
  XOR U37600 ( .A(n37162), .B(n37163), .Z(n26492) );
  XNOR U37601 ( .A(n26488), .B(n26490), .Z(n37163) );
  XNOR U37602 ( .A(q[1]), .B(DB[1486]), .Z(n26490) );
  XNOR U37603 ( .A(q[4]), .B(DB[1489]), .Z(n26488) );
  IV U37604 ( .A(n26487), .Z(n37162) );
  XNOR U37605 ( .A(n26485), .B(n37164), .Z(n26487) );
  XNOR U37606 ( .A(q[3]), .B(DB[1488]), .Z(n37164) );
  XNOR U37607 ( .A(q[2]), .B(DB[1487]), .Z(n26485) );
  XOR U37608 ( .A(n37165), .B(n26383), .Z(n26311) );
  XOR U37609 ( .A(n37166), .B(n26375), .Z(n26383) );
  XOR U37610 ( .A(n37167), .B(n26364), .Z(n26375) );
  XNOR U37611 ( .A(q[14]), .B(DB[1514]), .Z(n26364) );
  IV U37612 ( .A(n26363), .Z(n37167) );
  XNOR U37613 ( .A(n26361), .B(n37168), .Z(n26363) );
  XNOR U37614 ( .A(q[13]), .B(DB[1513]), .Z(n37168) );
  XNOR U37615 ( .A(q[12]), .B(DB[1512]), .Z(n26361) );
  IV U37616 ( .A(n26374), .Z(n37166) );
  XOR U37617 ( .A(n37169), .B(n37170), .Z(n26374) );
  XNOR U37618 ( .A(n26370), .B(n26372), .Z(n37170) );
  XNOR U37619 ( .A(q[8]), .B(DB[1508]), .Z(n26372) );
  XNOR U37620 ( .A(q[11]), .B(DB[1511]), .Z(n26370) );
  IV U37621 ( .A(n26369), .Z(n37169) );
  XNOR U37622 ( .A(n26367), .B(n37171), .Z(n26369) );
  XNOR U37623 ( .A(q[10]), .B(DB[1510]), .Z(n37171) );
  XNOR U37624 ( .A(q[9]), .B(DB[1509]), .Z(n26367) );
  IV U37625 ( .A(n26382), .Z(n37165) );
  XOR U37626 ( .A(n37172), .B(n37173), .Z(n26382) );
  XNOR U37627 ( .A(n26399), .B(n26380), .Z(n37173) );
  XNOR U37628 ( .A(q[0]), .B(DB[1500]), .Z(n26380) );
  XOR U37629 ( .A(n37174), .B(n26388), .Z(n26399) );
  XNOR U37630 ( .A(q[7]), .B(DB[1507]), .Z(n26388) );
  IV U37631 ( .A(n26387), .Z(n37174) );
  XNOR U37632 ( .A(n26385), .B(n37175), .Z(n26387) );
  XNOR U37633 ( .A(q[6]), .B(DB[1506]), .Z(n37175) );
  XNOR U37634 ( .A(q[5]), .B(DB[1505]), .Z(n26385) );
  IV U37635 ( .A(n26398), .Z(n37172) );
  XOR U37636 ( .A(n37176), .B(n37177), .Z(n26398) );
  XNOR U37637 ( .A(n26394), .B(n26396), .Z(n37177) );
  XNOR U37638 ( .A(q[1]), .B(DB[1501]), .Z(n26396) );
  XNOR U37639 ( .A(q[4]), .B(DB[1504]), .Z(n26394) );
  IV U37640 ( .A(n26393), .Z(n37176) );
  XNOR U37641 ( .A(n26391), .B(n37178), .Z(n26393) );
  XNOR U37642 ( .A(q[3]), .B(DB[1503]), .Z(n37178) );
  XNOR U37643 ( .A(q[2]), .B(DB[1502]), .Z(n26391) );
  XOR U37644 ( .A(n37179), .B(n26289), .Z(n26217) );
  XOR U37645 ( .A(n37180), .B(n26281), .Z(n26289) );
  XOR U37646 ( .A(n37181), .B(n26270), .Z(n26281) );
  XNOR U37647 ( .A(q[14]), .B(DB[1529]), .Z(n26270) );
  IV U37648 ( .A(n26269), .Z(n37181) );
  XNOR U37649 ( .A(n26267), .B(n37182), .Z(n26269) );
  XNOR U37650 ( .A(q[13]), .B(DB[1528]), .Z(n37182) );
  XNOR U37651 ( .A(q[12]), .B(DB[1527]), .Z(n26267) );
  IV U37652 ( .A(n26280), .Z(n37180) );
  XOR U37653 ( .A(n37183), .B(n37184), .Z(n26280) );
  XNOR U37654 ( .A(n26276), .B(n26278), .Z(n37184) );
  XNOR U37655 ( .A(q[8]), .B(DB[1523]), .Z(n26278) );
  XNOR U37656 ( .A(q[11]), .B(DB[1526]), .Z(n26276) );
  IV U37657 ( .A(n26275), .Z(n37183) );
  XNOR U37658 ( .A(n26273), .B(n37185), .Z(n26275) );
  XNOR U37659 ( .A(q[10]), .B(DB[1525]), .Z(n37185) );
  XNOR U37660 ( .A(q[9]), .B(DB[1524]), .Z(n26273) );
  IV U37661 ( .A(n26288), .Z(n37179) );
  XOR U37662 ( .A(n37186), .B(n37187), .Z(n26288) );
  XNOR U37663 ( .A(n26305), .B(n26286), .Z(n37187) );
  XNOR U37664 ( .A(q[0]), .B(DB[1515]), .Z(n26286) );
  XOR U37665 ( .A(n37188), .B(n26294), .Z(n26305) );
  XNOR U37666 ( .A(q[7]), .B(DB[1522]), .Z(n26294) );
  IV U37667 ( .A(n26293), .Z(n37188) );
  XNOR U37668 ( .A(n26291), .B(n37189), .Z(n26293) );
  XNOR U37669 ( .A(q[6]), .B(DB[1521]), .Z(n37189) );
  XNOR U37670 ( .A(q[5]), .B(DB[1520]), .Z(n26291) );
  IV U37671 ( .A(n26304), .Z(n37186) );
  XOR U37672 ( .A(n37190), .B(n37191), .Z(n26304) );
  XNOR U37673 ( .A(n26300), .B(n26302), .Z(n37191) );
  XNOR U37674 ( .A(q[1]), .B(DB[1516]), .Z(n26302) );
  XNOR U37675 ( .A(q[4]), .B(DB[1519]), .Z(n26300) );
  IV U37676 ( .A(n26299), .Z(n37190) );
  XNOR U37677 ( .A(n26297), .B(n37192), .Z(n26299) );
  XNOR U37678 ( .A(q[3]), .B(DB[1518]), .Z(n37192) );
  XNOR U37679 ( .A(q[2]), .B(DB[1517]), .Z(n26297) );
  XOR U37680 ( .A(n37193), .B(n26195), .Z(n26123) );
  XOR U37681 ( .A(n37194), .B(n26187), .Z(n26195) );
  XOR U37682 ( .A(n37195), .B(n26176), .Z(n26187) );
  XNOR U37683 ( .A(q[14]), .B(DB[1544]), .Z(n26176) );
  IV U37684 ( .A(n26175), .Z(n37195) );
  XNOR U37685 ( .A(n26173), .B(n37196), .Z(n26175) );
  XNOR U37686 ( .A(q[13]), .B(DB[1543]), .Z(n37196) );
  XNOR U37687 ( .A(q[12]), .B(DB[1542]), .Z(n26173) );
  IV U37688 ( .A(n26186), .Z(n37194) );
  XOR U37689 ( .A(n37197), .B(n37198), .Z(n26186) );
  XNOR U37690 ( .A(n26182), .B(n26184), .Z(n37198) );
  XNOR U37691 ( .A(q[8]), .B(DB[1538]), .Z(n26184) );
  XNOR U37692 ( .A(q[11]), .B(DB[1541]), .Z(n26182) );
  IV U37693 ( .A(n26181), .Z(n37197) );
  XNOR U37694 ( .A(n26179), .B(n37199), .Z(n26181) );
  XNOR U37695 ( .A(q[10]), .B(DB[1540]), .Z(n37199) );
  XNOR U37696 ( .A(q[9]), .B(DB[1539]), .Z(n26179) );
  IV U37697 ( .A(n26194), .Z(n37193) );
  XOR U37698 ( .A(n37200), .B(n37201), .Z(n26194) );
  XNOR U37699 ( .A(n26211), .B(n26192), .Z(n37201) );
  XNOR U37700 ( .A(q[0]), .B(DB[1530]), .Z(n26192) );
  XOR U37701 ( .A(n37202), .B(n26200), .Z(n26211) );
  XNOR U37702 ( .A(q[7]), .B(DB[1537]), .Z(n26200) );
  IV U37703 ( .A(n26199), .Z(n37202) );
  XNOR U37704 ( .A(n26197), .B(n37203), .Z(n26199) );
  XNOR U37705 ( .A(q[6]), .B(DB[1536]), .Z(n37203) );
  XNOR U37706 ( .A(q[5]), .B(DB[1535]), .Z(n26197) );
  IV U37707 ( .A(n26210), .Z(n37200) );
  XOR U37708 ( .A(n37204), .B(n37205), .Z(n26210) );
  XNOR U37709 ( .A(n26206), .B(n26208), .Z(n37205) );
  XNOR U37710 ( .A(q[1]), .B(DB[1531]), .Z(n26208) );
  XNOR U37711 ( .A(q[4]), .B(DB[1534]), .Z(n26206) );
  IV U37712 ( .A(n26205), .Z(n37204) );
  XNOR U37713 ( .A(n26203), .B(n37206), .Z(n26205) );
  XNOR U37714 ( .A(q[3]), .B(DB[1533]), .Z(n37206) );
  XNOR U37715 ( .A(q[2]), .B(DB[1532]), .Z(n26203) );
  XOR U37716 ( .A(n37207), .B(n26101), .Z(n26029) );
  XOR U37717 ( .A(n37208), .B(n26093), .Z(n26101) );
  XOR U37718 ( .A(n37209), .B(n26082), .Z(n26093) );
  XNOR U37719 ( .A(q[14]), .B(DB[1559]), .Z(n26082) );
  IV U37720 ( .A(n26081), .Z(n37209) );
  XNOR U37721 ( .A(n26079), .B(n37210), .Z(n26081) );
  XNOR U37722 ( .A(q[13]), .B(DB[1558]), .Z(n37210) );
  XNOR U37723 ( .A(q[12]), .B(DB[1557]), .Z(n26079) );
  IV U37724 ( .A(n26092), .Z(n37208) );
  XOR U37725 ( .A(n37211), .B(n37212), .Z(n26092) );
  XNOR U37726 ( .A(n26088), .B(n26090), .Z(n37212) );
  XNOR U37727 ( .A(q[8]), .B(DB[1553]), .Z(n26090) );
  XNOR U37728 ( .A(q[11]), .B(DB[1556]), .Z(n26088) );
  IV U37729 ( .A(n26087), .Z(n37211) );
  XNOR U37730 ( .A(n26085), .B(n37213), .Z(n26087) );
  XNOR U37731 ( .A(q[10]), .B(DB[1555]), .Z(n37213) );
  XNOR U37732 ( .A(q[9]), .B(DB[1554]), .Z(n26085) );
  IV U37733 ( .A(n26100), .Z(n37207) );
  XOR U37734 ( .A(n37214), .B(n37215), .Z(n26100) );
  XNOR U37735 ( .A(n26117), .B(n26098), .Z(n37215) );
  XNOR U37736 ( .A(q[0]), .B(DB[1545]), .Z(n26098) );
  XOR U37737 ( .A(n37216), .B(n26106), .Z(n26117) );
  XNOR U37738 ( .A(q[7]), .B(DB[1552]), .Z(n26106) );
  IV U37739 ( .A(n26105), .Z(n37216) );
  XNOR U37740 ( .A(n26103), .B(n37217), .Z(n26105) );
  XNOR U37741 ( .A(q[6]), .B(DB[1551]), .Z(n37217) );
  XNOR U37742 ( .A(q[5]), .B(DB[1550]), .Z(n26103) );
  IV U37743 ( .A(n26116), .Z(n37214) );
  XOR U37744 ( .A(n37218), .B(n37219), .Z(n26116) );
  XNOR U37745 ( .A(n26112), .B(n26114), .Z(n37219) );
  XNOR U37746 ( .A(q[1]), .B(DB[1546]), .Z(n26114) );
  XNOR U37747 ( .A(q[4]), .B(DB[1549]), .Z(n26112) );
  IV U37748 ( .A(n26111), .Z(n37218) );
  XNOR U37749 ( .A(n26109), .B(n37220), .Z(n26111) );
  XNOR U37750 ( .A(q[3]), .B(DB[1548]), .Z(n37220) );
  XNOR U37751 ( .A(q[2]), .B(DB[1547]), .Z(n26109) );
  XOR U37752 ( .A(n37221), .B(n26007), .Z(n25935) );
  XOR U37753 ( .A(n37222), .B(n25999), .Z(n26007) );
  XOR U37754 ( .A(n37223), .B(n25988), .Z(n25999) );
  XNOR U37755 ( .A(q[14]), .B(DB[1574]), .Z(n25988) );
  IV U37756 ( .A(n25987), .Z(n37223) );
  XNOR U37757 ( .A(n25985), .B(n37224), .Z(n25987) );
  XNOR U37758 ( .A(q[13]), .B(DB[1573]), .Z(n37224) );
  XNOR U37759 ( .A(q[12]), .B(DB[1572]), .Z(n25985) );
  IV U37760 ( .A(n25998), .Z(n37222) );
  XOR U37761 ( .A(n37225), .B(n37226), .Z(n25998) );
  XNOR U37762 ( .A(n25994), .B(n25996), .Z(n37226) );
  XNOR U37763 ( .A(q[8]), .B(DB[1568]), .Z(n25996) );
  XNOR U37764 ( .A(q[11]), .B(DB[1571]), .Z(n25994) );
  IV U37765 ( .A(n25993), .Z(n37225) );
  XNOR U37766 ( .A(n25991), .B(n37227), .Z(n25993) );
  XNOR U37767 ( .A(q[10]), .B(DB[1570]), .Z(n37227) );
  XNOR U37768 ( .A(q[9]), .B(DB[1569]), .Z(n25991) );
  IV U37769 ( .A(n26006), .Z(n37221) );
  XOR U37770 ( .A(n37228), .B(n37229), .Z(n26006) );
  XNOR U37771 ( .A(n26023), .B(n26004), .Z(n37229) );
  XNOR U37772 ( .A(q[0]), .B(DB[1560]), .Z(n26004) );
  XOR U37773 ( .A(n37230), .B(n26012), .Z(n26023) );
  XNOR U37774 ( .A(q[7]), .B(DB[1567]), .Z(n26012) );
  IV U37775 ( .A(n26011), .Z(n37230) );
  XNOR U37776 ( .A(n26009), .B(n37231), .Z(n26011) );
  XNOR U37777 ( .A(q[6]), .B(DB[1566]), .Z(n37231) );
  XNOR U37778 ( .A(q[5]), .B(DB[1565]), .Z(n26009) );
  IV U37779 ( .A(n26022), .Z(n37228) );
  XOR U37780 ( .A(n37232), .B(n37233), .Z(n26022) );
  XNOR U37781 ( .A(n26018), .B(n26020), .Z(n37233) );
  XNOR U37782 ( .A(q[1]), .B(DB[1561]), .Z(n26020) );
  XNOR U37783 ( .A(q[4]), .B(DB[1564]), .Z(n26018) );
  IV U37784 ( .A(n26017), .Z(n37232) );
  XNOR U37785 ( .A(n26015), .B(n37234), .Z(n26017) );
  XNOR U37786 ( .A(q[3]), .B(DB[1563]), .Z(n37234) );
  XNOR U37787 ( .A(q[2]), .B(DB[1562]), .Z(n26015) );
  XOR U37788 ( .A(n37235), .B(n25913), .Z(n25841) );
  XOR U37789 ( .A(n37236), .B(n25905), .Z(n25913) );
  XOR U37790 ( .A(n37237), .B(n25894), .Z(n25905) );
  XNOR U37791 ( .A(q[14]), .B(DB[1589]), .Z(n25894) );
  IV U37792 ( .A(n25893), .Z(n37237) );
  XNOR U37793 ( .A(n25891), .B(n37238), .Z(n25893) );
  XNOR U37794 ( .A(q[13]), .B(DB[1588]), .Z(n37238) );
  XNOR U37795 ( .A(q[12]), .B(DB[1587]), .Z(n25891) );
  IV U37796 ( .A(n25904), .Z(n37236) );
  XOR U37797 ( .A(n37239), .B(n37240), .Z(n25904) );
  XNOR U37798 ( .A(n25900), .B(n25902), .Z(n37240) );
  XNOR U37799 ( .A(q[8]), .B(DB[1583]), .Z(n25902) );
  XNOR U37800 ( .A(q[11]), .B(DB[1586]), .Z(n25900) );
  IV U37801 ( .A(n25899), .Z(n37239) );
  XNOR U37802 ( .A(n25897), .B(n37241), .Z(n25899) );
  XNOR U37803 ( .A(q[10]), .B(DB[1585]), .Z(n37241) );
  XNOR U37804 ( .A(q[9]), .B(DB[1584]), .Z(n25897) );
  IV U37805 ( .A(n25912), .Z(n37235) );
  XOR U37806 ( .A(n37242), .B(n37243), .Z(n25912) );
  XNOR U37807 ( .A(n25929), .B(n25910), .Z(n37243) );
  XNOR U37808 ( .A(q[0]), .B(DB[1575]), .Z(n25910) );
  XOR U37809 ( .A(n37244), .B(n25918), .Z(n25929) );
  XNOR U37810 ( .A(q[7]), .B(DB[1582]), .Z(n25918) );
  IV U37811 ( .A(n25917), .Z(n37244) );
  XNOR U37812 ( .A(n25915), .B(n37245), .Z(n25917) );
  XNOR U37813 ( .A(q[6]), .B(DB[1581]), .Z(n37245) );
  XNOR U37814 ( .A(q[5]), .B(DB[1580]), .Z(n25915) );
  IV U37815 ( .A(n25928), .Z(n37242) );
  XOR U37816 ( .A(n37246), .B(n37247), .Z(n25928) );
  XNOR U37817 ( .A(n25924), .B(n25926), .Z(n37247) );
  XNOR U37818 ( .A(q[1]), .B(DB[1576]), .Z(n25926) );
  XNOR U37819 ( .A(q[4]), .B(DB[1579]), .Z(n25924) );
  IV U37820 ( .A(n25923), .Z(n37246) );
  XNOR U37821 ( .A(n25921), .B(n37248), .Z(n25923) );
  XNOR U37822 ( .A(q[3]), .B(DB[1578]), .Z(n37248) );
  XNOR U37823 ( .A(q[2]), .B(DB[1577]), .Z(n25921) );
  XOR U37824 ( .A(n37249), .B(n25819), .Z(n25747) );
  XOR U37825 ( .A(n37250), .B(n25811), .Z(n25819) );
  XOR U37826 ( .A(n37251), .B(n25800), .Z(n25811) );
  XNOR U37827 ( .A(q[14]), .B(DB[1604]), .Z(n25800) );
  IV U37828 ( .A(n25799), .Z(n37251) );
  XNOR U37829 ( .A(n25797), .B(n37252), .Z(n25799) );
  XNOR U37830 ( .A(q[13]), .B(DB[1603]), .Z(n37252) );
  XNOR U37831 ( .A(q[12]), .B(DB[1602]), .Z(n25797) );
  IV U37832 ( .A(n25810), .Z(n37250) );
  XOR U37833 ( .A(n37253), .B(n37254), .Z(n25810) );
  XNOR U37834 ( .A(n25806), .B(n25808), .Z(n37254) );
  XNOR U37835 ( .A(q[8]), .B(DB[1598]), .Z(n25808) );
  XNOR U37836 ( .A(q[11]), .B(DB[1601]), .Z(n25806) );
  IV U37837 ( .A(n25805), .Z(n37253) );
  XNOR U37838 ( .A(n25803), .B(n37255), .Z(n25805) );
  XNOR U37839 ( .A(q[10]), .B(DB[1600]), .Z(n37255) );
  XNOR U37840 ( .A(q[9]), .B(DB[1599]), .Z(n25803) );
  IV U37841 ( .A(n25818), .Z(n37249) );
  XOR U37842 ( .A(n37256), .B(n37257), .Z(n25818) );
  XNOR U37843 ( .A(n25835), .B(n25816), .Z(n37257) );
  XNOR U37844 ( .A(q[0]), .B(DB[1590]), .Z(n25816) );
  XOR U37845 ( .A(n37258), .B(n25824), .Z(n25835) );
  XNOR U37846 ( .A(q[7]), .B(DB[1597]), .Z(n25824) );
  IV U37847 ( .A(n25823), .Z(n37258) );
  XNOR U37848 ( .A(n25821), .B(n37259), .Z(n25823) );
  XNOR U37849 ( .A(q[6]), .B(DB[1596]), .Z(n37259) );
  XNOR U37850 ( .A(q[5]), .B(DB[1595]), .Z(n25821) );
  IV U37851 ( .A(n25834), .Z(n37256) );
  XOR U37852 ( .A(n37260), .B(n37261), .Z(n25834) );
  XNOR U37853 ( .A(n25830), .B(n25832), .Z(n37261) );
  XNOR U37854 ( .A(q[1]), .B(DB[1591]), .Z(n25832) );
  XNOR U37855 ( .A(q[4]), .B(DB[1594]), .Z(n25830) );
  IV U37856 ( .A(n25829), .Z(n37260) );
  XNOR U37857 ( .A(n25827), .B(n37262), .Z(n25829) );
  XNOR U37858 ( .A(q[3]), .B(DB[1593]), .Z(n37262) );
  XNOR U37859 ( .A(q[2]), .B(DB[1592]), .Z(n25827) );
  XOR U37860 ( .A(n37263), .B(n25725), .Z(n25653) );
  XOR U37861 ( .A(n37264), .B(n25717), .Z(n25725) );
  XOR U37862 ( .A(n37265), .B(n25706), .Z(n25717) );
  XNOR U37863 ( .A(q[14]), .B(DB[1619]), .Z(n25706) );
  IV U37864 ( .A(n25705), .Z(n37265) );
  XNOR U37865 ( .A(n25703), .B(n37266), .Z(n25705) );
  XNOR U37866 ( .A(q[13]), .B(DB[1618]), .Z(n37266) );
  XNOR U37867 ( .A(q[12]), .B(DB[1617]), .Z(n25703) );
  IV U37868 ( .A(n25716), .Z(n37264) );
  XOR U37869 ( .A(n37267), .B(n37268), .Z(n25716) );
  XNOR U37870 ( .A(n25712), .B(n25714), .Z(n37268) );
  XNOR U37871 ( .A(q[8]), .B(DB[1613]), .Z(n25714) );
  XNOR U37872 ( .A(q[11]), .B(DB[1616]), .Z(n25712) );
  IV U37873 ( .A(n25711), .Z(n37267) );
  XNOR U37874 ( .A(n25709), .B(n37269), .Z(n25711) );
  XNOR U37875 ( .A(q[10]), .B(DB[1615]), .Z(n37269) );
  XNOR U37876 ( .A(q[9]), .B(DB[1614]), .Z(n25709) );
  IV U37877 ( .A(n25724), .Z(n37263) );
  XOR U37878 ( .A(n37270), .B(n37271), .Z(n25724) );
  XNOR U37879 ( .A(n25741), .B(n25722), .Z(n37271) );
  XNOR U37880 ( .A(q[0]), .B(DB[1605]), .Z(n25722) );
  XOR U37881 ( .A(n37272), .B(n25730), .Z(n25741) );
  XNOR U37882 ( .A(q[7]), .B(DB[1612]), .Z(n25730) );
  IV U37883 ( .A(n25729), .Z(n37272) );
  XNOR U37884 ( .A(n25727), .B(n37273), .Z(n25729) );
  XNOR U37885 ( .A(q[6]), .B(DB[1611]), .Z(n37273) );
  XNOR U37886 ( .A(q[5]), .B(DB[1610]), .Z(n25727) );
  IV U37887 ( .A(n25740), .Z(n37270) );
  XOR U37888 ( .A(n37274), .B(n37275), .Z(n25740) );
  XNOR U37889 ( .A(n25736), .B(n25738), .Z(n37275) );
  XNOR U37890 ( .A(q[1]), .B(DB[1606]), .Z(n25738) );
  XNOR U37891 ( .A(q[4]), .B(DB[1609]), .Z(n25736) );
  IV U37892 ( .A(n25735), .Z(n37274) );
  XNOR U37893 ( .A(n25733), .B(n37276), .Z(n25735) );
  XNOR U37894 ( .A(q[3]), .B(DB[1608]), .Z(n37276) );
  XNOR U37895 ( .A(q[2]), .B(DB[1607]), .Z(n25733) );
  XOR U37896 ( .A(n37277), .B(n25631), .Z(n25559) );
  XOR U37897 ( .A(n37278), .B(n25623), .Z(n25631) );
  XOR U37898 ( .A(n37279), .B(n25612), .Z(n25623) );
  XNOR U37899 ( .A(q[14]), .B(DB[1634]), .Z(n25612) );
  IV U37900 ( .A(n25611), .Z(n37279) );
  XNOR U37901 ( .A(n25609), .B(n37280), .Z(n25611) );
  XNOR U37902 ( .A(q[13]), .B(DB[1633]), .Z(n37280) );
  XNOR U37903 ( .A(q[12]), .B(DB[1632]), .Z(n25609) );
  IV U37904 ( .A(n25622), .Z(n37278) );
  XOR U37905 ( .A(n37281), .B(n37282), .Z(n25622) );
  XNOR U37906 ( .A(n25618), .B(n25620), .Z(n37282) );
  XNOR U37907 ( .A(q[8]), .B(DB[1628]), .Z(n25620) );
  XNOR U37908 ( .A(q[11]), .B(DB[1631]), .Z(n25618) );
  IV U37909 ( .A(n25617), .Z(n37281) );
  XNOR U37910 ( .A(n25615), .B(n37283), .Z(n25617) );
  XNOR U37911 ( .A(q[10]), .B(DB[1630]), .Z(n37283) );
  XNOR U37912 ( .A(q[9]), .B(DB[1629]), .Z(n25615) );
  IV U37913 ( .A(n25630), .Z(n37277) );
  XOR U37914 ( .A(n37284), .B(n37285), .Z(n25630) );
  XNOR U37915 ( .A(n25647), .B(n25628), .Z(n37285) );
  XNOR U37916 ( .A(q[0]), .B(DB[1620]), .Z(n25628) );
  XOR U37917 ( .A(n37286), .B(n25636), .Z(n25647) );
  XNOR U37918 ( .A(q[7]), .B(DB[1627]), .Z(n25636) );
  IV U37919 ( .A(n25635), .Z(n37286) );
  XNOR U37920 ( .A(n25633), .B(n37287), .Z(n25635) );
  XNOR U37921 ( .A(q[6]), .B(DB[1626]), .Z(n37287) );
  XNOR U37922 ( .A(q[5]), .B(DB[1625]), .Z(n25633) );
  IV U37923 ( .A(n25646), .Z(n37284) );
  XOR U37924 ( .A(n37288), .B(n37289), .Z(n25646) );
  XNOR U37925 ( .A(n25642), .B(n25644), .Z(n37289) );
  XNOR U37926 ( .A(q[1]), .B(DB[1621]), .Z(n25644) );
  XNOR U37927 ( .A(q[4]), .B(DB[1624]), .Z(n25642) );
  IV U37928 ( .A(n25641), .Z(n37288) );
  XNOR U37929 ( .A(n25639), .B(n37290), .Z(n25641) );
  XNOR U37930 ( .A(q[3]), .B(DB[1623]), .Z(n37290) );
  XNOR U37931 ( .A(q[2]), .B(DB[1622]), .Z(n25639) );
  XOR U37932 ( .A(n37291), .B(n25537), .Z(n25465) );
  XOR U37933 ( .A(n37292), .B(n25529), .Z(n25537) );
  XOR U37934 ( .A(n37293), .B(n25518), .Z(n25529) );
  XNOR U37935 ( .A(q[14]), .B(DB[1649]), .Z(n25518) );
  IV U37936 ( .A(n25517), .Z(n37293) );
  XNOR U37937 ( .A(n25515), .B(n37294), .Z(n25517) );
  XNOR U37938 ( .A(q[13]), .B(DB[1648]), .Z(n37294) );
  XNOR U37939 ( .A(q[12]), .B(DB[1647]), .Z(n25515) );
  IV U37940 ( .A(n25528), .Z(n37292) );
  XOR U37941 ( .A(n37295), .B(n37296), .Z(n25528) );
  XNOR U37942 ( .A(n25524), .B(n25526), .Z(n37296) );
  XNOR U37943 ( .A(q[8]), .B(DB[1643]), .Z(n25526) );
  XNOR U37944 ( .A(q[11]), .B(DB[1646]), .Z(n25524) );
  IV U37945 ( .A(n25523), .Z(n37295) );
  XNOR U37946 ( .A(n25521), .B(n37297), .Z(n25523) );
  XNOR U37947 ( .A(q[10]), .B(DB[1645]), .Z(n37297) );
  XNOR U37948 ( .A(q[9]), .B(DB[1644]), .Z(n25521) );
  IV U37949 ( .A(n25536), .Z(n37291) );
  XOR U37950 ( .A(n37298), .B(n37299), .Z(n25536) );
  XNOR U37951 ( .A(n25553), .B(n25534), .Z(n37299) );
  XNOR U37952 ( .A(q[0]), .B(DB[1635]), .Z(n25534) );
  XOR U37953 ( .A(n37300), .B(n25542), .Z(n25553) );
  XNOR U37954 ( .A(q[7]), .B(DB[1642]), .Z(n25542) );
  IV U37955 ( .A(n25541), .Z(n37300) );
  XNOR U37956 ( .A(n25539), .B(n37301), .Z(n25541) );
  XNOR U37957 ( .A(q[6]), .B(DB[1641]), .Z(n37301) );
  XNOR U37958 ( .A(q[5]), .B(DB[1640]), .Z(n25539) );
  IV U37959 ( .A(n25552), .Z(n37298) );
  XOR U37960 ( .A(n37302), .B(n37303), .Z(n25552) );
  XNOR U37961 ( .A(n25548), .B(n25550), .Z(n37303) );
  XNOR U37962 ( .A(q[1]), .B(DB[1636]), .Z(n25550) );
  XNOR U37963 ( .A(q[4]), .B(DB[1639]), .Z(n25548) );
  IV U37964 ( .A(n25547), .Z(n37302) );
  XNOR U37965 ( .A(n25545), .B(n37304), .Z(n25547) );
  XNOR U37966 ( .A(q[3]), .B(DB[1638]), .Z(n37304) );
  XNOR U37967 ( .A(q[2]), .B(DB[1637]), .Z(n25545) );
  XOR U37968 ( .A(n37305), .B(n25443), .Z(n25371) );
  XOR U37969 ( .A(n37306), .B(n25435), .Z(n25443) );
  XOR U37970 ( .A(n37307), .B(n25424), .Z(n25435) );
  XNOR U37971 ( .A(q[14]), .B(DB[1664]), .Z(n25424) );
  IV U37972 ( .A(n25423), .Z(n37307) );
  XNOR U37973 ( .A(n25421), .B(n37308), .Z(n25423) );
  XNOR U37974 ( .A(q[13]), .B(DB[1663]), .Z(n37308) );
  XNOR U37975 ( .A(q[12]), .B(DB[1662]), .Z(n25421) );
  IV U37976 ( .A(n25434), .Z(n37306) );
  XOR U37977 ( .A(n37309), .B(n37310), .Z(n25434) );
  XNOR U37978 ( .A(n25430), .B(n25432), .Z(n37310) );
  XNOR U37979 ( .A(q[8]), .B(DB[1658]), .Z(n25432) );
  XNOR U37980 ( .A(q[11]), .B(DB[1661]), .Z(n25430) );
  IV U37981 ( .A(n25429), .Z(n37309) );
  XNOR U37982 ( .A(n25427), .B(n37311), .Z(n25429) );
  XNOR U37983 ( .A(q[10]), .B(DB[1660]), .Z(n37311) );
  XNOR U37984 ( .A(q[9]), .B(DB[1659]), .Z(n25427) );
  IV U37985 ( .A(n25442), .Z(n37305) );
  XOR U37986 ( .A(n37312), .B(n37313), .Z(n25442) );
  XNOR U37987 ( .A(n25459), .B(n25440), .Z(n37313) );
  XNOR U37988 ( .A(q[0]), .B(DB[1650]), .Z(n25440) );
  XOR U37989 ( .A(n37314), .B(n25448), .Z(n25459) );
  XNOR U37990 ( .A(q[7]), .B(DB[1657]), .Z(n25448) );
  IV U37991 ( .A(n25447), .Z(n37314) );
  XNOR U37992 ( .A(n25445), .B(n37315), .Z(n25447) );
  XNOR U37993 ( .A(q[6]), .B(DB[1656]), .Z(n37315) );
  XNOR U37994 ( .A(q[5]), .B(DB[1655]), .Z(n25445) );
  IV U37995 ( .A(n25458), .Z(n37312) );
  XOR U37996 ( .A(n37316), .B(n37317), .Z(n25458) );
  XNOR U37997 ( .A(n25454), .B(n25456), .Z(n37317) );
  XNOR U37998 ( .A(q[1]), .B(DB[1651]), .Z(n25456) );
  XNOR U37999 ( .A(q[4]), .B(DB[1654]), .Z(n25454) );
  IV U38000 ( .A(n25453), .Z(n37316) );
  XNOR U38001 ( .A(n25451), .B(n37318), .Z(n25453) );
  XNOR U38002 ( .A(q[3]), .B(DB[1653]), .Z(n37318) );
  XNOR U38003 ( .A(q[2]), .B(DB[1652]), .Z(n25451) );
  XOR U38004 ( .A(n37319), .B(n25349), .Z(n25277) );
  XOR U38005 ( .A(n37320), .B(n25341), .Z(n25349) );
  XOR U38006 ( .A(n37321), .B(n25330), .Z(n25341) );
  XNOR U38007 ( .A(q[14]), .B(DB[1679]), .Z(n25330) );
  IV U38008 ( .A(n25329), .Z(n37321) );
  XNOR U38009 ( .A(n25327), .B(n37322), .Z(n25329) );
  XNOR U38010 ( .A(q[13]), .B(DB[1678]), .Z(n37322) );
  XNOR U38011 ( .A(q[12]), .B(DB[1677]), .Z(n25327) );
  IV U38012 ( .A(n25340), .Z(n37320) );
  XOR U38013 ( .A(n37323), .B(n37324), .Z(n25340) );
  XNOR U38014 ( .A(n25336), .B(n25338), .Z(n37324) );
  XNOR U38015 ( .A(q[8]), .B(DB[1673]), .Z(n25338) );
  XNOR U38016 ( .A(q[11]), .B(DB[1676]), .Z(n25336) );
  IV U38017 ( .A(n25335), .Z(n37323) );
  XNOR U38018 ( .A(n25333), .B(n37325), .Z(n25335) );
  XNOR U38019 ( .A(q[10]), .B(DB[1675]), .Z(n37325) );
  XNOR U38020 ( .A(q[9]), .B(DB[1674]), .Z(n25333) );
  IV U38021 ( .A(n25348), .Z(n37319) );
  XOR U38022 ( .A(n37326), .B(n37327), .Z(n25348) );
  XNOR U38023 ( .A(n25365), .B(n25346), .Z(n37327) );
  XNOR U38024 ( .A(q[0]), .B(DB[1665]), .Z(n25346) );
  XOR U38025 ( .A(n37328), .B(n25354), .Z(n25365) );
  XNOR U38026 ( .A(q[7]), .B(DB[1672]), .Z(n25354) );
  IV U38027 ( .A(n25353), .Z(n37328) );
  XNOR U38028 ( .A(n25351), .B(n37329), .Z(n25353) );
  XNOR U38029 ( .A(q[6]), .B(DB[1671]), .Z(n37329) );
  XNOR U38030 ( .A(q[5]), .B(DB[1670]), .Z(n25351) );
  IV U38031 ( .A(n25364), .Z(n37326) );
  XOR U38032 ( .A(n37330), .B(n37331), .Z(n25364) );
  XNOR U38033 ( .A(n25360), .B(n25362), .Z(n37331) );
  XNOR U38034 ( .A(q[1]), .B(DB[1666]), .Z(n25362) );
  XNOR U38035 ( .A(q[4]), .B(DB[1669]), .Z(n25360) );
  IV U38036 ( .A(n25359), .Z(n37330) );
  XNOR U38037 ( .A(n25357), .B(n37332), .Z(n25359) );
  XNOR U38038 ( .A(q[3]), .B(DB[1668]), .Z(n37332) );
  XNOR U38039 ( .A(q[2]), .B(DB[1667]), .Z(n25357) );
  XOR U38040 ( .A(n37333), .B(n25255), .Z(n25183) );
  XOR U38041 ( .A(n37334), .B(n25247), .Z(n25255) );
  XOR U38042 ( .A(n37335), .B(n25236), .Z(n25247) );
  XNOR U38043 ( .A(q[14]), .B(DB[1694]), .Z(n25236) );
  IV U38044 ( .A(n25235), .Z(n37335) );
  XNOR U38045 ( .A(n25233), .B(n37336), .Z(n25235) );
  XNOR U38046 ( .A(q[13]), .B(DB[1693]), .Z(n37336) );
  XNOR U38047 ( .A(q[12]), .B(DB[1692]), .Z(n25233) );
  IV U38048 ( .A(n25246), .Z(n37334) );
  XOR U38049 ( .A(n37337), .B(n37338), .Z(n25246) );
  XNOR U38050 ( .A(n25242), .B(n25244), .Z(n37338) );
  XNOR U38051 ( .A(q[8]), .B(DB[1688]), .Z(n25244) );
  XNOR U38052 ( .A(q[11]), .B(DB[1691]), .Z(n25242) );
  IV U38053 ( .A(n25241), .Z(n37337) );
  XNOR U38054 ( .A(n25239), .B(n37339), .Z(n25241) );
  XNOR U38055 ( .A(q[10]), .B(DB[1690]), .Z(n37339) );
  XNOR U38056 ( .A(q[9]), .B(DB[1689]), .Z(n25239) );
  IV U38057 ( .A(n25254), .Z(n37333) );
  XOR U38058 ( .A(n37340), .B(n37341), .Z(n25254) );
  XNOR U38059 ( .A(n25271), .B(n25252), .Z(n37341) );
  XNOR U38060 ( .A(q[0]), .B(DB[1680]), .Z(n25252) );
  XOR U38061 ( .A(n37342), .B(n25260), .Z(n25271) );
  XNOR U38062 ( .A(q[7]), .B(DB[1687]), .Z(n25260) );
  IV U38063 ( .A(n25259), .Z(n37342) );
  XNOR U38064 ( .A(n25257), .B(n37343), .Z(n25259) );
  XNOR U38065 ( .A(q[6]), .B(DB[1686]), .Z(n37343) );
  XNOR U38066 ( .A(q[5]), .B(DB[1685]), .Z(n25257) );
  IV U38067 ( .A(n25270), .Z(n37340) );
  XOR U38068 ( .A(n37344), .B(n37345), .Z(n25270) );
  XNOR U38069 ( .A(n25266), .B(n25268), .Z(n37345) );
  XNOR U38070 ( .A(q[1]), .B(DB[1681]), .Z(n25268) );
  XNOR U38071 ( .A(q[4]), .B(DB[1684]), .Z(n25266) );
  IV U38072 ( .A(n25265), .Z(n37344) );
  XNOR U38073 ( .A(n25263), .B(n37346), .Z(n25265) );
  XNOR U38074 ( .A(q[3]), .B(DB[1683]), .Z(n37346) );
  XNOR U38075 ( .A(q[2]), .B(DB[1682]), .Z(n25263) );
  XOR U38076 ( .A(n37347), .B(n25161), .Z(n25089) );
  XOR U38077 ( .A(n37348), .B(n25153), .Z(n25161) );
  XOR U38078 ( .A(n37349), .B(n25142), .Z(n25153) );
  XNOR U38079 ( .A(q[14]), .B(DB[1709]), .Z(n25142) );
  IV U38080 ( .A(n25141), .Z(n37349) );
  XNOR U38081 ( .A(n25139), .B(n37350), .Z(n25141) );
  XNOR U38082 ( .A(q[13]), .B(DB[1708]), .Z(n37350) );
  XNOR U38083 ( .A(q[12]), .B(DB[1707]), .Z(n25139) );
  IV U38084 ( .A(n25152), .Z(n37348) );
  XOR U38085 ( .A(n37351), .B(n37352), .Z(n25152) );
  XNOR U38086 ( .A(n25148), .B(n25150), .Z(n37352) );
  XNOR U38087 ( .A(q[8]), .B(DB[1703]), .Z(n25150) );
  XNOR U38088 ( .A(q[11]), .B(DB[1706]), .Z(n25148) );
  IV U38089 ( .A(n25147), .Z(n37351) );
  XNOR U38090 ( .A(n25145), .B(n37353), .Z(n25147) );
  XNOR U38091 ( .A(q[10]), .B(DB[1705]), .Z(n37353) );
  XNOR U38092 ( .A(q[9]), .B(DB[1704]), .Z(n25145) );
  IV U38093 ( .A(n25160), .Z(n37347) );
  XOR U38094 ( .A(n37354), .B(n37355), .Z(n25160) );
  XNOR U38095 ( .A(n25177), .B(n25158), .Z(n37355) );
  XNOR U38096 ( .A(q[0]), .B(DB[1695]), .Z(n25158) );
  XOR U38097 ( .A(n37356), .B(n25166), .Z(n25177) );
  XNOR U38098 ( .A(q[7]), .B(DB[1702]), .Z(n25166) );
  IV U38099 ( .A(n25165), .Z(n37356) );
  XNOR U38100 ( .A(n25163), .B(n37357), .Z(n25165) );
  XNOR U38101 ( .A(q[6]), .B(DB[1701]), .Z(n37357) );
  XNOR U38102 ( .A(q[5]), .B(DB[1700]), .Z(n25163) );
  IV U38103 ( .A(n25176), .Z(n37354) );
  XOR U38104 ( .A(n37358), .B(n37359), .Z(n25176) );
  XNOR U38105 ( .A(n25172), .B(n25174), .Z(n37359) );
  XNOR U38106 ( .A(q[1]), .B(DB[1696]), .Z(n25174) );
  XNOR U38107 ( .A(q[4]), .B(DB[1699]), .Z(n25172) );
  IV U38108 ( .A(n25171), .Z(n37358) );
  XNOR U38109 ( .A(n25169), .B(n37360), .Z(n25171) );
  XNOR U38110 ( .A(q[3]), .B(DB[1698]), .Z(n37360) );
  XNOR U38111 ( .A(q[2]), .B(DB[1697]), .Z(n25169) );
  XOR U38112 ( .A(n37361), .B(n25067), .Z(n24995) );
  XOR U38113 ( .A(n37362), .B(n25059), .Z(n25067) );
  XOR U38114 ( .A(n37363), .B(n25048), .Z(n25059) );
  XNOR U38115 ( .A(q[14]), .B(DB[1724]), .Z(n25048) );
  IV U38116 ( .A(n25047), .Z(n37363) );
  XNOR U38117 ( .A(n25045), .B(n37364), .Z(n25047) );
  XNOR U38118 ( .A(q[13]), .B(DB[1723]), .Z(n37364) );
  XNOR U38119 ( .A(q[12]), .B(DB[1722]), .Z(n25045) );
  IV U38120 ( .A(n25058), .Z(n37362) );
  XOR U38121 ( .A(n37365), .B(n37366), .Z(n25058) );
  XNOR U38122 ( .A(n25054), .B(n25056), .Z(n37366) );
  XNOR U38123 ( .A(q[8]), .B(DB[1718]), .Z(n25056) );
  XNOR U38124 ( .A(q[11]), .B(DB[1721]), .Z(n25054) );
  IV U38125 ( .A(n25053), .Z(n37365) );
  XNOR U38126 ( .A(n25051), .B(n37367), .Z(n25053) );
  XNOR U38127 ( .A(q[10]), .B(DB[1720]), .Z(n37367) );
  XNOR U38128 ( .A(q[9]), .B(DB[1719]), .Z(n25051) );
  IV U38129 ( .A(n25066), .Z(n37361) );
  XOR U38130 ( .A(n37368), .B(n37369), .Z(n25066) );
  XNOR U38131 ( .A(n25083), .B(n25064), .Z(n37369) );
  XNOR U38132 ( .A(q[0]), .B(DB[1710]), .Z(n25064) );
  XOR U38133 ( .A(n37370), .B(n25072), .Z(n25083) );
  XNOR U38134 ( .A(q[7]), .B(DB[1717]), .Z(n25072) );
  IV U38135 ( .A(n25071), .Z(n37370) );
  XNOR U38136 ( .A(n25069), .B(n37371), .Z(n25071) );
  XNOR U38137 ( .A(q[6]), .B(DB[1716]), .Z(n37371) );
  XNOR U38138 ( .A(q[5]), .B(DB[1715]), .Z(n25069) );
  IV U38139 ( .A(n25082), .Z(n37368) );
  XOR U38140 ( .A(n37372), .B(n37373), .Z(n25082) );
  XNOR U38141 ( .A(n25078), .B(n25080), .Z(n37373) );
  XNOR U38142 ( .A(q[1]), .B(DB[1711]), .Z(n25080) );
  XNOR U38143 ( .A(q[4]), .B(DB[1714]), .Z(n25078) );
  IV U38144 ( .A(n25077), .Z(n37372) );
  XNOR U38145 ( .A(n25075), .B(n37374), .Z(n25077) );
  XNOR U38146 ( .A(q[3]), .B(DB[1713]), .Z(n37374) );
  XNOR U38147 ( .A(q[2]), .B(DB[1712]), .Z(n25075) );
  XOR U38148 ( .A(n37375), .B(n24973), .Z(n24901) );
  XOR U38149 ( .A(n37376), .B(n24965), .Z(n24973) );
  XOR U38150 ( .A(n37377), .B(n24954), .Z(n24965) );
  XNOR U38151 ( .A(q[14]), .B(DB[1739]), .Z(n24954) );
  IV U38152 ( .A(n24953), .Z(n37377) );
  XNOR U38153 ( .A(n24951), .B(n37378), .Z(n24953) );
  XNOR U38154 ( .A(q[13]), .B(DB[1738]), .Z(n37378) );
  XNOR U38155 ( .A(q[12]), .B(DB[1737]), .Z(n24951) );
  IV U38156 ( .A(n24964), .Z(n37376) );
  XOR U38157 ( .A(n37379), .B(n37380), .Z(n24964) );
  XNOR U38158 ( .A(n24960), .B(n24962), .Z(n37380) );
  XNOR U38159 ( .A(q[8]), .B(DB[1733]), .Z(n24962) );
  XNOR U38160 ( .A(q[11]), .B(DB[1736]), .Z(n24960) );
  IV U38161 ( .A(n24959), .Z(n37379) );
  XNOR U38162 ( .A(n24957), .B(n37381), .Z(n24959) );
  XNOR U38163 ( .A(q[10]), .B(DB[1735]), .Z(n37381) );
  XNOR U38164 ( .A(q[9]), .B(DB[1734]), .Z(n24957) );
  IV U38165 ( .A(n24972), .Z(n37375) );
  XOR U38166 ( .A(n37382), .B(n37383), .Z(n24972) );
  XNOR U38167 ( .A(n24989), .B(n24970), .Z(n37383) );
  XNOR U38168 ( .A(q[0]), .B(DB[1725]), .Z(n24970) );
  XOR U38169 ( .A(n37384), .B(n24978), .Z(n24989) );
  XNOR U38170 ( .A(q[7]), .B(DB[1732]), .Z(n24978) );
  IV U38171 ( .A(n24977), .Z(n37384) );
  XNOR U38172 ( .A(n24975), .B(n37385), .Z(n24977) );
  XNOR U38173 ( .A(q[6]), .B(DB[1731]), .Z(n37385) );
  XNOR U38174 ( .A(q[5]), .B(DB[1730]), .Z(n24975) );
  IV U38175 ( .A(n24988), .Z(n37382) );
  XOR U38176 ( .A(n37386), .B(n37387), .Z(n24988) );
  XNOR U38177 ( .A(n24984), .B(n24986), .Z(n37387) );
  XNOR U38178 ( .A(q[1]), .B(DB[1726]), .Z(n24986) );
  XNOR U38179 ( .A(q[4]), .B(DB[1729]), .Z(n24984) );
  IV U38180 ( .A(n24983), .Z(n37386) );
  XNOR U38181 ( .A(n24981), .B(n37388), .Z(n24983) );
  XNOR U38182 ( .A(q[3]), .B(DB[1728]), .Z(n37388) );
  XNOR U38183 ( .A(q[2]), .B(DB[1727]), .Z(n24981) );
  XOR U38184 ( .A(n37389), .B(n24879), .Z(n24807) );
  XOR U38185 ( .A(n37390), .B(n24871), .Z(n24879) );
  XOR U38186 ( .A(n37391), .B(n24860), .Z(n24871) );
  XNOR U38187 ( .A(q[14]), .B(DB[1754]), .Z(n24860) );
  IV U38188 ( .A(n24859), .Z(n37391) );
  XNOR U38189 ( .A(n24857), .B(n37392), .Z(n24859) );
  XNOR U38190 ( .A(q[13]), .B(DB[1753]), .Z(n37392) );
  XNOR U38191 ( .A(q[12]), .B(DB[1752]), .Z(n24857) );
  IV U38192 ( .A(n24870), .Z(n37390) );
  XOR U38193 ( .A(n37393), .B(n37394), .Z(n24870) );
  XNOR U38194 ( .A(n24866), .B(n24868), .Z(n37394) );
  XNOR U38195 ( .A(q[8]), .B(DB[1748]), .Z(n24868) );
  XNOR U38196 ( .A(q[11]), .B(DB[1751]), .Z(n24866) );
  IV U38197 ( .A(n24865), .Z(n37393) );
  XNOR U38198 ( .A(n24863), .B(n37395), .Z(n24865) );
  XNOR U38199 ( .A(q[10]), .B(DB[1750]), .Z(n37395) );
  XNOR U38200 ( .A(q[9]), .B(DB[1749]), .Z(n24863) );
  IV U38201 ( .A(n24878), .Z(n37389) );
  XOR U38202 ( .A(n37396), .B(n37397), .Z(n24878) );
  XNOR U38203 ( .A(n24895), .B(n24876), .Z(n37397) );
  XNOR U38204 ( .A(q[0]), .B(DB[1740]), .Z(n24876) );
  XOR U38205 ( .A(n37398), .B(n24884), .Z(n24895) );
  XNOR U38206 ( .A(q[7]), .B(DB[1747]), .Z(n24884) );
  IV U38207 ( .A(n24883), .Z(n37398) );
  XNOR U38208 ( .A(n24881), .B(n37399), .Z(n24883) );
  XNOR U38209 ( .A(q[6]), .B(DB[1746]), .Z(n37399) );
  XNOR U38210 ( .A(q[5]), .B(DB[1745]), .Z(n24881) );
  IV U38211 ( .A(n24894), .Z(n37396) );
  XOR U38212 ( .A(n37400), .B(n37401), .Z(n24894) );
  XNOR U38213 ( .A(n24890), .B(n24892), .Z(n37401) );
  XNOR U38214 ( .A(q[1]), .B(DB[1741]), .Z(n24892) );
  XNOR U38215 ( .A(q[4]), .B(DB[1744]), .Z(n24890) );
  IV U38216 ( .A(n24889), .Z(n37400) );
  XNOR U38217 ( .A(n24887), .B(n37402), .Z(n24889) );
  XNOR U38218 ( .A(q[3]), .B(DB[1743]), .Z(n37402) );
  XNOR U38219 ( .A(q[2]), .B(DB[1742]), .Z(n24887) );
  XOR U38220 ( .A(n37403), .B(n24785), .Z(n24713) );
  XOR U38221 ( .A(n37404), .B(n24777), .Z(n24785) );
  XOR U38222 ( .A(n37405), .B(n24766), .Z(n24777) );
  XNOR U38223 ( .A(q[14]), .B(DB[1769]), .Z(n24766) );
  IV U38224 ( .A(n24765), .Z(n37405) );
  XNOR U38225 ( .A(n24763), .B(n37406), .Z(n24765) );
  XNOR U38226 ( .A(q[13]), .B(DB[1768]), .Z(n37406) );
  XNOR U38227 ( .A(q[12]), .B(DB[1767]), .Z(n24763) );
  IV U38228 ( .A(n24776), .Z(n37404) );
  XOR U38229 ( .A(n37407), .B(n37408), .Z(n24776) );
  XNOR U38230 ( .A(n24772), .B(n24774), .Z(n37408) );
  XNOR U38231 ( .A(q[8]), .B(DB[1763]), .Z(n24774) );
  XNOR U38232 ( .A(q[11]), .B(DB[1766]), .Z(n24772) );
  IV U38233 ( .A(n24771), .Z(n37407) );
  XNOR U38234 ( .A(n24769), .B(n37409), .Z(n24771) );
  XNOR U38235 ( .A(q[10]), .B(DB[1765]), .Z(n37409) );
  XNOR U38236 ( .A(q[9]), .B(DB[1764]), .Z(n24769) );
  IV U38237 ( .A(n24784), .Z(n37403) );
  XOR U38238 ( .A(n37410), .B(n37411), .Z(n24784) );
  XNOR U38239 ( .A(n24801), .B(n24782), .Z(n37411) );
  XNOR U38240 ( .A(q[0]), .B(DB[1755]), .Z(n24782) );
  XOR U38241 ( .A(n37412), .B(n24790), .Z(n24801) );
  XNOR U38242 ( .A(q[7]), .B(DB[1762]), .Z(n24790) );
  IV U38243 ( .A(n24789), .Z(n37412) );
  XNOR U38244 ( .A(n24787), .B(n37413), .Z(n24789) );
  XNOR U38245 ( .A(q[6]), .B(DB[1761]), .Z(n37413) );
  XNOR U38246 ( .A(q[5]), .B(DB[1760]), .Z(n24787) );
  IV U38247 ( .A(n24800), .Z(n37410) );
  XOR U38248 ( .A(n37414), .B(n37415), .Z(n24800) );
  XNOR U38249 ( .A(n24796), .B(n24798), .Z(n37415) );
  XNOR U38250 ( .A(q[1]), .B(DB[1756]), .Z(n24798) );
  XNOR U38251 ( .A(q[4]), .B(DB[1759]), .Z(n24796) );
  IV U38252 ( .A(n24795), .Z(n37414) );
  XNOR U38253 ( .A(n24793), .B(n37416), .Z(n24795) );
  XNOR U38254 ( .A(q[3]), .B(DB[1758]), .Z(n37416) );
  XNOR U38255 ( .A(q[2]), .B(DB[1757]), .Z(n24793) );
  XOR U38256 ( .A(n37417), .B(n24691), .Z(n24619) );
  XOR U38257 ( .A(n37418), .B(n24683), .Z(n24691) );
  XOR U38258 ( .A(n37419), .B(n24672), .Z(n24683) );
  XNOR U38259 ( .A(q[14]), .B(DB[1784]), .Z(n24672) );
  IV U38260 ( .A(n24671), .Z(n37419) );
  XNOR U38261 ( .A(n24669), .B(n37420), .Z(n24671) );
  XNOR U38262 ( .A(q[13]), .B(DB[1783]), .Z(n37420) );
  XNOR U38263 ( .A(q[12]), .B(DB[1782]), .Z(n24669) );
  IV U38264 ( .A(n24682), .Z(n37418) );
  XOR U38265 ( .A(n37421), .B(n37422), .Z(n24682) );
  XNOR U38266 ( .A(n24678), .B(n24680), .Z(n37422) );
  XNOR U38267 ( .A(q[8]), .B(DB[1778]), .Z(n24680) );
  XNOR U38268 ( .A(q[11]), .B(DB[1781]), .Z(n24678) );
  IV U38269 ( .A(n24677), .Z(n37421) );
  XNOR U38270 ( .A(n24675), .B(n37423), .Z(n24677) );
  XNOR U38271 ( .A(q[10]), .B(DB[1780]), .Z(n37423) );
  XNOR U38272 ( .A(q[9]), .B(DB[1779]), .Z(n24675) );
  IV U38273 ( .A(n24690), .Z(n37417) );
  XOR U38274 ( .A(n37424), .B(n37425), .Z(n24690) );
  XNOR U38275 ( .A(n24707), .B(n24688), .Z(n37425) );
  XNOR U38276 ( .A(q[0]), .B(DB[1770]), .Z(n24688) );
  XOR U38277 ( .A(n37426), .B(n24696), .Z(n24707) );
  XNOR U38278 ( .A(q[7]), .B(DB[1777]), .Z(n24696) );
  IV U38279 ( .A(n24695), .Z(n37426) );
  XNOR U38280 ( .A(n24693), .B(n37427), .Z(n24695) );
  XNOR U38281 ( .A(q[6]), .B(DB[1776]), .Z(n37427) );
  XNOR U38282 ( .A(q[5]), .B(DB[1775]), .Z(n24693) );
  IV U38283 ( .A(n24706), .Z(n37424) );
  XOR U38284 ( .A(n37428), .B(n37429), .Z(n24706) );
  XNOR U38285 ( .A(n24702), .B(n24704), .Z(n37429) );
  XNOR U38286 ( .A(q[1]), .B(DB[1771]), .Z(n24704) );
  XNOR U38287 ( .A(q[4]), .B(DB[1774]), .Z(n24702) );
  IV U38288 ( .A(n24701), .Z(n37428) );
  XNOR U38289 ( .A(n24699), .B(n37430), .Z(n24701) );
  XNOR U38290 ( .A(q[3]), .B(DB[1773]), .Z(n37430) );
  XNOR U38291 ( .A(q[2]), .B(DB[1772]), .Z(n24699) );
  XOR U38292 ( .A(n37431), .B(n24597), .Z(n24525) );
  XOR U38293 ( .A(n37432), .B(n24589), .Z(n24597) );
  XOR U38294 ( .A(n37433), .B(n24578), .Z(n24589) );
  XNOR U38295 ( .A(q[14]), .B(DB[1799]), .Z(n24578) );
  IV U38296 ( .A(n24577), .Z(n37433) );
  XNOR U38297 ( .A(n24575), .B(n37434), .Z(n24577) );
  XNOR U38298 ( .A(q[13]), .B(DB[1798]), .Z(n37434) );
  XNOR U38299 ( .A(q[12]), .B(DB[1797]), .Z(n24575) );
  IV U38300 ( .A(n24588), .Z(n37432) );
  XOR U38301 ( .A(n37435), .B(n37436), .Z(n24588) );
  XNOR U38302 ( .A(n24584), .B(n24586), .Z(n37436) );
  XNOR U38303 ( .A(q[8]), .B(DB[1793]), .Z(n24586) );
  XNOR U38304 ( .A(q[11]), .B(DB[1796]), .Z(n24584) );
  IV U38305 ( .A(n24583), .Z(n37435) );
  XNOR U38306 ( .A(n24581), .B(n37437), .Z(n24583) );
  XNOR U38307 ( .A(q[10]), .B(DB[1795]), .Z(n37437) );
  XNOR U38308 ( .A(q[9]), .B(DB[1794]), .Z(n24581) );
  IV U38309 ( .A(n24596), .Z(n37431) );
  XOR U38310 ( .A(n37438), .B(n37439), .Z(n24596) );
  XNOR U38311 ( .A(n24613), .B(n24594), .Z(n37439) );
  XNOR U38312 ( .A(q[0]), .B(DB[1785]), .Z(n24594) );
  XOR U38313 ( .A(n37440), .B(n24602), .Z(n24613) );
  XNOR U38314 ( .A(q[7]), .B(DB[1792]), .Z(n24602) );
  IV U38315 ( .A(n24601), .Z(n37440) );
  XNOR U38316 ( .A(n24599), .B(n37441), .Z(n24601) );
  XNOR U38317 ( .A(q[6]), .B(DB[1791]), .Z(n37441) );
  XNOR U38318 ( .A(q[5]), .B(DB[1790]), .Z(n24599) );
  IV U38319 ( .A(n24612), .Z(n37438) );
  XOR U38320 ( .A(n37442), .B(n37443), .Z(n24612) );
  XNOR U38321 ( .A(n24608), .B(n24610), .Z(n37443) );
  XNOR U38322 ( .A(q[1]), .B(DB[1786]), .Z(n24610) );
  XNOR U38323 ( .A(q[4]), .B(DB[1789]), .Z(n24608) );
  IV U38324 ( .A(n24607), .Z(n37442) );
  XNOR U38325 ( .A(n24605), .B(n37444), .Z(n24607) );
  XNOR U38326 ( .A(q[3]), .B(DB[1788]), .Z(n37444) );
  XNOR U38327 ( .A(q[2]), .B(DB[1787]), .Z(n24605) );
  XOR U38328 ( .A(n37445), .B(n24503), .Z(n24431) );
  XOR U38329 ( .A(n37446), .B(n24495), .Z(n24503) );
  XOR U38330 ( .A(n37447), .B(n24484), .Z(n24495) );
  XNOR U38331 ( .A(q[14]), .B(DB[1814]), .Z(n24484) );
  IV U38332 ( .A(n24483), .Z(n37447) );
  XNOR U38333 ( .A(n24481), .B(n37448), .Z(n24483) );
  XNOR U38334 ( .A(q[13]), .B(DB[1813]), .Z(n37448) );
  XNOR U38335 ( .A(q[12]), .B(DB[1812]), .Z(n24481) );
  IV U38336 ( .A(n24494), .Z(n37446) );
  XOR U38337 ( .A(n37449), .B(n37450), .Z(n24494) );
  XNOR U38338 ( .A(n24490), .B(n24492), .Z(n37450) );
  XNOR U38339 ( .A(q[8]), .B(DB[1808]), .Z(n24492) );
  XNOR U38340 ( .A(q[11]), .B(DB[1811]), .Z(n24490) );
  IV U38341 ( .A(n24489), .Z(n37449) );
  XNOR U38342 ( .A(n24487), .B(n37451), .Z(n24489) );
  XNOR U38343 ( .A(q[10]), .B(DB[1810]), .Z(n37451) );
  XNOR U38344 ( .A(q[9]), .B(DB[1809]), .Z(n24487) );
  IV U38345 ( .A(n24502), .Z(n37445) );
  XOR U38346 ( .A(n37452), .B(n37453), .Z(n24502) );
  XNOR U38347 ( .A(n24519), .B(n24500), .Z(n37453) );
  XNOR U38348 ( .A(q[0]), .B(DB[1800]), .Z(n24500) );
  XOR U38349 ( .A(n37454), .B(n24508), .Z(n24519) );
  XNOR U38350 ( .A(q[7]), .B(DB[1807]), .Z(n24508) );
  IV U38351 ( .A(n24507), .Z(n37454) );
  XNOR U38352 ( .A(n24505), .B(n37455), .Z(n24507) );
  XNOR U38353 ( .A(q[6]), .B(DB[1806]), .Z(n37455) );
  XNOR U38354 ( .A(q[5]), .B(DB[1805]), .Z(n24505) );
  IV U38355 ( .A(n24518), .Z(n37452) );
  XOR U38356 ( .A(n37456), .B(n37457), .Z(n24518) );
  XNOR U38357 ( .A(n24514), .B(n24516), .Z(n37457) );
  XNOR U38358 ( .A(q[1]), .B(DB[1801]), .Z(n24516) );
  XNOR U38359 ( .A(q[4]), .B(DB[1804]), .Z(n24514) );
  IV U38360 ( .A(n24513), .Z(n37456) );
  XNOR U38361 ( .A(n24511), .B(n37458), .Z(n24513) );
  XNOR U38362 ( .A(q[3]), .B(DB[1803]), .Z(n37458) );
  XNOR U38363 ( .A(q[2]), .B(DB[1802]), .Z(n24511) );
  XOR U38364 ( .A(n37459), .B(n24409), .Z(n24337) );
  XOR U38365 ( .A(n37460), .B(n24401), .Z(n24409) );
  XOR U38366 ( .A(n37461), .B(n24390), .Z(n24401) );
  XNOR U38367 ( .A(q[14]), .B(DB[1829]), .Z(n24390) );
  IV U38368 ( .A(n24389), .Z(n37461) );
  XNOR U38369 ( .A(n24387), .B(n37462), .Z(n24389) );
  XNOR U38370 ( .A(q[13]), .B(DB[1828]), .Z(n37462) );
  XNOR U38371 ( .A(q[12]), .B(DB[1827]), .Z(n24387) );
  IV U38372 ( .A(n24400), .Z(n37460) );
  XOR U38373 ( .A(n37463), .B(n37464), .Z(n24400) );
  XNOR U38374 ( .A(n24396), .B(n24398), .Z(n37464) );
  XNOR U38375 ( .A(q[8]), .B(DB[1823]), .Z(n24398) );
  XNOR U38376 ( .A(q[11]), .B(DB[1826]), .Z(n24396) );
  IV U38377 ( .A(n24395), .Z(n37463) );
  XNOR U38378 ( .A(n24393), .B(n37465), .Z(n24395) );
  XNOR U38379 ( .A(q[10]), .B(DB[1825]), .Z(n37465) );
  XNOR U38380 ( .A(q[9]), .B(DB[1824]), .Z(n24393) );
  IV U38381 ( .A(n24408), .Z(n37459) );
  XOR U38382 ( .A(n37466), .B(n37467), .Z(n24408) );
  XNOR U38383 ( .A(n24425), .B(n24406), .Z(n37467) );
  XNOR U38384 ( .A(q[0]), .B(DB[1815]), .Z(n24406) );
  XOR U38385 ( .A(n37468), .B(n24414), .Z(n24425) );
  XNOR U38386 ( .A(q[7]), .B(DB[1822]), .Z(n24414) );
  IV U38387 ( .A(n24413), .Z(n37468) );
  XNOR U38388 ( .A(n24411), .B(n37469), .Z(n24413) );
  XNOR U38389 ( .A(q[6]), .B(DB[1821]), .Z(n37469) );
  XNOR U38390 ( .A(q[5]), .B(DB[1820]), .Z(n24411) );
  IV U38391 ( .A(n24424), .Z(n37466) );
  XOR U38392 ( .A(n37470), .B(n37471), .Z(n24424) );
  XNOR U38393 ( .A(n24420), .B(n24422), .Z(n37471) );
  XNOR U38394 ( .A(q[1]), .B(DB[1816]), .Z(n24422) );
  XNOR U38395 ( .A(q[4]), .B(DB[1819]), .Z(n24420) );
  IV U38396 ( .A(n24419), .Z(n37470) );
  XNOR U38397 ( .A(n24417), .B(n37472), .Z(n24419) );
  XNOR U38398 ( .A(q[3]), .B(DB[1818]), .Z(n37472) );
  XNOR U38399 ( .A(q[2]), .B(DB[1817]), .Z(n24417) );
  XOR U38400 ( .A(n37473), .B(n24315), .Z(n24243) );
  XOR U38401 ( .A(n37474), .B(n24307), .Z(n24315) );
  XOR U38402 ( .A(n37475), .B(n24296), .Z(n24307) );
  XNOR U38403 ( .A(q[14]), .B(DB[1844]), .Z(n24296) );
  IV U38404 ( .A(n24295), .Z(n37475) );
  XNOR U38405 ( .A(n24293), .B(n37476), .Z(n24295) );
  XNOR U38406 ( .A(q[13]), .B(DB[1843]), .Z(n37476) );
  XNOR U38407 ( .A(q[12]), .B(DB[1842]), .Z(n24293) );
  IV U38408 ( .A(n24306), .Z(n37474) );
  XOR U38409 ( .A(n37477), .B(n37478), .Z(n24306) );
  XNOR U38410 ( .A(n24302), .B(n24304), .Z(n37478) );
  XNOR U38411 ( .A(q[8]), .B(DB[1838]), .Z(n24304) );
  XNOR U38412 ( .A(q[11]), .B(DB[1841]), .Z(n24302) );
  IV U38413 ( .A(n24301), .Z(n37477) );
  XNOR U38414 ( .A(n24299), .B(n37479), .Z(n24301) );
  XNOR U38415 ( .A(q[10]), .B(DB[1840]), .Z(n37479) );
  XNOR U38416 ( .A(q[9]), .B(DB[1839]), .Z(n24299) );
  IV U38417 ( .A(n24314), .Z(n37473) );
  XOR U38418 ( .A(n37480), .B(n37481), .Z(n24314) );
  XNOR U38419 ( .A(n24331), .B(n24312), .Z(n37481) );
  XNOR U38420 ( .A(q[0]), .B(DB[1830]), .Z(n24312) );
  XOR U38421 ( .A(n37482), .B(n24320), .Z(n24331) );
  XNOR U38422 ( .A(q[7]), .B(DB[1837]), .Z(n24320) );
  IV U38423 ( .A(n24319), .Z(n37482) );
  XNOR U38424 ( .A(n24317), .B(n37483), .Z(n24319) );
  XNOR U38425 ( .A(q[6]), .B(DB[1836]), .Z(n37483) );
  XNOR U38426 ( .A(q[5]), .B(DB[1835]), .Z(n24317) );
  IV U38427 ( .A(n24330), .Z(n37480) );
  XOR U38428 ( .A(n37484), .B(n37485), .Z(n24330) );
  XNOR U38429 ( .A(n24326), .B(n24328), .Z(n37485) );
  XNOR U38430 ( .A(q[1]), .B(DB[1831]), .Z(n24328) );
  XNOR U38431 ( .A(q[4]), .B(DB[1834]), .Z(n24326) );
  IV U38432 ( .A(n24325), .Z(n37484) );
  XNOR U38433 ( .A(n24323), .B(n37486), .Z(n24325) );
  XNOR U38434 ( .A(q[3]), .B(DB[1833]), .Z(n37486) );
  XNOR U38435 ( .A(q[2]), .B(DB[1832]), .Z(n24323) );
  XOR U38436 ( .A(n37487), .B(n24221), .Z(n24149) );
  XOR U38437 ( .A(n37488), .B(n24213), .Z(n24221) );
  XOR U38438 ( .A(n37489), .B(n24202), .Z(n24213) );
  XNOR U38439 ( .A(q[14]), .B(DB[1859]), .Z(n24202) );
  IV U38440 ( .A(n24201), .Z(n37489) );
  XNOR U38441 ( .A(n24199), .B(n37490), .Z(n24201) );
  XNOR U38442 ( .A(q[13]), .B(DB[1858]), .Z(n37490) );
  XNOR U38443 ( .A(q[12]), .B(DB[1857]), .Z(n24199) );
  IV U38444 ( .A(n24212), .Z(n37488) );
  XOR U38445 ( .A(n37491), .B(n37492), .Z(n24212) );
  XNOR U38446 ( .A(n24208), .B(n24210), .Z(n37492) );
  XNOR U38447 ( .A(q[8]), .B(DB[1853]), .Z(n24210) );
  XNOR U38448 ( .A(q[11]), .B(DB[1856]), .Z(n24208) );
  IV U38449 ( .A(n24207), .Z(n37491) );
  XNOR U38450 ( .A(n24205), .B(n37493), .Z(n24207) );
  XNOR U38451 ( .A(q[10]), .B(DB[1855]), .Z(n37493) );
  XNOR U38452 ( .A(q[9]), .B(DB[1854]), .Z(n24205) );
  IV U38453 ( .A(n24220), .Z(n37487) );
  XOR U38454 ( .A(n37494), .B(n37495), .Z(n24220) );
  XNOR U38455 ( .A(n24237), .B(n24218), .Z(n37495) );
  XNOR U38456 ( .A(q[0]), .B(DB[1845]), .Z(n24218) );
  XOR U38457 ( .A(n37496), .B(n24226), .Z(n24237) );
  XNOR U38458 ( .A(q[7]), .B(DB[1852]), .Z(n24226) );
  IV U38459 ( .A(n24225), .Z(n37496) );
  XNOR U38460 ( .A(n24223), .B(n37497), .Z(n24225) );
  XNOR U38461 ( .A(q[6]), .B(DB[1851]), .Z(n37497) );
  XNOR U38462 ( .A(q[5]), .B(DB[1850]), .Z(n24223) );
  IV U38463 ( .A(n24236), .Z(n37494) );
  XOR U38464 ( .A(n37498), .B(n37499), .Z(n24236) );
  XNOR U38465 ( .A(n24232), .B(n24234), .Z(n37499) );
  XNOR U38466 ( .A(q[1]), .B(DB[1846]), .Z(n24234) );
  XNOR U38467 ( .A(q[4]), .B(DB[1849]), .Z(n24232) );
  IV U38468 ( .A(n24231), .Z(n37498) );
  XNOR U38469 ( .A(n24229), .B(n37500), .Z(n24231) );
  XNOR U38470 ( .A(q[3]), .B(DB[1848]), .Z(n37500) );
  XNOR U38471 ( .A(q[2]), .B(DB[1847]), .Z(n24229) );
  XOR U38472 ( .A(n37501), .B(n24127), .Z(n24055) );
  XOR U38473 ( .A(n37502), .B(n24119), .Z(n24127) );
  XOR U38474 ( .A(n37503), .B(n24108), .Z(n24119) );
  XNOR U38475 ( .A(q[14]), .B(DB[1874]), .Z(n24108) );
  IV U38476 ( .A(n24107), .Z(n37503) );
  XNOR U38477 ( .A(n24105), .B(n37504), .Z(n24107) );
  XNOR U38478 ( .A(q[13]), .B(DB[1873]), .Z(n37504) );
  XNOR U38479 ( .A(q[12]), .B(DB[1872]), .Z(n24105) );
  IV U38480 ( .A(n24118), .Z(n37502) );
  XOR U38481 ( .A(n37505), .B(n37506), .Z(n24118) );
  XNOR U38482 ( .A(n24114), .B(n24116), .Z(n37506) );
  XNOR U38483 ( .A(q[8]), .B(DB[1868]), .Z(n24116) );
  XNOR U38484 ( .A(q[11]), .B(DB[1871]), .Z(n24114) );
  IV U38485 ( .A(n24113), .Z(n37505) );
  XNOR U38486 ( .A(n24111), .B(n37507), .Z(n24113) );
  XNOR U38487 ( .A(q[10]), .B(DB[1870]), .Z(n37507) );
  XNOR U38488 ( .A(q[9]), .B(DB[1869]), .Z(n24111) );
  IV U38489 ( .A(n24126), .Z(n37501) );
  XOR U38490 ( .A(n37508), .B(n37509), .Z(n24126) );
  XNOR U38491 ( .A(n24143), .B(n24124), .Z(n37509) );
  XNOR U38492 ( .A(q[0]), .B(DB[1860]), .Z(n24124) );
  XOR U38493 ( .A(n37510), .B(n24132), .Z(n24143) );
  XNOR U38494 ( .A(q[7]), .B(DB[1867]), .Z(n24132) );
  IV U38495 ( .A(n24131), .Z(n37510) );
  XNOR U38496 ( .A(n24129), .B(n37511), .Z(n24131) );
  XNOR U38497 ( .A(q[6]), .B(DB[1866]), .Z(n37511) );
  XNOR U38498 ( .A(q[5]), .B(DB[1865]), .Z(n24129) );
  IV U38499 ( .A(n24142), .Z(n37508) );
  XOR U38500 ( .A(n37512), .B(n37513), .Z(n24142) );
  XNOR U38501 ( .A(n24138), .B(n24140), .Z(n37513) );
  XNOR U38502 ( .A(q[1]), .B(DB[1861]), .Z(n24140) );
  XNOR U38503 ( .A(q[4]), .B(DB[1864]), .Z(n24138) );
  IV U38504 ( .A(n24137), .Z(n37512) );
  XNOR U38505 ( .A(n24135), .B(n37514), .Z(n24137) );
  XNOR U38506 ( .A(q[3]), .B(DB[1863]), .Z(n37514) );
  XNOR U38507 ( .A(q[2]), .B(DB[1862]), .Z(n24135) );
  XOR U38508 ( .A(n37515), .B(n24033), .Z(n23961) );
  XOR U38509 ( .A(n37516), .B(n24025), .Z(n24033) );
  XOR U38510 ( .A(n37517), .B(n24014), .Z(n24025) );
  XNOR U38511 ( .A(q[14]), .B(DB[1889]), .Z(n24014) );
  IV U38512 ( .A(n24013), .Z(n37517) );
  XNOR U38513 ( .A(n24011), .B(n37518), .Z(n24013) );
  XNOR U38514 ( .A(q[13]), .B(DB[1888]), .Z(n37518) );
  XNOR U38515 ( .A(q[12]), .B(DB[1887]), .Z(n24011) );
  IV U38516 ( .A(n24024), .Z(n37516) );
  XOR U38517 ( .A(n37519), .B(n37520), .Z(n24024) );
  XNOR U38518 ( .A(n24020), .B(n24022), .Z(n37520) );
  XNOR U38519 ( .A(q[8]), .B(DB[1883]), .Z(n24022) );
  XNOR U38520 ( .A(q[11]), .B(DB[1886]), .Z(n24020) );
  IV U38521 ( .A(n24019), .Z(n37519) );
  XNOR U38522 ( .A(n24017), .B(n37521), .Z(n24019) );
  XNOR U38523 ( .A(q[10]), .B(DB[1885]), .Z(n37521) );
  XNOR U38524 ( .A(q[9]), .B(DB[1884]), .Z(n24017) );
  IV U38525 ( .A(n24032), .Z(n37515) );
  XOR U38526 ( .A(n37522), .B(n37523), .Z(n24032) );
  XNOR U38527 ( .A(n24049), .B(n24030), .Z(n37523) );
  XNOR U38528 ( .A(q[0]), .B(DB[1875]), .Z(n24030) );
  XOR U38529 ( .A(n37524), .B(n24038), .Z(n24049) );
  XNOR U38530 ( .A(q[7]), .B(DB[1882]), .Z(n24038) );
  IV U38531 ( .A(n24037), .Z(n37524) );
  XNOR U38532 ( .A(n24035), .B(n37525), .Z(n24037) );
  XNOR U38533 ( .A(q[6]), .B(DB[1881]), .Z(n37525) );
  XNOR U38534 ( .A(q[5]), .B(DB[1880]), .Z(n24035) );
  IV U38535 ( .A(n24048), .Z(n37522) );
  XOR U38536 ( .A(n37526), .B(n37527), .Z(n24048) );
  XNOR U38537 ( .A(n24044), .B(n24046), .Z(n37527) );
  XNOR U38538 ( .A(q[1]), .B(DB[1876]), .Z(n24046) );
  XNOR U38539 ( .A(q[4]), .B(DB[1879]), .Z(n24044) );
  IV U38540 ( .A(n24043), .Z(n37526) );
  XNOR U38541 ( .A(n24041), .B(n37528), .Z(n24043) );
  XNOR U38542 ( .A(q[3]), .B(DB[1878]), .Z(n37528) );
  XNOR U38543 ( .A(q[2]), .B(DB[1877]), .Z(n24041) );
  XOR U38544 ( .A(n37529), .B(n23939), .Z(n23867) );
  XOR U38545 ( .A(n37530), .B(n23931), .Z(n23939) );
  XOR U38546 ( .A(n37531), .B(n23920), .Z(n23931) );
  XNOR U38547 ( .A(q[14]), .B(DB[1904]), .Z(n23920) );
  IV U38548 ( .A(n23919), .Z(n37531) );
  XNOR U38549 ( .A(n23917), .B(n37532), .Z(n23919) );
  XNOR U38550 ( .A(q[13]), .B(DB[1903]), .Z(n37532) );
  XNOR U38551 ( .A(q[12]), .B(DB[1902]), .Z(n23917) );
  IV U38552 ( .A(n23930), .Z(n37530) );
  XOR U38553 ( .A(n37533), .B(n37534), .Z(n23930) );
  XNOR U38554 ( .A(n23926), .B(n23928), .Z(n37534) );
  XNOR U38555 ( .A(q[8]), .B(DB[1898]), .Z(n23928) );
  XNOR U38556 ( .A(q[11]), .B(DB[1901]), .Z(n23926) );
  IV U38557 ( .A(n23925), .Z(n37533) );
  XNOR U38558 ( .A(n23923), .B(n37535), .Z(n23925) );
  XNOR U38559 ( .A(q[10]), .B(DB[1900]), .Z(n37535) );
  XNOR U38560 ( .A(q[9]), .B(DB[1899]), .Z(n23923) );
  IV U38561 ( .A(n23938), .Z(n37529) );
  XOR U38562 ( .A(n37536), .B(n37537), .Z(n23938) );
  XNOR U38563 ( .A(n23955), .B(n23936), .Z(n37537) );
  XNOR U38564 ( .A(q[0]), .B(DB[1890]), .Z(n23936) );
  XOR U38565 ( .A(n37538), .B(n23944), .Z(n23955) );
  XNOR U38566 ( .A(q[7]), .B(DB[1897]), .Z(n23944) );
  IV U38567 ( .A(n23943), .Z(n37538) );
  XNOR U38568 ( .A(n23941), .B(n37539), .Z(n23943) );
  XNOR U38569 ( .A(q[6]), .B(DB[1896]), .Z(n37539) );
  XNOR U38570 ( .A(q[5]), .B(DB[1895]), .Z(n23941) );
  IV U38571 ( .A(n23954), .Z(n37536) );
  XOR U38572 ( .A(n37540), .B(n37541), .Z(n23954) );
  XNOR U38573 ( .A(n23950), .B(n23952), .Z(n37541) );
  XNOR U38574 ( .A(q[1]), .B(DB[1891]), .Z(n23952) );
  XNOR U38575 ( .A(q[4]), .B(DB[1894]), .Z(n23950) );
  IV U38576 ( .A(n23949), .Z(n37540) );
  XNOR U38577 ( .A(n23947), .B(n37542), .Z(n23949) );
  XNOR U38578 ( .A(q[3]), .B(DB[1893]), .Z(n37542) );
  XNOR U38579 ( .A(q[2]), .B(DB[1892]), .Z(n23947) );
  XOR U38580 ( .A(n37543), .B(n23845), .Z(n23773) );
  XOR U38581 ( .A(n37544), .B(n23837), .Z(n23845) );
  XOR U38582 ( .A(n37545), .B(n23826), .Z(n23837) );
  XNOR U38583 ( .A(q[14]), .B(DB[1919]), .Z(n23826) );
  IV U38584 ( .A(n23825), .Z(n37545) );
  XNOR U38585 ( .A(n23823), .B(n37546), .Z(n23825) );
  XNOR U38586 ( .A(q[13]), .B(DB[1918]), .Z(n37546) );
  XNOR U38587 ( .A(q[12]), .B(DB[1917]), .Z(n23823) );
  IV U38588 ( .A(n23836), .Z(n37544) );
  XOR U38589 ( .A(n37547), .B(n37548), .Z(n23836) );
  XNOR U38590 ( .A(n23832), .B(n23834), .Z(n37548) );
  XNOR U38591 ( .A(q[8]), .B(DB[1913]), .Z(n23834) );
  XNOR U38592 ( .A(q[11]), .B(DB[1916]), .Z(n23832) );
  IV U38593 ( .A(n23831), .Z(n37547) );
  XNOR U38594 ( .A(n23829), .B(n37549), .Z(n23831) );
  XNOR U38595 ( .A(q[10]), .B(DB[1915]), .Z(n37549) );
  XNOR U38596 ( .A(q[9]), .B(DB[1914]), .Z(n23829) );
  IV U38597 ( .A(n23844), .Z(n37543) );
  XOR U38598 ( .A(n37550), .B(n37551), .Z(n23844) );
  XNOR U38599 ( .A(n23861), .B(n23842), .Z(n37551) );
  XNOR U38600 ( .A(q[0]), .B(DB[1905]), .Z(n23842) );
  XOR U38601 ( .A(n37552), .B(n23850), .Z(n23861) );
  XNOR U38602 ( .A(q[7]), .B(DB[1912]), .Z(n23850) );
  IV U38603 ( .A(n23849), .Z(n37552) );
  XNOR U38604 ( .A(n23847), .B(n37553), .Z(n23849) );
  XNOR U38605 ( .A(q[6]), .B(DB[1911]), .Z(n37553) );
  XNOR U38606 ( .A(q[5]), .B(DB[1910]), .Z(n23847) );
  IV U38607 ( .A(n23860), .Z(n37550) );
  XOR U38608 ( .A(n37554), .B(n37555), .Z(n23860) );
  XNOR U38609 ( .A(n23856), .B(n23858), .Z(n37555) );
  XNOR U38610 ( .A(q[1]), .B(DB[1906]), .Z(n23858) );
  XNOR U38611 ( .A(q[4]), .B(DB[1909]), .Z(n23856) );
  IV U38612 ( .A(n23855), .Z(n37554) );
  XNOR U38613 ( .A(n23853), .B(n37556), .Z(n23855) );
  XNOR U38614 ( .A(q[3]), .B(DB[1908]), .Z(n37556) );
  XNOR U38615 ( .A(q[2]), .B(DB[1907]), .Z(n23853) );
  XOR U38616 ( .A(n37557), .B(n23751), .Z(n23679) );
  XOR U38617 ( .A(n37558), .B(n23743), .Z(n23751) );
  XOR U38618 ( .A(n37559), .B(n23732), .Z(n23743) );
  XNOR U38619 ( .A(q[14]), .B(DB[1934]), .Z(n23732) );
  IV U38620 ( .A(n23731), .Z(n37559) );
  XNOR U38621 ( .A(n23729), .B(n37560), .Z(n23731) );
  XNOR U38622 ( .A(q[13]), .B(DB[1933]), .Z(n37560) );
  XNOR U38623 ( .A(q[12]), .B(DB[1932]), .Z(n23729) );
  IV U38624 ( .A(n23742), .Z(n37558) );
  XOR U38625 ( .A(n37561), .B(n37562), .Z(n23742) );
  XNOR U38626 ( .A(n23738), .B(n23740), .Z(n37562) );
  XNOR U38627 ( .A(q[8]), .B(DB[1928]), .Z(n23740) );
  XNOR U38628 ( .A(q[11]), .B(DB[1931]), .Z(n23738) );
  IV U38629 ( .A(n23737), .Z(n37561) );
  XNOR U38630 ( .A(n23735), .B(n37563), .Z(n23737) );
  XNOR U38631 ( .A(q[10]), .B(DB[1930]), .Z(n37563) );
  XNOR U38632 ( .A(q[9]), .B(DB[1929]), .Z(n23735) );
  IV U38633 ( .A(n23750), .Z(n37557) );
  XOR U38634 ( .A(n37564), .B(n37565), .Z(n23750) );
  XNOR U38635 ( .A(n23767), .B(n23748), .Z(n37565) );
  XNOR U38636 ( .A(q[0]), .B(DB[1920]), .Z(n23748) );
  XOR U38637 ( .A(n37566), .B(n23756), .Z(n23767) );
  XNOR U38638 ( .A(q[7]), .B(DB[1927]), .Z(n23756) );
  IV U38639 ( .A(n23755), .Z(n37566) );
  XNOR U38640 ( .A(n23753), .B(n37567), .Z(n23755) );
  XNOR U38641 ( .A(q[6]), .B(DB[1926]), .Z(n37567) );
  XNOR U38642 ( .A(q[5]), .B(DB[1925]), .Z(n23753) );
  IV U38643 ( .A(n23766), .Z(n37564) );
  XOR U38644 ( .A(n37568), .B(n37569), .Z(n23766) );
  XNOR U38645 ( .A(n23762), .B(n23764), .Z(n37569) );
  XNOR U38646 ( .A(q[1]), .B(DB[1921]), .Z(n23764) );
  XNOR U38647 ( .A(q[4]), .B(DB[1924]), .Z(n23762) );
  IV U38648 ( .A(n23761), .Z(n37568) );
  XNOR U38649 ( .A(n23759), .B(n37570), .Z(n23761) );
  XNOR U38650 ( .A(q[3]), .B(DB[1923]), .Z(n37570) );
  XNOR U38651 ( .A(q[2]), .B(DB[1922]), .Z(n23759) );
  XOR U38652 ( .A(n37571), .B(n23657), .Z(n23585) );
  XOR U38653 ( .A(n37572), .B(n23649), .Z(n23657) );
  XOR U38654 ( .A(n37573), .B(n23638), .Z(n23649) );
  XNOR U38655 ( .A(q[14]), .B(DB[1949]), .Z(n23638) );
  IV U38656 ( .A(n23637), .Z(n37573) );
  XNOR U38657 ( .A(n23635), .B(n37574), .Z(n23637) );
  XNOR U38658 ( .A(q[13]), .B(DB[1948]), .Z(n37574) );
  XNOR U38659 ( .A(q[12]), .B(DB[1947]), .Z(n23635) );
  IV U38660 ( .A(n23648), .Z(n37572) );
  XOR U38661 ( .A(n37575), .B(n37576), .Z(n23648) );
  XNOR U38662 ( .A(n23644), .B(n23646), .Z(n37576) );
  XNOR U38663 ( .A(q[8]), .B(DB[1943]), .Z(n23646) );
  XNOR U38664 ( .A(q[11]), .B(DB[1946]), .Z(n23644) );
  IV U38665 ( .A(n23643), .Z(n37575) );
  XNOR U38666 ( .A(n23641), .B(n37577), .Z(n23643) );
  XNOR U38667 ( .A(q[10]), .B(DB[1945]), .Z(n37577) );
  XNOR U38668 ( .A(q[9]), .B(DB[1944]), .Z(n23641) );
  IV U38669 ( .A(n23656), .Z(n37571) );
  XOR U38670 ( .A(n37578), .B(n37579), .Z(n23656) );
  XNOR U38671 ( .A(n23673), .B(n23654), .Z(n37579) );
  XNOR U38672 ( .A(q[0]), .B(DB[1935]), .Z(n23654) );
  XOR U38673 ( .A(n37580), .B(n23662), .Z(n23673) );
  XNOR U38674 ( .A(q[7]), .B(DB[1942]), .Z(n23662) );
  IV U38675 ( .A(n23661), .Z(n37580) );
  XNOR U38676 ( .A(n23659), .B(n37581), .Z(n23661) );
  XNOR U38677 ( .A(q[6]), .B(DB[1941]), .Z(n37581) );
  XNOR U38678 ( .A(q[5]), .B(DB[1940]), .Z(n23659) );
  IV U38679 ( .A(n23672), .Z(n37578) );
  XOR U38680 ( .A(n37582), .B(n37583), .Z(n23672) );
  XNOR U38681 ( .A(n23668), .B(n23670), .Z(n37583) );
  XNOR U38682 ( .A(q[1]), .B(DB[1936]), .Z(n23670) );
  XNOR U38683 ( .A(q[4]), .B(DB[1939]), .Z(n23668) );
  IV U38684 ( .A(n23667), .Z(n37582) );
  XNOR U38685 ( .A(n23665), .B(n37584), .Z(n23667) );
  XNOR U38686 ( .A(q[3]), .B(DB[1938]), .Z(n37584) );
  XNOR U38687 ( .A(q[2]), .B(DB[1937]), .Z(n23665) );
  XOR U38688 ( .A(n37585), .B(n23563), .Z(n23491) );
  XOR U38689 ( .A(n37586), .B(n23555), .Z(n23563) );
  XOR U38690 ( .A(n37587), .B(n23544), .Z(n23555) );
  XNOR U38691 ( .A(q[14]), .B(DB[1964]), .Z(n23544) );
  IV U38692 ( .A(n23543), .Z(n37587) );
  XNOR U38693 ( .A(n23541), .B(n37588), .Z(n23543) );
  XNOR U38694 ( .A(q[13]), .B(DB[1963]), .Z(n37588) );
  XNOR U38695 ( .A(q[12]), .B(DB[1962]), .Z(n23541) );
  IV U38696 ( .A(n23554), .Z(n37586) );
  XOR U38697 ( .A(n37589), .B(n37590), .Z(n23554) );
  XNOR U38698 ( .A(n23550), .B(n23552), .Z(n37590) );
  XNOR U38699 ( .A(q[8]), .B(DB[1958]), .Z(n23552) );
  XNOR U38700 ( .A(q[11]), .B(DB[1961]), .Z(n23550) );
  IV U38701 ( .A(n23549), .Z(n37589) );
  XNOR U38702 ( .A(n23547), .B(n37591), .Z(n23549) );
  XNOR U38703 ( .A(q[10]), .B(DB[1960]), .Z(n37591) );
  XNOR U38704 ( .A(q[9]), .B(DB[1959]), .Z(n23547) );
  IV U38705 ( .A(n23562), .Z(n37585) );
  XOR U38706 ( .A(n37592), .B(n37593), .Z(n23562) );
  XNOR U38707 ( .A(n23579), .B(n23560), .Z(n37593) );
  XNOR U38708 ( .A(q[0]), .B(DB[1950]), .Z(n23560) );
  XOR U38709 ( .A(n37594), .B(n23568), .Z(n23579) );
  XNOR U38710 ( .A(q[7]), .B(DB[1957]), .Z(n23568) );
  IV U38711 ( .A(n23567), .Z(n37594) );
  XNOR U38712 ( .A(n23565), .B(n37595), .Z(n23567) );
  XNOR U38713 ( .A(q[6]), .B(DB[1956]), .Z(n37595) );
  XNOR U38714 ( .A(q[5]), .B(DB[1955]), .Z(n23565) );
  IV U38715 ( .A(n23578), .Z(n37592) );
  XOR U38716 ( .A(n37596), .B(n37597), .Z(n23578) );
  XNOR U38717 ( .A(n23574), .B(n23576), .Z(n37597) );
  XNOR U38718 ( .A(q[1]), .B(DB[1951]), .Z(n23576) );
  XNOR U38719 ( .A(q[4]), .B(DB[1954]), .Z(n23574) );
  IV U38720 ( .A(n23573), .Z(n37596) );
  XNOR U38721 ( .A(n23571), .B(n37598), .Z(n23573) );
  XNOR U38722 ( .A(q[3]), .B(DB[1953]), .Z(n37598) );
  XNOR U38723 ( .A(q[2]), .B(DB[1952]), .Z(n23571) );
  XOR U38724 ( .A(n37599), .B(n23469), .Z(n23397) );
  XOR U38725 ( .A(n37600), .B(n23461), .Z(n23469) );
  XOR U38726 ( .A(n37601), .B(n23450), .Z(n23461) );
  XNOR U38727 ( .A(q[14]), .B(DB[1979]), .Z(n23450) );
  IV U38728 ( .A(n23449), .Z(n37601) );
  XNOR U38729 ( .A(n23447), .B(n37602), .Z(n23449) );
  XNOR U38730 ( .A(q[13]), .B(DB[1978]), .Z(n37602) );
  XNOR U38731 ( .A(q[12]), .B(DB[1977]), .Z(n23447) );
  IV U38732 ( .A(n23460), .Z(n37600) );
  XOR U38733 ( .A(n37603), .B(n37604), .Z(n23460) );
  XNOR U38734 ( .A(n23456), .B(n23458), .Z(n37604) );
  XNOR U38735 ( .A(q[8]), .B(DB[1973]), .Z(n23458) );
  XNOR U38736 ( .A(q[11]), .B(DB[1976]), .Z(n23456) );
  IV U38737 ( .A(n23455), .Z(n37603) );
  XNOR U38738 ( .A(n23453), .B(n37605), .Z(n23455) );
  XNOR U38739 ( .A(q[10]), .B(DB[1975]), .Z(n37605) );
  XNOR U38740 ( .A(q[9]), .B(DB[1974]), .Z(n23453) );
  IV U38741 ( .A(n23468), .Z(n37599) );
  XOR U38742 ( .A(n37606), .B(n37607), .Z(n23468) );
  XNOR U38743 ( .A(n23485), .B(n23466), .Z(n37607) );
  XNOR U38744 ( .A(q[0]), .B(DB[1965]), .Z(n23466) );
  XOR U38745 ( .A(n37608), .B(n23474), .Z(n23485) );
  XNOR U38746 ( .A(q[7]), .B(DB[1972]), .Z(n23474) );
  IV U38747 ( .A(n23473), .Z(n37608) );
  XNOR U38748 ( .A(n23471), .B(n37609), .Z(n23473) );
  XNOR U38749 ( .A(q[6]), .B(DB[1971]), .Z(n37609) );
  XNOR U38750 ( .A(q[5]), .B(DB[1970]), .Z(n23471) );
  IV U38751 ( .A(n23484), .Z(n37606) );
  XOR U38752 ( .A(n37610), .B(n37611), .Z(n23484) );
  XNOR U38753 ( .A(n23480), .B(n23482), .Z(n37611) );
  XNOR U38754 ( .A(q[1]), .B(DB[1966]), .Z(n23482) );
  XNOR U38755 ( .A(q[4]), .B(DB[1969]), .Z(n23480) );
  IV U38756 ( .A(n23479), .Z(n37610) );
  XNOR U38757 ( .A(n23477), .B(n37612), .Z(n23479) );
  XNOR U38758 ( .A(q[3]), .B(DB[1968]), .Z(n37612) );
  XNOR U38759 ( .A(q[2]), .B(DB[1967]), .Z(n23477) );
  XOR U38760 ( .A(n37613), .B(n23375), .Z(n23303) );
  XOR U38761 ( .A(n37614), .B(n23367), .Z(n23375) );
  XOR U38762 ( .A(n37615), .B(n23356), .Z(n23367) );
  XNOR U38763 ( .A(q[14]), .B(DB[1994]), .Z(n23356) );
  IV U38764 ( .A(n23355), .Z(n37615) );
  XNOR U38765 ( .A(n23353), .B(n37616), .Z(n23355) );
  XNOR U38766 ( .A(q[13]), .B(DB[1993]), .Z(n37616) );
  XNOR U38767 ( .A(q[12]), .B(DB[1992]), .Z(n23353) );
  IV U38768 ( .A(n23366), .Z(n37614) );
  XOR U38769 ( .A(n37617), .B(n37618), .Z(n23366) );
  XNOR U38770 ( .A(n23362), .B(n23364), .Z(n37618) );
  XNOR U38771 ( .A(q[8]), .B(DB[1988]), .Z(n23364) );
  XNOR U38772 ( .A(q[11]), .B(DB[1991]), .Z(n23362) );
  IV U38773 ( .A(n23361), .Z(n37617) );
  XNOR U38774 ( .A(n23359), .B(n37619), .Z(n23361) );
  XNOR U38775 ( .A(q[10]), .B(DB[1990]), .Z(n37619) );
  XNOR U38776 ( .A(q[9]), .B(DB[1989]), .Z(n23359) );
  IV U38777 ( .A(n23374), .Z(n37613) );
  XOR U38778 ( .A(n37620), .B(n37621), .Z(n23374) );
  XNOR U38779 ( .A(n23391), .B(n23372), .Z(n37621) );
  XNOR U38780 ( .A(q[0]), .B(DB[1980]), .Z(n23372) );
  XOR U38781 ( .A(n37622), .B(n23380), .Z(n23391) );
  XNOR U38782 ( .A(q[7]), .B(DB[1987]), .Z(n23380) );
  IV U38783 ( .A(n23379), .Z(n37622) );
  XNOR U38784 ( .A(n23377), .B(n37623), .Z(n23379) );
  XNOR U38785 ( .A(q[6]), .B(DB[1986]), .Z(n37623) );
  XNOR U38786 ( .A(q[5]), .B(DB[1985]), .Z(n23377) );
  IV U38787 ( .A(n23390), .Z(n37620) );
  XOR U38788 ( .A(n37624), .B(n37625), .Z(n23390) );
  XNOR U38789 ( .A(n23386), .B(n23388), .Z(n37625) );
  XNOR U38790 ( .A(q[1]), .B(DB[1981]), .Z(n23388) );
  XNOR U38791 ( .A(q[4]), .B(DB[1984]), .Z(n23386) );
  IV U38792 ( .A(n23385), .Z(n37624) );
  XNOR U38793 ( .A(n23383), .B(n37626), .Z(n23385) );
  XNOR U38794 ( .A(q[3]), .B(DB[1983]), .Z(n37626) );
  XNOR U38795 ( .A(q[2]), .B(DB[1982]), .Z(n23383) );
  XOR U38796 ( .A(n37627), .B(n23281), .Z(n23209) );
  XOR U38797 ( .A(n37628), .B(n23273), .Z(n23281) );
  XOR U38798 ( .A(n37629), .B(n23262), .Z(n23273) );
  XNOR U38799 ( .A(q[14]), .B(DB[2009]), .Z(n23262) );
  IV U38800 ( .A(n23261), .Z(n37629) );
  XNOR U38801 ( .A(n23259), .B(n37630), .Z(n23261) );
  XNOR U38802 ( .A(q[13]), .B(DB[2008]), .Z(n37630) );
  XNOR U38803 ( .A(q[12]), .B(DB[2007]), .Z(n23259) );
  IV U38804 ( .A(n23272), .Z(n37628) );
  XOR U38805 ( .A(n37631), .B(n37632), .Z(n23272) );
  XNOR U38806 ( .A(n23268), .B(n23270), .Z(n37632) );
  XNOR U38807 ( .A(q[8]), .B(DB[2003]), .Z(n23270) );
  XNOR U38808 ( .A(q[11]), .B(DB[2006]), .Z(n23268) );
  IV U38809 ( .A(n23267), .Z(n37631) );
  XNOR U38810 ( .A(n23265), .B(n37633), .Z(n23267) );
  XNOR U38811 ( .A(q[10]), .B(DB[2005]), .Z(n37633) );
  XNOR U38812 ( .A(q[9]), .B(DB[2004]), .Z(n23265) );
  IV U38813 ( .A(n23280), .Z(n37627) );
  XOR U38814 ( .A(n37634), .B(n37635), .Z(n23280) );
  XNOR U38815 ( .A(n23297), .B(n23278), .Z(n37635) );
  XNOR U38816 ( .A(q[0]), .B(DB[1995]), .Z(n23278) );
  XOR U38817 ( .A(n37636), .B(n23286), .Z(n23297) );
  XNOR U38818 ( .A(q[7]), .B(DB[2002]), .Z(n23286) );
  IV U38819 ( .A(n23285), .Z(n37636) );
  XNOR U38820 ( .A(n23283), .B(n37637), .Z(n23285) );
  XNOR U38821 ( .A(q[6]), .B(DB[2001]), .Z(n37637) );
  XNOR U38822 ( .A(q[5]), .B(DB[2000]), .Z(n23283) );
  IV U38823 ( .A(n23296), .Z(n37634) );
  XOR U38824 ( .A(n37638), .B(n37639), .Z(n23296) );
  XNOR U38825 ( .A(n23292), .B(n23294), .Z(n37639) );
  XNOR U38826 ( .A(q[1]), .B(DB[1996]), .Z(n23294) );
  XNOR U38827 ( .A(q[4]), .B(DB[1999]), .Z(n23292) );
  IV U38828 ( .A(n23291), .Z(n37638) );
  XNOR U38829 ( .A(n23289), .B(n37640), .Z(n23291) );
  XNOR U38830 ( .A(q[3]), .B(DB[1998]), .Z(n37640) );
  XNOR U38831 ( .A(q[2]), .B(DB[1997]), .Z(n23289) );
  XOR U38832 ( .A(n37641), .B(n23187), .Z(n23115) );
  XOR U38833 ( .A(n37642), .B(n23179), .Z(n23187) );
  XOR U38834 ( .A(n37643), .B(n23168), .Z(n23179) );
  XNOR U38835 ( .A(q[14]), .B(DB[2024]), .Z(n23168) );
  IV U38836 ( .A(n23167), .Z(n37643) );
  XNOR U38837 ( .A(n23165), .B(n37644), .Z(n23167) );
  XNOR U38838 ( .A(q[13]), .B(DB[2023]), .Z(n37644) );
  XNOR U38839 ( .A(q[12]), .B(DB[2022]), .Z(n23165) );
  IV U38840 ( .A(n23178), .Z(n37642) );
  XOR U38841 ( .A(n37645), .B(n37646), .Z(n23178) );
  XNOR U38842 ( .A(n23174), .B(n23176), .Z(n37646) );
  XNOR U38843 ( .A(q[8]), .B(DB[2018]), .Z(n23176) );
  XNOR U38844 ( .A(q[11]), .B(DB[2021]), .Z(n23174) );
  IV U38845 ( .A(n23173), .Z(n37645) );
  XNOR U38846 ( .A(n23171), .B(n37647), .Z(n23173) );
  XNOR U38847 ( .A(q[10]), .B(DB[2020]), .Z(n37647) );
  XNOR U38848 ( .A(q[9]), .B(DB[2019]), .Z(n23171) );
  IV U38849 ( .A(n23186), .Z(n37641) );
  XOR U38850 ( .A(n37648), .B(n37649), .Z(n23186) );
  XNOR U38851 ( .A(n23203), .B(n23184), .Z(n37649) );
  XNOR U38852 ( .A(q[0]), .B(DB[2010]), .Z(n23184) );
  XOR U38853 ( .A(n37650), .B(n23192), .Z(n23203) );
  XNOR U38854 ( .A(q[7]), .B(DB[2017]), .Z(n23192) );
  IV U38855 ( .A(n23191), .Z(n37650) );
  XNOR U38856 ( .A(n23189), .B(n37651), .Z(n23191) );
  XNOR U38857 ( .A(q[6]), .B(DB[2016]), .Z(n37651) );
  XNOR U38858 ( .A(q[5]), .B(DB[2015]), .Z(n23189) );
  IV U38859 ( .A(n23202), .Z(n37648) );
  XOR U38860 ( .A(n37652), .B(n37653), .Z(n23202) );
  XNOR U38861 ( .A(n23198), .B(n23200), .Z(n37653) );
  XNOR U38862 ( .A(q[1]), .B(DB[2011]), .Z(n23200) );
  XNOR U38863 ( .A(q[4]), .B(DB[2014]), .Z(n23198) );
  IV U38864 ( .A(n23197), .Z(n37652) );
  XNOR U38865 ( .A(n23195), .B(n37654), .Z(n23197) );
  XNOR U38866 ( .A(q[3]), .B(DB[2013]), .Z(n37654) );
  XNOR U38867 ( .A(q[2]), .B(DB[2012]), .Z(n23195) );
  XOR U38868 ( .A(n37655), .B(n23093), .Z(n23021) );
  XOR U38869 ( .A(n37656), .B(n23085), .Z(n23093) );
  XOR U38870 ( .A(n37657), .B(n23074), .Z(n23085) );
  XNOR U38871 ( .A(q[14]), .B(DB[2039]), .Z(n23074) );
  IV U38872 ( .A(n23073), .Z(n37657) );
  XNOR U38873 ( .A(n23071), .B(n37658), .Z(n23073) );
  XNOR U38874 ( .A(q[13]), .B(DB[2038]), .Z(n37658) );
  XNOR U38875 ( .A(q[12]), .B(DB[2037]), .Z(n23071) );
  IV U38876 ( .A(n23084), .Z(n37656) );
  XOR U38877 ( .A(n37659), .B(n37660), .Z(n23084) );
  XNOR U38878 ( .A(n23080), .B(n23082), .Z(n37660) );
  XNOR U38879 ( .A(q[8]), .B(DB[2033]), .Z(n23082) );
  XNOR U38880 ( .A(q[11]), .B(DB[2036]), .Z(n23080) );
  IV U38881 ( .A(n23079), .Z(n37659) );
  XNOR U38882 ( .A(n23077), .B(n37661), .Z(n23079) );
  XNOR U38883 ( .A(q[10]), .B(DB[2035]), .Z(n37661) );
  XNOR U38884 ( .A(q[9]), .B(DB[2034]), .Z(n23077) );
  IV U38885 ( .A(n23092), .Z(n37655) );
  XOR U38886 ( .A(n37662), .B(n37663), .Z(n23092) );
  XNOR U38887 ( .A(n23109), .B(n23090), .Z(n37663) );
  XNOR U38888 ( .A(q[0]), .B(DB[2025]), .Z(n23090) );
  XOR U38889 ( .A(n37664), .B(n23098), .Z(n23109) );
  XNOR U38890 ( .A(q[7]), .B(DB[2032]), .Z(n23098) );
  IV U38891 ( .A(n23097), .Z(n37664) );
  XNOR U38892 ( .A(n23095), .B(n37665), .Z(n23097) );
  XNOR U38893 ( .A(q[6]), .B(DB[2031]), .Z(n37665) );
  XNOR U38894 ( .A(q[5]), .B(DB[2030]), .Z(n23095) );
  IV U38895 ( .A(n23108), .Z(n37662) );
  XOR U38896 ( .A(n37666), .B(n37667), .Z(n23108) );
  XNOR U38897 ( .A(n23104), .B(n23106), .Z(n37667) );
  XNOR U38898 ( .A(q[1]), .B(DB[2026]), .Z(n23106) );
  XNOR U38899 ( .A(q[4]), .B(DB[2029]), .Z(n23104) );
  IV U38900 ( .A(n23103), .Z(n37666) );
  XNOR U38901 ( .A(n23101), .B(n37668), .Z(n23103) );
  XNOR U38902 ( .A(q[3]), .B(DB[2028]), .Z(n37668) );
  XNOR U38903 ( .A(q[2]), .B(DB[2027]), .Z(n23101) );
  XOR U38904 ( .A(n37669), .B(n22999), .Z(n22927) );
  XOR U38905 ( .A(n37670), .B(n22991), .Z(n22999) );
  XOR U38906 ( .A(n37671), .B(n22980), .Z(n22991) );
  XNOR U38907 ( .A(q[14]), .B(DB[2054]), .Z(n22980) );
  IV U38908 ( .A(n22979), .Z(n37671) );
  XNOR U38909 ( .A(n22977), .B(n37672), .Z(n22979) );
  XNOR U38910 ( .A(q[13]), .B(DB[2053]), .Z(n37672) );
  XNOR U38911 ( .A(q[12]), .B(DB[2052]), .Z(n22977) );
  IV U38912 ( .A(n22990), .Z(n37670) );
  XOR U38913 ( .A(n37673), .B(n37674), .Z(n22990) );
  XNOR U38914 ( .A(n22986), .B(n22988), .Z(n37674) );
  XNOR U38915 ( .A(q[8]), .B(DB[2048]), .Z(n22988) );
  XNOR U38916 ( .A(q[11]), .B(DB[2051]), .Z(n22986) );
  IV U38917 ( .A(n22985), .Z(n37673) );
  XNOR U38918 ( .A(n22983), .B(n37675), .Z(n22985) );
  XNOR U38919 ( .A(q[10]), .B(DB[2050]), .Z(n37675) );
  XNOR U38920 ( .A(q[9]), .B(DB[2049]), .Z(n22983) );
  IV U38921 ( .A(n22998), .Z(n37669) );
  XOR U38922 ( .A(n37676), .B(n37677), .Z(n22998) );
  XNOR U38923 ( .A(n23015), .B(n22996), .Z(n37677) );
  XNOR U38924 ( .A(q[0]), .B(DB[2040]), .Z(n22996) );
  XOR U38925 ( .A(n37678), .B(n23004), .Z(n23015) );
  XNOR U38926 ( .A(q[7]), .B(DB[2047]), .Z(n23004) );
  IV U38927 ( .A(n23003), .Z(n37678) );
  XNOR U38928 ( .A(n23001), .B(n37679), .Z(n23003) );
  XNOR U38929 ( .A(q[6]), .B(DB[2046]), .Z(n37679) );
  XNOR U38930 ( .A(q[5]), .B(DB[2045]), .Z(n23001) );
  IV U38931 ( .A(n23014), .Z(n37676) );
  XOR U38932 ( .A(n37680), .B(n37681), .Z(n23014) );
  XNOR U38933 ( .A(n23010), .B(n23012), .Z(n37681) );
  XNOR U38934 ( .A(q[1]), .B(DB[2041]), .Z(n23012) );
  XNOR U38935 ( .A(q[4]), .B(DB[2044]), .Z(n23010) );
  IV U38936 ( .A(n23009), .Z(n37680) );
  XNOR U38937 ( .A(n23007), .B(n37682), .Z(n23009) );
  XNOR U38938 ( .A(q[3]), .B(DB[2043]), .Z(n37682) );
  XNOR U38939 ( .A(q[2]), .B(DB[2042]), .Z(n23007) );
  XOR U38940 ( .A(n37683), .B(n22905), .Z(n22833) );
  XOR U38941 ( .A(n37684), .B(n22897), .Z(n22905) );
  XOR U38942 ( .A(n37685), .B(n22886), .Z(n22897) );
  XNOR U38943 ( .A(q[14]), .B(DB[2069]), .Z(n22886) );
  IV U38944 ( .A(n22885), .Z(n37685) );
  XNOR U38945 ( .A(n22883), .B(n37686), .Z(n22885) );
  XNOR U38946 ( .A(q[13]), .B(DB[2068]), .Z(n37686) );
  XNOR U38947 ( .A(q[12]), .B(DB[2067]), .Z(n22883) );
  IV U38948 ( .A(n22896), .Z(n37684) );
  XOR U38949 ( .A(n37687), .B(n37688), .Z(n22896) );
  XNOR U38950 ( .A(n22892), .B(n22894), .Z(n37688) );
  XNOR U38951 ( .A(q[8]), .B(DB[2063]), .Z(n22894) );
  XNOR U38952 ( .A(q[11]), .B(DB[2066]), .Z(n22892) );
  IV U38953 ( .A(n22891), .Z(n37687) );
  XNOR U38954 ( .A(n22889), .B(n37689), .Z(n22891) );
  XNOR U38955 ( .A(q[10]), .B(DB[2065]), .Z(n37689) );
  XNOR U38956 ( .A(q[9]), .B(DB[2064]), .Z(n22889) );
  IV U38957 ( .A(n22904), .Z(n37683) );
  XOR U38958 ( .A(n37690), .B(n37691), .Z(n22904) );
  XNOR U38959 ( .A(n22921), .B(n22902), .Z(n37691) );
  XNOR U38960 ( .A(q[0]), .B(DB[2055]), .Z(n22902) );
  XOR U38961 ( .A(n37692), .B(n22910), .Z(n22921) );
  XNOR U38962 ( .A(q[7]), .B(DB[2062]), .Z(n22910) );
  IV U38963 ( .A(n22909), .Z(n37692) );
  XNOR U38964 ( .A(n22907), .B(n37693), .Z(n22909) );
  XNOR U38965 ( .A(q[6]), .B(DB[2061]), .Z(n37693) );
  XNOR U38966 ( .A(q[5]), .B(DB[2060]), .Z(n22907) );
  IV U38967 ( .A(n22920), .Z(n37690) );
  XOR U38968 ( .A(n37694), .B(n37695), .Z(n22920) );
  XNOR U38969 ( .A(n22916), .B(n22918), .Z(n37695) );
  XNOR U38970 ( .A(q[1]), .B(DB[2056]), .Z(n22918) );
  XNOR U38971 ( .A(q[4]), .B(DB[2059]), .Z(n22916) );
  IV U38972 ( .A(n22915), .Z(n37694) );
  XNOR U38973 ( .A(n22913), .B(n37696), .Z(n22915) );
  XNOR U38974 ( .A(q[3]), .B(DB[2058]), .Z(n37696) );
  XNOR U38975 ( .A(q[2]), .B(DB[2057]), .Z(n22913) );
  XOR U38976 ( .A(n37697), .B(n22811), .Z(n22739) );
  XOR U38977 ( .A(n37698), .B(n22803), .Z(n22811) );
  XOR U38978 ( .A(n37699), .B(n22792), .Z(n22803) );
  XNOR U38979 ( .A(q[14]), .B(DB[2084]), .Z(n22792) );
  IV U38980 ( .A(n22791), .Z(n37699) );
  XNOR U38981 ( .A(n22789), .B(n37700), .Z(n22791) );
  XNOR U38982 ( .A(q[13]), .B(DB[2083]), .Z(n37700) );
  XNOR U38983 ( .A(q[12]), .B(DB[2082]), .Z(n22789) );
  IV U38984 ( .A(n22802), .Z(n37698) );
  XOR U38985 ( .A(n37701), .B(n37702), .Z(n22802) );
  XNOR U38986 ( .A(n22798), .B(n22800), .Z(n37702) );
  XNOR U38987 ( .A(q[8]), .B(DB[2078]), .Z(n22800) );
  XNOR U38988 ( .A(q[11]), .B(DB[2081]), .Z(n22798) );
  IV U38989 ( .A(n22797), .Z(n37701) );
  XNOR U38990 ( .A(n22795), .B(n37703), .Z(n22797) );
  XNOR U38991 ( .A(q[10]), .B(DB[2080]), .Z(n37703) );
  XNOR U38992 ( .A(q[9]), .B(DB[2079]), .Z(n22795) );
  IV U38993 ( .A(n22810), .Z(n37697) );
  XOR U38994 ( .A(n37704), .B(n37705), .Z(n22810) );
  XNOR U38995 ( .A(n22827), .B(n22808), .Z(n37705) );
  XNOR U38996 ( .A(q[0]), .B(DB[2070]), .Z(n22808) );
  XOR U38997 ( .A(n37706), .B(n22816), .Z(n22827) );
  XNOR U38998 ( .A(q[7]), .B(DB[2077]), .Z(n22816) );
  IV U38999 ( .A(n22815), .Z(n37706) );
  XNOR U39000 ( .A(n22813), .B(n37707), .Z(n22815) );
  XNOR U39001 ( .A(q[6]), .B(DB[2076]), .Z(n37707) );
  XNOR U39002 ( .A(q[5]), .B(DB[2075]), .Z(n22813) );
  IV U39003 ( .A(n22826), .Z(n37704) );
  XOR U39004 ( .A(n37708), .B(n37709), .Z(n22826) );
  XNOR U39005 ( .A(n22822), .B(n22824), .Z(n37709) );
  XNOR U39006 ( .A(q[1]), .B(DB[2071]), .Z(n22824) );
  XNOR U39007 ( .A(q[4]), .B(DB[2074]), .Z(n22822) );
  IV U39008 ( .A(n22821), .Z(n37708) );
  XNOR U39009 ( .A(n22819), .B(n37710), .Z(n22821) );
  XNOR U39010 ( .A(q[3]), .B(DB[2073]), .Z(n37710) );
  XNOR U39011 ( .A(q[2]), .B(DB[2072]), .Z(n22819) );
  XOR U39012 ( .A(n37711), .B(n22717), .Z(n22645) );
  XOR U39013 ( .A(n37712), .B(n22709), .Z(n22717) );
  XOR U39014 ( .A(n37713), .B(n22698), .Z(n22709) );
  XNOR U39015 ( .A(q[14]), .B(DB[2099]), .Z(n22698) );
  IV U39016 ( .A(n22697), .Z(n37713) );
  XNOR U39017 ( .A(n22695), .B(n37714), .Z(n22697) );
  XNOR U39018 ( .A(q[13]), .B(DB[2098]), .Z(n37714) );
  XNOR U39019 ( .A(q[12]), .B(DB[2097]), .Z(n22695) );
  IV U39020 ( .A(n22708), .Z(n37712) );
  XOR U39021 ( .A(n37715), .B(n37716), .Z(n22708) );
  XNOR U39022 ( .A(n22704), .B(n22706), .Z(n37716) );
  XNOR U39023 ( .A(q[8]), .B(DB[2093]), .Z(n22706) );
  XNOR U39024 ( .A(q[11]), .B(DB[2096]), .Z(n22704) );
  IV U39025 ( .A(n22703), .Z(n37715) );
  XNOR U39026 ( .A(n22701), .B(n37717), .Z(n22703) );
  XNOR U39027 ( .A(q[10]), .B(DB[2095]), .Z(n37717) );
  XNOR U39028 ( .A(q[9]), .B(DB[2094]), .Z(n22701) );
  IV U39029 ( .A(n22716), .Z(n37711) );
  XOR U39030 ( .A(n37718), .B(n37719), .Z(n22716) );
  XNOR U39031 ( .A(n22733), .B(n22714), .Z(n37719) );
  XNOR U39032 ( .A(q[0]), .B(DB[2085]), .Z(n22714) );
  XOR U39033 ( .A(n37720), .B(n22722), .Z(n22733) );
  XNOR U39034 ( .A(q[7]), .B(DB[2092]), .Z(n22722) );
  IV U39035 ( .A(n22721), .Z(n37720) );
  XNOR U39036 ( .A(n22719), .B(n37721), .Z(n22721) );
  XNOR U39037 ( .A(q[6]), .B(DB[2091]), .Z(n37721) );
  XNOR U39038 ( .A(q[5]), .B(DB[2090]), .Z(n22719) );
  IV U39039 ( .A(n22732), .Z(n37718) );
  XOR U39040 ( .A(n37722), .B(n37723), .Z(n22732) );
  XNOR U39041 ( .A(n22728), .B(n22730), .Z(n37723) );
  XNOR U39042 ( .A(q[1]), .B(DB[2086]), .Z(n22730) );
  XNOR U39043 ( .A(q[4]), .B(DB[2089]), .Z(n22728) );
  IV U39044 ( .A(n22727), .Z(n37722) );
  XNOR U39045 ( .A(n22725), .B(n37724), .Z(n22727) );
  XNOR U39046 ( .A(q[3]), .B(DB[2088]), .Z(n37724) );
  XNOR U39047 ( .A(q[2]), .B(DB[2087]), .Z(n22725) );
  XOR U39048 ( .A(n37725), .B(n22623), .Z(n22551) );
  XOR U39049 ( .A(n37726), .B(n22615), .Z(n22623) );
  XOR U39050 ( .A(n37727), .B(n22604), .Z(n22615) );
  XNOR U39051 ( .A(q[14]), .B(DB[2114]), .Z(n22604) );
  IV U39052 ( .A(n22603), .Z(n37727) );
  XNOR U39053 ( .A(n22601), .B(n37728), .Z(n22603) );
  XNOR U39054 ( .A(q[13]), .B(DB[2113]), .Z(n37728) );
  XNOR U39055 ( .A(q[12]), .B(DB[2112]), .Z(n22601) );
  IV U39056 ( .A(n22614), .Z(n37726) );
  XOR U39057 ( .A(n37729), .B(n37730), .Z(n22614) );
  XNOR U39058 ( .A(n22610), .B(n22612), .Z(n37730) );
  XNOR U39059 ( .A(q[8]), .B(DB[2108]), .Z(n22612) );
  XNOR U39060 ( .A(q[11]), .B(DB[2111]), .Z(n22610) );
  IV U39061 ( .A(n22609), .Z(n37729) );
  XNOR U39062 ( .A(n22607), .B(n37731), .Z(n22609) );
  XNOR U39063 ( .A(q[10]), .B(DB[2110]), .Z(n37731) );
  XNOR U39064 ( .A(q[9]), .B(DB[2109]), .Z(n22607) );
  IV U39065 ( .A(n22622), .Z(n37725) );
  XOR U39066 ( .A(n37732), .B(n37733), .Z(n22622) );
  XNOR U39067 ( .A(n22639), .B(n22620), .Z(n37733) );
  XNOR U39068 ( .A(q[0]), .B(DB[2100]), .Z(n22620) );
  XOR U39069 ( .A(n37734), .B(n22628), .Z(n22639) );
  XNOR U39070 ( .A(q[7]), .B(DB[2107]), .Z(n22628) );
  IV U39071 ( .A(n22627), .Z(n37734) );
  XNOR U39072 ( .A(n22625), .B(n37735), .Z(n22627) );
  XNOR U39073 ( .A(q[6]), .B(DB[2106]), .Z(n37735) );
  XNOR U39074 ( .A(q[5]), .B(DB[2105]), .Z(n22625) );
  IV U39075 ( .A(n22638), .Z(n37732) );
  XOR U39076 ( .A(n37736), .B(n37737), .Z(n22638) );
  XNOR U39077 ( .A(n22634), .B(n22636), .Z(n37737) );
  XNOR U39078 ( .A(q[1]), .B(DB[2101]), .Z(n22636) );
  XNOR U39079 ( .A(q[4]), .B(DB[2104]), .Z(n22634) );
  IV U39080 ( .A(n22633), .Z(n37736) );
  XNOR U39081 ( .A(n22631), .B(n37738), .Z(n22633) );
  XNOR U39082 ( .A(q[3]), .B(DB[2103]), .Z(n37738) );
  XNOR U39083 ( .A(q[2]), .B(DB[2102]), .Z(n22631) );
  XOR U39084 ( .A(n37739), .B(n22529), .Z(n22457) );
  XOR U39085 ( .A(n37740), .B(n22521), .Z(n22529) );
  XOR U39086 ( .A(n37741), .B(n22510), .Z(n22521) );
  XNOR U39087 ( .A(q[14]), .B(DB[2129]), .Z(n22510) );
  IV U39088 ( .A(n22509), .Z(n37741) );
  XNOR U39089 ( .A(n22507), .B(n37742), .Z(n22509) );
  XNOR U39090 ( .A(q[13]), .B(DB[2128]), .Z(n37742) );
  XNOR U39091 ( .A(q[12]), .B(DB[2127]), .Z(n22507) );
  IV U39092 ( .A(n22520), .Z(n37740) );
  XOR U39093 ( .A(n37743), .B(n37744), .Z(n22520) );
  XNOR U39094 ( .A(n22516), .B(n22518), .Z(n37744) );
  XNOR U39095 ( .A(q[8]), .B(DB[2123]), .Z(n22518) );
  XNOR U39096 ( .A(q[11]), .B(DB[2126]), .Z(n22516) );
  IV U39097 ( .A(n22515), .Z(n37743) );
  XNOR U39098 ( .A(n22513), .B(n37745), .Z(n22515) );
  XNOR U39099 ( .A(q[10]), .B(DB[2125]), .Z(n37745) );
  XNOR U39100 ( .A(q[9]), .B(DB[2124]), .Z(n22513) );
  IV U39101 ( .A(n22528), .Z(n37739) );
  XOR U39102 ( .A(n37746), .B(n37747), .Z(n22528) );
  XNOR U39103 ( .A(n22545), .B(n22526), .Z(n37747) );
  XNOR U39104 ( .A(q[0]), .B(DB[2115]), .Z(n22526) );
  XOR U39105 ( .A(n37748), .B(n22534), .Z(n22545) );
  XNOR U39106 ( .A(q[7]), .B(DB[2122]), .Z(n22534) );
  IV U39107 ( .A(n22533), .Z(n37748) );
  XNOR U39108 ( .A(n22531), .B(n37749), .Z(n22533) );
  XNOR U39109 ( .A(q[6]), .B(DB[2121]), .Z(n37749) );
  XNOR U39110 ( .A(q[5]), .B(DB[2120]), .Z(n22531) );
  IV U39111 ( .A(n22544), .Z(n37746) );
  XOR U39112 ( .A(n37750), .B(n37751), .Z(n22544) );
  XNOR U39113 ( .A(n22540), .B(n22542), .Z(n37751) );
  XNOR U39114 ( .A(q[1]), .B(DB[2116]), .Z(n22542) );
  XNOR U39115 ( .A(q[4]), .B(DB[2119]), .Z(n22540) );
  IV U39116 ( .A(n22539), .Z(n37750) );
  XNOR U39117 ( .A(n22537), .B(n37752), .Z(n22539) );
  XNOR U39118 ( .A(q[3]), .B(DB[2118]), .Z(n37752) );
  XNOR U39119 ( .A(q[2]), .B(DB[2117]), .Z(n22537) );
  XOR U39120 ( .A(n37753), .B(n22435), .Z(n22363) );
  XOR U39121 ( .A(n37754), .B(n22427), .Z(n22435) );
  XOR U39122 ( .A(n37755), .B(n22416), .Z(n22427) );
  XNOR U39123 ( .A(q[14]), .B(DB[2144]), .Z(n22416) );
  IV U39124 ( .A(n22415), .Z(n37755) );
  XNOR U39125 ( .A(n22413), .B(n37756), .Z(n22415) );
  XNOR U39126 ( .A(q[13]), .B(DB[2143]), .Z(n37756) );
  XNOR U39127 ( .A(q[12]), .B(DB[2142]), .Z(n22413) );
  IV U39128 ( .A(n22426), .Z(n37754) );
  XOR U39129 ( .A(n37757), .B(n37758), .Z(n22426) );
  XNOR U39130 ( .A(n22422), .B(n22424), .Z(n37758) );
  XNOR U39131 ( .A(q[8]), .B(DB[2138]), .Z(n22424) );
  XNOR U39132 ( .A(q[11]), .B(DB[2141]), .Z(n22422) );
  IV U39133 ( .A(n22421), .Z(n37757) );
  XNOR U39134 ( .A(n22419), .B(n37759), .Z(n22421) );
  XNOR U39135 ( .A(q[10]), .B(DB[2140]), .Z(n37759) );
  XNOR U39136 ( .A(q[9]), .B(DB[2139]), .Z(n22419) );
  IV U39137 ( .A(n22434), .Z(n37753) );
  XOR U39138 ( .A(n37760), .B(n37761), .Z(n22434) );
  XNOR U39139 ( .A(n22451), .B(n22432), .Z(n37761) );
  XNOR U39140 ( .A(q[0]), .B(DB[2130]), .Z(n22432) );
  XOR U39141 ( .A(n37762), .B(n22440), .Z(n22451) );
  XNOR U39142 ( .A(q[7]), .B(DB[2137]), .Z(n22440) );
  IV U39143 ( .A(n22439), .Z(n37762) );
  XNOR U39144 ( .A(n22437), .B(n37763), .Z(n22439) );
  XNOR U39145 ( .A(q[6]), .B(DB[2136]), .Z(n37763) );
  XNOR U39146 ( .A(q[5]), .B(DB[2135]), .Z(n22437) );
  IV U39147 ( .A(n22450), .Z(n37760) );
  XOR U39148 ( .A(n37764), .B(n37765), .Z(n22450) );
  XNOR U39149 ( .A(n22446), .B(n22448), .Z(n37765) );
  XNOR U39150 ( .A(q[1]), .B(DB[2131]), .Z(n22448) );
  XNOR U39151 ( .A(q[4]), .B(DB[2134]), .Z(n22446) );
  IV U39152 ( .A(n22445), .Z(n37764) );
  XNOR U39153 ( .A(n22443), .B(n37766), .Z(n22445) );
  XNOR U39154 ( .A(q[3]), .B(DB[2133]), .Z(n37766) );
  XNOR U39155 ( .A(q[2]), .B(DB[2132]), .Z(n22443) );
  XOR U39156 ( .A(n37767), .B(n22341), .Z(n22269) );
  XOR U39157 ( .A(n37768), .B(n22333), .Z(n22341) );
  XOR U39158 ( .A(n37769), .B(n22322), .Z(n22333) );
  XNOR U39159 ( .A(q[14]), .B(DB[2159]), .Z(n22322) );
  IV U39160 ( .A(n22321), .Z(n37769) );
  XNOR U39161 ( .A(n22319), .B(n37770), .Z(n22321) );
  XNOR U39162 ( .A(q[13]), .B(DB[2158]), .Z(n37770) );
  XNOR U39163 ( .A(q[12]), .B(DB[2157]), .Z(n22319) );
  IV U39164 ( .A(n22332), .Z(n37768) );
  XOR U39165 ( .A(n37771), .B(n37772), .Z(n22332) );
  XNOR U39166 ( .A(n22328), .B(n22330), .Z(n37772) );
  XNOR U39167 ( .A(q[8]), .B(DB[2153]), .Z(n22330) );
  XNOR U39168 ( .A(q[11]), .B(DB[2156]), .Z(n22328) );
  IV U39169 ( .A(n22327), .Z(n37771) );
  XNOR U39170 ( .A(n22325), .B(n37773), .Z(n22327) );
  XNOR U39171 ( .A(q[10]), .B(DB[2155]), .Z(n37773) );
  XNOR U39172 ( .A(q[9]), .B(DB[2154]), .Z(n22325) );
  IV U39173 ( .A(n22340), .Z(n37767) );
  XOR U39174 ( .A(n37774), .B(n37775), .Z(n22340) );
  XNOR U39175 ( .A(n22357), .B(n22338), .Z(n37775) );
  XNOR U39176 ( .A(q[0]), .B(DB[2145]), .Z(n22338) );
  XOR U39177 ( .A(n37776), .B(n22346), .Z(n22357) );
  XNOR U39178 ( .A(q[7]), .B(DB[2152]), .Z(n22346) );
  IV U39179 ( .A(n22345), .Z(n37776) );
  XNOR U39180 ( .A(n22343), .B(n37777), .Z(n22345) );
  XNOR U39181 ( .A(q[6]), .B(DB[2151]), .Z(n37777) );
  XNOR U39182 ( .A(q[5]), .B(DB[2150]), .Z(n22343) );
  IV U39183 ( .A(n22356), .Z(n37774) );
  XOR U39184 ( .A(n37778), .B(n37779), .Z(n22356) );
  XNOR U39185 ( .A(n22352), .B(n22354), .Z(n37779) );
  XNOR U39186 ( .A(q[1]), .B(DB[2146]), .Z(n22354) );
  XNOR U39187 ( .A(q[4]), .B(DB[2149]), .Z(n22352) );
  IV U39188 ( .A(n22351), .Z(n37778) );
  XNOR U39189 ( .A(n22349), .B(n37780), .Z(n22351) );
  XNOR U39190 ( .A(q[3]), .B(DB[2148]), .Z(n37780) );
  XNOR U39191 ( .A(q[2]), .B(DB[2147]), .Z(n22349) );
  XOR U39192 ( .A(n37781), .B(n22247), .Z(n22175) );
  XOR U39193 ( .A(n37782), .B(n22239), .Z(n22247) );
  XOR U39194 ( .A(n37783), .B(n22228), .Z(n22239) );
  XNOR U39195 ( .A(q[14]), .B(DB[2174]), .Z(n22228) );
  IV U39196 ( .A(n22227), .Z(n37783) );
  XNOR U39197 ( .A(n22225), .B(n37784), .Z(n22227) );
  XNOR U39198 ( .A(q[13]), .B(DB[2173]), .Z(n37784) );
  XNOR U39199 ( .A(q[12]), .B(DB[2172]), .Z(n22225) );
  IV U39200 ( .A(n22238), .Z(n37782) );
  XOR U39201 ( .A(n37785), .B(n37786), .Z(n22238) );
  XNOR U39202 ( .A(n22234), .B(n22236), .Z(n37786) );
  XNOR U39203 ( .A(q[8]), .B(DB[2168]), .Z(n22236) );
  XNOR U39204 ( .A(q[11]), .B(DB[2171]), .Z(n22234) );
  IV U39205 ( .A(n22233), .Z(n37785) );
  XNOR U39206 ( .A(n22231), .B(n37787), .Z(n22233) );
  XNOR U39207 ( .A(q[10]), .B(DB[2170]), .Z(n37787) );
  XNOR U39208 ( .A(q[9]), .B(DB[2169]), .Z(n22231) );
  IV U39209 ( .A(n22246), .Z(n37781) );
  XOR U39210 ( .A(n37788), .B(n37789), .Z(n22246) );
  XNOR U39211 ( .A(n22263), .B(n22244), .Z(n37789) );
  XNOR U39212 ( .A(q[0]), .B(DB[2160]), .Z(n22244) );
  XOR U39213 ( .A(n37790), .B(n22252), .Z(n22263) );
  XNOR U39214 ( .A(q[7]), .B(DB[2167]), .Z(n22252) );
  IV U39215 ( .A(n22251), .Z(n37790) );
  XNOR U39216 ( .A(n22249), .B(n37791), .Z(n22251) );
  XNOR U39217 ( .A(q[6]), .B(DB[2166]), .Z(n37791) );
  XNOR U39218 ( .A(q[5]), .B(DB[2165]), .Z(n22249) );
  IV U39219 ( .A(n22262), .Z(n37788) );
  XOR U39220 ( .A(n37792), .B(n37793), .Z(n22262) );
  XNOR U39221 ( .A(n22258), .B(n22260), .Z(n37793) );
  XNOR U39222 ( .A(q[1]), .B(DB[2161]), .Z(n22260) );
  XNOR U39223 ( .A(q[4]), .B(DB[2164]), .Z(n22258) );
  IV U39224 ( .A(n22257), .Z(n37792) );
  XNOR U39225 ( .A(n22255), .B(n37794), .Z(n22257) );
  XNOR U39226 ( .A(q[3]), .B(DB[2163]), .Z(n37794) );
  XNOR U39227 ( .A(q[2]), .B(DB[2162]), .Z(n22255) );
  XOR U39228 ( .A(n37795), .B(n22153), .Z(n22081) );
  XOR U39229 ( .A(n37796), .B(n22145), .Z(n22153) );
  XOR U39230 ( .A(n37797), .B(n22134), .Z(n22145) );
  XNOR U39231 ( .A(q[14]), .B(DB[2189]), .Z(n22134) );
  IV U39232 ( .A(n22133), .Z(n37797) );
  XNOR U39233 ( .A(n22131), .B(n37798), .Z(n22133) );
  XNOR U39234 ( .A(q[13]), .B(DB[2188]), .Z(n37798) );
  XNOR U39235 ( .A(q[12]), .B(DB[2187]), .Z(n22131) );
  IV U39236 ( .A(n22144), .Z(n37796) );
  XOR U39237 ( .A(n37799), .B(n37800), .Z(n22144) );
  XNOR U39238 ( .A(n22140), .B(n22142), .Z(n37800) );
  XNOR U39239 ( .A(q[8]), .B(DB[2183]), .Z(n22142) );
  XNOR U39240 ( .A(q[11]), .B(DB[2186]), .Z(n22140) );
  IV U39241 ( .A(n22139), .Z(n37799) );
  XNOR U39242 ( .A(n22137), .B(n37801), .Z(n22139) );
  XNOR U39243 ( .A(q[10]), .B(DB[2185]), .Z(n37801) );
  XNOR U39244 ( .A(q[9]), .B(DB[2184]), .Z(n22137) );
  IV U39245 ( .A(n22152), .Z(n37795) );
  XOR U39246 ( .A(n37802), .B(n37803), .Z(n22152) );
  XNOR U39247 ( .A(n22169), .B(n22150), .Z(n37803) );
  XNOR U39248 ( .A(q[0]), .B(DB[2175]), .Z(n22150) );
  XOR U39249 ( .A(n37804), .B(n22158), .Z(n22169) );
  XNOR U39250 ( .A(q[7]), .B(DB[2182]), .Z(n22158) );
  IV U39251 ( .A(n22157), .Z(n37804) );
  XNOR U39252 ( .A(n22155), .B(n37805), .Z(n22157) );
  XNOR U39253 ( .A(q[6]), .B(DB[2181]), .Z(n37805) );
  XNOR U39254 ( .A(q[5]), .B(DB[2180]), .Z(n22155) );
  IV U39255 ( .A(n22168), .Z(n37802) );
  XOR U39256 ( .A(n37806), .B(n37807), .Z(n22168) );
  XNOR U39257 ( .A(n22164), .B(n22166), .Z(n37807) );
  XNOR U39258 ( .A(q[1]), .B(DB[2176]), .Z(n22166) );
  XNOR U39259 ( .A(q[4]), .B(DB[2179]), .Z(n22164) );
  IV U39260 ( .A(n22163), .Z(n37806) );
  XNOR U39261 ( .A(n22161), .B(n37808), .Z(n22163) );
  XNOR U39262 ( .A(q[3]), .B(DB[2178]), .Z(n37808) );
  XNOR U39263 ( .A(q[2]), .B(DB[2177]), .Z(n22161) );
  XOR U39264 ( .A(n37809), .B(n22059), .Z(n21987) );
  XOR U39265 ( .A(n37810), .B(n22051), .Z(n22059) );
  XOR U39266 ( .A(n37811), .B(n22040), .Z(n22051) );
  XNOR U39267 ( .A(q[14]), .B(DB[2204]), .Z(n22040) );
  IV U39268 ( .A(n22039), .Z(n37811) );
  XNOR U39269 ( .A(n22037), .B(n37812), .Z(n22039) );
  XNOR U39270 ( .A(q[13]), .B(DB[2203]), .Z(n37812) );
  XNOR U39271 ( .A(q[12]), .B(DB[2202]), .Z(n22037) );
  IV U39272 ( .A(n22050), .Z(n37810) );
  XOR U39273 ( .A(n37813), .B(n37814), .Z(n22050) );
  XNOR U39274 ( .A(n22046), .B(n22048), .Z(n37814) );
  XNOR U39275 ( .A(q[8]), .B(DB[2198]), .Z(n22048) );
  XNOR U39276 ( .A(q[11]), .B(DB[2201]), .Z(n22046) );
  IV U39277 ( .A(n22045), .Z(n37813) );
  XNOR U39278 ( .A(n22043), .B(n37815), .Z(n22045) );
  XNOR U39279 ( .A(q[10]), .B(DB[2200]), .Z(n37815) );
  XNOR U39280 ( .A(q[9]), .B(DB[2199]), .Z(n22043) );
  IV U39281 ( .A(n22058), .Z(n37809) );
  XOR U39282 ( .A(n37816), .B(n37817), .Z(n22058) );
  XNOR U39283 ( .A(n22075), .B(n22056), .Z(n37817) );
  XNOR U39284 ( .A(q[0]), .B(DB[2190]), .Z(n22056) );
  XOR U39285 ( .A(n37818), .B(n22064), .Z(n22075) );
  XNOR U39286 ( .A(q[7]), .B(DB[2197]), .Z(n22064) );
  IV U39287 ( .A(n22063), .Z(n37818) );
  XNOR U39288 ( .A(n22061), .B(n37819), .Z(n22063) );
  XNOR U39289 ( .A(q[6]), .B(DB[2196]), .Z(n37819) );
  XNOR U39290 ( .A(q[5]), .B(DB[2195]), .Z(n22061) );
  IV U39291 ( .A(n22074), .Z(n37816) );
  XOR U39292 ( .A(n37820), .B(n37821), .Z(n22074) );
  XNOR U39293 ( .A(n22070), .B(n22072), .Z(n37821) );
  XNOR U39294 ( .A(q[1]), .B(DB[2191]), .Z(n22072) );
  XNOR U39295 ( .A(q[4]), .B(DB[2194]), .Z(n22070) );
  IV U39296 ( .A(n22069), .Z(n37820) );
  XNOR U39297 ( .A(n22067), .B(n37822), .Z(n22069) );
  XNOR U39298 ( .A(q[3]), .B(DB[2193]), .Z(n37822) );
  XNOR U39299 ( .A(q[2]), .B(DB[2192]), .Z(n22067) );
  XOR U39300 ( .A(n37823), .B(n21965), .Z(n21893) );
  XOR U39301 ( .A(n37824), .B(n21957), .Z(n21965) );
  XOR U39302 ( .A(n37825), .B(n21946), .Z(n21957) );
  XNOR U39303 ( .A(q[14]), .B(DB[2219]), .Z(n21946) );
  IV U39304 ( .A(n21945), .Z(n37825) );
  XNOR U39305 ( .A(n21943), .B(n37826), .Z(n21945) );
  XNOR U39306 ( .A(q[13]), .B(DB[2218]), .Z(n37826) );
  XNOR U39307 ( .A(q[12]), .B(DB[2217]), .Z(n21943) );
  IV U39308 ( .A(n21956), .Z(n37824) );
  XOR U39309 ( .A(n37827), .B(n37828), .Z(n21956) );
  XNOR U39310 ( .A(n21952), .B(n21954), .Z(n37828) );
  XNOR U39311 ( .A(q[8]), .B(DB[2213]), .Z(n21954) );
  XNOR U39312 ( .A(q[11]), .B(DB[2216]), .Z(n21952) );
  IV U39313 ( .A(n21951), .Z(n37827) );
  XNOR U39314 ( .A(n21949), .B(n37829), .Z(n21951) );
  XNOR U39315 ( .A(q[10]), .B(DB[2215]), .Z(n37829) );
  XNOR U39316 ( .A(q[9]), .B(DB[2214]), .Z(n21949) );
  IV U39317 ( .A(n21964), .Z(n37823) );
  XOR U39318 ( .A(n37830), .B(n37831), .Z(n21964) );
  XNOR U39319 ( .A(n21981), .B(n21962), .Z(n37831) );
  XNOR U39320 ( .A(q[0]), .B(DB[2205]), .Z(n21962) );
  XOR U39321 ( .A(n37832), .B(n21970), .Z(n21981) );
  XNOR U39322 ( .A(q[7]), .B(DB[2212]), .Z(n21970) );
  IV U39323 ( .A(n21969), .Z(n37832) );
  XNOR U39324 ( .A(n21967), .B(n37833), .Z(n21969) );
  XNOR U39325 ( .A(q[6]), .B(DB[2211]), .Z(n37833) );
  XNOR U39326 ( .A(q[5]), .B(DB[2210]), .Z(n21967) );
  IV U39327 ( .A(n21980), .Z(n37830) );
  XOR U39328 ( .A(n37834), .B(n37835), .Z(n21980) );
  XNOR U39329 ( .A(n21976), .B(n21978), .Z(n37835) );
  XNOR U39330 ( .A(q[1]), .B(DB[2206]), .Z(n21978) );
  XNOR U39331 ( .A(q[4]), .B(DB[2209]), .Z(n21976) );
  IV U39332 ( .A(n21975), .Z(n37834) );
  XNOR U39333 ( .A(n21973), .B(n37836), .Z(n21975) );
  XNOR U39334 ( .A(q[3]), .B(DB[2208]), .Z(n37836) );
  XNOR U39335 ( .A(q[2]), .B(DB[2207]), .Z(n21973) );
  XOR U39336 ( .A(n37837), .B(n21871), .Z(n21799) );
  XOR U39337 ( .A(n37838), .B(n21863), .Z(n21871) );
  XOR U39338 ( .A(n37839), .B(n21852), .Z(n21863) );
  XNOR U39339 ( .A(q[14]), .B(DB[2234]), .Z(n21852) );
  IV U39340 ( .A(n21851), .Z(n37839) );
  XNOR U39341 ( .A(n21849), .B(n37840), .Z(n21851) );
  XNOR U39342 ( .A(q[13]), .B(DB[2233]), .Z(n37840) );
  XNOR U39343 ( .A(q[12]), .B(DB[2232]), .Z(n21849) );
  IV U39344 ( .A(n21862), .Z(n37838) );
  XOR U39345 ( .A(n37841), .B(n37842), .Z(n21862) );
  XNOR U39346 ( .A(n21858), .B(n21860), .Z(n37842) );
  XNOR U39347 ( .A(q[8]), .B(DB[2228]), .Z(n21860) );
  XNOR U39348 ( .A(q[11]), .B(DB[2231]), .Z(n21858) );
  IV U39349 ( .A(n21857), .Z(n37841) );
  XNOR U39350 ( .A(n21855), .B(n37843), .Z(n21857) );
  XNOR U39351 ( .A(q[10]), .B(DB[2230]), .Z(n37843) );
  XNOR U39352 ( .A(q[9]), .B(DB[2229]), .Z(n21855) );
  IV U39353 ( .A(n21870), .Z(n37837) );
  XOR U39354 ( .A(n37844), .B(n37845), .Z(n21870) );
  XNOR U39355 ( .A(n21887), .B(n21868), .Z(n37845) );
  XNOR U39356 ( .A(q[0]), .B(DB[2220]), .Z(n21868) );
  XOR U39357 ( .A(n37846), .B(n21876), .Z(n21887) );
  XNOR U39358 ( .A(q[7]), .B(DB[2227]), .Z(n21876) );
  IV U39359 ( .A(n21875), .Z(n37846) );
  XNOR U39360 ( .A(n21873), .B(n37847), .Z(n21875) );
  XNOR U39361 ( .A(q[6]), .B(DB[2226]), .Z(n37847) );
  XNOR U39362 ( .A(q[5]), .B(DB[2225]), .Z(n21873) );
  IV U39363 ( .A(n21886), .Z(n37844) );
  XOR U39364 ( .A(n37848), .B(n37849), .Z(n21886) );
  XNOR U39365 ( .A(n21882), .B(n21884), .Z(n37849) );
  XNOR U39366 ( .A(q[1]), .B(DB[2221]), .Z(n21884) );
  XNOR U39367 ( .A(q[4]), .B(DB[2224]), .Z(n21882) );
  IV U39368 ( .A(n21881), .Z(n37848) );
  XNOR U39369 ( .A(n21879), .B(n37850), .Z(n21881) );
  XNOR U39370 ( .A(q[3]), .B(DB[2223]), .Z(n37850) );
  XNOR U39371 ( .A(q[2]), .B(DB[2222]), .Z(n21879) );
  XOR U39372 ( .A(n37851), .B(n21777), .Z(n21705) );
  XOR U39373 ( .A(n37852), .B(n21769), .Z(n21777) );
  XOR U39374 ( .A(n37853), .B(n21758), .Z(n21769) );
  XNOR U39375 ( .A(q[14]), .B(DB[2249]), .Z(n21758) );
  IV U39376 ( .A(n21757), .Z(n37853) );
  XNOR U39377 ( .A(n21755), .B(n37854), .Z(n21757) );
  XNOR U39378 ( .A(q[13]), .B(DB[2248]), .Z(n37854) );
  XNOR U39379 ( .A(q[12]), .B(DB[2247]), .Z(n21755) );
  IV U39380 ( .A(n21768), .Z(n37852) );
  XOR U39381 ( .A(n37855), .B(n37856), .Z(n21768) );
  XNOR U39382 ( .A(n21764), .B(n21766), .Z(n37856) );
  XNOR U39383 ( .A(q[8]), .B(DB[2243]), .Z(n21766) );
  XNOR U39384 ( .A(q[11]), .B(DB[2246]), .Z(n21764) );
  IV U39385 ( .A(n21763), .Z(n37855) );
  XNOR U39386 ( .A(n21761), .B(n37857), .Z(n21763) );
  XNOR U39387 ( .A(q[10]), .B(DB[2245]), .Z(n37857) );
  XNOR U39388 ( .A(q[9]), .B(DB[2244]), .Z(n21761) );
  IV U39389 ( .A(n21776), .Z(n37851) );
  XOR U39390 ( .A(n37858), .B(n37859), .Z(n21776) );
  XNOR U39391 ( .A(n21793), .B(n21774), .Z(n37859) );
  XNOR U39392 ( .A(q[0]), .B(DB[2235]), .Z(n21774) );
  XOR U39393 ( .A(n37860), .B(n21782), .Z(n21793) );
  XNOR U39394 ( .A(q[7]), .B(DB[2242]), .Z(n21782) );
  IV U39395 ( .A(n21781), .Z(n37860) );
  XNOR U39396 ( .A(n21779), .B(n37861), .Z(n21781) );
  XNOR U39397 ( .A(q[6]), .B(DB[2241]), .Z(n37861) );
  XNOR U39398 ( .A(q[5]), .B(DB[2240]), .Z(n21779) );
  IV U39399 ( .A(n21792), .Z(n37858) );
  XOR U39400 ( .A(n37862), .B(n37863), .Z(n21792) );
  XNOR U39401 ( .A(n21788), .B(n21790), .Z(n37863) );
  XNOR U39402 ( .A(q[1]), .B(DB[2236]), .Z(n21790) );
  XNOR U39403 ( .A(q[4]), .B(DB[2239]), .Z(n21788) );
  IV U39404 ( .A(n21787), .Z(n37862) );
  XNOR U39405 ( .A(n21785), .B(n37864), .Z(n21787) );
  XNOR U39406 ( .A(q[3]), .B(DB[2238]), .Z(n37864) );
  XNOR U39407 ( .A(q[2]), .B(DB[2237]), .Z(n21785) );
  XOR U39408 ( .A(n37865), .B(n21683), .Z(n21611) );
  XOR U39409 ( .A(n37866), .B(n21675), .Z(n21683) );
  XOR U39410 ( .A(n37867), .B(n21664), .Z(n21675) );
  XNOR U39411 ( .A(q[14]), .B(DB[2264]), .Z(n21664) );
  IV U39412 ( .A(n21663), .Z(n37867) );
  XNOR U39413 ( .A(n21661), .B(n37868), .Z(n21663) );
  XNOR U39414 ( .A(q[13]), .B(DB[2263]), .Z(n37868) );
  XNOR U39415 ( .A(q[12]), .B(DB[2262]), .Z(n21661) );
  IV U39416 ( .A(n21674), .Z(n37866) );
  XOR U39417 ( .A(n37869), .B(n37870), .Z(n21674) );
  XNOR U39418 ( .A(n21670), .B(n21672), .Z(n37870) );
  XNOR U39419 ( .A(q[8]), .B(DB[2258]), .Z(n21672) );
  XNOR U39420 ( .A(q[11]), .B(DB[2261]), .Z(n21670) );
  IV U39421 ( .A(n21669), .Z(n37869) );
  XNOR U39422 ( .A(n21667), .B(n37871), .Z(n21669) );
  XNOR U39423 ( .A(q[10]), .B(DB[2260]), .Z(n37871) );
  XNOR U39424 ( .A(q[9]), .B(DB[2259]), .Z(n21667) );
  IV U39425 ( .A(n21682), .Z(n37865) );
  XOR U39426 ( .A(n37872), .B(n37873), .Z(n21682) );
  XNOR U39427 ( .A(n21699), .B(n21680), .Z(n37873) );
  XNOR U39428 ( .A(q[0]), .B(DB[2250]), .Z(n21680) );
  XOR U39429 ( .A(n37874), .B(n21688), .Z(n21699) );
  XNOR U39430 ( .A(q[7]), .B(DB[2257]), .Z(n21688) );
  IV U39431 ( .A(n21687), .Z(n37874) );
  XNOR U39432 ( .A(n21685), .B(n37875), .Z(n21687) );
  XNOR U39433 ( .A(q[6]), .B(DB[2256]), .Z(n37875) );
  XNOR U39434 ( .A(q[5]), .B(DB[2255]), .Z(n21685) );
  IV U39435 ( .A(n21698), .Z(n37872) );
  XOR U39436 ( .A(n37876), .B(n37877), .Z(n21698) );
  XNOR U39437 ( .A(n21694), .B(n21696), .Z(n37877) );
  XNOR U39438 ( .A(q[1]), .B(DB[2251]), .Z(n21696) );
  XNOR U39439 ( .A(q[4]), .B(DB[2254]), .Z(n21694) );
  IV U39440 ( .A(n21693), .Z(n37876) );
  XNOR U39441 ( .A(n21691), .B(n37878), .Z(n21693) );
  XNOR U39442 ( .A(q[3]), .B(DB[2253]), .Z(n37878) );
  XNOR U39443 ( .A(q[2]), .B(DB[2252]), .Z(n21691) );
  XOR U39444 ( .A(n37879), .B(n21589), .Z(n21517) );
  XOR U39445 ( .A(n37880), .B(n21581), .Z(n21589) );
  XOR U39446 ( .A(n37881), .B(n21570), .Z(n21581) );
  XNOR U39447 ( .A(q[14]), .B(DB[2279]), .Z(n21570) );
  IV U39448 ( .A(n21569), .Z(n37881) );
  XNOR U39449 ( .A(n21567), .B(n37882), .Z(n21569) );
  XNOR U39450 ( .A(q[13]), .B(DB[2278]), .Z(n37882) );
  XNOR U39451 ( .A(q[12]), .B(DB[2277]), .Z(n21567) );
  IV U39452 ( .A(n21580), .Z(n37880) );
  XOR U39453 ( .A(n37883), .B(n37884), .Z(n21580) );
  XNOR U39454 ( .A(n21576), .B(n21578), .Z(n37884) );
  XNOR U39455 ( .A(q[8]), .B(DB[2273]), .Z(n21578) );
  XNOR U39456 ( .A(q[11]), .B(DB[2276]), .Z(n21576) );
  IV U39457 ( .A(n21575), .Z(n37883) );
  XNOR U39458 ( .A(n21573), .B(n37885), .Z(n21575) );
  XNOR U39459 ( .A(q[10]), .B(DB[2275]), .Z(n37885) );
  XNOR U39460 ( .A(q[9]), .B(DB[2274]), .Z(n21573) );
  IV U39461 ( .A(n21588), .Z(n37879) );
  XOR U39462 ( .A(n37886), .B(n37887), .Z(n21588) );
  XNOR U39463 ( .A(n21605), .B(n21586), .Z(n37887) );
  XNOR U39464 ( .A(q[0]), .B(DB[2265]), .Z(n21586) );
  XOR U39465 ( .A(n37888), .B(n21594), .Z(n21605) );
  XNOR U39466 ( .A(q[7]), .B(DB[2272]), .Z(n21594) );
  IV U39467 ( .A(n21593), .Z(n37888) );
  XNOR U39468 ( .A(n21591), .B(n37889), .Z(n21593) );
  XNOR U39469 ( .A(q[6]), .B(DB[2271]), .Z(n37889) );
  XNOR U39470 ( .A(q[5]), .B(DB[2270]), .Z(n21591) );
  IV U39471 ( .A(n21604), .Z(n37886) );
  XOR U39472 ( .A(n37890), .B(n37891), .Z(n21604) );
  XNOR U39473 ( .A(n21600), .B(n21602), .Z(n37891) );
  XNOR U39474 ( .A(q[1]), .B(DB[2266]), .Z(n21602) );
  XNOR U39475 ( .A(q[4]), .B(DB[2269]), .Z(n21600) );
  IV U39476 ( .A(n21599), .Z(n37890) );
  XNOR U39477 ( .A(n21597), .B(n37892), .Z(n21599) );
  XNOR U39478 ( .A(q[3]), .B(DB[2268]), .Z(n37892) );
  XNOR U39479 ( .A(q[2]), .B(DB[2267]), .Z(n21597) );
  XOR U39480 ( .A(n37893), .B(n21495), .Z(n21423) );
  XOR U39481 ( .A(n37894), .B(n21487), .Z(n21495) );
  XOR U39482 ( .A(n37895), .B(n21476), .Z(n21487) );
  XNOR U39483 ( .A(q[14]), .B(DB[2294]), .Z(n21476) );
  IV U39484 ( .A(n21475), .Z(n37895) );
  XNOR U39485 ( .A(n21473), .B(n37896), .Z(n21475) );
  XNOR U39486 ( .A(q[13]), .B(DB[2293]), .Z(n37896) );
  XNOR U39487 ( .A(q[12]), .B(DB[2292]), .Z(n21473) );
  IV U39488 ( .A(n21486), .Z(n37894) );
  XOR U39489 ( .A(n37897), .B(n37898), .Z(n21486) );
  XNOR U39490 ( .A(n21482), .B(n21484), .Z(n37898) );
  XNOR U39491 ( .A(q[8]), .B(DB[2288]), .Z(n21484) );
  XNOR U39492 ( .A(q[11]), .B(DB[2291]), .Z(n21482) );
  IV U39493 ( .A(n21481), .Z(n37897) );
  XNOR U39494 ( .A(n21479), .B(n37899), .Z(n21481) );
  XNOR U39495 ( .A(q[10]), .B(DB[2290]), .Z(n37899) );
  XNOR U39496 ( .A(q[9]), .B(DB[2289]), .Z(n21479) );
  IV U39497 ( .A(n21494), .Z(n37893) );
  XOR U39498 ( .A(n37900), .B(n37901), .Z(n21494) );
  XNOR U39499 ( .A(n21511), .B(n21492), .Z(n37901) );
  XNOR U39500 ( .A(q[0]), .B(DB[2280]), .Z(n21492) );
  XOR U39501 ( .A(n37902), .B(n21500), .Z(n21511) );
  XNOR U39502 ( .A(q[7]), .B(DB[2287]), .Z(n21500) );
  IV U39503 ( .A(n21499), .Z(n37902) );
  XNOR U39504 ( .A(n21497), .B(n37903), .Z(n21499) );
  XNOR U39505 ( .A(q[6]), .B(DB[2286]), .Z(n37903) );
  XNOR U39506 ( .A(q[5]), .B(DB[2285]), .Z(n21497) );
  IV U39507 ( .A(n21510), .Z(n37900) );
  XOR U39508 ( .A(n37904), .B(n37905), .Z(n21510) );
  XNOR U39509 ( .A(n21506), .B(n21508), .Z(n37905) );
  XNOR U39510 ( .A(q[1]), .B(DB[2281]), .Z(n21508) );
  XNOR U39511 ( .A(q[4]), .B(DB[2284]), .Z(n21506) );
  IV U39512 ( .A(n21505), .Z(n37904) );
  XNOR U39513 ( .A(n21503), .B(n37906), .Z(n21505) );
  XNOR U39514 ( .A(q[3]), .B(DB[2283]), .Z(n37906) );
  XNOR U39515 ( .A(q[2]), .B(DB[2282]), .Z(n21503) );
  XOR U39516 ( .A(n37907), .B(n21401), .Z(n21329) );
  XOR U39517 ( .A(n37908), .B(n21393), .Z(n21401) );
  XOR U39518 ( .A(n37909), .B(n21382), .Z(n21393) );
  XNOR U39519 ( .A(q[14]), .B(DB[2309]), .Z(n21382) );
  IV U39520 ( .A(n21381), .Z(n37909) );
  XNOR U39521 ( .A(n21379), .B(n37910), .Z(n21381) );
  XNOR U39522 ( .A(q[13]), .B(DB[2308]), .Z(n37910) );
  XNOR U39523 ( .A(q[12]), .B(DB[2307]), .Z(n21379) );
  IV U39524 ( .A(n21392), .Z(n37908) );
  XOR U39525 ( .A(n37911), .B(n37912), .Z(n21392) );
  XNOR U39526 ( .A(n21388), .B(n21390), .Z(n37912) );
  XNOR U39527 ( .A(q[8]), .B(DB[2303]), .Z(n21390) );
  XNOR U39528 ( .A(q[11]), .B(DB[2306]), .Z(n21388) );
  IV U39529 ( .A(n21387), .Z(n37911) );
  XNOR U39530 ( .A(n21385), .B(n37913), .Z(n21387) );
  XNOR U39531 ( .A(q[10]), .B(DB[2305]), .Z(n37913) );
  XNOR U39532 ( .A(q[9]), .B(DB[2304]), .Z(n21385) );
  IV U39533 ( .A(n21400), .Z(n37907) );
  XOR U39534 ( .A(n37914), .B(n37915), .Z(n21400) );
  XNOR U39535 ( .A(n21417), .B(n21398), .Z(n37915) );
  XNOR U39536 ( .A(q[0]), .B(DB[2295]), .Z(n21398) );
  XOR U39537 ( .A(n37916), .B(n21406), .Z(n21417) );
  XNOR U39538 ( .A(q[7]), .B(DB[2302]), .Z(n21406) );
  IV U39539 ( .A(n21405), .Z(n37916) );
  XNOR U39540 ( .A(n21403), .B(n37917), .Z(n21405) );
  XNOR U39541 ( .A(q[6]), .B(DB[2301]), .Z(n37917) );
  XNOR U39542 ( .A(q[5]), .B(DB[2300]), .Z(n21403) );
  IV U39543 ( .A(n21416), .Z(n37914) );
  XOR U39544 ( .A(n37918), .B(n37919), .Z(n21416) );
  XNOR U39545 ( .A(n21412), .B(n21414), .Z(n37919) );
  XNOR U39546 ( .A(q[1]), .B(DB[2296]), .Z(n21414) );
  XNOR U39547 ( .A(q[4]), .B(DB[2299]), .Z(n21412) );
  IV U39548 ( .A(n21411), .Z(n37918) );
  XNOR U39549 ( .A(n21409), .B(n37920), .Z(n21411) );
  XNOR U39550 ( .A(q[3]), .B(DB[2298]), .Z(n37920) );
  XNOR U39551 ( .A(q[2]), .B(DB[2297]), .Z(n21409) );
  XOR U39552 ( .A(n37921), .B(n21307), .Z(n21235) );
  XOR U39553 ( .A(n37922), .B(n21299), .Z(n21307) );
  XOR U39554 ( .A(n37923), .B(n21288), .Z(n21299) );
  XNOR U39555 ( .A(q[14]), .B(DB[2324]), .Z(n21288) );
  IV U39556 ( .A(n21287), .Z(n37923) );
  XNOR U39557 ( .A(n21285), .B(n37924), .Z(n21287) );
  XNOR U39558 ( .A(q[13]), .B(DB[2323]), .Z(n37924) );
  XNOR U39559 ( .A(q[12]), .B(DB[2322]), .Z(n21285) );
  IV U39560 ( .A(n21298), .Z(n37922) );
  XOR U39561 ( .A(n37925), .B(n37926), .Z(n21298) );
  XNOR U39562 ( .A(n21294), .B(n21296), .Z(n37926) );
  XNOR U39563 ( .A(q[8]), .B(DB[2318]), .Z(n21296) );
  XNOR U39564 ( .A(q[11]), .B(DB[2321]), .Z(n21294) );
  IV U39565 ( .A(n21293), .Z(n37925) );
  XNOR U39566 ( .A(n21291), .B(n37927), .Z(n21293) );
  XNOR U39567 ( .A(q[10]), .B(DB[2320]), .Z(n37927) );
  XNOR U39568 ( .A(q[9]), .B(DB[2319]), .Z(n21291) );
  IV U39569 ( .A(n21306), .Z(n37921) );
  XOR U39570 ( .A(n37928), .B(n37929), .Z(n21306) );
  XNOR U39571 ( .A(n21323), .B(n21304), .Z(n37929) );
  XNOR U39572 ( .A(q[0]), .B(DB[2310]), .Z(n21304) );
  XOR U39573 ( .A(n37930), .B(n21312), .Z(n21323) );
  XNOR U39574 ( .A(q[7]), .B(DB[2317]), .Z(n21312) );
  IV U39575 ( .A(n21311), .Z(n37930) );
  XNOR U39576 ( .A(n21309), .B(n37931), .Z(n21311) );
  XNOR U39577 ( .A(q[6]), .B(DB[2316]), .Z(n37931) );
  XNOR U39578 ( .A(q[5]), .B(DB[2315]), .Z(n21309) );
  IV U39579 ( .A(n21322), .Z(n37928) );
  XOR U39580 ( .A(n37932), .B(n37933), .Z(n21322) );
  XNOR U39581 ( .A(n21318), .B(n21320), .Z(n37933) );
  XNOR U39582 ( .A(q[1]), .B(DB[2311]), .Z(n21320) );
  XNOR U39583 ( .A(q[4]), .B(DB[2314]), .Z(n21318) );
  IV U39584 ( .A(n21317), .Z(n37932) );
  XNOR U39585 ( .A(n21315), .B(n37934), .Z(n21317) );
  XNOR U39586 ( .A(q[3]), .B(DB[2313]), .Z(n37934) );
  XNOR U39587 ( .A(q[2]), .B(DB[2312]), .Z(n21315) );
  XOR U39588 ( .A(n37935), .B(n21213), .Z(n21141) );
  XOR U39589 ( .A(n37936), .B(n21205), .Z(n21213) );
  XOR U39590 ( .A(n37937), .B(n21194), .Z(n21205) );
  XNOR U39591 ( .A(q[14]), .B(DB[2339]), .Z(n21194) );
  IV U39592 ( .A(n21193), .Z(n37937) );
  XNOR U39593 ( .A(n21191), .B(n37938), .Z(n21193) );
  XNOR U39594 ( .A(q[13]), .B(DB[2338]), .Z(n37938) );
  XNOR U39595 ( .A(q[12]), .B(DB[2337]), .Z(n21191) );
  IV U39596 ( .A(n21204), .Z(n37936) );
  XOR U39597 ( .A(n37939), .B(n37940), .Z(n21204) );
  XNOR U39598 ( .A(n21200), .B(n21202), .Z(n37940) );
  XNOR U39599 ( .A(q[8]), .B(DB[2333]), .Z(n21202) );
  XNOR U39600 ( .A(q[11]), .B(DB[2336]), .Z(n21200) );
  IV U39601 ( .A(n21199), .Z(n37939) );
  XNOR U39602 ( .A(n21197), .B(n37941), .Z(n21199) );
  XNOR U39603 ( .A(q[10]), .B(DB[2335]), .Z(n37941) );
  XNOR U39604 ( .A(q[9]), .B(DB[2334]), .Z(n21197) );
  IV U39605 ( .A(n21212), .Z(n37935) );
  XOR U39606 ( .A(n37942), .B(n37943), .Z(n21212) );
  XNOR U39607 ( .A(n21229), .B(n21210), .Z(n37943) );
  XNOR U39608 ( .A(q[0]), .B(DB[2325]), .Z(n21210) );
  XOR U39609 ( .A(n37944), .B(n21218), .Z(n21229) );
  XNOR U39610 ( .A(q[7]), .B(DB[2332]), .Z(n21218) );
  IV U39611 ( .A(n21217), .Z(n37944) );
  XNOR U39612 ( .A(n21215), .B(n37945), .Z(n21217) );
  XNOR U39613 ( .A(q[6]), .B(DB[2331]), .Z(n37945) );
  XNOR U39614 ( .A(q[5]), .B(DB[2330]), .Z(n21215) );
  IV U39615 ( .A(n21228), .Z(n37942) );
  XOR U39616 ( .A(n37946), .B(n37947), .Z(n21228) );
  XNOR U39617 ( .A(n21224), .B(n21226), .Z(n37947) );
  XNOR U39618 ( .A(q[1]), .B(DB[2326]), .Z(n21226) );
  XNOR U39619 ( .A(q[4]), .B(DB[2329]), .Z(n21224) );
  IV U39620 ( .A(n21223), .Z(n37946) );
  XNOR U39621 ( .A(n21221), .B(n37948), .Z(n21223) );
  XNOR U39622 ( .A(q[3]), .B(DB[2328]), .Z(n37948) );
  XNOR U39623 ( .A(q[2]), .B(DB[2327]), .Z(n21221) );
  XOR U39624 ( .A(n37949), .B(n21119), .Z(n21047) );
  XOR U39625 ( .A(n37950), .B(n21111), .Z(n21119) );
  XOR U39626 ( .A(n37951), .B(n21100), .Z(n21111) );
  XNOR U39627 ( .A(q[14]), .B(DB[2354]), .Z(n21100) );
  IV U39628 ( .A(n21099), .Z(n37951) );
  XNOR U39629 ( .A(n21097), .B(n37952), .Z(n21099) );
  XNOR U39630 ( .A(q[13]), .B(DB[2353]), .Z(n37952) );
  XNOR U39631 ( .A(q[12]), .B(DB[2352]), .Z(n21097) );
  IV U39632 ( .A(n21110), .Z(n37950) );
  XOR U39633 ( .A(n37953), .B(n37954), .Z(n21110) );
  XNOR U39634 ( .A(n21106), .B(n21108), .Z(n37954) );
  XNOR U39635 ( .A(q[8]), .B(DB[2348]), .Z(n21108) );
  XNOR U39636 ( .A(q[11]), .B(DB[2351]), .Z(n21106) );
  IV U39637 ( .A(n21105), .Z(n37953) );
  XNOR U39638 ( .A(n21103), .B(n37955), .Z(n21105) );
  XNOR U39639 ( .A(q[10]), .B(DB[2350]), .Z(n37955) );
  XNOR U39640 ( .A(q[9]), .B(DB[2349]), .Z(n21103) );
  IV U39641 ( .A(n21118), .Z(n37949) );
  XOR U39642 ( .A(n37956), .B(n37957), .Z(n21118) );
  XNOR U39643 ( .A(n21135), .B(n21116), .Z(n37957) );
  XNOR U39644 ( .A(q[0]), .B(DB[2340]), .Z(n21116) );
  XOR U39645 ( .A(n37958), .B(n21124), .Z(n21135) );
  XNOR U39646 ( .A(q[7]), .B(DB[2347]), .Z(n21124) );
  IV U39647 ( .A(n21123), .Z(n37958) );
  XNOR U39648 ( .A(n21121), .B(n37959), .Z(n21123) );
  XNOR U39649 ( .A(q[6]), .B(DB[2346]), .Z(n37959) );
  XNOR U39650 ( .A(q[5]), .B(DB[2345]), .Z(n21121) );
  IV U39651 ( .A(n21134), .Z(n37956) );
  XOR U39652 ( .A(n37960), .B(n37961), .Z(n21134) );
  XNOR U39653 ( .A(n21130), .B(n21132), .Z(n37961) );
  XNOR U39654 ( .A(q[1]), .B(DB[2341]), .Z(n21132) );
  XNOR U39655 ( .A(q[4]), .B(DB[2344]), .Z(n21130) );
  IV U39656 ( .A(n21129), .Z(n37960) );
  XNOR U39657 ( .A(n21127), .B(n37962), .Z(n21129) );
  XNOR U39658 ( .A(q[3]), .B(DB[2343]), .Z(n37962) );
  XNOR U39659 ( .A(q[2]), .B(DB[2342]), .Z(n21127) );
  XOR U39660 ( .A(n37963), .B(n21025), .Z(n20953) );
  XOR U39661 ( .A(n37964), .B(n21017), .Z(n21025) );
  XOR U39662 ( .A(n37965), .B(n21006), .Z(n21017) );
  XNOR U39663 ( .A(q[14]), .B(DB[2369]), .Z(n21006) );
  IV U39664 ( .A(n21005), .Z(n37965) );
  XNOR U39665 ( .A(n21003), .B(n37966), .Z(n21005) );
  XNOR U39666 ( .A(q[13]), .B(DB[2368]), .Z(n37966) );
  XNOR U39667 ( .A(q[12]), .B(DB[2367]), .Z(n21003) );
  IV U39668 ( .A(n21016), .Z(n37964) );
  XOR U39669 ( .A(n37967), .B(n37968), .Z(n21016) );
  XNOR U39670 ( .A(n21012), .B(n21014), .Z(n37968) );
  XNOR U39671 ( .A(q[8]), .B(DB[2363]), .Z(n21014) );
  XNOR U39672 ( .A(q[11]), .B(DB[2366]), .Z(n21012) );
  IV U39673 ( .A(n21011), .Z(n37967) );
  XNOR U39674 ( .A(n21009), .B(n37969), .Z(n21011) );
  XNOR U39675 ( .A(q[10]), .B(DB[2365]), .Z(n37969) );
  XNOR U39676 ( .A(q[9]), .B(DB[2364]), .Z(n21009) );
  IV U39677 ( .A(n21024), .Z(n37963) );
  XOR U39678 ( .A(n37970), .B(n37971), .Z(n21024) );
  XNOR U39679 ( .A(n21041), .B(n21022), .Z(n37971) );
  XNOR U39680 ( .A(q[0]), .B(DB[2355]), .Z(n21022) );
  XOR U39681 ( .A(n37972), .B(n21030), .Z(n21041) );
  XNOR U39682 ( .A(q[7]), .B(DB[2362]), .Z(n21030) );
  IV U39683 ( .A(n21029), .Z(n37972) );
  XNOR U39684 ( .A(n21027), .B(n37973), .Z(n21029) );
  XNOR U39685 ( .A(q[6]), .B(DB[2361]), .Z(n37973) );
  XNOR U39686 ( .A(q[5]), .B(DB[2360]), .Z(n21027) );
  IV U39687 ( .A(n21040), .Z(n37970) );
  XOR U39688 ( .A(n37974), .B(n37975), .Z(n21040) );
  XNOR U39689 ( .A(n21036), .B(n21038), .Z(n37975) );
  XNOR U39690 ( .A(q[1]), .B(DB[2356]), .Z(n21038) );
  XNOR U39691 ( .A(q[4]), .B(DB[2359]), .Z(n21036) );
  IV U39692 ( .A(n21035), .Z(n37974) );
  XNOR U39693 ( .A(n21033), .B(n37976), .Z(n21035) );
  XNOR U39694 ( .A(q[3]), .B(DB[2358]), .Z(n37976) );
  XNOR U39695 ( .A(q[2]), .B(DB[2357]), .Z(n21033) );
  XOR U39696 ( .A(n37977), .B(n20931), .Z(n20859) );
  XOR U39697 ( .A(n37978), .B(n20923), .Z(n20931) );
  XOR U39698 ( .A(n37979), .B(n20912), .Z(n20923) );
  XNOR U39699 ( .A(q[14]), .B(DB[2384]), .Z(n20912) );
  IV U39700 ( .A(n20911), .Z(n37979) );
  XNOR U39701 ( .A(n20909), .B(n37980), .Z(n20911) );
  XNOR U39702 ( .A(q[13]), .B(DB[2383]), .Z(n37980) );
  XNOR U39703 ( .A(q[12]), .B(DB[2382]), .Z(n20909) );
  IV U39704 ( .A(n20922), .Z(n37978) );
  XOR U39705 ( .A(n37981), .B(n37982), .Z(n20922) );
  XNOR U39706 ( .A(n20918), .B(n20920), .Z(n37982) );
  XNOR U39707 ( .A(q[8]), .B(DB[2378]), .Z(n20920) );
  XNOR U39708 ( .A(q[11]), .B(DB[2381]), .Z(n20918) );
  IV U39709 ( .A(n20917), .Z(n37981) );
  XNOR U39710 ( .A(n20915), .B(n37983), .Z(n20917) );
  XNOR U39711 ( .A(q[10]), .B(DB[2380]), .Z(n37983) );
  XNOR U39712 ( .A(q[9]), .B(DB[2379]), .Z(n20915) );
  IV U39713 ( .A(n20930), .Z(n37977) );
  XOR U39714 ( .A(n37984), .B(n37985), .Z(n20930) );
  XNOR U39715 ( .A(n20947), .B(n20928), .Z(n37985) );
  XNOR U39716 ( .A(q[0]), .B(DB[2370]), .Z(n20928) );
  XOR U39717 ( .A(n37986), .B(n20936), .Z(n20947) );
  XNOR U39718 ( .A(q[7]), .B(DB[2377]), .Z(n20936) );
  IV U39719 ( .A(n20935), .Z(n37986) );
  XNOR U39720 ( .A(n20933), .B(n37987), .Z(n20935) );
  XNOR U39721 ( .A(q[6]), .B(DB[2376]), .Z(n37987) );
  XNOR U39722 ( .A(q[5]), .B(DB[2375]), .Z(n20933) );
  IV U39723 ( .A(n20946), .Z(n37984) );
  XOR U39724 ( .A(n37988), .B(n37989), .Z(n20946) );
  XNOR U39725 ( .A(n20942), .B(n20944), .Z(n37989) );
  XNOR U39726 ( .A(q[1]), .B(DB[2371]), .Z(n20944) );
  XNOR U39727 ( .A(q[4]), .B(DB[2374]), .Z(n20942) );
  IV U39728 ( .A(n20941), .Z(n37988) );
  XNOR U39729 ( .A(n20939), .B(n37990), .Z(n20941) );
  XNOR U39730 ( .A(q[3]), .B(DB[2373]), .Z(n37990) );
  XNOR U39731 ( .A(q[2]), .B(DB[2372]), .Z(n20939) );
  XOR U39732 ( .A(n37991), .B(n20837), .Z(n20765) );
  XOR U39733 ( .A(n37992), .B(n20829), .Z(n20837) );
  XOR U39734 ( .A(n37993), .B(n20818), .Z(n20829) );
  XNOR U39735 ( .A(q[14]), .B(DB[2399]), .Z(n20818) );
  IV U39736 ( .A(n20817), .Z(n37993) );
  XNOR U39737 ( .A(n20815), .B(n37994), .Z(n20817) );
  XNOR U39738 ( .A(q[13]), .B(DB[2398]), .Z(n37994) );
  XNOR U39739 ( .A(q[12]), .B(DB[2397]), .Z(n20815) );
  IV U39740 ( .A(n20828), .Z(n37992) );
  XOR U39741 ( .A(n37995), .B(n37996), .Z(n20828) );
  XNOR U39742 ( .A(n20824), .B(n20826), .Z(n37996) );
  XNOR U39743 ( .A(q[8]), .B(DB[2393]), .Z(n20826) );
  XNOR U39744 ( .A(q[11]), .B(DB[2396]), .Z(n20824) );
  IV U39745 ( .A(n20823), .Z(n37995) );
  XNOR U39746 ( .A(n20821), .B(n37997), .Z(n20823) );
  XNOR U39747 ( .A(q[10]), .B(DB[2395]), .Z(n37997) );
  XNOR U39748 ( .A(q[9]), .B(DB[2394]), .Z(n20821) );
  IV U39749 ( .A(n20836), .Z(n37991) );
  XOR U39750 ( .A(n37998), .B(n37999), .Z(n20836) );
  XNOR U39751 ( .A(n20853), .B(n20834), .Z(n37999) );
  XNOR U39752 ( .A(q[0]), .B(DB[2385]), .Z(n20834) );
  XOR U39753 ( .A(n38000), .B(n20842), .Z(n20853) );
  XNOR U39754 ( .A(q[7]), .B(DB[2392]), .Z(n20842) );
  IV U39755 ( .A(n20841), .Z(n38000) );
  XNOR U39756 ( .A(n20839), .B(n38001), .Z(n20841) );
  XNOR U39757 ( .A(q[6]), .B(DB[2391]), .Z(n38001) );
  XNOR U39758 ( .A(q[5]), .B(DB[2390]), .Z(n20839) );
  IV U39759 ( .A(n20852), .Z(n37998) );
  XOR U39760 ( .A(n38002), .B(n38003), .Z(n20852) );
  XNOR U39761 ( .A(n20848), .B(n20850), .Z(n38003) );
  XNOR U39762 ( .A(q[1]), .B(DB[2386]), .Z(n20850) );
  XNOR U39763 ( .A(q[4]), .B(DB[2389]), .Z(n20848) );
  IV U39764 ( .A(n20847), .Z(n38002) );
  XNOR U39765 ( .A(n20845), .B(n38004), .Z(n20847) );
  XNOR U39766 ( .A(q[3]), .B(DB[2388]), .Z(n38004) );
  XNOR U39767 ( .A(q[2]), .B(DB[2387]), .Z(n20845) );
  XOR U39768 ( .A(n38005), .B(n20743), .Z(n20671) );
  XOR U39769 ( .A(n38006), .B(n20735), .Z(n20743) );
  XOR U39770 ( .A(n38007), .B(n20724), .Z(n20735) );
  XNOR U39771 ( .A(q[14]), .B(DB[2414]), .Z(n20724) );
  IV U39772 ( .A(n20723), .Z(n38007) );
  XNOR U39773 ( .A(n20721), .B(n38008), .Z(n20723) );
  XNOR U39774 ( .A(q[13]), .B(DB[2413]), .Z(n38008) );
  XNOR U39775 ( .A(q[12]), .B(DB[2412]), .Z(n20721) );
  IV U39776 ( .A(n20734), .Z(n38006) );
  XOR U39777 ( .A(n38009), .B(n38010), .Z(n20734) );
  XNOR U39778 ( .A(n20730), .B(n20732), .Z(n38010) );
  XNOR U39779 ( .A(q[8]), .B(DB[2408]), .Z(n20732) );
  XNOR U39780 ( .A(q[11]), .B(DB[2411]), .Z(n20730) );
  IV U39781 ( .A(n20729), .Z(n38009) );
  XNOR U39782 ( .A(n20727), .B(n38011), .Z(n20729) );
  XNOR U39783 ( .A(q[10]), .B(DB[2410]), .Z(n38011) );
  XNOR U39784 ( .A(q[9]), .B(DB[2409]), .Z(n20727) );
  IV U39785 ( .A(n20742), .Z(n38005) );
  XOR U39786 ( .A(n38012), .B(n38013), .Z(n20742) );
  XNOR U39787 ( .A(n20759), .B(n20740), .Z(n38013) );
  XNOR U39788 ( .A(q[0]), .B(DB[2400]), .Z(n20740) );
  XOR U39789 ( .A(n38014), .B(n20748), .Z(n20759) );
  XNOR U39790 ( .A(q[7]), .B(DB[2407]), .Z(n20748) );
  IV U39791 ( .A(n20747), .Z(n38014) );
  XNOR U39792 ( .A(n20745), .B(n38015), .Z(n20747) );
  XNOR U39793 ( .A(q[6]), .B(DB[2406]), .Z(n38015) );
  XNOR U39794 ( .A(q[5]), .B(DB[2405]), .Z(n20745) );
  IV U39795 ( .A(n20758), .Z(n38012) );
  XOR U39796 ( .A(n38016), .B(n38017), .Z(n20758) );
  XNOR U39797 ( .A(n20754), .B(n20756), .Z(n38017) );
  XNOR U39798 ( .A(q[1]), .B(DB[2401]), .Z(n20756) );
  XNOR U39799 ( .A(q[4]), .B(DB[2404]), .Z(n20754) );
  IV U39800 ( .A(n20753), .Z(n38016) );
  XNOR U39801 ( .A(n20751), .B(n38018), .Z(n20753) );
  XNOR U39802 ( .A(q[3]), .B(DB[2403]), .Z(n38018) );
  XNOR U39803 ( .A(q[2]), .B(DB[2402]), .Z(n20751) );
  XOR U39804 ( .A(n38019), .B(n20649), .Z(n20577) );
  XOR U39805 ( .A(n38020), .B(n20641), .Z(n20649) );
  XOR U39806 ( .A(n38021), .B(n20630), .Z(n20641) );
  XNOR U39807 ( .A(q[14]), .B(DB[2429]), .Z(n20630) );
  IV U39808 ( .A(n20629), .Z(n38021) );
  XNOR U39809 ( .A(n20627), .B(n38022), .Z(n20629) );
  XNOR U39810 ( .A(q[13]), .B(DB[2428]), .Z(n38022) );
  XNOR U39811 ( .A(q[12]), .B(DB[2427]), .Z(n20627) );
  IV U39812 ( .A(n20640), .Z(n38020) );
  XOR U39813 ( .A(n38023), .B(n38024), .Z(n20640) );
  XNOR U39814 ( .A(n20636), .B(n20638), .Z(n38024) );
  XNOR U39815 ( .A(q[8]), .B(DB[2423]), .Z(n20638) );
  XNOR U39816 ( .A(q[11]), .B(DB[2426]), .Z(n20636) );
  IV U39817 ( .A(n20635), .Z(n38023) );
  XNOR U39818 ( .A(n20633), .B(n38025), .Z(n20635) );
  XNOR U39819 ( .A(q[10]), .B(DB[2425]), .Z(n38025) );
  XNOR U39820 ( .A(q[9]), .B(DB[2424]), .Z(n20633) );
  IV U39821 ( .A(n20648), .Z(n38019) );
  XOR U39822 ( .A(n38026), .B(n38027), .Z(n20648) );
  XNOR U39823 ( .A(n20665), .B(n20646), .Z(n38027) );
  XNOR U39824 ( .A(q[0]), .B(DB[2415]), .Z(n20646) );
  XOR U39825 ( .A(n38028), .B(n20654), .Z(n20665) );
  XNOR U39826 ( .A(q[7]), .B(DB[2422]), .Z(n20654) );
  IV U39827 ( .A(n20653), .Z(n38028) );
  XNOR U39828 ( .A(n20651), .B(n38029), .Z(n20653) );
  XNOR U39829 ( .A(q[6]), .B(DB[2421]), .Z(n38029) );
  XNOR U39830 ( .A(q[5]), .B(DB[2420]), .Z(n20651) );
  IV U39831 ( .A(n20664), .Z(n38026) );
  XOR U39832 ( .A(n38030), .B(n38031), .Z(n20664) );
  XNOR U39833 ( .A(n20660), .B(n20662), .Z(n38031) );
  XNOR U39834 ( .A(q[1]), .B(DB[2416]), .Z(n20662) );
  XNOR U39835 ( .A(q[4]), .B(DB[2419]), .Z(n20660) );
  IV U39836 ( .A(n20659), .Z(n38030) );
  XNOR U39837 ( .A(n20657), .B(n38032), .Z(n20659) );
  XNOR U39838 ( .A(q[3]), .B(DB[2418]), .Z(n38032) );
  XNOR U39839 ( .A(q[2]), .B(DB[2417]), .Z(n20657) );
  XOR U39840 ( .A(n38033), .B(n20555), .Z(n20483) );
  XOR U39841 ( .A(n38034), .B(n20547), .Z(n20555) );
  XOR U39842 ( .A(n38035), .B(n20536), .Z(n20547) );
  XNOR U39843 ( .A(q[14]), .B(DB[2444]), .Z(n20536) );
  IV U39844 ( .A(n20535), .Z(n38035) );
  XNOR U39845 ( .A(n20533), .B(n38036), .Z(n20535) );
  XNOR U39846 ( .A(q[13]), .B(DB[2443]), .Z(n38036) );
  XNOR U39847 ( .A(q[12]), .B(DB[2442]), .Z(n20533) );
  IV U39848 ( .A(n20546), .Z(n38034) );
  XOR U39849 ( .A(n38037), .B(n38038), .Z(n20546) );
  XNOR U39850 ( .A(n20542), .B(n20544), .Z(n38038) );
  XNOR U39851 ( .A(q[8]), .B(DB[2438]), .Z(n20544) );
  XNOR U39852 ( .A(q[11]), .B(DB[2441]), .Z(n20542) );
  IV U39853 ( .A(n20541), .Z(n38037) );
  XNOR U39854 ( .A(n20539), .B(n38039), .Z(n20541) );
  XNOR U39855 ( .A(q[10]), .B(DB[2440]), .Z(n38039) );
  XNOR U39856 ( .A(q[9]), .B(DB[2439]), .Z(n20539) );
  IV U39857 ( .A(n20554), .Z(n38033) );
  XOR U39858 ( .A(n38040), .B(n38041), .Z(n20554) );
  XNOR U39859 ( .A(n20571), .B(n20552), .Z(n38041) );
  XNOR U39860 ( .A(q[0]), .B(DB[2430]), .Z(n20552) );
  XOR U39861 ( .A(n38042), .B(n20560), .Z(n20571) );
  XNOR U39862 ( .A(q[7]), .B(DB[2437]), .Z(n20560) );
  IV U39863 ( .A(n20559), .Z(n38042) );
  XNOR U39864 ( .A(n20557), .B(n38043), .Z(n20559) );
  XNOR U39865 ( .A(q[6]), .B(DB[2436]), .Z(n38043) );
  XNOR U39866 ( .A(q[5]), .B(DB[2435]), .Z(n20557) );
  IV U39867 ( .A(n20570), .Z(n38040) );
  XOR U39868 ( .A(n38044), .B(n38045), .Z(n20570) );
  XNOR U39869 ( .A(n20566), .B(n20568), .Z(n38045) );
  XNOR U39870 ( .A(q[1]), .B(DB[2431]), .Z(n20568) );
  XNOR U39871 ( .A(q[4]), .B(DB[2434]), .Z(n20566) );
  IV U39872 ( .A(n20565), .Z(n38044) );
  XNOR U39873 ( .A(n20563), .B(n38046), .Z(n20565) );
  XNOR U39874 ( .A(q[3]), .B(DB[2433]), .Z(n38046) );
  XNOR U39875 ( .A(q[2]), .B(DB[2432]), .Z(n20563) );
  XOR U39876 ( .A(n38047), .B(n20461), .Z(n20389) );
  XOR U39877 ( .A(n38048), .B(n20453), .Z(n20461) );
  XOR U39878 ( .A(n38049), .B(n20442), .Z(n20453) );
  XNOR U39879 ( .A(q[14]), .B(DB[2459]), .Z(n20442) );
  IV U39880 ( .A(n20441), .Z(n38049) );
  XNOR U39881 ( .A(n20439), .B(n38050), .Z(n20441) );
  XNOR U39882 ( .A(q[13]), .B(DB[2458]), .Z(n38050) );
  XNOR U39883 ( .A(q[12]), .B(DB[2457]), .Z(n20439) );
  IV U39884 ( .A(n20452), .Z(n38048) );
  XOR U39885 ( .A(n38051), .B(n38052), .Z(n20452) );
  XNOR U39886 ( .A(n20448), .B(n20450), .Z(n38052) );
  XNOR U39887 ( .A(q[8]), .B(DB[2453]), .Z(n20450) );
  XNOR U39888 ( .A(q[11]), .B(DB[2456]), .Z(n20448) );
  IV U39889 ( .A(n20447), .Z(n38051) );
  XNOR U39890 ( .A(n20445), .B(n38053), .Z(n20447) );
  XNOR U39891 ( .A(q[10]), .B(DB[2455]), .Z(n38053) );
  XNOR U39892 ( .A(q[9]), .B(DB[2454]), .Z(n20445) );
  IV U39893 ( .A(n20460), .Z(n38047) );
  XOR U39894 ( .A(n38054), .B(n38055), .Z(n20460) );
  XNOR U39895 ( .A(n20477), .B(n20458), .Z(n38055) );
  XNOR U39896 ( .A(q[0]), .B(DB[2445]), .Z(n20458) );
  XOR U39897 ( .A(n38056), .B(n20466), .Z(n20477) );
  XNOR U39898 ( .A(q[7]), .B(DB[2452]), .Z(n20466) );
  IV U39899 ( .A(n20465), .Z(n38056) );
  XNOR U39900 ( .A(n20463), .B(n38057), .Z(n20465) );
  XNOR U39901 ( .A(q[6]), .B(DB[2451]), .Z(n38057) );
  XNOR U39902 ( .A(q[5]), .B(DB[2450]), .Z(n20463) );
  IV U39903 ( .A(n20476), .Z(n38054) );
  XOR U39904 ( .A(n38058), .B(n38059), .Z(n20476) );
  XNOR U39905 ( .A(n20472), .B(n20474), .Z(n38059) );
  XNOR U39906 ( .A(q[1]), .B(DB[2446]), .Z(n20474) );
  XNOR U39907 ( .A(q[4]), .B(DB[2449]), .Z(n20472) );
  IV U39908 ( .A(n20471), .Z(n38058) );
  XNOR U39909 ( .A(n20469), .B(n38060), .Z(n20471) );
  XNOR U39910 ( .A(q[3]), .B(DB[2448]), .Z(n38060) );
  XNOR U39911 ( .A(q[2]), .B(DB[2447]), .Z(n20469) );
  XOR U39912 ( .A(n38061), .B(n20367), .Z(n20295) );
  XOR U39913 ( .A(n38062), .B(n20359), .Z(n20367) );
  XOR U39914 ( .A(n38063), .B(n20348), .Z(n20359) );
  XNOR U39915 ( .A(q[14]), .B(DB[2474]), .Z(n20348) );
  IV U39916 ( .A(n20347), .Z(n38063) );
  XNOR U39917 ( .A(n20345), .B(n38064), .Z(n20347) );
  XNOR U39918 ( .A(q[13]), .B(DB[2473]), .Z(n38064) );
  XNOR U39919 ( .A(q[12]), .B(DB[2472]), .Z(n20345) );
  IV U39920 ( .A(n20358), .Z(n38062) );
  XOR U39921 ( .A(n38065), .B(n38066), .Z(n20358) );
  XNOR U39922 ( .A(n20354), .B(n20356), .Z(n38066) );
  XNOR U39923 ( .A(q[8]), .B(DB[2468]), .Z(n20356) );
  XNOR U39924 ( .A(q[11]), .B(DB[2471]), .Z(n20354) );
  IV U39925 ( .A(n20353), .Z(n38065) );
  XNOR U39926 ( .A(n20351), .B(n38067), .Z(n20353) );
  XNOR U39927 ( .A(q[10]), .B(DB[2470]), .Z(n38067) );
  XNOR U39928 ( .A(q[9]), .B(DB[2469]), .Z(n20351) );
  IV U39929 ( .A(n20366), .Z(n38061) );
  XOR U39930 ( .A(n38068), .B(n38069), .Z(n20366) );
  XNOR U39931 ( .A(n20383), .B(n20364), .Z(n38069) );
  XNOR U39932 ( .A(q[0]), .B(DB[2460]), .Z(n20364) );
  XOR U39933 ( .A(n38070), .B(n20372), .Z(n20383) );
  XNOR U39934 ( .A(q[7]), .B(DB[2467]), .Z(n20372) );
  IV U39935 ( .A(n20371), .Z(n38070) );
  XNOR U39936 ( .A(n20369), .B(n38071), .Z(n20371) );
  XNOR U39937 ( .A(q[6]), .B(DB[2466]), .Z(n38071) );
  XNOR U39938 ( .A(q[5]), .B(DB[2465]), .Z(n20369) );
  IV U39939 ( .A(n20382), .Z(n38068) );
  XOR U39940 ( .A(n38072), .B(n38073), .Z(n20382) );
  XNOR U39941 ( .A(n20378), .B(n20380), .Z(n38073) );
  XNOR U39942 ( .A(q[1]), .B(DB[2461]), .Z(n20380) );
  XNOR U39943 ( .A(q[4]), .B(DB[2464]), .Z(n20378) );
  IV U39944 ( .A(n20377), .Z(n38072) );
  XNOR U39945 ( .A(n20375), .B(n38074), .Z(n20377) );
  XNOR U39946 ( .A(q[3]), .B(DB[2463]), .Z(n38074) );
  XNOR U39947 ( .A(q[2]), .B(DB[2462]), .Z(n20375) );
  XOR U39948 ( .A(n38075), .B(n20273), .Z(n20201) );
  XOR U39949 ( .A(n38076), .B(n20265), .Z(n20273) );
  XOR U39950 ( .A(n38077), .B(n20254), .Z(n20265) );
  XNOR U39951 ( .A(q[14]), .B(DB[2489]), .Z(n20254) );
  IV U39952 ( .A(n20253), .Z(n38077) );
  XNOR U39953 ( .A(n20251), .B(n38078), .Z(n20253) );
  XNOR U39954 ( .A(q[13]), .B(DB[2488]), .Z(n38078) );
  XNOR U39955 ( .A(q[12]), .B(DB[2487]), .Z(n20251) );
  IV U39956 ( .A(n20264), .Z(n38076) );
  XOR U39957 ( .A(n38079), .B(n38080), .Z(n20264) );
  XNOR U39958 ( .A(n20260), .B(n20262), .Z(n38080) );
  XNOR U39959 ( .A(q[8]), .B(DB[2483]), .Z(n20262) );
  XNOR U39960 ( .A(q[11]), .B(DB[2486]), .Z(n20260) );
  IV U39961 ( .A(n20259), .Z(n38079) );
  XNOR U39962 ( .A(n20257), .B(n38081), .Z(n20259) );
  XNOR U39963 ( .A(q[10]), .B(DB[2485]), .Z(n38081) );
  XNOR U39964 ( .A(q[9]), .B(DB[2484]), .Z(n20257) );
  IV U39965 ( .A(n20272), .Z(n38075) );
  XOR U39966 ( .A(n38082), .B(n38083), .Z(n20272) );
  XNOR U39967 ( .A(n20289), .B(n20270), .Z(n38083) );
  XNOR U39968 ( .A(q[0]), .B(DB[2475]), .Z(n20270) );
  XOR U39969 ( .A(n38084), .B(n20278), .Z(n20289) );
  XNOR U39970 ( .A(q[7]), .B(DB[2482]), .Z(n20278) );
  IV U39971 ( .A(n20277), .Z(n38084) );
  XNOR U39972 ( .A(n20275), .B(n38085), .Z(n20277) );
  XNOR U39973 ( .A(q[6]), .B(DB[2481]), .Z(n38085) );
  XNOR U39974 ( .A(q[5]), .B(DB[2480]), .Z(n20275) );
  IV U39975 ( .A(n20288), .Z(n38082) );
  XOR U39976 ( .A(n38086), .B(n38087), .Z(n20288) );
  XNOR U39977 ( .A(n20284), .B(n20286), .Z(n38087) );
  XNOR U39978 ( .A(q[1]), .B(DB[2476]), .Z(n20286) );
  XNOR U39979 ( .A(q[4]), .B(DB[2479]), .Z(n20284) );
  IV U39980 ( .A(n20283), .Z(n38086) );
  XNOR U39981 ( .A(n20281), .B(n38088), .Z(n20283) );
  XNOR U39982 ( .A(q[3]), .B(DB[2478]), .Z(n38088) );
  XNOR U39983 ( .A(q[2]), .B(DB[2477]), .Z(n20281) );
  XOR U39984 ( .A(n38089), .B(n20179), .Z(n20107) );
  XOR U39985 ( .A(n38090), .B(n20171), .Z(n20179) );
  XOR U39986 ( .A(n38091), .B(n20160), .Z(n20171) );
  XNOR U39987 ( .A(q[14]), .B(DB[2504]), .Z(n20160) );
  IV U39988 ( .A(n20159), .Z(n38091) );
  XNOR U39989 ( .A(n20157), .B(n38092), .Z(n20159) );
  XNOR U39990 ( .A(q[13]), .B(DB[2503]), .Z(n38092) );
  XNOR U39991 ( .A(q[12]), .B(DB[2502]), .Z(n20157) );
  IV U39992 ( .A(n20170), .Z(n38090) );
  XOR U39993 ( .A(n38093), .B(n38094), .Z(n20170) );
  XNOR U39994 ( .A(n20166), .B(n20168), .Z(n38094) );
  XNOR U39995 ( .A(q[8]), .B(DB[2498]), .Z(n20168) );
  XNOR U39996 ( .A(q[11]), .B(DB[2501]), .Z(n20166) );
  IV U39997 ( .A(n20165), .Z(n38093) );
  XNOR U39998 ( .A(n20163), .B(n38095), .Z(n20165) );
  XNOR U39999 ( .A(q[10]), .B(DB[2500]), .Z(n38095) );
  XNOR U40000 ( .A(q[9]), .B(DB[2499]), .Z(n20163) );
  IV U40001 ( .A(n20178), .Z(n38089) );
  XOR U40002 ( .A(n38096), .B(n38097), .Z(n20178) );
  XNOR U40003 ( .A(n20195), .B(n20176), .Z(n38097) );
  XNOR U40004 ( .A(q[0]), .B(DB[2490]), .Z(n20176) );
  XOR U40005 ( .A(n38098), .B(n20184), .Z(n20195) );
  XNOR U40006 ( .A(q[7]), .B(DB[2497]), .Z(n20184) );
  IV U40007 ( .A(n20183), .Z(n38098) );
  XNOR U40008 ( .A(n20181), .B(n38099), .Z(n20183) );
  XNOR U40009 ( .A(q[6]), .B(DB[2496]), .Z(n38099) );
  XNOR U40010 ( .A(q[5]), .B(DB[2495]), .Z(n20181) );
  IV U40011 ( .A(n20194), .Z(n38096) );
  XOR U40012 ( .A(n38100), .B(n38101), .Z(n20194) );
  XNOR U40013 ( .A(n20190), .B(n20192), .Z(n38101) );
  XNOR U40014 ( .A(q[1]), .B(DB[2491]), .Z(n20192) );
  XNOR U40015 ( .A(q[4]), .B(DB[2494]), .Z(n20190) );
  IV U40016 ( .A(n20189), .Z(n38100) );
  XNOR U40017 ( .A(n20187), .B(n38102), .Z(n20189) );
  XNOR U40018 ( .A(q[3]), .B(DB[2493]), .Z(n38102) );
  XNOR U40019 ( .A(q[2]), .B(DB[2492]), .Z(n20187) );
  XOR U40020 ( .A(n38103), .B(n20085), .Z(n20013) );
  XOR U40021 ( .A(n38104), .B(n20077), .Z(n20085) );
  XOR U40022 ( .A(n38105), .B(n20066), .Z(n20077) );
  XNOR U40023 ( .A(q[14]), .B(DB[2519]), .Z(n20066) );
  IV U40024 ( .A(n20065), .Z(n38105) );
  XNOR U40025 ( .A(n20063), .B(n38106), .Z(n20065) );
  XNOR U40026 ( .A(q[13]), .B(DB[2518]), .Z(n38106) );
  XNOR U40027 ( .A(q[12]), .B(DB[2517]), .Z(n20063) );
  IV U40028 ( .A(n20076), .Z(n38104) );
  XOR U40029 ( .A(n38107), .B(n38108), .Z(n20076) );
  XNOR U40030 ( .A(n20072), .B(n20074), .Z(n38108) );
  XNOR U40031 ( .A(q[8]), .B(DB[2513]), .Z(n20074) );
  XNOR U40032 ( .A(q[11]), .B(DB[2516]), .Z(n20072) );
  IV U40033 ( .A(n20071), .Z(n38107) );
  XNOR U40034 ( .A(n20069), .B(n38109), .Z(n20071) );
  XNOR U40035 ( .A(q[10]), .B(DB[2515]), .Z(n38109) );
  XNOR U40036 ( .A(q[9]), .B(DB[2514]), .Z(n20069) );
  IV U40037 ( .A(n20084), .Z(n38103) );
  XOR U40038 ( .A(n38110), .B(n38111), .Z(n20084) );
  XNOR U40039 ( .A(n20101), .B(n20082), .Z(n38111) );
  XNOR U40040 ( .A(q[0]), .B(DB[2505]), .Z(n20082) );
  XOR U40041 ( .A(n38112), .B(n20090), .Z(n20101) );
  XNOR U40042 ( .A(q[7]), .B(DB[2512]), .Z(n20090) );
  IV U40043 ( .A(n20089), .Z(n38112) );
  XNOR U40044 ( .A(n20087), .B(n38113), .Z(n20089) );
  XNOR U40045 ( .A(q[6]), .B(DB[2511]), .Z(n38113) );
  XNOR U40046 ( .A(q[5]), .B(DB[2510]), .Z(n20087) );
  IV U40047 ( .A(n20100), .Z(n38110) );
  XOR U40048 ( .A(n38114), .B(n38115), .Z(n20100) );
  XNOR U40049 ( .A(n20096), .B(n20098), .Z(n38115) );
  XNOR U40050 ( .A(q[1]), .B(DB[2506]), .Z(n20098) );
  XNOR U40051 ( .A(q[4]), .B(DB[2509]), .Z(n20096) );
  IV U40052 ( .A(n20095), .Z(n38114) );
  XNOR U40053 ( .A(n20093), .B(n38116), .Z(n20095) );
  XNOR U40054 ( .A(q[3]), .B(DB[2508]), .Z(n38116) );
  XNOR U40055 ( .A(q[2]), .B(DB[2507]), .Z(n20093) );
  XOR U40056 ( .A(n38117), .B(n19991), .Z(n19919) );
  XOR U40057 ( .A(n38118), .B(n19983), .Z(n19991) );
  XOR U40058 ( .A(n38119), .B(n19972), .Z(n19983) );
  XNOR U40059 ( .A(q[14]), .B(DB[2534]), .Z(n19972) );
  IV U40060 ( .A(n19971), .Z(n38119) );
  XNOR U40061 ( .A(n19969), .B(n38120), .Z(n19971) );
  XNOR U40062 ( .A(q[13]), .B(DB[2533]), .Z(n38120) );
  XNOR U40063 ( .A(q[12]), .B(DB[2532]), .Z(n19969) );
  IV U40064 ( .A(n19982), .Z(n38118) );
  XOR U40065 ( .A(n38121), .B(n38122), .Z(n19982) );
  XNOR U40066 ( .A(n19978), .B(n19980), .Z(n38122) );
  XNOR U40067 ( .A(q[8]), .B(DB[2528]), .Z(n19980) );
  XNOR U40068 ( .A(q[11]), .B(DB[2531]), .Z(n19978) );
  IV U40069 ( .A(n19977), .Z(n38121) );
  XNOR U40070 ( .A(n19975), .B(n38123), .Z(n19977) );
  XNOR U40071 ( .A(q[10]), .B(DB[2530]), .Z(n38123) );
  XNOR U40072 ( .A(q[9]), .B(DB[2529]), .Z(n19975) );
  IV U40073 ( .A(n19990), .Z(n38117) );
  XOR U40074 ( .A(n38124), .B(n38125), .Z(n19990) );
  XNOR U40075 ( .A(n20007), .B(n19988), .Z(n38125) );
  XNOR U40076 ( .A(q[0]), .B(DB[2520]), .Z(n19988) );
  XOR U40077 ( .A(n38126), .B(n19996), .Z(n20007) );
  XNOR U40078 ( .A(q[7]), .B(DB[2527]), .Z(n19996) );
  IV U40079 ( .A(n19995), .Z(n38126) );
  XNOR U40080 ( .A(n19993), .B(n38127), .Z(n19995) );
  XNOR U40081 ( .A(q[6]), .B(DB[2526]), .Z(n38127) );
  XNOR U40082 ( .A(q[5]), .B(DB[2525]), .Z(n19993) );
  IV U40083 ( .A(n20006), .Z(n38124) );
  XOR U40084 ( .A(n38128), .B(n38129), .Z(n20006) );
  XNOR U40085 ( .A(n20002), .B(n20004), .Z(n38129) );
  XNOR U40086 ( .A(q[1]), .B(DB[2521]), .Z(n20004) );
  XNOR U40087 ( .A(q[4]), .B(DB[2524]), .Z(n20002) );
  IV U40088 ( .A(n20001), .Z(n38128) );
  XNOR U40089 ( .A(n19999), .B(n38130), .Z(n20001) );
  XNOR U40090 ( .A(q[3]), .B(DB[2523]), .Z(n38130) );
  XNOR U40091 ( .A(q[2]), .B(DB[2522]), .Z(n19999) );
  XOR U40092 ( .A(n38131), .B(n19897), .Z(n19825) );
  XOR U40093 ( .A(n38132), .B(n19889), .Z(n19897) );
  XOR U40094 ( .A(n38133), .B(n19878), .Z(n19889) );
  XNOR U40095 ( .A(q[14]), .B(DB[2549]), .Z(n19878) );
  IV U40096 ( .A(n19877), .Z(n38133) );
  XNOR U40097 ( .A(n19875), .B(n38134), .Z(n19877) );
  XNOR U40098 ( .A(q[13]), .B(DB[2548]), .Z(n38134) );
  XNOR U40099 ( .A(q[12]), .B(DB[2547]), .Z(n19875) );
  IV U40100 ( .A(n19888), .Z(n38132) );
  XOR U40101 ( .A(n38135), .B(n38136), .Z(n19888) );
  XNOR U40102 ( .A(n19884), .B(n19886), .Z(n38136) );
  XNOR U40103 ( .A(q[8]), .B(DB[2543]), .Z(n19886) );
  XNOR U40104 ( .A(q[11]), .B(DB[2546]), .Z(n19884) );
  IV U40105 ( .A(n19883), .Z(n38135) );
  XNOR U40106 ( .A(n19881), .B(n38137), .Z(n19883) );
  XNOR U40107 ( .A(q[10]), .B(DB[2545]), .Z(n38137) );
  XNOR U40108 ( .A(q[9]), .B(DB[2544]), .Z(n19881) );
  IV U40109 ( .A(n19896), .Z(n38131) );
  XOR U40110 ( .A(n38138), .B(n38139), .Z(n19896) );
  XNOR U40111 ( .A(n19913), .B(n19894), .Z(n38139) );
  XNOR U40112 ( .A(q[0]), .B(DB[2535]), .Z(n19894) );
  XOR U40113 ( .A(n38140), .B(n19902), .Z(n19913) );
  XNOR U40114 ( .A(q[7]), .B(DB[2542]), .Z(n19902) );
  IV U40115 ( .A(n19901), .Z(n38140) );
  XNOR U40116 ( .A(n19899), .B(n38141), .Z(n19901) );
  XNOR U40117 ( .A(q[6]), .B(DB[2541]), .Z(n38141) );
  XNOR U40118 ( .A(q[5]), .B(DB[2540]), .Z(n19899) );
  IV U40119 ( .A(n19912), .Z(n38138) );
  XOR U40120 ( .A(n38142), .B(n38143), .Z(n19912) );
  XNOR U40121 ( .A(n19908), .B(n19910), .Z(n38143) );
  XNOR U40122 ( .A(q[1]), .B(DB[2536]), .Z(n19910) );
  XNOR U40123 ( .A(q[4]), .B(DB[2539]), .Z(n19908) );
  IV U40124 ( .A(n19907), .Z(n38142) );
  XNOR U40125 ( .A(n19905), .B(n38144), .Z(n19907) );
  XNOR U40126 ( .A(q[3]), .B(DB[2538]), .Z(n38144) );
  XNOR U40127 ( .A(q[2]), .B(DB[2537]), .Z(n19905) );
  XOR U40128 ( .A(n38145), .B(n19803), .Z(n19731) );
  XOR U40129 ( .A(n38146), .B(n19795), .Z(n19803) );
  XOR U40130 ( .A(n38147), .B(n19784), .Z(n19795) );
  XNOR U40131 ( .A(q[14]), .B(DB[2564]), .Z(n19784) );
  IV U40132 ( .A(n19783), .Z(n38147) );
  XNOR U40133 ( .A(n19781), .B(n38148), .Z(n19783) );
  XNOR U40134 ( .A(q[13]), .B(DB[2563]), .Z(n38148) );
  XNOR U40135 ( .A(q[12]), .B(DB[2562]), .Z(n19781) );
  IV U40136 ( .A(n19794), .Z(n38146) );
  XOR U40137 ( .A(n38149), .B(n38150), .Z(n19794) );
  XNOR U40138 ( .A(n19790), .B(n19792), .Z(n38150) );
  XNOR U40139 ( .A(q[8]), .B(DB[2558]), .Z(n19792) );
  XNOR U40140 ( .A(q[11]), .B(DB[2561]), .Z(n19790) );
  IV U40141 ( .A(n19789), .Z(n38149) );
  XNOR U40142 ( .A(n19787), .B(n38151), .Z(n19789) );
  XNOR U40143 ( .A(q[10]), .B(DB[2560]), .Z(n38151) );
  XNOR U40144 ( .A(q[9]), .B(DB[2559]), .Z(n19787) );
  IV U40145 ( .A(n19802), .Z(n38145) );
  XOR U40146 ( .A(n38152), .B(n38153), .Z(n19802) );
  XNOR U40147 ( .A(n19819), .B(n19800), .Z(n38153) );
  XNOR U40148 ( .A(q[0]), .B(DB[2550]), .Z(n19800) );
  XOR U40149 ( .A(n38154), .B(n19808), .Z(n19819) );
  XNOR U40150 ( .A(q[7]), .B(DB[2557]), .Z(n19808) );
  IV U40151 ( .A(n19807), .Z(n38154) );
  XNOR U40152 ( .A(n19805), .B(n38155), .Z(n19807) );
  XNOR U40153 ( .A(q[6]), .B(DB[2556]), .Z(n38155) );
  XNOR U40154 ( .A(q[5]), .B(DB[2555]), .Z(n19805) );
  IV U40155 ( .A(n19818), .Z(n38152) );
  XOR U40156 ( .A(n38156), .B(n38157), .Z(n19818) );
  XNOR U40157 ( .A(n19814), .B(n19816), .Z(n38157) );
  XNOR U40158 ( .A(q[1]), .B(DB[2551]), .Z(n19816) );
  XNOR U40159 ( .A(q[4]), .B(DB[2554]), .Z(n19814) );
  IV U40160 ( .A(n19813), .Z(n38156) );
  XNOR U40161 ( .A(n19811), .B(n38158), .Z(n19813) );
  XNOR U40162 ( .A(q[3]), .B(DB[2553]), .Z(n38158) );
  XNOR U40163 ( .A(q[2]), .B(DB[2552]), .Z(n19811) );
  XOR U40164 ( .A(n38159), .B(n19709), .Z(n19637) );
  XOR U40165 ( .A(n38160), .B(n19701), .Z(n19709) );
  XOR U40166 ( .A(n38161), .B(n19690), .Z(n19701) );
  XNOR U40167 ( .A(q[14]), .B(DB[2579]), .Z(n19690) );
  IV U40168 ( .A(n19689), .Z(n38161) );
  XNOR U40169 ( .A(n19687), .B(n38162), .Z(n19689) );
  XNOR U40170 ( .A(q[13]), .B(DB[2578]), .Z(n38162) );
  XNOR U40171 ( .A(q[12]), .B(DB[2577]), .Z(n19687) );
  IV U40172 ( .A(n19700), .Z(n38160) );
  XOR U40173 ( .A(n38163), .B(n38164), .Z(n19700) );
  XNOR U40174 ( .A(n19696), .B(n19698), .Z(n38164) );
  XNOR U40175 ( .A(q[8]), .B(DB[2573]), .Z(n19698) );
  XNOR U40176 ( .A(q[11]), .B(DB[2576]), .Z(n19696) );
  IV U40177 ( .A(n19695), .Z(n38163) );
  XNOR U40178 ( .A(n19693), .B(n38165), .Z(n19695) );
  XNOR U40179 ( .A(q[10]), .B(DB[2575]), .Z(n38165) );
  XNOR U40180 ( .A(q[9]), .B(DB[2574]), .Z(n19693) );
  IV U40181 ( .A(n19708), .Z(n38159) );
  XOR U40182 ( .A(n38166), .B(n38167), .Z(n19708) );
  XNOR U40183 ( .A(n19725), .B(n19706), .Z(n38167) );
  XNOR U40184 ( .A(q[0]), .B(DB[2565]), .Z(n19706) );
  XOR U40185 ( .A(n38168), .B(n19714), .Z(n19725) );
  XNOR U40186 ( .A(q[7]), .B(DB[2572]), .Z(n19714) );
  IV U40187 ( .A(n19713), .Z(n38168) );
  XNOR U40188 ( .A(n19711), .B(n38169), .Z(n19713) );
  XNOR U40189 ( .A(q[6]), .B(DB[2571]), .Z(n38169) );
  XNOR U40190 ( .A(q[5]), .B(DB[2570]), .Z(n19711) );
  IV U40191 ( .A(n19724), .Z(n38166) );
  XOR U40192 ( .A(n38170), .B(n38171), .Z(n19724) );
  XNOR U40193 ( .A(n19720), .B(n19722), .Z(n38171) );
  XNOR U40194 ( .A(q[1]), .B(DB[2566]), .Z(n19722) );
  XNOR U40195 ( .A(q[4]), .B(DB[2569]), .Z(n19720) );
  IV U40196 ( .A(n19719), .Z(n38170) );
  XNOR U40197 ( .A(n19717), .B(n38172), .Z(n19719) );
  XNOR U40198 ( .A(q[3]), .B(DB[2568]), .Z(n38172) );
  XNOR U40199 ( .A(q[2]), .B(DB[2567]), .Z(n19717) );
  XOR U40200 ( .A(n38173), .B(n19615), .Z(n19543) );
  XOR U40201 ( .A(n38174), .B(n19607), .Z(n19615) );
  XOR U40202 ( .A(n38175), .B(n19596), .Z(n19607) );
  XNOR U40203 ( .A(q[14]), .B(DB[2594]), .Z(n19596) );
  IV U40204 ( .A(n19595), .Z(n38175) );
  XNOR U40205 ( .A(n19593), .B(n38176), .Z(n19595) );
  XNOR U40206 ( .A(q[13]), .B(DB[2593]), .Z(n38176) );
  XNOR U40207 ( .A(q[12]), .B(DB[2592]), .Z(n19593) );
  IV U40208 ( .A(n19606), .Z(n38174) );
  XOR U40209 ( .A(n38177), .B(n38178), .Z(n19606) );
  XNOR U40210 ( .A(n19602), .B(n19604), .Z(n38178) );
  XNOR U40211 ( .A(q[8]), .B(DB[2588]), .Z(n19604) );
  XNOR U40212 ( .A(q[11]), .B(DB[2591]), .Z(n19602) );
  IV U40213 ( .A(n19601), .Z(n38177) );
  XNOR U40214 ( .A(n19599), .B(n38179), .Z(n19601) );
  XNOR U40215 ( .A(q[10]), .B(DB[2590]), .Z(n38179) );
  XNOR U40216 ( .A(q[9]), .B(DB[2589]), .Z(n19599) );
  IV U40217 ( .A(n19614), .Z(n38173) );
  XOR U40218 ( .A(n38180), .B(n38181), .Z(n19614) );
  XNOR U40219 ( .A(n19631), .B(n19612), .Z(n38181) );
  XNOR U40220 ( .A(q[0]), .B(DB[2580]), .Z(n19612) );
  XOR U40221 ( .A(n38182), .B(n19620), .Z(n19631) );
  XNOR U40222 ( .A(q[7]), .B(DB[2587]), .Z(n19620) );
  IV U40223 ( .A(n19619), .Z(n38182) );
  XNOR U40224 ( .A(n19617), .B(n38183), .Z(n19619) );
  XNOR U40225 ( .A(q[6]), .B(DB[2586]), .Z(n38183) );
  XNOR U40226 ( .A(q[5]), .B(DB[2585]), .Z(n19617) );
  IV U40227 ( .A(n19630), .Z(n38180) );
  XOR U40228 ( .A(n38184), .B(n38185), .Z(n19630) );
  XNOR U40229 ( .A(n19626), .B(n19628), .Z(n38185) );
  XNOR U40230 ( .A(q[1]), .B(DB[2581]), .Z(n19628) );
  XNOR U40231 ( .A(q[4]), .B(DB[2584]), .Z(n19626) );
  IV U40232 ( .A(n19625), .Z(n38184) );
  XNOR U40233 ( .A(n19623), .B(n38186), .Z(n19625) );
  XNOR U40234 ( .A(q[3]), .B(DB[2583]), .Z(n38186) );
  XNOR U40235 ( .A(q[2]), .B(DB[2582]), .Z(n19623) );
  XOR U40236 ( .A(n38187), .B(n19521), .Z(n19449) );
  XOR U40237 ( .A(n38188), .B(n19513), .Z(n19521) );
  XOR U40238 ( .A(n38189), .B(n19502), .Z(n19513) );
  XNOR U40239 ( .A(q[14]), .B(DB[2609]), .Z(n19502) );
  IV U40240 ( .A(n19501), .Z(n38189) );
  XNOR U40241 ( .A(n19499), .B(n38190), .Z(n19501) );
  XNOR U40242 ( .A(q[13]), .B(DB[2608]), .Z(n38190) );
  XNOR U40243 ( .A(q[12]), .B(DB[2607]), .Z(n19499) );
  IV U40244 ( .A(n19512), .Z(n38188) );
  XOR U40245 ( .A(n38191), .B(n38192), .Z(n19512) );
  XNOR U40246 ( .A(n19508), .B(n19510), .Z(n38192) );
  XNOR U40247 ( .A(q[8]), .B(DB[2603]), .Z(n19510) );
  XNOR U40248 ( .A(q[11]), .B(DB[2606]), .Z(n19508) );
  IV U40249 ( .A(n19507), .Z(n38191) );
  XNOR U40250 ( .A(n19505), .B(n38193), .Z(n19507) );
  XNOR U40251 ( .A(q[10]), .B(DB[2605]), .Z(n38193) );
  XNOR U40252 ( .A(q[9]), .B(DB[2604]), .Z(n19505) );
  IV U40253 ( .A(n19520), .Z(n38187) );
  XOR U40254 ( .A(n38194), .B(n38195), .Z(n19520) );
  XNOR U40255 ( .A(n19537), .B(n19518), .Z(n38195) );
  XNOR U40256 ( .A(q[0]), .B(DB[2595]), .Z(n19518) );
  XOR U40257 ( .A(n38196), .B(n19526), .Z(n19537) );
  XNOR U40258 ( .A(q[7]), .B(DB[2602]), .Z(n19526) );
  IV U40259 ( .A(n19525), .Z(n38196) );
  XNOR U40260 ( .A(n19523), .B(n38197), .Z(n19525) );
  XNOR U40261 ( .A(q[6]), .B(DB[2601]), .Z(n38197) );
  XNOR U40262 ( .A(q[5]), .B(DB[2600]), .Z(n19523) );
  IV U40263 ( .A(n19536), .Z(n38194) );
  XOR U40264 ( .A(n38198), .B(n38199), .Z(n19536) );
  XNOR U40265 ( .A(n19532), .B(n19534), .Z(n38199) );
  XNOR U40266 ( .A(q[1]), .B(DB[2596]), .Z(n19534) );
  XNOR U40267 ( .A(q[4]), .B(DB[2599]), .Z(n19532) );
  IV U40268 ( .A(n19531), .Z(n38198) );
  XNOR U40269 ( .A(n19529), .B(n38200), .Z(n19531) );
  XNOR U40270 ( .A(q[3]), .B(DB[2598]), .Z(n38200) );
  XNOR U40271 ( .A(q[2]), .B(DB[2597]), .Z(n19529) );
  XOR U40272 ( .A(n38201), .B(n19427), .Z(n19355) );
  XOR U40273 ( .A(n38202), .B(n19419), .Z(n19427) );
  XOR U40274 ( .A(n38203), .B(n19408), .Z(n19419) );
  XNOR U40275 ( .A(q[14]), .B(DB[2624]), .Z(n19408) );
  IV U40276 ( .A(n19407), .Z(n38203) );
  XNOR U40277 ( .A(n19405), .B(n38204), .Z(n19407) );
  XNOR U40278 ( .A(q[13]), .B(DB[2623]), .Z(n38204) );
  XNOR U40279 ( .A(q[12]), .B(DB[2622]), .Z(n19405) );
  IV U40280 ( .A(n19418), .Z(n38202) );
  XOR U40281 ( .A(n38205), .B(n38206), .Z(n19418) );
  XNOR U40282 ( .A(n19414), .B(n19416), .Z(n38206) );
  XNOR U40283 ( .A(q[8]), .B(DB[2618]), .Z(n19416) );
  XNOR U40284 ( .A(q[11]), .B(DB[2621]), .Z(n19414) );
  IV U40285 ( .A(n19413), .Z(n38205) );
  XNOR U40286 ( .A(n19411), .B(n38207), .Z(n19413) );
  XNOR U40287 ( .A(q[10]), .B(DB[2620]), .Z(n38207) );
  XNOR U40288 ( .A(q[9]), .B(DB[2619]), .Z(n19411) );
  IV U40289 ( .A(n19426), .Z(n38201) );
  XOR U40290 ( .A(n38208), .B(n38209), .Z(n19426) );
  XNOR U40291 ( .A(n19443), .B(n19424), .Z(n38209) );
  XNOR U40292 ( .A(q[0]), .B(DB[2610]), .Z(n19424) );
  XOR U40293 ( .A(n38210), .B(n19432), .Z(n19443) );
  XNOR U40294 ( .A(q[7]), .B(DB[2617]), .Z(n19432) );
  IV U40295 ( .A(n19431), .Z(n38210) );
  XNOR U40296 ( .A(n19429), .B(n38211), .Z(n19431) );
  XNOR U40297 ( .A(q[6]), .B(DB[2616]), .Z(n38211) );
  XNOR U40298 ( .A(q[5]), .B(DB[2615]), .Z(n19429) );
  IV U40299 ( .A(n19442), .Z(n38208) );
  XOR U40300 ( .A(n38212), .B(n38213), .Z(n19442) );
  XNOR U40301 ( .A(n19438), .B(n19440), .Z(n38213) );
  XNOR U40302 ( .A(q[1]), .B(DB[2611]), .Z(n19440) );
  XNOR U40303 ( .A(q[4]), .B(DB[2614]), .Z(n19438) );
  IV U40304 ( .A(n19437), .Z(n38212) );
  XNOR U40305 ( .A(n19435), .B(n38214), .Z(n19437) );
  XNOR U40306 ( .A(q[3]), .B(DB[2613]), .Z(n38214) );
  XNOR U40307 ( .A(q[2]), .B(DB[2612]), .Z(n19435) );
  XOR U40308 ( .A(n38215), .B(n19333), .Z(n19261) );
  XOR U40309 ( .A(n38216), .B(n19325), .Z(n19333) );
  XOR U40310 ( .A(n38217), .B(n19314), .Z(n19325) );
  XNOR U40311 ( .A(q[14]), .B(DB[2639]), .Z(n19314) );
  IV U40312 ( .A(n19313), .Z(n38217) );
  XNOR U40313 ( .A(n19311), .B(n38218), .Z(n19313) );
  XNOR U40314 ( .A(q[13]), .B(DB[2638]), .Z(n38218) );
  XNOR U40315 ( .A(q[12]), .B(DB[2637]), .Z(n19311) );
  IV U40316 ( .A(n19324), .Z(n38216) );
  XOR U40317 ( .A(n38219), .B(n38220), .Z(n19324) );
  XNOR U40318 ( .A(n19320), .B(n19322), .Z(n38220) );
  XNOR U40319 ( .A(q[8]), .B(DB[2633]), .Z(n19322) );
  XNOR U40320 ( .A(q[11]), .B(DB[2636]), .Z(n19320) );
  IV U40321 ( .A(n19319), .Z(n38219) );
  XNOR U40322 ( .A(n19317), .B(n38221), .Z(n19319) );
  XNOR U40323 ( .A(q[10]), .B(DB[2635]), .Z(n38221) );
  XNOR U40324 ( .A(q[9]), .B(DB[2634]), .Z(n19317) );
  IV U40325 ( .A(n19332), .Z(n38215) );
  XOR U40326 ( .A(n38222), .B(n38223), .Z(n19332) );
  XNOR U40327 ( .A(n19349), .B(n19330), .Z(n38223) );
  XNOR U40328 ( .A(q[0]), .B(DB[2625]), .Z(n19330) );
  XOR U40329 ( .A(n38224), .B(n19338), .Z(n19349) );
  XNOR U40330 ( .A(q[7]), .B(DB[2632]), .Z(n19338) );
  IV U40331 ( .A(n19337), .Z(n38224) );
  XNOR U40332 ( .A(n19335), .B(n38225), .Z(n19337) );
  XNOR U40333 ( .A(q[6]), .B(DB[2631]), .Z(n38225) );
  XNOR U40334 ( .A(q[5]), .B(DB[2630]), .Z(n19335) );
  IV U40335 ( .A(n19348), .Z(n38222) );
  XOR U40336 ( .A(n38226), .B(n38227), .Z(n19348) );
  XNOR U40337 ( .A(n19344), .B(n19346), .Z(n38227) );
  XNOR U40338 ( .A(q[1]), .B(DB[2626]), .Z(n19346) );
  XNOR U40339 ( .A(q[4]), .B(DB[2629]), .Z(n19344) );
  IV U40340 ( .A(n19343), .Z(n38226) );
  XNOR U40341 ( .A(n19341), .B(n38228), .Z(n19343) );
  XNOR U40342 ( .A(q[3]), .B(DB[2628]), .Z(n38228) );
  XNOR U40343 ( .A(q[2]), .B(DB[2627]), .Z(n19341) );
  XOR U40344 ( .A(n38229), .B(n19239), .Z(n19167) );
  XOR U40345 ( .A(n38230), .B(n19231), .Z(n19239) );
  XOR U40346 ( .A(n38231), .B(n19220), .Z(n19231) );
  XNOR U40347 ( .A(q[14]), .B(DB[2654]), .Z(n19220) );
  IV U40348 ( .A(n19219), .Z(n38231) );
  XNOR U40349 ( .A(n19217), .B(n38232), .Z(n19219) );
  XNOR U40350 ( .A(q[13]), .B(DB[2653]), .Z(n38232) );
  XNOR U40351 ( .A(q[12]), .B(DB[2652]), .Z(n19217) );
  IV U40352 ( .A(n19230), .Z(n38230) );
  XOR U40353 ( .A(n38233), .B(n38234), .Z(n19230) );
  XNOR U40354 ( .A(n19226), .B(n19228), .Z(n38234) );
  XNOR U40355 ( .A(q[8]), .B(DB[2648]), .Z(n19228) );
  XNOR U40356 ( .A(q[11]), .B(DB[2651]), .Z(n19226) );
  IV U40357 ( .A(n19225), .Z(n38233) );
  XNOR U40358 ( .A(n19223), .B(n38235), .Z(n19225) );
  XNOR U40359 ( .A(q[10]), .B(DB[2650]), .Z(n38235) );
  XNOR U40360 ( .A(q[9]), .B(DB[2649]), .Z(n19223) );
  IV U40361 ( .A(n19238), .Z(n38229) );
  XOR U40362 ( .A(n38236), .B(n38237), .Z(n19238) );
  XNOR U40363 ( .A(n19255), .B(n19236), .Z(n38237) );
  XNOR U40364 ( .A(q[0]), .B(DB[2640]), .Z(n19236) );
  XOR U40365 ( .A(n38238), .B(n19244), .Z(n19255) );
  XNOR U40366 ( .A(q[7]), .B(DB[2647]), .Z(n19244) );
  IV U40367 ( .A(n19243), .Z(n38238) );
  XNOR U40368 ( .A(n19241), .B(n38239), .Z(n19243) );
  XNOR U40369 ( .A(q[6]), .B(DB[2646]), .Z(n38239) );
  XNOR U40370 ( .A(q[5]), .B(DB[2645]), .Z(n19241) );
  IV U40371 ( .A(n19254), .Z(n38236) );
  XOR U40372 ( .A(n38240), .B(n38241), .Z(n19254) );
  XNOR U40373 ( .A(n19250), .B(n19252), .Z(n38241) );
  XNOR U40374 ( .A(q[1]), .B(DB[2641]), .Z(n19252) );
  XNOR U40375 ( .A(q[4]), .B(DB[2644]), .Z(n19250) );
  IV U40376 ( .A(n19249), .Z(n38240) );
  XNOR U40377 ( .A(n19247), .B(n38242), .Z(n19249) );
  XNOR U40378 ( .A(q[3]), .B(DB[2643]), .Z(n38242) );
  XNOR U40379 ( .A(q[2]), .B(DB[2642]), .Z(n19247) );
  XOR U40380 ( .A(n38243), .B(n19145), .Z(n19073) );
  XOR U40381 ( .A(n38244), .B(n19137), .Z(n19145) );
  XOR U40382 ( .A(n38245), .B(n19126), .Z(n19137) );
  XNOR U40383 ( .A(q[14]), .B(DB[2669]), .Z(n19126) );
  IV U40384 ( .A(n19125), .Z(n38245) );
  XNOR U40385 ( .A(n19123), .B(n38246), .Z(n19125) );
  XNOR U40386 ( .A(q[13]), .B(DB[2668]), .Z(n38246) );
  XNOR U40387 ( .A(q[12]), .B(DB[2667]), .Z(n19123) );
  IV U40388 ( .A(n19136), .Z(n38244) );
  XOR U40389 ( .A(n38247), .B(n38248), .Z(n19136) );
  XNOR U40390 ( .A(n19132), .B(n19134), .Z(n38248) );
  XNOR U40391 ( .A(q[8]), .B(DB[2663]), .Z(n19134) );
  XNOR U40392 ( .A(q[11]), .B(DB[2666]), .Z(n19132) );
  IV U40393 ( .A(n19131), .Z(n38247) );
  XNOR U40394 ( .A(n19129), .B(n38249), .Z(n19131) );
  XNOR U40395 ( .A(q[10]), .B(DB[2665]), .Z(n38249) );
  XNOR U40396 ( .A(q[9]), .B(DB[2664]), .Z(n19129) );
  IV U40397 ( .A(n19144), .Z(n38243) );
  XOR U40398 ( .A(n38250), .B(n38251), .Z(n19144) );
  XNOR U40399 ( .A(n19161), .B(n19142), .Z(n38251) );
  XNOR U40400 ( .A(q[0]), .B(DB[2655]), .Z(n19142) );
  XOR U40401 ( .A(n38252), .B(n19150), .Z(n19161) );
  XNOR U40402 ( .A(q[7]), .B(DB[2662]), .Z(n19150) );
  IV U40403 ( .A(n19149), .Z(n38252) );
  XNOR U40404 ( .A(n19147), .B(n38253), .Z(n19149) );
  XNOR U40405 ( .A(q[6]), .B(DB[2661]), .Z(n38253) );
  XNOR U40406 ( .A(q[5]), .B(DB[2660]), .Z(n19147) );
  IV U40407 ( .A(n19160), .Z(n38250) );
  XOR U40408 ( .A(n38254), .B(n38255), .Z(n19160) );
  XNOR U40409 ( .A(n19156), .B(n19158), .Z(n38255) );
  XNOR U40410 ( .A(q[1]), .B(DB[2656]), .Z(n19158) );
  XNOR U40411 ( .A(q[4]), .B(DB[2659]), .Z(n19156) );
  IV U40412 ( .A(n19155), .Z(n38254) );
  XNOR U40413 ( .A(n19153), .B(n38256), .Z(n19155) );
  XNOR U40414 ( .A(q[3]), .B(DB[2658]), .Z(n38256) );
  XNOR U40415 ( .A(q[2]), .B(DB[2657]), .Z(n19153) );
  XOR U40416 ( .A(n38257), .B(n19051), .Z(n18979) );
  XOR U40417 ( .A(n38258), .B(n19043), .Z(n19051) );
  XOR U40418 ( .A(n38259), .B(n19032), .Z(n19043) );
  XNOR U40419 ( .A(q[14]), .B(DB[2684]), .Z(n19032) );
  IV U40420 ( .A(n19031), .Z(n38259) );
  XNOR U40421 ( .A(n19029), .B(n38260), .Z(n19031) );
  XNOR U40422 ( .A(q[13]), .B(DB[2683]), .Z(n38260) );
  XNOR U40423 ( .A(q[12]), .B(DB[2682]), .Z(n19029) );
  IV U40424 ( .A(n19042), .Z(n38258) );
  XOR U40425 ( .A(n38261), .B(n38262), .Z(n19042) );
  XNOR U40426 ( .A(n19038), .B(n19040), .Z(n38262) );
  XNOR U40427 ( .A(q[8]), .B(DB[2678]), .Z(n19040) );
  XNOR U40428 ( .A(q[11]), .B(DB[2681]), .Z(n19038) );
  IV U40429 ( .A(n19037), .Z(n38261) );
  XNOR U40430 ( .A(n19035), .B(n38263), .Z(n19037) );
  XNOR U40431 ( .A(q[10]), .B(DB[2680]), .Z(n38263) );
  XNOR U40432 ( .A(q[9]), .B(DB[2679]), .Z(n19035) );
  IV U40433 ( .A(n19050), .Z(n38257) );
  XOR U40434 ( .A(n38264), .B(n38265), .Z(n19050) );
  XNOR U40435 ( .A(n19067), .B(n19048), .Z(n38265) );
  XNOR U40436 ( .A(q[0]), .B(DB[2670]), .Z(n19048) );
  XOR U40437 ( .A(n38266), .B(n19056), .Z(n19067) );
  XNOR U40438 ( .A(q[7]), .B(DB[2677]), .Z(n19056) );
  IV U40439 ( .A(n19055), .Z(n38266) );
  XNOR U40440 ( .A(n19053), .B(n38267), .Z(n19055) );
  XNOR U40441 ( .A(q[6]), .B(DB[2676]), .Z(n38267) );
  XNOR U40442 ( .A(q[5]), .B(DB[2675]), .Z(n19053) );
  IV U40443 ( .A(n19066), .Z(n38264) );
  XOR U40444 ( .A(n38268), .B(n38269), .Z(n19066) );
  XNOR U40445 ( .A(n19062), .B(n19064), .Z(n38269) );
  XNOR U40446 ( .A(q[1]), .B(DB[2671]), .Z(n19064) );
  XNOR U40447 ( .A(q[4]), .B(DB[2674]), .Z(n19062) );
  IV U40448 ( .A(n19061), .Z(n38268) );
  XNOR U40449 ( .A(n19059), .B(n38270), .Z(n19061) );
  XNOR U40450 ( .A(q[3]), .B(DB[2673]), .Z(n38270) );
  XNOR U40451 ( .A(q[2]), .B(DB[2672]), .Z(n19059) );
  XOR U40452 ( .A(n38271), .B(n18957), .Z(n18885) );
  XOR U40453 ( .A(n38272), .B(n18949), .Z(n18957) );
  XOR U40454 ( .A(n38273), .B(n18938), .Z(n18949) );
  XNOR U40455 ( .A(q[14]), .B(DB[2699]), .Z(n18938) );
  IV U40456 ( .A(n18937), .Z(n38273) );
  XNOR U40457 ( .A(n18935), .B(n38274), .Z(n18937) );
  XNOR U40458 ( .A(q[13]), .B(DB[2698]), .Z(n38274) );
  XNOR U40459 ( .A(q[12]), .B(DB[2697]), .Z(n18935) );
  IV U40460 ( .A(n18948), .Z(n38272) );
  XOR U40461 ( .A(n38275), .B(n38276), .Z(n18948) );
  XNOR U40462 ( .A(n18944), .B(n18946), .Z(n38276) );
  XNOR U40463 ( .A(q[8]), .B(DB[2693]), .Z(n18946) );
  XNOR U40464 ( .A(q[11]), .B(DB[2696]), .Z(n18944) );
  IV U40465 ( .A(n18943), .Z(n38275) );
  XNOR U40466 ( .A(n18941), .B(n38277), .Z(n18943) );
  XNOR U40467 ( .A(q[10]), .B(DB[2695]), .Z(n38277) );
  XNOR U40468 ( .A(q[9]), .B(DB[2694]), .Z(n18941) );
  IV U40469 ( .A(n18956), .Z(n38271) );
  XOR U40470 ( .A(n38278), .B(n38279), .Z(n18956) );
  XNOR U40471 ( .A(n18973), .B(n18954), .Z(n38279) );
  XNOR U40472 ( .A(q[0]), .B(DB[2685]), .Z(n18954) );
  XOR U40473 ( .A(n38280), .B(n18962), .Z(n18973) );
  XNOR U40474 ( .A(q[7]), .B(DB[2692]), .Z(n18962) );
  IV U40475 ( .A(n18961), .Z(n38280) );
  XNOR U40476 ( .A(n18959), .B(n38281), .Z(n18961) );
  XNOR U40477 ( .A(q[6]), .B(DB[2691]), .Z(n38281) );
  XNOR U40478 ( .A(q[5]), .B(DB[2690]), .Z(n18959) );
  IV U40479 ( .A(n18972), .Z(n38278) );
  XOR U40480 ( .A(n38282), .B(n38283), .Z(n18972) );
  XNOR U40481 ( .A(n18968), .B(n18970), .Z(n38283) );
  XNOR U40482 ( .A(q[1]), .B(DB[2686]), .Z(n18970) );
  XNOR U40483 ( .A(q[4]), .B(DB[2689]), .Z(n18968) );
  IV U40484 ( .A(n18967), .Z(n38282) );
  XNOR U40485 ( .A(n18965), .B(n38284), .Z(n18967) );
  XNOR U40486 ( .A(q[3]), .B(DB[2688]), .Z(n38284) );
  XNOR U40487 ( .A(q[2]), .B(DB[2687]), .Z(n18965) );
  XOR U40488 ( .A(n38285), .B(n18863), .Z(n18791) );
  XOR U40489 ( .A(n38286), .B(n18855), .Z(n18863) );
  XOR U40490 ( .A(n38287), .B(n18844), .Z(n18855) );
  XNOR U40491 ( .A(q[14]), .B(DB[2714]), .Z(n18844) );
  IV U40492 ( .A(n18843), .Z(n38287) );
  XNOR U40493 ( .A(n18841), .B(n38288), .Z(n18843) );
  XNOR U40494 ( .A(q[13]), .B(DB[2713]), .Z(n38288) );
  XNOR U40495 ( .A(q[12]), .B(DB[2712]), .Z(n18841) );
  IV U40496 ( .A(n18854), .Z(n38286) );
  XOR U40497 ( .A(n38289), .B(n38290), .Z(n18854) );
  XNOR U40498 ( .A(n18850), .B(n18852), .Z(n38290) );
  XNOR U40499 ( .A(q[8]), .B(DB[2708]), .Z(n18852) );
  XNOR U40500 ( .A(q[11]), .B(DB[2711]), .Z(n18850) );
  IV U40501 ( .A(n18849), .Z(n38289) );
  XNOR U40502 ( .A(n18847), .B(n38291), .Z(n18849) );
  XNOR U40503 ( .A(q[10]), .B(DB[2710]), .Z(n38291) );
  XNOR U40504 ( .A(q[9]), .B(DB[2709]), .Z(n18847) );
  IV U40505 ( .A(n18862), .Z(n38285) );
  XOR U40506 ( .A(n38292), .B(n38293), .Z(n18862) );
  XNOR U40507 ( .A(n18879), .B(n18860), .Z(n38293) );
  XNOR U40508 ( .A(q[0]), .B(DB[2700]), .Z(n18860) );
  XOR U40509 ( .A(n38294), .B(n18868), .Z(n18879) );
  XNOR U40510 ( .A(q[7]), .B(DB[2707]), .Z(n18868) );
  IV U40511 ( .A(n18867), .Z(n38294) );
  XNOR U40512 ( .A(n18865), .B(n38295), .Z(n18867) );
  XNOR U40513 ( .A(q[6]), .B(DB[2706]), .Z(n38295) );
  XNOR U40514 ( .A(q[5]), .B(DB[2705]), .Z(n18865) );
  IV U40515 ( .A(n18878), .Z(n38292) );
  XOR U40516 ( .A(n38296), .B(n38297), .Z(n18878) );
  XNOR U40517 ( .A(n18874), .B(n18876), .Z(n38297) );
  XNOR U40518 ( .A(q[1]), .B(DB[2701]), .Z(n18876) );
  XNOR U40519 ( .A(q[4]), .B(DB[2704]), .Z(n18874) );
  IV U40520 ( .A(n18873), .Z(n38296) );
  XNOR U40521 ( .A(n18871), .B(n38298), .Z(n18873) );
  XNOR U40522 ( .A(q[3]), .B(DB[2703]), .Z(n38298) );
  XNOR U40523 ( .A(q[2]), .B(DB[2702]), .Z(n18871) );
  XOR U40524 ( .A(n38299), .B(n18769), .Z(n18697) );
  XOR U40525 ( .A(n38300), .B(n18761), .Z(n18769) );
  XOR U40526 ( .A(n38301), .B(n18750), .Z(n18761) );
  XNOR U40527 ( .A(q[14]), .B(DB[2729]), .Z(n18750) );
  IV U40528 ( .A(n18749), .Z(n38301) );
  XNOR U40529 ( .A(n18747), .B(n38302), .Z(n18749) );
  XNOR U40530 ( .A(q[13]), .B(DB[2728]), .Z(n38302) );
  XNOR U40531 ( .A(q[12]), .B(DB[2727]), .Z(n18747) );
  IV U40532 ( .A(n18760), .Z(n38300) );
  XOR U40533 ( .A(n38303), .B(n38304), .Z(n18760) );
  XNOR U40534 ( .A(n18756), .B(n18758), .Z(n38304) );
  XNOR U40535 ( .A(q[8]), .B(DB[2723]), .Z(n18758) );
  XNOR U40536 ( .A(q[11]), .B(DB[2726]), .Z(n18756) );
  IV U40537 ( .A(n18755), .Z(n38303) );
  XNOR U40538 ( .A(n18753), .B(n38305), .Z(n18755) );
  XNOR U40539 ( .A(q[10]), .B(DB[2725]), .Z(n38305) );
  XNOR U40540 ( .A(q[9]), .B(DB[2724]), .Z(n18753) );
  IV U40541 ( .A(n18768), .Z(n38299) );
  XOR U40542 ( .A(n38306), .B(n38307), .Z(n18768) );
  XNOR U40543 ( .A(n18785), .B(n18766), .Z(n38307) );
  XNOR U40544 ( .A(q[0]), .B(DB[2715]), .Z(n18766) );
  XOR U40545 ( .A(n38308), .B(n18774), .Z(n18785) );
  XNOR U40546 ( .A(q[7]), .B(DB[2722]), .Z(n18774) );
  IV U40547 ( .A(n18773), .Z(n38308) );
  XNOR U40548 ( .A(n18771), .B(n38309), .Z(n18773) );
  XNOR U40549 ( .A(q[6]), .B(DB[2721]), .Z(n38309) );
  XNOR U40550 ( .A(q[5]), .B(DB[2720]), .Z(n18771) );
  IV U40551 ( .A(n18784), .Z(n38306) );
  XOR U40552 ( .A(n38310), .B(n38311), .Z(n18784) );
  XNOR U40553 ( .A(n18780), .B(n18782), .Z(n38311) );
  XNOR U40554 ( .A(q[1]), .B(DB[2716]), .Z(n18782) );
  XNOR U40555 ( .A(q[4]), .B(DB[2719]), .Z(n18780) );
  IV U40556 ( .A(n18779), .Z(n38310) );
  XNOR U40557 ( .A(n18777), .B(n38312), .Z(n18779) );
  XNOR U40558 ( .A(q[3]), .B(DB[2718]), .Z(n38312) );
  XNOR U40559 ( .A(q[2]), .B(DB[2717]), .Z(n18777) );
  XOR U40560 ( .A(n38313), .B(n18675), .Z(n18603) );
  XOR U40561 ( .A(n38314), .B(n18667), .Z(n18675) );
  XOR U40562 ( .A(n38315), .B(n18656), .Z(n18667) );
  XNOR U40563 ( .A(q[14]), .B(DB[2744]), .Z(n18656) );
  IV U40564 ( .A(n18655), .Z(n38315) );
  XNOR U40565 ( .A(n18653), .B(n38316), .Z(n18655) );
  XNOR U40566 ( .A(q[13]), .B(DB[2743]), .Z(n38316) );
  XNOR U40567 ( .A(q[12]), .B(DB[2742]), .Z(n18653) );
  IV U40568 ( .A(n18666), .Z(n38314) );
  XOR U40569 ( .A(n38317), .B(n38318), .Z(n18666) );
  XNOR U40570 ( .A(n18662), .B(n18664), .Z(n38318) );
  XNOR U40571 ( .A(q[8]), .B(DB[2738]), .Z(n18664) );
  XNOR U40572 ( .A(q[11]), .B(DB[2741]), .Z(n18662) );
  IV U40573 ( .A(n18661), .Z(n38317) );
  XNOR U40574 ( .A(n18659), .B(n38319), .Z(n18661) );
  XNOR U40575 ( .A(q[10]), .B(DB[2740]), .Z(n38319) );
  XNOR U40576 ( .A(q[9]), .B(DB[2739]), .Z(n18659) );
  IV U40577 ( .A(n18674), .Z(n38313) );
  XOR U40578 ( .A(n38320), .B(n38321), .Z(n18674) );
  XNOR U40579 ( .A(n18691), .B(n18672), .Z(n38321) );
  XNOR U40580 ( .A(q[0]), .B(DB[2730]), .Z(n18672) );
  XOR U40581 ( .A(n38322), .B(n18680), .Z(n18691) );
  XNOR U40582 ( .A(q[7]), .B(DB[2737]), .Z(n18680) );
  IV U40583 ( .A(n18679), .Z(n38322) );
  XNOR U40584 ( .A(n18677), .B(n38323), .Z(n18679) );
  XNOR U40585 ( .A(q[6]), .B(DB[2736]), .Z(n38323) );
  XNOR U40586 ( .A(q[5]), .B(DB[2735]), .Z(n18677) );
  IV U40587 ( .A(n18690), .Z(n38320) );
  XOR U40588 ( .A(n38324), .B(n38325), .Z(n18690) );
  XNOR U40589 ( .A(n18686), .B(n18688), .Z(n38325) );
  XNOR U40590 ( .A(q[1]), .B(DB[2731]), .Z(n18688) );
  XNOR U40591 ( .A(q[4]), .B(DB[2734]), .Z(n18686) );
  IV U40592 ( .A(n18685), .Z(n38324) );
  XNOR U40593 ( .A(n18683), .B(n38326), .Z(n18685) );
  XNOR U40594 ( .A(q[3]), .B(DB[2733]), .Z(n38326) );
  XNOR U40595 ( .A(q[2]), .B(DB[2732]), .Z(n18683) );
  XOR U40596 ( .A(n38327), .B(n18581), .Z(n18509) );
  XOR U40597 ( .A(n38328), .B(n18573), .Z(n18581) );
  XOR U40598 ( .A(n38329), .B(n18562), .Z(n18573) );
  XNOR U40599 ( .A(q[14]), .B(DB[2759]), .Z(n18562) );
  IV U40600 ( .A(n18561), .Z(n38329) );
  XNOR U40601 ( .A(n18559), .B(n38330), .Z(n18561) );
  XNOR U40602 ( .A(q[13]), .B(DB[2758]), .Z(n38330) );
  XNOR U40603 ( .A(q[12]), .B(DB[2757]), .Z(n18559) );
  IV U40604 ( .A(n18572), .Z(n38328) );
  XOR U40605 ( .A(n38331), .B(n38332), .Z(n18572) );
  XNOR U40606 ( .A(n18568), .B(n18570), .Z(n38332) );
  XNOR U40607 ( .A(q[8]), .B(DB[2753]), .Z(n18570) );
  XNOR U40608 ( .A(q[11]), .B(DB[2756]), .Z(n18568) );
  IV U40609 ( .A(n18567), .Z(n38331) );
  XNOR U40610 ( .A(n18565), .B(n38333), .Z(n18567) );
  XNOR U40611 ( .A(q[10]), .B(DB[2755]), .Z(n38333) );
  XNOR U40612 ( .A(q[9]), .B(DB[2754]), .Z(n18565) );
  IV U40613 ( .A(n18580), .Z(n38327) );
  XOR U40614 ( .A(n38334), .B(n38335), .Z(n18580) );
  XNOR U40615 ( .A(n18597), .B(n18578), .Z(n38335) );
  XNOR U40616 ( .A(q[0]), .B(DB[2745]), .Z(n18578) );
  XOR U40617 ( .A(n38336), .B(n18586), .Z(n18597) );
  XNOR U40618 ( .A(q[7]), .B(DB[2752]), .Z(n18586) );
  IV U40619 ( .A(n18585), .Z(n38336) );
  XNOR U40620 ( .A(n18583), .B(n38337), .Z(n18585) );
  XNOR U40621 ( .A(q[6]), .B(DB[2751]), .Z(n38337) );
  XNOR U40622 ( .A(q[5]), .B(DB[2750]), .Z(n18583) );
  IV U40623 ( .A(n18596), .Z(n38334) );
  XOR U40624 ( .A(n38338), .B(n38339), .Z(n18596) );
  XNOR U40625 ( .A(n18592), .B(n18594), .Z(n38339) );
  XNOR U40626 ( .A(q[1]), .B(DB[2746]), .Z(n18594) );
  XNOR U40627 ( .A(q[4]), .B(DB[2749]), .Z(n18592) );
  IV U40628 ( .A(n18591), .Z(n38338) );
  XNOR U40629 ( .A(n18589), .B(n38340), .Z(n18591) );
  XNOR U40630 ( .A(q[3]), .B(DB[2748]), .Z(n38340) );
  XNOR U40631 ( .A(q[2]), .B(DB[2747]), .Z(n18589) );
  XOR U40632 ( .A(n38341), .B(n18487), .Z(n18415) );
  XOR U40633 ( .A(n38342), .B(n18479), .Z(n18487) );
  XOR U40634 ( .A(n38343), .B(n18468), .Z(n18479) );
  XNOR U40635 ( .A(q[14]), .B(DB[2774]), .Z(n18468) );
  IV U40636 ( .A(n18467), .Z(n38343) );
  XNOR U40637 ( .A(n18465), .B(n38344), .Z(n18467) );
  XNOR U40638 ( .A(q[13]), .B(DB[2773]), .Z(n38344) );
  XNOR U40639 ( .A(q[12]), .B(DB[2772]), .Z(n18465) );
  IV U40640 ( .A(n18478), .Z(n38342) );
  XOR U40641 ( .A(n38345), .B(n38346), .Z(n18478) );
  XNOR U40642 ( .A(n18474), .B(n18476), .Z(n38346) );
  XNOR U40643 ( .A(q[8]), .B(DB[2768]), .Z(n18476) );
  XNOR U40644 ( .A(q[11]), .B(DB[2771]), .Z(n18474) );
  IV U40645 ( .A(n18473), .Z(n38345) );
  XNOR U40646 ( .A(n18471), .B(n38347), .Z(n18473) );
  XNOR U40647 ( .A(q[10]), .B(DB[2770]), .Z(n38347) );
  XNOR U40648 ( .A(q[9]), .B(DB[2769]), .Z(n18471) );
  IV U40649 ( .A(n18486), .Z(n38341) );
  XOR U40650 ( .A(n38348), .B(n38349), .Z(n18486) );
  XNOR U40651 ( .A(n18503), .B(n18484), .Z(n38349) );
  XNOR U40652 ( .A(q[0]), .B(DB[2760]), .Z(n18484) );
  XOR U40653 ( .A(n38350), .B(n18492), .Z(n18503) );
  XNOR U40654 ( .A(q[7]), .B(DB[2767]), .Z(n18492) );
  IV U40655 ( .A(n18491), .Z(n38350) );
  XNOR U40656 ( .A(n18489), .B(n38351), .Z(n18491) );
  XNOR U40657 ( .A(q[6]), .B(DB[2766]), .Z(n38351) );
  XNOR U40658 ( .A(q[5]), .B(DB[2765]), .Z(n18489) );
  IV U40659 ( .A(n18502), .Z(n38348) );
  XOR U40660 ( .A(n38352), .B(n38353), .Z(n18502) );
  XNOR U40661 ( .A(n18498), .B(n18500), .Z(n38353) );
  XNOR U40662 ( .A(q[1]), .B(DB[2761]), .Z(n18500) );
  XNOR U40663 ( .A(q[4]), .B(DB[2764]), .Z(n18498) );
  IV U40664 ( .A(n18497), .Z(n38352) );
  XNOR U40665 ( .A(n18495), .B(n38354), .Z(n18497) );
  XNOR U40666 ( .A(q[3]), .B(DB[2763]), .Z(n38354) );
  XNOR U40667 ( .A(q[2]), .B(DB[2762]), .Z(n18495) );
  XOR U40668 ( .A(n38355), .B(n18393), .Z(n18321) );
  XOR U40669 ( .A(n38356), .B(n18385), .Z(n18393) );
  XOR U40670 ( .A(n38357), .B(n18374), .Z(n18385) );
  XNOR U40671 ( .A(q[14]), .B(DB[2789]), .Z(n18374) );
  IV U40672 ( .A(n18373), .Z(n38357) );
  XNOR U40673 ( .A(n18371), .B(n38358), .Z(n18373) );
  XNOR U40674 ( .A(q[13]), .B(DB[2788]), .Z(n38358) );
  XNOR U40675 ( .A(q[12]), .B(DB[2787]), .Z(n18371) );
  IV U40676 ( .A(n18384), .Z(n38356) );
  XOR U40677 ( .A(n38359), .B(n38360), .Z(n18384) );
  XNOR U40678 ( .A(n18380), .B(n18382), .Z(n38360) );
  XNOR U40679 ( .A(q[8]), .B(DB[2783]), .Z(n18382) );
  XNOR U40680 ( .A(q[11]), .B(DB[2786]), .Z(n18380) );
  IV U40681 ( .A(n18379), .Z(n38359) );
  XNOR U40682 ( .A(n18377), .B(n38361), .Z(n18379) );
  XNOR U40683 ( .A(q[10]), .B(DB[2785]), .Z(n38361) );
  XNOR U40684 ( .A(q[9]), .B(DB[2784]), .Z(n18377) );
  IV U40685 ( .A(n18392), .Z(n38355) );
  XOR U40686 ( .A(n38362), .B(n38363), .Z(n18392) );
  XNOR U40687 ( .A(n18409), .B(n18390), .Z(n38363) );
  XNOR U40688 ( .A(q[0]), .B(DB[2775]), .Z(n18390) );
  XOR U40689 ( .A(n38364), .B(n18398), .Z(n18409) );
  XNOR U40690 ( .A(q[7]), .B(DB[2782]), .Z(n18398) );
  IV U40691 ( .A(n18397), .Z(n38364) );
  XNOR U40692 ( .A(n18395), .B(n38365), .Z(n18397) );
  XNOR U40693 ( .A(q[6]), .B(DB[2781]), .Z(n38365) );
  XNOR U40694 ( .A(q[5]), .B(DB[2780]), .Z(n18395) );
  IV U40695 ( .A(n18408), .Z(n38362) );
  XOR U40696 ( .A(n38366), .B(n38367), .Z(n18408) );
  XNOR U40697 ( .A(n18404), .B(n18406), .Z(n38367) );
  XNOR U40698 ( .A(q[1]), .B(DB[2776]), .Z(n18406) );
  XNOR U40699 ( .A(q[4]), .B(DB[2779]), .Z(n18404) );
  IV U40700 ( .A(n18403), .Z(n38366) );
  XNOR U40701 ( .A(n18401), .B(n38368), .Z(n18403) );
  XNOR U40702 ( .A(q[3]), .B(DB[2778]), .Z(n38368) );
  XNOR U40703 ( .A(q[2]), .B(DB[2777]), .Z(n18401) );
  XOR U40704 ( .A(n38369), .B(n18299), .Z(n18227) );
  XOR U40705 ( .A(n38370), .B(n18291), .Z(n18299) );
  XOR U40706 ( .A(n38371), .B(n18280), .Z(n18291) );
  XNOR U40707 ( .A(q[14]), .B(DB[2804]), .Z(n18280) );
  IV U40708 ( .A(n18279), .Z(n38371) );
  XNOR U40709 ( .A(n18277), .B(n38372), .Z(n18279) );
  XNOR U40710 ( .A(q[13]), .B(DB[2803]), .Z(n38372) );
  XNOR U40711 ( .A(q[12]), .B(DB[2802]), .Z(n18277) );
  IV U40712 ( .A(n18290), .Z(n38370) );
  XOR U40713 ( .A(n38373), .B(n38374), .Z(n18290) );
  XNOR U40714 ( .A(n18286), .B(n18288), .Z(n38374) );
  XNOR U40715 ( .A(q[8]), .B(DB[2798]), .Z(n18288) );
  XNOR U40716 ( .A(q[11]), .B(DB[2801]), .Z(n18286) );
  IV U40717 ( .A(n18285), .Z(n38373) );
  XNOR U40718 ( .A(n18283), .B(n38375), .Z(n18285) );
  XNOR U40719 ( .A(q[10]), .B(DB[2800]), .Z(n38375) );
  XNOR U40720 ( .A(q[9]), .B(DB[2799]), .Z(n18283) );
  IV U40721 ( .A(n18298), .Z(n38369) );
  XOR U40722 ( .A(n38376), .B(n38377), .Z(n18298) );
  XNOR U40723 ( .A(n18315), .B(n18296), .Z(n38377) );
  XNOR U40724 ( .A(q[0]), .B(DB[2790]), .Z(n18296) );
  XOR U40725 ( .A(n38378), .B(n18304), .Z(n18315) );
  XNOR U40726 ( .A(q[7]), .B(DB[2797]), .Z(n18304) );
  IV U40727 ( .A(n18303), .Z(n38378) );
  XNOR U40728 ( .A(n18301), .B(n38379), .Z(n18303) );
  XNOR U40729 ( .A(q[6]), .B(DB[2796]), .Z(n38379) );
  XNOR U40730 ( .A(q[5]), .B(DB[2795]), .Z(n18301) );
  IV U40731 ( .A(n18314), .Z(n38376) );
  XOR U40732 ( .A(n38380), .B(n38381), .Z(n18314) );
  XNOR U40733 ( .A(n18310), .B(n18312), .Z(n38381) );
  XNOR U40734 ( .A(q[1]), .B(DB[2791]), .Z(n18312) );
  XNOR U40735 ( .A(q[4]), .B(DB[2794]), .Z(n18310) );
  IV U40736 ( .A(n18309), .Z(n38380) );
  XNOR U40737 ( .A(n18307), .B(n38382), .Z(n18309) );
  XNOR U40738 ( .A(q[3]), .B(DB[2793]), .Z(n38382) );
  XNOR U40739 ( .A(q[2]), .B(DB[2792]), .Z(n18307) );
  XOR U40740 ( .A(n38383), .B(n18205), .Z(n18133) );
  XOR U40741 ( .A(n38384), .B(n18197), .Z(n18205) );
  XOR U40742 ( .A(n38385), .B(n18186), .Z(n18197) );
  XNOR U40743 ( .A(q[14]), .B(DB[2819]), .Z(n18186) );
  IV U40744 ( .A(n18185), .Z(n38385) );
  XNOR U40745 ( .A(n18183), .B(n38386), .Z(n18185) );
  XNOR U40746 ( .A(q[13]), .B(DB[2818]), .Z(n38386) );
  XNOR U40747 ( .A(q[12]), .B(DB[2817]), .Z(n18183) );
  IV U40748 ( .A(n18196), .Z(n38384) );
  XOR U40749 ( .A(n38387), .B(n38388), .Z(n18196) );
  XNOR U40750 ( .A(n18192), .B(n18194), .Z(n38388) );
  XNOR U40751 ( .A(q[8]), .B(DB[2813]), .Z(n18194) );
  XNOR U40752 ( .A(q[11]), .B(DB[2816]), .Z(n18192) );
  IV U40753 ( .A(n18191), .Z(n38387) );
  XNOR U40754 ( .A(n18189), .B(n38389), .Z(n18191) );
  XNOR U40755 ( .A(q[10]), .B(DB[2815]), .Z(n38389) );
  XNOR U40756 ( .A(q[9]), .B(DB[2814]), .Z(n18189) );
  IV U40757 ( .A(n18204), .Z(n38383) );
  XOR U40758 ( .A(n38390), .B(n38391), .Z(n18204) );
  XNOR U40759 ( .A(n18221), .B(n18202), .Z(n38391) );
  XNOR U40760 ( .A(q[0]), .B(DB[2805]), .Z(n18202) );
  XOR U40761 ( .A(n38392), .B(n18210), .Z(n18221) );
  XNOR U40762 ( .A(q[7]), .B(DB[2812]), .Z(n18210) );
  IV U40763 ( .A(n18209), .Z(n38392) );
  XNOR U40764 ( .A(n18207), .B(n38393), .Z(n18209) );
  XNOR U40765 ( .A(q[6]), .B(DB[2811]), .Z(n38393) );
  XNOR U40766 ( .A(q[5]), .B(DB[2810]), .Z(n18207) );
  IV U40767 ( .A(n18220), .Z(n38390) );
  XOR U40768 ( .A(n38394), .B(n38395), .Z(n18220) );
  XNOR U40769 ( .A(n18216), .B(n18218), .Z(n38395) );
  XNOR U40770 ( .A(q[1]), .B(DB[2806]), .Z(n18218) );
  XNOR U40771 ( .A(q[4]), .B(DB[2809]), .Z(n18216) );
  IV U40772 ( .A(n18215), .Z(n38394) );
  XNOR U40773 ( .A(n18213), .B(n38396), .Z(n18215) );
  XNOR U40774 ( .A(q[3]), .B(DB[2808]), .Z(n38396) );
  XNOR U40775 ( .A(q[2]), .B(DB[2807]), .Z(n18213) );
  XOR U40776 ( .A(n38397), .B(n18111), .Z(n18039) );
  XOR U40777 ( .A(n38398), .B(n18103), .Z(n18111) );
  XOR U40778 ( .A(n38399), .B(n18092), .Z(n18103) );
  XNOR U40779 ( .A(q[14]), .B(DB[2834]), .Z(n18092) );
  IV U40780 ( .A(n18091), .Z(n38399) );
  XNOR U40781 ( .A(n18089), .B(n38400), .Z(n18091) );
  XNOR U40782 ( .A(q[13]), .B(DB[2833]), .Z(n38400) );
  XNOR U40783 ( .A(q[12]), .B(DB[2832]), .Z(n18089) );
  IV U40784 ( .A(n18102), .Z(n38398) );
  XOR U40785 ( .A(n38401), .B(n38402), .Z(n18102) );
  XNOR U40786 ( .A(n18098), .B(n18100), .Z(n38402) );
  XNOR U40787 ( .A(q[8]), .B(DB[2828]), .Z(n18100) );
  XNOR U40788 ( .A(q[11]), .B(DB[2831]), .Z(n18098) );
  IV U40789 ( .A(n18097), .Z(n38401) );
  XNOR U40790 ( .A(n18095), .B(n38403), .Z(n18097) );
  XNOR U40791 ( .A(q[10]), .B(DB[2830]), .Z(n38403) );
  XNOR U40792 ( .A(q[9]), .B(DB[2829]), .Z(n18095) );
  IV U40793 ( .A(n18110), .Z(n38397) );
  XOR U40794 ( .A(n38404), .B(n38405), .Z(n18110) );
  XNOR U40795 ( .A(n18127), .B(n18108), .Z(n38405) );
  XNOR U40796 ( .A(q[0]), .B(DB[2820]), .Z(n18108) );
  XOR U40797 ( .A(n38406), .B(n18116), .Z(n18127) );
  XNOR U40798 ( .A(q[7]), .B(DB[2827]), .Z(n18116) );
  IV U40799 ( .A(n18115), .Z(n38406) );
  XNOR U40800 ( .A(n18113), .B(n38407), .Z(n18115) );
  XNOR U40801 ( .A(q[6]), .B(DB[2826]), .Z(n38407) );
  XNOR U40802 ( .A(q[5]), .B(DB[2825]), .Z(n18113) );
  IV U40803 ( .A(n18126), .Z(n38404) );
  XOR U40804 ( .A(n38408), .B(n38409), .Z(n18126) );
  XNOR U40805 ( .A(n18122), .B(n18124), .Z(n38409) );
  XNOR U40806 ( .A(q[1]), .B(DB[2821]), .Z(n18124) );
  XNOR U40807 ( .A(q[4]), .B(DB[2824]), .Z(n18122) );
  IV U40808 ( .A(n18121), .Z(n38408) );
  XNOR U40809 ( .A(n18119), .B(n38410), .Z(n18121) );
  XNOR U40810 ( .A(q[3]), .B(DB[2823]), .Z(n38410) );
  XNOR U40811 ( .A(q[2]), .B(DB[2822]), .Z(n18119) );
  XOR U40812 ( .A(n38411), .B(n18017), .Z(n17945) );
  XOR U40813 ( .A(n38412), .B(n18009), .Z(n18017) );
  XOR U40814 ( .A(n38413), .B(n17998), .Z(n18009) );
  XNOR U40815 ( .A(q[14]), .B(DB[2849]), .Z(n17998) );
  IV U40816 ( .A(n17997), .Z(n38413) );
  XNOR U40817 ( .A(n17995), .B(n38414), .Z(n17997) );
  XNOR U40818 ( .A(q[13]), .B(DB[2848]), .Z(n38414) );
  XNOR U40819 ( .A(q[12]), .B(DB[2847]), .Z(n17995) );
  IV U40820 ( .A(n18008), .Z(n38412) );
  XOR U40821 ( .A(n38415), .B(n38416), .Z(n18008) );
  XNOR U40822 ( .A(n18004), .B(n18006), .Z(n38416) );
  XNOR U40823 ( .A(q[8]), .B(DB[2843]), .Z(n18006) );
  XNOR U40824 ( .A(q[11]), .B(DB[2846]), .Z(n18004) );
  IV U40825 ( .A(n18003), .Z(n38415) );
  XNOR U40826 ( .A(n18001), .B(n38417), .Z(n18003) );
  XNOR U40827 ( .A(q[10]), .B(DB[2845]), .Z(n38417) );
  XNOR U40828 ( .A(q[9]), .B(DB[2844]), .Z(n18001) );
  IV U40829 ( .A(n18016), .Z(n38411) );
  XOR U40830 ( .A(n38418), .B(n38419), .Z(n18016) );
  XNOR U40831 ( .A(n18033), .B(n18014), .Z(n38419) );
  XNOR U40832 ( .A(q[0]), .B(DB[2835]), .Z(n18014) );
  XOR U40833 ( .A(n38420), .B(n18022), .Z(n18033) );
  XNOR U40834 ( .A(q[7]), .B(DB[2842]), .Z(n18022) );
  IV U40835 ( .A(n18021), .Z(n38420) );
  XNOR U40836 ( .A(n18019), .B(n38421), .Z(n18021) );
  XNOR U40837 ( .A(q[6]), .B(DB[2841]), .Z(n38421) );
  XNOR U40838 ( .A(q[5]), .B(DB[2840]), .Z(n18019) );
  IV U40839 ( .A(n18032), .Z(n38418) );
  XOR U40840 ( .A(n38422), .B(n38423), .Z(n18032) );
  XNOR U40841 ( .A(n18028), .B(n18030), .Z(n38423) );
  XNOR U40842 ( .A(q[1]), .B(DB[2836]), .Z(n18030) );
  XNOR U40843 ( .A(q[4]), .B(DB[2839]), .Z(n18028) );
  IV U40844 ( .A(n18027), .Z(n38422) );
  XNOR U40845 ( .A(n18025), .B(n38424), .Z(n18027) );
  XNOR U40846 ( .A(q[3]), .B(DB[2838]), .Z(n38424) );
  XNOR U40847 ( .A(q[2]), .B(DB[2837]), .Z(n18025) );
  XOR U40848 ( .A(n38425), .B(n17923), .Z(n17851) );
  XOR U40849 ( .A(n38426), .B(n17915), .Z(n17923) );
  XOR U40850 ( .A(n38427), .B(n17904), .Z(n17915) );
  XNOR U40851 ( .A(q[14]), .B(DB[2864]), .Z(n17904) );
  IV U40852 ( .A(n17903), .Z(n38427) );
  XNOR U40853 ( .A(n17901), .B(n38428), .Z(n17903) );
  XNOR U40854 ( .A(q[13]), .B(DB[2863]), .Z(n38428) );
  XNOR U40855 ( .A(q[12]), .B(DB[2862]), .Z(n17901) );
  IV U40856 ( .A(n17914), .Z(n38426) );
  XOR U40857 ( .A(n38429), .B(n38430), .Z(n17914) );
  XNOR U40858 ( .A(n17910), .B(n17912), .Z(n38430) );
  XNOR U40859 ( .A(q[8]), .B(DB[2858]), .Z(n17912) );
  XNOR U40860 ( .A(q[11]), .B(DB[2861]), .Z(n17910) );
  IV U40861 ( .A(n17909), .Z(n38429) );
  XNOR U40862 ( .A(n17907), .B(n38431), .Z(n17909) );
  XNOR U40863 ( .A(q[10]), .B(DB[2860]), .Z(n38431) );
  XNOR U40864 ( .A(q[9]), .B(DB[2859]), .Z(n17907) );
  IV U40865 ( .A(n17922), .Z(n38425) );
  XOR U40866 ( .A(n38432), .B(n38433), .Z(n17922) );
  XNOR U40867 ( .A(n17939), .B(n17920), .Z(n38433) );
  XNOR U40868 ( .A(q[0]), .B(DB[2850]), .Z(n17920) );
  XOR U40869 ( .A(n38434), .B(n17928), .Z(n17939) );
  XNOR U40870 ( .A(q[7]), .B(DB[2857]), .Z(n17928) );
  IV U40871 ( .A(n17927), .Z(n38434) );
  XNOR U40872 ( .A(n17925), .B(n38435), .Z(n17927) );
  XNOR U40873 ( .A(q[6]), .B(DB[2856]), .Z(n38435) );
  XNOR U40874 ( .A(q[5]), .B(DB[2855]), .Z(n17925) );
  IV U40875 ( .A(n17938), .Z(n38432) );
  XOR U40876 ( .A(n38436), .B(n38437), .Z(n17938) );
  XNOR U40877 ( .A(n17934), .B(n17936), .Z(n38437) );
  XNOR U40878 ( .A(q[1]), .B(DB[2851]), .Z(n17936) );
  XNOR U40879 ( .A(q[4]), .B(DB[2854]), .Z(n17934) );
  IV U40880 ( .A(n17933), .Z(n38436) );
  XNOR U40881 ( .A(n17931), .B(n38438), .Z(n17933) );
  XNOR U40882 ( .A(q[3]), .B(DB[2853]), .Z(n38438) );
  XNOR U40883 ( .A(q[2]), .B(DB[2852]), .Z(n17931) );
  XOR U40884 ( .A(n38439), .B(n17829), .Z(n17757) );
  XOR U40885 ( .A(n38440), .B(n17821), .Z(n17829) );
  XOR U40886 ( .A(n38441), .B(n17810), .Z(n17821) );
  XNOR U40887 ( .A(q[14]), .B(DB[2879]), .Z(n17810) );
  IV U40888 ( .A(n17809), .Z(n38441) );
  XNOR U40889 ( .A(n17807), .B(n38442), .Z(n17809) );
  XNOR U40890 ( .A(q[13]), .B(DB[2878]), .Z(n38442) );
  XNOR U40891 ( .A(q[12]), .B(DB[2877]), .Z(n17807) );
  IV U40892 ( .A(n17820), .Z(n38440) );
  XOR U40893 ( .A(n38443), .B(n38444), .Z(n17820) );
  XNOR U40894 ( .A(n17816), .B(n17818), .Z(n38444) );
  XNOR U40895 ( .A(q[8]), .B(DB[2873]), .Z(n17818) );
  XNOR U40896 ( .A(q[11]), .B(DB[2876]), .Z(n17816) );
  IV U40897 ( .A(n17815), .Z(n38443) );
  XNOR U40898 ( .A(n17813), .B(n38445), .Z(n17815) );
  XNOR U40899 ( .A(q[10]), .B(DB[2875]), .Z(n38445) );
  XNOR U40900 ( .A(q[9]), .B(DB[2874]), .Z(n17813) );
  IV U40901 ( .A(n17828), .Z(n38439) );
  XOR U40902 ( .A(n38446), .B(n38447), .Z(n17828) );
  XNOR U40903 ( .A(n17845), .B(n17826), .Z(n38447) );
  XNOR U40904 ( .A(q[0]), .B(DB[2865]), .Z(n17826) );
  XOR U40905 ( .A(n38448), .B(n17834), .Z(n17845) );
  XNOR U40906 ( .A(q[7]), .B(DB[2872]), .Z(n17834) );
  IV U40907 ( .A(n17833), .Z(n38448) );
  XNOR U40908 ( .A(n17831), .B(n38449), .Z(n17833) );
  XNOR U40909 ( .A(q[6]), .B(DB[2871]), .Z(n38449) );
  XNOR U40910 ( .A(q[5]), .B(DB[2870]), .Z(n17831) );
  IV U40911 ( .A(n17844), .Z(n38446) );
  XOR U40912 ( .A(n38450), .B(n38451), .Z(n17844) );
  XNOR U40913 ( .A(n17840), .B(n17842), .Z(n38451) );
  XNOR U40914 ( .A(q[1]), .B(DB[2866]), .Z(n17842) );
  XNOR U40915 ( .A(q[4]), .B(DB[2869]), .Z(n17840) );
  IV U40916 ( .A(n17839), .Z(n38450) );
  XNOR U40917 ( .A(n17837), .B(n38452), .Z(n17839) );
  XNOR U40918 ( .A(q[3]), .B(DB[2868]), .Z(n38452) );
  XNOR U40919 ( .A(q[2]), .B(DB[2867]), .Z(n17837) );
  XOR U40920 ( .A(n38453), .B(n17735), .Z(n17663) );
  XOR U40921 ( .A(n38454), .B(n17727), .Z(n17735) );
  XOR U40922 ( .A(n38455), .B(n17716), .Z(n17727) );
  XNOR U40923 ( .A(q[14]), .B(DB[2894]), .Z(n17716) );
  IV U40924 ( .A(n17715), .Z(n38455) );
  XNOR U40925 ( .A(n17713), .B(n38456), .Z(n17715) );
  XNOR U40926 ( .A(q[13]), .B(DB[2893]), .Z(n38456) );
  XNOR U40927 ( .A(q[12]), .B(DB[2892]), .Z(n17713) );
  IV U40928 ( .A(n17726), .Z(n38454) );
  XOR U40929 ( .A(n38457), .B(n38458), .Z(n17726) );
  XNOR U40930 ( .A(n17722), .B(n17724), .Z(n38458) );
  XNOR U40931 ( .A(q[8]), .B(DB[2888]), .Z(n17724) );
  XNOR U40932 ( .A(q[11]), .B(DB[2891]), .Z(n17722) );
  IV U40933 ( .A(n17721), .Z(n38457) );
  XNOR U40934 ( .A(n17719), .B(n38459), .Z(n17721) );
  XNOR U40935 ( .A(q[10]), .B(DB[2890]), .Z(n38459) );
  XNOR U40936 ( .A(q[9]), .B(DB[2889]), .Z(n17719) );
  IV U40937 ( .A(n17734), .Z(n38453) );
  XOR U40938 ( .A(n38460), .B(n38461), .Z(n17734) );
  XNOR U40939 ( .A(n17751), .B(n17732), .Z(n38461) );
  XNOR U40940 ( .A(q[0]), .B(DB[2880]), .Z(n17732) );
  XOR U40941 ( .A(n38462), .B(n17740), .Z(n17751) );
  XNOR U40942 ( .A(q[7]), .B(DB[2887]), .Z(n17740) );
  IV U40943 ( .A(n17739), .Z(n38462) );
  XNOR U40944 ( .A(n17737), .B(n38463), .Z(n17739) );
  XNOR U40945 ( .A(q[6]), .B(DB[2886]), .Z(n38463) );
  XNOR U40946 ( .A(q[5]), .B(DB[2885]), .Z(n17737) );
  IV U40947 ( .A(n17750), .Z(n38460) );
  XOR U40948 ( .A(n38464), .B(n38465), .Z(n17750) );
  XNOR U40949 ( .A(n17746), .B(n17748), .Z(n38465) );
  XNOR U40950 ( .A(q[1]), .B(DB[2881]), .Z(n17748) );
  XNOR U40951 ( .A(q[4]), .B(DB[2884]), .Z(n17746) );
  IV U40952 ( .A(n17745), .Z(n38464) );
  XNOR U40953 ( .A(n17743), .B(n38466), .Z(n17745) );
  XNOR U40954 ( .A(q[3]), .B(DB[2883]), .Z(n38466) );
  XNOR U40955 ( .A(q[2]), .B(DB[2882]), .Z(n17743) );
  XOR U40956 ( .A(n38467), .B(n17641), .Z(n17569) );
  XOR U40957 ( .A(n38468), .B(n17633), .Z(n17641) );
  XOR U40958 ( .A(n38469), .B(n17622), .Z(n17633) );
  XNOR U40959 ( .A(q[14]), .B(DB[2909]), .Z(n17622) );
  IV U40960 ( .A(n17621), .Z(n38469) );
  XNOR U40961 ( .A(n17619), .B(n38470), .Z(n17621) );
  XNOR U40962 ( .A(q[13]), .B(DB[2908]), .Z(n38470) );
  XNOR U40963 ( .A(q[12]), .B(DB[2907]), .Z(n17619) );
  IV U40964 ( .A(n17632), .Z(n38468) );
  XOR U40965 ( .A(n38471), .B(n38472), .Z(n17632) );
  XNOR U40966 ( .A(n17628), .B(n17630), .Z(n38472) );
  XNOR U40967 ( .A(q[8]), .B(DB[2903]), .Z(n17630) );
  XNOR U40968 ( .A(q[11]), .B(DB[2906]), .Z(n17628) );
  IV U40969 ( .A(n17627), .Z(n38471) );
  XNOR U40970 ( .A(n17625), .B(n38473), .Z(n17627) );
  XNOR U40971 ( .A(q[10]), .B(DB[2905]), .Z(n38473) );
  XNOR U40972 ( .A(q[9]), .B(DB[2904]), .Z(n17625) );
  IV U40973 ( .A(n17640), .Z(n38467) );
  XOR U40974 ( .A(n38474), .B(n38475), .Z(n17640) );
  XNOR U40975 ( .A(n17657), .B(n17638), .Z(n38475) );
  XNOR U40976 ( .A(q[0]), .B(DB[2895]), .Z(n17638) );
  XOR U40977 ( .A(n38476), .B(n17646), .Z(n17657) );
  XNOR U40978 ( .A(q[7]), .B(DB[2902]), .Z(n17646) );
  IV U40979 ( .A(n17645), .Z(n38476) );
  XNOR U40980 ( .A(n17643), .B(n38477), .Z(n17645) );
  XNOR U40981 ( .A(q[6]), .B(DB[2901]), .Z(n38477) );
  XNOR U40982 ( .A(q[5]), .B(DB[2900]), .Z(n17643) );
  IV U40983 ( .A(n17656), .Z(n38474) );
  XOR U40984 ( .A(n38478), .B(n38479), .Z(n17656) );
  XNOR U40985 ( .A(n17652), .B(n17654), .Z(n38479) );
  XNOR U40986 ( .A(q[1]), .B(DB[2896]), .Z(n17654) );
  XNOR U40987 ( .A(q[4]), .B(DB[2899]), .Z(n17652) );
  IV U40988 ( .A(n17651), .Z(n38478) );
  XNOR U40989 ( .A(n17649), .B(n38480), .Z(n17651) );
  XNOR U40990 ( .A(q[3]), .B(DB[2898]), .Z(n38480) );
  XNOR U40991 ( .A(q[2]), .B(DB[2897]), .Z(n17649) );
  XOR U40992 ( .A(n38481), .B(n17547), .Z(n17475) );
  XOR U40993 ( .A(n38482), .B(n17539), .Z(n17547) );
  XOR U40994 ( .A(n38483), .B(n17528), .Z(n17539) );
  XNOR U40995 ( .A(q[14]), .B(DB[2924]), .Z(n17528) );
  IV U40996 ( .A(n17527), .Z(n38483) );
  XNOR U40997 ( .A(n17525), .B(n38484), .Z(n17527) );
  XNOR U40998 ( .A(q[13]), .B(DB[2923]), .Z(n38484) );
  XNOR U40999 ( .A(q[12]), .B(DB[2922]), .Z(n17525) );
  IV U41000 ( .A(n17538), .Z(n38482) );
  XOR U41001 ( .A(n38485), .B(n38486), .Z(n17538) );
  XNOR U41002 ( .A(n17534), .B(n17536), .Z(n38486) );
  XNOR U41003 ( .A(q[8]), .B(DB[2918]), .Z(n17536) );
  XNOR U41004 ( .A(q[11]), .B(DB[2921]), .Z(n17534) );
  IV U41005 ( .A(n17533), .Z(n38485) );
  XNOR U41006 ( .A(n17531), .B(n38487), .Z(n17533) );
  XNOR U41007 ( .A(q[10]), .B(DB[2920]), .Z(n38487) );
  XNOR U41008 ( .A(q[9]), .B(DB[2919]), .Z(n17531) );
  IV U41009 ( .A(n17546), .Z(n38481) );
  XOR U41010 ( .A(n38488), .B(n38489), .Z(n17546) );
  XNOR U41011 ( .A(n17563), .B(n17544), .Z(n38489) );
  XNOR U41012 ( .A(q[0]), .B(DB[2910]), .Z(n17544) );
  XOR U41013 ( .A(n38490), .B(n17552), .Z(n17563) );
  XNOR U41014 ( .A(q[7]), .B(DB[2917]), .Z(n17552) );
  IV U41015 ( .A(n17551), .Z(n38490) );
  XNOR U41016 ( .A(n17549), .B(n38491), .Z(n17551) );
  XNOR U41017 ( .A(q[6]), .B(DB[2916]), .Z(n38491) );
  XNOR U41018 ( .A(q[5]), .B(DB[2915]), .Z(n17549) );
  IV U41019 ( .A(n17562), .Z(n38488) );
  XOR U41020 ( .A(n38492), .B(n38493), .Z(n17562) );
  XNOR U41021 ( .A(n17558), .B(n17560), .Z(n38493) );
  XNOR U41022 ( .A(q[1]), .B(DB[2911]), .Z(n17560) );
  XNOR U41023 ( .A(q[4]), .B(DB[2914]), .Z(n17558) );
  IV U41024 ( .A(n17557), .Z(n38492) );
  XNOR U41025 ( .A(n17555), .B(n38494), .Z(n17557) );
  XNOR U41026 ( .A(q[3]), .B(DB[2913]), .Z(n38494) );
  XNOR U41027 ( .A(q[2]), .B(DB[2912]), .Z(n17555) );
  XOR U41028 ( .A(n38495), .B(n17453), .Z(n17381) );
  XOR U41029 ( .A(n38496), .B(n17445), .Z(n17453) );
  XOR U41030 ( .A(n38497), .B(n17434), .Z(n17445) );
  XNOR U41031 ( .A(q[14]), .B(DB[2939]), .Z(n17434) );
  IV U41032 ( .A(n17433), .Z(n38497) );
  XNOR U41033 ( .A(n17431), .B(n38498), .Z(n17433) );
  XNOR U41034 ( .A(q[13]), .B(DB[2938]), .Z(n38498) );
  XNOR U41035 ( .A(q[12]), .B(DB[2937]), .Z(n17431) );
  IV U41036 ( .A(n17444), .Z(n38496) );
  XOR U41037 ( .A(n38499), .B(n38500), .Z(n17444) );
  XNOR U41038 ( .A(n17440), .B(n17442), .Z(n38500) );
  XNOR U41039 ( .A(q[8]), .B(DB[2933]), .Z(n17442) );
  XNOR U41040 ( .A(q[11]), .B(DB[2936]), .Z(n17440) );
  IV U41041 ( .A(n17439), .Z(n38499) );
  XNOR U41042 ( .A(n17437), .B(n38501), .Z(n17439) );
  XNOR U41043 ( .A(q[10]), .B(DB[2935]), .Z(n38501) );
  XNOR U41044 ( .A(q[9]), .B(DB[2934]), .Z(n17437) );
  IV U41045 ( .A(n17452), .Z(n38495) );
  XOR U41046 ( .A(n38502), .B(n38503), .Z(n17452) );
  XNOR U41047 ( .A(n17469), .B(n17450), .Z(n38503) );
  XNOR U41048 ( .A(q[0]), .B(DB[2925]), .Z(n17450) );
  XOR U41049 ( .A(n38504), .B(n17458), .Z(n17469) );
  XNOR U41050 ( .A(q[7]), .B(DB[2932]), .Z(n17458) );
  IV U41051 ( .A(n17457), .Z(n38504) );
  XNOR U41052 ( .A(n17455), .B(n38505), .Z(n17457) );
  XNOR U41053 ( .A(q[6]), .B(DB[2931]), .Z(n38505) );
  XNOR U41054 ( .A(q[5]), .B(DB[2930]), .Z(n17455) );
  IV U41055 ( .A(n17468), .Z(n38502) );
  XOR U41056 ( .A(n38506), .B(n38507), .Z(n17468) );
  XNOR U41057 ( .A(n17464), .B(n17466), .Z(n38507) );
  XNOR U41058 ( .A(q[1]), .B(DB[2926]), .Z(n17466) );
  XNOR U41059 ( .A(q[4]), .B(DB[2929]), .Z(n17464) );
  IV U41060 ( .A(n17463), .Z(n38506) );
  XNOR U41061 ( .A(n17461), .B(n38508), .Z(n17463) );
  XNOR U41062 ( .A(q[3]), .B(DB[2928]), .Z(n38508) );
  XNOR U41063 ( .A(q[2]), .B(DB[2927]), .Z(n17461) );
  XOR U41064 ( .A(n38509), .B(n17359), .Z(n17287) );
  XOR U41065 ( .A(n38510), .B(n17351), .Z(n17359) );
  XOR U41066 ( .A(n38511), .B(n17340), .Z(n17351) );
  XNOR U41067 ( .A(q[14]), .B(DB[2954]), .Z(n17340) );
  IV U41068 ( .A(n17339), .Z(n38511) );
  XNOR U41069 ( .A(n17337), .B(n38512), .Z(n17339) );
  XNOR U41070 ( .A(q[13]), .B(DB[2953]), .Z(n38512) );
  XNOR U41071 ( .A(q[12]), .B(DB[2952]), .Z(n17337) );
  IV U41072 ( .A(n17350), .Z(n38510) );
  XOR U41073 ( .A(n38513), .B(n38514), .Z(n17350) );
  XNOR U41074 ( .A(n17346), .B(n17348), .Z(n38514) );
  XNOR U41075 ( .A(q[8]), .B(DB[2948]), .Z(n17348) );
  XNOR U41076 ( .A(q[11]), .B(DB[2951]), .Z(n17346) );
  IV U41077 ( .A(n17345), .Z(n38513) );
  XNOR U41078 ( .A(n17343), .B(n38515), .Z(n17345) );
  XNOR U41079 ( .A(q[10]), .B(DB[2950]), .Z(n38515) );
  XNOR U41080 ( .A(q[9]), .B(DB[2949]), .Z(n17343) );
  IV U41081 ( .A(n17358), .Z(n38509) );
  XOR U41082 ( .A(n38516), .B(n38517), .Z(n17358) );
  XNOR U41083 ( .A(n17375), .B(n17356), .Z(n38517) );
  XNOR U41084 ( .A(q[0]), .B(DB[2940]), .Z(n17356) );
  XOR U41085 ( .A(n38518), .B(n17364), .Z(n17375) );
  XNOR U41086 ( .A(q[7]), .B(DB[2947]), .Z(n17364) );
  IV U41087 ( .A(n17363), .Z(n38518) );
  XNOR U41088 ( .A(n17361), .B(n38519), .Z(n17363) );
  XNOR U41089 ( .A(q[6]), .B(DB[2946]), .Z(n38519) );
  XNOR U41090 ( .A(q[5]), .B(DB[2945]), .Z(n17361) );
  IV U41091 ( .A(n17374), .Z(n38516) );
  XOR U41092 ( .A(n38520), .B(n38521), .Z(n17374) );
  XNOR U41093 ( .A(n17370), .B(n17372), .Z(n38521) );
  XNOR U41094 ( .A(q[1]), .B(DB[2941]), .Z(n17372) );
  XNOR U41095 ( .A(q[4]), .B(DB[2944]), .Z(n17370) );
  IV U41096 ( .A(n17369), .Z(n38520) );
  XNOR U41097 ( .A(n17367), .B(n38522), .Z(n17369) );
  XNOR U41098 ( .A(q[3]), .B(DB[2943]), .Z(n38522) );
  XNOR U41099 ( .A(q[2]), .B(DB[2942]), .Z(n17367) );
  XOR U41100 ( .A(n38523), .B(n17265), .Z(n17193) );
  XOR U41101 ( .A(n38524), .B(n17257), .Z(n17265) );
  XOR U41102 ( .A(n38525), .B(n17246), .Z(n17257) );
  XNOR U41103 ( .A(q[14]), .B(DB[2969]), .Z(n17246) );
  IV U41104 ( .A(n17245), .Z(n38525) );
  XNOR U41105 ( .A(n17243), .B(n38526), .Z(n17245) );
  XNOR U41106 ( .A(q[13]), .B(DB[2968]), .Z(n38526) );
  XNOR U41107 ( .A(q[12]), .B(DB[2967]), .Z(n17243) );
  IV U41108 ( .A(n17256), .Z(n38524) );
  XOR U41109 ( .A(n38527), .B(n38528), .Z(n17256) );
  XNOR U41110 ( .A(n17252), .B(n17254), .Z(n38528) );
  XNOR U41111 ( .A(q[8]), .B(DB[2963]), .Z(n17254) );
  XNOR U41112 ( .A(q[11]), .B(DB[2966]), .Z(n17252) );
  IV U41113 ( .A(n17251), .Z(n38527) );
  XNOR U41114 ( .A(n17249), .B(n38529), .Z(n17251) );
  XNOR U41115 ( .A(q[10]), .B(DB[2965]), .Z(n38529) );
  XNOR U41116 ( .A(q[9]), .B(DB[2964]), .Z(n17249) );
  IV U41117 ( .A(n17264), .Z(n38523) );
  XOR U41118 ( .A(n38530), .B(n38531), .Z(n17264) );
  XNOR U41119 ( .A(n17281), .B(n17262), .Z(n38531) );
  XNOR U41120 ( .A(q[0]), .B(DB[2955]), .Z(n17262) );
  XOR U41121 ( .A(n38532), .B(n17270), .Z(n17281) );
  XNOR U41122 ( .A(q[7]), .B(DB[2962]), .Z(n17270) );
  IV U41123 ( .A(n17269), .Z(n38532) );
  XNOR U41124 ( .A(n17267), .B(n38533), .Z(n17269) );
  XNOR U41125 ( .A(q[6]), .B(DB[2961]), .Z(n38533) );
  XNOR U41126 ( .A(q[5]), .B(DB[2960]), .Z(n17267) );
  IV U41127 ( .A(n17280), .Z(n38530) );
  XOR U41128 ( .A(n38534), .B(n38535), .Z(n17280) );
  XNOR U41129 ( .A(n17276), .B(n17278), .Z(n38535) );
  XNOR U41130 ( .A(q[1]), .B(DB[2956]), .Z(n17278) );
  XNOR U41131 ( .A(q[4]), .B(DB[2959]), .Z(n17276) );
  IV U41132 ( .A(n17275), .Z(n38534) );
  XNOR U41133 ( .A(n17273), .B(n38536), .Z(n17275) );
  XNOR U41134 ( .A(q[3]), .B(DB[2958]), .Z(n38536) );
  XNOR U41135 ( .A(q[2]), .B(DB[2957]), .Z(n17273) );
  XOR U41136 ( .A(n38537), .B(n17171), .Z(n17099) );
  XOR U41137 ( .A(n38538), .B(n17163), .Z(n17171) );
  XOR U41138 ( .A(n38539), .B(n17152), .Z(n17163) );
  XNOR U41139 ( .A(q[14]), .B(DB[2984]), .Z(n17152) );
  IV U41140 ( .A(n17151), .Z(n38539) );
  XNOR U41141 ( .A(n17149), .B(n38540), .Z(n17151) );
  XNOR U41142 ( .A(q[13]), .B(DB[2983]), .Z(n38540) );
  XNOR U41143 ( .A(q[12]), .B(DB[2982]), .Z(n17149) );
  IV U41144 ( .A(n17162), .Z(n38538) );
  XOR U41145 ( .A(n38541), .B(n38542), .Z(n17162) );
  XNOR U41146 ( .A(n17158), .B(n17160), .Z(n38542) );
  XNOR U41147 ( .A(q[8]), .B(DB[2978]), .Z(n17160) );
  XNOR U41148 ( .A(q[11]), .B(DB[2981]), .Z(n17158) );
  IV U41149 ( .A(n17157), .Z(n38541) );
  XNOR U41150 ( .A(n17155), .B(n38543), .Z(n17157) );
  XNOR U41151 ( .A(q[10]), .B(DB[2980]), .Z(n38543) );
  XNOR U41152 ( .A(q[9]), .B(DB[2979]), .Z(n17155) );
  IV U41153 ( .A(n17170), .Z(n38537) );
  XOR U41154 ( .A(n38544), .B(n38545), .Z(n17170) );
  XNOR U41155 ( .A(n17187), .B(n17168), .Z(n38545) );
  XNOR U41156 ( .A(q[0]), .B(DB[2970]), .Z(n17168) );
  XOR U41157 ( .A(n38546), .B(n17176), .Z(n17187) );
  XNOR U41158 ( .A(q[7]), .B(DB[2977]), .Z(n17176) );
  IV U41159 ( .A(n17175), .Z(n38546) );
  XNOR U41160 ( .A(n17173), .B(n38547), .Z(n17175) );
  XNOR U41161 ( .A(q[6]), .B(DB[2976]), .Z(n38547) );
  XNOR U41162 ( .A(q[5]), .B(DB[2975]), .Z(n17173) );
  IV U41163 ( .A(n17186), .Z(n38544) );
  XOR U41164 ( .A(n38548), .B(n38549), .Z(n17186) );
  XNOR U41165 ( .A(n17182), .B(n17184), .Z(n38549) );
  XNOR U41166 ( .A(q[1]), .B(DB[2971]), .Z(n17184) );
  XNOR U41167 ( .A(q[4]), .B(DB[2974]), .Z(n17182) );
  IV U41168 ( .A(n17181), .Z(n38548) );
  XNOR U41169 ( .A(n17179), .B(n38550), .Z(n17181) );
  XNOR U41170 ( .A(q[3]), .B(DB[2973]), .Z(n38550) );
  XNOR U41171 ( .A(q[2]), .B(DB[2972]), .Z(n17179) );
  XOR U41172 ( .A(n38551), .B(n17077), .Z(n17005) );
  XOR U41173 ( .A(n38552), .B(n17069), .Z(n17077) );
  XOR U41174 ( .A(n38553), .B(n17058), .Z(n17069) );
  XNOR U41175 ( .A(q[14]), .B(DB[2999]), .Z(n17058) );
  IV U41176 ( .A(n17057), .Z(n38553) );
  XNOR U41177 ( .A(n17055), .B(n38554), .Z(n17057) );
  XNOR U41178 ( .A(q[13]), .B(DB[2998]), .Z(n38554) );
  XNOR U41179 ( .A(q[12]), .B(DB[2997]), .Z(n17055) );
  IV U41180 ( .A(n17068), .Z(n38552) );
  XOR U41181 ( .A(n38555), .B(n38556), .Z(n17068) );
  XNOR U41182 ( .A(n17064), .B(n17066), .Z(n38556) );
  XNOR U41183 ( .A(q[8]), .B(DB[2993]), .Z(n17066) );
  XNOR U41184 ( .A(q[11]), .B(DB[2996]), .Z(n17064) );
  IV U41185 ( .A(n17063), .Z(n38555) );
  XNOR U41186 ( .A(n17061), .B(n38557), .Z(n17063) );
  XNOR U41187 ( .A(q[10]), .B(DB[2995]), .Z(n38557) );
  XNOR U41188 ( .A(q[9]), .B(DB[2994]), .Z(n17061) );
  IV U41189 ( .A(n17076), .Z(n38551) );
  XOR U41190 ( .A(n38558), .B(n38559), .Z(n17076) );
  XNOR U41191 ( .A(n17093), .B(n17074), .Z(n38559) );
  XNOR U41192 ( .A(q[0]), .B(DB[2985]), .Z(n17074) );
  XOR U41193 ( .A(n38560), .B(n17082), .Z(n17093) );
  XNOR U41194 ( .A(q[7]), .B(DB[2992]), .Z(n17082) );
  IV U41195 ( .A(n17081), .Z(n38560) );
  XNOR U41196 ( .A(n17079), .B(n38561), .Z(n17081) );
  XNOR U41197 ( .A(q[6]), .B(DB[2991]), .Z(n38561) );
  XNOR U41198 ( .A(q[5]), .B(DB[2990]), .Z(n17079) );
  IV U41199 ( .A(n17092), .Z(n38558) );
  XOR U41200 ( .A(n38562), .B(n38563), .Z(n17092) );
  XNOR U41201 ( .A(n17088), .B(n17090), .Z(n38563) );
  XNOR U41202 ( .A(q[1]), .B(DB[2986]), .Z(n17090) );
  XNOR U41203 ( .A(q[4]), .B(DB[2989]), .Z(n17088) );
  IV U41204 ( .A(n17087), .Z(n38562) );
  XNOR U41205 ( .A(n17085), .B(n38564), .Z(n17087) );
  XNOR U41206 ( .A(q[3]), .B(DB[2988]), .Z(n38564) );
  XNOR U41207 ( .A(q[2]), .B(DB[2987]), .Z(n17085) );
  XOR U41208 ( .A(n38565), .B(n16983), .Z(n16911) );
  XOR U41209 ( .A(n38566), .B(n16975), .Z(n16983) );
  XOR U41210 ( .A(n38567), .B(n16964), .Z(n16975) );
  XNOR U41211 ( .A(q[14]), .B(DB[3014]), .Z(n16964) );
  IV U41212 ( .A(n16963), .Z(n38567) );
  XNOR U41213 ( .A(n16961), .B(n38568), .Z(n16963) );
  XNOR U41214 ( .A(q[13]), .B(DB[3013]), .Z(n38568) );
  XNOR U41215 ( .A(q[12]), .B(DB[3012]), .Z(n16961) );
  IV U41216 ( .A(n16974), .Z(n38566) );
  XOR U41217 ( .A(n38569), .B(n38570), .Z(n16974) );
  XNOR U41218 ( .A(n16970), .B(n16972), .Z(n38570) );
  XNOR U41219 ( .A(q[8]), .B(DB[3008]), .Z(n16972) );
  XNOR U41220 ( .A(q[11]), .B(DB[3011]), .Z(n16970) );
  IV U41221 ( .A(n16969), .Z(n38569) );
  XNOR U41222 ( .A(n16967), .B(n38571), .Z(n16969) );
  XNOR U41223 ( .A(q[10]), .B(DB[3010]), .Z(n38571) );
  XNOR U41224 ( .A(q[9]), .B(DB[3009]), .Z(n16967) );
  IV U41225 ( .A(n16982), .Z(n38565) );
  XOR U41226 ( .A(n38572), .B(n38573), .Z(n16982) );
  XNOR U41227 ( .A(n16999), .B(n16980), .Z(n38573) );
  XNOR U41228 ( .A(q[0]), .B(DB[3000]), .Z(n16980) );
  XOR U41229 ( .A(n38574), .B(n16988), .Z(n16999) );
  XNOR U41230 ( .A(q[7]), .B(DB[3007]), .Z(n16988) );
  IV U41231 ( .A(n16987), .Z(n38574) );
  XNOR U41232 ( .A(n16985), .B(n38575), .Z(n16987) );
  XNOR U41233 ( .A(q[6]), .B(DB[3006]), .Z(n38575) );
  XNOR U41234 ( .A(q[5]), .B(DB[3005]), .Z(n16985) );
  IV U41235 ( .A(n16998), .Z(n38572) );
  XOR U41236 ( .A(n38576), .B(n38577), .Z(n16998) );
  XNOR U41237 ( .A(n16994), .B(n16996), .Z(n38577) );
  XNOR U41238 ( .A(q[1]), .B(DB[3001]), .Z(n16996) );
  XNOR U41239 ( .A(q[4]), .B(DB[3004]), .Z(n16994) );
  IV U41240 ( .A(n16993), .Z(n38576) );
  XNOR U41241 ( .A(n16991), .B(n38578), .Z(n16993) );
  XNOR U41242 ( .A(q[3]), .B(DB[3003]), .Z(n38578) );
  XNOR U41243 ( .A(q[2]), .B(DB[3002]), .Z(n16991) );
  XOR U41244 ( .A(n38579), .B(n16889), .Z(n16817) );
  XOR U41245 ( .A(n38580), .B(n16881), .Z(n16889) );
  XOR U41246 ( .A(n38581), .B(n16870), .Z(n16881) );
  XNOR U41247 ( .A(q[14]), .B(DB[3029]), .Z(n16870) );
  IV U41248 ( .A(n16869), .Z(n38581) );
  XNOR U41249 ( .A(n16867), .B(n38582), .Z(n16869) );
  XNOR U41250 ( .A(q[13]), .B(DB[3028]), .Z(n38582) );
  XNOR U41251 ( .A(q[12]), .B(DB[3027]), .Z(n16867) );
  IV U41252 ( .A(n16880), .Z(n38580) );
  XOR U41253 ( .A(n38583), .B(n38584), .Z(n16880) );
  XNOR U41254 ( .A(n16876), .B(n16878), .Z(n38584) );
  XNOR U41255 ( .A(q[8]), .B(DB[3023]), .Z(n16878) );
  XNOR U41256 ( .A(q[11]), .B(DB[3026]), .Z(n16876) );
  IV U41257 ( .A(n16875), .Z(n38583) );
  XNOR U41258 ( .A(n16873), .B(n38585), .Z(n16875) );
  XNOR U41259 ( .A(q[10]), .B(DB[3025]), .Z(n38585) );
  XNOR U41260 ( .A(q[9]), .B(DB[3024]), .Z(n16873) );
  IV U41261 ( .A(n16888), .Z(n38579) );
  XOR U41262 ( .A(n38586), .B(n38587), .Z(n16888) );
  XNOR U41263 ( .A(n16905), .B(n16886), .Z(n38587) );
  XNOR U41264 ( .A(q[0]), .B(DB[3015]), .Z(n16886) );
  XOR U41265 ( .A(n38588), .B(n16894), .Z(n16905) );
  XNOR U41266 ( .A(q[7]), .B(DB[3022]), .Z(n16894) );
  IV U41267 ( .A(n16893), .Z(n38588) );
  XNOR U41268 ( .A(n16891), .B(n38589), .Z(n16893) );
  XNOR U41269 ( .A(q[6]), .B(DB[3021]), .Z(n38589) );
  XNOR U41270 ( .A(q[5]), .B(DB[3020]), .Z(n16891) );
  IV U41271 ( .A(n16904), .Z(n38586) );
  XOR U41272 ( .A(n38590), .B(n38591), .Z(n16904) );
  XNOR U41273 ( .A(n16900), .B(n16902), .Z(n38591) );
  XNOR U41274 ( .A(q[1]), .B(DB[3016]), .Z(n16902) );
  XNOR U41275 ( .A(q[4]), .B(DB[3019]), .Z(n16900) );
  IV U41276 ( .A(n16899), .Z(n38590) );
  XNOR U41277 ( .A(n16897), .B(n38592), .Z(n16899) );
  XNOR U41278 ( .A(q[3]), .B(DB[3018]), .Z(n38592) );
  XNOR U41279 ( .A(q[2]), .B(DB[3017]), .Z(n16897) );
  XOR U41280 ( .A(n38593), .B(n16795), .Z(n16723) );
  XOR U41281 ( .A(n38594), .B(n16787), .Z(n16795) );
  XOR U41282 ( .A(n38595), .B(n16776), .Z(n16787) );
  XNOR U41283 ( .A(q[14]), .B(DB[3044]), .Z(n16776) );
  IV U41284 ( .A(n16775), .Z(n38595) );
  XNOR U41285 ( .A(n16773), .B(n38596), .Z(n16775) );
  XNOR U41286 ( .A(q[13]), .B(DB[3043]), .Z(n38596) );
  XNOR U41287 ( .A(q[12]), .B(DB[3042]), .Z(n16773) );
  IV U41288 ( .A(n16786), .Z(n38594) );
  XOR U41289 ( .A(n38597), .B(n38598), .Z(n16786) );
  XNOR U41290 ( .A(n16782), .B(n16784), .Z(n38598) );
  XNOR U41291 ( .A(q[8]), .B(DB[3038]), .Z(n16784) );
  XNOR U41292 ( .A(q[11]), .B(DB[3041]), .Z(n16782) );
  IV U41293 ( .A(n16781), .Z(n38597) );
  XNOR U41294 ( .A(n16779), .B(n38599), .Z(n16781) );
  XNOR U41295 ( .A(q[10]), .B(DB[3040]), .Z(n38599) );
  XNOR U41296 ( .A(q[9]), .B(DB[3039]), .Z(n16779) );
  IV U41297 ( .A(n16794), .Z(n38593) );
  XOR U41298 ( .A(n38600), .B(n38601), .Z(n16794) );
  XNOR U41299 ( .A(n16811), .B(n16792), .Z(n38601) );
  XNOR U41300 ( .A(q[0]), .B(DB[3030]), .Z(n16792) );
  XOR U41301 ( .A(n38602), .B(n16800), .Z(n16811) );
  XNOR U41302 ( .A(q[7]), .B(DB[3037]), .Z(n16800) );
  IV U41303 ( .A(n16799), .Z(n38602) );
  XNOR U41304 ( .A(n16797), .B(n38603), .Z(n16799) );
  XNOR U41305 ( .A(q[6]), .B(DB[3036]), .Z(n38603) );
  XNOR U41306 ( .A(q[5]), .B(DB[3035]), .Z(n16797) );
  IV U41307 ( .A(n16810), .Z(n38600) );
  XOR U41308 ( .A(n38604), .B(n38605), .Z(n16810) );
  XNOR U41309 ( .A(n16806), .B(n16808), .Z(n38605) );
  XNOR U41310 ( .A(q[1]), .B(DB[3031]), .Z(n16808) );
  XNOR U41311 ( .A(q[4]), .B(DB[3034]), .Z(n16806) );
  IV U41312 ( .A(n16805), .Z(n38604) );
  XNOR U41313 ( .A(n16803), .B(n38606), .Z(n16805) );
  XNOR U41314 ( .A(q[3]), .B(DB[3033]), .Z(n38606) );
  XNOR U41315 ( .A(q[2]), .B(DB[3032]), .Z(n16803) );
  XOR U41316 ( .A(n38607), .B(n16701), .Z(n16629) );
  XOR U41317 ( .A(n38608), .B(n16693), .Z(n16701) );
  XOR U41318 ( .A(n38609), .B(n16682), .Z(n16693) );
  XNOR U41319 ( .A(q[14]), .B(DB[3059]), .Z(n16682) );
  IV U41320 ( .A(n16681), .Z(n38609) );
  XNOR U41321 ( .A(n16679), .B(n38610), .Z(n16681) );
  XNOR U41322 ( .A(q[13]), .B(DB[3058]), .Z(n38610) );
  XNOR U41323 ( .A(q[12]), .B(DB[3057]), .Z(n16679) );
  IV U41324 ( .A(n16692), .Z(n38608) );
  XOR U41325 ( .A(n38611), .B(n38612), .Z(n16692) );
  XNOR U41326 ( .A(n16688), .B(n16690), .Z(n38612) );
  XNOR U41327 ( .A(q[8]), .B(DB[3053]), .Z(n16690) );
  XNOR U41328 ( .A(q[11]), .B(DB[3056]), .Z(n16688) );
  IV U41329 ( .A(n16687), .Z(n38611) );
  XNOR U41330 ( .A(n16685), .B(n38613), .Z(n16687) );
  XNOR U41331 ( .A(q[10]), .B(DB[3055]), .Z(n38613) );
  XNOR U41332 ( .A(q[9]), .B(DB[3054]), .Z(n16685) );
  IV U41333 ( .A(n16700), .Z(n38607) );
  XOR U41334 ( .A(n38614), .B(n38615), .Z(n16700) );
  XNOR U41335 ( .A(n16717), .B(n16698), .Z(n38615) );
  XNOR U41336 ( .A(q[0]), .B(DB[3045]), .Z(n16698) );
  XOR U41337 ( .A(n38616), .B(n16706), .Z(n16717) );
  XNOR U41338 ( .A(q[7]), .B(DB[3052]), .Z(n16706) );
  IV U41339 ( .A(n16705), .Z(n38616) );
  XNOR U41340 ( .A(n16703), .B(n38617), .Z(n16705) );
  XNOR U41341 ( .A(q[6]), .B(DB[3051]), .Z(n38617) );
  XNOR U41342 ( .A(q[5]), .B(DB[3050]), .Z(n16703) );
  IV U41343 ( .A(n16716), .Z(n38614) );
  XOR U41344 ( .A(n38618), .B(n38619), .Z(n16716) );
  XNOR U41345 ( .A(n16712), .B(n16714), .Z(n38619) );
  XNOR U41346 ( .A(q[1]), .B(DB[3046]), .Z(n16714) );
  XNOR U41347 ( .A(q[4]), .B(DB[3049]), .Z(n16712) );
  IV U41348 ( .A(n16711), .Z(n38618) );
  XNOR U41349 ( .A(n16709), .B(n38620), .Z(n16711) );
  XNOR U41350 ( .A(q[3]), .B(DB[3048]), .Z(n38620) );
  XNOR U41351 ( .A(q[2]), .B(DB[3047]), .Z(n16709) );
  XOR U41352 ( .A(n38621), .B(n16607), .Z(n16535) );
  XOR U41353 ( .A(n38622), .B(n16599), .Z(n16607) );
  XOR U41354 ( .A(n38623), .B(n16588), .Z(n16599) );
  XNOR U41355 ( .A(q[14]), .B(DB[3074]), .Z(n16588) );
  IV U41356 ( .A(n16587), .Z(n38623) );
  XNOR U41357 ( .A(n16585), .B(n38624), .Z(n16587) );
  XNOR U41358 ( .A(q[13]), .B(DB[3073]), .Z(n38624) );
  XNOR U41359 ( .A(q[12]), .B(DB[3072]), .Z(n16585) );
  IV U41360 ( .A(n16598), .Z(n38622) );
  XOR U41361 ( .A(n38625), .B(n38626), .Z(n16598) );
  XNOR U41362 ( .A(n16594), .B(n16596), .Z(n38626) );
  XNOR U41363 ( .A(q[8]), .B(DB[3068]), .Z(n16596) );
  XNOR U41364 ( .A(q[11]), .B(DB[3071]), .Z(n16594) );
  IV U41365 ( .A(n16593), .Z(n38625) );
  XNOR U41366 ( .A(n16591), .B(n38627), .Z(n16593) );
  XNOR U41367 ( .A(q[10]), .B(DB[3070]), .Z(n38627) );
  XNOR U41368 ( .A(q[9]), .B(DB[3069]), .Z(n16591) );
  IV U41369 ( .A(n16606), .Z(n38621) );
  XOR U41370 ( .A(n38628), .B(n38629), .Z(n16606) );
  XNOR U41371 ( .A(n16623), .B(n16604), .Z(n38629) );
  XNOR U41372 ( .A(q[0]), .B(DB[3060]), .Z(n16604) );
  XOR U41373 ( .A(n38630), .B(n16612), .Z(n16623) );
  XNOR U41374 ( .A(q[7]), .B(DB[3067]), .Z(n16612) );
  IV U41375 ( .A(n16611), .Z(n38630) );
  XNOR U41376 ( .A(n16609), .B(n38631), .Z(n16611) );
  XNOR U41377 ( .A(q[6]), .B(DB[3066]), .Z(n38631) );
  XNOR U41378 ( .A(q[5]), .B(DB[3065]), .Z(n16609) );
  IV U41379 ( .A(n16622), .Z(n38628) );
  XOR U41380 ( .A(n38632), .B(n38633), .Z(n16622) );
  XNOR U41381 ( .A(n16618), .B(n16620), .Z(n38633) );
  XNOR U41382 ( .A(q[1]), .B(DB[3061]), .Z(n16620) );
  XNOR U41383 ( .A(q[4]), .B(DB[3064]), .Z(n16618) );
  IV U41384 ( .A(n16617), .Z(n38632) );
  XNOR U41385 ( .A(n16615), .B(n38634), .Z(n16617) );
  XNOR U41386 ( .A(q[3]), .B(DB[3063]), .Z(n38634) );
  XNOR U41387 ( .A(q[2]), .B(DB[3062]), .Z(n16615) );
  XOR U41388 ( .A(n38635), .B(n16513), .Z(n16441) );
  XOR U41389 ( .A(n38636), .B(n16505), .Z(n16513) );
  XOR U41390 ( .A(n38637), .B(n16494), .Z(n16505) );
  XNOR U41391 ( .A(q[14]), .B(DB[3089]), .Z(n16494) );
  IV U41392 ( .A(n16493), .Z(n38637) );
  XNOR U41393 ( .A(n16491), .B(n38638), .Z(n16493) );
  XNOR U41394 ( .A(q[13]), .B(DB[3088]), .Z(n38638) );
  XNOR U41395 ( .A(q[12]), .B(DB[3087]), .Z(n16491) );
  IV U41396 ( .A(n16504), .Z(n38636) );
  XOR U41397 ( .A(n38639), .B(n38640), .Z(n16504) );
  XNOR U41398 ( .A(n16500), .B(n16502), .Z(n38640) );
  XNOR U41399 ( .A(q[8]), .B(DB[3083]), .Z(n16502) );
  XNOR U41400 ( .A(q[11]), .B(DB[3086]), .Z(n16500) );
  IV U41401 ( .A(n16499), .Z(n38639) );
  XNOR U41402 ( .A(n16497), .B(n38641), .Z(n16499) );
  XNOR U41403 ( .A(q[10]), .B(DB[3085]), .Z(n38641) );
  XNOR U41404 ( .A(q[9]), .B(DB[3084]), .Z(n16497) );
  IV U41405 ( .A(n16512), .Z(n38635) );
  XOR U41406 ( .A(n38642), .B(n38643), .Z(n16512) );
  XNOR U41407 ( .A(n16529), .B(n16510), .Z(n38643) );
  XNOR U41408 ( .A(q[0]), .B(DB[3075]), .Z(n16510) );
  XOR U41409 ( .A(n38644), .B(n16518), .Z(n16529) );
  XNOR U41410 ( .A(q[7]), .B(DB[3082]), .Z(n16518) );
  IV U41411 ( .A(n16517), .Z(n38644) );
  XNOR U41412 ( .A(n16515), .B(n38645), .Z(n16517) );
  XNOR U41413 ( .A(q[6]), .B(DB[3081]), .Z(n38645) );
  XNOR U41414 ( .A(q[5]), .B(DB[3080]), .Z(n16515) );
  IV U41415 ( .A(n16528), .Z(n38642) );
  XOR U41416 ( .A(n38646), .B(n38647), .Z(n16528) );
  XNOR U41417 ( .A(n16524), .B(n16526), .Z(n38647) );
  XNOR U41418 ( .A(q[1]), .B(DB[3076]), .Z(n16526) );
  XNOR U41419 ( .A(q[4]), .B(DB[3079]), .Z(n16524) );
  IV U41420 ( .A(n16523), .Z(n38646) );
  XNOR U41421 ( .A(n16521), .B(n38648), .Z(n16523) );
  XNOR U41422 ( .A(q[3]), .B(DB[3078]), .Z(n38648) );
  XNOR U41423 ( .A(q[2]), .B(DB[3077]), .Z(n16521) );
  XOR U41424 ( .A(n38649), .B(n16419), .Z(n16347) );
  XOR U41425 ( .A(n38650), .B(n16411), .Z(n16419) );
  XOR U41426 ( .A(n38651), .B(n16400), .Z(n16411) );
  XNOR U41427 ( .A(q[14]), .B(DB[3104]), .Z(n16400) );
  IV U41428 ( .A(n16399), .Z(n38651) );
  XNOR U41429 ( .A(n16397), .B(n38652), .Z(n16399) );
  XNOR U41430 ( .A(q[13]), .B(DB[3103]), .Z(n38652) );
  XNOR U41431 ( .A(q[12]), .B(DB[3102]), .Z(n16397) );
  IV U41432 ( .A(n16410), .Z(n38650) );
  XOR U41433 ( .A(n38653), .B(n38654), .Z(n16410) );
  XNOR U41434 ( .A(n16406), .B(n16408), .Z(n38654) );
  XNOR U41435 ( .A(q[8]), .B(DB[3098]), .Z(n16408) );
  XNOR U41436 ( .A(q[11]), .B(DB[3101]), .Z(n16406) );
  IV U41437 ( .A(n16405), .Z(n38653) );
  XNOR U41438 ( .A(n16403), .B(n38655), .Z(n16405) );
  XNOR U41439 ( .A(q[10]), .B(DB[3100]), .Z(n38655) );
  XNOR U41440 ( .A(q[9]), .B(DB[3099]), .Z(n16403) );
  IV U41441 ( .A(n16418), .Z(n38649) );
  XOR U41442 ( .A(n38656), .B(n38657), .Z(n16418) );
  XNOR U41443 ( .A(n16435), .B(n16416), .Z(n38657) );
  XNOR U41444 ( .A(q[0]), .B(DB[3090]), .Z(n16416) );
  XOR U41445 ( .A(n38658), .B(n16424), .Z(n16435) );
  XNOR U41446 ( .A(q[7]), .B(DB[3097]), .Z(n16424) );
  IV U41447 ( .A(n16423), .Z(n38658) );
  XNOR U41448 ( .A(n16421), .B(n38659), .Z(n16423) );
  XNOR U41449 ( .A(q[6]), .B(DB[3096]), .Z(n38659) );
  XNOR U41450 ( .A(q[5]), .B(DB[3095]), .Z(n16421) );
  IV U41451 ( .A(n16434), .Z(n38656) );
  XOR U41452 ( .A(n38660), .B(n38661), .Z(n16434) );
  XNOR U41453 ( .A(n16430), .B(n16432), .Z(n38661) );
  XNOR U41454 ( .A(q[1]), .B(DB[3091]), .Z(n16432) );
  XNOR U41455 ( .A(q[4]), .B(DB[3094]), .Z(n16430) );
  IV U41456 ( .A(n16429), .Z(n38660) );
  XNOR U41457 ( .A(n16427), .B(n38662), .Z(n16429) );
  XNOR U41458 ( .A(q[3]), .B(DB[3093]), .Z(n38662) );
  XNOR U41459 ( .A(q[2]), .B(DB[3092]), .Z(n16427) );
  XOR U41460 ( .A(n38663), .B(n16325), .Z(n16253) );
  XOR U41461 ( .A(n38664), .B(n16317), .Z(n16325) );
  XOR U41462 ( .A(n38665), .B(n16306), .Z(n16317) );
  XNOR U41463 ( .A(q[14]), .B(DB[3119]), .Z(n16306) );
  IV U41464 ( .A(n16305), .Z(n38665) );
  XNOR U41465 ( .A(n16303), .B(n38666), .Z(n16305) );
  XNOR U41466 ( .A(q[13]), .B(DB[3118]), .Z(n38666) );
  XNOR U41467 ( .A(q[12]), .B(DB[3117]), .Z(n16303) );
  IV U41468 ( .A(n16316), .Z(n38664) );
  XOR U41469 ( .A(n38667), .B(n38668), .Z(n16316) );
  XNOR U41470 ( .A(n16312), .B(n16314), .Z(n38668) );
  XNOR U41471 ( .A(q[8]), .B(DB[3113]), .Z(n16314) );
  XNOR U41472 ( .A(q[11]), .B(DB[3116]), .Z(n16312) );
  IV U41473 ( .A(n16311), .Z(n38667) );
  XNOR U41474 ( .A(n16309), .B(n38669), .Z(n16311) );
  XNOR U41475 ( .A(q[10]), .B(DB[3115]), .Z(n38669) );
  XNOR U41476 ( .A(q[9]), .B(DB[3114]), .Z(n16309) );
  IV U41477 ( .A(n16324), .Z(n38663) );
  XOR U41478 ( .A(n38670), .B(n38671), .Z(n16324) );
  XNOR U41479 ( .A(n16341), .B(n16322), .Z(n38671) );
  XNOR U41480 ( .A(q[0]), .B(DB[3105]), .Z(n16322) );
  XOR U41481 ( .A(n38672), .B(n16330), .Z(n16341) );
  XNOR U41482 ( .A(q[7]), .B(DB[3112]), .Z(n16330) );
  IV U41483 ( .A(n16329), .Z(n38672) );
  XNOR U41484 ( .A(n16327), .B(n38673), .Z(n16329) );
  XNOR U41485 ( .A(q[6]), .B(DB[3111]), .Z(n38673) );
  XNOR U41486 ( .A(q[5]), .B(DB[3110]), .Z(n16327) );
  IV U41487 ( .A(n16340), .Z(n38670) );
  XOR U41488 ( .A(n38674), .B(n38675), .Z(n16340) );
  XNOR U41489 ( .A(n16336), .B(n16338), .Z(n38675) );
  XNOR U41490 ( .A(q[1]), .B(DB[3106]), .Z(n16338) );
  XNOR U41491 ( .A(q[4]), .B(DB[3109]), .Z(n16336) );
  IV U41492 ( .A(n16335), .Z(n38674) );
  XNOR U41493 ( .A(n16333), .B(n38676), .Z(n16335) );
  XNOR U41494 ( .A(q[3]), .B(DB[3108]), .Z(n38676) );
  XNOR U41495 ( .A(q[2]), .B(DB[3107]), .Z(n16333) );
  XOR U41496 ( .A(n38677), .B(n16231), .Z(n16159) );
  XOR U41497 ( .A(n38678), .B(n16223), .Z(n16231) );
  XOR U41498 ( .A(n38679), .B(n16212), .Z(n16223) );
  XNOR U41499 ( .A(q[14]), .B(DB[3134]), .Z(n16212) );
  IV U41500 ( .A(n16211), .Z(n38679) );
  XNOR U41501 ( .A(n16209), .B(n38680), .Z(n16211) );
  XNOR U41502 ( .A(q[13]), .B(DB[3133]), .Z(n38680) );
  XNOR U41503 ( .A(q[12]), .B(DB[3132]), .Z(n16209) );
  IV U41504 ( .A(n16222), .Z(n38678) );
  XOR U41505 ( .A(n38681), .B(n38682), .Z(n16222) );
  XNOR U41506 ( .A(n16218), .B(n16220), .Z(n38682) );
  XNOR U41507 ( .A(q[8]), .B(DB[3128]), .Z(n16220) );
  XNOR U41508 ( .A(q[11]), .B(DB[3131]), .Z(n16218) );
  IV U41509 ( .A(n16217), .Z(n38681) );
  XNOR U41510 ( .A(n16215), .B(n38683), .Z(n16217) );
  XNOR U41511 ( .A(q[10]), .B(DB[3130]), .Z(n38683) );
  XNOR U41512 ( .A(q[9]), .B(DB[3129]), .Z(n16215) );
  IV U41513 ( .A(n16230), .Z(n38677) );
  XOR U41514 ( .A(n38684), .B(n38685), .Z(n16230) );
  XNOR U41515 ( .A(n16247), .B(n16228), .Z(n38685) );
  XNOR U41516 ( .A(q[0]), .B(DB[3120]), .Z(n16228) );
  XOR U41517 ( .A(n38686), .B(n16236), .Z(n16247) );
  XNOR U41518 ( .A(q[7]), .B(DB[3127]), .Z(n16236) );
  IV U41519 ( .A(n16235), .Z(n38686) );
  XNOR U41520 ( .A(n16233), .B(n38687), .Z(n16235) );
  XNOR U41521 ( .A(q[6]), .B(DB[3126]), .Z(n38687) );
  XNOR U41522 ( .A(q[5]), .B(DB[3125]), .Z(n16233) );
  IV U41523 ( .A(n16246), .Z(n38684) );
  XOR U41524 ( .A(n38688), .B(n38689), .Z(n16246) );
  XNOR U41525 ( .A(n16242), .B(n16244), .Z(n38689) );
  XNOR U41526 ( .A(q[1]), .B(DB[3121]), .Z(n16244) );
  XNOR U41527 ( .A(q[4]), .B(DB[3124]), .Z(n16242) );
  IV U41528 ( .A(n16241), .Z(n38688) );
  XNOR U41529 ( .A(n16239), .B(n38690), .Z(n16241) );
  XNOR U41530 ( .A(q[3]), .B(DB[3123]), .Z(n38690) );
  XNOR U41531 ( .A(q[2]), .B(DB[3122]), .Z(n16239) );
  XOR U41532 ( .A(n38691), .B(n16137), .Z(n16065) );
  XOR U41533 ( .A(n38692), .B(n16129), .Z(n16137) );
  XOR U41534 ( .A(n38693), .B(n16118), .Z(n16129) );
  XNOR U41535 ( .A(q[14]), .B(DB[3149]), .Z(n16118) );
  IV U41536 ( .A(n16117), .Z(n38693) );
  XNOR U41537 ( .A(n16115), .B(n38694), .Z(n16117) );
  XNOR U41538 ( .A(q[13]), .B(DB[3148]), .Z(n38694) );
  XNOR U41539 ( .A(q[12]), .B(DB[3147]), .Z(n16115) );
  IV U41540 ( .A(n16128), .Z(n38692) );
  XOR U41541 ( .A(n38695), .B(n38696), .Z(n16128) );
  XNOR U41542 ( .A(n16124), .B(n16126), .Z(n38696) );
  XNOR U41543 ( .A(q[8]), .B(DB[3143]), .Z(n16126) );
  XNOR U41544 ( .A(q[11]), .B(DB[3146]), .Z(n16124) );
  IV U41545 ( .A(n16123), .Z(n38695) );
  XNOR U41546 ( .A(n16121), .B(n38697), .Z(n16123) );
  XNOR U41547 ( .A(q[10]), .B(DB[3145]), .Z(n38697) );
  XNOR U41548 ( .A(q[9]), .B(DB[3144]), .Z(n16121) );
  IV U41549 ( .A(n16136), .Z(n38691) );
  XOR U41550 ( .A(n38698), .B(n38699), .Z(n16136) );
  XNOR U41551 ( .A(n16153), .B(n16134), .Z(n38699) );
  XNOR U41552 ( .A(q[0]), .B(DB[3135]), .Z(n16134) );
  XOR U41553 ( .A(n38700), .B(n16142), .Z(n16153) );
  XNOR U41554 ( .A(q[7]), .B(DB[3142]), .Z(n16142) );
  IV U41555 ( .A(n16141), .Z(n38700) );
  XNOR U41556 ( .A(n16139), .B(n38701), .Z(n16141) );
  XNOR U41557 ( .A(q[6]), .B(DB[3141]), .Z(n38701) );
  XNOR U41558 ( .A(q[5]), .B(DB[3140]), .Z(n16139) );
  IV U41559 ( .A(n16152), .Z(n38698) );
  XOR U41560 ( .A(n38702), .B(n38703), .Z(n16152) );
  XNOR U41561 ( .A(n16148), .B(n16150), .Z(n38703) );
  XNOR U41562 ( .A(q[1]), .B(DB[3136]), .Z(n16150) );
  XNOR U41563 ( .A(q[4]), .B(DB[3139]), .Z(n16148) );
  IV U41564 ( .A(n16147), .Z(n38702) );
  XNOR U41565 ( .A(n16145), .B(n38704), .Z(n16147) );
  XNOR U41566 ( .A(q[3]), .B(DB[3138]), .Z(n38704) );
  XNOR U41567 ( .A(q[2]), .B(DB[3137]), .Z(n16145) );
  XOR U41568 ( .A(n38705), .B(n16043), .Z(n15971) );
  XOR U41569 ( .A(n38706), .B(n16035), .Z(n16043) );
  XOR U41570 ( .A(n38707), .B(n16024), .Z(n16035) );
  XNOR U41571 ( .A(q[14]), .B(DB[3164]), .Z(n16024) );
  IV U41572 ( .A(n16023), .Z(n38707) );
  XNOR U41573 ( .A(n16021), .B(n38708), .Z(n16023) );
  XNOR U41574 ( .A(q[13]), .B(DB[3163]), .Z(n38708) );
  XNOR U41575 ( .A(q[12]), .B(DB[3162]), .Z(n16021) );
  IV U41576 ( .A(n16034), .Z(n38706) );
  XOR U41577 ( .A(n38709), .B(n38710), .Z(n16034) );
  XNOR U41578 ( .A(n16030), .B(n16032), .Z(n38710) );
  XNOR U41579 ( .A(q[8]), .B(DB[3158]), .Z(n16032) );
  XNOR U41580 ( .A(q[11]), .B(DB[3161]), .Z(n16030) );
  IV U41581 ( .A(n16029), .Z(n38709) );
  XNOR U41582 ( .A(n16027), .B(n38711), .Z(n16029) );
  XNOR U41583 ( .A(q[10]), .B(DB[3160]), .Z(n38711) );
  XNOR U41584 ( .A(q[9]), .B(DB[3159]), .Z(n16027) );
  IV U41585 ( .A(n16042), .Z(n38705) );
  XOR U41586 ( .A(n38712), .B(n38713), .Z(n16042) );
  XNOR U41587 ( .A(n16059), .B(n16040), .Z(n38713) );
  XNOR U41588 ( .A(q[0]), .B(DB[3150]), .Z(n16040) );
  XOR U41589 ( .A(n38714), .B(n16048), .Z(n16059) );
  XNOR U41590 ( .A(q[7]), .B(DB[3157]), .Z(n16048) );
  IV U41591 ( .A(n16047), .Z(n38714) );
  XNOR U41592 ( .A(n16045), .B(n38715), .Z(n16047) );
  XNOR U41593 ( .A(q[6]), .B(DB[3156]), .Z(n38715) );
  XNOR U41594 ( .A(q[5]), .B(DB[3155]), .Z(n16045) );
  IV U41595 ( .A(n16058), .Z(n38712) );
  XOR U41596 ( .A(n38716), .B(n38717), .Z(n16058) );
  XNOR U41597 ( .A(n16054), .B(n16056), .Z(n38717) );
  XNOR U41598 ( .A(q[1]), .B(DB[3151]), .Z(n16056) );
  XNOR U41599 ( .A(q[4]), .B(DB[3154]), .Z(n16054) );
  IV U41600 ( .A(n16053), .Z(n38716) );
  XNOR U41601 ( .A(n16051), .B(n38718), .Z(n16053) );
  XNOR U41602 ( .A(q[3]), .B(DB[3153]), .Z(n38718) );
  XNOR U41603 ( .A(q[2]), .B(DB[3152]), .Z(n16051) );
  XOR U41604 ( .A(n38719), .B(n15949), .Z(n15877) );
  XOR U41605 ( .A(n38720), .B(n15941), .Z(n15949) );
  XOR U41606 ( .A(n38721), .B(n15930), .Z(n15941) );
  XNOR U41607 ( .A(q[14]), .B(DB[3179]), .Z(n15930) );
  IV U41608 ( .A(n15929), .Z(n38721) );
  XNOR U41609 ( .A(n15927), .B(n38722), .Z(n15929) );
  XNOR U41610 ( .A(q[13]), .B(DB[3178]), .Z(n38722) );
  XNOR U41611 ( .A(q[12]), .B(DB[3177]), .Z(n15927) );
  IV U41612 ( .A(n15940), .Z(n38720) );
  XOR U41613 ( .A(n38723), .B(n38724), .Z(n15940) );
  XNOR U41614 ( .A(n15936), .B(n15938), .Z(n38724) );
  XNOR U41615 ( .A(q[8]), .B(DB[3173]), .Z(n15938) );
  XNOR U41616 ( .A(q[11]), .B(DB[3176]), .Z(n15936) );
  IV U41617 ( .A(n15935), .Z(n38723) );
  XNOR U41618 ( .A(n15933), .B(n38725), .Z(n15935) );
  XNOR U41619 ( .A(q[10]), .B(DB[3175]), .Z(n38725) );
  XNOR U41620 ( .A(q[9]), .B(DB[3174]), .Z(n15933) );
  IV U41621 ( .A(n15948), .Z(n38719) );
  XOR U41622 ( .A(n38726), .B(n38727), .Z(n15948) );
  XNOR U41623 ( .A(n15965), .B(n15946), .Z(n38727) );
  XNOR U41624 ( .A(q[0]), .B(DB[3165]), .Z(n15946) );
  XOR U41625 ( .A(n38728), .B(n15954), .Z(n15965) );
  XNOR U41626 ( .A(q[7]), .B(DB[3172]), .Z(n15954) );
  IV U41627 ( .A(n15953), .Z(n38728) );
  XNOR U41628 ( .A(n15951), .B(n38729), .Z(n15953) );
  XNOR U41629 ( .A(q[6]), .B(DB[3171]), .Z(n38729) );
  XNOR U41630 ( .A(q[5]), .B(DB[3170]), .Z(n15951) );
  IV U41631 ( .A(n15964), .Z(n38726) );
  XOR U41632 ( .A(n38730), .B(n38731), .Z(n15964) );
  XNOR U41633 ( .A(n15960), .B(n15962), .Z(n38731) );
  XNOR U41634 ( .A(q[1]), .B(DB[3166]), .Z(n15962) );
  XNOR U41635 ( .A(q[4]), .B(DB[3169]), .Z(n15960) );
  IV U41636 ( .A(n15959), .Z(n38730) );
  XNOR U41637 ( .A(n15957), .B(n38732), .Z(n15959) );
  XNOR U41638 ( .A(q[3]), .B(DB[3168]), .Z(n38732) );
  XNOR U41639 ( .A(q[2]), .B(DB[3167]), .Z(n15957) );
  XOR U41640 ( .A(n38733), .B(n15855), .Z(n15783) );
  XOR U41641 ( .A(n38734), .B(n15847), .Z(n15855) );
  XOR U41642 ( .A(n38735), .B(n15836), .Z(n15847) );
  XNOR U41643 ( .A(q[14]), .B(DB[3194]), .Z(n15836) );
  IV U41644 ( .A(n15835), .Z(n38735) );
  XNOR U41645 ( .A(n15833), .B(n38736), .Z(n15835) );
  XNOR U41646 ( .A(q[13]), .B(DB[3193]), .Z(n38736) );
  XNOR U41647 ( .A(q[12]), .B(DB[3192]), .Z(n15833) );
  IV U41648 ( .A(n15846), .Z(n38734) );
  XOR U41649 ( .A(n38737), .B(n38738), .Z(n15846) );
  XNOR U41650 ( .A(n15842), .B(n15844), .Z(n38738) );
  XNOR U41651 ( .A(q[8]), .B(DB[3188]), .Z(n15844) );
  XNOR U41652 ( .A(q[11]), .B(DB[3191]), .Z(n15842) );
  IV U41653 ( .A(n15841), .Z(n38737) );
  XNOR U41654 ( .A(n15839), .B(n38739), .Z(n15841) );
  XNOR U41655 ( .A(q[10]), .B(DB[3190]), .Z(n38739) );
  XNOR U41656 ( .A(q[9]), .B(DB[3189]), .Z(n15839) );
  IV U41657 ( .A(n15854), .Z(n38733) );
  XOR U41658 ( .A(n38740), .B(n38741), .Z(n15854) );
  XNOR U41659 ( .A(n15871), .B(n15852), .Z(n38741) );
  XNOR U41660 ( .A(q[0]), .B(DB[3180]), .Z(n15852) );
  XOR U41661 ( .A(n38742), .B(n15860), .Z(n15871) );
  XNOR U41662 ( .A(q[7]), .B(DB[3187]), .Z(n15860) );
  IV U41663 ( .A(n15859), .Z(n38742) );
  XNOR U41664 ( .A(n15857), .B(n38743), .Z(n15859) );
  XNOR U41665 ( .A(q[6]), .B(DB[3186]), .Z(n38743) );
  XNOR U41666 ( .A(q[5]), .B(DB[3185]), .Z(n15857) );
  IV U41667 ( .A(n15870), .Z(n38740) );
  XOR U41668 ( .A(n38744), .B(n38745), .Z(n15870) );
  XNOR U41669 ( .A(n15866), .B(n15868), .Z(n38745) );
  XNOR U41670 ( .A(q[1]), .B(DB[3181]), .Z(n15868) );
  XNOR U41671 ( .A(q[4]), .B(DB[3184]), .Z(n15866) );
  IV U41672 ( .A(n15865), .Z(n38744) );
  XNOR U41673 ( .A(n15863), .B(n38746), .Z(n15865) );
  XNOR U41674 ( .A(q[3]), .B(DB[3183]), .Z(n38746) );
  XNOR U41675 ( .A(q[2]), .B(DB[3182]), .Z(n15863) );
  XOR U41676 ( .A(n38747), .B(n15761), .Z(n15689) );
  XOR U41677 ( .A(n38748), .B(n15753), .Z(n15761) );
  XOR U41678 ( .A(n38749), .B(n15742), .Z(n15753) );
  XNOR U41679 ( .A(q[14]), .B(DB[3209]), .Z(n15742) );
  IV U41680 ( .A(n15741), .Z(n38749) );
  XNOR U41681 ( .A(n15739), .B(n38750), .Z(n15741) );
  XNOR U41682 ( .A(q[13]), .B(DB[3208]), .Z(n38750) );
  XNOR U41683 ( .A(q[12]), .B(DB[3207]), .Z(n15739) );
  IV U41684 ( .A(n15752), .Z(n38748) );
  XOR U41685 ( .A(n38751), .B(n38752), .Z(n15752) );
  XNOR U41686 ( .A(n15748), .B(n15750), .Z(n38752) );
  XNOR U41687 ( .A(q[8]), .B(DB[3203]), .Z(n15750) );
  XNOR U41688 ( .A(q[11]), .B(DB[3206]), .Z(n15748) );
  IV U41689 ( .A(n15747), .Z(n38751) );
  XNOR U41690 ( .A(n15745), .B(n38753), .Z(n15747) );
  XNOR U41691 ( .A(q[10]), .B(DB[3205]), .Z(n38753) );
  XNOR U41692 ( .A(q[9]), .B(DB[3204]), .Z(n15745) );
  IV U41693 ( .A(n15760), .Z(n38747) );
  XOR U41694 ( .A(n38754), .B(n38755), .Z(n15760) );
  XNOR U41695 ( .A(n15777), .B(n15758), .Z(n38755) );
  XNOR U41696 ( .A(q[0]), .B(DB[3195]), .Z(n15758) );
  XOR U41697 ( .A(n38756), .B(n15766), .Z(n15777) );
  XNOR U41698 ( .A(q[7]), .B(DB[3202]), .Z(n15766) );
  IV U41699 ( .A(n15765), .Z(n38756) );
  XNOR U41700 ( .A(n15763), .B(n38757), .Z(n15765) );
  XNOR U41701 ( .A(q[6]), .B(DB[3201]), .Z(n38757) );
  XNOR U41702 ( .A(q[5]), .B(DB[3200]), .Z(n15763) );
  IV U41703 ( .A(n15776), .Z(n38754) );
  XOR U41704 ( .A(n38758), .B(n38759), .Z(n15776) );
  XNOR U41705 ( .A(n15772), .B(n15774), .Z(n38759) );
  XNOR U41706 ( .A(q[1]), .B(DB[3196]), .Z(n15774) );
  XNOR U41707 ( .A(q[4]), .B(DB[3199]), .Z(n15772) );
  IV U41708 ( .A(n15771), .Z(n38758) );
  XNOR U41709 ( .A(n15769), .B(n38760), .Z(n15771) );
  XNOR U41710 ( .A(q[3]), .B(DB[3198]), .Z(n38760) );
  XNOR U41711 ( .A(q[2]), .B(DB[3197]), .Z(n15769) );
  XOR U41712 ( .A(n38761), .B(n15667), .Z(n15595) );
  XOR U41713 ( .A(n38762), .B(n15659), .Z(n15667) );
  XOR U41714 ( .A(n38763), .B(n15648), .Z(n15659) );
  XNOR U41715 ( .A(q[14]), .B(DB[3224]), .Z(n15648) );
  IV U41716 ( .A(n15647), .Z(n38763) );
  XNOR U41717 ( .A(n15645), .B(n38764), .Z(n15647) );
  XNOR U41718 ( .A(q[13]), .B(DB[3223]), .Z(n38764) );
  XNOR U41719 ( .A(q[12]), .B(DB[3222]), .Z(n15645) );
  IV U41720 ( .A(n15658), .Z(n38762) );
  XOR U41721 ( .A(n38765), .B(n38766), .Z(n15658) );
  XNOR U41722 ( .A(n15654), .B(n15656), .Z(n38766) );
  XNOR U41723 ( .A(q[8]), .B(DB[3218]), .Z(n15656) );
  XNOR U41724 ( .A(q[11]), .B(DB[3221]), .Z(n15654) );
  IV U41725 ( .A(n15653), .Z(n38765) );
  XNOR U41726 ( .A(n15651), .B(n38767), .Z(n15653) );
  XNOR U41727 ( .A(q[10]), .B(DB[3220]), .Z(n38767) );
  XNOR U41728 ( .A(q[9]), .B(DB[3219]), .Z(n15651) );
  IV U41729 ( .A(n15666), .Z(n38761) );
  XOR U41730 ( .A(n38768), .B(n38769), .Z(n15666) );
  XNOR U41731 ( .A(n15683), .B(n15664), .Z(n38769) );
  XNOR U41732 ( .A(q[0]), .B(DB[3210]), .Z(n15664) );
  XOR U41733 ( .A(n38770), .B(n15672), .Z(n15683) );
  XNOR U41734 ( .A(q[7]), .B(DB[3217]), .Z(n15672) );
  IV U41735 ( .A(n15671), .Z(n38770) );
  XNOR U41736 ( .A(n15669), .B(n38771), .Z(n15671) );
  XNOR U41737 ( .A(q[6]), .B(DB[3216]), .Z(n38771) );
  XNOR U41738 ( .A(q[5]), .B(DB[3215]), .Z(n15669) );
  IV U41739 ( .A(n15682), .Z(n38768) );
  XOR U41740 ( .A(n38772), .B(n38773), .Z(n15682) );
  XNOR U41741 ( .A(n15678), .B(n15680), .Z(n38773) );
  XNOR U41742 ( .A(q[1]), .B(DB[3211]), .Z(n15680) );
  XNOR U41743 ( .A(q[4]), .B(DB[3214]), .Z(n15678) );
  IV U41744 ( .A(n15677), .Z(n38772) );
  XNOR U41745 ( .A(n15675), .B(n38774), .Z(n15677) );
  XNOR U41746 ( .A(q[3]), .B(DB[3213]), .Z(n38774) );
  XNOR U41747 ( .A(q[2]), .B(DB[3212]), .Z(n15675) );
  XOR U41748 ( .A(n38775), .B(n15573), .Z(n15501) );
  XOR U41749 ( .A(n38776), .B(n15565), .Z(n15573) );
  XOR U41750 ( .A(n38777), .B(n15554), .Z(n15565) );
  XNOR U41751 ( .A(q[14]), .B(DB[3239]), .Z(n15554) );
  IV U41752 ( .A(n15553), .Z(n38777) );
  XNOR U41753 ( .A(n15551), .B(n38778), .Z(n15553) );
  XNOR U41754 ( .A(q[13]), .B(DB[3238]), .Z(n38778) );
  XNOR U41755 ( .A(q[12]), .B(DB[3237]), .Z(n15551) );
  IV U41756 ( .A(n15564), .Z(n38776) );
  XOR U41757 ( .A(n38779), .B(n38780), .Z(n15564) );
  XNOR U41758 ( .A(n15560), .B(n15562), .Z(n38780) );
  XNOR U41759 ( .A(q[8]), .B(DB[3233]), .Z(n15562) );
  XNOR U41760 ( .A(q[11]), .B(DB[3236]), .Z(n15560) );
  IV U41761 ( .A(n15559), .Z(n38779) );
  XNOR U41762 ( .A(n15557), .B(n38781), .Z(n15559) );
  XNOR U41763 ( .A(q[10]), .B(DB[3235]), .Z(n38781) );
  XNOR U41764 ( .A(q[9]), .B(DB[3234]), .Z(n15557) );
  IV U41765 ( .A(n15572), .Z(n38775) );
  XOR U41766 ( .A(n38782), .B(n38783), .Z(n15572) );
  XNOR U41767 ( .A(n15589), .B(n15570), .Z(n38783) );
  XNOR U41768 ( .A(q[0]), .B(DB[3225]), .Z(n15570) );
  XOR U41769 ( .A(n38784), .B(n15578), .Z(n15589) );
  XNOR U41770 ( .A(q[7]), .B(DB[3232]), .Z(n15578) );
  IV U41771 ( .A(n15577), .Z(n38784) );
  XNOR U41772 ( .A(n15575), .B(n38785), .Z(n15577) );
  XNOR U41773 ( .A(q[6]), .B(DB[3231]), .Z(n38785) );
  XNOR U41774 ( .A(q[5]), .B(DB[3230]), .Z(n15575) );
  IV U41775 ( .A(n15588), .Z(n38782) );
  XOR U41776 ( .A(n38786), .B(n38787), .Z(n15588) );
  XNOR U41777 ( .A(n15584), .B(n15586), .Z(n38787) );
  XNOR U41778 ( .A(q[1]), .B(DB[3226]), .Z(n15586) );
  XNOR U41779 ( .A(q[4]), .B(DB[3229]), .Z(n15584) );
  IV U41780 ( .A(n15583), .Z(n38786) );
  XNOR U41781 ( .A(n15581), .B(n38788), .Z(n15583) );
  XNOR U41782 ( .A(q[3]), .B(DB[3228]), .Z(n38788) );
  XNOR U41783 ( .A(q[2]), .B(DB[3227]), .Z(n15581) );
  XOR U41784 ( .A(n38789), .B(n15479), .Z(n15407) );
  XOR U41785 ( .A(n38790), .B(n15471), .Z(n15479) );
  XOR U41786 ( .A(n38791), .B(n15460), .Z(n15471) );
  XNOR U41787 ( .A(q[14]), .B(DB[3254]), .Z(n15460) );
  IV U41788 ( .A(n15459), .Z(n38791) );
  XNOR U41789 ( .A(n15457), .B(n38792), .Z(n15459) );
  XNOR U41790 ( .A(q[13]), .B(DB[3253]), .Z(n38792) );
  XNOR U41791 ( .A(q[12]), .B(DB[3252]), .Z(n15457) );
  IV U41792 ( .A(n15470), .Z(n38790) );
  XOR U41793 ( .A(n38793), .B(n38794), .Z(n15470) );
  XNOR U41794 ( .A(n15466), .B(n15468), .Z(n38794) );
  XNOR U41795 ( .A(q[8]), .B(DB[3248]), .Z(n15468) );
  XNOR U41796 ( .A(q[11]), .B(DB[3251]), .Z(n15466) );
  IV U41797 ( .A(n15465), .Z(n38793) );
  XNOR U41798 ( .A(n15463), .B(n38795), .Z(n15465) );
  XNOR U41799 ( .A(q[10]), .B(DB[3250]), .Z(n38795) );
  XNOR U41800 ( .A(q[9]), .B(DB[3249]), .Z(n15463) );
  IV U41801 ( .A(n15478), .Z(n38789) );
  XOR U41802 ( .A(n38796), .B(n38797), .Z(n15478) );
  XNOR U41803 ( .A(n15495), .B(n15476), .Z(n38797) );
  XNOR U41804 ( .A(q[0]), .B(DB[3240]), .Z(n15476) );
  XOR U41805 ( .A(n38798), .B(n15484), .Z(n15495) );
  XNOR U41806 ( .A(q[7]), .B(DB[3247]), .Z(n15484) );
  IV U41807 ( .A(n15483), .Z(n38798) );
  XNOR U41808 ( .A(n15481), .B(n38799), .Z(n15483) );
  XNOR U41809 ( .A(q[6]), .B(DB[3246]), .Z(n38799) );
  XNOR U41810 ( .A(q[5]), .B(DB[3245]), .Z(n15481) );
  IV U41811 ( .A(n15494), .Z(n38796) );
  XOR U41812 ( .A(n38800), .B(n38801), .Z(n15494) );
  XNOR U41813 ( .A(n15490), .B(n15492), .Z(n38801) );
  XNOR U41814 ( .A(q[1]), .B(DB[3241]), .Z(n15492) );
  XNOR U41815 ( .A(q[4]), .B(DB[3244]), .Z(n15490) );
  IV U41816 ( .A(n15489), .Z(n38800) );
  XNOR U41817 ( .A(n15487), .B(n38802), .Z(n15489) );
  XNOR U41818 ( .A(q[3]), .B(DB[3243]), .Z(n38802) );
  XNOR U41819 ( .A(q[2]), .B(DB[3242]), .Z(n15487) );
  XOR U41820 ( .A(n38803), .B(n15385), .Z(n15313) );
  XOR U41821 ( .A(n38804), .B(n15377), .Z(n15385) );
  XOR U41822 ( .A(n38805), .B(n15366), .Z(n15377) );
  XNOR U41823 ( .A(q[14]), .B(DB[3269]), .Z(n15366) );
  IV U41824 ( .A(n15365), .Z(n38805) );
  XNOR U41825 ( .A(n15363), .B(n38806), .Z(n15365) );
  XNOR U41826 ( .A(q[13]), .B(DB[3268]), .Z(n38806) );
  XNOR U41827 ( .A(q[12]), .B(DB[3267]), .Z(n15363) );
  IV U41828 ( .A(n15376), .Z(n38804) );
  XOR U41829 ( .A(n38807), .B(n38808), .Z(n15376) );
  XNOR U41830 ( .A(n15372), .B(n15374), .Z(n38808) );
  XNOR U41831 ( .A(q[8]), .B(DB[3263]), .Z(n15374) );
  XNOR U41832 ( .A(q[11]), .B(DB[3266]), .Z(n15372) );
  IV U41833 ( .A(n15371), .Z(n38807) );
  XNOR U41834 ( .A(n15369), .B(n38809), .Z(n15371) );
  XNOR U41835 ( .A(q[10]), .B(DB[3265]), .Z(n38809) );
  XNOR U41836 ( .A(q[9]), .B(DB[3264]), .Z(n15369) );
  IV U41837 ( .A(n15384), .Z(n38803) );
  XOR U41838 ( .A(n38810), .B(n38811), .Z(n15384) );
  XNOR U41839 ( .A(n15401), .B(n15382), .Z(n38811) );
  XNOR U41840 ( .A(q[0]), .B(DB[3255]), .Z(n15382) );
  XOR U41841 ( .A(n38812), .B(n15390), .Z(n15401) );
  XNOR U41842 ( .A(q[7]), .B(DB[3262]), .Z(n15390) );
  IV U41843 ( .A(n15389), .Z(n38812) );
  XNOR U41844 ( .A(n15387), .B(n38813), .Z(n15389) );
  XNOR U41845 ( .A(q[6]), .B(DB[3261]), .Z(n38813) );
  XNOR U41846 ( .A(q[5]), .B(DB[3260]), .Z(n15387) );
  IV U41847 ( .A(n15400), .Z(n38810) );
  XOR U41848 ( .A(n38814), .B(n38815), .Z(n15400) );
  XNOR U41849 ( .A(n15396), .B(n15398), .Z(n38815) );
  XNOR U41850 ( .A(q[1]), .B(DB[3256]), .Z(n15398) );
  XNOR U41851 ( .A(q[4]), .B(DB[3259]), .Z(n15396) );
  IV U41852 ( .A(n15395), .Z(n38814) );
  XNOR U41853 ( .A(n15393), .B(n38816), .Z(n15395) );
  XNOR U41854 ( .A(q[3]), .B(DB[3258]), .Z(n38816) );
  XNOR U41855 ( .A(q[2]), .B(DB[3257]), .Z(n15393) );
  XOR U41856 ( .A(n38817), .B(n15291), .Z(n15219) );
  XOR U41857 ( .A(n38818), .B(n15283), .Z(n15291) );
  XOR U41858 ( .A(n38819), .B(n15272), .Z(n15283) );
  XNOR U41859 ( .A(q[14]), .B(DB[3284]), .Z(n15272) );
  IV U41860 ( .A(n15271), .Z(n38819) );
  XNOR U41861 ( .A(n15269), .B(n38820), .Z(n15271) );
  XNOR U41862 ( .A(q[13]), .B(DB[3283]), .Z(n38820) );
  XNOR U41863 ( .A(q[12]), .B(DB[3282]), .Z(n15269) );
  IV U41864 ( .A(n15282), .Z(n38818) );
  XOR U41865 ( .A(n38821), .B(n38822), .Z(n15282) );
  XNOR U41866 ( .A(n15278), .B(n15280), .Z(n38822) );
  XNOR U41867 ( .A(q[8]), .B(DB[3278]), .Z(n15280) );
  XNOR U41868 ( .A(q[11]), .B(DB[3281]), .Z(n15278) );
  IV U41869 ( .A(n15277), .Z(n38821) );
  XNOR U41870 ( .A(n15275), .B(n38823), .Z(n15277) );
  XNOR U41871 ( .A(q[10]), .B(DB[3280]), .Z(n38823) );
  XNOR U41872 ( .A(q[9]), .B(DB[3279]), .Z(n15275) );
  IV U41873 ( .A(n15290), .Z(n38817) );
  XOR U41874 ( .A(n38824), .B(n38825), .Z(n15290) );
  XNOR U41875 ( .A(n15307), .B(n15288), .Z(n38825) );
  XNOR U41876 ( .A(q[0]), .B(DB[3270]), .Z(n15288) );
  XOR U41877 ( .A(n38826), .B(n15296), .Z(n15307) );
  XNOR U41878 ( .A(q[7]), .B(DB[3277]), .Z(n15296) );
  IV U41879 ( .A(n15295), .Z(n38826) );
  XNOR U41880 ( .A(n15293), .B(n38827), .Z(n15295) );
  XNOR U41881 ( .A(q[6]), .B(DB[3276]), .Z(n38827) );
  XNOR U41882 ( .A(q[5]), .B(DB[3275]), .Z(n15293) );
  IV U41883 ( .A(n15306), .Z(n38824) );
  XOR U41884 ( .A(n38828), .B(n38829), .Z(n15306) );
  XNOR U41885 ( .A(n15302), .B(n15304), .Z(n38829) );
  XNOR U41886 ( .A(q[1]), .B(DB[3271]), .Z(n15304) );
  XNOR U41887 ( .A(q[4]), .B(DB[3274]), .Z(n15302) );
  IV U41888 ( .A(n15301), .Z(n38828) );
  XNOR U41889 ( .A(n15299), .B(n38830), .Z(n15301) );
  XNOR U41890 ( .A(q[3]), .B(DB[3273]), .Z(n38830) );
  XNOR U41891 ( .A(q[2]), .B(DB[3272]), .Z(n15299) );
  XOR U41892 ( .A(n38831), .B(n15197), .Z(n15125) );
  XOR U41893 ( .A(n38832), .B(n15189), .Z(n15197) );
  XOR U41894 ( .A(n38833), .B(n15178), .Z(n15189) );
  XNOR U41895 ( .A(q[14]), .B(DB[3299]), .Z(n15178) );
  IV U41896 ( .A(n15177), .Z(n38833) );
  XNOR U41897 ( .A(n15175), .B(n38834), .Z(n15177) );
  XNOR U41898 ( .A(q[13]), .B(DB[3298]), .Z(n38834) );
  XNOR U41899 ( .A(q[12]), .B(DB[3297]), .Z(n15175) );
  IV U41900 ( .A(n15188), .Z(n38832) );
  XOR U41901 ( .A(n38835), .B(n38836), .Z(n15188) );
  XNOR U41902 ( .A(n15184), .B(n15186), .Z(n38836) );
  XNOR U41903 ( .A(q[8]), .B(DB[3293]), .Z(n15186) );
  XNOR U41904 ( .A(q[11]), .B(DB[3296]), .Z(n15184) );
  IV U41905 ( .A(n15183), .Z(n38835) );
  XNOR U41906 ( .A(n15181), .B(n38837), .Z(n15183) );
  XNOR U41907 ( .A(q[10]), .B(DB[3295]), .Z(n38837) );
  XNOR U41908 ( .A(q[9]), .B(DB[3294]), .Z(n15181) );
  IV U41909 ( .A(n15196), .Z(n38831) );
  XOR U41910 ( .A(n38838), .B(n38839), .Z(n15196) );
  XNOR U41911 ( .A(n15213), .B(n15194), .Z(n38839) );
  XNOR U41912 ( .A(q[0]), .B(DB[3285]), .Z(n15194) );
  XOR U41913 ( .A(n38840), .B(n15202), .Z(n15213) );
  XNOR U41914 ( .A(q[7]), .B(DB[3292]), .Z(n15202) );
  IV U41915 ( .A(n15201), .Z(n38840) );
  XNOR U41916 ( .A(n15199), .B(n38841), .Z(n15201) );
  XNOR U41917 ( .A(q[6]), .B(DB[3291]), .Z(n38841) );
  XNOR U41918 ( .A(q[5]), .B(DB[3290]), .Z(n15199) );
  IV U41919 ( .A(n15212), .Z(n38838) );
  XOR U41920 ( .A(n38842), .B(n38843), .Z(n15212) );
  XNOR U41921 ( .A(n15208), .B(n15210), .Z(n38843) );
  XNOR U41922 ( .A(q[1]), .B(DB[3286]), .Z(n15210) );
  XNOR U41923 ( .A(q[4]), .B(DB[3289]), .Z(n15208) );
  IV U41924 ( .A(n15207), .Z(n38842) );
  XNOR U41925 ( .A(n15205), .B(n38844), .Z(n15207) );
  XNOR U41926 ( .A(q[3]), .B(DB[3288]), .Z(n38844) );
  XNOR U41927 ( .A(q[2]), .B(DB[3287]), .Z(n15205) );
  XOR U41928 ( .A(n38845), .B(n15103), .Z(n15031) );
  XOR U41929 ( .A(n38846), .B(n15095), .Z(n15103) );
  XOR U41930 ( .A(n38847), .B(n15084), .Z(n15095) );
  XNOR U41931 ( .A(q[14]), .B(DB[3314]), .Z(n15084) );
  IV U41932 ( .A(n15083), .Z(n38847) );
  XNOR U41933 ( .A(n15081), .B(n38848), .Z(n15083) );
  XNOR U41934 ( .A(q[13]), .B(DB[3313]), .Z(n38848) );
  XNOR U41935 ( .A(q[12]), .B(DB[3312]), .Z(n15081) );
  IV U41936 ( .A(n15094), .Z(n38846) );
  XOR U41937 ( .A(n38849), .B(n38850), .Z(n15094) );
  XNOR U41938 ( .A(n15090), .B(n15092), .Z(n38850) );
  XNOR U41939 ( .A(q[8]), .B(DB[3308]), .Z(n15092) );
  XNOR U41940 ( .A(q[11]), .B(DB[3311]), .Z(n15090) );
  IV U41941 ( .A(n15089), .Z(n38849) );
  XNOR U41942 ( .A(n15087), .B(n38851), .Z(n15089) );
  XNOR U41943 ( .A(q[10]), .B(DB[3310]), .Z(n38851) );
  XNOR U41944 ( .A(q[9]), .B(DB[3309]), .Z(n15087) );
  IV U41945 ( .A(n15102), .Z(n38845) );
  XOR U41946 ( .A(n38852), .B(n38853), .Z(n15102) );
  XNOR U41947 ( .A(n15119), .B(n15100), .Z(n38853) );
  XNOR U41948 ( .A(q[0]), .B(DB[3300]), .Z(n15100) );
  XOR U41949 ( .A(n38854), .B(n15108), .Z(n15119) );
  XNOR U41950 ( .A(q[7]), .B(DB[3307]), .Z(n15108) );
  IV U41951 ( .A(n15107), .Z(n38854) );
  XNOR U41952 ( .A(n15105), .B(n38855), .Z(n15107) );
  XNOR U41953 ( .A(q[6]), .B(DB[3306]), .Z(n38855) );
  XNOR U41954 ( .A(q[5]), .B(DB[3305]), .Z(n15105) );
  IV U41955 ( .A(n15118), .Z(n38852) );
  XOR U41956 ( .A(n38856), .B(n38857), .Z(n15118) );
  XNOR U41957 ( .A(n15114), .B(n15116), .Z(n38857) );
  XNOR U41958 ( .A(q[1]), .B(DB[3301]), .Z(n15116) );
  XNOR U41959 ( .A(q[4]), .B(DB[3304]), .Z(n15114) );
  IV U41960 ( .A(n15113), .Z(n38856) );
  XNOR U41961 ( .A(n15111), .B(n38858), .Z(n15113) );
  XNOR U41962 ( .A(q[3]), .B(DB[3303]), .Z(n38858) );
  XNOR U41963 ( .A(q[2]), .B(DB[3302]), .Z(n15111) );
  XOR U41964 ( .A(n38859), .B(n15009), .Z(n14937) );
  XOR U41965 ( .A(n38860), .B(n15001), .Z(n15009) );
  XOR U41966 ( .A(n38861), .B(n14990), .Z(n15001) );
  XNOR U41967 ( .A(q[14]), .B(DB[3329]), .Z(n14990) );
  IV U41968 ( .A(n14989), .Z(n38861) );
  XNOR U41969 ( .A(n14987), .B(n38862), .Z(n14989) );
  XNOR U41970 ( .A(q[13]), .B(DB[3328]), .Z(n38862) );
  XNOR U41971 ( .A(q[12]), .B(DB[3327]), .Z(n14987) );
  IV U41972 ( .A(n15000), .Z(n38860) );
  XOR U41973 ( .A(n38863), .B(n38864), .Z(n15000) );
  XNOR U41974 ( .A(n14996), .B(n14998), .Z(n38864) );
  XNOR U41975 ( .A(q[8]), .B(DB[3323]), .Z(n14998) );
  XNOR U41976 ( .A(q[11]), .B(DB[3326]), .Z(n14996) );
  IV U41977 ( .A(n14995), .Z(n38863) );
  XNOR U41978 ( .A(n14993), .B(n38865), .Z(n14995) );
  XNOR U41979 ( .A(q[10]), .B(DB[3325]), .Z(n38865) );
  XNOR U41980 ( .A(q[9]), .B(DB[3324]), .Z(n14993) );
  IV U41981 ( .A(n15008), .Z(n38859) );
  XOR U41982 ( .A(n38866), .B(n38867), .Z(n15008) );
  XNOR U41983 ( .A(n15025), .B(n15006), .Z(n38867) );
  XNOR U41984 ( .A(q[0]), .B(DB[3315]), .Z(n15006) );
  XOR U41985 ( .A(n38868), .B(n15014), .Z(n15025) );
  XNOR U41986 ( .A(q[7]), .B(DB[3322]), .Z(n15014) );
  IV U41987 ( .A(n15013), .Z(n38868) );
  XNOR U41988 ( .A(n15011), .B(n38869), .Z(n15013) );
  XNOR U41989 ( .A(q[6]), .B(DB[3321]), .Z(n38869) );
  XNOR U41990 ( .A(q[5]), .B(DB[3320]), .Z(n15011) );
  IV U41991 ( .A(n15024), .Z(n38866) );
  XOR U41992 ( .A(n38870), .B(n38871), .Z(n15024) );
  XNOR U41993 ( .A(n15020), .B(n15022), .Z(n38871) );
  XNOR U41994 ( .A(q[1]), .B(DB[3316]), .Z(n15022) );
  XNOR U41995 ( .A(q[4]), .B(DB[3319]), .Z(n15020) );
  IV U41996 ( .A(n15019), .Z(n38870) );
  XNOR U41997 ( .A(n15017), .B(n38872), .Z(n15019) );
  XNOR U41998 ( .A(q[3]), .B(DB[3318]), .Z(n38872) );
  XNOR U41999 ( .A(q[2]), .B(DB[3317]), .Z(n15017) );
  XOR U42000 ( .A(n38873), .B(n14915), .Z(n14843) );
  XOR U42001 ( .A(n38874), .B(n14907), .Z(n14915) );
  XOR U42002 ( .A(n38875), .B(n14896), .Z(n14907) );
  XNOR U42003 ( .A(q[14]), .B(DB[3344]), .Z(n14896) );
  IV U42004 ( .A(n14895), .Z(n38875) );
  XNOR U42005 ( .A(n14893), .B(n38876), .Z(n14895) );
  XNOR U42006 ( .A(q[13]), .B(DB[3343]), .Z(n38876) );
  XNOR U42007 ( .A(q[12]), .B(DB[3342]), .Z(n14893) );
  IV U42008 ( .A(n14906), .Z(n38874) );
  XOR U42009 ( .A(n38877), .B(n38878), .Z(n14906) );
  XNOR U42010 ( .A(n14902), .B(n14904), .Z(n38878) );
  XNOR U42011 ( .A(q[8]), .B(DB[3338]), .Z(n14904) );
  XNOR U42012 ( .A(q[11]), .B(DB[3341]), .Z(n14902) );
  IV U42013 ( .A(n14901), .Z(n38877) );
  XNOR U42014 ( .A(n14899), .B(n38879), .Z(n14901) );
  XNOR U42015 ( .A(q[10]), .B(DB[3340]), .Z(n38879) );
  XNOR U42016 ( .A(q[9]), .B(DB[3339]), .Z(n14899) );
  IV U42017 ( .A(n14914), .Z(n38873) );
  XOR U42018 ( .A(n38880), .B(n38881), .Z(n14914) );
  XNOR U42019 ( .A(n14931), .B(n14912), .Z(n38881) );
  XNOR U42020 ( .A(q[0]), .B(DB[3330]), .Z(n14912) );
  XOR U42021 ( .A(n38882), .B(n14920), .Z(n14931) );
  XNOR U42022 ( .A(q[7]), .B(DB[3337]), .Z(n14920) );
  IV U42023 ( .A(n14919), .Z(n38882) );
  XNOR U42024 ( .A(n14917), .B(n38883), .Z(n14919) );
  XNOR U42025 ( .A(q[6]), .B(DB[3336]), .Z(n38883) );
  XNOR U42026 ( .A(q[5]), .B(DB[3335]), .Z(n14917) );
  IV U42027 ( .A(n14930), .Z(n38880) );
  XOR U42028 ( .A(n38884), .B(n38885), .Z(n14930) );
  XNOR U42029 ( .A(n14926), .B(n14928), .Z(n38885) );
  XNOR U42030 ( .A(q[1]), .B(DB[3331]), .Z(n14928) );
  XNOR U42031 ( .A(q[4]), .B(DB[3334]), .Z(n14926) );
  IV U42032 ( .A(n14925), .Z(n38884) );
  XNOR U42033 ( .A(n14923), .B(n38886), .Z(n14925) );
  XNOR U42034 ( .A(q[3]), .B(DB[3333]), .Z(n38886) );
  XNOR U42035 ( .A(q[2]), .B(DB[3332]), .Z(n14923) );
  XOR U42036 ( .A(n38887), .B(n14821), .Z(n14749) );
  XOR U42037 ( .A(n38888), .B(n14813), .Z(n14821) );
  XOR U42038 ( .A(n38889), .B(n14802), .Z(n14813) );
  XNOR U42039 ( .A(q[14]), .B(DB[3359]), .Z(n14802) );
  IV U42040 ( .A(n14801), .Z(n38889) );
  XNOR U42041 ( .A(n14799), .B(n38890), .Z(n14801) );
  XNOR U42042 ( .A(q[13]), .B(DB[3358]), .Z(n38890) );
  XNOR U42043 ( .A(q[12]), .B(DB[3357]), .Z(n14799) );
  IV U42044 ( .A(n14812), .Z(n38888) );
  XOR U42045 ( .A(n38891), .B(n38892), .Z(n14812) );
  XNOR U42046 ( .A(n14808), .B(n14810), .Z(n38892) );
  XNOR U42047 ( .A(q[8]), .B(DB[3353]), .Z(n14810) );
  XNOR U42048 ( .A(q[11]), .B(DB[3356]), .Z(n14808) );
  IV U42049 ( .A(n14807), .Z(n38891) );
  XNOR U42050 ( .A(n14805), .B(n38893), .Z(n14807) );
  XNOR U42051 ( .A(q[10]), .B(DB[3355]), .Z(n38893) );
  XNOR U42052 ( .A(q[9]), .B(DB[3354]), .Z(n14805) );
  IV U42053 ( .A(n14820), .Z(n38887) );
  XOR U42054 ( .A(n38894), .B(n38895), .Z(n14820) );
  XNOR U42055 ( .A(n14837), .B(n14818), .Z(n38895) );
  XNOR U42056 ( .A(q[0]), .B(DB[3345]), .Z(n14818) );
  XOR U42057 ( .A(n38896), .B(n14826), .Z(n14837) );
  XNOR U42058 ( .A(q[7]), .B(DB[3352]), .Z(n14826) );
  IV U42059 ( .A(n14825), .Z(n38896) );
  XNOR U42060 ( .A(n14823), .B(n38897), .Z(n14825) );
  XNOR U42061 ( .A(q[6]), .B(DB[3351]), .Z(n38897) );
  XNOR U42062 ( .A(q[5]), .B(DB[3350]), .Z(n14823) );
  IV U42063 ( .A(n14836), .Z(n38894) );
  XOR U42064 ( .A(n38898), .B(n38899), .Z(n14836) );
  XNOR U42065 ( .A(n14832), .B(n14834), .Z(n38899) );
  XNOR U42066 ( .A(q[1]), .B(DB[3346]), .Z(n14834) );
  XNOR U42067 ( .A(q[4]), .B(DB[3349]), .Z(n14832) );
  IV U42068 ( .A(n14831), .Z(n38898) );
  XNOR U42069 ( .A(n14829), .B(n38900), .Z(n14831) );
  XNOR U42070 ( .A(q[3]), .B(DB[3348]), .Z(n38900) );
  XNOR U42071 ( .A(q[2]), .B(DB[3347]), .Z(n14829) );
  XOR U42072 ( .A(n38901), .B(n14727), .Z(n14655) );
  XOR U42073 ( .A(n38902), .B(n14719), .Z(n14727) );
  XOR U42074 ( .A(n38903), .B(n14708), .Z(n14719) );
  XNOR U42075 ( .A(q[14]), .B(DB[3374]), .Z(n14708) );
  IV U42076 ( .A(n14707), .Z(n38903) );
  XNOR U42077 ( .A(n14705), .B(n38904), .Z(n14707) );
  XNOR U42078 ( .A(q[13]), .B(DB[3373]), .Z(n38904) );
  XNOR U42079 ( .A(q[12]), .B(DB[3372]), .Z(n14705) );
  IV U42080 ( .A(n14718), .Z(n38902) );
  XOR U42081 ( .A(n38905), .B(n38906), .Z(n14718) );
  XNOR U42082 ( .A(n14714), .B(n14716), .Z(n38906) );
  XNOR U42083 ( .A(q[8]), .B(DB[3368]), .Z(n14716) );
  XNOR U42084 ( .A(q[11]), .B(DB[3371]), .Z(n14714) );
  IV U42085 ( .A(n14713), .Z(n38905) );
  XNOR U42086 ( .A(n14711), .B(n38907), .Z(n14713) );
  XNOR U42087 ( .A(q[10]), .B(DB[3370]), .Z(n38907) );
  XNOR U42088 ( .A(q[9]), .B(DB[3369]), .Z(n14711) );
  IV U42089 ( .A(n14726), .Z(n38901) );
  XOR U42090 ( .A(n38908), .B(n38909), .Z(n14726) );
  XNOR U42091 ( .A(n14743), .B(n14724), .Z(n38909) );
  XNOR U42092 ( .A(q[0]), .B(DB[3360]), .Z(n14724) );
  XOR U42093 ( .A(n38910), .B(n14732), .Z(n14743) );
  XNOR U42094 ( .A(q[7]), .B(DB[3367]), .Z(n14732) );
  IV U42095 ( .A(n14731), .Z(n38910) );
  XNOR U42096 ( .A(n14729), .B(n38911), .Z(n14731) );
  XNOR U42097 ( .A(q[6]), .B(DB[3366]), .Z(n38911) );
  XNOR U42098 ( .A(q[5]), .B(DB[3365]), .Z(n14729) );
  IV U42099 ( .A(n14742), .Z(n38908) );
  XOR U42100 ( .A(n38912), .B(n38913), .Z(n14742) );
  XNOR U42101 ( .A(n14738), .B(n14740), .Z(n38913) );
  XNOR U42102 ( .A(q[1]), .B(DB[3361]), .Z(n14740) );
  XNOR U42103 ( .A(q[4]), .B(DB[3364]), .Z(n14738) );
  IV U42104 ( .A(n14737), .Z(n38912) );
  XNOR U42105 ( .A(n14735), .B(n38914), .Z(n14737) );
  XNOR U42106 ( .A(q[3]), .B(DB[3363]), .Z(n38914) );
  XNOR U42107 ( .A(q[2]), .B(DB[3362]), .Z(n14735) );
  XOR U42108 ( .A(n38915), .B(n14633), .Z(n14561) );
  XOR U42109 ( .A(n38916), .B(n14625), .Z(n14633) );
  XOR U42110 ( .A(n38917), .B(n14614), .Z(n14625) );
  XNOR U42111 ( .A(q[14]), .B(DB[3389]), .Z(n14614) );
  IV U42112 ( .A(n14613), .Z(n38917) );
  XNOR U42113 ( .A(n14611), .B(n38918), .Z(n14613) );
  XNOR U42114 ( .A(q[13]), .B(DB[3388]), .Z(n38918) );
  XNOR U42115 ( .A(q[12]), .B(DB[3387]), .Z(n14611) );
  IV U42116 ( .A(n14624), .Z(n38916) );
  XOR U42117 ( .A(n38919), .B(n38920), .Z(n14624) );
  XNOR U42118 ( .A(n14620), .B(n14622), .Z(n38920) );
  XNOR U42119 ( .A(q[8]), .B(DB[3383]), .Z(n14622) );
  XNOR U42120 ( .A(q[11]), .B(DB[3386]), .Z(n14620) );
  IV U42121 ( .A(n14619), .Z(n38919) );
  XNOR U42122 ( .A(n14617), .B(n38921), .Z(n14619) );
  XNOR U42123 ( .A(q[10]), .B(DB[3385]), .Z(n38921) );
  XNOR U42124 ( .A(q[9]), .B(DB[3384]), .Z(n14617) );
  IV U42125 ( .A(n14632), .Z(n38915) );
  XOR U42126 ( .A(n38922), .B(n38923), .Z(n14632) );
  XNOR U42127 ( .A(n14649), .B(n14630), .Z(n38923) );
  XNOR U42128 ( .A(q[0]), .B(DB[3375]), .Z(n14630) );
  XOR U42129 ( .A(n38924), .B(n14638), .Z(n14649) );
  XNOR U42130 ( .A(q[7]), .B(DB[3382]), .Z(n14638) );
  IV U42131 ( .A(n14637), .Z(n38924) );
  XNOR U42132 ( .A(n14635), .B(n38925), .Z(n14637) );
  XNOR U42133 ( .A(q[6]), .B(DB[3381]), .Z(n38925) );
  XNOR U42134 ( .A(q[5]), .B(DB[3380]), .Z(n14635) );
  IV U42135 ( .A(n14648), .Z(n38922) );
  XOR U42136 ( .A(n38926), .B(n38927), .Z(n14648) );
  XNOR U42137 ( .A(n14644), .B(n14646), .Z(n38927) );
  XNOR U42138 ( .A(q[1]), .B(DB[3376]), .Z(n14646) );
  XNOR U42139 ( .A(q[4]), .B(DB[3379]), .Z(n14644) );
  IV U42140 ( .A(n14643), .Z(n38926) );
  XNOR U42141 ( .A(n14641), .B(n38928), .Z(n14643) );
  XNOR U42142 ( .A(q[3]), .B(DB[3378]), .Z(n38928) );
  XNOR U42143 ( .A(q[2]), .B(DB[3377]), .Z(n14641) );
  XOR U42144 ( .A(n38929), .B(n14539), .Z(n14467) );
  XOR U42145 ( .A(n38930), .B(n14531), .Z(n14539) );
  XOR U42146 ( .A(n38931), .B(n14520), .Z(n14531) );
  XNOR U42147 ( .A(q[14]), .B(DB[3404]), .Z(n14520) );
  IV U42148 ( .A(n14519), .Z(n38931) );
  XNOR U42149 ( .A(n14517), .B(n38932), .Z(n14519) );
  XNOR U42150 ( .A(q[13]), .B(DB[3403]), .Z(n38932) );
  XNOR U42151 ( .A(q[12]), .B(DB[3402]), .Z(n14517) );
  IV U42152 ( .A(n14530), .Z(n38930) );
  XOR U42153 ( .A(n38933), .B(n38934), .Z(n14530) );
  XNOR U42154 ( .A(n14526), .B(n14528), .Z(n38934) );
  XNOR U42155 ( .A(q[8]), .B(DB[3398]), .Z(n14528) );
  XNOR U42156 ( .A(q[11]), .B(DB[3401]), .Z(n14526) );
  IV U42157 ( .A(n14525), .Z(n38933) );
  XNOR U42158 ( .A(n14523), .B(n38935), .Z(n14525) );
  XNOR U42159 ( .A(q[10]), .B(DB[3400]), .Z(n38935) );
  XNOR U42160 ( .A(q[9]), .B(DB[3399]), .Z(n14523) );
  IV U42161 ( .A(n14538), .Z(n38929) );
  XOR U42162 ( .A(n38936), .B(n38937), .Z(n14538) );
  XNOR U42163 ( .A(n14555), .B(n14536), .Z(n38937) );
  XNOR U42164 ( .A(q[0]), .B(DB[3390]), .Z(n14536) );
  XOR U42165 ( .A(n38938), .B(n14544), .Z(n14555) );
  XNOR U42166 ( .A(q[7]), .B(DB[3397]), .Z(n14544) );
  IV U42167 ( .A(n14543), .Z(n38938) );
  XNOR U42168 ( .A(n14541), .B(n38939), .Z(n14543) );
  XNOR U42169 ( .A(q[6]), .B(DB[3396]), .Z(n38939) );
  XNOR U42170 ( .A(q[5]), .B(DB[3395]), .Z(n14541) );
  IV U42171 ( .A(n14554), .Z(n38936) );
  XOR U42172 ( .A(n38940), .B(n38941), .Z(n14554) );
  XNOR U42173 ( .A(n14550), .B(n14552), .Z(n38941) );
  XNOR U42174 ( .A(q[1]), .B(DB[3391]), .Z(n14552) );
  XNOR U42175 ( .A(q[4]), .B(DB[3394]), .Z(n14550) );
  IV U42176 ( .A(n14549), .Z(n38940) );
  XNOR U42177 ( .A(n14547), .B(n38942), .Z(n14549) );
  XNOR U42178 ( .A(q[3]), .B(DB[3393]), .Z(n38942) );
  XNOR U42179 ( .A(q[2]), .B(DB[3392]), .Z(n14547) );
  XOR U42180 ( .A(n38943), .B(n14445), .Z(n14373) );
  XOR U42181 ( .A(n38944), .B(n14437), .Z(n14445) );
  XOR U42182 ( .A(n38945), .B(n14426), .Z(n14437) );
  XNOR U42183 ( .A(q[14]), .B(DB[3419]), .Z(n14426) );
  IV U42184 ( .A(n14425), .Z(n38945) );
  XNOR U42185 ( .A(n14423), .B(n38946), .Z(n14425) );
  XNOR U42186 ( .A(q[13]), .B(DB[3418]), .Z(n38946) );
  XNOR U42187 ( .A(q[12]), .B(DB[3417]), .Z(n14423) );
  IV U42188 ( .A(n14436), .Z(n38944) );
  XOR U42189 ( .A(n38947), .B(n38948), .Z(n14436) );
  XNOR U42190 ( .A(n14432), .B(n14434), .Z(n38948) );
  XNOR U42191 ( .A(q[8]), .B(DB[3413]), .Z(n14434) );
  XNOR U42192 ( .A(q[11]), .B(DB[3416]), .Z(n14432) );
  IV U42193 ( .A(n14431), .Z(n38947) );
  XNOR U42194 ( .A(n14429), .B(n38949), .Z(n14431) );
  XNOR U42195 ( .A(q[10]), .B(DB[3415]), .Z(n38949) );
  XNOR U42196 ( .A(q[9]), .B(DB[3414]), .Z(n14429) );
  IV U42197 ( .A(n14444), .Z(n38943) );
  XOR U42198 ( .A(n38950), .B(n38951), .Z(n14444) );
  XNOR U42199 ( .A(n14461), .B(n14442), .Z(n38951) );
  XNOR U42200 ( .A(q[0]), .B(DB[3405]), .Z(n14442) );
  XOR U42201 ( .A(n38952), .B(n14450), .Z(n14461) );
  XNOR U42202 ( .A(q[7]), .B(DB[3412]), .Z(n14450) );
  IV U42203 ( .A(n14449), .Z(n38952) );
  XNOR U42204 ( .A(n14447), .B(n38953), .Z(n14449) );
  XNOR U42205 ( .A(q[6]), .B(DB[3411]), .Z(n38953) );
  XNOR U42206 ( .A(q[5]), .B(DB[3410]), .Z(n14447) );
  IV U42207 ( .A(n14460), .Z(n38950) );
  XOR U42208 ( .A(n38954), .B(n38955), .Z(n14460) );
  XNOR U42209 ( .A(n14456), .B(n14458), .Z(n38955) );
  XNOR U42210 ( .A(q[1]), .B(DB[3406]), .Z(n14458) );
  XNOR U42211 ( .A(q[4]), .B(DB[3409]), .Z(n14456) );
  IV U42212 ( .A(n14455), .Z(n38954) );
  XNOR U42213 ( .A(n14453), .B(n38956), .Z(n14455) );
  XNOR U42214 ( .A(q[3]), .B(DB[3408]), .Z(n38956) );
  XNOR U42215 ( .A(q[2]), .B(DB[3407]), .Z(n14453) );
  XOR U42216 ( .A(n38957), .B(n14351), .Z(n14279) );
  XOR U42217 ( .A(n38958), .B(n14343), .Z(n14351) );
  XOR U42218 ( .A(n38959), .B(n14332), .Z(n14343) );
  XNOR U42219 ( .A(q[14]), .B(DB[3434]), .Z(n14332) );
  IV U42220 ( .A(n14331), .Z(n38959) );
  XNOR U42221 ( .A(n14329), .B(n38960), .Z(n14331) );
  XNOR U42222 ( .A(q[13]), .B(DB[3433]), .Z(n38960) );
  XNOR U42223 ( .A(q[12]), .B(DB[3432]), .Z(n14329) );
  IV U42224 ( .A(n14342), .Z(n38958) );
  XOR U42225 ( .A(n38961), .B(n38962), .Z(n14342) );
  XNOR U42226 ( .A(n14338), .B(n14340), .Z(n38962) );
  XNOR U42227 ( .A(q[8]), .B(DB[3428]), .Z(n14340) );
  XNOR U42228 ( .A(q[11]), .B(DB[3431]), .Z(n14338) );
  IV U42229 ( .A(n14337), .Z(n38961) );
  XNOR U42230 ( .A(n14335), .B(n38963), .Z(n14337) );
  XNOR U42231 ( .A(q[10]), .B(DB[3430]), .Z(n38963) );
  XNOR U42232 ( .A(q[9]), .B(DB[3429]), .Z(n14335) );
  IV U42233 ( .A(n14350), .Z(n38957) );
  XOR U42234 ( .A(n38964), .B(n38965), .Z(n14350) );
  XNOR U42235 ( .A(n14367), .B(n14348), .Z(n38965) );
  XNOR U42236 ( .A(q[0]), .B(DB[3420]), .Z(n14348) );
  XOR U42237 ( .A(n38966), .B(n14356), .Z(n14367) );
  XNOR U42238 ( .A(q[7]), .B(DB[3427]), .Z(n14356) );
  IV U42239 ( .A(n14355), .Z(n38966) );
  XNOR U42240 ( .A(n14353), .B(n38967), .Z(n14355) );
  XNOR U42241 ( .A(q[6]), .B(DB[3426]), .Z(n38967) );
  XNOR U42242 ( .A(q[5]), .B(DB[3425]), .Z(n14353) );
  IV U42243 ( .A(n14366), .Z(n38964) );
  XOR U42244 ( .A(n38968), .B(n38969), .Z(n14366) );
  XNOR U42245 ( .A(n14362), .B(n14364), .Z(n38969) );
  XNOR U42246 ( .A(q[1]), .B(DB[3421]), .Z(n14364) );
  XNOR U42247 ( .A(q[4]), .B(DB[3424]), .Z(n14362) );
  IV U42248 ( .A(n14361), .Z(n38968) );
  XNOR U42249 ( .A(n14359), .B(n38970), .Z(n14361) );
  XNOR U42250 ( .A(q[3]), .B(DB[3423]), .Z(n38970) );
  XNOR U42251 ( .A(q[2]), .B(DB[3422]), .Z(n14359) );
  XOR U42252 ( .A(n38971), .B(n14257), .Z(n14185) );
  XOR U42253 ( .A(n38972), .B(n14249), .Z(n14257) );
  XOR U42254 ( .A(n38973), .B(n14238), .Z(n14249) );
  XNOR U42255 ( .A(q[14]), .B(DB[3449]), .Z(n14238) );
  IV U42256 ( .A(n14237), .Z(n38973) );
  XNOR U42257 ( .A(n14235), .B(n38974), .Z(n14237) );
  XNOR U42258 ( .A(q[13]), .B(DB[3448]), .Z(n38974) );
  XNOR U42259 ( .A(q[12]), .B(DB[3447]), .Z(n14235) );
  IV U42260 ( .A(n14248), .Z(n38972) );
  XOR U42261 ( .A(n38975), .B(n38976), .Z(n14248) );
  XNOR U42262 ( .A(n14244), .B(n14246), .Z(n38976) );
  XNOR U42263 ( .A(q[8]), .B(DB[3443]), .Z(n14246) );
  XNOR U42264 ( .A(q[11]), .B(DB[3446]), .Z(n14244) );
  IV U42265 ( .A(n14243), .Z(n38975) );
  XNOR U42266 ( .A(n14241), .B(n38977), .Z(n14243) );
  XNOR U42267 ( .A(q[10]), .B(DB[3445]), .Z(n38977) );
  XNOR U42268 ( .A(q[9]), .B(DB[3444]), .Z(n14241) );
  IV U42269 ( .A(n14256), .Z(n38971) );
  XOR U42270 ( .A(n38978), .B(n38979), .Z(n14256) );
  XNOR U42271 ( .A(n14273), .B(n14254), .Z(n38979) );
  XNOR U42272 ( .A(q[0]), .B(DB[3435]), .Z(n14254) );
  XOR U42273 ( .A(n38980), .B(n14262), .Z(n14273) );
  XNOR U42274 ( .A(q[7]), .B(DB[3442]), .Z(n14262) );
  IV U42275 ( .A(n14261), .Z(n38980) );
  XNOR U42276 ( .A(n14259), .B(n38981), .Z(n14261) );
  XNOR U42277 ( .A(q[6]), .B(DB[3441]), .Z(n38981) );
  XNOR U42278 ( .A(q[5]), .B(DB[3440]), .Z(n14259) );
  IV U42279 ( .A(n14272), .Z(n38978) );
  XOR U42280 ( .A(n38982), .B(n38983), .Z(n14272) );
  XNOR U42281 ( .A(n14268), .B(n14270), .Z(n38983) );
  XNOR U42282 ( .A(q[1]), .B(DB[3436]), .Z(n14270) );
  XNOR U42283 ( .A(q[4]), .B(DB[3439]), .Z(n14268) );
  IV U42284 ( .A(n14267), .Z(n38982) );
  XNOR U42285 ( .A(n14265), .B(n38984), .Z(n14267) );
  XNOR U42286 ( .A(q[3]), .B(DB[3438]), .Z(n38984) );
  XNOR U42287 ( .A(q[2]), .B(DB[3437]), .Z(n14265) );
  XOR U42288 ( .A(n38985), .B(n14163), .Z(n14091) );
  XOR U42289 ( .A(n38986), .B(n14155), .Z(n14163) );
  XOR U42290 ( .A(n38987), .B(n14144), .Z(n14155) );
  XNOR U42291 ( .A(q[14]), .B(DB[3464]), .Z(n14144) );
  IV U42292 ( .A(n14143), .Z(n38987) );
  XNOR U42293 ( .A(n14141), .B(n38988), .Z(n14143) );
  XNOR U42294 ( .A(q[13]), .B(DB[3463]), .Z(n38988) );
  XNOR U42295 ( .A(q[12]), .B(DB[3462]), .Z(n14141) );
  IV U42296 ( .A(n14154), .Z(n38986) );
  XOR U42297 ( .A(n38989), .B(n38990), .Z(n14154) );
  XNOR U42298 ( .A(n14150), .B(n14152), .Z(n38990) );
  XNOR U42299 ( .A(q[8]), .B(DB[3458]), .Z(n14152) );
  XNOR U42300 ( .A(q[11]), .B(DB[3461]), .Z(n14150) );
  IV U42301 ( .A(n14149), .Z(n38989) );
  XNOR U42302 ( .A(n14147), .B(n38991), .Z(n14149) );
  XNOR U42303 ( .A(q[10]), .B(DB[3460]), .Z(n38991) );
  XNOR U42304 ( .A(q[9]), .B(DB[3459]), .Z(n14147) );
  IV U42305 ( .A(n14162), .Z(n38985) );
  XOR U42306 ( .A(n38992), .B(n38993), .Z(n14162) );
  XNOR U42307 ( .A(n14179), .B(n14160), .Z(n38993) );
  XNOR U42308 ( .A(q[0]), .B(DB[3450]), .Z(n14160) );
  XOR U42309 ( .A(n38994), .B(n14168), .Z(n14179) );
  XNOR U42310 ( .A(q[7]), .B(DB[3457]), .Z(n14168) );
  IV U42311 ( .A(n14167), .Z(n38994) );
  XNOR U42312 ( .A(n14165), .B(n38995), .Z(n14167) );
  XNOR U42313 ( .A(q[6]), .B(DB[3456]), .Z(n38995) );
  XNOR U42314 ( .A(q[5]), .B(DB[3455]), .Z(n14165) );
  IV U42315 ( .A(n14178), .Z(n38992) );
  XOR U42316 ( .A(n38996), .B(n38997), .Z(n14178) );
  XNOR U42317 ( .A(n14174), .B(n14176), .Z(n38997) );
  XNOR U42318 ( .A(q[1]), .B(DB[3451]), .Z(n14176) );
  XNOR U42319 ( .A(q[4]), .B(DB[3454]), .Z(n14174) );
  IV U42320 ( .A(n14173), .Z(n38996) );
  XNOR U42321 ( .A(n14171), .B(n38998), .Z(n14173) );
  XNOR U42322 ( .A(q[3]), .B(DB[3453]), .Z(n38998) );
  XNOR U42323 ( .A(q[2]), .B(DB[3452]), .Z(n14171) );
  XOR U42324 ( .A(n38999), .B(n14069), .Z(n13997) );
  XOR U42325 ( .A(n39000), .B(n14061), .Z(n14069) );
  XOR U42326 ( .A(n39001), .B(n14050), .Z(n14061) );
  XNOR U42327 ( .A(q[14]), .B(DB[3479]), .Z(n14050) );
  IV U42328 ( .A(n14049), .Z(n39001) );
  XNOR U42329 ( .A(n14047), .B(n39002), .Z(n14049) );
  XNOR U42330 ( .A(q[13]), .B(DB[3478]), .Z(n39002) );
  XNOR U42331 ( .A(q[12]), .B(DB[3477]), .Z(n14047) );
  IV U42332 ( .A(n14060), .Z(n39000) );
  XOR U42333 ( .A(n39003), .B(n39004), .Z(n14060) );
  XNOR U42334 ( .A(n14056), .B(n14058), .Z(n39004) );
  XNOR U42335 ( .A(q[8]), .B(DB[3473]), .Z(n14058) );
  XNOR U42336 ( .A(q[11]), .B(DB[3476]), .Z(n14056) );
  IV U42337 ( .A(n14055), .Z(n39003) );
  XNOR U42338 ( .A(n14053), .B(n39005), .Z(n14055) );
  XNOR U42339 ( .A(q[10]), .B(DB[3475]), .Z(n39005) );
  XNOR U42340 ( .A(q[9]), .B(DB[3474]), .Z(n14053) );
  IV U42341 ( .A(n14068), .Z(n38999) );
  XOR U42342 ( .A(n39006), .B(n39007), .Z(n14068) );
  XNOR U42343 ( .A(n14085), .B(n14066), .Z(n39007) );
  XNOR U42344 ( .A(q[0]), .B(DB[3465]), .Z(n14066) );
  XOR U42345 ( .A(n39008), .B(n14074), .Z(n14085) );
  XNOR U42346 ( .A(q[7]), .B(DB[3472]), .Z(n14074) );
  IV U42347 ( .A(n14073), .Z(n39008) );
  XNOR U42348 ( .A(n14071), .B(n39009), .Z(n14073) );
  XNOR U42349 ( .A(q[6]), .B(DB[3471]), .Z(n39009) );
  XNOR U42350 ( .A(q[5]), .B(DB[3470]), .Z(n14071) );
  IV U42351 ( .A(n14084), .Z(n39006) );
  XOR U42352 ( .A(n39010), .B(n39011), .Z(n14084) );
  XNOR U42353 ( .A(n14080), .B(n14082), .Z(n39011) );
  XNOR U42354 ( .A(q[1]), .B(DB[3466]), .Z(n14082) );
  XNOR U42355 ( .A(q[4]), .B(DB[3469]), .Z(n14080) );
  IV U42356 ( .A(n14079), .Z(n39010) );
  XNOR U42357 ( .A(n14077), .B(n39012), .Z(n14079) );
  XNOR U42358 ( .A(q[3]), .B(DB[3468]), .Z(n39012) );
  XNOR U42359 ( .A(q[2]), .B(DB[3467]), .Z(n14077) );
  XOR U42360 ( .A(n39013), .B(n13975), .Z(n13903) );
  XOR U42361 ( .A(n39014), .B(n13967), .Z(n13975) );
  XOR U42362 ( .A(n39015), .B(n13956), .Z(n13967) );
  XNOR U42363 ( .A(q[14]), .B(DB[3494]), .Z(n13956) );
  IV U42364 ( .A(n13955), .Z(n39015) );
  XNOR U42365 ( .A(n13953), .B(n39016), .Z(n13955) );
  XNOR U42366 ( .A(q[13]), .B(DB[3493]), .Z(n39016) );
  XNOR U42367 ( .A(q[12]), .B(DB[3492]), .Z(n13953) );
  IV U42368 ( .A(n13966), .Z(n39014) );
  XOR U42369 ( .A(n39017), .B(n39018), .Z(n13966) );
  XNOR U42370 ( .A(n13962), .B(n13964), .Z(n39018) );
  XNOR U42371 ( .A(q[8]), .B(DB[3488]), .Z(n13964) );
  XNOR U42372 ( .A(q[11]), .B(DB[3491]), .Z(n13962) );
  IV U42373 ( .A(n13961), .Z(n39017) );
  XNOR U42374 ( .A(n13959), .B(n39019), .Z(n13961) );
  XNOR U42375 ( .A(q[10]), .B(DB[3490]), .Z(n39019) );
  XNOR U42376 ( .A(q[9]), .B(DB[3489]), .Z(n13959) );
  IV U42377 ( .A(n13974), .Z(n39013) );
  XOR U42378 ( .A(n39020), .B(n39021), .Z(n13974) );
  XNOR U42379 ( .A(n13991), .B(n13972), .Z(n39021) );
  XNOR U42380 ( .A(q[0]), .B(DB[3480]), .Z(n13972) );
  XOR U42381 ( .A(n39022), .B(n13980), .Z(n13991) );
  XNOR U42382 ( .A(q[7]), .B(DB[3487]), .Z(n13980) );
  IV U42383 ( .A(n13979), .Z(n39022) );
  XNOR U42384 ( .A(n13977), .B(n39023), .Z(n13979) );
  XNOR U42385 ( .A(q[6]), .B(DB[3486]), .Z(n39023) );
  XNOR U42386 ( .A(q[5]), .B(DB[3485]), .Z(n13977) );
  IV U42387 ( .A(n13990), .Z(n39020) );
  XOR U42388 ( .A(n39024), .B(n39025), .Z(n13990) );
  XNOR U42389 ( .A(n13986), .B(n13988), .Z(n39025) );
  XNOR U42390 ( .A(q[1]), .B(DB[3481]), .Z(n13988) );
  XNOR U42391 ( .A(q[4]), .B(DB[3484]), .Z(n13986) );
  IV U42392 ( .A(n13985), .Z(n39024) );
  XNOR U42393 ( .A(n13983), .B(n39026), .Z(n13985) );
  XNOR U42394 ( .A(q[3]), .B(DB[3483]), .Z(n39026) );
  XNOR U42395 ( .A(q[2]), .B(DB[3482]), .Z(n13983) );
  XOR U42396 ( .A(n39027), .B(n13881), .Z(n13809) );
  XOR U42397 ( .A(n39028), .B(n13873), .Z(n13881) );
  XOR U42398 ( .A(n39029), .B(n13862), .Z(n13873) );
  XNOR U42399 ( .A(q[14]), .B(DB[3509]), .Z(n13862) );
  IV U42400 ( .A(n13861), .Z(n39029) );
  XNOR U42401 ( .A(n13859), .B(n39030), .Z(n13861) );
  XNOR U42402 ( .A(q[13]), .B(DB[3508]), .Z(n39030) );
  XNOR U42403 ( .A(q[12]), .B(DB[3507]), .Z(n13859) );
  IV U42404 ( .A(n13872), .Z(n39028) );
  XOR U42405 ( .A(n39031), .B(n39032), .Z(n13872) );
  XNOR U42406 ( .A(n13868), .B(n13870), .Z(n39032) );
  XNOR U42407 ( .A(q[8]), .B(DB[3503]), .Z(n13870) );
  XNOR U42408 ( .A(q[11]), .B(DB[3506]), .Z(n13868) );
  IV U42409 ( .A(n13867), .Z(n39031) );
  XNOR U42410 ( .A(n13865), .B(n39033), .Z(n13867) );
  XNOR U42411 ( .A(q[10]), .B(DB[3505]), .Z(n39033) );
  XNOR U42412 ( .A(q[9]), .B(DB[3504]), .Z(n13865) );
  IV U42413 ( .A(n13880), .Z(n39027) );
  XOR U42414 ( .A(n39034), .B(n39035), .Z(n13880) );
  XNOR U42415 ( .A(n13897), .B(n13878), .Z(n39035) );
  XNOR U42416 ( .A(q[0]), .B(DB[3495]), .Z(n13878) );
  XOR U42417 ( .A(n39036), .B(n13886), .Z(n13897) );
  XNOR U42418 ( .A(q[7]), .B(DB[3502]), .Z(n13886) );
  IV U42419 ( .A(n13885), .Z(n39036) );
  XNOR U42420 ( .A(n13883), .B(n39037), .Z(n13885) );
  XNOR U42421 ( .A(q[6]), .B(DB[3501]), .Z(n39037) );
  XNOR U42422 ( .A(q[5]), .B(DB[3500]), .Z(n13883) );
  IV U42423 ( .A(n13896), .Z(n39034) );
  XOR U42424 ( .A(n39038), .B(n39039), .Z(n13896) );
  XNOR U42425 ( .A(n13892), .B(n13894), .Z(n39039) );
  XNOR U42426 ( .A(q[1]), .B(DB[3496]), .Z(n13894) );
  XNOR U42427 ( .A(q[4]), .B(DB[3499]), .Z(n13892) );
  IV U42428 ( .A(n13891), .Z(n39038) );
  XNOR U42429 ( .A(n13889), .B(n39040), .Z(n13891) );
  XNOR U42430 ( .A(q[3]), .B(DB[3498]), .Z(n39040) );
  XNOR U42431 ( .A(q[2]), .B(DB[3497]), .Z(n13889) );
  XOR U42432 ( .A(n39041), .B(n13787), .Z(n13715) );
  XOR U42433 ( .A(n39042), .B(n13779), .Z(n13787) );
  XOR U42434 ( .A(n39043), .B(n13768), .Z(n13779) );
  XNOR U42435 ( .A(q[14]), .B(DB[3524]), .Z(n13768) );
  IV U42436 ( .A(n13767), .Z(n39043) );
  XNOR U42437 ( .A(n13765), .B(n39044), .Z(n13767) );
  XNOR U42438 ( .A(q[13]), .B(DB[3523]), .Z(n39044) );
  XNOR U42439 ( .A(q[12]), .B(DB[3522]), .Z(n13765) );
  IV U42440 ( .A(n13778), .Z(n39042) );
  XOR U42441 ( .A(n39045), .B(n39046), .Z(n13778) );
  XNOR U42442 ( .A(n13774), .B(n13776), .Z(n39046) );
  XNOR U42443 ( .A(q[8]), .B(DB[3518]), .Z(n13776) );
  XNOR U42444 ( .A(q[11]), .B(DB[3521]), .Z(n13774) );
  IV U42445 ( .A(n13773), .Z(n39045) );
  XNOR U42446 ( .A(n13771), .B(n39047), .Z(n13773) );
  XNOR U42447 ( .A(q[10]), .B(DB[3520]), .Z(n39047) );
  XNOR U42448 ( .A(q[9]), .B(DB[3519]), .Z(n13771) );
  IV U42449 ( .A(n13786), .Z(n39041) );
  XOR U42450 ( .A(n39048), .B(n39049), .Z(n13786) );
  XNOR U42451 ( .A(n13803), .B(n13784), .Z(n39049) );
  XNOR U42452 ( .A(q[0]), .B(DB[3510]), .Z(n13784) );
  XOR U42453 ( .A(n39050), .B(n13792), .Z(n13803) );
  XNOR U42454 ( .A(q[7]), .B(DB[3517]), .Z(n13792) );
  IV U42455 ( .A(n13791), .Z(n39050) );
  XNOR U42456 ( .A(n13789), .B(n39051), .Z(n13791) );
  XNOR U42457 ( .A(q[6]), .B(DB[3516]), .Z(n39051) );
  XNOR U42458 ( .A(q[5]), .B(DB[3515]), .Z(n13789) );
  IV U42459 ( .A(n13802), .Z(n39048) );
  XOR U42460 ( .A(n39052), .B(n39053), .Z(n13802) );
  XNOR U42461 ( .A(n13798), .B(n13800), .Z(n39053) );
  XNOR U42462 ( .A(q[1]), .B(DB[3511]), .Z(n13800) );
  XNOR U42463 ( .A(q[4]), .B(DB[3514]), .Z(n13798) );
  IV U42464 ( .A(n13797), .Z(n39052) );
  XNOR U42465 ( .A(n13795), .B(n39054), .Z(n13797) );
  XNOR U42466 ( .A(q[3]), .B(DB[3513]), .Z(n39054) );
  XNOR U42467 ( .A(q[2]), .B(DB[3512]), .Z(n13795) );
  XOR U42468 ( .A(n39055), .B(n13693), .Z(n13621) );
  XOR U42469 ( .A(n39056), .B(n13685), .Z(n13693) );
  XOR U42470 ( .A(n39057), .B(n13674), .Z(n13685) );
  XNOR U42471 ( .A(q[14]), .B(DB[3539]), .Z(n13674) );
  IV U42472 ( .A(n13673), .Z(n39057) );
  XNOR U42473 ( .A(n13671), .B(n39058), .Z(n13673) );
  XNOR U42474 ( .A(q[13]), .B(DB[3538]), .Z(n39058) );
  XNOR U42475 ( .A(q[12]), .B(DB[3537]), .Z(n13671) );
  IV U42476 ( .A(n13684), .Z(n39056) );
  XOR U42477 ( .A(n39059), .B(n39060), .Z(n13684) );
  XNOR U42478 ( .A(n13680), .B(n13682), .Z(n39060) );
  XNOR U42479 ( .A(q[8]), .B(DB[3533]), .Z(n13682) );
  XNOR U42480 ( .A(q[11]), .B(DB[3536]), .Z(n13680) );
  IV U42481 ( .A(n13679), .Z(n39059) );
  XNOR U42482 ( .A(n13677), .B(n39061), .Z(n13679) );
  XNOR U42483 ( .A(q[10]), .B(DB[3535]), .Z(n39061) );
  XNOR U42484 ( .A(q[9]), .B(DB[3534]), .Z(n13677) );
  IV U42485 ( .A(n13692), .Z(n39055) );
  XOR U42486 ( .A(n39062), .B(n39063), .Z(n13692) );
  XNOR U42487 ( .A(n13709), .B(n13690), .Z(n39063) );
  XNOR U42488 ( .A(q[0]), .B(DB[3525]), .Z(n13690) );
  XOR U42489 ( .A(n39064), .B(n13698), .Z(n13709) );
  XNOR U42490 ( .A(q[7]), .B(DB[3532]), .Z(n13698) );
  IV U42491 ( .A(n13697), .Z(n39064) );
  XNOR U42492 ( .A(n13695), .B(n39065), .Z(n13697) );
  XNOR U42493 ( .A(q[6]), .B(DB[3531]), .Z(n39065) );
  XNOR U42494 ( .A(q[5]), .B(DB[3530]), .Z(n13695) );
  IV U42495 ( .A(n13708), .Z(n39062) );
  XOR U42496 ( .A(n39066), .B(n39067), .Z(n13708) );
  XNOR U42497 ( .A(n13704), .B(n13706), .Z(n39067) );
  XNOR U42498 ( .A(q[1]), .B(DB[3526]), .Z(n13706) );
  XNOR U42499 ( .A(q[4]), .B(DB[3529]), .Z(n13704) );
  IV U42500 ( .A(n13703), .Z(n39066) );
  XNOR U42501 ( .A(n13701), .B(n39068), .Z(n13703) );
  XNOR U42502 ( .A(q[3]), .B(DB[3528]), .Z(n39068) );
  XNOR U42503 ( .A(q[2]), .B(DB[3527]), .Z(n13701) );
  XOR U42504 ( .A(n39069), .B(n13599), .Z(n13527) );
  XOR U42505 ( .A(n39070), .B(n13591), .Z(n13599) );
  XOR U42506 ( .A(n39071), .B(n13580), .Z(n13591) );
  XNOR U42507 ( .A(q[14]), .B(DB[3554]), .Z(n13580) );
  IV U42508 ( .A(n13579), .Z(n39071) );
  XNOR U42509 ( .A(n13577), .B(n39072), .Z(n13579) );
  XNOR U42510 ( .A(q[13]), .B(DB[3553]), .Z(n39072) );
  XNOR U42511 ( .A(q[12]), .B(DB[3552]), .Z(n13577) );
  IV U42512 ( .A(n13590), .Z(n39070) );
  XOR U42513 ( .A(n39073), .B(n39074), .Z(n13590) );
  XNOR U42514 ( .A(n13586), .B(n13588), .Z(n39074) );
  XNOR U42515 ( .A(q[8]), .B(DB[3548]), .Z(n13588) );
  XNOR U42516 ( .A(q[11]), .B(DB[3551]), .Z(n13586) );
  IV U42517 ( .A(n13585), .Z(n39073) );
  XNOR U42518 ( .A(n13583), .B(n39075), .Z(n13585) );
  XNOR U42519 ( .A(q[10]), .B(DB[3550]), .Z(n39075) );
  XNOR U42520 ( .A(q[9]), .B(DB[3549]), .Z(n13583) );
  IV U42521 ( .A(n13598), .Z(n39069) );
  XOR U42522 ( .A(n39076), .B(n39077), .Z(n13598) );
  XNOR U42523 ( .A(n13615), .B(n13596), .Z(n39077) );
  XNOR U42524 ( .A(q[0]), .B(DB[3540]), .Z(n13596) );
  XOR U42525 ( .A(n39078), .B(n13604), .Z(n13615) );
  XNOR U42526 ( .A(q[7]), .B(DB[3547]), .Z(n13604) );
  IV U42527 ( .A(n13603), .Z(n39078) );
  XNOR U42528 ( .A(n13601), .B(n39079), .Z(n13603) );
  XNOR U42529 ( .A(q[6]), .B(DB[3546]), .Z(n39079) );
  XNOR U42530 ( .A(q[5]), .B(DB[3545]), .Z(n13601) );
  IV U42531 ( .A(n13614), .Z(n39076) );
  XOR U42532 ( .A(n39080), .B(n39081), .Z(n13614) );
  XNOR U42533 ( .A(n13610), .B(n13612), .Z(n39081) );
  XNOR U42534 ( .A(q[1]), .B(DB[3541]), .Z(n13612) );
  XNOR U42535 ( .A(q[4]), .B(DB[3544]), .Z(n13610) );
  IV U42536 ( .A(n13609), .Z(n39080) );
  XNOR U42537 ( .A(n13607), .B(n39082), .Z(n13609) );
  XNOR U42538 ( .A(q[3]), .B(DB[3543]), .Z(n39082) );
  XNOR U42539 ( .A(q[2]), .B(DB[3542]), .Z(n13607) );
  XOR U42540 ( .A(n39083), .B(n13505), .Z(n13433) );
  XOR U42541 ( .A(n39084), .B(n13497), .Z(n13505) );
  XOR U42542 ( .A(n39085), .B(n13486), .Z(n13497) );
  XNOR U42543 ( .A(q[14]), .B(DB[3569]), .Z(n13486) );
  IV U42544 ( .A(n13485), .Z(n39085) );
  XNOR U42545 ( .A(n13483), .B(n39086), .Z(n13485) );
  XNOR U42546 ( .A(q[13]), .B(DB[3568]), .Z(n39086) );
  XNOR U42547 ( .A(q[12]), .B(DB[3567]), .Z(n13483) );
  IV U42548 ( .A(n13496), .Z(n39084) );
  XOR U42549 ( .A(n39087), .B(n39088), .Z(n13496) );
  XNOR U42550 ( .A(n13492), .B(n13494), .Z(n39088) );
  XNOR U42551 ( .A(q[8]), .B(DB[3563]), .Z(n13494) );
  XNOR U42552 ( .A(q[11]), .B(DB[3566]), .Z(n13492) );
  IV U42553 ( .A(n13491), .Z(n39087) );
  XNOR U42554 ( .A(n13489), .B(n39089), .Z(n13491) );
  XNOR U42555 ( .A(q[10]), .B(DB[3565]), .Z(n39089) );
  XNOR U42556 ( .A(q[9]), .B(DB[3564]), .Z(n13489) );
  IV U42557 ( .A(n13504), .Z(n39083) );
  XOR U42558 ( .A(n39090), .B(n39091), .Z(n13504) );
  XNOR U42559 ( .A(n13521), .B(n13502), .Z(n39091) );
  XNOR U42560 ( .A(q[0]), .B(DB[3555]), .Z(n13502) );
  XOR U42561 ( .A(n39092), .B(n13510), .Z(n13521) );
  XNOR U42562 ( .A(q[7]), .B(DB[3562]), .Z(n13510) );
  IV U42563 ( .A(n13509), .Z(n39092) );
  XNOR U42564 ( .A(n13507), .B(n39093), .Z(n13509) );
  XNOR U42565 ( .A(q[6]), .B(DB[3561]), .Z(n39093) );
  XNOR U42566 ( .A(q[5]), .B(DB[3560]), .Z(n13507) );
  IV U42567 ( .A(n13520), .Z(n39090) );
  XOR U42568 ( .A(n39094), .B(n39095), .Z(n13520) );
  XNOR U42569 ( .A(n13516), .B(n13518), .Z(n39095) );
  XNOR U42570 ( .A(q[1]), .B(DB[3556]), .Z(n13518) );
  XNOR U42571 ( .A(q[4]), .B(DB[3559]), .Z(n13516) );
  IV U42572 ( .A(n13515), .Z(n39094) );
  XNOR U42573 ( .A(n13513), .B(n39096), .Z(n13515) );
  XNOR U42574 ( .A(q[3]), .B(DB[3558]), .Z(n39096) );
  XNOR U42575 ( .A(q[2]), .B(DB[3557]), .Z(n13513) );
  XOR U42576 ( .A(n39097), .B(n13411), .Z(n13339) );
  XOR U42577 ( .A(n39098), .B(n13403), .Z(n13411) );
  XOR U42578 ( .A(n39099), .B(n13392), .Z(n13403) );
  XNOR U42579 ( .A(q[14]), .B(DB[3584]), .Z(n13392) );
  IV U42580 ( .A(n13391), .Z(n39099) );
  XNOR U42581 ( .A(n13389), .B(n39100), .Z(n13391) );
  XNOR U42582 ( .A(q[13]), .B(DB[3583]), .Z(n39100) );
  XNOR U42583 ( .A(q[12]), .B(DB[3582]), .Z(n13389) );
  IV U42584 ( .A(n13402), .Z(n39098) );
  XOR U42585 ( .A(n39101), .B(n39102), .Z(n13402) );
  XNOR U42586 ( .A(n13398), .B(n13400), .Z(n39102) );
  XNOR U42587 ( .A(q[8]), .B(DB[3578]), .Z(n13400) );
  XNOR U42588 ( .A(q[11]), .B(DB[3581]), .Z(n13398) );
  IV U42589 ( .A(n13397), .Z(n39101) );
  XNOR U42590 ( .A(n13395), .B(n39103), .Z(n13397) );
  XNOR U42591 ( .A(q[10]), .B(DB[3580]), .Z(n39103) );
  XNOR U42592 ( .A(q[9]), .B(DB[3579]), .Z(n13395) );
  IV U42593 ( .A(n13410), .Z(n39097) );
  XOR U42594 ( .A(n39104), .B(n39105), .Z(n13410) );
  XNOR U42595 ( .A(n13427), .B(n13408), .Z(n39105) );
  XNOR U42596 ( .A(q[0]), .B(DB[3570]), .Z(n13408) );
  XOR U42597 ( .A(n39106), .B(n13416), .Z(n13427) );
  XNOR U42598 ( .A(q[7]), .B(DB[3577]), .Z(n13416) );
  IV U42599 ( .A(n13415), .Z(n39106) );
  XNOR U42600 ( .A(n13413), .B(n39107), .Z(n13415) );
  XNOR U42601 ( .A(q[6]), .B(DB[3576]), .Z(n39107) );
  XNOR U42602 ( .A(q[5]), .B(DB[3575]), .Z(n13413) );
  IV U42603 ( .A(n13426), .Z(n39104) );
  XOR U42604 ( .A(n39108), .B(n39109), .Z(n13426) );
  XNOR U42605 ( .A(n13422), .B(n13424), .Z(n39109) );
  XNOR U42606 ( .A(q[1]), .B(DB[3571]), .Z(n13424) );
  XNOR U42607 ( .A(q[4]), .B(DB[3574]), .Z(n13422) );
  IV U42608 ( .A(n13421), .Z(n39108) );
  XNOR U42609 ( .A(n13419), .B(n39110), .Z(n13421) );
  XNOR U42610 ( .A(q[3]), .B(DB[3573]), .Z(n39110) );
  XNOR U42611 ( .A(q[2]), .B(DB[3572]), .Z(n13419) );
  XOR U42612 ( .A(n39111), .B(n13317), .Z(n13245) );
  XOR U42613 ( .A(n39112), .B(n13309), .Z(n13317) );
  XOR U42614 ( .A(n39113), .B(n13298), .Z(n13309) );
  XNOR U42615 ( .A(q[14]), .B(DB[3599]), .Z(n13298) );
  IV U42616 ( .A(n13297), .Z(n39113) );
  XNOR U42617 ( .A(n13295), .B(n39114), .Z(n13297) );
  XNOR U42618 ( .A(q[13]), .B(DB[3598]), .Z(n39114) );
  XNOR U42619 ( .A(q[12]), .B(DB[3597]), .Z(n13295) );
  IV U42620 ( .A(n13308), .Z(n39112) );
  XOR U42621 ( .A(n39115), .B(n39116), .Z(n13308) );
  XNOR U42622 ( .A(n13304), .B(n13306), .Z(n39116) );
  XNOR U42623 ( .A(q[8]), .B(DB[3593]), .Z(n13306) );
  XNOR U42624 ( .A(q[11]), .B(DB[3596]), .Z(n13304) );
  IV U42625 ( .A(n13303), .Z(n39115) );
  XNOR U42626 ( .A(n13301), .B(n39117), .Z(n13303) );
  XNOR U42627 ( .A(q[10]), .B(DB[3595]), .Z(n39117) );
  XNOR U42628 ( .A(q[9]), .B(DB[3594]), .Z(n13301) );
  IV U42629 ( .A(n13316), .Z(n39111) );
  XOR U42630 ( .A(n39118), .B(n39119), .Z(n13316) );
  XNOR U42631 ( .A(n13333), .B(n13314), .Z(n39119) );
  XNOR U42632 ( .A(q[0]), .B(DB[3585]), .Z(n13314) );
  XOR U42633 ( .A(n39120), .B(n13322), .Z(n13333) );
  XNOR U42634 ( .A(q[7]), .B(DB[3592]), .Z(n13322) );
  IV U42635 ( .A(n13321), .Z(n39120) );
  XNOR U42636 ( .A(n13319), .B(n39121), .Z(n13321) );
  XNOR U42637 ( .A(q[6]), .B(DB[3591]), .Z(n39121) );
  XNOR U42638 ( .A(q[5]), .B(DB[3590]), .Z(n13319) );
  IV U42639 ( .A(n13332), .Z(n39118) );
  XOR U42640 ( .A(n39122), .B(n39123), .Z(n13332) );
  XNOR U42641 ( .A(n13328), .B(n13330), .Z(n39123) );
  XNOR U42642 ( .A(q[1]), .B(DB[3586]), .Z(n13330) );
  XNOR U42643 ( .A(q[4]), .B(DB[3589]), .Z(n13328) );
  IV U42644 ( .A(n13327), .Z(n39122) );
  XNOR U42645 ( .A(n13325), .B(n39124), .Z(n13327) );
  XNOR U42646 ( .A(q[3]), .B(DB[3588]), .Z(n39124) );
  XNOR U42647 ( .A(q[2]), .B(DB[3587]), .Z(n13325) );
  XOR U42648 ( .A(n39125), .B(n13223), .Z(n13151) );
  XOR U42649 ( .A(n39126), .B(n13215), .Z(n13223) );
  XOR U42650 ( .A(n39127), .B(n13204), .Z(n13215) );
  XNOR U42651 ( .A(q[14]), .B(DB[3614]), .Z(n13204) );
  IV U42652 ( .A(n13203), .Z(n39127) );
  XNOR U42653 ( .A(n13201), .B(n39128), .Z(n13203) );
  XNOR U42654 ( .A(q[13]), .B(DB[3613]), .Z(n39128) );
  XNOR U42655 ( .A(q[12]), .B(DB[3612]), .Z(n13201) );
  IV U42656 ( .A(n13214), .Z(n39126) );
  XOR U42657 ( .A(n39129), .B(n39130), .Z(n13214) );
  XNOR U42658 ( .A(n13210), .B(n13212), .Z(n39130) );
  XNOR U42659 ( .A(q[8]), .B(DB[3608]), .Z(n13212) );
  XNOR U42660 ( .A(q[11]), .B(DB[3611]), .Z(n13210) );
  IV U42661 ( .A(n13209), .Z(n39129) );
  XNOR U42662 ( .A(n13207), .B(n39131), .Z(n13209) );
  XNOR U42663 ( .A(q[10]), .B(DB[3610]), .Z(n39131) );
  XNOR U42664 ( .A(q[9]), .B(DB[3609]), .Z(n13207) );
  IV U42665 ( .A(n13222), .Z(n39125) );
  XOR U42666 ( .A(n39132), .B(n39133), .Z(n13222) );
  XNOR U42667 ( .A(n13239), .B(n13220), .Z(n39133) );
  XNOR U42668 ( .A(q[0]), .B(DB[3600]), .Z(n13220) );
  XOR U42669 ( .A(n39134), .B(n13228), .Z(n13239) );
  XNOR U42670 ( .A(q[7]), .B(DB[3607]), .Z(n13228) );
  IV U42671 ( .A(n13227), .Z(n39134) );
  XNOR U42672 ( .A(n13225), .B(n39135), .Z(n13227) );
  XNOR U42673 ( .A(q[6]), .B(DB[3606]), .Z(n39135) );
  XNOR U42674 ( .A(q[5]), .B(DB[3605]), .Z(n13225) );
  IV U42675 ( .A(n13238), .Z(n39132) );
  XOR U42676 ( .A(n39136), .B(n39137), .Z(n13238) );
  XNOR U42677 ( .A(n13234), .B(n13236), .Z(n39137) );
  XNOR U42678 ( .A(q[1]), .B(DB[3601]), .Z(n13236) );
  XNOR U42679 ( .A(q[4]), .B(DB[3604]), .Z(n13234) );
  IV U42680 ( .A(n13233), .Z(n39136) );
  XNOR U42681 ( .A(n13231), .B(n39138), .Z(n13233) );
  XNOR U42682 ( .A(q[3]), .B(DB[3603]), .Z(n39138) );
  XNOR U42683 ( .A(q[2]), .B(DB[3602]), .Z(n13231) );
  XOR U42684 ( .A(n39139), .B(n13129), .Z(n13057) );
  XOR U42685 ( .A(n39140), .B(n13121), .Z(n13129) );
  XOR U42686 ( .A(n39141), .B(n13110), .Z(n13121) );
  XNOR U42687 ( .A(q[14]), .B(DB[3629]), .Z(n13110) );
  IV U42688 ( .A(n13109), .Z(n39141) );
  XNOR U42689 ( .A(n13107), .B(n39142), .Z(n13109) );
  XNOR U42690 ( .A(q[13]), .B(DB[3628]), .Z(n39142) );
  XNOR U42691 ( .A(q[12]), .B(DB[3627]), .Z(n13107) );
  IV U42692 ( .A(n13120), .Z(n39140) );
  XOR U42693 ( .A(n39143), .B(n39144), .Z(n13120) );
  XNOR U42694 ( .A(n13116), .B(n13118), .Z(n39144) );
  XNOR U42695 ( .A(q[8]), .B(DB[3623]), .Z(n13118) );
  XNOR U42696 ( .A(q[11]), .B(DB[3626]), .Z(n13116) );
  IV U42697 ( .A(n13115), .Z(n39143) );
  XNOR U42698 ( .A(n13113), .B(n39145), .Z(n13115) );
  XNOR U42699 ( .A(q[10]), .B(DB[3625]), .Z(n39145) );
  XNOR U42700 ( .A(q[9]), .B(DB[3624]), .Z(n13113) );
  IV U42701 ( .A(n13128), .Z(n39139) );
  XOR U42702 ( .A(n39146), .B(n39147), .Z(n13128) );
  XNOR U42703 ( .A(n13145), .B(n13126), .Z(n39147) );
  XNOR U42704 ( .A(q[0]), .B(DB[3615]), .Z(n13126) );
  XOR U42705 ( .A(n39148), .B(n13134), .Z(n13145) );
  XNOR U42706 ( .A(q[7]), .B(DB[3622]), .Z(n13134) );
  IV U42707 ( .A(n13133), .Z(n39148) );
  XNOR U42708 ( .A(n13131), .B(n39149), .Z(n13133) );
  XNOR U42709 ( .A(q[6]), .B(DB[3621]), .Z(n39149) );
  XNOR U42710 ( .A(q[5]), .B(DB[3620]), .Z(n13131) );
  IV U42711 ( .A(n13144), .Z(n39146) );
  XOR U42712 ( .A(n39150), .B(n39151), .Z(n13144) );
  XNOR U42713 ( .A(n13140), .B(n13142), .Z(n39151) );
  XNOR U42714 ( .A(q[1]), .B(DB[3616]), .Z(n13142) );
  XNOR U42715 ( .A(q[4]), .B(DB[3619]), .Z(n13140) );
  IV U42716 ( .A(n13139), .Z(n39150) );
  XNOR U42717 ( .A(n13137), .B(n39152), .Z(n13139) );
  XNOR U42718 ( .A(q[3]), .B(DB[3618]), .Z(n39152) );
  XNOR U42719 ( .A(q[2]), .B(DB[3617]), .Z(n13137) );
  XOR U42720 ( .A(n39153), .B(n13035), .Z(n12963) );
  XOR U42721 ( .A(n39154), .B(n13027), .Z(n13035) );
  XOR U42722 ( .A(n39155), .B(n13016), .Z(n13027) );
  XNOR U42723 ( .A(q[14]), .B(DB[3644]), .Z(n13016) );
  IV U42724 ( .A(n13015), .Z(n39155) );
  XNOR U42725 ( .A(n13013), .B(n39156), .Z(n13015) );
  XNOR U42726 ( .A(q[13]), .B(DB[3643]), .Z(n39156) );
  XNOR U42727 ( .A(q[12]), .B(DB[3642]), .Z(n13013) );
  IV U42728 ( .A(n13026), .Z(n39154) );
  XOR U42729 ( .A(n39157), .B(n39158), .Z(n13026) );
  XNOR U42730 ( .A(n13022), .B(n13024), .Z(n39158) );
  XNOR U42731 ( .A(q[8]), .B(DB[3638]), .Z(n13024) );
  XNOR U42732 ( .A(q[11]), .B(DB[3641]), .Z(n13022) );
  IV U42733 ( .A(n13021), .Z(n39157) );
  XNOR U42734 ( .A(n13019), .B(n39159), .Z(n13021) );
  XNOR U42735 ( .A(q[10]), .B(DB[3640]), .Z(n39159) );
  XNOR U42736 ( .A(q[9]), .B(DB[3639]), .Z(n13019) );
  IV U42737 ( .A(n13034), .Z(n39153) );
  XOR U42738 ( .A(n39160), .B(n39161), .Z(n13034) );
  XNOR U42739 ( .A(n13051), .B(n13032), .Z(n39161) );
  XNOR U42740 ( .A(q[0]), .B(DB[3630]), .Z(n13032) );
  XOR U42741 ( .A(n39162), .B(n13040), .Z(n13051) );
  XNOR U42742 ( .A(q[7]), .B(DB[3637]), .Z(n13040) );
  IV U42743 ( .A(n13039), .Z(n39162) );
  XNOR U42744 ( .A(n13037), .B(n39163), .Z(n13039) );
  XNOR U42745 ( .A(q[6]), .B(DB[3636]), .Z(n39163) );
  XNOR U42746 ( .A(q[5]), .B(DB[3635]), .Z(n13037) );
  IV U42747 ( .A(n13050), .Z(n39160) );
  XOR U42748 ( .A(n39164), .B(n39165), .Z(n13050) );
  XNOR U42749 ( .A(n13046), .B(n13048), .Z(n39165) );
  XNOR U42750 ( .A(q[1]), .B(DB[3631]), .Z(n13048) );
  XNOR U42751 ( .A(q[4]), .B(DB[3634]), .Z(n13046) );
  IV U42752 ( .A(n13045), .Z(n39164) );
  XNOR U42753 ( .A(n13043), .B(n39166), .Z(n13045) );
  XNOR U42754 ( .A(q[3]), .B(DB[3633]), .Z(n39166) );
  XNOR U42755 ( .A(q[2]), .B(DB[3632]), .Z(n13043) );
  XOR U42756 ( .A(n39167), .B(n12941), .Z(n12869) );
  XOR U42757 ( .A(n39168), .B(n12933), .Z(n12941) );
  XOR U42758 ( .A(n39169), .B(n12922), .Z(n12933) );
  XNOR U42759 ( .A(q[14]), .B(DB[3659]), .Z(n12922) );
  IV U42760 ( .A(n12921), .Z(n39169) );
  XNOR U42761 ( .A(n12919), .B(n39170), .Z(n12921) );
  XNOR U42762 ( .A(q[13]), .B(DB[3658]), .Z(n39170) );
  XNOR U42763 ( .A(q[12]), .B(DB[3657]), .Z(n12919) );
  IV U42764 ( .A(n12932), .Z(n39168) );
  XOR U42765 ( .A(n39171), .B(n39172), .Z(n12932) );
  XNOR U42766 ( .A(n12928), .B(n12930), .Z(n39172) );
  XNOR U42767 ( .A(q[8]), .B(DB[3653]), .Z(n12930) );
  XNOR U42768 ( .A(q[11]), .B(DB[3656]), .Z(n12928) );
  IV U42769 ( .A(n12927), .Z(n39171) );
  XNOR U42770 ( .A(n12925), .B(n39173), .Z(n12927) );
  XNOR U42771 ( .A(q[10]), .B(DB[3655]), .Z(n39173) );
  XNOR U42772 ( .A(q[9]), .B(DB[3654]), .Z(n12925) );
  IV U42773 ( .A(n12940), .Z(n39167) );
  XOR U42774 ( .A(n39174), .B(n39175), .Z(n12940) );
  XNOR U42775 ( .A(n12957), .B(n12938), .Z(n39175) );
  XNOR U42776 ( .A(q[0]), .B(DB[3645]), .Z(n12938) );
  XOR U42777 ( .A(n39176), .B(n12946), .Z(n12957) );
  XNOR U42778 ( .A(q[7]), .B(DB[3652]), .Z(n12946) );
  IV U42779 ( .A(n12945), .Z(n39176) );
  XNOR U42780 ( .A(n12943), .B(n39177), .Z(n12945) );
  XNOR U42781 ( .A(q[6]), .B(DB[3651]), .Z(n39177) );
  XNOR U42782 ( .A(q[5]), .B(DB[3650]), .Z(n12943) );
  IV U42783 ( .A(n12956), .Z(n39174) );
  XOR U42784 ( .A(n39178), .B(n39179), .Z(n12956) );
  XNOR U42785 ( .A(n12952), .B(n12954), .Z(n39179) );
  XNOR U42786 ( .A(q[1]), .B(DB[3646]), .Z(n12954) );
  XNOR U42787 ( .A(q[4]), .B(DB[3649]), .Z(n12952) );
  IV U42788 ( .A(n12951), .Z(n39178) );
  XNOR U42789 ( .A(n12949), .B(n39180), .Z(n12951) );
  XNOR U42790 ( .A(q[3]), .B(DB[3648]), .Z(n39180) );
  XNOR U42791 ( .A(q[2]), .B(DB[3647]), .Z(n12949) );
  XOR U42792 ( .A(n39181), .B(n12847), .Z(n12775) );
  XOR U42793 ( .A(n39182), .B(n12839), .Z(n12847) );
  XOR U42794 ( .A(n39183), .B(n12828), .Z(n12839) );
  XNOR U42795 ( .A(q[14]), .B(DB[3674]), .Z(n12828) );
  IV U42796 ( .A(n12827), .Z(n39183) );
  XNOR U42797 ( .A(n12825), .B(n39184), .Z(n12827) );
  XNOR U42798 ( .A(q[13]), .B(DB[3673]), .Z(n39184) );
  XNOR U42799 ( .A(q[12]), .B(DB[3672]), .Z(n12825) );
  IV U42800 ( .A(n12838), .Z(n39182) );
  XOR U42801 ( .A(n39185), .B(n39186), .Z(n12838) );
  XNOR U42802 ( .A(n12834), .B(n12836), .Z(n39186) );
  XNOR U42803 ( .A(q[8]), .B(DB[3668]), .Z(n12836) );
  XNOR U42804 ( .A(q[11]), .B(DB[3671]), .Z(n12834) );
  IV U42805 ( .A(n12833), .Z(n39185) );
  XNOR U42806 ( .A(n12831), .B(n39187), .Z(n12833) );
  XNOR U42807 ( .A(q[10]), .B(DB[3670]), .Z(n39187) );
  XNOR U42808 ( .A(q[9]), .B(DB[3669]), .Z(n12831) );
  IV U42809 ( .A(n12846), .Z(n39181) );
  XOR U42810 ( .A(n39188), .B(n39189), .Z(n12846) );
  XNOR U42811 ( .A(n12863), .B(n12844), .Z(n39189) );
  XNOR U42812 ( .A(q[0]), .B(DB[3660]), .Z(n12844) );
  XOR U42813 ( .A(n39190), .B(n12852), .Z(n12863) );
  XNOR U42814 ( .A(q[7]), .B(DB[3667]), .Z(n12852) );
  IV U42815 ( .A(n12851), .Z(n39190) );
  XNOR U42816 ( .A(n12849), .B(n39191), .Z(n12851) );
  XNOR U42817 ( .A(q[6]), .B(DB[3666]), .Z(n39191) );
  XNOR U42818 ( .A(q[5]), .B(DB[3665]), .Z(n12849) );
  IV U42819 ( .A(n12862), .Z(n39188) );
  XOR U42820 ( .A(n39192), .B(n39193), .Z(n12862) );
  XNOR U42821 ( .A(n12858), .B(n12860), .Z(n39193) );
  XNOR U42822 ( .A(q[1]), .B(DB[3661]), .Z(n12860) );
  XNOR U42823 ( .A(q[4]), .B(DB[3664]), .Z(n12858) );
  IV U42824 ( .A(n12857), .Z(n39192) );
  XNOR U42825 ( .A(n12855), .B(n39194), .Z(n12857) );
  XNOR U42826 ( .A(q[3]), .B(DB[3663]), .Z(n39194) );
  XNOR U42827 ( .A(q[2]), .B(DB[3662]), .Z(n12855) );
  XOR U42828 ( .A(n39195), .B(n12753), .Z(n12681) );
  XOR U42829 ( .A(n39196), .B(n12745), .Z(n12753) );
  XOR U42830 ( .A(n39197), .B(n12734), .Z(n12745) );
  XNOR U42831 ( .A(q[14]), .B(DB[3689]), .Z(n12734) );
  IV U42832 ( .A(n12733), .Z(n39197) );
  XNOR U42833 ( .A(n12731), .B(n39198), .Z(n12733) );
  XNOR U42834 ( .A(q[13]), .B(DB[3688]), .Z(n39198) );
  XNOR U42835 ( .A(q[12]), .B(DB[3687]), .Z(n12731) );
  IV U42836 ( .A(n12744), .Z(n39196) );
  XOR U42837 ( .A(n39199), .B(n39200), .Z(n12744) );
  XNOR U42838 ( .A(n12740), .B(n12742), .Z(n39200) );
  XNOR U42839 ( .A(q[8]), .B(DB[3683]), .Z(n12742) );
  XNOR U42840 ( .A(q[11]), .B(DB[3686]), .Z(n12740) );
  IV U42841 ( .A(n12739), .Z(n39199) );
  XNOR U42842 ( .A(n12737), .B(n39201), .Z(n12739) );
  XNOR U42843 ( .A(q[10]), .B(DB[3685]), .Z(n39201) );
  XNOR U42844 ( .A(q[9]), .B(DB[3684]), .Z(n12737) );
  IV U42845 ( .A(n12752), .Z(n39195) );
  XOR U42846 ( .A(n39202), .B(n39203), .Z(n12752) );
  XNOR U42847 ( .A(n12769), .B(n12750), .Z(n39203) );
  XNOR U42848 ( .A(q[0]), .B(DB[3675]), .Z(n12750) );
  XOR U42849 ( .A(n39204), .B(n12758), .Z(n12769) );
  XNOR U42850 ( .A(q[7]), .B(DB[3682]), .Z(n12758) );
  IV U42851 ( .A(n12757), .Z(n39204) );
  XNOR U42852 ( .A(n12755), .B(n39205), .Z(n12757) );
  XNOR U42853 ( .A(q[6]), .B(DB[3681]), .Z(n39205) );
  XNOR U42854 ( .A(q[5]), .B(DB[3680]), .Z(n12755) );
  IV U42855 ( .A(n12768), .Z(n39202) );
  XOR U42856 ( .A(n39206), .B(n39207), .Z(n12768) );
  XNOR U42857 ( .A(n12764), .B(n12766), .Z(n39207) );
  XNOR U42858 ( .A(q[1]), .B(DB[3676]), .Z(n12766) );
  XNOR U42859 ( .A(q[4]), .B(DB[3679]), .Z(n12764) );
  IV U42860 ( .A(n12763), .Z(n39206) );
  XNOR U42861 ( .A(n12761), .B(n39208), .Z(n12763) );
  XNOR U42862 ( .A(q[3]), .B(DB[3678]), .Z(n39208) );
  XNOR U42863 ( .A(q[2]), .B(DB[3677]), .Z(n12761) );
  XOR U42864 ( .A(n39209), .B(n12659), .Z(n12587) );
  XOR U42865 ( .A(n39210), .B(n12651), .Z(n12659) );
  XOR U42866 ( .A(n39211), .B(n12640), .Z(n12651) );
  XNOR U42867 ( .A(q[14]), .B(DB[3704]), .Z(n12640) );
  IV U42868 ( .A(n12639), .Z(n39211) );
  XNOR U42869 ( .A(n12637), .B(n39212), .Z(n12639) );
  XNOR U42870 ( .A(q[13]), .B(DB[3703]), .Z(n39212) );
  XNOR U42871 ( .A(q[12]), .B(DB[3702]), .Z(n12637) );
  IV U42872 ( .A(n12650), .Z(n39210) );
  XOR U42873 ( .A(n39213), .B(n39214), .Z(n12650) );
  XNOR U42874 ( .A(n12646), .B(n12648), .Z(n39214) );
  XNOR U42875 ( .A(q[8]), .B(DB[3698]), .Z(n12648) );
  XNOR U42876 ( .A(q[11]), .B(DB[3701]), .Z(n12646) );
  IV U42877 ( .A(n12645), .Z(n39213) );
  XNOR U42878 ( .A(n12643), .B(n39215), .Z(n12645) );
  XNOR U42879 ( .A(q[10]), .B(DB[3700]), .Z(n39215) );
  XNOR U42880 ( .A(q[9]), .B(DB[3699]), .Z(n12643) );
  IV U42881 ( .A(n12658), .Z(n39209) );
  XOR U42882 ( .A(n39216), .B(n39217), .Z(n12658) );
  XNOR U42883 ( .A(n12675), .B(n12656), .Z(n39217) );
  XNOR U42884 ( .A(q[0]), .B(DB[3690]), .Z(n12656) );
  XOR U42885 ( .A(n39218), .B(n12664), .Z(n12675) );
  XNOR U42886 ( .A(q[7]), .B(DB[3697]), .Z(n12664) );
  IV U42887 ( .A(n12663), .Z(n39218) );
  XNOR U42888 ( .A(n12661), .B(n39219), .Z(n12663) );
  XNOR U42889 ( .A(q[6]), .B(DB[3696]), .Z(n39219) );
  XNOR U42890 ( .A(q[5]), .B(DB[3695]), .Z(n12661) );
  IV U42891 ( .A(n12674), .Z(n39216) );
  XOR U42892 ( .A(n39220), .B(n39221), .Z(n12674) );
  XNOR U42893 ( .A(n12670), .B(n12672), .Z(n39221) );
  XNOR U42894 ( .A(q[1]), .B(DB[3691]), .Z(n12672) );
  XNOR U42895 ( .A(q[4]), .B(DB[3694]), .Z(n12670) );
  IV U42896 ( .A(n12669), .Z(n39220) );
  XNOR U42897 ( .A(n12667), .B(n39222), .Z(n12669) );
  XNOR U42898 ( .A(q[3]), .B(DB[3693]), .Z(n39222) );
  XNOR U42899 ( .A(q[2]), .B(DB[3692]), .Z(n12667) );
  XOR U42900 ( .A(n39223), .B(n12565), .Z(n12493) );
  XOR U42901 ( .A(n39224), .B(n12557), .Z(n12565) );
  XOR U42902 ( .A(n39225), .B(n12546), .Z(n12557) );
  XNOR U42903 ( .A(q[14]), .B(DB[3719]), .Z(n12546) );
  IV U42904 ( .A(n12545), .Z(n39225) );
  XNOR U42905 ( .A(n12543), .B(n39226), .Z(n12545) );
  XNOR U42906 ( .A(q[13]), .B(DB[3718]), .Z(n39226) );
  XNOR U42907 ( .A(q[12]), .B(DB[3717]), .Z(n12543) );
  IV U42908 ( .A(n12556), .Z(n39224) );
  XOR U42909 ( .A(n39227), .B(n39228), .Z(n12556) );
  XNOR U42910 ( .A(n12552), .B(n12554), .Z(n39228) );
  XNOR U42911 ( .A(q[8]), .B(DB[3713]), .Z(n12554) );
  XNOR U42912 ( .A(q[11]), .B(DB[3716]), .Z(n12552) );
  IV U42913 ( .A(n12551), .Z(n39227) );
  XNOR U42914 ( .A(n12549), .B(n39229), .Z(n12551) );
  XNOR U42915 ( .A(q[10]), .B(DB[3715]), .Z(n39229) );
  XNOR U42916 ( .A(q[9]), .B(DB[3714]), .Z(n12549) );
  IV U42917 ( .A(n12564), .Z(n39223) );
  XOR U42918 ( .A(n39230), .B(n39231), .Z(n12564) );
  XNOR U42919 ( .A(n12581), .B(n12562), .Z(n39231) );
  XNOR U42920 ( .A(q[0]), .B(DB[3705]), .Z(n12562) );
  XOR U42921 ( .A(n39232), .B(n12570), .Z(n12581) );
  XNOR U42922 ( .A(q[7]), .B(DB[3712]), .Z(n12570) );
  IV U42923 ( .A(n12569), .Z(n39232) );
  XNOR U42924 ( .A(n12567), .B(n39233), .Z(n12569) );
  XNOR U42925 ( .A(q[6]), .B(DB[3711]), .Z(n39233) );
  XNOR U42926 ( .A(q[5]), .B(DB[3710]), .Z(n12567) );
  IV U42927 ( .A(n12580), .Z(n39230) );
  XOR U42928 ( .A(n39234), .B(n39235), .Z(n12580) );
  XNOR U42929 ( .A(n12576), .B(n12578), .Z(n39235) );
  XNOR U42930 ( .A(q[1]), .B(DB[3706]), .Z(n12578) );
  XNOR U42931 ( .A(q[4]), .B(DB[3709]), .Z(n12576) );
  IV U42932 ( .A(n12575), .Z(n39234) );
  XNOR U42933 ( .A(n12573), .B(n39236), .Z(n12575) );
  XNOR U42934 ( .A(q[3]), .B(DB[3708]), .Z(n39236) );
  XNOR U42935 ( .A(q[2]), .B(DB[3707]), .Z(n12573) );
  XOR U42936 ( .A(n39237), .B(n12471), .Z(n12399) );
  XOR U42937 ( .A(n39238), .B(n12463), .Z(n12471) );
  XOR U42938 ( .A(n39239), .B(n12452), .Z(n12463) );
  XNOR U42939 ( .A(q[14]), .B(DB[3734]), .Z(n12452) );
  IV U42940 ( .A(n12451), .Z(n39239) );
  XNOR U42941 ( .A(n12449), .B(n39240), .Z(n12451) );
  XNOR U42942 ( .A(q[13]), .B(DB[3733]), .Z(n39240) );
  XNOR U42943 ( .A(q[12]), .B(DB[3732]), .Z(n12449) );
  IV U42944 ( .A(n12462), .Z(n39238) );
  XOR U42945 ( .A(n39241), .B(n39242), .Z(n12462) );
  XNOR U42946 ( .A(n12458), .B(n12460), .Z(n39242) );
  XNOR U42947 ( .A(q[8]), .B(DB[3728]), .Z(n12460) );
  XNOR U42948 ( .A(q[11]), .B(DB[3731]), .Z(n12458) );
  IV U42949 ( .A(n12457), .Z(n39241) );
  XNOR U42950 ( .A(n12455), .B(n39243), .Z(n12457) );
  XNOR U42951 ( .A(q[10]), .B(DB[3730]), .Z(n39243) );
  XNOR U42952 ( .A(q[9]), .B(DB[3729]), .Z(n12455) );
  IV U42953 ( .A(n12470), .Z(n39237) );
  XOR U42954 ( .A(n39244), .B(n39245), .Z(n12470) );
  XNOR U42955 ( .A(n12487), .B(n12468), .Z(n39245) );
  XNOR U42956 ( .A(q[0]), .B(DB[3720]), .Z(n12468) );
  XOR U42957 ( .A(n39246), .B(n12476), .Z(n12487) );
  XNOR U42958 ( .A(q[7]), .B(DB[3727]), .Z(n12476) );
  IV U42959 ( .A(n12475), .Z(n39246) );
  XNOR U42960 ( .A(n12473), .B(n39247), .Z(n12475) );
  XNOR U42961 ( .A(q[6]), .B(DB[3726]), .Z(n39247) );
  XNOR U42962 ( .A(q[5]), .B(DB[3725]), .Z(n12473) );
  IV U42963 ( .A(n12486), .Z(n39244) );
  XOR U42964 ( .A(n39248), .B(n39249), .Z(n12486) );
  XNOR U42965 ( .A(n12482), .B(n12484), .Z(n39249) );
  XNOR U42966 ( .A(q[1]), .B(DB[3721]), .Z(n12484) );
  XNOR U42967 ( .A(q[4]), .B(DB[3724]), .Z(n12482) );
  IV U42968 ( .A(n12481), .Z(n39248) );
  XNOR U42969 ( .A(n12479), .B(n39250), .Z(n12481) );
  XNOR U42970 ( .A(q[3]), .B(DB[3723]), .Z(n39250) );
  XNOR U42971 ( .A(q[2]), .B(DB[3722]), .Z(n12479) );
  XOR U42972 ( .A(n39251), .B(n12377), .Z(n12305) );
  XOR U42973 ( .A(n39252), .B(n12369), .Z(n12377) );
  XOR U42974 ( .A(n39253), .B(n12358), .Z(n12369) );
  XNOR U42975 ( .A(q[14]), .B(DB[3749]), .Z(n12358) );
  IV U42976 ( .A(n12357), .Z(n39253) );
  XNOR U42977 ( .A(n12355), .B(n39254), .Z(n12357) );
  XNOR U42978 ( .A(q[13]), .B(DB[3748]), .Z(n39254) );
  XNOR U42979 ( .A(q[12]), .B(DB[3747]), .Z(n12355) );
  IV U42980 ( .A(n12368), .Z(n39252) );
  XOR U42981 ( .A(n39255), .B(n39256), .Z(n12368) );
  XNOR U42982 ( .A(n12364), .B(n12366), .Z(n39256) );
  XNOR U42983 ( .A(q[8]), .B(DB[3743]), .Z(n12366) );
  XNOR U42984 ( .A(q[11]), .B(DB[3746]), .Z(n12364) );
  IV U42985 ( .A(n12363), .Z(n39255) );
  XNOR U42986 ( .A(n12361), .B(n39257), .Z(n12363) );
  XNOR U42987 ( .A(q[10]), .B(DB[3745]), .Z(n39257) );
  XNOR U42988 ( .A(q[9]), .B(DB[3744]), .Z(n12361) );
  IV U42989 ( .A(n12376), .Z(n39251) );
  XOR U42990 ( .A(n39258), .B(n39259), .Z(n12376) );
  XNOR U42991 ( .A(n12393), .B(n12374), .Z(n39259) );
  XNOR U42992 ( .A(q[0]), .B(DB[3735]), .Z(n12374) );
  XOR U42993 ( .A(n39260), .B(n12382), .Z(n12393) );
  XNOR U42994 ( .A(q[7]), .B(DB[3742]), .Z(n12382) );
  IV U42995 ( .A(n12381), .Z(n39260) );
  XNOR U42996 ( .A(n12379), .B(n39261), .Z(n12381) );
  XNOR U42997 ( .A(q[6]), .B(DB[3741]), .Z(n39261) );
  XNOR U42998 ( .A(q[5]), .B(DB[3740]), .Z(n12379) );
  IV U42999 ( .A(n12392), .Z(n39258) );
  XOR U43000 ( .A(n39262), .B(n39263), .Z(n12392) );
  XNOR U43001 ( .A(n12388), .B(n12390), .Z(n39263) );
  XNOR U43002 ( .A(q[1]), .B(DB[3736]), .Z(n12390) );
  XNOR U43003 ( .A(q[4]), .B(DB[3739]), .Z(n12388) );
  IV U43004 ( .A(n12387), .Z(n39262) );
  XNOR U43005 ( .A(n12385), .B(n39264), .Z(n12387) );
  XNOR U43006 ( .A(q[3]), .B(DB[3738]), .Z(n39264) );
  XNOR U43007 ( .A(q[2]), .B(DB[3737]), .Z(n12385) );
  XOR U43008 ( .A(n39265), .B(n12283), .Z(n12211) );
  XOR U43009 ( .A(n39266), .B(n12275), .Z(n12283) );
  XOR U43010 ( .A(n39267), .B(n12264), .Z(n12275) );
  XNOR U43011 ( .A(q[14]), .B(DB[3764]), .Z(n12264) );
  IV U43012 ( .A(n12263), .Z(n39267) );
  XNOR U43013 ( .A(n12261), .B(n39268), .Z(n12263) );
  XNOR U43014 ( .A(q[13]), .B(DB[3763]), .Z(n39268) );
  XNOR U43015 ( .A(q[12]), .B(DB[3762]), .Z(n12261) );
  IV U43016 ( .A(n12274), .Z(n39266) );
  XOR U43017 ( .A(n39269), .B(n39270), .Z(n12274) );
  XNOR U43018 ( .A(n12270), .B(n12272), .Z(n39270) );
  XNOR U43019 ( .A(q[8]), .B(DB[3758]), .Z(n12272) );
  XNOR U43020 ( .A(q[11]), .B(DB[3761]), .Z(n12270) );
  IV U43021 ( .A(n12269), .Z(n39269) );
  XNOR U43022 ( .A(n12267), .B(n39271), .Z(n12269) );
  XNOR U43023 ( .A(q[10]), .B(DB[3760]), .Z(n39271) );
  XNOR U43024 ( .A(q[9]), .B(DB[3759]), .Z(n12267) );
  IV U43025 ( .A(n12282), .Z(n39265) );
  XOR U43026 ( .A(n39272), .B(n39273), .Z(n12282) );
  XNOR U43027 ( .A(n12299), .B(n12280), .Z(n39273) );
  XNOR U43028 ( .A(q[0]), .B(DB[3750]), .Z(n12280) );
  XOR U43029 ( .A(n39274), .B(n12288), .Z(n12299) );
  XNOR U43030 ( .A(q[7]), .B(DB[3757]), .Z(n12288) );
  IV U43031 ( .A(n12287), .Z(n39274) );
  XNOR U43032 ( .A(n12285), .B(n39275), .Z(n12287) );
  XNOR U43033 ( .A(q[6]), .B(DB[3756]), .Z(n39275) );
  XNOR U43034 ( .A(q[5]), .B(DB[3755]), .Z(n12285) );
  IV U43035 ( .A(n12298), .Z(n39272) );
  XOR U43036 ( .A(n39276), .B(n39277), .Z(n12298) );
  XNOR U43037 ( .A(n12294), .B(n12296), .Z(n39277) );
  XNOR U43038 ( .A(q[1]), .B(DB[3751]), .Z(n12296) );
  XNOR U43039 ( .A(q[4]), .B(DB[3754]), .Z(n12294) );
  IV U43040 ( .A(n12293), .Z(n39276) );
  XNOR U43041 ( .A(n12291), .B(n39278), .Z(n12293) );
  XNOR U43042 ( .A(q[3]), .B(DB[3753]), .Z(n39278) );
  XNOR U43043 ( .A(q[2]), .B(DB[3752]), .Z(n12291) );
  XOR U43044 ( .A(n39279), .B(n12189), .Z(n12117) );
  XOR U43045 ( .A(n39280), .B(n12181), .Z(n12189) );
  XOR U43046 ( .A(n39281), .B(n12170), .Z(n12181) );
  XNOR U43047 ( .A(q[14]), .B(DB[3779]), .Z(n12170) );
  IV U43048 ( .A(n12169), .Z(n39281) );
  XNOR U43049 ( .A(n12167), .B(n39282), .Z(n12169) );
  XNOR U43050 ( .A(q[13]), .B(DB[3778]), .Z(n39282) );
  XNOR U43051 ( .A(q[12]), .B(DB[3777]), .Z(n12167) );
  IV U43052 ( .A(n12180), .Z(n39280) );
  XOR U43053 ( .A(n39283), .B(n39284), .Z(n12180) );
  XNOR U43054 ( .A(n12176), .B(n12178), .Z(n39284) );
  XNOR U43055 ( .A(q[8]), .B(DB[3773]), .Z(n12178) );
  XNOR U43056 ( .A(q[11]), .B(DB[3776]), .Z(n12176) );
  IV U43057 ( .A(n12175), .Z(n39283) );
  XNOR U43058 ( .A(n12173), .B(n39285), .Z(n12175) );
  XNOR U43059 ( .A(q[10]), .B(DB[3775]), .Z(n39285) );
  XNOR U43060 ( .A(q[9]), .B(DB[3774]), .Z(n12173) );
  IV U43061 ( .A(n12188), .Z(n39279) );
  XOR U43062 ( .A(n39286), .B(n39287), .Z(n12188) );
  XNOR U43063 ( .A(n12205), .B(n12186), .Z(n39287) );
  XNOR U43064 ( .A(q[0]), .B(DB[3765]), .Z(n12186) );
  XOR U43065 ( .A(n39288), .B(n12194), .Z(n12205) );
  XNOR U43066 ( .A(q[7]), .B(DB[3772]), .Z(n12194) );
  IV U43067 ( .A(n12193), .Z(n39288) );
  XNOR U43068 ( .A(n12191), .B(n39289), .Z(n12193) );
  XNOR U43069 ( .A(q[6]), .B(DB[3771]), .Z(n39289) );
  XNOR U43070 ( .A(q[5]), .B(DB[3770]), .Z(n12191) );
  IV U43071 ( .A(n12204), .Z(n39286) );
  XOR U43072 ( .A(n39290), .B(n39291), .Z(n12204) );
  XNOR U43073 ( .A(n12200), .B(n12202), .Z(n39291) );
  XNOR U43074 ( .A(q[1]), .B(DB[3766]), .Z(n12202) );
  XNOR U43075 ( .A(q[4]), .B(DB[3769]), .Z(n12200) );
  IV U43076 ( .A(n12199), .Z(n39290) );
  XNOR U43077 ( .A(n12197), .B(n39292), .Z(n12199) );
  XNOR U43078 ( .A(q[3]), .B(DB[3768]), .Z(n39292) );
  XNOR U43079 ( .A(q[2]), .B(DB[3767]), .Z(n12197) );
  XOR U43080 ( .A(n39293), .B(n12095), .Z(n12023) );
  XOR U43081 ( .A(n39294), .B(n12087), .Z(n12095) );
  XOR U43082 ( .A(n39295), .B(n12076), .Z(n12087) );
  XNOR U43083 ( .A(q[14]), .B(DB[3794]), .Z(n12076) );
  IV U43084 ( .A(n12075), .Z(n39295) );
  XNOR U43085 ( .A(n12073), .B(n39296), .Z(n12075) );
  XNOR U43086 ( .A(q[13]), .B(DB[3793]), .Z(n39296) );
  XNOR U43087 ( .A(q[12]), .B(DB[3792]), .Z(n12073) );
  IV U43088 ( .A(n12086), .Z(n39294) );
  XOR U43089 ( .A(n39297), .B(n39298), .Z(n12086) );
  XNOR U43090 ( .A(n12082), .B(n12084), .Z(n39298) );
  XNOR U43091 ( .A(q[8]), .B(DB[3788]), .Z(n12084) );
  XNOR U43092 ( .A(q[11]), .B(DB[3791]), .Z(n12082) );
  IV U43093 ( .A(n12081), .Z(n39297) );
  XNOR U43094 ( .A(n12079), .B(n39299), .Z(n12081) );
  XNOR U43095 ( .A(q[10]), .B(DB[3790]), .Z(n39299) );
  XNOR U43096 ( .A(q[9]), .B(DB[3789]), .Z(n12079) );
  IV U43097 ( .A(n12094), .Z(n39293) );
  XOR U43098 ( .A(n39300), .B(n39301), .Z(n12094) );
  XNOR U43099 ( .A(n12111), .B(n12092), .Z(n39301) );
  XNOR U43100 ( .A(q[0]), .B(DB[3780]), .Z(n12092) );
  XOR U43101 ( .A(n39302), .B(n12100), .Z(n12111) );
  XNOR U43102 ( .A(q[7]), .B(DB[3787]), .Z(n12100) );
  IV U43103 ( .A(n12099), .Z(n39302) );
  XNOR U43104 ( .A(n12097), .B(n39303), .Z(n12099) );
  XNOR U43105 ( .A(q[6]), .B(DB[3786]), .Z(n39303) );
  XNOR U43106 ( .A(q[5]), .B(DB[3785]), .Z(n12097) );
  IV U43107 ( .A(n12110), .Z(n39300) );
  XOR U43108 ( .A(n39304), .B(n39305), .Z(n12110) );
  XNOR U43109 ( .A(n12106), .B(n12108), .Z(n39305) );
  XNOR U43110 ( .A(q[1]), .B(DB[3781]), .Z(n12108) );
  XNOR U43111 ( .A(q[4]), .B(DB[3784]), .Z(n12106) );
  IV U43112 ( .A(n12105), .Z(n39304) );
  XNOR U43113 ( .A(n12103), .B(n39306), .Z(n12105) );
  XNOR U43114 ( .A(q[3]), .B(DB[3783]), .Z(n39306) );
  XNOR U43115 ( .A(q[2]), .B(DB[3782]), .Z(n12103) );
  XOR U43116 ( .A(n39307), .B(n12001), .Z(n11929) );
  XOR U43117 ( .A(n39308), .B(n11993), .Z(n12001) );
  XOR U43118 ( .A(n39309), .B(n11982), .Z(n11993) );
  XNOR U43119 ( .A(q[14]), .B(DB[3809]), .Z(n11982) );
  IV U43120 ( .A(n11981), .Z(n39309) );
  XNOR U43121 ( .A(n11979), .B(n39310), .Z(n11981) );
  XNOR U43122 ( .A(q[13]), .B(DB[3808]), .Z(n39310) );
  XNOR U43123 ( .A(q[12]), .B(DB[3807]), .Z(n11979) );
  IV U43124 ( .A(n11992), .Z(n39308) );
  XOR U43125 ( .A(n39311), .B(n39312), .Z(n11992) );
  XNOR U43126 ( .A(n11988), .B(n11990), .Z(n39312) );
  XNOR U43127 ( .A(q[8]), .B(DB[3803]), .Z(n11990) );
  XNOR U43128 ( .A(q[11]), .B(DB[3806]), .Z(n11988) );
  IV U43129 ( .A(n11987), .Z(n39311) );
  XNOR U43130 ( .A(n11985), .B(n39313), .Z(n11987) );
  XNOR U43131 ( .A(q[10]), .B(DB[3805]), .Z(n39313) );
  XNOR U43132 ( .A(q[9]), .B(DB[3804]), .Z(n11985) );
  IV U43133 ( .A(n12000), .Z(n39307) );
  XOR U43134 ( .A(n39314), .B(n39315), .Z(n12000) );
  XNOR U43135 ( .A(n12017), .B(n11998), .Z(n39315) );
  XNOR U43136 ( .A(q[0]), .B(DB[3795]), .Z(n11998) );
  XOR U43137 ( .A(n39316), .B(n12006), .Z(n12017) );
  XNOR U43138 ( .A(q[7]), .B(DB[3802]), .Z(n12006) );
  IV U43139 ( .A(n12005), .Z(n39316) );
  XNOR U43140 ( .A(n12003), .B(n39317), .Z(n12005) );
  XNOR U43141 ( .A(q[6]), .B(DB[3801]), .Z(n39317) );
  XNOR U43142 ( .A(q[5]), .B(DB[3800]), .Z(n12003) );
  IV U43143 ( .A(n12016), .Z(n39314) );
  XOR U43144 ( .A(n39318), .B(n39319), .Z(n12016) );
  XNOR U43145 ( .A(n12012), .B(n12014), .Z(n39319) );
  XNOR U43146 ( .A(q[1]), .B(DB[3796]), .Z(n12014) );
  XNOR U43147 ( .A(q[4]), .B(DB[3799]), .Z(n12012) );
  IV U43148 ( .A(n12011), .Z(n39318) );
  XNOR U43149 ( .A(n12009), .B(n39320), .Z(n12011) );
  XNOR U43150 ( .A(q[3]), .B(DB[3798]), .Z(n39320) );
  XNOR U43151 ( .A(q[2]), .B(DB[3797]), .Z(n12009) );
  XOR U43152 ( .A(n39321), .B(n11907), .Z(n11833) );
  XOR U43153 ( .A(n39322), .B(n11899), .Z(n11907) );
  XOR U43154 ( .A(n39323), .B(n11888), .Z(n11899) );
  XNOR U43155 ( .A(q[14]), .B(DB[3824]), .Z(n11888) );
  IV U43156 ( .A(n11887), .Z(n39323) );
  XNOR U43157 ( .A(n11885), .B(n39324), .Z(n11887) );
  XNOR U43158 ( .A(q[13]), .B(DB[3823]), .Z(n39324) );
  XOR U43159 ( .A(q[12]), .B(n8665), .Z(n11885) );
  IV U43160 ( .A(DB[3822]), .Z(n8665) );
  IV U43161 ( .A(n11898), .Z(n39322) );
  XOR U43162 ( .A(n39325), .B(n39326), .Z(n11898) );
  XNOR U43163 ( .A(n11894), .B(n11896), .Z(n39326) );
  XNOR U43164 ( .A(q[8]), .B(DB[3818]), .Z(n11896) );
  XOR U43165 ( .A(q[11]), .B(n9431), .Z(n11894) );
  IV U43166 ( .A(DB[3821]), .Z(n9431) );
  IV U43167 ( .A(n11893), .Z(n39325) );
  XNOR U43168 ( .A(n11891), .B(n39327), .Z(n11893) );
  XNOR U43169 ( .A(q[10]), .B(DB[3820]), .Z(n39327) );
  XNOR U43170 ( .A(q[9]), .B(DB[3819]), .Z(n11891) );
  IV U43171 ( .A(n11906), .Z(n39321) );
  XOR U43172 ( .A(n39328), .B(n39329), .Z(n11906) );
  XNOR U43173 ( .A(n11923), .B(n11904), .Z(n39329) );
  XNOR U43174 ( .A(q[0]), .B(DB[3810]), .Z(n11904) );
  XOR U43175 ( .A(n39330), .B(n11912), .Z(n11923) );
  XNOR U43176 ( .A(q[7]), .B(DB[3817]), .Z(n11912) );
  IV U43177 ( .A(n11911), .Z(n39330) );
  XNOR U43178 ( .A(n11909), .B(n39331), .Z(n11911) );
  XNOR U43179 ( .A(q[6]), .B(DB[3816]), .Z(n39331) );
  XNOR U43180 ( .A(q[5]), .B(DB[3815]), .Z(n11909) );
  IV U43181 ( .A(n11922), .Z(n39328) );
  XOR U43182 ( .A(n39332), .B(n39333), .Z(n11922) );
  XNOR U43183 ( .A(n11918), .B(n11920), .Z(n39333) );
  XNOR U43184 ( .A(q[1]), .B(DB[3811]), .Z(n11920) );
  XNOR U43185 ( .A(q[4]), .B(DB[3814]), .Z(n11918) );
  IV U43186 ( .A(n11917), .Z(n39332) );
  XNOR U43187 ( .A(n11915), .B(n39334), .Z(n11917) );
  XNOR U43188 ( .A(q[3]), .B(DB[3813]), .Z(n39334) );
  XNOR U43189 ( .A(q[2]), .B(DB[3812]), .Z(n11915) );
endmodule

