
module sum_N16384_CC512 ( clk, rst, a, b, c );
  input [31:0] a;
  input [31:0] b;
  output [31:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        carry_on) );
  XOR U4 ( .A(n2), .B(n3), .Z(carry_on_d) );
  ANDN U5 ( .B(n4), .A(n5), .Z(n2) );
  XOR U6 ( .A(b[31]), .B(n3), .Z(n4) );
  XNOR U7 ( .A(b[9]), .B(n6), .Z(c[9]) );
  XNOR U8 ( .A(b[8]), .B(n7), .Z(c[8]) );
  XNOR U9 ( .A(b[7]), .B(n8), .Z(c[7]) );
  XNOR U10 ( .A(b[6]), .B(n9), .Z(c[6]) );
  XNOR U11 ( .A(b[5]), .B(n10), .Z(c[5]) );
  XNOR U12 ( .A(b[4]), .B(n11), .Z(c[4]) );
  XNOR U13 ( .A(b[3]), .B(n12), .Z(c[3]) );
  XNOR U14 ( .A(b[31]), .B(n5), .Z(c[31]) );
  XNOR U15 ( .A(a[31]), .B(n3), .Z(n5) );
  XNOR U16 ( .A(n13), .B(n14), .Z(n3) );
  ANDN U17 ( .B(n15), .A(n16), .Z(n13) );
  XNOR U18 ( .A(b[30]), .B(n14), .Z(n15) );
  XNOR U19 ( .A(b[30]), .B(n16), .Z(c[30]) );
  XNOR U20 ( .A(a[30]), .B(n17), .Z(n16) );
  IV U21 ( .A(n14), .Z(n17) );
  XOR U22 ( .A(n18), .B(n19), .Z(n14) );
  ANDN U23 ( .B(n20), .A(n21), .Z(n18) );
  XNOR U24 ( .A(b[29]), .B(n19), .Z(n20) );
  XNOR U25 ( .A(b[2]), .B(n22), .Z(c[2]) );
  XNOR U26 ( .A(b[29]), .B(n21), .Z(c[29]) );
  XNOR U27 ( .A(a[29]), .B(n23), .Z(n21) );
  IV U28 ( .A(n19), .Z(n23) );
  XOR U29 ( .A(n24), .B(n25), .Z(n19) );
  ANDN U30 ( .B(n26), .A(n27), .Z(n24) );
  XNOR U31 ( .A(b[28]), .B(n25), .Z(n26) );
  XNOR U32 ( .A(b[28]), .B(n27), .Z(c[28]) );
  XNOR U33 ( .A(a[28]), .B(n28), .Z(n27) );
  IV U34 ( .A(n25), .Z(n28) );
  XOR U35 ( .A(n29), .B(n30), .Z(n25) );
  ANDN U36 ( .B(n31), .A(n32), .Z(n29) );
  XNOR U37 ( .A(b[27]), .B(n30), .Z(n31) );
  XNOR U38 ( .A(b[27]), .B(n32), .Z(c[27]) );
  XNOR U39 ( .A(a[27]), .B(n33), .Z(n32) );
  IV U40 ( .A(n30), .Z(n33) );
  XOR U41 ( .A(n34), .B(n35), .Z(n30) );
  ANDN U42 ( .B(n36), .A(n37), .Z(n34) );
  XNOR U43 ( .A(b[26]), .B(n35), .Z(n36) );
  XNOR U44 ( .A(b[26]), .B(n37), .Z(c[26]) );
  XNOR U45 ( .A(a[26]), .B(n38), .Z(n37) );
  IV U46 ( .A(n35), .Z(n38) );
  XOR U47 ( .A(n39), .B(n40), .Z(n35) );
  ANDN U48 ( .B(n41), .A(n42), .Z(n39) );
  XNOR U49 ( .A(b[25]), .B(n40), .Z(n41) );
  XNOR U50 ( .A(b[25]), .B(n42), .Z(c[25]) );
  XNOR U51 ( .A(a[25]), .B(n43), .Z(n42) );
  IV U52 ( .A(n40), .Z(n43) );
  XOR U53 ( .A(n44), .B(n45), .Z(n40) );
  ANDN U54 ( .B(n46), .A(n47), .Z(n44) );
  XNOR U55 ( .A(b[24]), .B(n45), .Z(n46) );
  XNOR U56 ( .A(b[24]), .B(n47), .Z(c[24]) );
  XNOR U57 ( .A(a[24]), .B(n48), .Z(n47) );
  IV U58 ( .A(n45), .Z(n48) );
  XOR U59 ( .A(n49), .B(n50), .Z(n45) );
  ANDN U60 ( .B(n51), .A(n52), .Z(n49) );
  XNOR U61 ( .A(b[23]), .B(n50), .Z(n51) );
  XNOR U62 ( .A(b[23]), .B(n52), .Z(c[23]) );
  XNOR U63 ( .A(a[23]), .B(n53), .Z(n52) );
  IV U64 ( .A(n50), .Z(n53) );
  XOR U65 ( .A(n54), .B(n55), .Z(n50) );
  ANDN U66 ( .B(n56), .A(n57), .Z(n54) );
  XNOR U67 ( .A(b[22]), .B(n55), .Z(n56) );
  XNOR U68 ( .A(b[22]), .B(n57), .Z(c[22]) );
  XNOR U69 ( .A(a[22]), .B(n58), .Z(n57) );
  IV U70 ( .A(n55), .Z(n58) );
  XOR U71 ( .A(n59), .B(n60), .Z(n55) );
  ANDN U72 ( .B(n61), .A(n62), .Z(n59) );
  XNOR U73 ( .A(b[21]), .B(n60), .Z(n61) );
  XNOR U74 ( .A(b[21]), .B(n62), .Z(c[21]) );
  XNOR U75 ( .A(a[21]), .B(n63), .Z(n62) );
  IV U76 ( .A(n60), .Z(n63) );
  XOR U77 ( .A(n64), .B(n65), .Z(n60) );
  ANDN U78 ( .B(n66), .A(n67), .Z(n64) );
  XNOR U79 ( .A(b[20]), .B(n65), .Z(n66) );
  XNOR U80 ( .A(b[20]), .B(n67), .Z(c[20]) );
  XNOR U81 ( .A(a[20]), .B(n68), .Z(n67) );
  IV U82 ( .A(n65), .Z(n68) );
  XOR U83 ( .A(n69), .B(n70), .Z(n65) );
  ANDN U84 ( .B(n71), .A(n72), .Z(n69) );
  XNOR U85 ( .A(b[19]), .B(n70), .Z(n71) );
  XNOR U86 ( .A(b[1]), .B(n73), .Z(c[1]) );
  XNOR U87 ( .A(b[19]), .B(n72), .Z(c[19]) );
  XNOR U88 ( .A(a[19]), .B(n74), .Z(n72) );
  IV U89 ( .A(n70), .Z(n74) );
  XOR U90 ( .A(n75), .B(n76), .Z(n70) );
  ANDN U91 ( .B(n77), .A(n78), .Z(n75) );
  XNOR U92 ( .A(b[18]), .B(n76), .Z(n77) );
  XNOR U93 ( .A(b[18]), .B(n78), .Z(c[18]) );
  XNOR U94 ( .A(a[18]), .B(n79), .Z(n78) );
  IV U95 ( .A(n76), .Z(n79) );
  XOR U96 ( .A(n80), .B(n81), .Z(n76) );
  ANDN U97 ( .B(n82), .A(n83), .Z(n80) );
  XNOR U98 ( .A(b[17]), .B(n81), .Z(n82) );
  XNOR U99 ( .A(b[17]), .B(n83), .Z(c[17]) );
  XNOR U100 ( .A(a[17]), .B(n84), .Z(n83) );
  IV U101 ( .A(n81), .Z(n84) );
  XOR U102 ( .A(n85), .B(n86), .Z(n81) );
  ANDN U103 ( .B(n87), .A(n88), .Z(n85) );
  XNOR U104 ( .A(b[16]), .B(n86), .Z(n87) );
  XNOR U105 ( .A(b[16]), .B(n88), .Z(c[16]) );
  XNOR U106 ( .A(a[16]), .B(n89), .Z(n88) );
  IV U107 ( .A(n86), .Z(n89) );
  XOR U108 ( .A(n90), .B(n91), .Z(n86) );
  ANDN U109 ( .B(n92), .A(n93), .Z(n90) );
  XNOR U110 ( .A(b[15]), .B(n91), .Z(n92) );
  XNOR U111 ( .A(b[15]), .B(n93), .Z(c[15]) );
  XNOR U112 ( .A(a[15]), .B(n94), .Z(n93) );
  IV U113 ( .A(n91), .Z(n94) );
  XOR U114 ( .A(n95), .B(n96), .Z(n91) );
  ANDN U115 ( .B(n97), .A(n98), .Z(n95) );
  XNOR U116 ( .A(b[14]), .B(n96), .Z(n97) );
  XNOR U117 ( .A(b[14]), .B(n98), .Z(c[14]) );
  XNOR U118 ( .A(a[14]), .B(n99), .Z(n98) );
  IV U119 ( .A(n96), .Z(n99) );
  XOR U120 ( .A(n100), .B(n101), .Z(n96) );
  ANDN U121 ( .B(n102), .A(n103), .Z(n100) );
  XNOR U122 ( .A(b[13]), .B(n101), .Z(n102) );
  XNOR U123 ( .A(b[13]), .B(n103), .Z(c[13]) );
  XNOR U124 ( .A(a[13]), .B(n104), .Z(n103) );
  IV U125 ( .A(n101), .Z(n104) );
  XOR U126 ( .A(n105), .B(n106), .Z(n101) );
  ANDN U127 ( .B(n107), .A(n108), .Z(n105) );
  XNOR U128 ( .A(b[12]), .B(n106), .Z(n107) );
  XNOR U129 ( .A(b[12]), .B(n108), .Z(c[12]) );
  XNOR U130 ( .A(a[12]), .B(n109), .Z(n108) );
  IV U131 ( .A(n106), .Z(n109) );
  XOR U132 ( .A(n110), .B(n111), .Z(n106) );
  ANDN U133 ( .B(n112), .A(n113), .Z(n110) );
  XNOR U134 ( .A(b[11]), .B(n111), .Z(n112) );
  XNOR U135 ( .A(b[11]), .B(n113), .Z(c[11]) );
  XNOR U136 ( .A(a[11]), .B(n114), .Z(n113) );
  IV U137 ( .A(n111), .Z(n114) );
  XOR U138 ( .A(n115), .B(n116), .Z(n111) );
  ANDN U139 ( .B(n117), .A(n118), .Z(n115) );
  XNOR U140 ( .A(b[10]), .B(n116), .Z(n117) );
  XNOR U141 ( .A(b[10]), .B(n118), .Z(c[10]) );
  XNOR U142 ( .A(a[10]), .B(n119), .Z(n118) );
  IV U143 ( .A(n116), .Z(n119) );
  XOR U144 ( .A(n120), .B(n121), .Z(n116) );
  ANDN U145 ( .B(n122), .A(n6), .Z(n120) );
  XNOR U146 ( .A(a[9]), .B(n123), .Z(n6) );
  IV U147 ( .A(n121), .Z(n123) );
  XNOR U148 ( .A(b[9]), .B(n121), .Z(n122) );
  XOR U149 ( .A(n124), .B(n125), .Z(n121) );
  ANDN U150 ( .B(n126), .A(n7), .Z(n124) );
  XNOR U151 ( .A(a[8]), .B(n127), .Z(n7) );
  IV U152 ( .A(n125), .Z(n127) );
  XNOR U153 ( .A(b[8]), .B(n125), .Z(n126) );
  XOR U154 ( .A(n128), .B(n129), .Z(n125) );
  ANDN U155 ( .B(n130), .A(n8), .Z(n128) );
  XNOR U156 ( .A(a[7]), .B(n131), .Z(n8) );
  IV U157 ( .A(n129), .Z(n131) );
  XNOR U158 ( .A(b[7]), .B(n129), .Z(n130) );
  XOR U159 ( .A(n132), .B(n133), .Z(n129) );
  ANDN U160 ( .B(n134), .A(n9), .Z(n132) );
  XNOR U161 ( .A(a[6]), .B(n135), .Z(n9) );
  IV U162 ( .A(n133), .Z(n135) );
  XNOR U163 ( .A(b[6]), .B(n133), .Z(n134) );
  XOR U164 ( .A(n136), .B(n137), .Z(n133) );
  ANDN U165 ( .B(n138), .A(n10), .Z(n136) );
  XNOR U166 ( .A(a[5]), .B(n139), .Z(n10) );
  IV U167 ( .A(n137), .Z(n139) );
  XNOR U168 ( .A(b[5]), .B(n137), .Z(n138) );
  XOR U169 ( .A(n140), .B(n141), .Z(n137) );
  ANDN U170 ( .B(n142), .A(n11), .Z(n140) );
  XNOR U171 ( .A(a[4]), .B(n143), .Z(n11) );
  IV U172 ( .A(n141), .Z(n143) );
  XNOR U173 ( .A(b[4]), .B(n141), .Z(n142) );
  XOR U174 ( .A(n144), .B(n145), .Z(n141) );
  ANDN U175 ( .B(n146), .A(n12), .Z(n144) );
  XNOR U176 ( .A(a[3]), .B(n147), .Z(n12) );
  IV U177 ( .A(n145), .Z(n147) );
  XNOR U178 ( .A(b[3]), .B(n145), .Z(n146) );
  XOR U179 ( .A(n148), .B(n149), .Z(n145) );
  ANDN U180 ( .B(n150), .A(n22), .Z(n148) );
  XNOR U181 ( .A(a[2]), .B(n151), .Z(n22) );
  IV U182 ( .A(n149), .Z(n151) );
  XNOR U183 ( .A(b[2]), .B(n149), .Z(n150) );
  XOR U184 ( .A(n152), .B(n153), .Z(n149) );
  ANDN U185 ( .B(n154), .A(n73), .Z(n152) );
  XNOR U186 ( .A(a[1]), .B(n155), .Z(n73) );
  IV U187 ( .A(n153), .Z(n155) );
  XNOR U188 ( .A(b[1]), .B(n153), .Z(n154) );
  XOR U189 ( .A(carry_on), .B(n156), .Z(n153) );
  NANDN U190 ( .A(n157), .B(n158), .Z(n156) );
  XOR U191 ( .A(carry_on), .B(b[0]), .Z(n158) );
  XNOR U192 ( .A(b[0]), .B(n157), .Z(c[0]) );
  XNOR U193 ( .A(a[0]), .B(carry_on), .Z(n157) );
endmodule

