
module sum_N262144_CC4096 ( clk, rst, a, b, c );
  input [63:0] a;
  input [63:0] b;
  output [63:0] c;
  input clk, rst;
  wire   carry_on, carry_on_d, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
         n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141,
         n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256;

  DFF carry_on_reg ( .D(carry_on_d), .CLK(clk), .RST(rst), .I(1'b0), .Q(
        carry_on) );
  XOR U4 ( .A(a[3]), .B(n246), .Z(n108) );
  XOR U5 ( .A(a[6]), .B(n237), .Z(n9) );
  XOR U6 ( .A(a[9]), .B(n228), .Z(n6) );
  XOR U7 ( .A(a[12]), .B(n216), .Z(n218) );
  XOR U8 ( .A(a[15]), .B(n204), .Z(n206) );
  XOR U9 ( .A(a[18]), .B(n192), .Z(n194) );
  XOR U10 ( .A(a[21]), .B(n179), .Z(n181) );
  XOR U11 ( .A(a[24]), .B(n167), .Z(n169) );
  XOR U12 ( .A(a[27]), .B(n155), .Z(n157) );
  XOR U13 ( .A(a[30]), .B(n142), .Z(n144) );
  XOR U14 ( .A(a[33]), .B(n130), .Z(n132) );
  XOR U15 ( .A(a[36]), .B(n118), .Z(n120) );
  XOR U16 ( .A(a[39]), .B(n105), .Z(n107) );
  XOR U17 ( .A(a[42]), .B(n93), .Z(n95) );
  XOR U18 ( .A(a[45]), .B(n81), .Z(n83) );
  XOR U19 ( .A(a[48]), .B(n69), .Z(n71) );
  XOR U20 ( .A(a[51]), .B(n56), .Z(n58) );
  XOR U21 ( .A(a[54]), .B(n44), .Z(n46) );
  XOR U22 ( .A(a[57]), .B(n32), .Z(n34) );
  XOR U23 ( .A(a[60]), .B(n19), .Z(n21) );
  XOR U24 ( .A(a[1]), .B(n252), .Z(n190) );
  XOR U25 ( .A(a[4]), .B(n243), .Z(n67) );
  XOR U26 ( .A(a[7]), .B(n234), .Z(n8) );
  XOR U27 ( .A(a[10]), .B(n224), .Z(n226) );
  XOR U28 ( .A(a[13]), .B(n212), .Z(n214) );
  XOR U29 ( .A(a[16]), .B(n200), .Z(n202) );
  XOR U30 ( .A(a[19]), .B(n187), .Z(n189) );
  XOR U31 ( .A(a[22]), .B(n175), .Z(n177) );
  XOR U32 ( .A(a[25]), .B(n163), .Z(n165) );
  XOR U33 ( .A(a[28]), .B(n151), .Z(n153) );
  XOR U34 ( .A(a[31]), .B(n138), .Z(n140) );
  XOR U35 ( .A(a[34]), .B(n126), .Z(n128) );
  XOR U36 ( .A(a[37]), .B(n114), .Z(n116) );
  XOR U37 ( .A(a[40]), .B(n101), .Z(n103) );
  XOR U38 ( .A(a[43]), .B(n89), .Z(n91) );
  XOR U39 ( .A(a[46]), .B(n77), .Z(n79) );
  XOR U40 ( .A(a[49]), .B(n64), .Z(n66) );
  XOR U41 ( .A(a[52]), .B(n52), .Z(n54) );
  XOR U42 ( .A(a[55]), .B(n40), .Z(n42) );
  XOR U43 ( .A(a[58]), .B(n28), .Z(n30) );
  XOR U44 ( .A(a[61]), .B(n15), .Z(n17) );
  XOR U45 ( .A(a[2]), .B(n249), .Z(n149) );
  XOR U46 ( .A(a[5]), .B(n240), .Z(n26) );
  XOR U47 ( .A(a[8]), .B(n231), .Z(n7) );
  XOR U48 ( .A(a[11]), .B(n220), .Z(n222) );
  XOR U49 ( .A(a[14]), .B(n208), .Z(n210) );
  XOR U50 ( .A(a[17]), .B(n196), .Z(n198) );
  XOR U51 ( .A(a[20]), .B(n183), .Z(n185) );
  XOR U52 ( .A(a[23]), .B(n171), .Z(n173) );
  XOR U53 ( .A(a[26]), .B(n159), .Z(n161) );
  XOR U54 ( .A(a[29]), .B(n146), .Z(n148) );
  XOR U55 ( .A(a[32]), .B(n134), .Z(n136) );
  XOR U56 ( .A(a[35]), .B(n122), .Z(n124) );
  XOR U57 ( .A(a[38]), .B(n110), .Z(n112) );
  XOR U58 ( .A(a[41]), .B(n97), .Z(n99) );
  XOR U59 ( .A(a[44]), .B(n85), .Z(n87) );
  XOR U60 ( .A(a[47]), .B(n73), .Z(n75) );
  XOR U61 ( .A(a[50]), .B(n60), .Z(n62) );
  XOR U62 ( .A(a[53]), .B(n48), .Z(n50) );
  XOR U63 ( .A(a[56]), .B(n36), .Z(n38) );
  XOR U64 ( .A(a[59]), .B(n23), .Z(n25) );
  XOR U65 ( .A(a[62]), .B(n11), .Z(n13) );
  XOR U66 ( .A(n2), .B(n3), .Z(carry_on_d) );
  ANDN U67 ( .B(n4), .A(n5), .Z(n2) );
  XOR U68 ( .A(b[63]), .B(n3), .Z(n4) );
  XNOR U69 ( .A(b[9]), .B(n6), .Z(c[9]) );
  XNOR U70 ( .A(b[8]), .B(n7), .Z(c[8]) );
  XNOR U71 ( .A(b[7]), .B(n8), .Z(c[7]) );
  XNOR U72 ( .A(b[6]), .B(n9), .Z(c[6]) );
  XNOR U73 ( .A(b[63]), .B(n5), .Z(c[63]) );
  XNOR U74 ( .A(a[63]), .B(n3), .Z(n5) );
  XNOR U75 ( .A(n10), .B(n11), .Z(n3) );
  ANDN U76 ( .B(n12), .A(n13), .Z(n10) );
  XNOR U77 ( .A(b[62]), .B(n11), .Z(n12) );
  XNOR U78 ( .A(b[62]), .B(n13), .Z(c[62]) );
  XOR U79 ( .A(n14), .B(n15), .Z(n11) );
  ANDN U80 ( .B(n16), .A(n17), .Z(n14) );
  XNOR U81 ( .A(b[61]), .B(n15), .Z(n16) );
  XNOR U82 ( .A(b[61]), .B(n17), .Z(c[61]) );
  XOR U83 ( .A(n18), .B(n19), .Z(n15) );
  ANDN U84 ( .B(n20), .A(n21), .Z(n18) );
  XNOR U85 ( .A(b[60]), .B(n19), .Z(n20) );
  XNOR U86 ( .A(b[60]), .B(n21), .Z(c[60]) );
  XOR U87 ( .A(n22), .B(n23), .Z(n19) );
  ANDN U88 ( .B(n24), .A(n25), .Z(n22) );
  XNOR U89 ( .A(b[59]), .B(n23), .Z(n24) );
  XNOR U90 ( .A(b[5]), .B(n26), .Z(c[5]) );
  XNOR U91 ( .A(b[59]), .B(n25), .Z(c[59]) );
  XOR U92 ( .A(n27), .B(n28), .Z(n23) );
  ANDN U93 ( .B(n29), .A(n30), .Z(n27) );
  XNOR U94 ( .A(b[58]), .B(n28), .Z(n29) );
  XNOR U95 ( .A(b[58]), .B(n30), .Z(c[58]) );
  XOR U96 ( .A(n31), .B(n32), .Z(n28) );
  ANDN U97 ( .B(n33), .A(n34), .Z(n31) );
  XNOR U98 ( .A(b[57]), .B(n32), .Z(n33) );
  XNOR U99 ( .A(b[57]), .B(n34), .Z(c[57]) );
  XOR U100 ( .A(n35), .B(n36), .Z(n32) );
  ANDN U101 ( .B(n37), .A(n38), .Z(n35) );
  XNOR U102 ( .A(b[56]), .B(n36), .Z(n37) );
  XNOR U103 ( .A(b[56]), .B(n38), .Z(c[56]) );
  XOR U104 ( .A(n39), .B(n40), .Z(n36) );
  ANDN U105 ( .B(n41), .A(n42), .Z(n39) );
  XNOR U106 ( .A(b[55]), .B(n40), .Z(n41) );
  XNOR U107 ( .A(b[55]), .B(n42), .Z(c[55]) );
  XOR U108 ( .A(n43), .B(n44), .Z(n40) );
  ANDN U109 ( .B(n45), .A(n46), .Z(n43) );
  XNOR U110 ( .A(b[54]), .B(n44), .Z(n45) );
  XNOR U111 ( .A(b[54]), .B(n46), .Z(c[54]) );
  XOR U112 ( .A(n47), .B(n48), .Z(n44) );
  ANDN U113 ( .B(n49), .A(n50), .Z(n47) );
  XNOR U114 ( .A(b[53]), .B(n48), .Z(n49) );
  XNOR U115 ( .A(b[53]), .B(n50), .Z(c[53]) );
  XOR U116 ( .A(n51), .B(n52), .Z(n48) );
  ANDN U117 ( .B(n53), .A(n54), .Z(n51) );
  XNOR U118 ( .A(b[52]), .B(n52), .Z(n53) );
  XNOR U119 ( .A(b[52]), .B(n54), .Z(c[52]) );
  XOR U120 ( .A(n55), .B(n56), .Z(n52) );
  ANDN U121 ( .B(n57), .A(n58), .Z(n55) );
  XNOR U122 ( .A(b[51]), .B(n56), .Z(n57) );
  XNOR U123 ( .A(b[51]), .B(n58), .Z(c[51]) );
  XOR U124 ( .A(n59), .B(n60), .Z(n56) );
  ANDN U125 ( .B(n61), .A(n62), .Z(n59) );
  XNOR U126 ( .A(b[50]), .B(n60), .Z(n61) );
  XNOR U127 ( .A(b[50]), .B(n62), .Z(c[50]) );
  XOR U128 ( .A(n63), .B(n64), .Z(n60) );
  ANDN U129 ( .B(n65), .A(n66), .Z(n63) );
  XNOR U130 ( .A(b[49]), .B(n64), .Z(n65) );
  XNOR U131 ( .A(b[4]), .B(n67), .Z(c[4]) );
  XNOR U132 ( .A(b[49]), .B(n66), .Z(c[49]) );
  XOR U133 ( .A(n68), .B(n69), .Z(n64) );
  ANDN U134 ( .B(n70), .A(n71), .Z(n68) );
  XNOR U135 ( .A(b[48]), .B(n69), .Z(n70) );
  XNOR U136 ( .A(b[48]), .B(n71), .Z(c[48]) );
  XOR U137 ( .A(n72), .B(n73), .Z(n69) );
  ANDN U138 ( .B(n74), .A(n75), .Z(n72) );
  XNOR U139 ( .A(b[47]), .B(n73), .Z(n74) );
  XNOR U140 ( .A(b[47]), .B(n75), .Z(c[47]) );
  XOR U141 ( .A(n76), .B(n77), .Z(n73) );
  ANDN U142 ( .B(n78), .A(n79), .Z(n76) );
  XNOR U143 ( .A(b[46]), .B(n77), .Z(n78) );
  XNOR U144 ( .A(b[46]), .B(n79), .Z(c[46]) );
  XOR U145 ( .A(n80), .B(n81), .Z(n77) );
  ANDN U146 ( .B(n82), .A(n83), .Z(n80) );
  XNOR U147 ( .A(b[45]), .B(n81), .Z(n82) );
  XNOR U148 ( .A(b[45]), .B(n83), .Z(c[45]) );
  XOR U149 ( .A(n84), .B(n85), .Z(n81) );
  ANDN U150 ( .B(n86), .A(n87), .Z(n84) );
  XNOR U151 ( .A(b[44]), .B(n85), .Z(n86) );
  XNOR U152 ( .A(b[44]), .B(n87), .Z(c[44]) );
  XOR U153 ( .A(n88), .B(n89), .Z(n85) );
  ANDN U154 ( .B(n90), .A(n91), .Z(n88) );
  XNOR U155 ( .A(b[43]), .B(n89), .Z(n90) );
  XNOR U156 ( .A(b[43]), .B(n91), .Z(c[43]) );
  XOR U157 ( .A(n92), .B(n93), .Z(n89) );
  ANDN U158 ( .B(n94), .A(n95), .Z(n92) );
  XNOR U159 ( .A(b[42]), .B(n93), .Z(n94) );
  XNOR U160 ( .A(b[42]), .B(n95), .Z(c[42]) );
  XOR U161 ( .A(n96), .B(n97), .Z(n93) );
  ANDN U162 ( .B(n98), .A(n99), .Z(n96) );
  XNOR U163 ( .A(b[41]), .B(n97), .Z(n98) );
  XNOR U164 ( .A(b[41]), .B(n99), .Z(c[41]) );
  XOR U165 ( .A(n100), .B(n101), .Z(n97) );
  ANDN U166 ( .B(n102), .A(n103), .Z(n100) );
  XNOR U167 ( .A(b[40]), .B(n101), .Z(n102) );
  XNOR U168 ( .A(b[40]), .B(n103), .Z(c[40]) );
  XOR U169 ( .A(n104), .B(n105), .Z(n101) );
  ANDN U170 ( .B(n106), .A(n107), .Z(n104) );
  XNOR U171 ( .A(b[39]), .B(n105), .Z(n106) );
  XNOR U172 ( .A(b[3]), .B(n108), .Z(c[3]) );
  XNOR U173 ( .A(b[39]), .B(n107), .Z(c[39]) );
  XOR U174 ( .A(n109), .B(n110), .Z(n105) );
  ANDN U175 ( .B(n111), .A(n112), .Z(n109) );
  XNOR U176 ( .A(b[38]), .B(n110), .Z(n111) );
  XNOR U177 ( .A(b[38]), .B(n112), .Z(c[38]) );
  XOR U178 ( .A(n113), .B(n114), .Z(n110) );
  ANDN U179 ( .B(n115), .A(n116), .Z(n113) );
  XNOR U180 ( .A(b[37]), .B(n114), .Z(n115) );
  XNOR U181 ( .A(b[37]), .B(n116), .Z(c[37]) );
  XOR U182 ( .A(n117), .B(n118), .Z(n114) );
  ANDN U183 ( .B(n119), .A(n120), .Z(n117) );
  XNOR U184 ( .A(b[36]), .B(n118), .Z(n119) );
  XNOR U185 ( .A(b[36]), .B(n120), .Z(c[36]) );
  XOR U186 ( .A(n121), .B(n122), .Z(n118) );
  ANDN U187 ( .B(n123), .A(n124), .Z(n121) );
  XNOR U188 ( .A(b[35]), .B(n122), .Z(n123) );
  XNOR U189 ( .A(b[35]), .B(n124), .Z(c[35]) );
  XOR U190 ( .A(n125), .B(n126), .Z(n122) );
  ANDN U191 ( .B(n127), .A(n128), .Z(n125) );
  XNOR U192 ( .A(b[34]), .B(n126), .Z(n127) );
  XNOR U193 ( .A(b[34]), .B(n128), .Z(c[34]) );
  XOR U194 ( .A(n129), .B(n130), .Z(n126) );
  ANDN U195 ( .B(n131), .A(n132), .Z(n129) );
  XNOR U196 ( .A(b[33]), .B(n130), .Z(n131) );
  XNOR U197 ( .A(b[33]), .B(n132), .Z(c[33]) );
  XOR U198 ( .A(n133), .B(n134), .Z(n130) );
  ANDN U199 ( .B(n135), .A(n136), .Z(n133) );
  XNOR U200 ( .A(b[32]), .B(n134), .Z(n135) );
  XNOR U201 ( .A(b[32]), .B(n136), .Z(c[32]) );
  XOR U202 ( .A(n137), .B(n138), .Z(n134) );
  ANDN U203 ( .B(n139), .A(n140), .Z(n137) );
  XNOR U204 ( .A(b[31]), .B(n138), .Z(n139) );
  XNOR U205 ( .A(b[31]), .B(n140), .Z(c[31]) );
  XOR U206 ( .A(n141), .B(n142), .Z(n138) );
  ANDN U207 ( .B(n143), .A(n144), .Z(n141) );
  XNOR U208 ( .A(b[30]), .B(n142), .Z(n143) );
  XNOR U209 ( .A(b[30]), .B(n144), .Z(c[30]) );
  XOR U210 ( .A(n145), .B(n146), .Z(n142) );
  ANDN U211 ( .B(n147), .A(n148), .Z(n145) );
  XNOR U212 ( .A(b[29]), .B(n146), .Z(n147) );
  XNOR U213 ( .A(b[2]), .B(n149), .Z(c[2]) );
  XNOR U214 ( .A(b[29]), .B(n148), .Z(c[29]) );
  XOR U215 ( .A(n150), .B(n151), .Z(n146) );
  ANDN U216 ( .B(n152), .A(n153), .Z(n150) );
  XNOR U217 ( .A(b[28]), .B(n151), .Z(n152) );
  XNOR U218 ( .A(b[28]), .B(n153), .Z(c[28]) );
  XOR U219 ( .A(n154), .B(n155), .Z(n151) );
  ANDN U220 ( .B(n156), .A(n157), .Z(n154) );
  XNOR U221 ( .A(b[27]), .B(n155), .Z(n156) );
  XNOR U222 ( .A(b[27]), .B(n157), .Z(c[27]) );
  XOR U223 ( .A(n158), .B(n159), .Z(n155) );
  ANDN U224 ( .B(n160), .A(n161), .Z(n158) );
  XNOR U225 ( .A(b[26]), .B(n159), .Z(n160) );
  XNOR U226 ( .A(b[26]), .B(n161), .Z(c[26]) );
  XOR U227 ( .A(n162), .B(n163), .Z(n159) );
  ANDN U228 ( .B(n164), .A(n165), .Z(n162) );
  XNOR U229 ( .A(b[25]), .B(n163), .Z(n164) );
  XNOR U230 ( .A(b[25]), .B(n165), .Z(c[25]) );
  XOR U231 ( .A(n166), .B(n167), .Z(n163) );
  ANDN U232 ( .B(n168), .A(n169), .Z(n166) );
  XNOR U233 ( .A(b[24]), .B(n167), .Z(n168) );
  XNOR U234 ( .A(b[24]), .B(n169), .Z(c[24]) );
  XOR U235 ( .A(n170), .B(n171), .Z(n167) );
  ANDN U236 ( .B(n172), .A(n173), .Z(n170) );
  XNOR U237 ( .A(b[23]), .B(n171), .Z(n172) );
  XNOR U238 ( .A(b[23]), .B(n173), .Z(c[23]) );
  XOR U239 ( .A(n174), .B(n175), .Z(n171) );
  ANDN U240 ( .B(n176), .A(n177), .Z(n174) );
  XNOR U241 ( .A(b[22]), .B(n175), .Z(n176) );
  XNOR U242 ( .A(b[22]), .B(n177), .Z(c[22]) );
  XOR U243 ( .A(n178), .B(n179), .Z(n175) );
  ANDN U244 ( .B(n180), .A(n181), .Z(n178) );
  XNOR U245 ( .A(b[21]), .B(n179), .Z(n180) );
  XNOR U246 ( .A(b[21]), .B(n181), .Z(c[21]) );
  XOR U247 ( .A(n182), .B(n183), .Z(n179) );
  ANDN U248 ( .B(n184), .A(n185), .Z(n182) );
  XNOR U249 ( .A(b[20]), .B(n183), .Z(n184) );
  XNOR U250 ( .A(b[20]), .B(n185), .Z(c[20]) );
  XOR U251 ( .A(n186), .B(n187), .Z(n183) );
  ANDN U252 ( .B(n188), .A(n189), .Z(n186) );
  XNOR U253 ( .A(b[19]), .B(n187), .Z(n188) );
  XNOR U254 ( .A(b[1]), .B(n190), .Z(c[1]) );
  XNOR U255 ( .A(b[19]), .B(n189), .Z(c[19]) );
  XOR U256 ( .A(n191), .B(n192), .Z(n187) );
  ANDN U257 ( .B(n193), .A(n194), .Z(n191) );
  XNOR U258 ( .A(b[18]), .B(n192), .Z(n193) );
  XNOR U259 ( .A(b[18]), .B(n194), .Z(c[18]) );
  XOR U260 ( .A(n195), .B(n196), .Z(n192) );
  ANDN U261 ( .B(n197), .A(n198), .Z(n195) );
  XNOR U262 ( .A(b[17]), .B(n196), .Z(n197) );
  XNOR U263 ( .A(b[17]), .B(n198), .Z(c[17]) );
  XOR U264 ( .A(n199), .B(n200), .Z(n196) );
  ANDN U265 ( .B(n201), .A(n202), .Z(n199) );
  XNOR U266 ( .A(b[16]), .B(n200), .Z(n201) );
  XNOR U267 ( .A(b[16]), .B(n202), .Z(c[16]) );
  XOR U268 ( .A(n203), .B(n204), .Z(n200) );
  ANDN U269 ( .B(n205), .A(n206), .Z(n203) );
  XNOR U270 ( .A(b[15]), .B(n204), .Z(n205) );
  XNOR U271 ( .A(b[15]), .B(n206), .Z(c[15]) );
  XOR U272 ( .A(n207), .B(n208), .Z(n204) );
  ANDN U273 ( .B(n209), .A(n210), .Z(n207) );
  XNOR U274 ( .A(b[14]), .B(n208), .Z(n209) );
  XNOR U275 ( .A(b[14]), .B(n210), .Z(c[14]) );
  XOR U276 ( .A(n211), .B(n212), .Z(n208) );
  ANDN U277 ( .B(n213), .A(n214), .Z(n211) );
  XNOR U278 ( .A(b[13]), .B(n212), .Z(n213) );
  XNOR U279 ( .A(b[13]), .B(n214), .Z(c[13]) );
  XOR U280 ( .A(n215), .B(n216), .Z(n212) );
  ANDN U281 ( .B(n217), .A(n218), .Z(n215) );
  XNOR U282 ( .A(b[12]), .B(n216), .Z(n217) );
  XNOR U283 ( .A(b[12]), .B(n218), .Z(c[12]) );
  XOR U284 ( .A(n219), .B(n220), .Z(n216) );
  ANDN U285 ( .B(n221), .A(n222), .Z(n219) );
  XNOR U286 ( .A(b[11]), .B(n220), .Z(n221) );
  XNOR U287 ( .A(b[11]), .B(n222), .Z(c[11]) );
  XOR U288 ( .A(n223), .B(n224), .Z(n220) );
  ANDN U289 ( .B(n225), .A(n226), .Z(n223) );
  XNOR U290 ( .A(b[10]), .B(n224), .Z(n225) );
  XNOR U291 ( .A(b[10]), .B(n226), .Z(c[10]) );
  XOR U292 ( .A(n227), .B(n228), .Z(n224) );
  ANDN U293 ( .B(n229), .A(n6), .Z(n227) );
  XNOR U294 ( .A(b[9]), .B(n228), .Z(n229) );
  XOR U295 ( .A(n230), .B(n231), .Z(n228) );
  ANDN U296 ( .B(n232), .A(n7), .Z(n230) );
  XNOR U297 ( .A(b[8]), .B(n231), .Z(n232) );
  XOR U298 ( .A(n233), .B(n234), .Z(n231) );
  ANDN U299 ( .B(n235), .A(n8), .Z(n233) );
  XNOR U300 ( .A(b[7]), .B(n234), .Z(n235) );
  XOR U301 ( .A(n236), .B(n237), .Z(n234) );
  ANDN U302 ( .B(n238), .A(n9), .Z(n236) );
  XNOR U303 ( .A(b[6]), .B(n237), .Z(n238) );
  XOR U304 ( .A(n239), .B(n240), .Z(n237) );
  ANDN U305 ( .B(n241), .A(n26), .Z(n239) );
  XNOR U306 ( .A(b[5]), .B(n240), .Z(n241) );
  XOR U307 ( .A(n242), .B(n243), .Z(n240) );
  ANDN U308 ( .B(n244), .A(n67), .Z(n242) );
  XNOR U309 ( .A(b[4]), .B(n243), .Z(n244) );
  XOR U310 ( .A(n245), .B(n246), .Z(n243) );
  ANDN U311 ( .B(n247), .A(n108), .Z(n245) );
  XNOR U312 ( .A(b[3]), .B(n246), .Z(n247) );
  XOR U313 ( .A(n248), .B(n249), .Z(n246) );
  ANDN U314 ( .B(n250), .A(n149), .Z(n248) );
  XNOR U315 ( .A(b[2]), .B(n249), .Z(n250) );
  XOR U316 ( .A(n251), .B(n252), .Z(n249) );
  ANDN U317 ( .B(n253), .A(n190), .Z(n251) );
  XNOR U318 ( .A(b[1]), .B(n252), .Z(n253) );
  XOR U319 ( .A(carry_on), .B(n254), .Z(n252) );
  NANDN U320 ( .A(n255), .B(n256), .Z(n254) );
  XOR U321 ( .A(carry_on), .B(b[0]), .Z(n256) );
  XNOR U322 ( .A(b[0]), .B(n255), .Z(c[0]) );
  XNOR U323 ( .A(a[0]), .B(carry_on), .Z(n255) );
endmodule

