
module mult_N1024_CC1024 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [0:0] b;
  output [2047:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118;
  wire   [2047:0] sreg;

  DFF \sreg_reg[2046]  ( .D(c[2047]), .CLK(clk), .RST(rst), .Q(sreg[2046]) );
  DFF \sreg_reg[2045]  ( .D(c[2046]), .CLK(clk), .RST(rst), .Q(sreg[2045]) );
  DFF \sreg_reg[2044]  ( .D(c[2045]), .CLK(clk), .RST(rst), .Q(sreg[2044]) );
  DFF \sreg_reg[2043]  ( .D(c[2044]), .CLK(clk), .RST(rst), .Q(sreg[2043]) );
  DFF \sreg_reg[2042]  ( .D(c[2043]), .CLK(clk), .RST(rst), .Q(sreg[2042]) );
  DFF \sreg_reg[2041]  ( .D(c[2042]), .CLK(clk), .RST(rst), .Q(sreg[2041]) );
  DFF \sreg_reg[2040]  ( .D(c[2041]), .CLK(clk), .RST(rst), .Q(sreg[2040]) );
  DFF \sreg_reg[2039]  ( .D(c[2040]), .CLK(clk), .RST(rst), .Q(sreg[2039]) );
  DFF \sreg_reg[2038]  ( .D(c[2039]), .CLK(clk), .RST(rst), .Q(sreg[2038]) );
  DFF \sreg_reg[2037]  ( .D(c[2038]), .CLK(clk), .RST(rst), .Q(sreg[2037]) );
  DFF \sreg_reg[2036]  ( .D(c[2037]), .CLK(clk), .RST(rst), .Q(sreg[2036]) );
  DFF \sreg_reg[2035]  ( .D(c[2036]), .CLK(clk), .RST(rst), .Q(sreg[2035]) );
  DFF \sreg_reg[2034]  ( .D(c[2035]), .CLK(clk), .RST(rst), .Q(sreg[2034]) );
  DFF \sreg_reg[2033]  ( .D(c[2034]), .CLK(clk), .RST(rst), .Q(sreg[2033]) );
  DFF \sreg_reg[2032]  ( .D(c[2033]), .CLK(clk), .RST(rst), .Q(sreg[2032]) );
  DFF \sreg_reg[2031]  ( .D(c[2032]), .CLK(clk), .RST(rst), .Q(sreg[2031]) );
  DFF \sreg_reg[2030]  ( .D(c[2031]), .CLK(clk), .RST(rst), .Q(sreg[2030]) );
  DFF \sreg_reg[2029]  ( .D(c[2030]), .CLK(clk), .RST(rst), .Q(sreg[2029]) );
  DFF \sreg_reg[2028]  ( .D(c[2029]), .CLK(clk), .RST(rst), .Q(sreg[2028]) );
  DFF \sreg_reg[2027]  ( .D(c[2028]), .CLK(clk), .RST(rst), .Q(sreg[2027]) );
  DFF \sreg_reg[2026]  ( .D(c[2027]), .CLK(clk), .RST(rst), .Q(sreg[2026]) );
  DFF \sreg_reg[2025]  ( .D(c[2026]), .CLK(clk), .RST(rst), .Q(sreg[2025]) );
  DFF \sreg_reg[2024]  ( .D(c[2025]), .CLK(clk), .RST(rst), .Q(sreg[2024]) );
  DFF \sreg_reg[2023]  ( .D(c[2024]), .CLK(clk), .RST(rst), .Q(sreg[2023]) );
  DFF \sreg_reg[2022]  ( .D(c[2023]), .CLK(clk), .RST(rst), .Q(sreg[2022]) );
  DFF \sreg_reg[2021]  ( .D(c[2022]), .CLK(clk), .RST(rst), .Q(sreg[2021]) );
  DFF \sreg_reg[2020]  ( .D(c[2021]), .CLK(clk), .RST(rst), .Q(sreg[2020]) );
  DFF \sreg_reg[2019]  ( .D(c[2020]), .CLK(clk), .RST(rst), .Q(sreg[2019]) );
  DFF \sreg_reg[2018]  ( .D(c[2019]), .CLK(clk), .RST(rst), .Q(sreg[2018]) );
  DFF \sreg_reg[2017]  ( .D(c[2018]), .CLK(clk), .RST(rst), .Q(sreg[2017]) );
  DFF \sreg_reg[2016]  ( .D(c[2017]), .CLK(clk), .RST(rst), .Q(sreg[2016]) );
  DFF \sreg_reg[2015]  ( .D(c[2016]), .CLK(clk), .RST(rst), .Q(sreg[2015]) );
  DFF \sreg_reg[2014]  ( .D(c[2015]), .CLK(clk), .RST(rst), .Q(sreg[2014]) );
  DFF \sreg_reg[2013]  ( .D(c[2014]), .CLK(clk), .RST(rst), .Q(sreg[2013]) );
  DFF \sreg_reg[2012]  ( .D(c[2013]), .CLK(clk), .RST(rst), .Q(sreg[2012]) );
  DFF \sreg_reg[2011]  ( .D(c[2012]), .CLK(clk), .RST(rst), .Q(sreg[2011]) );
  DFF \sreg_reg[2010]  ( .D(c[2011]), .CLK(clk), .RST(rst), .Q(sreg[2010]) );
  DFF \sreg_reg[2009]  ( .D(c[2010]), .CLK(clk), .RST(rst), .Q(sreg[2009]) );
  DFF \sreg_reg[2008]  ( .D(c[2009]), .CLK(clk), .RST(rst), .Q(sreg[2008]) );
  DFF \sreg_reg[2007]  ( .D(c[2008]), .CLK(clk), .RST(rst), .Q(sreg[2007]) );
  DFF \sreg_reg[2006]  ( .D(c[2007]), .CLK(clk), .RST(rst), .Q(sreg[2006]) );
  DFF \sreg_reg[2005]  ( .D(c[2006]), .CLK(clk), .RST(rst), .Q(sreg[2005]) );
  DFF \sreg_reg[2004]  ( .D(c[2005]), .CLK(clk), .RST(rst), .Q(sreg[2004]) );
  DFF \sreg_reg[2003]  ( .D(c[2004]), .CLK(clk), .RST(rst), .Q(sreg[2003]) );
  DFF \sreg_reg[2002]  ( .D(c[2003]), .CLK(clk), .RST(rst), .Q(sreg[2002]) );
  DFF \sreg_reg[2001]  ( .D(c[2002]), .CLK(clk), .RST(rst), .Q(sreg[2001]) );
  DFF \sreg_reg[2000]  ( .D(c[2001]), .CLK(clk), .RST(rst), .Q(sreg[2000]) );
  DFF \sreg_reg[1999]  ( .D(c[2000]), .CLK(clk), .RST(rst), .Q(sreg[1999]) );
  DFF \sreg_reg[1998]  ( .D(c[1999]), .CLK(clk), .RST(rst), .Q(sreg[1998]) );
  DFF \sreg_reg[1997]  ( .D(c[1998]), .CLK(clk), .RST(rst), .Q(sreg[1997]) );
  DFF \sreg_reg[1996]  ( .D(c[1997]), .CLK(clk), .RST(rst), .Q(sreg[1996]) );
  DFF \sreg_reg[1995]  ( .D(c[1996]), .CLK(clk), .RST(rst), .Q(sreg[1995]) );
  DFF \sreg_reg[1994]  ( .D(c[1995]), .CLK(clk), .RST(rst), .Q(sreg[1994]) );
  DFF \sreg_reg[1993]  ( .D(c[1994]), .CLK(clk), .RST(rst), .Q(sreg[1993]) );
  DFF \sreg_reg[1992]  ( .D(c[1993]), .CLK(clk), .RST(rst), .Q(sreg[1992]) );
  DFF \sreg_reg[1991]  ( .D(c[1992]), .CLK(clk), .RST(rst), .Q(sreg[1991]) );
  DFF \sreg_reg[1990]  ( .D(c[1991]), .CLK(clk), .RST(rst), .Q(sreg[1990]) );
  DFF \sreg_reg[1989]  ( .D(c[1990]), .CLK(clk), .RST(rst), .Q(sreg[1989]) );
  DFF \sreg_reg[1988]  ( .D(c[1989]), .CLK(clk), .RST(rst), .Q(sreg[1988]) );
  DFF \sreg_reg[1987]  ( .D(c[1988]), .CLK(clk), .RST(rst), .Q(sreg[1987]) );
  DFF \sreg_reg[1986]  ( .D(c[1987]), .CLK(clk), .RST(rst), .Q(sreg[1986]) );
  DFF \sreg_reg[1985]  ( .D(c[1986]), .CLK(clk), .RST(rst), .Q(sreg[1985]) );
  DFF \sreg_reg[1984]  ( .D(c[1985]), .CLK(clk), .RST(rst), .Q(sreg[1984]) );
  DFF \sreg_reg[1983]  ( .D(c[1984]), .CLK(clk), .RST(rst), .Q(sreg[1983]) );
  DFF \sreg_reg[1982]  ( .D(c[1983]), .CLK(clk), .RST(rst), .Q(sreg[1982]) );
  DFF \sreg_reg[1981]  ( .D(c[1982]), .CLK(clk), .RST(rst), .Q(sreg[1981]) );
  DFF \sreg_reg[1980]  ( .D(c[1981]), .CLK(clk), .RST(rst), .Q(sreg[1980]) );
  DFF \sreg_reg[1979]  ( .D(c[1980]), .CLK(clk), .RST(rst), .Q(sreg[1979]) );
  DFF \sreg_reg[1978]  ( .D(c[1979]), .CLK(clk), .RST(rst), .Q(sreg[1978]) );
  DFF \sreg_reg[1977]  ( .D(c[1978]), .CLK(clk), .RST(rst), .Q(sreg[1977]) );
  DFF \sreg_reg[1976]  ( .D(c[1977]), .CLK(clk), .RST(rst), .Q(sreg[1976]) );
  DFF \sreg_reg[1975]  ( .D(c[1976]), .CLK(clk), .RST(rst), .Q(sreg[1975]) );
  DFF \sreg_reg[1974]  ( .D(c[1975]), .CLK(clk), .RST(rst), .Q(sreg[1974]) );
  DFF \sreg_reg[1973]  ( .D(c[1974]), .CLK(clk), .RST(rst), .Q(sreg[1973]) );
  DFF \sreg_reg[1972]  ( .D(c[1973]), .CLK(clk), .RST(rst), .Q(sreg[1972]) );
  DFF \sreg_reg[1971]  ( .D(c[1972]), .CLK(clk), .RST(rst), .Q(sreg[1971]) );
  DFF \sreg_reg[1970]  ( .D(c[1971]), .CLK(clk), .RST(rst), .Q(sreg[1970]) );
  DFF \sreg_reg[1969]  ( .D(c[1970]), .CLK(clk), .RST(rst), .Q(sreg[1969]) );
  DFF \sreg_reg[1968]  ( .D(c[1969]), .CLK(clk), .RST(rst), .Q(sreg[1968]) );
  DFF \sreg_reg[1967]  ( .D(c[1968]), .CLK(clk), .RST(rst), .Q(sreg[1967]) );
  DFF \sreg_reg[1966]  ( .D(c[1967]), .CLK(clk), .RST(rst), .Q(sreg[1966]) );
  DFF \sreg_reg[1965]  ( .D(c[1966]), .CLK(clk), .RST(rst), .Q(sreg[1965]) );
  DFF \sreg_reg[1964]  ( .D(c[1965]), .CLK(clk), .RST(rst), .Q(sreg[1964]) );
  DFF \sreg_reg[1963]  ( .D(c[1964]), .CLK(clk), .RST(rst), .Q(sreg[1963]) );
  DFF \sreg_reg[1962]  ( .D(c[1963]), .CLK(clk), .RST(rst), .Q(sreg[1962]) );
  DFF \sreg_reg[1961]  ( .D(c[1962]), .CLK(clk), .RST(rst), .Q(sreg[1961]) );
  DFF \sreg_reg[1960]  ( .D(c[1961]), .CLK(clk), .RST(rst), .Q(sreg[1960]) );
  DFF \sreg_reg[1959]  ( .D(c[1960]), .CLK(clk), .RST(rst), .Q(sreg[1959]) );
  DFF \sreg_reg[1958]  ( .D(c[1959]), .CLK(clk), .RST(rst), .Q(sreg[1958]) );
  DFF \sreg_reg[1957]  ( .D(c[1958]), .CLK(clk), .RST(rst), .Q(sreg[1957]) );
  DFF \sreg_reg[1956]  ( .D(c[1957]), .CLK(clk), .RST(rst), .Q(sreg[1956]) );
  DFF \sreg_reg[1955]  ( .D(c[1956]), .CLK(clk), .RST(rst), .Q(sreg[1955]) );
  DFF \sreg_reg[1954]  ( .D(c[1955]), .CLK(clk), .RST(rst), .Q(sreg[1954]) );
  DFF \sreg_reg[1953]  ( .D(c[1954]), .CLK(clk), .RST(rst), .Q(sreg[1953]) );
  DFF \sreg_reg[1952]  ( .D(c[1953]), .CLK(clk), .RST(rst), .Q(sreg[1952]) );
  DFF \sreg_reg[1951]  ( .D(c[1952]), .CLK(clk), .RST(rst), .Q(sreg[1951]) );
  DFF \sreg_reg[1950]  ( .D(c[1951]), .CLK(clk), .RST(rst), .Q(sreg[1950]) );
  DFF \sreg_reg[1949]  ( .D(c[1950]), .CLK(clk), .RST(rst), .Q(sreg[1949]) );
  DFF \sreg_reg[1948]  ( .D(c[1949]), .CLK(clk), .RST(rst), .Q(sreg[1948]) );
  DFF \sreg_reg[1947]  ( .D(c[1948]), .CLK(clk), .RST(rst), .Q(sreg[1947]) );
  DFF \sreg_reg[1946]  ( .D(c[1947]), .CLK(clk), .RST(rst), .Q(sreg[1946]) );
  DFF \sreg_reg[1945]  ( .D(c[1946]), .CLK(clk), .RST(rst), .Q(sreg[1945]) );
  DFF \sreg_reg[1944]  ( .D(c[1945]), .CLK(clk), .RST(rst), .Q(sreg[1944]) );
  DFF \sreg_reg[1943]  ( .D(c[1944]), .CLK(clk), .RST(rst), .Q(sreg[1943]) );
  DFF \sreg_reg[1942]  ( .D(c[1943]), .CLK(clk), .RST(rst), .Q(sreg[1942]) );
  DFF \sreg_reg[1941]  ( .D(c[1942]), .CLK(clk), .RST(rst), .Q(sreg[1941]) );
  DFF \sreg_reg[1940]  ( .D(c[1941]), .CLK(clk), .RST(rst), .Q(sreg[1940]) );
  DFF \sreg_reg[1939]  ( .D(c[1940]), .CLK(clk), .RST(rst), .Q(sreg[1939]) );
  DFF \sreg_reg[1938]  ( .D(c[1939]), .CLK(clk), .RST(rst), .Q(sreg[1938]) );
  DFF \sreg_reg[1937]  ( .D(c[1938]), .CLK(clk), .RST(rst), .Q(sreg[1937]) );
  DFF \sreg_reg[1936]  ( .D(c[1937]), .CLK(clk), .RST(rst), .Q(sreg[1936]) );
  DFF \sreg_reg[1935]  ( .D(c[1936]), .CLK(clk), .RST(rst), .Q(sreg[1935]) );
  DFF \sreg_reg[1934]  ( .D(c[1935]), .CLK(clk), .RST(rst), .Q(sreg[1934]) );
  DFF \sreg_reg[1933]  ( .D(c[1934]), .CLK(clk), .RST(rst), .Q(sreg[1933]) );
  DFF \sreg_reg[1932]  ( .D(c[1933]), .CLK(clk), .RST(rst), .Q(sreg[1932]) );
  DFF \sreg_reg[1931]  ( .D(c[1932]), .CLK(clk), .RST(rst), .Q(sreg[1931]) );
  DFF \sreg_reg[1930]  ( .D(c[1931]), .CLK(clk), .RST(rst), .Q(sreg[1930]) );
  DFF \sreg_reg[1929]  ( .D(c[1930]), .CLK(clk), .RST(rst), .Q(sreg[1929]) );
  DFF \sreg_reg[1928]  ( .D(c[1929]), .CLK(clk), .RST(rst), .Q(sreg[1928]) );
  DFF \sreg_reg[1927]  ( .D(c[1928]), .CLK(clk), .RST(rst), .Q(sreg[1927]) );
  DFF \sreg_reg[1926]  ( .D(c[1927]), .CLK(clk), .RST(rst), .Q(sreg[1926]) );
  DFF \sreg_reg[1925]  ( .D(c[1926]), .CLK(clk), .RST(rst), .Q(sreg[1925]) );
  DFF \sreg_reg[1924]  ( .D(c[1925]), .CLK(clk), .RST(rst), .Q(sreg[1924]) );
  DFF \sreg_reg[1923]  ( .D(c[1924]), .CLK(clk), .RST(rst), .Q(sreg[1923]) );
  DFF \sreg_reg[1922]  ( .D(c[1923]), .CLK(clk), .RST(rst), .Q(sreg[1922]) );
  DFF \sreg_reg[1921]  ( .D(c[1922]), .CLK(clk), .RST(rst), .Q(sreg[1921]) );
  DFF \sreg_reg[1920]  ( .D(c[1921]), .CLK(clk), .RST(rst), .Q(sreg[1920]) );
  DFF \sreg_reg[1919]  ( .D(c[1920]), .CLK(clk), .RST(rst), .Q(sreg[1919]) );
  DFF \sreg_reg[1918]  ( .D(c[1919]), .CLK(clk), .RST(rst), .Q(sreg[1918]) );
  DFF \sreg_reg[1917]  ( .D(c[1918]), .CLK(clk), .RST(rst), .Q(sreg[1917]) );
  DFF \sreg_reg[1916]  ( .D(c[1917]), .CLK(clk), .RST(rst), .Q(sreg[1916]) );
  DFF \sreg_reg[1915]  ( .D(c[1916]), .CLK(clk), .RST(rst), .Q(sreg[1915]) );
  DFF \sreg_reg[1914]  ( .D(c[1915]), .CLK(clk), .RST(rst), .Q(sreg[1914]) );
  DFF \sreg_reg[1913]  ( .D(c[1914]), .CLK(clk), .RST(rst), .Q(sreg[1913]) );
  DFF \sreg_reg[1912]  ( .D(c[1913]), .CLK(clk), .RST(rst), .Q(sreg[1912]) );
  DFF \sreg_reg[1911]  ( .D(c[1912]), .CLK(clk), .RST(rst), .Q(sreg[1911]) );
  DFF \sreg_reg[1910]  ( .D(c[1911]), .CLK(clk), .RST(rst), .Q(sreg[1910]) );
  DFF \sreg_reg[1909]  ( .D(c[1910]), .CLK(clk), .RST(rst), .Q(sreg[1909]) );
  DFF \sreg_reg[1908]  ( .D(c[1909]), .CLK(clk), .RST(rst), .Q(sreg[1908]) );
  DFF \sreg_reg[1907]  ( .D(c[1908]), .CLK(clk), .RST(rst), .Q(sreg[1907]) );
  DFF \sreg_reg[1906]  ( .D(c[1907]), .CLK(clk), .RST(rst), .Q(sreg[1906]) );
  DFF \sreg_reg[1905]  ( .D(c[1906]), .CLK(clk), .RST(rst), .Q(sreg[1905]) );
  DFF \sreg_reg[1904]  ( .D(c[1905]), .CLK(clk), .RST(rst), .Q(sreg[1904]) );
  DFF \sreg_reg[1903]  ( .D(c[1904]), .CLK(clk), .RST(rst), .Q(sreg[1903]) );
  DFF \sreg_reg[1902]  ( .D(c[1903]), .CLK(clk), .RST(rst), .Q(sreg[1902]) );
  DFF \sreg_reg[1901]  ( .D(c[1902]), .CLK(clk), .RST(rst), .Q(sreg[1901]) );
  DFF \sreg_reg[1900]  ( .D(c[1901]), .CLK(clk), .RST(rst), .Q(sreg[1900]) );
  DFF \sreg_reg[1899]  ( .D(c[1900]), .CLK(clk), .RST(rst), .Q(sreg[1899]) );
  DFF \sreg_reg[1898]  ( .D(c[1899]), .CLK(clk), .RST(rst), .Q(sreg[1898]) );
  DFF \sreg_reg[1897]  ( .D(c[1898]), .CLK(clk), .RST(rst), .Q(sreg[1897]) );
  DFF \sreg_reg[1896]  ( .D(c[1897]), .CLK(clk), .RST(rst), .Q(sreg[1896]) );
  DFF \sreg_reg[1895]  ( .D(c[1896]), .CLK(clk), .RST(rst), .Q(sreg[1895]) );
  DFF \sreg_reg[1894]  ( .D(c[1895]), .CLK(clk), .RST(rst), .Q(sreg[1894]) );
  DFF \sreg_reg[1893]  ( .D(c[1894]), .CLK(clk), .RST(rst), .Q(sreg[1893]) );
  DFF \sreg_reg[1892]  ( .D(c[1893]), .CLK(clk), .RST(rst), .Q(sreg[1892]) );
  DFF \sreg_reg[1891]  ( .D(c[1892]), .CLK(clk), .RST(rst), .Q(sreg[1891]) );
  DFF \sreg_reg[1890]  ( .D(c[1891]), .CLK(clk), .RST(rst), .Q(sreg[1890]) );
  DFF \sreg_reg[1889]  ( .D(c[1890]), .CLK(clk), .RST(rst), .Q(sreg[1889]) );
  DFF \sreg_reg[1888]  ( .D(c[1889]), .CLK(clk), .RST(rst), .Q(sreg[1888]) );
  DFF \sreg_reg[1887]  ( .D(c[1888]), .CLK(clk), .RST(rst), .Q(sreg[1887]) );
  DFF \sreg_reg[1886]  ( .D(c[1887]), .CLK(clk), .RST(rst), .Q(sreg[1886]) );
  DFF \sreg_reg[1885]  ( .D(c[1886]), .CLK(clk), .RST(rst), .Q(sreg[1885]) );
  DFF \sreg_reg[1884]  ( .D(c[1885]), .CLK(clk), .RST(rst), .Q(sreg[1884]) );
  DFF \sreg_reg[1883]  ( .D(c[1884]), .CLK(clk), .RST(rst), .Q(sreg[1883]) );
  DFF \sreg_reg[1882]  ( .D(c[1883]), .CLK(clk), .RST(rst), .Q(sreg[1882]) );
  DFF \sreg_reg[1881]  ( .D(c[1882]), .CLK(clk), .RST(rst), .Q(sreg[1881]) );
  DFF \sreg_reg[1880]  ( .D(c[1881]), .CLK(clk), .RST(rst), .Q(sreg[1880]) );
  DFF \sreg_reg[1879]  ( .D(c[1880]), .CLK(clk), .RST(rst), .Q(sreg[1879]) );
  DFF \sreg_reg[1878]  ( .D(c[1879]), .CLK(clk), .RST(rst), .Q(sreg[1878]) );
  DFF \sreg_reg[1877]  ( .D(c[1878]), .CLK(clk), .RST(rst), .Q(sreg[1877]) );
  DFF \sreg_reg[1876]  ( .D(c[1877]), .CLK(clk), .RST(rst), .Q(sreg[1876]) );
  DFF \sreg_reg[1875]  ( .D(c[1876]), .CLK(clk), .RST(rst), .Q(sreg[1875]) );
  DFF \sreg_reg[1874]  ( .D(c[1875]), .CLK(clk), .RST(rst), .Q(sreg[1874]) );
  DFF \sreg_reg[1873]  ( .D(c[1874]), .CLK(clk), .RST(rst), .Q(sreg[1873]) );
  DFF \sreg_reg[1872]  ( .D(c[1873]), .CLK(clk), .RST(rst), .Q(sreg[1872]) );
  DFF \sreg_reg[1871]  ( .D(c[1872]), .CLK(clk), .RST(rst), .Q(sreg[1871]) );
  DFF \sreg_reg[1870]  ( .D(c[1871]), .CLK(clk), .RST(rst), .Q(sreg[1870]) );
  DFF \sreg_reg[1869]  ( .D(c[1870]), .CLK(clk), .RST(rst), .Q(sreg[1869]) );
  DFF \sreg_reg[1868]  ( .D(c[1869]), .CLK(clk), .RST(rst), .Q(sreg[1868]) );
  DFF \sreg_reg[1867]  ( .D(c[1868]), .CLK(clk), .RST(rst), .Q(sreg[1867]) );
  DFF \sreg_reg[1866]  ( .D(c[1867]), .CLK(clk), .RST(rst), .Q(sreg[1866]) );
  DFF \sreg_reg[1865]  ( .D(c[1866]), .CLK(clk), .RST(rst), .Q(sreg[1865]) );
  DFF \sreg_reg[1864]  ( .D(c[1865]), .CLK(clk), .RST(rst), .Q(sreg[1864]) );
  DFF \sreg_reg[1863]  ( .D(c[1864]), .CLK(clk), .RST(rst), .Q(sreg[1863]) );
  DFF \sreg_reg[1862]  ( .D(c[1863]), .CLK(clk), .RST(rst), .Q(sreg[1862]) );
  DFF \sreg_reg[1861]  ( .D(c[1862]), .CLK(clk), .RST(rst), .Q(sreg[1861]) );
  DFF \sreg_reg[1860]  ( .D(c[1861]), .CLK(clk), .RST(rst), .Q(sreg[1860]) );
  DFF \sreg_reg[1859]  ( .D(c[1860]), .CLK(clk), .RST(rst), .Q(sreg[1859]) );
  DFF \sreg_reg[1858]  ( .D(c[1859]), .CLK(clk), .RST(rst), .Q(sreg[1858]) );
  DFF \sreg_reg[1857]  ( .D(c[1858]), .CLK(clk), .RST(rst), .Q(sreg[1857]) );
  DFF \sreg_reg[1856]  ( .D(c[1857]), .CLK(clk), .RST(rst), .Q(sreg[1856]) );
  DFF \sreg_reg[1855]  ( .D(c[1856]), .CLK(clk), .RST(rst), .Q(sreg[1855]) );
  DFF \sreg_reg[1854]  ( .D(c[1855]), .CLK(clk), .RST(rst), .Q(sreg[1854]) );
  DFF \sreg_reg[1853]  ( .D(c[1854]), .CLK(clk), .RST(rst), .Q(sreg[1853]) );
  DFF \sreg_reg[1852]  ( .D(c[1853]), .CLK(clk), .RST(rst), .Q(sreg[1852]) );
  DFF \sreg_reg[1851]  ( .D(c[1852]), .CLK(clk), .RST(rst), .Q(sreg[1851]) );
  DFF \sreg_reg[1850]  ( .D(c[1851]), .CLK(clk), .RST(rst), .Q(sreg[1850]) );
  DFF \sreg_reg[1849]  ( .D(c[1850]), .CLK(clk), .RST(rst), .Q(sreg[1849]) );
  DFF \sreg_reg[1848]  ( .D(c[1849]), .CLK(clk), .RST(rst), .Q(sreg[1848]) );
  DFF \sreg_reg[1847]  ( .D(c[1848]), .CLK(clk), .RST(rst), .Q(sreg[1847]) );
  DFF \sreg_reg[1846]  ( .D(c[1847]), .CLK(clk), .RST(rst), .Q(sreg[1846]) );
  DFF \sreg_reg[1845]  ( .D(c[1846]), .CLK(clk), .RST(rst), .Q(sreg[1845]) );
  DFF \sreg_reg[1844]  ( .D(c[1845]), .CLK(clk), .RST(rst), .Q(sreg[1844]) );
  DFF \sreg_reg[1843]  ( .D(c[1844]), .CLK(clk), .RST(rst), .Q(sreg[1843]) );
  DFF \sreg_reg[1842]  ( .D(c[1843]), .CLK(clk), .RST(rst), .Q(sreg[1842]) );
  DFF \sreg_reg[1841]  ( .D(c[1842]), .CLK(clk), .RST(rst), .Q(sreg[1841]) );
  DFF \sreg_reg[1840]  ( .D(c[1841]), .CLK(clk), .RST(rst), .Q(sreg[1840]) );
  DFF \sreg_reg[1839]  ( .D(c[1840]), .CLK(clk), .RST(rst), .Q(sreg[1839]) );
  DFF \sreg_reg[1838]  ( .D(c[1839]), .CLK(clk), .RST(rst), .Q(sreg[1838]) );
  DFF \sreg_reg[1837]  ( .D(c[1838]), .CLK(clk), .RST(rst), .Q(sreg[1837]) );
  DFF \sreg_reg[1836]  ( .D(c[1837]), .CLK(clk), .RST(rst), .Q(sreg[1836]) );
  DFF \sreg_reg[1835]  ( .D(c[1836]), .CLK(clk), .RST(rst), .Q(sreg[1835]) );
  DFF \sreg_reg[1834]  ( .D(c[1835]), .CLK(clk), .RST(rst), .Q(sreg[1834]) );
  DFF \sreg_reg[1833]  ( .D(c[1834]), .CLK(clk), .RST(rst), .Q(sreg[1833]) );
  DFF \sreg_reg[1832]  ( .D(c[1833]), .CLK(clk), .RST(rst), .Q(sreg[1832]) );
  DFF \sreg_reg[1831]  ( .D(c[1832]), .CLK(clk), .RST(rst), .Q(sreg[1831]) );
  DFF \sreg_reg[1830]  ( .D(c[1831]), .CLK(clk), .RST(rst), .Q(sreg[1830]) );
  DFF \sreg_reg[1829]  ( .D(c[1830]), .CLK(clk), .RST(rst), .Q(sreg[1829]) );
  DFF \sreg_reg[1828]  ( .D(c[1829]), .CLK(clk), .RST(rst), .Q(sreg[1828]) );
  DFF \sreg_reg[1827]  ( .D(c[1828]), .CLK(clk), .RST(rst), .Q(sreg[1827]) );
  DFF \sreg_reg[1826]  ( .D(c[1827]), .CLK(clk), .RST(rst), .Q(sreg[1826]) );
  DFF \sreg_reg[1825]  ( .D(c[1826]), .CLK(clk), .RST(rst), .Q(sreg[1825]) );
  DFF \sreg_reg[1824]  ( .D(c[1825]), .CLK(clk), .RST(rst), .Q(sreg[1824]) );
  DFF \sreg_reg[1823]  ( .D(c[1824]), .CLK(clk), .RST(rst), .Q(sreg[1823]) );
  DFF \sreg_reg[1822]  ( .D(c[1823]), .CLK(clk), .RST(rst), .Q(sreg[1822]) );
  DFF \sreg_reg[1821]  ( .D(c[1822]), .CLK(clk), .RST(rst), .Q(sreg[1821]) );
  DFF \sreg_reg[1820]  ( .D(c[1821]), .CLK(clk), .RST(rst), .Q(sreg[1820]) );
  DFF \sreg_reg[1819]  ( .D(c[1820]), .CLK(clk), .RST(rst), .Q(sreg[1819]) );
  DFF \sreg_reg[1818]  ( .D(c[1819]), .CLK(clk), .RST(rst), .Q(sreg[1818]) );
  DFF \sreg_reg[1817]  ( .D(c[1818]), .CLK(clk), .RST(rst), .Q(sreg[1817]) );
  DFF \sreg_reg[1816]  ( .D(c[1817]), .CLK(clk), .RST(rst), .Q(sreg[1816]) );
  DFF \sreg_reg[1815]  ( .D(c[1816]), .CLK(clk), .RST(rst), .Q(sreg[1815]) );
  DFF \sreg_reg[1814]  ( .D(c[1815]), .CLK(clk), .RST(rst), .Q(sreg[1814]) );
  DFF \sreg_reg[1813]  ( .D(c[1814]), .CLK(clk), .RST(rst), .Q(sreg[1813]) );
  DFF \sreg_reg[1812]  ( .D(c[1813]), .CLK(clk), .RST(rst), .Q(sreg[1812]) );
  DFF \sreg_reg[1811]  ( .D(c[1812]), .CLK(clk), .RST(rst), .Q(sreg[1811]) );
  DFF \sreg_reg[1810]  ( .D(c[1811]), .CLK(clk), .RST(rst), .Q(sreg[1810]) );
  DFF \sreg_reg[1809]  ( .D(c[1810]), .CLK(clk), .RST(rst), .Q(sreg[1809]) );
  DFF \sreg_reg[1808]  ( .D(c[1809]), .CLK(clk), .RST(rst), .Q(sreg[1808]) );
  DFF \sreg_reg[1807]  ( .D(c[1808]), .CLK(clk), .RST(rst), .Q(sreg[1807]) );
  DFF \sreg_reg[1806]  ( .D(c[1807]), .CLK(clk), .RST(rst), .Q(sreg[1806]) );
  DFF \sreg_reg[1805]  ( .D(c[1806]), .CLK(clk), .RST(rst), .Q(sreg[1805]) );
  DFF \sreg_reg[1804]  ( .D(c[1805]), .CLK(clk), .RST(rst), .Q(sreg[1804]) );
  DFF \sreg_reg[1803]  ( .D(c[1804]), .CLK(clk), .RST(rst), .Q(sreg[1803]) );
  DFF \sreg_reg[1802]  ( .D(c[1803]), .CLK(clk), .RST(rst), .Q(sreg[1802]) );
  DFF \sreg_reg[1801]  ( .D(c[1802]), .CLK(clk), .RST(rst), .Q(sreg[1801]) );
  DFF \sreg_reg[1800]  ( .D(c[1801]), .CLK(clk), .RST(rst), .Q(sreg[1800]) );
  DFF \sreg_reg[1799]  ( .D(c[1800]), .CLK(clk), .RST(rst), .Q(sreg[1799]) );
  DFF \sreg_reg[1798]  ( .D(c[1799]), .CLK(clk), .RST(rst), .Q(sreg[1798]) );
  DFF \sreg_reg[1797]  ( .D(c[1798]), .CLK(clk), .RST(rst), .Q(sreg[1797]) );
  DFF \sreg_reg[1796]  ( .D(c[1797]), .CLK(clk), .RST(rst), .Q(sreg[1796]) );
  DFF \sreg_reg[1795]  ( .D(c[1796]), .CLK(clk), .RST(rst), .Q(sreg[1795]) );
  DFF \sreg_reg[1794]  ( .D(c[1795]), .CLK(clk), .RST(rst), .Q(sreg[1794]) );
  DFF \sreg_reg[1793]  ( .D(c[1794]), .CLK(clk), .RST(rst), .Q(sreg[1793]) );
  DFF \sreg_reg[1792]  ( .D(c[1793]), .CLK(clk), .RST(rst), .Q(sreg[1792]) );
  DFF \sreg_reg[1791]  ( .D(c[1792]), .CLK(clk), .RST(rst), .Q(sreg[1791]) );
  DFF \sreg_reg[1790]  ( .D(c[1791]), .CLK(clk), .RST(rst), .Q(sreg[1790]) );
  DFF \sreg_reg[1789]  ( .D(c[1790]), .CLK(clk), .RST(rst), .Q(sreg[1789]) );
  DFF \sreg_reg[1788]  ( .D(c[1789]), .CLK(clk), .RST(rst), .Q(sreg[1788]) );
  DFF \sreg_reg[1787]  ( .D(c[1788]), .CLK(clk), .RST(rst), .Q(sreg[1787]) );
  DFF \sreg_reg[1786]  ( .D(c[1787]), .CLK(clk), .RST(rst), .Q(sreg[1786]) );
  DFF \sreg_reg[1785]  ( .D(c[1786]), .CLK(clk), .RST(rst), .Q(sreg[1785]) );
  DFF \sreg_reg[1784]  ( .D(c[1785]), .CLK(clk), .RST(rst), .Q(sreg[1784]) );
  DFF \sreg_reg[1783]  ( .D(c[1784]), .CLK(clk), .RST(rst), .Q(sreg[1783]) );
  DFF \sreg_reg[1782]  ( .D(c[1783]), .CLK(clk), .RST(rst), .Q(sreg[1782]) );
  DFF \sreg_reg[1781]  ( .D(c[1782]), .CLK(clk), .RST(rst), .Q(sreg[1781]) );
  DFF \sreg_reg[1780]  ( .D(c[1781]), .CLK(clk), .RST(rst), .Q(sreg[1780]) );
  DFF \sreg_reg[1779]  ( .D(c[1780]), .CLK(clk), .RST(rst), .Q(sreg[1779]) );
  DFF \sreg_reg[1778]  ( .D(c[1779]), .CLK(clk), .RST(rst), .Q(sreg[1778]) );
  DFF \sreg_reg[1777]  ( .D(c[1778]), .CLK(clk), .RST(rst), .Q(sreg[1777]) );
  DFF \sreg_reg[1776]  ( .D(c[1777]), .CLK(clk), .RST(rst), .Q(sreg[1776]) );
  DFF \sreg_reg[1775]  ( .D(c[1776]), .CLK(clk), .RST(rst), .Q(sreg[1775]) );
  DFF \sreg_reg[1774]  ( .D(c[1775]), .CLK(clk), .RST(rst), .Q(sreg[1774]) );
  DFF \sreg_reg[1773]  ( .D(c[1774]), .CLK(clk), .RST(rst), .Q(sreg[1773]) );
  DFF \sreg_reg[1772]  ( .D(c[1773]), .CLK(clk), .RST(rst), .Q(sreg[1772]) );
  DFF \sreg_reg[1771]  ( .D(c[1772]), .CLK(clk), .RST(rst), .Q(sreg[1771]) );
  DFF \sreg_reg[1770]  ( .D(c[1771]), .CLK(clk), .RST(rst), .Q(sreg[1770]) );
  DFF \sreg_reg[1769]  ( .D(c[1770]), .CLK(clk), .RST(rst), .Q(sreg[1769]) );
  DFF \sreg_reg[1768]  ( .D(c[1769]), .CLK(clk), .RST(rst), .Q(sreg[1768]) );
  DFF \sreg_reg[1767]  ( .D(c[1768]), .CLK(clk), .RST(rst), .Q(sreg[1767]) );
  DFF \sreg_reg[1766]  ( .D(c[1767]), .CLK(clk), .RST(rst), .Q(sreg[1766]) );
  DFF \sreg_reg[1765]  ( .D(c[1766]), .CLK(clk), .RST(rst), .Q(sreg[1765]) );
  DFF \sreg_reg[1764]  ( .D(c[1765]), .CLK(clk), .RST(rst), .Q(sreg[1764]) );
  DFF \sreg_reg[1763]  ( .D(c[1764]), .CLK(clk), .RST(rst), .Q(sreg[1763]) );
  DFF \sreg_reg[1762]  ( .D(c[1763]), .CLK(clk), .RST(rst), .Q(sreg[1762]) );
  DFF \sreg_reg[1761]  ( .D(c[1762]), .CLK(clk), .RST(rst), .Q(sreg[1761]) );
  DFF \sreg_reg[1760]  ( .D(c[1761]), .CLK(clk), .RST(rst), .Q(sreg[1760]) );
  DFF \sreg_reg[1759]  ( .D(c[1760]), .CLK(clk), .RST(rst), .Q(sreg[1759]) );
  DFF \sreg_reg[1758]  ( .D(c[1759]), .CLK(clk), .RST(rst), .Q(sreg[1758]) );
  DFF \sreg_reg[1757]  ( .D(c[1758]), .CLK(clk), .RST(rst), .Q(sreg[1757]) );
  DFF \sreg_reg[1756]  ( .D(c[1757]), .CLK(clk), .RST(rst), .Q(sreg[1756]) );
  DFF \sreg_reg[1755]  ( .D(c[1756]), .CLK(clk), .RST(rst), .Q(sreg[1755]) );
  DFF \sreg_reg[1754]  ( .D(c[1755]), .CLK(clk), .RST(rst), .Q(sreg[1754]) );
  DFF \sreg_reg[1753]  ( .D(c[1754]), .CLK(clk), .RST(rst), .Q(sreg[1753]) );
  DFF \sreg_reg[1752]  ( .D(c[1753]), .CLK(clk), .RST(rst), .Q(sreg[1752]) );
  DFF \sreg_reg[1751]  ( .D(c[1752]), .CLK(clk), .RST(rst), .Q(sreg[1751]) );
  DFF \sreg_reg[1750]  ( .D(c[1751]), .CLK(clk), .RST(rst), .Q(sreg[1750]) );
  DFF \sreg_reg[1749]  ( .D(c[1750]), .CLK(clk), .RST(rst), .Q(sreg[1749]) );
  DFF \sreg_reg[1748]  ( .D(c[1749]), .CLK(clk), .RST(rst), .Q(sreg[1748]) );
  DFF \sreg_reg[1747]  ( .D(c[1748]), .CLK(clk), .RST(rst), .Q(sreg[1747]) );
  DFF \sreg_reg[1746]  ( .D(c[1747]), .CLK(clk), .RST(rst), .Q(sreg[1746]) );
  DFF \sreg_reg[1745]  ( .D(c[1746]), .CLK(clk), .RST(rst), .Q(sreg[1745]) );
  DFF \sreg_reg[1744]  ( .D(c[1745]), .CLK(clk), .RST(rst), .Q(sreg[1744]) );
  DFF \sreg_reg[1743]  ( .D(c[1744]), .CLK(clk), .RST(rst), .Q(sreg[1743]) );
  DFF \sreg_reg[1742]  ( .D(c[1743]), .CLK(clk), .RST(rst), .Q(sreg[1742]) );
  DFF \sreg_reg[1741]  ( .D(c[1742]), .CLK(clk), .RST(rst), .Q(sreg[1741]) );
  DFF \sreg_reg[1740]  ( .D(c[1741]), .CLK(clk), .RST(rst), .Q(sreg[1740]) );
  DFF \sreg_reg[1739]  ( .D(c[1740]), .CLK(clk), .RST(rst), .Q(sreg[1739]) );
  DFF \sreg_reg[1738]  ( .D(c[1739]), .CLK(clk), .RST(rst), .Q(sreg[1738]) );
  DFF \sreg_reg[1737]  ( .D(c[1738]), .CLK(clk), .RST(rst), .Q(sreg[1737]) );
  DFF \sreg_reg[1736]  ( .D(c[1737]), .CLK(clk), .RST(rst), .Q(sreg[1736]) );
  DFF \sreg_reg[1735]  ( .D(c[1736]), .CLK(clk), .RST(rst), .Q(sreg[1735]) );
  DFF \sreg_reg[1734]  ( .D(c[1735]), .CLK(clk), .RST(rst), .Q(sreg[1734]) );
  DFF \sreg_reg[1733]  ( .D(c[1734]), .CLK(clk), .RST(rst), .Q(sreg[1733]) );
  DFF \sreg_reg[1732]  ( .D(c[1733]), .CLK(clk), .RST(rst), .Q(sreg[1732]) );
  DFF \sreg_reg[1731]  ( .D(c[1732]), .CLK(clk), .RST(rst), .Q(sreg[1731]) );
  DFF \sreg_reg[1730]  ( .D(c[1731]), .CLK(clk), .RST(rst), .Q(sreg[1730]) );
  DFF \sreg_reg[1729]  ( .D(c[1730]), .CLK(clk), .RST(rst), .Q(sreg[1729]) );
  DFF \sreg_reg[1728]  ( .D(c[1729]), .CLK(clk), .RST(rst), .Q(sreg[1728]) );
  DFF \sreg_reg[1727]  ( .D(c[1728]), .CLK(clk), .RST(rst), .Q(sreg[1727]) );
  DFF \sreg_reg[1726]  ( .D(c[1727]), .CLK(clk), .RST(rst), .Q(sreg[1726]) );
  DFF \sreg_reg[1725]  ( .D(c[1726]), .CLK(clk), .RST(rst), .Q(sreg[1725]) );
  DFF \sreg_reg[1724]  ( .D(c[1725]), .CLK(clk), .RST(rst), .Q(sreg[1724]) );
  DFF \sreg_reg[1723]  ( .D(c[1724]), .CLK(clk), .RST(rst), .Q(sreg[1723]) );
  DFF \sreg_reg[1722]  ( .D(c[1723]), .CLK(clk), .RST(rst), .Q(sreg[1722]) );
  DFF \sreg_reg[1721]  ( .D(c[1722]), .CLK(clk), .RST(rst), .Q(sreg[1721]) );
  DFF \sreg_reg[1720]  ( .D(c[1721]), .CLK(clk), .RST(rst), .Q(sreg[1720]) );
  DFF \sreg_reg[1719]  ( .D(c[1720]), .CLK(clk), .RST(rst), .Q(sreg[1719]) );
  DFF \sreg_reg[1718]  ( .D(c[1719]), .CLK(clk), .RST(rst), .Q(sreg[1718]) );
  DFF \sreg_reg[1717]  ( .D(c[1718]), .CLK(clk), .RST(rst), .Q(sreg[1717]) );
  DFF \sreg_reg[1716]  ( .D(c[1717]), .CLK(clk), .RST(rst), .Q(sreg[1716]) );
  DFF \sreg_reg[1715]  ( .D(c[1716]), .CLK(clk), .RST(rst), .Q(sreg[1715]) );
  DFF \sreg_reg[1714]  ( .D(c[1715]), .CLK(clk), .RST(rst), .Q(sreg[1714]) );
  DFF \sreg_reg[1713]  ( .D(c[1714]), .CLK(clk), .RST(rst), .Q(sreg[1713]) );
  DFF \sreg_reg[1712]  ( .D(c[1713]), .CLK(clk), .RST(rst), .Q(sreg[1712]) );
  DFF \sreg_reg[1711]  ( .D(c[1712]), .CLK(clk), .RST(rst), .Q(sreg[1711]) );
  DFF \sreg_reg[1710]  ( .D(c[1711]), .CLK(clk), .RST(rst), .Q(sreg[1710]) );
  DFF \sreg_reg[1709]  ( .D(c[1710]), .CLK(clk), .RST(rst), .Q(sreg[1709]) );
  DFF \sreg_reg[1708]  ( .D(c[1709]), .CLK(clk), .RST(rst), .Q(sreg[1708]) );
  DFF \sreg_reg[1707]  ( .D(c[1708]), .CLK(clk), .RST(rst), .Q(sreg[1707]) );
  DFF \sreg_reg[1706]  ( .D(c[1707]), .CLK(clk), .RST(rst), .Q(sreg[1706]) );
  DFF \sreg_reg[1705]  ( .D(c[1706]), .CLK(clk), .RST(rst), .Q(sreg[1705]) );
  DFF \sreg_reg[1704]  ( .D(c[1705]), .CLK(clk), .RST(rst), .Q(sreg[1704]) );
  DFF \sreg_reg[1703]  ( .D(c[1704]), .CLK(clk), .RST(rst), .Q(sreg[1703]) );
  DFF \sreg_reg[1702]  ( .D(c[1703]), .CLK(clk), .RST(rst), .Q(sreg[1702]) );
  DFF \sreg_reg[1701]  ( .D(c[1702]), .CLK(clk), .RST(rst), .Q(sreg[1701]) );
  DFF \sreg_reg[1700]  ( .D(c[1701]), .CLK(clk), .RST(rst), .Q(sreg[1700]) );
  DFF \sreg_reg[1699]  ( .D(c[1700]), .CLK(clk), .RST(rst), .Q(sreg[1699]) );
  DFF \sreg_reg[1698]  ( .D(c[1699]), .CLK(clk), .RST(rst), .Q(sreg[1698]) );
  DFF \sreg_reg[1697]  ( .D(c[1698]), .CLK(clk), .RST(rst), .Q(sreg[1697]) );
  DFF \sreg_reg[1696]  ( .D(c[1697]), .CLK(clk), .RST(rst), .Q(sreg[1696]) );
  DFF \sreg_reg[1695]  ( .D(c[1696]), .CLK(clk), .RST(rst), .Q(sreg[1695]) );
  DFF \sreg_reg[1694]  ( .D(c[1695]), .CLK(clk), .RST(rst), .Q(sreg[1694]) );
  DFF \sreg_reg[1693]  ( .D(c[1694]), .CLK(clk), .RST(rst), .Q(sreg[1693]) );
  DFF \sreg_reg[1692]  ( .D(c[1693]), .CLK(clk), .RST(rst), .Q(sreg[1692]) );
  DFF \sreg_reg[1691]  ( .D(c[1692]), .CLK(clk), .RST(rst), .Q(sreg[1691]) );
  DFF \sreg_reg[1690]  ( .D(c[1691]), .CLK(clk), .RST(rst), .Q(sreg[1690]) );
  DFF \sreg_reg[1689]  ( .D(c[1690]), .CLK(clk), .RST(rst), .Q(sreg[1689]) );
  DFF \sreg_reg[1688]  ( .D(c[1689]), .CLK(clk), .RST(rst), .Q(sreg[1688]) );
  DFF \sreg_reg[1687]  ( .D(c[1688]), .CLK(clk), .RST(rst), .Q(sreg[1687]) );
  DFF \sreg_reg[1686]  ( .D(c[1687]), .CLK(clk), .RST(rst), .Q(sreg[1686]) );
  DFF \sreg_reg[1685]  ( .D(c[1686]), .CLK(clk), .RST(rst), .Q(sreg[1685]) );
  DFF \sreg_reg[1684]  ( .D(c[1685]), .CLK(clk), .RST(rst), .Q(sreg[1684]) );
  DFF \sreg_reg[1683]  ( .D(c[1684]), .CLK(clk), .RST(rst), .Q(sreg[1683]) );
  DFF \sreg_reg[1682]  ( .D(c[1683]), .CLK(clk), .RST(rst), .Q(sreg[1682]) );
  DFF \sreg_reg[1681]  ( .D(c[1682]), .CLK(clk), .RST(rst), .Q(sreg[1681]) );
  DFF \sreg_reg[1680]  ( .D(c[1681]), .CLK(clk), .RST(rst), .Q(sreg[1680]) );
  DFF \sreg_reg[1679]  ( .D(c[1680]), .CLK(clk), .RST(rst), .Q(sreg[1679]) );
  DFF \sreg_reg[1678]  ( .D(c[1679]), .CLK(clk), .RST(rst), .Q(sreg[1678]) );
  DFF \sreg_reg[1677]  ( .D(c[1678]), .CLK(clk), .RST(rst), .Q(sreg[1677]) );
  DFF \sreg_reg[1676]  ( .D(c[1677]), .CLK(clk), .RST(rst), .Q(sreg[1676]) );
  DFF \sreg_reg[1675]  ( .D(c[1676]), .CLK(clk), .RST(rst), .Q(sreg[1675]) );
  DFF \sreg_reg[1674]  ( .D(c[1675]), .CLK(clk), .RST(rst), .Q(sreg[1674]) );
  DFF \sreg_reg[1673]  ( .D(c[1674]), .CLK(clk), .RST(rst), .Q(sreg[1673]) );
  DFF \sreg_reg[1672]  ( .D(c[1673]), .CLK(clk), .RST(rst), .Q(sreg[1672]) );
  DFF \sreg_reg[1671]  ( .D(c[1672]), .CLK(clk), .RST(rst), .Q(sreg[1671]) );
  DFF \sreg_reg[1670]  ( .D(c[1671]), .CLK(clk), .RST(rst), .Q(sreg[1670]) );
  DFF \sreg_reg[1669]  ( .D(c[1670]), .CLK(clk), .RST(rst), .Q(sreg[1669]) );
  DFF \sreg_reg[1668]  ( .D(c[1669]), .CLK(clk), .RST(rst), .Q(sreg[1668]) );
  DFF \sreg_reg[1667]  ( .D(c[1668]), .CLK(clk), .RST(rst), .Q(sreg[1667]) );
  DFF \sreg_reg[1666]  ( .D(c[1667]), .CLK(clk), .RST(rst), .Q(sreg[1666]) );
  DFF \sreg_reg[1665]  ( .D(c[1666]), .CLK(clk), .RST(rst), .Q(sreg[1665]) );
  DFF \sreg_reg[1664]  ( .D(c[1665]), .CLK(clk), .RST(rst), .Q(sreg[1664]) );
  DFF \sreg_reg[1663]  ( .D(c[1664]), .CLK(clk), .RST(rst), .Q(sreg[1663]) );
  DFF \sreg_reg[1662]  ( .D(c[1663]), .CLK(clk), .RST(rst), .Q(sreg[1662]) );
  DFF \sreg_reg[1661]  ( .D(c[1662]), .CLK(clk), .RST(rst), .Q(sreg[1661]) );
  DFF \sreg_reg[1660]  ( .D(c[1661]), .CLK(clk), .RST(rst), .Q(sreg[1660]) );
  DFF \sreg_reg[1659]  ( .D(c[1660]), .CLK(clk), .RST(rst), .Q(sreg[1659]) );
  DFF \sreg_reg[1658]  ( .D(c[1659]), .CLK(clk), .RST(rst), .Q(sreg[1658]) );
  DFF \sreg_reg[1657]  ( .D(c[1658]), .CLK(clk), .RST(rst), .Q(sreg[1657]) );
  DFF \sreg_reg[1656]  ( .D(c[1657]), .CLK(clk), .RST(rst), .Q(sreg[1656]) );
  DFF \sreg_reg[1655]  ( .D(c[1656]), .CLK(clk), .RST(rst), .Q(sreg[1655]) );
  DFF \sreg_reg[1654]  ( .D(c[1655]), .CLK(clk), .RST(rst), .Q(sreg[1654]) );
  DFF \sreg_reg[1653]  ( .D(c[1654]), .CLK(clk), .RST(rst), .Q(sreg[1653]) );
  DFF \sreg_reg[1652]  ( .D(c[1653]), .CLK(clk), .RST(rst), .Q(sreg[1652]) );
  DFF \sreg_reg[1651]  ( .D(c[1652]), .CLK(clk), .RST(rst), .Q(sreg[1651]) );
  DFF \sreg_reg[1650]  ( .D(c[1651]), .CLK(clk), .RST(rst), .Q(sreg[1650]) );
  DFF \sreg_reg[1649]  ( .D(c[1650]), .CLK(clk), .RST(rst), .Q(sreg[1649]) );
  DFF \sreg_reg[1648]  ( .D(c[1649]), .CLK(clk), .RST(rst), .Q(sreg[1648]) );
  DFF \sreg_reg[1647]  ( .D(c[1648]), .CLK(clk), .RST(rst), .Q(sreg[1647]) );
  DFF \sreg_reg[1646]  ( .D(c[1647]), .CLK(clk), .RST(rst), .Q(sreg[1646]) );
  DFF \sreg_reg[1645]  ( .D(c[1646]), .CLK(clk), .RST(rst), .Q(sreg[1645]) );
  DFF \sreg_reg[1644]  ( .D(c[1645]), .CLK(clk), .RST(rst), .Q(sreg[1644]) );
  DFF \sreg_reg[1643]  ( .D(c[1644]), .CLK(clk), .RST(rst), .Q(sreg[1643]) );
  DFF \sreg_reg[1642]  ( .D(c[1643]), .CLK(clk), .RST(rst), .Q(sreg[1642]) );
  DFF \sreg_reg[1641]  ( .D(c[1642]), .CLK(clk), .RST(rst), .Q(sreg[1641]) );
  DFF \sreg_reg[1640]  ( .D(c[1641]), .CLK(clk), .RST(rst), .Q(sreg[1640]) );
  DFF \sreg_reg[1639]  ( .D(c[1640]), .CLK(clk), .RST(rst), .Q(sreg[1639]) );
  DFF \sreg_reg[1638]  ( .D(c[1639]), .CLK(clk), .RST(rst), .Q(sreg[1638]) );
  DFF \sreg_reg[1637]  ( .D(c[1638]), .CLK(clk), .RST(rst), .Q(sreg[1637]) );
  DFF \sreg_reg[1636]  ( .D(c[1637]), .CLK(clk), .RST(rst), .Q(sreg[1636]) );
  DFF \sreg_reg[1635]  ( .D(c[1636]), .CLK(clk), .RST(rst), .Q(sreg[1635]) );
  DFF \sreg_reg[1634]  ( .D(c[1635]), .CLK(clk), .RST(rst), .Q(sreg[1634]) );
  DFF \sreg_reg[1633]  ( .D(c[1634]), .CLK(clk), .RST(rst), .Q(sreg[1633]) );
  DFF \sreg_reg[1632]  ( .D(c[1633]), .CLK(clk), .RST(rst), .Q(sreg[1632]) );
  DFF \sreg_reg[1631]  ( .D(c[1632]), .CLK(clk), .RST(rst), .Q(sreg[1631]) );
  DFF \sreg_reg[1630]  ( .D(c[1631]), .CLK(clk), .RST(rst), .Q(sreg[1630]) );
  DFF \sreg_reg[1629]  ( .D(c[1630]), .CLK(clk), .RST(rst), .Q(sreg[1629]) );
  DFF \sreg_reg[1628]  ( .D(c[1629]), .CLK(clk), .RST(rst), .Q(sreg[1628]) );
  DFF \sreg_reg[1627]  ( .D(c[1628]), .CLK(clk), .RST(rst), .Q(sreg[1627]) );
  DFF \sreg_reg[1626]  ( .D(c[1627]), .CLK(clk), .RST(rst), .Q(sreg[1626]) );
  DFF \sreg_reg[1625]  ( .D(c[1626]), .CLK(clk), .RST(rst), .Q(sreg[1625]) );
  DFF \sreg_reg[1624]  ( .D(c[1625]), .CLK(clk), .RST(rst), .Q(sreg[1624]) );
  DFF \sreg_reg[1623]  ( .D(c[1624]), .CLK(clk), .RST(rst), .Q(sreg[1623]) );
  DFF \sreg_reg[1622]  ( .D(c[1623]), .CLK(clk), .RST(rst), .Q(sreg[1622]) );
  DFF \sreg_reg[1621]  ( .D(c[1622]), .CLK(clk), .RST(rst), .Q(sreg[1621]) );
  DFF \sreg_reg[1620]  ( .D(c[1621]), .CLK(clk), .RST(rst), .Q(sreg[1620]) );
  DFF \sreg_reg[1619]  ( .D(c[1620]), .CLK(clk), .RST(rst), .Q(sreg[1619]) );
  DFF \sreg_reg[1618]  ( .D(c[1619]), .CLK(clk), .RST(rst), .Q(sreg[1618]) );
  DFF \sreg_reg[1617]  ( .D(c[1618]), .CLK(clk), .RST(rst), .Q(sreg[1617]) );
  DFF \sreg_reg[1616]  ( .D(c[1617]), .CLK(clk), .RST(rst), .Q(sreg[1616]) );
  DFF \sreg_reg[1615]  ( .D(c[1616]), .CLK(clk), .RST(rst), .Q(sreg[1615]) );
  DFF \sreg_reg[1614]  ( .D(c[1615]), .CLK(clk), .RST(rst), .Q(sreg[1614]) );
  DFF \sreg_reg[1613]  ( .D(c[1614]), .CLK(clk), .RST(rst), .Q(sreg[1613]) );
  DFF \sreg_reg[1612]  ( .D(c[1613]), .CLK(clk), .RST(rst), .Q(sreg[1612]) );
  DFF \sreg_reg[1611]  ( .D(c[1612]), .CLK(clk), .RST(rst), .Q(sreg[1611]) );
  DFF \sreg_reg[1610]  ( .D(c[1611]), .CLK(clk), .RST(rst), .Q(sreg[1610]) );
  DFF \sreg_reg[1609]  ( .D(c[1610]), .CLK(clk), .RST(rst), .Q(sreg[1609]) );
  DFF \sreg_reg[1608]  ( .D(c[1609]), .CLK(clk), .RST(rst), .Q(sreg[1608]) );
  DFF \sreg_reg[1607]  ( .D(c[1608]), .CLK(clk), .RST(rst), .Q(sreg[1607]) );
  DFF \sreg_reg[1606]  ( .D(c[1607]), .CLK(clk), .RST(rst), .Q(sreg[1606]) );
  DFF \sreg_reg[1605]  ( .D(c[1606]), .CLK(clk), .RST(rst), .Q(sreg[1605]) );
  DFF \sreg_reg[1604]  ( .D(c[1605]), .CLK(clk), .RST(rst), .Q(sreg[1604]) );
  DFF \sreg_reg[1603]  ( .D(c[1604]), .CLK(clk), .RST(rst), .Q(sreg[1603]) );
  DFF \sreg_reg[1602]  ( .D(c[1603]), .CLK(clk), .RST(rst), .Q(sreg[1602]) );
  DFF \sreg_reg[1601]  ( .D(c[1602]), .CLK(clk), .RST(rst), .Q(sreg[1601]) );
  DFF \sreg_reg[1600]  ( .D(c[1601]), .CLK(clk), .RST(rst), .Q(sreg[1600]) );
  DFF \sreg_reg[1599]  ( .D(c[1600]), .CLK(clk), .RST(rst), .Q(sreg[1599]) );
  DFF \sreg_reg[1598]  ( .D(c[1599]), .CLK(clk), .RST(rst), .Q(sreg[1598]) );
  DFF \sreg_reg[1597]  ( .D(c[1598]), .CLK(clk), .RST(rst), .Q(sreg[1597]) );
  DFF \sreg_reg[1596]  ( .D(c[1597]), .CLK(clk), .RST(rst), .Q(sreg[1596]) );
  DFF \sreg_reg[1595]  ( .D(c[1596]), .CLK(clk), .RST(rst), .Q(sreg[1595]) );
  DFF \sreg_reg[1594]  ( .D(c[1595]), .CLK(clk), .RST(rst), .Q(sreg[1594]) );
  DFF \sreg_reg[1593]  ( .D(c[1594]), .CLK(clk), .RST(rst), .Q(sreg[1593]) );
  DFF \sreg_reg[1592]  ( .D(c[1593]), .CLK(clk), .RST(rst), .Q(sreg[1592]) );
  DFF \sreg_reg[1591]  ( .D(c[1592]), .CLK(clk), .RST(rst), .Q(sreg[1591]) );
  DFF \sreg_reg[1590]  ( .D(c[1591]), .CLK(clk), .RST(rst), .Q(sreg[1590]) );
  DFF \sreg_reg[1589]  ( .D(c[1590]), .CLK(clk), .RST(rst), .Q(sreg[1589]) );
  DFF \sreg_reg[1588]  ( .D(c[1589]), .CLK(clk), .RST(rst), .Q(sreg[1588]) );
  DFF \sreg_reg[1587]  ( .D(c[1588]), .CLK(clk), .RST(rst), .Q(sreg[1587]) );
  DFF \sreg_reg[1586]  ( .D(c[1587]), .CLK(clk), .RST(rst), .Q(sreg[1586]) );
  DFF \sreg_reg[1585]  ( .D(c[1586]), .CLK(clk), .RST(rst), .Q(sreg[1585]) );
  DFF \sreg_reg[1584]  ( .D(c[1585]), .CLK(clk), .RST(rst), .Q(sreg[1584]) );
  DFF \sreg_reg[1583]  ( .D(c[1584]), .CLK(clk), .RST(rst), .Q(sreg[1583]) );
  DFF \sreg_reg[1582]  ( .D(c[1583]), .CLK(clk), .RST(rst), .Q(sreg[1582]) );
  DFF \sreg_reg[1581]  ( .D(c[1582]), .CLK(clk), .RST(rst), .Q(sreg[1581]) );
  DFF \sreg_reg[1580]  ( .D(c[1581]), .CLK(clk), .RST(rst), .Q(sreg[1580]) );
  DFF \sreg_reg[1579]  ( .D(c[1580]), .CLK(clk), .RST(rst), .Q(sreg[1579]) );
  DFF \sreg_reg[1578]  ( .D(c[1579]), .CLK(clk), .RST(rst), .Q(sreg[1578]) );
  DFF \sreg_reg[1577]  ( .D(c[1578]), .CLK(clk), .RST(rst), .Q(sreg[1577]) );
  DFF \sreg_reg[1576]  ( .D(c[1577]), .CLK(clk), .RST(rst), .Q(sreg[1576]) );
  DFF \sreg_reg[1575]  ( .D(c[1576]), .CLK(clk), .RST(rst), .Q(sreg[1575]) );
  DFF \sreg_reg[1574]  ( .D(c[1575]), .CLK(clk), .RST(rst), .Q(sreg[1574]) );
  DFF \sreg_reg[1573]  ( .D(c[1574]), .CLK(clk), .RST(rst), .Q(sreg[1573]) );
  DFF \sreg_reg[1572]  ( .D(c[1573]), .CLK(clk), .RST(rst), .Q(sreg[1572]) );
  DFF \sreg_reg[1571]  ( .D(c[1572]), .CLK(clk), .RST(rst), .Q(sreg[1571]) );
  DFF \sreg_reg[1570]  ( .D(c[1571]), .CLK(clk), .RST(rst), .Q(sreg[1570]) );
  DFF \sreg_reg[1569]  ( .D(c[1570]), .CLK(clk), .RST(rst), .Q(sreg[1569]) );
  DFF \sreg_reg[1568]  ( .D(c[1569]), .CLK(clk), .RST(rst), .Q(sreg[1568]) );
  DFF \sreg_reg[1567]  ( .D(c[1568]), .CLK(clk), .RST(rst), .Q(sreg[1567]) );
  DFF \sreg_reg[1566]  ( .D(c[1567]), .CLK(clk), .RST(rst), .Q(sreg[1566]) );
  DFF \sreg_reg[1565]  ( .D(c[1566]), .CLK(clk), .RST(rst), .Q(sreg[1565]) );
  DFF \sreg_reg[1564]  ( .D(c[1565]), .CLK(clk), .RST(rst), .Q(sreg[1564]) );
  DFF \sreg_reg[1563]  ( .D(c[1564]), .CLK(clk), .RST(rst), .Q(sreg[1563]) );
  DFF \sreg_reg[1562]  ( .D(c[1563]), .CLK(clk), .RST(rst), .Q(sreg[1562]) );
  DFF \sreg_reg[1561]  ( .D(c[1562]), .CLK(clk), .RST(rst), .Q(sreg[1561]) );
  DFF \sreg_reg[1560]  ( .D(c[1561]), .CLK(clk), .RST(rst), .Q(sreg[1560]) );
  DFF \sreg_reg[1559]  ( .D(c[1560]), .CLK(clk), .RST(rst), .Q(sreg[1559]) );
  DFF \sreg_reg[1558]  ( .D(c[1559]), .CLK(clk), .RST(rst), .Q(sreg[1558]) );
  DFF \sreg_reg[1557]  ( .D(c[1558]), .CLK(clk), .RST(rst), .Q(sreg[1557]) );
  DFF \sreg_reg[1556]  ( .D(c[1557]), .CLK(clk), .RST(rst), .Q(sreg[1556]) );
  DFF \sreg_reg[1555]  ( .D(c[1556]), .CLK(clk), .RST(rst), .Q(sreg[1555]) );
  DFF \sreg_reg[1554]  ( .D(c[1555]), .CLK(clk), .RST(rst), .Q(sreg[1554]) );
  DFF \sreg_reg[1553]  ( .D(c[1554]), .CLK(clk), .RST(rst), .Q(sreg[1553]) );
  DFF \sreg_reg[1552]  ( .D(c[1553]), .CLK(clk), .RST(rst), .Q(sreg[1552]) );
  DFF \sreg_reg[1551]  ( .D(c[1552]), .CLK(clk), .RST(rst), .Q(sreg[1551]) );
  DFF \sreg_reg[1550]  ( .D(c[1551]), .CLK(clk), .RST(rst), .Q(sreg[1550]) );
  DFF \sreg_reg[1549]  ( .D(c[1550]), .CLK(clk), .RST(rst), .Q(sreg[1549]) );
  DFF \sreg_reg[1548]  ( .D(c[1549]), .CLK(clk), .RST(rst), .Q(sreg[1548]) );
  DFF \sreg_reg[1547]  ( .D(c[1548]), .CLK(clk), .RST(rst), .Q(sreg[1547]) );
  DFF \sreg_reg[1546]  ( .D(c[1547]), .CLK(clk), .RST(rst), .Q(sreg[1546]) );
  DFF \sreg_reg[1545]  ( .D(c[1546]), .CLK(clk), .RST(rst), .Q(sreg[1545]) );
  DFF \sreg_reg[1544]  ( .D(c[1545]), .CLK(clk), .RST(rst), .Q(sreg[1544]) );
  DFF \sreg_reg[1543]  ( .D(c[1544]), .CLK(clk), .RST(rst), .Q(sreg[1543]) );
  DFF \sreg_reg[1542]  ( .D(c[1543]), .CLK(clk), .RST(rst), .Q(sreg[1542]) );
  DFF \sreg_reg[1541]  ( .D(c[1542]), .CLK(clk), .RST(rst), .Q(sreg[1541]) );
  DFF \sreg_reg[1540]  ( .D(c[1541]), .CLK(clk), .RST(rst), .Q(sreg[1540]) );
  DFF \sreg_reg[1539]  ( .D(c[1540]), .CLK(clk), .RST(rst), .Q(sreg[1539]) );
  DFF \sreg_reg[1538]  ( .D(c[1539]), .CLK(clk), .RST(rst), .Q(sreg[1538]) );
  DFF \sreg_reg[1537]  ( .D(c[1538]), .CLK(clk), .RST(rst), .Q(sreg[1537]) );
  DFF \sreg_reg[1536]  ( .D(c[1537]), .CLK(clk), .RST(rst), .Q(sreg[1536]) );
  DFF \sreg_reg[1535]  ( .D(c[1536]), .CLK(clk), .RST(rst), .Q(sreg[1535]) );
  DFF \sreg_reg[1534]  ( .D(c[1535]), .CLK(clk), .RST(rst), .Q(sreg[1534]) );
  DFF \sreg_reg[1533]  ( .D(c[1534]), .CLK(clk), .RST(rst), .Q(sreg[1533]) );
  DFF \sreg_reg[1532]  ( .D(c[1533]), .CLK(clk), .RST(rst), .Q(sreg[1532]) );
  DFF \sreg_reg[1531]  ( .D(c[1532]), .CLK(clk), .RST(rst), .Q(sreg[1531]) );
  DFF \sreg_reg[1530]  ( .D(c[1531]), .CLK(clk), .RST(rst), .Q(sreg[1530]) );
  DFF \sreg_reg[1529]  ( .D(c[1530]), .CLK(clk), .RST(rst), .Q(sreg[1529]) );
  DFF \sreg_reg[1528]  ( .D(c[1529]), .CLK(clk), .RST(rst), .Q(sreg[1528]) );
  DFF \sreg_reg[1527]  ( .D(c[1528]), .CLK(clk), .RST(rst), .Q(sreg[1527]) );
  DFF \sreg_reg[1526]  ( .D(c[1527]), .CLK(clk), .RST(rst), .Q(sreg[1526]) );
  DFF \sreg_reg[1525]  ( .D(c[1526]), .CLK(clk), .RST(rst), .Q(sreg[1525]) );
  DFF \sreg_reg[1524]  ( .D(c[1525]), .CLK(clk), .RST(rst), .Q(sreg[1524]) );
  DFF \sreg_reg[1523]  ( .D(c[1524]), .CLK(clk), .RST(rst), .Q(sreg[1523]) );
  DFF \sreg_reg[1522]  ( .D(c[1523]), .CLK(clk), .RST(rst), .Q(sreg[1522]) );
  DFF \sreg_reg[1521]  ( .D(c[1522]), .CLK(clk), .RST(rst), .Q(sreg[1521]) );
  DFF \sreg_reg[1520]  ( .D(c[1521]), .CLK(clk), .RST(rst), .Q(sreg[1520]) );
  DFF \sreg_reg[1519]  ( .D(c[1520]), .CLK(clk), .RST(rst), .Q(sreg[1519]) );
  DFF \sreg_reg[1518]  ( .D(c[1519]), .CLK(clk), .RST(rst), .Q(sreg[1518]) );
  DFF \sreg_reg[1517]  ( .D(c[1518]), .CLK(clk), .RST(rst), .Q(sreg[1517]) );
  DFF \sreg_reg[1516]  ( .D(c[1517]), .CLK(clk), .RST(rst), .Q(sreg[1516]) );
  DFF \sreg_reg[1515]  ( .D(c[1516]), .CLK(clk), .RST(rst), .Q(sreg[1515]) );
  DFF \sreg_reg[1514]  ( .D(c[1515]), .CLK(clk), .RST(rst), .Q(sreg[1514]) );
  DFF \sreg_reg[1513]  ( .D(c[1514]), .CLK(clk), .RST(rst), .Q(sreg[1513]) );
  DFF \sreg_reg[1512]  ( .D(c[1513]), .CLK(clk), .RST(rst), .Q(sreg[1512]) );
  DFF \sreg_reg[1511]  ( .D(c[1512]), .CLK(clk), .RST(rst), .Q(sreg[1511]) );
  DFF \sreg_reg[1510]  ( .D(c[1511]), .CLK(clk), .RST(rst), .Q(sreg[1510]) );
  DFF \sreg_reg[1509]  ( .D(c[1510]), .CLK(clk), .RST(rst), .Q(sreg[1509]) );
  DFF \sreg_reg[1508]  ( .D(c[1509]), .CLK(clk), .RST(rst), .Q(sreg[1508]) );
  DFF \sreg_reg[1507]  ( .D(c[1508]), .CLK(clk), .RST(rst), .Q(sreg[1507]) );
  DFF \sreg_reg[1506]  ( .D(c[1507]), .CLK(clk), .RST(rst), .Q(sreg[1506]) );
  DFF \sreg_reg[1505]  ( .D(c[1506]), .CLK(clk), .RST(rst), .Q(sreg[1505]) );
  DFF \sreg_reg[1504]  ( .D(c[1505]), .CLK(clk), .RST(rst), .Q(sreg[1504]) );
  DFF \sreg_reg[1503]  ( .D(c[1504]), .CLK(clk), .RST(rst), .Q(sreg[1503]) );
  DFF \sreg_reg[1502]  ( .D(c[1503]), .CLK(clk), .RST(rst), .Q(sreg[1502]) );
  DFF \sreg_reg[1501]  ( .D(c[1502]), .CLK(clk), .RST(rst), .Q(sreg[1501]) );
  DFF \sreg_reg[1500]  ( .D(c[1501]), .CLK(clk), .RST(rst), .Q(sreg[1500]) );
  DFF \sreg_reg[1499]  ( .D(c[1500]), .CLK(clk), .RST(rst), .Q(sreg[1499]) );
  DFF \sreg_reg[1498]  ( .D(c[1499]), .CLK(clk), .RST(rst), .Q(sreg[1498]) );
  DFF \sreg_reg[1497]  ( .D(c[1498]), .CLK(clk), .RST(rst), .Q(sreg[1497]) );
  DFF \sreg_reg[1496]  ( .D(c[1497]), .CLK(clk), .RST(rst), .Q(sreg[1496]) );
  DFF \sreg_reg[1495]  ( .D(c[1496]), .CLK(clk), .RST(rst), .Q(sreg[1495]) );
  DFF \sreg_reg[1494]  ( .D(c[1495]), .CLK(clk), .RST(rst), .Q(sreg[1494]) );
  DFF \sreg_reg[1493]  ( .D(c[1494]), .CLK(clk), .RST(rst), .Q(sreg[1493]) );
  DFF \sreg_reg[1492]  ( .D(c[1493]), .CLK(clk), .RST(rst), .Q(sreg[1492]) );
  DFF \sreg_reg[1491]  ( .D(c[1492]), .CLK(clk), .RST(rst), .Q(sreg[1491]) );
  DFF \sreg_reg[1490]  ( .D(c[1491]), .CLK(clk), .RST(rst), .Q(sreg[1490]) );
  DFF \sreg_reg[1489]  ( .D(c[1490]), .CLK(clk), .RST(rst), .Q(sreg[1489]) );
  DFF \sreg_reg[1488]  ( .D(c[1489]), .CLK(clk), .RST(rst), .Q(sreg[1488]) );
  DFF \sreg_reg[1487]  ( .D(c[1488]), .CLK(clk), .RST(rst), .Q(sreg[1487]) );
  DFF \sreg_reg[1486]  ( .D(c[1487]), .CLK(clk), .RST(rst), .Q(sreg[1486]) );
  DFF \sreg_reg[1485]  ( .D(c[1486]), .CLK(clk), .RST(rst), .Q(sreg[1485]) );
  DFF \sreg_reg[1484]  ( .D(c[1485]), .CLK(clk), .RST(rst), .Q(sreg[1484]) );
  DFF \sreg_reg[1483]  ( .D(c[1484]), .CLK(clk), .RST(rst), .Q(sreg[1483]) );
  DFF \sreg_reg[1482]  ( .D(c[1483]), .CLK(clk), .RST(rst), .Q(sreg[1482]) );
  DFF \sreg_reg[1481]  ( .D(c[1482]), .CLK(clk), .RST(rst), .Q(sreg[1481]) );
  DFF \sreg_reg[1480]  ( .D(c[1481]), .CLK(clk), .RST(rst), .Q(sreg[1480]) );
  DFF \sreg_reg[1479]  ( .D(c[1480]), .CLK(clk), .RST(rst), .Q(sreg[1479]) );
  DFF \sreg_reg[1478]  ( .D(c[1479]), .CLK(clk), .RST(rst), .Q(sreg[1478]) );
  DFF \sreg_reg[1477]  ( .D(c[1478]), .CLK(clk), .RST(rst), .Q(sreg[1477]) );
  DFF \sreg_reg[1476]  ( .D(c[1477]), .CLK(clk), .RST(rst), .Q(sreg[1476]) );
  DFF \sreg_reg[1475]  ( .D(c[1476]), .CLK(clk), .RST(rst), .Q(sreg[1475]) );
  DFF \sreg_reg[1474]  ( .D(c[1475]), .CLK(clk), .RST(rst), .Q(sreg[1474]) );
  DFF \sreg_reg[1473]  ( .D(c[1474]), .CLK(clk), .RST(rst), .Q(sreg[1473]) );
  DFF \sreg_reg[1472]  ( .D(c[1473]), .CLK(clk), .RST(rst), .Q(sreg[1472]) );
  DFF \sreg_reg[1471]  ( .D(c[1472]), .CLK(clk), .RST(rst), .Q(sreg[1471]) );
  DFF \sreg_reg[1470]  ( .D(c[1471]), .CLK(clk), .RST(rst), .Q(sreg[1470]) );
  DFF \sreg_reg[1469]  ( .D(c[1470]), .CLK(clk), .RST(rst), .Q(sreg[1469]) );
  DFF \sreg_reg[1468]  ( .D(c[1469]), .CLK(clk), .RST(rst), .Q(sreg[1468]) );
  DFF \sreg_reg[1467]  ( .D(c[1468]), .CLK(clk), .RST(rst), .Q(sreg[1467]) );
  DFF \sreg_reg[1466]  ( .D(c[1467]), .CLK(clk), .RST(rst), .Q(sreg[1466]) );
  DFF \sreg_reg[1465]  ( .D(c[1466]), .CLK(clk), .RST(rst), .Q(sreg[1465]) );
  DFF \sreg_reg[1464]  ( .D(c[1465]), .CLK(clk), .RST(rst), .Q(sreg[1464]) );
  DFF \sreg_reg[1463]  ( .D(c[1464]), .CLK(clk), .RST(rst), .Q(sreg[1463]) );
  DFF \sreg_reg[1462]  ( .D(c[1463]), .CLK(clk), .RST(rst), .Q(sreg[1462]) );
  DFF \sreg_reg[1461]  ( .D(c[1462]), .CLK(clk), .RST(rst), .Q(sreg[1461]) );
  DFF \sreg_reg[1460]  ( .D(c[1461]), .CLK(clk), .RST(rst), .Q(sreg[1460]) );
  DFF \sreg_reg[1459]  ( .D(c[1460]), .CLK(clk), .RST(rst), .Q(sreg[1459]) );
  DFF \sreg_reg[1458]  ( .D(c[1459]), .CLK(clk), .RST(rst), .Q(sreg[1458]) );
  DFF \sreg_reg[1457]  ( .D(c[1458]), .CLK(clk), .RST(rst), .Q(sreg[1457]) );
  DFF \sreg_reg[1456]  ( .D(c[1457]), .CLK(clk), .RST(rst), .Q(sreg[1456]) );
  DFF \sreg_reg[1455]  ( .D(c[1456]), .CLK(clk), .RST(rst), .Q(sreg[1455]) );
  DFF \sreg_reg[1454]  ( .D(c[1455]), .CLK(clk), .RST(rst), .Q(sreg[1454]) );
  DFF \sreg_reg[1453]  ( .D(c[1454]), .CLK(clk), .RST(rst), .Q(sreg[1453]) );
  DFF \sreg_reg[1452]  ( .D(c[1453]), .CLK(clk), .RST(rst), .Q(sreg[1452]) );
  DFF \sreg_reg[1451]  ( .D(c[1452]), .CLK(clk), .RST(rst), .Q(sreg[1451]) );
  DFF \sreg_reg[1450]  ( .D(c[1451]), .CLK(clk), .RST(rst), .Q(sreg[1450]) );
  DFF \sreg_reg[1449]  ( .D(c[1450]), .CLK(clk), .RST(rst), .Q(sreg[1449]) );
  DFF \sreg_reg[1448]  ( .D(c[1449]), .CLK(clk), .RST(rst), .Q(sreg[1448]) );
  DFF \sreg_reg[1447]  ( .D(c[1448]), .CLK(clk), .RST(rst), .Q(sreg[1447]) );
  DFF \sreg_reg[1446]  ( .D(c[1447]), .CLK(clk), .RST(rst), .Q(sreg[1446]) );
  DFF \sreg_reg[1445]  ( .D(c[1446]), .CLK(clk), .RST(rst), .Q(sreg[1445]) );
  DFF \sreg_reg[1444]  ( .D(c[1445]), .CLK(clk), .RST(rst), .Q(sreg[1444]) );
  DFF \sreg_reg[1443]  ( .D(c[1444]), .CLK(clk), .RST(rst), .Q(sreg[1443]) );
  DFF \sreg_reg[1442]  ( .D(c[1443]), .CLK(clk), .RST(rst), .Q(sreg[1442]) );
  DFF \sreg_reg[1441]  ( .D(c[1442]), .CLK(clk), .RST(rst), .Q(sreg[1441]) );
  DFF \sreg_reg[1440]  ( .D(c[1441]), .CLK(clk), .RST(rst), .Q(sreg[1440]) );
  DFF \sreg_reg[1439]  ( .D(c[1440]), .CLK(clk), .RST(rst), .Q(sreg[1439]) );
  DFF \sreg_reg[1438]  ( .D(c[1439]), .CLK(clk), .RST(rst), .Q(sreg[1438]) );
  DFF \sreg_reg[1437]  ( .D(c[1438]), .CLK(clk), .RST(rst), .Q(sreg[1437]) );
  DFF \sreg_reg[1436]  ( .D(c[1437]), .CLK(clk), .RST(rst), .Q(sreg[1436]) );
  DFF \sreg_reg[1435]  ( .D(c[1436]), .CLK(clk), .RST(rst), .Q(sreg[1435]) );
  DFF \sreg_reg[1434]  ( .D(c[1435]), .CLK(clk), .RST(rst), .Q(sreg[1434]) );
  DFF \sreg_reg[1433]  ( .D(c[1434]), .CLK(clk), .RST(rst), .Q(sreg[1433]) );
  DFF \sreg_reg[1432]  ( .D(c[1433]), .CLK(clk), .RST(rst), .Q(sreg[1432]) );
  DFF \sreg_reg[1431]  ( .D(c[1432]), .CLK(clk), .RST(rst), .Q(sreg[1431]) );
  DFF \sreg_reg[1430]  ( .D(c[1431]), .CLK(clk), .RST(rst), .Q(sreg[1430]) );
  DFF \sreg_reg[1429]  ( .D(c[1430]), .CLK(clk), .RST(rst), .Q(sreg[1429]) );
  DFF \sreg_reg[1428]  ( .D(c[1429]), .CLK(clk), .RST(rst), .Q(sreg[1428]) );
  DFF \sreg_reg[1427]  ( .D(c[1428]), .CLK(clk), .RST(rst), .Q(sreg[1427]) );
  DFF \sreg_reg[1426]  ( .D(c[1427]), .CLK(clk), .RST(rst), .Q(sreg[1426]) );
  DFF \sreg_reg[1425]  ( .D(c[1426]), .CLK(clk), .RST(rst), .Q(sreg[1425]) );
  DFF \sreg_reg[1424]  ( .D(c[1425]), .CLK(clk), .RST(rst), .Q(sreg[1424]) );
  DFF \sreg_reg[1423]  ( .D(c[1424]), .CLK(clk), .RST(rst), .Q(sreg[1423]) );
  DFF \sreg_reg[1422]  ( .D(c[1423]), .CLK(clk), .RST(rst), .Q(sreg[1422]) );
  DFF \sreg_reg[1421]  ( .D(c[1422]), .CLK(clk), .RST(rst), .Q(sreg[1421]) );
  DFF \sreg_reg[1420]  ( .D(c[1421]), .CLK(clk), .RST(rst), .Q(sreg[1420]) );
  DFF \sreg_reg[1419]  ( .D(c[1420]), .CLK(clk), .RST(rst), .Q(sreg[1419]) );
  DFF \sreg_reg[1418]  ( .D(c[1419]), .CLK(clk), .RST(rst), .Q(sreg[1418]) );
  DFF \sreg_reg[1417]  ( .D(c[1418]), .CLK(clk), .RST(rst), .Q(sreg[1417]) );
  DFF \sreg_reg[1416]  ( .D(c[1417]), .CLK(clk), .RST(rst), .Q(sreg[1416]) );
  DFF \sreg_reg[1415]  ( .D(c[1416]), .CLK(clk), .RST(rst), .Q(sreg[1415]) );
  DFF \sreg_reg[1414]  ( .D(c[1415]), .CLK(clk), .RST(rst), .Q(sreg[1414]) );
  DFF \sreg_reg[1413]  ( .D(c[1414]), .CLK(clk), .RST(rst), .Q(sreg[1413]) );
  DFF \sreg_reg[1412]  ( .D(c[1413]), .CLK(clk), .RST(rst), .Q(sreg[1412]) );
  DFF \sreg_reg[1411]  ( .D(c[1412]), .CLK(clk), .RST(rst), .Q(sreg[1411]) );
  DFF \sreg_reg[1410]  ( .D(c[1411]), .CLK(clk), .RST(rst), .Q(sreg[1410]) );
  DFF \sreg_reg[1409]  ( .D(c[1410]), .CLK(clk), .RST(rst), .Q(sreg[1409]) );
  DFF \sreg_reg[1408]  ( .D(c[1409]), .CLK(clk), .RST(rst), .Q(sreg[1408]) );
  DFF \sreg_reg[1407]  ( .D(c[1408]), .CLK(clk), .RST(rst), .Q(sreg[1407]) );
  DFF \sreg_reg[1406]  ( .D(c[1407]), .CLK(clk), .RST(rst), .Q(sreg[1406]) );
  DFF \sreg_reg[1405]  ( .D(c[1406]), .CLK(clk), .RST(rst), .Q(sreg[1405]) );
  DFF \sreg_reg[1404]  ( .D(c[1405]), .CLK(clk), .RST(rst), .Q(sreg[1404]) );
  DFF \sreg_reg[1403]  ( .D(c[1404]), .CLK(clk), .RST(rst), .Q(sreg[1403]) );
  DFF \sreg_reg[1402]  ( .D(c[1403]), .CLK(clk), .RST(rst), .Q(sreg[1402]) );
  DFF \sreg_reg[1401]  ( .D(c[1402]), .CLK(clk), .RST(rst), .Q(sreg[1401]) );
  DFF \sreg_reg[1400]  ( .D(c[1401]), .CLK(clk), .RST(rst), .Q(sreg[1400]) );
  DFF \sreg_reg[1399]  ( .D(c[1400]), .CLK(clk), .RST(rst), .Q(sreg[1399]) );
  DFF \sreg_reg[1398]  ( .D(c[1399]), .CLK(clk), .RST(rst), .Q(sreg[1398]) );
  DFF \sreg_reg[1397]  ( .D(c[1398]), .CLK(clk), .RST(rst), .Q(sreg[1397]) );
  DFF \sreg_reg[1396]  ( .D(c[1397]), .CLK(clk), .RST(rst), .Q(sreg[1396]) );
  DFF \sreg_reg[1395]  ( .D(c[1396]), .CLK(clk), .RST(rst), .Q(sreg[1395]) );
  DFF \sreg_reg[1394]  ( .D(c[1395]), .CLK(clk), .RST(rst), .Q(sreg[1394]) );
  DFF \sreg_reg[1393]  ( .D(c[1394]), .CLK(clk), .RST(rst), .Q(sreg[1393]) );
  DFF \sreg_reg[1392]  ( .D(c[1393]), .CLK(clk), .RST(rst), .Q(sreg[1392]) );
  DFF \sreg_reg[1391]  ( .D(c[1392]), .CLK(clk), .RST(rst), .Q(sreg[1391]) );
  DFF \sreg_reg[1390]  ( .D(c[1391]), .CLK(clk), .RST(rst), .Q(sreg[1390]) );
  DFF \sreg_reg[1389]  ( .D(c[1390]), .CLK(clk), .RST(rst), .Q(sreg[1389]) );
  DFF \sreg_reg[1388]  ( .D(c[1389]), .CLK(clk), .RST(rst), .Q(sreg[1388]) );
  DFF \sreg_reg[1387]  ( .D(c[1388]), .CLK(clk), .RST(rst), .Q(sreg[1387]) );
  DFF \sreg_reg[1386]  ( .D(c[1387]), .CLK(clk), .RST(rst), .Q(sreg[1386]) );
  DFF \sreg_reg[1385]  ( .D(c[1386]), .CLK(clk), .RST(rst), .Q(sreg[1385]) );
  DFF \sreg_reg[1384]  ( .D(c[1385]), .CLK(clk), .RST(rst), .Q(sreg[1384]) );
  DFF \sreg_reg[1383]  ( .D(c[1384]), .CLK(clk), .RST(rst), .Q(sreg[1383]) );
  DFF \sreg_reg[1382]  ( .D(c[1383]), .CLK(clk), .RST(rst), .Q(sreg[1382]) );
  DFF \sreg_reg[1381]  ( .D(c[1382]), .CLK(clk), .RST(rst), .Q(sreg[1381]) );
  DFF \sreg_reg[1380]  ( .D(c[1381]), .CLK(clk), .RST(rst), .Q(sreg[1380]) );
  DFF \sreg_reg[1379]  ( .D(c[1380]), .CLK(clk), .RST(rst), .Q(sreg[1379]) );
  DFF \sreg_reg[1378]  ( .D(c[1379]), .CLK(clk), .RST(rst), .Q(sreg[1378]) );
  DFF \sreg_reg[1377]  ( .D(c[1378]), .CLK(clk), .RST(rst), .Q(sreg[1377]) );
  DFF \sreg_reg[1376]  ( .D(c[1377]), .CLK(clk), .RST(rst), .Q(sreg[1376]) );
  DFF \sreg_reg[1375]  ( .D(c[1376]), .CLK(clk), .RST(rst), .Q(sreg[1375]) );
  DFF \sreg_reg[1374]  ( .D(c[1375]), .CLK(clk), .RST(rst), .Q(sreg[1374]) );
  DFF \sreg_reg[1373]  ( .D(c[1374]), .CLK(clk), .RST(rst), .Q(sreg[1373]) );
  DFF \sreg_reg[1372]  ( .D(c[1373]), .CLK(clk), .RST(rst), .Q(sreg[1372]) );
  DFF \sreg_reg[1371]  ( .D(c[1372]), .CLK(clk), .RST(rst), .Q(sreg[1371]) );
  DFF \sreg_reg[1370]  ( .D(c[1371]), .CLK(clk), .RST(rst), .Q(sreg[1370]) );
  DFF \sreg_reg[1369]  ( .D(c[1370]), .CLK(clk), .RST(rst), .Q(sreg[1369]) );
  DFF \sreg_reg[1368]  ( .D(c[1369]), .CLK(clk), .RST(rst), .Q(sreg[1368]) );
  DFF \sreg_reg[1367]  ( .D(c[1368]), .CLK(clk), .RST(rst), .Q(sreg[1367]) );
  DFF \sreg_reg[1366]  ( .D(c[1367]), .CLK(clk), .RST(rst), .Q(sreg[1366]) );
  DFF \sreg_reg[1365]  ( .D(c[1366]), .CLK(clk), .RST(rst), .Q(sreg[1365]) );
  DFF \sreg_reg[1364]  ( .D(c[1365]), .CLK(clk), .RST(rst), .Q(sreg[1364]) );
  DFF \sreg_reg[1363]  ( .D(c[1364]), .CLK(clk), .RST(rst), .Q(sreg[1363]) );
  DFF \sreg_reg[1362]  ( .D(c[1363]), .CLK(clk), .RST(rst), .Q(sreg[1362]) );
  DFF \sreg_reg[1361]  ( .D(c[1362]), .CLK(clk), .RST(rst), .Q(sreg[1361]) );
  DFF \sreg_reg[1360]  ( .D(c[1361]), .CLK(clk), .RST(rst), .Q(sreg[1360]) );
  DFF \sreg_reg[1359]  ( .D(c[1360]), .CLK(clk), .RST(rst), .Q(sreg[1359]) );
  DFF \sreg_reg[1358]  ( .D(c[1359]), .CLK(clk), .RST(rst), .Q(sreg[1358]) );
  DFF \sreg_reg[1357]  ( .D(c[1358]), .CLK(clk), .RST(rst), .Q(sreg[1357]) );
  DFF \sreg_reg[1356]  ( .D(c[1357]), .CLK(clk), .RST(rst), .Q(sreg[1356]) );
  DFF \sreg_reg[1355]  ( .D(c[1356]), .CLK(clk), .RST(rst), .Q(sreg[1355]) );
  DFF \sreg_reg[1354]  ( .D(c[1355]), .CLK(clk), .RST(rst), .Q(sreg[1354]) );
  DFF \sreg_reg[1353]  ( .D(c[1354]), .CLK(clk), .RST(rst), .Q(sreg[1353]) );
  DFF \sreg_reg[1352]  ( .D(c[1353]), .CLK(clk), .RST(rst), .Q(sreg[1352]) );
  DFF \sreg_reg[1351]  ( .D(c[1352]), .CLK(clk), .RST(rst), .Q(sreg[1351]) );
  DFF \sreg_reg[1350]  ( .D(c[1351]), .CLK(clk), .RST(rst), .Q(sreg[1350]) );
  DFF \sreg_reg[1349]  ( .D(c[1350]), .CLK(clk), .RST(rst), .Q(sreg[1349]) );
  DFF \sreg_reg[1348]  ( .D(c[1349]), .CLK(clk), .RST(rst), .Q(sreg[1348]) );
  DFF \sreg_reg[1347]  ( .D(c[1348]), .CLK(clk), .RST(rst), .Q(sreg[1347]) );
  DFF \sreg_reg[1346]  ( .D(c[1347]), .CLK(clk), .RST(rst), .Q(sreg[1346]) );
  DFF \sreg_reg[1345]  ( .D(c[1346]), .CLK(clk), .RST(rst), .Q(sreg[1345]) );
  DFF \sreg_reg[1344]  ( .D(c[1345]), .CLK(clk), .RST(rst), .Q(sreg[1344]) );
  DFF \sreg_reg[1343]  ( .D(c[1344]), .CLK(clk), .RST(rst), .Q(sreg[1343]) );
  DFF \sreg_reg[1342]  ( .D(c[1343]), .CLK(clk), .RST(rst), .Q(sreg[1342]) );
  DFF \sreg_reg[1341]  ( .D(c[1342]), .CLK(clk), .RST(rst), .Q(sreg[1341]) );
  DFF \sreg_reg[1340]  ( .D(c[1341]), .CLK(clk), .RST(rst), .Q(sreg[1340]) );
  DFF \sreg_reg[1339]  ( .D(c[1340]), .CLK(clk), .RST(rst), .Q(sreg[1339]) );
  DFF \sreg_reg[1338]  ( .D(c[1339]), .CLK(clk), .RST(rst), .Q(sreg[1338]) );
  DFF \sreg_reg[1337]  ( .D(c[1338]), .CLK(clk), .RST(rst), .Q(sreg[1337]) );
  DFF \sreg_reg[1336]  ( .D(c[1337]), .CLK(clk), .RST(rst), .Q(sreg[1336]) );
  DFF \sreg_reg[1335]  ( .D(c[1336]), .CLK(clk), .RST(rst), .Q(sreg[1335]) );
  DFF \sreg_reg[1334]  ( .D(c[1335]), .CLK(clk), .RST(rst), .Q(sreg[1334]) );
  DFF \sreg_reg[1333]  ( .D(c[1334]), .CLK(clk), .RST(rst), .Q(sreg[1333]) );
  DFF \sreg_reg[1332]  ( .D(c[1333]), .CLK(clk), .RST(rst), .Q(sreg[1332]) );
  DFF \sreg_reg[1331]  ( .D(c[1332]), .CLK(clk), .RST(rst), .Q(sreg[1331]) );
  DFF \sreg_reg[1330]  ( .D(c[1331]), .CLK(clk), .RST(rst), .Q(sreg[1330]) );
  DFF \sreg_reg[1329]  ( .D(c[1330]), .CLK(clk), .RST(rst), .Q(sreg[1329]) );
  DFF \sreg_reg[1328]  ( .D(c[1329]), .CLK(clk), .RST(rst), .Q(sreg[1328]) );
  DFF \sreg_reg[1327]  ( .D(c[1328]), .CLK(clk), .RST(rst), .Q(sreg[1327]) );
  DFF \sreg_reg[1326]  ( .D(c[1327]), .CLK(clk), .RST(rst), .Q(sreg[1326]) );
  DFF \sreg_reg[1325]  ( .D(c[1326]), .CLK(clk), .RST(rst), .Q(sreg[1325]) );
  DFF \sreg_reg[1324]  ( .D(c[1325]), .CLK(clk), .RST(rst), .Q(sreg[1324]) );
  DFF \sreg_reg[1323]  ( .D(c[1324]), .CLK(clk), .RST(rst), .Q(sreg[1323]) );
  DFF \sreg_reg[1322]  ( .D(c[1323]), .CLK(clk), .RST(rst), .Q(sreg[1322]) );
  DFF \sreg_reg[1321]  ( .D(c[1322]), .CLK(clk), .RST(rst), .Q(sreg[1321]) );
  DFF \sreg_reg[1320]  ( .D(c[1321]), .CLK(clk), .RST(rst), .Q(sreg[1320]) );
  DFF \sreg_reg[1319]  ( .D(c[1320]), .CLK(clk), .RST(rst), .Q(sreg[1319]) );
  DFF \sreg_reg[1318]  ( .D(c[1319]), .CLK(clk), .RST(rst), .Q(sreg[1318]) );
  DFF \sreg_reg[1317]  ( .D(c[1318]), .CLK(clk), .RST(rst), .Q(sreg[1317]) );
  DFF \sreg_reg[1316]  ( .D(c[1317]), .CLK(clk), .RST(rst), .Q(sreg[1316]) );
  DFF \sreg_reg[1315]  ( .D(c[1316]), .CLK(clk), .RST(rst), .Q(sreg[1315]) );
  DFF \sreg_reg[1314]  ( .D(c[1315]), .CLK(clk), .RST(rst), .Q(sreg[1314]) );
  DFF \sreg_reg[1313]  ( .D(c[1314]), .CLK(clk), .RST(rst), .Q(sreg[1313]) );
  DFF \sreg_reg[1312]  ( .D(c[1313]), .CLK(clk), .RST(rst), .Q(sreg[1312]) );
  DFF \sreg_reg[1311]  ( .D(c[1312]), .CLK(clk), .RST(rst), .Q(sreg[1311]) );
  DFF \sreg_reg[1310]  ( .D(c[1311]), .CLK(clk), .RST(rst), .Q(sreg[1310]) );
  DFF \sreg_reg[1309]  ( .D(c[1310]), .CLK(clk), .RST(rst), .Q(sreg[1309]) );
  DFF \sreg_reg[1308]  ( .D(c[1309]), .CLK(clk), .RST(rst), .Q(sreg[1308]) );
  DFF \sreg_reg[1307]  ( .D(c[1308]), .CLK(clk), .RST(rst), .Q(sreg[1307]) );
  DFF \sreg_reg[1306]  ( .D(c[1307]), .CLK(clk), .RST(rst), .Q(sreg[1306]) );
  DFF \sreg_reg[1305]  ( .D(c[1306]), .CLK(clk), .RST(rst), .Q(sreg[1305]) );
  DFF \sreg_reg[1304]  ( .D(c[1305]), .CLK(clk), .RST(rst), .Q(sreg[1304]) );
  DFF \sreg_reg[1303]  ( .D(c[1304]), .CLK(clk), .RST(rst), .Q(sreg[1303]) );
  DFF \sreg_reg[1302]  ( .D(c[1303]), .CLK(clk), .RST(rst), .Q(sreg[1302]) );
  DFF \sreg_reg[1301]  ( .D(c[1302]), .CLK(clk), .RST(rst), .Q(sreg[1301]) );
  DFF \sreg_reg[1300]  ( .D(c[1301]), .CLK(clk), .RST(rst), .Q(sreg[1300]) );
  DFF \sreg_reg[1299]  ( .D(c[1300]), .CLK(clk), .RST(rst), .Q(sreg[1299]) );
  DFF \sreg_reg[1298]  ( .D(c[1299]), .CLK(clk), .RST(rst), .Q(sreg[1298]) );
  DFF \sreg_reg[1297]  ( .D(c[1298]), .CLK(clk), .RST(rst), .Q(sreg[1297]) );
  DFF \sreg_reg[1296]  ( .D(c[1297]), .CLK(clk), .RST(rst), .Q(sreg[1296]) );
  DFF \sreg_reg[1295]  ( .D(c[1296]), .CLK(clk), .RST(rst), .Q(sreg[1295]) );
  DFF \sreg_reg[1294]  ( .D(c[1295]), .CLK(clk), .RST(rst), .Q(sreg[1294]) );
  DFF \sreg_reg[1293]  ( .D(c[1294]), .CLK(clk), .RST(rst), .Q(sreg[1293]) );
  DFF \sreg_reg[1292]  ( .D(c[1293]), .CLK(clk), .RST(rst), .Q(sreg[1292]) );
  DFF \sreg_reg[1291]  ( .D(c[1292]), .CLK(clk), .RST(rst), .Q(sreg[1291]) );
  DFF \sreg_reg[1290]  ( .D(c[1291]), .CLK(clk), .RST(rst), .Q(sreg[1290]) );
  DFF \sreg_reg[1289]  ( .D(c[1290]), .CLK(clk), .RST(rst), .Q(sreg[1289]) );
  DFF \sreg_reg[1288]  ( .D(c[1289]), .CLK(clk), .RST(rst), .Q(sreg[1288]) );
  DFF \sreg_reg[1287]  ( .D(c[1288]), .CLK(clk), .RST(rst), .Q(sreg[1287]) );
  DFF \sreg_reg[1286]  ( .D(c[1287]), .CLK(clk), .RST(rst), .Q(sreg[1286]) );
  DFF \sreg_reg[1285]  ( .D(c[1286]), .CLK(clk), .RST(rst), .Q(sreg[1285]) );
  DFF \sreg_reg[1284]  ( .D(c[1285]), .CLK(clk), .RST(rst), .Q(sreg[1284]) );
  DFF \sreg_reg[1283]  ( .D(c[1284]), .CLK(clk), .RST(rst), .Q(sreg[1283]) );
  DFF \sreg_reg[1282]  ( .D(c[1283]), .CLK(clk), .RST(rst), .Q(sreg[1282]) );
  DFF \sreg_reg[1281]  ( .D(c[1282]), .CLK(clk), .RST(rst), .Q(sreg[1281]) );
  DFF \sreg_reg[1280]  ( .D(c[1281]), .CLK(clk), .RST(rst), .Q(sreg[1280]) );
  DFF \sreg_reg[1279]  ( .D(c[1280]), .CLK(clk), .RST(rst), .Q(sreg[1279]) );
  DFF \sreg_reg[1278]  ( .D(c[1279]), .CLK(clk), .RST(rst), .Q(sreg[1278]) );
  DFF \sreg_reg[1277]  ( .D(c[1278]), .CLK(clk), .RST(rst), .Q(sreg[1277]) );
  DFF \sreg_reg[1276]  ( .D(c[1277]), .CLK(clk), .RST(rst), .Q(sreg[1276]) );
  DFF \sreg_reg[1275]  ( .D(c[1276]), .CLK(clk), .RST(rst), .Q(sreg[1275]) );
  DFF \sreg_reg[1274]  ( .D(c[1275]), .CLK(clk), .RST(rst), .Q(sreg[1274]) );
  DFF \sreg_reg[1273]  ( .D(c[1274]), .CLK(clk), .RST(rst), .Q(sreg[1273]) );
  DFF \sreg_reg[1272]  ( .D(c[1273]), .CLK(clk), .RST(rst), .Q(sreg[1272]) );
  DFF \sreg_reg[1271]  ( .D(c[1272]), .CLK(clk), .RST(rst), .Q(sreg[1271]) );
  DFF \sreg_reg[1270]  ( .D(c[1271]), .CLK(clk), .RST(rst), .Q(sreg[1270]) );
  DFF \sreg_reg[1269]  ( .D(c[1270]), .CLK(clk), .RST(rst), .Q(sreg[1269]) );
  DFF \sreg_reg[1268]  ( .D(c[1269]), .CLK(clk), .RST(rst), .Q(sreg[1268]) );
  DFF \sreg_reg[1267]  ( .D(c[1268]), .CLK(clk), .RST(rst), .Q(sreg[1267]) );
  DFF \sreg_reg[1266]  ( .D(c[1267]), .CLK(clk), .RST(rst), .Q(sreg[1266]) );
  DFF \sreg_reg[1265]  ( .D(c[1266]), .CLK(clk), .RST(rst), .Q(sreg[1265]) );
  DFF \sreg_reg[1264]  ( .D(c[1265]), .CLK(clk), .RST(rst), .Q(sreg[1264]) );
  DFF \sreg_reg[1263]  ( .D(c[1264]), .CLK(clk), .RST(rst), .Q(sreg[1263]) );
  DFF \sreg_reg[1262]  ( .D(c[1263]), .CLK(clk), .RST(rst), .Q(sreg[1262]) );
  DFF \sreg_reg[1261]  ( .D(c[1262]), .CLK(clk), .RST(rst), .Q(sreg[1261]) );
  DFF \sreg_reg[1260]  ( .D(c[1261]), .CLK(clk), .RST(rst), .Q(sreg[1260]) );
  DFF \sreg_reg[1259]  ( .D(c[1260]), .CLK(clk), .RST(rst), .Q(sreg[1259]) );
  DFF \sreg_reg[1258]  ( .D(c[1259]), .CLK(clk), .RST(rst), .Q(sreg[1258]) );
  DFF \sreg_reg[1257]  ( .D(c[1258]), .CLK(clk), .RST(rst), .Q(sreg[1257]) );
  DFF \sreg_reg[1256]  ( .D(c[1257]), .CLK(clk), .RST(rst), .Q(sreg[1256]) );
  DFF \sreg_reg[1255]  ( .D(c[1256]), .CLK(clk), .RST(rst), .Q(sreg[1255]) );
  DFF \sreg_reg[1254]  ( .D(c[1255]), .CLK(clk), .RST(rst), .Q(sreg[1254]) );
  DFF \sreg_reg[1253]  ( .D(c[1254]), .CLK(clk), .RST(rst), .Q(sreg[1253]) );
  DFF \sreg_reg[1252]  ( .D(c[1253]), .CLK(clk), .RST(rst), .Q(sreg[1252]) );
  DFF \sreg_reg[1251]  ( .D(c[1252]), .CLK(clk), .RST(rst), .Q(sreg[1251]) );
  DFF \sreg_reg[1250]  ( .D(c[1251]), .CLK(clk), .RST(rst), .Q(sreg[1250]) );
  DFF \sreg_reg[1249]  ( .D(c[1250]), .CLK(clk), .RST(rst), .Q(sreg[1249]) );
  DFF \sreg_reg[1248]  ( .D(c[1249]), .CLK(clk), .RST(rst), .Q(sreg[1248]) );
  DFF \sreg_reg[1247]  ( .D(c[1248]), .CLK(clk), .RST(rst), .Q(sreg[1247]) );
  DFF \sreg_reg[1246]  ( .D(c[1247]), .CLK(clk), .RST(rst), .Q(sreg[1246]) );
  DFF \sreg_reg[1245]  ( .D(c[1246]), .CLK(clk), .RST(rst), .Q(sreg[1245]) );
  DFF \sreg_reg[1244]  ( .D(c[1245]), .CLK(clk), .RST(rst), .Q(sreg[1244]) );
  DFF \sreg_reg[1243]  ( .D(c[1244]), .CLK(clk), .RST(rst), .Q(sreg[1243]) );
  DFF \sreg_reg[1242]  ( .D(c[1243]), .CLK(clk), .RST(rst), .Q(sreg[1242]) );
  DFF \sreg_reg[1241]  ( .D(c[1242]), .CLK(clk), .RST(rst), .Q(sreg[1241]) );
  DFF \sreg_reg[1240]  ( .D(c[1241]), .CLK(clk), .RST(rst), .Q(sreg[1240]) );
  DFF \sreg_reg[1239]  ( .D(c[1240]), .CLK(clk), .RST(rst), .Q(sreg[1239]) );
  DFF \sreg_reg[1238]  ( .D(c[1239]), .CLK(clk), .RST(rst), .Q(sreg[1238]) );
  DFF \sreg_reg[1237]  ( .D(c[1238]), .CLK(clk), .RST(rst), .Q(sreg[1237]) );
  DFF \sreg_reg[1236]  ( .D(c[1237]), .CLK(clk), .RST(rst), .Q(sreg[1236]) );
  DFF \sreg_reg[1235]  ( .D(c[1236]), .CLK(clk), .RST(rst), .Q(sreg[1235]) );
  DFF \sreg_reg[1234]  ( .D(c[1235]), .CLK(clk), .RST(rst), .Q(sreg[1234]) );
  DFF \sreg_reg[1233]  ( .D(c[1234]), .CLK(clk), .RST(rst), .Q(sreg[1233]) );
  DFF \sreg_reg[1232]  ( .D(c[1233]), .CLK(clk), .RST(rst), .Q(sreg[1232]) );
  DFF \sreg_reg[1231]  ( .D(c[1232]), .CLK(clk), .RST(rst), .Q(sreg[1231]) );
  DFF \sreg_reg[1230]  ( .D(c[1231]), .CLK(clk), .RST(rst), .Q(sreg[1230]) );
  DFF \sreg_reg[1229]  ( .D(c[1230]), .CLK(clk), .RST(rst), .Q(sreg[1229]) );
  DFF \sreg_reg[1228]  ( .D(c[1229]), .CLK(clk), .RST(rst), .Q(sreg[1228]) );
  DFF \sreg_reg[1227]  ( .D(c[1228]), .CLK(clk), .RST(rst), .Q(sreg[1227]) );
  DFF \sreg_reg[1226]  ( .D(c[1227]), .CLK(clk), .RST(rst), .Q(sreg[1226]) );
  DFF \sreg_reg[1225]  ( .D(c[1226]), .CLK(clk), .RST(rst), .Q(sreg[1225]) );
  DFF \sreg_reg[1224]  ( .D(c[1225]), .CLK(clk), .RST(rst), .Q(sreg[1224]) );
  DFF \sreg_reg[1223]  ( .D(c[1224]), .CLK(clk), .RST(rst), .Q(sreg[1223]) );
  DFF \sreg_reg[1222]  ( .D(c[1223]), .CLK(clk), .RST(rst), .Q(sreg[1222]) );
  DFF \sreg_reg[1221]  ( .D(c[1222]), .CLK(clk), .RST(rst), .Q(sreg[1221]) );
  DFF \sreg_reg[1220]  ( .D(c[1221]), .CLK(clk), .RST(rst), .Q(sreg[1220]) );
  DFF \sreg_reg[1219]  ( .D(c[1220]), .CLK(clk), .RST(rst), .Q(sreg[1219]) );
  DFF \sreg_reg[1218]  ( .D(c[1219]), .CLK(clk), .RST(rst), .Q(sreg[1218]) );
  DFF \sreg_reg[1217]  ( .D(c[1218]), .CLK(clk), .RST(rst), .Q(sreg[1217]) );
  DFF \sreg_reg[1216]  ( .D(c[1217]), .CLK(clk), .RST(rst), .Q(sreg[1216]) );
  DFF \sreg_reg[1215]  ( .D(c[1216]), .CLK(clk), .RST(rst), .Q(sreg[1215]) );
  DFF \sreg_reg[1214]  ( .D(c[1215]), .CLK(clk), .RST(rst), .Q(sreg[1214]) );
  DFF \sreg_reg[1213]  ( .D(c[1214]), .CLK(clk), .RST(rst), .Q(sreg[1213]) );
  DFF \sreg_reg[1212]  ( .D(c[1213]), .CLK(clk), .RST(rst), .Q(sreg[1212]) );
  DFF \sreg_reg[1211]  ( .D(c[1212]), .CLK(clk), .RST(rst), .Q(sreg[1211]) );
  DFF \sreg_reg[1210]  ( .D(c[1211]), .CLK(clk), .RST(rst), .Q(sreg[1210]) );
  DFF \sreg_reg[1209]  ( .D(c[1210]), .CLK(clk), .RST(rst), .Q(sreg[1209]) );
  DFF \sreg_reg[1208]  ( .D(c[1209]), .CLK(clk), .RST(rst), .Q(sreg[1208]) );
  DFF \sreg_reg[1207]  ( .D(c[1208]), .CLK(clk), .RST(rst), .Q(sreg[1207]) );
  DFF \sreg_reg[1206]  ( .D(c[1207]), .CLK(clk), .RST(rst), .Q(sreg[1206]) );
  DFF \sreg_reg[1205]  ( .D(c[1206]), .CLK(clk), .RST(rst), .Q(sreg[1205]) );
  DFF \sreg_reg[1204]  ( .D(c[1205]), .CLK(clk), .RST(rst), .Q(sreg[1204]) );
  DFF \sreg_reg[1203]  ( .D(c[1204]), .CLK(clk), .RST(rst), .Q(sreg[1203]) );
  DFF \sreg_reg[1202]  ( .D(c[1203]), .CLK(clk), .RST(rst), .Q(sreg[1202]) );
  DFF \sreg_reg[1201]  ( .D(c[1202]), .CLK(clk), .RST(rst), .Q(sreg[1201]) );
  DFF \sreg_reg[1200]  ( .D(c[1201]), .CLK(clk), .RST(rst), .Q(sreg[1200]) );
  DFF \sreg_reg[1199]  ( .D(c[1200]), .CLK(clk), .RST(rst), .Q(sreg[1199]) );
  DFF \sreg_reg[1198]  ( .D(c[1199]), .CLK(clk), .RST(rst), .Q(sreg[1198]) );
  DFF \sreg_reg[1197]  ( .D(c[1198]), .CLK(clk), .RST(rst), .Q(sreg[1197]) );
  DFF \sreg_reg[1196]  ( .D(c[1197]), .CLK(clk), .RST(rst), .Q(sreg[1196]) );
  DFF \sreg_reg[1195]  ( .D(c[1196]), .CLK(clk), .RST(rst), .Q(sreg[1195]) );
  DFF \sreg_reg[1194]  ( .D(c[1195]), .CLK(clk), .RST(rst), .Q(sreg[1194]) );
  DFF \sreg_reg[1193]  ( .D(c[1194]), .CLK(clk), .RST(rst), .Q(sreg[1193]) );
  DFF \sreg_reg[1192]  ( .D(c[1193]), .CLK(clk), .RST(rst), .Q(sreg[1192]) );
  DFF \sreg_reg[1191]  ( .D(c[1192]), .CLK(clk), .RST(rst), .Q(sreg[1191]) );
  DFF \sreg_reg[1190]  ( .D(c[1191]), .CLK(clk), .RST(rst), .Q(sreg[1190]) );
  DFF \sreg_reg[1189]  ( .D(c[1190]), .CLK(clk), .RST(rst), .Q(sreg[1189]) );
  DFF \sreg_reg[1188]  ( .D(c[1189]), .CLK(clk), .RST(rst), .Q(sreg[1188]) );
  DFF \sreg_reg[1187]  ( .D(c[1188]), .CLK(clk), .RST(rst), .Q(sreg[1187]) );
  DFF \sreg_reg[1186]  ( .D(c[1187]), .CLK(clk), .RST(rst), .Q(sreg[1186]) );
  DFF \sreg_reg[1185]  ( .D(c[1186]), .CLK(clk), .RST(rst), .Q(sreg[1185]) );
  DFF \sreg_reg[1184]  ( .D(c[1185]), .CLK(clk), .RST(rst), .Q(sreg[1184]) );
  DFF \sreg_reg[1183]  ( .D(c[1184]), .CLK(clk), .RST(rst), .Q(sreg[1183]) );
  DFF \sreg_reg[1182]  ( .D(c[1183]), .CLK(clk), .RST(rst), .Q(sreg[1182]) );
  DFF \sreg_reg[1181]  ( .D(c[1182]), .CLK(clk), .RST(rst), .Q(sreg[1181]) );
  DFF \sreg_reg[1180]  ( .D(c[1181]), .CLK(clk), .RST(rst), .Q(sreg[1180]) );
  DFF \sreg_reg[1179]  ( .D(c[1180]), .CLK(clk), .RST(rst), .Q(sreg[1179]) );
  DFF \sreg_reg[1178]  ( .D(c[1179]), .CLK(clk), .RST(rst), .Q(sreg[1178]) );
  DFF \sreg_reg[1177]  ( .D(c[1178]), .CLK(clk), .RST(rst), .Q(sreg[1177]) );
  DFF \sreg_reg[1176]  ( .D(c[1177]), .CLK(clk), .RST(rst), .Q(sreg[1176]) );
  DFF \sreg_reg[1175]  ( .D(c[1176]), .CLK(clk), .RST(rst), .Q(sreg[1175]) );
  DFF \sreg_reg[1174]  ( .D(c[1175]), .CLK(clk), .RST(rst), .Q(sreg[1174]) );
  DFF \sreg_reg[1173]  ( .D(c[1174]), .CLK(clk), .RST(rst), .Q(sreg[1173]) );
  DFF \sreg_reg[1172]  ( .D(c[1173]), .CLK(clk), .RST(rst), .Q(sreg[1172]) );
  DFF \sreg_reg[1171]  ( .D(c[1172]), .CLK(clk), .RST(rst), .Q(sreg[1171]) );
  DFF \sreg_reg[1170]  ( .D(c[1171]), .CLK(clk), .RST(rst), .Q(sreg[1170]) );
  DFF \sreg_reg[1169]  ( .D(c[1170]), .CLK(clk), .RST(rst), .Q(sreg[1169]) );
  DFF \sreg_reg[1168]  ( .D(c[1169]), .CLK(clk), .RST(rst), .Q(sreg[1168]) );
  DFF \sreg_reg[1167]  ( .D(c[1168]), .CLK(clk), .RST(rst), .Q(sreg[1167]) );
  DFF \sreg_reg[1166]  ( .D(c[1167]), .CLK(clk), .RST(rst), .Q(sreg[1166]) );
  DFF \sreg_reg[1165]  ( .D(c[1166]), .CLK(clk), .RST(rst), .Q(sreg[1165]) );
  DFF \sreg_reg[1164]  ( .D(c[1165]), .CLK(clk), .RST(rst), .Q(sreg[1164]) );
  DFF \sreg_reg[1163]  ( .D(c[1164]), .CLK(clk), .RST(rst), .Q(sreg[1163]) );
  DFF \sreg_reg[1162]  ( .D(c[1163]), .CLK(clk), .RST(rst), .Q(sreg[1162]) );
  DFF \sreg_reg[1161]  ( .D(c[1162]), .CLK(clk), .RST(rst), .Q(sreg[1161]) );
  DFF \sreg_reg[1160]  ( .D(c[1161]), .CLK(clk), .RST(rst), .Q(sreg[1160]) );
  DFF \sreg_reg[1159]  ( .D(c[1160]), .CLK(clk), .RST(rst), .Q(sreg[1159]) );
  DFF \sreg_reg[1158]  ( .D(c[1159]), .CLK(clk), .RST(rst), .Q(sreg[1158]) );
  DFF \sreg_reg[1157]  ( .D(c[1158]), .CLK(clk), .RST(rst), .Q(sreg[1157]) );
  DFF \sreg_reg[1156]  ( .D(c[1157]), .CLK(clk), .RST(rst), .Q(sreg[1156]) );
  DFF \sreg_reg[1155]  ( .D(c[1156]), .CLK(clk), .RST(rst), .Q(sreg[1155]) );
  DFF \sreg_reg[1154]  ( .D(c[1155]), .CLK(clk), .RST(rst), .Q(sreg[1154]) );
  DFF \sreg_reg[1153]  ( .D(c[1154]), .CLK(clk), .RST(rst), .Q(sreg[1153]) );
  DFF \sreg_reg[1152]  ( .D(c[1153]), .CLK(clk), .RST(rst), .Q(sreg[1152]) );
  DFF \sreg_reg[1151]  ( .D(c[1152]), .CLK(clk), .RST(rst), .Q(sreg[1151]) );
  DFF \sreg_reg[1150]  ( .D(c[1151]), .CLK(clk), .RST(rst), .Q(sreg[1150]) );
  DFF \sreg_reg[1149]  ( .D(c[1150]), .CLK(clk), .RST(rst), .Q(sreg[1149]) );
  DFF \sreg_reg[1148]  ( .D(c[1149]), .CLK(clk), .RST(rst), .Q(sreg[1148]) );
  DFF \sreg_reg[1147]  ( .D(c[1148]), .CLK(clk), .RST(rst), .Q(sreg[1147]) );
  DFF \sreg_reg[1146]  ( .D(c[1147]), .CLK(clk), .RST(rst), .Q(sreg[1146]) );
  DFF \sreg_reg[1145]  ( .D(c[1146]), .CLK(clk), .RST(rst), .Q(sreg[1145]) );
  DFF \sreg_reg[1144]  ( .D(c[1145]), .CLK(clk), .RST(rst), .Q(sreg[1144]) );
  DFF \sreg_reg[1143]  ( .D(c[1144]), .CLK(clk), .RST(rst), .Q(sreg[1143]) );
  DFF \sreg_reg[1142]  ( .D(c[1143]), .CLK(clk), .RST(rst), .Q(sreg[1142]) );
  DFF \sreg_reg[1141]  ( .D(c[1142]), .CLK(clk), .RST(rst), .Q(sreg[1141]) );
  DFF \sreg_reg[1140]  ( .D(c[1141]), .CLK(clk), .RST(rst), .Q(sreg[1140]) );
  DFF \sreg_reg[1139]  ( .D(c[1140]), .CLK(clk), .RST(rst), .Q(sreg[1139]) );
  DFF \sreg_reg[1138]  ( .D(c[1139]), .CLK(clk), .RST(rst), .Q(sreg[1138]) );
  DFF \sreg_reg[1137]  ( .D(c[1138]), .CLK(clk), .RST(rst), .Q(sreg[1137]) );
  DFF \sreg_reg[1136]  ( .D(c[1137]), .CLK(clk), .RST(rst), .Q(sreg[1136]) );
  DFF \sreg_reg[1135]  ( .D(c[1136]), .CLK(clk), .RST(rst), .Q(sreg[1135]) );
  DFF \sreg_reg[1134]  ( .D(c[1135]), .CLK(clk), .RST(rst), .Q(sreg[1134]) );
  DFF \sreg_reg[1133]  ( .D(c[1134]), .CLK(clk), .RST(rst), .Q(sreg[1133]) );
  DFF \sreg_reg[1132]  ( .D(c[1133]), .CLK(clk), .RST(rst), .Q(sreg[1132]) );
  DFF \sreg_reg[1131]  ( .D(c[1132]), .CLK(clk), .RST(rst), .Q(sreg[1131]) );
  DFF \sreg_reg[1130]  ( .D(c[1131]), .CLK(clk), .RST(rst), .Q(sreg[1130]) );
  DFF \sreg_reg[1129]  ( .D(c[1130]), .CLK(clk), .RST(rst), .Q(sreg[1129]) );
  DFF \sreg_reg[1128]  ( .D(c[1129]), .CLK(clk), .RST(rst), .Q(sreg[1128]) );
  DFF \sreg_reg[1127]  ( .D(c[1128]), .CLK(clk), .RST(rst), .Q(sreg[1127]) );
  DFF \sreg_reg[1126]  ( .D(c[1127]), .CLK(clk), .RST(rst), .Q(sreg[1126]) );
  DFF \sreg_reg[1125]  ( .D(c[1126]), .CLK(clk), .RST(rst), .Q(sreg[1125]) );
  DFF \sreg_reg[1124]  ( .D(c[1125]), .CLK(clk), .RST(rst), .Q(sreg[1124]) );
  DFF \sreg_reg[1123]  ( .D(c[1124]), .CLK(clk), .RST(rst), .Q(sreg[1123]) );
  DFF \sreg_reg[1122]  ( .D(c[1123]), .CLK(clk), .RST(rst), .Q(sreg[1122]) );
  DFF \sreg_reg[1121]  ( .D(c[1122]), .CLK(clk), .RST(rst), .Q(sreg[1121]) );
  DFF \sreg_reg[1120]  ( .D(c[1121]), .CLK(clk), .RST(rst), .Q(sreg[1120]) );
  DFF \sreg_reg[1119]  ( .D(c[1120]), .CLK(clk), .RST(rst), .Q(sreg[1119]) );
  DFF \sreg_reg[1118]  ( .D(c[1119]), .CLK(clk), .RST(rst), .Q(sreg[1118]) );
  DFF \sreg_reg[1117]  ( .D(c[1118]), .CLK(clk), .RST(rst), .Q(sreg[1117]) );
  DFF \sreg_reg[1116]  ( .D(c[1117]), .CLK(clk), .RST(rst), .Q(sreg[1116]) );
  DFF \sreg_reg[1115]  ( .D(c[1116]), .CLK(clk), .RST(rst), .Q(sreg[1115]) );
  DFF \sreg_reg[1114]  ( .D(c[1115]), .CLK(clk), .RST(rst), .Q(sreg[1114]) );
  DFF \sreg_reg[1113]  ( .D(c[1114]), .CLK(clk), .RST(rst), .Q(sreg[1113]) );
  DFF \sreg_reg[1112]  ( .D(c[1113]), .CLK(clk), .RST(rst), .Q(sreg[1112]) );
  DFF \sreg_reg[1111]  ( .D(c[1112]), .CLK(clk), .RST(rst), .Q(sreg[1111]) );
  DFF \sreg_reg[1110]  ( .D(c[1111]), .CLK(clk), .RST(rst), .Q(sreg[1110]) );
  DFF \sreg_reg[1109]  ( .D(c[1110]), .CLK(clk), .RST(rst), .Q(sreg[1109]) );
  DFF \sreg_reg[1108]  ( .D(c[1109]), .CLK(clk), .RST(rst), .Q(sreg[1108]) );
  DFF \sreg_reg[1107]  ( .D(c[1108]), .CLK(clk), .RST(rst), .Q(sreg[1107]) );
  DFF \sreg_reg[1106]  ( .D(c[1107]), .CLK(clk), .RST(rst), .Q(sreg[1106]) );
  DFF \sreg_reg[1105]  ( .D(c[1106]), .CLK(clk), .RST(rst), .Q(sreg[1105]) );
  DFF \sreg_reg[1104]  ( .D(c[1105]), .CLK(clk), .RST(rst), .Q(sreg[1104]) );
  DFF \sreg_reg[1103]  ( .D(c[1104]), .CLK(clk), .RST(rst), .Q(sreg[1103]) );
  DFF \sreg_reg[1102]  ( .D(c[1103]), .CLK(clk), .RST(rst), .Q(sreg[1102]) );
  DFF \sreg_reg[1101]  ( .D(c[1102]), .CLK(clk), .RST(rst), .Q(sreg[1101]) );
  DFF \sreg_reg[1100]  ( .D(c[1101]), .CLK(clk), .RST(rst), .Q(sreg[1100]) );
  DFF \sreg_reg[1099]  ( .D(c[1100]), .CLK(clk), .RST(rst), .Q(sreg[1099]) );
  DFF \sreg_reg[1098]  ( .D(c[1099]), .CLK(clk), .RST(rst), .Q(sreg[1098]) );
  DFF \sreg_reg[1097]  ( .D(c[1098]), .CLK(clk), .RST(rst), .Q(sreg[1097]) );
  DFF \sreg_reg[1096]  ( .D(c[1097]), .CLK(clk), .RST(rst), .Q(sreg[1096]) );
  DFF \sreg_reg[1095]  ( .D(c[1096]), .CLK(clk), .RST(rst), .Q(sreg[1095]) );
  DFF \sreg_reg[1094]  ( .D(c[1095]), .CLK(clk), .RST(rst), .Q(sreg[1094]) );
  DFF \sreg_reg[1093]  ( .D(c[1094]), .CLK(clk), .RST(rst), .Q(sreg[1093]) );
  DFF \sreg_reg[1092]  ( .D(c[1093]), .CLK(clk), .RST(rst), .Q(sreg[1092]) );
  DFF \sreg_reg[1091]  ( .D(c[1092]), .CLK(clk), .RST(rst), .Q(sreg[1091]) );
  DFF \sreg_reg[1090]  ( .D(c[1091]), .CLK(clk), .RST(rst), .Q(sreg[1090]) );
  DFF \sreg_reg[1089]  ( .D(c[1090]), .CLK(clk), .RST(rst), .Q(sreg[1089]) );
  DFF \sreg_reg[1088]  ( .D(c[1089]), .CLK(clk), .RST(rst), .Q(sreg[1088]) );
  DFF \sreg_reg[1087]  ( .D(c[1088]), .CLK(clk), .RST(rst), .Q(sreg[1087]) );
  DFF \sreg_reg[1086]  ( .D(c[1087]), .CLK(clk), .RST(rst), .Q(sreg[1086]) );
  DFF \sreg_reg[1085]  ( .D(c[1086]), .CLK(clk), .RST(rst), .Q(sreg[1085]) );
  DFF \sreg_reg[1084]  ( .D(c[1085]), .CLK(clk), .RST(rst), .Q(sreg[1084]) );
  DFF \sreg_reg[1083]  ( .D(c[1084]), .CLK(clk), .RST(rst), .Q(sreg[1083]) );
  DFF \sreg_reg[1082]  ( .D(c[1083]), .CLK(clk), .RST(rst), .Q(sreg[1082]) );
  DFF \sreg_reg[1081]  ( .D(c[1082]), .CLK(clk), .RST(rst), .Q(sreg[1081]) );
  DFF \sreg_reg[1080]  ( .D(c[1081]), .CLK(clk), .RST(rst), .Q(sreg[1080]) );
  DFF \sreg_reg[1079]  ( .D(c[1080]), .CLK(clk), .RST(rst), .Q(sreg[1079]) );
  DFF \sreg_reg[1078]  ( .D(c[1079]), .CLK(clk), .RST(rst), .Q(sreg[1078]) );
  DFF \sreg_reg[1077]  ( .D(c[1078]), .CLK(clk), .RST(rst), .Q(sreg[1077]) );
  DFF \sreg_reg[1076]  ( .D(c[1077]), .CLK(clk), .RST(rst), .Q(sreg[1076]) );
  DFF \sreg_reg[1075]  ( .D(c[1076]), .CLK(clk), .RST(rst), .Q(sreg[1075]) );
  DFF \sreg_reg[1074]  ( .D(c[1075]), .CLK(clk), .RST(rst), .Q(sreg[1074]) );
  DFF \sreg_reg[1073]  ( .D(c[1074]), .CLK(clk), .RST(rst), .Q(sreg[1073]) );
  DFF \sreg_reg[1072]  ( .D(c[1073]), .CLK(clk), .RST(rst), .Q(sreg[1072]) );
  DFF \sreg_reg[1071]  ( .D(c[1072]), .CLK(clk), .RST(rst), .Q(sreg[1071]) );
  DFF \sreg_reg[1070]  ( .D(c[1071]), .CLK(clk), .RST(rst), .Q(sreg[1070]) );
  DFF \sreg_reg[1069]  ( .D(c[1070]), .CLK(clk), .RST(rst), .Q(sreg[1069]) );
  DFF \sreg_reg[1068]  ( .D(c[1069]), .CLK(clk), .RST(rst), .Q(sreg[1068]) );
  DFF \sreg_reg[1067]  ( .D(c[1068]), .CLK(clk), .RST(rst), .Q(sreg[1067]) );
  DFF \sreg_reg[1066]  ( .D(c[1067]), .CLK(clk), .RST(rst), .Q(sreg[1066]) );
  DFF \sreg_reg[1065]  ( .D(c[1066]), .CLK(clk), .RST(rst), .Q(sreg[1065]) );
  DFF \sreg_reg[1064]  ( .D(c[1065]), .CLK(clk), .RST(rst), .Q(sreg[1064]) );
  DFF \sreg_reg[1063]  ( .D(c[1064]), .CLK(clk), .RST(rst), .Q(sreg[1063]) );
  DFF \sreg_reg[1062]  ( .D(c[1063]), .CLK(clk), .RST(rst), .Q(sreg[1062]) );
  DFF \sreg_reg[1061]  ( .D(c[1062]), .CLK(clk), .RST(rst), .Q(sreg[1061]) );
  DFF \sreg_reg[1060]  ( .D(c[1061]), .CLK(clk), .RST(rst), .Q(sreg[1060]) );
  DFF \sreg_reg[1059]  ( .D(c[1060]), .CLK(clk), .RST(rst), .Q(sreg[1059]) );
  DFF \sreg_reg[1058]  ( .D(c[1059]), .CLK(clk), .RST(rst), .Q(sreg[1058]) );
  DFF \sreg_reg[1057]  ( .D(c[1058]), .CLK(clk), .RST(rst), .Q(sreg[1057]) );
  DFF \sreg_reg[1056]  ( .D(c[1057]), .CLK(clk), .RST(rst), .Q(sreg[1056]) );
  DFF \sreg_reg[1055]  ( .D(c[1056]), .CLK(clk), .RST(rst), .Q(sreg[1055]) );
  DFF \sreg_reg[1054]  ( .D(c[1055]), .CLK(clk), .RST(rst), .Q(sreg[1054]) );
  DFF \sreg_reg[1053]  ( .D(c[1054]), .CLK(clk), .RST(rst), .Q(sreg[1053]) );
  DFF \sreg_reg[1052]  ( .D(c[1053]), .CLK(clk), .RST(rst), .Q(sreg[1052]) );
  DFF \sreg_reg[1051]  ( .D(c[1052]), .CLK(clk), .RST(rst), .Q(sreg[1051]) );
  DFF \sreg_reg[1050]  ( .D(c[1051]), .CLK(clk), .RST(rst), .Q(sreg[1050]) );
  DFF \sreg_reg[1049]  ( .D(c[1050]), .CLK(clk), .RST(rst), .Q(sreg[1049]) );
  DFF \sreg_reg[1048]  ( .D(c[1049]), .CLK(clk), .RST(rst), .Q(sreg[1048]) );
  DFF \sreg_reg[1047]  ( .D(c[1048]), .CLK(clk), .RST(rst), .Q(sreg[1047]) );
  DFF \sreg_reg[1046]  ( .D(c[1047]), .CLK(clk), .RST(rst), .Q(sreg[1046]) );
  DFF \sreg_reg[1045]  ( .D(c[1046]), .CLK(clk), .RST(rst), .Q(sreg[1045]) );
  DFF \sreg_reg[1044]  ( .D(c[1045]), .CLK(clk), .RST(rst), .Q(sreg[1044]) );
  DFF \sreg_reg[1043]  ( .D(c[1044]), .CLK(clk), .RST(rst), .Q(sreg[1043]) );
  DFF \sreg_reg[1042]  ( .D(c[1043]), .CLK(clk), .RST(rst), .Q(sreg[1042]) );
  DFF \sreg_reg[1041]  ( .D(c[1042]), .CLK(clk), .RST(rst), .Q(sreg[1041]) );
  DFF \sreg_reg[1040]  ( .D(c[1041]), .CLK(clk), .RST(rst), .Q(sreg[1040]) );
  DFF \sreg_reg[1039]  ( .D(c[1040]), .CLK(clk), .RST(rst), .Q(sreg[1039]) );
  DFF \sreg_reg[1038]  ( .D(c[1039]), .CLK(clk), .RST(rst), .Q(sreg[1038]) );
  DFF \sreg_reg[1037]  ( .D(c[1038]), .CLK(clk), .RST(rst), .Q(sreg[1037]) );
  DFF \sreg_reg[1036]  ( .D(c[1037]), .CLK(clk), .RST(rst), .Q(sreg[1036]) );
  DFF \sreg_reg[1035]  ( .D(c[1036]), .CLK(clk), .RST(rst), .Q(sreg[1035]) );
  DFF \sreg_reg[1034]  ( .D(c[1035]), .CLK(clk), .RST(rst), .Q(sreg[1034]) );
  DFF \sreg_reg[1033]  ( .D(c[1034]), .CLK(clk), .RST(rst), .Q(sreg[1033]) );
  DFF \sreg_reg[1032]  ( .D(c[1033]), .CLK(clk), .RST(rst), .Q(sreg[1032]) );
  DFF \sreg_reg[1031]  ( .D(c[1032]), .CLK(clk), .RST(rst), .Q(sreg[1031]) );
  DFF \sreg_reg[1030]  ( .D(c[1031]), .CLK(clk), .RST(rst), .Q(sreg[1030]) );
  DFF \sreg_reg[1029]  ( .D(c[1030]), .CLK(clk), .RST(rst), .Q(sreg[1029]) );
  DFF \sreg_reg[1028]  ( .D(c[1029]), .CLK(clk), .RST(rst), .Q(sreg[1028]) );
  DFF \sreg_reg[1027]  ( .D(c[1028]), .CLK(clk), .RST(rst), .Q(sreg[1027]) );
  DFF \sreg_reg[1026]  ( .D(c[1027]), .CLK(clk), .RST(rst), .Q(sreg[1026]) );
  DFF \sreg_reg[1025]  ( .D(c[1026]), .CLK(clk), .RST(rst), .Q(sreg[1025]) );
  DFF \sreg_reg[1024]  ( .D(c[1025]), .CLK(clk), .RST(rst), .Q(sreg[1024]) );
  DFF \sreg_reg[1023]  ( .D(c[1024]), .CLK(clk), .RST(rst), .Q(sreg[1023]) );
  DFF \sreg_reg[1022]  ( .D(c[1023]), .CLK(clk), .RST(rst), .Q(c[1022]) );
  DFF \sreg_reg[1021]  ( .D(c[1022]), .CLK(clk), .RST(rst), .Q(c[1021]) );
  DFF \sreg_reg[1020]  ( .D(c[1021]), .CLK(clk), .RST(rst), .Q(c[1020]) );
  DFF \sreg_reg[1019]  ( .D(c[1020]), .CLK(clk), .RST(rst), .Q(c[1019]) );
  DFF \sreg_reg[1018]  ( .D(c[1019]), .CLK(clk), .RST(rst), .Q(c[1018]) );
  DFF \sreg_reg[1017]  ( .D(c[1018]), .CLK(clk), .RST(rst), .Q(c[1017]) );
  DFF \sreg_reg[1016]  ( .D(c[1017]), .CLK(clk), .RST(rst), .Q(c[1016]) );
  DFF \sreg_reg[1015]  ( .D(c[1016]), .CLK(clk), .RST(rst), .Q(c[1015]) );
  DFF \sreg_reg[1014]  ( .D(c[1015]), .CLK(clk), .RST(rst), .Q(c[1014]) );
  DFF \sreg_reg[1013]  ( .D(c[1014]), .CLK(clk), .RST(rst), .Q(c[1013]) );
  DFF \sreg_reg[1012]  ( .D(c[1013]), .CLK(clk), .RST(rst), .Q(c[1012]) );
  DFF \sreg_reg[1011]  ( .D(c[1012]), .CLK(clk), .RST(rst), .Q(c[1011]) );
  DFF \sreg_reg[1010]  ( .D(c[1011]), .CLK(clk), .RST(rst), .Q(c[1010]) );
  DFF \sreg_reg[1009]  ( .D(c[1010]), .CLK(clk), .RST(rst), .Q(c[1009]) );
  DFF \sreg_reg[1008]  ( .D(c[1009]), .CLK(clk), .RST(rst), .Q(c[1008]) );
  DFF \sreg_reg[1007]  ( .D(c[1008]), .CLK(clk), .RST(rst), .Q(c[1007]) );
  DFF \sreg_reg[1006]  ( .D(c[1007]), .CLK(clk), .RST(rst), .Q(c[1006]) );
  DFF \sreg_reg[1005]  ( .D(c[1006]), .CLK(clk), .RST(rst), .Q(c[1005]) );
  DFF \sreg_reg[1004]  ( .D(c[1005]), .CLK(clk), .RST(rst), .Q(c[1004]) );
  DFF \sreg_reg[1003]  ( .D(c[1004]), .CLK(clk), .RST(rst), .Q(c[1003]) );
  DFF \sreg_reg[1002]  ( .D(c[1003]), .CLK(clk), .RST(rst), .Q(c[1002]) );
  DFF \sreg_reg[1001]  ( .D(c[1002]), .CLK(clk), .RST(rst), .Q(c[1001]) );
  DFF \sreg_reg[1000]  ( .D(c[1001]), .CLK(clk), .RST(rst), .Q(c[1000]) );
  DFF \sreg_reg[999]  ( .D(c[1000]), .CLK(clk), .RST(rst), .Q(c[999]) );
  DFF \sreg_reg[998]  ( .D(c[999]), .CLK(clk), .RST(rst), .Q(c[998]) );
  DFF \sreg_reg[997]  ( .D(c[998]), .CLK(clk), .RST(rst), .Q(c[997]) );
  DFF \sreg_reg[996]  ( .D(c[997]), .CLK(clk), .RST(rst), .Q(c[996]) );
  DFF \sreg_reg[995]  ( .D(c[996]), .CLK(clk), .RST(rst), .Q(c[995]) );
  DFF \sreg_reg[994]  ( .D(c[995]), .CLK(clk), .RST(rst), .Q(c[994]) );
  DFF \sreg_reg[993]  ( .D(c[994]), .CLK(clk), .RST(rst), .Q(c[993]) );
  DFF \sreg_reg[992]  ( .D(c[993]), .CLK(clk), .RST(rst), .Q(c[992]) );
  DFF \sreg_reg[991]  ( .D(c[992]), .CLK(clk), .RST(rst), .Q(c[991]) );
  DFF \sreg_reg[990]  ( .D(c[991]), .CLK(clk), .RST(rst), .Q(c[990]) );
  DFF \sreg_reg[989]  ( .D(c[990]), .CLK(clk), .RST(rst), .Q(c[989]) );
  DFF \sreg_reg[988]  ( .D(c[989]), .CLK(clk), .RST(rst), .Q(c[988]) );
  DFF \sreg_reg[987]  ( .D(c[988]), .CLK(clk), .RST(rst), .Q(c[987]) );
  DFF \sreg_reg[986]  ( .D(c[987]), .CLK(clk), .RST(rst), .Q(c[986]) );
  DFF \sreg_reg[985]  ( .D(c[986]), .CLK(clk), .RST(rst), .Q(c[985]) );
  DFF \sreg_reg[984]  ( .D(c[985]), .CLK(clk), .RST(rst), .Q(c[984]) );
  DFF \sreg_reg[983]  ( .D(c[984]), .CLK(clk), .RST(rst), .Q(c[983]) );
  DFF \sreg_reg[982]  ( .D(c[983]), .CLK(clk), .RST(rst), .Q(c[982]) );
  DFF \sreg_reg[981]  ( .D(c[982]), .CLK(clk), .RST(rst), .Q(c[981]) );
  DFF \sreg_reg[980]  ( .D(c[981]), .CLK(clk), .RST(rst), .Q(c[980]) );
  DFF \sreg_reg[979]  ( .D(c[980]), .CLK(clk), .RST(rst), .Q(c[979]) );
  DFF \sreg_reg[978]  ( .D(c[979]), .CLK(clk), .RST(rst), .Q(c[978]) );
  DFF \sreg_reg[977]  ( .D(c[978]), .CLK(clk), .RST(rst), .Q(c[977]) );
  DFF \sreg_reg[976]  ( .D(c[977]), .CLK(clk), .RST(rst), .Q(c[976]) );
  DFF \sreg_reg[975]  ( .D(c[976]), .CLK(clk), .RST(rst), .Q(c[975]) );
  DFF \sreg_reg[974]  ( .D(c[975]), .CLK(clk), .RST(rst), .Q(c[974]) );
  DFF \sreg_reg[973]  ( .D(c[974]), .CLK(clk), .RST(rst), .Q(c[973]) );
  DFF \sreg_reg[972]  ( .D(c[973]), .CLK(clk), .RST(rst), .Q(c[972]) );
  DFF \sreg_reg[971]  ( .D(c[972]), .CLK(clk), .RST(rst), .Q(c[971]) );
  DFF \sreg_reg[970]  ( .D(c[971]), .CLK(clk), .RST(rst), .Q(c[970]) );
  DFF \sreg_reg[969]  ( .D(c[970]), .CLK(clk), .RST(rst), .Q(c[969]) );
  DFF \sreg_reg[968]  ( .D(c[969]), .CLK(clk), .RST(rst), .Q(c[968]) );
  DFF \sreg_reg[967]  ( .D(c[968]), .CLK(clk), .RST(rst), .Q(c[967]) );
  DFF \sreg_reg[966]  ( .D(c[967]), .CLK(clk), .RST(rst), .Q(c[966]) );
  DFF \sreg_reg[965]  ( .D(c[966]), .CLK(clk), .RST(rst), .Q(c[965]) );
  DFF \sreg_reg[964]  ( .D(c[965]), .CLK(clk), .RST(rst), .Q(c[964]) );
  DFF \sreg_reg[963]  ( .D(c[964]), .CLK(clk), .RST(rst), .Q(c[963]) );
  DFF \sreg_reg[962]  ( .D(c[963]), .CLK(clk), .RST(rst), .Q(c[962]) );
  DFF \sreg_reg[961]  ( .D(c[962]), .CLK(clk), .RST(rst), .Q(c[961]) );
  DFF \sreg_reg[960]  ( .D(c[961]), .CLK(clk), .RST(rst), .Q(c[960]) );
  DFF \sreg_reg[959]  ( .D(c[960]), .CLK(clk), .RST(rst), .Q(c[959]) );
  DFF \sreg_reg[958]  ( .D(c[959]), .CLK(clk), .RST(rst), .Q(c[958]) );
  DFF \sreg_reg[957]  ( .D(c[958]), .CLK(clk), .RST(rst), .Q(c[957]) );
  DFF \sreg_reg[956]  ( .D(c[957]), .CLK(clk), .RST(rst), .Q(c[956]) );
  DFF \sreg_reg[955]  ( .D(c[956]), .CLK(clk), .RST(rst), .Q(c[955]) );
  DFF \sreg_reg[954]  ( .D(c[955]), .CLK(clk), .RST(rst), .Q(c[954]) );
  DFF \sreg_reg[953]  ( .D(c[954]), .CLK(clk), .RST(rst), .Q(c[953]) );
  DFF \sreg_reg[952]  ( .D(c[953]), .CLK(clk), .RST(rst), .Q(c[952]) );
  DFF \sreg_reg[951]  ( .D(c[952]), .CLK(clk), .RST(rst), .Q(c[951]) );
  DFF \sreg_reg[950]  ( .D(c[951]), .CLK(clk), .RST(rst), .Q(c[950]) );
  DFF \sreg_reg[949]  ( .D(c[950]), .CLK(clk), .RST(rst), .Q(c[949]) );
  DFF \sreg_reg[948]  ( .D(c[949]), .CLK(clk), .RST(rst), .Q(c[948]) );
  DFF \sreg_reg[947]  ( .D(c[948]), .CLK(clk), .RST(rst), .Q(c[947]) );
  DFF \sreg_reg[946]  ( .D(c[947]), .CLK(clk), .RST(rst), .Q(c[946]) );
  DFF \sreg_reg[945]  ( .D(c[946]), .CLK(clk), .RST(rst), .Q(c[945]) );
  DFF \sreg_reg[944]  ( .D(c[945]), .CLK(clk), .RST(rst), .Q(c[944]) );
  DFF \sreg_reg[943]  ( .D(c[944]), .CLK(clk), .RST(rst), .Q(c[943]) );
  DFF \sreg_reg[942]  ( .D(c[943]), .CLK(clk), .RST(rst), .Q(c[942]) );
  DFF \sreg_reg[941]  ( .D(c[942]), .CLK(clk), .RST(rst), .Q(c[941]) );
  DFF \sreg_reg[940]  ( .D(c[941]), .CLK(clk), .RST(rst), .Q(c[940]) );
  DFF \sreg_reg[939]  ( .D(c[940]), .CLK(clk), .RST(rst), .Q(c[939]) );
  DFF \sreg_reg[938]  ( .D(c[939]), .CLK(clk), .RST(rst), .Q(c[938]) );
  DFF \sreg_reg[937]  ( .D(c[938]), .CLK(clk), .RST(rst), .Q(c[937]) );
  DFF \sreg_reg[936]  ( .D(c[937]), .CLK(clk), .RST(rst), .Q(c[936]) );
  DFF \sreg_reg[935]  ( .D(c[936]), .CLK(clk), .RST(rst), .Q(c[935]) );
  DFF \sreg_reg[934]  ( .D(c[935]), .CLK(clk), .RST(rst), .Q(c[934]) );
  DFF \sreg_reg[933]  ( .D(c[934]), .CLK(clk), .RST(rst), .Q(c[933]) );
  DFF \sreg_reg[932]  ( .D(c[933]), .CLK(clk), .RST(rst), .Q(c[932]) );
  DFF \sreg_reg[931]  ( .D(c[932]), .CLK(clk), .RST(rst), .Q(c[931]) );
  DFF \sreg_reg[930]  ( .D(c[931]), .CLK(clk), .RST(rst), .Q(c[930]) );
  DFF \sreg_reg[929]  ( .D(c[930]), .CLK(clk), .RST(rst), .Q(c[929]) );
  DFF \sreg_reg[928]  ( .D(c[929]), .CLK(clk), .RST(rst), .Q(c[928]) );
  DFF \sreg_reg[927]  ( .D(c[928]), .CLK(clk), .RST(rst), .Q(c[927]) );
  DFF \sreg_reg[926]  ( .D(c[927]), .CLK(clk), .RST(rst), .Q(c[926]) );
  DFF \sreg_reg[925]  ( .D(c[926]), .CLK(clk), .RST(rst), .Q(c[925]) );
  DFF \sreg_reg[924]  ( .D(c[925]), .CLK(clk), .RST(rst), .Q(c[924]) );
  DFF \sreg_reg[923]  ( .D(c[924]), .CLK(clk), .RST(rst), .Q(c[923]) );
  DFF \sreg_reg[922]  ( .D(c[923]), .CLK(clk), .RST(rst), .Q(c[922]) );
  DFF \sreg_reg[921]  ( .D(c[922]), .CLK(clk), .RST(rst), .Q(c[921]) );
  DFF \sreg_reg[920]  ( .D(c[921]), .CLK(clk), .RST(rst), .Q(c[920]) );
  DFF \sreg_reg[919]  ( .D(c[920]), .CLK(clk), .RST(rst), .Q(c[919]) );
  DFF \sreg_reg[918]  ( .D(c[919]), .CLK(clk), .RST(rst), .Q(c[918]) );
  DFF \sreg_reg[917]  ( .D(c[918]), .CLK(clk), .RST(rst), .Q(c[917]) );
  DFF \sreg_reg[916]  ( .D(c[917]), .CLK(clk), .RST(rst), .Q(c[916]) );
  DFF \sreg_reg[915]  ( .D(c[916]), .CLK(clk), .RST(rst), .Q(c[915]) );
  DFF \sreg_reg[914]  ( .D(c[915]), .CLK(clk), .RST(rst), .Q(c[914]) );
  DFF \sreg_reg[913]  ( .D(c[914]), .CLK(clk), .RST(rst), .Q(c[913]) );
  DFF \sreg_reg[912]  ( .D(c[913]), .CLK(clk), .RST(rst), .Q(c[912]) );
  DFF \sreg_reg[911]  ( .D(c[912]), .CLK(clk), .RST(rst), .Q(c[911]) );
  DFF \sreg_reg[910]  ( .D(c[911]), .CLK(clk), .RST(rst), .Q(c[910]) );
  DFF \sreg_reg[909]  ( .D(c[910]), .CLK(clk), .RST(rst), .Q(c[909]) );
  DFF \sreg_reg[908]  ( .D(c[909]), .CLK(clk), .RST(rst), .Q(c[908]) );
  DFF \sreg_reg[907]  ( .D(c[908]), .CLK(clk), .RST(rst), .Q(c[907]) );
  DFF \sreg_reg[906]  ( .D(c[907]), .CLK(clk), .RST(rst), .Q(c[906]) );
  DFF \sreg_reg[905]  ( .D(c[906]), .CLK(clk), .RST(rst), .Q(c[905]) );
  DFF \sreg_reg[904]  ( .D(c[905]), .CLK(clk), .RST(rst), .Q(c[904]) );
  DFF \sreg_reg[903]  ( .D(c[904]), .CLK(clk), .RST(rst), .Q(c[903]) );
  DFF \sreg_reg[902]  ( .D(c[903]), .CLK(clk), .RST(rst), .Q(c[902]) );
  DFF \sreg_reg[901]  ( .D(c[902]), .CLK(clk), .RST(rst), .Q(c[901]) );
  DFF \sreg_reg[900]  ( .D(c[901]), .CLK(clk), .RST(rst), .Q(c[900]) );
  DFF \sreg_reg[899]  ( .D(c[900]), .CLK(clk), .RST(rst), .Q(c[899]) );
  DFF \sreg_reg[898]  ( .D(c[899]), .CLK(clk), .RST(rst), .Q(c[898]) );
  DFF \sreg_reg[897]  ( .D(c[898]), .CLK(clk), .RST(rst), .Q(c[897]) );
  DFF \sreg_reg[896]  ( .D(c[897]), .CLK(clk), .RST(rst), .Q(c[896]) );
  DFF \sreg_reg[895]  ( .D(c[896]), .CLK(clk), .RST(rst), .Q(c[895]) );
  DFF \sreg_reg[894]  ( .D(c[895]), .CLK(clk), .RST(rst), .Q(c[894]) );
  DFF \sreg_reg[893]  ( .D(c[894]), .CLK(clk), .RST(rst), .Q(c[893]) );
  DFF \sreg_reg[892]  ( .D(c[893]), .CLK(clk), .RST(rst), .Q(c[892]) );
  DFF \sreg_reg[891]  ( .D(c[892]), .CLK(clk), .RST(rst), .Q(c[891]) );
  DFF \sreg_reg[890]  ( .D(c[891]), .CLK(clk), .RST(rst), .Q(c[890]) );
  DFF \sreg_reg[889]  ( .D(c[890]), .CLK(clk), .RST(rst), .Q(c[889]) );
  DFF \sreg_reg[888]  ( .D(c[889]), .CLK(clk), .RST(rst), .Q(c[888]) );
  DFF \sreg_reg[887]  ( .D(c[888]), .CLK(clk), .RST(rst), .Q(c[887]) );
  DFF \sreg_reg[886]  ( .D(c[887]), .CLK(clk), .RST(rst), .Q(c[886]) );
  DFF \sreg_reg[885]  ( .D(c[886]), .CLK(clk), .RST(rst), .Q(c[885]) );
  DFF \sreg_reg[884]  ( .D(c[885]), .CLK(clk), .RST(rst), .Q(c[884]) );
  DFF \sreg_reg[883]  ( .D(c[884]), .CLK(clk), .RST(rst), .Q(c[883]) );
  DFF \sreg_reg[882]  ( .D(c[883]), .CLK(clk), .RST(rst), .Q(c[882]) );
  DFF \sreg_reg[881]  ( .D(c[882]), .CLK(clk), .RST(rst), .Q(c[881]) );
  DFF \sreg_reg[880]  ( .D(c[881]), .CLK(clk), .RST(rst), .Q(c[880]) );
  DFF \sreg_reg[879]  ( .D(c[880]), .CLK(clk), .RST(rst), .Q(c[879]) );
  DFF \sreg_reg[878]  ( .D(c[879]), .CLK(clk), .RST(rst), .Q(c[878]) );
  DFF \sreg_reg[877]  ( .D(c[878]), .CLK(clk), .RST(rst), .Q(c[877]) );
  DFF \sreg_reg[876]  ( .D(c[877]), .CLK(clk), .RST(rst), .Q(c[876]) );
  DFF \sreg_reg[875]  ( .D(c[876]), .CLK(clk), .RST(rst), .Q(c[875]) );
  DFF \sreg_reg[874]  ( .D(c[875]), .CLK(clk), .RST(rst), .Q(c[874]) );
  DFF \sreg_reg[873]  ( .D(c[874]), .CLK(clk), .RST(rst), .Q(c[873]) );
  DFF \sreg_reg[872]  ( .D(c[873]), .CLK(clk), .RST(rst), .Q(c[872]) );
  DFF \sreg_reg[871]  ( .D(c[872]), .CLK(clk), .RST(rst), .Q(c[871]) );
  DFF \sreg_reg[870]  ( .D(c[871]), .CLK(clk), .RST(rst), .Q(c[870]) );
  DFF \sreg_reg[869]  ( .D(c[870]), .CLK(clk), .RST(rst), .Q(c[869]) );
  DFF \sreg_reg[868]  ( .D(c[869]), .CLK(clk), .RST(rst), .Q(c[868]) );
  DFF \sreg_reg[867]  ( .D(c[868]), .CLK(clk), .RST(rst), .Q(c[867]) );
  DFF \sreg_reg[866]  ( .D(c[867]), .CLK(clk), .RST(rst), .Q(c[866]) );
  DFF \sreg_reg[865]  ( .D(c[866]), .CLK(clk), .RST(rst), .Q(c[865]) );
  DFF \sreg_reg[864]  ( .D(c[865]), .CLK(clk), .RST(rst), .Q(c[864]) );
  DFF \sreg_reg[863]  ( .D(c[864]), .CLK(clk), .RST(rst), .Q(c[863]) );
  DFF \sreg_reg[862]  ( .D(c[863]), .CLK(clk), .RST(rst), .Q(c[862]) );
  DFF \sreg_reg[861]  ( .D(c[862]), .CLK(clk), .RST(rst), .Q(c[861]) );
  DFF \sreg_reg[860]  ( .D(c[861]), .CLK(clk), .RST(rst), .Q(c[860]) );
  DFF \sreg_reg[859]  ( .D(c[860]), .CLK(clk), .RST(rst), .Q(c[859]) );
  DFF \sreg_reg[858]  ( .D(c[859]), .CLK(clk), .RST(rst), .Q(c[858]) );
  DFF \sreg_reg[857]  ( .D(c[858]), .CLK(clk), .RST(rst), .Q(c[857]) );
  DFF \sreg_reg[856]  ( .D(c[857]), .CLK(clk), .RST(rst), .Q(c[856]) );
  DFF \sreg_reg[855]  ( .D(c[856]), .CLK(clk), .RST(rst), .Q(c[855]) );
  DFF \sreg_reg[854]  ( .D(c[855]), .CLK(clk), .RST(rst), .Q(c[854]) );
  DFF \sreg_reg[853]  ( .D(c[854]), .CLK(clk), .RST(rst), .Q(c[853]) );
  DFF \sreg_reg[852]  ( .D(c[853]), .CLK(clk), .RST(rst), .Q(c[852]) );
  DFF \sreg_reg[851]  ( .D(c[852]), .CLK(clk), .RST(rst), .Q(c[851]) );
  DFF \sreg_reg[850]  ( .D(c[851]), .CLK(clk), .RST(rst), .Q(c[850]) );
  DFF \sreg_reg[849]  ( .D(c[850]), .CLK(clk), .RST(rst), .Q(c[849]) );
  DFF \sreg_reg[848]  ( .D(c[849]), .CLK(clk), .RST(rst), .Q(c[848]) );
  DFF \sreg_reg[847]  ( .D(c[848]), .CLK(clk), .RST(rst), .Q(c[847]) );
  DFF \sreg_reg[846]  ( .D(c[847]), .CLK(clk), .RST(rst), .Q(c[846]) );
  DFF \sreg_reg[845]  ( .D(c[846]), .CLK(clk), .RST(rst), .Q(c[845]) );
  DFF \sreg_reg[844]  ( .D(c[845]), .CLK(clk), .RST(rst), .Q(c[844]) );
  DFF \sreg_reg[843]  ( .D(c[844]), .CLK(clk), .RST(rst), .Q(c[843]) );
  DFF \sreg_reg[842]  ( .D(c[843]), .CLK(clk), .RST(rst), .Q(c[842]) );
  DFF \sreg_reg[841]  ( .D(c[842]), .CLK(clk), .RST(rst), .Q(c[841]) );
  DFF \sreg_reg[840]  ( .D(c[841]), .CLK(clk), .RST(rst), .Q(c[840]) );
  DFF \sreg_reg[839]  ( .D(c[840]), .CLK(clk), .RST(rst), .Q(c[839]) );
  DFF \sreg_reg[838]  ( .D(c[839]), .CLK(clk), .RST(rst), .Q(c[838]) );
  DFF \sreg_reg[837]  ( .D(c[838]), .CLK(clk), .RST(rst), .Q(c[837]) );
  DFF \sreg_reg[836]  ( .D(c[837]), .CLK(clk), .RST(rst), .Q(c[836]) );
  DFF \sreg_reg[835]  ( .D(c[836]), .CLK(clk), .RST(rst), .Q(c[835]) );
  DFF \sreg_reg[834]  ( .D(c[835]), .CLK(clk), .RST(rst), .Q(c[834]) );
  DFF \sreg_reg[833]  ( .D(c[834]), .CLK(clk), .RST(rst), .Q(c[833]) );
  DFF \sreg_reg[832]  ( .D(c[833]), .CLK(clk), .RST(rst), .Q(c[832]) );
  DFF \sreg_reg[831]  ( .D(c[832]), .CLK(clk), .RST(rst), .Q(c[831]) );
  DFF \sreg_reg[830]  ( .D(c[831]), .CLK(clk), .RST(rst), .Q(c[830]) );
  DFF \sreg_reg[829]  ( .D(c[830]), .CLK(clk), .RST(rst), .Q(c[829]) );
  DFF \sreg_reg[828]  ( .D(c[829]), .CLK(clk), .RST(rst), .Q(c[828]) );
  DFF \sreg_reg[827]  ( .D(c[828]), .CLK(clk), .RST(rst), .Q(c[827]) );
  DFF \sreg_reg[826]  ( .D(c[827]), .CLK(clk), .RST(rst), .Q(c[826]) );
  DFF \sreg_reg[825]  ( .D(c[826]), .CLK(clk), .RST(rst), .Q(c[825]) );
  DFF \sreg_reg[824]  ( .D(c[825]), .CLK(clk), .RST(rst), .Q(c[824]) );
  DFF \sreg_reg[823]  ( .D(c[824]), .CLK(clk), .RST(rst), .Q(c[823]) );
  DFF \sreg_reg[822]  ( .D(c[823]), .CLK(clk), .RST(rst), .Q(c[822]) );
  DFF \sreg_reg[821]  ( .D(c[822]), .CLK(clk), .RST(rst), .Q(c[821]) );
  DFF \sreg_reg[820]  ( .D(c[821]), .CLK(clk), .RST(rst), .Q(c[820]) );
  DFF \sreg_reg[819]  ( .D(c[820]), .CLK(clk), .RST(rst), .Q(c[819]) );
  DFF \sreg_reg[818]  ( .D(c[819]), .CLK(clk), .RST(rst), .Q(c[818]) );
  DFF \sreg_reg[817]  ( .D(c[818]), .CLK(clk), .RST(rst), .Q(c[817]) );
  DFF \sreg_reg[816]  ( .D(c[817]), .CLK(clk), .RST(rst), .Q(c[816]) );
  DFF \sreg_reg[815]  ( .D(c[816]), .CLK(clk), .RST(rst), .Q(c[815]) );
  DFF \sreg_reg[814]  ( .D(c[815]), .CLK(clk), .RST(rst), .Q(c[814]) );
  DFF \sreg_reg[813]  ( .D(c[814]), .CLK(clk), .RST(rst), .Q(c[813]) );
  DFF \sreg_reg[812]  ( .D(c[813]), .CLK(clk), .RST(rst), .Q(c[812]) );
  DFF \sreg_reg[811]  ( .D(c[812]), .CLK(clk), .RST(rst), .Q(c[811]) );
  DFF \sreg_reg[810]  ( .D(c[811]), .CLK(clk), .RST(rst), .Q(c[810]) );
  DFF \sreg_reg[809]  ( .D(c[810]), .CLK(clk), .RST(rst), .Q(c[809]) );
  DFF \sreg_reg[808]  ( .D(c[809]), .CLK(clk), .RST(rst), .Q(c[808]) );
  DFF \sreg_reg[807]  ( .D(c[808]), .CLK(clk), .RST(rst), .Q(c[807]) );
  DFF \sreg_reg[806]  ( .D(c[807]), .CLK(clk), .RST(rst), .Q(c[806]) );
  DFF \sreg_reg[805]  ( .D(c[806]), .CLK(clk), .RST(rst), .Q(c[805]) );
  DFF \sreg_reg[804]  ( .D(c[805]), .CLK(clk), .RST(rst), .Q(c[804]) );
  DFF \sreg_reg[803]  ( .D(c[804]), .CLK(clk), .RST(rst), .Q(c[803]) );
  DFF \sreg_reg[802]  ( .D(c[803]), .CLK(clk), .RST(rst), .Q(c[802]) );
  DFF \sreg_reg[801]  ( .D(c[802]), .CLK(clk), .RST(rst), .Q(c[801]) );
  DFF \sreg_reg[800]  ( .D(c[801]), .CLK(clk), .RST(rst), .Q(c[800]) );
  DFF \sreg_reg[799]  ( .D(c[800]), .CLK(clk), .RST(rst), .Q(c[799]) );
  DFF \sreg_reg[798]  ( .D(c[799]), .CLK(clk), .RST(rst), .Q(c[798]) );
  DFF \sreg_reg[797]  ( .D(c[798]), .CLK(clk), .RST(rst), .Q(c[797]) );
  DFF \sreg_reg[796]  ( .D(c[797]), .CLK(clk), .RST(rst), .Q(c[796]) );
  DFF \sreg_reg[795]  ( .D(c[796]), .CLK(clk), .RST(rst), .Q(c[795]) );
  DFF \sreg_reg[794]  ( .D(c[795]), .CLK(clk), .RST(rst), .Q(c[794]) );
  DFF \sreg_reg[793]  ( .D(c[794]), .CLK(clk), .RST(rst), .Q(c[793]) );
  DFF \sreg_reg[792]  ( .D(c[793]), .CLK(clk), .RST(rst), .Q(c[792]) );
  DFF \sreg_reg[791]  ( .D(c[792]), .CLK(clk), .RST(rst), .Q(c[791]) );
  DFF \sreg_reg[790]  ( .D(c[791]), .CLK(clk), .RST(rst), .Q(c[790]) );
  DFF \sreg_reg[789]  ( .D(c[790]), .CLK(clk), .RST(rst), .Q(c[789]) );
  DFF \sreg_reg[788]  ( .D(c[789]), .CLK(clk), .RST(rst), .Q(c[788]) );
  DFF \sreg_reg[787]  ( .D(c[788]), .CLK(clk), .RST(rst), .Q(c[787]) );
  DFF \sreg_reg[786]  ( .D(c[787]), .CLK(clk), .RST(rst), .Q(c[786]) );
  DFF \sreg_reg[785]  ( .D(c[786]), .CLK(clk), .RST(rst), .Q(c[785]) );
  DFF \sreg_reg[784]  ( .D(c[785]), .CLK(clk), .RST(rst), .Q(c[784]) );
  DFF \sreg_reg[783]  ( .D(c[784]), .CLK(clk), .RST(rst), .Q(c[783]) );
  DFF \sreg_reg[782]  ( .D(c[783]), .CLK(clk), .RST(rst), .Q(c[782]) );
  DFF \sreg_reg[781]  ( .D(c[782]), .CLK(clk), .RST(rst), .Q(c[781]) );
  DFF \sreg_reg[780]  ( .D(c[781]), .CLK(clk), .RST(rst), .Q(c[780]) );
  DFF \sreg_reg[779]  ( .D(c[780]), .CLK(clk), .RST(rst), .Q(c[779]) );
  DFF \sreg_reg[778]  ( .D(c[779]), .CLK(clk), .RST(rst), .Q(c[778]) );
  DFF \sreg_reg[777]  ( .D(c[778]), .CLK(clk), .RST(rst), .Q(c[777]) );
  DFF \sreg_reg[776]  ( .D(c[777]), .CLK(clk), .RST(rst), .Q(c[776]) );
  DFF \sreg_reg[775]  ( .D(c[776]), .CLK(clk), .RST(rst), .Q(c[775]) );
  DFF \sreg_reg[774]  ( .D(c[775]), .CLK(clk), .RST(rst), .Q(c[774]) );
  DFF \sreg_reg[773]  ( .D(c[774]), .CLK(clk), .RST(rst), .Q(c[773]) );
  DFF \sreg_reg[772]  ( .D(c[773]), .CLK(clk), .RST(rst), .Q(c[772]) );
  DFF \sreg_reg[771]  ( .D(c[772]), .CLK(clk), .RST(rst), .Q(c[771]) );
  DFF \sreg_reg[770]  ( .D(c[771]), .CLK(clk), .RST(rst), .Q(c[770]) );
  DFF \sreg_reg[769]  ( .D(c[770]), .CLK(clk), .RST(rst), .Q(c[769]) );
  DFF \sreg_reg[768]  ( .D(c[769]), .CLK(clk), .RST(rst), .Q(c[768]) );
  DFF \sreg_reg[767]  ( .D(c[768]), .CLK(clk), .RST(rst), .Q(c[767]) );
  DFF \sreg_reg[766]  ( .D(c[767]), .CLK(clk), .RST(rst), .Q(c[766]) );
  DFF \sreg_reg[765]  ( .D(c[766]), .CLK(clk), .RST(rst), .Q(c[765]) );
  DFF \sreg_reg[764]  ( .D(c[765]), .CLK(clk), .RST(rst), .Q(c[764]) );
  DFF \sreg_reg[763]  ( .D(c[764]), .CLK(clk), .RST(rst), .Q(c[763]) );
  DFF \sreg_reg[762]  ( .D(c[763]), .CLK(clk), .RST(rst), .Q(c[762]) );
  DFF \sreg_reg[761]  ( .D(c[762]), .CLK(clk), .RST(rst), .Q(c[761]) );
  DFF \sreg_reg[760]  ( .D(c[761]), .CLK(clk), .RST(rst), .Q(c[760]) );
  DFF \sreg_reg[759]  ( .D(c[760]), .CLK(clk), .RST(rst), .Q(c[759]) );
  DFF \sreg_reg[758]  ( .D(c[759]), .CLK(clk), .RST(rst), .Q(c[758]) );
  DFF \sreg_reg[757]  ( .D(c[758]), .CLK(clk), .RST(rst), .Q(c[757]) );
  DFF \sreg_reg[756]  ( .D(c[757]), .CLK(clk), .RST(rst), .Q(c[756]) );
  DFF \sreg_reg[755]  ( .D(c[756]), .CLK(clk), .RST(rst), .Q(c[755]) );
  DFF \sreg_reg[754]  ( .D(c[755]), .CLK(clk), .RST(rst), .Q(c[754]) );
  DFF \sreg_reg[753]  ( .D(c[754]), .CLK(clk), .RST(rst), .Q(c[753]) );
  DFF \sreg_reg[752]  ( .D(c[753]), .CLK(clk), .RST(rst), .Q(c[752]) );
  DFF \sreg_reg[751]  ( .D(c[752]), .CLK(clk), .RST(rst), .Q(c[751]) );
  DFF \sreg_reg[750]  ( .D(c[751]), .CLK(clk), .RST(rst), .Q(c[750]) );
  DFF \sreg_reg[749]  ( .D(c[750]), .CLK(clk), .RST(rst), .Q(c[749]) );
  DFF \sreg_reg[748]  ( .D(c[749]), .CLK(clk), .RST(rst), .Q(c[748]) );
  DFF \sreg_reg[747]  ( .D(c[748]), .CLK(clk), .RST(rst), .Q(c[747]) );
  DFF \sreg_reg[746]  ( .D(c[747]), .CLK(clk), .RST(rst), .Q(c[746]) );
  DFF \sreg_reg[745]  ( .D(c[746]), .CLK(clk), .RST(rst), .Q(c[745]) );
  DFF \sreg_reg[744]  ( .D(c[745]), .CLK(clk), .RST(rst), .Q(c[744]) );
  DFF \sreg_reg[743]  ( .D(c[744]), .CLK(clk), .RST(rst), .Q(c[743]) );
  DFF \sreg_reg[742]  ( .D(c[743]), .CLK(clk), .RST(rst), .Q(c[742]) );
  DFF \sreg_reg[741]  ( .D(c[742]), .CLK(clk), .RST(rst), .Q(c[741]) );
  DFF \sreg_reg[740]  ( .D(c[741]), .CLK(clk), .RST(rst), .Q(c[740]) );
  DFF \sreg_reg[739]  ( .D(c[740]), .CLK(clk), .RST(rst), .Q(c[739]) );
  DFF \sreg_reg[738]  ( .D(c[739]), .CLK(clk), .RST(rst), .Q(c[738]) );
  DFF \sreg_reg[737]  ( .D(c[738]), .CLK(clk), .RST(rst), .Q(c[737]) );
  DFF \sreg_reg[736]  ( .D(c[737]), .CLK(clk), .RST(rst), .Q(c[736]) );
  DFF \sreg_reg[735]  ( .D(c[736]), .CLK(clk), .RST(rst), .Q(c[735]) );
  DFF \sreg_reg[734]  ( .D(c[735]), .CLK(clk), .RST(rst), .Q(c[734]) );
  DFF \sreg_reg[733]  ( .D(c[734]), .CLK(clk), .RST(rst), .Q(c[733]) );
  DFF \sreg_reg[732]  ( .D(c[733]), .CLK(clk), .RST(rst), .Q(c[732]) );
  DFF \sreg_reg[731]  ( .D(c[732]), .CLK(clk), .RST(rst), .Q(c[731]) );
  DFF \sreg_reg[730]  ( .D(c[731]), .CLK(clk), .RST(rst), .Q(c[730]) );
  DFF \sreg_reg[729]  ( .D(c[730]), .CLK(clk), .RST(rst), .Q(c[729]) );
  DFF \sreg_reg[728]  ( .D(c[729]), .CLK(clk), .RST(rst), .Q(c[728]) );
  DFF \sreg_reg[727]  ( .D(c[728]), .CLK(clk), .RST(rst), .Q(c[727]) );
  DFF \sreg_reg[726]  ( .D(c[727]), .CLK(clk), .RST(rst), .Q(c[726]) );
  DFF \sreg_reg[725]  ( .D(c[726]), .CLK(clk), .RST(rst), .Q(c[725]) );
  DFF \sreg_reg[724]  ( .D(c[725]), .CLK(clk), .RST(rst), .Q(c[724]) );
  DFF \sreg_reg[723]  ( .D(c[724]), .CLK(clk), .RST(rst), .Q(c[723]) );
  DFF \sreg_reg[722]  ( .D(c[723]), .CLK(clk), .RST(rst), .Q(c[722]) );
  DFF \sreg_reg[721]  ( .D(c[722]), .CLK(clk), .RST(rst), .Q(c[721]) );
  DFF \sreg_reg[720]  ( .D(c[721]), .CLK(clk), .RST(rst), .Q(c[720]) );
  DFF \sreg_reg[719]  ( .D(c[720]), .CLK(clk), .RST(rst), .Q(c[719]) );
  DFF \sreg_reg[718]  ( .D(c[719]), .CLK(clk), .RST(rst), .Q(c[718]) );
  DFF \sreg_reg[717]  ( .D(c[718]), .CLK(clk), .RST(rst), .Q(c[717]) );
  DFF \sreg_reg[716]  ( .D(c[717]), .CLK(clk), .RST(rst), .Q(c[716]) );
  DFF \sreg_reg[715]  ( .D(c[716]), .CLK(clk), .RST(rst), .Q(c[715]) );
  DFF \sreg_reg[714]  ( .D(c[715]), .CLK(clk), .RST(rst), .Q(c[714]) );
  DFF \sreg_reg[713]  ( .D(c[714]), .CLK(clk), .RST(rst), .Q(c[713]) );
  DFF \sreg_reg[712]  ( .D(c[713]), .CLK(clk), .RST(rst), .Q(c[712]) );
  DFF \sreg_reg[711]  ( .D(c[712]), .CLK(clk), .RST(rst), .Q(c[711]) );
  DFF \sreg_reg[710]  ( .D(c[711]), .CLK(clk), .RST(rst), .Q(c[710]) );
  DFF \sreg_reg[709]  ( .D(c[710]), .CLK(clk), .RST(rst), .Q(c[709]) );
  DFF \sreg_reg[708]  ( .D(c[709]), .CLK(clk), .RST(rst), .Q(c[708]) );
  DFF \sreg_reg[707]  ( .D(c[708]), .CLK(clk), .RST(rst), .Q(c[707]) );
  DFF \sreg_reg[706]  ( .D(c[707]), .CLK(clk), .RST(rst), .Q(c[706]) );
  DFF \sreg_reg[705]  ( .D(c[706]), .CLK(clk), .RST(rst), .Q(c[705]) );
  DFF \sreg_reg[704]  ( .D(c[705]), .CLK(clk), .RST(rst), .Q(c[704]) );
  DFF \sreg_reg[703]  ( .D(c[704]), .CLK(clk), .RST(rst), .Q(c[703]) );
  DFF \sreg_reg[702]  ( .D(c[703]), .CLK(clk), .RST(rst), .Q(c[702]) );
  DFF \sreg_reg[701]  ( .D(c[702]), .CLK(clk), .RST(rst), .Q(c[701]) );
  DFF \sreg_reg[700]  ( .D(c[701]), .CLK(clk), .RST(rst), .Q(c[700]) );
  DFF \sreg_reg[699]  ( .D(c[700]), .CLK(clk), .RST(rst), .Q(c[699]) );
  DFF \sreg_reg[698]  ( .D(c[699]), .CLK(clk), .RST(rst), .Q(c[698]) );
  DFF \sreg_reg[697]  ( .D(c[698]), .CLK(clk), .RST(rst), .Q(c[697]) );
  DFF \sreg_reg[696]  ( .D(c[697]), .CLK(clk), .RST(rst), .Q(c[696]) );
  DFF \sreg_reg[695]  ( .D(c[696]), .CLK(clk), .RST(rst), .Q(c[695]) );
  DFF \sreg_reg[694]  ( .D(c[695]), .CLK(clk), .RST(rst), .Q(c[694]) );
  DFF \sreg_reg[693]  ( .D(c[694]), .CLK(clk), .RST(rst), .Q(c[693]) );
  DFF \sreg_reg[692]  ( .D(c[693]), .CLK(clk), .RST(rst), .Q(c[692]) );
  DFF \sreg_reg[691]  ( .D(c[692]), .CLK(clk), .RST(rst), .Q(c[691]) );
  DFF \sreg_reg[690]  ( .D(c[691]), .CLK(clk), .RST(rst), .Q(c[690]) );
  DFF \sreg_reg[689]  ( .D(c[690]), .CLK(clk), .RST(rst), .Q(c[689]) );
  DFF \sreg_reg[688]  ( .D(c[689]), .CLK(clk), .RST(rst), .Q(c[688]) );
  DFF \sreg_reg[687]  ( .D(c[688]), .CLK(clk), .RST(rst), .Q(c[687]) );
  DFF \sreg_reg[686]  ( .D(c[687]), .CLK(clk), .RST(rst), .Q(c[686]) );
  DFF \sreg_reg[685]  ( .D(c[686]), .CLK(clk), .RST(rst), .Q(c[685]) );
  DFF \sreg_reg[684]  ( .D(c[685]), .CLK(clk), .RST(rst), .Q(c[684]) );
  DFF \sreg_reg[683]  ( .D(c[684]), .CLK(clk), .RST(rst), .Q(c[683]) );
  DFF \sreg_reg[682]  ( .D(c[683]), .CLK(clk), .RST(rst), .Q(c[682]) );
  DFF \sreg_reg[681]  ( .D(c[682]), .CLK(clk), .RST(rst), .Q(c[681]) );
  DFF \sreg_reg[680]  ( .D(c[681]), .CLK(clk), .RST(rst), .Q(c[680]) );
  DFF \sreg_reg[679]  ( .D(c[680]), .CLK(clk), .RST(rst), .Q(c[679]) );
  DFF \sreg_reg[678]  ( .D(c[679]), .CLK(clk), .RST(rst), .Q(c[678]) );
  DFF \sreg_reg[677]  ( .D(c[678]), .CLK(clk), .RST(rst), .Q(c[677]) );
  DFF \sreg_reg[676]  ( .D(c[677]), .CLK(clk), .RST(rst), .Q(c[676]) );
  DFF \sreg_reg[675]  ( .D(c[676]), .CLK(clk), .RST(rst), .Q(c[675]) );
  DFF \sreg_reg[674]  ( .D(c[675]), .CLK(clk), .RST(rst), .Q(c[674]) );
  DFF \sreg_reg[673]  ( .D(c[674]), .CLK(clk), .RST(rst), .Q(c[673]) );
  DFF \sreg_reg[672]  ( .D(c[673]), .CLK(clk), .RST(rst), .Q(c[672]) );
  DFF \sreg_reg[671]  ( .D(c[672]), .CLK(clk), .RST(rst), .Q(c[671]) );
  DFF \sreg_reg[670]  ( .D(c[671]), .CLK(clk), .RST(rst), .Q(c[670]) );
  DFF \sreg_reg[669]  ( .D(c[670]), .CLK(clk), .RST(rst), .Q(c[669]) );
  DFF \sreg_reg[668]  ( .D(c[669]), .CLK(clk), .RST(rst), .Q(c[668]) );
  DFF \sreg_reg[667]  ( .D(c[668]), .CLK(clk), .RST(rst), .Q(c[667]) );
  DFF \sreg_reg[666]  ( .D(c[667]), .CLK(clk), .RST(rst), .Q(c[666]) );
  DFF \sreg_reg[665]  ( .D(c[666]), .CLK(clk), .RST(rst), .Q(c[665]) );
  DFF \sreg_reg[664]  ( .D(c[665]), .CLK(clk), .RST(rst), .Q(c[664]) );
  DFF \sreg_reg[663]  ( .D(c[664]), .CLK(clk), .RST(rst), .Q(c[663]) );
  DFF \sreg_reg[662]  ( .D(c[663]), .CLK(clk), .RST(rst), .Q(c[662]) );
  DFF \sreg_reg[661]  ( .D(c[662]), .CLK(clk), .RST(rst), .Q(c[661]) );
  DFF \sreg_reg[660]  ( .D(c[661]), .CLK(clk), .RST(rst), .Q(c[660]) );
  DFF \sreg_reg[659]  ( .D(c[660]), .CLK(clk), .RST(rst), .Q(c[659]) );
  DFF \sreg_reg[658]  ( .D(c[659]), .CLK(clk), .RST(rst), .Q(c[658]) );
  DFF \sreg_reg[657]  ( .D(c[658]), .CLK(clk), .RST(rst), .Q(c[657]) );
  DFF \sreg_reg[656]  ( .D(c[657]), .CLK(clk), .RST(rst), .Q(c[656]) );
  DFF \sreg_reg[655]  ( .D(c[656]), .CLK(clk), .RST(rst), .Q(c[655]) );
  DFF \sreg_reg[654]  ( .D(c[655]), .CLK(clk), .RST(rst), .Q(c[654]) );
  DFF \sreg_reg[653]  ( .D(c[654]), .CLK(clk), .RST(rst), .Q(c[653]) );
  DFF \sreg_reg[652]  ( .D(c[653]), .CLK(clk), .RST(rst), .Q(c[652]) );
  DFF \sreg_reg[651]  ( .D(c[652]), .CLK(clk), .RST(rst), .Q(c[651]) );
  DFF \sreg_reg[650]  ( .D(c[651]), .CLK(clk), .RST(rst), .Q(c[650]) );
  DFF \sreg_reg[649]  ( .D(c[650]), .CLK(clk), .RST(rst), .Q(c[649]) );
  DFF \sreg_reg[648]  ( .D(c[649]), .CLK(clk), .RST(rst), .Q(c[648]) );
  DFF \sreg_reg[647]  ( .D(c[648]), .CLK(clk), .RST(rst), .Q(c[647]) );
  DFF \sreg_reg[646]  ( .D(c[647]), .CLK(clk), .RST(rst), .Q(c[646]) );
  DFF \sreg_reg[645]  ( .D(c[646]), .CLK(clk), .RST(rst), .Q(c[645]) );
  DFF \sreg_reg[644]  ( .D(c[645]), .CLK(clk), .RST(rst), .Q(c[644]) );
  DFF \sreg_reg[643]  ( .D(c[644]), .CLK(clk), .RST(rst), .Q(c[643]) );
  DFF \sreg_reg[642]  ( .D(c[643]), .CLK(clk), .RST(rst), .Q(c[642]) );
  DFF \sreg_reg[641]  ( .D(c[642]), .CLK(clk), .RST(rst), .Q(c[641]) );
  DFF \sreg_reg[640]  ( .D(c[641]), .CLK(clk), .RST(rst), .Q(c[640]) );
  DFF \sreg_reg[639]  ( .D(c[640]), .CLK(clk), .RST(rst), .Q(c[639]) );
  DFF \sreg_reg[638]  ( .D(c[639]), .CLK(clk), .RST(rst), .Q(c[638]) );
  DFF \sreg_reg[637]  ( .D(c[638]), .CLK(clk), .RST(rst), .Q(c[637]) );
  DFF \sreg_reg[636]  ( .D(c[637]), .CLK(clk), .RST(rst), .Q(c[636]) );
  DFF \sreg_reg[635]  ( .D(c[636]), .CLK(clk), .RST(rst), .Q(c[635]) );
  DFF \sreg_reg[634]  ( .D(c[635]), .CLK(clk), .RST(rst), .Q(c[634]) );
  DFF \sreg_reg[633]  ( .D(c[634]), .CLK(clk), .RST(rst), .Q(c[633]) );
  DFF \sreg_reg[632]  ( .D(c[633]), .CLK(clk), .RST(rst), .Q(c[632]) );
  DFF \sreg_reg[631]  ( .D(c[632]), .CLK(clk), .RST(rst), .Q(c[631]) );
  DFF \sreg_reg[630]  ( .D(c[631]), .CLK(clk), .RST(rst), .Q(c[630]) );
  DFF \sreg_reg[629]  ( .D(c[630]), .CLK(clk), .RST(rst), .Q(c[629]) );
  DFF \sreg_reg[628]  ( .D(c[629]), .CLK(clk), .RST(rst), .Q(c[628]) );
  DFF \sreg_reg[627]  ( .D(c[628]), .CLK(clk), .RST(rst), .Q(c[627]) );
  DFF \sreg_reg[626]  ( .D(c[627]), .CLK(clk), .RST(rst), .Q(c[626]) );
  DFF \sreg_reg[625]  ( .D(c[626]), .CLK(clk), .RST(rst), .Q(c[625]) );
  DFF \sreg_reg[624]  ( .D(c[625]), .CLK(clk), .RST(rst), .Q(c[624]) );
  DFF \sreg_reg[623]  ( .D(c[624]), .CLK(clk), .RST(rst), .Q(c[623]) );
  DFF \sreg_reg[622]  ( .D(c[623]), .CLK(clk), .RST(rst), .Q(c[622]) );
  DFF \sreg_reg[621]  ( .D(c[622]), .CLK(clk), .RST(rst), .Q(c[621]) );
  DFF \sreg_reg[620]  ( .D(c[621]), .CLK(clk), .RST(rst), .Q(c[620]) );
  DFF \sreg_reg[619]  ( .D(c[620]), .CLK(clk), .RST(rst), .Q(c[619]) );
  DFF \sreg_reg[618]  ( .D(c[619]), .CLK(clk), .RST(rst), .Q(c[618]) );
  DFF \sreg_reg[617]  ( .D(c[618]), .CLK(clk), .RST(rst), .Q(c[617]) );
  DFF \sreg_reg[616]  ( .D(c[617]), .CLK(clk), .RST(rst), .Q(c[616]) );
  DFF \sreg_reg[615]  ( .D(c[616]), .CLK(clk), .RST(rst), .Q(c[615]) );
  DFF \sreg_reg[614]  ( .D(c[615]), .CLK(clk), .RST(rst), .Q(c[614]) );
  DFF \sreg_reg[613]  ( .D(c[614]), .CLK(clk), .RST(rst), .Q(c[613]) );
  DFF \sreg_reg[612]  ( .D(c[613]), .CLK(clk), .RST(rst), .Q(c[612]) );
  DFF \sreg_reg[611]  ( .D(c[612]), .CLK(clk), .RST(rst), .Q(c[611]) );
  DFF \sreg_reg[610]  ( .D(c[611]), .CLK(clk), .RST(rst), .Q(c[610]) );
  DFF \sreg_reg[609]  ( .D(c[610]), .CLK(clk), .RST(rst), .Q(c[609]) );
  DFF \sreg_reg[608]  ( .D(c[609]), .CLK(clk), .RST(rst), .Q(c[608]) );
  DFF \sreg_reg[607]  ( .D(c[608]), .CLK(clk), .RST(rst), .Q(c[607]) );
  DFF \sreg_reg[606]  ( .D(c[607]), .CLK(clk), .RST(rst), .Q(c[606]) );
  DFF \sreg_reg[605]  ( .D(c[606]), .CLK(clk), .RST(rst), .Q(c[605]) );
  DFF \sreg_reg[604]  ( .D(c[605]), .CLK(clk), .RST(rst), .Q(c[604]) );
  DFF \sreg_reg[603]  ( .D(c[604]), .CLK(clk), .RST(rst), .Q(c[603]) );
  DFF \sreg_reg[602]  ( .D(c[603]), .CLK(clk), .RST(rst), .Q(c[602]) );
  DFF \sreg_reg[601]  ( .D(c[602]), .CLK(clk), .RST(rst), .Q(c[601]) );
  DFF \sreg_reg[600]  ( .D(c[601]), .CLK(clk), .RST(rst), .Q(c[600]) );
  DFF \sreg_reg[599]  ( .D(c[600]), .CLK(clk), .RST(rst), .Q(c[599]) );
  DFF \sreg_reg[598]  ( .D(c[599]), .CLK(clk), .RST(rst), .Q(c[598]) );
  DFF \sreg_reg[597]  ( .D(c[598]), .CLK(clk), .RST(rst), .Q(c[597]) );
  DFF \sreg_reg[596]  ( .D(c[597]), .CLK(clk), .RST(rst), .Q(c[596]) );
  DFF \sreg_reg[595]  ( .D(c[596]), .CLK(clk), .RST(rst), .Q(c[595]) );
  DFF \sreg_reg[594]  ( .D(c[595]), .CLK(clk), .RST(rst), .Q(c[594]) );
  DFF \sreg_reg[593]  ( .D(c[594]), .CLK(clk), .RST(rst), .Q(c[593]) );
  DFF \sreg_reg[592]  ( .D(c[593]), .CLK(clk), .RST(rst), .Q(c[592]) );
  DFF \sreg_reg[591]  ( .D(c[592]), .CLK(clk), .RST(rst), .Q(c[591]) );
  DFF \sreg_reg[590]  ( .D(c[591]), .CLK(clk), .RST(rst), .Q(c[590]) );
  DFF \sreg_reg[589]  ( .D(c[590]), .CLK(clk), .RST(rst), .Q(c[589]) );
  DFF \sreg_reg[588]  ( .D(c[589]), .CLK(clk), .RST(rst), .Q(c[588]) );
  DFF \sreg_reg[587]  ( .D(c[588]), .CLK(clk), .RST(rst), .Q(c[587]) );
  DFF \sreg_reg[586]  ( .D(c[587]), .CLK(clk), .RST(rst), .Q(c[586]) );
  DFF \sreg_reg[585]  ( .D(c[586]), .CLK(clk), .RST(rst), .Q(c[585]) );
  DFF \sreg_reg[584]  ( .D(c[585]), .CLK(clk), .RST(rst), .Q(c[584]) );
  DFF \sreg_reg[583]  ( .D(c[584]), .CLK(clk), .RST(rst), .Q(c[583]) );
  DFF \sreg_reg[582]  ( .D(c[583]), .CLK(clk), .RST(rst), .Q(c[582]) );
  DFF \sreg_reg[581]  ( .D(c[582]), .CLK(clk), .RST(rst), .Q(c[581]) );
  DFF \sreg_reg[580]  ( .D(c[581]), .CLK(clk), .RST(rst), .Q(c[580]) );
  DFF \sreg_reg[579]  ( .D(c[580]), .CLK(clk), .RST(rst), .Q(c[579]) );
  DFF \sreg_reg[578]  ( .D(c[579]), .CLK(clk), .RST(rst), .Q(c[578]) );
  DFF \sreg_reg[577]  ( .D(c[578]), .CLK(clk), .RST(rst), .Q(c[577]) );
  DFF \sreg_reg[576]  ( .D(c[577]), .CLK(clk), .RST(rst), .Q(c[576]) );
  DFF \sreg_reg[575]  ( .D(c[576]), .CLK(clk), .RST(rst), .Q(c[575]) );
  DFF \sreg_reg[574]  ( .D(c[575]), .CLK(clk), .RST(rst), .Q(c[574]) );
  DFF \sreg_reg[573]  ( .D(c[574]), .CLK(clk), .RST(rst), .Q(c[573]) );
  DFF \sreg_reg[572]  ( .D(c[573]), .CLK(clk), .RST(rst), .Q(c[572]) );
  DFF \sreg_reg[571]  ( .D(c[572]), .CLK(clk), .RST(rst), .Q(c[571]) );
  DFF \sreg_reg[570]  ( .D(c[571]), .CLK(clk), .RST(rst), .Q(c[570]) );
  DFF \sreg_reg[569]  ( .D(c[570]), .CLK(clk), .RST(rst), .Q(c[569]) );
  DFF \sreg_reg[568]  ( .D(c[569]), .CLK(clk), .RST(rst), .Q(c[568]) );
  DFF \sreg_reg[567]  ( .D(c[568]), .CLK(clk), .RST(rst), .Q(c[567]) );
  DFF \sreg_reg[566]  ( .D(c[567]), .CLK(clk), .RST(rst), .Q(c[566]) );
  DFF \sreg_reg[565]  ( .D(c[566]), .CLK(clk), .RST(rst), .Q(c[565]) );
  DFF \sreg_reg[564]  ( .D(c[565]), .CLK(clk), .RST(rst), .Q(c[564]) );
  DFF \sreg_reg[563]  ( .D(c[564]), .CLK(clk), .RST(rst), .Q(c[563]) );
  DFF \sreg_reg[562]  ( .D(c[563]), .CLK(clk), .RST(rst), .Q(c[562]) );
  DFF \sreg_reg[561]  ( .D(c[562]), .CLK(clk), .RST(rst), .Q(c[561]) );
  DFF \sreg_reg[560]  ( .D(c[561]), .CLK(clk), .RST(rst), .Q(c[560]) );
  DFF \sreg_reg[559]  ( .D(c[560]), .CLK(clk), .RST(rst), .Q(c[559]) );
  DFF \sreg_reg[558]  ( .D(c[559]), .CLK(clk), .RST(rst), .Q(c[558]) );
  DFF \sreg_reg[557]  ( .D(c[558]), .CLK(clk), .RST(rst), .Q(c[557]) );
  DFF \sreg_reg[556]  ( .D(c[557]), .CLK(clk), .RST(rst), .Q(c[556]) );
  DFF \sreg_reg[555]  ( .D(c[556]), .CLK(clk), .RST(rst), .Q(c[555]) );
  DFF \sreg_reg[554]  ( .D(c[555]), .CLK(clk), .RST(rst), .Q(c[554]) );
  DFF \sreg_reg[553]  ( .D(c[554]), .CLK(clk), .RST(rst), .Q(c[553]) );
  DFF \sreg_reg[552]  ( .D(c[553]), .CLK(clk), .RST(rst), .Q(c[552]) );
  DFF \sreg_reg[551]  ( .D(c[552]), .CLK(clk), .RST(rst), .Q(c[551]) );
  DFF \sreg_reg[550]  ( .D(c[551]), .CLK(clk), .RST(rst), .Q(c[550]) );
  DFF \sreg_reg[549]  ( .D(c[550]), .CLK(clk), .RST(rst), .Q(c[549]) );
  DFF \sreg_reg[548]  ( .D(c[549]), .CLK(clk), .RST(rst), .Q(c[548]) );
  DFF \sreg_reg[547]  ( .D(c[548]), .CLK(clk), .RST(rst), .Q(c[547]) );
  DFF \sreg_reg[546]  ( .D(c[547]), .CLK(clk), .RST(rst), .Q(c[546]) );
  DFF \sreg_reg[545]  ( .D(c[546]), .CLK(clk), .RST(rst), .Q(c[545]) );
  DFF \sreg_reg[544]  ( .D(c[545]), .CLK(clk), .RST(rst), .Q(c[544]) );
  DFF \sreg_reg[543]  ( .D(c[544]), .CLK(clk), .RST(rst), .Q(c[543]) );
  DFF \sreg_reg[542]  ( .D(c[543]), .CLK(clk), .RST(rst), .Q(c[542]) );
  DFF \sreg_reg[541]  ( .D(c[542]), .CLK(clk), .RST(rst), .Q(c[541]) );
  DFF \sreg_reg[540]  ( .D(c[541]), .CLK(clk), .RST(rst), .Q(c[540]) );
  DFF \sreg_reg[539]  ( .D(c[540]), .CLK(clk), .RST(rst), .Q(c[539]) );
  DFF \sreg_reg[538]  ( .D(c[539]), .CLK(clk), .RST(rst), .Q(c[538]) );
  DFF \sreg_reg[537]  ( .D(c[538]), .CLK(clk), .RST(rst), .Q(c[537]) );
  DFF \sreg_reg[536]  ( .D(c[537]), .CLK(clk), .RST(rst), .Q(c[536]) );
  DFF \sreg_reg[535]  ( .D(c[536]), .CLK(clk), .RST(rst), .Q(c[535]) );
  DFF \sreg_reg[534]  ( .D(c[535]), .CLK(clk), .RST(rst), .Q(c[534]) );
  DFF \sreg_reg[533]  ( .D(c[534]), .CLK(clk), .RST(rst), .Q(c[533]) );
  DFF \sreg_reg[532]  ( .D(c[533]), .CLK(clk), .RST(rst), .Q(c[532]) );
  DFF \sreg_reg[531]  ( .D(c[532]), .CLK(clk), .RST(rst), .Q(c[531]) );
  DFF \sreg_reg[530]  ( .D(c[531]), .CLK(clk), .RST(rst), .Q(c[530]) );
  DFF \sreg_reg[529]  ( .D(c[530]), .CLK(clk), .RST(rst), .Q(c[529]) );
  DFF \sreg_reg[528]  ( .D(c[529]), .CLK(clk), .RST(rst), .Q(c[528]) );
  DFF \sreg_reg[527]  ( .D(c[528]), .CLK(clk), .RST(rst), .Q(c[527]) );
  DFF \sreg_reg[526]  ( .D(c[527]), .CLK(clk), .RST(rst), .Q(c[526]) );
  DFF \sreg_reg[525]  ( .D(c[526]), .CLK(clk), .RST(rst), .Q(c[525]) );
  DFF \sreg_reg[524]  ( .D(c[525]), .CLK(clk), .RST(rst), .Q(c[524]) );
  DFF \sreg_reg[523]  ( .D(c[524]), .CLK(clk), .RST(rst), .Q(c[523]) );
  DFF \sreg_reg[522]  ( .D(c[523]), .CLK(clk), .RST(rst), .Q(c[522]) );
  DFF \sreg_reg[521]  ( .D(c[522]), .CLK(clk), .RST(rst), .Q(c[521]) );
  DFF \sreg_reg[520]  ( .D(c[521]), .CLK(clk), .RST(rst), .Q(c[520]) );
  DFF \sreg_reg[519]  ( .D(c[520]), .CLK(clk), .RST(rst), .Q(c[519]) );
  DFF \sreg_reg[518]  ( .D(c[519]), .CLK(clk), .RST(rst), .Q(c[518]) );
  DFF \sreg_reg[517]  ( .D(c[518]), .CLK(clk), .RST(rst), .Q(c[517]) );
  DFF \sreg_reg[516]  ( .D(c[517]), .CLK(clk), .RST(rst), .Q(c[516]) );
  DFF \sreg_reg[515]  ( .D(c[516]), .CLK(clk), .RST(rst), .Q(c[515]) );
  DFF \sreg_reg[514]  ( .D(c[515]), .CLK(clk), .RST(rst), .Q(c[514]) );
  DFF \sreg_reg[513]  ( .D(c[514]), .CLK(clk), .RST(rst), .Q(c[513]) );
  DFF \sreg_reg[512]  ( .D(c[513]), .CLK(clk), .RST(rst), .Q(c[512]) );
  DFF \sreg_reg[511]  ( .D(c[512]), .CLK(clk), .RST(rst), .Q(c[511]) );
  DFF \sreg_reg[510]  ( .D(c[511]), .CLK(clk), .RST(rst), .Q(c[510]) );
  DFF \sreg_reg[509]  ( .D(c[510]), .CLK(clk), .RST(rst), .Q(c[509]) );
  DFF \sreg_reg[508]  ( .D(c[509]), .CLK(clk), .RST(rst), .Q(c[508]) );
  DFF \sreg_reg[507]  ( .D(c[508]), .CLK(clk), .RST(rst), .Q(c[507]) );
  DFF \sreg_reg[506]  ( .D(c[507]), .CLK(clk), .RST(rst), .Q(c[506]) );
  DFF \sreg_reg[505]  ( .D(c[506]), .CLK(clk), .RST(rst), .Q(c[505]) );
  DFF \sreg_reg[504]  ( .D(c[505]), .CLK(clk), .RST(rst), .Q(c[504]) );
  DFF \sreg_reg[503]  ( .D(c[504]), .CLK(clk), .RST(rst), .Q(c[503]) );
  DFF \sreg_reg[502]  ( .D(c[503]), .CLK(clk), .RST(rst), .Q(c[502]) );
  DFF \sreg_reg[501]  ( .D(c[502]), .CLK(clk), .RST(rst), .Q(c[501]) );
  DFF \sreg_reg[500]  ( .D(c[501]), .CLK(clk), .RST(rst), .Q(c[500]) );
  DFF \sreg_reg[499]  ( .D(c[500]), .CLK(clk), .RST(rst), .Q(c[499]) );
  DFF \sreg_reg[498]  ( .D(c[499]), .CLK(clk), .RST(rst), .Q(c[498]) );
  DFF \sreg_reg[497]  ( .D(c[498]), .CLK(clk), .RST(rst), .Q(c[497]) );
  DFF \sreg_reg[496]  ( .D(c[497]), .CLK(clk), .RST(rst), .Q(c[496]) );
  DFF \sreg_reg[495]  ( .D(c[496]), .CLK(clk), .RST(rst), .Q(c[495]) );
  DFF \sreg_reg[494]  ( .D(c[495]), .CLK(clk), .RST(rst), .Q(c[494]) );
  DFF \sreg_reg[493]  ( .D(c[494]), .CLK(clk), .RST(rst), .Q(c[493]) );
  DFF \sreg_reg[492]  ( .D(c[493]), .CLK(clk), .RST(rst), .Q(c[492]) );
  DFF \sreg_reg[491]  ( .D(c[492]), .CLK(clk), .RST(rst), .Q(c[491]) );
  DFF \sreg_reg[490]  ( .D(c[491]), .CLK(clk), .RST(rst), .Q(c[490]) );
  DFF \sreg_reg[489]  ( .D(c[490]), .CLK(clk), .RST(rst), .Q(c[489]) );
  DFF \sreg_reg[488]  ( .D(c[489]), .CLK(clk), .RST(rst), .Q(c[488]) );
  DFF \sreg_reg[487]  ( .D(c[488]), .CLK(clk), .RST(rst), .Q(c[487]) );
  DFF \sreg_reg[486]  ( .D(c[487]), .CLK(clk), .RST(rst), .Q(c[486]) );
  DFF \sreg_reg[485]  ( .D(c[486]), .CLK(clk), .RST(rst), .Q(c[485]) );
  DFF \sreg_reg[484]  ( .D(c[485]), .CLK(clk), .RST(rst), .Q(c[484]) );
  DFF \sreg_reg[483]  ( .D(c[484]), .CLK(clk), .RST(rst), .Q(c[483]) );
  DFF \sreg_reg[482]  ( .D(c[483]), .CLK(clk), .RST(rst), .Q(c[482]) );
  DFF \sreg_reg[481]  ( .D(c[482]), .CLK(clk), .RST(rst), .Q(c[481]) );
  DFF \sreg_reg[480]  ( .D(c[481]), .CLK(clk), .RST(rst), .Q(c[480]) );
  DFF \sreg_reg[479]  ( .D(c[480]), .CLK(clk), .RST(rst), .Q(c[479]) );
  DFF \sreg_reg[478]  ( .D(c[479]), .CLK(clk), .RST(rst), .Q(c[478]) );
  DFF \sreg_reg[477]  ( .D(c[478]), .CLK(clk), .RST(rst), .Q(c[477]) );
  DFF \sreg_reg[476]  ( .D(c[477]), .CLK(clk), .RST(rst), .Q(c[476]) );
  DFF \sreg_reg[475]  ( .D(c[476]), .CLK(clk), .RST(rst), .Q(c[475]) );
  DFF \sreg_reg[474]  ( .D(c[475]), .CLK(clk), .RST(rst), .Q(c[474]) );
  DFF \sreg_reg[473]  ( .D(c[474]), .CLK(clk), .RST(rst), .Q(c[473]) );
  DFF \sreg_reg[472]  ( .D(c[473]), .CLK(clk), .RST(rst), .Q(c[472]) );
  DFF \sreg_reg[471]  ( .D(c[472]), .CLK(clk), .RST(rst), .Q(c[471]) );
  DFF \sreg_reg[470]  ( .D(c[471]), .CLK(clk), .RST(rst), .Q(c[470]) );
  DFF \sreg_reg[469]  ( .D(c[470]), .CLK(clk), .RST(rst), .Q(c[469]) );
  DFF \sreg_reg[468]  ( .D(c[469]), .CLK(clk), .RST(rst), .Q(c[468]) );
  DFF \sreg_reg[467]  ( .D(c[468]), .CLK(clk), .RST(rst), .Q(c[467]) );
  DFF \sreg_reg[466]  ( .D(c[467]), .CLK(clk), .RST(rst), .Q(c[466]) );
  DFF \sreg_reg[465]  ( .D(c[466]), .CLK(clk), .RST(rst), .Q(c[465]) );
  DFF \sreg_reg[464]  ( .D(c[465]), .CLK(clk), .RST(rst), .Q(c[464]) );
  DFF \sreg_reg[463]  ( .D(c[464]), .CLK(clk), .RST(rst), .Q(c[463]) );
  DFF \sreg_reg[462]  ( .D(c[463]), .CLK(clk), .RST(rst), .Q(c[462]) );
  DFF \sreg_reg[461]  ( .D(c[462]), .CLK(clk), .RST(rst), .Q(c[461]) );
  DFF \sreg_reg[460]  ( .D(c[461]), .CLK(clk), .RST(rst), .Q(c[460]) );
  DFF \sreg_reg[459]  ( .D(c[460]), .CLK(clk), .RST(rst), .Q(c[459]) );
  DFF \sreg_reg[458]  ( .D(c[459]), .CLK(clk), .RST(rst), .Q(c[458]) );
  DFF \sreg_reg[457]  ( .D(c[458]), .CLK(clk), .RST(rst), .Q(c[457]) );
  DFF \sreg_reg[456]  ( .D(c[457]), .CLK(clk), .RST(rst), .Q(c[456]) );
  DFF \sreg_reg[455]  ( .D(c[456]), .CLK(clk), .RST(rst), .Q(c[455]) );
  DFF \sreg_reg[454]  ( .D(c[455]), .CLK(clk), .RST(rst), .Q(c[454]) );
  DFF \sreg_reg[453]  ( .D(c[454]), .CLK(clk), .RST(rst), .Q(c[453]) );
  DFF \sreg_reg[452]  ( .D(c[453]), .CLK(clk), .RST(rst), .Q(c[452]) );
  DFF \sreg_reg[451]  ( .D(c[452]), .CLK(clk), .RST(rst), .Q(c[451]) );
  DFF \sreg_reg[450]  ( .D(c[451]), .CLK(clk), .RST(rst), .Q(c[450]) );
  DFF \sreg_reg[449]  ( .D(c[450]), .CLK(clk), .RST(rst), .Q(c[449]) );
  DFF \sreg_reg[448]  ( .D(c[449]), .CLK(clk), .RST(rst), .Q(c[448]) );
  DFF \sreg_reg[447]  ( .D(c[448]), .CLK(clk), .RST(rst), .Q(c[447]) );
  DFF \sreg_reg[446]  ( .D(c[447]), .CLK(clk), .RST(rst), .Q(c[446]) );
  DFF \sreg_reg[445]  ( .D(c[446]), .CLK(clk), .RST(rst), .Q(c[445]) );
  DFF \sreg_reg[444]  ( .D(c[445]), .CLK(clk), .RST(rst), .Q(c[444]) );
  DFF \sreg_reg[443]  ( .D(c[444]), .CLK(clk), .RST(rst), .Q(c[443]) );
  DFF \sreg_reg[442]  ( .D(c[443]), .CLK(clk), .RST(rst), .Q(c[442]) );
  DFF \sreg_reg[441]  ( .D(c[442]), .CLK(clk), .RST(rst), .Q(c[441]) );
  DFF \sreg_reg[440]  ( .D(c[441]), .CLK(clk), .RST(rst), .Q(c[440]) );
  DFF \sreg_reg[439]  ( .D(c[440]), .CLK(clk), .RST(rst), .Q(c[439]) );
  DFF \sreg_reg[438]  ( .D(c[439]), .CLK(clk), .RST(rst), .Q(c[438]) );
  DFF \sreg_reg[437]  ( .D(c[438]), .CLK(clk), .RST(rst), .Q(c[437]) );
  DFF \sreg_reg[436]  ( .D(c[437]), .CLK(clk), .RST(rst), .Q(c[436]) );
  DFF \sreg_reg[435]  ( .D(c[436]), .CLK(clk), .RST(rst), .Q(c[435]) );
  DFF \sreg_reg[434]  ( .D(c[435]), .CLK(clk), .RST(rst), .Q(c[434]) );
  DFF \sreg_reg[433]  ( .D(c[434]), .CLK(clk), .RST(rst), .Q(c[433]) );
  DFF \sreg_reg[432]  ( .D(c[433]), .CLK(clk), .RST(rst), .Q(c[432]) );
  DFF \sreg_reg[431]  ( .D(c[432]), .CLK(clk), .RST(rst), .Q(c[431]) );
  DFF \sreg_reg[430]  ( .D(c[431]), .CLK(clk), .RST(rst), .Q(c[430]) );
  DFF \sreg_reg[429]  ( .D(c[430]), .CLK(clk), .RST(rst), .Q(c[429]) );
  DFF \sreg_reg[428]  ( .D(c[429]), .CLK(clk), .RST(rst), .Q(c[428]) );
  DFF \sreg_reg[427]  ( .D(c[428]), .CLK(clk), .RST(rst), .Q(c[427]) );
  DFF \sreg_reg[426]  ( .D(c[427]), .CLK(clk), .RST(rst), .Q(c[426]) );
  DFF \sreg_reg[425]  ( .D(c[426]), .CLK(clk), .RST(rst), .Q(c[425]) );
  DFF \sreg_reg[424]  ( .D(c[425]), .CLK(clk), .RST(rst), .Q(c[424]) );
  DFF \sreg_reg[423]  ( .D(c[424]), .CLK(clk), .RST(rst), .Q(c[423]) );
  DFF \sreg_reg[422]  ( .D(c[423]), .CLK(clk), .RST(rst), .Q(c[422]) );
  DFF \sreg_reg[421]  ( .D(c[422]), .CLK(clk), .RST(rst), .Q(c[421]) );
  DFF \sreg_reg[420]  ( .D(c[421]), .CLK(clk), .RST(rst), .Q(c[420]) );
  DFF \sreg_reg[419]  ( .D(c[420]), .CLK(clk), .RST(rst), .Q(c[419]) );
  DFF \sreg_reg[418]  ( .D(c[419]), .CLK(clk), .RST(rst), .Q(c[418]) );
  DFF \sreg_reg[417]  ( .D(c[418]), .CLK(clk), .RST(rst), .Q(c[417]) );
  DFF \sreg_reg[416]  ( .D(c[417]), .CLK(clk), .RST(rst), .Q(c[416]) );
  DFF \sreg_reg[415]  ( .D(c[416]), .CLK(clk), .RST(rst), .Q(c[415]) );
  DFF \sreg_reg[414]  ( .D(c[415]), .CLK(clk), .RST(rst), .Q(c[414]) );
  DFF \sreg_reg[413]  ( .D(c[414]), .CLK(clk), .RST(rst), .Q(c[413]) );
  DFF \sreg_reg[412]  ( .D(c[413]), .CLK(clk), .RST(rst), .Q(c[412]) );
  DFF \sreg_reg[411]  ( .D(c[412]), .CLK(clk), .RST(rst), .Q(c[411]) );
  DFF \sreg_reg[410]  ( .D(c[411]), .CLK(clk), .RST(rst), .Q(c[410]) );
  DFF \sreg_reg[409]  ( .D(c[410]), .CLK(clk), .RST(rst), .Q(c[409]) );
  DFF \sreg_reg[408]  ( .D(c[409]), .CLK(clk), .RST(rst), .Q(c[408]) );
  DFF \sreg_reg[407]  ( .D(c[408]), .CLK(clk), .RST(rst), .Q(c[407]) );
  DFF \sreg_reg[406]  ( .D(c[407]), .CLK(clk), .RST(rst), .Q(c[406]) );
  DFF \sreg_reg[405]  ( .D(c[406]), .CLK(clk), .RST(rst), .Q(c[405]) );
  DFF \sreg_reg[404]  ( .D(c[405]), .CLK(clk), .RST(rst), .Q(c[404]) );
  DFF \sreg_reg[403]  ( .D(c[404]), .CLK(clk), .RST(rst), .Q(c[403]) );
  DFF \sreg_reg[402]  ( .D(c[403]), .CLK(clk), .RST(rst), .Q(c[402]) );
  DFF \sreg_reg[401]  ( .D(c[402]), .CLK(clk), .RST(rst), .Q(c[401]) );
  DFF \sreg_reg[400]  ( .D(c[401]), .CLK(clk), .RST(rst), .Q(c[400]) );
  DFF \sreg_reg[399]  ( .D(c[400]), .CLK(clk), .RST(rst), .Q(c[399]) );
  DFF \sreg_reg[398]  ( .D(c[399]), .CLK(clk), .RST(rst), .Q(c[398]) );
  DFF \sreg_reg[397]  ( .D(c[398]), .CLK(clk), .RST(rst), .Q(c[397]) );
  DFF \sreg_reg[396]  ( .D(c[397]), .CLK(clk), .RST(rst), .Q(c[396]) );
  DFF \sreg_reg[395]  ( .D(c[396]), .CLK(clk), .RST(rst), .Q(c[395]) );
  DFF \sreg_reg[394]  ( .D(c[395]), .CLK(clk), .RST(rst), .Q(c[394]) );
  DFF \sreg_reg[393]  ( .D(c[394]), .CLK(clk), .RST(rst), .Q(c[393]) );
  DFF \sreg_reg[392]  ( .D(c[393]), .CLK(clk), .RST(rst), .Q(c[392]) );
  DFF \sreg_reg[391]  ( .D(c[392]), .CLK(clk), .RST(rst), .Q(c[391]) );
  DFF \sreg_reg[390]  ( .D(c[391]), .CLK(clk), .RST(rst), .Q(c[390]) );
  DFF \sreg_reg[389]  ( .D(c[390]), .CLK(clk), .RST(rst), .Q(c[389]) );
  DFF \sreg_reg[388]  ( .D(c[389]), .CLK(clk), .RST(rst), .Q(c[388]) );
  DFF \sreg_reg[387]  ( .D(c[388]), .CLK(clk), .RST(rst), .Q(c[387]) );
  DFF \sreg_reg[386]  ( .D(c[387]), .CLK(clk), .RST(rst), .Q(c[386]) );
  DFF \sreg_reg[385]  ( .D(c[386]), .CLK(clk), .RST(rst), .Q(c[385]) );
  DFF \sreg_reg[384]  ( .D(c[385]), .CLK(clk), .RST(rst), .Q(c[384]) );
  DFF \sreg_reg[383]  ( .D(c[384]), .CLK(clk), .RST(rst), .Q(c[383]) );
  DFF \sreg_reg[382]  ( .D(c[383]), .CLK(clk), .RST(rst), .Q(c[382]) );
  DFF \sreg_reg[381]  ( .D(c[382]), .CLK(clk), .RST(rst), .Q(c[381]) );
  DFF \sreg_reg[380]  ( .D(c[381]), .CLK(clk), .RST(rst), .Q(c[380]) );
  DFF \sreg_reg[379]  ( .D(c[380]), .CLK(clk), .RST(rst), .Q(c[379]) );
  DFF \sreg_reg[378]  ( .D(c[379]), .CLK(clk), .RST(rst), .Q(c[378]) );
  DFF \sreg_reg[377]  ( .D(c[378]), .CLK(clk), .RST(rst), .Q(c[377]) );
  DFF \sreg_reg[376]  ( .D(c[377]), .CLK(clk), .RST(rst), .Q(c[376]) );
  DFF \sreg_reg[375]  ( .D(c[376]), .CLK(clk), .RST(rst), .Q(c[375]) );
  DFF \sreg_reg[374]  ( .D(c[375]), .CLK(clk), .RST(rst), .Q(c[374]) );
  DFF \sreg_reg[373]  ( .D(c[374]), .CLK(clk), .RST(rst), .Q(c[373]) );
  DFF \sreg_reg[372]  ( .D(c[373]), .CLK(clk), .RST(rst), .Q(c[372]) );
  DFF \sreg_reg[371]  ( .D(c[372]), .CLK(clk), .RST(rst), .Q(c[371]) );
  DFF \sreg_reg[370]  ( .D(c[371]), .CLK(clk), .RST(rst), .Q(c[370]) );
  DFF \sreg_reg[369]  ( .D(c[370]), .CLK(clk), .RST(rst), .Q(c[369]) );
  DFF \sreg_reg[368]  ( .D(c[369]), .CLK(clk), .RST(rst), .Q(c[368]) );
  DFF \sreg_reg[367]  ( .D(c[368]), .CLK(clk), .RST(rst), .Q(c[367]) );
  DFF \sreg_reg[366]  ( .D(c[367]), .CLK(clk), .RST(rst), .Q(c[366]) );
  DFF \sreg_reg[365]  ( .D(c[366]), .CLK(clk), .RST(rst), .Q(c[365]) );
  DFF \sreg_reg[364]  ( .D(c[365]), .CLK(clk), .RST(rst), .Q(c[364]) );
  DFF \sreg_reg[363]  ( .D(c[364]), .CLK(clk), .RST(rst), .Q(c[363]) );
  DFF \sreg_reg[362]  ( .D(c[363]), .CLK(clk), .RST(rst), .Q(c[362]) );
  DFF \sreg_reg[361]  ( .D(c[362]), .CLK(clk), .RST(rst), .Q(c[361]) );
  DFF \sreg_reg[360]  ( .D(c[361]), .CLK(clk), .RST(rst), .Q(c[360]) );
  DFF \sreg_reg[359]  ( .D(c[360]), .CLK(clk), .RST(rst), .Q(c[359]) );
  DFF \sreg_reg[358]  ( .D(c[359]), .CLK(clk), .RST(rst), .Q(c[358]) );
  DFF \sreg_reg[357]  ( .D(c[358]), .CLK(clk), .RST(rst), .Q(c[357]) );
  DFF \sreg_reg[356]  ( .D(c[357]), .CLK(clk), .RST(rst), .Q(c[356]) );
  DFF \sreg_reg[355]  ( .D(c[356]), .CLK(clk), .RST(rst), .Q(c[355]) );
  DFF \sreg_reg[354]  ( .D(c[355]), .CLK(clk), .RST(rst), .Q(c[354]) );
  DFF \sreg_reg[353]  ( .D(c[354]), .CLK(clk), .RST(rst), .Q(c[353]) );
  DFF \sreg_reg[352]  ( .D(c[353]), .CLK(clk), .RST(rst), .Q(c[352]) );
  DFF \sreg_reg[351]  ( .D(c[352]), .CLK(clk), .RST(rst), .Q(c[351]) );
  DFF \sreg_reg[350]  ( .D(c[351]), .CLK(clk), .RST(rst), .Q(c[350]) );
  DFF \sreg_reg[349]  ( .D(c[350]), .CLK(clk), .RST(rst), .Q(c[349]) );
  DFF \sreg_reg[348]  ( .D(c[349]), .CLK(clk), .RST(rst), .Q(c[348]) );
  DFF \sreg_reg[347]  ( .D(c[348]), .CLK(clk), .RST(rst), .Q(c[347]) );
  DFF \sreg_reg[346]  ( .D(c[347]), .CLK(clk), .RST(rst), .Q(c[346]) );
  DFF \sreg_reg[345]  ( .D(c[346]), .CLK(clk), .RST(rst), .Q(c[345]) );
  DFF \sreg_reg[344]  ( .D(c[345]), .CLK(clk), .RST(rst), .Q(c[344]) );
  DFF \sreg_reg[343]  ( .D(c[344]), .CLK(clk), .RST(rst), .Q(c[343]) );
  DFF \sreg_reg[342]  ( .D(c[343]), .CLK(clk), .RST(rst), .Q(c[342]) );
  DFF \sreg_reg[341]  ( .D(c[342]), .CLK(clk), .RST(rst), .Q(c[341]) );
  DFF \sreg_reg[340]  ( .D(c[341]), .CLK(clk), .RST(rst), .Q(c[340]) );
  DFF \sreg_reg[339]  ( .D(c[340]), .CLK(clk), .RST(rst), .Q(c[339]) );
  DFF \sreg_reg[338]  ( .D(c[339]), .CLK(clk), .RST(rst), .Q(c[338]) );
  DFF \sreg_reg[337]  ( .D(c[338]), .CLK(clk), .RST(rst), .Q(c[337]) );
  DFF \sreg_reg[336]  ( .D(c[337]), .CLK(clk), .RST(rst), .Q(c[336]) );
  DFF \sreg_reg[335]  ( .D(c[336]), .CLK(clk), .RST(rst), .Q(c[335]) );
  DFF \sreg_reg[334]  ( .D(c[335]), .CLK(clk), .RST(rst), .Q(c[334]) );
  DFF \sreg_reg[333]  ( .D(c[334]), .CLK(clk), .RST(rst), .Q(c[333]) );
  DFF \sreg_reg[332]  ( .D(c[333]), .CLK(clk), .RST(rst), .Q(c[332]) );
  DFF \sreg_reg[331]  ( .D(c[332]), .CLK(clk), .RST(rst), .Q(c[331]) );
  DFF \sreg_reg[330]  ( .D(c[331]), .CLK(clk), .RST(rst), .Q(c[330]) );
  DFF \sreg_reg[329]  ( .D(c[330]), .CLK(clk), .RST(rst), .Q(c[329]) );
  DFF \sreg_reg[328]  ( .D(c[329]), .CLK(clk), .RST(rst), .Q(c[328]) );
  DFF \sreg_reg[327]  ( .D(c[328]), .CLK(clk), .RST(rst), .Q(c[327]) );
  DFF \sreg_reg[326]  ( .D(c[327]), .CLK(clk), .RST(rst), .Q(c[326]) );
  DFF \sreg_reg[325]  ( .D(c[326]), .CLK(clk), .RST(rst), .Q(c[325]) );
  DFF \sreg_reg[324]  ( .D(c[325]), .CLK(clk), .RST(rst), .Q(c[324]) );
  DFF \sreg_reg[323]  ( .D(c[324]), .CLK(clk), .RST(rst), .Q(c[323]) );
  DFF \sreg_reg[322]  ( .D(c[323]), .CLK(clk), .RST(rst), .Q(c[322]) );
  DFF \sreg_reg[321]  ( .D(c[322]), .CLK(clk), .RST(rst), .Q(c[321]) );
  DFF \sreg_reg[320]  ( .D(c[321]), .CLK(clk), .RST(rst), .Q(c[320]) );
  DFF \sreg_reg[319]  ( .D(c[320]), .CLK(clk), .RST(rst), .Q(c[319]) );
  DFF \sreg_reg[318]  ( .D(c[319]), .CLK(clk), .RST(rst), .Q(c[318]) );
  DFF \sreg_reg[317]  ( .D(c[318]), .CLK(clk), .RST(rst), .Q(c[317]) );
  DFF \sreg_reg[316]  ( .D(c[317]), .CLK(clk), .RST(rst), .Q(c[316]) );
  DFF \sreg_reg[315]  ( .D(c[316]), .CLK(clk), .RST(rst), .Q(c[315]) );
  DFF \sreg_reg[314]  ( .D(c[315]), .CLK(clk), .RST(rst), .Q(c[314]) );
  DFF \sreg_reg[313]  ( .D(c[314]), .CLK(clk), .RST(rst), .Q(c[313]) );
  DFF \sreg_reg[312]  ( .D(c[313]), .CLK(clk), .RST(rst), .Q(c[312]) );
  DFF \sreg_reg[311]  ( .D(c[312]), .CLK(clk), .RST(rst), .Q(c[311]) );
  DFF \sreg_reg[310]  ( .D(c[311]), .CLK(clk), .RST(rst), .Q(c[310]) );
  DFF \sreg_reg[309]  ( .D(c[310]), .CLK(clk), .RST(rst), .Q(c[309]) );
  DFF \sreg_reg[308]  ( .D(c[309]), .CLK(clk), .RST(rst), .Q(c[308]) );
  DFF \sreg_reg[307]  ( .D(c[308]), .CLK(clk), .RST(rst), .Q(c[307]) );
  DFF \sreg_reg[306]  ( .D(c[307]), .CLK(clk), .RST(rst), .Q(c[306]) );
  DFF \sreg_reg[305]  ( .D(c[306]), .CLK(clk), .RST(rst), .Q(c[305]) );
  DFF \sreg_reg[304]  ( .D(c[305]), .CLK(clk), .RST(rst), .Q(c[304]) );
  DFF \sreg_reg[303]  ( .D(c[304]), .CLK(clk), .RST(rst), .Q(c[303]) );
  DFF \sreg_reg[302]  ( .D(c[303]), .CLK(clk), .RST(rst), .Q(c[302]) );
  DFF \sreg_reg[301]  ( .D(c[302]), .CLK(clk), .RST(rst), .Q(c[301]) );
  DFF \sreg_reg[300]  ( .D(c[301]), .CLK(clk), .RST(rst), .Q(c[300]) );
  DFF \sreg_reg[299]  ( .D(c[300]), .CLK(clk), .RST(rst), .Q(c[299]) );
  DFF \sreg_reg[298]  ( .D(c[299]), .CLK(clk), .RST(rst), .Q(c[298]) );
  DFF \sreg_reg[297]  ( .D(c[298]), .CLK(clk), .RST(rst), .Q(c[297]) );
  DFF \sreg_reg[296]  ( .D(c[297]), .CLK(clk), .RST(rst), .Q(c[296]) );
  DFF \sreg_reg[295]  ( .D(c[296]), .CLK(clk), .RST(rst), .Q(c[295]) );
  DFF \sreg_reg[294]  ( .D(c[295]), .CLK(clk), .RST(rst), .Q(c[294]) );
  DFF \sreg_reg[293]  ( .D(c[294]), .CLK(clk), .RST(rst), .Q(c[293]) );
  DFF \sreg_reg[292]  ( .D(c[293]), .CLK(clk), .RST(rst), .Q(c[292]) );
  DFF \sreg_reg[291]  ( .D(c[292]), .CLK(clk), .RST(rst), .Q(c[291]) );
  DFF \sreg_reg[290]  ( .D(c[291]), .CLK(clk), .RST(rst), .Q(c[290]) );
  DFF \sreg_reg[289]  ( .D(c[290]), .CLK(clk), .RST(rst), .Q(c[289]) );
  DFF \sreg_reg[288]  ( .D(c[289]), .CLK(clk), .RST(rst), .Q(c[288]) );
  DFF \sreg_reg[287]  ( .D(c[288]), .CLK(clk), .RST(rst), .Q(c[287]) );
  DFF \sreg_reg[286]  ( .D(c[287]), .CLK(clk), .RST(rst), .Q(c[286]) );
  DFF \sreg_reg[285]  ( .D(c[286]), .CLK(clk), .RST(rst), .Q(c[285]) );
  DFF \sreg_reg[284]  ( .D(c[285]), .CLK(clk), .RST(rst), .Q(c[284]) );
  DFF \sreg_reg[283]  ( .D(c[284]), .CLK(clk), .RST(rst), .Q(c[283]) );
  DFF \sreg_reg[282]  ( .D(c[283]), .CLK(clk), .RST(rst), .Q(c[282]) );
  DFF \sreg_reg[281]  ( .D(c[282]), .CLK(clk), .RST(rst), .Q(c[281]) );
  DFF \sreg_reg[280]  ( .D(c[281]), .CLK(clk), .RST(rst), .Q(c[280]) );
  DFF \sreg_reg[279]  ( .D(c[280]), .CLK(clk), .RST(rst), .Q(c[279]) );
  DFF \sreg_reg[278]  ( .D(c[279]), .CLK(clk), .RST(rst), .Q(c[278]) );
  DFF \sreg_reg[277]  ( .D(c[278]), .CLK(clk), .RST(rst), .Q(c[277]) );
  DFF \sreg_reg[276]  ( .D(c[277]), .CLK(clk), .RST(rst), .Q(c[276]) );
  DFF \sreg_reg[275]  ( .D(c[276]), .CLK(clk), .RST(rst), .Q(c[275]) );
  DFF \sreg_reg[274]  ( .D(c[275]), .CLK(clk), .RST(rst), .Q(c[274]) );
  DFF \sreg_reg[273]  ( .D(c[274]), .CLK(clk), .RST(rst), .Q(c[273]) );
  DFF \sreg_reg[272]  ( .D(c[273]), .CLK(clk), .RST(rst), .Q(c[272]) );
  DFF \sreg_reg[271]  ( .D(c[272]), .CLK(clk), .RST(rst), .Q(c[271]) );
  DFF \sreg_reg[270]  ( .D(c[271]), .CLK(clk), .RST(rst), .Q(c[270]) );
  DFF \sreg_reg[269]  ( .D(c[270]), .CLK(clk), .RST(rst), .Q(c[269]) );
  DFF \sreg_reg[268]  ( .D(c[269]), .CLK(clk), .RST(rst), .Q(c[268]) );
  DFF \sreg_reg[267]  ( .D(c[268]), .CLK(clk), .RST(rst), .Q(c[267]) );
  DFF \sreg_reg[266]  ( .D(c[267]), .CLK(clk), .RST(rst), .Q(c[266]) );
  DFF \sreg_reg[265]  ( .D(c[266]), .CLK(clk), .RST(rst), .Q(c[265]) );
  DFF \sreg_reg[264]  ( .D(c[265]), .CLK(clk), .RST(rst), .Q(c[264]) );
  DFF \sreg_reg[263]  ( .D(c[264]), .CLK(clk), .RST(rst), .Q(c[263]) );
  DFF \sreg_reg[262]  ( .D(c[263]), .CLK(clk), .RST(rst), .Q(c[262]) );
  DFF \sreg_reg[261]  ( .D(c[262]), .CLK(clk), .RST(rst), .Q(c[261]) );
  DFF \sreg_reg[260]  ( .D(c[261]), .CLK(clk), .RST(rst), .Q(c[260]) );
  DFF \sreg_reg[259]  ( .D(c[260]), .CLK(clk), .RST(rst), .Q(c[259]) );
  DFF \sreg_reg[258]  ( .D(c[259]), .CLK(clk), .RST(rst), .Q(c[258]) );
  DFF \sreg_reg[257]  ( .D(c[258]), .CLK(clk), .RST(rst), .Q(c[257]) );
  DFF \sreg_reg[256]  ( .D(c[257]), .CLK(clk), .RST(rst), .Q(c[256]) );
  DFF \sreg_reg[255]  ( .D(c[256]), .CLK(clk), .RST(rst), .Q(c[255]) );
  DFF \sreg_reg[254]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[254]) );
  DFF \sreg_reg[253]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[253]) );
  DFF \sreg_reg[252]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[252]) );
  DFF \sreg_reg[251]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[251]) );
  DFF \sreg_reg[250]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[250]) );
  DFF \sreg_reg[249]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[249]) );
  DFF \sreg_reg[248]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[248]) );
  DFF \sreg_reg[247]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[247]) );
  DFF \sreg_reg[246]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[246]) );
  DFF \sreg_reg[245]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[245]) );
  DFF \sreg_reg[244]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[244]) );
  DFF \sreg_reg[243]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[243]) );
  DFF \sreg_reg[242]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[242]) );
  DFF \sreg_reg[241]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[241]) );
  DFF \sreg_reg[240]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[240]) );
  DFF \sreg_reg[239]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[238]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[237]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[236]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[235]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[234]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[233]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[232]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[231]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[230]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[229]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[228]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[227]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[226]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[225]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[224]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[223]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[222]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[221]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[220]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[219]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[218]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[217]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[216]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[215]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[214]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[213]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[212]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[211]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[210]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[209]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[208]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[207]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[206]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[205]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[204]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[203]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[202]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[201]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[200]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[199]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[198]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[197]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[196]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[195]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[194]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[193]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[192]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[191]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[190]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[189]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[188]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[187]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[186]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[185]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[184]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[183]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[182]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[181]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[180]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[179]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[178]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[177]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[176]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[175]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[174]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[173]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[172]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[171]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[170]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[169]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[168]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[167]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[166]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[165]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[164]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[163]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[162]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[161]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[160]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[159]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[158]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[157]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[156]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[155]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[154]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[153]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[152]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[151]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[150]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[149]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[148]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[147]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[146]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[145]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[144]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[143]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[142]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[141]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[140]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[139]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[138]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[137]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[136]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[135]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[134]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[133]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[132]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[131]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[130]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[129]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[128]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[127]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[126]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[125]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[124]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[123]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[3]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[2]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[1]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U4 ( .A(b[0]), .B(a[0]), .Z(n1) );
  XNOR U5 ( .A(n1), .B(sreg[1023]), .Z(c[1023]) );
  NAND U6 ( .A(b[0]), .B(a[1]), .Z(n6) );
  XOR U7 ( .A(n6), .B(sreg[1024]), .Z(n2) );
  NANDN U8 ( .A(n1), .B(sreg[1023]), .Z(n3) );
  NAND U9 ( .A(n2), .B(n3), .Z(n5) );
  XOR U10 ( .A(a[1]), .B(sreg[1024]), .Z(n4) );
  ANDN U11 ( .B(n4), .A(n3), .Z(n7) );
  ANDN U12 ( .B(n5), .A(n7), .Z(c[1024]) );
  NAND U13 ( .A(b[0]), .B(a[2]), .Z(n9) );
  XOR U14 ( .A(sreg[1025]), .B(n9), .Z(n11) );
  NANDN U15 ( .A(n6), .B(sreg[1024]), .Z(n8) );
  ANDN U16 ( .B(n8), .A(n7), .Z(n10) );
  XOR U17 ( .A(n11), .B(n10), .Z(c[1025]) );
  NAND U18 ( .A(b[0]), .B(a[3]), .Z(n14) );
  XOR U19 ( .A(sreg[1026]), .B(n14), .Z(n16) );
  NANDN U20 ( .A(n9), .B(sreg[1025]), .Z(n13) );
  OR U21 ( .A(n11), .B(n10), .Z(n12) );
  AND U22 ( .A(n13), .B(n12), .Z(n15) );
  XOR U23 ( .A(n16), .B(n15), .Z(c[1026]) );
  NAND U24 ( .A(b[0]), .B(a[4]), .Z(n19) );
  XOR U25 ( .A(sreg[1027]), .B(n19), .Z(n21) );
  NANDN U26 ( .A(n14), .B(sreg[1026]), .Z(n18) );
  OR U27 ( .A(n16), .B(n15), .Z(n17) );
  AND U28 ( .A(n18), .B(n17), .Z(n20) );
  XOR U29 ( .A(n21), .B(n20), .Z(c[1027]) );
  NAND U30 ( .A(b[0]), .B(a[5]), .Z(n24) );
  XOR U31 ( .A(sreg[1028]), .B(n24), .Z(n26) );
  NANDN U32 ( .A(n19), .B(sreg[1027]), .Z(n23) );
  OR U33 ( .A(n21), .B(n20), .Z(n22) );
  AND U34 ( .A(n23), .B(n22), .Z(n25) );
  XOR U35 ( .A(n26), .B(n25), .Z(c[1028]) );
  NAND U36 ( .A(b[0]), .B(a[6]), .Z(n29) );
  XOR U37 ( .A(sreg[1029]), .B(n29), .Z(n31) );
  NANDN U38 ( .A(n24), .B(sreg[1028]), .Z(n28) );
  OR U39 ( .A(n26), .B(n25), .Z(n27) );
  AND U40 ( .A(n28), .B(n27), .Z(n30) );
  XOR U41 ( .A(n31), .B(n30), .Z(c[1029]) );
  NAND U42 ( .A(b[0]), .B(a[7]), .Z(n34) );
  XOR U43 ( .A(sreg[1030]), .B(n34), .Z(n36) );
  NANDN U44 ( .A(n29), .B(sreg[1029]), .Z(n33) );
  OR U45 ( .A(n31), .B(n30), .Z(n32) );
  AND U46 ( .A(n33), .B(n32), .Z(n35) );
  XOR U47 ( .A(n36), .B(n35), .Z(c[1030]) );
  NAND U48 ( .A(b[0]), .B(a[8]), .Z(n39) );
  XOR U49 ( .A(sreg[1031]), .B(n39), .Z(n41) );
  NANDN U50 ( .A(n34), .B(sreg[1030]), .Z(n38) );
  OR U51 ( .A(n36), .B(n35), .Z(n37) );
  AND U52 ( .A(n38), .B(n37), .Z(n40) );
  XOR U53 ( .A(n41), .B(n40), .Z(c[1031]) );
  NAND U54 ( .A(b[0]), .B(a[9]), .Z(n44) );
  XOR U55 ( .A(sreg[1032]), .B(n44), .Z(n46) );
  NANDN U56 ( .A(n39), .B(sreg[1031]), .Z(n43) );
  OR U57 ( .A(n41), .B(n40), .Z(n42) );
  AND U58 ( .A(n43), .B(n42), .Z(n45) );
  XOR U59 ( .A(n46), .B(n45), .Z(c[1032]) );
  NAND U60 ( .A(b[0]), .B(a[10]), .Z(n49) );
  XOR U61 ( .A(sreg[1033]), .B(n49), .Z(n51) );
  NANDN U62 ( .A(n44), .B(sreg[1032]), .Z(n48) );
  OR U63 ( .A(n46), .B(n45), .Z(n47) );
  AND U64 ( .A(n48), .B(n47), .Z(n50) );
  XOR U65 ( .A(n51), .B(n50), .Z(c[1033]) );
  NAND U66 ( .A(b[0]), .B(a[11]), .Z(n54) );
  XOR U67 ( .A(sreg[1034]), .B(n54), .Z(n56) );
  NANDN U68 ( .A(n49), .B(sreg[1033]), .Z(n53) );
  OR U69 ( .A(n51), .B(n50), .Z(n52) );
  AND U70 ( .A(n53), .B(n52), .Z(n55) );
  XOR U71 ( .A(n56), .B(n55), .Z(c[1034]) );
  NAND U72 ( .A(b[0]), .B(a[12]), .Z(n59) );
  XOR U73 ( .A(sreg[1035]), .B(n59), .Z(n61) );
  NANDN U74 ( .A(n54), .B(sreg[1034]), .Z(n58) );
  OR U75 ( .A(n56), .B(n55), .Z(n57) );
  AND U76 ( .A(n58), .B(n57), .Z(n60) );
  XOR U77 ( .A(n61), .B(n60), .Z(c[1035]) );
  NAND U78 ( .A(b[0]), .B(a[13]), .Z(n64) );
  XOR U79 ( .A(sreg[1036]), .B(n64), .Z(n66) );
  NANDN U80 ( .A(n59), .B(sreg[1035]), .Z(n63) );
  OR U81 ( .A(n61), .B(n60), .Z(n62) );
  AND U82 ( .A(n63), .B(n62), .Z(n65) );
  XOR U83 ( .A(n66), .B(n65), .Z(c[1036]) );
  NAND U84 ( .A(b[0]), .B(a[14]), .Z(n69) );
  XOR U85 ( .A(sreg[1037]), .B(n69), .Z(n71) );
  NANDN U86 ( .A(n64), .B(sreg[1036]), .Z(n68) );
  OR U87 ( .A(n66), .B(n65), .Z(n67) );
  AND U88 ( .A(n68), .B(n67), .Z(n70) );
  XOR U89 ( .A(n71), .B(n70), .Z(c[1037]) );
  NAND U90 ( .A(b[0]), .B(a[15]), .Z(n74) );
  XOR U91 ( .A(sreg[1038]), .B(n74), .Z(n76) );
  NANDN U92 ( .A(n69), .B(sreg[1037]), .Z(n73) );
  OR U93 ( .A(n71), .B(n70), .Z(n72) );
  AND U94 ( .A(n73), .B(n72), .Z(n75) );
  XOR U95 ( .A(n76), .B(n75), .Z(c[1038]) );
  NAND U96 ( .A(b[0]), .B(a[16]), .Z(n79) );
  XOR U97 ( .A(sreg[1039]), .B(n79), .Z(n81) );
  NANDN U98 ( .A(n74), .B(sreg[1038]), .Z(n78) );
  OR U99 ( .A(n76), .B(n75), .Z(n77) );
  AND U100 ( .A(n78), .B(n77), .Z(n80) );
  XOR U101 ( .A(n81), .B(n80), .Z(c[1039]) );
  NAND U102 ( .A(b[0]), .B(a[17]), .Z(n84) );
  XOR U103 ( .A(sreg[1040]), .B(n84), .Z(n86) );
  NANDN U104 ( .A(n79), .B(sreg[1039]), .Z(n83) );
  OR U105 ( .A(n81), .B(n80), .Z(n82) );
  AND U106 ( .A(n83), .B(n82), .Z(n85) );
  XOR U107 ( .A(n86), .B(n85), .Z(c[1040]) );
  NAND U108 ( .A(b[0]), .B(a[18]), .Z(n89) );
  XOR U109 ( .A(sreg[1041]), .B(n89), .Z(n91) );
  NANDN U110 ( .A(n84), .B(sreg[1040]), .Z(n88) );
  OR U111 ( .A(n86), .B(n85), .Z(n87) );
  AND U112 ( .A(n88), .B(n87), .Z(n90) );
  XOR U113 ( .A(n91), .B(n90), .Z(c[1041]) );
  NAND U114 ( .A(b[0]), .B(a[19]), .Z(n94) );
  XOR U115 ( .A(sreg[1042]), .B(n94), .Z(n96) );
  NANDN U116 ( .A(n89), .B(sreg[1041]), .Z(n93) );
  OR U117 ( .A(n91), .B(n90), .Z(n92) );
  AND U118 ( .A(n93), .B(n92), .Z(n95) );
  XOR U119 ( .A(n96), .B(n95), .Z(c[1042]) );
  NAND U120 ( .A(b[0]), .B(a[20]), .Z(n99) );
  XOR U121 ( .A(sreg[1043]), .B(n99), .Z(n101) );
  NANDN U122 ( .A(n94), .B(sreg[1042]), .Z(n98) );
  OR U123 ( .A(n96), .B(n95), .Z(n97) );
  AND U124 ( .A(n98), .B(n97), .Z(n100) );
  XOR U125 ( .A(n101), .B(n100), .Z(c[1043]) );
  NAND U126 ( .A(b[0]), .B(a[21]), .Z(n104) );
  XOR U127 ( .A(sreg[1044]), .B(n104), .Z(n106) );
  NANDN U128 ( .A(n99), .B(sreg[1043]), .Z(n103) );
  OR U129 ( .A(n101), .B(n100), .Z(n102) );
  AND U130 ( .A(n103), .B(n102), .Z(n105) );
  XOR U131 ( .A(n106), .B(n105), .Z(c[1044]) );
  NAND U132 ( .A(b[0]), .B(a[22]), .Z(n109) );
  XOR U133 ( .A(sreg[1045]), .B(n109), .Z(n111) );
  NANDN U134 ( .A(n104), .B(sreg[1044]), .Z(n108) );
  OR U135 ( .A(n106), .B(n105), .Z(n107) );
  AND U136 ( .A(n108), .B(n107), .Z(n110) );
  XOR U137 ( .A(n111), .B(n110), .Z(c[1045]) );
  NAND U138 ( .A(b[0]), .B(a[23]), .Z(n114) );
  XOR U139 ( .A(sreg[1046]), .B(n114), .Z(n116) );
  NANDN U140 ( .A(n109), .B(sreg[1045]), .Z(n113) );
  OR U141 ( .A(n111), .B(n110), .Z(n112) );
  AND U142 ( .A(n113), .B(n112), .Z(n115) );
  XOR U143 ( .A(n116), .B(n115), .Z(c[1046]) );
  NAND U144 ( .A(b[0]), .B(a[24]), .Z(n119) );
  XOR U145 ( .A(sreg[1047]), .B(n119), .Z(n121) );
  NANDN U146 ( .A(n114), .B(sreg[1046]), .Z(n118) );
  OR U147 ( .A(n116), .B(n115), .Z(n117) );
  AND U148 ( .A(n118), .B(n117), .Z(n120) );
  XOR U149 ( .A(n121), .B(n120), .Z(c[1047]) );
  NAND U150 ( .A(b[0]), .B(a[25]), .Z(n124) );
  XOR U151 ( .A(sreg[1048]), .B(n124), .Z(n126) );
  NANDN U152 ( .A(n119), .B(sreg[1047]), .Z(n123) );
  OR U153 ( .A(n121), .B(n120), .Z(n122) );
  AND U154 ( .A(n123), .B(n122), .Z(n125) );
  XOR U155 ( .A(n126), .B(n125), .Z(c[1048]) );
  NAND U156 ( .A(b[0]), .B(a[26]), .Z(n129) );
  XOR U157 ( .A(sreg[1049]), .B(n129), .Z(n131) );
  NANDN U158 ( .A(n124), .B(sreg[1048]), .Z(n128) );
  OR U159 ( .A(n126), .B(n125), .Z(n127) );
  AND U160 ( .A(n128), .B(n127), .Z(n130) );
  XOR U161 ( .A(n131), .B(n130), .Z(c[1049]) );
  NAND U162 ( .A(b[0]), .B(a[27]), .Z(n134) );
  XOR U163 ( .A(sreg[1050]), .B(n134), .Z(n136) );
  NANDN U164 ( .A(n129), .B(sreg[1049]), .Z(n133) );
  OR U165 ( .A(n131), .B(n130), .Z(n132) );
  AND U166 ( .A(n133), .B(n132), .Z(n135) );
  XOR U167 ( .A(n136), .B(n135), .Z(c[1050]) );
  NAND U168 ( .A(b[0]), .B(a[28]), .Z(n139) );
  XOR U169 ( .A(sreg[1051]), .B(n139), .Z(n141) );
  NANDN U170 ( .A(n134), .B(sreg[1050]), .Z(n138) );
  OR U171 ( .A(n136), .B(n135), .Z(n137) );
  AND U172 ( .A(n138), .B(n137), .Z(n140) );
  XOR U173 ( .A(n141), .B(n140), .Z(c[1051]) );
  NAND U174 ( .A(b[0]), .B(a[29]), .Z(n144) );
  XOR U175 ( .A(sreg[1052]), .B(n144), .Z(n146) );
  NANDN U176 ( .A(n139), .B(sreg[1051]), .Z(n143) );
  OR U177 ( .A(n141), .B(n140), .Z(n142) );
  AND U178 ( .A(n143), .B(n142), .Z(n145) );
  XOR U179 ( .A(n146), .B(n145), .Z(c[1052]) );
  NAND U180 ( .A(b[0]), .B(a[30]), .Z(n149) );
  XOR U181 ( .A(sreg[1053]), .B(n149), .Z(n151) );
  NANDN U182 ( .A(n144), .B(sreg[1052]), .Z(n148) );
  OR U183 ( .A(n146), .B(n145), .Z(n147) );
  AND U184 ( .A(n148), .B(n147), .Z(n150) );
  XOR U185 ( .A(n151), .B(n150), .Z(c[1053]) );
  NAND U186 ( .A(b[0]), .B(a[31]), .Z(n154) );
  XOR U187 ( .A(sreg[1054]), .B(n154), .Z(n156) );
  NANDN U188 ( .A(n149), .B(sreg[1053]), .Z(n153) );
  OR U189 ( .A(n151), .B(n150), .Z(n152) );
  AND U190 ( .A(n153), .B(n152), .Z(n155) );
  XOR U191 ( .A(n156), .B(n155), .Z(c[1054]) );
  NAND U192 ( .A(b[0]), .B(a[32]), .Z(n159) );
  XOR U193 ( .A(sreg[1055]), .B(n159), .Z(n161) );
  NANDN U194 ( .A(n154), .B(sreg[1054]), .Z(n158) );
  OR U195 ( .A(n156), .B(n155), .Z(n157) );
  AND U196 ( .A(n158), .B(n157), .Z(n160) );
  XOR U197 ( .A(n161), .B(n160), .Z(c[1055]) );
  NAND U198 ( .A(b[0]), .B(a[33]), .Z(n164) );
  XOR U199 ( .A(sreg[1056]), .B(n164), .Z(n166) );
  NANDN U200 ( .A(n159), .B(sreg[1055]), .Z(n163) );
  OR U201 ( .A(n161), .B(n160), .Z(n162) );
  AND U202 ( .A(n163), .B(n162), .Z(n165) );
  XOR U203 ( .A(n166), .B(n165), .Z(c[1056]) );
  NAND U204 ( .A(b[0]), .B(a[34]), .Z(n169) );
  XOR U205 ( .A(sreg[1057]), .B(n169), .Z(n171) );
  NANDN U206 ( .A(n164), .B(sreg[1056]), .Z(n168) );
  OR U207 ( .A(n166), .B(n165), .Z(n167) );
  AND U208 ( .A(n168), .B(n167), .Z(n170) );
  XOR U209 ( .A(n171), .B(n170), .Z(c[1057]) );
  NAND U210 ( .A(b[0]), .B(a[35]), .Z(n174) );
  XOR U211 ( .A(sreg[1058]), .B(n174), .Z(n176) );
  NANDN U212 ( .A(n169), .B(sreg[1057]), .Z(n173) );
  OR U213 ( .A(n171), .B(n170), .Z(n172) );
  AND U214 ( .A(n173), .B(n172), .Z(n175) );
  XOR U215 ( .A(n176), .B(n175), .Z(c[1058]) );
  NAND U216 ( .A(b[0]), .B(a[36]), .Z(n179) );
  XOR U217 ( .A(sreg[1059]), .B(n179), .Z(n181) );
  NANDN U218 ( .A(n174), .B(sreg[1058]), .Z(n178) );
  OR U219 ( .A(n176), .B(n175), .Z(n177) );
  AND U220 ( .A(n178), .B(n177), .Z(n180) );
  XOR U221 ( .A(n181), .B(n180), .Z(c[1059]) );
  NAND U222 ( .A(b[0]), .B(a[37]), .Z(n184) );
  XOR U223 ( .A(sreg[1060]), .B(n184), .Z(n186) );
  NANDN U224 ( .A(n179), .B(sreg[1059]), .Z(n183) );
  OR U225 ( .A(n181), .B(n180), .Z(n182) );
  AND U226 ( .A(n183), .B(n182), .Z(n185) );
  XOR U227 ( .A(n186), .B(n185), .Z(c[1060]) );
  NAND U228 ( .A(b[0]), .B(a[38]), .Z(n189) );
  XOR U229 ( .A(sreg[1061]), .B(n189), .Z(n191) );
  NANDN U230 ( .A(n184), .B(sreg[1060]), .Z(n188) );
  OR U231 ( .A(n186), .B(n185), .Z(n187) );
  AND U232 ( .A(n188), .B(n187), .Z(n190) );
  XOR U233 ( .A(n191), .B(n190), .Z(c[1061]) );
  NAND U234 ( .A(b[0]), .B(a[39]), .Z(n194) );
  XOR U235 ( .A(sreg[1062]), .B(n194), .Z(n196) );
  NANDN U236 ( .A(n189), .B(sreg[1061]), .Z(n193) );
  OR U237 ( .A(n191), .B(n190), .Z(n192) );
  AND U238 ( .A(n193), .B(n192), .Z(n195) );
  XOR U239 ( .A(n196), .B(n195), .Z(c[1062]) );
  NAND U240 ( .A(b[0]), .B(a[40]), .Z(n199) );
  XOR U241 ( .A(sreg[1063]), .B(n199), .Z(n201) );
  NANDN U242 ( .A(n194), .B(sreg[1062]), .Z(n198) );
  OR U243 ( .A(n196), .B(n195), .Z(n197) );
  AND U244 ( .A(n198), .B(n197), .Z(n200) );
  XOR U245 ( .A(n201), .B(n200), .Z(c[1063]) );
  NAND U246 ( .A(b[0]), .B(a[41]), .Z(n204) );
  XOR U247 ( .A(sreg[1064]), .B(n204), .Z(n206) );
  NANDN U248 ( .A(n199), .B(sreg[1063]), .Z(n203) );
  OR U249 ( .A(n201), .B(n200), .Z(n202) );
  AND U250 ( .A(n203), .B(n202), .Z(n205) );
  XOR U251 ( .A(n206), .B(n205), .Z(c[1064]) );
  NAND U252 ( .A(b[0]), .B(a[42]), .Z(n209) );
  XOR U253 ( .A(sreg[1065]), .B(n209), .Z(n211) );
  NANDN U254 ( .A(n204), .B(sreg[1064]), .Z(n208) );
  OR U255 ( .A(n206), .B(n205), .Z(n207) );
  AND U256 ( .A(n208), .B(n207), .Z(n210) );
  XOR U257 ( .A(n211), .B(n210), .Z(c[1065]) );
  NAND U258 ( .A(b[0]), .B(a[43]), .Z(n214) );
  XOR U259 ( .A(sreg[1066]), .B(n214), .Z(n216) );
  NANDN U260 ( .A(n209), .B(sreg[1065]), .Z(n213) );
  OR U261 ( .A(n211), .B(n210), .Z(n212) );
  AND U262 ( .A(n213), .B(n212), .Z(n215) );
  XOR U263 ( .A(n216), .B(n215), .Z(c[1066]) );
  NAND U264 ( .A(b[0]), .B(a[44]), .Z(n219) );
  XOR U265 ( .A(sreg[1067]), .B(n219), .Z(n221) );
  NANDN U266 ( .A(n214), .B(sreg[1066]), .Z(n218) );
  OR U267 ( .A(n216), .B(n215), .Z(n217) );
  AND U268 ( .A(n218), .B(n217), .Z(n220) );
  XOR U269 ( .A(n221), .B(n220), .Z(c[1067]) );
  NAND U270 ( .A(b[0]), .B(a[45]), .Z(n224) );
  XOR U271 ( .A(sreg[1068]), .B(n224), .Z(n226) );
  NANDN U272 ( .A(n219), .B(sreg[1067]), .Z(n223) );
  OR U273 ( .A(n221), .B(n220), .Z(n222) );
  AND U274 ( .A(n223), .B(n222), .Z(n225) );
  XOR U275 ( .A(n226), .B(n225), .Z(c[1068]) );
  NAND U276 ( .A(b[0]), .B(a[46]), .Z(n229) );
  XOR U277 ( .A(sreg[1069]), .B(n229), .Z(n231) );
  NANDN U278 ( .A(n224), .B(sreg[1068]), .Z(n228) );
  OR U279 ( .A(n226), .B(n225), .Z(n227) );
  AND U280 ( .A(n228), .B(n227), .Z(n230) );
  XOR U281 ( .A(n231), .B(n230), .Z(c[1069]) );
  NAND U282 ( .A(b[0]), .B(a[47]), .Z(n234) );
  XOR U283 ( .A(sreg[1070]), .B(n234), .Z(n236) );
  NANDN U284 ( .A(n229), .B(sreg[1069]), .Z(n233) );
  OR U285 ( .A(n231), .B(n230), .Z(n232) );
  AND U286 ( .A(n233), .B(n232), .Z(n235) );
  XOR U287 ( .A(n236), .B(n235), .Z(c[1070]) );
  NAND U288 ( .A(b[0]), .B(a[48]), .Z(n239) );
  XOR U289 ( .A(sreg[1071]), .B(n239), .Z(n241) );
  NANDN U290 ( .A(n234), .B(sreg[1070]), .Z(n238) );
  OR U291 ( .A(n236), .B(n235), .Z(n237) );
  AND U292 ( .A(n238), .B(n237), .Z(n240) );
  XOR U293 ( .A(n241), .B(n240), .Z(c[1071]) );
  NAND U294 ( .A(b[0]), .B(a[49]), .Z(n244) );
  XOR U295 ( .A(sreg[1072]), .B(n244), .Z(n246) );
  NANDN U296 ( .A(n239), .B(sreg[1071]), .Z(n243) );
  OR U297 ( .A(n241), .B(n240), .Z(n242) );
  AND U298 ( .A(n243), .B(n242), .Z(n245) );
  XOR U299 ( .A(n246), .B(n245), .Z(c[1072]) );
  NAND U300 ( .A(b[0]), .B(a[50]), .Z(n249) );
  XOR U301 ( .A(sreg[1073]), .B(n249), .Z(n251) );
  NANDN U302 ( .A(n244), .B(sreg[1072]), .Z(n248) );
  OR U303 ( .A(n246), .B(n245), .Z(n247) );
  AND U304 ( .A(n248), .B(n247), .Z(n250) );
  XOR U305 ( .A(n251), .B(n250), .Z(c[1073]) );
  NAND U306 ( .A(b[0]), .B(a[51]), .Z(n254) );
  XOR U307 ( .A(sreg[1074]), .B(n254), .Z(n256) );
  NANDN U308 ( .A(n249), .B(sreg[1073]), .Z(n253) );
  OR U309 ( .A(n251), .B(n250), .Z(n252) );
  AND U310 ( .A(n253), .B(n252), .Z(n255) );
  XOR U311 ( .A(n256), .B(n255), .Z(c[1074]) );
  NAND U312 ( .A(b[0]), .B(a[52]), .Z(n259) );
  XOR U313 ( .A(sreg[1075]), .B(n259), .Z(n261) );
  NANDN U314 ( .A(n254), .B(sreg[1074]), .Z(n258) );
  OR U315 ( .A(n256), .B(n255), .Z(n257) );
  AND U316 ( .A(n258), .B(n257), .Z(n260) );
  XOR U317 ( .A(n261), .B(n260), .Z(c[1075]) );
  NAND U318 ( .A(b[0]), .B(a[53]), .Z(n264) );
  XOR U319 ( .A(sreg[1076]), .B(n264), .Z(n266) );
  NANDN U320 ( .A(n259), .B(sreg[1075]), .Z(n263) );
  OR U321 ( .A(n261), .B(n260), .Z(n262) );
  AND U322 ( .A(n263), .B(n262), .Z(n265) );
  XOR U323 ( .A(n266), .B(n265), .Z(c[1076]) );
  NAND U324 ( .A(b[0]), .B(a[54]), .Z(n269) );
  XOR U325 ( .A(sreg[1077]), .B(n269), .Z(n271) );
  NANDN U326 ( .A(n264), .B(sreg[1076]), .Z(n268) );
  OR U327 ( .A(n266), .B(n265), .Z(n267) );
  AND U328 ( .A(n268), .B(n267), .Z(n270) );
  XOR U329 ( .A(n271), .B(n270), .Z(c[1077]) );
  NAND U330 ( .A(b[0]), .B(a[55]), .Z(n274) );
  XOR U331 ( .A(sreg[1078]), .B(n274), .Z(n276) );
  NANDN U332 ( .A(n269), .B(sreg[1077]), .Z(n273) );
  OR U333 ( .A(n271), .B(n270), .Z(n272) );
  AND U334 ( .A(n273), .B(n272), .Z(n275) );
  XOR U335 ( .A(n276), .B(n275), .Z(c[1078]) );
  NAND U336 ( .A(b[0]), .B(a[56]), .Z(n279) );
  XOR U337 ( .A(sreg[1079]), .B(n279), .Z(n281) );
  NANDN U338 ( .A(n274), .B(sreg[1078]), .Z(n278) );
  OR U339 ( .A(n276), .B(n275), .Z(n277) );
  AND U340 ( .A(n278), .B(n277), .Z(n280) );
  XOR U341 ( .A(n281), .B(n280), .Z(c[1079]) );
  NAND U342 ( .A(b[0]), .B(a[57]), .Z(n284) );
  XOR U343 ( .A(sreg[1080]), .B(n284), .Z(n286) );
  NANDN U344 ( .A(n279), .B(sreg[1079]), .Z(n283) );
  OR U345 ( .A(n281), .B(n280), .Z(n282) );
  AND U346 ( .A(n283), .B(n282), .Z(n285) );
  XOR U347 ( .A(n286), .B(n285), .Z(c[1080]) );
  NAND U348 ( .A(b[0]), .B(a[58]), .Z(n289) );
  XOR U349 ( .A(sreg[1081]), .B(n289), .Z(n291) );
  NANDN U350 ( .A(n284), .B(sreg[1080]), .Z(n288) );
  OR U351 ( .A(n286), .B(n285), .Z(n287) );
  AND U352 ( .A(n288), .B(n287), .Z(n290) );
  XOR U353 ( .A(n291), .B(n290), .Z(c[1081]) );
  NAND U354 ( .A(b[0]), .B(a[59]), .Z(n294) );
  XOR U355 ( .A(sreg[1082]), .B(n294), .Z(n296) );
  NANDN U356 ( .A(n289), .B(sreg[1081]), .Z(n293) );
  OR U357 ( .A(n291), .B(n290), .Z(n292) );
  AND U358 ( .A(n293), .B(n292), .Z(n295) );
  XOR U359 ( .A(n296), .B(n295), .Z(c[1082]) );
  NAND U360 ( .A(b[0]), .B(a[60]), .Z(n299) );
  XOR U361 ( .A(sreg[1083]), .B(n299), .Z(n301) );
  NANDN U362 ( .A(n294), .B(sreg[1082]), .Z(n298) );
  OR U363 ( .A(n296), .B(n295), .Z(n297) );
  AND U364 ( .A(n298), .B(n297), .Z(n300) );
  XOR U365 ( .A(n301), .B(n300), .Z(c[1083]) );
  NAND U366 ( .A(b[0]), .B(a[61]), .Z(n304) );
  XOR U367 ( .A(sreg[1084]), .B(n304), .Z(n306) );
  NANDN U368 ( .A(n299), .B(sreg[1083]), .Z(n303) );
  OR U369 ( .A(n301), .B(n300), .Z(n302) );
  AND U370 ( .A(n303), .B(n302), .Z(n305) );
  XOR U371 ( .A(n306), .B(n305), .Z(c[1084]) );
  NAND U372 ( .A(b[0]), .B(a[62]), .Z(n309) );
  XOR U373 ( .A(sreg[1085]), .B(n309), .Z(n311) );
  NANDN U374 ( .A(n304), .B(sreg[1084]), .Z(n308) );
  OR U375 ( .A(n306), .B(n305), .Z(n307) );
  AND U376 ( .A(n308), .B(n307), .Z(n310) );
  XOR U377 ( .A(n311), .B(n310), .Z(c[1085]) );
  NAND U378 ( .A(b[0]), .B(a[63]), .Z(n314) );
  XOR U379 ( .A(sreg[1086]), .B(n314), .Z(n316) );
  NANDN U380 ( .A(n309), .B(sreg[1085]), .Z(n313) );
  OR U381 ( .A(n311), .B(n310), .Z(n312) );
  AND U382 ( .A(n313), .B(n312), .Z(n315) );
  XOR U383 ( .A(n316), .B(n315), .Z(c[1086]) );
  NAND U384 ( .A(b[0]), .B(a[64]), .Z(n319) );
  XOR U385 ( .A(sreg[1087]), .B(n319), .Z(n321) );
  NANDN U386 ( .A(n314), .B(sreg[1086]), .Z(n318) );
  OR U387 ( .A(n316), .B(n315), .Z(n317) );
  AND U388 ( .A(n318), .B(n317), .Z(n320) );
  XOR U389 ( .A(n321), .B(n320), .Z(c[1087]) );
  NAND U390 ( .A(b[0]), .B(a[65]), .Z(n324) );
  XOR U391 ( .A(sreg[1088]), .B(n324), .Z(n326) );
  NANDN U392 ( .A(n319), .B(sreg[1087]), .Z(n323) );
  OR U393 ( .A(n321), .B(n320), .Z(n322) );
  AND U394 ( .A(n323), .B(n322), .Z(n325) );
  XOR U395 ( .A(n326), .B(n325), .Z(c[1088]) );
  NAND U396 ( .A(b[0]), .B(a[66]), .Z(n329) );
  XOR U397 ( .A(sreg[1089]), .B(n329), .Z(n331) );
  NANDN U398 ( .A(n324), .B(sreg[1088]), .Z(n328) );
  OR U399 ( .A(n326), .B(n325), .Z(n327) );
  AND U400 ( .A(n328), .B(n327), .Z(n330) );
  XOR U401 ( .A(n331), .B(n330), .Z(c[1089]) );
  NAND U402 ( .A(b[0]), .B(a[67]), .Z(n334) );
  XOR U403 ( .A(sreg[1090]), .B(n334), .Z(n336) );
  NANDN U404 ( .A(n329), .B(sreg[1089]), .Z(n333) );
  OR U405 ( .A(n331), .B(n330), .Z(n332) );
  AND U406 ( .A(n333), .B(n332), .Z(n335) );
  XOR U407 ( .A(n336), .B(n335), .Z(c[1090]) );
  NAND U408 ( .A(b[0]), .B(a[68]), .Z(n339) );
  XOR U409 ( .A(sreg[1091]), .B(n339), .Z(n341) );
  NANDN U410 ( .A(n334), .B(sreg[1090]), .Z(n338) );
  OR U411 ( .A(n336), .B(n335), .Z(n337) );
  AND U412 ( .A(n338), .B(n337), .Z(n340) );
  XOR U413 ( .A(n341), .B(n340), .Z(c[1091]) );
  NAND U414 ( .A(b[0]), .B(a[69]), .Z(n344) );
  XOR U415 ( .A(sreg[1092]), .B(n344), .Z(n346) );
  NANDN U416 ( .A(n339), .B(sreg[1091]), .Z(n343) );
  OR U417 ( .A(n341), .B(n340), .Z(n342) );
  AND U418 ( .A(n343), .B(n342), .Z(n345) );
  XOR U419 ( .A(n346), .B(n345), .Z(c[1092]) );
  NAND U420 ( .A(b[0]), .B(a[70]), .Z(n349) );
  XOR U421 ( .A(sreg[1093]), .B(n349), .Z(n351) );
  NANDN U422 ( .A(n344), .B(sreg[1092]), .Z(n348) );
  OR U423 ( .A(n346), .B(n345), .Z(n347) );
  AND U424 ( .A(n348), .B(n347), .Z(n350) );
  XOR U425 ( .A(n351), .B(n350), .Z(c[1093]) );
  NAND U426 ( .A(b[0]), .B(a[71]), .Z(n354) );
  XOR U427 ( .A(sreg[1094]), .B(n354), .Z(n356) );
  NANDN U428 ( .A(n349), .B(sreg[1093]), .Z(n353) );
  OR U429 ( .A(n351), .B(n350), .Z(n352) );
  AND U430 ( .A(n353), .B(n352), .Z(n355) );
  XOR U431 ( .A(n356), .B(n355), .Z(c[1094]) );
  NAND U432 ( .A(b[0]), .B(a[72]), .Z(n359) );
  XOR U433 ( .A(sreg[1095]), .B(n359), .Z(n361) );
  NANDN U434 ( .A(n354), .B(sreg[1094]), .Z(n358) );
  OR U435 ( .A(n356), .B(n355), .Z(n357) );
  AND U436 ( .A(n358), .B(n357), .Z(n360) );
  XOR U437 ( .A(n361), .B(n360), .Z(c[1095]) );
  NAND U438 ( .A(b[0]), .B(a[73]), .Z(n364) );
  XOR U439 ( .A(sreg[1096]), .B(n364), .Z(n366) );
  NANDN U440 ( .A(n359), .B(sreg[1095]), .Z(n363) );
  OR U441 ( .A(n361), .B(n360), .Z(n362) );
  AND U442 ( .A(n363), .B(n362), .Z(n365) );
  XOR U443 ( .A(n366), .B(n365), .Z(c[1096]) );
  NAND U444 ( .A(b[0]), .B(a[74]), .Z(n369) );
  XOR U445 ( .A(sreg[1097]), .B(n369), .Z(n371) );
  NANDN U446 ( .A(n364), .B(sreg[1096]), .Z(n368) );
  OR U447 ( .A(n366), .B(n365), .Z(n367) );
  AND U448 ( .A(n368), .B(n367), .Z(n370) );
  XOR U449 ( .A(n371), .B(n370), .Z(c[1097]) );
  NAND U450 ( .A(b[0]), .B(a[75]), .Z(n374) );
  XOR U451 ( .A(sreg[1098]), .B(n374), .Z(n376) );
  NANDN U452 ( .A(n369), .B(sreg[1097]), .Z(n373) );
  OR U453 ( .A(n371), .B(n370), .Z(n372) );
  AND U454 ( .A(n373), .B(n372), .Z(n375) );
  XOR U455 ( .A(n376), .B(n375), .Z(c[1098]) );
  NAND U456 ( .A(b[0]), .B(a[76]), .Z(n379) );
  XOR U457 ( .A(sreg[1099]), .B(n379), .Z(n381) );
  NANDN U458 ( .A(n374), .B(sreg[1098]), .Z(n378) );
  OR U459 ( .A(n376), .B(n375), .Z(n377) );
  AND U460 ( .A(n378), .B(n377), .Z(n380) );
  XOR U461 ( .A(n381), .B(n380), .Z(c[1099]) );
  NAND U462 ( .A(b[0]), .B(a[77]), .Z(n384) );
  XOR U463 ( .A(sreg[1100]), .B(n384), .Z(n386) );
  NANDN U464 ( .A(n379), .B(sreg[1099]), .Z(n383) );
  OR U465 ( .A(n381), .B(n380), .Z(n382) );
  AND U466 ( .A(n383), .B(n382), .Z(n385) );
  XOR U467 ( .A(n386), .B(n385), .Z(c[1100]) );
  NAND U468 ( .A(b[0]), .B(a[78]), .Z(n389) );
  XOR U469 ( .A(sreg[1101]), .B(n389), .Z(n391) );
  NANDN U470 ( .A(n384), .B(sreg[1100]), .Z(n388) );
  OR U471 ( .A(n386), .B(n385), .Z(n387) );
  AND U472 ( .A(n388), .B(n387), .Z(n390) );
  XOR U473 ( .A(n391), .B(n390), .Z(c[1101]) );
  NAND U474 ( .A(b[0]), .B(a[79]), .Z(n394) );
  XOR U475 ( .A(sreg[1102]), .B(n394), .Z(n396) );
  NANDN U476 ( .A(n389), .B(sreg[1101]), .Z(n393) );
  OR U477 ( .A(n391), .B(n390), .Z(n392) );
  AND U478 ( .A(n393), .B(n392), .Z(n395) );
  XOR U479 ( .A(n396), .B(n395), .Z(c[1102]) );
  NAND U480 ( .A(b[0]), .B(a[80]), .Z(n399) );
  XOR U481 ( .A(sreg[1103]), .B(n399), .Z(n401) );
  NANDN U482 ( .A(n394), .B(sreg[1102]), .Z(n398) );
  OR U483 ( .A(n396), .B(n395), .Z(n397) );
  AND U484 ( .A(n398), .B(n397), .Z(n400) );
  XOR U485 ( .A(n401), .B(n400), .Z(c[1103]) );
  NAND U486 ( .A(b[0]), .B(a[81]), .Z(n404) );
  XOR U487 ( .A(sreg[1104]), .B(n404), .Z(n406) );
  NANDN U488 ( .A(n399), .B(sreg[1103]), .Z(n403) );
  OR U489 ( .A(n401), .B(n400), .Z(n402) );
  AND U490 ( .A(n403), .B(n402), .Z(n405) );
  XOR U491 ( .A(n406), .B(n405), .Z(c[1104]) );
  NAND U492 ( .A(b[0]), .B(a[82]), .Z(n409) );
  XOR U493 ( .A(sreg[1105]), .B(n409), .Z(n411) );
  NANDN U494 ( .A(n404), .B(sreg[1104]), .Z(n408) );
  OR U495 ( .A(n406), .B(n405), .Z(n407) );
  AND U496 ( .A(n408), .B(n407), .Z(n410) );
  XOR U497 ( .A(n411), .B(n410), .Z(c[1105]) );
  NAND U498 ( .A(b[0]), .B(a[83]), .Z(n414) );
  XOR U499 ( .A(sreg[1106]), .B(n414), .Z(n416) );
  NANDN U500 ( .A(n409), .B(sreg[1105]), .Z(n413) );
  OR U501 ( .A(n411), .B(n410), .Z(n412) );
  AND U502 ( .A(n413), .B(n412), .Z(n415) );
  XOR U503 ( .A(n416), .B(n415), .Z(c[1106]) );
  NAND U504 ( .A(b[0]), .B(a[84]), .Z(n419) );
  XOR U505 ( .A(sreg[1107]), .B(n419), .Z(n421) );
  NANDN U506 ( .A(n414), .B(sreg[1106]), .Z(n418) );
  OR U507 ( .A(n416), .B(n415), .Z(n417) );
  AND U508 ( .A(n418), .B(n417), .Z(n420) );
  XOR U509 ( .A(n421), .B(n420), .Z(c[1107]) );
  NAND U510 ( .A(b[0]), .B(a[85]), .Z(n424) );
  XOR U511 ( .A(sreg[1108]), .B(n424), .Z(n426) );
  NANDN U512 ( .A(n419), .B(sreg[1107]), .Z(n423) );
  OR U513 ( .A(n421), .B(n420), .Z(n422) );
  AND U514 ( .A(n423), .B(n422), .Z(n425) );
  XOR U515 ( .A(n426), .B(n425), .Z(c[1108]) );
  NAND U516 ( .A(b[0]), .B(a[86]), .Z(n429) );
  XOR U517 ( .A(sreg[1109]), .B(n429), .Z(n431) );
  NANDN U518 ( .A(n424), .B(sreg[1108]), .Z(n428) );
  OR U519 ( .A(n426), .B(n425), .Z(n427) );
  AND U520 ( .A(n428), .B(n427), .Z(n430) );
  XOR U521 ( .A(n431), .B(n430), .Z(c[1109]) );
  NAND U522 ( .A(b[0]), .B(a[87]), .Z(n434) );
  XOR U523 ( .A(sreg[1110]), .B(n434), .Z(n436) );
  NANDN U524 ( .A(n429), .B(sreg[1109]), .Z(n433) );
  OR U525 ( .A(n431), .B(n430), .Z(n432) );
  AND U526 ( .A(n433), .B(n432), .Z(n435) );
  XOR U527 ( .A(n436), .B(n435), .Z(c[1110]) );
  NAND U528 ( .A(b[0]), .B(a[88]), .Z(n439) );
  XOR U529 ( .A(sreg[1111]), .B(n439), .Z(n441) );
  NANDN U530 ( .A(n434), .B(sreg[1110]), .Z(n438) );
  OR U531 ( .A(n436), .B(n435), .Z(n437) );
  AND U532 ( .A(n438), .B(n437), .Z(n440) );
  XOR U533 ( .A(n441), .B(n440), .Z(c[1111]) );
  NAND U534 ( .A(b[0]), .B(a[89]), .Z(n444) );
  XOR U535 ( .A(sreg[1112]), .B(n444), .Z(n446) );
  NANDN U536 ( .A(n439), .B(sreg[1111]), .Z(n443) );
  OR U537 ( .A(n441), .B(n440), .Z(n442) );
  AND U538 ( .A(n443), .B(n442), .Z(n445) );
  XOR U539 ( .A(n446), .B(n445), .Z(c[1112]) );
  NAND U540 ( .A(b[0]), .B(a[90]), .Z(n449) );
  XOR U541 ( .A(sreg[1113]), .B(n449), .Z(n451) );
  NANDN U542 ( .A(n444), .B(sreg[1112]), .Z(n448) );
  OR U543 ( .A(n446), .B(n445), .Z(n447) );
  AND U544 ( .A(n448), .B(n447), .Z(n450) );
  XOR U545 ( .A(n451), .B(n450), .Z(c[1113]) );
  NAND U546 ( .A(b[0]), .B(a[91]), .Z(n454) );
  XOR U547 ( .A(sreg[1114]), .B(n454), .Z(n456) );
  NANDN U548 ( .A(n449), .B(sreg[1113]), .Z(n453) );
  OR U549 ( .A(n451), .B(n450), .Z(n452) );
  AND U550 ( .A(n453), .B(n452), .Z(n455) );
  XOR U551 ( .A(n456), .B(n455), .Z(c[1114]) );
  NAND U552 ( .A(b[0]), .B(a[92]), .Z(n459) );
  XOR U553 ( .A(sreg[1115]), .B(n459), .Z(n461) );
  NANDN U554 ( .A(n454), .B(sreg[1114]), .Z(n458) );
  OR U555 ( .A(n456), .B(n455), .Z(n457) );
  AND U556 ( .A(n458), .B(n457), .Z(n460) );
  XOR U557 ( .A(n461), .B(n460), .Z(c[1115]) );
  NAND U558 ( .A(b[0]), .B(a[93]), .Z(n464) );
  XOR U559 ( .A(sreg[1116]), .B(n464), .Z(n466) );
  NANDN U560 ( .A(n459), .B(sreg[1115]), .Z(n463) );
  OR U561 ( .A(n461), .B(n460), .Z(n462) );
  AND U562 ( .A(n463), .B(n462), .Z(n465) );
  XOR U563 ( .A(n466), .B(n465), .Z(c[1116]) );
  NAND U564 ( .A(b[0]), .B(a[94]), .Z(n469) );
  XOR U565 ( .A(sreg[1117]), .B(n469), .Z(n471) );
  NANDN U566 ( .A(n464), .B(sreg[1116]), .Z(n468) );
  OR U567 ( .A(n466), .B(n465), .Z(n467) );
  AND U568 ( .A(n468), .B(n467), .Z(n470) );
  XOR U569 ( .A(n471), .B(n470), .Z(c[1117]) );
  NAND U570 ( .A(b[0]), .B(a[95]), .Z(n474) );
  XOR U571 ( .A(sreg[1118]), .B(n474), .Z(n476) );
  NANDN U572 ( .A(n469), .B(sreg[1117]), .Z(n473) );
  OR U573 ( .A(n471), .B(n470), .Z(n472) );
  AND U574 ( .A(n473), .B(n472), .Z(n475) );
  XOR U575 ( .A(n476), .B(n475), .Z(c[1118]) );
  NAND U576 ( .A(b[0]), .B(a[96]), .Z(n479) );
  XOR U577 ( .A(sreg[1119]), .B(n479), .Z(n481) );
  NANDN U578 ( .A(n474), .B(sreg[1118]), .Z(n478) );
  OR U579 ( .A(n476), .B(n475), .Z(n477) );
  AND U580 ( .A(n478), .B(n477), .Z(n480) );
  XOR U581 ( .A(n481), .B(n480), .Z(c[1119]) );
  NAND U582 ( .A(b[0]), .B(a[97]), .Z(n484) );
  XOR U583 ( .A(sreg[1120]), .B(n484), .Z(n486) );
  NANDN U584 ( .A(n479), .B(sreg[1119]), .Z(n483) );
  OR U585 ( .A(n481), .B(n480), .Z(n482) );
  AND U586 ( .A(n483), .B(n482), .Z(n485) );
  XOR U587 ( .A(n486), .B(n485), .Z(c[1120]) );
  NAND U588 ( .A(b[0]), .B(a[98]), .Z(n489) );
  XOR U589 ( .A(sreg[1121]), .B(n489), .Z(n491) );
  NANDN U590 ( .A(n484), .B(sreg[1120]), .Z(n488) );
  OR U591 ( .A(n486), .B(n485), .Z(n487) );
  AND U592 ( .A(n488), .B(n487), .Z(n490) );
  XOR U593 ( .A(n491), .B(n490), .Z(c[1121]) );
  NAND U594 ( .A(b[0]), .B(a[99]), .Z(n494) );
  XOR U595 ( .A(sreg[1122]), .B(n494), .Z(n496) );
  NANDN U596 ( .A(n489), .B(sreg[1121]), .Z(n493) );
  OR U597 ( .A(n491), .B(n490), .Z(n492) );
  AND U598 ( .A(n493), .B(n492), .Z(n495) );
  XOR U599 ( .A(n496), .B(n495), .Z(c[1122]) );
  NAND U600 ( .A(b[0]), .B(a[100]), .Z(n499) );
  XOR U601 ( .A(sreg[1123]), .B(n499), .Z(n501) );
  NANDN U602 ( .A(n494), .B(sreg[1122]), .Z(n498) );
  OR U603 ( .A(n496), .B(n495), .Z(n497) );
  AND U604 ( .A(n498), .B(n497), .Z(n500) );
  XOR U605 ( .A(n501), .B(n500), .Z(c[1123]) );
  NAND U606 ( .A(b[0]), .B(a[101]), .Z(n504) );
  XOR U607 ( .A(sreg[1124]), .B(n504), .Z(n506) );
  NANDN U608 ( .A(n499), .B(sreg[1123]), .Z(n503) );
  OR U609 ( .A(n501), .B(n500), .Z(n502) );
  AND U610 ( .A(n503), .B(n502), .Z(n505) );
  XOR U611 ( .A(n506), .B(n505), .Z(c[1124]) );
  NAND U612 ( .A(b[0]), .B(a[102]), .Z(n509) );
  XOR U613 ( .A(sreg[1125]), .B(n509), .Z(n511) );
  NANDN U614 ( .A(n504), .B(sreg[1124]), .Z(n508) );
  OR U615 ( .A(n506), .B(n505), .Z(n507) );
  AND U616 ( .A(n508), .B(n507), .Z(n510) );
  XOR U617 ( .A(n511), .B(n510), .Z(c[1125]) );
  NAND U618 ( .A(b[0]), .B(a[103]), .Z(n514) );
  XOR U619 ( .A(sreg[1126]), .B(n514), .Z(n516) );
  NANDN U620 ( .A(n509), .B(sreg[1125]), .Z(n513) );
  OR U621 ( .A(n511), .B(n510), .Z(n512) );
  AND U622 ( .A(n513), .B(n512), .Z(n515) );
  XOR U623 ( .A(n516), .B(n515), .Z(c[1126]) );
  NAND U624 ( .A(b[0]), .B(a[104]), .Z(n519) );
  XOR U625 ( .A(sreg[1127]), .B(n519), .Z(n521) );
  NANDN U626 ( .A(n514), .B(sreg[1126]), .Z(n518) );
  OR U627 ( .A(n516), .B(n515), .Z(n517) );
  AND U628 ( .A(n518), .B(n517), .Z(n520) );
  XOR U629 ( .A(n521), .B(n520), .Z(c[1127]) );
  NAND U630 ( .A(b[0]), .B(a[105]), .Z(n524) );
  XOR U631 ( .A(sreg[1128]), .B(n524), .Z(n526) );
  NANDN U632 ( .A(n519), .B(sreg[1127]), .Z(n523) );
  OR U633 ( .A(n521), .B(n520), .Z(n522) );
  AND U634 ( .A(n523), .B(n522), .Z(n525) );
  XOR U635 ( .A(n526), .B(n525), .Z(c[1128]) );
  NAND U636 ( .A(b[0]), .B(a[106]), .Z(n529) );
  XOR U637 ( .A(sreg[1129]), .B(n529), .Z(n531) );
  NANDN U638 ( .A(n524), .B(sreg[1128]), .Z(n528) );
  OR U639 ( .A(n526), .B(n525), .Z(n527) );
  AND U640 ( .A(n528), .B(n527), .Z(n530) );
  XOR U641 ( .A(n531), .B(n530), .Z(c[1129]) );
  NAND U642 ( .A(b[0]), .B(a[107]), .Z(n534) );
  XOR U643 ( .A(sreg[1130]), .B(n534), .Z(n536) );
  NANDN U644 ( .A(n529), .B(sreg[1129]), .Z(n533) );
  OR U645 ( .A(n531), .B(n530), .Z(n532) );
  AND U646 ( .A(n533), .B(n532), .Z(n535) );
  XOR U647 ( .A(n536), .B(n535), .Z(c[1130]) );
  NAND U648 ( .A(b[0]), .B(a[108]), .Z(n539) );
  XOR U649 ( .A(sreg[1131]), .B(n539), .Z(n541) );
  NANDN U650 ( .A(n534), .B(sreg[1130]), .Z(n538) );
  OR U651 ( .A(n536), .B(n535), .Z(n537) );
  AND U652 ( .A(n538), .B(n537), .Z(n540) );
  XOR U653 ( .A(n541), .B(n540), .Z(c[1131]) );
  NAND U654 ( .A(b[0]), .B(a[109]), .Z(n544) );
  XOR U655 ( .A(sreg[1132]), .B(n544), .Z(n546) );
  NANDN U656 ( .A(n539), .B(sreg[1131]), .Z(n543) );
  OR U657 ( .A(n541), .B(n540), .Z(n542) );
  AND U658 ( .A(n543), .B(n542), .Z(n545) );
  XOR U659 ( .A(n546), .B(n545), .Z(c[1132]) );
  NAND U660 ( .A(b[0]), .B(a[110]), .Z(n549) );
  XOR U661 ( .A(sreg[1133]), .B(n549), .Z(n551) );
  NANDN U662 ( .A(n544), .B(sreg[1132]), .Z(n548) );
  OR U663 ( .A(n546), .B(n545), .Z(n547) );
  AND U664 ( .A(n548), .B(n547), .Z(n550) );
  XOR U665 ( .A(n551), .B(n550), .Z(c[1133]) );
  NAND U666 ( .A(b[0]), .B(a[111]), .Z(n554) );
  XOR U667 ( .A(sreg[1134]), .B(n554), .Z(n556) );
  NANDN U668 ( .A(n549), .B(sreg[1133]), .Z(n553) );
  OR U669 ( .A(n551), .B(n550), .Z(n552) );
  AND U670 ( .A(n553), .B(n552), .Z(n555) );
  XOR U671 ( .A(n556), .B(n555), .Z(c[1134]) );
  NAND U672 ( .A(b[0]), .B(a[112]), .Z(n559) );
  XOR U673 ( .A(sreg[1135]), .B(n559), .Z(n561) );
  NANDN U674 ( .A(n554), .B(sreg[1134]), .Z(n558) );
  OR U675 ( .A(n556), .B(n555), .Z(n557) );
  AND U676 ( .A(n558), .B(n557), .Z(n560) );
  XOR U677 ( .A(n561), .B(n560), .Z(c[1135]) );
  NAND U678 ( .A(b[0]), .B(a[113]), .Z(n564) );
  XOR U679 ( .A(sreg[1136]), .B(n564), .Z(n566) );
  NANDN U680 ( .A(n559), .B(sreg[1135]), .Z(n563) );
  OR U681 ( .A(n561), .B(n560), .Z(n562) );
  AND U682 ( .A(n563), .B(n562), .Z(n565) );
  XOR U683 ( .A(n566), .B(n565), .Z(c[1136]) );
  NAND U684 ( .A(b[0]), .B(a[114]), .Z(n569) );
  XOR U685 ( .A(sreg[1137]), .B(n569), .Z(n571) );
  NANDN U686 ( .A(n564), .B(sreg[1136]), .Z(n568) );
  OR U687 ( .A(n566), .B(n565), .Z(n567) );
  AND U688 ( .A(n568), .B(n567), .Z(n570) );
  XOR U689 ( .A(n571), .B(n570), .Z(c[1137]) );
  NAND U690 ( .A(b[0]), .B(a[115]), .Z(n574) );
  XOR U691 ( .A(sreg[1138]), .B(n574), .Z(n576) );
  NANDN U692 ( .A(n569), .B(sreg[1137]), .Z(n573) );
  OR U693 ( .A(n571), .B(n570), .Z(n572) );
  AND U694 ( .A(n573), .B(n572), .Z(n575) );
  XOR U695 ( .A(n576), .B(n575), .Z(c[1138]) );
  NAND U696 ( .A(b[0]), .B(a[116]), .Z(n579) );
  XOR U697 ( .A(sreg[1139]), .B(n579), .Z(n581) );
  NANDN U698 ( .A(n574), .B(sreg[1138]), .Z(n578) );
  OR U699 ( .A(n576), .B(n575), .Z(n577) );
  AND U700 ( .A(n578), .B(n577), .Z(n580) );
  XOR U701 ( .A(n581), .B(n580), .Z(c[1139]) );
  NAND U702 ( .A(b[0]), .B(a[117]), .Z(n584) );
  XOR U703 ( .A(sreg[1140]), .B(n584), .Z(n586) );
  NANDN U704 ( .A(n579), .B(sreg[1139]), .Z(n583) );
  OR U705 ( .A(n581), .B(n580), .Z(n582) );
  AND U706 ( .A(n583), .B(n582), .Z(n585) );
  XOR U707 ( .A(n586), .B(n585), .Z(c[1140]) );
  NAND U708 ( .A(b[0]), .B(a[118]), .Z(n589) );
  XOR U709 ( .A(sreg[1141]), .B(n589), .Z(n591) );
  NANDN U710 ( .A(n584), .B(sreg[1140]), .Z(n588) );
  OR U711 ( .A(n586), .B(n585), .Z(n587) );
  AND U712 ( .A(n588), .B(n587), .Z(n590) );
  XOR U713 ( .A(n591), .B(n590), .Z(c[1141]) );
  NAND U714 ( .A(b[0]), .B(a[119]), .Z(n594) );
  XOR U715 ( .A(sreg[1142]), .B(n594), .Z(n596) );
  NANDN U716 ( .A(n589), .B(sreg[1141]), .Z(n593) );
  OR U717 ( .A(n591), .B(n590), .Z(n592) );
  AND U718 ( .A(n593), .B(n592), .Z(n595) );
  XOR U719 ( .A(n596), .B(n595), .Z(c[1142]) );
  NAND U720 ( .A(b[0]), .B(a[120]), .Z(n599) );
  XOR U721 ( .A(sreg[1143]), .B(n599), .Z(n601) );
  NANDN U722 ( .A(n594), .B(sreg[1142]), .Z(n598) );
  OR U723 ( .A(n596), .B(n595), .Z(n597) );
  AND U724 ( .A(n598), .B(n597), .Z(n600) );
  XOR U725 ( .A(n601), .B(n600), .Z(c[1143]) );
  NAND U726 ( .A(b[0]), .B(a[121]), .Z(n604) );
  XOR U727 ( .A(sreg[1144]), .B(n604), .Z(n606) );
  NANDN U728 ( .A(n599), .B(sreg[1143]), .Z(n603) );
  OR U729 ( .A(n601), .B(n600), .Z(n602) );
  AND U730 ( .A(n603), .B(n602), .Z(n605) );
  XOR U731 ( .A(n606), .B(n605), .Z(c[1144]) );
  NAND U732 ( .A(b[0]), .B(a[122]), .Z(n609) );
  XOR U733 ( .A(sreg[1145]), .B(n609), .Z(n611) );
  NANDN U734 ( .A(n604), .B(sreg[1144]), .Z(n608) );
  OR U735 ( .A(n606), .B(n605), .Z(n607) );
  AND U736 ( .A(n608), .B(n607), .Z(n610) );
  XOR U737 ( .A(n611), .B(n610), .Z(c[1145]) );
  NAND U738 ( .A(b[0]), .B(a[123]), .Z(n614) );
  XOR U739 ( .A(sreg[1146]), .B(n614), .Z(n616) );
  NANDN U740 ( .A(n609), .B(sreg[1145]), .Z(n613) );
  OR U741 ( .A(n611), .B(n610), .Z(n612) );
  AND U742 ( .A(n613), .B(n612), .Z(n615) );
  XOR U743 ( .A(n616), .B(n615), .Z(c[1146]) );
  NAND U744 ( .A(b[0]), .B(a[124]), .Z(n619) );
  XOR U745 ( .A(sreg[1147]), .B(n619), .Z(n621) );
  NANDN U746 ( .A(n614), .B(sreg[1146]), .Z(n618) );
  OR U747 ( .A(n616), .B(n615), .Z(n617) );
  AND U748 ( .A(n618), .B(n617), .Z(n620) );
  XOR U749 ( .A(n621), .B(n620), .Z(c[1147]) );
  NAND U750 ( .A(b[0]), .B(a[125]), .Z(n624) );
  XOR U751 ( .A(sreg[1148]), .B(n624), .Z(n626) );
  NANDN U752 ( .A(n619), .B(sreg[1147]), .Z(n623) );
  OR U753 ( .A(n621), .B(n620), .Z(n622) );
  AND U754 ( .A(n623), .B(n622), .Z(n625) );
  XOR U755 ( .A(n626), .B(n625), .Z(c[1148]) );
  NAND U756 ( .A(b[0]), .B(a[126]), .Z(n629) );
  XOR U757 ( .A(sreg[1149]), .B(n629), .Z(n631) );
  NANDN U758 ( .A(n624), .B(sreg[1148]), .Z(n628) );
  OR U759 ( .A(n626), .B(n625), .Z(n627) );
  AND U760 ( .A(n628), .B(n627), .Z(n630) );
  XOR U761 ( .A(n631), .B(n630), .Z(c[1149]) );
  NAND U762 ( .A(b[0]), .B(a[127]), .Z(n634) );
  XOR U763 ( .A(sreg[1150]), .B(n634), .Z(n636) );
  NANDN U764 ( .A(n629), .B(sreg[1149]), .Z(n633) );
  OR U765 ( .A(n631), .B(n630), .Z(n632) );
  AND U766 ( .A(n633), .B(n632), .Z(n635) );
  XOR U767 ( .A(n636), .B(n635), .Z(c[1150]) );
  NAND U768 ( .A(b[0]), .B(a[128]), .Z(n639) );
  XOR U769 ( .A(sreg[1151]), .B(n639), .Z(n641) );
  NANDN U770 ( .A(n634), .B(sreg[1150]), .Z(n638) );
  OR U771 ( .A(n636), .B(n635), .Z(n637) );
  AND U772 ( .A(n638), .B(n637), .Z(n640) );
  XOR U773 ( .A(n641), .B(n640), .Z(c[1151]) );
  NAND U774 ( .A(b[0]), .B(a[129]), .Z(n644) );
  XOR U775 ( .A(sreg[1152]), .B(n644), .Z(n646) );
  NANDN U776 ( .A(n639), .B(sreg[1151]), .Z(n643) );
  OR U777 ( .A(n641), .B(n640), .Z(n642) );
  AND U778 ( .A(n643), .B(n642), .Z(n645) );
  XOR U779 ( .A(n646), .B(n645), .Z(c[1152]) );
  NAND U780 ( .A(b[0]), .B(a[130]), .Z(n649) );
  XOR U781 ( .A(sreg[1153]), .B(n649), .Z(n651) );
  NANDN U782 ( .A(n644), .B(sreg[1152]), .Z(n648) );
  OR U783 ( .A(n646), .B(n645), .Z(n647) );
  AND U784 ( .A(n648), .B(n647), .Z(n650) );
  XOR U785 ( .A(n651), .B(n650), .Z(c[1153]) );
  NAND U786 ( .A(b[0]), .B(a[131]), .Z(n654) );
  XOR U787 ( .A(sreg[1154]), .B(n654), .Z(n656) );
  NANDN U788 ( .A(n649), .B(sreg[1153]), .Z(n653) );
  OR U789 ( .A(n651), .B(n650), .Z(n652) );
  AND U790 ( .A(n653), .B(n652), .Z(n655) );
  XOR U791 ( .A(n656), .B(n655), .Z(c[1154]) );
  NAND U792 ( .A(b[0]), .B(a[132]), .Z(n659) );
  XOR U793 ( .A(sreg[1155]), .B(n659), .Z(n661) );
  NANDN U794 ( .A(n654), .B(sreg[1154]), .Z(n658) );
  OR U795 ( .A(n656), .B(n655), .Z(n657) );
  AND U796 ( .A(n658), .B(n657), .Z(n660) );
  XOR U797 ( .A(n661), .B(n660), .Z(c[1155]) );
  NAND U798 ( .A(b[0]), .B(a[133]), .Z(n664) );
  XOR U799 ( .A(sreg[1156]), .B(n664), .Z(n666) );
  NANDN U800 ( .A(n659), .B(sreg[1155]), .Z(n663) );
  OR U801 ( .A(n661), .B(n660), .Z(n662) );
  AND U802 ( .A(n663), .B(n662), .Z(n665) );
  XOR U803 ( .A(n666), .B(n665), .Z(c[1156]) );
  NAND U804 ( .A(b[0]), .B(a[134]), .Z(n669) );
  XOR U805 ( .A(sreg[1157]), .B(n669), .Z(n671) );
  NANDN U806 ( .A(n664), .B(sreg[1156]), .Z(n668) );
  OR U807 ( .A(n666), .B(n665), .Z(n667) );
  AND U808 ( .A(n668), .B(n667), .Z(n670) );
  XOR U809 ( .A(n671), .B(n670), .Z(c[1157]) );
  NAND U810 ( .A(b[0]), .B(a[135]), .Z(n674) );
  XOR U811 ( .A(sreg[1158]), .B(n674), .Z(n676) );
  NANDN U812 ( .A(n669), .B(sreg[1157]), .Z(n673) );
  OR U813 ( .A(n671), .B(n670), .Z(n672) );
  AND U814 ( .A(n673), .B(n672), .Z(n675) );
  XOR U815 ( .A(n676), .B(n675), .Z(c[1158]) );
  NAND U816 ( .A(b[0]), .B(a[136]), .Z(n679) );
  XOR U817 ( .A(sreg[1159]), .B(n679), .Z(n681) );
  NANDN U818 ( .A(n674), .B(sreg[1158]), .Z(n678) );
  OR U819 ( .A(n676), .B(n675), .Z(n677) );
  AND U820 ( .A(n678), .B(n677), .Z(n680) );
  XOR U821 ( .A(n681), .B(n680), .Z(c[1159]) );
  NAND U822 ( .A(b[0]), .B(a[137]), .Z(n684) );
  XOR U823 ( .A(sreg[1160]), .B(n684), .Z(n686) );
  NANDN U824 ( .A(n679), .B(sreg[1159]), .Z(n683) );
  OR U825 ( .A(n681), .B(n680), .Z(n682) );
  AND U826 ( .A(n683), .B(n682), .Z(n685) );
  XOR U827 ( .A(n686), .B(n685), .Z(c[1160]) );
  NAND U828 ( .A(b[0]), .B(a[138]), .Z(n689) );
  XOR U829 ( .A(sreg[1161]), .B(n689), .Z(n691) );
  NANDN U830 ( .A(n684), .B(sreg[1160]), .Z(n688) );
  OR U831 ( .A(n686), .B(n685), .Z(n687) );
  AND U832 ( .A(n688), .B(n687), .Z(n690) );
  XOR U833 ( .A(n691), .B(n690), .Z(c[1161]) );
  NAND U834 ( .A(b[0]), .B(a[139]), .Z(n694) );
  XOR U835 ( .A(sreg[1162]), .B(n694), .Z(n696) );
  NANDN U836 ( .A(n689), .B(sreg[1161]), .Z(n693) );
  OR U837 ( .A(n691), .B(n690), .Z(n692) );
  AND U838 ( .A(n693), .B(n692), .Z(n695) );
  XOR U839 ( .A(n696), .B(n695), .Z(c[1162]) );
  NAND U840 ( .A(b[0]), .B(a[140]), .Z(n699) );
  XOR U841 ( .A(sreg[1163]), .B(n699), .Z(n701) );
  NANDN U842 ( .A(n694), .B(sreg[1162]), .Z(n698) );
  OR U843 ( .A(n696), .B(n695), .Z(n697) );
  AND U844 ( .A(n698), .B(n697), .Z(n700) );
  XOR U845 ( .A(n701), .B(n700), .Z(c[1163]) );
  NAND U846 ( .A(b[0]), .B(a[141]), .Z(n704) );
  XOR U847 ( .A(sreg[1164]), .B(n704), .Z(n706) );
  NANDN U848 ( .A(n699), .B(sreg[1163]), .Z(n703) );
  OR U849 ( .A(n701), .B(n700), .Z(n702) );
  AND U850 ( .A(n703), .B(n702), .Z(n705) );
  XOR U851 ( .A(n706), .B(n705), .Z(c[1164]) );
  NAND U852 ( .A(b[0]), .B(a[142]), .Z(n709) );
  XOR U853 ( .A(sreg[1165]), .B(n709), .Z(n711) );
  NANDN U854 ( .A(n704), .B(sreg[1164]), .Z(n708) );
  OR U855 ( .A(n706), .B(n705), .Z(n707) );
  AND U856 ( .A(n708), .B(n707), .Z(n710) );
  XOR U857 ( .A(n711), .B(n710), .Z(c[1165]) );
  NAND U858 ( .A(b[0]), .B(a[143]), .Z(n714) );
  XOR U859 ( .A(sreg[1166]), .B(n714), .Z(n716) );
  NANDN U860 ( .A(n709), .B(sreg[1165]), .Z(n713) );
  OR U861 ( .A(n711), .B(n710), .Z(n712) );
  AND U862 ( .A(n713), .B(n712), .Z(n715) );
  XOR U863 ( .A(n716), .B(n715), .Z(c[1166]) );
  NAND U864 ( .A(b[0]), .B(a[144]), .Z(n719) );
  XOR U865 ( .A(sreg[1167]), .B(n719), .Z(n721) );
  NANDN U866 ( .A(n714), .B(sreg[1166]), .Z(n718) );
  OR U867 ( .A(n716), .B(n715), .Z(n717) );
  AND U868 ( .A(n718), .B(n717), .Z(n720) );
  XOR U869 ( .A(n721), .B(n720), .Z(c[1167]) );
  NAND U870 ( .A(b[0]), .B(a[145]), .Z(n724) );
  XOR U871 ( .A(sreg[1168]), .B(n724), .Z(n726) );
  NANDN U872 ( .A(n719), .B(sreg[1167]), .Z(n723) );
  OR U873 ( .A(n721), .B(n720), .Z(n722) );
  AND U874 ( .A(n723), .B(n722), .Z(n725) );
  XOR U875 ( .A(n726), .B(n725), .Z(c[1168]) );
  NAND U876 ( .A(b[0]), .B(a[146]), .Z(n729) );
  XOR U877 ( .A(sreg[1169]), .B(n729), .Z(n731) );
  NANDN U878 ( .A(n724), .B(sreg[1168]), .Z(n728) );
  OR U879 ( .A(n726), .B(n725), .Z(n727) );
  AND U880 ( .A(n728), .B(n727), .Z(n730) );
  XOR U881 ( .A(n731), .B(n730), .Z(c[1169]) );
  NAND U882 ( .A(b[0]), .B(a[147]), .Z(n734) );
  XOR U883 ( .A(sreg[1170]), .B(n734), .Z(n736) );
  NANDN U884 ( .A(n729), .B(sreg[1169]), .Z(n733) );
  OR U885 ( .A(n731), .B(n730), .Z(n732) );
  AND U886 ( .A(n733), .B(n732), .Z(n735) );
  XOR U887 ( .A(n736), .B(n735), .Z(c[1170]) );
  NAND U888 ( .A(b[0]), .B(a[148]), .Z(n739) );
  XOR U889 ( .A(sreg[1171]), .B(n739), .Z(n741) );
  NANDN U890 ( .A(n734), .B(sreg[1170]), .Z(n738) );
  OR U891 ( .A(n736), .B(n735), .Z(n737) );
  AND U892 ( .A(n738), .B(n737), .Z(n740) );
  XOR U893 ( .A(n741), .B(n740), .Z(c[1171]) );
  NAND U894 ( .A(b[0]), .B(a[149]), .Z(n744) );
  XOR U895 ( .A(sreg[1172]), .B(n744), .Z(n746) );
  NANDN U896 ( .A(n739), .B(sreg[1171]), .Z(n743) );
  OR U897 ( .A(n741), .B(n740), .Z(n742) );
  AND U898 ( .A(n743), .B(n742), .Z(n745) );
  XOR U899 ( .A(n746), .B(n745), .Z(c[1172]) );
  NAND U900 ( .A(b[0]), .B(a[150]), .Z(n749) );
  XOR U901 ( .A(sreg[1173]), .B(n749), .Z(n751) );
  NANDN U902 ( .A(n744), .B(sreg[1172]), .Z(n748) );
  OR U903 ( .A(n746), .B(n745), .Z(n747) );
  AND U904 ( .A(n748), .B(n747), .Z(n750) );
  XOR U905 ( .A(n751), .B(n750), .Z(c[1173]) );
  NAND U906 ( .A(b[0]), .B(a[151]), .Z(n754) );
  XOR U907 ( .A(sreg[1174]), .B(n754), .Z(n756) );
  NANDN U908 ( .A(n749), .B(sreg[1173]), .Z(n753) );
  OR U909 ( .A(n751), .B(n750), .Z(n752) );
  AND U910 ( .A(n753), .B(n752), .Z(n755) );
  XOR U911 ( .A(n756), .B(n755), .Z(c[1174]) );
  NAND U912 ( .A(b[0]), .B(a[152]), .Z(n759) );
  XOR U913 ( .A(sreg[1175]), .B(n759), .Z(n761) );
  NANDN U914 ( .A(n754), .B(sreg[1174]), .Z(n758) );
  OR U915 ( .A(n756), .B(n755), .Z(n757) );
  AND U916 ( .A(n758), .B(n757), .Z(n760) );
  XOR U917 ( .A(n761), .B(n760), .Z(c[1175]) );
  NAND U918 ( .A(b[0]), .B(a[153]), .Z(n764) );
  XOR U919 ( .A(sreg[1176]), .B(n764), .Z(n766) );
  NANDN U920 ( .A(n759), .B(sreg[1175]), .Z(n763) );
  OR U921 ( .A(n761), .B(n760), .Z(n762) );
  AND U922 ( .A(n763), .B(n762), .Z(n765) );
  XOR U923 ( .A(n766), .B(n765), .Z(c[1176]) );
  NAND U924 ( .A(b[0]), .B(a[154]), .Z(n769) );
  XOR U925 ( .A(sreg[1177]), .B(n769), .Z(n771) );
  NANDN U926 ( .A(n764), .B(sreg[1176]), .Z(n768) );
  OR U927 ( .A(n766), .B(n765), .Z(n767) );
  AND U928 ( .A(n768), .B(n767), .Z(n770) );
  XOR U929 ( .A(n771), .B(n770), .Z(c[1177]) );
  NAND U930 ( .A(b[0]), .B(a[155]), .Z(n774) );
  XOR U931 ( .A(sreg[1178]), .B(n774), .Z(n776) );
  NANDN U932 ( .A(n769), .B(sreg[1177]), .Z(n773) );
  OR U933 ( .A(n771), .B(n770), .Z(n772) );
  AND U934 ( .A(n773), .B(n772), .Z(n775) );
  XOR U935 ( .A(n776), .B(n775), .Z(c[1178]) );
  NAND U936 ( .A(b[0]), .B(a[156]), .Z(n779) );
  XOR U937 ( .A(sreg[1179]), .B(n779), .Z(n781) );
  NANDN U938 ( .A(n774), .B(sreg[1178]), .Z(n778) );
  OR U939 ( .A(n776), .B(n775), .Z(n777) );
  AND U940 ( .A(n778), .B(n777), .Z(n780) );
  XOR U941 ( .A(n781), .B(n780), .Z(c[1179]) );
  NAND U942 ( .A(b[0]), .B(a[157]), .Z(n784) );
  XOR U943 ( .A(sreg[1180]), .B(n784), .Z(n786) );
  NANDN U944 ( .A(n779), .B(sreg[1179]), .Z(n783) );
  OR U945 ( .A(n781), .B(n780), .Z(n782) );
  AND U946 ( .A(n783), .B(n782), .Z(n785) );
  XOR U947 ( .A(n786), .B(n785), .Z(c[1180]) );
  NAND U948 ( .A(b[0]), .B(a[158]), .Z(n789) );
  XOR U949 ( .A(sreg[1181]), .B(n789), .Z(n791) );
  NANDN U950 ( .A(n784), .B(sreg[1180]), .Z(n788) );
  OR U951 ( .A(n786), .B(n785), .Z(n787) );
  AND U952 ( .A(n788), .B(n787), .Z(n790) );
  XOR U953 ( .A(n791), .B(n790), .Z(c[1181]) );
  NAND U954 ( .A(b[0]), .B(a[159]), .Z(n794) );
  XOR U955 ( .A(sreg[1182]), .B(n794), .Z(n796) );
  NANDN U956 ( .A(n789), .B(sreg[1181]), .Z(n793) );
  OR U957 ( .A(n791), .B(n790), .Z(n792) );
  AND U958 ( .A(n793), .B(n792), .Z(n795) );
  XOR U959 ( .A(n796), .B(n795), .Z(c[1182]) );
  NAND U960 ( .A(b[0]), .B(a[160]), .Z(n799) );
  XOR U961 ( .A(sreg[1183]), .B(n799), .Z(n801) );
  NANDN U962 ( .A(n794), .B(sreg[1182]), .Z(n798) );
  OR U963 ( .A(n796), .B(n795), .Z(n797) );
  AND U964 ( .A(n798), .B(n797), .Z(n800) );
  XOR U965 ( .A(n801), .B(n800), .Z(c[1183]) );
  NAND U966 ( .A(b[0]), .B(a[161]), .Z(n804) );
  XOR U967 ( .A(sreg[1184]), .B(n804), .Z(n806) );
  NANDN U968 ( .A(n799), .B(sreg[1183]), .Z(n803) );
  OR U969 ( .A(n801), .B(n800), .Z(n802) );
  AND U970 ( .A(n803), .B(n802), .Z(n805) );
  XOR U971 ( .A(n806), .B(n805), .Z(c[1184]) );
  NAND U972 ( .A(b[0]), .B(a[162]), .Z(n809) );
  XOR U973 ( .A(sreg[1185]), .B(n809), .Z(n811) );
  NANDN U974 ( .A(n804), .B(sreg[1184]), .Z(n808) );
  OR U975 ( .A(n806), .B(n805), .Z(n807) );
  AND U976 ( .A(n808), .B(n807), .Z(n810) );
  XOR U977 ( .A(n811), .B(n810), .Z(c[1185]) );
  NAND U978 ( .A(b[0]), .B(a[163]), .Z(n814) );
  XOR U979 ( .A(sreg[1186]), .B(n814), .Z(n816) );
  NANDN U980 ( .A(n809), .B(sreg[1185]), .Z(n813) );
  OR U981 ( .A(n811), .B(n810), .Z(n812) );
  AND U982 ( .A(n813), .B(n812), .Z(n815) );
  XOR U983 ( .A(n816), .B(n815), .Z(c[1186]) );
  NAND U984 ( .A(b[0]), .B(a[164]), .Z(n819) );
  XOR U985 ( .A(sreg[1187]), .B(n819), .Z(n821) );
  NANDN U986 ( .A(n814), .B(sreg[1186]), .Z(n818) );
  OR U987 ( .A(n816), .B(n815), .Z(n817) );
  AND U988 ( .A(n818), .B(n817), .Z(n820) );
  XOR U989 ( .A(n821), .B(n820), .Z(c[1187]) );
  NAND U990 ( .A(b[0]), .B(a[165]), .Z(n824) );
  XOR U991 ( .A(sreg[1188]), .B(n824), .Z(n826) );
  NANDN U992 ( .A(n819), .B(sreg[1187]), .Z(n823) );
  OR U993 ( .A(n821), .B(n820), .Z(n822) );
  AND U994 ( .A(n823), .B(n822), .Z(n825) );
  XOR U995 ( .A(n826), .B(n825), .Z(c[1188]) );
  NAND U996 ( .A(b[0]), .B(a[166]), .Z(n829) );
  XOR U997 ( .A(sreg[1189]), .B(n829), .Z(n831) );
  NANDN U998 ( .A(n824), .B(sreg[1188]), .Z(n828) );
  OR U999 ( .A(n826), .B(n825), .Z(n827) );
  AND U1000 ( .A(n828), .B(n827), .Z(n830) );
  XOR U1001 ( .A(n831), .B(n830), .Z(c[1189]) );
  NAND U1002 ( .A(b[0]), .B(a[167]), .Z(n834) );
  XOR U1003 ( .A(sreg[1190]), .B(n834), .Z(n836) );
  NANDN U1004 ( .A(n829), .B(sreg[1189]), .Z(n833) );
  OR U1005 ( .A(n831), .B(n830), .Z(n832) );
  AND U1006 ( .A(n833), .B(n832), .Z(n835) );
  XOR U1007 ( .A(n836), .B(n835), .Z(c[1190]) );
  NAND U1008 ( .A(b[0]), .B(a[168]), .Z(n839) );
  XOR U1009 ( .A(sreg[1191]), .B(n839), .Z(n841) );
  NANDN U1010 ( .A(n834), .B(sreg[1190]), .Z(n838) );
  OR U1011 ( .A(n836), .B(n835), .Z(n837) );
  AND U1012 ( .A(n838), .B(n837), .Z(n840) );
  XOR U1013 ( .A(n841), .B(n840), .Z(c[1191]) );
  NAND U1014 ( .A(b[0]), .B(a[169]), .Z(n844) );
  XOR U1015 ( .A(sreg[1192]), .B(n844), .Z(n846) );
  NANDN U1016 ( .A(n839), .B(sreg[1191]), .Z(n843) );
  OR U1017 ( .A(n841), .B(n840), .Z(n842) );
  AND U1018 ( .A(n843), .B(n842), .Z(n845) );
  XOR U1019 ( .A(n846), .B(n845), .Z(c[1192]) );
  NAND U1020 ( .A(b[0]), .B(a[170]), .Z(n849) );
  XOR U1021 ( .A(sreg[1193]), .B(n849), .Z(n851) );
  NANDN U1022 ( .A(n844), .B(sreg[1192]), .Z(n848) );
  OR U1023 ( .A(n846), .B(n845), .Z(n847) );
  AND U1024 ( .A(n848), .B(n847), .Z(n850) );
  XOR U1025 ( .A(n851), .B(n850), .Z(c[1193]) );
  NAND U1026 ( .A(b[0]), .B(a[171]), .Z(n854) );
  XOR U1027 ( .A(sreg[1194]), .B(n854), .Z(n856) );
  NANDN U1028 ( .A(n849), .B(sreg[1193]), .Z(n853) );
  OR U1029 ( .A(n851), .B(n850), .Z(n852) );
  AND U1030 ( .A(n853), .B(n852), .Z(n855) );
  XOR U1031 ( .A(n856), .B(n855), .Z(c[1194]) );
  NAND U1032 ( .A(b[0]), .B(a[172]), .Z(n859) );
  XOR U1033 ( .A(sreg[1195]), .B(n859), .Z(n861) );
  NANDN U1034 ( .A(n854), .B(sreg[1194]), .Z(n858) );
  OR U1035 ( .A(n856), .B(n855), .Z(n857) );
  AND U1036 ( .A(n858), .B(n857), .Z(n860) );
  XOR U1037 ( .A(n861), .B(n860), .Z(c[1195]) );
  NAND U1038 ( .A(b[0]), .B(a[173]), .Z(n864) );
  XOR U1039 ( .A(sreg[1196]), .B(n864), .Z(n866) );
  NANDN U1040 ( .A(n859), .B(sreg[1195]), .Z(n863) );
  OR U1041 ( .A(n861), .B(n860), .Z(n862) );
  AND U1042 ( .A(n863), .B(n862), .Z(n865) );
  XOR U1043 ( .A(n866), .B(n865), .Z(c[1196]) );
  NAND U1044 ( .A(b[0]), .B(a[174]), .Z(n869) );
  XOR U1045 ( .A(sreg[1197]), .B(n869), .Z(n871) );
  NANDN U1046 ( .A(n864), .B(sreg[1196]), .Z(n868) );
  OR U1047 ( .A(n866), .B(n865), .Z(n867) );
  AND U1048 ( .A(n868), .B(n867), .Z(n870) );
  XOR U1049 ( .A(n871), .B(n870), .Z(c[1197]) );
  NAND U1050 ( .A(b[0]), .B(a[175]), .Z(n874) );
  XOR U1051 ( .A(sreg[1198]), .B(n874), .Z(n876) );
  NANDN U1052 ( .A(n869), .B(sreg[1197]), .Z(n873) );
  OR U1053 ( .A(n871), .B(n870), .Z(n872) );
  AND U1054 ( .A(n873), .B(n872), .Z(n875) );
  XOR U1055 ( .A(n876), .B(n875), .Z(c[1198]) );
  NAND U1056 ( .A(b[0]), .B(a[176]), .Z(n879) );
  XOR U1057 ( .A(sreg[1199]), .B(n879), .Z(n881) );
  NANDN U1058 ( .A(n874), .B(sreg[1198]), .Z(n878) );
  OR U1059 ( .A(n876), .B(n875), .Z(n877) );
  AND U1060 ( .A(n878), .B(n877), .Z(n880) );
  XOR U1061 ( .A(n881), .B(n880), .Z(c[1199]) );
  NAND U1062 ( .A(b[0]), .B(a[177]), .Z(n884) );
  XOR U1063 ( .A(sreg[1200]), .B(n884), .Z(n886) );
  NANDN U1064 ( .A(n879), .B(sreg[1199]), .Z(n883) );
  OR U1065 ( .A(n881), .B(n880), .Z(n882) );
  AND U1066 ( .A(n883), .B(n882), .Z(n885) );
  XOR U1067 ( .A(n886), .B(n885), .Z(c[1200]) );
  NAND U1068 ( .A(b[0]), .B(a[178]), .Z(n889) );
  XOR U1069 ( .A(sreg[1201]), .B(n889), .Z(n891) );
  NANDN U1070 ( .A(n884), .B(sreg[1200]), .Z(n888) );
  OR U1071 ( .A(n886), .B(n885), .Z(n887) );
  AND U1072 ( .A(n888), .B(n887), .Z(n890) );
  XOR U1073 ( .A(n891), .B(n890), .Z(c[1201]) );
  NAND U1074 ( .A(b[0]), .B(a[179]), .Z(n894) );
  XOR U1075 ( .A(sreg[1202]), .B(n894), .Z(n896) );
  NANDN U1076 ( .A(n889), .B(sreg[1201]), .Z(n893) );
  OR U1077 ( .A(n891), .B(n890), .Z(n892) );
  AND U1078 ( .A(n893), .B(n892), .Z(n895) );
  XOR U1079 ( .A(n896), .B(n895), .Z(c[1202]) );
  NAND U1080 ( .A(b[0]), .B(a[180]), .Z(n899) );
  XOR U1081 ( .A(sreg[1203]), .B(n899), .Z(n901) );
  NANDN U1082 ( .A(n894), .B(sreg[1202]), .Z(n898) );
  OR U1083 ( .A(n896), .B(n895), .Z(n897) );
  AND U1084 ( .A(n898), .B(n897), .Z(n900) );
  XOR U1085 ( .A(n901), .B(n900), .Z(c[1203]) );
  NAND U1086 ( .A(b[0]), .B(a[181]), .Z(n904) );
  XOR U1087 ( .A(sreg[1204]), .B(n904), .Z(n906) );
  NANDN U1088 ( .A(n899), .B(sreg[1203]), .Z(n903) );
  OR U1089 ( .A(n901), .B(n900), .Z(n902) );
  AND U1090 ( .A(n903), .B(n902), .Z(n905) );
  XOR U1091 ( .A(n906), .B(n905), .Z(c[1204]) );
  NAND U1092 ( .A(b[0]), .B(a[182]), .Z(n909) );
  XOR U1093 ( .A(sreg[1205]), .B(n909), .Z(n911) );
  NANDN U1094 ( .A(n904), .B(sreg[1204]), .Z(n908) );
  OR U1095 ( .A(n906), .B(n905), .Z(n907) );
  AND U1096 ( .A(n908), .B(n907), .Z(n910) );
  XOR U1097 ( .A(n911), .B(n910), .Z(c[1205]) );
  NAND U1098 ( .A(b[0]), .B(a[183]), .Z(n914) );
  XOR U1099 ( .A(sreg[1206]), .B(n914), .Z(n916) );
  NANDN U1100 ( .A(n909), .B(sreg[1205]), .Z(n913) );
  OR U1101 ( .A(n911), .B(n910), .Z(n912) );
  AND U1102 ( .A(n913), .B(n912), .Z(n915) );
  XOR U1103 ( .A(n916), .B(n915), .Z(c[1206]) );
  NAND U1104 ( .A(b[0]), .B(a[184]), .Z(n919) );
  XOR U1105 ( .A(sreg[1207]), .B(n919), .Z(n921) );
  NANDN U1106 ( .A(n914), .B(sreg[1206]), .Z(n918) );
  OR U1107 ( .A(n916), .B(n915), .Z(n917) );
  AND U1108 ( .A(n918), .B(n917), .Z(n920) );
  XOR U1109 ( .A(n921), .B(n920), .Z(c[1207]) );
  NAND U1110 ( .A(b[0]), .B(a[185]), .Z(n924) );
  XOR U1111 ( .A(sreg[1208]), .B(n924), .Z(n926) );
  NANDN U1112 ( .A(n919), .B(sreg[1207]), .Z(n923) );
  OR U1113 ( .A(n921), .B(n920), .Z(n922) );
  AND U1114 ( .A(n923), .B(n922), .Z(n925) );
  XOR U1115 ( .A(n926), .B(n925), .Z(c[1208]) );
  NAND U1116 ( .A(b[0]), .B(a[186]), .Z(n929) );
  XOR U1117 ( .A(sreg[1209]), .B(n929), .Z(n931) );
  NANDN U1118 ( .A(n924), .B(sreg[1208]), .Z(n928) );
  OR U1119 ( .A(n926), .B(n925), .Z(n927) );
  AND U1120 ( .A(n928), .B(n927), .Z(n930) );
  XOR U1121 ( .A(n931), .B(n930), .Z(c[1209]) );
  NAND U1122 ( .A(b[0]), .B(a[187]), .Z(n934) );
  XOR U1123 ( .A(sreg[1210]), .B(n934), .Z(n936) );
  NANDN U1124 ( .A(n929), .B(sreg[1209]), .Z(n933) );
  OR U1125 ( .A(n931), .B(n930), .Z(n932) );
  AND U1126 ( .A(n933), .B(n932), .Z(n935) );
  XOR U1127 ( .A(n936), .B(n935), .Z(c[1210]) );
  NAND U1128 ( .A(b[0]), .B(a[188]), .Z(n939) );
  XOR U1129 ( .A(sreg[1211]), .B(n939), .Z(n941) );
  NANDN U1130 ( .A(n934), .B(sreg[1210]), .Z(n938) );
  OR U1131 ( .A(n936), .B(n935), .Z(n937) );
  AND U1132 ( .A(n938), .B(n937), .Z(n940) );
  XOR U1133 ( .A(n941), .B(n940), .Z(c[1211]) );
  NAND U1134 ( .A(b[0]), .B(a[189]), .Z(n944) );
  XOR U1135 ( .A(sreg[1212]), .B(n944), .Z(n946) );
  NANDN U1136 ( .A(n939), .B(sreg[1211]), .Z(n943) );
  OR U1137 ( .A(n941), .B(n940), .Z(n942) );
  AND U1138 ( .A(n943), .B(n942), .Z(n945) );
  XOR U1139 ( .A(n946), .B(n945), .Z(c[1212]) );
  NAND U1140 ( .A(b[0]), .B(a[190]), .Z(n949) );
  XOR U1141 ( .A(sreg[1213]), .B(n949), .Z(n951) );
  NANDN U1142 ( .A(n944), .B(sreg[1212]), .Z(n948) );
  OR U1143 ( .A(n946), .B(n945), .Z(n947) );
  AND U1144 ( .A(n948), .B(n947), .Z(n950) );
  XOR U1145 ( .A(n951), .B(n950), .Z(c[1213]) );
  NAND U1146 ( .A(b[0]), .B(a[191]), .Z(n954) );
  XOR U1147 ( .A(sreg[1214]), .B(n954), .Z(n956) );
  NANDN U1148 ( .A(n949), .B(sreg[1213]), .Z(n953) );
  OR U1149 ( .A(n951), .B(n950), .Z(n952) );
  AND U1150 ( .A(n953), .B(n952), .Z(n955) );
  XOR U1151 ( .A(n956), .B(n955), .Z(c[1214]) );
  NAND U1152 ( .A(b[0]), .B(a[192]), .Z(n959) );
  XOR U1153 ( .A(sreg[1215]), .B(n959), .Z(n961) );
  NANDN U1154 ( .A(n954), .B(sreg[1214]), .Z(n958) );
  OR U1155 ( .A(n956), .B(n955), .Z(n957) );
  AND U1156 ( .A(n958), .B(n957), .Z(n960) );
  XOR U1157 ( .A(n961), .B(n960), .Z(c[1215]) );
  NAND U1158 ( .A(b[0]), .B(a[193]), .Z(n964) );
  XOR U1159 ( .A(sreg[1216]), .B(n964), .Z(n966) );
  NANDN U1160 ( .A(n959), .B(sreg[1215]), .Z(n963) );
  OR U1161 ( .A(n961), .B(n960), .Z(n962) );
  AND U1162 ( .A(n963), .B(n962), .Z(n965) );
  XOR U1163 ( .A(n966), .B(n965), .Z(c[1216]) );
  NAND U1164 ( .A(b[0]), .B(a[194]), .Z(n969) );
  XOR U1165 ( .A(sreg[1217]), .B(n969), .Z(n971) );
  NANDN U1166 ( .A(n964), .B(sreg[1216]), .Z(n968) );
  OR U1167 ( .A(n966), .B(n965), .Z(n967) );
  AND U1168 ( .A(n968), .B(n967), .Z(n970) );
  XOR U1169 ( .A(n971), .B(n970), .Z(c[1217]) );
  NAND U1170 ( .A(b[0]), .B(a[195]), .Z(n974) );
  XOR U1171 ( .A(sreg[1218]), .B(n974), .Z(n976) );
  NANDN U1172 ( .A(n969), .B(sreg[1217]), .Z(n973) );
  OR U1173 ( .A(n971), .B(n970), .Z(n972) );
  AND U1174 ( .A(n973), .B(n972), .Z(n975) );
  XOR U1175 ( .A(n976), .B(n975), .Z(c[1218]) );
  NAND U1176 ( .A(b[0]), .B(a[196]), .Z(n979) );
  XOR U1177 ( .A(sreg[1219]), .B(n979), .Z(n981) );
  NANDN U1178 ( .A(n974), .B(sreg[1218]), .Z(n978) );
  OR U1179 ( .A(n976), .B(n975), .Z(n977) );
  AND U1180 ( .A(n978), .B(n977), .Z(n980) );
  XOR U1181 ( .A(n981), .B(n980), .Z(c[1219]) );
  NAND U1182 ( .A(b[0]), .B(a[197]), .Z(n984) );
  XOR U1183 ( .A(sreg[1220]), .B(n984), .Z(n986) );
  NANDN U1184 ( .A(n979), .B(sreg[1219]), .Z(n983) );
  OR U1185 ( .A(n981), .B(n980), .Z(n982) );
  AND U1186 ( .A(n983), .B(n982), .Z(n985) );
  XOR U1187 ( .A(n986), .B(n985), .Z(c[1220]) );
  NAND U1188 ( .A(b[0]), .B(a[198]), .Z(n989) );
  XOR U1189 ( .A(sreg[1221]), .B(n989), .Z(n991) );
  NANDN U1190 ( .A(n984), .B(sreg[1220]), .Z(n988) );
  OR U1191 ( .A(n986), .B(n985), .Z(n987) );
  AND U1192 ( .A(n988), .B(n987), .Z(n990) );
  XOR U1193 ( .A(n991), .B(n990), .Z(c[1221]) );
  NAND U1194 ( .A(b[0]), .B(a[199]), .Z(n994) );
  XOR U1195 ( .A(sreg[1222]), .B(n994), .Z(n996) );
  NANDN U1196 ( .A(n989), .B(sreg[1221]), .Z(n993) );
  OR U1197 ( .A(n991), .B(n990), .Z(n992) );
  AND U1198 ( .A(n993), .B(n992), .Z(n995) );
  XOR U1199 ( .A(n996), .B(n995), .Z(c[1222]) );
  NAND U1200 ( .A(b[0]), .B(a[200]), .Z(n999) );
  XOR U1201 ( .A(sreg[1223]), .B(n999), .Z(n1001) );
  NANDN U1202 ( .A(n994), .B(sreg[1222]), .Z(n998) );
  OR U1203 ( .A(n996), .B(n995), .Z(n997) );
  AND U1204 ( .A(n998), .B(n997), .Z(n1000) );
  XOR U1205 ( .A(n1001), .B(n1000), .Z(c[1223]) );
  NAND U1206 ( .A(b[0]), .B(a[201]), .Z(n1004) );
  XOR U1207 ( .A(sreg[1224]), .B(n1004), .Z(n1006) );
  NANDN U1208 ( .A(n999), .B(sreg[1223]), .Z(n1003) );
  OR U1209 ( .A(n1001), .B(n1000), .Z(n1002) );
  AND U1210 ( .A(n1003), .B(n1002), .Z(n1005) );
  XOR U1211 ( .A(n1006), .B(n1005), .Z(c[1224]) );
  NAND U1212 ( .A(b[0]), .B(a[202]), .Z(n1009) );
  XOR U1213 ( .A(sreg[1225]), .B(n1009), .Z(n1011) );
  NANDN U1214 ( .A(n1004), .B(sreg[1224]), .Z(n1008) );
  OR U1215 ( .A(n1006), .B(n1005), .Z(n1007) );
  AND U1216 ( .A(n1008), .B(n1007), .Z(n1010) );
  XOR U1217 ( .A(n1011), .B(n1010), .Z(c[1225]) );
  NAND U1218 ( .A(b[0]), .B(a[203]), .Z(n1014) );
  XOR U1219 ( .A(sreg[1226]), .B(n1014), .Z(n1016) );
  NANDN U1220 ( .A(n1009), .B(sreg[1225]), .Z(n1013) );
  OR U1221 ( .A(n1011), .B(n1010), .Z(n1012) );
  AND U1222 ( .A(n1013), .B(n1012), .Z(n1015) );
  XOR U1223 ( .A(n1016), .B(n1015), .Z(c[1226]) );
  NAND U1224 ( .A(b[0]), .B(a[204]), .Z(n1019) );
  XOR U1225 ( .A(sreg[1227]), .B(n1019), .Z(n1021) );
  NANDN U1226 ( .A(n1014), .B(sreg[1226]), .Z(n1018) );
  OR U1227 ( .A(n1016), .B(n1015), .Z(n1017) );
  AND U1228 ( .A(n1018), .B(n1017), .Z(n1020) );
  XOR U1229 ( .A(n1021), .B(n1020), .Z(c[1227]) );
  NAND U1230 ( .A(b[0]), .B(a[205]), .Z(n1024) );
  XOR U1231 ( .A(sreg[1228]), .B(n1024), .Z(n1026) );
  NANDN U1232 ( .A(n1019), .B(sreg[1227]), .Z(n1023) );
  OR U1233 ( .A(n1021), .B(n1020), .Z(n1022) );
  AND U1234 ( .A(n1023), .B(n1022), .Z(n1025) );
  XOR U1235 ( .A(n1026), .B(n1025), .Z(c[1228]) );
  NAND U1236 ( .A(b[0]), .B(a[206]), .Z(n1029) );
  XOR U1237 ( .A(sreg[1229]), .B(n1029), .Z(n1031) );
  NANDN U1238 ( .A(n1024), .B(sreg[1228]), .Z(n1028) );
  OR U1239 ( .A(n1026), .B(n1025), .Z(n1027) );
  AND U1240 ( .A(n1028), .B(n1027), .Z(n1030) );
  XOR U1241 ( .A(n1031), .B(n1030), .Z(c[1229]) );
  NAND U1242 ( .A(b[0]), .B(a[207]), .Z(n1034) );
  XOR U1243 ( .A(sreg[1230]), .B(n1034), .Z(n1036) );
  NANDN U1244 ( .A(n1029), .B(sreg[1229]), .Z(n1033) );
  OR U1245 ( .A(n1031), .B(n1030), .Z(n1032) );
  AND U1246 ( .A(n1033), .B(n1032), .Z(n1035) );
  XOR U1247 ( .A(n1036), .B(n1035), .Z(c[1230]) );
  NAND U1248 ( .A(b[0]), .B(a[208]), .Z(n1039) );
  XOR U1249 ( .A(sreg[1231]), .B(n1039), .Z(n1041) );
  NANDN U1250 ( .A(n1034), .B(sreg[1230]), .Z(n1038) );
  OR U1251 ( .A(n1036), .B(n1035), .Z(n1037) );
  AND U1252 ( .A(n1038), .B(n1037), .Z(n1040) );
  XOR U1253 ( .A(n1041), .B(n1040), .Z(c[1231]) );
  NAND U1254 ( .A(b[0]), .B(a[209]), .Z(n1044) );
  XOR U1255 ( .A(sreg[1232]), .B(n1044), .Z(n1046) );
  NANDN U1256 ( .A(n1039), .B(sreg[1231]), .Z(n1043) );
  OR U1257 ( .A(n1041), .B(n1040), .Z(n1042) );
  AND U1258 ( .A(n1043), .B(n1042), .Z(n1045) );
  XOR U1259 ( .A(n1046), .B(n1045), .Z(c[1232]) );
  NAND U1260 ( .A(b[0]), .B(a[210]), .Z(n1049) );
  XOR U1261 ( .A(sreg[1233]), .B(n1049), .Z(n1051) );
  NANDN U1262 ( .A(n1044), .B(sreg[1232]), .Z(n1048) );
  OR U1263 ( .A(n1046), .B(n1045), .Z(n1047) );
  AND U1264 ( .A(n1048), .B(n1047), .Z(n1050) );
  XOR U1265 ( .A(n1051), .B(n1050), .Z(c[1233]) );
  NAND U1266 ( .A(b[0]), .B(a[211]), .Z(n1054) );
  XOR U1267 ( .A(sreg[1234]), .B(n1054), .Z(n1056) );
  NANDN U1268 ( .A(n1049), .B(sreg[1233]), .Z(n1053) );
  OR U1269 ( .A(n1051), .B(n1050), .Z(n1052) );
  AND U1270 ( .A(n1053), .B(n1052), .Z(n1055) );
  XOR U1271 ( .A(n1056), .B(n1055), .Z(c[1234]) );
  NAND U1272 ( .A(b[0]), .B(a[212]), .Z(n1059) );
  XOR U1273 ( .A(sreg[1235]), .B(n1059), .Z(n1061) );
  NANDN U1274 ( .A(n1054), .B(sreg[1234]), .Z(n1058) );
  OR U1275 ( .A(n1056), .B(n1055), .Z(n1057) );
  AND U1276 ( .A(n1058), .B(n1057), .Z(n1060) );
  XOR U1277 ( .A(n1061), .B(n1060), .Z(c[1235]) );
  NAND U1278 ( .A(b[0]), .B(a[213]), .Z(n1064) );
  XOR U1279 ( .A(sreg[1236]), .B(n1064), .Z(n1066) );
  NANDN U1280 ( .A(n1059), .B(sreg[1235]), .Z(n1063) );
  OR U1281 ( .A(n1061), .B(n1060), .Z(n1062) );
  AND U1282 ( .A(n1063), .B(n1062), .Z(n1065) );
  XOR U1283 ( .A(n1066), .B(n1065), .Z(c[1236]) );
  NAND U1284 ( .A(b[0]), .B(a[214]), .Z(n1069) );
  XOR U1285 ( .A(sreg[1237]), .B(n1069), .Z(n1071) );
  NANDN U1286 ( .A(n1064), .B(sreg[1236]), .Z(n1068) );
  OR U1287 ( .A(n1066), .B(n1065), .Z(n1067) );
  AND U1288 ( .A(n1068), .B(n1067), .Z(n1070) );
  XOR U1289 ( .A(n1071), .B(n1070), .Z(c[1237]) );
  NAND U1290 ( .A(b[0]), .B(a[215]), .Z(n1074) );
  XOR U1291 ( .A(sreg[1238]), .B(n1074), .Z(n1076) );
  NANDN U1292 ( .A(n1069), .B(sreg[1237]), .Z(n1073) );
  OR U1293 ( .A(n1071), .B(n1070), .Z(n1072) );
  AND U1294 ( .A(n1073), .B(n1072), .Z(n1075) );
  XOR U1295 ( .A(n1076), .B(n1075), .Z(c[1238]) );
  NAND U1296 ( .A(b[0]), .B(a[216]), .Z(n1079) );
  XOR U1297 ( .A(sreg[1239]), .B(n1079), .Z(n1081) );
  NANDN U1298 ( .A(n1074), .B(sreg[1238]), .Z(n1078) );
  OR U1299 ( .A(n1076), .B(n1075), .Z(n1077) );
  AND U1300 ( .A(n1078), .B(n1077), .Z(n1080) );
  XOR U1301 ( .A(n1081), .B(n1080), .Z(c[1239]) );
  NAND U1302 ( .A(b[0]), .B(a[217]), .Z(n1084) );
  XOR U1303 ( .A(sreg[1240]), .B(n1084), .Z(n1086) );
  NANDN U1304 ( .A(n1079), .B(sreg[1239]), .Z(n1083) );
  OR U1305 ( .A(n1081), .B(n1080), .Z(n1082) );
  AND U1306 ( .A(n1083), .B(n1082), .Z(n1085) );
  XOR U1307 ( .A(n1086), .B(n1085), .Z(c[1240]) );
  NAND U1308 ( .A(b[0]), .B(a[218]), .Z(n1089) );
  XOR U1309 ( .A(sreg[1241]), .B(n1089), .Z(n1091) );
  NANDN U1310 ( .A(n1084), .B(sreg[1240]), .Z(n1088) );
  OR U1311 ( .A(n1086), .B(n1085), .Z(n1087) );
  AND U1312 ( .A(n1088), .B(n1087), .Z(n1090) );
  XOR U1313 ( .A(n1091), .B(n1090), .Z(c[1241]) );
  NAND U1314 ( .A(b[0]), .B(a[219]), .Z(n1094) );
  XOR U1315 ( .A(sreg[1242]), .B(n1094), .Z(n1096) );
  NANDN U1316 ( .A(n1089), .B(sreg[1241]), .Z(n1093) );
  OR U1317 ( .A(n1091), .B(n1090), .Z(n1092) );
  AND U1318 ( .A(n1093), .B(n1092), .Z(n1095) );
  XOR U1319 ( .A(n1096), .B(n1095), .Z(c[1242]) );
  NAND U1320 ( .A(b[0]), .B(a[220]), .Z(n1099) );
  XOR U1321 ( .A(sreg[1243]), .B(n1099), .Z(n1101) );
  NANDN U1322 ( .A(n1094), .B(sreg[1242]), .Z(n1098) );
  OR U1323 ( .A(n1096), .B(n1095), .Z(n1097) );
  AND U1324 ( .A(n1098), .B(n1097), .Z(n1100) );
  XOR U1325 ( .A(n1101), .B(n1100), .Z(c[1243]) );
  NAND U1326 ( .A(b[0]), .B(a[221]), .Z(n1104) );
  XOR U1327 ( .A(sreg[1244]), .B(n1104), .Z(n1106) );
  NANDN U1328 ( .A(n1099), .B(sreg[1243]), .Z(n1103) );
  OR U1329 ( .A(n1101), .B(n1100), .Z(n1102) );
  AND U1330 ( .A(n1103), .B(n1102), .Z(n1105) );
  XOR U1331 ( .A(n1106), .B(n1105), .Z(c[1244]) );
  NAND U1332 ( .A(b[0]), .B(a[222]), .Z(n1109) );
  XOR U1333 ( .A(sreg[1245]), .B(n1109), .Z(n1111) );
  NANDN U1334 ( .A(n1104), .B(sreg[1244]), .Z(n1108) );
  OR U1335 ( .A(n1106), .B(n1105), .Z(n1107) );
  AND U1336 ( .A(n1108), .B(n1107), .Z(n1110) );
  XOR U1337 ( .A(n1111), .B(n1110), .Z(c[1245]) );
  NAND U1338 ( .A(b[0]), .B(a[223]), .Z(n1114) );
  XOR U1339 ( .A(sreg[1246]), .B(n1114), .Z(n1116) );
  NANDN U1340 ( .A(n1109), .B(sreg[1245]), .Z(n1113) );
  OR U1341 ( .A(n1111), .B(n1110), .Z(n1112) );
  AND U1342 ( .A(n1113), .B(n1112), .Z(n1115) );
  XOR U1343 ( .A(n1116), .B(n1115), .Z(c[1246]) );
  NAND U1344 ( .A(b[0]), .B(a[224]), .Z(n1119) );
  XOR U1345 ( .A(sreg[1247]), .B(n1119), .Z(n1121) );
  NANDN U1346 ( .A(n1114), .B(sreg[1246]), .Z(n1118) );
  OR U1347 ( .A(n1116), .B(n1115), .Z(n1117) );
  AND U1348 ( .A(n1118), .B(n1117), .Z(n1120) );
  XOR U1349 ( .A(n1121), .B(n1120), .Z(c[1247]) );
  NAND U1350 ( .A(b[0]), .B(a[225]), .Z(n1124) );
  XOR U1351 ( .A(sreg[1248]), .B(n1124), .Z(n1126) );
  NANDN U1352 ( .A(n1119), .B(sreg[1247]), .Z(n1123) );
  OR U1353 ( .A(n1121), .B(n1120), .Z(n1122) );
  AND U1354 ( .A(n1123), .B(n1122), .Z(n1125) );
  XOR U1355 ( .A(n1126), .B(n1125), .Z(c[1248]) );
  NAND U1356 ( .A(b[0]), .B(a[226]), .Z(n1129) );
  XOR U1357 ( .A(sreg[1249]), .B(n1129), .Z(n1131) );
  NANDN U1358 ( .A(n1124), .B(sreg[1248]), .Z(n1128) );
  OR U1359 ( .A(n1126), .B(n1125), .Z(n1127) );
  AND U1360 ( .A(n1128), .B(n1127), .Z(n1130) );
  XOR U1361 ( .A(n1131), .B(n1130), .Z(c[1249]) );
  NAND U1362 ( .A(b[0]), .B(a[227]), .Z(n1134) );
  XOR U1363 ( .A(sreg[1250]), .B(n1134), .Z(n1136) );
  NANDN U1364 ( .A(n1129), .B(sreg[1249]), .Z(n1133) );
  OR U1365 ( .A(n1131), .B(n1130), .Z(n1132) );
  AND U1366 ( .A(n1133), .B(n1132), .Z(n1135) );
  XOR U1367 ( .A(n1136), .B(n1135), .Z(c[1250]) );
  NAND U1368 ( .A(b[0]), .B(a[228]), .Z(n1139) );
  XOR U1369 ( .A(sreg[1251]), .B(n1139), .Z(n1141) );
  NANDN U1370 ( .A(n1134), .B(sreg[1250]), .Z(n1138) );
  OR U1371 ( .A(n1136), .B(n1135), .Z(n1137) );
  AND U1372 ( .A(n1138), .B(n1137), .Z(n1140) );
  XOR U1373 ( .A(n1141), .B(n1140), .Z(c[1251]) );
  NAND U1374 ( .A(b[0]), .B(a[229]), .Z(n1144) );
  XOR U1375 ( .A(sreg[1252]), .B(n1144), .Z(n1146) );
  NANDN U1376 ( .A(n1139), .B(sreg[1251]), .Z(n1143) );
  OR U1377 ( .A(n1141), .B(n1140), .Z(n1142) );
  AND U1378 ( .A(n1143), .B(n1142), .Z(n1145) );
  XOR U1379 ( .A(n1146), .B(n1145), .Z(c[1252]) );
  NAND U1380 ( .A(b[0]), .B(a[230]), .Z(n1149) );
  XOR U1381 ( .A(sreg[1253]), .B(n1149), .Z(n1151) );
  NANDN U1382 ( .A(n1144), .B(sreg[1252]), .Z(n1148) );
  OR U1383 ( .A(n1146), .B(n1145), .Z(n1147) );
  AND U1384 ( .A(n1148), .B(n1147), .Z(n1150) );
  XOR U1385 ( .A(n1151), .B(n1150), .Z(c[1253]) );
  NAND U1386 ( .A(b[0]), .B(a[231]), .Z(n1154) );
  XOR U1387 ( .A(sreg[1254]), .B(n1154), .Z(n1156) );
  NANDN U1388 ( .A(n1149), .B(sreg[1253]), .Z(n1153) );
  OR U1389 ( .A(n1151), .B(n1150), .Z(n1152) );
  AND U1390 ( .A(n1153), .B(n1152), .Z(n1155) );
  XOR U1391 ( .A(n1156), .B(n1155), .Z(c[1254]) );
  NAND U1392 ( .A(b[0]), .B(a[232]), .Z(n1159) );
  XOR U1393 ( .A(sreg[1255]), .B(n1159), .Z(n1161) );
  NANDN U1394 ( .A(n1154), .B(sreg[1254]), .Z(n1158) );
  OR U1395 ( .A(n1156), .B(n1155), .Z(n1157) );
  AND U1396 ( .A(n1158), .B(n1157), .Z(n1160) );
  XOR U1397 ( .A(n1161), .B(n1160), .Z(c[1255]) );
  NAND U1398 ( .A(b[0]), .B(a[233]), .Z(n1164) );
  XOR U1399 ( .A(sreg[1256]), .B(n1164), .Z(n1166) );
  NANDN U1400 ( .A(n1159), .B(sreg[1255]), .Z(n1163) );
  OR U1401 ( .A(n1161), .B(n1160), .Z(n1162) );
  AND U1402 ( .A(n1163), .B(n1162), .Z(n1165) );
  XOR U1403 ( .A(n1166), .B(n1165), .Z(c[1256]) );
  NAND U1404 ( .A(b[0]), .B(a[234]), .Z(n1169) );
  XOR U1405 ( .A(sreg[1257]), .B(n1169), .Z(n1171) );
  NANDN U1406 ( .A(n1164), .B(sreg[1256]), .Z(n1168) );
  OR U1407 ( .A(n1166), .B(n1165), .Z(n1167) );
  AND U1408 ( .A(n1168), .B(n1167), .Z(n1170) );
  XOR U1409 ( .A(n1171), .B(n1170), .Z(c[1257]) );
  NAND U1410 ( .A(b[0]), .B(a[235]), .Z(n1174) );
  XOR U1411 ( .A(sreg[1258]), .B(n1174), .Z(n1176) );
  NANDN U1412 ( .A(n1169), .B(sreg[1257]), .Z(n1173) );
  OR U1413 ( .A(n1171), .B(n1170), .Z(n1172) );
  AND U1414 ( .A(n1173), .B(n1172), .Z(n1175) );
  XOR U1415 ( .A(n1176), .B(n1175), .Z(c[1258]) );
  NAND U1416 ( .A(b[0]), .B(a[236]), .Z(n1179) );
  XOR U1417 ( .A(sreg[1259]), .B(n1179), .Z(n1181) );
  NANDN U1418 ( .A(n1174), .B(sreg[1258]), .Z(n1178) );
  OR U1419 ( .A(n1176), .B(n1175), .Z(n1177) );
  AND U1420 ( .A(n1178), .B(n1177), .Z(n1180) );
  XOR U1421 ( .A(n1181), .B(n1180), .Z(c[1259]) );
  NAND U1422 ( .A(b[0]), .B(a[237]), .Z(n1184) );
  XOR U1423 ( .A(sreg[1260]), .B(n1184), .Z(n1186) );
  NANDN U1424 ( .A(n1179), .B(sreg[1259]), .Z(n1183) );
  OR U1425 ( .A(n1181), .B(n1180), .Z(n1182) );
  AND U1426 ( .A(n1183), .B(n1182), .Z(n1185) );
  XOR U1427 ( .A(n1186), .B(n1185), .Z(c[1260]) );
  NAND U1428 ( .A(b[0]), .B(a[238]), .Z(n1189) );
  XOR U1429 ( .A(sreg[1261]), .B(n1189), .Z(n1191) );
  NANDN U1430 ( .A(n1184), .B(sreg[1260]), .Z(n1188) );
  OR U1431 ( .A(n1186), .B(n1185), .Z(n1187) );
  AND U1432 ( .A(n1188), .B(n1187), .Z(n1190) );
  XOR U1433 ( .A(n1191), .B(n1190), .Z(c[1261]) );
  NAND U1434 ( .A(b[0]), .B(a[239]), .Z(n1194) );
  XOR U1435 ( .A(sreg[1262]), .B(n1194), .Z(n1196) );
  NANDN U1436 ( .A(n1189), .B(sreg[1261]), .Z(n1193) );
  OR U1437 ( .A(n1191), .B(n1190), .Z(n1192) );
  AND U1438 ( .A(n1193), .B(n1192), .Z(n1195) );
  XOR U1439 ( .A(n1196), .B(n1195), .Z(c[1262]) );
  NAND U1440 ( .A(b[0]), .B(a[240]), .Z(n1199) );
  XOR U1441 ( .A(sreg[1263]), .B(n1199), .Z(n1201) );
  NANDN U1442 ( .A(n1194), .B(sreg[1262]), .Z(n1198) );
  OR U1443 ( .A(n1196), .B(n1195), .Z(n1197) );
  AND U1444 ( .A(n1198), .B(n1197), .Z(n1200) );
  XOR U1445 ( .A(n1201), .B(n1200), .Z(c[1263]) );
  NAND U1446 ( .A(b[0]), .B(a[241]), .Z(n1204) );
  XOR U1447 ( .A(sreg[1264]), .B(n1204), .Z(n1206) );
  NANDN U1448 ( .A(n1199), .B(sreg[1263]), .Z(n1203) );
  OR U1449 ( .A(n1201), .B(n1200), .Z(n1202) );
  AND U1450 ( .A(n1203), .B(n1202), .Z(n1205) );
  XOR U1451 ( .A(n1206), .B(n1205), .Z(c[1264]) );
  NAND U1452 ( .A(b[0]), .B(a[242]), .Z(n1209) );
  XOR U1453 ( .A(sreg[1265]), .B(n1209), .Z(n1211) );
  NANDN U1454 ( .A(n1204), .B(sreg[1264]), .Z(n1208) );
  OR U1455 ( .A(n1206), .B(n1205), .Z(n1207) );
  AND U1456 ( .A(n1208), .B(n1207), .Z(n1210) );
  XOR U1457 ( .A(n1211), .B(n1210), .Z(c[1265]) );
  NAND U1458 ( .A(b[0]), .B(a[243]), .Z(n1214) );
  XOR U1459 ( .A(sreg[1266]), .B(n1214), .Z(n1216) );
  NANDN U1460 ( .A(n1209), .B(sreg[1265]), .Z(n1213) );
  OR U1461 ( .A(n1211), .B(n1210), .Z(n1212) );
  AND U1462 ( .A(n1213), .B(n1212), .Z(n1215) );
  XOR U1463 ( .A(n1216), .B(n1215), .Z(c[1266]) );
  NAND U1464 ( .A(b[0]), .B(a[244]), .Z(n1219) );
  XOR U1465 ( .A(sreg[1267]), .B(n1219), .Z(n1221) );
  NANDN U1466 ( .A(n1214), .B(sreg[1266]), .Z(n1218) );
  OR U1467 ( .A(n1216), .B(n1215), .Z(n1217) );
  AND U1468 ( .A(n1218), .B(n1217), .Z(n1220) );
  XOR U1469 ( .A(n1221), .B(n1220), .Z(c[1267]) );
  NAND U1470 ( .A(b[0]), .B(a[245]), .Z(n1224) );
  XOR U1471 ( .A(sreg[1268]), .B(n1224), .Z(n1226) );
  NANDN U1472 ( .A(n1219), .B(sreg[1267]), .Z(n1223) );
  OR U1473 ( .A(n1221), .B(n1220), .Z(n1222) );
  AND U1474 ( .A(n1223), .B(n1222), .Z(n1225) );
  XOR U1475 ( .A(n1226), .B(n1225), .Z(c[1268]) );
  NAND U1476 ( .A(b[0]), .B(a[246]), .Z(n1229) );
  XOR U1477 ( .A(sreg[1269]), .B(n1229), .Z(n1231) );
  NANDN U1478 ( .A(n1224), .B(sreg[1268]), .Z(n1228) );
  OR U1479 ( .A(n1226), .B(n1225), .Z(n1227) );
  AND U1480 ( .A(n1228), .B(n1227), .Z(n1230) );
  XOR U1481 ( .A(n1231), .B(n1230), .Z(c[1269]) );
  NAND U1482 ( .A(b[0]), .B(a[247]), .Z(n1234) );
  XOR U1483 ( .A(sreg[1270]), .B(n1234), .Z(n1236) );
  NANDN U1484 ( .A(n1229), .B(sreg[1269]), .Z(n1233) );
  OR U1485 ( .A(n1231), .B(n1230), .Z(n1232) );
  AND U1486 ( .A(n1233), .B(n1232), .Z(n1235) );
  XOR U1487 ( .A(n1236), .B(n1235), .Z(c[1270]) );
  NAND U1488 ( .A(b[0]), .B(a[248]), .Z(n1239) );
  XOR U1489 ( .A(sreg[1271]), .B(n1239), .Z(n1241) );
  NANDN U1490 ( .A(n1234), .B(sreg[1270]), .Z(n1238) );
  OR U1491 ( .A(n1236), .B(n1235), .Z(n1237) );
  AND U1492 ( .A(n1238), .B(n1237), .Z(n1240) );
  XOR U1493 ( .A(n1241), .B(n1240), .Z(c[1271]) );
  NAND U1494 ( .A(b[0]), .B(a[249]), .Z(n1244) );
  XOR U1495 ( .A(sreg[1272]), .B(n1244), .Z(n1246) );
  NANDN U1496 ( .A(n1239), .B(sreg[1271]), .Z(n1243) );
  OR U1497 ( .A(n1241), .B(n1240), .Z(n1242) );
  AND U1498 ( .A(n1243), .B(n1242), .Z(n1245) );
  XOR U1499 ( .A(n1246), .B(n1245), .Z(c[1272]) );
  NAND U1500 ( .A(b[0]), .B(a[250]), .Z(n1249) );
  XOR U1501 ( .A(sreg[1273]), .B(n1249), .Z(n1251) );
  NANDN U1502 ( .A(n1244), .B(sreg[1272]), .Z(n1248) );
  OR U1503 ( .A(n1246), .B(n1245), .Z(n1247) );
  AND U1504 ( .A(n1248), .B(n1247), .Z(n1250) );
  XOR U1505 ( .A(n1251), .B(n1250), .Z(c[1273]) );
  NAND U1506 ( .A(b[0]), .B(a[251]), .Z(n1254) );
  XOR U1507 ( .A(sreg[1274]), .B(n1254), .Z(n1256) );
  NANDN U1508 ( .A(n1249), .B(sreg[1273]), .Z(n1253) );
  OR U1509 ( .A(n1251), .B(n1250), .Z(n1252) );
  AND U1510 ( .A(n1253), .B(n1252), .Z(n1255) );
  XOR U1511 ( .A(n1256), .B(n1255), .Z(c[1274]) );
  NAND U1512 ( .A(b[0]), .B(a[252]), .Z(n1259) );
  XOR U1513 ( .A(sreg[1275]), .B(n1259), .Z(n1261) );
  NANDN U1514 ( .A(n1254), .B(sreg[1274]), .Z(n1258) );
  OR U1515 ( .A(n1256), .B(n1255), .Z(n1257) );
  AND U1516 ( .A(n1258), .B(n1257), .Z(n1260) );
  XOR U1517 ( .A(n1261), .B(n1260), .Z(c[1275]) );
  NAND U1518 ( .A(b[0]), .B(a[253]), .Z(n1264) );
  XOR U1519 ( .A(sreg[1276]), .B(n1264), .Z(n1266) );
  NANDN U1520 ( .A(n1259), .B(sreg[1275]), .Z(n1263) );
  OR U1521 ( .A(n1261), .B(n1260), .Z(n1262) );
  AND U1522 ( .A(n1263), .B(n1262), .Z(n1265) );
  XOR U1523 ( .A(n1266), .B(n1265), .Z(c[1276]) );
  NAND U1524 ( .A(b[0]), .B(a[254]), .Z(n1269) );
  XOR U1525 ( .A(sreg[1277]), .B(n1269), .Z(n1271) );
  NANDN U1526 ( .A(n1264), .B(sreg[1276]), .Z(n1268) );
  OR U1527 ( .A(n1266), .B(n1265), .Z(n1267) );
  AND U1528 ( .A(n1268), .B(n1267), .Z(n1270) );
  XOR U1529 ( .A(n1271), .B(n1270), .Z(c[1277]) );
  NAND U1530 ( .A(b[0]), .B(a[255]), .Z(n1274) );
  XOR U1531 ( .A(sreg[1278]), .B(n1274), .Z(n1276) );
  NANDN U1532 ( .A(n1269), .B(sreg[1277]), .Z(n1273) );
  OR U1533 ( .A(n1271), .B(n1270), .Z(n1272) );
  AND U1534 ( .A(n1273), .B(n1272), .Z(n1275) );
  XOR U1535 ( .A(n1276), .B(n1275), .Z(c[1278]) );
  NAND U1536 ( .A(b[0]), .B(a[256]), .Z(n1279) );
  XOR U1537 ( .A(sreg[1279]), .B(n1279), .Z(n1281) );
  NANDN U1538 ( .A(n1274), .B(sreg[1278]), .Z(n1278) );
  OR U1539 ( .A(n1276), .B(n1275), .Z(n1277) );
  AND U1540 ( .A(n1278), .B(n1277), .Z(n1280) );
  XOR U1541 ( .A(n1281), .B(n1280), .Z(c[1279]) );
  NAND U1542 ( .A(b[0]), .B(a[257]), .Z(n1284) );
  XOR U1543 ( .A(sreg[1280]), .B(n1284), .Z(n1286) );
  NANDN U1544 ( .A(n1279), .B(sreg[1279]), .Z(n1283) );
  OR U1545 ( .A(n1281), .B(n1280), .Z(n1282) );
  AND U1546 ( .A(n1283), .B(n1282), .Z(n1285) );
  XOR U1547 ( .A(n1286), .B(n1285), .Z(c[1280]) );
  NAND U1548 ( .A(b[0]), .B(a[258]), .Z(n1289) );
  XOR U1549 ( .A(sreg[1281]), .B(n1289), .Z(n1291) );
  NANDN U1550 ( .A(n1284), .B(sreg[1280]), .Z(n1288) );
  OR U1551 ( .A(n1286), .B(n1285), .Z(n1287) );
  AND U1552 ( .A(n1288), .B(n1287), .Z(n1290) );
  XOR U1553 ( .A(n1291), .B(n1290), .Z(c[1281]) );
  NAND U1554 ( .A(b[0]), .B(a[259]), .Z(n1294) );
  XOR U1555 ( .A(sreg[1282]), .B(n1294), .Z(n1296) );
  NANDN U1556 ( .A(n1289), .B(sreg[1281]), .Z(n1293) );
  OR U1557 ( .A(n1291), .B(n1290), .Z(n1292) );
  AND U1558 ( .A(n1293), .B(n1292), .Z(n1295) );
  XOR U1559 ( .A(n1296), .B(n1295), .Z(c[1282]) );
  NAND U1560 ( .A(b[0]), .B(a[260]), .Z(n1299) );
  XOR U1561 ( .A(sreg[1283]), .B(n1299), .Z(n1301) );
  NANDN U1562 ( .A(n1294), .B(sreg[1282]), .Z(n1298) );
  OR U1563 ( .A(n1296), .B(n1295), .Z(n1297) );
  AND U1564 ( .A(n1298), .B(n1297), .Z(n1300) );
  XOR U1565 ( .A(n1301), .B(n1300), .Z(c[1283]) );
  NAND U1566 ( .A(b[0]), .B(a[261]), .Z(n1304) );
  XOR U1567 ( .A(sreg[1284]), .B(n1304), .Z(n1306) );
  NANDN U1568 ( .A(n1299), .B(sreg[1283]), .Z(n1303) );
  OR U1569 ( .A(n1301), .B(n1300), .Z(n1302) );
  AND U1570 ( .A(n1303), .B(n1302), .Z(n1305) );
  XOR U1571 ( .A(n1306), .B(n1305), .Z(c[1284]) );
  NAND U1572 ( .A(b[0]), .B(a[262]), .Z(n1309) );
  XOR U1573 ( .A(sreg[1285]), .B(n1309), .Z(n1311) );
  NANDN U1574 ( .A(n1304), .B(sreg[1284]), .Z(n1308) );
  OR U1575 ( .A(n1306), .B(n1305), .Z(n1307) );
  AND U1576 ( .A(n1308), .B(n1307), .Z(n1310) );
  XOR U1577 ( .A(n1311), .B(n1310), .Z(c[1285]) );
  NAND U1578 ( .A(b[0]), .B(a[263]), .Z(n1314) );
  XOR U1579 ( .A(sreg[1286]), .B(n1314), .Z(n1316) );
  NANDN U1580 ( .A(n1309), .B(sreg[1285]), .Z(n1313) );
  OR U1581 ( .A(n1311), .B(n1310), .Z(n1312) );
  AND U1582 ( .A(n1313), .B(n1312), .Z(n1315) );
  XOR U1583 ( .A(n1316), .B(n1315), .Z(c[1286]) );
  NAND U1584 ( .A(b[0]), .B(a[264]), .Z(n1319) );
  XOR U1585 ( .A(sreg[1287]), .B(n1319), .Z(n1321) );
  NANDN U1586 ( .A(n1314), .B(sreg[1286]), .Z(n1318) );
  OR U1587 ( .A(n1316), .B(n1315), .Z(n1317) );
  AND U1588 ( .A(n1318), .B(n1317), .Z(n1320) );
  XOR U1589 ( .A(n1321), .B(n1320), .Z(c[1287]) );
  NAND U1590 ( .A(b[0]), .B(a[265]), .Z(n1324) );
  XOR U1591 ( .A(sreg[1288]), .B(n1324), .Z(n1326) );
  NANDN U1592 ( .A(n1319), .B(sreg[1287]), .Z(n1323) );
  OR U1593 ( .A(n1321), .B(n1320), .Z(n1322) );
  AND U1594 ( .A(n1323), .B(n1322), .Z(n1325) );
  XOR U1595 ( .A(n1326), .B(n1325), .Z(c[1288]) );
  NAND U1596 ( .A(b[0]), .B(a[266]), .Z(n1329) );
  XOR U1597 ( .A(sreg[1289]), .B(n1329), .Z(n1331) );
  NANDN U1598 ( .A(n1324), .B(sreg[1288]), .Z(n1328) );
  OR U1599 ( .A(n1326), .B(n1325), .Z(n1327) );
  AND U1600 ( .A(n1328), .B(n1327), .Z(n1330) );
  XOR U1601 ( .A(n1331), .B(n1330), .Z(c[1289]) );
  NAND U1602 ( .A(b[0]), .B(a[267]), .Z(n1334) );
  XOR U1603 ( .A(sreg[1290]), .B(n1334), .Z(n1336) );
  NANDN U1604 ( .A(n1329), .B(sreg[1289]), .Z(n1333) );
  OR U1605 ( .A(n1331), .B(n1330), .Z(n1332) );
  AND U1606 ( .A(n1333), .B(n1332), .Z(n1335) );
  XOR U1607 ( .A(n1336), .B(n1335), .Z(c[1290]) );
  NAND U1608 ( .A(b[0]), .B(a[268]), .Z(n1339) );
  XOR U1609 ( .A(sreg[1291]), .B(n1339), .Z(n1341) );
  NANDN U1610 ( .A(n1334), .B(sreg[1290]), .Z(n1338) );
  OR U1611 ( .A(n1336), .B(n1335), .Z(n1337) );
  AND U1612 ( .A(n1338), .B(n1337), .Z(n1340) );
  XOR U1613 ( .A(n1341), .B(n1340), .Z(c[1291]) );
  NAND U1614 ( .A(b[0]), .B(a[269]), .Z(n1344) );
  XOR U1615 ( .A(sreg[1292]), .B(n1344), .Z(n1346) );
  NANDN U1616 ( .A(n1339), .B(sreg[1291]), .Z(n1343) );
  OR U1617 ( .A(n1341), .B(n1340), .Z(n1342) );
  AND U1618 ( .A(n1343), .B(n1342), .Z(n1345) );
  XOR U1619 ( .A(n1346), .B(n1345), .Z(c[1292]) );
  NAND U1620 ( .A(b[0]), .B(a[270]), .Z(n1349) );
  XOR U1621 ( .A(sreg[1293]), .B(n1349), .Z(n1351) );
  NANDN U1622 ( .A(n1344), .B(sreg[1292]), .Z(n1348) );
  OR U1623 ( .A(n1346), .B(n1345), .Z(n1347) );
  AND U1624 ( .A(n1348), .B(n1347), .Z(n1350) );
  XOR U1625 ( .A(n1351), .B(n1350), .Z(c[1293]) );
  NAND U1626 ( .A(b[0]), .B(a[271]), .Z(n1354) );
  XOR U1627 ( .A(sreg[1294]), .B(n1354), .Z(n1356) );
  NANDN U1628 ( .A(n1349), .B(sreg[1293]), .Z(n1353) );
  OR U1629 ( .A(n1351), .B(n1350), .Z(n1352) );
  AND U1630 ( .A(n1353), .B(n1352), .Z(n1355) );
  XOR U1631 ( .A(n1356), .B(n1355), .Z(c[1294]) );
  NAND U1632 ( .A(b[0]), .B(a[272]), .Z(n1359) );
  XOR U1633 ( .A(sreg[1295]), .B(n1359), .Z(n1361) );
  NANDN U1634 ( .A(n1354), .B(sreg[1294]), .Z(n1358) );
  OR U1635 ( .A(n1356), .B(n1355), .Z(n1357) );
  AND U1636 ( .A(n1358), .B(n1357), .Z(n1360) );
  XOR U1637 ( .A(n1361), .B(n1360), .Z(c[1295]) );
  NAND U1638 ( .A(b[0]), .B(a[273]), .Z(n1364) );
  XOR U1639 ( .A(sreg[1296]), .B(n1364), .Z(n1366) );
  NANDN U1640 ( .A(n1359), .B(sreg[1295]), .Z(n1363) );
  OR U1641 ( .A(n1361), .B(n1360), .Z(n1362) );
  AND U1642 ( .A(n1363), .B(n1362), .Z(n1365) );
  XOR U1643 ( .A(n1366), .B(n1365), .Z(c[1296]) );
  NAND U1644 ( .A(b[0]), .B(a[274]), .Z(n1369) );
  XOR U1645 ( .A(sreg[1297]), .B(n1369), .Z(n1371) );
  NANDN U1646 ( .A(n1364), .B(sreg[1296]), .Z(n1368) );
  OR U1647 ( .A(n1366), .B(n1365), .Z(n1367) );
  AND U1648 ( .A(n1368), .B(n1367), .Z(n1370) );
  XOR U1649 ( .A(n1371), .B(n1370), .Z(c[1297]) );
  NAND U1650 ( .A(b[0]), .B(a[275]), .Z(n1374) );
  XOR U1651 ( .A(sreg[1298]), .B(n1374), .Z(n1376) );
  NANDN U1652 ( .A(n1369), .B(sreg[1297]), .Z(n1373) );
  OR U1653 ( .A(n1371), .B(n1370), .Z(n1372) );
  AND U1654 ( .A(n1373), .B(n1372), .Z(n1375) );
  XOR U1655 ( .A(n1376), .B(n1375), .Z(c[1298]) );
  NAND U1656 ( .A(b[0]), .B(a[276]), .Z(n1379) );
  XOR U1657 ( .A(sreg[1299]), .B(n1379), .Z(n1381) );
  NANDN U1658 ( .A(n1374), .B(sreg[1298]), .Z(n1378) );
  OR U1659 ( .A(n1376), .B(n1375), .Z(n1377) );
  AND U1660 ( .A(n1378), .B(n1377), .Z(n1380) );
  XOR U1661 ( .A(n1381), .B(n1380), .Z(c[1299]) );
  NAND U1662 ( .A(b[0]), .B(a[277]), .Z(n1384) );
  XOR U1663 ( .A(sreg[1300]), .B(n1384), .Z(n1386) );
  NANDN U1664 ( .A(n1379), .B(sreg[1299]), .Z(n1383) );
  OR U1665 ( .A(n1381), .B(n1380), .Z(n1382) );
  AND U1666 ( .A(n1383), .B(n1382), .Z(n1385) );
  XOR U1667 ( .A(n1386), .B(n1385), .Z(c[1300]) );
  NAND U1668 ( .A(b[0]), .B(a[278]), .Z(n1389) );
  XOR U1669 ( .A(sreg[1301]), .B(n1389), .Z(n1391) );
  NANDN U1670 ( .A(n1384), .B(sreg[1300]), .Z(n1388) );
  OR U1671 ( .A(n1386), .B(n1385), .Z(n1387) );
  AND U1672 ( .A(n1388), .B(n1387), .Z(n1390) );
  XOR U1673 ( .A(n1391), .B(n1390), .Z(c[1301]) );
  NAND U1674 ( .A(b[0]), .B(a[279]), .Z(n1394) );
  XOR U1675 ( .A(sreg[1302]), .B(n1394), .Z(n1396) );
  NANDN U1676 ( .A(n1389), .B(sreg[1301]), .Z(n1393) );
  OR U1677 ( .A(n1391), .B(n1390), .Z(n1392) );
  AND U1678 ( .A(n1393), .B(n1392), .Z(n1395) );
  XOR U1679 ( .A(n1396), .B(n1395), .Z(c[1302]) );
  NAND U1680 ( .A(b[0]), .B(a[280]), .Z(n1399) );
  XOR U1681 ( .A(sreg[1303]), .B(n1399), .Z(n1401) );
  NANDN U1682 ( .A(n1394), .B(sreg[1302]), .Z(n1398) );
  OR U1683 ( .A(n1396), .B(n1395), .Z(n1397) );
  AND U1684 ( .A(n1398), .B(n1397), .Z(n1400) );
  XOR U1685 ( .A(n1401), .B(n1400), .Z(c[1303]) );
  NAND U1686 ( .A(b[0]), .B(a[281]), .Z(n1404) );
  XOR U1687 ( .A(sreg[1304]), .B(n1404), .Z(n1406) );
  NANDN U1688 ( .A(n1399), .B(sreg[1303]), .Z(n1403) );
  OR U1689 ( .A(n1401), .B(n1400), .Z(n1402) );
  AND U1690 ( .A(n1403), .B(n1402), .Z(n1405) );
  XOR U1691 ( .A(n1406), .B(n1405), .Z(c[1304]) );
  NAND U1692 ( .A(b[0]), .B(a[282]), .Z(n1409) );
  XOR U1693 ( .A(sreg[1305]), .B(n1409), .Z(n1411) );
  NANDN U1694 ( .A(n1404), .B(sreg[1304]), .Z(n1408) );
  OR U1695 ( .A(n1406), .B(n1405), .Z(n1407) );
  AND U1696 ( .A(n1408), .B(n1407), .Z(n1410) );
  XOR U1697 ( .A(n1411), .B(n1410), .Z(c[1305]) );
  NAND U1698 ( .A(b[0]), .B(a[283]), .Z(n1414) );
  XOR U1699 ( .A(sreg[1306]), .B(n1414), .Z(n1416) );
  NANDN U1700 ( .A(n1409), .B(sreg[1305]), .Z(n1413) );
  OR U1701 ( .A(n1411), .B(n1410), .Z(n1412) );
  AND U1702 ( .A(n1413), .B(n1412), .Z(n1415) );
  XOR U1703 ( .A(n1416), .B(n1415), .Z(c[1306]) );
  NAND U1704 ( .A(b[0]), .B(a[284]), .Z(n1419) );
  XOR U1705 ( .A(sreg[1307]), .B(n1419), .Z(n1421) );
  NANDN U1706 ( .A(n1414), .B(sreg[1306]), .Z(n1418) );
  OR U1707 ( .A(n1416), .B(n1415), .Z(n1417) );
  AND U1708 ( .A(n1418), .B(n1417), .Z(n1420) );
  XOR U1709 ( .A(n1421), .B(n1420), .Z(c[1307]) );
  NAND U1710 ( .A(b[0]), .B(a[285]), .Z(n1424) );
  XOR U1711 ( .A(sreg[1308]), .B(n1424), .Z(n1426) );
  NANDN U1712 ( .A(n1419), .B(sreg[1307]), .Z(n1423) );
  OR U1713 ( .A(n1421), .B(n1420), .Z(n1422) );
  AND U1714 ( .A(n1423), .B(n1422), .Z(n1425) );
  XOR U1715 ( .A(n1426), .B(n1425), .Z(c[1308]) );
  NAND U1716 ( .A(b[0]), .B(a[286]), .Z(n1429) );
  XOR U1717 ( .A(sreg[1309]), .B(n1429), .Z(n1431) );
  NANDN U1718 ( .A(n1424), .B(sreg[1308]), .Z(n1428) );
  OR U1719 ( .A(n1426), .B(n1425), .Z(n1427) );
  AND U1720 ( .A(n1428), .B(n1427), .Z(n1430) );
  XOR U1721 ( .A(n1431), .B(n1430), .Z(c[1309]) );
  NAND U1722 ( .A(b[0]), .B(a[287]), .Z(n1434) );
  XOR U1723 ( .A(sreg[1310]), .B(n1434), .Z(n1436) );
  NANDN U1724 ( .A(n1429), .B(sreg[1309]), .Z(n1433) );
  OR U1725 ( .A(n1431), .B(n1430), .Z(n1432) );
  AND U1726 ( .A(n1433), .B(n1432), .Z(n1435) );
  XOR U1727 ( .A(n1436), .B(n1435), .Z(c[1310]) );
  NAND U1728 ( .A(b[0]), .B(a[288]), .Z(n1439) );
  XOR U1729 ( .A(sreg[1311]), .B(n1439), .Z(n1441) );
  NANDN U1730 ( .A(n1434), .B(sreg[1310]), .Z(n1438) );
  OR U1731 ( .A(n1436), .B(n1435), .Z(n1437) );
  AND U1732 ( .A(n1438), .B(n1437), .Z(n1440) );
  XOR U1733 ( .A(n1441), .B(n1440), .Z(c[1311]) );
  NAND U1734 ( .A(b[0]), .B(a[289]), .Z(n1444) );
  XOR U1735 ( .A(sreg[1312]), .B(n1444), .Z(n1446) );
  NANDN U1736 ( .A(n1439), .B(sreg[1311]), .Z(n1443) );
  OR U1737 ( .A(n1441), .B(n1440), .Z(n1442) );
  AND U1738 ( .A(n1443), .B(n1442), .Z(n1445) );
  XOR U1739 ( .A(n1446), .B(n1445), .Z(c[1312]) );
  NAND U1740 ( .A(b[0]), .B(a[290]), .Z(n1449) );
  XOR U1741 ( .A(sreg[1313]), .B(n1449), .Z(n1451) );
  NANDN U1742 ( .A(n1444), .B(sreg[1312]), .Z(n1448) );
  OR U1743 ( .A(n1446), .B(n1445), .Z(n1447) );
  AND U1744 ( .A(n1448), .B(n1447), .Z(n1450) );
  XOR U1745 ( .A(n1451), .B(n1450), .Z(c[1313]) );
  NAND U1746 ( .A(b[0]), .B(a[291]), .Z(n1454) );
  XOR U1747 ( .A(sreg[1314]), .B(n1454), .Z(n1456) );
  NANDN U1748 ( .A(n1449), .B(sreg[1313]), .Z(n1453) );
  OR U1749 ( .A(n1451), .B(n1450), .Z(n1452) );
  AND U1750 ( .A(n1453), .B(n1452), .Z(n1455) );
  XOR U1751 ( .A(n1456), .B(n1455), .Z(c[1314]) );
  NAND U1752 ( .A(b[0]), .B(a[292]), .Z(n1459) );
  XOR U1753 ( .A(sreg[1315]), .B(n1459), .Z(n1461) );
  NANDN U1754 ( .A(n1454), .B(sreg[1314]), .Z(n1458) );
  OR U1755 ( .A(n1456), .B(n1455), .Z(n1457) );
  AND U1756 ( .A(n1458), .B(n1457), .Z(n1460) );
  XOR U1757 ( .A(n1461), .B(n1460), .Z(c[1315]) );
  NAND U1758 ( .A(b[0]), .B(a[293]), .Z(n1464) );
  XOR U1759 ( .A(sreg[1316]), .B(n1464), .Z(n1466) );
  NANDN U1760 ( .A(n1459), .B(sreg[1315]), .Z(n1463) );
  OR U1761 ( .A(n1461), .B(n1460), .Z(n1462) );
  AND U1762 ( .A(n1463), .B(n1462), .Z(n1465) );
  XOR U1763 ( .A(n1466), .B(n1465), .Z(c[1316]) );
  NAND U1764 ( .A(b[0]), .B(a[294]), .Z(n1469) );
  XOR U1765 ( .A(sreg[1317]), .B(n1469), .Z(n1471) );
  NANDN U1766 ( .A(n1464), .B(sreg[1316]), .Z(n1468) );
  OR U1767 ( .A(n1466), .B(n1465), .Z(n1467) );
  AND U1768 ( .A(n1468), .B(n1467), .Z(n1470) );
  XOR U1769 ( .A(n1471), .B(n1470), .Z(c[1317]) );
  NAND U1770 ( .A(b[0]), .B(a[295]), .Z(n1474) );
  XOR U1771 ( .A(sreg[1318]), .B(n1474), .Z(n1476) );
  NANDN U1772 ( .A(n1469), .B(sreg[1317]), .Z(n1473) );
  OR U1773 ( .A(n1471), .B(n1470), .Z(n1472) );
  AND U1774 ( .A(n1473), .B(n1472), .Z(n1475) );
  XOR U1775 ( .A(n1476), .B(n1475), .Z(c[1318]) );
  NAND U1776 ( .A(b[0]), .B(a[296]), .Z(n1479) );
  XOR U1777 ( .A(sreg[1319]), .B(n1479), .Z(n1481) );
  NANDN U1778 ( .A(n1474), .B(sreg[1318]), .Z(n1478) );
  OR U1779 ( .A(n1476), .B(n1475), .Z(n1477) );
  AND U1780 ( .A(n1478), .B(n1477), .Z(n1480) );
  XOR U1781 ( .A(n1481), .B(n1480), .Z(c[1319]) );
  NAND U1782 ( .A(b[0]), .B(a[297]), .Z(n1484) );
  XOR U1783 ( .A(sreg[1320]), .B(n1484), .Z(n1486) );
  NANDN U1784 ( .A(n1479), .B(sreg[1319]), .Z(n1483) );
  OR U1785 ( .A(n1481), .B(n1480), .Z(n1482) );
  AND U1786 ( .A(n1483), .B(n1482), .Z(n1485) );
  XOR U1787 ( .A(n1486), .B(n1485), .Z(c[1320]) );
  NAND U1788 ( .A(b[0]), .B(a[298]), .Z(n1489) );
  XOR U1789 ( .A(sreg[1321]), .B(n1489), .Z(n1491) );
  NANDN U1790 ( .A(n1484), .B(sreg[1320]), .Z(n1488) );
  OR U1791 ( .A(n1486), .B(n1485), .Z(n1487) );
  AND U1792 ( .A(n1488), .B(n1487), .Z(n1490) );
  XOR U1793 ( .A(n1491), .B(n1490), .Z(c[1321]) );
  NAND U1794 ( .A(b[0]), .B(a[299]), .Z(n1494) );
  XOR U1795 ( .A(sreg[1322]), .B(n1494), .Z(n1496) );
  NANDN U1796 ( .A(n1489), .B(sreg[1321]), .Z(n1493) );
  OR U1797 ( .A(n1491), .B(n1490), .Z(n1492) );
  AND U1798 ( .A(n1493), .B(n1492), .Z(n1495) );
  XOR U1799 ( .A(n1496), .B(n1495), .Z(c[1322]) );
  NAND U1800 ( .A(b[0]), .B(a[300]), .Z(n1499) );
  XOR U1801 ( .A(sreg[1323]), .B(n1499), .Z(n1501) );
  NANDN U1802 ( .A(n1494), .B(sreg[1322]), .Z(n1498) );
  OR U1803 ( .A(n1496), .B(n1495), .Z(n1497) );
  AND U1804 ( .A(n1498), .B(n1497), .Z(n1500) );
  XOR U1805 ( .A(n1501), .B(n1500), .Z(c[1323]) );
  NAND U1806 ( .A(b[0]), .B(a[301]), .Z(n1504) );
  XOR U1807 ( .A(sreg[1324]), .B(n1504), .Z(n1506) );
  NANDN U1808 ( .A(n1499), .B(sreg[1323]), .Z(n1503) );
  OR U1809 ( .A(n1501), .B(n1500), .Z(n1502) );
  AND U1810 ( .A(n1503), .B(n1502), .Z(n1505) );
  XOR U1811 ( .A(n1506), .B(n1505), .Z(c[1324]) );
  NAND U1812 ( .A(b[0]), .B(a[302]), .Z(n1509) );
  XOR U1813 ( .A(sreg[1325]), .B(n1509), .Z(n1511) );
  NANDN U1814 ( .A(n1504), .B(sreg[1324]), .Z(n1508) );
  OR U1815 ( .A(n1506), .B(n1505), .Z(n1507) );
  AND U1816 ( .A(n1508), .B(n1507), .Z(n1510) );
  XOR U1817 ( .A(n1511), .B(n1510), .Z(c[1325]) );
  NAND U1818 ( .A(b[0]), .B(a[303]), .Z(n1514) );
  XOR U1819 ( .A(sreg[1326]), .B(n1514), .Z(n1516) );
  NANDN U1820 ( .A(n1509), .B(sreg[1325]), .Z(n1513) );
  OR U1821 ( .A(n1511), .B(n1510), .Z(n1512) );
  AND U1822 ( .A(n1513), .B(n1512), .Z(n1515) );
  XOR U1823 ( .A(n1516), .B(n1515), .Z(c[1326]) );
  NAND U1824 ( .A(b[0]), .B(a[304]), .Z(n1519) );
  XOR U1825 ( .A(sreg[1327]), .B(n1519), .Z(n1521) );
  NANDN U1826 ( .A(n1514), .B(sreg[1326]), .Z(n1518) );
  OR U1827 ( .A(n1516), .B(n1515), .Z(n1517) );
  AND U1828 ( .A(n1518), .B(n1517), .Z(n1520) );
  XOR U1829 ( .A(n1521), .B(n1520), .Z(c[1327]) );
  NAND U1830 ( .A(b[0]), .B(a[305]), .Z(n1524) );
  XOR U1831 ( .A(sreg[1328]), .B(n1524), .Z(n1526) );
  NANDN U1832 ( .A(n1519), .B(sreg[1327]), .Z(n1523) );
  OR U1833 ( .A(n1521), .B(n1520), .Z(n1522) );
  AND U1834 ( .A(n1523), .B(n1522), .Z(n1525) );
  XOR U1835 ( .A(n1526), .B(n1525), .Z(c[1328]) );
  NAND U1836 ( .A(b[0]), .B(a[306]), .Z(n1529) );
  XOR U1837 ( .A(sreg[1329]), .B(n1529), .Z(n1531) );
  NANDN U1838 ( .A(n1524), .B(sreg[1328]), .Z(n1528) );
  OR U1839 ( .A(n1526), .B(n1525), .Z(n1527) );
  AND U1840 ( .A(n1528), .B(n1527), .Z(n1530) );
  XOR U1841 ( .A(n1531), .B(n1530), .Z(c[1329]) );
  NAND U1842 ( .A(b[0]), .B(a[307]), .Z(n1534) );
  XOR U1843 ( .A(sreg[1330]), .B(n1534), .Z(n1536) );
  NANDN U1844 ( .A(n1529), .B(sreg[1329]), .Z(n1533) );
  OR U1845 ( .A(n1531), .B(n1530), .Z(n1532) );
  AND U1846 ( .A(n1533), .B(n1532), .Z(n1535) );
  XOR U1847 ( .A(n1536), .B(n1535), .Z(c[1330]) );
  NAND U1848 ( .A(b[0]), .B(a[308]), .Z(n1539) );
  XOR U1849 ( .A(sreg[1331]), .B(n1539), .Z(n1541) );
  NANDN U1850 ( .A(n1534), .B(sreg[1330]), .Z(n1538) );
  OR U1851 ( .A(n1536), .B(n1535), .Z(n1537) );
  AND U1852 ( .A(n1538), .B(n1537), .Z(n1540) );
  XOR U1853 ( .A(n1541), .B(n1540), .Z(c[1331]) );
  NAND U1854 ( .A(b[0]), .B(a[309]), .Z(n1544) );
  XOR U1855 ( .A(sreg[1332]), .B(n1544), .Z(n1546) );
  NANDN U1856 ( .A(n1539), .B(sreg[1331]), .Z(n1543) );
  OR U1857 ( .A(n1541), .B(n1540), .Z(n1542) );
  AND U1858 ( .A(n1543), .B(n1542), .Z(n1545) );
  XOR U1859 ( .A(n1546), .B(n1545), .Z(c[1332]) );
  NAND U1860 ( .A(b[0]), .B(a[310]), .Z(n1549) );
  XOR U1861 ( .A(sreg[1333]), .B(n1549), .Z(n1551) );
  NANDN U1862 ( .A(n1544), .B(sreg[1332]), .Z(n1548) );
  OR U1863 ( .A(n1546), .B(n1545), .Z(n1547) );
  AND U1864 ( .A(n1548), .B(n1547), .Z(n1550) );
  XOR U1865 ( .A(n1551), .B(n1550), .Z(c[1333]) );
  NAND U1866 ( .A(b[0]), .B(a[311]), .Z(n1554) );
  XOR U1867 ( .A(sreg[1334]), .B(n1554), .Z(n1556) );
  NANDN U1868 ( .A(n1549), .B(sreg[1333]), .Z(n1553) );
  OR U1869 ( .A(n1551), .B(n1550), .Z(n1552) );
  AND U1870 ( .A(n1553), .B(n1552), .Z(n1555) );
  XOR U1871 ( .A(n1556), .B(n1555), .Z(c[1334]) );
  NAND U1872 ( .A(b[0]), .B(a[312]), .Z(n1559) );
  XOR U1873 ( .A(sreg[1335]), .B(n1559), .Z(n1561) );
  NANDN U1874 ( .A(n1554), .B(sreg[1334]), .Z(n1558) );
  OR U1875 ( .A(n1556), .B(n1555), .Z(n1557) );
  AND U1876 ( .A(n1558), .B(n1557), .Z(n1560) );
  XOR U1877 ( .A(n1561), .B(n1560), .Z(c[1335]) );
  NAND U1878 ( .A(b[0]), .B(a[313]), .Z(n1564) );
  XOR U1879 ( .A(sreg[1336]), .B(n1564), .Z(n1566) );
  NANDN U1880 ( .A(n1559), .B(sreg[1335]), .Z(n1563) );
  OR U1881 ( .A(n1561), .B(n1560), .Z(n1562) );
  AND U1882 ( .A(n1563), .B(n1562), .Z(n1565) );
  XOR U1883 ( .A(n1566), .B(n1565), .Z(c[1336]) );
  NAND U1884 ( .A(b[0]), .B(a[314]), .Z(n1569) );
  XOR U1885 ( .A(sreg[1337]), .B(n1569), .Z(n1571) );
  NANDN U1886 ( .A(n1564), .B(sreg[1336]), .Z(n1568) );
  OR U1887 ( .A(n1566), .B(n1565), .Z(n1567) );
  AND U1888 ( .A(n1568), .B(n1567), .Z(n1570) );
  XOR U1889 ( .A(n1571), .B(n1570), .Z(c[1337]) );
  NAND U1890 ( .A(b[0]), .B(a[315]), .Z(n1574) );
  XOR U1891 ( .A(sreg[1338]), .B(n1574), .Z(n1576) );
  NANDN U1892 ( .A(n1569), .B(sreg[1337]), .Z(n1573) );
  OR U1893 ( .A(n1571), .B(n1570), .Z(n1572) );
  AND U1894 ( .A(n1573), .B(n1572), .Z(n1575) );
  XOR U1895 ( .A(n1576), .B(n1575), .Z(c[1338]) );
  NAND U1896 ( .A(b[0]), .B(a[316]), .Z(n1579) );
  XOR U1897 ( .A(sreg[1339]), .B(n1579), .Z(n1581) );
  NANDN U1898 ( .A(n1574), .B(sreg[1338]), .Z(n1578) );
  OR U1899 ( .A(n1576), .B(n1575), .Z(n1577) );
  AND U1900 ( .A(n1578), .B(n1577), .Z(n1580) );
  XOR U1901 ( .A(n1581), .B(n1580), .Z(c[1339]) );
  NAND U1902 ( .A(b[0]), .B(a[317]), .Z(n1584) );
  XOR U1903 ( .A(sreg[1340]), .B(n1584), .Z(n1586) );
  NANDN U1904 ( .A(n1579), .B(sreg[1339]), .Z(n1583) );
  OR U1905 ( .A(n1581), .B(n1580), .Z(n1582) );
  AND U1906 ( .A(n1583), .B(n1582), .Z(n1585) );
  XOR U1907 ( .A(n1586), .B(n1585), .Z(c[1340]) );
  NAND U1908 ( .A(b[0]), .B(a[318]), .Z(n1589) );
  XOR U1909 ( .A(sreg[1341]), .B(n1589), .Z(n1591) );
  NANDN U1910 ( .A(n1584), .B(sreg[1340]), .Z(n1588) );
  OR U1911 ( .A(n1586), .B(n1585), .Z(n1587) );
  AND U1912 ( .A(n1588), .B(n1587), .Z(n1590) );
  XOR U1913 ( .A(n1591), .B(n1590), .Z(c[1341]) );
  NAND U1914 ( .A(b[0]), .B(a[319]), .Z(n1594) );
  XOR U1915 ( .A(sreg[1342]), .B(n1594), .Z(n1596) );
  NANDN U1916 ( .A(n1589), .B(sreg[1341]), .Z(n1593) );
  OR U1917 ( .A(n1591), .B(n1590), .Z(n1592) );
  AND U1918 ( .A(n1593), .B(n1592), .Z(n1595) );
  XOR U1919 ( .A(n1596), .B(n1595), .Z(c[1342]) );
  NAND U1920 ( .A(b[0]), .B(a[320]), .Z(n1599) );
  XOR U1921 ( .A(sreg[1343]), .B(n1599), .Z(n1601) );
  NANDN U1922 ( .A(n1594), .B(sreg[1342]), .Z(n1598) );
  OR U1923 ( .A(n1596), .B(n1595), .Z(n1597) );
  AND U1924 ( .A(n1598), .B(n1597), .Z(n1600) );
  XOR U1925 ( .A(n1601), .B(n1600), .Z(c[1343]) );
  NAND U1926 ( .A(b[0]), .B(a[321]), .Z(n1604) );
  XOR U1927 ( .A(sreg[1344]), .B(n1604), .Z(n1606) );
  NANDN U1928 ( .A(n1599), .B(sreg[1343]), .Z(n1603) );
  OR U1929 ( .A(n1601), .B(n1600), .Z(n1602) );
  AND U1930 ( .A(n1603), .B(n1602), .Z(n1605) );
  XOR U1931 ( .A(n1606), .B(n1605), .Z(c[1344]) );
  NAND U1932 ( .A(b[0]), .B(a[322]), .Z(n1609) );
  XOR U1933 ( .A(sreg[1345]), .B(n1609), .Z(n1611) );
  NANDN U1934 ( .A(n1604), .B(sreg[1344]), .Z(n1608) );
  OR U1935 ( .A(n1606), .B(n1605), .Z(n1607) );
  AND U1936 ( .A(n1608), .B(n1607), .Z(n1610) );
  XOR U1937 ( .A(n1611), .B(n1610), .Z(c[1345]) );
  NAND U1938 ( .A(b[0]), .B(a[323]), .Z(n1614) );
  XOR U1939 ( .A(sreg[1346]), .B(n1614), .Z(n1616) );
  NANDN U1940 ( .A(n1609), .B(sreg[1345]), .Z(n1613) );
  OR U1941 ( .A(n1611), .B(n1610), .Z(n1612) );
  AND U1942 ( .A(n1613), .B(n1612), .Z(n1615) );
  XOR U1943 ( .A(n1616), .B(n1615), .Z(c[1346]) );
  NAND U1944 ( .A(b[0]), .B(a[324]), .Z(n1619) );
  XOR U1945 ( .A(sreg[1347]), .B(n1619), .Z(n1621) );
  NANDN U1946 ( .A(n1614), .B(sreg[1346]), .Z(n1618) );
  OR U1947 ( .A(n1616), .B(n1615), .Z(n1617) );
  AND U1948 ( .A(n1618), .B(n1617), .Z(n1620) );
  XOR U1949 ( .A(n1621), .B(n1620), .Z(c[1347]) );
  NAND U1950 ( .A(b[0]), .B(a[325]), .Z(n1624) );
  XOR U1951 ( .A(sreg[1348]), .B(n1624), .Z(n1626) );
  NANDN U1952 ( .A(n1619), .B(sreg[1347]), .Z(n1623) );
  OR U1953 ( .A(n1621), .B(n1620), .Z(n1622) );
  AND U1954 ( .A(n1623), .B(n1622), .Z(n1625) );
  XOR U1955 ( .A(n1626), .B(n1625), .Z(c[1348]) );
  NAND U1956 ( .A(b[0]), .B(a[326]), .Z(n1629) );
  XOR U1957 ( .A(sreg[1349]), .B(n1629), .Z(n1631) );
  NANDN U1958 ( .A(n1624), .B(sreg[1348]), .Z(n1628) );
  OR U1959 ( .A(n1626), .B(n1625), .Z(n1627) );
  AND U1960 ( .A(n1628), .B(n1627), .Z(n1630) );
  XOR U1961 ( .A(n1631), .B(n1630), .Z(c[1349]) );
  NAND U1962 ( .A(b[0]), .B(a[327]), .Z(n1634) );
  XOR U1963 ( .A(sreg[1350]), .B(n1634), .Z(n1636) );
  NANDN U1964 ( .A(n1629), .B(sreg[1349]), .Z(n1633) );
  OR U1965 ( .A(n1631), .B(n1630), .Z(n1632) );
  AND U1966 ( .A(n1633), .B(n1632), .Z(n1635) );
  XOR U1967 ( .A(n1636), .B(n1635), .Z(c[1350]) );
  NAND U1968 ( .A(b[0]), .B(a[328]), .Z(n1639) );
  XOR U1969 ( .A(sreg[1351]), .B(n1639), .Z(n1641) );
  NANDN U1970 ( .A(n1634), .B(sreg[1350]), .Z(n1638) );
  OR U1971 ( .A(n1636), .B(n1635), .Z(n1637) );
  AND U1972 ( .A(n1638), .B(n1637), .Z(n1640) );
  XOR U1973 ( .A(n1641), .B(n1640), .Z(c[1351]) );
  NAND U1974 ( .A(b[0]), .B(a[329]), .Z(n1644) );
  XOR U1975 ( .A(sreg[1352]), .B(n1644), .Z(n1646) );
  NANDN U1976 ( .A(n1639), .B(sreg[1351]), .Z(n1643) );
  OR U1977 ( .A(n1641), .B(n1640), .Z(n1642) );
  AND U1978 ( .A(n1643), .B(n1642), .Z(n1645) );
  XOR U1979 ( .A(n1646), .B(n1645), .Z(c[1352]) );
  NAND U1980 ( .A(b[0]), .B(a[330]), .Z(n1649) );
  XOR U1981 ( .A(sreg[1353]), .B(n1649), .Z(n1651) );
  NANDN U1982 ( .A(n1644), .B(sreg[1352]), .Z(n1648) );
  OR U1983 ( .A(n1646), .B(n1645), .Z(n1647) );
  AND U1984 ( .A(n1648), .B(n1647), .Z(n1650) );
  XOR U1985 ( .A(n1651), .B(n1650), .Z(c[1353]) );
  NAND U1986 ( .A(b[0]), .B(a[331]), .Z(n1654) );
  XOR U1987 ( .A(sreg[1354]), .B(n1654), .Z(n1656) );
  NANDN U1988 ( .A(n1649), .B(sreg[1353]), .Z(n1653) );
  OR U1989 ( .A(n1651), .B(n1650), .Z(n1652) );
  AND U1990 ( .A(n1653), .B(n1652), .Z(n1655) );
  XOR U1991 ( .A(n1656), .B(n1655), .Z(c[1354]) );
  NAND U1992 ( .A(b[0]), .B(a[332]), .Z(n1659) );
  XOR U1993 ( .A(sreg[1355]), .B(n1659), .Z(n1661) );
  NANDN U1994 ( .A(n1654), .B(sreg[1354]), .Z(n1658) );
  OR U1995 ( .A(n1656), .B(n1655), .Z(n1657) );
  AND U1996 ( .A(n1658), .B(n1657), .Z(n1660) );
  XOR U1997 ( .A(n1661), .B(n1660), .Z(c[1355]) );
  NAND U1998 ( .A(b[0]), .B(a[333]), .Z(n1664) );
  XOR U1999 ( .A(sreg[1356]), .B(n1664), .Z(n1666) );
  NANDN U2000 ( .A(n1659), .B(sreg[1355]), .Z(n1663) );
  OR U2001 ( .A(n1661), .B(n1660), .Z(n1662) );
  AND U2002 ( .A(n1663), .B(n1662), .Z(n1665) );
  XOR U2003 ( .A(n1666), .B(n1665), .Z(c[1356]) );
  NAND U2004 ( .A(b[0]), .B(a[334]), .Z(n1669) );
  XOR U2005 ( .A(sreg[1357]), .B(n1669), .Z(n1671) );
  NANDN U2006 ( .A(n1664), .B(sreg[1356]), .Z(n1668) );
  OR U2007 ( .A(n1666), .B(n1665), .Z(n1667) );
  AND U2008 ( .A(n1668), .B(n1667), .Z(n1670) );
  XOR U2009 ( .A(n1671), .B(n1670), .Z(c[1357]) );
  NAND U2010 ( .A(b[0]), .B(a[335]), .Z(n1674) );
  XOR U2011 ( .A(sreg[1358]), .B(n1674), .Z(n1676) );
  NANDN U2012 ( .A(n1669), .B(sreg[1357]), .Z(n1673) );
  OR U2013 ( .A(n1671), .B(n1670), .Z(n1672) );
  AND U2014 ( .A(n1673), .B(n1672), .Z(n1675) );
  XOR U2015 ( .A(n1676), .B(n1675), .Z(c[1358]) );
  NAND U2016 ( .A(b[0]), .B(a[336]), .Z(n1679) );
  XOR U2017 ( .A(sreg[1359]), .B(n1679), .Z(n1681) );
  NANDN U2018 ( .A(n1674), .B(sreg[1358]), .Z(n1678) );
  OR U2019 ( .A(n1676), .B(n1675), .Z(n1677) );
  AND U2020 ( .A(n1678), .B(n1677), .Z(n1680) );
  XOR U2021 ( .A(n1681), .B(n1680), .Z(c[1359]) );
  NAND U2022 ( .A(b[0]), .B(a[337]), .Z(n1684) );
  XOR U2023 ( .A(sreg[1360]), .B(n1684), .Z(n1686) );
  NANDN U2024 ( .A(n1679), .B(sreg[1359]), .Z(n1683) );
  OR U2025 ( .A(n1681), .B(n1680), .Z(n1682) );
  AND U2026 ( .A(n1683), .B(n1682), .Z(n1685) );
  XOR U2027 ( .A(n1686), .B(n1685), .Z(c[1360]) );
  NAND U2028 ( .A(b[0]), .B(a[338]), .Z(n1689) );
  XOR U2029 ( .A(sreg[1361]), .B(n1689), .Z(n1691) );
  NANDN U2030 ( .A(n1684), .B(sreg[1360]), .Z(n1688) );
  OR U2031 ( .A(n1686), .B(n1685), .Z(n1687) );
  AND U2032 ( .A(n1688), .B(n1687), .Z(n1690) );
  XOR U2033 ( .A(n1691), .B(n1690), .Z(c[1361]) );
  NAND U2034 ( .A(b[0]), .B(a[339]), .Z(n1694) );
  XOR U2035 ( .A(sreg[1362]), .B(n1694), .Z(n1696) );
  NANDN U2036 ( .A(n1689), .B(sreg[1361]), .Z(n1693) );
  OR U2037 ( .A(n1691), .B(n1690), .Z(n1692) );
  AND U2038 ( .A(n1693), .B(n1692), .Z(n1695) );
  XOR U2039 ( .A(n1696), .B(n1695), .Z(c[1362]) );
  NAND U2040 ( .A(b[0]), .B(a[340]), .Z(n1699) );
  XOR U2041 ( .A(sreg[1363]), .B(n1699), .Z(n1701) );
  NANDN U2042 ( .A(n1694), .B(sreg[1362]), .Z(n1698) );
  OR U2043 ( .A(n1696), .B(n1695), .Z(n1697) );
  AND U2044 ( .A(n1698), .B(n1697), .Z(n1700) );
  XOR U2045 ( .A(n1701), .B(n1700), .Z(c[1363]) );
  NAND U2046 ( .A(b[0]), .B(a[341]), .Z(n1704) );
  XOR U2047 ( .A(sreg[1364]), .B(n1704), .Z(n1706) );
  NANDN U2048 ( .A(n1699), .B(sreg[1363]), .Z(n1703) );
  OR U2049 ( .A(n1701), .B(n1700), .Z(n1702) );
  AND U2050 ( .A(n1703), .B(n1702), .Z(n1705) );
  XOR U2051 ( .A(n1706), .B(n1705), .Z(c[1364]) );
  NAND U2052 ( .A(b[0]), .B(a[342]), .Z(n1709) );
  XOR U2053 ( .A(sreg[1365]), .B(n1709), .Z(n1711) );
  NANDN U2054 ( .A(n1704), .B(sreg[1364]), .Z(n1708) );
  OR U2055 ( .A(n1706), .B(n1705), .Z(n1707) );
  AND U2056 ( .A(n1708), .B(n1707), .Z(n1710) );
  XOR U2057 ( .A(n1711), .B(n1710), .Z(c[1365]) );
  NAND U2058 ( .A(b[0]), .B(a[343]), .Z(n1714) );
  XOR U2059 ( .A(sreg[1366]), .B(n1714), .Z(n1716) );
  NANDN U2060 ( .A(n1709), .B(sreg[1365]), .Z(n1713) );
  OR U2061 ( .A(n1711), .B(n1710), .Z(n1712) );
  AND U2062 ( .A(n1713), .B(n1712), .Z(n1715) );
  XOR U2063 ( .A(n1716), .B(n1715), .Z(c[1366]) );
  NAND U2064 ( .A(b[0]), .B(a[344]), .Z(n1719) );
  XOR U2065 ( .A(sreg[1367]), .B(n1719), .Z(n1721) );
  NANDN U2066 ( .A(n1714), .B(sreg[1366]), .Z(n1718) );
  OR U2067 ( .A(n1716), .B(n1715), .Z(n1717) );
  AND U2068 ( .A(n1718), .B(n1717), .Z(n1720) );
  XOR U2069 ( .A(n1721), .B(n1720), .Z(c[1367]) );
  NAND U2070 ( .A(b[0]), .B(a[345]), .Z(n1724) );
  XOR U2071 ( .A(sreg[1368]), .B(n1724), .Z(n1726) );
  NANDN U2072 ( .A(n1719), .B(sreg[1367]), .Z(n1723) );
  OR U2073 ( .A(n1721), .B(n1720), .Z(n1722) );
  AND U2074 ( .A(n1723), .B(n1722), .Z(n1725) );
  XOR U2075 ( .A(n1726), .B(n1725), .Z(c[1368]) );
  NAND U2076 ( .A(b[0]), .B(a[346]), .Z(n1729) );
  XOR U2077 ( .A(sreg[1369]), .B(n1729), .Z(n1731) );
  NANDN U2078 ( .A(n1724), .B(sreg[1368]), .Z(n1728) );
  OR U2079 ( .A(n1726), .B(n1725), .Z(n1727) );
  AND U2080 ( .A(n1728), .B(n1727), .Z(n1730) );
  XOR U2081 ( .A(n1731), .B(n1730), .Z(c[1369]) );
  NAND U2082 ( .A(b[0]), .B(a[347]), .Z(n1734) );
  XOR U2083 ( .A(sreg[1370]), .B(n1734), .Z(n1736) );
  NANDN U2084 ( .A(n1729), .B(sreg[1369]), .Z(n1733) );
  OR U2085 ( .A(n1731), .B(n1730), .Z(n1732) );
  AND U2086 ( .A(n1733), .B(n1732), .Z(n1735) );
  XOR U2087 ( .A(n1736), .B(n1735), .Z(c[1370]) );
  NAND U2088 ( .A(b[0]), .B(a[348]), .Z(n1739) );
  XOR U2089 ( .A(sreg[1371]), .B(n1739), .Z(n1741) );
  NANDN U2090 ( .A(n1734), .B(sreg[1370]), .Z(n1738) );
  OR U2091 ( .A(n1736), .B(n1735), .Z(n1737) );
  AND U2092 ( .A(n1738), .B(n1737), .Z(n1740) );
  XOR U2093 ( .A(n1741), .B(n1740), .Z(c[1371]) );
  NAND U2094 ( .A(b[0]), .B(a[349]), .Z(n1744) );
  XOR U2095 ( .A(sreg[1372]), .B(n1744), .Z(n1746) );
  NANDN U2096 ( .A(n1739), .B(sreg[1371]), .Z(n1743) );
  OR U2097 ( .A(n1741), .B(n1740), .Z(n1742) );
  AND U2098 ( .A(n1743), .B(n1742), .Z(n1745) );
  XOR U2099 ( .A(n1746), .B(n1745), .Z(c[1372]) );
  NAND U2100 ( .A(b[0]), .B(a[350]), .Z(n1749) );
  XOR U2101 ( .A(sreg[1373]), .B(n1749), .Z(n1751) );
  NANDN U2102 ( .A(n1744), .B(sreg[1372]), .Z(n1748) );
  OR U2103 ( .A(n1746), .B(n1745), .Z(n1747) );
  AND U2104 ( .A(n1748), .B(n1747), .Z(n1750) );
  XOR U2105 ( .A(n1751), .B(n1750), .Z(c[1373]) );
  NAND U2106 ( .A(b[0]), .B(a[351]), .Z(n1754) );
  XOR U2107 ( .A(sreg[1374]), .B(n1754), .Z(n1756) );
  NANDN U2108 ( .A(n1749), .B(sreg[1373]), .Z(n1753) );
  OR U2109 ( .A(n1751), .B(n1750), .Z(n1752) );
  AND U2110 ( .A(n1753), .B(n1752), .Z(n1755) );
  XOR U2111 ( .A(n1756), .B(n1755), .Z(c[1374]) );
  NAND U2112 ( .A(b[0]), .B(a[352]), .Z(n1759) );
  XOR U2113 ( .A(sreg[1375]), .B(n1759), .Z(n1761) );
  NANDN U2114 ( .A(n1754), .B(sreg[1374]), .Z(n1758) );
  OR U2115 ( .A(n1756), .B(n1755), .Z(n1757) );
  AND U2116 ( .A(n1758), .B(n1757), .Z(n1760) );
  XOR U2117 ( .A(n1761), .B(n1760), .Z(c[1375]) );
  NAND U2118 ( .A(b[0]), .B(a[353]), .Z(n1764) );
  XOR U2119 ( .A(sreg[1376]), .B(n1764), .Z(n1766) );
  NANDN U2120 ( .A(n1759), .B(sreg[1375]), .Z(n1763) );
  OR U2121 ( .A(n1761), .B(n1760), .Z(n1762) );
  AND U2122 ( .A(n1763), .B(n1762), .Z(n1765) );
  XOR U2123 ( .A(n1766), .B(n1765), .Z(c[1376]) );
  NAND U2124 ( .A(b[0]), .B(a[354]), .Z(n1769) );
  XOR U2125 ( .A(sreg[1377]), .B(n1769), .Z(n1771) );
  NANDN U2126 ( .A(n1764), .B(sreg[1376]), .Z(n1768) );
  OR U2127 ( .A(n1766), .B(n1765), .Z(n1767) );
  AND U2128 ( .A(n1768), .B(n1767), .Z(n1770) );
  XOR U2129 ( .A(n1771), .B(n1770), .Z(c[1377]) );
  NAND U2130 ( .A(b[0]), .B(a[355]), .Z(n1774) );
  XOR U2131 ( .A(sreg[1378]), .B(n1774), .Z(n1776) );
  NANDN U2132 ( .A(n1769), .B(sreg[1377]), .Z(n1773) );
  OR U2133 ( .A(n1771), .B(n1770), .Z(n1772) );
  AND U2134 ( .A(n1773), .B(n1772), .Z(n1775) );
  XOR U2135 ( .A(n1776), .B(n1775), .Z(c[1378]) );
  NAND U2136 ( .A(b[0]), .B(a[356]), .Z(n1779) );
  XOR U2137 ( .A(sreg[1379]), .B(n1779), .Z(n1781) );
  NANDN U2138 ( .A(n1774), .B(sreg[1378]), .Z(n1778) );
  OR U2139 ( .A(n1776), .B(n1775), .Z(n1777) );
  AND U2140 ( .A(n1778), .B(n1777), .Z(n1780) );
  XOR U2141 ( .A(n1781), .B(n1780), .Z(c[1379]) );
  NAND U2142 ( .A(b[0]), .B(a[357]), .Z(n1784) );
  XOR U2143 ( .A(sreg[1380]), .B(n1784), .Z(n1786) );
  NANDN U2144 ( .A(n1779), .B(sreg[1379]), .Z(n1783) );
  OR U2145 ( .A(n1781), .B(n1780), .Z(n1782) );
  AND U2146 ( .A(n1783), .B(n1782), .Z(n1785) );
  XOR U2147 ( .A(n1786), .B(n1785), .Z(c[1380]) );
  NAND U2148 ( .A(b[0]), .B(a[358]), .Z(n1789) );
  XOR U2149 ( .A(sreg[1381]), .B(n1789), .Z(n1791) );
  NANDN U2150 ( .A(n1784), .B(sreg[1380]), .Z(n1788) );
  OR U2151 ( .A(n1786), .B(n1785), .Z(n1787) );
  AND U2152 ( .A(n1788), .B(n1787), .Z(n1790) );
  XOR U2153 ( .A(n1791), .B(n1790), .Z(c[1381]) );
  NAND U2154 ( .A(b[0]), .B(a[359]), .Z(n1794) );
  XOR U2155 ( .A(sreg[1382]), .B(n1794), .Z(n1796) );
  NANDN U2156 ( .A(n1789), .B(sreg[1381]), .Z(n1793) );
  OR U2157 ( .A(n1791), .B(n1790), .Z(n1792) );
  AND U2158 ( .A(n1793), .B(n1792), .Z(n1795) );
  XOR U2159 ( .A(n1796), .B(n1795), .Z(c[1382]) );
  NAND U2160 ( .A(b[0]), .B(a[360]), .Z(n1799) );
  XOR U2161 ( .A(sreg[1383]), .B(n1799), .Z(n1801) );
  NANDN U2162 ( .A(n1794), .B(sreg[1382]), .Z(n1798) );
  OR U2163 ( .A(n1796), .B(n1795), .Z(n1797) );
  AND U2164 ( .A(n1798), .B(n1797), .Z(n1800) );
  XOR U2165 ( .A(n1801), .B(n1800), .Z(c[1383]) );
  NAND U2166 ( .A(b[0]), .B(a[361]), .Z(n1804) );
  XOR U2167 ( .A(sreg[1384]), .B(n1804), .Z(n1806) );
  NANDN U2168 ( .A(n1799), .B(sreg[1383]), .Z(n1803) );
  OR U2169 ( .A(n1801), .B(n1800), .Z(n1802) );
  AND U2170 ( .A(n1803), .B(n1802), .Z(n1805) );
  XOR U2171 ( .A(n1806), .B(n1805), .Z(c[1384]) );
  NAND U2172 ( .A(b[0]), .B(a[362]), .Z(n1809) );
  XOR U2173 ( .A(sreg[1385]), .B(n1809), .Z(n1811) );
  NANDN U2174 ( .A(n1804), .B(sreg[1384]), .Z(n1808) );
  OR U2175 ( .A(n1806), .B(n1805), .Z(n1807) );
  AND U2176 ( .A(n1808), .B(n1807), .Z(n1810) );
  XOR U2177 ( .A(n1811), .B(n1810), .Z(c[1385]) );
  NAND U2178 ( .A(b[0]), .B(a[363]), .Z(n1814) );
  XOR U2179 ( .A(sreg[1386]), .B(n1814), .Z(n1816) );
  NANDN U2180 ( .A(n1809), .B(sreg[1385]), .Z(n1813) );
  OR U2181 ( .A(n1811), .B(n1810), .Z(n1812) );
  AND U2182 ( .A(n1813), .B(n1812), .Z(n1815) );
  XOR U2183 ( .A(n1816), .B(n1815), .Z(c[1386]) );
  NAND U2184 ( .A(b[0]), .B(a[364]), .Z(n1819) );
  XOR U2185 ( .A(sreg[1387]), .B(n1819), .Z(n1821) );
  NANDN U2186 ( .A(n1814), .B(sreg[1386]), .Z(n1818) );
  OR U2187 ( .A(n1816), .B(n1815), .Z(n1817) );
  AND U2188 ( .A(n1818), .B(n1817), .Z(n1820) );
  XOR U2189 ( .A(n1821), .B(n1820), .Z(c[1387]) );
  NAND U2190 ( .A(b[0]), .B(a[365]), .Z(n1824) );
  XOR U2191 ( .A(sreg[1388]), .B(n1824), .Z(n1826) );
  NANDN U2192 ( .A(n1819), .B(sreg[1387]), .Z(n1823) );
  OR U2193 ( .A(n1821), .B(n1820), .Z(n1822) );
  AND U2194 ( .A(n1823), .B(n1822), .Z(n1825) );
  XOR U2195 ( .A(n1826), .B(n1825), .Z(c[1388]) );
  NAND U2196 ( .A(b[0]), .B(a[366]), .Z(n1829) );
  XOR U2197 ( .A(sreg[1389]), .B(n1829), .Z(n1831) );
  NANDN U2198 ( .A(n1824), .B(sreg[1388]), .Z(n1828) );
  OR U2199 ( .A(n1826), .B(n1825), .Z(n1827) );
  AND U2200 ( .A(n1828), .B(n1827), .Z(n1830) );
  XOR U2201 ( .A(n1831), .B(n1830), .Z(c[1389]) );
  NAND U2202 ( .A(b[0]), .B(a[367]), .Z(n1834) );
  XOR U2203 ( .A(sreg[1390]), .B(n1834), .Z(n1836) );
  NANDN U2204 ( .A(n1829), .B(sreg[1389]), .Z(n1833) );
  OR U2205 ( .A(n1831), .B(n1830), .Z(n1832) );
  AND U2206 ( .A(n1833), .B(n1832), .Z(n1835) );
  XOR U2207 ( .A(n1836), .B(n1835), .Z(c[1390]) );
  NAND U2208 ( .A(b[0]), .B(a[368]), .Z(n1839) );
  XOR U2209 ( .A(sreg[1391]), .B(n1839), .Z(n1841) );
  NANDN U2210 ( .A(n1834), .B(sreg[1390]), .Z(n1838) );
  OR U2211 ( .A(n1836), .B(n1835), .Z(n1837) );
  AND U2212 ( .A(n1838), .B(n1837), .Z(n1840) );
  XOR U2213 ( .A(n1841), .B(n1840), .Z(c[1391]) );
  NAND U2214 ( .A(b[0]), .B(a[369]), .Z(n1844) );
  XOR U2215 ( .A(sreg[1392]), .B(n1844), .Z(n1846) );
  NANDN U2216 ( .A(n1839), .B(sreg[1391]), .Z(n1843) );
  OR U2217 ( .A(n1841), .B(n1840), .Z(n1842) );
  AND U2218 ( .A(n1843), .B(n1842), .Z(n1845) );
  XOR U2219 ( .A(n1846), .B(n1845), .Z(c[1392]) );
  NAND U2220 ( .A(b[0]), .B(a[370]), .Z(n1849) );
  XOR U2221 ( .A(sreg[1393]), .B(n1849), .Z(n1851) );
  NANDN U2222 ( .A(n1844), .B(sreg[1392]), .Z(n1848) );
  OR U2223 ( .A(n1846), .B(n1845), .Z(n1847) );
  AND U2224 ( .A(n1848), .B(n1847), .Z(n1850) );
  XOR U2225 ( .A(n1851), .B(n1850), .Z(c[1393]) );
  NAND U2226 ( .A(b[0]), .B(a[371]), .Z(n1854) );
  XOR U2227 ( .A(sreg[1394]), .B(n1854), .Z(n1856) );
  NANDN U2228 ( .A(n1849), .B(sreg[1393]), .Z(n1853) );
  OR U2229 ( .A(n1851), .B(n1850), .Z(n1852) );
  AND U2230 ( .A(n1853), .B(n1852), .Z(n1855) );
  XOR U2231 ( .A(n1856), .B(n1855), .Z(c[1394]) );
  NAND U2232 ( .A(b[0]), .B(a[372]), .Z(n1859) );
  XOR U2233 ( .A(sreg[1395]), .B(n1859), .Z(n1861) );
  NANDN U2234 ( .A(n1854), .B(sreg[1394]), .Z(n1858) );
  OR U2235 ( .A(n1856), .B(n1855), .Z(n1857) );
  AND U2236 ( .A(n1858), .B(n1857), .Z(n1860) );
  XOR U2237 ( .A(n1861), .B(n1860), .Z(c[1395]) );
  NAND U2238 ( .A(b[0]), .B(a[373]), .Z(n1864) );
  XOR U2239 ( .A(sreg[1396]), .B(n1864), .Z(n1866) );
  NANDN U2240 ( .A(n1859), .B(sreg[1395]), .Z(n1863) );
  OR U2241 ( .A(n1861), .B(n1860), .Z(n1862) );
  AND U2242 ( .A(n1863), .B(n1862), .Z(n1865) );
  XOR U2243 ( .A(n1866), .B(n1865), .Z(c[1396]) );
  NAND U2244 ( .A(b[0]), .B(a[374]), .Z(n1869) );
  XOR U2245 ( .A(sreg[1397]), .B(n1869), .Z(n1871) );
  NANDN U2246 ( .A(n1864), .B(sreg[1396]), .Z(n1868) );
  OR U2247 ( .A(n1866), .B(n1865), .Z(n1867) );
  AND U2248 ( .A(n1868), .B(n1867), .Z(n1870) );
  XOR U2249 ( .A(n1871), .B(n1870), .Z(c[1397]) );
  NAND U2250 ( .A(b[0]), .B(a[375]), .Z(n1874) );
  XOR U2251 ( .A(sreg[1398]), .B(n1874), .Z(n1876) );
  NANDN U2252 ( .A(n1869), .B(sreg[1397]), .Z(n1873) );
  OR U2253 ( .A(n1871), .B(n1870), .Z(n1872) );
  AND U2254 ( .A(n1873), .B(n1872), .Z(n1875) );
  XOR U2255 ( .A(n1876), .B(n1875), .Z(c[1398]) );
  NAND U2256 ( .A(b[0]), .B(a[376]), .Z(n1879) );
  XOR U2257 ( .A(sreg[1399]), .B(n1879), .Z(n1881) );
  NANDN U2258 ( .A(n1874), .B(sreg[1398]), .Z(n1878) );
  OR U2259 ( .A(n1876), .B(n1875), .Z(n1877) );
  AND U2260 ( .A(n1878), .B(n1877), .Z(n1880) );
  XOR U2261 ( .A(n1881), .B(n1880), .Z(c[1399]) );
  NAND U2262 ( .A(b[0]), .B(a[377]), .Z(n1884) );
  XOR U2263 ( .A(sreg[1400]), .B(n1884), .Z(n1886) );
  NANDN U2264 ( .A(n1879), .B(sreg[1399]), .Z(n1883) );
  OR U2265 ( .A(n1881), .B(n1880), .Z(n1882) );
  AND U2266 ( .A(n1883), .B(n1882), .Z(n1885) );
  XOR U2267 ( .A(n1886), .B(n1885), .Z(c[1400]) );
  NAND U2268 ( .A(b[0]), .B(a[378]), .Z(n1889) );
  XOR U2269 ( .A(sreg[1401]), .B(n1889), .Z(n1891) );
  NANDN U2270 ( .A(n1884), .B(sreg[1400]), .Z(n1888) );
  OR U2271 ( .A(n1886), .B(n1885), .Z(n1887) );
  AND U2272 ( .A(n1888), .B(n1887), .Z(n1890) );
  XOR U2273 ( .A(n1891), .B(n1890), .Z(c[1401]) );
  NAND U2274 ( .A(b[0]), .B(a[379]), .Z(n1894) );
  XOR U2275 ( .A(sreg[1402]), .B(n1894), .Z(n1896) );
  NANDN U2276 ( .A(n1889), .B(sreg[1401]), .Z(n1893) );
  OR U2277 ( .A(n1891), .B(n1890), .Z(n1892) );
  AND U2278 ( .A(n1893), .B(n1892), .Z(n1895) );
  XOR U2279 ( .A(n1896), .B(n1895), .Z(c[1402]) );
  NAND U2280 ( .A(b[0]), .B(a[380]), .Z(n1899) );
  XOR U2281 ( .A(sreg[1403]), .B(n1899), .Z(n1901) );
  NANDN U2282 ( .A(n1894), .B(sreg[1402]), .Z(n1898) );
  OR U2283 ( .A(n1896), .B(n1895), .Z(n1897) );
  AND U2284 ( .A(n1898), .B(n1897), .Z(n1900) );
  XOR U2285 ( .A(n1901), .B(n1900), .Z(c[1403]) );
  NAND U2286 ( .A(b[0]), .B(a[381]), .Z(n1904) );
  XOR U2287 ( .A(sreg[1404]), .B(n1904), .Z(n1906) );
  NANDN U2288 ( .A(n1899), .B(sreg[1403]), .Z(n1903) );
  OR U2289 ( .A(n1901), .B(n1900), .Z(n1902) );
  AND U2290 ( .A(n1903), .B(n1902), .Z(n1905) );
  XOR U2291 ( .A(n1906), .B(n1905), .Z(c[1404]) );
  NAND U2292 ( .A(b[0]), .B(a[382]), .Z(n1909) );
  XOR U2293 ( .A(sreg[1405]), .B(n1909), .Z(n1911) );
  NANDN U2294 ( .A(n1904), .B(sreg[1404]), .Z(n1908) );
  OR U2295 ( .A(n1906), .B(n1905), .Z(n1907) );
  AND U2296 ( .A(n1908), .B(n1907), .Z(n1910) );
  XOR U2297 ( .A(n1911), .B(n1910), .Z(c[1405]) );
  NAND U2298 ( .A(b[0]), .B(a[383]), .Z(n1914) );
  XOR U2299 ( .A(sreg[1406]), .B(n1914), .Z(n1916) );
  NANDN U2300 ( .A(n1909), .B(sreg[1405]), .Z(n1913) );
  OR U2301 ( .A(n1911), .B(n1910), .Z(n1912) );
  AND U2302 ( .A(n1913), .B(n1912), .Z(n1915) );
  XOR U2303 ( .A(n1916), .B(n1915), .Z(c[1406]) );
  NAND U2304 ( .A(b[0]), .B(a[384]), .Z(n1919) );
  XOR U2305 ( .A(sreg[1407]), .B(n1919), .Z(n1921) );
  NANDN U2306 ( .A(n1914), .B(sreg[1406]), .Z(n1918) );
  OR U2307 ( .A(n1916), .B(n1915), .Z(n1917) );
  AND U2308 ( .A(n1918), .B(n1917), .Z(n1920) );
  XOR U2309 ( .A(n1921), .B(n1920), .Z(c[1407]) );
  NAND U2310 ( .A(b[0]), .B(a[385]), .Z(n1924) );
  XOR U2311 ( .A(sreg[1408]), .B(n1924), .Z(n1926) );
  NANDN U2312 ( .A(n1919), .B(sreg[1407]), .Z(n1923) );
  OR U2313 ( .A(n1921), .B(n1920), .Z(n1922) );
  AND U2314 ( .A(n1923), .B(n1922), .Z(n1925) );
  XOR U2315 ( .A(n1926), .B(n1925), .Z(c[1408]) );
  NAND U2316 ( .A(b[0]), .B(a[386]), .Z(n1929) );
  XOR U2317 ( .A(sreg[1409]), .B(n1929), .Z(n1931) );
  NANDN U2318 ( .A(n1924), .B(sreg[1408]), .Z(n1928) );
  OR U2319 ( .A(n1926), .B(n1925), .Z(n1927) );
  AND U2320 ( .A(n1928), .B(n1927), .Z(n1930) );
  XOR U2321 ( .A(n1931), .B(n1930), .Z(c[1409]) );
  NAND U2322 ( .A(b[0]), .B(a[387]), .Z(n1934) );
  XOR U2323 ( .A(sreg[1410]), .B(n1934), .Z(n1936) );
  NANDN U2324 ( .A(n1929), .B(sreg[1409]), .Z(n1933) );
  OR U2325 ( .A(n1931), .B(n1930), .Z(n1932) );
  AND U2326 ( .A(n1933), .B(n1932), .Z(n1935) );
  XOR U2327 ( .A(n1936), .B(n1935), .Z(c[1410]) );
  NAND U2328 ( .A(b[0]), .B(a[388]), .Z(n1939) );
  XOR U2329 ( .A(sreg[1411]), .B(n1939), .Z(n1941) );
  NANDN U2330 ( .A(n1934), .B(sreg[1410]), .Z(n1938) );
  OR U2331 ( .A(n1936), .B(n1935), .Z(n1937) );
  AND U2332 ( .A(n1938), .B(n1937), .Z(n1940) );
  XOR U2333 ( .A(n1941), .B(n1940), .Z(c[1411]) );
  NAND U2334 ( .A(b[0]), .B(a[389]), .Z(n1944) );
  XOR U2335 ( .A(sreg[1412]), .B(n1944), .Z(n1946) );
  NANDN U2336 ( .A(n1939), .B(sreg[1411]), .Z(n1943) );
  OR U2337 ( .A(n1941), .B(n1940), .Z(n1942) );
  AND U2338 ( .A(n1943), .B(n1942), .Z(n1945) );
  XOR U2339 ( .A(n1946), .B(n1945), .Z(c[1412]) );
  NAND U2340 ( .A(b[0]), .B(a[390]), .Z(n1949) );
  XOR U2341 ( .A(sreg[1413]), .B(n1949), .Z(n1951) );
  NANDN U2342 ( .A(n1944), .B(sreg[1412]), .Z(n1948) );
  OR U2343 ( .A(n1946), .B(n1945), .Z(n1947) );
  AND U2344 ( .A(n1948), .B(n1947), .Z(n1950) );
  XOR U2345 ( .A(n1951), .B(n1950), .Z(c[1413]) );
  NAND U2346 ( .A(b[0]), .B(a[391]), .Z(n1954) );
  XOR U2347 ( .A(sreg[1414]), .B(n1954), .Z(n1956) );
  NANDN U2348 ( .A(n1949), .B(sreg[1413]), .Z(n1953) );
  OR U2349 ( .A(n1951), .B(n1950), .Z(n1952) );
  AND U2350 ( .A(n1953), .B(n1952), .Z(n1955) );
  XOR U2351 ( .A(n1956), .B(n1955), .Z(c[1414]) );
  NAND U2352 ( .A(b[0]), .B(a[392]), .Z(n1959) );
  XOR U2353 ( .A(sreg[1415]), .B(n1959), .Z(n1961) );
  NANDN U2354 ( .A(n1954), .B(sreg[1414]), .Z(n1958) );
  OR U2355 ( .A(n1956), .B(n1955), .Z(n1957) );
  AND U2356 ( .A(n1958), .B(n1957), .Z(n1960) );
  XOR U2357 ( .A(n1961), .B(n1960), .Z(c[1415]) );
  NAND U2358 ( .A(b[0]), .B(a[393]), .Z(n1964) );
  XOR U2359 ( .A(sreg[1416]), .B(n1964), .Z(n1966) );
  NANDN U2360 ( .A(n1959), .B(sreg[1415]), .Z(n1963) );
  OR U2361 ( .A(n1961), .B(n1960), .Z(n1962) );
  AND U2362 ( .A(n1963), .B(n1962), .Z(n1965) );
  XOR U2363 ( .A(n1966), .B(n1965), .Z(c[1416]) );
  NAND U2364 ( .A(b[0]), .B(a[394]), .Z(n1969) );
  XOR U2365 ( .A(sreg[1417]), .B(n1969), .Z(n1971) );
  NANDN U2366 ( .A(n1964), .B(sreg[1416]), .Z(n1968) );
  OR U2367 ( .A(n1966), .B(n1965), .Z(n1967) );
  AND U2368 ( .A(n1968), .B(n1967), .Z(n1970) );
  XOR U2369 ( .A(n1971), .B(n1970), .Z(c[1417]) );
  NAND U2370 ( .A(b[0]), .B(a[395]), .Z(n1974) );
  XOR U2371 ( .A(sreg[1418]), .B(n1974), .Z(n1976) );
  NANDN U2372 ( .A(n1969), .B(sreg[1417]), .Z(n1973) );
  OR U2373 ( .A(n1971), .B(n1970), .Z(n1972) );
  AND U2374 ( .A(n1973), .B(n1972), .Z(n1975) );
  XOR U2375 ( .A(n1976), .B(n1975), .Z(c[1418]) );
  NAND U2376 ( .A(b[0]), .B(a[396]), .Z(n1979) );
  XOR U2377 ( .A(sreg[1419]), .B(n1979), .Z(n1981) );
  NANDN U2378 ( .A(n1974), .B(sreg[1418]), .Z(n1978) );
  OR U2379 ( .A(n1976), .B(n1975), .Z(n1977) );
  AND U2380 ( .A(n1978), .B(n1977), .Z(n1980) );
  XOR U2381 ( .A(n1981), .B(n1980), .Z(c[1419]) );
  NAND U2382 ( .A(b[0]), .B(a[397]), .Z(n1984) );
  XOR U2383 ( .A(sreg[1420]), .B(n1984), .Z(n1986) );
  NANDN U2384 ( .A(n1979), .B(sreg[1419]), .Z(n1983) );
  OR U2385 ( .A(n1981), .B(n1980), .Z(n1982) );
  AND U2386 ( .A(n1983), .B(n1982), .Z(n1985) );
  XOR U2387 ( .A(n1986), .B(n1985), .Z(c[1420]) );
  NAND U2388 ( .A(b[0]), .B(a[398]), .Z(n1989) );
  XOR U2389 ( .A(sreg[1421]), .B(n1989), .Z(n1991) );
  NANDN U2390 ( .A(n1984), .B(sreg[1420]), .Z(n1988) );
  OR U2391 ( .A(n1986), .B(n1985), .Z(n1987) );
  AND U2392 ( .A(n1988), .B(n1987), .Z(n1990) );
  XOR U2393 ( .A(n1991), .B(n1990), .Z(c[1421]) );
  NAND U2394 ( .A(b[0]), .B(a[399]), .Z(n1994) );
  XOR U2395 ( .A(sreg[1422]), .B(n1994), .Z(n1996) );
  NANDN U2396 ( .A(n1989), .B(sreg[1421]), .Z(n1993) );
  OR U2397 ( .A(n1991), .B(n1990), .Z(n1992) );
  AND U2398 ( .A(n1993), .B(n1992), .Z(n1995) );
  XOR U2399 ( .A(n1996), .B(n1995), .Z(c[1422]) );
  NAND U2400 ( .A(b[0]), .B(a[400]), .Z(n1999) );
  XOR U2401 ( .A(sreg[1423]), .B(n1999), .Z(n2001) );
  NANDN U2402 ( .A(n1994), .B(sreg[1422]), .Z(n1998) );
  OR U2403 ( .A(n1996), .B(n1995), .Z(n1997) );
  AND U2404 ( .A(n1998), .B(n1997), .Z(n2000) );
  XOR U2405 ( .A(n2001), .B(n2000), .Z(c[1423]) );
  NAND U2406 ( .A(b[0]), .B(a[401]), .Z(n2004) );
  XOR U2407 ( .A(sreg[1424]), .B(n2004), .Z(n2006) );
  NANDN U2408 ( .A(n1999), .B(sreg[1423]), .Z(n2003) );
  OR U2409 ( .A(n2001), .B(n2000), .Z(n2002) );
  AND U2410 ( .A(n2003), .B(n2002), .Z(n2005) );
  XOR U2411 ( .A(n2006), .B(n2005), .Z(c[1424]) );
  NAND U2412 ( .A(b[0]), .B(a[402]), .Z(n2009) );
  XOR U2413 ( .A(sreg[1425]), .B(n2009), .Z(n2011) );
  NANDN U2414 ( .A(n2004), .B(sreg[1424]), .Z(n2008) );
  OR U2415 ( .A(n2006), .B(n2005), .Z(n2007) );
  AND U2416 ( .A(n2008), .B(n2007), .Z(n2010) );
  XOR U2417 ( .A(n2011), .B(n2010), .Z(c[1425]) );
  NAND U2418 ( .A(b[0]), .B(a[403]), .Z(n2014) );
  XOR U2419 ( .A(sreg[1426]), .B(n2014), .Z(n2016) );
  NANDN U2420 ( .A(n2009), .B(sreg[1425]), .Z(n2013) );
  OR U2421 ( .A(n2011), .B(n2010), .Z(n2012) );
  AND U2422 ( .A(n2013), .B(n2012), .Z(n2015) );
  XOR U2423 ( .A(n2016), .B(n2015), .Z(c[1426]) );
  NAND U2424 ( .A(b[0]), .B(a[404]), .Z(n2019) );
  XOR U2425 ( .A(sreg[1427]), .B(n2019), .Z(n2021) );
  NANDN U2426 ( .A(n2014), .B(sreg[1426]), .Z(n2018) );
  OR U2427 ( .A(n2016), .B(n2015), .Z(n2017) );
  AND U2428 ( .A(n2018), .B(n2017), .Z(n2020) );
  XOR U2429 ( .A(n2021), .B(n2020), .Z(c[1427]) );
  NAND U2430 ( .A(b[0]), .B(a[405]), .Z(n2024) );
  XOR U2431 ( .A(sreg[1428]), .B(n2024), .Z(n2026) );
  NANDN U2432 ( .A(n2019), .B(sreg[1427]), .Z(n2023) );
  OR U2433 ( .A(n2021), .B(n2020), .Z(n2022) );
  AND U2434 ( .A(n2023), .B(n2022), .Z(n2025) );
  XOR U2435 ( .A(n2026), .B(n2025), .Z(c[1428]) );
  NAND U2436 ( .A(b[0]), .B(a[406]), .Z(n2029) );
  XOR U2437 ( .A(sreg[1429]), .B(n2029), .Z(n2031) );
  NANDN U2438 ( .A(n2024), .B(sreg[1428]), .Z(n2028) );
  OR U2439 ( .A(n2026), .B(n2025), .Z(n2027) );
  AND U2440 ( .A(n2028), .B(n2027), .Z(n2030) );
  XOR U2441 ( .A(n2031), .B(n2030), .Z(c[1429]) );
  NAND U2442 ( .A(b[0]), .B(a[407]), .Z(n2034) );
  XOR U2443 ( .A(sreg[1430]), .B(n2034), .Z(n2036) );
  NANDN U2444 ( .A(n2029), .B(sreg[1429]), .Z(n2033) );
  OR U2445 ( .A(n2031), .B(n2030), .Z(n2032) );
  AND U2446 ( .A(n2033), .B(n2032), .Z(n2035) );
  XOR U2447 ( .A(n2036), .B(n2035), .Z(c[1430]) );
  NAND U2448 ( .A(b[0]), .B(a[408]), .Z(n2039) );
  XOR U2449 ( .A(sreg[1431]), .B(n2039), .Z(n2041) );
  NANDN U2450 ( .A(n2034), .B(sreg[1430]), .Z(n2038) );
  OR U2451 ( .A(n2036), .B(n2035), .Z(n2037) );
  AND U2452 ( .A(n2038), .B(n2037), .Z(n2040) );
  XOR U2453 ( .A(n2041), .B(n2040), .Z(c[1431]) );
  NAND U2454 ( .A(b[0]), .B(a[409]), .Z(n2044) );
  XOR U2455 ( .A(sreg[1432]), .B(n2044), .Z(n2046) );
  NANDN U2456 ( .A(n2039), .B(sreg[1431]), .Z(n2043) );
  OR U2457 ( .A(n2041), .B(n2040), .Z(n2042) );
  AND U2458 ( .A(n2043), .B(n2042), .Z(n2045) );
  XOR U2459 ( .A(n2046), .B(n2045), .Z(c[1432]) );
  NAND U2460 ( .A(b[0]), .B(a[410]), .Z(n2049) );
  XOR U2461 ( .A(sreg[1433]), .B(n2049), .Z(n2051) );
  NANDN U2462 ( .A(n2044), .B(sreg[1432]), .Z(n2048) );
  OR U2463 ( .A(n2046), .B(n2045), .Z(n2047) );
  AND U2464 ( .A(n2048), .B(n2047), .Z(n2050) );
  XOR U2465 ( .A(n2051), .B(n2050), .Z(c[1433]) );
  NAND U2466 ( .A(b[0]), .B(a[411]), .Z(n2054) );
  XOR U2467 ( .A(sreg[1434]), .B(n2054), .Z(n2056) );
  NANDN U2468 ( .A(n2049), .B(sreg[1433]), .Z(n2053) );
  OR U2469 ( .A(n2051), .B(n2050), .Z(n2052) );
  AND U2470 ( .A(n2053), .B(n2052), .Z(n2055) );
  XOR U2471 ( .A(n2056), .B(n2055), .Z(c[1434]) );
  NAND U2472 ( .A(b[0]), .B(a[412]), .Z(n2059) );
  XOR U2473 ( .A(sreg[1435]), .B(n2059), .Z(n2061) );
  NANDN U2474 ( .A(n2054), .B(sreg[1434]), .Z(n2058) );
  OR U2475 ( .A(n2056), .B(n2055), .Z(n2057) );
  AND U2476 ( .A(n2058), .B(n2057), .Z(n2060) );
  XOR U2477 ( .A(n2061), .B(n2060), .Z(c[1435]) );
  NAND U2478 ( .A(b[0]), .B(a[413]), .Z(n2064) );
  XOR U2479 ( .A(sreg[1436]), .B(n2064), .Z(n2066) );
  NANDN U2480 ( .A(n2059), .B(sreg[1435]), .Z(n2063) );
  OR U2481 ( .A(n2061), .B(n2060), .Z(n2062) );
  AND U2482 ( .A(n2063), .B(n2062), .Z(n2065) );
  XOR U2483 ( .A(n2066), .B(n2065), .Z(c[1436]) );
  NAND U2484 ( .A(b[0]), .B(a[414]), .Z(n2069) );
  XOR U2485 ( .A(sreg[1437]), .B(n2069), .Z(n2071) );
  NANDN U2486 ( .A(n2064), .B(sreg[1436]), .Z(n2068) );
  OR U2487 ( .A(n2066), .B(n2065), .Z(n2067) );
  AND U2488 ( .A(n2068), .B(n2067), .Z(n2070) );
  XOR U2489 ( .A(n2071), .B(n2070), .Z(c[1437]) );
  NAND U2490 ( .A(b[0]), .B(a[415]), .Z(n2074) );
  XOR U2491 ( .A(sreg[1438]), .B(n2074), .Z(n2076) );
  NANDN U2492 ( .A(n2069), .B(sreg[1437]), .Z(n2073) );
  OR U2493 ( .A(n2071), .B(n2070), .Z(n2072) );
  AND U2494 ( .A(n2073), .B(n2072), .Z(n2075) );
  XOR U2495 ( .A(n2076), .B(n2075), .Z(c[1438]) );
  NAND U2496 ( .A(b[0]), .B(a[416]), .Z(n2079) );
  XOR U2497 ( .A(sreg[1439]), .B(n2079), .Z(n2081) );
  NANDN U2498 ( .A(n2074), .B(sreg[1438]), .Z(n2078) );
  OR U2499 ( .A(n2076), .B(n2075), .Z(n2077) );
  AND U2500 ( .A(n2078), .B(n2077), .Z(n2080) );
  XOR U2501 ( .A(n2081), .B(n2080), .Z(c[1439]) );
  NAND U2502 ( .A(b[0]), .B(a[417]), .Z(n2084) );
  XOR U2503 ( .A(sreg[1440]), .B(n2084), .Z(n2086) );
  NANDN U2504 ( .A(n2079), .B(sreg[1439]), .Z(n2083) );
  OR U2505 ( .A(n2081), .B(n2080), .Z(n2082) );
  AND U2506 ( .A(n2083), .B(n2082), .Z(n2085) );
  XOR U2507 ( .A(n2086), .B(n2085), .Z(c[1440]) );
  NAND U2508 ( .A(b[0]), .B(a[418]), .Z(n2089) );
  XOR U2509 ( .A(sreg[1441]), .B(n2089), .Z(n2091) );
  NANDN U2510 ( .A(n2084), .B(sreg[1440]), .Z(n2088) );
  OR U2511 ( .A(n2086), .B(n2085), .Z(n2087) );
  AND U2512 ( .A(n2088), .B(n2087), .Z(n2090) );
  XOR U2513 ( .A(n2091), .B(n2090), .Z(c[1441]) );
  NAND U2514 ( .A(b[0]), .B(a[419]), .Z(n2094) );
  XOR U2515 ( .A(sreg[1442]), .B(n2094), .Z(n2096) );
  NANDN U2516 ( .A(n2089), .B(sreg[1441]), .Z(n2093) );
  OR U2517 ( .A(n2091), .B(n2090), .Z(n2092) );
  AND U2518 ( .A(n2093), .B(n2092), .Z(n2095) );
  XOR U2519 ( .A(n2096), .B(n2095), .Z(c[1442]) );
  NAND U2520 ( .A(b[0]), .B(a[420]), .Z(n2099) );
  XOR U2521 ( .A(sreg[1443]), .B(n2099), .Z(n2101) );
  NANDN U2522 ( .A(n2094), .B(sreg[1442]), .Z(n2098) );
  OR U2523 ( .A(n2096), .B(n2095), .Z(n2097) );
  AND U2524 ( .A(n2098), .B(n2097), .Z(n2100) );
  XOR U2525 ( .A(n2101), .B(n2100), .Z(c[1443]) );
  NAND U2526 ( .A(b[0]), .B(a[421]), .Z(n2104) );
  XOR U2527 ( .A(sreg[1444]), .B(n2104), .Z(n2106) );
  NANDN U2528 ( .A(n2099), .B(sreg[1443]), .Z(n2103) );
  OR U2529 ( .A(n2101), .B(n2100), .Z(n2102) );
  AND U2530 ( .A(n2103), .B(n2102), .Z(n2105) );
  XOR U2531 ( .A(n2106), .B(n2105), .Z(c[1444]) );
  NAND U2532 ( .A(b[0]), .B(a[422]), .Z(n2109) );
  XOR U2533 ( .A(sreg[1445]), .B(n2109), .Z(n2111) );
  NANDN U2534 ( .A(n2104), .B(sreg[1444]), .Z(n2108) );
  OR U2535 ( .A(n2106), .B(n2105), .Z(n2107) );
  AND U2536 ( .A(n2108), .B(n2107), .Z(n2110) );
  XOR U2537 ( .A(n2111), .B(n2110), .Z(c[1445]) );
  NAND U2538 ( .A(b[0]), .B(a[423]), .Z(n2114) );
  XOR U2539 ( .A(sreg[1446]), .B(n2114), .Z(n2116) );
  NANDN U2540 ( .A(n2109), .B(sreg[1445]), .Z(n2113) );
  OR U2541 ( .A(n2111), .B(n2110), .Z(n2112) );
  AND U2542 ( .A(n2113), .B(n2112), .Z(n2115) );
  XOR U2543 ( .A(n2116), .B(n2115), .Z(c[1446]) );
  NAND U2544 ( .A(b[0]), .B(a[424]), .Z(n2119) );
  XOR U2545 ( .A(sreg[1447]), .B(n2119), .Z(n2121) );
  NANDN U2546 ( .A(n2114), .B(sreg[1446]), .Z(n2118) );
  OR U2547 ( .A(n2116), .B(n2115), .Z(n2117) );
  AND U2548 ( .A(n2118), .B(n2117), .Z(n2120) );
  XOR U2549 ( .A(n2121), .B(n2120), .Z(c[1447]) );
  NAND U2550 ( .A(b[0]), .B(a[425]), .Z(n2124) );
  XOR U2551 ( .A(sreg[1448]), .B(n2124), .Z(n2126) );
  NANDN U2552 ( .A(n2119), .B(sreg[1447]), .Z(n2123) );
  OR U2553 ( .A(n2121), .B(n2120), .Z(n2122) );
  AND U2554 ( .A(n2123), .B(n2122), .Z(n2125) );
  XOR U2555 ( .A(n2126), .B(n2125), .Z(c[1448]) );
  NAND U2556 ( .A(b[0]), .B(a[426]), .Z(n2129) );
  XOR U2557 ( .A(sreg[1449]), .B(n2129), .Z(n2131) );
  NANDN U2558 ( .A(n2124), .B(sreg[1448]), .Z(n2128) );
  OR U2559 ( .A(n2126), .B(n2125), .Z(n2127) );
  AND U2560 ( .A(n2128), .B(n2127), .Z(n2130) );
  XOR U2561 ( .A(n2131), .B(n2130), .Z(c[1449]) );
  NAND U2562 ( .A(b[0]), .B(a[427]), .Z(n2134) );
  XOR U2563 ( .A(sreg[1450]), .B(n2134), .Z(n2136) );
  NANDN U2564 ( .A(n2129), .B(sreg[1449]), .Z(n2133) );
  OR U2565 ( .A(n2131), .B(n2130), .Z(n2132) );
  AND U2566 ( .A(n2133), .B(n2132), .Z(n2135) );
  XOR U2567 ( .A(n2136), .B(n2135), .Z(c[1450]) );
  NAND U2568 ( .A(b[0]), .B(a[428]), .Z(n2139) );
  XOR U2569 ( .A(sreg[1451]), .B(n2139), .Z(n2141) );
  NANDN U2570 ( .A(n2134), .B(sreg[1450]), .Z(n2138) );
  OR U2571 ( .A(n2136), .B(n2135), .Z(n2137) );
  AND U2572 ( .A(n2138), .B(n2137), .Z(n2140) );
  XOR U2573 ( .A(n2141), .B(n2140), .Z(c[1451]) );
  NAND U2574 ( .A(b[0]), .B(a[429]), .Z(n2144) );
  XOR U2575 ( .A(sreg[1452]), .B(n2144), .Z(n2146) );
  NANDN U2576 ( .A(n2139), .B(sreg[1451]), .Z(n2143) );
  OR U2577 ( .A(n2141), .B(n2140), .Z(n2142) );
  AND U2578 ( .A(n2143), .B(n2142), .Z(n2145) );
  XOR U2579 ( .A(n2146), .B(n2145), .Z(c[1452]) );
  NAND U2580 ( .A(b[0]), .B(a[430]), .Z(n2149) );
  XOR U2581 ( .A(sreg[1453]), .B(n2149), .Z(n2151) );
  NANDN U2582 ( .A(n2144), .B(sreg[1452]), .Z(n2148) );
  OR U2583 ( .A(n2146), .B(n2145), .Z(n2147) );
  AND U2584 ( .A(n2148), .B(n2147), .Z(n2150) );
  XOR U2585 ( .A(n2151), .B(n2150), .Z(c[1453]) );
  NAND U2586 ( .A(b[0]), .B(a[431]), .Z(n2154) );
  XOR U2587 ( .A(sreg[1454]), .B(n2154), .Z(n2156) );
  NANDN U2588 ( .A(n2149), .B(sreg[1453]), .Z(n2153) );
  OR U2589 ( .A(n2151), .B(n2150), .Z(n2152) );
  AND U2590 ( .A(n2153), .B(n2152), .Z(n2155) );
  XOR U2591 ( .A(n2156), .B(n2155), .Z(c[1454]) );
  NAND U2592 ( .A(b[0]), .B(a[432]), .Z(n2159) );
  XOR U2593 ( .A(sreg[1455]), .B(n2159), .Z(n2161) );
  NANDN U2594 ( .A(n2154), .B(sreg[1454]), .Z(n2158) );
  OR U2595 ( .A(n2156), .B(n2155), .Z(n2157) );
  AND U2596 ( .A(n2158), .B(n2157), .Z(n2160) );
  XOR U2597 ( .A(n2161), .B(n2160), .Z(c[1455]) );
  NAND U2598 ( .A(b[0]), .B(a[433]), .Z(n2164) );
  XOR U2599 ( .A(sreg[1456]), .B(n2164), .Z(n2166) );
  NANDN U2600 ( .A(n2159), .B(sreg[1455]), .Z(n2163) );
  OR U2601 ( .A(n2161), .B(n2160), .Z(n2162) );
  AND U2602 ( .A(n2163), .B(n2162), .Z(n2165) );
  XOR U2603 ( .A(n2166), .B(n2165), .Z(c[1456]) );
  NAND U2604 ( .A(b[0]), .B(a[434]), .Z(n2169) );
  XOR U2605 ( .A(sreg[1457]), .B(n2169), .Z(n2171) );
  NANDN U2606 ( .A(n2164), .B(sreg[1456]), .Z(n2168) );
  OR U2607 ( .A(n2166), .B(n2165), .Z(n2167) );
  AND U2608 ( .A(n2168), .B(n2167), .Z(n2170) );
  XOR U2609 ( .A(n2171), .B(n2170), .Z(c[1457]) );
  NAND U2610 ( .A(b[0]), .B(a[435]), .Z(n2174) );
  XOR U2611 ( .A(sreg[1458]), .B(n2174), .Z(n2176) );
  NANDN U2612 ( .A(n2169), .B(sreg[1457]), .Z(n2173) );
  OR U2613 ( .A(n2171), .B(n2170), .Z(n2172) );
  AND U2614 ( .A(n2173), .B(n2172), .Z(n2175) );
  XOR U2615 ( .A(n2176), .B(n2175), .Z(c[1458]) );
  NAND U2616 ( .A(b[0]), .B(a[436]), .Z(n2179) );
  XOR U2617 ( .A(sreg[1459]), .B(n2179), .Z(n2181) );
  NANDN U2618 ( .A(n2174), .B(sreg[1458]), .Z(n2178) );
  OR U2619 ( .A(n2176), .B(n2175), .Z(n2177) );
  AND U2620 ( .A(n2178), .B(n2177), .Z(n2180) );
  XOR U2621 ( .A(n2181), .B(n2180), .Z(c[1459]) );
  NAND U2622 ( .A(b[0]), .B(a[437]), .Z(n2184) );
  XOR U2623 ( .A(sreg[1460]), .B(n2184), .Z(n2186) );
  NANDN U2624 ( .A(n2179), .B(sreg[1459]), .Z(n2183) );
  OR U2625 ( .A(n2181), .B(n2180), .Z(n2182) );
  AND U2626 ( .A(n2183), .B(n2182), .Z(n2185) );
  XOR U2627 ( .A(n2186), .B(n2185), .Z(c[1460]) );
  NAND U2628 ( .A(b[0]), .B(a[438]), .Z(n2189) );
  XOR U2629 ( .A(sreg[1461]), .B(n2189), .Z(n2191) );
  NANDN U2630 ( .A(n2184), .B(sreg[1460]), .Z(n2188) );
  OR U2631 ( .A(n2186), .B(n2185), .Z(n2187) );
  AND U2632 ( .A(n2188), .B(n2187), .Z(n2190) );
  XOR U2633 ( .A(n2191), .B(n2190), .Z(c[1461]) );
  NAND U2634 ( .A(b[0]), .B(a[439]), .Z(n2194) );
  XOR U2635 ( .A(sreg[1462]), .B(n2194), .Z(n2196) );
  NANDN U2636 ( .A(n2189), .B(sreg[1461]), .Z(n2193) );
  OR U2637 ( .A(n2191), .B(n2190), .Z(n2192) );
  AND U2638 ( .A(n2193), .B(n2192), .Z(n2195) );
  XOR U2639 ( .A(n2196), .B(n2195), .Z(c[1462]) );
  NAND U2640 ( .A(b[0]), .B(a[440]), .Z(n2199) );
  XOR U2641 ( .A(sreg[1463]), .B(n2199), .Z(n2201) );
  NANDN U2642 ( .A(n2194), .B(sreg[1462]), .Z(n2198) );
  OR U2643 ( .A(n2196), .B(n2195), .Z(n2197) );
  AND U2644 ( .A(n2198), .B(n2197), .Z(n2200) );
  XOR U2645 ( .A(n2201), .B(n2200), .Z(c[1463]) );
  NAND U2646 ( .A(b[0]), .B(a[441]), .Z(n2204) );
  XOR U2647 ( .A(sreg[1464]), .B(n2204), .Z(n2206) );
  NANDN U2648 ( .A(n2199), .B(sreg[1463]), .Z(n2203) );
  OR U2649 ( .A(n2201), .B(n2200), .Z(n2202) );
  AND U2650 ( .A(n2203), .B(n2202), .Z(n2205) );
  XOR U2651 ( .A(n2206), .B(n2205), .Z(c[1464]) );
  NAND U2652 ( .A(b[0]), .B(a[442]), .Z(n2209) );
  XOR U2653 ( .A(sreg[1465]), .B(n2209), .Z(n2211) );
  NANDN U2654 ( .A(n2204), .B(sreg[1464]), .Z(n2208) );
  OR U2655 ( .A(n2206), .B(n2205), .Z(n2207) );
  AND U2656 ( .A(n2208), .B(n2207), .Z(n2210) );
  XOR U2657 ( .A(n2211), .B(n2210), .Z(c[1465]) );
  NAND U2658 ( .A(b[0]), .B(a[443]), .Z(n2214) );
  XOR U2659 ( .A(sreg[1466]), .B(n2214), .Z(n2216) );
  NANDN U2660 ( .A(n2209), .B(sreg[1465]), .Z(n2213) );
  OR U2661 ( .A(n2211), .B(n2210), .Z(n2212) );
  AND U2662 ( .A(n2213), .B(n2212), .Z(n2215) );
  XOR U2663 ( .A(n2216), .B(n2215), .Z(c[1466]) );
  NAND U2664 ( .A(b[0]), .B(a[444]), .Z(n2219) );
  XOR U2665 ( .A(sreg[1467]), .B(n2219), .Z(n2221) );
  NANDN U2666 ( .A(n2214), .B(sreg[1466]), .Z(n2218) );
  OR U2667 ( .A(n2216), .B(n2215), .Z(n2217) );
  AND U2668 ( .A(n2218), .B(n2217), .Z(n2220) );
  XOR U2669 ( .A(n2221), .B(n2220), .Z(c[1467]) );
  NAND U2670 ( .A(b[0]), .B(a[445]), .Z(n2224) );
  XOR U2671 ( .A(sreg[1468]), .B(n2224), .Z(n2226) );
  NANDN U2672 ( .A(n2219), .B(sreg[1467]), .Z(n2223) );
  OR U2673 ( .A(n2221), .B(n2220), .Z(n2222) );
  AND U2674 ( .A(n2223), .B(n2222), .Z(n2225) );
  XOR U2675 ( .A(n2226), .B(n2225), .Z(c[1468]) );
  NAND U2676 ( .A(b[0]), .B(a[446]), .Z(n2229) );
  XOR U2677 ( .A(sreg[1469]), .B(n2229), .Z(n2231) );
  NANDN U2678 ( .A(n2224), .B(sreg[1468]), .Z(n2228) );
  OR U2679 ( .A(n2226), .B(n2225), .Z(n2227) );
  AND U2680 ( .A(n2228), .B(n2227), .Z(n2230) );
  XOR U2681 ( .A(n2231), .B(n2230), .Z(c[1469]) );
  NAND U2682 ( .A(b[0]), .B(a[447]), .Z(n2234) );
  XOR U2683 ( .A(sreg[1470]), .B(n2234), .Z(n2236) );
  NANDN U2684 ( .A(n2229), .B(sreg[1469]), .Z(n2233) );
  OR U2685 ( .A(n2231), .B(n2230), .Z(n2232) );
  AND U2686 ( .A(n2233), .B(n2232), .Z(n2235) );
  XOR U2687 ( .A(n2236), .B(n2235), .Z(c[1470]) );
  NAND U2688 ( .A(b[0]), .B(a[448]), .Z(n2239) );
  XOR U2689 ( .A(sreg[1471]), .B(n2239), .Z(n2241) );
  NANDN U2690 ( .A(n2234), .B(sreg[1470]), .Z(n2238) );
  OR U2691 ( .A(n2236), .B(n2235), .Z(n2237) );
  AND U2692 ( .A(n2238), .B(n2237), .Z(n2240) );
  XOR U2693 ( .A(n2241), .B(n2240), .Z(c[1471]) );
  NAND U2694 ( .A(b[0]), .B(a[449]), .Z(n2244) );
  XOR U2695 ( .A(sreg[1472]), .B(n2244), .Z(n2246) );
  NANDN U2696 ( .A(n2239), .B(sreg[1471]), .Z(n2243) );
  OR U2697 ( .A(n2241), .B(n2240), .Z(n2242) );
  AND U2698 ( .A(n2243), .B(n2242), .Z(n2245) );
  XOR U2699 ( .A(n2246), .B(n2245), .Z(c[1472]) );
  NAND U2700 ( .A(b[0]), .B(a[450]), .Z(n2249) );
  XOR U2701 ( .A(sreg[1473]), .B(n2249), .Z(n2251) );
  NANDN U2702 ( .A(n2244), .B(sreg[1472]), .Z(n2248) );
  OR U2703 ( .A(n2246), .B(n2245), .Z(n2247) );
  AND U2704 ( .A(n2248), .B(n2247), .Z(n2250) );
  XOR U2705 ( .A(n2251), .B(n2250), .Z(c[1473]) );
  NAND U2706 ( .A(b[0]), .B(a[451]), .Z(n2254) );
  XOR U2707 ( .A(sreg[1474]), .B(n2254), .Z(n2256) );
  NANDN U2708 ( .A(n2249), .B(sreg[1473]), .Z(n2253) );
  OR U2709 ( .A(n2251), .B(n2250), .Z(n2252) );
  AND U2710 ( .A(n2253), .B(n2252), .Z(n2255) );
  XOR U2711 ( .A(n2256), .B(n2255), .Z(c[1474]) );
  NAND U2712 ( .A(b[0]), .B(a[452]), .Z(n2259) );
  XOR U2713 ( .A(sreg[1475]), .B(n2259), .Z(n2261) );
  NANDN U2714 ( .A(n2254), .B(sreg[1474]), .Z(n2258) );
  OR U2715 ( .A(n2256), .B(n2255), .Z(n2257) );
  AND U2716 ( .A(n2258), .B(n2257), .Z(n2260) );
  XOR U2717 ( .A(n2261), .B(n2260), .Z(c[1475]) );
  NAND U2718 ( .A(b[0]), .B(a[453]), .Z(n2264) );
  XOR U2719 ( .A(sreg[1476]), .B(n2264), .Z(n2266) );
  NANDN U2720 ( .A(n2259), .B(sreg[1475]), .Z(n2263) );
  OR U2721 ( .A(n2261), .B(n2260), .Z(n2262) );
  AND U2722 ( .A(n2263), .B(n2262), .Z(n2265) );
  XOR U2723 ( .A(n2266), .B(n2265), .Z(c[1476]) );
  NAND U2724 ( .A(b[0]), .B(a[454]), .Z(n2269) );
  XOR U2725 ( .A(sreg[1477]), .B(n2269), .Z(n2271) );
  NANDN U2726 ( .A(n2264), .B(sreg[1476]), .Z(n2268) );
  OR U2727 ( .A(n2266), .B(n2265), .Z(n2267) );
  AND U2728 ( .A(n2268), .B(n2267), .Z(n2270) );
  XOR U2729 ( .A(n2271), .B(n2270), .Z(c[1477]) );
  NAND U2730 ( .A(b[0]), .B(a[455]), .Z(n2274) );
  XOR U2731 ( .A(sreg[1478]), .B(n2274), .Z(n2276) );
  NANDN U2732 ( .A(n2269), .B(sreg[1477]), .Z(n2273) );
  OR U2733 ( .A(n2271), .B(n2270), .Z(n2272) );
  AND U2734 ( .A(n2273), .B(n2272), .Z(n2275) );
  XOR U2735 ( .A(n2276), .B(n2275), .Z(c[1478]) );
  NAND U2736 ( .A(b[0]), .B(a[456]), .Z(n2279) );
  XOR U2737 ( .A(sreg[1479]), .B(n2279), .Z(n2281) );
  NANDN U2738 ( .A(n2274), .B(sreg[1478]), .Z(n2278) );
  OR U2739 ( .A(n2276), .B(n2275), .Z(n2277) );
  AND U2740 ( .A(n2278), .B(n2277), .Z(n2280) );
  XOR U2741 ( .A(n2281), .B(n2280), .Z(c[1479]) );
  NAND U2742 ( .A(b[0]), .B(a[457]), .Z(n2284) );
  XOR U2743 ( .A(sreg[1480]), .B(n2284), .Z(n2286) );
  NANDN U2744 ( .A(n2279), .B(sreg[1479]), .Z(n2283) );
  OR U2745 ( .A(n2281), .B(n2280), .Z(n2282) );
  AND U2746 ( .A(n2283), .B(n2282), .Z(n2285) );
  XOR U2747 ( .A(n2286), .B(n2285), .Z(c[1480]) );
  NAND U2748 ( .A(b[0]), .B(a[458]), .Z(n2289) );
  XOR U2749 ( .A(sreg[1481]), .B(n2289), .Z(n2291) );
  NANDN U2750 ( .A(n2284), .B(sreg[1480]), .Z(n2288) );
  OR U2751 ( .A(n2286), .B(n2285), .Z(n2287) );
  AND U2752 ( .A(n2288), .B(n2287), .Z(n2290) );
  XOR U2753 ( .A(n2291), .B(n2290), .Z(c[1481]) );
  NAND U2754 ( .A(b[0]), .B(a[459]), .Z(n2294) );
  XOR U2755 ( .A(sreg[1482]), .B(n2294), .Z(n2296) );
  NANDN U2756 ( .A(n2289), .B(sreg[1481]), .Z(n2293) );
  OR U2757 ( .A(n2291), .B(n2290), .Z(n2292) );
  AND U2758 ( .A(n2293), .B(n2292), .Z(n2295) );
  XOR U2759 ( .A(n2296), .B(n2295), .Z(c[1482]) );
  NAND U2760 ( .A(b[0]), .B(a[460]), .Z(n2299) );
  XOR U2761 ( .A(sreg[1483]), .B(n2299), .Z(n2301) );
  NANDN U2762 ( .A(n2294), .B(sreg[1482]), .Z(n2298) );
  OR U2763 ( .A(n2296), .B(n2295), .Z(n2297) );
  AND U2764 ( .A(n2298), .B(n2297), .Z(n2300) );
  XOR U2765 ( .A(n2301), .B(n2300), .Z(c[1483]) );
  NAND U2766 ( .A(b[0]), .B(a[461]), .Z(n2304) );
  XOR U2767 ( .A(sreg[1484]), .B(n2304), .Z(n2306) );
  NANDN U2768 ( .A(n2299), .B(sreg[1483]), .Z(n2303) );
  OR U2769 ( .A(n2301), .B(n2300), .Z(n2302) );
  AND U2770 ( .A(n2303), .B(n2302), .Z(n2305) );
  XOR U2771 ( .A(n2306), .B(n2305), .Z(c[1484]) );
  NAND U2772 ( .A(b[0]), .B(a[462]), .Z(n2309) );
  XOR U2773 ( .A(sreg[1485]), .B(n2309), .Z(n2311) );
  NANDN U2774 ( .A(n2304), .B(sreg[1484]), .Z(n2308) );
  OR U2775 ( .A(n2306), .B(n2305), .Z(n2307) );
  AND U2776 ( .A(n2308), .B(n2307), .Z(n2310) );
  XOR U2777 ( .A(n2311), .B(n2310), .Z(c[1485]) );
  NAND U2778 ( .A(b[0]), .B(a[463]), .Z(n2314) );
  XOR U2779 ( .A(sreg[1486]), .B(n2314), .Z(n2316) );
  NANDN U2780 ( .A(n2309), .B(sreg[1485]), .Z(n2313) );
  OR U2781 ( .A(n2311), .B(n2310), .Z(n2312) );
  AND U2782 ( .A(n2313), .B(n2312), .Z(n2315) );
  XOR U2783 ( .A(n2316), .B(n2315), .Z(c[1486]) );
  NAND U2784 ( .A(b[0]), .B(a[464]), .Z(n2319) );
  XOR U2785 ( .A(sreg[1487]), .B(n2319), .Z(n2321) );
  NANDN U2786 ( .A(n2314), .B(sreg[1486]), .Z(n2318) );
  OR U2787 ( .A(n2316), .B(n2315), .Z(n2317) );
  AND U2788 ( .A(n2318), .B(n2317), .Z(n2320) );
  XOR U2789 ( .A(n2321), .B(n2320), .Z(c[1487]) );
  NAND U2790 ( .A(b[0]), .B(a[465]), .Z(n2324) );
  XOR U2791 ( .A(sreg[1488]), .B(n2324), .Z(n2326) );
  NANDN U2792 ( .A(n2319), .B(sreg[1487]), .Z(n2323) );
  OR U2793 ( .A(n2321), .B(n2320), .Z(n2322) );
  AND U2794 ( .A(n2323), .B(n2322), .Z(n2325) );
  XOR U2795 ( .A(n2326), .B(n2325), .Z(c[1488]) );
  NAND U2796 ( .A(b[0]), .B(a[466]), .Z(n2329) );
  XOR U2797 ( .A(sreg[1489]), .B(n2329), .Z(n2331) );
  NANDN U2798 ( .A(n2324), .B(sreg[1488]), .Z(n2328) );
  OR U2799 ( .A(n2326), .B(n2325), .Z(n2327) );
  AND U2800 ( .A(n2328), .B(n2327), .Z(n2330) );
  XOR U2801 ( .A(n2331), .B(n2330), .Z(c[1489]) );
  NAND U2802 ( .A(b[0]), .B(a[467]), .Z(n2334) );
  XOR U2803 ( .A(sreg[1490]), .B(n2334), .Z(n2336) );
  NANDN U2804 ( .A(n2329), .B(sreg[1489]), .Z(n2333) );
  OR U2805 ( .A(n2331), .B(n2330), .Z(n2332) );
  AND U2806 ( .A(n2333), .B(n2332), .Z(n2335) );
  XOR U2807 ( .A(n2336), .B(n2335), .Z(c[1490]) );
  NAND U2808 ( .A(b[0]), .B(a[468]), .Z(n2339) );
  XOR U2809 ( .A(sreg[1491]), .B(n2339), .Z(n2341) );
  NANDN U2810 ( .A(n2334), .B(sreg[1490]), .Z(n2338) );
  OR U2811 ( .A(n2336), .B(n2335), .Z(n2337) );
  AND U2812 ( .A(n2338), .B(n2337), .Z(n2340) );
  XOR U2813 ( .A(n2341), .B(n2340), .Z(c[1491]) );
  NAND U2814 ( .A(b[0]), .B(a[469]), .Z(n2344) );
  XOR U2815 ( .A(sreg[1492]), .B(n2344), .Z(n2346) );
  NANDN U2816 ( .A(n2339), .B(sreg[1491]), .Z(n2343) );
  OR U2817 ( .A(n2341), .B(n2340), .Z(n2342) );
  AND U2818 ( .A(n2343), .B(n2342), .Z(n2345) );
  XOR U2819 ( .A(n2346), .B(n2345), .Z(c[1492]) );
  NAND U2820 ( .A(b[0]), .B(a[470]), .Z(n2349) );
  XOR U2821 ( .A(sreg[1493]), .B(n2349), .Z(n2351) );
  NANDN U2822 ( .A(n2344), .B(sreg[1492]), .Z(n2348) );
  OR U2823 ( .A(n2346), .B(n2345), .Z(n2347) );
  AND U2824 ( .A(n2348), .B(n2347), .Z(n2350) );
  XOR U2825 ( .A(n2351), .B(n2350), .Z(c[1493]) );
  NAND U2826 ( .A(b[0]), .B(a[471]), .Z(n2354) );
  XOR U2827 ( .A(sreg[1494]), .B(n2354), .Z(n2356) );
  NANDN U2828 ( .A(n2349), .B(sreg[1493]), .Z(n2353) );
  OR U2829 ( .A(n2351), .B(n2350), .Z(n2352) );
  AND U2830 ( .A(n2353), .B(n2352), .Z(n2355) );
  XOR U2831 ( .A(n2356), .B(n2355), .Z(c[1494]) );
  NAND U2832 ( .A(b[0]), .B(a[472]), .Z(n2359) );
  XOR U2833 ( .A(sreg[1495]), .B(n2359), .Z(n2361) );
  NANDN U2834 ( .A(n2354), .B(sreg[1494]), .Z(n2358) );
  OR U2835 ( .A(n2356), .B(n2355), .Z(n2357) );
  AND U2836 ( .A(n2358), .B(n2357), .Z(n2360) );
  XOR U2837 ( .A(n2361), .B(n2360), .Z(c[1495]) );
  NAND U2838 ( .A(b[0]), .B(a[473]), .Z(n2364) );
  XOR U2839 ( .A(sreg[1496]), .B(n2364), .Z(n2366) );
  NANDN U2840 ( .A(n2359), .B(sreg[1495]), .Z(n2363) );
  OR U2841 ( .A(n2361), .B(n2360), .Z(n2362) );
  AND U2842 ( .A(n2363), .B(n2362), .Z(n2365) );
  XOR U2843 ( .A(n2366), .B(n2365), .Z(c[1496]) );
  NAND U2844 ( .A(b[0]), .B(a[474]), .Z(n2369) );
  XOR U2845 ( .A(sreg[1497]), .B(n2369), .Z(n2371) );
  NANDN U2846 ( .A(n2364), .B(sreg[1496]), .Z(n2368) );
  OR U2847 ( .A(n2366), .B(n2365), .Z(n2367) );
  AND U2848 ( .A(n2368), .B(n2367), .Z(n2370) );
  XOR U2849 ( .A(n2371), .B(n2370), .Z(c[1497]) );
  NAND U2850 ( .A(b[0]), .B(a[475]), .Z(n2374) );
  XOR U2851 ( .A(sreg[1498]), .B(n2374), .Z(n2376) );
  NANDN U2852 ( .A(n2369), .B(sreg[1497]), .Z(n2373) );
  OR U2853 ( .A(n2371), .B(n2370), .Z(n2372) );
  AND U2854 ( .A(n2373), .B(n2372), .Z(n2375) );
  XOR U2855 ( .A(n2376), .B(n2375), .Z(c[1498]) );
  NAND U2856 ( .A(b[0]), .B(a[476]), .Z(n2379) );
  XOR U2857 ( .A(sreg[1499]), .B(n2379), .Z(n2381) );
  NANDN U2858 ( .A(n2374), .B(sreg[1498]), .Z(n2378) );
  OR U2859 ( .A(n2376), .B(n2375), .Z(n2377) );
  AND U2860 ( .A(n2378), .B(n2377), .Z(n2380) );
  XOR U2861 ( .A(n2381), .B(n2380), .Z(c[1499]) );
  NAND U2862 ( .A(b[0]), .B(a[477]), .Z(n2384) );
  XOR U2863 ( .A(sreg[1500]), .B(n2384), .Z(n2386) );
  NANDN U2864 ( .A(n2379), .B(sreg[1499]), .Z(n2383) );
  OR U2865 ( .A(n2381), .B(n2380), .Z(n2382) );
  AND U2866 ( .A(n2383), .B(n2382), .Z(n2385) );
  XOR U2867 ( .A(n2386), .B(n2385), .Z(c[1500]) );
  NAND U2868 ( .A(b[0]), .B(a[478]), .Z(n2389) );
  XOR U2869 ( .A(sreg[1501]), .B(n2389), .Z(n2391) );
  NANDN U2870 ( .A(n2384), .B(sreg[1500]), .Z(n2388) );
  OR U2871 ( .A(n2386), .B(n2385), .Z(n2387) );
  AND U2872 ( .A(n2388), .B(n2387), .Z(n2390) );
  XOR U2873 ( .A(n2391), .B(n2390), .Z(c[1501]) );
  NAND U2874 ( .A(b[0]), .B(a[479]), .Z(n2394) );
  XOR U2875 ( .A(sreg[1502]), .B(n2394), .Z(n2396) );
  NANDN U2876 ( .A(n2389), .B(sreg[1501]), .Z(n2393) );
  OR U2877 ( .A(n2391), .B(n2390), .Z(n2392) );
  AND U2878 ( .A(n2393), .B(n2392), .Z(n2395) );
  XOR U2879 ( .A(n2396), .B(n2395), .Z(c[1502]) );
  NAND U2880 ( .A(b[0]), .B(a[480]), .Z(n2399) );
  XOR U2881 ( .A(sreg[1503]), .B(n2399), .Z(n2401) );
  NANDN U2882 ( .A(n2394), .B(sreg[1502]), .Z(n2398) );
  OR U2883 ( .A(n2396), .B(n2395), .Z(n2397) );
  AND U2884 ( .A(n2398), .B(n2397), .Z(n2400) );
  XOR U2885 ( .A(n2401), .B(n2400), .Z(c[1503]) );
  NAND U2886 ( .A(b[0]), .B(a[481]), .Z(n2404) );
  XOR U2887 ( .A(sreg[1504]), .B(n2404), .Z(n2406) );
  NANDN U2888 ( .A(n2399), .B(sreg[1503]), .Z(n2403) );
  OR U2889 ( .A(n2401), .B(n2400), .Z(n2402) );
  AND U2890 ( .A(n2403), .B(n2402), .Z(n2405) );
  XOR U2891 ( .A(n2406), .B(n2405), .Z(c[1504]) );
  NAND U2892 ( .A(b[0]), .B(a[482]), .Z(n2409) );
  XOR U2893 ( .A(sreg[1505]), .B(n2409), .Z(n2411) );
  NANDN U2894 ( .A(n2404), .B(sreg[1504]), .Z(n2408) );
  OR U2895 ( .A(n2406), .B(n2405), .Z(n2407) );
  AND U2896 ( .A(n2408), .B(n2407), .Z(n2410) );
  XOR U2897 ( .A(n2411), .B(n2410), .Z(c[1505]) );
  NAND U2898 ( .A(b[0]), .B(a[483]), .Z(n2414) );
  XOR U2899 ( .A(sreg[1506]), .B(n2414), .Z(n2416) );
  NANDN U2900 ( .A(n2409), .B(sreg[1505]), .Z(n2413) );
  OR U2901 ( .A(n2411), .B(n2410), .Z(n2412) );
  AND U2902 ( .A(n2413), .B(n2412), .Z(n2415) );
  XOR U2903 ( .A(n2416), .B(n2415), .Z(c[1506]) );
  NAND U2904 ( .A(b[0]), .B(a[484]), .Z(n2419) );
  XOR U2905 ( .A(sreg[1507]), .B(n2419), .Z(n2421) );
  NANDN U2906 ( .A(n2414), .B(sreg[1506]), .Z(n2418) );
  OR U2907 ( .A(n2416), .B(n2415), .Z(n2417) );
  AND U2908 ( .A(n2418), .B(n2417), .Z(n2420) );
  XOR U2909 ( .A(n2421), .B(n2420), .Z(c[1507]) );
  NAND U2910 ( .A(b[0]), .B(a[485]), .Z(n2424) );
  XOR U2911 ( .A(sreg[1508]), .B(n2424), .Z(n2426) );
  NANDN U2912 ( .A(n2419), .B(sreg[1507]), .Z(n2423) );
  OR U2913 ( .A(n2421), .B(n2420), .Z(n2422) );
  AND U2914 ( .A(n2423), .B(n2422), .Z(n2425) );
  XOR U2915 ( .A(n2426), .B(n2425), .Z(c[1508]) );
  NAND U2916 ( .A(b[0]), .B(a[486]), .Z(n2429) );
  XOR U2917 ( .A(sreg[1509]), .B(n2429), .Z(n2431) );
  NANDN U2918 ( .A(n2424), .B(sreg[1508]), .Z(n2428) );
  OR U2919 ( .A(n2426), .B(n2425), .Z(n2427) );
  AND U2920 ( .A(n2428), .B(n2427), .Z(n2430) );
  XOR U2921 ( .A(n2431), .B(n2430), .Z(c[1509]) );
  NAND U2922 ( .A(b[0]), .B(a[487]), .Z(n2434) );
  XOR U2923 ( .A(sreg[1510]), .B(n2434), .Z(n2436) );
  NANDN U2924 ( .A(n2429), .B(sreg[1509]), .Z(n2433) );
  OR U2925 ( .A(n2431), .B(n2430), .Z(n2432) );
  AND U2926 ( .A(n2433), .B(n2432), .Z(n2435) );
  XOR U2927 ( .A(n2436), .B(n2435), .Z(c[1510]) );
  NAND U2928 ( .A(b[0]), .B(a[488]), .Z(n2439) );
  XOR U2929 ( .A(sreg[1511]), .B(n2439), .Z(n2441) );
  NANDN U2930 ( .A(n2434), .B(sreg[1510]), .Z(n2438) );
  OR U2931 ( .A(n2436), .B(n2435), .Z(n2437) );
  AND U2932 ( .A(n2438), .B(n2437), .Z(n2440) );
  XOR U2933 ( .A(n2441), .B(n2440), .Z(c[1511]) );
  NAND U2934 ( .A(b[0]), .B(a[489]), .Z(n2444) );
  XOR U2935 ( .A(sreg[1512]), .B(n2444), .Z(n2446) );
  NANDN U2936 ( .A(n2439), .B(sreg[1511]), .Z(n2443) );
  OR U2937 ( .A(n2441), .B(n2440), .Z(n2442) );
  AND U2938 ( .A(n2443), .B(n2442), .Z(n2445) );
  XOR U2939 ( .A(n2446), .B(n2445), .Z(c[1512]) );
  NAND U2940 ( .A(b[0]), .B(a[490]), .Z(n2449) );
  XOR U2941 ( .A(sreg[1513]), .B(n2449), .Z(n2451) );
  NANDN U2942 ( .A(n2444), .B(sreg[1512]), .Z(n2448) );
  OR U2943 ( .A(n2446), .B(n2445), .Z(n2447) );
  AND U2944 ( .A(n2448), .B(n2447), .Z(n2450) );
  XOR U2945 ( .A(n2451), .B(n2450), .Z(c[1513]) );
  NAND U2946 ( .A(b[0]), .B(a[491]), .Z(n2454) );
  XOR U2947 ( .A(sreg[1514]), .B(n2454), .Z(n2456) );
  NANDN U2948 ( .A(n2449), .B(sreg[1513]), .Z(n2453) );
  OR U2949 ( .A(n2451), .B(n2450), .Z(n2452) );
  AND U2950 ( .A(n2453), .B(n2452), .Z(n2455) );
  XOR U2951 ( .A(n2456), .B(n2455), .Z(c[1514]) );
  NAND U2952 ( .A(b[0]), .B(a[492]), .Z(n2459) );
  XOR U2953 ( .A(sreg[1515]), .B(n2459), .Z(n2461) );
  NANDN U2954 ( .A(n2454), .B(sreg[1514]), .Z(n2458) );
  OR U2955 ( .A(n2456), .B(n2455), .Z(n2457) );
  AND U2956 ( .A(n2458), .B(n2457), .Z(n2460) );
  XOR U2957 ( .A(n2461), .B(n2460), .Z(c[1515]) );
  NAND U2958 ( .A(b[0]), .B(a[493]), .Z(n2464) );
  XOR U2959 ( .A(sreg[1516]), .B(n2464), .Z(n2466) );
  NANDN U2960 ( .A(n2459), .B(sreg[1515]), .Z(n2463) );
  OR U2961 ( .A(n2461), .B(n2460), .Z(n2462) );
  AND U2962 ( .A(n2463), .B(n2462), .Z(n2465) );
  XOR U2963 ( .A(n2466), .B(n2465), .Z(c[1516]) );
  NAND U2964 ( .A(b[0]), .B(a[494]), .Z(n2469) );
  XOR U2965 ( .A(sreg[1517]), .B(n2469), .Z(n2471) );
  NANDN U2966 ( .A(n2464), .B(sreg[1516]), .Z(n2468) );
  OR U2967 ( .A(n2466), .B(n2465), .Z(n2467) );
  AND U2968 ( .A(n2468), .B(n2467), .Z(n2470) );
  XOR U2969 ( .A(n2471), .B(n2470), .Z(c[1517]) );
  NAND U2970 ( .A(b[0]), .B(a[495]), .Z(n2474) );
  XOR U2971 ( .A(sreg[1518]), .B(n2474), .Z(n2476) );
  NANDN U2972 ( .A(n2469), .B(sreg[1517]), .Z(n2473) );
  OR U2973 ( .A(n2471), .B(n2470), .Z(n2472) );
  AND U2974 ( .A(n2473), .B(n2472), .Z(n2475) );
  XOR U2975 ( .A(n2476), .B(n2475), .Z(c[1518]) );
  NAND U2976 ( .A(b[0]), .B(a[496]), .Z(n2479) );
  XOR U2977 ( .A(sreg[1519]), .B(n2479), .Z(n2481) );
  NANDN U2978 ( .A(n2474), .B(sreg[1518]), .Z(n2478) );
  OR U2979 ( .A(n2476), .B(n2475), .Z(n2477) );
  AND U2980 ( .A(n2478), .B(n2477), .Z(n2480) );
  XOR U2981 ( .A(n2481), .B(n2480), .Z(c[1519]) );
  NAND U2982 ( .A(b[0]), .B(a[497]), .Z(n2484) );
  XOR U2983 ( .A(sreg[1520]), .B(n2484), .Z(n2486) );
  NANDN U2984 ( .A(n2479), .B(sreg[1519]), .Z(n2483) );
  OR U2985 ( .A(n2481), .B(n2480), .Z(n2482) );
  AND U2986 ( .A(n2483), .B(n2482), .Z(n2485) );
  XOR U2987 ( .A(n2486), .B(n2485), .Z(c[1520]) );
  NAND U2988 ( .A(b[0]), .B(a[498]), .Z(n2489) );
  XOR U2989 ( .A(sreg[1521]), .B(n2489), .Z(n2491) );
  NANDN U2990 ( .A(n2484), .B(sreg[1520]), .Z(n2488) );
  OR U2991 ( .A(n2486), .B(n2485), .Z(n2487) );
  AND U2992 ( .A(n2488), .B(n2487), .Z(n2490) );
  XOR U2993 ( .A(n2491), .B(n2490), .Z(c[1521]) );
  NAND U2994 ( .A(b[0]), .B(a[499]), .Z(n2494) );
  XOR U2995 ( .A(sreg[1522]), .B(n2494), .Z(n2496) );
  NANDN U2996 ( .A(n2489), .B(sreg[1521]), .Z(n2493) );
  OR U2997 ( .A(n2491), .B(n2490), .Z(n2492) );
  AND U2998 ( .A(n2493), .B(n2492), .Z(n2495) );
  XOR U2999 ( .A(n2496), .B(n2495), .Z(c[1522]) );
  NAND U3000 ( .A(b[0]), .B(a[500]), .Z(n2499) );
  XOR U3001 ( .A(sreg[1523]), .B(n2499), .Z(n2501) );
  NANDN U3002 ( .A(n2494), .B(sreg[1522]), .Z(n2498) );
  OR U3003 ( .A(n2496), .B(n2495), .Z(n2497) );
  AND U3004 ( .A(n2498), .B(n2497), .Z(n2500) );
  XOR U3005 ( .A(n2501), .B(n2500), .Z(c[1523]) );
  NAND U3006 ( .A(b[0]), .B(a[501]), .Z(n2504) );
  XOR U3007 ( .A(sreg[1524]), .B(n2504), .Z(n2506) );
  NANDN U3008 ( .A(n2499), .B(sreg[1523]), .Z(n2503) );
  OR U3009 ( .A(n2501), .B(n2500), .Z(n2502) );
  AND U3010 ( .A(n2503), .B(n2502), .Z(n2505) );
  XOR U3011 ( .A(n2506), .B(n2505), .Z(c[1524]) );
  NAND U3012 ( .A(b[0]), .B(a[502]), .Z(n2509) );
  XOR U3013 ( .A(sreg[1525]), .B(n2509), .Z(n2511) );
  NANDN U3014 ( .A(n2504), .B(sreg[1524]), .Z(n2508) );
  OR U3015 ( .A(n2506), .B(n2505), .Z(n2507) );
  AND U3016 ( .A(n2508), .B(n2507), .Z(n2510) );
  XOR U3017 ( .A(n2511), .B(n2510), .Z(c[1525]) );
  NAND U3018 ( .A(b[0]), .B(a[503]), .Z(n2514) );
  XOR U3019 ( .A(sreg[1526]), .B(n2514), .Z(n2516) );
  NANDN U3020 ( .A(n2509), .B(sreg[1525]), .Z(n2513) );
  OR U3021 ( .A(n2511), .B(n2510), .Z(n2512) );
  AND U3022 ( .A(n2513), .B(n2512), .Z(n2515) );
  XOR U3023 ( .A(n2516), .B(n2515), .Z(c[1526]) );
  NAND U3024 ( .A(b[0]), .B(a[504]), .Z(n2519) );
  XOR U3025 ( .A(sreg[1527]), .B(n2519), .Z(n2521) );
  NANDN U3026 ( .A(n2514), .B(sreg[1526]), .Z(n2518) );
  OR U3027 ( .A(n2516), .B(n2515), .Z(n2517) );
  AND U3028 ( .A(n2518), .B(n2517), .Z(n2520) );
  XOR U3029 ( .A(n2521), .B(n2520), .Z(c[1527]) );
  NAND U3030 ( .A(b[0]), .B(a[505]), .Z(n2524) );
  XOR U3031 ( .A(sreg[1528]), .B(n2524), .Z(n2526) );
  NANDN U3032 ( .A(n2519), .B(sreg[1527]), .Z(n2523) );
  OR U3033 ( .A(n2521), .B(n2520), .Z(n2522) );
  AND U3034 ( .A(n2523), .B(n2522), .Z(n2525) );
  XOR U3035 ( .A(n2526), .B(n2525), .Z(c[1528]) );
  NAND U3036 ( .A(b[0]), .B(a[506]), .Z(n2529) );
  XOR U3037 ( .A(sreg[1529]), .B(n2529), .Z(n2531) );
  NANDN U3038 ( .A(n2524), .B(sreg[1528]), .Z(n2528) );
  OR U3039 ( .A(n2526), .B(n2525), .Z(n2527) );
  AND U3040 ( .A(n2528), .B(n2527), .Z(n2530) );
  XOR U3041 ( .A(n2531), .B(n2530), .Z(c[1529]) );
  NAND U3042 ( .A(b[0]), .B(a[507]), .Z(n2534) );
  XOR U3043 ( .A(sreg[1530]), .B(n2534), .Z(n2536) );
  NANDN U3044 ( .A(n2529), .B(sreg[1529]), .Z(n2533) );
  OR U3045 ( .A(n2531), .B(n2530), .Z(n2532) );
  AND U3046 ( .A(n2533), .B(n2532), .Z(n2535) );
  XOR U3047 ( .A(n2536), .B(n2535), .Z(c[1530]) );
  NAND U3048 ( .A(b[0]), .B(a[508]), .Z(n2539) );
  XOR U3049 ( .A(sreg[1531]), .B(n2539), .Z(n2541) );
  NANDN U3050 ( .A(n2534), .B(sreg[1530]), .Z(n2538) );
  OR U3051 ( .A(n2536), .B(n2535), .Z(n2537) );
  AND U3052 ( .A(n2538), .B(n2537), .Z(n2540) );
  XOR U3053 ( .A(n2541), .B(n2540), .Z(c[1531]) );
  NAND U3054 ( .A(b[0]), .B(a[509]), .Z(n2544) );
  XOR U3055 ( .A(sreg[1532]), .B(n2544), .Z(n2546) );
  NANDN U3056 ( .A(n2539), .B(sreg[1531]), .Z(n2543) );
  OR U3057 ( .A(n2541), .B(n2540), .Z(n2542) );
  AND U3058 ( .A(n2543), .B(n2542), .Z(n2545) );
  XOR U3059 ( .A(n2546), .B(n2545), .Z(c[1532]) );
  NAND U3060 ( .A(b[0]), .B(a[510]), .Z(n2549) );
  XOR U3061 ( .A(sreg[1533]), .B(n2549), .Z(n2551) );
  NANDN U3062 ( .A(n2544), .B(sreg[1532]), .Z(n2548) );
  OR U3063 ( .A(n2546), .B(n2545), .Z(n2547) );
  AND U3064 ( .A(n2548), .B(n2547), .Z(n2550) );
  XOR U3065 ( .A(n2551), .B(n2550), .Z(c[1533]) );
  NAND U3066 ( .A(b[0]), .B(a[511]), .Z(n2554) );
  XOR U3067 ( .A(sreg[1534]), .B(n2554), .Z(n2556) );
  NANDN U3068 ( .A(n2549), .B(sreg[1533]), .Z(n2553) );
  OR U3069 ( .A(n2551), .B(n2550), .Z(n2552) );
  AND U3070 ( .A(n2553), .B(n2552), .Z(n2555) );
  XOR U3071 ( .A(n2556), .B(n2555), .Z(c[1534]) );
  NAND U3072 ( .A(b[0]), .B(a[512]), .Z(n2559) );
  XOR U3073 ( .A(sreg[1535]), .B(n2559), .Z(n2561) );
  NANDN U3074 ( .A(n2554), .B(sreg[1534]), .Z(n2558) );
  OR U3075 ( .A(n2556), .B(n2555), .Z(n2557) );
  AND U3076 ( .A(n2558), .B(n2557), .Z(n2560) );
  XOR U3077 ( .A(n2561), .B(n2560), .Z(c[1535]) );
  NAND U3078 ( .A(b[0]), .B(a[513]), .Z(n2564) );
  XOR U3079 ( .A(sreg[1536]), .B(n2564), .Z(n2566) );
  NANDN U3080 ( .A(n2559), .B(sreg[1535]), .Z(n2563) );
  OR U3081 ( .A(n2561), .B(n2560), .Z(n2562) );
  AND U3082 ( .A(n2563), .B(n2562), .Z(n2565) );
  XOR U3083 ( .A(n2566), .B(n2565), .Z(c[1536]) );
  NAND U3084 ( .A(b[0]), .B(a[514]), .Z(n2569) );
  XOR U3085 ( .A(sreg[1537]), .B(n2569), .Z(n2571) );
  NANDN U3086 ( .A(n2564), .B(sreg[1536]), .Z(n2568) );
  OR U3087 ( .A(n2566), .B(n2565), .Z(n2567) );
  AND U3088 ( .A(n2568), .B(n2567), .Z(n2570) );
  XOR U3089 ( .A(n2571), .B(n2570), .Z(c[1537]) );
  NAND U3090 ( .A(b[0]), .B(a[515]), .Z(n2574) );
  XOR U3091 ( .A(sreg[1538]), .B(n2574), .Z(n2576) );
  NANDN U3092 ( .A(n2569), .B(sreg[1537]), .Z(n2573) );
  OR U3093 ( .A(n2571), .B(n2570), .Z(n2572) );
  AND U3094 ( .A(n2573), .B(n2572), .Z(n2575) );
  XOR U3095 ( .A(n2576), .B(n2575), .Z(c[1538]) );
  NAND U3096 ( .A(b[0]), .B(a[516]), .Z(n2579) );
  XOR U3097 ( .A(sreg[1539]), .B(n2579), .Z(n2581) );
  NANDN U3098 ( .A(n2574), .B(sreg[1538]), .Z(n2578) );
  OR U3099 ( .A(n2576), .B(n2575), .Z(n2577) );
  AND U3100 ( .A(n2578), .B(n2577), .Z(n2580) );
  XOR U3101 ( .A(n2581), .B(n2580), .Z(c[1539]) );
  NAND U3102 ( .A(b[0]), .B(a[517]), .Z(n2584) );
  XOR U3103 ( .A(sreg[1540]), .B(n2584), .Z(n2586) );
  NANDN U3104 ( .A(n2579), .B(sreg[1539]), .Z(n2583) );
  OR U3105 ( .A(n2581), .B(n2580), .Z(n2582) );
  AND U3106 ( .A(n2583), .B(n2582), .Z(n2585) );
  XOR U3107 ( .A(n2586), .B(n2585), .Z(c[1540]) );
  NAND U3108 ( .A(b[0]), .B(a[518]), .Z(n2589) );
  XOR U3109 ( .A(sreg[1541]), .B(n2589), .Z(n2591) );
  NANDN U3110 ( .A(n2584), .B(sreg[1540]), .Z(n2588) );
  OR U3111 ( .A(n2586), .B(n2585), .Z(n2587) );
  AND U3112 ( .A(n2588), .B(n2587), .Z(n2590) );
  XOR U3113 ( .A(n2591), .B(n2590), .Z(c[1541]) );
  NAND U3114 ( .A(b[0]), .B(a[519]), .Z(n2594) );
  XOR U3115 ( .A(sreg[1542]), .B(n2594), .Z(n2596) );
  NANDN U3116 ( .A(n2589), .B(sreg[1541]), .Z(n2593) );
  OR U3117 ( .A(n2591), .B(n2590), .Z(n2592) );
  AND U3118 ( .A(n2593), .B(n2592), .Z(n2595) );
  XOR U3119 ( .A(n2596), .B(n2595), .Z(c[1542]) );
  NAND U3120 ( .A(b[0]), .B(a[520]), .Z(n2599) );
  XOR U3121 ( .A(sreg[1543]), .B(n2599), .Z(n2601) );
  NANDN U3122 ( .A(n2594), .B(sreg[1542]), .Z(n2598) );
  OR U3123 ( .A(n2596), .B(n2595), .Z(n2597) );
  AND U3124 ( .A(n2598), .B(n2597), .Z(n2600) );
  XOR U3125 ( .A(n2601), .B(n2600), .Z(c[1543]) );
  NAND U3126 ( .A(b[0]), .B(a[521]), .Z(n2604) );
  XOR U3127 ( .A(sreg[1544]), .B(n2604), .Z(n2606) );
  NANDN U3128 ( .A(n2599), .B(sreg[1543]), .Z(n2603) );
  OR U3129 ( .A(n2601), .B(n2600), .Z(n2602) );
  AND U3130 ( .A(n2603), .B(n2602), .Z(n2605) );
  XOR U3131 ( .A(n2606), .B(n2605), .Z(c[1544]) );
  NAND U3132 ( .A(b[0]), .B(a[522]), .Z(n2609) );
  XOR U3133 ( .A(sreg[1545]), .B(n2609), .Z(n2611) );
  NANDN U3134 ( .A(n2604), .B(sreg[1544]), .Z(n2608) );
  OR U3135 ( .A(n2606), .B(n2605), .Z(n2607) );
  AND U3136 ( .A(n2608), .B(n2607), .Z(n2610) );
  XOR U3137 ( .A(n2611), .B(n2610), .Z(c[1545]) );
  NAND U3138 ( .A(b[0]), .B(a[523]), .Z(n2614) );
  XOR U3139 ( .A(sreg[1546]), .B(n2614), .Z(n2616) );
  NANDN U3140 ( .A(n2609), .B(sreg[1545]), .Z(n2613) );
  OR U3141 ( .A(n2611), .B(n2610), .Z(n2612) );
  AND U3142 ( .A(n2613), .B(n2612), .Z(n2615) );
  XOR U3143 ( .A(n2616), .B(n2615), .Z(c[1546]) );
  NAND U3144 ( .A(b[0]), .B(a[524]), .Z(n2619) );
  XOR U3145 ( .A(sreg[1547]), .B(n2619), .Z(n2621) );
  NANDN U3146 ( .A(n2614), .B(sreg[1546]), .Z(n2618) );
  OR U3147 ( .A(n2616), .B(n2615), .Z(n2617) );
  AND U3148 ( .A(n2618), .B(n2617), .Z(n2620) );
  XOR U3149 ( .A(n2621), .B(n2620), .Z(c[1547]) );
  NAND U3150 ( .A(b[0]), .B(a[525]), .Z(n2624) );
  XOR U3151 ( .A(sreg[1548]), .B(n2624), .Z(n2626) );
  NANDN U3152 ( .A(n2619), .B(sreg[1547]), .Z(n2623) );
  OR U3153 ( .A(n2621), .B(n2620), .Z(n2622) );
  AND U3154 ( .A(n2623), .B(n2622), .Z(n2625) );
  XOR U3155 ( .A(n2626), .B(n2625), .Z(c[1548]) );
  NAND U3156 ( .A(b[0]), .B(a[526]), .Z(n2629) );
  XOR U3157 ( .A(sreg[1549]), .B(n2629), .Z(n2631) );
  NANDN U3158 ( .A(n2624), .B(sreg[1548]), .Z(n2628) );
  OR U3159 ( .A(n2626), .B(n2625), .Z(n2627) );
  AND U3160 ( .A(n2628), .B(n2627), .Z(n2630) );
  XOR U3161 ( .A(n2631), .B(n2630), .Z(c[1549]) );
  NAND U3162 ( .A(b[0]), .B(a[527]), .Z(n2634) );
  XOR U3163 ( .A(sreg[1550]), .B(n2634), .Z(n2636) );
  NANDN U3164 ( .A(n2629), .B(sreg[1549]), .Z(n2633) );
  OR U3165 ( .A(n2631), .B(n2630), .Z(n2632) );
  AND U3166 ( .A(n2633), .B(n2632), .Z(n2635) );
  XOR U3167 ( .A(n2636), .B(n2635), .Z(c[1550]) );
  NAND U3168 ( .A(b[0]), .B(a[528]), .Z(n2639) );
  XOR U3169 ( .A(sreg[1551]), .B(n2639), .Z(n2641) );
  NANDN U3170 ( .A(n2634), .B(sreg[1550]), .Z(n2638) );
  OR U3171 ( .A(n2636), .B(n2635), .Z(n2637) );
  AND U3172 ( .A(n2638), .B(n2637), .Z(n2640) );
  XOR U3173 ( .A(n2641), .B(n2640), .Z(c[1551]) );
  NAND U3174 ( .A(b[0]), .B(a[529]), .Z(n2644) );
  XOR U3175 ( .A(sreg[1552]), .B(n2644), .Z(n2646) );
  NANDN U3176 ( .A(n2639), .B(sreg[1551]), .Z(n2643) );
  OR U3177 ( .A(n2641), .B(n2640), .Z(n2642) );
  AND U3178 ( .A(n2643), .B(n2642), .Z(n2645) );
  XOR U3179 ( .A(n2646), .B(n2645), .Z(c[1552]) );
  NAND U3180 ( .A(b[0]), .B(a[530]), .Z(n2649) );
  XOR U3181 ( .A(sreg[1553]), .B(n2649), .Z(n2651) );
  NANDN U3182 ( .A(n2644), .B(sreg[1552]), .Z(n2648) );
  OR U3183 ( .A(n2646), .B(n2645), .Z(n2647) );
  AND U3184 ( .A(n2648), .B(n2647), .Z(n2650) );
  XOR U3185 ( .A(n2651), .B(n2650), .Z(c[1553]) );
  NAND U3186 ( .A(b[0]), .B(a[531]), .Z(n2654) );
  XOR U3187 ( .A(sreg[1554]), .B(n2654), .Z(n2656) );
  NANDN U3188 ( .A(n2649), .B(sreg[1553]), .Z(n2653) );
  OR U3189 ( .A(n2651), .B(n2650), .Z(n2652) );
  AND U3190 ( .A(n2653), .B(n2652), .Z(n2655) );
  XOR U3191 ( .A(n2656), .B(n2655), .Z(c[1554]) );
  NAND U3192 ( .A(b[0]), .B(a[532]), .Z(n2659) );
  XOR U3193 ( .A(sreg[1555]), .B(n2659), .Z(n2661) );
  NANDN U3194 ( .A(n2654), .B(sreg[1554]), .Z(n2658) );
  OR U3195 ( .A(n2656), .B(n2655), .Z(n2657) );
  AND U3196 ( .A(n2658), .B(n2657), .Z(n2660) );
  XOR U3197 ( .A(n2661), .B(n2660), .Z(c[1555]) );
  NAND U3198 ( .A(b[0]), .B(a[533]), .Z(n2664) );
  XOR U3199 ( .A(sreg[1556]), .B(n2664), .Z(n2666) );
  NANDN U3200 ( .A(n2659), .B(sreg[1555]), .Z(n2663) );
  OR U3201 ( .A(n2661), .B(n2660), .Z(n2662) );
  AND U3202 ( .A(n2663), .B(n2662), .Z(n2665) );
  XOR U3203 ( .A(n2666), .B(n2665), .Z(c[1556]) );
  NAND U3204 ( .A(b[0]), .B(a[534]), .Z(n2669) );
  XOR U3205 ( .A(sreg[1557]), .B(n2669), .Z(n2671) );
  NANDN U3206 ( .A(n2664), .B(sreg[1556]), .Z(n2668) );
  OR U3207 ( .A(n2666), .B(n2665), .Z(n2667) );
  AND U3208 ( .A(n2668), .B(n2667), .Z(n2670) );
  XOR U3209 ( .A(n2671), .B(n2670), .Z(c[1557]) );
  NAND U3210 ( .A(b[0]), .B(a[535]), .Z(n2674) );
  XOR U3211 ( .A(sreg[1558]), .B(n2674), .Z(n2676) );
  NANDN U3212 ( .A(n2669), .B(sreg[1557]), .Z(n2673) );
  OR U3213 ( .A(n2671), .B(n2670), .Z(n2672) );
  AND U3214 ( .A(n2673), .B(n2672), .Z(n2675) );
  XOR U3215 ( .A(n2676), .B(n2675), .Z(c[1558]) );
  NAND U3216 ( .A(b[0]), .B(a[536]), .Z(n2679) );
  XOR U3217 ( .A(sreg[1559]), .B(n2679), .Z(n2681) );
  NANDN U3218 ( .A(n2674), .B(sreg[1558]), .Z(n2678) );
  OR U3219 ( .A(n2676), .B(n2675), .Z(n2677) );
  AND U3220 ( .A(n2678), .B(n2677), .Z(n2680) );
  XOR U3221 ( .A(n2681), .B(n2680), .Z(c[1559]) );
  NAND U3222 ( .A(b[0]), .B(a[537]), .Z(n2684) );
  XOR U3223 ( .A(sreg[1560]), .B(n2684), .Z(n2686) );
  NANDN U3224 ( .A(n2679), .B(sreg[1559]), .Z(n2683) );
  OR U3225 ( .A(n2681), .B(n2680), .Z(n2682) );
  AND U3226 ( .A(n2683), .B(n2682), .Z(n2685) );
  XOR U3227 ( .A(n2686), .B(n2685), .Z(c[1560]) );
  NAND U3228 ( .A(b[0]), .B(a[538]), .Z(n2689) );
  XOR U3229 ( .A(sreg[1561]), .B(n2689), .Z(n2691) );
  NANDN U3230 ( .A(n2684), .B(sreg[1560]), .Z(n2688) );
  OR U3231 ( .A(n2686), .B(n2685), .Z(n2687) );
  AND U3232 ( .A(n2688), .B(n2687), .Z(n2690) );
  XOR U3233 ( .A(n2691), .B(n2690), .Z(c[1561]) );
  NAND U3234 ( .A(b[0]), .B(a[539]), .Z(n2694) );
  XOR U3235 ( .A(sreg[1562]), .B(n2694), .Z(n2696) );
  NANDN U3236 ( .A(n2689), .B(sreg[1561]), .Z(n2693) );
  OR U3237 ( .A(n2691), .B(n2690), .Z(n2692) );
  AND U3238 ( .A(n2693), .B(n2692), .Z(n2695) );
  XOR U3239 ( .A(n2696), .B(n2695), .Z(c[1562]) );
  NAND U3240 ( .A(b[0]), .B(a[540]), .Z(n2699) );
  XOR U3241 ( .A(sreg[1563]), .B(n2699), .Z(n2701) );
  NANDN U3242 ( .A(n2694), .B(sreg[1562]), .Z(n2698) );
  OR U3243 ( .A(n2696), .B(n2695), .Z(n2697) );
  AND U3244 ( .A(n2698), .B(n2697), .Z(n2700) );
  XOR U3245 ( .A(n2701), .B(n2700), .Z(c[1563]) );
  NAND U3246 ( .A(b[0]), .B(a[541]), .Z(n2704) );
  XOR U3247 ( .A(sreg[1564]), .B(n2704), .Z(n2706) );
  NANDN U3248 ( .A(n2699), .B(sreg[1563]), .Z(n2703) );
  OR U3249 ( .A(n2701), .B(n2700), .Z(n2702) );
  AND U3250 ( .A(n2703), .B(n2702), .Z(n2705) );
  XOR U3251 ( .A(n2706), .B(n2705), .Z(c[1564]) );
  NAND U3252 ( .A(b[0]), .B(a[542]), .Z(n2709) );
  XOR U3253 ( .A(sreg[1565]), .B(n2709), .Z(n2711) );
  NANDN U3254 ( .A(n2704), .B(sreg[1564]), .Z(n2708) );
  OR U3255 ( .A(n2706), .B(n2705), .Z(n2707) );
  AND U3256 ( .A(n2708), .B(n2707), .Z(n2710) );
  XOR U3257 ( .A(n2711), .B(n2710), .Z(c[1565]) );
  NAND U3258 ( .A(b[0]), .B(a[543]), .Z(n2714) );
  XOR U3259 ( .A(sreg[1566]), .B(n2714), .Z(n2716) );
  NANDN U3260 ( .A(n2709), .B(sreg[1565]), .Z(n2713) );
  OR U3261 ( .A(n2711), .B(n2710), .Z(n2712) );
  AND U3262 ( .A(n2713), .B(n2712), .Z(n2715) );
  XOR U3263 ( .A(n2716), .B(n2715), .Z(c[1566]) );
  NAND U3264 ( .A(b[0]), .B(a[544]), .Z(n2719) );
  XOR U3265 ( .A(sreg[1567]), .B(n2719), .Z(n2721) );
  NANDN U3266 ( .A(n2714), .B(sreg[1566]), .Z(n2718) );
  OR U3267 ( .A(n2716), .B(n2715), .Z(n2717) );
  AND U3268 ( .A(n2718), .B(n2717), .Z(n2720) );
  XOR U3269 ( .A(n2721), .B(n2720), .Z(c[1567]) );
  NAND U3270 ( .A(b[0]), .B(a[545]), .Z(n2724) );
  XOR U3271 ( .A(sreg[1568]), .B(n2724), .Z(n2726) );
  NANDN U3272 ( .A(n2719), .B(sreg[1567]), .Z(n2723) );
  OR U3273 ( .A(n2721), .B(n2720), .Z(n2722) );
  AND U3274 ( .A(n2723), .B(n2722), .Z(n2725) );
  XOR U3275 ( .A(n2726), .B(n2725), .Z(c[1568]) );
  NAND U3276 ( .A(b[0]), .B(a[546]), .Z(n2729) );
  XOR U3277 ( .A(sreg[1569]), .B(n2729), .Z(n2731) );
  NANDN U3278 ( .A(n2724), .B(sreg[1568]), .Z(n2728) );
  OR U3279 ( .A(n2726), .B(n2725), .Z(n2727) );
  AND U3280 ( .A(n2728), .B(n2727), .Z(n2730) );
  XOR U3281 ( .A(n2731), .B(n2730), .Z(c[1569]) );
  NAND U3282 ( .A(b[0]), .B(a[547]), .Z(n2734) );
  XOR U3283 ( .A(sreg[1570]), .B(n2734), .Z(n2736) );
  NANDN U3284 ( .A(n2729), .B(sreg[1569]), .Z(n2733) );
  OR U3285 ( .A(n2731), .B(n2730), .Z(n2732) );
  AND U3286 ( .A(n2733), .B(n2732), .Z(n2735) );
  XOR U3287 ( .A(n2736), .B(n2735), .Z(c[1570]) );
  NAND U3288 ( .A(b[0]), .B(a[548]), .Z(n2739) );
  XOR U3289 ( .A(sreg[1571]), .B(n2739), .Z(n2741) );
  NANDN U3290 ( .A(n2734), .B(sreg[1570]), .Z(n2738) );
  OR U3291 ( .A(n2736), .B(n2735), .Z(n2737) );
  AND U3292 ( .A(n2738), .B(n2737), .Z(n2740) );
  XOR U3293 ( .A(n2741), .B(n2740), .Z(c[1571]) );
  NAND U3294 ( .A(b[0]), .B(a[549]), .Z(n2744) );
  XOR U3295 ( .A(sreg[1572]), .B(n2744), .Z(n2746) );
  NANDN U3296 ( .A(n2739), .B(sreg[1571]), .Z(n2743) );
  OR U3297 ( .A(n2741), .B(n2740), .Z(n2742) );
  AND U3298 ( .A(n2743), .B(n2742), .Z(n2745) );
  XOR U3299 ( .A(n2746), .B(n2745), .Z(c[1572]) );
  NAND U3300 ( .A(b[0]), .B(a[550]), .Z(n2749) );
  XOR U3301 ( .A(sreg[1573]), .B(n2749), .Z(n2751) );
  NANDN U3302 ( .A(n2744), .B(sreg[1572]), .Z(n2748) );
  OR U3303 ( .A(n2746), .B(n2745), .Z(n2747) );
  AND U3304 ( .A(n2748), .B(n2747), .Z(n2750) );
  XOR U3305 ( .A(n2751), .B(n2750), .Z(c[1573]) );
  NAND U3306 ( .A(b[0]), .B(a[551]), .Z(n2754) );
  XOR U3307 ( .A(sreg[1574]), .B(n2754), .Z(n2756) );
  NANDN U3308 ( .A(n2749), .B(sreg[1573]), .Z(n2753) );
  OR U3309 ( .A(n2751), .B(n2750), .Z(n2752) );
  AND U3310 ( .A(n2753), .B(n2752), .Z(n2755) );
  XOR U3311 ( .A(n2756), .B(n2755), .Z(c[1574]) );
  NAND U3312 ( .A(b[0]), .B(a[552]), .Z(n2759) );
  XOR U3313 ( .A(sreg[1575]), .B(n2759), .Z(n2761) );
  NANDN U3314 ( .A(n2754), .B(sreg[1574]), .Z(n2758) );
  OR U3315 ( .A(n2756), .B(n2755), .Z(n2757) );
  AND U3316 ( .A(n2758), .B(n2757), .Z(n2760) );
  XOR U3317 ( .A(n2761), .B(n2760), .Z(c[1575]) );
  NAND U3318 ( .A(b[0]), .B(a[553]), .Z(n2764) );
  XOR U3319 ( .A(sreg[1576]), .B(n2764), .Z(n2766) );
  NANDN U3320 ( .A(n2759), .B(sreg[1575]), .Z(n2763) );
  OR U3321 ( .A(n2761), .B(n2760), .Z(n2762) );
  AND U3322 ( .A(n2763), .B(n2762), .Z(n2765) );
  XOR U3323 ( .A(n2766), .B(n2765), .Z(c[1576]) );
  NAND U3324 ( .A(b[0]), .B(a[554]), .Z(n2769) );
  XOR U3325 ( .A(sreg[1577]), .B(n2769), .Z(n2771) );
  NANDN U3326 ( .A(n2764), .B(sreg[1576]), .Z(n2768) );
  OR U3327 ( .A(n2766), .B(n2765), .Z(n2767) );
  AND U3328 ( .A(n2768), .B(n2767), .Z(n2770) );
  XOR U3329 ( .A(n2771), .B(n2770), .Z(c[1577]) );
  NAND U3330 ( .A(b[0]), .B(a[555]), .Z(n2774) );
  XOR U3331 ( .A(sreg[1578]), .B(n2774), .Z(n2776) );
  NANDN U3332 ( .A(n2769), .B(sreg[1577]), .Z(n2773) );
  OR U3333 ( .A(n2771), .B(n2770), .Z(n2772) );
  AND U3334 ( .A(n2773), .B(n2772), .Z(n2775) );
  XOR U3335 ( .A(n2776), .B(n2775), .Z(c[1578]) );
  NAND U3336 ( .A(b[0]), .B(a[556]), .Z(n2779) );
  XOR U3337 ( .A(sreg[1579]), .B(n2779), .Z(n2781) );
  NANDN U3338 ( .A(n2774), .B(sreg[1578]), .Z(n2778) );
  OR U3339 ( .A(n2776), .B(n2775), .Z(n2777) );
  AND U3340 ( .A(n2778), .B(n2777), .Z(n2780) );
  XOR U3341 ( .A(n2781), .B(n2780), .Z(c[1579]) );
  NAND U3342 ( .A(b[0]), .B(a[557]), .Z(n2784) );
  XOR U3343 ( .A(sreg[1580]), .B(n2784), .Z(n2786) );
  NANDN U3344 ( .A(n2779), .B(sreg[1579]), .Z(n2783) );
  OR U3345 ( .A(n2781), .B(n2780), .Z(n2782) );
  AND U3346 ( .A(n2783), .B(n2782), .Z(n2785) );
  XOR U3347 ( .A(n2786), .B(n2785), .Z(c[1580]) );
  NAND U3348 ( .A(b[0]), .B(a[558]), .Z(n2789) );
  XOR U3349 ( .A(sreg[1581]), .B(n2789), .Z(n2791) );
  NANDN U3350 ( .A(n2784), .B(sreg[1580]), .Z(n2788) );
  OR U3351 ( .A(n2786), .B(n2785), .Z(n2787) );
  AND U3352 ( .A(n2788), .B(n2787), .Z(n2790) );
  XOR U3353 ( .A(n2791), .B(n2790), .Z(c[1581]) );
  NAND U3354 ( .A(b[0]), .B(a[559]), .Z(n2794) );
  XOR U3355 ( .A(sreg[1582]), .B(n2794), .Z(n2796) );
  NANDN U3356 ( .A(n2789), .B(sreg[1581]), .Z(n2793) );
  OR U3357 ( .A(n2791), .B(n2790), .Z(n2792) );
  AND U3358 ( .A(n2793), .B(n2792), .Z(n2795) );
  XOR U3359 ( .A(n2796), .B(n2795), .Z(c[1582]) );
  NAND U3360 ( .A(b[0]), .B(a[560]), .Z(n2799) );
  XOR U3361 ( .A(sreg[1583]), .B(n2799), .Z(n2801) );
  NANDN U3362 ( .A(n2794), .B(sreg[1582]), .Z(n2798) );
  OR U3363 ( .A(n2796), .B(n2795), .Z(n2797) );
  AND U3364 ( .A(n2798), .B(n2797), .Z(n2800) );
  XOR U3365 ( .A(n2801), .B(n2800), .Z(c[1583]) );
  NAND U3366 ( .A(b[0]), .B(a[561]), .Z(n2804) );
  XOR U3367 ( .A(sreg[1584]), .B(n2804), .Z(n2806) );
  NANDN U3368 ( .A(n2799), .B(sreg[1583]), .Z(n2803) );
  OR U3369 ( .A(n2801), .B(n2800), .Z(n2802) );
  AND U3370 ( .A(n2803), .B(n2802), .Z(n2805) );
  XOR U3371 ( .A(n2806), .B(n2805), .Z(c[1584]) );
  NAND U3372 ( .A(b[0]), .B(a[562]), .Z(n2809) );
  XOR U3373 ( .A(sreg[1585]), .B(n2809), .Z(n2811) );
  NANDN U3374 ( .A(n2804), .B(sreg[1584]), .Z(n2808) );
  OR U3375 ( .A(n2806), .B(n2805), .Z(n2807) );
  AND U3376 ( .A(n2808), .B(n2807), .Z(n2810) );
  XOR U3377 ( .A(n2811), .B(n2810), .Z(c[1585]) );
  NAND U3378 ( .A(b[0]), .B(a[563]), .Z(n2814) );
  XOR U3379 ( .A(sreg[1586]), .B(n2814), .Z(n2816) );
  NANDN U3380 ( .A(n2809), .B(sreg[1585]), .Z(n2813) );
  OR U3381 ( .A(n2811), .B(n2810), .Z(n2812) );
  AND U3382 ( .A(n2813), .B(n2812), .Z(n2815) );
  XOR U3383 ( .A(n2816), .B(n2815), .Z(c[1586]) );
  NAND U3384 ( .A(b[0]), .B(a[564]), .Z(n2819) );
  XOR U3385 ( .A(sreg[1587]), .B(n2819), .Z(n2821) );
  NANDN U3386 ( .A(n2814), .B(sreg[1586]), .Z(n2818) );
  OR U3387 ( .A(n2816), .B(n2815), .Z(n2817) );
  AND U3388 ( .A(n2818), .B(n2817), .Z(n2820) );
  XOR U3389 ( .A(n2821), .B(n2820), .Z(c[1587]) );
  NAND U3390 ( .A(b[0]), .B(a[565]), .Z(n2824) );
  XOR U3391 ( .A(sreg[1588]), .B(n2824), .Z(n2826) );
  NANDN U3392 ( .A(n2819), .B(sreg[1587]), .Z(n2823) );
  OR U3393 ( .A(n2821), .B(n2820), .Z(n2822) );
  AND U3394 ( .A(n2823), .B(n2822), .Z(n2825) );
  XOR U3395 ( .A(n2826), .B(n2825), .Z(c[1588]) );
  NAND U3396 ( .A(b[0]), .B(a[566]), .Z(n2829) );
  XOR U3397 ( .A(sreg[1589]), .B(n2829), .Z(n2831) );
  NANDN U3398 ( .A(n2824), .B(sreg[1588]), .Z(n2828) );
  OR U3399 ( .A(n2826), .B(n2825), .Z(n2827) );
  AND U3400 ( .A(n2828), .B(n2827), .Z(n2830) );
  XOR U3401 ( .A(n2831), .B(n2830), .Z(c[1589]) );
  NAND U3402 ( .A(b[0]), .B(a[567]), .Z(n2834) );
  XOR U3403 ( .A(sreg[1590]), .B(n2834), .Z(n2836) );
  NANDN U3404 ( .A(n2829), .B(sreg[1589]), .Z(n2833) );
  OR U3405 ( .A(n2831), .B(n2830), .Z(n2832) );
  AND U3406 ( .A(n2833), .B(n2832), .Z(n2835) );
  XOR U3407 ( .A(n2836), .B(n2835), .Z(c[1590]) );
  NAND U3408 ( .A(b[0]), .B(a[568]), .Z(n2839) );
  XOR U3409 ( .A(sreg[1591]), .B(n2839), .Z(n2841) );
  NANDN U3410 ( .A(n2834), .B(sreg[1590]), .Z(n2838) );
  OR U3411 ( .A(n2836), .B(n2835), .Z(n2837) );
  AND U3412 ( .A(n2838), .B(n2837), .Z(n2840) );
  XOR U3413 ( .A(n2841), .B(n2840), .Z(c[1591]) );
  NAND U3414 ( .A(b[0]), .B(a[569]), .Z(n2844) );
  XOR U3415 ( .A(sreg[1592]), .B(n2844), .Z(n2846) );
  NANDN U3416 ( .A(n2839), .B(sreg[1591]), .Z(n2843) );
  OR U3417 ( .A(n2841), .B(n2840), .Z(n2842) );
  AND U3418 ( .A(n2843), .B(n2842), .Z(n2845) );
  XOR U3419 ( .A(n2846), .B(n2845), .Z(c[1592]) );
  NAND U3420 ( .A(b[0]), .B(a[570]), .Z(n2849) );
  XOR U3421 ( .A(sreg[1593]), .B(n2849), .Z(n2851) );
  NANDN U3422 ( .A(n2844), .B(sreg[1592]), .Z(n2848) );
  OR U3423 ( .A(n2846), .B(n2845), .Z(n2847) );
  AND U3424 ( .A(n2848), .B(n2847), .Z(n2850) );
  XOR U3425 ( .A(n2851), .B(n2850), .Z(c[1593]) );
  NAND U3426 ( .A(b[0]), .B(a[571]), .Z(n2854) );
  XOR U3427 ( .A(sreg[1594]), .B(n2854), .Z(n2856) );
  NANDN U3428 ( .A(n2849), .B(sreg[1593]), .Z(n2853) );
  OR U3429 ( .A(n2851), .B(n2850), .Z(n2852) );
  AND U3430 ( .A(n2853), .B(n2852), .Z(n2855) );
  XOR U3431 ( .A(n2856), .B(n2855), .Z(c[1594]) );
  NAND U3432 ( .A(b[0]), .B(a[572]), .Z(n2859) );
  XOR U3433 ( .A(sreg[1595]), .B(n2859), .Z(n2861) );
  NANDN U3434 ( .A(n2854), .B(sreg[1594]), .Z(n2858) );
  OR U3435 ( .A(n2856), .B(n2855), .Z(n2857) );
  AND U3436 ( .A(n2858), .B(n2857), .Z(n2860) );
  XOR U3437 ( .A(n2861), .B(n2860), .Z(c[1595]) );
  NAND U3438 ( .A(b[0]), .B(a[573]), .Z(n2864) );
  XOR U3439 ( .A(sreg[1596]), .B(n2864), .Z(n2866) );
  NANDN U3440 ( .A(n2859), .B(sreg[1595]), .Z(n2863) );
  OR U3441 ( .A(n2861), .B(n2860), .Z(n2862) );
  AND U3442 ( .A(n2863), .B(n2862), .Z(n2865) );
  XOR U3443 ( .A(n2866), .B(n2865), .Z(c[1596]) );
  NAND U3444 ( .A(b[0]), .B(a[574]), .Z(n2869) );
  XOR U3445 ( .A(sreg[1597]), .B(n2869), .Z(n2871) );
  NANDN U3446 ( .A(n2864), .B(sreg[1596]), .Z(n2868) );
  OR U3447 ( .A(n2866), .B(n2865), .Z(n2867) );
  AND U3448 ( .A(n2868), .B(n2867), .Z(n2870) );
  XOR U3449 ( .A(n2871), .B(n2870), .Z(c[1597]) );
  NAND U3450 ( .A(b[0]), .B(a[575]), .Z(n2874) );
  XOR U3451 ( .A(sreg[1598]), .B(n2874), .Z(n2876) );
  NANDN U3452 ( .A(n2869), .B(sreg[1597]), .Z(n2873) );
  OR U3453 ( .A(n2871), .B(n2870), .Z(n2872) );
  AND U3454 ( .A(n2873), .B(n2872), .Z(n2875) );
  XOR U3455 ( .A(n2876), .B(n2875), .Z(c[1598]) );
  NAND U3456 ( .A(b[0]), .B(a[576]), .Z(n2879) );
  XOR U3457 ( .A(sreg[1599]), .B(n2879), .Z(n2881) );
  NANDN U3458 ( .A(n2874), .B(sreg[1598]), .Z(n2878) );
  OR U3459 ( .A(n2876), .B(n2875), .Z(n2877) );
  AND U3460 ( .A(n2878), .B(n2877), .Z(n2880) );
  XOR U3461 ( .A(n2881), .B(n2880), .Z(c[1599]) );
  NAND U3462 ( .A(b[0]), .B(a[577]), .Z(n2884) );
  XOR U3463 ( .A(sreg[1600]), .B(n2884), .Z(n2886) );
  NANDN U3464 ( .A(n2879), .B(sreg[1599]), .Z(n2883) );
  OR U3465 ( .A(n2881), .B(n2880), .Z(n2882) );
  AND U3466 ( .A(n2883), .B(n2882), .Z(n2885) );
  XOR U3467 ( .A(n2886), .B(n2885), .Z(c[1600]) );
  NAND U3468 ( .A(b[0]), .B(a[578]), .Z(n2889) );
  XOR U3469 ( .A(sreg[1601]), .B(n2889), .Z(n2891) );
  NANDN U3470 ( .A(n2884), .B(sreg[1600]), .Z(n2888) );
  OR U3471 ( .A(n2886), .B(n2885), .Z(n2887) );
  AND U3472 ( .A(n2888), .B(n2887), .Z(n2890) );
  XOR U3473 ( .A(n2891), .B(n2890), .Z(c[1601]) );
  NAND U3474 ( .A(b[0]), .B(a[579]), .Z(n2894) );
  XOR U3475 ( .A(sreg[1602]), .B(n2894), .Z(n2896) );
  NANDN U3476 ( .A(n2889), .B(sreg[1601]), .Z(n2893) );
  OR U3477 ( .A(n2891), .B(n2890), .Z(n2892) );
  AND U3478 ( .A(n2893), .B(n2892), .Z(n2895) );
  XOR U3479 ( .A(n2896), .B(n2895), .Z(c[1602]) );
  NAND U3480 ( .A(b[0]), .B(a[580]), .Z(n2899) );
  XOR U3481 ( .A(sreg[1603]), .B(n2899), .Z(n2901) );
  NANDN U3482 ( .A(n2894), .B(sreg[1602]), .Z(n2898) );
  OR U3483 ( .A(n2896), .B(n2895), .Z(n2897) );
  AND U3484 ( .A(n2898), .B(n2897), .Z(n2900) );
  XOR U3485 ( .A(n2901), .B(n2900), .Z(c[1603]) );
  NAND U3486 ( .A(b[0]), .B(a[581]), .Z(n2904) );
  XOR U3487 ( .A(sreg[1604]), .B(n2904), .Z(n2906) );
  NANDN U3488 ( .A(n2899), .B(sreg[1603]), .Z(n2903) );
  OR U3489 ( .A(n2901), .B(n2900), .Z(n2902) );
  AND U3490 ( .A(n2903), .B(n2902), .Z(n2905) );
  XOR U3491 ( .A(n2906), .B(n2905), .Z(c[1604]) );
  NAND U3492 ( .A(b[0]), .B(a[582]), .Z(n2909) );
  XOR U3493 ( .A(sreg[1605]), .B(n2909), .Z(n2911) );
  NANDN U3494 ( .A(n2904), .B(sreg[1604]), .Z(n2908) );
  OR U3495 ( .A(n2906), .B(n2905), .Z(n2907) );
  AND U3496 ( .A(n2908), .B(n2907), .Z(n2910) );
  XOR U3497 ( .A(n2911), .B(n2910), .Z(c[1605]) );
  NAND U3498 ( .A(b[0]), .B(a[583]), .Z(n2914) );
  XOR U3499 ( .A(sreg[1606]), .B(n2914), .Z(n2916) );
  NANDN U3500 ( .A(n2909), .B(sreg[1605]), .Z(n2913) );
  OR U3501 ( .A(n2911), .B(n2910), .Z(n2912) );
  AND U3502 ( .A(n2913), .B(n2912), .Z(n2915) );
  XOR U3503 ( .A(n2916), .B(n2915), .Z(c[1606]) );
  NAND U3504 ( .A(b[0]), .B(a[584]), .Z(n2919) );
  XOR U3505 ( .A(sreg[1607]), .B(n2919), .Z(n2921) );
  NANDN U3506 ( .A(n2914), .B(sreg[1606]), .Z(n2918) );
  OR U3507 ( .A(n2916), .B(n2915), .Z(n2917) );
  AND U3508 ( .A(n2918), .B(n2917), .Z(n2920) );
  XOR U3509 ( .A(n2921), .B(n2920), .Z(c[1607]) );
  NAND U3510 ( .A(b[0]), .B(a[585]), .Z(n2924) );
  XOR U3511 ( .A(sreg[1608]), .B(n2924), .Z(n2926) );
  NANDN U3512 ( .A(n2919), .B(sreg[1607]), .Z(n2923) );
  OR U3513 ( .A(n2921), .B(n2920), .Z(n2922) );
  AND U3514 ( .A(n2923), .B(n2922), .Z(n2925) );
  XOR U3515 ( .A(n2926), .B(n2925), .Z(c[1608]) );
  NAND U3516 ( .A(b[0]), .B(a[586]), .Z(n2929) );
  XOR U3517 ( .A(sreg[1609]), .B(n2929), .Z(n2931) );
  NANDN U3518 ( .A(n2924), .B(sreg[1608]), .Z(n2928) );
  OR U3519 ( .A(n2926), .B(n2925), .Z(n2927) );
  AND U3520 ( .A(n2928), .B(n2927), .Z(n2930) );
  XOR U3521 ( .A(n2931), .B(n2930), .Z(c[1609]) );
  NAND U3522 ( .A(b[0]), .B(a[587]), .Z(n2934) );
  XOR U3523 ( .A(sreg[1610]), .B(n2934), .Z(n2936) );
  NANDN U3524 ( .A(n2929), .B(sreg[1609]), .Z(n2933) );
  OR U3525 ( .A(n2931), .B(n2930), .Z(n2932) );
  AND U3526 ( .A(n2933), .B(n2932), .Z(n2935) );
  XOR U3527 ( .A(n2936), .B(n2935), .Z(c[1610]) );
  NAND U3528 ( .A(b[0]), .B(a[588]), .Z(n2939) );
  XOR U3529 ( .A(sreg[1611]), .B(n2939), .Z(n2941) );
  NANDN U3530 ( .A(n2934), .B(sreg[1610]), .Z(n2938) );
  OR U3531 ( .A(n2936), .B(n2935), .Z(n2937) );
  AND U3532 ( .A(n2938), .B(n2937), .Z(n2940) );
  XOR U3533 ( .A(n2941), .B(n2940), .Z(c[1611]) );
  NAND U3534 ( .A(b[0]), .B(a[589]), .Z(n2944) );
  XOR U3535 ( .A(sreg[1612]), .B(n2944), .Z(n2946) );
  NANDN U3536 ( .A(n2939), .B(sreg[1611]), .Z(n2943) );
  OR U3537 ( .A(n2941), .B(n2940), .Z(n2942) );
  AND U3538 ( .A(n2943), .B(n2942), .Z(n2945) );
  XOR U3539 ( .A(n2946), .B(n2945), .Z(c[1612]) );
  NAND U3540 ( .A(b[0]), .B(a[590]), .Z(n2949) );
  XOR U3541 ( .A(sreg[1613]), .B(n2949), .Z(n2951) );
  NANDN U3542 ( .A(n2944), .B(sreg[1612]), .Z(n2948) );
  OR U3543 ( .A(n2946), .B(n2945), .Z(n2947) );
  AND U3544 ( .A(n2948), .B(n2947), .Z(n2950) );
  XOR U3545 ( .A(n2951), .B(n2950), .Z(c[1613]) );
  NAND U3546 ( .A(b[0]), .B(a[591]), .Z(n2954) );
  XOR U3547 ( .A(sreg[1614]), .B(n2954), .Z(n2956) );
  NANDN U3548 ( .A(n2949), .B(sreg[1613]), .Z(n2953) );
  OR U3549 ( .A(n2951), .B(n2950), .Z(n2952) );
  AND U3550 ( .A(n2953), .B(n2952), .Z(n2955) );
  XOR U3551 ( .A(n2956), .B(n2955), .Z(c[1614]) );
  NAND U3552 ( .A(b[0]), .B(a[592]), .Z(n2959) );
  XOR U3553 ( .A(sreg[1615]), .B(n2959), .Z(n2961) );
  NANDN U3554 ( .A(n2954), .B(sreg[1614]), .Z(n2958) );
  OR U3555 ( .A(n2956), .B(n2955), .Z(n2957) );
  AND U3556 ( .A(n2958), .B(n2957), .Z(n2960) );
  XOR U3557 ( .A(n2961), .B(n2960), .Z(c[1615]) );
  NAND U3558 ( .A(b[0]), .B(a[593]), .Z(n2964) );
  XOR U3559 ( .A(sreg[1616]), .B(n2964), .Z(n2966) );
  NANDN U3560 ( .A(n2959), .B(sreg[1615]), .Z(n2963) );
  OR U3561 ( .A(n2961), .B(n2960), .Z(n2962) );
  AND U3562 ( .A(n2963), .B(n2962), .Z(n2965) );
  XOR U3563 ( .A(n2966), .B(n2965), .Z(c[1616]) );
  NAND U3564 ( .A(b[0]), .B(a[594]), .Z(n2969) );
  XOR U3565 ( .A(sreg[1617]), .B(n2969), .Z(n2971) );
  NANDN U3566 ( .A(n2964), .B(sreg[1616]), .Z(n2968) );
  OR U3567 ( .A(n2966), .B(n2965), .Z(n2967) );
  AND U3568 ( .A(n2968), .B(n2967), .Z(n2970) );
  XOR U3569 ( .A(n2971), .B(n2970), .Z(c[1617]) );
  NAND U3570 ( .A(b[0]), .B(a[595]), .Z(n2974) );
  XOR U3571 ( .A(sreg[1618]), .B(n2974), .Z(n2976) );
  NANDN U3572 ( .A(n2969), .B(sreg[1617]), .Z(n2973) );
  OR U3573 ( .A(n2971), .B(n2970), .Z(n2972) );
  AND U3574 ( .A(n2973), .B(n2972), .Z(n2975) );
  XOR U3575 ( .A(n2976), .B(n2975), .Z(c[1618]) );
  NAND U3576 ( .A(b[0]), .B(a[596]), .Z(n2979) );
  XOR U3577 ( .A(sreg[1619]), .B(n2979), .Z(n2981) );
  NANDN U3578 ( .A(n2974), .B(sreg[1618]), .Z(n2978) );
  OR U3579 ( .A(n2976), .B(n2975), .Z(n2977) );
  AND U3580 ( .A(n2978), .B(n2977), .Z(n2980) );
  XOR U3581 ( .A(n2981), .B(n2980), .Z(c[1619]) );
  NAND U3582 ( .A(b[0]), .B(a[597]), .Z(n2984) );
  XOR U3583 ( .A(sreg[1620]), .B(n2984), .Z(n2986) );
  NANDN U3584 ( .A(n2979), .B(sreg[1619]), .Z(n2983) );
  OR U3585 ( .A(n2981), .B(n2980), .Z(n2982) );
  AND U3586 ( .A(n2983), .B(n2982), .Z(n2985) );
  XOR U3587 ( .A(n2986), .B(n2985), .Z(c[1620]) );
  NAND U3588 ( .A(b[0]), .B(a[598]), .Z(n2989) );
  XOR U3589 ( .A(sreg[1621]), .B(n2989), .Z(n2991) );
  NANDN U3590 ( .A(n2984), .B(sreg[1620]), .Z(n2988) );
  OR U3591 ( .A(n2986), .B(n2985), .Z(n2987) );
  AND U3592 ( .A(n2988), .B(n2987), .Z(n2990) );
  XOR U3593 ( .A(n2991), .B(n2990), .Z(c[1621]) );
  NAND U3594 ( .A(b[0]), .B(a[599]), .Z(n2994) );
  XOR U3595 ( .A(sreg[1622]), .B(n2994), .Z(n2996) );
  NANDN U3596 ( .A(n2989), .B(sreg[1621]), .Z(n2993) );
  OR U3597 ( .A(n2991), .B(n2990), .Z(n2992) );
  AND U3598 ( .A(n2993), .B(n2992), .Z(n2995) );
  XOR U3599 ( .A(n2996), .B(n2995), .Z(c[1622]) );
  NAND U3600 ( .A(b[0]), .B(a[600]), .Z(n2999) );
  XOR U3601 ( .A(sreg[1623]), .B(n2999), .Z(n3001) );
  NANDN U3602 ( .A(n2994), .B(sreg[1622]), .Z(n2998) );
  OR U3603 ( .A(n2996), .B(n2995), .Z(n2997) );
  AND U3604 ( .A(n2998), .B(n2997), .Z(n3000) );
  XOR U3605 ( .A(n3001), .B(n3000), .Z(c[1623]) );
  NAND U3606 ( .A(b[0]), .B(a[601]), .Z(n3004) );
  XOR U3607 ( .A(sreg[1624]), .B(n3004), .Z(n3006) );
  NANDN U3608 ( .A(n2999), .B(sreg[1623]), .Z(n3003) );
  OR U3609 ( .A(n3001), .B(n3000), .Z(n3002) );
  AND U3610 ( .A(n3003), .B(n3002), .Z(n3005) );
  XOR U3611 ( .A(n3006), .B(n3005), .Z(c[1624]) );
  NAND U3612 ( .A(b[0]), .B(a[602]), .Z(n3009) );
  XOR U3613 ( .A(sreg[1625]), .B(n3009), .Z(n3011) );
  NANDN U3614 ( .A(n3004), .B(sreg[1624]), .Z(n3008) );
  OR U3615 ( .A(n3006), .B(n3005), .Z(n3007) );
  AND U3616 ( .A(n3008), .B(n3007), .Z(n3010) );
  XOR U3617 ( .A(n3011), .B(n3010), .Z(c[1625]) );
  NAND U3618 ( .A(b[0]), .B(a[603]), .Z(n3014) );
  XOR U3619 ( .A(sreg[1626]), .B(n3014), .Z(n3016) );
  NANDN U3620 ( .A(n3009), .B(sreg[1625]), .Z(n3013) );
  OR U3621 ( .A(n3011), .B(n3010), .Z(n3012) );
  AND U3622 ( .A(n3013), .B(n3012), .Z(n3015) );
  XOR U3623 ( .A(n3016), .B(n3015), .Z(c[1626]) );
  NAND U3624 ( .A(b[0]), .B(a[604]), .Z(n3019) );
  XOR U3625 ( .A(sreg[1627]), .B(n3019), .Z(n3021) );
  NANDN U3626 ( .A(n3014), .B(sreg[1626]), .Z(n3018) );
  OR U3627 ( .A(n3016), .B(n3015), .Z(n3017) );
  AND U3628 ( .A(n3018), .B(n3017), .Z(n3020) );
  XOR U3629 ( .A(n3021), .B(n3020), .Z(c[1627]) );
  NAND U3630 ( .A(b[0]), .B(a[605]), .Z(n3024) );
  XOR U3631 ( .A(sreg[1628]), .B(n3024), .Z(n3026) );
  NANDN U3632 ( .A(n3019), .B(sreg[1627]), .Z(n3023) );
  OR U3633 ( .A(n3021), .B(n3020), .Z(n3022) );
  AND U3634 ( .A(n3023), .B(n3022), .Z(n3025) );
  XOR U3635 ( .A(n3026), .B(n3025), .Z(c[1628]) );
  NAND U3636 ( .A(b[0]), .B(a[606]), .Z(n3029) );
  XOR U3637 ( .A(sreg[1629]), .B(n3029), .Z(n3031) );
  NANDN U3638 ( .A(n3024), .B(sreg[1628]), .Z(n3028) );
  OR U3639 ( .A(n3026), .B(n3025), .Z(n3027) );
  AND U3640 ( .A(n3028), .B(n3027), .Z(n3030) );
  XOR U3641 ( .A(n3031), .B(n3030), .Z(c[1629]) );
  NAND U3642 ( .A(b[0]), .B(a[607]), .Z(n3034) );
  XOR U3643 ( .A(sreg[1630]), .B(n3034), .Z(n3036) );
  NANDN U3644 ( .A(n3029), .B(sreg[1629]), .Z(n3033) );
  OR U3645 ( .A(n3031), .B(n3030), .Z(n3032) );
  AND U3646 ( .A(n3033), .B(n3032), .Z(n3035) );
  XOR U3647 ( .A(n3036), .B(n3035), .Z(c[1630]) );
  NAND U3648 ( .A(b[0]), .B(a[608]), .Z(n3039) );
  XOR U3649 ( .A(sreg[1631]), .B(n3039), .Z(n3041) );
  NANDN U3650 ( .A(n3034), .B(sreg[1630]), .Z(n3038) );
  OR U3651 ( .A(n3036), .B(n3035), .Z(n3037) );
  AND U3652 ( .A(n3038), .B(n3037), .Z(n3040) );
  XOR U3653 ( .A(n3041), .B(n3040), .Z(c[1631]) );
  NAND U3654 ( .A(b[0]), .B(a[609]), .Z(n3044) );
  XOR U3655 ( .A(sreg[1632]), .B(n3044), .Z(n3046) );
  NANDN U3656 ( .A(n3039), .B(sreg[1631]), .Z(n3043) );
  OR U3657 ( .A(n3041), .B(n3040), .Z(n3042) );
  AND U3658 ( .A(n3043), .B(n3042), .Z(n3045) );
  XOR U3659 ( .A(n3046), .B(n3045), .Z(c[1632]) );
  NAND U3660 ( .A(b[0]), .B(a[610]), .Z(n3049) );
  XOR U3661 ( .A(sreg[1633]), .B(n3049), .Z(n3051) );
  NANDN U3662 ( .A(n3044), .B(sreg[1632]), .Z(n3048) );
  OR U3663 ( .A(n3046), .B(n3045), .Z(n3047) );
  AND U3664 ( .A(n3048), .B(n3047), .Z(n3050) );
  XOR U3665 ( .A(n3051), .B(n3050), .Z(c[1633]) );
  NAND U3666 ( .A(b[0]), .B(a[611]), .Z(n3054) );
  XOR U3667 ( .A(sreg[1634]), .B(n3054), .Z(n3056) );
  NANDN U3668 ( .A(n3049), .B(sreg[1633]), .Z(n3053) );
  OR U3669 ( .A(n3051), .B(n3050), .Z(n3052) );
  AND U3670 ( .A(n3053), .B(n3052), .Z(n3055) );
  XOR U3671 ( .A(n3056), .B(n3055), .Z(c[1634]) );
  NAND U3672 ( .A(b[0]), .B(a[612]), .Z(n3059) );
  XOR U3673 ( .A(sreg[1635]), .B(n3059), .Z(n3061) );
  NANDN U3674 ( .A(n3054), .B(sreg[1634]), .Z(n3058) );
  OR U3675 ( .A(n3056), .B(n3055), .Z(n3057) );
  AND U3676 ( .A(n3058), .B(n3057), .Z(n3060) );
  XOR U3677 ( .A(n3061), .B(n3060), .Z(c[1635]) );
  NAND U3678 ( .A(b[0]), .B(a[613]), .Z(n3064) );
  XOR U3679 ( .A(sreg[1636]), .B(n3064), .Z(n3066) );
  NANDN U3680 ( .A(n3059), .B(sreg[1635]), .Z(n3063) );
  OR U3681 ( .A(n3061), .B(n3060), .Z(n3062) );
  AND U3682 ( .A(n3063), .B(n3062), .Z(n3065) );
  XOR U3683 ( .A(n3066), .B(n3065), .Z(c[1636]) );
  NAND U3684 ( .A(b[0]), .B(a[614]), .Z(n3069) );
  XOR U3685 ( .A(sreg[1637]), .B(n3069), .Z(n3071) );
  NANDN U3686 ( .A(n3064), .B(sreg[1636]), .Z(n3068) );
  OR U3687 ( .A(n3066), .B(n3065), .Z(n3067) );
  AND U3688 ( .A(n3068), .B(n3067), .Z(n3070) );
  XOR U3689 ( .A(n3071), .B(n3070), .Z(c[1637]) );
  NAND U3690 ( .A(b[0]), .B(a[615]), .Z(n3074) );
  XOR U3691 ( .A(sreg[1638]), .B(n3074), .Z(n3076) );
  NANDN U3692 ( .A(n3069), .B(sreg[1637]), .Z(n3073) );
  OR U3693 ( .A(n3071), .B(n3070), .Z(n3072) );
  AND U3694 ( .A(n3073), .B(n3072), .Z(n3075) );
  XOR U3695 ( .A(n3076), .B(n3075), .Z(c[1638]) );
  NAND U3696 ( .A(b[0]), .B(a[616]), .Z(n3079) );
  XOR U3697 ( .A(sreg[1639]), .B(n3079), .Z(n3081) );
  NANDN U3698 ( .A(n3074), .B(sreg[1638]), .Z(n3078) );
  OR U3699 ( .A(n3076), .B(n3075), .Z(n3077) );
  AND U3700 ( .A(n3078), .B(n3077), .Z(n3080) );
  XOR U3701 ( .A(n3081), .B(n3080), .Z(c[1639]) );
  NAND U3702 ( .A(b[0]), .B(a[617]), .Z(n3084) );
  XOR U3703 ( .A(sreg[1640]), .B(n3084), .Z(n3086) );
  NANDN U3704 ( .A(n3079), .B(sreg[1639]), .Z(n3083) );
  OR U3705 ( .A(n3081), .B(n3080), .Z(n3082) );
  AND U3706 ( .A(n3083), .B(n3082), .Z(n3085) );
  XOR U3707 ( .A(n3086), .B(n3085), .Z(c[1640]) );
  NAND U3708 ( .A(b[0]), .B(a[618]), .Z(n3089) );
  XOR U3709 ( .A(sreg[1641]), .B(n3089), .Z(n3091) );
  NANDN U3710 ( .A(n3084), .B(sreg[1640]), .Z(n3088) );
  OR U3711 ( .A(n3086), .B(n3085), .Z(n3087) );
  AND U3712 ( .A(n3088), .B(n3087), .Z(n3090) );
  XOR U3713 ( .A(n3091), .B(n3090), .Z(c[1641]) );
  NAND U3714 ( .A(b[0]), .B(a[619]), .Z(n3094) );
  XOR U3715 ( .A(sreg[1642]), .B(n3094), .Z(n3096) );
  NANDN U3716 ( .A(n3089), .B(sreg[1641]), .Z(n3093) );
  OR U3717 ( .A(n3091), .B(n3090), .Z(n3092) );
  AND U3718 ( .A(n3093), .B(n3092), .Z(n3095) );
  XOR U3719 ( .A(n3096), .B(n3095), .Z(c[1642]) );
  NAND U3720 ( .A(b[0]), .B(a[620]), .Z(n3099) );
  XOR U3721 ( .A(sreg[1643]), .B(n3099), .Z(n3101) );
  NANDN U3722 ( .A(n3094), .B(sreg[1642]), .Z(n3098) );
  OR U3723 ( .A(n3096), .B(n3095), .Z(n3097) );
  AND U3724 ( .A(n3098), .B(n3097), .Z(n3100) );
  XOR U3725 ( .A(n3101), .B(n3100), .Z(c[1643]) );
  NAND U3726 ( .A(b[0]), .B(a[621]), .Z(n3104) );
  XOR U3727 ( .A(sreg[1644]), .B(n3104), .Z(n3106) );
  NANDN U3728 ( .A(n3099), .B(sreg[1643]), .Z(n3103) );
  OR U3729 ( .A(n3101), .B(n3100), .Z(n3102) );
  AND U3730 ( .A(n3103), .B(n3102), .Z(n3105) );
  XOR U3731 ( .A(n3106), .B(n3105), .Z(c[1644]) );
  NAND U3732 ( .A(b[0]), .B(a[622]), .Z(n3109) );
  XOR U3733 ( .A(sreg[1645]), .B(n3109), .Z(n3111) );
  NANDN U3734 ( .A(n3104), .B(sreg[1644]), .Z(n3108) );
  OR U3735 ( .A(n3106), .B(n3105), .Z(n3107) );
  AND U3736 ( .A(n3108), .B(n3107), .Z(n3110) );
  XOR U3737 ( .A(n3111), .B(n3110), .Z(c[1645]) );
  NAND U3738 ( .A(b[0]), .B(a[623]), .Z(n3114) );
  XOR U3739 ( .A(sreg[1646]), .B(n3114), .Z(n3116) );
  NANDN U3740 ( .A(n3109), .B(sreg[1645]), .Z(n3113) );
  OR U3741 ( .A(n3111), .B(n3110), .Z(n3112) );
  AND U3742 ( .A(n3113), .B(n3112), .Z(n3115) );
  XOR U3743 ( .A(n3116), .B(n3115), .Z(c[1646]) );
  NAND U3744 ( .A(b[0]), .B(a[624]), .Z(n3119) );
  XOR U3745 ( .A(sreg[1647]), .B(n3119), .Z(n3121) );
  NANDN U3746 ( .A(n3114), .B(sreg[1646]), .Z(n3118) );
  OR U3747 ( .A(n3116), .B(n3115), .Z(n3117) );
  AND U3748 ( .A(n3118), .B(n3117), .Z(n3120) );
  XOR U3749 ( .A(n3121), .B(n3120), .Z(c[1647]) );
  NAND U3750 ( .A(b[0]), .B(a[625]), .Z(n3124) );
  XOR U3751 ( .A(sreg[1648]), .B(n3124), .Z(n3126) );
  NANDN U3752 ( .A(n3119), .B(sreg[1647]), .Z(n3123) );
  OR U3753 ( .A(n3121), .B(n3120), .Z(n3122) );
  AND U3754 ( .A(n3123), .B(n3122), .Z(n3125) );
  XOR U3755 ( .A(n3126), .B(n3125), .Z(c[1648]) );
  NAND U3756 ( .A(b[0]), .B(a[626]), .Z(n3129) );
  XOR U3757 ( .A(sreg[1649]), .B(n3129), .Z(n3131) );
  NANDN U3758 ( .A(n3124), .B(sreg[1648]), .Z(n3128) );
  OR U3759 ( .A(n3126), .B(n3125), .Z(n3127) );
  AND U3760 ( .A(n3128), .B(n3127), .Z(n3130) );
  XOR U3761 ( .A(n3131), .B(n3130), .Z(c[1649]) );
  NAND U3762 ( .A(b[0]), .B(a[627]), .Z(n3134) );
  XOR U3763 ( .A(sreg[1650]), .B(n3134), .Z(n3136) );
  NANDN U3764 ( .A(n3129), .B(sreg[1649]), .Z(n3133) );
  OR U3765 ( .A(n3131), .B(n3130), .Z(n3132) );
  AND U3766 ( .A(n3133), .B(n3132), .Z(n3135) );
  XOR U3767 ( .A(n3136), .B(n3135), .Z(c[1650]) );
  NAND U3768 ( .A(b[0]), .B(a[628]), .Z(n3139) );
  XOR U3769 ( .A(sreg[1651]), .B(n3139), .Z(n3141) );
  NANDN U3770 ( .A(n3134), .B(sreg[1650]), .Z(n3138) );
  OR U3771 ( .A(n3136), .B(n3135), .Z(n3137) );
  AND U3772 ( .A(n3138), .B(n3137), .Z(n3140) );
  XOR U3773 ( .A(n3141), .B(n3140), .Z(c[1651]) );
  NAND U3774 ( .A(b[0]), .B(a[629]), .Z(n3144) );
  XOR U3775 ( .A(sreg[1652]), .B(n3144), .Z(n3146) );
  NANDN U3776 ( .A(n3139), .B(sreg[1651]), .Z(n3143) );
  OR U3777 ( .A(n3141), .B(n3140), .Z(n3142) );
  AND U3778 ( .A(n3143), .B(n3142), .Z(n3145) );
  XOR U3779 ( .A(n3146), .B(n3145), .Z(c[1652]) );
  NAND U3780 ( .A(b[0]), .B(a[630]), .Z(n3149) );
  XOR U3781 ( .A(sreg[1653]), .B(n3149), .Z(n3151) );
  NANDN U3782 ( .A(n3144), .B(sreg[1652]), .Z(n3148) );
  OR U3783 ( .A(n3146), .B(n3145), .Z(n3147) );
  AND U3784 ( .A(n3148), .B(n3147), .Z(n3150) );
  XOR U3785 ( .A(n3151), .B(n3150), .Z(c[1653]) );
  NAND U3786 ( .A(b[0]), .B(a[631]), .Z(n3154) );
  XOR U3787 ( .A(sreg[1654]), .B(n3154), .Z(n3156) );
  NANDN U3788 ( .A(n3149), .B(sreg[1653]), .Z(n3153) );
  OR U3789 ( .A(n3151), .B(n3150), .Z(n3152) );
  AND U3790 ( .A(n3153), .B(n3152), .Z(n3155) );
  XOR U3791 ( .A(n3156), .B(n3155), .Z(c[1654]) );
  NAND U3792 ( .A(b[0]), .B(a[632]), .Z(n3159) );
  XOR U3793 ( .A(sreg[1655]), .B(n3159), .Z(n3161) );
  NANDN U3794 ( .A(n3154), .B(sreg[1654]), .Z(n3158) );
  OR U3795 ( .A(n3156), .B(n3155), .Z(n3157) );
  AND U3796 ( .A(n3158), .B(n3157), .Z(n3160) );
  XOR U3797 ( .A(n3161), .B(n3160), .Z(c[1655]) );
  NAND U3798 ( .A(b[0]), .B(a[633]), .Z(n3164) );
  XOR U3799 ( .A(sreg[1656]), .B(n3164), .Z(n3166) );
  NANDN U3800 ( .A(n3159), .B(sreg[1655]), .Z(n3163) );
  OR U3801 ( .A(n3161), .B(n3160), .Z(n3162) );
  AND U3802 ( .A(n3163), .B(n3162), .Z(n3165) );
  XOR U3803 ( .A(n3166), .B(n3165), .Z(c[1656]) );
  NAND U3804 ( .A(b[0]), .B(a[634]), .Z(n3169) );
  XOR U3805 ( .A(sreg[1657]), .B(n3169), .Z(n3171) );
  NANDN U3806 ( .A(n3164), .B(sreg[1656]), .Z(n3168) );
  OR U3807 ( .A(n3166), .B(n3165), .Z(n3167) );
  AND U3808 ( .A(n3168), .B(n3167), .Z(n3170) );
  XOR U3809 ( .A(n3171), .B(n3170), .Z(c[1657]) );
  NAND U3810 ( .A(b[0]), .B(a[635]), .Z(n3174) );
  XOR U3811 ( .A(sreg[1658]), .B(n3174), .Z(n3176) );
  NANDN U3812 ( .A(n3169), .B(sreg[1657]), .Z(n3173) );
  OR U3813 ( .A(n3171), .B(n3170), .Z(n3172) );
  AND U3814 ( .A(n3173), .B(n3172), .Z(n3175) );
  XOR U3815 ( .A(n3176), .B(n3175), .Z(c[1658]) );
  NAND U3816 ( .A(b[0]), .B(a[636]), .Z(n3179) );
  XOR U3817 ( .A(sreg[1659]), .B(n3179), .Z(n3181) );
  NANDN U3818 ( .A(n3174), .B(sreg[1658]), .Z(n3178) );
  OR U3819 ( .A(n3176), .B(n3175), .Z(n3177) );
  AND U3820 ( .A(n3178), .B(n3177), .Z(n3180) );
  XOR U3821 ( .A(n3181), .B(n3180), .Z(c[1659]) );
  NAND U3822 ( .A(b[0]), .B(a[637]), .Z(n3184) );
  XOR U3823 ( .A(sreg[1660]), .B(n3184), .Z(n3186) );
  NANDN U3824 ( .A(n3179), .B(sreg[1659]), .Z(n3183) );
  OR U3825 ( .A(n3181), .B(n3180), .Z(n3182) );
  AND U3826 ( .A(n3183), .B(n3182), .Z(n3185) );
  XOR U3827 ( .A(n3186), .B(n3185), .Z(c[1660]) );
  NAND U3828 ( .A(b[0]), .B(a[638]), .Z(n3189) );
  XOR U3829 ( .A(sreg[1661]), .B(n3189), .Z(n3191) );
  NANDN U3830 ( .A(n3184), .B(sreg[1660]), .Z(n3188) );
  OR U3831 ( .A(n3186), .B(n3185), .Z(n3187) );
  AND U3832 ( .A(n3188), .B(n3187), .Z(n3190) );
  XOR U3833 ( .A(n3191), .B(n3190), .Z(c[1661]) );
  NAND U3834 ( .A(b[0]), .B(a[639]), .Z(n3194) );
  XOR U3835 ( .A(sreg[1662]), .B(n3194), .Z(n3196) );
  NANDN U3836 ( .A(n3189), .B(sreg[1661]), .Z(n3193) );
  OR U3837 ( .A(n3191), .B(n3190), .Z(n3192) );
  AND U3838 ( .A(n3193), .B(n3192), .Z(n3195) );
  XOR U3839 ( .A(n3196), .B(n3195), .Z(c[1662]) );
  NAND U3840 ( .A(b[0]), .B(a[640]), .Z(n3199) );
  XOR U3841 ( .A(sreg[1663]), .B(n3199), .Z(n3201) );
  NANDN U3842 ( .A(n3194), .B(sreg[1662]), .Z(n3198) );
  OR U3843 ( .A(n3196), .B(n3195), .Z(n3197) );
  AND U3844 ( .A(n3198), .B(n3197), .Z(n3200) );
  XOR U3845 ( .A(n3201), .B(n3200), .Z(c[1663]) );
  NAND U3846 ( .A(b[0]), .B(a[641]), .Z(n3204) );
  XOR U3847 ( .A(sreg[1664]), .B(n3204), .Z(n3206) );
  NANDN U3848 ( .A(n3199), .B(sreg[1663]), .Z(n3203) );
  OR U3849 ( .A(n3201), .B(n3200), .Z(n3202) );
  AND U3850 ( .A(n3203), .B(n3202), .Z(n3205) );
  XOR U3851 ( .A(n3206), .B(n3205), .Z(c[1664]) );
  NAND U3852 ( .A(b[0]), .B(a[642]), .Z(n3209) );
  XOR U3853 ( .A(sreg[1665]), .B(n3209), .Z(n3211) );
  NANDN U3854 ( .A(n3204), .B(sreg[1664]), .Z(n3208) );
  OR U3855 ( .A(n3206), .B(n3205), .Z(n3207) );
  AND U3856 ( .A(n3208), .B(n3207), .Z(n3210) );
  XOR U3857 ( .A(n3211), .B(n3210), .Z(c[1665]) );
  NAND U3858 ( .A(b[0]), .B(a[643]), .Z(n3214) );
  XOR U3859 ( .A(sreg[1666]), .B(n3214), .Z(n3216) );
  NANDN U3860 ( .A(n3209), .B(sreg[1665]), .Z(n3213) );
  OR U3861 ( .A(n3211), .B(n3210), .Z(n3212) );
  AND U3862 ( .A(n3213), .B(n3212), .Z(n3215) );
  XOR U3863 ( .A(n3216), .B(n3215), .Z(c[1666]) );
  NAND U3864 ( .A(b[0]), .B(a[644]), .Z(n3219) );
  XOR U3865 ( .A(sreg[1667]), .B(n3219), .Z(n3221) );
  NANDN U3866 ( .A(n3214), .B(sreg[1666]), .Z(n3218) );
  OR U3867 ( .A(n3216), .B(n3215), .Z(n3217) );
  AND U3868 ( .A(n3218), .B(n3217), .Z(n3220) );
  XOR U3869 ( .A(n3221), .B(n3220), .Z(c[1667]) );
  NAND U3870 ( .A(b[0]), .B(a[645]), .Z(n3224) );
  XOR U3871 ( .A(sreg[1668]), .B(n3224), .Z(n3226) );
  NANDN U3872 ( .A(n3219), .B(sreg[1667]), .Z(n3223) );
  OR U3873 ( .A(n3221), .B(n3220), .Z(n3222) );
  AND U3874 ( .A(n3223), .B(n3222), .Z(n3225) );
  XOR U3875 ( .A(n3226), .B(n3225), .Z(c[1668]) );
  NAND U3876 ( .A(b[0]), .B(a[646]), .Z(n3229) );
  XOR U3877 ( .A(sreg[1669]), .B(n3229), .Z(n3231) );
  NANDN U3878 ( .A(n3224), .B(sreg[1668]), .Z(n3228) );
  OR U3879 ( .A(n3226), .B(n3225), .Z(n3227) );
  AND U3880 ( .A(n3228), .B(n3227), .Z(n3230) );
  XOR U3881 ( .A(n3231), .B(n3230), .Z(c[1669]) );
  NAND U3882 ( .A(b[0]), .B(a[647]), .Z(n3234) );
  XOR U3883 ( .A(sreg[1670]), .B(n3234), .Z(n3236) );
  NANDN U3884 ( .A(n3229), .B(sreg[1669]), .Z(n3233) );
  OR U3885 ( .A(n3231), .B(n3230), .Z(n3232) );
  AND U3886 ( .A(n3233), .B(n3232), .Z(n3235) );
  XOR U3887 ( .A(n3236), .B(n3235), .Z(c[1670]) );
  NAND U3888 ( .A(b[0]), .B(a[648]), .Z(n3239) );
  XOR U3889 ( .A(sreg[1671]), .B(n3239), .Z(n3241) );
  NANDN U3890 ( .A(n3234), .B(sreg[1670]), .Z(n3238) );
  OR U3891 ( .A(n3236), .B(n3235), .Z(n3237) );
  AND U3892 ( .A(n3238), .B(n3237), .Z(n3240) );
  XOR U3893 ( .A(n3241), .B(n3240), .Z(c[1671]) );
  NAND U3894 ( .A(b[0]), .B(a[649]), .Z(n3244) );
  XOR U3895 ( .A(sreg[1672]), .B(n3244), .Z(n3246) );
  NANDN U3896 ( .A(n3239), .B(sreg[1671]), .Z(n3243) );
  OR U3897 ( .A(n3241), .B(n3240), .Z(n3242) );
  AND U3898 ( .A(n3243), .B(n3242), .Z(n3245) );
  XOR U3899 ( .A(n3246), .B(n3245), .Z(c[1672]) );
  NAND U3900 ( .A(b[0]), .B(a[650]), .Z(n3249) );
  XOR U3901 ( .A(sreg[1673]), .B(n3249), .Z(n3251) );
  NANDN U3902 ( .A(n3244), .B(sreg[1672]), .Z(n3248) );
  OR U3903 ( .A(n3246), .B(n3245), .Z(n3247) );
  AND U3904 ( .A(n3248), .B(n3247), .Z(n3250) );
  XOR U3905 ( .A(n3251), .B(n3250), .Z(c[1673]) );
  NAND U3906 ( .A(b[0]), .B(a[651]), .Z(n3254) );
  XOR U3907 ( .A(sreg[1674]), .B(n3254), .Z(n3256) );
  NANDN U3908 ( .A(n3249), .B(sreg[1673]), .Z(n3253) );
  OR U3909 ( .A(n3251), .B(n3250), .Z(n3252) );
  AND U3910 ( .A(n3253), .B(n3252), .Z(n3255) );
  XOR U3911 ( .A(n3256), .B(n3255), .Z(c[1674]) );
  NAND U3912 ( .A(b[0]), .B(a[652]), .Z(n3259) );
  XOR U3913 ( .A(sreg[1675]), .B(n3259), .Z(n3261) );
  NANDN U3914 ( .A(n3254), .B(sreg[1674]), .Z(n3258) );
  OR U3915 ( .A(n3256), .B(n3255), .Z(n3257) );
  AND U3916 ( .A(n3258), .B(n3257), .Z(n3260) );
  XOR U3917 ( .A(n3261), .B(n3260), .Z(c[1675]) );
  NAND U3918 ( .A(b[0]), .B(a[653]), .Z(n3264) );
  XOR U3919 ( .A(sreg[1676]), .B(n3264), .Z(n3266) );
  NANDN U3920 ( .A(n3259), .B(sreg[1675]), .Z(n3263) );
  OR U3921 ( .A(n3261), .B(n3260), .Z(n3262) );
  AND U3922 ( .A(n3263), .B(n3262), .Z(n3265) );
  XOR U3923 ( .A(n3266), .B(n3265), .Z(c[1676]) );
  NAND U3924 ( .A(b[0]), .B(a[654]), .Z(n3269) );
  XOR U3925 ( .A(sreg[1677]), .B(n3269), .Z(n3271) );
  NANDN U3926 ( .A(n3264), .B(sreg[1676]), .Z(n3268) );
  OR U3927 ( .A(n3266), .B(n3265), .Z(n3267) );
  AND U3928 ( .A(n3268), .B(n3267), .Z(n3270) );
  XOR U3929 ( .A(n3271), .B(n3270), .Z(c[1677]) );
  NAND U3930 ( .A(b[0]), .B(a[655]), .Z(n3274) );
  XOR U3931 ( .A(sreg[1678]), .B(n3274), .Z(n3276) );
  NANDN U3932 ( .A(n3269), .B(sreg[1677]), .Z(n3273) );
  OR U3933 ( .A(n3271), .B(n3270), .Z(n3272) );
  AND U3934 ( .A(n3273), .B(n3272), .Z(n3275) );
  XOR U3935 ( .A(n3276), .B(n3275), .Z(c[1678]) );
  NAND U3936 ( .A(b[0]), .B(a[656]), .Z(n3279) );
  XOR U3937 ( .A(sreg[1679]), .B(n3279), .Z(n3281) );
  NANDN U3938 ( .A(n3274), .B(sreg[1678]), .Z(n3278) );
  OR U3939 ( .A(n3276), .B(n3275), .Z(n3277) );
  AND U3940 ( .A(n3278), .B(n3277), .Z(n3280) );
  XOR U3941 ( .A(n3281), .B(n3280), .Z(c[1679]) );
  NAND U3942 ( .A(b[0]), .B(a[657]), .Z(n3284) );
  XOR U3943 ( .A(sreg[1680]), .B(n3284), .Z(n3286) );
  NANDN U3944 ( .A(n3279), .B(sreg[1679]), .Z(n3283) );
  OR U3945 ( .A(n3281), .B(n3280), .Z(n3282) );
  AND U3946 ( .A(n3283), .B(n3282), .Z(n3285) );
  XOR U3947 ( .A(n3286), .B(n3285), .Z(c[1680]) );
  NAND U3948 ( .A(b[0]), .B(a[658]), .Z(n3289) );
  XOR U3949 ( .A(sreg[1681]), .B(n3289), .Z(n3291) );
  NANDN U3950 ( .A(n3284), .B(sreg[1680]), .Z(n3288) );
  OR U3951 ( .A(n3286), .B(n3285), .Z(n3287) );
  AND U3952 ( .A(n3288), .B(n3287), .Z(n3290) );
  XOR U3953 ( .A(n3291), .B(n3290), .Z(c[1681]) );
  NAND U3954 ( .A(b[0]), .B(a[659]), .Z(n3294) );
  XOR U3955 ( .A(sreg[1682]), .B(n3294), .Z(n3296) );
  NANDN U3956 ( .A(n3289), .B(sreg[1681]), .Z(n3293) );
  OR U3957 ( .A(n3291), .B(n3290), .Z(n3292) );
  AND U3958 ( .A(n3293), .B(n3292), .Z(n3295) );
  XOR U3959 ( .A(n3296), .B(n3295), .Z(c[1682]) );
  NAND U3960 ( .A(b[0]), .B(a[660]), .Z(n3299) );
  XOR U3961 ( .A(sreg[1683]), .B(n3299), .Z(n3301) );
  NANDN U3962 ( .A(n3294), .B(sreg[1682]), .Z(n3298) );
  OR U3963 ( .A(n3296), .B(n3295), .Z(n3297) );
  AND U3964 ( .A(n3298), .B(n3297), .Z(n3300) );
  XOR U3965 ( .A(n3301), .B(n3300), .Z(c[1683]) );
  NAND U3966 ( .A(b[0]), .B(a[661]), .Z(n3304) );
  XOR U3967 ( .A(sreg[1684]), .B(n3304), .Z(n3306) );
  NANDN U3968 ( .A(n3299), .B(sreg[1683]), .Z(n3303) );
  OR U3969 ( .A(n3301), .B(n3300), .Z(n3302) );
  AND U3970 ( .A(n3303), .B(n3302), .Z(n3305) );
  XOR U3971 ( .A(n3306), .B(n3305), .Z(c[1684]) );
  NAND U3972 ( .A(b[0]), .B(a[662]), .Z(n3309) );
  XOR U3973 ( .A(sreg[1685]), .B(n3309), .Z(n3311) );
  NANDN U3974 ( .A(n3304), .B(sreg[1684]), .Z(n3308) );
  OR U3975 ( .A(n3306), .B(n3305), .Z(n3307) );
  AND U3976 ( .A(n3308), .B(n3307), .Z(n3310) );
  XOR U3977 ( .A(n3311), .B(n3310), .Z(c[1685]) );
  NAND U3978 ( .A(b[0]), .B(a[663]), .Z(n3314) );
  XOR U3979 ( .A(sreg[1686]), .B(n3314), .Z(n3316) );
  NANDN U3980 ( .A(n3309), .B(sreg[1685]), .Z(n3313) );
  OR U3981 ( .A(n3311), .B(n3310), .Z(n3312) );
  AND U3982 ( .A(n3313), .B(n3312), .Z(n3315) );
  XOR U3983 ( .A(n3316), .B(n3315), .Z(c[1686]) );
  NAND U3984 ( .A(b[0]), .B(a[664]), .Z(n3319) );
  XOR U3985 ( .A(sreg[1687]), .B(n3319), .Z(n3321) );
  NANDN U3986 ( .A(n3314), .B(sreg[1686]), .Z(n3318) );
  OR U3987 ( .A(n3316), .B(n3315), .Z(n3317) );
  AND U3988 ( .A(n3318), .B(n3317), .Z(n3320) );
  XOR U3989 ( .A(n3321), .B(n3320), .Z(c[1687]) );
  NAND U3990 ( .A(b[0]), .B(a[665]), .Z(n3324) );
  XOR U3991 ( .A(sreg[1688]), .B(n3324), .Z(n3326) );
  NANDN U3992 ( .A(n3319), .B(sreg[1687]), .Z(n3323) );
  OR U3993 ( .A(n3321), .B(n3320), .Z(n3322) );
  AND U3994 ( .A(n3323), .B(n3322), .Z(n3325) );
  XOR U3995 ( .A(n3326), .B(n3325), .Z(c[1688]) );
  NAND U3996 ( .A(b[0]), .B(a[666]), .Z(n3329) );
  XOR U3997 ( .A(sreg[1689]), .B(n3329), .Z(n3331) );
  NANDN U3998 ( .A(n3324), .B(sreg[1688]), .Z(n3328) );
  OR U3999 ( .A(n3326), .B(n3325), .Z(n3327) );
  AND U4000 ( .A(n3328), .B(n3327), .Z(n3330) );
  XOR U4001 ( .A(n3331), .B(n3330), .Z(c[1689]) );
  NAND U4002 ( .A(b[0]), .B(a[667]), .Z(n3334) );
  XOR U4003 ( .A(sreg[1690]), .B(n3334), .Z(n3336) );
  NANDN U4004 ( .A(n3329), .B(sreg[1689]), .Z(n3333) );
  OR U4005 ( .A(n3331), .B(n3330), .Z(n3332) );
  AND U4006 ( .A(n3333), .B(n3332), .Z(n3335) );
  XOR U4007 ( .A(n3336), .B(n3335), .Z(c[1690]) );
  NAND U4008 ( .A(b[0]), .B(a[668]), .Z(n3339) );
  XOR U4009 ( .A(sreg[1691]), .B(n3339), .Z(n3341) );
  NANDN U4010 ( .A(n3334), .B(sreg[1690]), .Z(n3338) );
  OR U4011 ( .A(n3336), .B(n3335), .Z(n3337) );
  AND U4012 ( .A(n3338), .B(n3337), .Z(n3340) );
  XOR U4013 ( .A(n3341), .B(n3340), .Z(c[1691]) );
  NAND U4014 ( .A(b[0]), .B(a[669]), .Z(n3344) );
  XOR U4015 ( .A(sreg[1692]), .B(n3344), .Z(n3346) );
  NANDN U4016 ( .A(n3339), .B(sreg[1691]), .Z(n3343) );
  OR U4017 ( .A(n3341), .B(n3340), .Z(n3342) );
  AND U4018 ( .A(n3343), .B(n3342), .Z(n3345) );
  XOR U4019 ( .A(n3346), .B(n3345), .Z(c[1692]) );
  NAND U4020 ( .A(b[0]), .B(a[670]), .Z(n3349) );
  XOR U4021 ( .A(sreg[1693]), .B(n3349), .Z(n3351) );
  NANDN U4022 ( .A(n3344), .B(sreg[1692]), .Z(n3348) );
  OR U4023 ( .A(n3346), .B(n3345), .Z(n3347) );
  AND U4024 ( .A(n3348), .B(n3347), .Z(n3350) );
  XOR U4025 ( .A(n3351), .B(n3350), .Z(c[1693]) );
  NAND U4026 ( .A(b[0]), .B(a[671]), .Z(n3354) );
  XOR U4027 ( .A(sreg[1694]), .B(n3354), .Z(n3356) );
  NANDN U4028 ( .A(n3349), .B(sreg[1693]), .Z(n3353) );
  OR U4029 ( .A(n3351), .B(n3350), .Z(n3352) );
  AND U4030 ( .A(n3353), .B(n3352), .Z(n3355) );
  XOR U4031 ( .A(n3356), .B(n3355), .Z(c[1694]) );
  NAND U4032 ( .A(b[0]), .B(a[672]), .Z(n3359) );
  XOR U4033 ( .A(sreg[1695]), .B(n3359), .Z(n3361) );
  NANDN U4034 ( .A(n3354), .B(sreg[1694]), .Z(n3358) );
  OR U4035 ( .A(n3356), .B(n3355), .Z(n3357) );
  AND U4036 ( .A(n3358), .B(n3357), .Z(n3360) );
  XOR U4037 ( .A(n3361), .B(n3360), .Z(c[1695]) );
  NAND U4038 ( .A(b[0]), .B(a[673]), .Z(n3364) );
  XOR U4039 ( .A(sreg[1696]), .B(n3364), .Z(n3366) );
  NANDN U4040 ( .A(n3359), .B(sreg[1695]), .Z(n3363) );
  OR U4041 ( .A(n3361), .B(n3360), .Z(n3362) );
  AND U4042 ( .A(n3363), .B(n3362), .Z(n3365) );
  XOR U4043 ( .A(n3366), .B(n3365), .Z(c[1696]) );
  NAND U4044 ( .A(b[0]), .B(a[674]), .Z(n3369) );
  XOR U4045 ( .A(sreg[1697]), .B(n3369), .Z(n3371) );
  NANDN U4046 ( .A(n3364), .B(sreg[1696]), .Z(n3368) );
  OR U4047 ( .A(n3366), .B(n3365), .Z(n3367) );
  AND U4048 ( .A(n3368), .B(n3367), .Z(n3370) );
  XOR U4049 ( .A(n3371), .B(n3370), .Z(c[1697]) );
  NAND U4050 ( .A(b[0]), .B(a[675]), .Z(n3374) );
  XOR U4051 ( .A(sreg[1698]), .B(n3374), .Z(n3376) );
  NANDN U4052 ( .A(n3369), .B(sreg[1697]), .Z(n3373) );
  OR U4053 ( .A(n3371), .B(n3370), .Z(n3372) );
  AND U4054 ( .A(n3373), .B(n3372), .Z(n3375) );
  XOR U4055 ( .A(n3376), .B(n3375), .Z(c[1698]) );
  NAND U4056 ( .A(b[0]), .B(a[676]), .Z(n3379) );
  XOR U4057 ( .A(sreg[1699]), .B(n3379), .Z(n3381) );
  NANDN U4058 ( .A(n3374), .B(sreg[1698]), .Z(n3378) );
  OR U4059 ( .A(n3376), .B(n3375), .Z(n3377) );
  AND U4060 ( .A(n3378), .B(n3377), .Z(n3380) );
  XOR U4061 ( .A(n3381), .B(n3380), .Z(c[1699]) );
  NAND U4062 ( .A(b[0]), .B(a[677]), .Z(n3384) );
  XOR U4063 ( .A(sreg[1700]), .B(n3384), .Z(n3386) );
  NANDN U4064 ( .A(n3379), .B(sreg[1699]), .Z(n3383) );
  OR U4065 ( .A(n3381), .B(n3380), .Z(n3382) );
  AND U4066 ( .A(n3383), .B(n3382), .Z(n3385) );
  XOR U4067 ( .A(n3386), .B(n3385), .Z(c[1700]) );
  NAND U4068 ( .A(b[0]), .B(a[678]), .Z(n3389) );
  XOR U4069 ( .A(sreg[1701]), .B(n3389), .Z(n3391) );
  NANDN U4070 ( .A(n3384), .B(sreg[1700]), .Z(n3388) );
  OR U4071 ( .A(n3386), .B(n3385), .Z(n3387) );
  AND U4072 ( .A(n3388), .B(n3387), .Z(n3390) );
  XOR U4073 ( .A(n3391), .B(n3390), .Z(c[1701]) );
  NAND U4074 ( .A(b[0]), .B(a[679]), .Z(n3394) );
  XOR U4075 ( .A(sreg[1702]), .B(n3394), .Z(n3396) );
  NANDN U4076 ( .A(n3389), .B(sreg[1701]), .Z(n3393) );
  OR U4077 ( .A(n3391), .B(n3390), .Z(n3392) );
  AND U4078 ( .A(n3393), .B(n3392), .Z(n3395) );
  XOR U4079 ( .A(n3396), .B(n3395), .Z(c[1702]) );
  NAND U4080 ( .A(b[0]), .B(a[680]), .Z(n3399) );
  XOR U4081 ( .A(sreg[1703]), .B(n3399), .Z(n3401) );
  NANDN U4082 ( .A(n3394), .B(sreg[1702]), .Z(n3398) );
  OR U4083 ( .A(n3396), .B(n3395), .Z(n3397) );
  AND U4084 ( .A(n3398), .B(n3397), .Z(n3400) );
  XOR U4085 ( .A(n3401), .B(n3400), .Z(c[1703]) );
  NAND U4086 ( .A(b[0]), .B(a[681]), .Z(n3404) );
  XOR U4087 ( .A(sreg[1704]), .B(n3404), .Z(n3406) );
  NANDN U4088 ( .A(n3399), .B(sreg[1703]), .Z(n3403) );
  OR U4089 ( .A(n3401), .B(n3400), .Z(n3402) );
  AND U4090 ( .A(n3403), .B(n3402), .Z(n3405) );
  XOR U4091 ( .A(n3406), .B(n3405), .Z(c[1704]) );
  NAND U4092 ( .A(b[0]), .B(a[682]), .Z(n3409) );
  XOR U4093 ( .A(sreg[1705]), .B(n3409), .Z(n3411) );
  NANDN U4094 ( .A(n3404), .B(sreg[1704]), .Z(n3408) );
  OR U4095 ( .A(n3406), .B(n3405), .Z(n3407) );
  AND U4096 ( .A(n3408), .B(n3407), .Z(n3410) );
  XOR U4097 ( .A(n3411), .B(n3410), .Z(c[1705]) );
  NAND U4098 ( .A(b[0]), .B(a[683]), .Z(n3414) );
  XOR U4099 ( .A(sreg[1706]), .B(n3414), .Z(n3416) );
  NANDN U4100 ( .A(n3409), .B(sreg[1705]), .Z(n3413) );
  OR U4101 ( .A(n3411), .B(n3410), .Z(n3412) );
  AND U4102 ( .A(n3413), .B(n3412), .Z(n3415) );
  XOR U4103 ( .A(n3416), .B(n3415), .Z(c[1706]) );
  NAND U4104 ( .A(b[0]), .B(a[684]), .Z(n3419) );
  XOR U4105 ( .A(sreg[1707]), .B(n3419), .Z(n3421) );
  NANDN U4106 ( .A(n3414), .B(sreg[1706]), .Z(n3418) );
  OR U4107 ( .A(n3416), .B(n3415), .Z(n3417) );
  AND U4108 ( .A(n3418), .B(n3417), .Z(n3420) );
  XOR U4109 ( .A(n3421), .B(n3420), .Z(c[1707]) );
  NAND U4110 ( .A(b[0]), .B(a[685]), .Z(n3424) );
  XOR U4111 ( .A(sreg[1708]), .B(n3424), .Z(n3426) );
  NANDN U4112 ( .A(n3419), .B(sreg[1707]), .Z(n3423) );
  OR U4113 ( .A(n3421), .B(n3420), .Z(n3422) );
  AND U4114 ( .A(n3423), .B(n3422), .Z(n3425) );
  XOR U4115 ( .A(n3426), .B(n3425), .Z(c[1708]) );
  NAND U4116 ( .A(b[0]), .B(a[686]), .Z(n3429) );
  XOR U4117 ( .A(sreg[1709]), .B(n3429), .Z(n3431) );
  NANDN U4118 ( .A(n3424), .B(sreg[1708]), .Z(n3428) );
  OR U4119 ( .A(n3426), .B(n3425), .Z(n3427) );
  AND U4120 ( .A(n3428), .B(n3427), .Z(n3430) );
  XOR U4121 ( .A(n3431), .B(n3430), .Z(c[1709]) );
  NAND U4122 ( .A(b[0]), .B(a[687]), .Z(n3434) );
  XOR U4123 ( .A(sreg[1710]), .B(n3434), .Z(n3436) );
  NANDN U4124 ( .A(n3429), .B(sreg[1709]), .Z(n3433) );
  OR U4125 ( .A(n3431), .B(n3430), .Z(n3432) );
  AND U4126 ( .A(n3433), .B(n3432), .Z(n3435) );
  XOR U4127 ( .A(n3436), .B(n3435), .Z(c[1710]) );
  NAND U4128 ( .A(b[0]), .B(a[688]), .Z(n3439) );
  XOR U4129 ( .A(sreg[1711]), .B(n3439), .Z(n3441) );
  NANDN U4130 ( .A(n3434), .B(sreg[1710]), .Z(n3438) );
  OR U4131 ( .A(n3436), .B(n3435), .Z(n3437) );
  AND U4132 ( .A(n3438), .B(n3437), .Z(n3440) );
  XOR U4133 ( .A(n3441), .B(n3440), .Z(c[1711]) );
  NAND U4134 ( .A(b[0]), .B(a[689]), .Z(n3444) );
  XOR U4135 ( .A(sreg[1712]), .B(n3444), .Z(n3446) );
  NANDN U4136 ( .A(n3439), .B(sreg[1711]), .Z(n3443) );
  OR U4137 ( .A(n3441), .B(n3440), .Z(n3442) );
  AND U4138 ( .A(n3443), .B(n3442), .Z(n3445) );
  XOR U4139 ( .A(n3446), .B(n3445), .Z(c[1712]) );
  NAND U4140 ( .A(b[0]), .B(a[690]), .Z(n3449) );
  XOR U4141 ( .A(sreg[1713]), .B(n3449), .Z(n3451) );
  NANDN U4142 ( .A(n3444), .B(sreg[1712]), .Z(n3448) );
  OR U4143 ( .A(n3446), .B(n3445), .Z(n3447) );
  AND U4144 ( .A(n3448), .B(n3447), .Z(n3450) );
  XOR U4145 ( .A(n3451), .B(n3450), .Z(c[1713]) );
  NAND U4146 ( .A(b[0]), .B(a[691]), .Z(n3454) );
  XOR U4147 ( .A(sreg[1714]), .B(n3454), .Z(n3456) );
  NANDN U4148 ( .A(n3449), .B(sreg[1713]), .Z(n3453) );
  OR U4149 ( .A(n3451), .B(n3450), .Z(n3452) );
  AND U4150 ( .A(n3453), .B(n3452), .Z(n3455) );
  XOR U4151 ( .A(n3456), .B(n3455), .Z(c[1714]) );
  NAND U4152 ( .A(b[0]), .B(a[692]), .Z(n3459) );
  XOR U4153 ( .A(sreg[1715]), .B(n3459), .Z(n3461) );
  NANDN U4154 ( .A(n3454), .B(sreg[1714]), .Z(n3458) );
  OR U4155 ( .A(n3456), .B(n3455), .Z(n3457) );
  AND U4156 ( .A(n3458), .B(n3457), .Z(n3460) );
  XOR U4157 ( .A(n3461), .B(n3460), .Z(c[1715]) );
  NAND U4158 ( .A(b[0]), .B(a[693]), .Z(n3464) );
  XOR U4159 ( .A(sreg[1716]), .B(n3464), .Z(n3466) );
  NANDN U4160 ( .A(n3459), .B(sreg[1715]), .Z(n3463) );
  OR U4161 ( .A(n3461), .B(n3460), .Z(n3462) );
  AND U4162 ( .A(n3463), .B(n3462), .Z(n3465) );
  XOR U4163 ( .A(n3466), .B(n3465), .Z(c[1716]) );
  NAND U4164 ( .A(b[0]), .B(a[694]), .Z(n3469) );
  XOR U4165 ( .A(sreg[1717]), .B(n3469), .Z(n3471) );
  NANDN U4166 ( .A(n3464), .B(sreg[1716]), .Z(n3468) );
  OR U4167 ( .A(n3466), .B(n3465), .Z(n3467) );
  AND U4168 ( .A(n3468), .B(n3467), .Z(n3470) );
  XOR U4169 ( .A(n3471), .B(n3470), .Z(c[1717]) );
  NAND U4170 ( .A(b[0]), .B(a[695]), .Z(n3474) );
  XOR U4171 ( .A(sreg[1718]), .B(n3474), .Z(n3476) );
  NANDN U4172 ( .A(n3469), .B(sreg[1717]), .Z(n3473) );
  OR U4173 ( .A(n3471), .B(n3470), .Z(n3472) );
  AND U4174 ( .A(n3473), .B(n3472), .Z(n3475) );
  XOR U4175 ( .A(n3476), .B(n3475), .Z(c[1718]) );
  NAND U4176 ( .A(b[0]), .B(a[696]), .Z(n3479) );
  XOR U4177 ( .A(sreg[1719]), .B(n3479), .Z(n3481) );
  NANDN U4178 ( .A(n3474), .B(sreg[1718]), .Z(n3478) );
  OR U4179 ( .A(n3476), .B(n3475), .Z(n3477) );
  AND U4180 ( .A(n3478), .B(n3477), .Z(n3480) );
  XOR U4181 ( .A(n3481), .B(n3480), .Z(c[1719]) );
  NAND U4182 ( .A(b[0]), .B(a[697]), .Z(n3484) );
  XOR U4183 ( .A(sreg[1720]), .B(n3484), .Z(n3486) );
  NANDN U4184 ( .A(n3479), .B(sreg[1719]), .Z(n3483) );
  OR U4185 ( .A(n3481), .B(n3480), .Z(n3482) );
  AND U4186 ( .A(n3483), .B(n3482), .Z(n3485) );
  XOR U4187 ( .A(n3486), .B(n3485), .Z(c[1720]) );
  NAND U4188 ( .A(b[0]), .B(a[698]), .Z(n3489) );
  XOR U4189 ( .A(sreg[1721]), .B(n3489), .Z(n3491) );
  NANDN U4190 ( .A(n3484), .B(sreg[1720]), .Z(n3488) );
  OR U4191 ( .A(n3486), .B(n3485), .Z(n3487) );
  AND U4192 ( .A(n3488), .B(n3487), .Z(n3490) );
  XOR U4193 ( .A(n3491), .B(n3490), .Z(c[1721]) );
  NAND U4194 ( .A(b[0]), .B(a[699]), .Z(n3494) );
  XOR U4195 ( .A(sreg[1722]), .B(n3494), .Z(n3496) );
  NANDN U4196 ( .A(n3489), .B(sreg[1721]), .Z(n3493) );
  OR U4197 ( .A(n3491), .B(n3490), .Z(n3492) );
  AND U4198 ( .A(n3493), .B(n3492), .Z(n3495) );
  XOR U4199 ( .A(n3496), .B(n3495), .Z(c[1722]) );
  NAND U4200 ( .A(b[0]), .B(a[700]), .Z(n3499) );
  XOR U4201 ( .A(sreg[1723]), .B(n3499), .Z(n3501) );
  NANDN U4202 ( .A(n3494), .B(sreg[1722]), .Z(n3498) );
  OR U4203 ( .A(n3496), .B(n3495), .Z(n3497) );
  AND U4204 ( .A(n3498), .B(n3497), .Z(n3500) );
  XOR U4205 ( .A(n3501), .B(n3500), .Z(c[1723]) );
  NAND U4206 ( .A(b[0]), .B(a[701]), .Z(n3504) );
  XOR U4207 ( .A(sreg[1724]), .B(n3504), .Z(n3506) );
  NANDN U4208 ( .A(n3499), .B(sreg[1723]), .Z(n3503) );
  OR U4209 ( .A(n3501), .B(n3500), .Z(n3502) );
  AND U4210 ( .A(n3503), .B(n3502), .Z(n3505) );
  XOR U4211 ( .A(n3506), .B(n3505), .Z(c[1724]) );
  NAND U4212 ( .A(b[0]), .B(a[702]), .Z(n3509) );
  XOR U4213 ( .A(sreg[1725]), .B(n3509), .Z(n3511) );
  NANDN U4214 ( .A(n3504), .B(sreg[1724]), .Z(n3508) );
  OR U4215 ( .A(n3506), .B(n3505), .Z(n3507) );
  AND U4216 ( .A(n3508), .B(n3507), .Z(n3510) );
  XOR U4217 ( .A(n3511), .B(n3510), .Z(c[1725]) );
  NAND U4218 ( .A(b[0]), .B(a[703]), .Z(n3514) );
  XOR U4219 ( .A(sreg[1726]), .B(n3514), .Z(n3516) );
  NANDN U4220 ( .A(n3509), .B(sreg[1725]), .Z(n3513) );
  OR U4221 ( .A(n3511), .B(n3510), .Z(n3512) );
  AND U4222 ( .A(n3513), .B(n3512), .Z(n3515) );
  XOR U4223 ( .A(n3516), .B(n3515), .Z(c[1726]) );
  NAND U4224 ( .A(b[0]), .B(a[704]), .Z(n3519) );
  XOR U4225 ( .A(sreg[1727]), .B(n3519), .Z(n3521) );
  NANDN U4226 ( .A(n3514), .B(sreg[1726]), .Z(n3518) );
  OR U4227 ( .A(n3516), .B(n3515), .Z(n3517) );
  AND U4228 ( .A(n3518), .B(n3517), .Z(n3520) );
  XOR U4229 ( .A(n3521), .B(n3520), .Z(c[1727]) );
  NAND U4230 ( .A(b[0]), .B(a[705]), .Z(n3524) );
  XOR U4231 ( .A(sreg[1728]), .B(n3524), .Z(n3526) );
  NANDN U4232 ( .A(n3519), .B(sreg[1727]), .Z(n3523) );
  OR U4233 ( .A(n3521), .B(n3520), .Z(n3522) );
  AND U4234 ( .A(n3523), .B(n3522), .Z(n3525) );
  XOR U4235 ( .A(n3526), .B(n3525), .Z(c[1728]) );
  NAND U4236 ( .A(b[0]), .B(a[706]), .Z(n3529) );
  XOR U4237 ( .A(sreg[1729]), .B(n3529), .Z(n3531) );
  NANDN U4238 ( .A(n3524), .B(sreg[1728]), .Z(n3528) );
  OR U4239 ( .A(n3526), .B(n3525), .Z(n3527) );
  AND U4240 ( .A(n3528), .B(n3527), .Z(n3530) );
  XOR U4241 ( .A(n3531), .B(n3530), .Z(c[1729]) );
  NAND U4242 ( .A(b[0]), .B(a[707]), .Z(n3534) );
  XOR U4243 ( .A(sreg[1730]), .B(n3534), .Z(n3536) );
  NANDN U4244 ( .A(n3529), .B(sreg[1729]), .Z(n3533) );
  OR U4245 ( .A(n3531), .B(n3530), .Z(n3532) );
  AND U4246 ( .A(n3533), .B(n3532), .Z(n3535) );
  XOR U4247 ( .A(n3536), .B(n3535), .Z(c[1730]) );
  NAND U4248 ( .A(b[0]), .B(a[708]), .Z(n3539) );
  XOR U4249 ( .A(sreg[1731]), .B(n3539), .Z(n3541) );
  NANDN U4250 ( .A(n3534), .B(sreg[1730]), .Z(n3538) );
  OR U4251 ( .A(n3536), .B(n3535), .Z(n3537) );
  AND U4252 ( .A(n3538), .B(n3537), .Z(n3540) );
  XOR U4253 ( .A(n3541), .B(n3540), .Z(c[1731]) );
  NAND U4254 ( .A(b[0]), .B(a[709]), .Z(n3544) );
  XOR U4255 ( .A(sreg[1732]), .B(n3544), .Z(n3546) );
  NANDN U4256 ( .A(n3539), .B(sreg[1731]), .Z(n3543) );
  OR U4257 ( .A(n3541), .B(n3540), .Z(n3542) );
  AND U4258 ( .A(n3543), .B(n3542), .Z(n3545) );
  XOR U4259 ( .A(n3546), .B(n3545), .Z(c[1732]) );
  NAND U4260 ( .A(b[0]), .B(a[710]), .Z(n3549) );
  XOR U4261 ( .A(sreg[1733]), .B(n3549), .Z(n3551) );
  NANDN U4262 ( .A(n3544), .B(sreg[1732]), .Z(n3548) );
  OR U4263 ( .A(n3546), .B(n3545), .Z(n3547) );
  AND U4264 ( .A(n3548), .B(n3547), .Z(n3550) );
  XOR U4265 ( .A(n3551), .B(n3550), .Z(c[1733]) );
  NAND U4266 ( .A(b[0]), .B(a[711]), .Z(n3554) );
  XOR U4267 ( .A(sreg[1734]), .B(n3554), .Z(n3556) );
  NANDN U4268 ( .A(n3549), .B(sreg[1733]), .Z(n3553) );
  OR U4269 ( .A(n3551), .B(n3550), .Z(n3552) );
  AND U4270 ( .A(n3553), .B(n3552), .Z(n3555) );
  XOR U4271 ( .A(n3556), .B(n3555), .Z(c[1734]) );
  NAND U4272 ( .A(b[0]), .B(a[712]), .Z(n3559) );
  XOR U4273 ( .A(sreg[1735]), .B(n3559), .Z(n3561) );
  NANDN U4274 ( .A(n3554), .B(sreg[1734]), .Z(n3558) );
  OR U4275 ( .A(n3556), .B(n3555), .Z(n3557) );
  AND U4276 ( .A(n3558), .B(n3557), .Z(n3560) );
  XOR U4277 ( .A(n3561), .B(n3560), .Z(c[1735]) );
  NAND U4278 ( .A(b[0]), .B(a[713]), .Z(n3564) );
  XOR U4279 ( .A(sreg[1736]), .B(n3564), .Z(n3566) );
  NANDN U4280 ( .A(n3559), .B(sreg[1735]), .Z(n3563) );
  OR U4281 ( .A(n3561), .B(n3560), .Z(n3562) );
  AND U4282 ( .A(n3563), .B(n3562), .Z(n3565) );
  XOR U4283 ( .A(n3566), .B(n3565), .Z(c[1736]) );
  NAND U4284 ( .A(b[0]), .B(a[714]), .Z(n3569) );
  XOR U4285 ( .A(sreg[1737]), .B(n3569), .Z(n3571) );
  NANDN U4286 ( .A(n3564), .B(sreg[1736]), .Z(n3568) );
  OR U4287 ( .A(n3566), .B(n3565), .Z(n3567) );
  AND U4288 ( .A(n3568), .B(n3567), .Z(n3570) );
  XOR U4289 ( .A(n3571), .B(n3570), .Z(c[1737]) );
  NAND U4290 ( .A(b[0]), .B(a[715]), .Z(n3574) );
  XOR U4291 ( .A(sreg[1738]), .B(n3574), .Z(n3576) );
  NANDN U4292 ( .A(n3569), .B(sreg[1737]), .Z(n3573) );
  OR U4293 ( .A(n3571), .B(n3570), .Z(n3572) );
  AND U4294 ( .A(n3573), .B(n3572), .Z(n3575) );
  XOR U4295 ( .A(n3576), .B(n3575), .Z(c[1738]) );
  NAND U4296 ( .A(b[0]), .B(a[716]), .Z(n3579) );
  XOR U4297 ( .A(sreg[1739]), .B(n3579), .Z(n3581) );
  NANDN U4298 ( .A(n3574), .B(sreg[1738]), .Z(n3578) );
  OR U4299 ( .A(n3576), .B(n3575), .Z(n3577) );
  AND U4300 ( .A(n3578), .B(n3577), .Z(n3580) );
  XOR U4301 ( .A(n3581), .B(n3580), .Z(c[1739]) );
  NAND U4302 ( .A(b[0]), .B(a[717]), .Z(n3584) );
  XOR U4303 ( .A(sreg[1740]), .B(n3584), .Z(n3586) );
  NANDN U4304 ( .A(n3579), .B(sreg[1739]), .Z(n3583) );
  OR U4305 ( .A(n3581), .B(n3580), .Z(n3582) );
  AND U4306 ( .A(n3583), .B(n3582), .Z(n3585) );
  XOR U4307 ( .A(n3586), .B(n3585), .Z(c[1740]) );
  NAND U4308 ( .A(b[0]), .B(a[718]), .Z(n3589) );
  XOR U4309 ( .A(sreg[1741]), .B(n3589), .Z(n3591) );
  NANDN U4310 ( .A(n3584), .B(sreg[1740]), .Z(n3588) );
  OR U4311 ( .A(n3586), .B(n3585), .Z(n3587) );
  AND U4312 ( .A(n3588), .B(n3587), .Z(n3590) );
  XOR U4313 ( .A(n3591), .B(n3590), .Z(c[1741]) );
  NAND U4314 ( .A(b[0]), .B(a[719]), .Z(n3594) );
  XOR U4315 ( .A(sreg[1742]), .B(n3594), .Z(n3596) );
  NANDN U4316 ( .A(n3589), .B(sreg[1741]), .Z(n3593) );
  OR U4317 ( .A(n3591), .B(n3590), .Z(n3592) );
  AND U4318 ( .A(n3593), .B(n3592), .Z(n3595) );
  XOR U4319 ( .A(n3596), .B(n3595), .Z(c[1742]) );
  NAND U4320 ( .A(b[0]), .B(a[720]), .Z(n3599) );
  XOR U4321 ( .A(sreg[1743]), .B(n3599), .Z(n3601) );
  NANDN U4322 ( .A(n3594), .B(sreg[1742]), .Z(n3598) );
  OR U4323 ( .A(n3596), .B(n3595), .Z(n3597) );
  AND U4324 ( .A(n3598), .B(n3597), .Z(n3600) );
  XOR U4325 ( .A(n3601), .B(n3600), .Z(c[1743]) );
  NAND U4326 ( .A(b[0]), .B(a[721]), .Z(n3604) );
  XOR U4327 ( .A(sreg[1744]), .B(n3604), .Z(n3606) );
  NANDN U4328 ( .A(n3599), .B(sreg[1743]), .Z(n3603) );
  OR U4329 ( .A(n3601), .B(n3600), .Z(n3602) );
  AND U4330 ( .A(n3603), .B(n3602), .Z(n3605) );
  XOR U4331 ( .A(n3606), .B(n3605), .Z(c[1744]) );
  NAND U4332 ( .A(b[0]), .B(a[722]), .Z(n3609) );
  XOR U4333 ( .A(sreg[1745]), .B(n3609), .Z(n3611) );
  NANDN U4334 ( .A(n3604), .B(sreg[1744]), .Z(n3608) );
  OR U4335 ( .A(n3606), .B(n3605), .Z(n3607) );
  AND U4336 ( .A(n3608), .B(n3607), .Z(n3610) );
  XOR U4337 ( .A(n3611), .B(n3610), .Z(c[1745]) );
  NAND U4338 ( .A(b[0]), .B(a[723]), .Z(n3614) );
  XOR U4339 ( .A(sreg[1746]), .B(n3614), .Z(n3616) );
  NANDN U4340 ( .A(n3609), .B(sreg[1745]), .Z(n3613) );
  OR U4341 ( .A(n3611), .B(n3610), .Z(n3612) );
  AND U4342 ( .A(n3613), .B(n3612), .Z(n3615) );
  XOR U4343 ( .A(n3616), .B(n3615), .Z(c[1746]) );
  NAND U4344 ( .A(b[0]), .B(a[724]), .Z(n3619) );
  XOR U4345 ( .A(sreg[1747]), .B(n3619), .Z(n3621) );
  NANDN U4346 ( .A(n3614), .B(sreg[1746]), .Z(n3618) );
  OR U4347 ( .A(n3616), .B(n3615), .Z(n3617) );
  AND U4348 ( .A(n3618), .B(n3617), .Z(n3620) );
  XOR U4349 ( .A(n3621), .B(n3620), .Z(c[1747]) );
  NAND U4350 ( .A(b[0]), .B(a[725]), .Z(n3624) );
  XOR U4351 ( .A(sreg[1748]), .B(n3624), .Z(n3626) );
  NANDN U4352 ( .A(n3619), .B(sreg[1747]), .Z(n3623) );
  OR U4353 ( .A(n3621), .B(n3620), .Z(n3622) );
  AND U4354 ( .A(n3623), .B(n3622), .Z(n3625) );
  XOR U4355 ( .A(n3626), .B(n3625), .Z(c[1748]) );
  NAND U4356 ( .A(b[0]), .B(a[726]), .Z(n3629) );
  XOR U4357 ( .A(sreg[1749]), .B(n3629), .Z(n3631) );
  NANDN U4358 ( .A(n3624), .B(sreg[1748]), .Z(n3628) );
  OR U4359 ( .A(n3626), .B(n3625), .Z(n3627) );
  AND U4360 ( .A(n3628), .B(n3627), .Z(n3630) );
  XOR U4361 ( .A(n3631), .B(n3630), .Z(c[1749]) );
  NAND U4362 ( .A(b[0]), .B(a[727]), .Z(n3634) );
  XOR U4363 ( .A(sreg[1750]), .B(n3634), .Z(n3636) );
  NANDN U4364 ( .A(n3629), .B(sreg[1749]), .Z(n3633) );
  OR U4365 ( .A(n3631), .B(n3630), .Z(n3632) );
  AND U4366 ( .A(n3633), .B(n3632), .Z(n3635) );
  XOR U4367 ( .A(n3636), .B(n3635), .Z(c[1750]) );
  NAND U4368 ( .A(b[0]), .B(a[728]), .Z(n3639) );
  XOR U4369 ( .A(sreg[1751]), .B(n3639), .Z(n3641) );
  NANDN U4370 ( .A(n3634), .B(sreg[1750]), .Z(n3638) );
  OR U4371 ( .A(n3636), .B(n3635), .Z(n3637) );
  AND U4372 ( .A(n3638), .B(n3637), .Z(n3640) );
  XOR U4373 ( .A(n3641), .B(n3640), .Z(c[1751]) );
  NAND U4374 ( .A(b[0]), .B(a[729]), .Z(n3644) );
  XOR U4375 ( .A(sreg[1752]), .B(n3644), .Z(n3646) );
  NANDN U4376 ( .A(n3639), .B(sreg[1751]), .Z(n3643) );
  OR U4377 ( .A(n3641), .B(n3640), .Z(n3642) );
  AND U4378 ( .A(n3643), .B(n3642), .Z(n3645) );
  XOR U4379 ( .A(n3646), .B(n3645), .Z(c[1752]) );
  NAND U4380 ( .A(b[0]), .B(a[730]), .Z(n3649) );
  XOR U4381 ( .A(sreg[1753]), .B(n3649), .Z(n3651) );
  NANDN U4382 ( .A(n3644), .B(sreg[1752]), .Z(n3648) );
  OR U4383 ( .A(n3646), .B(n3645), .Z(n3647) );
  AND U4384 ( .A(n3648), .B(n3647), .Z(n3650) );
  XOR U4385 ( .A(n3651), .B(n3650), .Z(c[1753]) );
  NAND U4386 ( .A(b[0]), .B(a[731]), .Z(n3654) );
  XOR U4387 ( .A(sreg[1754]), .B(n3654), .Z(n3656) );
  NANDN U4388 ( .A(n3649), .B(sreg[1753]), .Z(n3653) );
  OR U4389 ( .A(n3651), .B(n3650), .Z(n3652) );
  AND U4390 ( .A(n3653), .B(n3652), .Z(n3655) );
  XOR U4391 ( .A(n3656), .B(n3655), .Z(c[1754]) );
  NAND U4392 ( .A(b[0]), .B(a[732]), .Z(n3659) );
  XOR U4393 ( .A(sreg[1755]), .B(n3659), .Z(n3661) );
  NANDN U4394 ( .A(n3654), .B(sreg[1754]), .Z(n3658) );
  OR U4395 ( .A(n3656), .B(n3655), .Z(n3657) );
  AND U4396 ( .A(n3658), .B(n3657), .Z(n3660) );
  XOR U4397 ( .A(n3661), .B(n3660), .Z(c[1755]) );
  NAND U4398 ( .A(b[0]), .B(a[733]), .Z(n3664) );
  XOR U4399 ( .A(sreg[1756]), .B(n3664), .Z(n3666) );
  NANDN U4400 ( .A(n3659), .B(sreg[1755]), .Z(n3663) );
  OR U4401 ( .A(n3661), .B(n3660), .Z(n3662) );
  AND U4402 ( .A(n3663), .B(n3662), .Z(n3665) );
  XOR U4403 ( .A(n3666), .B(n3665), .Z(c[1756]) );
  NAND U4404 ( .A(b[0]), .B(a[734]), .Z(n3669) );
  XOR U4405 ( .A(sreg[1757]), .B(n3669), .Z(n3671) );
  NANDN U4406 ( .A(n3664), .B(sreg[1756]), .Z(n3668) );
  OR U4407 ( .A(n3666), .B(n3665), .Z(n3667) );
  AND U4408 ( .A(n3668), .B(n3667), .Z(n3670) );
  XOR U4409 ( .A(n3671), .B(n3670), .Z(c[1757]) );
  NAND U4410 ( .A(b[0]), .B(a[735]), .Z(n3674) );
  XOR U4411 ( .A(sreg[1758]), .B(n3674), .Z(n3676) );
  NANDN U4412 ( .A(n3669), .B(sreg[1757]), .Z(n3673) );
  OR U4413 ( .A(n3671), .B(n3670), .Z(n3672) );
  AND U4414 ( .A(n3673), .B(n3672), .Z(n3675) );
  XOR U4415 ( .A(n3676), .B(n3675), .Z(c[1758]) );
  NAND U4416 ( .A(b[0]), .B(a[736]), .Z(n3679) );
  XOR U4417 ( .A(sreg[1759]), .B(n3679), .Z(n3681) );
  NANDN U4418 ( .A(n3674), .B(sreg[1758]), .Z(n3678) );
  OR U4419 ( .A(n3676), .B(n3675), .Z(n3677) );
  AND U4420 ( .A(n3678), .B(n3677), .Z(n3680) );
  XOR U4421 ( .A(n3681), .B(n3680), .Z(c[1759]) );
  NAND U4422 ( .A(b[0]), .B(a[737]), .Z(n3684) );
  XOR U4423 ( .A(sreg[1760]), .B(n3684), .Z(n3686) );
  NANDN U4424 ( .A(n3679), .B(sreg[1759]), .Z(n3683) );
  OR U4425 ( .A(n3681), .B(n3680), .Z(n3682) );
  AND U4426 ( .A(n3683), .B(n3682), .Z(n3685) );
  XOR U4427 ( .A(n3686), .B(n3685), .Z(c[1760]) );
  NAND U4428 ( .A(b[0]), .B(a[738]), .Z(n3689) );
  XOR U4429 ( .A(sreg[1761]), .B(n3689), .Z(n3691) );
  NANDN U4430 ( .A(n3684), .B(sreg[1760]), .Z(n3688) );
  OR U4431 ( .A(n3686), .B(n3685), .Z(n3687) );
  AND U4432 ( .A(n3688), .B(n3687), .Z(n3690) );
  XOR U4433 ( .A(n3691), .B(n3690), .Z(c[1761]) );
  NAND U4434 ( .A(b[0]), .B(a[739]), .Z(n3694) );
  XOR U4435 ( .A(sreg[1762]), .B(n3694), .Z(n3696) );
  NANDN U4436 ( .A(n3689), .B(sreg[1761]), .Z(n3693) );
  OR U4437 ( .A(n3691), .B(n3690), .Z(n3692) );
  AND U4438 ( .A(n3693), .B(n3692), .Z(n3695) );
  XOR U4439 ( .A(n3696), .B(n3695), .Z(c[1762]) );
  NAND U4440 ( .A(b[0]), .B(a[740]), .Z(n3699) );
  XOR U4441 ( .A(sreg[1763]), .B(n3699), .Z(n3701) );
  NANDN U4442 ( .A(n3694), .B(sreg[1762]), .Z(n3698) );
  OR U4443 ( .A(n3696), .B(n3695), .Z(n3697) );
  AND U4444 ( .A(n3698), .B(n3697), .Z(n3700) );
  XOR U4445 ( .A(n3701), .B(n3700), .Z(c[1763]) );
  NAND U4446 ( .A(b[0]), .B(a[741]), .Z(n3704) );
  XOR U4447 ( .A(sreg[1764]), .B(n3704), .Z(n3706) );
  NANDN U4448 ( .A(n3699), .B(sreg[1763]), .Z(n3703) );
  OR U4449 ( .A(n3701), .B(n3700), .Z(n3702) );
  AND U4450 ( .A(n3703), .B(n3702), .Z(n3705) );
  XOR U4451 ( .A(n3706), .B(n3705), .Z(c[1764]) );
  NAND U4452 ( .A(b[0]), .B(a[742]), .Z(n3709) );
  XOR U4453 ( .A(sreg[1765]), .B(n3709), .Z(n3711) );
  NANDN U4454 ( .A(n3704), .B(sreg[1764]), .Z(n3708) );
  OR U4455 ( .A(n3706), .B(n3705), .Z(n3707) );
  AND U4456 ( .A(n3708), .B(n3707), .Z(n3710) );
  XOR U4457 ( .A(n3711), .B(n3710), .Z(c[1765]) );
  NAND U4458 ( .A(b[0]), .B(a[743]), .Z(n3714) );
  XOR U4459 ( .A(sreg[1766]), .B(n3714), .Z(n3716) );
  NANDN U4460 ( .A(n3709), .B(sreg[1765]), .Z(n3713) );
  OR U4461 ( .A(n3711), .B(n3710), .Z(n3712) );
  AND U4462 ( .A(n3713), .B(n3712), .Z(n3715) );
  XOR U4463 ( .A(n3716), .B(n3715), .Z(c[1766]) );
  NAND U4464 ( .A(b[0]), .B(a[744]), .Z(n3719) );
  XOR U4465 ( .A(sreg[1767]), .B(n3719), .Z(n3721) );
  NANDN U4466 ( .A(n3714), .B(sreg[1766]), .Z(n3718) );
  OR U4467 ( .A(n3716), .B(n3715), .Z(n3717) );
  AND U4468 ( .A(n3718), .B(n3717), .Z(n3720) );
  XOR U4469 ( .A(n3721), .B(n3720), .Z(c[1767]) );
  NAND U4470 ( .A(b[0]), .B(a[745]), .Z(n3724) );
  XOR U4471 ( .A(sreg[1768]), .B(n3724), .Z(n3726) );
  NANDN U4472 ( .A(n3719), .B(sreg[1767]), .Z(n3723) );
  OR U4473 ( .A(n3721), .B(n3720), .Z(n3722) );
  AND U4474 ( .A(n3723), .B(n3722), .Z(n3725) );
  XOR U4475 ( .A(n3726), .B(n3725), .Z(c[1768]) );
  NAND U4476 ( .A(b[0]), .B(a[746]), .Z(n3729) );
  XOR U4477 ( .A(sreg[1769]), .B(n3729), .Z(n3731) );
  NANDN U4478 ( .A(n3724), .B(sreg[1768]), .Z(n3728) );
  OR U4479 ( .A(n3726), .B(n3725), .Z(n3727) );
  AND U4480 ( .A(n3728), .B(n3727), .Z(n3730) );
  XOR U4481 ( .A(n3731), .B(n3730), .Z(c[1769]) );
  NAND U4482 ( .A(b[0]), .B(a[747]), .Z(n3734) );
  XOR U4483 ( .A(sreg[1770]), .B(n3734), .Z(n3736) );
  NANDN U4484 ( .A(n3729), .B(sreg[1769]), .Z(n3733) );
  OR U4485 ( .A(n3731), .B(n3730), .Z(n3732) );
  AND U4486 ( .A(n3733), .B(n3732), .Z(n3735) );
  XOR U4487 ( .A(n3736), .B(n3735), .Z(c[1770]) );
  NAND U4488 ( .A(b[0]), .B(a[748]), .Z(n3739) );
  XOR U4489 ( .A(sreg[1771]), .B(n3739), .Z(n3741) );
  NANDN U4490 ( .A(n3734), .B(sreg[1770]), .Z(n3738) );
  OR U4491 ( .A(n3736), .B(n3735), .Z(n3737) );
  AND U4492 ( .A(n3738), .B(n3737), .Z(n3740) );
  XOR U4493 ( .A(n3741), .B(n3740), .Z(c[1771]) );
  NAND U4494 ( .A(b[0]), .B(a[749]), .Z(n3744) );
  XOR U4495 ( .A(sreg[1772]), .B(n3744), .Z(n3746) );
  NANDN U4496 ( .A(n3739), .B(sreg[1771]), .Z(n3743) );
  OR U4497 ( .A(n3741), .B(n3740), .Z(n3742) );
  AND U4498 ( .A(n3743), .B(n3742), .Z(n3745) );
  XOR U4499 ( .A(n3746), .B(n3745), .Z(c[1772]) );
  NAND U4500 ( .A(b[0]), .B(a[750]), .Z(n3749) );
  XOR U4501 ( .A(sreg[1773]), .B(n3749), .Z(n3751) );
  NANDN U4502 ( .A(n3744), .B(sreg[1772]), .Z(n3748) );
  OR U4503 ( .A(n3746), .B(n3745), .Z(n3747) );
  AND U4504 ( .A(n3748), .B(n3747), .Z(n3750) );
  XOR U4505 ( .A(n3751), .B(n3750), .Z(c[1773]) );
  NAND U4506 ( .A(b[0]), .B(a[751]), .Z(n3754) );
  XOR U4507 ( .A(sreg[1774]), .B(n3754), .Z(n3756) );
  NANDN U4508 ( .A(n3749), .B(sreg[1773]), .Z(n3753) );
  OR U4509 ( .A(n3751), .B(n3750), .Z(n3752) );
  AND U4510 ( .A(n3753), .B(n3752), .Z(n3755) );
  XOR U4511 ( .A(n3756), .B(n3755), .Z(c[1774]) );
  NAND U4512 ( .A(b[0]), .B(a[752]), .Z(n3759) );
  XOR U4513 ( .A(sreg[1775]), .B(n3759), .Z(n3761) );
  NANDN U4514 ( .A(n3754), .B(sreg[1774]), .Z(n3758) );
  OR U4515 ( .A(n3756), .B(n3755), .Z(n3757) );
  AND U4516 ( .A(n3758), .B(n3757), .Z(n3760) );
  XOR U4517 ( .A(n3761), .B(n3760), .Z(c[1775]) );
  NAND U4518 ( .A(b[0]), .B(a[753]), .Z(n3764) );
  XOR U4519 ( .A(sreg[1776]), .B(n3764), .Z(n3766) );
  NANDN U4520 ( .A(n3759), .B(sreg[1775]), .Z(n3763) );
  OR U4521 ( .A(n3761), .B(n3760), .Z(n3762) );
  AND U4522 ( .A(n3763), .B(n3762), .Z(n3765) );
  XOR U4523 ( .A(n3766), .B(n3765), .Z(c[1776]) );
  NAND U4524 ( .A(b[0]), .B(a[754]), .Z(n3769) );
  XOR U4525 ( .A(sreg[1777]), .B(n3769), .Z(n3771) );
  NANDN U4526 ( .A(n3764), .B(sreg[1776]), .Z(n3768) );
  OR U4527 ( .A(n3766), .B(n3765), .Z(n3767) );
  AND U4528 ( .A(n3768), .B(n3767), .Z(n3770) );
  XOR U4529 ( .A(n3771), .B(n3770), .Z(c[1777]) );
  NAND U4530 ( .A(b[0]), .B(a[755]), .Z(n3774) );
  XOR U4531 ( .A(sreg[1778]), .B(n3774), .Z(n3776) );
  NANDN U4532 ( .A(n3769), .B(sreg[1777]), .Z(n3773) );
  OR U4533 ( .A(n3771), .B(n3770), .Z(n3772) );
  AND U4534 ( .A(n3773), .B(n3772), .Z(n3775) );
  XOR U4535 ( .A(n3776), .B(n3775), .Z(c[1778]) );
  NAND U4536 ( .A(b[0]), .B(a[756]), .Z(n3779) );
  XOR U4537 ( .A(sreg[1779]), .B(n3779), .Z(n3781) );
  NANDN U4538 ( .A(n3774), .B(sreg[1778]), .Z(n3778) );
  OR U4539 ( .A(n3776), .B(n3775), .Z(n3777) );
  AND U4540 ( .A(n3778), .B(n3777), .Z(n3780) );
  XOR U4541 ( .A(n3781), .B(n3780), .Z(c[1779]) );
  NAND U4542 ( .A(b[0]), .B(a[757]), .Z(n3784) );
  XOR U4543 ( .A(sreg[1780]), .B(n3784), .Z(n3786) );
  NANDN U4544 ( .A(n3779), .B(sreg[1779]), .Z(n3783) );
  OR U4545 ( .A(n3781), .B(n3780), .Z(n3782) );
  AND U4546 ( .A(n3783), .B(n3782), .Z(n3785) );
  XOR U4547 ( .A(n3786), .B(n3785), .Z(c[1780]) );
  NAND U4548 ( .A(b[0]), .B(a[758]), .Z(n3789) );
  XOR U4549 ( .A(sreg[1781]), .B(n3789), .Z(n3791) );
  NANDN U4550 ( .A(n3784), .B(sreg[1780]), .Z(n3788) );
  OR U4551 ( .A(n3786), .B(n3785), .Z(n3787) );
  AND U4552 ( .A(n3788), .B(n3787), .Z(n3790) );
  XOR U4553 ( .A(n3791), .B(n3790), .Z(c[1781]) );
  NAND U4554 ( .A(b[0]), .B(a[759]), .Z(n3794) );
  XOR U4555 ( .A(sreg[1782]), .B(n3794), .Z(n3796) );
  NANDN U4556 ( .A(n3789), .B(sreg[1781]), .Z(n3793) );
  OR U4557 ( .A(n3791), .B(n3790), .Z(n3792) );
  AND U4558 ( .A(n3793), .B(n3792), .Z(n3795) );
  XOR U4559 ( .A(n3796), .B(n3795), .Z(c[1782]) );
  NAND U4560 ( .A(b[0]), .B(a[760]), .Z(n3799) );
  XOR U4561 ( .A(sreg[1783]), .B(n3799), .Z(n3801) );
  NANDN U4562 ( .A(n3794), .B(sreg[1782]), .Z(n3798) );
  OR U4563 ( .A(n3796), .B(n3795), .Z(n3797) );
  AND U4564 ( .A(n3798), .B(n3797), .Z(n3800) );
  XOR U4565 ( .A(n3801), .B(n3800), .Z(c[1783]) );
  NAND U4566 ( .A(b[0]), .B(a[761]), .Z(n3804) );
  XOR U4567 ( .A(sreg[1784]), .B(n3804), .Z(n3806) );
  NANDN U4568 ( .A(n3799), .B(sreg[1783]), .Z(n3803) );
  OR U4569 ( .A(n3801), .B(n3800), .Z(n3802) );
  AND U4570 ( .A(n3803), .B(n3802), .Z(n3805) );
  XOR U4571 ( .A(n3806), .B(n3805), .Z(c[1784]) );
  NAND U4572 ( .A(b[0]), .B(a[762]), .Z(n3809) );
  XOR U4573 ( .A(sreg[1785]), .B(n3809), .Z(n3811) );
  NANDN U4574 ( .A(n3804), .B(sreg[1784]), .Z(n3808) );
  OR U4575 ( .A(n3806), .B(n3805), .Z(n3807) );
  AND U4576 ( .A(n3808), .B(n3807), .Z(n3810) );
  XOR U4577 ( .A(n3811), .B(n3810), .Z(c[1785]) );
  NAND U4578 ( .A(b[0]), .B(a[763]), .Z(n3814) );
  XOR U4579 ( .A(sreg[1786]), .B(n3814), .Z(n3816) );
  NANDN U4580 ( .A(n3809), .B(sreg[1785]), .Z(n3813) );
  OR U4581 ( .A(n3811), .B(n3810), .Z(n3812) );
  AND U4582 ( .A(n3813), .B(n3812), .Z(n3815) );
  XOR U4583 ( .A(n3816), .B(n3815), .Z(c[1786]) );
  NAND U4584 ( .A(b[0]), .B(a[764]), .Z(n3819) );
  XOR U4585 ( .A(sreg[1787]), .B(n3819), .Z(n3821) );
  NANDN U4586 ( .A(n3814), .B(sreg[1786]), .Z(n3818) );
  OR U4587 ( .A(n3816), .B(n3815), .Z(n3817) );
  AND U4588 ( .A(n3818), .B(n3817), .Z(n3820) );
  XOR U4589 ( .A(n3821), .B(n3820), .Z(c[1787]) );
  NAND U4590 ( .A(b[0]), .B(a[765]), .Z(n3824) );
  XOR U4591 ( .A(sreg[1788]), .B(n3824), .Z(n3826) );
  NANDN U4592 ( .A(n3819), .B(sreg[1787]), .Z(n3823) );
  OR U4593 ( .A(n3821), .B(n3820), .Z(n3822) );
  AND U4594 ( .A(n3823), .B(n3822), .Z(n3825) );
  XOR U4595 ( .A(n3826), .B(n3825), .Z(c[1788]) );
  NAND U4596 ( .A(b[0]), .B(a[766]), .Z(n3829) );
  XOR U4597 ( .A(sreg[1789]), .B(n3829), .Z(n3831) );
  NANDN U4598 ( .A(n3824), .B(sreg[1788]), .Z(n3828) );
  OR U4599 ( .A(n3826), .B(n3825), .Z(n3827) );
  AND U4600 ( .A(n3828), .B(n3827), .Z(n3830) );
  XOR U4601 ( .A(n3831), .B(n3830), .Z(c[1789]) );
  NAND U4602 ( .A(b[0]), .B(a[767]), .Z(n3834) );
  XOR U4603 ( .A(sreg[1790]), .B(n3834), .Z(n3836) );
  NANDN U4604 ( .A(n3829), .B(sreg[1789]), .Z(n3833) );
  OR U4605 ( .A(n3831), .B(n3830), .Z(n3832) );
  AND U4606 ( .A(n3833), .B(n3832), .Z(n3835) );
  XOR U4607 ( .A(n3836), .B(n3835), .Z(c[1790]) );
  NAND U4608 ( .A(b[0]), .B(a[768]), .Z(n3839) );
  XOR U4609 ( .A(sreg[1791]), .B(n3839), .Z(n3841) );
  NANDN U4610 ( .A(n3834), .B(sreg[1790]), .Z(n3838) );
  OR U4611 ( .A(n3836), .B(n3835), .Z(n3837) );
  AND U4612 ( .A(n3838), .B(n3837), .Z(n3840) );
  XOR U4613 ( .A(n3841), .B(n3840), .Z(c[1791]) );
  NAND U4614 ( .A(b[0]), .B(a[769]), .Z(n3844) );
  XOR U4615 ( .A(sreg[1792]), .B(n3844), .Z(n3846) );
  NANDN U4616 ( .A(n3839), .B(sreg[1791]), .Z(n3843) );
  OR U4617 ( .A(n3841), .B(n3840), .Z(n3842) );
  AND U4618 ( .A(n3843), .B(n3842), .Z(n3845) );
  XOR U4619 ( .A(n3846), .B(n3845), .Z(c[1792]) );
  NAND U4620 ( .A(b[0]), .B(a[770]), .Z(n3849) );
  XOR U4621 ( .A(sreg[1793]), .B(n3849), .Z(n3851) );
  NANDN U4622 ( .A(n3844), .B(sreg[1792]), .Z(n3848) );
  OR U4623 ( .A(n3846), .B(n3845), .Z(n3847) );
  AND U4624 ( .A(n3848), .B(n3847), .Z(n3850) );
  XOR U4625 ( .A(n3851), .B(n3850), .Z(c[1793]) );
  NAND U4626 ( .A(b[0]), .B(a[771]), .Z(n3854) );
  XOR U4627 ( .A(sreg[1794]), .B(n3854), .Z(n3856) );
  NANDN U4628 ( .A(n3849), .B(sreg[1793]), .Z(n3853) );
  OR U4629 ( .A(n3851), .B(n3850), .Z(n3852) );
  AND U4630 ( .A(n3853), .B(n3852), .Z(n3855) );
  XOR U4631 ( .A(n3856), .B(n3855), .Z(c[1794]) );
  NAND U4632 ( .A(b[0]), .B(a[772]), .Z(n3859) );
  XOR U4633 ( .A(sreg[1795]), .B(n3859), .Z(n3861) );
  NANDN U4634 ( .A(n3854), .B(sreg[1794]), .Z(n3858) );
  OR U4635 ( .A(n3856), .B(n3855), .Z(n3857) );
  AND U4636 ( .A(n3858), .B(n3857), .Z(n3860) );
  XOR U4637 ( .A(n3861), .B(n3860), .Z(c[1795]) );
  NAND U4638 ( .A(b[0]), .B(a[773]), .Z(n3864) );
  XOR U4639 ( .A(sreg[1796]), .B(n3864), .Z(n3866) );
  NANDN U4640 ( .A(n3859), .B(sreg[1795]), .Z(n3863) );
  OR U4641 ( .A(n3861), .B(n3860), .Z(n3862) );
  AND U4642 ( .A(n3863), .B(n3862), .Z(n3865) );
  XOR U4643 ( .A(n3866), .B(n3865), .Z(c[1796]) );
  NAND U4644 ( .A(b[0]), .B(a[774]), .Z(n3869) );
  XOR U4645 ( .A(sreg[1797]), .B(n3869), .Z(n3871) );
  NANDN U4646 ( .A(n3864), .B(sreg[1796]), .Z(n3868) );
  OR U4647 ( .A(n3866), .B(n3865), .Z(n3867) );
  AND U4648 ( .A(n3868), .B(n3867), .Z(n3870) );
  XOR U4649 ( .A(n3871), .B(n3870), .Z(c[1797]) );
  NAND U4650 ( .A(b[0]), .B(a[775]), .Z(n3874) );
  XOR U4651 ( .A(sreg[1798]), .B(n3874), .Z(n3876) );
  NANDN U4652 ( .A(n3869), .B(sreg[1797]), .Z(n3873) );
  OR U4653 ( .A(n3871), .B(n3870), .Z(n3872) );
  AND U4654 ( .A(n3873), .B(n3872), .Z(n3875) );
  XOR U4655 ( .A(n3876), .B(n3875), .Z(c[1798]) );
  NAND U4656 ( .A(b[0]), .B(a[776]), .Z(n3879) );
  XOR U4657 ( .A(sreg[1799]), .B(n3879), .Z(n3881) );
  NANDN U4658 ( .A(n3874), .B(sreg[1798]), .Z(n3878) );
  OR U4659 ( .A(n3876), .B(n3875), .Z(n3877) );
  AND U4660 ( .A(n3878), .B(n3877), .Z(n3880) );
  XOR U4661 ( .A(n3881), .B(n3880), .Z(c[1799]) );
  NAND U4662 ( .A(b[0]), .B(a[777]), .Z(n3884) );
  XOR U4663 ( .A(sreg[1800]), .B(n3884), .Z(n3886) );
  NANDN U4664 ( .A(n3879), .B(sreg[1799]), .Z(n3883) );
  OR U4665 ( .A(n3881), .B(n3880), .Z(n3882) );
  AND U4666 ( .A(n3883), .B(n3882), .Z(n3885) );
  XOR U4667 ( .A(n3886), .B(n3885), .Z(c[1800]) );
  NAND U4668 ( .A(b[0]), .B(a[778]), .Z(n3889) );
  XOR U4669 ( .A(sreg[1801]), .B(n3889), .Z(n3891) );
  NANDN U4670 ( .A(n3884), .B(sreg[1800]), .Z(n3888) );
  OR U4671 ( .A(n3886), .B(n3885), .Z(n3887) );
  AND U4672 ( .A(n3888), .B(n3887), .Z(n3890) );
  XOR U4673 ( .A(n3891), .B(n3890), .Z(c[1801]) );
  NAND U4674 ( .A(b[0]), .B(a[779]), .Z(n3894) );
  XOR U4675 ( .A(sreg[1802]), .B(n3894), .Z(n3896) );
  NANDN U4676 ( .A(n3889), .B(sreg[1801]), .Z(n3893) );
  OR U4677 ( .A(n3891), .B(n3890), .Z(n3892) );
  AND U4678 ( .A(n3893), .B(n3892), .Z(n3895) );
  XOR U4679 ( .A(n3896), .B(n3895), .Z(c[1802]) );
  NAND U4680 ( .A(b[0]), .B(a[780]), .Z(n3899) );
  XOR U4681 ( .A(sreg[1803]), .B(n3899), .Z(n3901) );
  NANDN U4682 ( .A(n3894), .B(sreg[1802]), .Z(n3898) );
  OR U4683 ( .A(n3896), .B(n3895), .Z(n3897) );
  AND U4684 ( .A(n3898), .B(n3897), .Z(n3900) );
  XOR U4685 ( .A(n3901), .B(n3900), .Z(c[1803]) );
  NAND U4686 ( .A(b[0]), .B(a[781]), .Z(n3904) );
  XOR U4687 ( .A(sreg[1804]), .B(n3904), .Z(n3906) );
  NANDN U4688 ( .A(n3899), .B(sreg[1803]), .Z(n3903) );
  OR U4689 ( .A(n3901), .B(n3900), .Z(n3902) );
  AND U4690 ( .A(n3903), .B(n3902), .Z(n3905) );
  XOR U4691 ( .A(n3906), .B(n3905), .Z(c[1804]) );
  NAND U4692 ( .A(b[0]), .B(a[782]), .Z(n3909) );
  XOR U4693 ( .A(sreg[1805]), .B(n3909), .Z(n3911) );
  NANDN U4694 ( .A(n3904), .B(sreg[1804]), .Z(n3908) );
  OR U4695 ( .A(n3906), .B(n3905), .Z(n3907) );
  AND U4696 ( .A(n3908), .B(n3907), .Z(n3910) );
  XOR U4697 ( .A(n3911), .B(n3910), .Z(c[1805]) );
  NAND U4698 ( .A(b[0]), .B(a[783]), .Z(n3914) );
  XOR U4699 ( .A(sreg[1806]), .B(n3914), .Z(n3916) );
  NANDN U4700 ( .A(n3909), .B(sreg[1805]), .Z(n3913) );
  OR U4701 ( .A(n3911), .B(n3910), .Z(n3912) );
  AND U4702 ( .A(n3913), .B(n3912), .Z(n3915) );
  XOR U4703 ( .A(n3916), .B(n3915), .Z(c[1806]) );
  NAND U4704 ( .A(b[0]), .B(a[784]), .Z(n3919) );
  XOR U4705 ( .A(sreg[1807]), .B(n3919), .Z(n3921) );
  NANDN U4706 ( .A(n3914), .B(sreg[1806]), .Z(n3918) );
  OR U4707 ( .A(n3916), .B(n3915), .Z(n3917) );
  AND U4708 ( .A(n3918), .B(n3917), .Z(n3920) );
  XOR U4709 ( .A(n3921), .B(n3920), .Z(c[1807]) );
  NAND U4710 ( .A(b[0]), .B(a[785]), .Z(n3924) );
  XOR U4711 ( .A(sreg[1808]), .B(n3924), .Z(n3926) );
  NANDN U4712 ( .A(n3919), .B(sreg[1807]), .Z(n3923) );
  OR U4713 ( .A(n3921), .B(n3920), .Z(n3922) );
  AND U4714 ( .A(n3923), .B(n3922), .Z(n3925) );
  XOR U4715 ( .A(n3926), .B(n3925), .Z(c[1808]) );
  NAND U4716 ( .A(b[0]), .B(a[786]), .Z(n3929) );
  XOR U4717 ( .A(sreg[1809]), .B(n3929), .Z(n3931) );
  NANDN U4718 ( .A(n3924), .B(sreg[1808]), .Z(n3928) );
  OR U4719 ( .A(n3926), .B(n3925), .Z(n3927) );
  AND U4720 ( .A(n3928), .B(n3927), .Z(n3930) );
  XOR U4721 ( .A(n3931), .B(n3930), .Z(c[1809]) );
  NAND U4722 ( .A(b[0]), .B(a[787]), .Z(n3934) );
  XOR U4723 ( .A(sreg[1810]), .B(n3934), .Z(n3936) );
  NANDN U4724 ( .A(n3929), .B(sreg[1809]), .Z(n3933) );
  OR U4725 ( .A(n3931), .B(n3930), .Z(n3932) );
  AND U4726 ( .A(n3933), .B(n3932), .Z(n3935) );
  XOR U4727 ( .A(n3936), .B(n3935), .Z(c[1810]) );
  NAND U4728 ( .A(b[0]), .B(a[788]), .Z(n3939) );
  XOR U4729 ( .A(sreg[1811]), .B(n3939), .Z(n3941) );
  NANDN U4730 ( .A(n3934), .B(sreg[1810]), .Z(n3938) );
  OR U4731 ( .A(n3936), .B(n3935), .Z(n3937) );
  AND U4732 ( .A(n3938), .B(n3937), .Z(n3940) );
  XOR U4733 ( .A(n3941), .B(n3940), .Z(c[1811]) );
  NAND U4734 ( .A(b[0]), .B(a[789]), .Z(n3944) );
  XOR U4735 ( .A(sreg[1812]), .B(n3944), .Z(n3946) );
  NANDN U4736 ( .A(n3939), .B(sreg[1811]), .Z(n3943) );
  OR U4737 ( .A(n3941), .B(n3940), .Z(n3942) );
  AND U4738 ( .A(n3943), .B(n3942), .Z(n3945) );
  XOR U4739 ( .A(n3946), .B(n3945), .Z(c[1812]) );
  NAND U4740 ( .A(b[0]), .B(a[790]), .Z(n3949) );
  XOR U4741 ( .A(sreg[1813]), .B(n3949), .Z(n3951) );
  NANDN U4742 ( .A(n3944), .B(sreg[1812]), .Z(n3948) );
  OR U4743 ( .A(n3946), .B(n3945), .Z(n3947) );
  AND U4744 ( .A(n3948), .B(n3947), .Z(n3950) );
  XOR U4745 ( .A(n3951), .B(n3950), .Z(c[1813]) );
  NAND U4746 ( .A(b[0]), .B(a[791]), .Z(n3954) );
  XOR U4747 ( .A(sreg[1814]), .B(n3954), .Z(n3956) );
  NANDN U4748 ( .A(n3949), .B(sreg[1813]), .Z(n3953) );
  OR U4749 ( .A(n3951), .B(n3950), .Z(n3952) );
  AND U4750 ( .A(n3953), .B(n3952), .Z(n3955) );
  XOR U4751 ( .A(n3956), .B(n3955), .Z(c[1814]) );
  NAND U4752 ( .A(b[0]), .B(a[792]), .Z(n3959) );
  XOR U4753 ( .A(sreg[1815]), .B(n3959), .Z(n3961) );
  NANDN U4754 ( .A(n3954), .B(sreg[1814]), .Z(n3958) );
  OR U4755 ( .A(n3956), .B(n3955), .Z(n3957) );
  AND U4756 ( .A(n3958), .B(n3957), .Z(n3960) );
  XOR U4757 ( .A(n3961), .B(n3960), .Z(c[1815]) );
  NAND U4758 ( .A(b[0]), .B(a[793]), .Z(n3964) );
  XOR U4759 ( .A(sreg[1816]), .B(n3964), .Z(n3966) );
  NANDN U4760 ( .A(n3959), .B(sreg[1815]), .Z(n3963) );
  OR U4761 ( .A(n3961), .B(n3960), .Z(n3962) );
  AND U4762 ( .A(n3963), .B(n3962), .Z(n3965) );
  XOR U4763 ( .A(n3966), .B(n3965), .Z(c[1816]) );
  NAND U4764 ( .A(b[0]), .B(a[794]), .Z(n3969) );
  XOR U4765 ( .A(sreg[1817]), .B(n3969), .Z(n3971) );
  NANDN U4766 ( .A(n3964), .B(sreg[1816]), .Z(n3968) );
  OR U4767 ( .A(n3966), .B(n3965), .Z(n3967) );
  AND U4768 ( .A(n3968), .B(n3967), .Z(n3970) );
  XOR U4769 ( .A(n3971), .B(n3970), .Z(c[1817]) );
  NAND U4770 ( .A(b[0]), .B(a[795]), .Z(n3974) );
  XOR U4771 ( .A(sreg[1818]), .B(n3974), .Z(n3976) );
  NANDN U4772 ( .A(n3969), .B(sreg[1817]), .Z(n3973) );
  OR U4773 ( .A(n3971), .B(n3970), .Z(n3972) );
  AND U4774 ( .A(n3973), .B(n3972), .Z(n3975) );
  XOR U4775 ( .A(n3976), .B(n3975), .Z(c[1818]) );
  NAND U4776 ( .A(b[0]), .B(a[796]), .Z(n3979) );
  XOR U4777 ( .A(sreg[1819]), .B(n3979), .Z(n3981) );
  NANDN U4778 ( .A(n3974), .B(sreg[1818]), .Z(n3978) );
  OR U4779 ( .A(n3976), .B(n3975), .Z(n3977) );
  AND U4780 ( .A(n3978), .B(n3977), .Z(n3980) );
  XOR U4781 ( .A(n3981), .B(n3980), .Z(c[1819]) );
  NAND U4782 ( .A(b[0]), .B(a[797]), .Z(n3984) );
  XOR U4783 ( .A(sreg[1820]), .B(n3984), .Z(n3986) );
  NANDN U4784 ( .A(n3979), .B(sreg[1819]), .Z(n3983) );
  OR U4785 ( .A(n3981), .B(n3980), .Z(n3982) );
  AND U4786 ( .A(n3983), .B(n3982), .Z(n3985) );
  XOR U4787 ( .A(n3986), .B(n3985), .Z(c[1820]) );
  NAND U4788 ( .A(b[0]), .B(a[798]), .Z(n3989) );
  XOR U4789 ( .A(sreg[1821]), .B(n3989), .Z(n3991) );
  NANDN U4790 ( .A(n3984), .B(sreg[1820]), .Z(n3988) );
  OR U4791 ( .A(n3986), .B(n3985), .Z(n3987) );
  AND U4792 ( .A(n3988), .B(n3987), .Z(n3990) );
  XOR U4793 ( .A(n3991), .B(n3990), .Z(c[1821]) );
  NAND U4794 ( .A(b[0]), .B(a[799]), .Z(n3994) );
  XOR U4795 ( .A(sreg[1822]), .B(n3994), .Z(n3996) );
  NANDN U4796 ( .A(n3989), .B(sreg[1821]), .Z(n3993) );
  OR U4797 ( .A(n3991), .B(n3990), .Z(n3992) );
  AND U4798 ( .A(n3993), .B(n3992), .Z(n3995) );
  XOR U4799 ( .A(n3996), .B(n3995), .Z(c[1822]) );
  NAND U4800 ( .A(b[0]), .B(a[800]), .Z(n3999) );
  XOR U4801 ( .A(sreg[1823]), .B(n3999), .Z(n4001) );
  NANDN U4802 ( .A(n3994), .B(sreg[1822]), .Z(n3998) );
  OR U4803 ( .A(n3996), .B(n3995), .Z(n3997) );
  AND U4804 ( .A(n3998), .B(n3997), .Z(n4000) );
  XOR U4805 ( .A(n4001), .B(n4000), .Z(c[1823]) );
  NAND U4806 ( .A(b[0]), .B(a[801]), .Z(n4004) );
  XOR U4807 ( .A(sreg[1824]), .B(n4004), .Z(n4006) );
  NANDN U4808 ( .A(n3999), .B(sreg[1823]), .Z(n4003) );
  OR U4809 ( .A(n4001), .B(n4000), .Z(n4002) );
  AND U4810 ( .A(n4003), .B(n4002), .Z(n4005) );
  XOR U4811 ( .A(n4006), .B(n4005), .Z(c[1824]) );
  NAND U4812 ( .A(b[0]), .B(a[802]), .Z(n4009) );
  XOR U4813 ( .A(sreg[1825]), .B(n4009), .Z(n4011) );
  NANDN U4814 ( .A(n4004), .B(sreg[1824]), .Z(n4008) );
  OR U4815 ( .A(n4006), .B(n4005), .Z(n4007) );
  AND U4816 ( .A(n4008), .B(n4007), .Z(n4010) );
  XOR U4817 ( .A(n4011), .B(n4010), .Z(c[1825]) );
  NAND U4818 ( .A(b[0]), .B(a[803]), .Z(n4014) );
  XOR U4819 ( .A(sreg[1826]), .B(n4014), .Z(n4016) );
  NANDN U4820 ( .A(n4009), .B(sreg[1825]), .Z(n4013) );
  OR U4821 ( .A(n4011), .B(n4010), .Z(n4012) );
  AND U4822 ( .A(n4013), .B(n4012), .Z(n4015) );
  XOR U4823 ( .A(n4016), .B(n4015), .Z(c[1826]) );
  NAND U4824 ( .A(b[0]), .B(a[804]), .Z(n4019) );
  XOR U4825 ( .A(sreg[1827]), .B(n4019), .Z(n4021) );
  NANDN U4826 ( .A(n4014), .B(sreg[1826]), .Z(n4018) );
  OR U4827 ( .A(n4016), .B(n4015), .Z(n4017) );
  AND U4828 ( .A(n4018), .B(n4017), .Z(n4020) );
  XOR U4829 ( .A(n4021), .B(n4020), .Z(c[1827]) );
  NAND U4830 ( .A(b[0]), .B(a[805]), .Z(n4024) );
  XOR U4831 ( .A(sreg[1828]), .B(n4024), .Z(n4026) );
  NANDN U4832 ( .A(n4019), .B(sreg[1827]), .Z(n4023) );
  OR U4833 ( .A(n4021), .B(n4020), .Z(n4022) );
  AND U4834 ( .A(n4023), .B(n4022), .Z(n4025) );
  XOR U4835 ( .A(n4026), .B(n4025), .Z(c[1828]) );
  NAND U4836 ( .A(b[0]), .B(a[806]), .Z(n4029) );
  XOR U4837 ( .A(sreg[1829]), .B(n4029), .Z(n4031) );
  NANDN U4838 ( .A(n4024), .B(sreg[1828]), .Z(n4028) );
  OR U4839 ( .A(n4026), .B(n4025), .Z(n4027) );
  AND U4840 ( .A(n4028), .B(n4027), .Z(n4030) );
  XOR U4841 ( .A(n4031), .B(n4030), .Z(c[1829]) );
  NAND U4842 ( .A(b[0]), .B(a[807]), .Z(n4034) );
  XOR U4843 ( .A(sreg[1830]), .B(n4034), .Z(n4036) );
  NANDN U4844 ( .A(n4029), .B(sreg[1829]), .Z(n4033) );
  OR U4845 ( .A(n4031), .B(n4030), .Z(n4032) );
  AND U4846 ( .A(n4033), .B(n4032), .Z(n4035) );
  XOR U4847 ( .A(n4036), .B(n4035), .Z(c[1830]) );
  NAND U4848 ( .A(b[0]), .B(a[808]), .Z(n4039) );
  XOR U4849 ( .A(sreg[1831]), .B(n4039), .Z(n4041) );
  NANDN U4850 ( .A(n4034), .B(sreg[1830]), .Z(n4038) );
  OR U4851 ( .A(n4036), .B(n4035), .Z(n4037) );
  AND U4852 ( .A(n4038), .B(n4037), .Z(n4040) );
  XOR U4853 ( .A(n4041), .B(n4040), .Z(c[1831]) );
  NAND U4854 ( .A(b[0]), .B(a[809]), .Z(n4044) );
  XOR U4855 ( .A(sreg[1832]), .B(n4044), .Z(n4046) );
  NANDN U4856 ( .A(n4039), .B(sreg[1831]), .Z(n4043) );
  OR U4857 ( .A(n4041), .B(n4040), .Z(n4042) );
  AND U4858 ( .A(n4043), .B(n4042), .Z(n4045) );
  XOR U4859 ( .A(n4046), .B(n4045), .Z(c[1832]) );
  NAND U4860 ( .A(b[0]), .B(a[810]), .Z(n4049) );
  XOR U4861 ( .A(sreg[1833]), .B(n4049), .Z(n4051) );
  NANDN U4862 ( .A(n4044), .B(sreg[1832]), .Z(n4048) );
  OR U4863 ( .A(n4046), .B(n4045), .Z(n4047) );
  AND U4864 ( .A(n4048), .B(n4047), .Z(n4050) );
  XOR U4865 ( .A(n4051), .B(n4050), .Z(c[1833]) );
  NAND U4866 ( .A(b[0]), .B(a[811]), .Z(n4054) );
  XOR U4867 ( .A(sreg[1834]), .B(n4054), .Z(n4056) );
  NANDN U4868 ( .A(n4049), .B(sreg[1833]), .Z(n4053) );
  OR U4869 ( .A(n4051), .B(n4050), .Z(n4052) );
  AND U4870 ( .A(n4053), .B(n4052), .Z(n4055) );
  XOR U4871 ( .A(n4056), .B(n4055), .Z(c[1834]) );
  NAND U4872 ( .A(b[0]), .B(a[812]), .Z(n4059) );
  XOR U4873 ( .A(sreg[1835]), .B(n4059), .Z(n4061) );
  NANDN U4874 ( .A(n4054), .B(sreg[1834]), .Z(n4058) );
  OR U4875 ( .A(n4056), .B(n4055), .Z(n4057) );
  AND U4876 ( .A(n4058), .B(n4057), .Z(n4060) );
  XOR U4877 ( .A(n4061), .B(n4060), .Z(c[1835]) );
  NAND U4878 ( .A(b[0]), .B(a[813]), .Z(n4064) );
  XOR U4879 ( .A(sreg[1836]), .B(n4064), .Z(n4066) );
  NANDN U4880 ( .A(n4059), .B(sreg[1835]), .Z(n4063) );
  OR U4881 ( .A(n4061), .B(n4060), .Z(n4062) );
  AND U4882 ( .A(n4063), .B(n4062), .Z(n4065) );
  XOR U4883 ( .A(n4066), .B(n4065), .Z(c[1836]) );
  NAND U4884 ( .A(b[0]), .B(a[814]), .Z(n4069) );
  XOR U4885 ( .A(sreg[1837]), .B(n4069), .Z(n4071) );
  NANDN U4886 ( .A(n4064), .B(sreg[1836]), .Z(n4068) );
  OR U4887 ( .A(n4066), .B(n4065), .Z(n4067) );
  AND U4888 ( .A(n4068), .B(n4067), .Z(n4070) );
  XOR U4889 ( .A(n4071), .B(n4070), .Z(c[1837]) );
  NAND U4890 ( .A(b[0]), .B(a[815]), .Z(n4074) );
  XOR U4891 ( .A(sreg[1838]), .B(n4074), .Z(n4076) );
  NANDN U4892 ( .A(n4069), .B(sreg[1837]), .Z(n4073) );
  OR U4893 ( .A(n4071), .B(n4070), .Z(n4072) );
  AND U4894 ( .A(n4073), .B(n4072), .Z(n4075) );
  XOR U4895 ( .A(n4076), .B(n4075), .Z(c[1838]) );
  NAND U4896 ( .A(b[0]), .B(a[816]), .Z(n4079) );
  XOR U4897 ( .A(sreg[1839]), .B(n4079), .Z(n4081) );
  NANDN U4898 ( .A(n4074), .B(sreg[1838]), .Z(n4078) );
  OR U4899 ( .A(n4076), .B(n4075), .Z(n4077) );
  AND U4900 ( .A(n4078), .B(n4077), .Z(n4080) );
  XOR U4901 ( .A(n4081), .B(n4080), .Z(c[1839]) );
  NAND U4902 ( .A(b[0]), .B(a[817]), .Z(n4084) );
  XOR U4903 ( .A(sreg[1840]), .B(n4084), .Z(n4086) );
  NANDN U4904 ( .A(n4079), .B(sreg[1839]), .Z(n4083) );
  OR U4905 ( .A(n4081), .B(n4080), .Z(n4082) );
  AND U4906 ( .A(n4083), .B(n4082), .Z(n4085) );
  XOR U4907 ( .A(n4086), .B(n4085), .Z(c[1840]) );
  NAND U4908 ( .A(b[0]), .B(a[818]), .Z(n4089) );
  XOR U4909 ( .A(sreg[1841]), .B(n4089), .Z(n4091) );
  NANDN U4910 ( .A(n4084), .B(sreg[1840]), .Z(n4088) );
  OR U4911 ( .A(n4086), .B(n4085), .Z(n4087) );
  AND U4912 ( .A(n4088), .B(n4087), .Z(n4090) );
  XOR U4913 ( .A(n4091), .B(n4090), .Z(c[1841]) );
  NAND U4914 ( .A(b[0]), .B(a[819]), .Z(n4094) );
  XOR U4915 ( .A(sreg[1842]), .B(n4094), .Z(n4096) );
  NANDN U4916 ( .A(n4089), .B(sreg[1841]), .Z(n4093) );
  OR U4917 ( .A(n4091), .B(n4090), .Z(n4092) );
  AND U4918 ( .A(n4093), .B(n4092), .Z(n4095) );
  XOR U4919 ( .A(n4096), .B(n4095), .Z(c[1842]) );
  NAND U4920 ( .A(b[0]), .B(a[820]), .Z(n4099) );
  XOR U4921 ( .A(sreg[1843]), .B(n4099), .Z(n4101) );
  NANDN U4922 ( .A(n4094), .B(sreg[1842]), .Z(n4098) );
  OR U4923 ( .A(n4096), .B(n4095), .Z(n4097) );
  AND U4924 ( .A(n4098), .B(n4097), .Z(n4100) );
  XOR U4925 ( .A(n4101), .B(n4100), .Z(c[1843]) );
  NAND U4926 ( .A(b[0]), .B(a[821]), .Z(n4104) );
  XOR U4927 ( .A(sreg[1844]), .B(n4104), .Z(n4106) );
  NANDN U4928 ( .A(n4099), .B(sreg[1843]), .Z(n4103) );
  OR U4929 ( .A(n4101), .B(n4100), .Z(n4102) );
  AND U4930 ( .A(n4103), .B(n4102), .Z(n4105) );
  XOR U4931 ( .A(n4106), .B(n4105), .Z(c[1844]) );
  NAND U4932 ( .A(b[0]), .B(a[822]), .Z(n4109) );
  XOR U4933 ( .A(sreg[1845]), .B(n4109), .Z(n4111) );
  NANDN U4934 ( .A(n4104), .B(sreg[1844]), .Z(n4108) );
  OR U4935 ( .A(n4106), .B(n4105), .Z(n4107) );
  AND U4936 ( .A(n4108), .B(n4107), .Z(n4110) );
  XOR U4937 ( .A(n4111), .B(n4110), .Z(c[1845]) );
  NAND U4938 ( .A(b[0]), .B(a[823]), .Z(n4114) );
  XOR U4939 ( .A(sreg[1846]), .B(n4114), .Z(n4116) );
  NANDN U4940 ( .A(n4109), .B(sreg[1845]), .Z(n4113) );
  OR U4941 ( .A(n4111), .B(n4110), .Z(n4112) );
  AND U4942 ( .A(n4113), .B(n4112), .Z(n4115) );
  XOR U4943 ( .A(n4116), .B(n4115), .Z(c[1846]) );
  NAND U4944 ( .A(b[0]), .B(a[824]), .Z(n4119) );
  XOR U4945 ( .A(sreg[1847]), .B(n4119), .Z(n4121) );
  NANDN U4946 ( .A(n4114), .B(sreg[1846]), .Z(n4118) );
  OR U4947 ( .A(n4116), .B(n4115), .Z(n4117) );
  AND U4948 ( .A(n4118), .B(n4117), .Z(n4120) );
  XOR U4949 ( .A(n4121), .B(n4120), .Z(c[1847]) );
  NAND U4950 ( .A(b[0]), .B(a[825]), .Z(n4124) );
  XOR U4951 ( .A(sreg[1848]), .B(n4124), .Z(n4126) );
  NANDN U4952 ( .A(n4119), .B(sreg[1847]), .Z(n4123) );
  OR U4953 ( .A(n4121), .B(n4120), .Z(n4122) );
  AND U4954 ( .A(n4123), .B(n4122), .Z(n4125) );
  XOR U4955 ( .A(n4126), .B(n4125), .Z(c[1848]) );
  NAND U4956 ( .A(b[0]), .B(a[826]), .Z(n4129) );
  XOR U4957 ( .A(sreg[1849]), .B(n4129), .Z(n4131) );
  NANDN U4958 ( .A(n4124), .B(sreg[1848]), .Z(n4128) );
  OR U4959 ( .A(n4126), .B(n4125), .Z(n4127) );
  AND U4960 ( .A(n4128), .B(n4127), .Z(n4130) );
  XOR U4961 ( .A(n4131), .B(n4130), .Z(c[1849]) );
  NAND U4962 ( .A(b[0]), .B(a[827]), .Z(n4134) );
  XOR U4963 ( .A(sreg[1850]), .B(n4134), .Z(n4136) );
  NANDN U4964 ( .A(n4129), .B(sreg[1849]), .Z(n4133) );
  OR U4965 ( .A(n4131), .B(n4130), .Z(n4132) );
  AND U4966 ( .A(n4133), .B(n4132), .Z(n4135) );
  XOR U4967 ( .A(n4136), .B(n4135), .Z(c[1850]) );
  NAND U4968 ( .A(b[0]), .B(a[828]), .Z(n4139) );
  XOR U4969 ( .A(sreg[1851]), .B(n4139), .Z(n4141) );
  NANDN U4970 ( .A(n4134), .B(sreg[1850]), .Z(n4138) );
  OR U4971 ( .A(n4136), .B(n4135), .Z(n4137) );
  AND U4972 ( .A(n4138), .B(n4137), .Z(n4140) );
  XOR U4973 ( .A(n4141), .B(n4140), .Z(c[1851]) );
  NAND U4974 ( .A(b[0]), .B(a[829]), .Z(n4144) );
  XOR U4975 ( .A(sreg[1852]), .B(n4144), .Z(n4146) );
  NANDN U4976 ( .A(n4139), .B(sreg[1851]), .Z(n4143) );
  OR U4977 ( .A(n4141), .B(n4140), .Z(n4142) );
  AND U4978 ( .A(n4143), .B(n4142), .Z(n4145) );
  XOR U4979 ( .A(n4146), .B(n4145), .Z(c[1852]) );
  NAND U4980 ( .A(b[0]), .B(a[830]), .Z(n4149) );
  XOR U4981 ( .A(sreg[1853]), .B(n4149), .Z(n4151) );
  NANDN U4982 ( .A(n4144), .B(sreg[1852]), .Z(n4148) );
  OR U4983 ( .A(n4146), .B(n4145), .Z(n4147) );
  AND U4984 ( .A(n4148), .B(n4147), .Z(n4150) );
  XOR U4985 ( .A(n4151), .B(n4150), .Z(c[1853]) );
  NAND U4986 ( .A(b[0]), .B(a[831]), .Z(n4154) );
  XOR U4987 ( .A(sreg[1854]), .B(n4154), .Z(n4156) );
  NANDN U4988 ( .A(n4149), .B(sreg[1853]), .Z(n4153) );
  OR U4989 ( .A(n4151), .B(n4150), .Z(n4152) );
  AND U4990 ( .A(n4153), .B(n4152), .Z(n4155) );
  XOR U4991 ( .A(n4156), .B(n4155), .Z(c[1854]) );
  NAND U4992 ( .A(b[0]), .B(a[832]), .Z(n4159) );
  XOR U4993 ( .A(sreg[1855]), .B(n4159), .Z(n4161) );
  NANDN U4994 ( .A(n4154), .B(sreg[1854]), .Z(n4158) );
  OR U4995 ( .A(n4156), .B(n4155), .Z(n4157) );
  AND U4996 ( .A(n4158), .B(n4157), .Z(n4160) );
  XOR U4997 ( .A(n4161), .B(n4160), .Z(c[1855]) );
  NAND U4998 ( .A(b[0]), .B(a[833]), .Z(n4164) );
  XOR U4999 ( .A(sreg[1856]), .B(n4164), .Z(n4166) );
  NANDN U5000 ( .A(n4159), .B(sreg[1855]), .Z(n4163) );
  OR U5001 ( .A(n4161), .B(n4160), .Z(n4162) );
  AND U5002 ( .A(n4163), .B(n4162), .Z(n4165) );
  XOR U5003 ( .A(n4166), .B(n4165), .Z(c[1856]) );
  NAND U5004 ( .A(b[0]), .B(a[834]), .Z(n4169) );
  XOR U5005 ( .A(sreg[1857]), .B(n4169), .Z(n4171) );
  NANDN U5006 ( .A(n4164), .B(sreg[1856]), .Z(n4168) );
  OR U5007 ( .A(n4166), .B(n4165), .Z(n4167) );
  AND U5008 ( .A(n4168), .B(n4167), .Z(n4170) );
  XOR U5009 ( .A(n4171), .B(n4170), .Z(c[1857]) );
  NAND U5010 ( .A(b[0]), .B(a[835]), .Z(n4174) );
  XOR U5011 ( .A(sreg[1858]), .B(n4174), .Z(n4176) );
  NANDN U5012 ( .A(n4169), .B(sreg[1857]), .Z(n4173) );
  OR U5013 ( .A(n4171), .B(n4170), .Z(n4172) );
  AND U5014 ( .A(n4173), .B(n4172), .Z(n4175) );
  XOR U5015 ( .A(n4176), .B(n4175), .Z(c[1858]) );
  NAND U5016 ( .A(b[0]), .B(a[836]), .Z(n4179) );
  XOR U5017 ( .A(sreg[1859]), .B(n4179), .Z(n4181) );
  NANDN U5018 ( .A(n4174), .B(sreg[1858]), .Z(n4178) );
  OR U5019 ( .A(n4176), .B(n4175), .Z(n4177) );
  AND U5020 ( .A(n4178), .B(n4177), .Z(n4180) );
  XOR U5021 ( .A(n4181), .B(n4180), .Z(c[1859]) );
  NAND U5022 ( .A(b[0]), .B(a[837]), .Z(n4184) );
  XOR U5023 ( .A(sreg[1860]), .B(n4184), .Z(n4186) );
  NANDN U5024 ( .A(n4179), .B(sreg[1859]), .Z(n4183) );
  OR U5025 ( .A(n4181), .B(n4180), .Z(n4182) );
  AND U5026 ( .A(n4183), .B(n4182), .Z(n4185) );
  XOR U5027 ( .A(n4186), .B(n4185), .Z(c[1860]) );
  NAND U5028 ( .A(b[0]), .B(a[838]), .Z(n4189) );
  XOR U5029 ( .A(sreg[1861]), .B(n4189), .Z(n4191) );
  NANDN U5030 ( .A(n4184), .B(sreg[1860]), .Z(n4188) );
  OR U5031 ( .A(n4186), .B(n4185), .Z(n4187) );
  AND U5032 ( .A(n4188), .B(n4187), .Z(n4190) );
  XOR U5033 ( .A(n4191), .B(n4190), .Z(c[1861]) );
  NAND U5034 ( .A(b[0]), .B(a[839]), .Z(n4194) );
  XOR U5035 ( .A(sreg[1862]), .B(n4194), .Z(n4196) );
  NANDN U5036 ( .A(n4189), .B(sreg[1861]), .Z(n4193) );
  OR U5037 ( .A(n4191), .B(n4190), .Z(n4192) );
  AND U5038 ( .A(n4193), .B(n4192), .Z(n4195) );
  XOR U5039 ( .A(n4196), .B(n4195), .Z(c[1862]) );
  NAND U5040 ( .A(b[0]), .B(a[840]), .Z(n4199) );
  XOR U5041 ( .A(sreg[1863]), .B(n4199), .Z(n4201) );
  NANDN U5042 ( .A(n4194), .B(sreg[1862]), .Z(n4198) );
  OR U5043 ( .A(n4196), .B(n4195), .Z(n4197) );
  AND U5044 ( .A(n4198), .B(n4197), .Z(n4200) );
  XOR U5045 ( .A(n4201), .B(n4200), .Z(c[1863]) );
  NAND U5046 ( .A(b[0]), .B(a[841]), .Z(n4204) );
  XOR U5047 ( .A(sreg[1864]), .B(n4204), .Z(n4206) );
  NANDN U5048 ( .A(n4199), .B(sreg[1863]), .Z(n4203) );
  OR U5049 ( .A(n4201), .B(n4200), .Z(n4202) );
  AND U5050 ( .A(n4203), .B(n4202), .Z(n4205) );
  XOR U5051 ( .A(n4206), .B(n4205), .Z(c[1864]) );
  NAND U5052 ( .A(b[0]), .B(a[842]), .Z(n4209) );
  XOR U5053 ( .A(sreg[1865]), .B(n4209), .Z(n4211) );
  NANDN U5054 ( .A(n4204), .B(sreg[1864]), .Z(n4208) );
  OR U5055 ( .A(n4206), .B(n4205), .Z(n4207) );
  AND U5056 ( .A(n4208), .B(n4207), .Z(n4210) );
  XOR U5057 ( .A(n4211), .B(n4210), .Z(c[1865]) );
  NAND U5058 ( .A(b[0]), .B(a[843]), .Z(n4214) );
  XOR U5059 ( .A(sreg[1866]), .B(n4214), .Z(n4216) );
  NANDN U5060 ( .A(n4209), .B(sreg[1865]), .Z(n4213) );
  OR U5061 ( .A(n4211), .B(n4210), .Z(n4212) );
  AND U5062 ( .A(n4213), .B(n4212), .Z(n4215) );
  XOR U5063 ( .A(n4216), .B(n4215), .Z(c[1866]) );
  NAND U5064 ( .A(b[0]), .B(a[844]), .Z(n4219) );
  XOR U5065 ( .A(sreg[1867]), .B(n4219), .Z(n4221) );
  NANDN U5066 ( .A(n4214), .B(sreg[1866]), .Z(n4218) );
  OR U5067 ( .A(n4216), .B(n4215), .Z(n4217) );
  AND U5068 ( .A(n4218), .B(n4217), .Z(n4220) );
  XOR U5069 ( .A(n4221), .B(n4220), .Z(c[1867]) );
  NAND U5070 ( .A(b[0]), .B(a[845]), .Z(n4224) );
  XOR U5071 ( .A(sreg[1868]), .B(n4224), .Z(n4226) );
  NANDN U5072 ( .A(n4219), .B(sreg[1867]), .Z(n4223) );
  OR U5073 ( .A(n4221), .B(n4220), .Z(n4222) );
  AND U5074 ( .A(n4223), .B(n4222), .Z(n4225) );
  XOR U5075 ( .A(n4226), .B(n4225), .Z(c[1868]) );
  NAND U5076 ( .A(b[0]), .B(a[846]), .Z(n4229) );
  XOR U5077 ( .A(sreg[1869]), .B(n4229), .Z(n4231) );
  NANDN U5078 ( .A(n4224), .B(sreg[1868]), .Z(n4228) );
  OR U5079 ( .A(n4226), .B(n4225), .Z(n4227) );
  AND U5080 ( .A(n4228), .B(n4227), .Z(n4230) );
  XOR U5081 ( .A(n4231), .B(n4230), .Z(c[1869]) );
  NAND U5082 ( .A(b[0]), .B(a[847]), .Z(n4234) );
  XOR U5083 ( .A(sreg[1870]), .B(n4234), .Z(n4236) );
  NANDN U5084 ( .A(n4229), .B(sreg[1869]), .Z(n4233) );
  OR U5085 ( .A(n4231), .B(n4230), .Z(n4232) );
  AND U5086 ( .A(n4233), .B(n4232), .Z(n4235) );
  XOR U5087 ( .A(n4236), .B(n4235), .Z(c[1870]) );
  NAND U5088 ( .A(b[0]), .B(a[848]), .Z(n4239) );
  XOR U5089 ( .A(sreg[1871]), .B(n4239), .Z(n4241) );
  NANDN U5090 ( .A(n4234), .B(sreg[1870]), .Z(n4238) );
  OR U5091 ( .A(n4236), .B(n4235), .Z(n4237) );
  AND U5092 ( .A(n4238), .B(n4237), .Z(n4240) );
  XOR U5093 ( .A(n4241), .B(n4240), .Z(c[1871]) );
  NAND U5094 ( .A(b[0]), .B(a[849]), .Z(n4244) );
  XOR U5095 ( .A(sreg[1872]), .B(n4244), .Z(n4246) );
  NANDN U5096 ( .A(n4239), .B(sreg[1871]), .Z(n4243) );
  OR U5097 ( .A(n4241), .B(n4240), .Z(n4242) );
  AND U5098 ( .A(n4243), .B(n4242), .Z(n4245) );
  XOR U5099 ( .A(n4246), .B(n4245), .Z(c[1872]) );
  NAND U5100 ( .A(b[0]), .B(a[850]), .Z(n4249) );
  XOR U5101 ( .A(sreg[1873]), .B(n4249), .Z(n4251) );
  NANDN U5102 ( .A(n4244), .B(sreg[1872]), .Z(n4248) );
  OR U5103 ( .A(n4246), .B(n4245), .Z(n4247) );
  AND U5104 ( .A(n4248), .B(n4247), .Z(n4250) );
  XOR U5105 ( .A(n4251), .B(n4250), .Z(c[1873]) );
  NAND U5106 ( .A(b[0]), .B(a[851]), .Z(n4254) );
  XOR U5107 ( .A(sreg[1874]), .B(n4254), .Z(n4256) );
  NANDN U5108 ( .A(n4249), .B(sreg[1873]), .Z(n4253) );
  OR U5109 ( .A(n4251), .B(n4250), .Z(n4252) );
  AND U5110 ( .A(n4253), .B(n4252), .Z(n4255) );
  XOR U5111 ( .A(n4256), .B(n4255), .Z(c[1874]) );
  NAND U5112 ( .A(b[0]), .B(a[852]), .Z(n4259) );
  XOR U5113 ( .A(sreg[1875]), .B(n4259), .Z(n4261) );
  NANDN U5114 ( .A(n4254), .B(sreg[1874]), .Z(n4258) );
  OR U5115 ( .A(n4256), .B(n4255), .Z(n4257) );
  AND U5116 ( .A(n4258), .B(n4257), .Z(n4260) );
  XOR U5117 ( .A(n4261), .B(n4260), .Z(c[1875]) );
  NAND U5118 ( .A(b[0]), .B(a[853]), .Z(n4264) );
  XOR U5119 ( .A(sreg[1876]), .B(n4264), .Z(n4266) );
  NANDN U5120 ( .A(n4259), .B(sreg[1875]), .Z(n4263) );
  OR U5121 ( .A(n4261), .B(n4260), .Z(n4262) );
  AND U5122 ( .A(n4263), .B(n4262), .Z(n4265) );
  XOR U5123 ( .A(n4266), .B(n4265), .Z(c[1876]) );
  NAND U5124 ( .A(b[0]), .B(a[854]), .Z(n4269) );
  XOR U5125 ( .A(sreg[1877]), .B(n4269), .Z(n4271) );
  NANDN U5126 ( .A(n4264), .B(sreg[1876]), .Z(n4268) );
  OR U5127 ( .A(n4266), .B(n4265), .Z(n4267) );
  AND U5128 ( .A(n4268), .B(n4267), .Z(n4270) );
  XOR U5129 ( .A(n4271), .B(n4270), .Z(c[1877]) );
  NAND U5130 ( .A(b[0]), .B(a[855]), .Z(n4274) );
  XOR U5131 ( .A(sreg[1878]), .B(n4274), .Z(n4276) );
  NANDN U5132 ( .A(n4269), .B(sreg[1877]), .Z(n4273) );
  OR U5133 ( .A(n4271), .B(n4270), .Z(n4272) );
  AND U5134 ( .A(n4273), .B(n4272), .Z(n4275) );
  XOR U5135 ( .A(n4276), .B(n4275), .Z(c[1878]) );
  NAND U5136 ( .A(b[0]), .B(a[856]), .Z(n4279) );
  XOR U5137 ( .A(sreg[1879]), .B(n4279), .Z(n4281) );
  NANDN U5138 ( .A(n4274), .B(sreg[1878]), .Z(n4278) );
  OR U5139 ( .A(n4276), .B(n4275), .Z(n4277) );
  AND U5140 ( .A(n4278), .B(n4277), .Z(n4280) );
  XOR U5141 ( .A(n4281), .B(n4280), .Z(c[1879]) );
  NAND U5142 ( .A(b[0]), .B(a[857]), .Z(n4284) );
  XOR U5143 ( .A(sreg[1880]), .B(n4284), .Z(n4286) );
  NANDN U5144 ( .A(n4279), .B(sreg[1879]), .Z(n4283) );
  OR U5145 ( .A(n4281), .B(n4280), .Z(n4282) );
  AND U5146 ( .A(n4283), .B(n4282), .Z(n4285) );
  XOR U5147 ( .A(n4286), .B(n4285), .Z(c[1880]) );
  NAND U5148 ( .A(b[0]), .B(a[858]), .Z(n4289) );
  XOR U5149 ( .A(sreg[1881]), .B(n4289), .Z(n4291) );
  NANDN U5150 ( .A(n4284), .B(sreg[1880]), .Z(n4288) );
  OR U5151 ( .A(n4286), .B(n4285), .Z(n4287) );
  AND U5152 ( .A(n4288), .B(n4287), .Z(n4290) );
  XOR U5153 ( .A(n4291), .B(n4290), .Z(c[1881]) );
  NAND U5154 ( .A(b[0]), .B(a[859]), .Z(n4294) );
  XOR U5155 ( .A(sreg[1882]), .B(n4294), .Z(n4296) );
  NANDN U5156 ( .A(n4289), .B(sreg[1881]), .Z(n4293) );
  OR U5157 ( .A(n4291), .B(n4290), .Z(n4292) );
  AND U5158 ( .A(n4293), .B(n4292), .Z(n4295) );
  XOR U5159 ( .A(n4296), .B(n4295), .Z(c[1882]) );
  NAND U5160 ( .A(b[0]), .B(a[860]), .Z(n4299) );
  XOR U5161 ( .A(sreg[1883]), .B(n4299), .Z(n4301) );
  NANDN U5162 ( .A(n4294), .B(sreg[1882]), .Z(n4298) );
  OR U5163 ( .A(n4296), .B(n4295), .Z(n4297) );
  AND U5164 ( .A(n4298), .B(n4297), .Z(n4300) );
  XOR U5165 ( .A(n4301), .B(n4300), .Z(c[1883]) );
  NAND U5166 ( .A(b[0]), .B(a[861]), .Z(n4304) );
  XOR U5167 ( .A(sreg[1884]), .B(n4304), .Z(n4306) );
  NANDN U5168 ( .A(n4299), .B(sreg[1883]), .Z(n4303) );
  OR U5169 ( .A(n4301), .B(n4300), .Z(n4302) );
  AND U5170 ( .A(n4303), .B(n4302), .Z(n4305) );
  XOR U5171 ( .A(n4306), .B(n4305), .Z(c[1884]) );
  NAND U5172 ( .A(b[0]), .B(a[862]), .Z(n4309) );
  XOR U5173 ( .A(sreg[1885]), .B(n4309), .Z(n4311) );
  NANDN U5174 ( .A(n4304), .B(sreg[1884]), .Z(n4308) );
  OR U5175 ( .A(n4306), .B(n4305), .Z(n4307) );
  AND U5176 ( .A(n4308), .B(n4307), .Z(n4310) );
  XOR U5177 ( .A(n4311), .B(n4310), .Z(c[1885]) );
  NAND U5178 ( .A(b[0]), .B(a[863]), .Z(n4314) );
  XOR U5179 ( .A(sreg[1886]), .B(n4314), .Z(n4316) );
  NANDN U5180 ( .A(n4309), .B(sreg[1885]), .Z(n4313) );
  OR U5181 ( .A(n4311), .B(n4310), .Z(n4312) );
  AND U5182 ( .A(n4313), .B(n4312), .Z(n4315) );
  XOR U5183 ( .A(n4316), .B(n4315), .Z(c[1886]) );
  NAND U5184 ( .A(b[0]), .B(a[864]), .Z(n4319) );
  XOR U5185 ( .A(sreg[1887]), .B(n4319), .Z(n4321) );
  NANDN U5186 ( .A(n4314), .B(sreg[1886]), .Z(n4318) );
  OR U5187 ( .A(n4316), .B(n4315), .Z(n4317) );
  AND U5188 ( .A(n4318), .B(n4317), .Z(n4320) );
  XOR U5189 ( .A(n4321), .B(n4320), .Z(c[1887]) );
  NAND U5190 ( .A(b[0]), .B(a[865]), .Z(n4324) );
  XOR U5191 ( .A(sreg[1888]), .B(n4324), .Z(n4326) );
  NANDN U5192 ( .A(n4319), .B(sreg[1887]), .Z(n4323) );
  OR U5193 ( .A(n4321), .B(n4320), .Z(n4322) );
  AND U5194 ( .A(n4323), .B(n4322), .Z(n4325) );
  XOR U5195 ( .A(n4326), .B(n4325), .Z(c[1888]) );
  NAND U5196 ( .A(b[0]), .B(a[866]), .Z(n4329) );
  XOR U5197 ( .A(sreg[1889]), .B(n4329), .Z(n4331) );
  NANDN U5198 ( .A(n4324), .B(sreg[1888]), .Z(n4328) );
  OR U5199 ( .A(n4326), .B(n4325), .Z(n4327) );
  AND U5200 ( .A(n4328), .B(n4327), .Z(n4330) );
  XOR U5201 ( .A(n4331), .B(n4330), .Z(c[1889]) );
  NAND U5202 ( .A(b[0]), .B(a[867]), .Z(n4334) );
  XOR U5203 ( .A(sreg[1890]), .B(n4334), .Z(n4336) );
  NANDN U5204 ( .A(n4329), .B(sreg[1889]), .Z(n4333) );
  OR U5205 ( .A(n4331), .B(n4330), .Z(n4332) );
  AND U5206 ( .A(n4333), .B(n4332), .Z(n4335) );
  XOR U5207 ( .A(n4336), .B(n4335), .Z(c[1890]) );
  NAND U5208 ( .A(b[0]), .B(a[868]), .Z(n4339) );
  XOR U5209 ( .A(sreg[1891]), .B(n4339), .Z(n4341) );
  NANDN U5210 ( .A(n4334), .B(sreg[1890]), .Z(n4338) );
  OR U5211 ( .A(n4336), .B(n4335), .Z(n4337) );
  AND U5212 ( .A(n4338), .B(n4337), .Z(n4340) );
  XOR U5213 ( .A(n4341), .B(n4340), .Z(c[1891]) );
  NAND U5214 ( .A(b[0]), .B(a[869]), .Z(n4344) );
  XOR U5215 ( .A(sreg[1892]), .B(n4344), .Z(n4346) );
  NANDN U5216 ( .A(n4339), .B(sreg[1891]), .Z(n4343) );
  OR U5217 ( .A(n4341), .B(n4340), .Z(n4342) );
  AND U5218 ( .A(n4343), .B(n4342), .Z(n4345) );
  XOR U5219 ( .A(n4346), .B(n4345), .Z(c[1892]) );
  NAND U5220 ( .A(b[0]), .B(a[870]), .Z(n4349) );
  XOR U5221 ( .A(sreg[1893]), .B(n4349), .Z(n4351) );
  NANDN U5222 ( .A(n4344), .B(sreg[1892]), .Z(n4348) );
  OR U5223 ( .A(n4346), .B(n4345), .Z(n4347) );
  AND U5224 ( .A(n4348), .B(n4347), .Z(n4350) );
  XOR U5225 ( .A(n4351), .B(n4350), .Z(c[1893]) );
  NAND U5226 ( .A(b[0]), .B(a[871]), .Z(n4354) );
  XOR U5227 ( .A(sreg[1894]), .B(n4354), .Z(n4356) );
  NANDN U5228 ( .A(n4349), .B(sreg[1893]), .Z(n4353) );
  OR U5229 ( .A(n4351), .B(n4350), .Z(n4352) );
  AND U5230 ( .A(n4353), .B(n4352), .Z(n4355) );
  XOR U5231 ( .A(n4356), .B(n4355), .Z(c[1894]) );
  NAND U5232 ( .A(b[0]), .B(a[872]), .Z(n4359) );
  XOR U5233 ( .A(sreg[1895]), .B(n4359), .Z(n4361) );
  NANDN U5234 ( .A(n4354), .B(sreg[1894]), .Z(n4358) );
  OR U5235 ( .A(n4356), .B(n4355), .Z(n4357) );
  AND U5236 ( .A(n4358), .B(n4357), .Z(n4360) );
  XOR U5237 ( .A(n4361), .B(n4360), .Z(c[1895]) );
  NAND U5238 ( .A(b[0]), .B(a[873]), .Z(n4364) );
  XOR U5239 ( .A(sreg[1896]), .B(n4364), .Z(n4366) );
  NANDN U5240 ( .A(n4359), .B(sreg[1895]), .Z(n4363) );
  OR U5241 ( .A(n4361), .B(n4360), .Z(n4362) );
  AND U5242 ( .A(n4363), .B(n4362), .Z(n4365) );
  XOR U5243 ( .A(n4366), .B(n4365), .Z(c[1896]) );
  NAND U5244 ( .A(b[0]), .B(a[874]), .Z(n4369) );
  XOR U5245 ( .A(sreg[1897]), .B(n4369), .Z(n4371) );
  NANDN U5246 ( .A(n4364), .B(sreg[1896]), .Z(n4368) );
  OR U5247 ( .A(n4366), .B(n4365), .Z(n4367) );
  AND U5248 ( .A(n4368), .B(n4367), .Z(n4370) );
  XOR U5249 ( .A(n4371), .B(n4370), .Z(c[1897]) );
  NAND U5250 ( .A(b[0]), .B(a[875]), .Z(n4374) );
  XOR U5251 ( .A(sreg[1898]), .B(n4374), .Z(n4376) );
  NANDN U5252 ( .A(n4369), .B(sreg[1897]), .Z(n4373) );
  OR U5253 ( .A(n4371), .B(n4370), .Z(n4372) );
  AND U5254 ( .A(n4373), .B(n4372), .Z(n4375) );
  XOR U5255 ( .A(n4376), .B(n4375), .Z(c[1898]) );
  NAND U5256 ( .A(b[0]), .B(a[876]), .Z(n4379) );
  XOR U5257 ( .A(sreg[1899]), .B(n4379), .Z(n4381) );
  NANDN U5258 ( .A(n4374), .B(sreg[1898]), .Z(n4378) );
  OR U5259 ( .A(n4376), .B(n4375), .Z(n4377) );
  AND U5260 ( .A(n4378), .B(n4377), .Z(n4380) );
  XOR U5261 ( .A(n4381), .B(n4380), .Z(c[1899]) );
  NAND U5262 ( .A(b[0]), .B(a[877]), .Z(n4384) );
  XOR U5263 ( .A(sreg[1900]), .B(n4384), .Z(n4386) );
  NANDN U5264 ( .A(n4379), .B(sreg[1899]), .Z(n4383) );
  OR U5265 ( .A(n4381), .B(n4380), .Z(n4382) );
  AND U5266 ( .A(n4383), .B(n4382), .Z(n4385) );
  XOR U5267 ( .A(n4386), .B(n4385), .Z(c[1900]) );
  NAND U5268 ( .A(b[0]), .B(a[878]), .Z(n4389) );
  XOR U5269 ( .A(sreg[1901]), .B(n4389), .Z(n4391) );
  NANDN U5270 ( .A(n4384), .B(sreg[1900]), .Z(n4388) );
  OR U5271 ( .A(n4386), .B(n4385), .Z(n4387) );
  AND U5272 ( .A(n4388), .B(n4387), .Z(n4390) );
  XOR U5273 ( .A(n4391), .B(n4390), .Z(c[1901]) );
  NAND U5274 ( .A(b[0]), .B(a[879]), .Z(n4394) );
  XOR U5275 ( .A(sreg[1902]), .B(n4394), .Z(n4396) );
  NANDN U5276 ( .A(n4389), .B(sreg[1901]), .Z(n4393) );
  OR U5277 ( .A(n4391), .B(n4390), .Z(n4392) );
  AND U5278 ( .A(n4393), .B(n4392), .Z(n4395) );
  XOR U5279 ( .A(n4396), .B(n4395), .Z(c[1902]) );
  NAND U5280 ( .A(b[0]), .B(a[880]), .Z(n4399) );
  XOR U5281 ( .A(sreg[1903]), .B(n4399), .Z(n4401) );
  NANDN U5282 ( .A(n4394), .B(sreg[1902]), .Z(n4398) );
  OR U5283 ( .A(n4396), .B(n4395), .Z(n4397) );
  AND U5284 ( .A(n4398), .B(n4397), .Z(n4400) );
  XOR U5285 ( .A(n4401), .B(n4400), .Z(c[1903]) );
  NAND U5286 ( .A(b[0]), .B(a[881]), .Z(n4404) );
  XOR U5287 ( .A(sreg[1904]), .B(n4404), .Z(n4406) );
  NANDN U5288 ( .A(n4399), .B(sreg[1903]), .Z(n4403) );
  OR U5289 ( .A(n4401), .B(n4400), .Z(n4402) );
  AND U5290 ( .A(n4403), .B(n4402), .Z(n4405) );
  XOR U5291 ( .A(n4406), .B(n4405), .Z(c[1904]) );
  NAND U5292 ( .A(b[0]), .B(a[882]), .Z(n4409) );
  XOR U5293 ( .A(sreg[1905]), .B(n4409), .Z(n4411) );
  NANDN U5294 ( .A(n4404), .B(sreg[1904]), .Z(n4408) );
  OR U5295 ( .A(n4406), .B(n4405), .Z(n4407) );
  AND U5296 ( .A(n4408), .B(n4407), .Z(n4410) );
  XOR U5297 ( .A(n4411), .B(n4410), .Z(c[1905]) );
  NAND U5298 ( .A(b[0]), .B(a[883]), .Z(n4414) );
  XOR U5299 ( .A(sreg[1906]), .B(n4414), .Z(n4416) );
  NANDN U5300 ( .A(n4409), .B(sreg[1905]), .Z(n4413) );
  OR U5301 ( .A(n4411), .B(n4410), .Z(n4412) );
  AND U5302 ( .A(n4413), .B(n4412), .Z(n4415) );
  XOR U5303 ( .A(n4416), .B(n4415), .Z(c[1906]) );
  NAND U5304 ( .A(b[0]), .B(a[884]), .Z(n4419) );
  XOR U5305 ( .A(sreg[1907]), .B(n4419), .Z(n4421) );
  NANDN U5306 ( .A(n4414), .B(sreg[1906]), .Z(n4418) );
  OR U5307 ( .A(n4416), .B(n4415), .Z(n4417) );
  AND U5308 ( .A(n4418), .B(n4417), .Z(n4420) );
  XOR U5309 ( .A(n4421), .B(n4420), .Z(c[1907]) );
  NAND U5310 ( .A(b[0]), .B(a[885]), .Z(n4424) );
  XOR U5311 ( .A(sreg[1908]), .B(n4424), .Z(n4426) );
  NANDN U5312 ( .A(n4419), .B(sreg[1907]), .Z(n4423) );
  OR U5313 ( .A(n4421), .B(n4420), .Z(n4422) );
  AND U5314 ( .A(n4423), .B(n4422), .Z(n4425) );
  XOR U5315 ( .A(n4426), .B(n4425), .Z(c[1908]) );
  NAND U5316 ( .A(b[0]), .B(a[886]), .Z(n4429) );
  XOR U5317 ( .A(sreg[1909]), .B(n4429), .Z(n4431) );
  NANDN U5318 ( .A(n4424), .B(sreg[1908]), .Z(n4428) );
  OR U5319 ( .A(n4426), .B(n4425), .Z(n4427) );
  AND U5320 ( .A(n4428), .B(n4427), .Z(n4430) );
  XOR U5321 ( .A(n4431), .B(n4430), .Z(c[1909]) );
  NAND U5322 ( .A(b[0]), .B(a[887]), .Z(n4434) );
  XOR U5323 ( .A(sreg[1910]), .B(n4434), .Z(n4436) );
  NANDN U5324 ( .A(n4429), .B(sreg[1909]), .Z(n4433) );
  OR U5325 ( .A(n4431), .B(n4430), .Z(n4432) );
  AND U5326 ( .A(n4433), .B(n4432), .Z(n4435) );
  XOR U5327 ( .A(n4436), .B(n4435), .Z(c[1910]) );
  NAND U5328 ( .A(b[0]), .B(a[888]), .Z(n4439) );
  XOR U5329 ( .A(sreg[1911]), .B(n4439), .Z(n4441) );
  NANDN U5330 ( .A(n4434), .B(sreg[1910]), .Z(n4438) );
  OR U5331 ( .A(n4436), .B(n4435), .Z(n4437) );
  AND U5332 ( .A(n4438), .B(n4437), .Z(n4440) );
  XOR U5333 ( .A(n4441), .B(n4440), .Z(c[1911]) );
  NAND U5334 ( .A(b[0]), .B(a[889]), .Z(n4444) );
  XOR U5335 ( .A(sreg[1912]), .B(n4444), .Z(n4446) );
  NANDN U5336 ( .A(n4439), .B(sreg[1911]), .Z(n4443) );
  OR U5337 ( .A(n4441), .B(n4440), .Z(n4442) );
  AND U5338 ( .A(n4443), .B(n4442), .Z(n4445) );
  XOR U5339 ( .A(n4446), .B(n4445), .Z(c[1912]) );
  NAND U5340 ( .A(b[0]), .B(a[890]), .Z(n4449) );
  XOR U5341 ( .A(sreg[1913]), .B(n4449), .Z(n4451) );
  NANDN U5342 ( .A(n4444), .B(sreg[1912]), .Z(n4448) );
  OR U5343 ( .A(n4446), .B(n4445), .Z(n4447) );
  AND U5344 ( .A(n4448), .B(n4447), .Z(n4450) );
  XOR U5345 ( .A(n4451), .B(n4450), .Z(c[1913]) );
  NAND U5346 ( .A(b[0]), .B(a[891]), .Z(n4454) );
  XOR U5347 ( .A(sreg[1914]), .B(n4454), .Z(n4456) );
  NANDN U5348 ( .A(n4449), .B(sreg[1913]), .Z(n4453) );
  OR U5349 ( .A(n4451), .B(n4450), .Z(n4452) );
  AND U5350 ( .A(n4453), .B(n4452), .Z(n4455) );
  XOR U5351 ( .A(n4456), .B(n4455), .Z(c[1914]) );
  NAND U5352 ( .A(b[0]), .B(a[892]), .Z(n4459) );
  XOR U5353 ( .A(sreg[1915]), .B(n4459), .Z(n4461) );
  NANDN U5354 ( .A(n4454), .B(sreg[1914]), .Z(n4458) );
  OR U5355 ( .A(n4456), .B(n4455), .Z(n4457) );
  AND U5356 ( .A(n4458), .B(n4457), .Z(n4460) );
  XOR U5357 ( .A(n4461), .B(n4460), .Z(c[1915]) );
  NAND U5358 ( .A(b[0]), .B(a[893]), .Z(n4464) );
  XOR U5359 ( .A(sreg[1916]), .B(n4464), .Z(n4466) );
  NANDN U5360 ( .A(n4459), .B(sreg[1915]), .Z(n4463) );
  OR U5361 ( .A(n4461), .B(n4460), .Z(n4462) );
  AND U5362 ( .A(n4463), .B(n4462), .Z(n4465) );
  XOR U5363 ( .A(n4466), .B(n4465), .Z(c[1916]) );
  NAND U5364 ( .A(b[0]), .B(a[894]), .Z(n4469) );
  XOR U5365 ( .A(sreg[1917]), .B(n4469), .Z(n4471) );
  NANDN U5366 ( .A(n4464), .B(sreg[1916]), .Z(n4468) );
  OR U5367 ( .A(n4466), .B(n4465), .Z(n4467) );
  AND U5368 ( .A(n4468), .B(n4467), .Z(n4470) );
  XOR U5369 ( .A(n4471), .B(n4470), .Z(c[1917]) );
  NAND U5370 ( .A(b[0]), .B(a[895]), .Z(n4474) );
  XOR U5371 ( .A(sreg[1918]), .B(n4474), .Z(n4476) );
  NANDN U5372 ( .A(n4469), .B(sreg[1917]), .Z(n4473) );
  OR U5373 ( .A(n4471), .B(n4470), .Z(n4472) );
  AND U5374 ( .A(n4473), .B(n4472), .Z(n4475) );
  XOR U5375 ( .A(n4476), .B(n4475), .Z(c[1918]) );
  NAND U5376 ( .A(b[0]), .B(a[896]), .Z(n4479) );
  XOR U5377 ( .A(sreg[1919]), .B(n4479), .Z(n4481) );
  NANDN U5378 ( .A(n4474), .B(sreg[1918]), .Z(n4478) );
  OR U5379 ( .A(n4476), .B(n4475), .Z(n4477) );
  AND U5380 ( .A(n4478), .B(n4477), .Z(n4480) );
  XOR U5381 ( .A(n4481), .B(n4480), .Z(c[1919]) );
  NAND U5382 ( .A(b[0]), .B(a[897]), .Z(n4484) );
  XOR U5383 ( .A(sreg[1920]), .B(n4484), .Z(n4486) );
  NANDN U5384 ( .A(n4479), .B(sreg[1919]), .Z(n4483) );
  OR U5385 ( .A(n4481), .B(n4480), .Z(n4482) );
  AND U5386 ( .A(n4483), .B(n4482), .Z(n4485) );
  XOR U5387 ( .A(n4486), .B(n4485), .Z(c[1920]) );
  NAND U5388 ( .A(b[0]), .B(a[898]), .Z(n4489) );
  XOR U5389 ( .A(sreg[1921]), .B(n4489), .Z(n4491) );
  NANDN U5390 ( .A(n4484), .B(sreg[1920]), .Z(n4488) );
  OR U5391 ( .A(n4486), .B(n4485), .Z(n4487) );
  AND U5392 ( .A(n4488), .B(n4487), .Z(n4490) );
  XOR U5393 ( .A(n4491), .B(n4490), .Z(c[1921]) );
  NAND U5394 ( .A(b[0]), .B(a[899]), .Z(n4494) );
  XOR U5395 ( .A(sreg[1922]), .B(n4494), .Z(n4496) );
  NANDN U5396 ( .A(n4489), .B(sreg[1921]), .Z(n4493) );
  OR U5397 ( .A(n4491), .B(n4490), .Z(n4492) );
  AND U5398 ( .A(n4493), .B(n4492), .Z(n4495) );
  XOR U5399 ( .A(n4496), .B(n4495), .Z(c[1922]) );
  NAND U5400 ( .A(b[0]), .B(a[900]), .Z(n4499) );
  XOR U5401 ( .A(sreg[1923]), .B(n4499), .Z(n4501) );
  NANDN U5402 ( .A(n4494), .B(sreg[1922]), .Z(n4498) );
  OR U5403 ( .A(n4496), .B(n4495), .Z(n4497) );
  AND U5404 ( .A(n4498), .B(n4497), .Z(n4500) );
  XOR U5405 ( .A(n4501), .B(n4500), .Z(c[1923]) );
  NAND U5406 ( .A(b[0]), .B(a[901]), .Z(n4504) );
  XOR U5407 ( .A(sreg[1924]), .B(n4504), .Z(n4506) );
  NANDN U5408 ( .A(n4499), .B(sreg[1923]), .Z(n4503) );
  OR U5409 ( .A(n4501), .B(n4500), .Z(n4502) );
  AND U5410 ( .A(n4503), .B(n4502), .Z(n4505) );
  XOR U5411 ( .A(n4506), .B(n4505), .Z(c[1924]) );
  NAND U5412 ( .A(b[0]), .B(a[902]), .Z(n4509) );
  XOR U5413 ( .A(sreg[1925]), .B(n4509), .Z(n4511) );
  NANDN U5414 ( .A(n4504), .B(sreg[1924]), .Z(n4508) );
  OR U5415 ( .A(n4506), .B(n4505), .Z(n4507) );
  AND U5416 ( .A(n4508), .B(n4507), .Z(n4510) );
  XOR U5417 ( .A(n4511), .B(n4510), .Z(c[1925]) );
  NAND U5418 ( .A(b[0]), .B(a[903]), .Z(n4514) );
  XOR U5419 ( .A(sreg[1926]), .B(n4514), .Z(n4516) );
  NANDN U5420 ( .A(n4509), .B(sreg[1925]), .Z(n4513) );
  OR U5421 ( .A(n4511), .B(n4510), .Z(n4512) );
  AND U5422 ( .A(n4513), .B(n4512), .Z(n4515) );
  XOR U5423 ( .A(n4516), .B(n4515), .Z(c[1926]) );
  NAND U5424 ( .A(b[0]), .B(a[904]), .Z(n4519) );
  XOR U5425 ( .A(sreg[1927]), .B(n4519), .Z(n4521) );
  NANDN U5426 ( .A(n4514), .B(sreg[1926]), .Z(n4518) );
  OR U5427 ( .A(n4516), .B(n4515), .Z(n4517) );
  AND U5428 ( .A(n4518), .B(n4517), .Z(n4520) );
  XOR U5429 ( .A(n4521), .B(n4520), .Z(c[1927]) );
  NAND U5430 ( .A(b[0]), .B(a[905]), .Z(n4524) );
  XOR U5431 ( .A(sreg[1928]), .B(n4524), .Z(n4526) );
  NANDN U5432 ( .A(n4519), .B(sreg[1927]), .Z(n4523) );
  OR U5433 ( .A(n4521), .B(n4520), .Z(n4522) );
  AND U5434 ( .A(n4523), .B(n4522), .Z(n4525) );
  XOR U5435 ( .A(n4526), .B(n4525), .Z(c[1928]) );
  NAND U5436 ( .A(b[0]), .B(a[906]), .Z(n4529) );
  XOR U5437 ( .A(sreg[1929]), .B(n4529), .Z(n4531) );
  NANDN U5438 ( .A(n4524), .B(sreg[1928]), .Z(n4528) );
  OR U5439 ( .A(n4526), .B(n4525), .Z(n4527) );
  AND U5440 ( .A(n4528), .B(n4527), .Z(n4530) );
  XOR U5441 ( .A(n4531), .B(n4530), .Z(c[1929]) );
  NAND U5442 ( .A(b[0]), .B(a[907]), .Z(n4534) );
  XOR U5443 ( .A(sreg[1930]), .B(n4534), .Z(n4536) );
  NANDN U5444 ( .A(n4529), .B(sreg[1929]), .Z(n4533) );
  OR U5445 ( .A(n4531), .B(n4530), .Z(n4532) );
  AND U5446 ( .A(n4533), .B(n4532), .Z(n4535) );
  XOR U5447 ( .A(n4536), .B(n4535), .Z(c[1930]) );
  NAND U5448 ( .A(b[0]), .B(a[908]), .Z(n4539) );
  XOR U5449 ( .A(sreg[1931]), .B(n4539), .Z(n4541) );
  NANDN U5450 ( .A(n4534), .B(sreg[1930]), .Z(n4538) );
  OR U5451 ( .A(n4536), .B(n4535), .Z(n4537) );
  AND U5452 ( .A(n4538), .B(n4537), .Z(n4540) );
  XOR U5453 ( .A(n4541), .B(n4540), .Z(c[1931]) );
  NAND U5454 ( .A(b[0]), .B(a[909]), .Z(n4544) );
  XOR U5455 ( .A(sreg[1932]), .B(n4544), .Z(n4546) );
  NANDN U5456 ( .A(n4539), .B(sreg[1931]), .Z(n4543) );
  OR U5457 ( .A(n4541), .B(n4540), .Z(n4542) );
  AND U5458 ( .A(n4543), .B(n4542), .Z(n4545) );
  XOR U5459 ( .A(n4546), .B(n4545), .Z(c[1932]) );
  NAND U5460 ( .A(b[0]), .B(a[910]), .Z(n4549) );
  XOR U5461 ( .A(sreg[1933]), .B(n4549), .Z(n4551) );
  NANDN U5462 ( .A(n4544), .B(sreg[1932]), .Z(n4548) );
  OR U5463 ( .A(n4546), .B(n4545), .Z(n4547) );
  AND U5464 ( .A(n4548), .B(n4547), .Z(n4550) );
  XOR U5465 ( .A(n4551), .B(n4550), .Z(c[1933]) );
  NAND U5466 ( .A(b[0]), .B(a[911]), .Z(n4554) );
  XOR U5467 ( .A(sreg[1934]), .B(n4554), .Z(n4556) );
  NANDN U5468 ( .A(n4549), .B(sreg[1933]), .Z(n4553) );
  OR U5469 ( .A(n4551), .B(n4550), .Z(n4552) );
  AND U5470 ( .A(n4553), .B(n4552), .Z(n4555) );
  XOR U5471 ( .A(n4556), .B(n4555), .Z(c[1934]) );
  NAND U5472 ( .A(b[0]), .B(a[912]), .Z(n4559) );
  XOR U5473 ( .A(sreg[1935]), .B(n4559), .Z(n4561) );
  NANDN U5474 ( .A(n4554), .B(sreg[1934]), .Z(n4558) );
  OR U5475 ( .A(n4556), .B(n4555), .Z(n4557) );
  AND U5476 ( .A(n4558), .B(n4557), .Z(n4560) );
  XOR U5477 ( .A(n4561), .B(n4560), .Z(c[1935]) );
  NAND U5478 ( .A(b[0]), .B(a[913]), .Z(n4564) );
  XOR U5479 ( .A(sreg[1936]), .B(n4564), .Z(n4566) );
  NANDN U5480 ( .A(n4559), .B(sreg[1935]), .Z(n4563) );
  OR U5481 ( .A(n4561), .B(n4560), .Z(n4562) );
  AND U5482 ( .A(n4563), .B(n4562), .Z(n4565) );
  XOR U5483 ( .A(n4566), .B(n4565), .Z(c[1936]) );
  NAND U5484 ( .A(b[0]), .B(a[914]), .Z(n4569) );
  XOR U5485 ( .A(sreg[1937]), .B(n4569), .Z(n4571) );
  NANDN U5486 ( .A(n4564), .B(sreg[1936]), .Z(n4568) );
  OR U5487 ( .A(n4566), .B(n4565), .Z(n4567) );
  AND U5488 ( .A(n4568), .B(n4567), .Z(n4570) );
  XOR U5489 ( .A(n4571), .B(n4570), .Z(c[1937]) );
  NAND U5490 ( .A(b[0]), .B(a[915]), .Z(n4574) );
  XOR U5491 ( .A(sreg[1938]), .B(n4574), .Z(n4576) );
  NANDN U5492 ( .A(n4569), .B(sreg[1937]), .Z(n4573) );
  OR U5493 ( .A(n4571), .B(n4570), .Z(n4572) );
  AND U5494 ( .A(n4573), .B(n4572), .Z(n4575) );
  XOR U5495 ( .A(n4576), .B(n4575), .Z(c[1938]) );
  NAND U5496 ( .A(b[0]), .B(a[916]), .Z(n4579) );
  XOR U5497 ( .A(sreg[1939]), .B(n4579), .Z(n4581) );
  NANDN U5498 ( .A(n4574), .B(sreg[1938]), .Z(n4578) );
  OR U5499 ( .A(n4576), .B(n4575), .Z(n4577) );
  AND U5500 ( .A(n4578), .B(n4577), .Z(n4580) );
  XOR U5501 ( .A(n4581), .B(n4580), .Z(c[1939]) );
  NAND U5502 ( .A(b[0]), .B(a[917]), .Z(n4584) );
  XOR U5503 ( .A(sreg[1940]), .B(n4584), .Z(n4586) );
  NANDN U5504 ( .A(n4579), .B(sreg[1939]), .Z(n4583) );
  OR U5505 ( .A(n4581), .B(n4580), .Z(n4582) );
  AND U5506 ( .A(n4583), .B(n4582), .Z(n4585) );
  XOR U5507 ( .A(n4586), .B(n4585), .Z(c[1940]) );
  NAND U5508 ( .A(b[0]), .B(a[918]), .Z(n4589) );
  XOR U5509 ( .A(sreg[1941]), .B(n4589), .Z(n4591) );
  NANDN U5510 ( .A(n4584), .B(sreg[1940]), .Z(n4588) );
  OR U5511 ( .A(n4586), .B(n4585), .Z(n4587) );
  AND U5512 ( .A(n4588), .B(n4587), .Z(n4590) );
  XOR U5513 ( .A(n4591), .B(n4590), .Z(c[1941]) );
  NAND U5514 ( .A(b[0]), .B(a[919]), .Z(n4594) );
  XOR U5515 ( .A(sreg[1942]), .B(n4594), .Z(n4596) );
  NANDN U5516 ( .A(n4589), .B(sreg[1941]), .Z(n4593) );
  OR U5517 ( .A(n4591), .B(n4590), .Z(n4592) );
  AND U5518 ( .A(n4593), .B(n4592), .Z(n4595) );
  XOR U5519 ( .A(n4596), .B(n4595), .Z(c[1942]) );
  NAND U5520 ( .A(b[0]), .B(a[920]), .Z(n4599) );
  XOR U5521 ( .A(sreg[1943]), .B(n4599), .Z(n4601) );
  NANDN U5522 ( .A(n4594), .B(sreg[1942]), .Z(n4598) );
  OR U5523 ( .A(n4596), .B(n4595), .Z(n4597) );
  AND U5524 ( .A(n4598), .B(n4597), .Z(n4600) );
  XOR U5525 ( .A(n4601), .B(n4600), .Z(c[1943]) );
  NAND U5526 ( .A(b[0]), .B(a[921]), .Z(n4604) );
  XOR U5527 ( .A(sreg[1944]), .B(n4604), .Z(n4606) );
  NANDN U5528 ( .A(n4599), .B(sreg[1943]), .Z(n4603) );
  OR U5529 ( .A(n4601), .B(n4600), .Z(n4602) );
  AND U5530 ( .A(n4603), .B(n4602), .Z(n4605) );
  XOR U5531 ( .A(n4606), .B(n4605), .Z(c[1944]) );
  NAND U5532 ( .A(b[0]), .B(a[922]), .Z(n4609) );
  XOR U5533 ( .A(sreg[1945]), .B(n4609), .Z(n4611) );
  NANDN U5534 ( .A(n4604), .B(sreg[1944]), .Z(n4608) );
  OR U5535 ( .A(n4606), .B(n4605), .Z(n4607) );
  AND U5536 ( .A(n4608), .B(n4607), .Z(n4610) );
  XOR U5537 ( .A(n4611), .B(n4610), .Z(c[1945]) );
  NAND U5538 ( .A(b[0]), .B(a[923]), .Z(n4614) );
  XOR U5539 ( .A(sreg[1946]), .B(n4614), .Z(n4616) );
  NANDN U5540 ( .A(n4609), .B(sreg[1945]), .Z(n4613) );
  OR U5541 ( .A(n4611), .B(n4610), .Z(n4612) );
  AND U5542 ( .A(n4613), .B(n4612), .Z(n4615) );
  XOR U5543 ( .A(n4616), .B(n4615), .Z(c[1946]) );
  NAND U5544 ( .A(b[0]), .B(a[924]), .Z(n4619) );
  XOR U5545 ( .A(sreg[1947]), .B(n4619), .Z(n4621) );
  NANDN U5546 ( .A(n4614), .B(sreg[1946]), .Z(n4618) );
  OR U5547 ( .A(n4616), .B(n4615), .Z(n4617) );
  AND U5548 ( .A(n4618), .B(n4617), .Z(n4620) );
  XOR U5549 ( .A(n4621), .B(n4620), .Z(c[1947]) );
  NAND U5550 ( .A(b[0]), .B(a[925]), .Z(n4624) );
  XOR U5551 ( .A(sreg[1948]), .B(n4624), .Z(n4626) );
  NANDN U5552 ( .A(n4619), .B(sreg[1947]), .Z(n4623) );
  OR U5553 ( .A(n4621), .B(n4620), .Z(n4622) );
  AND U5554 ( .A(n4623), .B(n4622), .Z(n4625) );
  XOR U5555 ( .A(n4626), .B(n4625), .Z(c[1948]) );
  NAND U5556 ( .A(b[0]), .B(a[926]), .Z(n4629) );
  XOR U5557 ( .A(sreg[1949]), .B(n4629), .Z(n4631) );
  NANDN U5558 ( .A(n4624), .B(sreg[1948]), .Z(n4628) );
  OR U5559 ( .A(n4626), .B(n4625), .Z(n4627) );
  AND U5560 ( .A(n4628), .B(n4627), .Z(n4630) );
  XOR U5561 ( .A(n4631), .B(n4630), .Z(c[1949]) );
  NAND U5562 ( .A(b[0]), .B(a[927]), .Z(n4634) );
  XOR U5563 ( .A(sreg[1950]), .B(n4634), .Z(n4636) );
  NANDN U5564 ( .A(n4629), .B(sreg[1949]), .Z(n4633) );
  OR U5565 ( .A(n4631), .B(n4630), .Z(n4632) );
  AND U5566 ( .A(n4633), .B(n4632), .Z(n4635) );
  XOR U5567 ( .A(n4636), .B(n4635), .Z(c[1950]) );
  NAND U5568 ( .A(b[0]), .B(a[928]), .Z(n4639) );
  XOR U5569 ( .A(sreg[1951]), .B(n4639), .Z(n4641) );
  NANDN U5570 ( .A(n4634), .B(sreg[1950]), .Z(n4638) );
  OR U5571 ( .A(n4636), .B(n4635), .Z(n4637) );
  AND U5572 ( .A(n4638), .B(n4637), .Z(n4640) );
  XOR U5573 ( .A(n4641), .B(n4640), .Z(c[1951]) );
  NAND U5574 ( .A(b[0]), .B(a[929]), .Z(n4644) );
  XOR U5575 ( .A(sreg[1952]), .B(n4644), .Z(n4646) );
  NANDN U5576 ( .A(n4639), .B(sreg[1951]), .Z(n4643) );
  OR U5577 ( .A(n4641), .B(n4640), .Z(n4642) );
  AND U5578 ( .A(n4643), .B(n4642), .Z(n4645) );
  XOR U5579 ( .A(n4646), .B(n4645), .Z(c[1952]) );
  NAND U5580 ( .A(b[0]), .B(a[930]), .Z(n4649) );
  XOR U5581 ( .A(sreg[1953]), .B(n4649), .Z(n4651) );
  NANDN U5582 ( .A(n4644), .B(sreg[1952]), .Z(n4648) );
  OR U5583 ( .A(n4646), .B(n4645), .Z(n4647) );
  AND U5584 ( .A(n4648), .B(n4647), .Z(n4650) );
  XOR U5585 ( .A(n4651), .B(n4650), .Z(c[1953]) );
  NAND U5586 ( .A(b[0]), .B(a[931]), .Z(n4654) );
  XOR U5587 ( .A(sreg[1954]), .B(n4654), .Z(n4656) );
  NANDN U5588 ( .A(n4649), .B(sreg[1953]), .Z(n4653) );
  OR U5589 ( .A(n4651), .B(n4650), .Z(n4652) );
  AND U5590 ( .A(n4653), .B(n4652), .Z(n4655) );
  XOR U5591 ( .A(n4656), .B(n4655), .Z(c[1954]) );
  NAND U5592 ( .A(b[0]), .B(a[932]), .Z(n4659) );
  XOR U5593 ( .A(sreg[1955]), .B(n4659), .Z(n4661) );
  NANDN U5594 ( .A(n4654), .B(sreg[1954]), .Z(n4658) );
  OR U5595 ( .A(n4656), .B(n4655), .Z(n4657) );
  AND U5596 ( .A(n4658), .B(n4657), .Z(n4660) );
  XOR U5597 ( .A(n4661), .B(n4660), .Z(c[1955]) );
  NAND U5598 ( .A(b[0]), .B(a[933]), .Z(n4664) );
  XOR U5599 ( .A(sreg[1956]), .B(n4664), .Z(n4666) );
  NANDN U5600 ( .A(n4659), .B(sreg[1955]), .Z(n4663) );
  OR U5601 ( .A(n4661), .B(n4660), .Z(n4662) );
  AND U5602 ( .A(n4663), .B(n4662), .Z(n4665) );
  XOR U5603 ( .A(n4666), .B(n4665), .Z(c[1956]) );
  NAND U5604 ( .A(b[0]), .B(a[934]), .Z(n4669) );
  XOR U5605 ( .A(sreg[1957]), .B(n4669), .Z(n4671) );
  NANDN U5606 ( .A(n4664), .B(sreg[1956]), .Z(n4668) );
  OR U5607 ( .A(n4666), .B(n4665), .Z(n4667) );
  AND U5608 ( .A(n4668), .B(n4667), .Z(n4670) );
  XOR U5609 ( .A(n4671), .B(n4670), .Z(c[1957]) );
  NAND U5610 ( .A(b[0]), .B(a[935]), .Z(n4674) );
  XOR U5611 ( .A(sreg[1958]), .B(n4674), .Z(n4676) );
  NANDN U5612 ( .A(n4669), .B(sreg[1957]), .Z(n4673) );
  OR U5613 ( .A(n4671), .B(n4670), .Z(n4672) );
  AND U5614 ( .A(n4673), .B(n4672), .Z(n4675) );
  XOR U5615 ( .A(n4676), .B(n4675), .Z(c[1958]) );
  NAND U5616 ( .A(b[0]), .B(a[936]), .Z(n4679) );
  XOR U5617 ( .A(sreg[1959]), .B(n4679), .Z(n4681) );
  NANDN U5618 ( .A(n4674), .B(sreg[1958]), .Z(n4678) );
  OR U5619 ( .A(n4676), .B(n4675), .Z(n4677) );
  AND U5620 ( .A(n4678), .B(n4677), .Z(n4680) );
  XOR U5621 ( .A(n4681), .B(n4680), .Z(c[1959]) );
  NAND U5622 ( .A(b[0]), .B(a[937]), .Z(n4684) );
  XOR U5623 ( .A(sreg[1960]), .B(n4684), .Z(n4686) );
  NANDN U5624 ( .A(n4679), .B(sreg[1959]), .Z(n4683) );
  OR U5625 ( .A(n4681), .B(n4680), .Z(n4682) );
  AND U5626 ( .A(n4683), .B(n4682), .Z(n4685) );
  XOR U5627 ( .A(n4686), .B(n4685), .Z(c[1960]) );
  NAND U5628 ( .A(b[0]), .B(a[938]), .Z(n4689) );
  XOR U5629 ( .A(sreg[1961]), .B(n4689), .Z(n4691) );
  NANDN U5630 ( .A(n4684), .B(sreg[1960]), .Z(n4688) );
  OR U5631 ( .A(n4686), .B(n4685), .Z(n4687) );
  AND U5632 ( .A(n4688), .B(n4687), .Z(n4690) );
  XOR U5633 ( .A(n4691), .B(n4690), .Z(c[1961]) );
  NAND U5634 ( .A(b[0]), .B(a[939]), .Z(n4694) );
  XOR U5635 ( .A(sreg[1962]), .B(n4694), .Z(n4696) );
  NANDN U5636 ( .A(n4689), .B(sreg[1961]), .Z(n4693) );
  OR U5637 ( .A(n4691), .B(n4690), .Z(n4692) );
  AND U5638 ( .A(n4693), .B(n4692), .Z(n4695) );
  XOR U5639 ( .A(n4696), .B(n4695), .Z(c[1962]) );
  NAND U5640 ( .A(b[0]), .B(a[940]), .Z(n4699) );
  XOR U5641 ( .A(sreg[1963]), .B(n4699), .Z(n4701) );
  NANDN U5642 ( .A(n4694), .B(sreg[1962]), .Z(n4698) );
  OR U5643 ( .A(n4696), .B(n4695), .Z(n4697) );
  AND U5644 ( .A(n4698), .B(n4697), .Z(n4700) );
  XOR U5645 ( .A(n4701), .B(n4700), .Z(c[1963]) );
  NAND U5646 ( .A(b[0]), .B(a[941]), .Z(n4704) );
  XOR U5647 ( .A(sreg[1964]), .B(n4704), .Z(n4706) );
  NANDN U5648 ( .A(n4699), .B(sreg[1963]), .Z(n4703) );
  OR U5649 ( .A(n4701), .B(n4700), .Z(n4702) );
  AND U5650 ( .A(n4703), .B(n4702), .Z(n4705) );
  XOR U5651 ( .A(n4706), .B(n4705), .Z(c[1964]) );
  NAND U5652 ( .A(b[0]), .B(a[942]), .Z(n4709) );
  XOR U5653 ( .A(sreg[1965]), .B(n4709), .Z(n4711) );
  NANDN U5654 ( .A(n4704), .B(sreg[1964]), .Z(n4708) );
  OR U5655 ( .A(n4706), .B(n4705), .Z(n4707) );
  AND U5656 ( .A(n4708), .B(n4707), .Z(n4710) );
  XOR U5657 ( .A(n4711), .B(n4710), .Z(c[1965]) );
  NAND U5658 ( .A(b[0]), .B(a[943]), .Z(n4714) );
  XOR U5659 ( .A(sreg[1966]), .B(n4714), .Z(n4716) );
  NANDN U5660 ( .A(n4709), .B(sreg[1965]), .Z(n4713) );
  OR U5661 ( .A(n4711), .B(n4710), .Z(n4712) );
  AND U5662 ( .A(n4713), .B(n4712), .Z(n4715) );
  XOR U5663 ( .A(n4716), .B(n4715), .Z(c[1966]) );
  NAND U5664 ( .A(b[0]), .B(a[944]), .Z(n4719) );
  XOR U5665 ( .A(sreg[1967]), .B(n4719), .Z(n4721) );
  NANDN U5666 ( .A(n4714), .B(sreg[1966]), .Z(n4718) );
  OR U5667 ( .A(n4716), .B(n4715), .Z(n4717) );
  AND U5668 ( .A(n4718), .B(n4717), .Z(n4720) );
  XOR U5669 ( .A(n4721), .B(n4720), .Z(c[1967]) );
  NAND U5670 ( .A(b[0]), .B(a[945]), .Z(n4724) );
  XOR U5671 ( .A(sreg[1968]), .B(n4724), .Z(n4726) );
  NANDN U5672 ( .A(n4719), .B(sreg[1967]), .Z(n4723) );
  OR U5673 ( .A(n4721), .B(n4720), .Z(n4722) );
  AND U5674 ( .A(n4723), .B(n4722), .Z(n4725) );
  XOR U5675 ( .A(n4726), .B(n4725), .Z(c[1968]) );
  NAND U5676 ( .A(b[0]), .B(a[946]), .Z(n4729) );
  XOR U5677 ( .A(sreg[1969]), .B(n4729), .Z(n4731) );
  NANDN U5678 ( .A(n4724), .B(sreg[1968]), .Z(n4728) );
  OR U5679 ( .A(n4726), .B(n4725), .Z(n4727) );
  AND U5680 ( .A(n4728), .B(n4727), .Z(n4730) );
  XOR U5681 ( .A(n4731), .B(n4730), .Z(c[1969]) );
  NAND U5682 ( .A(b[0]), .B(a[947]), .Z(n4734) );
  XOR U5683 ( .A(sreg[1970]), .B(n4734), .Z(n4736) );
  NANDN U5684 ( .A(n4729), .B(sreg[1969]), .Z(n4733) );
  OR U5685 ( .A(n4731), .B(n4730), .Z(n4732) );
  AND U5686 ( .A(n4733), .B(n4732), .Z(n4735) );
  XOR U5687 ( .A(n4736), .B(n4735), .Z(c[1970]) );
  NAND U5688 ( .A(b[0]), .B(a[948]), .Z(n4739) );
  XOR U5689 ( .A(sreg[1971]), .B(n4739), .Z(n4741) );
  NANDN U5690 ( .A(n4734), .B(sreg[1970]), .Z(n4738) );
  OR U5691 ( .A(n4736), .B(n4735), .Z(n4737) );
  AND U5692 ( .A(n4738), .B(n4737), .Z(n4740) );
  XOR U5693 ( .A(n4741), .B(n4740), .Z(c[1971]) );
  NAND U5694 ( .A(b[0]), .B(a[949]), .Z(n4744) );
  XOR U5695 ( .A(sreg[1972]), .B(n4744), .Z(n4746) );
  NANDN U5696 ( .A(n4739), .B(sreg[1971]), .Z(n4743) );
  OR U5697 ( .A(n4741), .B(n4740), .Z(n4742) );
  AND U5698 ( .A(n4743), .B(n4742), .Z(n4745) );
  XOR U5699 ( .A(n4746), .B(n4745), .Z(c[1972]) );
  NAND U5700 ( .A(b[0]), .B(a[950]), .Z(n4749) );
  XOR U5701 ( .A(sreg[1973]), .B(n4749), .Z(n4751) );
  NANDN U5702 ( .A(n4744), .B(sreg[1972]), .Z(n4748) );
  OR U5703 ( .A(n4746), .B(n4745), .Z(n4747) );
  AND U5704 ( .A(n4748), .B(n4747), .Z(n4750) );
  XOR U5705 ( .A(n4751), .B(n4750), .Z(c[1973]) );
  NAND U5706 ( .A(b[0]), .B(a[951]), .Z(n4754) );
  XOR U5707 ( .A(sreg[1974]), .B(n4754), .Z(n4756) );
  NANDN U5708 ( .A(n4749), .B(sreg[1973]), .Z(n4753) );
  OR U5709 ( .A(n4751), .B(n4750), .Z(n4752) );
  AND U5710 ( .A(n4753), .B(n4752), .Z(n4755) );
  XOR U5711 ( .A(n4756), .B(n4755), .Z(c[1974]) );
  NAND U5712 ( .A(b[0]), .B(a[952]), .Z(n4759) );
  XOR U5713 ( .A(sreg[1975]), .B(n4759), .Z(n4761) );
  NANDN U5714 ( .A(n4754), .B(sreg[1974]), .Z(n4758) );
  OR U5715 ( .A(n4756), .B(n4755), .Z(n4757) );
  AND U5716 ( .A(n4758), .B(n4757), .Z(n4760) );
  XOR U5717 ( .A(n4761), .B(n4760), .Z(c[1975]) );
  NAND U5718 ( .A(b[0]), .B(a[953]), .Z(n4764) );
  XOR U5719 ( .A(sreg[1976]), .B(n4764), .Z(n4766) );
  NANDN U5720 ( .A(n4759), .B(sreg[1975]), .Z(n4763) );
  OR U5721 ( .A(n4761), .B(n4760), .Z(n4762) );
  AND U5722 ( .A(n4763), .B(n4762), .Z(n4765) );
  XOR U5723 ( .A(n4766), .B(n4765), .Z(c[1976]) );
  NAND U5724 ( .A(b[0]), .B(a[954]), .Z(n4769) );
  XOR U5725 ( .A(sreg[1977]), .B(n4769), .Z(n4771) );
  NANDN U5726 ( .A(n4764), .B(sreg[1976]), .Z(n4768) );
  OR U5727 ( .A(n4766), .B(n4765), .Z(n4767) );
  AND U5728 ( .A(n4768), .B(n4767), .Z(n4770) );
  XOR U5729 ( .A(n4771), .B(n4770), .Z(c[1977]) );
  NAND U5730 ( .A(b[0]), .B(a[955]), .Z(n4774) );
  XOR U5731 ( .A(sreg[1978]), .B(n4774), .Z(n4776) );
  NANDN U5732 ( .A(n4769), .B(sreg[1977]), .Z(n4773) );
  OR U5733 ( .A(n4771), .B(n4770), .Z(n4772) );
  AND U5734 ( .A(n4773), .B(n4772), .Z(n4775) );
  XOR U5735 ( .A(n4776), .B(n4775), .Z(c[1978]) );
  NAND U5736 ( .A(b[0]), .B(a[956]), .Z(n4779) );
  XOR U5737 ( .A(sreg[1979]), .B(n4779), .Z(n4781) );
  NANDN U5738 ( .A(n4774), .B(sreg[1978]), .Z(n4778) );
  OR U5739 ( .A(n4776), .B(n4775), .Z(n4777) );
  AND U5740 ( .A(n4778), .B(n4777), .Z(n4780) );
  XOR U5741 ( .A(n4781), .B(n4780), .Z(c[1979]) );
  NAND U5742 ( .A(b[0]), .B(a[957]), .Z(n4784) );
  XOR U5743 ( .A(sreg[1980]), .B(n4784), .Z(n4786) );
  NANDN U5744 ( .A(n4779), .B(sreg[1979]), .Z(n4783) );
  OR U5745 ( .A(n4781), .B(n4780), .Z(n4782) );
  AND U5746 ( .A(n4783), .B(n4782), .Z(n4785) );
  XOR U5747 ( .A(n4786), .B(n4785), .Z(c[1980]) );
  NAND U5748 ( .A(b[0]), .B(a[958]), .Z(n4789) );
  XOR U5749 ( .A(sreg[1981]), .B(n4789), .Z(n4791) );
  NANDN U5750 ( .A(n4784), .B(sreg[1980]), .Z(n4788) );
  OR U5751 ( .A(n4786), .B(n4785), .Z(n4787) );
  AND U5752 ( .A(n4788), .B(n4787), .Z(n4790) );
  XOR U5753 ( .A(n4791), .B(n4790), .Z(c[1981]) );
  NAND U5754 ( .A(b[0]), .B(a[959]), .Z(n4794) );
  XOR U5755 ( .A(sreg[1982]), .B(n4794), .Z(n4796) );
  NANDN U5756 ( .A(n4789), .B(sreg[1981]), .Z(n4793) );
  OR U5757 ( .A(n4791), .B(n4790), .Z(n4792) );
  AND U5758 ( .A(n4793), .B(n4792), .Z(n4795) );
  XOR U5759 ( .A(n4796), .B(n4795), .Z(c[1982]) );
  NAND U5760 ( .A(b[0]), .B(a[960]), .Z(n4799) );
  XOR U5761 ( .A(sreg[1983]), .B(n4799), .Z(n4801) );
  NANDN U5762 ( .A(n4794), .B(sreg[1982]), .Z(n4798) );
  OR U5763 ( .A(n4796), .B(n4795), .Z(n4797) );
  AND U5764 ( .A(n4798), .B(n4797), .Z(n4800) );
  XOR U5765 ( .A(n4801), .B(n4800), .Z(c[1983]) );
  NAND U5766 ( .A(b[0]), .B(a[961]), .Z(n4804) );
  XOR U5767 ( .A(sreg[1984]), .B(n4804), .Z(n4806) );
  NANDN U5768 ( .A(n4799), .B(sreg[1983]), .Z(n4803) );
  OR U5769 ( .A(n4801), .B(n4800), .Z(n4802) );
  AND U5770 ( .A(n4803), .B(n4802), .Z(n4805) );
  XOR U5771 ( .A(n4806), .B(n4805), .Z(c[1984]) );
  NAND U5772 ( .A(b[0]), .B(a[962]), .Z(n4809) );
  XOR U5773 ( .A(sreg[1985]), .B(n4809), .Z(n4811) );
  NANDN U5774 ( .A(n4804), .B(sreg[1984]), .Z(n4808) );
  OR U5775 ( .A(n4806), .B(n4805), .Z(n4807) );
  AND U5776 ( .A(n4808), .B(n4807), .Z(n4810) );
  XOR U5777 ( .A(n4811), .B(n4810), .Z(c[1985]) );
  NAND U5778 ( .A(b[0]), .B(a[963]), .Z(n4814) );
  XOR U5779 ( .A(sreg[1986]), .B(n4814), .Z(n4816) );
  NANDN U5780 ( .A(n4809), .B(sreg[1985]), .Z(n4813) );
  OR U5781 ( .A(n4811), .B(n4810), .Z(n4812) );
  AND U5782 ( .A(n4813), .B(n4812), .Z(n4815) );
  XOR U5783 ( .A(n4816), .B(n4815), .Z(c[1986]) );
  NAND U5784 ( .A(b[0]), .B(a[964]), .Z(n4819) );
  XOR U5785 ( .A(sreg[1987]), .B(n4819), .Z(n4821) );
  NANDN U5786 ( .A(n4814), .B(sreg[1986]), .Z(n4818) );
  OR U5787 ( .A(n4816), .B(n4815), .Z(n4817) );
  AND U5788 ( .A(n4818), .B(n4817), .Z(n4820) );
  XOR U5789 ( .A(n4821), .B(n4820), .Z(c[1987]) );
  NAND U5790 ( .A(b[0]), .B(a[965]), .Z(n4824) );
  XOR U5791 ( .A(sreg[1988]), .B(n4824), .Z(n4826) );
  NANDN U5792 ( .A(n4819), .B(sreg[1987]), .Z(n4823) );
  OR U5793 ( .A(n4821), .B(n4820), .Z(n4822) );
  AND U5794 ( .A(n4823), .B(n4822), .Z(n4825) );
  XOR U5795 ( .A(n4826), .B(n4825), .Z(c[1988]) );
  NAND U5796 ( .A(b[0]), .B(a[966]), .Z(n4829) );
  XOR U5797 ( .A(sreg[1989]), .B(n4829), .Z(n4831) );
  NANDN U5798 ( .A(n4824), .B(sreg[1988]), .Z(n4828) );
  OR U5799 ( .A(n4826), .B(n4825), .Z(n4827) );
  AND U5800 ( .A(n4828), .B(n4827), .Z(n4830) );
  XOR U5801 ( .A(n4831), .B(n4830), .Z(c[1989]) );
  NAND U5802 ( .A(b[0]), .B(a[967]), .Z(n4834) );
  XOR U5803 ( .A(sreg[1990]), .B(n4834), .Z(n4836) );
  NANDN U5804 ( .A(n4829), .B(sreg[1989]), .Z(n4833) );
  OR U5805 ( .A(n4831), .B(n4830), .Z(n4832) );
  AND U5806 ( .A(n4833), .B(n4832), .Z(n4835) );
  XOR U5807 ( .A(n4836), .B(n4835), .Z(c[1990]) );
  NAND U5808 ( .A(b[0]), .B(a[968]), .Z(n4839) );
  XOR U5809 ( .A(sreg[1991]), .B(n4839), .Z(n4841) );
  NANDN U5810 ( .A(n4834), .B(sreg[1990]), .Z(n4838) );
  OR U5811 ( .A(n4836), .B(n4835), .Z(n4837) );
  AND U5812 ( .A(n4838), .B(n4837), .Z(n4840) );
  XOR U5813 ( .A(n4841), .B(n4840), .Z(c[1991]) );
  NAND U5814 ( .A(b[0]), .B(a[969]), .Z(n4844) );
  XOR U5815 ( .A(sreg[1992]), .B(n4844), .Z(n4846) );
  NANDN U5816 ( .A(n4839), .B(sreg[1991]), .Z(n4843) );
  OR U5817 ( .A(n4841), .B(n4840), .Z(n4842) );
  AND U5818 ( .A(n4843), .B(n4842), .Z(n4845) );
  XOR U5819 ( .A(n4846), .B(n4845), .Z(c[1992]) );
  NAND U5820 ( .A(b[0]), .B(a[970]), .Z(n4849) );
  XOR U5821 ( .A(sreg[1993]), .B(n4849), .Z(n4851) );
  NANDN U5822 ( .A(n4844), .B(sreg[1992]), .Z(n4848) );
  OR U5823 ( .A(n4846), .B(n4845), .Z(n4847) );
  AND U5824 ( .A(n4848), .B(n4847), .Z(n4850) );
  XOR U5825 ( .A(n4851), .B(n4850), .Z(c[1993]) );
  NAND U5826 ( .A(b[0]), .B(a[971]), .Z(n4854) );
  XOR U5827 ( .A(sreg[1994]), .B(n4854), .Z(n4856) );
  NANDN U5828 ( .A(n4849), .B(sreg[1993]), .Z(n4853) );
  OR U5829 ( .A(n4851), .B(n4850), .Z(n4852) );
  AND U5830 ( .A(n4853), .B(n4852), .Z(n4855) );
  XOR U5831 ( .A(n4856), .B(n4855), .Z(c[1994]) );
  NAND U5832 ( .A(b[0]), .B(a[972]), .Z(n4859) );
  XOR U5833 ( .A(sreg[1995]), .B(n4859), .Z(n4861) );
  NANDN U5834 ( .A(n4854), .B(sreg[1994]), .Z(n4858) );
  OR U5835 ( .A(n4856), .B(n4855), .Z(n4857) );
  AND U5836 ( .A(n4858), .B(n4857), .Z(n4860) );
  XOR U5837 ( .A(n4861), .B(n4860), .Z(c[1995]) );
  NAND U5838 ( .A(b[0]), .B(a[973]), .Z(n4864) );
  XOR U5839 ( .A(sreg[1996]), .B(n4864), .Z(n4866) );
  NANDN U5840 ( .A(n4859), .B(sreg[1995]), .Z(n4863) );
  OR U5841 ( .A(n4861), .B(n4860), .Z(n4862) );
  AND U5842 ( .A(n4863), .B(n4862), .Z(n4865) );
  XOR U5843 ( .A(n4866), .B(n4865), .Z(c[1996]) );
  NAND U5844 ( .A(b[0]), .B(a[974]), .Z(n4869) );
  XOR U5845 ( .A(sreg[1997]), .B(n4869), .Z(n4871) );
  NANDN U5846 ( .A(n4864), .B(sreg[1996]), .Z(n4868) );
  OR U5847 ( .A(n4866), .B(n4865), .Z(n4867) );
  AND U5848 ( .A(n4868), .B(n4867), .Z(n4870) );
  XOR U5849 ( .A(n4871), .B(n4870), .Z(c[1997]) );
  NAND U5850 ( .A(b[0]), .B(a[975]), .Z(n4874) );
  XOR U5851 ( .A(sreg[1998]), .B(n4874), .Z(n4876) );
  NANDN U5852 ( .A(n4869), .B(sreg[1997]), .Z(n4873) );
  OR U5853 ( .A(n4871), .B(n4870), .Z(n4872) );
  AND U5854 ( .A(n4873), .B(n4872), .Z(n4875) );
  XOR U5855 ( .A(n4876), .B(n4875), .Z(c[1998]) );
  NAND U5856 ( .A(b[0]), .B(a[976]), .Z(n4879) );
  XOR U5857 ( .A(sreg[1999]), .B(n4879), .Z(n4881) );
  NANDN U5858 ( .A(n4874), .B(sreg[1998]), .Z(n4878) );
  OR U5859 ( .A(n4876), .B(n4875), .Z(n4877) );
  AND U5860 ( .A(n4878), .B(n4877), .Z(n4880) );
  XOR U5861 ( .A(n4881), .B(n4880), .Z(c[1999]) );
  NAND U5862 ( .A(b[0]), .B(a[977]), .Z(n4884) );
  XOR U5863 ( .A(sreg[2000]), .B(n4884), .Z(n4886) );
  NANDN U5864 ( .A(n4879), .B(sreg[1999]), .Z(n4883) );
  OR U5865 ( .A(n4881), .B(n4880), .Z(n4882) );
  AND U5866 ( .A(n4883), .B(n4882), .Z(n4885) );
  XOR U5867 ( .A(n4886), .B(n4885), .Z(c[2000]) );
  NAND U5868 ( .A(b[0]), .B(a[978]), .Z(n4889) );
  XOR U5869 ( .A(sreg[2001]), .B(n4889), .Z(n4891) );
  NANDN U5870 ( .A(n4884), .B(sreg[2000]), .Z(n4888) );
  OR U5871 ( .A(n4886), .B(n4885), .Z(n4887) );
  AND U5872 ( .A(n4888), .B(n4887), .Z(n4890) );
  XOR U5873 ( .A(n4891), .B(n4890), .Z(c[2001]) );
  NAND U5874 ( .A(b[0]), .B(a[979]), .Z(n4894) );
  XOR U5875 ( .A(sreg[2002]), .B(n4894), .Z(n4896) );
  NANDN U5876 ( .A(n4889), .B(sreg[2001]), .Z(n4893) );
  OR U5877 ( .A(n4891), .B(n4890), .Z(n4892) );
  AND U5878 ( .A(n4893), .B(n4892), .Z(n4895) );
  XOR U5879 ( .A(n4896), .B(n4895), .Z(c[2002]) );
  NAND U5880 ( .A(b[0]), .B(a[980]), .Z(n4899) );
  XOR U5881 ( .A(sreg[2003]), .B(n4899), .Z(n4901) );
  NANDN U5882 ( .A(n4894), .B(sreg[2002]), .Z(n4898) );
  OR U5883 ( .A(n4896), .B(n4895), .Z(n4897) );
  AND U5884 ( .A(n4898), .B(n4897), .Z(n4900) );
  XOR U5885 ( .A(n4901), .B(n4900), .Z(c[2003]) );
  NAND U5886 ( .A(b[0]), .B(a[981]), .Z(n4904) );
  XOR U5887 ( .A(sreg[2004]), .B(n4904), .Z(n4906) );
  NANDN U5888 ( .A(n4899), .B(sreg[2003]), .Z(n4903) );
  OR U5889 ( .A(n4901), .B(n4900), .Z(n4902) );
  AND U5890 ( .A(n4903), .B(n4902), .Z(n4905) );
  XOR U5891 ( .A(n4906), .B(n4905), .Z(c[2004]) );
  NAND U5892 ( .A(b[0]), .B(a[982]), .Z(n4909) );
  XOR U5893 ( .A(sreg[2005]), .B(n4909), .Z(n4911) );
  NANDN U5894 ( .A(n4904), .B(sreg[2004]), .Z(n4908) );
  OR U5895 ( .A(n4906), .B(n4905), .Z(n4907) );
  AND U5896 ( .A(n4908), .B(n4907), .Z(n4910) );
  XOR U5897 ( .A(n4911), .B(n4910), .Z(c[2005]) );
  NAND U5898 ( .A(b[0]), .B(a[983]), .Z(n4914) );
  XOR U5899 ( .A(sreg[2006]), .B(n4914), .Z(n4916) );
  NANDN U5900 ( .A(n4909), .B(sreg[2005]), .Z(n4913) );
  OR U5901 ( .A(n4911), .B(n4910), .Z(n4912) );
  AND U5902 ( .A(n4913), .B(n4912), .Z(n4915) );
  XOR U5903 ( .A(n4916), .B(n4915), .Z(c[2006]) );
  NAND U5904 ( .A(b[0]), .B(a[984]), .Z(n4919) );
  XOR U5905 ( .A(sreg[2007]), .B(n4919), .Z(n4921) );
  NANDN U5906 ( .A(n4914), .B(sreg[2006]), .Z(n4918) );
  OR U5907 ( .A(n4916), .B(n4915), .Z(n4917) );
  AND U5908 ( .A(n4918), .B(n4917), .Z(n4920) );
  XOR U5909 ( .A(n4921), .B(n4920), .Z(c[2007]) );
  NAND U5910 ( .A(b[0]), .B(a[985]), .Z(n4924) );
  XOR U5911 ( .A(sreg[2008]), .B(n4924), .Z(n4926) );
  NANDN U5912 ( .A(n4919), .B(sreg[2007]), .Z(n4923) );
  OR U5913 ( .A(n4921), .B(n4920), .Z(n4922) );
  AND U5914 ( .A(n4923), .B(n4922), .Z(n4925) );
  XOR U5915 ( .A(n4926), .B(n4925), .Z(c[2008]) );
  NAND U5916 ( .A(b[0]), .B(a[986]), .Z(n4929) );
  XOR U5917 ( .A(sreg[2009]), .B(n4929), .Z(n4931) );
  NANDN U5918 ( .A(n4924), .B(sreg[2008]), .Z(n4928) );
  OR U5919 ( .A(n4926), .B(n4925), .Z(n4927) );
  AND U5920 ( .A(n4928), .B(n4927), .Z(n4930) );
  XOR U5921 ( .A(n4931), .B(n4930), .Z(c[2009]) );
  NAND U5922 ( .A(b[0]), .B(a[987]), .Z(n4934) );
  XOR U5923 ( .A(sreg[2010]), .B(n4934), .Z(n4936) );
  NANDN U5924 ( .A(n4929), .B(sreg[2009]), .Z(n4933) );
  OR U5925 ( .A(n4931), .B(n4930), .Z(n4932) );
  AND U5926 ( .A(n4933), .B(n4932), .Z(n4935) );
  XOR U5927 ( .A(n4936), .B(n4935), .Z(c[2010]) );
  NAND U5928 ( .A(b[0]), .B(a[988]), .Z(n4939) );
  XOR U5929 ( .A(sreg[2011]), .B(n4939), .Z(n4941) );
  NANDN U5930 ( .A(n4934), .B(sreg[2010]), .Z(n4938) );
  OR U5931 ( .A(n4936), .B(n4935), .Z(n4937) );
  AND U5932 ( .A(n4938), .B(n4937), .Z(n4940) );
  XOR U5933 ( .A(n4941), .B(n4940), .Z(c[2011]) );
  NAND U5934 ( .A(b[0]), .B(a[989]), .Z(n4944) );
  XOR U5935 ( .A(sreg[2012]), .B(n4944), .Z(n4946) );
  NANDN U5936 ( .A(n4939), .B(sreg[2011]), .Z(n4943) );
  OR U5937 ( .A(n4941), .B(n4940), .Z(n4942) );
  AND U5938 ( .A(n4943), .B(n4942), .Z(n4945) );
  XOR U5939 ( .A(n4946), .B(n4945), .Z(c[2012]) );
  NAND U5940 ( .A(b[0]), .B(a[990]), .Z(n4949) );
  XOR U5941 ( .A(sreg[2013]), .B(n4949), .Z(n4951) );
  NANDN U5942 ( .A(n4944), .B(sreg[2012]), .Z(n4948) );
  OR U5943 ( .A(n4946), .B(n4945), .Z(n4947) );
  AND U5944 ( .A(n4948), .B(n4947), .Z(n4950) );
  XOR U5945 ( .A(n4951), .B(n4950), .Z(c[2013]) );
  NAND U5946 ( .A(b[0]), .B(a[991]), .Z(n4954) );
  XOR U5947 ( .A(sreg[2014]), .B(n4954), .Z(n4956) );
  NANDN U5948 ( .A(n4949), .B(sreg[2013]), .Z(n4953) );
  OR U5949 ( .A(n4951), .B(n4950), .Z(n4952) );
  AND U5950 ( .A(n4953), .B(n4952), .Z(n4955) );
  XOR U5951 ( .A(n4956), .B(n4955), .Z(c[2014]) );
  NAND U5952 ( .A(b[0]), .B(a[992]), .Z(n4959) );
  XOR U5953 ( .A(sreg[2015]), .B(n4959), .Z(n4961) );
  NANDN U5954 ( .A(n4954), .B(sreg[2014]), .Z(n4958) );
  OR U5955 ( .A(n4956), .B(n4955), .Z(n4957) );
  AND U5956 ( .A(n4958), .B(n4957), .Z(n4960) );
  XOR U5957 ( .A(n4961), .B(n4960), .Z(c[2015]) );
  NAND U5958 ( .A(b[0]), .B(a[993]), .Z(n4964) );
  XOR U5959 ( .A(sreg[2016]), .B(n4964), .Z(n4966) );
  NANDN U5960 ( .A(n4959), .B(sreg[2015]), .Z(n4963) );
  OR U5961 ( .A(n4961), .B(n4960), .Z(n4962) );
  AND U5962 ( .A(n4963), .B(n4962), .Z(n4965) );
  XOR U5963 ( .A(n4966), .B(n4965), .Z(c[2016]) );
  NAND U5964 ( .A(b[0]), .B(a[994]), .Z(n4969) );
  XOR U5965 ( .A(sreg[2017]), .B(n4969), .Z(n4971) );
  NANDN U5966 ( .A(n4964), .B(sreg[2016]), .Z(n4968) );
  OR U5967 ( .A(n4966), .B(n4965), .Z(n4967) );
  AND U5968 ( .A(n4968), .B(n4967), .Z(n4970) );
  XOR U5969 ( .A(n4971), .B(n4970), .Z(c[2017]) );
  NAND U5970 ( .A(b[0]), .B(a[995]), .Z(n4974) );
  XOR U5971 ( .A(sreg[2018]), .B(n4974), .Z(n4976) );
  NANDN U5972 ( .A(n4969), .B(sreg[2017]), .Z(n4973) );
  OR U5973 ( .A(n4971), .B(n4970), .Z(n4972) );
  AND U5974 ( .A(n4973), .B(n4972), .Z(n4975) );
  XOR U5975 ( .A(n4976), .B(n4975), .Z(c[2018]) );
  NAND U5976 ( .A(b[0]), .B(a[996]), .Z(n4979) );
  XOR U5977 ( .A(sreg[2019]), .B(n4979), .Z(n4981) );
  NANDN U5978 ( .A(n4974), .B(sreg[2018]), .Z(n4978) );
  OR U5979 ( .A(n4976), .B(n4975), .Z(n4977) );
  AND U5980 ( .A(n4978), .B(n4977), .Z(n4980) );
  XOR U5981 ( .A(n4981), .B(n4980), .Z(c[2019]) );
  NAND U5982 ( .A(b[0]), .B(a[997]), .Z(n4984) );
  XOR U5983 ( .A(sreg[2020]), .B(n4984), .Z(n4986) );
  NANDN U5984 ( .A(n4979), .B(sreg[2019]), .Z(n4983) );
  OR U5985 ( .A(n4981), .B(n4980), .Z(n4982) );
  AND U5986 ( .A(n4983), .B(n4982), .Z(n4985) );
  XOR U5987 ( .A(n4986), .B(n4985), .Z(c[2020]) );
  NAND U5988 ( .A(b[0]), .B(a[998]), .Z(n4989) );
  XOR U5989 ( .A(sreg[2021]), .B(n4989), .Z(n4991) );
  NANDN U5990 ( .A(n4984), .B(sreg[2020]), .Z(n4988) );
  OR U5991 ( .A(n4986), .B(n4985), .Z(n4987) );
  AND U5992 ( .A(n4988), .B(n4987), .Z(n4990) );
  XOR U5993 ( .A(n4991), .B(n4990), .Z(c[2021]) );
  NAND U5994 ( .A(b[0]), .B(a[999]), .Z(n4994) );
  XOR U5995 ( .A(sreg[2022]), .B(n4994), .Z(n4996) );
  NANDN U5996 ( .A(n4989), .B(sreg[2021]), .Z(n4993) );
  OR U5997 ( .A(n4991), .B(n4990), .Z(n4992) );
  AND U5998 ( .A(n4993), .B(n4992), .Z(n4995) );
  XOR U5999 ( .A(n4996), .B(n4995), .Z(c[2022]) );
  NAND U6000 ( .A(b[0]), .B(a[1000]), .Z(n4999) );
  XOR U6001 ( .A(sreg[2023]), .B(n4999), .Z(n5001) );
  NANDN U6002 ( .A(n4994), .B(sreg[2022]), .Z(n4998) );
  OR U6003 ( .A(n4996), .B(n4995), .Z(n4997) );
  AND U6004 ( .A(n4998), .B(n4997), .Z(n5000) );
  XOR U6005 ( .A(n5001), .B(n5000), .Z(c[2023]) );
  NAND U6006 ( .A(b[0]), .B(a[1001]), .Z(n5004) );
  XOR U6007 ( .A(sreg[2024]), .B(n5004), .Z(n5006) );
  NANDN U6008 ( .A(n4999), .B(sreg[2023]), .Z(n5003) );
  OR U6009 ( .A(n5001), .B(n5000), .Z(n5002) );
  AND U6010 ( .A(n5003), .B(n5002), .Z(n5005) );
  XOR U6011 ( .A(n5006), .B(n5005), .Z(c[2024]) );
  NAND U6012 ( .A(b[0]), .B(a[1002]), .Z(n5009) );
  XOR U6013 ( .A(sreg[2025]), .B(n5009), .Z(n5011) );
  NANDN U6014 ( .A(n5004), .B(sreg[2024]), .Z(n5008) );
  OR U6015 ( .A(n5006), .B(n5005), .Z(n5007) );
  AND U6016 ( .A(n5008), .B(n5007), .Z(n5010) );
  XOR U6017 ( .A(n5011), .B(n5010), .Z(c[2025]) );
  NAND U6018 ( .A(b[0]), .B(a[1003]), .Z(n5014) );
  XOR U6019 ( .A(sreg[2026]), .B(n5014), .Z(n5016) );
  NANDN U6020 ( .A(n5009), .B(sreg[2025]), .Z(n5013) );
  OR U6021 ( .A(n5011), .B(n5010), .Z(n5012) );
  AND U6022 ( .A(n5013), .B(n5012), .Z(n5015) );
  XOR U6023 ( .A(n5016), .B(n5015), .Z(c[2026]) );
  NAND U6024 ( .A(b[0]), .B(a[1004]), .Z(n5019) );
  XOR U6025 ( .A(sreg[2027]), .B(n5019), .Z(n5021) );
  NANDN U6026 ( .A(n5014), .B(sreg[2026]), .Z(n5018) );
  OR U6027 ( .A(n5016), .B(n5015), .Z(n5017) );
  AND U6028 ( .A(n5018), .B(n5017), .Z(n5020) );
  XOR U6029 ( .A(n5021), .B(n5020), .Z(c[2027]) );
  NAND U6030 ( .A(b[0]), .B(a[1005]), .Z(n5024) );
  XOR U6031 ( .A(sreg[2028]), .B(n5024), .Z(n5026) );
  NANDN U6032 ( .A(n5019), .B(sreg[2027]), .Z(n5023) );
  OR U6033 ( .A(n5021), .B(n5020), .Z(n5022) );
  AND U6034 ( .A(n5023), .B(n5022), .Z(n5025) );
  XOR U6035 ( .A(n5026), .B(n5025), .Z(c[2028]) );
  NAND U6036 ( .A(b[0]), .B(a[1006]), .Z(n5029) );
  XOR U6037 ( .A(sreg[2029]), .B(n5029), .Z(n5031) );
  NANDN U6038 ( .A(n5024), .B(sreg[2028]), .Z(n5028) );
  OR U6039 ( .A(n5026), .B(n5025), .Z(n5027) );
  AND U6040 ( .A(n5028), .B(n5027), .Z(n5030) );
  XOR U6041 ( .A(n5031), .B(n5030), .Z(c[2029]) );
  NAND U6042 ( .A(b[0]), .B(a[1007]), .Z(n5034) );
  XOR U6043 ( .A(sreg[2030]), .B(n5034), .Z(n5036) );
  NANDN U6044 ( .A(n5029), .B(sreg[2029]), .Z(n5033) );
  OR U6045 ( .A(n5031), .B(n5030), .Z(n5032) );
  AND U6046 ( .A(n5033), .B(n5032), .Z(n5035) );
  XOR U6047 ( .A(n5036), .B(n5035), .Z(c[2030]) );
  NAND U6048 ( .A(b[0]), .B(a[1008]), .Z(n5039) );
  XOR U6049 ( .A(sreg[2031]), .B(n5039), .Z(n5041) );
  NANDN U6050 ( .A(n5034), .B(sreg[2030]), .Z(n5038) );
  OR U6051 ( .A(n5036), .B(n5035), .Z(n5037) );
  AND U6052 ( .A(n5038), .B(n5037), .Z(n5040) );
  XOR U6053 ( .A(n5041), .B(n5040), .Z(c[2031]) );
  NAND U6054 ( .A(b[0]), .B(a[1009]), .Z(n5044) );
  XOR U6055 ( .A(sreg[2032]), .B(n5044), .Z(n5046) );
  NANDN U6056 ( .A(n5039), .B(sreg[2031]), .Z(n5043) );
  OR U6057 ( .A(n5041), .B(n5040), .Z(n5042) );
  AND U6058 ( .A(n5043), .B(n5042), .Z(n5045) );
  XOR U6059 ( .A(n5046), .B(n5045), .Z(c[2032]) );
  NAND U6060 ( .A(b[0]), .B(a[1010]), .Z(n5049) );
  XOR U6061 ( .A(sreg[2033]), .B(n5049), .Z(n5051) );
  NANDN U6062 ( .A(n5044), .B(sreg[2032]), .Z(n5048) );
  OR U6063 ( .A(n5046), .B(n5045), .Z(n5047) );
  AND U6064 ( .A(n5048), .B(n5047), .Z(n5050) );
  XOR U6065 ( .A(n5051), .B(n5050), .Z(c[2033]) );
  NAND U6066 ( .A(b[0]), .B(a[1011]), .Z(n5054) );
  XOR U6067 ( .A(sreg[2034]), .B(n5054), .Z(n5056) );
  NANDN U6068 ( .A(n5049), .B(sreg[2033]), .Z(n5053) );
  OR U6069 ( .A(n5051), .B(n5050), .Z(n5052) );
  AND U6070 ( .A(n5053), .B(n5052), .Z(n5055) );
  XOR U6071 ( .A(n5056), .B(n5055), .Z(c[2034]) );
  NAND U6072 ( .A(b[0]), .B(a[1012]), .Z(n5059) );
  XOR U6073 ( .A(sreg[2035]), .B(n5059), .Z(n5061) );
  NANDN U6074 ( .A(n5054), .B(sreg[2034]), .Z(n5058) );
  OR U6075 ( .A(n5056), .B(n5055), .Z(n5057) );
  AND U6076 ( .A(n5058), .B(n5057), .Z(n5060) );
  XOR U6077 ( .A(n5061), .B(n5060), .Z(c[2035]) );
  NAND U6078 ( .A(b[0]), .B(a[1013]), .Z(n5064) );
  XOR U6079 ( .A(sreg[2036]), .B(n5064), .Z(n5066) );
  NANDN U6080 ( .A(n5059), .B(sreg[2035]), .Z(n5063) );
  OR U6081 ( .A(n5061), .B(n5060), .Z(n5062) );
  AND U6082 ( .A(n5063), .B(n5062), .Z(n5065) );
  XOR U6083 ( .A(n5066), .B(n5065), .Z(c[2036]) );
  NAND U6084 ( .A(b[0]), .B(a[1014]), .Z(n5069) );
  XOR U6085 ( .A(sreg[2037]), .B(n5069), .Z(n5071) );
  NANDN U6086 ( .A(n5064), .B(sreg[2036]), .Z(n5068) );
  OR U6087 ( .A(n5066), .B(n5065), .Z(n5067) );
  AND U6088 ( .A(n5068), .B(n5067), .Z(n5070) );
  XOR U6089 ( .A(n5071), .B(n5070), .Z(c[2037]) );
  NAND U6090 ( .A(b[0]), .B(a[1015]), .Z(n5074) );
  XOR U6091 ( .A(sreg[2038]), .B(n5074), .Z(n5076) );
  NANDN U6092 ( .A(n5069), .B(sreg[2037]), .Z(n5073) );
  OR U6093 ( .A(n5071), .B(n5070), .Z(n5072) );
  AND U6094 ( .A(n5073), .B(n5072), .Z(n5075) );
  XOR U6095 ( .A(n5076), .B(n5075), .Z(c[2038]) );
  NAND U6096 ( .A(b[0]), .B(a[1016]), .Z(n5079) );
  XOR U6097 ( .A(sreg[2039]), .B(n5079), .Z(n5081) );
  NANDN U6098 ( .A(n5074), .B(sreg[2038]), .Z(n5078) );
  OR U6099 ( .A(n5076), .B(n5075), .Z(n5077) );
  AND U6100 ( .A(n5078), .B(n5077), .Z(n5080) );
  XOR U6101 ( .A(n5081), .B(n5080), .Z(c[2039]) );
  NAND U6102 ( .A(b[0]), .B(a[1017]), .Z(n5084) );
  XOR U6103 ( .A(sreg[2040]), .B(n5084), .Z(n5086) );
  NANDN U6104 ( .A(n5079), .B(sreg[2039]), .Z(n5083) );
  OR U6105 ( .A(n5081), .B(n5080), .Z(n5082) );
  AND U6106 ( .A(n5083), .B(n5082), .Z(n5085) );
  XOR U6107 ( .A(n5086), .B(n5085), .Z(c[2040]) );
  NAND U6108 ( .A(b[0]), .B(a[1018]), .Z(n5089) );
  XOR U6109 ( .A(sreg[2041]), .B(n5089), .Z(n5091) );
  NANDN U6110 ( .A(n5084), .B(sreg[2040]), .Z(n5088) );
  OR U6111 ( .A(n5086), .B(n5085), .Z(n5087) );
  AND U6112 ( .A(n5088), .B(n5087), .Z(n5090) );
  XOR U6113 ( .A(n5091), .B(n5090), .Z(c[2041]) );
  NAND U6114 ( .A(b[0]), .B(a[1019]), .Z(n5094) );
  XOR U6115 ( .A(sreg[2042]), .B(n5094), .Z(n5096) );
  NANDN U6116 ( .A(n5089), .B(sreg[2041]), .Z(n5093) );
  OR U6117 ( .A(n5091), .B(n5090), .Z(n5092) );
  AND U6118 ( .A(n5093), .B(n5092), .Z(n5095) );
  XOR U6119 ( .A(n5096), .B(n5095), .Z(c[2042]) );
  NAND U6120 ( .A(b[0]), .B(a[1020]), .Z(n5099) );
  XOR U6121 ( .A(sreg[2043]), .B(n5099), .Z(n5101) );
  NANDN U6122 ( .A(n5094), .B(sreg[2042]), .Z(n5098) );
  OR U6123 ( .A(n5096), .B(n5095), .Z(n5097) );
  AND U6124 ( .A(n5098), .B(n5097), .Z(n5100) );
  XOR U6125 ( .A(n5101), .B(n5100), .Z(c[2043]) );
  NAND U6126 ( .A(b[0]), .B(a[1021]), .Z(n5104) );
  XOR U6127 ( .A(sreg[2044]), .B(n5104), .Z(n5106) );
  NANDN U6128 ( .A(n5099), .B(sreg[2043]), .Z(n5103) );
  OR U6129 ( .A(n5101), .B(n5100), .Z(n5102) );
  AND U6130 ( .A(n5103), .B(n5102), .Z(n5105) );
  XOR U6131 ( .A(n5106), .B(n5105), .Z(c[2044]) );
  NAND U6132 ( .A(b[0]), .B(a[1022]), .Z(n5109) );
  XOR U6133 ( .A(sreg[2045]), .B(n5109), .Z(n5111) );
  NANDN U6134 ( .A(n5104), .B(sreg[2044]), .Z(n5108) );
  OR U6135 ( .A(n5106), .B(n5105), .Z(n5107) );
  AND U6136 ( .A(n5108), .B(n5107), .Z(n5110) );
  XOR U6137 ( .A(n5111), .B(n5110), .Z(c[2045]) );
  NANDN U6138 ( .A(n5109), .B(sreg[2045]), .Z(n5113) );
  OR U6139 ( .A(n5111), .B(n5110), .Z(n5112) );
  NAND U6140 ( .A(n5113), .B(n5112), .Z(n5115) );
  NAND U6141 ( .A(b[0]), .B(a[1023]), .Z(n5114) );
  XOR U6142 ( .A(sreg[2046]), .B(n5114), .Z(n5116) );
  XNOR U6143 ( .A(n5115), .B(n5116), .Z(c[2046]) );
  NANDN U6144 ( .A(n5114), .B(sreg[2046]), .Z(n5118) );
  NANDN U6145 ( .A(n5116), .B(n5115), .Z(n5117) );
  NAND U6146 ( .A(n5118), .B(n5117), .Z(c[2047]) );
endmodule

