
module Shifter ( value, shift_amount, shift_func, c_shift );
  input [31:0] value;
  input [4:0] shift_amount;
  input [1:0] shift_func;
  output [31:0] c_shift;
  wire   N75, \sll_27/ML_int[5][16] , \sll_27/ML_int[5][17] ,
         \sll_27/ML_int[5][18] , \sll_27/ML_int[5][19] ,
         \sll_27/ML_int[5][20] , \sll_27/ML_int[5][21] ,
         \sll_27/ML_int[5][22] , \sll_27/ML_int[5][23] ,
         \sll_27/ML_int[5][24] , \sll_27/ML_int[5][25] ,
         \sll_27/ML_int[5][26] , \sll_27/ML_int[5][27] ,
         \sll_27/ML_int[5][28] , \sll_27/ML_int[5][29] ,
         \sll_27/ML_int[5][30] , \sll_27/ML_int[5][31] , \sll_27/ML_int[4][0] ,
         \sll_27/ML_int[4][1] , \sll_27/ML_int[4][2] , \sll_27/ML_int[4][3] ,
         \sll_27/ML_int[4][4] , \sll_27/ML_int[4][5] , \sll_27/ML_int[4][6] ,
         \sll_27/ML_int[4][7] , \sll_27/ML_int[4][8] , \sll_27/ML_int[4][9] ,
         \sll_27/ML_int[4][10] , \sll_27/ML_int[4][11] ,
         \sll_27/ML_int[4][12] , \sll_27/ML_int[4][13] ,
         \sll_27/ML_int[4][14] , \sll_27/ML_int[4][15] ,
         \sll_27/ML_int[4][16] , \sll_27/ML_int[4][17] ,
         \sll_27/ML_int[4][18] , \sll_27/ML_int[4][19] ,
         \sll_27/ML_int[4][20] , \sll_27/ML_int[4][21] ,
         \sll_27/ML_int[4][22] , \sll_27/ML_int[4][23] ,
         \sll_27/ML_int[4][24] , \sll_27/ML_int[4][25] ,
         \sll_27/ML_int[4][26] , \sll_27/ML_int[4][27] ,
         \sll_27/ML_int[4][28] , \sll_27/ML_int[4][29] ,
         \sll_27/ML_int[4][30] , \sll_27/ML_int[4][31] , \sll_27/ML_int[3][0] ,
         \sll_27/ML_int[3][1] , \sll_27/ML_int[3][2] , \sll_27/ML_int[3][3] ,
         \sll_27/ML_int[3][4] , \sll_27/ML_int[3][5] , \sll_27/ML_int[3][6] ,
         \sll_27/ML_int[3][7] , \sll_27/ML_int[3][8] , \sll_27/ML_int[3][9] ,
         \sll_27/ML_int[3][10] , \sll_27/ML_int[3][11] ,
         \sll_27/ML_int[3][12] , \sll_27/ML_int[3][13] ,
         \sll_27/ML_int[3][14] , \sll_27/ML_int[3][15] ,
         \sll_27/ML_int[3][16] , \sll_27/ML_int[3][17] ,
         \sll_27/ML_int[3][18] , \sll_27/ML_int[3][19] ,
         \sll_27/ML_int[3][20] , \sll_27/ML_int[3][21] ,
         \sll_27/ML_int[3][22] , \sll_27/ML_int[3][23] ,
         \sll_27/ML_int[3][24] , \sll_27/ML_int[3][25] ,
         \sll_27/ML_int[3][26] , \sll_27/ML_int[3][27] ,
         \sll_27/ML_int[3][28] , \sll_27/ML_int[3][29] ,
         \sll_27/ML_int[3][30] , \sll_27/ML_int[3][31] , \sll_27/ML_int[2][0] ,
         \sll_27/ML_int[2][1] , \sll_27/ML_int[2][2] , \sll_27/ML_int[2][3] ,
         \sll_27/ML_int[2][4] , \sll_27/ML_int[2][5] , \sll_27/ML_int[2][6] ,
         \sll_27/ML_int[2][7] , \sll_27/ML_int[2][8] , \sll_27/ML_int[2][9] ,
         \sll_27/ML_int[2][10] , \sll_27/ML_int[2][11] ,
         \sll_27/ML_int[2][12] , \sll_27/ML_int[2][13] ,
         \sll_27/ML_int[2][14] , \sll_27/ML_int[2][15] ,
         \sll_27/ML_int[2][16] , \sll_27/ML_int[2][17] ,
         \sll_27/ML_int[2][18] , \sll_27/ML_int[2][19] ,
         \sll_27/ML_int[2][20] , \sll_27/ML_int[2][21] ,
         \sll_27/ML_int[2][22] , \sll_27/ML_int[2][23] ,
         \sll_27/ML_int[2][24] , \sll_27/ML_int[2][25] ,
         \sll_27/ML_int[2][26] , \sll_27/ML_int[2][27] ,
         \sll_27/ML_int[2][28] , \sll_27/ML_int[2][29] ,
         \sll_27/ML_int[2][30] , \sll_27/ML_int[2][31] , \sll_27/ML_int[1][0] ,
         \sll_27/ML_int[1][1] , \sll_27/ML_int[1][2] , \sll_27/ML_int[1][3] ,
         \sll_27/ML_int[1][4] , \sll_27/ML_int[1][5] , \sll_27/ML_int[1][6] ,
         \sll_27/ML_int[1][7] , \sll_27/ML_int[1][8] , \sll_27/ML_int[1][9] ,
         \sll_27/ML_int[1][10] , \sll_27/ML_int[1][11] ,
         \sll_27/ML_int[1][12] , \sll_27/ML_int[1][13] ,
         \sll_27/ML_int[1][14] , \sll_27/ML_int[1][15] ,
         \sll_27/ML_int[1][16] , \sll_27/ML_int[1][17] ,
         \sll_27/ML_int[1][18] , \sll_27/ML_int[1][19] ,
         \sll_27/ML_int[1][20] , \sll_27/ML_int[1][21] ,
         \sll_27/ML_int[1][22] , \sll_27/ML_int[1][23] ,
         \sll_27/ML_int[1][24] , \sll_27/ML_int[1][25] ,
         \sll_27/ML_int[1][26] , \sll_27/ML_int[1][27] ,
         \sll_27/ML_int[1][28] , \sll_27/ML_int[1][29] ,
         \sll_27/ML_int[1][30] , \sll_27/ML_int[1][31] , n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067;
  assign N75 = value[31];

  MUX \sll_27/M1_0_1  ( .IN0(value[1]), .IN1(value[0]), .SEL(shift_amount[0]), 
        .F(\sll_27/ML_int[1][1] ) );
  MUX \sll_27/M1_0_2  ( .IN0(value[2]), .IN1(value[1]), .SEL(shift_amount[0]), 
        .F(\sll_27/ML_int[1][2] ) );
  MUX \sll_27/M1_0_3  ( .IN0(value[3]), .IN1(value[2]), .SEL(shift_amount[0]), 
        .F(\sll_27/ML_int[1][3] ) );
  MUX \sll_27/M1_0_4  ( .IN0(value[4]), .IN1(value[3]), .SEL(shift_amount[0]), 
        .F(\sll_27/ML_int[1][4] ) );
  MUX \sll_27/M1_0_5  ( .IN0(value[5]), .IN1(value[4]), .SEL(shift_amount[0]), 
        .F(\sll_27/ML_int[1][5] ) );
  MUX \sll_27/M1_0_6  ( .IN0(value[6]), .IN1(value[5]), .SEL(shift_amount[0]), 
        .F(\sll_27/ML_int[1][6] ) );
  MUX \sll_27/M1_0_7  ( .IN0(value[7]), .IN1(value[6]), .SEL(shift_amount[0]), 
        .F(\sll_27/ML_int[1][7] ) );
  MUX \sll_27/M1_0_8  ( .IN0(value[8]), .IN1(value[7]), .SEL(shift_amount[0]), 
        .F(\sll_27/ML_int[1][8] ) );
  MUX \sll_27/M1_0_9  ( .IN0(value[9]), .IN1(value[8]), .SEL(shift_amount[0]), 
        .F(\sll_27/ML_int[1][9] ) );
  MUX \sll_27/M1_0_10  ( .IN0(value[10]), .IN1(value[9]), .SEL(shift_amount[0]), .F(\sll_27/ML_int[1][10] ) );
  MUX \sll_27/M1_0_11  ( .IN0(value[11]), .IN1(value[10]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][11] ) );
  MUX \sll_27/M1_0_12  ( .IN0(value[12]), .IN1(value[11]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][12] ) );
  MUX \sll_27/M1_0_13  ( .IN0(value[13]), .IN1(value[12]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][13] ) );
  MUX \sll_27/M1_0_14  ( .IN0(value[14]), .IN1(value[13]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][14] ) );
  MUX \sll_27/M1_0_15  ( .IN0(value[15]), .IN1(value[14]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][15] ) );
  MUX \sll_27/M1_0_16  ( .IN0(value[16]), .IN1(value[15]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][16] ) );
  MUX \sll_27/M1_0_17  ( .IN0(value[17]), .IN1(value[16]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][17] ) );
  MUX \sll_27/M1_0_18  ( .IN0(value[18]), .IN1(value[17]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][18] ) );
  MUX \sll_27/M1_0_19  ( .IN0(value[19]), .IN1(value[18]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][19] ) );
  MUX \sll_27/M1_0_20  ( .IN0(value[20]), .IN1(value[19]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][20] ) );
  MUX \sll_27/M1_0_21  ( .IN0(value[21]), .IN1(value[20]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][21] ) );
  MUX \sll_27/M1_0_22  ( .IN0(value[22]), .IN1(value[21]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][22] ) );
  MUX \sll_27/M1_0_23  ( .IN0(value[23]), .IN1(value[22]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][23] ) );
  MUX \sll_27/M1_0_24  ( .IN0(value[24]), .IN1(value[23]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][24] ) );
  MUX \sll_27/M1_0_25  ( .IN0(value[25]), .IN1(value[24]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][25] ) );
  MUX \sll_27/M1_0_26  ( .IN0(value[26]), .IN1(value[25]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][26] ) );
  MUX \sll_27/M1_0_27  ( .IN0(value[27]), .IN1(value[26]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][27] ) );
  MUX \sll_27/M1_0_28  ( .IN0(value[28]), .IN1(value[27]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][28] ) );
  MUX \sll_27/M1_0_29  ( .IN0(value[29]), .IN1(value[28]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][29] ) );
  MUX \sll_27/M1_0_30  ( .IN0(value[30]), .IN1(value[29]), .SEL(
        shift_amount[0]), .F(\sll_27/ML_int[1][30] ) );
  MUX \sll_27/M1_0_31  ( .IN0(N75), .IN1(value[30]), .SEL(shift_amount[0]), 
        .F(\sll_27/ML_int[1][31] ) );
  MUX \sll_27/M1_1_2  ( .IN0(\sll_27/ML_int[1][2] ), .IN1(
        \sll_27/ML_int[1][0] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][2] ) );
  MUX \sll_27/M1_1_3  ( .IN0(\sll_27/ML_int[1][3] ), .IN1(
        \sll_27/ML_int[1][1] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][3] ) );
  MUX \sll_27/M1_1_4  ( .IN0(\sll_27/ML_int[1][4] ), .IN1(
        \sll_27/ML_int[1][2] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][4] ) );
  MUX \sll_27/M1_1_5  ( .IN0(\sll_27/ML_int[1][5] ), .IN1(
        \sll_27/ML_int[1][3] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][5] ) );
  MUX \sll_27/M1_1_6  ( .IN0(\sll_27/ML_int[1][6] ), .IN1(
        \sll_27/ML_int[1][4] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][6] ) );
  MUX \sll_27/M1_1_7  ( .IN0(\sll_27/ML_int[1][7] ), .IN1(
        \sll_27/ML_int[1][5] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][7] ) );
  MUX \sll_27/M1_1_8  ( .IN0(\sll_27/ML_int[1][8] ), .IN1(
        \sll_27/ML_int[1][6] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][8] ) );
  MUX \sll_27/M1_1_9  ( .IN0(\sll_27/ML_int[1][9] ), .IN1(
        \sll_27/ML_int[1][7] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][9] ) );
  MUX \sll_27/M1_1_10  ( .IN0(\sll_27/ML_int[1][10] ), .IN1(
        \sll_27/ML_int[1][8] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][10] ) );
  MUX \sll_27/M1_1_11  ( .IN0(\sll_27/ML_int[1][11] ), .IN1(
        \sll_27/ML_int[1][9] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][11] ) );
  MUX \sll_27/M1_1_12  ( .IN0(\sll_27/ML_int[1][12] ), .IN1(
        \sll_27/ML_int[1][10] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][12] ) );
  MUX \sll_27/M1_1_13  ( .IN0(\sll_27/ML_int[1][13] ), .IN1(
        \sll_27/ML_int[1][11] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][13] ) );
  MUX \sll_27/M1_1_14  ( .IN0(\sll_27/ML_int[1][14] ), .IN1(
        \sll_27/ML_int[1][12] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][14] ) );
  MUX \sll_27/M1_1_15  ( .IN0(\sll_27/ML_int[1][15] ), .IN1(
        \sll_27/ML_int[1][13] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][15] ) );
  MUX \sll_27/M1_1_16  ( .IN0(\sll_27/ML_int[1][16] ), .IN1(
        \sll_27/ML_int[1][14] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][16] ) );
  MUX \sll_27/M1_1_17  ( .IN0(\sll_27/ML_int[1][17] ), .IN1(
        \sll_27/ML_int[1][15] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][17] ) );
  MUX \sll_27/M1_1_18  ( .IN0(\sll_27/ML_int[1][18] ), .IN1(
        \sll_27/ML_int[1][16] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][18] ) );
  MUX \sll_27/M1_1_19  ( .IN0(\sll_27/ML_int[1][19] ), .IN1(
        \sll_27/ML_int[1][17] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][19] ) );
  MUX \sll_27/M1_1_20  ( .IN0(\sll_27/ML_int[1][20] ), .IN1(
        \sll_27/ML_int[1][18] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][20] ) );
  MUX \sll_27/M1_1_21  ( .IN0(\sll_27/ML_int[1][21] ), .IN1(
        \sll_27/ML_int[1][19] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][21] ) );
  MUX \sll_27/M1_1_22  ( .IN0(\sll_27/ML_int[1][22] ), .IN1(
        \sll_27/ML_int[1][20] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][22] ) );
  MUX \sll_27/M1_1_23  ( .IN0(\sll_27/ML_int[1][23] ), .IN1(
        \sll_27/ML_int[1][21] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][23] ) );
  MUX \sll_27/M1_1_24  ( .IN0(\sll_27/ML_int[1][24] ), .IN1(
        \sll_27/ML_int[1][22] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][24] ) );
  MUX \sll_27/M1_1_25  ( .IN0(\sll_27/ML_int[1][25] ), .IN1(
        \sll_27/ML_int[1][23] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][25] ) );
  MUX \sll_27/M1_1_26  ( .IN0(\sll_27/ML_int[1][26] ), .IN1(
        \sll_27/ML_int[1][24] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][26] ) );
  MUX \sll_27/M1_1_27  ( .IN0(\sll_27/ML_int[1][27] ), .IN1(
        \sll_27/ML_int[1][25] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][27] ) );
  MUX \sll_27/M1_1_28  ( .IN0(\sll_27/ML_int[1][28] ), .IN1(
        \sll_27/ML_int[1][26] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][28] ) );
  MUX \sll_27/M1_1_29  ( .IN0(\sll_27/ML_int[1][29] ), .IN1(
        \sll_27/ML_int[1][27] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][29] ) );
  MUX \sll_27/M1_1_30  ( .IN0(\sll_27/ML_int[1][30] ), .IN1(
        \sll_27/ML_int[1][28] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][30] ) );
  MUX \sll_27/M1_1_31  ( .IN0(\sll_27/ML_int[1][31] ), .IN1(
        \sll_27/ML_int[1][29] ), .SEL(shift_amount[1]), .F(
        \sll_27/ML_int[2][31] ) );
  MUX \sll_27/M1_2_4  ( .IN0(\sll_27/ML_int[2][4] ), .IN1(
        \sll_27/ML_int[2][0] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][4] ) );
  MUX \sll_27/M1_2_5  ( .IN0(\sll_27/ML_int[2][5] ), .IN1(
        \sll_27/ML_int[2][1] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][5] ) );
  MUX \sll_27/M1_2_6  ( .IN0(\sll_27/ML_int[2][6] ), .IN1(
        \sll_27/ML_int[2][2] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][6] ) );
  MUX \sll_27/M1_2_7  ( .IN0(\sll_27/ML_int[2][7] ), .IN1(
        \sll_27/ML_int[2][3] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][7] ) );
  MUX \sll_27/M1_2_8  ( .IN0(\sll_27/ML_int[2][8] ), .IN1(
        \sll_27/ML_int[2][4] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][8] ) );
  MUX \sll_27/M1_2_9  ( .IN0(\sll_27/ML_int[2][9] ), .IN1(
        \sll_27/ML_int[2][5] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][9] ) );
  MUX \sll_27/M1_2_10  ( .IN0(\sll_27/ML_int[2][10] ), .IN1(
        \sll_27/ML_int[2][6] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][10] ) );
  MUX \sll_27/M1_2_11  ( .IN0(\sll_27/ML_int[2][11] ), .IN1(
        \sll_27/ML_int[2][7] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][11] ) );
  MUX \sll_27/M1_2_12  ( .IN0(\sll_27/ML_int[2][12] ), .IN1(
        \sll_27/ML_int[2][8] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][12] ) );
  MUX \sll_27/M1_2_13  ( .IN0(\sll_27/ML_int[2][13] ), .IN1(
        \sll_27/ML_int[2][9] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][13] ) );
  MUX \sll_27/M1_2_14  ( .IN0(\sll_27/ML_int[2][14] ), .IN1(
        \sll_27/ML_int[2][10] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][14] ) );
  MUX \sll_27/M1_2_15  ( .IN0(\sll_27/ML_int[2][15] ), .IN1(
        \sll_27/ML_int[2][11] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][15] ) );
  MUX \sll_27/M1_2_16  ( .IN0(\sll_27/ML_int[2][16] ), .IN1(
        \sll_27/ML_int[2][12] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][16] ) );
  MUX \sll_27/M1_2_17  ( .IN0(\sll_27/ML_int[2][17] ), .IN1(
        \sll_27/ML_int[2][13] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][17] ) );
  MUX \sll_27/M1_2_18  ( .IN0(\sll_27/ML_int[2][18] ), .IN1(
        \sll_27/ML_int[2][14] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][18] ) );
  MUX \sll_27/M1_2_19  ( .IN0(\sll_27/ML_int[2][19] ), .IN1(
        \sll_27/ML_int[2][15] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][19] ) );
  MUX \sll_27/M1_2_20  ( .IN0(\sll_27/ML_int[2][20] ), .IN1(
        \sll_27/ML_int[2][16] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][20] ) );
  MUX \sll_27/M1_2_21  ( .IN0(\sll_27/ML_int[2][21] ), .IN1(
        \sll_27/ML_int[2][17] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][21] ) );
  MUX \sll_27/M1_2_22  ( .IN0(\sll_27/ML_int[2][22] ), .IN1(
        \sll_27/ML_int[2][18] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][22] ) );
  MUX \sll_27/M1_2_23  ( .IN0(\sll_27/ML_int[2][23] ), .IN1(
        \sll_27/ML_int[2][19] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][23] ) );
  MUX \sll_27/M1_2_24  ( .IN0(\sll_27/ML_int[2][24] ), .IN1(
        \sll_27/ML_int[2][20] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][24] ) );
  MUX \sll_27/M1_2_25  ( .IN0(\sll_27/ML_int[2][25] ), .IN1(
        \sll_27/ML_int[2][21] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][25] ) );
  MUX \sll_27/M1_2_26  ( .IN0(\sll_27/ML_int[2][26] ), .IN1(
        \sll_27/ML_int[2][22] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][26] ) );
  MUX \sll_27/M1_2_27  ( .IN0(\sll_27/ML_int[2][27] ), .IN1(
        \sll_27/ML_int[2][23] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][27] ) );
  MUX \sll_27/M1_2_28  ( .IN0(\sll_27/ML_int[2][28] ), .IN1(
        \sll_27/ML_int[2][24] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][28] ) );
  MUX \sll_27/M1_2_29  ( .IN0(\sll_27/ML_int[2][29] ), .IN1(
        \sll_27/ML_int[2][25] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][29] ) );
  MUX \sll_27/M1_2_30  ( .IN0(\sll_27/ML_int[2][30] ), .IN1(
        \sll_27/ML_int[2][26] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][30] ) );
  MUX \sll_27/M1_2_31  ( .IN0(\sll_27/ML_int[2][31] ), .IN1(
        \sll_27/ML_int[2][27] ), .SEL(shift_amount[2]), .F(
        \sll_27/ML_int[3][31] ) );
  MUX \sll_27/M1_3_8  ( .IN0(\sll_27/ML_int[3][8] ), .IN1(
        \sll_27/ML_int[3][0] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][8] ) );
  MUX \sll_27/M1_3_9  ( .IN0(\sll_27/ML_int[3][9] ), .IN1(
        \sll_27/ML_int[3][1] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][9] ) );
  MUX \sll_27/M1_3_10  ( .IN0(\sll_27/ML_int[3][10] ), .IN1(
        \sll_27/ML_int[3][2] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][10] ) );
  MUX \sll_27/M1_3_11  ( .IN0(\sll_27/ML_int[3][11] ), .IN1(
        \sll_27/ML_int[3][3] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][11] ) );
  MUX \sll_27/M1_3_12  ( .IN0(\sll_27/ML_int[3][12] ), .IN1(
        \sll_27/ML_int[3][4] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][12] ) );
  MUX \sll_27/M1_3_13  ( .IN0(\sll_27/ML_int[3][13] ), .IN1(
        \sll_27/ML_int[3][5] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][13] ) );
  MUX \sll_27/M1_3_14  ( .IN0(\sll_27/ML_int[3][14] ), .IN1(
        \sll_27/ML_int[3][6] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][14] ) );
  MUX \sll_27/M1_3_15  ( .IN0(\sll_27/ML_int[3][15] ), .IN1(
        \sll_27/ML_int[3][7] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][15] ) );
  MUX \sll_27/M1_3_16  ( .IN0(\sll_27/ML_int[3][16] ), .IN1(
        \sll_27/ML_int[3][8] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][16] ) );
  MUX \sll_27/M1_3_17  ( .IN0(\sll_27/ML_int[3][17] ), .IN1(
        \sll_27/ML_int[3][9] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][17] ) );
  MUX \sll_27/M1_3_18  ( .IN0(\sll_27/ML_int[3][18] ), .IN1(
        \sll_27/ML_int[3][10] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][18] ) );
  MUX \sll_27/M1_3_19  ( .IN0(\sll_27/ML_int[3][19] ), .IN1(
        \sll_27/ML_int[3][11] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][19] ) );
  MUX \sll_27/M1_3_20  ( .IN0(\sll_27/ML_int[3][20] ), .IN1(
        \sll_27/ML_int[3][12] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][20] ) );
  MUX \sll_27/M1_3_21  ( .IN0(\sll_27/ML_int[3][21] ), .IN1(
        \sll_27/ML_int[3][13] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][21] ) );
  MUX \sll_27/M1_3_22  ( .IN0(\sll_27/ML_int[3][22] ), .IN1(
        \sll_27/ML_int[3][14] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][22] ) );
  MUX \sll_27/M1_3_23  ( .IN0(\sll_27/ML_int[3][23] ), .IN1(
        \sll_27/ML_int[3][15] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][23] ) );
  MUX \sll_27/M1_3_24  ( .IN0(\sll_27/ML_int[3][24] ), .IN1(
        \sll_27/ML_int[3][16] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][24] ) );
  MUX \sll_27/M1_3_25  ( .IN0(\sll_27/ML_int[3][25] ), .IN1(
        \sll_27/ML_int[3][17] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][25] ) );
  MUX \sll_27/M1_3_26  ( .IN0(\sll_27/ML_int[3][26] ), .IN1(
        \sll_27/ML_int[3][18] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][26] ) );
  MUX \sll_27/M1_3_27  ( .IN0(\sll_27/ML_int[3][27] ), .IN1(
        \sll_27/ML_int[3][19] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][27] ) );
  MUX \sll_27/M1_3_28  ( .IN0(\sll_27/ML_int[3][28] ), .IN1(
        \sll_27/ML_int[3][20] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][28] ) );
  MUX \sll_27/M1_3_29  ( .IN0(\sll_27/ML_int[3][29] ), .IN1(
        \sll_27/ML_int[3][21] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][29] ) );
  MUX \sll_27/M1_3_30  ( .IN0(\sll_27/ML_int[3][30] ), .IN1(
        \sll_27/ML_int[3][22] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][30] ) );
  MUX \sll_27/M1_3_31  ( .IN0(\sll_27/ML_int[3][31] ), .IN1(
        \sll_27/ML_int[3][23] ), .SEL(shift_amount[3]), .F(
        \sll_27/ML_int[4][31] ) );
  MUX \sll_27/M1_4_16  ( .IN0(\sll_27/ML_int[4][16] ), .IN1(
        \sll_27/ML_int[4][0] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][16] ) );
  MUX \sll_27/M1_4_17  ( .IN0(\sll_27/ML_int[4][17] ), .IN1(
        \sll_27/ML_int[4][1] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][17] ) );
  MUX \sll_27/M1_4_18  ( .IN0(\sll_27/ML_int[4][18] ), .IN1(
        \sll_27/ML_int[4][2] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][18] ) );
  MUX \sll_27/M1_4_19  ( .IN0(\sll_27/ML_int[4][19] ), .IN1(
        \sll_27/ML_int[4][3] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][19] ) );
  MUX \sll_27/M1_4_20  ( .IN0(\sll_27/ML_int[4][20] ), .IN1(
        \sll_27/ML_int[4][4] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][20] ) );
  MUX \sll_27/M1_4_21  ( .IN0(\sll_27/ML_int[4][21] ), .IN1(
        \sll_27/ML_int[4][5] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][21] ) );
  MUX \sll_27/M1_4_22  ( .IN0(\sll_27/ML_int[4][22] ), .IN1(
        \sll_27/ML_int[4][6] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][22] ) );
  MUX \sll_27/M1_4_23  ( .IN0(\sll_27/ML_int[4][23] ), .IN1(
        \sll_27/ML_int[4][7] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][23] ) );
  MUX \sll_27/M1_4_24  ( .IN0(\sll_27/ML_int[4][24] ), .IN1(
        \sll_27/ML_int[4][8] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][24] ) );
  MUX \sll_27/M1_4_25  ( .IN0(\sll_27/ML_int[4][25] ), .IN1(
        \sll_27/ML_int[4][9] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][25] ) );
  MUX \sll_27/M1_4_26  ( .IN0(\sll_27/ML_int[4][26] ), .IN1(
        \sll_27/ML_int[4][10] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][26] ) );
  MUX \sll_27/M1_4_27  ( .IN0(\sll_27/ML_int[4][27] ), .IN1(
        \sll_27/ML_int[4][11] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][27] ) );
  MUX \sll_27/M1_4_28  ( .IN0(\sll_27/ML_int[4][28] ), .IN1(
        \sll_27/ML_int[4][12] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][28] ) );
  MUX \sll_27/M1_4_29  ( .IN0(\sll_27/ML_int[4][29] ), .IN1(
        \sll_27/ML_int[4][13] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][29] ) );
  MUX \sll_27/M1_4_30  ( .IN0(\sll_27/ML_int[4][30] ), .IN1(
        \sll_27/ML_int[4][14] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][30] ) );
  MUX \sll_27/M1_4_31  ( .IN0(\sll_27/ML_int[4][31] ), .IN1(
        \sll_27/ML_int[4][15] ), .SEL(shift_amount[4]), .F(
        \sll_27/ML_int[5][31] ) );
  NAND U173 ( .A(n144), .B(n145), .Z(c_shift[9]) );
  NAND U174 ( .A(n146), .B(\sll_27/ML_int[4][9] ), .Z(n145) );
  AND U175 ( .A(n147), .B(n148), .Z(n144) );
  NAND U176 ( .A(n149), .B(n150), .Z(n148) );
  NAND U177 ( .A(n151), .B(n152), .Z(n149) );
  AND U178 ( .A(n153), .B(n154), .Z(n152) );
  NAND U179 ( .A(n155), .B(n156), .Z(n154) );
  AND U180 ( .A(n157), .B(n158), .Z(n153) );
  OR U181 ( .A(n159), .B(n160), .Z(n158) );
  NANDN U182 ( .A(n161), .B(n162), .Z(n157) );
  AND U183 ( .A(n163), .B(n164), .Z(n151) );
  NAND U184 ( .A(n165), .B(n166), .Z(n164) );
  NAND U185 ( .A(n167), .B(n168), .Z(n163) );
  NAND U186 ( .A(n169), .B(n170), .Z(n147) );
  NAND U187 ( .A(n171), .B(n172), .Z(n169) );
  AND U188 ( .A(n173), .B(n174), .Z(n172) );
  NAND U189 ( .A(n175), .B(n156), .Z(n174) );
  AND U190 ( .A(n176), .B(n177), .Z(n173) );
  OR U191 ( .A(n178), .B(n160), .Z(n177) );
  NANDN U192 ( .A(n179), .B(n162), .Z(n176) );
  AND U193 ( .A(n180), .B(n181), .Z(n171) );
  NAND U194 ( .A(n182), .B(n166), .Z(n181) );
  NAND U195 ( .A(n183), .B(n168), .Z(n180) );
  NAND U196 ( .A(n184), .B(n185), .Z(c_shift[8]) );
  NAND U197 ( .A(n146), .B(\sll_27/ML_int[4][8] ), .Z(n185) );
  AND U198 ( .A(n186), .B(n187), .Z(n184) );
  NAND U199 ( .A(n188), .B(n150), .Z(n187) );
  NAND U200 ( .A(n189), .B(n190), .Z(n188) );
  AND U201 ( .A(n191), .B(n192), .Z(n190) );
  NAND U202 ( .A(n193), .B(n156), .Z(n192) );
  AND U203 ( .A(n194), .B(n195), .Z(n191) );
  OR U204 ( .A(n196), .B(n160), .Z(n195) );
  NANDN U205 ( .A(n197), .B(n162), .Z(n194) );
  AND U206 ( .A(n198), .B(n199), .Z(n189) );
  NAND U207 ( .A(n200), .B(n166), .Z(n199) );
  NAND U208 ( .A(n201), .B(n168), .Z(n198) );
  NAND U209 ( .A(n202), .B(n170), .Z(n186) );
  NAND U210 ( .A(n203), .B(n204), .Z(n202) );
  AND U211 ( .A(n205), .B(n206), .Z(n204) );
  NAND U212 ( .A(n207), .B(n156), .Z(n206) );
  AND U213 ( .A(n208), .B(n209), .Z(n205) );
  OR U214 ( .A(n210), .B(n160), .Z(n209) );
  NANDN U215 ( .A(n211), .B(n162), .Z(n208) );
  AND U216 ( .A(n212), .B(n213), .Z(n203) );
  NAND U217 ( .A(n214), .B(n166), .Z(n213) );
  NAND U218 ( .A(n215), .B(n168), .Z(n212) );
  NAND U219 ( .A(n216), .B(n217), .Z(c_shift[7]) );
  NAND U220 ( .A(n146), .B(\sll_27/ML_int[4][7] ), .Z(n217) );
  AND U221 ( .A(\sll_27/ML_int[3][7] ), .B(n218), .Z(\sll_27/ML_int[4][7] ) );
  AND U222 ( .A(n219), .B(n220), .Z(n216) );
  NAND U223 ( .A(n221), .B(n150), .Z(n220) );
  NAND U224 ( .A(n222), .B(n223), .Z(n221) );
  AND U225 ( .A(n224), .B(n225), .Z(n223) );
  NAND U226 ( .A(n226), .B(n156), .Z(n225) );
  AND U227 ( .A(n227), .B(n228), .Z(n224) );
  OR U228 ( .A(n229), .B(n160), .Z(n228) );
  NANDN U229 ( .A(n230), .B(n162), .Z(n227) );
  AND U230 ( .A(n231), .B(n232), .Z(n222) );
  NAND U231 ( .A(n233), .B(n166), .Z(n232) );
  NANDN U232 ( .A(n234), .B(n168), .Z(n231) );
  NAND U233 ( .A(n235), .B(n170), .Z(n219) );
  NAND U234 ( .A(n236), .B(n237), .Z(n235) );
  AND U235 ( .A(n238), .B(n239), .Z(n237) );
  NAND U236 ( .A(n240), .B(n156), .Z(n239) );
  AND U237 ( .A(n241), .B(n242), .Z(n238) );
  OR U238 ( .A(n243), .B(n160), .Z(n242) );
  NANDN U239 ( .A(n244), .B(n162), .Z(n241) );
  AND U240 ( .A(n245), .B(n246), .Z(n236) );
  NAND U241 ( .A(n247), .B(n166), .Z(n246) );
  NANDN U242 ( .A(n248), .B(n168), .Z(n245) );
  NAND U243 ( .A(n249), .B(n250), .Z(c_shift[6]) );
  NAND U244 ( .A(n146), .B(\sll_27/ML_int[4][6] ), .Z(n250) );
  AND U245 ( .A(\sll_27/ML_int[3][6] ), .B(n218), .Z(\sll_27/ML_int[4][6] ) );
  AND U246 ( .A(n251), .B(n252), .Z(n249) );
  NAND U247 ( .A(n253), .B(n150), .Z(n252) );
  NAND U248 ( .A(n254), .B(n255), .Z(n253) );
  AND U249 ( .A(n256), .B(n257), .Z(n255) );
  NAND U250 ( .A(n258), .B(n156), .Z(n257) );
  AND U251 ( .A(n259), .B(n260), .Z(n256) );
  OR U252 ( .A(n261), .B(n160), .Z(n260) );
  NANDN U253 ( .A(n262), .B(n162), .Z(n259) );
  AND U254 ( .A(n263), .B(n264), .Z(n254) );
  NAND U255 ( .A(n265), .B(n166), .Z(n264) );
  NANDN U256 ( .A(n266), .B(n168), .Z(n263) );
  NAND U257 ( .A(n267), .B(n170), .Z(n251) );
  NAND U258 ( .A(n268), .B(n269), .Z(n267) );
  AND U259 ( .A(n270), .B(n271), .Z(n269) );
  NAND U260 ( .A(n272), .B(n156), .Z(n271) );
  AND U261 ( .A(n273), .B(n274), .Z(n270) );
  OR U262 ( .A(n275), .B(n160), .Z(n274) );
  NANDN U263 ( .A(n276), .B(n162), .Z(n273) );
  AND U264 ( .A(n277), .B(n278), .Z(n268) );
  NAND U265 ( .A(n279), .B(n166), .Z(n278) );
  NANDN U266 ( .A(n280), .B(n168), .Z(n277) );
  NAND U267 ( .A(n281), .B(n282), .Z(c_shift[5]) );
  NAND U268 ( .A(n146), .B(\sll_27/ML_int[4][5] ), .Z(n282) );
  AND U269 ( .A(\sll_27/ML_int[3][5] ), .B(n218), .Z(\sll_27/ML_int[4][5] ) );
  AND U270 ( .A(n283), .B(n284), .Z(n281) );
  NAND U271 ( .A(n285), .B(n150), .Z(n284) );
  NAND U272 ( .A(n286), .B(n287), .Z(n285) );
  AND U273 ( .A(n288), .B(n289), .Z(n287) );
  NAND U274 ( .A(n165), .B(n156), .Z(n289) );
  AND U275 ( .A(n290), .B(n291), .Z(n288) );
  OR U276 ( .A(n292), .B(n160), .Z(n291) );
  NANDN U277 ( .A(n293), .B(n162), .Z(n290) );
  AND U278 ( .A(n294), .B(n295), .Z(n286) );
  NAND U279 ( .A(n167), .B(n166), .Z(n295) );
  NANDN U280 ( .A(n161), .B(n168), .Z(n294) );
  NAND U281 ( .A(n296), .B(n170), .Z(n283) );
  NAND U282 ( .A(n297), .B(n298), .Z(n296) );
  AND U283 ( .A(n299), .B(n300), .Z(n298) );
  NAND U284 ( .A(n182), .B(n156), .Z(n300) );
  AND U285 ( .A(n301), .B(n302), .Z(n299) );
  OR U286 ( .A(n303), .B(n160), .Z(n302) );
  NANDN U287 ( .A(n304), .B(n162), .Z(n301) );
  AND U288 ( .A(n305), .B(n306), .Z(n297) );
  NAND U289 ( .A(n183), .B(n166), .Z(n306) );
  NANDN U290 ( .A(n179), .B(n168), .Z(n305) );
  NAND U291 ( .A(n307), .B(n308), .Z(c_shift[4]) );
  NAND U292 ( .A(n146), .B(\sll_27/ML_int[4][4] ), .Z(n308) );
  AND U293 ( .A(\sll_27/ML_int[3][4] ), .B(n218), .Z(\sll_27/ML_int[4][4] ) );
  AND U294 ( .A(n309), .B(n310), .Z(n307) );
  NAND U295 ( .A(n311), .B(n150), .Z(n310) );
  NAND U296 ( .A(n312), .B(n313), .Z(n311) );
  AND U297 ( .A(n314), .B(n315), .Z(n313) );
  NAND U298 ( .A(n200), .B(n156), .Z(n315) );
  AND U299 ( .A(n316), .B(n317), .Z(n314) );
  OR U300 ( .A(n318), .B(n160), .Z(n317) );
  NANDN U301 ( .A(n319), .B(n162), .Z(n316) );
  AND U302 ( .A(n320), .B(n321), .Z(n312) );
  NAND U303 ( .A(n201), .B(n166), .Z(n321) );
  NANDN U304 ( .A(n197), .B(n168), .Z(n320) );
  NAND U305 ( .A(n322), .B(n170), .Z(n309) );
  NAND U306 ( .A(n323), .B(n324), .Z(n322) );
  AND U307 ( .A(n325), .B(n326), .Z(n324) );
  NAND U308 ( .A(n214), .B(n156), .Z(n326) );
  AND U309 ( .A(n327), .B(n328), .Z(n325) );
  OR U310 ( .A(n329), .B(n160), .Z(n328) );
  NANDN U311 ( .A(n330), .B(n162), .Z(n327) );
  AND U312 ( .A(n331), .B(n332), .Z(n323) );
  NAND U313 ( .A(n215), .B(n166), .Z(n332) );
  NANDN U314 ( .A(n211), .B(n168), .Z(n331) );
  NAND U315 ( .A(n333), .B(n334), .Z(c_shift[3]) );
  NAND U316 ( .A(n146), .B(\sll_27/ML_int[4][3] ), .Z(n334) );
  AND U317 ( .A(\sll_27/ML_int[3][3] ), .B(n218), .Z(\sll_27/ML_int[4][3] ) );
  AND U318 ( .A(\sll_27/ML_int[2][3] ), .B(n335), .Z(\sll_27/ML_int[3][3] ) );
  AND U319 ( .A(n336), .B(n337), .Z(n333) );
  NAND U320 ( .A(n338), .B(n150), .Z(n337) );
  NAND U321 ( .A(n339), .B(n340), .Z(n338) );
  AND U322 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U323 ( .A(n234), .B(n166), .Z(n342) );
  AND U324 ( .A(n343), .B(n344), .Z(n341) );
  OR U325 ( .A(n345), .B(n160), .Z(n344) );
  NANDN U326 ( .A(n230), .B(n168), .Z(n343) );
  AND U327 ( .A(n346), .B(n347), .Z(n230) );
  AND U328 ( .A(n348), .B(n349), .Z(n347) );
  NANDN U329 ( .A(n350), .B(value[7]), .Z(n349) );
  AND U330 ( .A(n351), .B(n352), .Z(n339) );
  NAND U331 ( .A(n353), .B(n162), .Z(n352) );
  NAND U332 ( .A(n354), .B(n355), .Z(n353) );
  AND U333 ( .A(n356), .B(n357), .Z(n355) );
  NANDN U334 ( .A(n350), .B(value[3]), .Z(n357) );
  NAND U335 ( .A(n233), .B(n156), .Z(n351) );
  NAND U336 ( .A(n358), .B(n170), .Z(n336) );
  NAND U337 ( .A(n359), .B(n360), .Z(n358) );
  AND U338 ( .A(n361), .B(n362), .Z(n360) );
  NANDN U339 ( .A(n248), .B(n166), .Z(n362) );
  AND U340 ( .A(n363), .B(n364), .Z(n361) );
  OR U341 ( .A(n365), .B(n160), .Z(n364) );
  NANDN U342 ( .A(n244), .B(n168), .Z(n363) );
  AND U343 ( .A(n346), .B(n366), .Z(n244) );
  AND U344 ( .A(n348), .B(n367), .Z(n366) );
  NANDN U345 ( .A(n368), .B(value[7]), .Z(n367) );
  NAND U346 ( .A(n369), .B(value[8]), .Z(n348) );
  AND U347 ( .A(n370), .B(n371), .Z(n346) );
  NAND U348 ( .A(n372), .B(value[10]), .Z(n371) );
  NAND U349 ( .A(n373), .B(value[9]), .Z(n370) );
  AND U350 ( .A(n374), .B(n375), .Z(n359) );
  NAND U351 ( .A(n376), .B(n162), .Z(n375) );
  NAND U352 ( .A(n354), .B(n377), .Z(n376) );
  AND U353 ( .A(n356), .B(n378), .Z(n377) );
  NANDN U354 ( .A(n368), .B(value[3]), .Z(n378) );
  NAND U355 ( .A(n369), .B(value[4]), .Z(n356) );
  AND U356 ( .A(n379), .B(n380), .Z(n354) );
  NAND U357 ( .A(n372), .B(value[6]), .Z(n380) );
  NAND U358 ( .A(n373), .B(value[5]), .Z(n379) );
  NAND U359 ( .A(n247), .B(n156), .Z(n374) );
  NAND U360 ( .A(n381), .B(n382), .Z(c_shift[31]) );
  NAND U361 ( .A(n383), .B(\sll_27/ML_int[5][31] ), .Z(n382) );
  AND U362 ( .A(n384), .B(n385), .Z(n381) );
  NANDN U363 ( .A(n386), .B(n150), .Z(n385) );
  NANDN U364 ( .A(n387), .B(n388), .Z(n384) );
  AND U365 ( .A(n162), .B(n170), .Z(n388) );
  NAND U366 ( .A(n389), .B(n390), .Z(c_shift[30]) );
  NAND U367 ( .A(n383), .B(\sll_27/ML_int[5][30] ), .Z(n390) );
  AND U368 ( .A(n391), .B(n392), .Z(n389) );
  NAND U369 ( .A(n393), .B(n150), .Z(n392) );
  NAND U370 ( .A(n394), .B(n395), .Z(n393) );
  OR U371 ( .A(n396), .B(shift_amount[4]), .Z(n394) );
  NAND U372 ( .A(n397), .B(n170), .Z(n391) );
  AND U373 ( .A(n398), .B(n162), .Z(n397) );
  NAND U374 ( .A(n399), .B(n400), .Z(c_shift[2]) );
  NAND U375 ( .A(n146), .B(\sll_27/ML_int[4][2] ), .Z(n400) );
  AND U376 ( .A(\sll_27/ML_int[3][2] ), .B(n218), .Z(\sll_27/ML_int[4][2] ) );
  AND U377 ( .A(\sll_27/ML_int[2][2] ), .B(n335), .Z(\sll_27/ML_int[3][2] ) );
  AND U378 ( .A(n401), .B(n402), .Z(n399) );
  NAND U379 ( .A(n403), .B(n150), .Z(n402) );
  NAND U380 ( .A(n404), .B(n405), .Z(n403) );
  AND U381 ( .A(n406), .B(n407), .Z(n405) );
  NANDN U382 ( .A(n266), .B(n166), .Z(n407) );
  AND U383 ( .A(n408), .B(n409), .Z(n406) );
  OR U384 ( .A(n410), .B(n160), .Z(n409) );
  NANDN U385 ( .A(n262), .B(n168), .Z(n408) );
  AND U386 ( .A(n411), .B(n412), .Z(n262) );
  AND U387 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U388 ( .A(n350), .B(value[6]), .Z(n414) );
  AND U389 ( .A(n415), .B(n416), .Z(n404) );
  NAND U390 ( .A(n417), .B(n162), .Z(n416) );
  NAND U391 ( .A(n418), .B(n419), .Z(n417) );
  AND U392 ( .A(n420), .B(n421), .Z(n419) );
  NANDN U393 ( .A(n350), .B(value[2]), .Z(n421) );
  NAND U394 ( .A(n265), .B(n156), .Z(n415) );
  NAND U395 ( .A(n422), .B(n170), .Z(n401) );
  NAND U396 ( .A(n423), .B(n424), .Z(n422) );
  AND U397 ( .A(n425), .B(n426), .Z(n424) );
  NANDN U398 ( .A(n280), .B(n166), .Z(n426) );
  AND U399 ( .A(n427), .B(n428), .Z(n425) );
  OR U400 ( .A(n429), .B(n160), .Z(n428) );
  NANDN U401 ( .A(n276), .B(n168), .Z(n427) );
  AND U402 ( .A(n411), .B(n430), .Z(n276) );
  AND U403 ( .A(n413), .B(n431), .Z(n430) );
  NANDN U404 ( .A(n368), .B(value[6]), .Z(n431) );
  NAND U405 ( .A(n369), .B(value[7]), .Z(n413) );
  AND U406 ( .A(n432), .B(n433), .Z(n411) );
  NAND U407 ( .A(n372), .B(value[9]), .Z(n433) );
  NAND U408 ( .A(n373), .B(value[8]), .Z(n432) );
  AND U409 ( .A(n434), .B(n435), .Z(n423) );
  NAND U410 ( .A(n436), .B(n162), .Z(n435) );
  NAND U411 ( .A(n418), .B(n437), .Z(n436) );
  AND U412 ( .A(n420), .B(n438), .Z(n437) );
  NANDN U413 ( .A(n368), .B(value[2]), .Z(n438) );
  NAND U414 ( .A(n369), .B(value[3]), .Z(n420) );
  AND U415 ( .A(n439), .B(n440), .Z(n418) );
  NAND U416 ( .A(n372), .B(value[5]), .Z(n440) );
  NAND U417 ( .A(n373), .B(value[4]), .Z(n439) );
  NAND U418 ( .A(n279), .B(n156), .Z(n434) );
  NAND U419 ( .A(n441), .B(n442), .Z(c_shift[29]) );
  NAND U420 ( .A(n383), .B(\sll_27/ML_int[5][29] ), .Z(n442) );
  AND U421 ( .A(n443), .B(n444), .Z(n441) );
  NAND U422 ( .A(n445), .B(n150), .Z(n444) );
  NAND U423 ( .A(n446), .B(n395), .Z(n445) );
  OR U424 ( .A(n447), .B(shift_amount[4]), .Z(n446) );
  NAND U425 ( .A(n448), .B(n170), .Z(n443) );
  AND U426 ( .A(n449), .B(n162), .Z(n448) );
  NAND U427 ( .A(n450), .B(n451), .Z(c_shift[28]) );
  NAND U428 ( .A(n383), .B(\sll_27/ML_int[5][28] ), .Z(n451) );
  AND U429 ( .A(n452), .B(n453), .Z(n450) );
  NAND U430 ( .A(n454), .B(n150), .Z(n453) );
  NAND U431 ( .A(n455), .B(n395), .Z(n454) );
  OR U432 ( .A(n456), .B(shift_amount[4]), .Z(n455) );
  NAND U433 ( .A(n457), .B(n170), .Z(n452) );
  AND U434 ( .A(n458), .B(n162), .Z(n457) );
  NAND U435 ( .A(n459), .B(n460), .Z(c_shift[27]) );
  NAND U436 ( .A(n383), .B(\sll_27/ML_int[5][27] ), .Z(n460) );
  AND U437 ( .A(n461), .B(n462), .Z(n459) );
  NAND U438 ( .A(n463), .B(n150), .Z(n462) );
  NAND U439 ( .A(n464), .B(n395), .Z(n463) );
  OR U440 ( .A(n465), .B(shift_amount[4]), .Z(n464) );
  NAND U441 ( .A(n466), .B(n467), .Z(n461) );
  ANDN U442 ( .B(n218), .A(shift_amount[4]), .Z(n467) );
  ANDN U443 ( .B(n170), .A(n468), .Z(n466) );
  NAND U444 ( .A(n469), .B(n470), .Z(c_shift[26]) );
  NAND U445 ( .A(n383), .B(\sll_27/ML_int[5][26] ), .Z(n470) );
  AND U446 ( .A(n471), .B(n472), .Z(n469) );
  NAND U447 ( .A(n473), .B(n150), .Z(n472) );
  NAND U448 ( .A(n474), .B(n395), .Z(n473) );
  OR U449 ( .A(n475), .B(shift_amount[4]), .Z(n474) );
  NAND U450 ( .A(n476), .B(n170), .Z(n471) );
  NOR U451 ( .A(shift_amount[4]), .B(n477), .Z(n476) );
  NAND U452 ( .A(n478), .B(n479), .Z(c_shift[25]) );
  NAND U453 ( .A(n383), .B(\sll_27/ML_int[5][25] ), .Z(n479) );
  AND U454 ( .A(n480), .B(n481), .Z(n478) );
  NAND U455 ( .A(n482), .B(n150), .Z(n481) );
  NAND U456 ( .A(n483), .B(n395), .Z(n482) );
  OR U457 ( .A(n159), .B(shift_amount[4]), .Z(n483) );
  AND U458 ( .A(n484), .B(n485), .Z(n159) );
  NAND U459 ( .A(n486), .B(n487), .Z(n485) );
  AND U460 ( .A(n488), .B(n489), .Z(n484) );
  NAND U461 ( .A(n490), .B(n491), .Z(n489) );
  NAND U462 ( .A(n492), .B(n170), .Z(n480) );
  NOR U463 ( .A(shift_amount[4]), .B(n178), .Z(n492) );
  AND U464 ( .A(n493), .B(n494), .Z(n178) );
  NAND U465 ( .A(n495), .B(n487), .Z(n494) );
  NAND U466 ( .A(n449), .B(n491), .Z(n493) );
  NAND U467 ( .A(n496), .B(n497), .Z(c_shift[24]) );
  NAND U468 ( .A(n383), .B(\sll_27/ML_int[5][24] ), .Z(n497) );
  AND U469 ( .A(n498), .B(n499), .Z(n496) );
  NAND U470 ( .A(n500), .B(n150), .Z(n499) );
  NAND U471 ( .A(n501), .B(n395), .Z(n500) );
  OR U472 ( .A(n196), .B(shift_amount[4]), .Z(n501) );
  AND U473 ( .A(n502), .B(n503), .Z(n196) );
  NAND U474 ( .A(n504), .B(n487), .Z(n503) );
  AND U475 ( .A(n488), .B(n505), .Z(n502) );
  NAND U476 ( .A(n506), .B(n491), .Z(n505) );
  NAND U477 ( .A(n507), .B(n170), .Z(n498) );
  NOR U478 ( .A(shift_amount[4]), .B(n210), .Z(n507) );
  AND U479 ( .A(n508), .B(n509), .Z(n210) );
  NAND U480 ( .A(n510), .B(n487), .Z(n509) );
  NAND U481 ( .A(n458), .B(n491), .Z(n508) );
  NAND U482 ( .A(n511), .B(n512), .Z(c_shift[23]) );
  NAND U483 ( .A(n383), .B(\sll_27/ML_int[5][23] ), .Z(n512) );
  AND U484 ( .A(n513), .B(n514), .Z(n511) );
  NAND U485 ( .A(n515), .B(n150), .Z(n514) );
  NAND U486 ( .A(n516), .B(n395), .Z(n515) );
  OR U487 ( .A(n229), .B(shift_amount[4]), .Z(n516) );
  AND U488 ( .A(n517), .B(n518), .Z(n229) );
  NAND U489 ( .A(n519), .B(n487), .Z(n518) );
  AND U490 ( .A(n488), .B(n520), .Z(n517) );
  NAND U491 ( .A(n521), .B(n491), .Z(n520) );
  NAND U492 ( .A(n522), .B(n170), .Z(n513) );
  NOR U493 ( .A(shift_amount[4]), .B(n243), .Z(n522) );
  AND U494 ( .A(n523), .B(n524), .Z(n243) );
  NAND U495 ( .A(n525), .B(n487), .Z(n524) );
  AND U496 ( .A(n526), .B(n527), .Z(n523) );
  NANDN U497 ( .A(n528), .B(n491), .Z(n527) );
  NANDN U498 ( .A(n387), .B(n529), .Z(n526) );
  NAND U499 ( .A(n530), .B(n531), .Z(c_shift[22]) );
  NAND U500 ( .A(n383), .B(\sll_27/ML_int[5][22] ), .Z(n531) );
  AND U501 ( .A(n532), .B(n533), .Z(n530) );
  NAND U502 ( .A(n534), .B(n150), .Z(n533) );
  NAND U503 ( .A(n535), .B(n395), .Z(n534) );
  OR U504 ( .A(n261), .B(shift_amount[4]), .Z(n535) );
  AND U505 ( .A(n536), .B(n537), .Z(n261) );
  AND U506 ( .A(n538), .B(n539), .Z(n537) );
  NAND U507 ( .A(n540), .B(n487), .Z(n539) );
  NAND U508 ( .A(n541), .B(n491), .Z(n538) );
  AND U509 ( .A(n542), .B(n543), .Z(n536) );
  NAND U510 ( .A(n544), .B(n529), .Z(n543) );
  NAND U511 ( .A(n545), .B(n170), .Z(n532) );
  NOR U512 ( .A(shift_amount[4]), .B(n275), .Z(n545) );
  AND U513 ( .A(n546), .B(n547), .Z(n275) );
  NAND U514 ( .A(n548), .B(n487), .Z(n547) );
  AND U515 ( .A(n549), .B(n550), .Z(n546) );
  NAND U516 ( .A(n551), .B(n491), .Z(n550) );
  NAND U517 ( .A(n398), .B(n529), .Z(n549) );
  NAND U518 ( .A(n552), .B(n553), .Z(c_shift[21]) );
  NAND U519 ( .A(n383), .B(\sll_27/ML_int[5][21] ), .Z(n553) );
  AND U520 ( .A(n554), .B(n555), .Z(n552) );
  NAND U521 ( .A(n556), .B(n150), .Z(n555) );
  NAND U522 ( .A(n557), .B(n395), .Z(n556) );
  OR U523 ( .A(n292), .B(shift_amount[4]), .Z(n557) );
  AND U524 ( .A(n558), .B(n559), .Z(n292) );
  AND U525 ( .A(n542), .B(n560), .Z(n559) );
  NAND U526 ( .A(n155), .B(n487), .Z(n560) );
  AND U527 ( .A(n561), .B(n562), .Z(n558) );
  NAND U528 ( .A(n486), .B(n491), .Z(n562) );
  NAND U529 ( .A(n490), .B(n529), .Z(n561) );
  NAND U530 ( .A(n563), .B(n170), .Z(n554) );
  NOR U531 ( .A(shift_amount[4]), .B(n303), .Z(n563) );
  AND U532 ( .A(n564), .B(n565), .Z(n303) );
  NAND U533 ( .A(n175), .B(n487), .Z(n565) );
  AND U534 ( .A(n566), .B(n567), .Z(n564) );
  NAND U535 ( .A(n495), .B(n491), .Z(n567) );
  NAND U536 ( .A(n449), .B(n529), .Z(n566) );
  NAND U537 ( .A(n568), .B(n569), .Z(c_shift[20]) );
  NAND U538 ( .A(n383), .B(\sll_27/ML_int[5][20] ), .Z(n569) );
  AND U539 ( .A(n570), .B(n571), .Z(n568) );
  NAND U540 ( .A(n572), .B(n150), .Z(n571) );
  NAND U541 ( .A(n573), .B(n395), .Z(n572) );
  OR U542 ( .A(n318), .B(shift_amount[4]), .Z(n573) );
  AND U543 ( .A(n574), .B(n575), .Z(n318) );
  AND U544 ( .A(n542), .B(n576), .Z(n575) );
  NAND U545 ( .A(n193), .B(n487), .Z(n576) );
  AND U546 ( .A(n577), .B(n578), .Z(n574) );
  NAND U547 ( .A(n504), .B(n491), .Z(n578) );
  NAND U548 ( .A(n506), .B(n529), .Z(n577) );
  NAND U549 ( .A(n579), .B(n170), .Z(n570) );
  NOR U550 ( .A(shift_amount[4]), .B(n329), .Z(n579) );
  AND U551 ( .A(n580), .B(n581), .Z(n329) );
  NAND U552 ( .A(n207), .B(n487), .Z(n581) );
  AND U553 ( .A(n582), .B(n583), .Z(n580) );
  NAND U554 ( .A(n510), .B(n491), .Z(n583) );
  NAND U555 ( .A(n458), .B(n529), .Z(n582) );
  NAND U556 ( .A(n584), .B(n585), .Z(c_shift[1]) );
  NAND U557 ( .A(n146), .B(\sll_27/ML_int[4][1] ), .Z(n585) );
  AND U558 ( .A(\sll_27/ML_int[3][1] ), .B(n218), .Z(\sll_27/ML_int[4][1] ) );
  AND U559 ( .A(\sll_27/ML_int[2][1] ), .B(n335), .Z(\sll_27/ML_int[3][1] ) );
  AND U560 ( .A(\sll_27/ML_int[1][1] ), .B(n586), .Z(\sll_27/ML_int[2][1] ) );
  AND U561 ( .A(n587), .B(n588), .Z(n584) );
  NAND U562 ( .A(n589), .B(n150), .Z(n588) );
  NAND U563 ( .A(n590), .B(n591), .Z(n589) );
  AND U564 ( .A(n592), .B(n593), .Z(n591) );
  NANDN U565 ( .A(n161), .B(n166), .Z(n593) );
  AND U566 ( .A(n594), .B(n595), .Z(n161) );
  AND U567 ( .A(n596), .B(n597), .Z(n595) );
  NANDN U568 ( .A(n350), .B(value[9]), .Z(n597) );
  AND U569 ( .A(n598), .B(n599), .Z(n592) );
  OR U570 ( .A(n600), .B(n160), .Z(n599) );
  NANDN U571 ( .A(n293), .B(n168), .Z(n598) );
  AND U572 ( .A(n601), .B(n602), .Z(n293) );
  AND U573 ( .A(n603), .B(n604), .Z(n602) );
  NANDN U574 ( .A(n350), .B(value[5]), .Z(n604) );
  AND U575 ( .A(n605), .B(n606), .Z(n590) );
  NAND U576 ( .A(n607), .B(n162), .Z(n606) );
  NAND U577 ( .A(n608), .B(n609), .Z(n607) );
  AND U578 ( .A(n610), .B(n611), .Z(n609) );
  NANDN U579 ( .A(n350), .B(value[1]), .Z(n611) );
  NAND U580 ( .A(n156), .B(n167), .Z(n605) );
  NAND U581 ( .A(n612), .B(n170), .Z(n587) );
  NAND U582 ( .A(n613), .B(n614), .Z(n612) );
  AND U583 ( .A(n615), .B(n616), .Z(n614) );
  NANDN U584 ( .A(n179), .B(n166), .Z(n616) );
  AND U585 ( .A(n594), .B(n617), .Z(n179) );
  AND U586 ( .A(n596), .B(n618), .Z(n617) );
  NANDN U587 ( .A(n368), .B(value[9]), .Z(n618) );
  NAND U588 ( .A(n369), .B(value[10]), .Z(n596) );
  AND U589 ( .A(n619), .B(n620), .Z(n594) );
  NAND U590 ( .A(n372), .B(value[12]), .Z(n620) );
  NAND U591 ( .A(n373), .B(value[11]), .Z(n619) );
  AND U592 ( .A(n621), .B(n622), .Z(n615) );
  OR U593 ( .A(n623), .B(n160), .Z(n622) );
  NANDN U594 ( .A(n304), .B(n168), .Z(n621) );
  AND U595 ( .A(n601), .B(n624), .Z(n304) );
  AND U596 ( .A(n603), .B(n625), .Z(n624) );
  NANDN U597 ( .A(n368), .B(value[5]), .Z(n625) );
  NAND U598 ( .A(n369), .B(value[6]), .Z(n603) );
  AND U599 ( .A(n626), .B(n627), .Z(n601) );
  NAND U600 ( .A(n372), .B(value[8]), .Z(n627) );
  NAND U601 ( .A(n373), .B(value[7]), .Z(n626) );
  AND U602 ( .A(n628), .B(n629), .Z(n613) );
  NAND U603 ( .A(n630), .B(n162), .Z(n629) );
  NAND U604 ( .A(n608), .B(n631), .Z(n630) );
  AND U605 ( .A(n610), .B(n632), .Z(n631) );
  NANDN U606 ( .A(n368), .B(value[1]), .Z(n632) );
  NAND U607 ( .A(n369), .B(value[2]), .Z(n610) );
  AND U608 ( .A(n633), .B(n634), .Z(n608) );
  NAND U609 ( .A(n372), .B(value[4]), .Z(n634) );
  NAND U610 ( .A(n373), .B(value[3]), .Z(n633) );
  NAND U611 ( .A(n156), .B(n183), .Z(n628) );
  NAND U612 ( .A(n635), .B(n636), .Z(c_shift[19]) );
  NAND U613 ( .A(n383), .B(\sll_27/ML_int[5][19] ), .Z(n636) );
  AND U614 ( .A(n637), .B(n638), .Z(n635) );
  NAND U615 ( .A(n639), .B(n150), .Z(n638) );
  NAND U616 ( .A(n640), .B(n395), .Z(n639) );
  OR U617 ( .A(n345), .B(shift_amount[4]), .Z(n640) );
  AND U618 ( .A(n641), .B(n642), .Z(n345) );
  AND U619 ( .A(n542), .B(n643), .Z(n642) );
  NAND U620 ( .A(n226), .B(n487), .Z(n643) );
  NANDN U621 ( .A(n488), .B(shift_amount[2]), .Z(n542) );
  AND U622 ( .A(n644), .B(n645), .Z(n641) );
  NAND U623 ( .A(n519), .B(n491), .Z(n645) );
  NAND U624 ( .A(n521), .B(n529), .Z(n644) );
  NAND U625 ( .A(n646), .B(n170), .Z(n637) );
  NOR U626 ( .A(shift_amount[4]), .B(n365), .Z(n646) );
  AND U627 ( .A(n647), .B(n648), .Z(n365) );
  OR U628 ( .A(n468), .B(n218), .Z(n648) );
  AND U629 ( .A(n649), .B(n650), .Z(n647) );
  NAND U630 ( .A(n240), .B(n487), .Z(n650) );
  NAND U631 ( .A(n525), .B(n491), .Z(n649) );
  NAND U632 ( .A(n651), .B(n652), .Z(c_shift[18]) );
  NAND U633 ( .A(n383), .B(\sll_27/ML_int[5][18] ), .Z(n652) );
  AND U634 ( .A(n653), .B(n654), .Z(n651) );
  NAND U635 ( .A(n655), .B(n150), .Z(n654) );
  NAND U636 ( .A(n656), .B(n395), .Z(n655) );
  OR U637 ( .A(n410), .B(shift_amount[4]), .Z(n656) );
  AND U638 ( .A(n657), .B(n658), .Z(n410) );
  AND U639 ( .A(n659), .B(n660), .Z(n658) );
  NAND U640 ( .A(n258), .B(n487), .Z(n660) );
  NAND U641 ( .A(n540), .B(n491), .Z(n659) );
  AND U642 ( .A(n661), .B(n662), .Z(n657) );
  NAND U643 ( .A(n541), .B(n529), .Z(n662) );
  NANDN U644 ( .A(n663), .B(n544), .Z(n661) );
  NAND U645 ( .A(n664), .B(n170), .Z(n653) );
  NOR U646 ( .A(shift_amount[4]), .B(n429), .Z(n664) );
  AND U647 ( .A(n665), .B(n666), .Z(n429) );
  AND U648 ( .A(n667), .B(n668), .Z(n666) );
  NAND U649 ( .A(n272), .B(n487), .Z(n668) );
  NAND U650 ( .A(n548), .B(n491), .Z(n667) );
  AND U651 ( .A(n669), .B(n670), .Z(n665) );
  NAND U652 ( .A(n551), .B(n529), .Z(n670) );
  NANDN U653 ( .A(n663), .B(n398), .Z(n669) );
  NAND U654 ( .A(n671), .B(n672), .Z(c_shift[17]) );
  NAND U655 ( .A(n383), .B(\sll_27/ML_int[5][17] ), .Z(n672) );
  AND U656 ( .A(n673), .B(n674), .Z(n671) );
  NAND U657 ( .A(n675), .B(n150), .Z(n674) );
  NAND U658 ( .A(n676), .B(n395), .Z(n675) );
  OR U659 ( .A(n600), .B(shift_amount[4]), .Z(n676) );
  AND U660 ( .A(n677), .B(n678), .Z(n600) );
  AND U661 ( .A(n679), .B(n680), .Z(n678) );
  NAND U662 ( .A(n487), .B(n165), .Z(n680) );
  NAND U663 ( .A(n491), .B(n155), .Z(n679) );
  AND U664 ( .A(n681), .B(n682), .Z(n677) );
  NAND U665 ( .A(n529), .B(n486), .Z(n682) );
  NANDN U666 ( .A(n663), .B(n490), .Z(n681) );
  NAND U667 ( .A(n683), .B(n170), .Z(n673) );
  NOR U668 ( .A(shift_amount[4]), .B(n623), .Z(n683) );
  AND U669 ( .A(n684), .B(n685), .Z(n623) );
  AND U670 ( .A(n686), .B(n687), .Z(n685) );
  NAND U671 ( .A(n487), .B(n182), .Z(n687) );
  NAND U672 ( .A(n491), .B(n175), .Z(n686) );
  AND U673 ( .A(n688), .B(n689), .Z(n684) );
  NAND U674 ( .A(n529), .B(n495), .Z(n689) );
  NANDN U675 ( .A(n663), .B(n449), .Z(n688) );
  NAND U676 ( .A(n690), .B(n691), .Z(c_shift[16]) );
  NAND U677 ( .A(n383), .B(\sll_27/ML_int[5][16] ), .Z(n691) );
  AND U678 ( .A(n692), .B(n693), .Z(n690) );
  NAND U679 ( .A(n694), .B(n150), .Z(n693) );
  NAND U680 ( .A(n695), .B(n395), .Z(n694) );
  OR U681 ( .A(n696), .B(shift_amount[4]), .Z(n695) );
  NAND U682 ( .A(n697), .B(n170), .Z(n692) );
  NOR U683 ( .A(shift_amount[4]), .B(n698), .Z(n697) );
  NAND U684 ( .A(n699), .B(n700), .Z(c_shift[15]) );
  NAND U685 ( .A(n146), .B(\sll_27/ML_int[4][15] ), .Z(n700) );
  AND U686 ( .A(n701), .B(n702), .Z(n699) );
  NAND U687 ( .A(n703), .B(n150), .Z(n702) );
  NAND U688 ( .A(n704), .B(n705), .Z(n703) );
  AND U689 ( .A(n706), .B(n707), .Z(n705) );
  NAND U690 ( .A(n168), .B(n226), .Z(n707) );
  AND U691 ( .A(n395), .B(n708), .Z(n706) );
  NAND U692 ( .A(n162), .B(n233), .Z(n708) );
  NAND U693 ( .A(N75), .B(shift_amount[4]), .Z(n395) );
  AND U694 ( .A(n709), .B(n710), .Z(n704) );
  NAND U695 ( .A(n166), .B(n519), .Z(n710) );
  NAND U696 ( .A(n521), .B(n156), .Z(n709) );
  NAND U697 ( .A(n711), .B(n170), .Z(n701) );
  NAND U698 ( .A(n712), .B(n713), .Z(n711) );
  AND U699 ( .A(n714), .B(n715), .Z(n713) );
  NAND U700 ( .A(n166), .B(n525), .Z(n715) );
  AND U701 ( .A(n716), .B(n717), .Z(n714) );
  NAND U702 ( .A(n162), .B(n247), .Z(n717) );
  NAND U703 ( .A(n168), .B(n240), .Z(n716) );
  AND U704 ( .A(n718), .B(n719), .Z(n712) );
  OR U705 ( .A(n720), .B(n387), .Z(n719) );
  NANDN U706 ( .A(n528), .B(n156), .Z(n718) );
  NAND U707 ( .A(n721), .B(n722), .Z(c_shift[14]) );
  NAND U708 ( .A(n146), .B(\sll_27/ML_int[4][14] ), .Z(n722) );
  AND U709 ( .A(n723), .B(n724), .Z(n721) );
  NAND U710 ( .A(n725), .B(n150), .Z(n724) );
  NAND U711 ( .A(n726), .B(n727), .Z(n725) );
  AND U712 ( .A(n728), .B(n729), .Z(n727) );
  NAND U713 ( .A(n541), .B(n156), .Z(n729) );
  AND U714 ( .A(n730), .B(n731), .Z(n728) );
  OR U715 ( .A(n396), .B(n160), .Z(n731) );
  AND U716 ( .A(n732), .B(n733), .Z(n396) );
  NAND U717 ( .A(n544), .B(n487), .Z(n732) );
  NAND U718 ( .A(n162), .B(n265), .Z(n730) );
  AND U719 ( .A(n734), .B(n735), .Z(n726) );
  NAND U720 ( .A(n166), .B(n540), .Z(n735) );
  NAND U721 ( .A(n168), .B(n258), .Z(n734) );
  NAND U722 ( .A(n736), .B(n170), .Z(n723) );
  NAND U723 ( .A(n737), .B(n738), .Z(n736) );
  AND U724 ( .A(n739), .B(n740), .Z(n738) );
  NAND U725 ( .A(n166), .B(n548), .Z(n740) );
  AND U726 ( .A(n741), .B(n742), .Z(n739) );
  NAND U727 ( .A(n162), .B(n279), .Z(n742) );
  NAND U728 ( .A(n168), .B(n272), .Z(n741) );
  AND U729 ( .A(n743), .B(n744), .Z(n737) );
  NANDN U730 ( .A(n720), .B(n398), .Z(n744) );
  NAND U731 ( .A(n551), .B(n156), .Z(n743) );
  NAND U732 ( .A(n745), .B(n746), .Z(c_shift[13]) );
  NAND U733 ( .A(n146), .B(\sll_27/ML_int[4][13] ), .Z(n746) );
  AND U734 ( .A(n747), .B(n748), .Z(n745) );
  NAND U735 ( .A(n749), .B(n150), .Z(n748) );
  NAND U736 ( .A(n750), .B(n751), .Z(n749) );
  AND U737 ( .A(n752), .B(n753), .Z(n751) );
  NAND U738 ( .A(n486), .B(n156), .Z(n753) );
  NAND U739 ( .A(n754), .B(n755), .Z(n486) );
  AND U740 ( .A(n756), .B(n757), .Z(n755) );
  NANDN U741 ( .A(n350), .B(value[25]), .Z(n757) );
  AND U742 ( .A(n758), .B(n759), .Z(n752) );
  OR U743 ( .A(n447), .B(n160), .Z(n759) );
  AND U744 ( .A(n760), .B(n733), .Z(n447) );
  IV U745 ( .A(n761), .Z(n733) );
  NAND U746 ( .A(n487), .B(n490), .Z(n760) );
  NAND U747 ( .A(n762), .B(n763), .Z(n490) );
  NANDN U748 ( .A(n386), .B(shift_amount[1]), .Z(n763) );
  AND U749 ( .A(n764), .B(n765), .Z(n762) );
  NANDN U750 ( .A(n350), .B(value[29]), .Z(n765) );
  NAND U751 ( .A(n167), .B(n162), .Z(n758) );
  NAND U752 ( .A(n766), .B(n767), .Z(n167) );
  AND U753 ( .A(n768), .B(n769), .Z(n767) );
  NANDN U754 ( .A(n350), .B(value[13]), .Z(n769) );
  AND U755 ( .A(n770), .B(n771), .Z(n750) );
  NAND U756 ( .A(n155), .B(n166), .Z(n771) );
  NAND U757 ( .A(n772), .B(n773), .Z(n155) );
  AND U758 ( .A(n774), .B(n775), .Z(n773) );
  NANDN U759 ( .A(n350), .B(value[21]), .Z(n775) );
  NAND U760 ( .A(n165), .B(n168), .Z(n770) );
  NAND U761 ( .A(n776), .B(n777), .Z(n165) );
  AND U762 ( .A(n778), .B(n779), .Z(n777) );
  NANDN U763 ( .A(n350), .B(value[17]), .Z(n779) );
  NAND U764 ( .A(n780), .B(n170), .Z(n747) );
  NAND U765 ( .A(n781), .B(n782), .Z(n780) );
  AND U766 ( .A(n783), .B(n784), .Z(n782) );
  NAND U767 ( .A(n175), .B(n166), .Z(n784) );
  NAND U768 ( .A(n772), .B(n785), .Z(n175) );
  AND U769 ( .A(n774), .B(n786), .Z(n785) );
  NANDN U770 ( .A(n368), .B(value[21]), .Z(n786) );
  NAND U771 ( .A(n369), .B(value[22]), .Z(n774) );
  AND U772 ( .A(n787), .B(n788), .Z(n772) );
  NAND U773 ( .A(n372), .B(value[24]), .Z(n788) );
  NAND U774 ( .A(n373), .B(value[23]), .Z(n787) );
  AND U775 ( .A(n789), .B(n790), .Z(n783) );
  NAND U776 ( .A(n183), .B(n162), .Z(n790) );
  NAND U777 ( .A(n766), .B(n791), .Z(n183) );
  AND U778 ( .A(n768), .B(n792), .Z(n791) );
  NANDN U779 ( .A(n368), .B(value[13]), .Z(n792) );
  NAND U780 ( .A(n369), .B(value[14]), .Z(n768) );
  AND U781 ( .A(n793), .B(n794), .Z(n766) );
  NAND U782 ( .A(n372), .B(value[16]), .Z(n794) );
  NAND U783 ( .A(n373), .B(value[15]), .Z(n793) );
  NAND U784 ( .A(n182), .B(n168), .Z(n789) );
  NAND U785 ( .A(n776), .B(n795), .Z(n182) );
  AND U786 ( .A(n778), .B(n796), .Z(n795) );
  NANDN U787 ( .A(n368), .B(value[17]), .Z(n796) );
  NAND U788 ( .A(n369), .B(value[18]), .Z(n778) );
  AND U789 ( .A(n797), .B(n798), .Z(n776) );
  NAND U790 ( .A(n372), .B(value[20]), .Z(n798) );
  NAND U791 ( .A(n373), .B(value[19]), .Z(n797) );
  AND U792 ( .A(n799), .B(n800), .Z(n781) );
  NANDN U793 ( .A(n720), .B(n449), .Z(n800) );
  NAND U794 ( .A(n801), .B(n802), .Z(n449) );
  NANDN U795 ( .A(n368), .B(value[29]), .Z(n802) );
  AND U796 ( .A(n803), .B(n764), .Z(n801) );
  NAND U797 ( .A(n369), .B(value[30]), .Z(n764) );
  NANDN U798 ( .A(n386), .B(n373), .Z(n803) );
  NAND U799 ( .A(n495), .B(n156), .Z(n799) );
  NAND U800 ( .A(n754), .B(n804), .Z(n495) );
  AND U801 ( .A(n756), .B(n805), .Z(n804) );
  NANDN U802 ( .A(n368), .B(value[25]), .Z(n805) );
  NAND U803 ( .A(n369), .B(value[26]), .Z(n756) );
  AND U804 ( .A(n806), .B(n807), .Z(n754) );
  NAND U805 ( .A(n372), .B(value[28]), .Z(n807) );
  NAND U806 ( .A(n373), .B(value[27]), .Z(n806) );
  NAND U807 ( .A(n808), .B(n809), .Z(c_shift[12]) );
  NAND U808 ( .A(n146), .B(\sll_27/ML_int[4][12] ), .Z(n809) );
  AND U809 ( .A(n810), .B(n811), .Z(n808) );
  NAND U810 ( .A(n812), .B(n150), .Z(n811) );
  NAND U811 ( .A(n813), .B(n814), .Z(n812) );
  AND U812 ( .A(n815), .B(n816), .Z(n814) );
  NAND U813 ( .A(n504), .B(n156), .Z(n816) );
  AND U814 ( .A(n817), .B(n818), .Z(n815) );
  OR U815 ( .A(n456), .B(n160), .Z(n818) );
  ANDN U816 ( .B(n819), .A(n761), .Z(n456) );
  NAND U817 ( .A(n487), .B(n506), .Z(n819) );
  NAND U818 ( .A(n162), .B(n201), .Z(n817) );
  AND U819 ( .A(n820), .B(n821), .Z(n813) );
  NAND U820 ( .A(n193), .B(n166), .Z(n821) );
  NAND U821 ( .A(n200), .B(n168), .Z(n820) );
  NAND U822 ( .A(n822), .B(n170), .Z(n810) );
  NAND U823 ( .A(n823), .B(n824), .Z(n822) );
  AND U824 ( .A(n825), .B(n826), .Z(n824) );
  NAND U825 ( .A(n207), .B(n166), .Z(n826) );
  AND U826 ( .A(n827), .B(n828), .Z(n825) );
  NAND U827 ( .A(n162), .B(n215), .Z(n828) );
  NAND U828 ( .A(n214), .B(n168), .Z(n827) );
  AND U829 ( .A(n829), .B(n830), .Z(n823) );
  NANDN U830 ( .A(n720), .B(n458), .Z(n830) );
  NANDN U831 ( .A(n160), .B(n487), .Z(n720) );
  NAND U832 ( .A(n510), .B(n156), .Z(n829) );
  NAND U833 ( .A(n831), .B(n832), .Z(c_shift[11]) );
  NAND U834 ( .A(n146), .B(\sll_27/ML_int[4][11] ), .Z(n832) );
  AND U835 ( .A(n833), .B(n834), .Z(n831) );
  NAND U836 ( .A(n835), .B(n150), .Z(n834) );
  NAND U837 ( .A(n836), .B(n837), .Z(n835) );
  AND U838 ( .A(n838), .B(n839), .Z(n837) );
  NAND U839 ( .A(n519), .B(n156), .Z(n839) );
  NAND U840 ( .A(n840), .B(n841), .Z(n519) );
  AND U841 ( .A(n842), .B(n843), .Z(n841) );
  NANDN U842 ( .A(n350), .B(value[23]), .Z(n843) );
  AND U843 ( .A(n844), .B(n845), .Z(n838) );
  OR U844 ( .A(n465), .B(n160), .Z(n845) );
  ANDN U845 ( .B(n846), .A(n761), .Z(n465) );
  NAND U846 ( .A(n847), .B(n488), .Z(n761) );
  NANDN U847 ( .A(n386), .B(shift_amount[2]), .Z(n847) );
  NAND U848 ( .A(n487), .B(n521), .Z(n846) );
  NAND U849 ( .A(n848), .B(n849), .Z(n521) );
  AND U850 ( .A(n850), .B(n851), .Z(n849) );
  NANDN U851 ( .A(n350), .B(value[27]), .Z(n851) );
  NANDN U852 ( .A(n234), .B(n162), .Z(n844) );
  AND U853 ( .A(n852), .B(n853), .Z(n234) );
  AND U854 ( .A(n854), .B(n855), .Z(n853) );
  NANDN U855 ( .A(n350), .B(value[11]), .Z(n855) );
  AND U856 ( .A(n856), .B(n857), .Z(n836) );
  NAND U857 ( .A(n226), .B(n166), .Z(n857) );
  NAND U858 ( .A(n858), .B(n859), .Z(n226) );
  AND U859 ( .A(n860), .B(n861), .Z(n859) );
  NANDN U860 ( .A(n350), .B(value[19]), .Z(n861) );
  NAND U861 ( .A(n233), .B(n168), .Z(n856) );
  NAND U862 ( .A(n862), .B(n863), .Z(n233) );
  AND U863 ( .A(n864), .B(n865), .Z(n863) );
  NANDN U864 ( .A(n350), .B(value[15]), .Z(n865) );
  NAND U865 ( .A(n866), .B(n170), .Z(n833) );
  NAND U866 ( .A(n867), .B(n868), .Z(n866) );
  AND U867 ( .A(n869), .B(n870), .Z(n868) );
  NAND U868 ( .A(n240), .B(n166), .Z(n870) );
  NAND U869 ( .A(n858), .B(n871), .Z(n240) );
  AND U870 ( .A(n860), .B(n872), .Z(n871) );
  NANDN U871 ( .A(n368), .B(value[19]), .Z(n872) );
  NAND U872 ( .A(n369), .B(value[20]), .Z(n860) );
  AND U873 ( .A(n873), .B(n874), .Z(n858) );
  NAND U874 ( .A(n372), .B(value[22]), .Z(n874) );
  NAND U875 ( .A(n373), .B(value[21]), .Z(n873) );
  AND U876 ( .A(n875), .B(n876), .Z(n869) );
  NANDN U877 ( .A(n248), .B(n162), .Z(n876) );
  AND U878 ( .A(n852), .B(n877), .Z(n248) );
  AND U879 ( .A(n854), .B(n878), .Z(n877) );
  NANDN U880 ( .A(n368), .B(value[11]), .Z(n878) );
  NAND U881 ( .A(n369), .B(value[12]), .Z(n854) );
  AND U882 ( .A(n879), .B(n880), .Z(n852) );
  NAND U883 ( .A(n372), .B(value[14]), .Z(n880) );
  NAND U884 ( .A(n373), .B(value[13]), .Z(n879) );
  NAND U885 ( .A(n247), .B(n168), .Z(n875) );
  NAND U886 ( .A(n862), .B(n881), .Z(n247) );
  AND U887 ( .A(n864), .B(n882), .Z(n881) );
  NANDN U888 ( .A(n368), .B(value[15]), .Z(n882) );
  NAND U889 ( .A(n369), .B(value[16]), .Z(n864) );
  AND U890 ( .A(n883), .B(n884), .Z(n862) );
  NAND U891 ( .A(n372), .B(value[18]), .Z(n884) );
  NAND U892 ( .A(n373), .B(value[17]), .Z(n883) );
  AND U893 ( .A(n885), .B(n886), .Z(n867) );
  NANDN U894 ( .A(n468), .B(n887), .Z(n886) );
  ANDN U895 ( .B(n218), .A(n160), .Z(n887) );
  MUX U896 ( .IN0(n528), .IN1(n387), .SEL(shift_amount[2]), .F(n468) );
  OR U897 ( .A(n368), .B(n386), .Z(n387) );
  AND U898 ( .A(n848), .B(n888), .Z(n528) );
  AND U899 ( .A(n850), .B(n889), .Z(n888) );
  NANDN U900 ( .A(n368), .B(value[27]), .Z(n889) );
  NAND U901 ( .A(n369), .B(value[28]), .Z(n850) );
  AND U902 ( .A(n890), .B(n891), .Z(n848) );
  NAND U903 ( .A(value[30]), .B(n372), .Z(n891) );
  NAND U904 ( .A(value[29]), .B(n373), .Z(n890) );
  NAND U905 ( .A(n525), .B(n156), .Z(n885) );
  NAND U906 ( .A(n840), .B(n892), .Z(n525) );
  AND U907 ( .A(n842), .B(n893), .Z(n892) );
  NANDN U908 ( .A(n368), .B(value[23]), .Z(n893) );
  NAND U909 ( .A(n369), .B(value[24]), .Z(n842) );
  AND U910 ( .A(n894), .B(n895), .Z(n840) );
  NAND U911 ( .A(value[26]), .B(n372), .Z(n895) );
  NAND U912 ( .A(value[25]), .B(n373), .Z(n894) );
  NAND U913 ( .A(n896), .B(n897), .Z(c_shift[10]) );
  NAND U914 ( .A(n146), .B(\sll_27/ML_int[4][10] ), .Z(n897) );
  AND U915 ( .A(n898), .B(n899), .Z(n896) );
  NAND U916 ( .A(n900), .B(n150), .Z(n899) );
  NAND U917 ( .A(n901), .B(n902), .Z(n900) );
  AND U918 ( .A(n903), .B(n904), .Z(n902) );
  NAND U919 ( .A(n540), .B(n156), .Z(n904) );
  NAND U920 ( .A(n905), .B(n906), .Z(n540) );
  AND U921 ( .A(n907), .B(n908), .Z(n906) );
  NANDN U922 ( .A(n350), .B(value[22]), .Z(n908) );
  AND U923 ( .A(n909), .B(n910), .Z(n903) );
  OR U924 ( .A(n475), .B(n160), .Z(n910) );
  AND U925 ( .A(n911), .B(n912), .Z(n475) );
  NAND U926 ( .A(n487), .B(n541), .Z(n912) );
  NAND U927 ( .A(n913), .B(n914), .Z(n541) );
  AND U928 ( .A(n915), .B(n916), .Z(n914) );
  NANDN U929 ( .A(n350), .B(value[26]), .Z(n916) );
  AND U930 ( .A(n488), .B(n917), .Z(n911) );
  NAND U931 ( .A(n544), .B(n491), .Z(n917) );
  MUX U932 ( .IN0(N75), .IN1(value[30]), .SEL(n918), .F(n544) );
  NAND U933 ( .A(N75), .B(shift_amount[3]), .Z(n488) );
  NANDN U934 ( .A(n266), .B(n162), .Z(n909) );
  AND U935 ( .A(n919), .B(n920), .Z(n266) );
  AND U936 ( .A(n921), .B(n922), .Z(n920) );
  NANDN U937 ( .A(n350), .B(value[10]), .Z(n922) );
  AND U938 ( .A(n923), .B(n924), .Z(n901) );
  NAND U939 ( .A(n258), .B(n166), .Z(n924) );
  NAND U940 ( .A(n925), .B(n926), .Z(n258) );
  AND U941 ( .A(n927), .B(n928), .Z(n926) );
  NANDN U942 ( .A(n350), .B(value[18]), .Z(n928) );
  NAND U943 ( .A(n265), .B(n168), .Z(n923) );
  NAND U944 ( .A(n929), .B(n930), .Z(n265) );
  AND U945 ( .A(n931), .B(n932), .Z(n930) );
  NANDN U946 ( .A(n350), .B(value[14]), .Z(n932) );
  NAND U947 ( .A(n933), .B(n170), .Z(n898) );
  NAND U948 ( .A(n934), .B(n935), .Z(n933) );
  AND U949 ( .A(n936), .B(n937), .Z(n935) );
  NAND U950 ( .A(n548), .B(n156), .Z(n937) );
  NAND U951 ( .A(n905), .B(n938), .Z(n548) );
  AND U952 ( .A(n907), .B(n939), .Z(n938) );
  NANDN U953 ( .A(n368), .B(value[22]), .Z(n939) );
  NAND U954 ( .A(n369), .B(value[23]), .Z(n907) );
  AND U955 ( .A(n940), .B(n941), .Z(n905) );
  NAND U956 ( .A(value[25]), .B(n372), .Z(n941) );
  NAND U957 ( .A(n373), .B(value[24]), .Z(n940) );
  AND U958 ( .A(n942), .B(n943), .Z(n936) );
  OR U959 ( .A(n477), .B(n160), .Z(n943) );
  AND U960 ( .A(n944), .B(n945), .Z(n477) );
  NAND U961 ( .A(n487), .B(n551), .Z(n945) );
  NAND U962 ( .A(n913), .B(n946), .Z(n551) );
  AND U963 ( .A(n915), .B(n947), .Z(n946) );
  NANDN U964 ( .A(n368), .B(value[26]), .Z(n947) );
  NAND U965 ( .A(n369), .B(value[27]), .Z(n915) );
  AND U966 ( .A(n948), .B(n949), .Z(n913) );
  NAND U967 ( .A(value[29]), .B(n372), .Z(n949) );
  NAND U968 ( .A(value[28]), .B(n373), .Z(n948) );
  NAND U969 ( .A(n398), .B(n491), .Z(n944) );
  NAND U970 ( .A(n950), .B(n951), .Z(n398) );
  NANDN U971 ( .A(n386), .B(n369), .Z(n951) );
  NANDN U972 ( .A(n368), .B(value[30]), .Z(n950) );
  NANDN U973 ( .A(n280), .B(n162), .Z(n942) );
  AND U974 ( .A(n919), .B(n952), .Z(n280) );
  AND U975 ( .A(n921), .B(n953), .Z(n952) );
  NANDN U976 ( .A(n368), .B(value[10]), .Z(n953) );
  NAND U977 ( .A(n369), .B(value[11]), .Z(n921) );
  AND U978 ( .A(n954), .B(n955), .Z(n919) );
  NAND U979 ( .A(n372), .B(value[13]), .Z(n955) );
  NAND U980 ( .A(n373), .B(value[12]), .Z(n954) );
  AND U981 ( .A(n956), .B(n957), .Z(n934) );
  NAND U982 ( .A(n272), .B(n166), .Z(n957) );
  NAND U983 ( .A(n925), .B(n958), .Z(n272) );
  AND U984 ( .A(n927), .B(n959), .Z(n958) );
  NANDN U985 ( .A(n368), .B(value[18]), .Z(n959) );
  NAND U986 ( .A(n369), .B(value[19]), .Z(n927) );
  AND U987 ( .A(n960), .B(n961), .Z(n925) );
  NAND U988 ( .A(n372), .B(value[21]), .Z(n961) );
  NAND U989 ( .A(n373), .B(value[20]), .Z(n960) );
  NAND U990 ( .A(n279), .B(n168), .Z(n956) );
  NAND U991 ( .A(n929), .B(n962), .Z(n279) );
  AND U992 ( .A(n931), .B(n963), .Z(n962) );
  NANDN U993 ( .A(n368), .B(value[14]), .Z(n963) );
  NAND U994 ( .A(n369), .B(value[15]), .Z(n931) );
  AND U995 ( .A(n964), .B(n965), .Z(n929) );
  NAND U996 ( .A(n372), .B(value[17]), .Z(n965) );
  NAND U997 ( .A(n373), .B(value[16]), .Z(n964) );
  NAND U998 ( .A(n966), .B(n967), .Z(c_shift[0]) );
  NAND U999 ( .A(n146), .B(\sll_27/ML_int[4][0] ), .Z(n967) );
  AND U1000 ( .A(\sll_27/ML_int[3][0] ), .B(n218), .Z(\sll_27/ML_int[4][0] )
         );
  AND U1001 ( .A(\sll_27/ML_int[2][0] ), .B(n335), .Z(\sll_27/ML_int[3][0] )
         );
  AND U1002 ( .A(\sll_27/ML_int[1][0] ), .B(n586), .Z(\sll_27/ML_int[2][0] )
         );
  AND U1003 ( .A(value[0]), .B(n968), .Z(\sll_27/ML_int[1][0] ) );
  ANDN U1004 ( .B(n383), .A(shift_amount[4]), .Z(n146) );
  ANDN U1005 ( .B(shift_func[0]), .A(shift_func[1]), .Z(n383) );
  AND U1006 ( .A(n969), .B(n970), .Z(n966) );
  NAND U1007 ( .A(n971), .B(n150), .Z(n970) );
  AND U1008 ( .A(shift_func[0]), .B(shift_func[1]), .Z(n150) );
  NAND U1009 ( .A(n972), .B(n973), .Z(n971) );
  AND U1010 ( .A(n974), .B(n975), .Z(n973) );
  NANDN U1011 ( .A(n197), .B(n166), .Z(n975) );
  AND U1012 ( .A(n976), .B(n977), .Z(n197) );
  AND U1013 ( .A(n978), .B(n979), .Z(n977) );
  NANDN U1014 ( .A(n350), .B(value[8]), .Z(n979) );
  AND U1015 ( .A(n980), .B(n981), .Z(n974) );
  OR U1016 ( .A(n696), .B(n160), .Z(n981) );
  AND U1017 ( .A(n982), .B(n983), .Z(n696) );
  AND U1018 ( .A(n984), .B(n985), .Z(n983) );
  NAND U1019 ( .A(n487), .B(n200), .Z(n985) );
  NAND U1020 ( .A(n986), .B(n987), .Z(n200) );
  AND U1021 ( .A(n988), .B(n989), .Z(n987) );
  NANDN U1022 ( .A(n350), .B(value[16]), .Z(n989) );
  NAND U1023 ( .A(n491), .B(n193), .Z(n984) );
  NAND U1024 ( .A(n990), .B(n991), .Z(n193) );
  AND U1025 ( .A(n992), .B(n993), .Z(n991) );
  NANDN U1026 ( .A(n350), .B(value[20]), .Z(n993) );
  AND U1027 ( .A(n994), .B(n995), .Z(n982) );
  NAND U1028 ( .A(n529), .B(n504), .Z(n995) );
  NAND U1029 ( .A(n996), .B(n997), .Z(n504) );
  AND U1030 ( .A(n998), .B(n999), .Z(n997) );
  NANDN U1031 ( .A(n350), .B(value[24]), .Z(n999) );
  NANDN U1032 ( .A(n663), .B(n506), .Z(n994) );
  NAND U1033 ( .A(n1000), .B(n1001), .Z(n506) );
  AND U1034 ( .A(n1002), .B(n1003), .Z(n1001) );
  NANDN U1035 ( .A(n350), .B(value[28]), .Z(n1003) );
  NANDN U1036 ( .A(n319), .B(n168), .Z(n980) );
  AND U1037 ( .A(n1004), .B(n1005), .Z(n319) );
  AND U1038 ( .A(n1006), .B(n1007), .Z(n1005) );
  NANDN U1039 ( .A(n350), .B(value[4]), .Z(n1007) );
  AND U1040 ( .A(n1008), .B(n1009), .Z(n972) );
  NAND U1041 ( .A(n1010), .B(n162), .Z(n1009) );
  NAND U1042 ( .A(n1011), .B(n1012), .Z(n1010) );
  AND U1043 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U1044 ( .A(n350), .B(value[0]), .Z(n1014) );
  NAND U1045 ( .A(n156), .B(n201), .Z(n1008) );
  NAND U1046 ( .A(n1015), .B(n1016), .Z(n201) );
  AND U1047 ( .A(n1017), .B(n1018), .Z(n1016) );
  NANDN U1048 ( .A(n350), .B(value[12]), .Z(n1018) );
  IV U1049 ( .A(n918), .Z(n350) );
  NOR U1050 ( .A(shift_amount[0]), .B(shift_amount[1]), .Z(n918) );
  NAND U1051 ( .A(n1019), .B(n170), .Z(n969) );
  ANDN U1052 ( .B(shift_func[1]), .A(shift_func[0]), .Z(n170) );
  NAND U1053 ( .A(n1020), .B(n1021), .Z(n1019) );
  AND U1054 ( .A(n1022), .B(n1023), .Z(n1021) );
  NANDN U1055 ( .A(n211), .B(n166), .Z(n1023) );
  NOR U1056 ( .A(shift_amount[2]), .B(n1024), .Z(n166) );
  AND U1057 ( .A(n976), .B(n1025), .Z(n211) );
  AND U1058 ( .A(n978), .B(n1026), .Z(n1025) );
  NANDN U1059 ( .A(n368), .B(value[8]), .Z(n1026) );
  NAND U1060 ( .A(n369), .B(value[9]), .Z(n978) );
  AND U1061 ( .A(n1027), .B(n1028), .Z(n976) );
  NAND U1062 ( .A(n372), .B(value[11]), .Z(n1028) );
  NAND U1063 ( .A(n373), .B(value[10]), .Z(n1027) );
  AND U1064 ( .A(n1029), .B(n1030), .Z(n1022) );
  OR U1065 ( .A(n698), .B(n160), .Z(n1030) );
  AND U1066 ( .A(n1031), .B(n1032), .Z(n698) );
  AND U1067 ( .A(n1033), .B(n1034), .Z(n1032) );
  NAND U1068 ( .A(n487), .B(n214), .Z(n1034) );
  NAND U1069 ( .A(n986), .B(n1035), .Z(n214) );
  AND U1070 ( .A(n988), .B(n1036), .Z(n1035) );
  NANDN U1071 ( .A(n368), .B(value[16]), .Z(n1036) );
  NAND U1072 ( .A(n369), .B(value[17]), .Z(n988) );
  AND U1073 ( .A(n1037), .B(n1038), .Z(n986) );
  NAND U1074 ( .A(n372), .B(value[19]), .Z(n1038) );
  NAND U1075 ( .A(n373), .B(value[18]), .Z(n1037) );
  NAND U1076 ( .A(n491), .B(n207), .Z(n1033) );
  NAND U1077 ( .A(n990), .B(n1039), .Z(n207) );
  AND U1078 ( .A(n992), .B(n1040), .Z(n1039) );
  NANDN U1079 ( .A(n368), .B(value[20]), .Z(n1040) );
  NAND U1080 ( .A(n369), .B(value[21]), .Z(n992) );
  AND U1081 ( .A(n1041), .B(n1042), .Z(n990) );
  NAND U1082 ( .A(n372), .B(value[23]), .Z(n1042) );
  NAND U1083 ( .A(n373), .B(value[22]), .Z(n1041) );
  AND U1084 ( .A(n1043), .B(n1044), .Z(n1031) );
  NAND U1085 ( .A(n529), .B(n510), .Z(n1044) );
  NAND U1086 ( .A(n996), .B(n1045), .Z(n510) );
  AND U1087 ( .A(n998), .B(n1046), .Z(n1045) );
  NANDN U1088 ( .A(n368), .B(value[24]), .Z(n1046) );
  NAND U1089 ( .A(n369), .B(value[25]), .Z(n998) );
  AND U1090 ( .A(n1047), .B(n1048), .Z(n996) );
  NAND U1091 ( .A(n372), .B(value[27]), .Z(n1048) );
  NAND U1092 ( .A(value[26]), .B(n373), .Z(n1047) );
  AND U1093 ( .A(shift_amount[3]), .B(n335), .Z(n529) );
  NANDN U1094 ( .A(n663), .B(n458), .Z(n1043) );
  NAND U1095 ( .A(n1000), .B(n1049), .Z(n458) );
  AND U1096 ( .A(n1002), .B(n1050), .Z(n1049) );
  NANDN U1097 ( .A(n368), .B(value[28]), .Z(n1050) );
  NAND U1098 ( .A(value[29]), .B(n369), .Z(n1002) );
  AND U1099 ( .A(n1051), .B(n1052), .Z(n1000) );
  NANDN U1100 ( .A(n386), .B(n372), .Z(n1052) );
  IV U1101 ( .A(N75), .Z(n386) );
  NAND U1102 ( .A(value[30]), .B(n373), .Z(n1051) );
  NANDN U1103 ( .A(n335), .B(shift_amount[3]), .Z(n663) );
  NANDN U1104 ( .A(n330), .B(n168), .Z(n1029) );
  AND U1105 ( .A(n491), .B(n160), .Z(n168) );
  ANDN U1106 ( .B(shift_amount[2]), .A(shift_amount[3]), .Z(n491) );
  AND U1107 ( .A(n1004), .B(n1053), .Z(n330) );
  AND U1108 ( .A(n1006), .B(n1054), .Z(n1053) );
  NANDN U1109 ( .A(n368), .B(value[4]), .Z(n1054) );
  NAND U1110 ( .A(n369), .B(value[5]), .Z(n1006) );
  AND U1111 ( .A(n1055), .B(n1056), .Z(n1004) );
  NAND U1112 ( .A(n372), .B(value[7]), .Z(n1056) );
  NAND U1113 ( .A(n373), .B(value[6]), .Z(n1055) );
  AND U1114 ( .A(n1057), .B(n1058), .Z(n1020) );
  NAND U1115 ( .A(n1059), .B(n162), .Z(n1058) );
  AND U1116 ( .A(n487), .B(n160), .Z(n162) );
  IV U1117 ( .A(shift_amount[4]), .Z(n160) );
  ANDN U1118 ( .B(n218), .A(shift_amount[2]), .Z(n487) );
  IV U1119 ( .A(shift_amount[3]), .Z(n218) );
  NAND U1120 ( .A(n1011), .B(n1060), .Z(n1059) );
  AND U1121 ( .A(n1013), .B(n1061), .Z(n1060) );
  NANDN U1122 ( .A(n368), .B(value[0]), .Z(n1061) );
  NAND U1123 ( .A(n369), .B(value[1]), .Z(n1013) );
  AND U1124 ( .A(n1062), .B(n1063), .Z(n1011) );
  NAND U1125 ( .A(n372), .B(value[3]), .Z(n1063) );
  NAND U1126 ( .A(n373), .B(value[2]), .Z(n1062) );
  NAND U1127 ( .A(n156), .B(n215), .Z(n1057) );
  NAND U1128 ( .A(n1015), .B(n1064), .Z(n215) );
  AND U1129 ( .A(n1017), .B(n1065), .Z(n1064) );
  NANDN U1130 ( .A(n368), .B(value[12]), .Z(n1065) );
  NANDN U1131 ( .A(shift_amount[0]), .B(n586), .Z(n368) );
  NAND U1132 ( .A(n369), .B(value[13]), .Z(n1017) );
  AND U1133 ( .A(shift_amount[0]), .B(n586), .Z(n369) );
  IV U1134 ( .A(shift_amount[1]), .Z(n586) );
  AND U1135 ( .A(n1066), .B(n1067), .Z(n1015) );
  NAND U1136 ( .A(n372), .B(value[15]), .Z(n1067) );
  AND U1137 ( .A(shift_amount[0]), .B(shift_amount[1]), .Z(n372) );
  NAND U1138 ( .A(n373), .B(value[14]), .Z(n1066) );
  AND U1139 ( .A(shift_amount[1]), .B(n968), .Z(n373) );
  IV U1140 ( .A(shift_amount[0]), .Z(n968) );
  NOR U1141 ( .A(n335), .B(n1024), .Z(n156) );
  NANDN U1142 ( .A(shift_amount[4]), .B(shift_amount[3]), .Z(n1024) );
  IV U1143 ( .A(shift_amount[2]), .Z(n335) );
endmodule

