
module mult_N64_CC2 ( clk, rst, a, b, c );
  input [63:0] a;
  input [31:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964;
  wire   [127:0] sreg;

  DFF \sreg_reg[95]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[94]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[93]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[92]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[91]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[90]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[89]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[88]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[87]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[86]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[85]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[84]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[83]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[82]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[81]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[80]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[79]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[78]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[77]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[76]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[75]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[74]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[73]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[72]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[71]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[70]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[69]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[68]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[67]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[66]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[65]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[64]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[63]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(sreg[63]) );
  DFF \sreg_reg[62]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(sreg[62]) );
  DFF \sreg_reg[61]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(sreg[61]) );
  DFF \sreg_reg[60]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(sreg[60]) );
  DFF \sreg_reg[59]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(sreg[59]) );
  DFF \sreg_reg[58]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(sreg[58]) );
  DFF \sreg_reg[57]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(sreg[57]) );
  DFF \sreg_reg[56]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(sreg[56]) );
  DFF \sreg_reg[55]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(sreg[55]) );
  DFF \sreg_reg[54]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(sreg[54]) );
  DFF \sreg_reg[53]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(sreg[53]) );
  DFF \sreg_reg[52]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(sreg[52]) );
  DFF \sreg_reg[51]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(sreg[51]) );
  DFF \sreg_reg[50]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(sreg[50]) );
  DFF \sreg_reg[49]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(sreg[49]) );
  DFF \sreg_reg[48]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(sreg[48]) );
  DFF \sreg_reg[47]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(sreg[47]) );
  DFF \sreg_reg[46]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(sreg[46]) );
  DFF \sreg_reg[45]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(sreg[45]) );
  DFF \sreg_reg[44]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(sreg[44]) );
  DFF \sreg_reg[43]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(sreg[43]) );
  DFF \sreg_reg[42]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(sreg[42]) );
  DFF \sreg_reg[41]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(sreg[41]) );
  DFF \sreg_reg[40]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(sreg[40]) );
  DFF \sreg_reg[39]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(sreg[39]) );
  DFF \sreg_reg[38]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(sreg[38]) );
  DFF \sreg_reg[37]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(sreg[37]) );
  DFF \sreg_reg[36]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(sreg[36]) );
  DFF \sreg_reg[35]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(sreg[35]) );
  DFF \sreg_reg[34]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(sreg[34]) );
  DFF \sreg_reg[33]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(sreg[33]) );
  DFF \sreg_reg[32]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(sreg[32]) );
  DFF \sreg_reg[31]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[0]) );
  ANDN U35 ( .B(n2616), .A(n320), .Z(n1) );
  AND U36 ( .A(n9706), .B(n1), .Z(n2) );
  NOR U37 ( .A(n320), .B(b[24]), .Z(n3) );
  NAND U38 ( .A(n3), .B(n319), .Z(n4) );
  NANDN U39 ( .A(n2), .B(n4), .Z(n1883) );
  XNOR U40 ( .A(n4339), .B(n4338), .Z(n4340) );
  XNOR U41 ( .A(n4970), .B(n4969), .Z(n4971) );
  XNOR U42 ( .A(n5817), .B(n5816), .Z(n5818) );
  XNOR U43 ( .A(n6114), .B(n6113), .Z(n6115) );
  XNOR U44 ( .A(n6262), .B(n6261), .Z(n6263) );
  XNOR U45 ( .A(n6447), .B(n6446), .Z(n6448) );
  OR U46 ( .A(n1072), .B(n1073), .Z(n1182) );
  ANDN U47 ( .B(n2616), .A(n318), .Z(n5) );
  AND U48 ( .A(n9493), .B(n5), .Z(n6) );
  NOR U49 ( .A(n318), .B(b[20]), .Z(n7) );
  NAND U50 ( .A(n7), .B(n9562), .Z(n8) );
  NANDN U51 ( .A(n6), .B(n8), .Z(n1413) );
  NAND U52 ( .A(n1900), .B(n1899), .Z(n9) );
  NANDN U53 ( .A(n1898), .B(n1897), .Z(n10) );
  NAND U54 ( .A(n9), .B(n10), .Z(n1954) );
  NAND U55 ( .A(n2448), .B(n2447), .Z(n11) );
  NANDN U56 ( .A(n2446), .B(n2445), .Z(n12) );
  NAND U57 ( .A(n11), .B(n12), .Z(n2641) );
  NAND U58 ( .A(n2893), .B(n2892), .Z(n13) );
  NANDN U59 ( .A(n2895), .B(n2894), .Z(n14) );
  AND U60 ( .A(n13), .B(n14), .Z(n3116) );
  NAND U61 ( .A(n3033), .B(n3032), .Z(n15) );
  NANDN U62 ( .A(n3035), .B(n3034), .Z(n16) );
  AND U63 ( .A(n15), .B(n16), .Z(n3206) );
  XNOR U64 ( .A(n3341), .B(n3342), .Z(n3344) );
  XNOR U65 ( .A(n3636), .B(n3637), .Z(n3639) );
  XNOR U66 ( .A(n4092), .B(n4093), .Z(n4095) );
  XNOR U67 ( .A(n4830), .B(n4831), .Z(n4833) );
  NAND U68 ( .A(n4966), .B(n4965), .Z(n17) );
  NANDN U69 ( .A(n4968), .B(n4967), .Z(n18) );
  AND U70 ( .A(n17), .B(n18), .Z(n5122) );
  XNOR U71 ( .A(n5419), .B(n5420), .Z(n5422) );
  NAND U72 ( .A(n6443), .B(n6442), .Z(n19) );
  NANDN U73 ( .A(n6445), .B(n6444), .Z(n20) );
  AND U74 ( .A(n19), .B(n20), .Z(n6600) );
  NANDN U75 ( .A(n2114), .B(n2113), .Z(n21) );
  NANDN U76 ( .A(n2112), .B(n2111), .Z(n22) );
  NAND U77 ( .A(n21), .B(n22), .Z(n2188) );
  NAND U78 ( .A(n978), .B(n977), .Z(n23) );
  NANDN U79 ( .A(n976), .B(n975), .Z(n24) );
  NAND U80 ( .A(n23), .B(n24), .Z(n1052) );
  NAND U81 ( .A(n1499), .B(n1500), .Z(n25) );
  NANDN U82 ( .A(n1498), .B(n1497), .Z(n26) );
  NAND U83 ( .A(n25), .B(n26), .Z(n1602) );
  NAND U84 ( .A(n2579), .B(n2578), .Z(n27) );
  NAND U85 ( .A(n2576), .B(n2577), .Z(n28) );
  NAND U86 ( .A(n27), .B(n28), .Z(n2844) );
  NAND U87 ( .A(n8074), .B(n8073), .Z(n29) );
  NANDN U88 ( .A(n8072), .B(n8071), .Z(n30) );
  NAND U89 ( .A(n29), .B(n30), .Z(n8111) );
  NAND U90 ( .A(n9549), .B(n9548), .Z(n31) );
  NANDN U91 ( .A(n9547), .B(n9546), .Z(n32) );
  NAND U92 ( .A(n31), .B(n32), .Z(n9604) );
  NAND U93 ( .A(n9607), .B(n9608), .Z(n33) );
  NANDN U94 ( .A(n9606), .B(n9605), .Z(n34) );
  NAND U95 ( .A(n33), .B(n34), .Z(n9646) );
  NANDN U96 ( .A(n7756), .B(b[3]), .Z(n35) );
  NANDN U97 ( .A(b[2]), .B(b[1]), .Z(n36) );
  NAND U98 ( .A(n35), .B(n36), .Z(n37) );
  NAND U99 ( .A(n7620), .B(n2616), .Z(n38) );
  NAND U100 ( .A(n38), .B(n37), .Z(n39) );
  NANDN U101 ( .A(n316), .B(n39), .Z(n360) );
  NAND U102 ( .A(n8222), .B(n8221), .Z(n40) );
  NANDN U103 ( .A(n8220), .B(n8219), .Z(n41) );
  AND U104 ( .A(n40), .B(n41), .Z(n8227) );
  NAND U105 ( .A(n7976), .B(n7975), .Z(n42) );
  XOR U106 ( .A(n7975), .B(n7976), .Z(n43) );
  NAND U107 ( .A(n43), .B(n7974), .Z(n44) );
  NAND U108 ( .A(n42), .B(n44), .Z(n8104) );
  NAND U109 ( .A(n8471), .B(n8470), .Z(n45) );
  NANDN U110 ( .A(n8469), .B(n8468), .Z(n46) );
  AND U111 ( .A(n45), .B(n46), .Z(n8579) );
  NAND U112 ( .A(n2516), .B(n2515), .Z(n47) );
  NANDN U113 ( .A(n2514), .B(n2513), .Z(n48) );
  AND U114 ( .A(n47), .B(n48), .Z(n2635) );
  XNOR U115 ( .A(n3173), .B(n3172), .Z(n3217) );
  XNOR U116 ( .A(n3454), .B(n3453), .Z(n3455) );
  XNOR U117 ( .A(n3898), .B(n3897), .Z(n3899) );
  XNOR U118 ( .A(n4192), .B(n4191), .Z(n4193) );
  XNOR U119 ( .A(n4636), .B(n4635), .Z(n4637) );
  XNOR U120 ( .A(n5235), .B(n5234), .Z(n5236) );
  XOR U121 ( .A(n6107), .B(n6108), .Z(n6109) );
  XOR U122 ( .A(n6101), .B(n6102), .Z(n6103) );
  XNOR U123 ( .A(n6264), .B(n6263), .Z(n6310) );
  NANDN U124 ( .A(n318), .B(n9669), .Z(n49) );
  ANDN U125 ( .B(n2616), .A(n9621), .Z(n50) );
  NANDN U126 ( .A(b[22]), .B(n49), .Z(n51) );
  NANDN U127 ( .A(n50), .B(n51), .Z(n52) );
  ANDN U128 ( .B(n52), .A(n319), .Z(n1640) );
  NAND U129 ( .A(n2028), .B(n2027), .Z(n53) );
  NANDN U130 ( .A(n2029), .B(n2030), .Z(n54) );
  AND U131 ( .A(n53), .B(n54), .Z(n2066) );
  NAND U132 ( .A(n2373), .B(n2372), .Z(n55) );
  NANDN U133 ( .A(n2371), .B(n2370), .Z(n56) );
  AND U134 ( .A(n55), .B(n56), .Z(n2469) );
  NAND U135 ( .A(n2407), .B(n2408), .Z(n57) );
  NANDN U136 ( .A(n2406), .B(n2405), .Z(n58) );
  NAND U137 ( .A(n57), .B(n58), .Z(n2474) );
  NAND U138 ( .A(n2641), .B(n2640), .Z(n59) );
  NANDN U139 ( .A(n2639), .B(n2638), .Z(n60) );
  NAND U140 ( .A(n59), .B(n60), .Z(n2744) );
  OR U141 ( .A(n2973), .B(n2974), .Z(n61) );
  NAND U142 ( .A(n2976), .B(n2975), .Z(n62) );
  NAND U143 ( .A(n61), .B(n62), .Z(n3005) );
  XOR U144 ( .A(n3783), .B(n3784), .Z(n3785) );
  XNOR U145 ( .A(n4533), .B(n4534), .Z(n4536) );
  XOR U146 ( .A(n5566), .B(n5567), .Z(n5568) );
  XOR U147 ( .A(n5703), .B(n5704), .Z(n5705) );
  XNOR U148 ( .A(n5999), .B(n6000), .Z(n6002) );
  XNOR U149 ( .A(n6297), .B(n6298), .Z(n6300) );
  XNOR U150 ( .A(n6700), .B(n6699), .Z(n6701) );
  NAND U151 ( .A(n1064), .B(n1065), .Z(n63) );
  NANDN U152 ( .A(n1063), .B(n1062), .Z(n64) );
  NAND U153 ( .A(n63), .B(n64), .Z(n1188) );
  NAND U154 ( .A(n1232), .B(n1231), .Z(n65) );
  NANDN U155 ( .A(n1230), .B(n1229), .Z(n66) );
  NAND U156 ( .A(n65), .B(n66), .Z(n1375) );
  NAND U157 ( .A(n1462), .B(n1461), .Z(n67) );
  NANDN U158 ( .A(n1460), .B(n1459), .Z(n68) );
  NAND U159 ( .A(n67), .B(n68), .Z(n1579) );
  NAND U160 ( .A(n2034), .B(n2033), .Z(n69) );
  NANDN U161 ( .A(n2032), .B(n2031), .Z(n70) );
  NAND U162 ( .A(n69), .B(n70), .Z(n2158) );
  NAND U163 ( .A(n3119), .B(n3118), .Z(n71) );
  NANDN U164 ( .A(n3117), .B(n3116), .Z(n72) );
  NAND U165 ( .A(n71), .B(n72), .Z(n3271) );
  NAND U166 ( .A(n3209), .B(n3208), .Z(n73) );
  NANDN U167 ( .A(n3207), .B(n3206), .Z(n74) );
  NAND U168 ( .A(n73), .B(n74), .Z(n3419) );
  NAND U169 ( .A(n3405), .B(n3404), .Z(n75) );
  NAND U170 ( .A(n3402), .B(n3403), .Z(n76) );
  NAND U171 ( .A(n75), .B(n76), .Z(n3562) );
  NAND U172 ( .A(n3699), .B(n3698), .Z(n77) );
  NAND U173 ( .A(n3696), .B(n3697), .Z(n78) );
  NAND U174 ( .A(n77), .B(n78), .Z(n3857) );
  NAND U175 ( .A(n4155), .B(n4154), .Z(n79) );
  NAND U176 ( .A(n4152), .B(n4153), .Z(n80) );
  NAND U177 ( .A(n79), .B(n80), .Z(n4300) );
  NAND U178 ( .A(n4893), .B(n4892), .Z(n81) );
  NAND U179 ( .A(n4890), .B(n4891), .Z(n82) );
  NAND U180 ( .A(n81), .B(n82), .Z(n4918) );
  XNOR U181 ( .A(n5189), .B(n5190), .Z(n5184) );
  NAND U182 ( .A(n5125), .B(n5124), .Z(n83) );
  NANDN U183 ( .A(n5123), .B(n5122), .Z(n84) );
  NAND U184 ( .A(n83), .B(n84), .Z(n5217) );
  NAND U185 ( .A(n5482), .B(n5481), .Z(n85) );
  NAND U186 ( .A(n5479), .B(n5480), .Z(n86) );
  NAND U187 ( .A(n85), .B(n86), .Z(n5507) );
  XNOR U188 ( .A(n6666), .B(n6667), .Z(n6661) );
  NAND U189 ( .A(n6603), .B(n6602), .Z(n87) );
  NANDN U190 ( .A(n6601), .B(n6600), .Z(n88) );
  NAND U191 ( .A(n87), .B(n88), .Z(n6812) );
  OR U192 ( .A(n6737), .B(n6738), .Z(n89) );
  NAND U193 ( .A(n6736), .B(n6735), .Z(n90) );
  NAND U194 ( .A(n89), .B(n90), .Z(n6951) );
  NAND U195 ( .A(n8058), .B(n8057), .Z(n91) );
  NANDN U196 ( .A(n8056), .B(n8055), .Z(n92) );
  AND U197 ( .A(n91), .B(n92), .Z(n8182) );
  NAND U198 ( .A(n8280), .B(n8279), .Z(n93) );
  NANDN U199 ( .A(n8278), .B(n8277), .Z(n94) );
  AND U200 ( .A(n93), .B(n94), .Z(n8378) );
  NANDN U201 ( .A(n922), .B(n921), .Z(n95) );
  NANDN U202 ( .A(n920), .B(n919), .Z(n96) );
  NAND U203 ( .A(n95), .B(n96), .Z(n970) );
  NAND U204 ( .A(n925), .B(n926), .Z(n97) );
  NANDN U205 ( .A(n924), .B(n923), .Z(n98) );
  NAND U206 ( .A(n97), .B(n98), .Z(n964) );
  NANDN U207 ( .A(n989), .B(n988), .Z(n99) );
  NANDN U208 ( .A(n991), .B(n990), .Z(n100) );
  NAND U209 ( .A(n99), .B(n100), .Z(n1055) );
  NAND U210 ( .A(n2144), .B(n2143), .Z(n101) );
  NANDN U211 ( .A(n2142), .B(n2141), .Z(n102) );
  AND U212 ( .A(n101), .B(n102), .Z(n2289) );
  NAND U213 ( .A(n6944), .B(n6943), .Z(n103) );
  NANDN U214 ( .A(n6942), .B(n6941), .Z(n104) );
  NAND U215 ( .A(n103), .B(n104), .Z(n7097) );
  NAND U216 ( .A(n8669), .B(n8668), .Z(n105) );
  NANDN U217 ( .A(n8667), .B(n8666), .Z(n106) );
  NAND U218 ( .A(n105), .B(n106), .Z(n8765) );
  NAND U219 ( .A(n8972), .B(n8971), .Z(n107) );
  NANDN U220 ( .A(n8970), .B(n8969), .Z(n108) );
  AND U221 ( .A(n107), .B(n108), .Z(n8994) );
  NAND U222 ( .A(n9310), .B(n9309), .Z(n109) );
  NANDN U223 ( .A(n9308), .B(n9307), .Z(n110) );
  NAND U224 ( .A(n109), .B(n110), .Z(n9328) );
  NAND U225 ( .A(n2844), .B(n2843), .Z(n111) );
  NANDN U226 ( .A(n2842), .B(n2841), .Z(n112) );
  NAND U227 ( .A(n111), .B(n112), .Z(n2851) );
  NAND U228 ( .A(n9226), .B(n9225), .Z(n113) );
  NANDN U229 ( .A(n9224), .B(n9223), .Z(n114) );
  NAND U230 ( .A(n113), .B(n114), .Z(n9255) );
  XOR U231 ( .A(n372), .B(n371), .Z(n115) );
  NANDN U232 ( .A(n373), .B(n115), .Z(n116) );
  NAND U233 ( .A(n372), .B(n371), .Z(n117) );
  AND U234 ( .A(n116), .B(n117), .Z(n398) );
  NAND U235 ( .A(n1601), .B(n1602), .Z(n118) );
  NANDN U236 ( .A(n1600), .B(n1599), .Z(n119) );
  NAND U237 ( .A(n118), .B(n119), .Z(n1694) );
  NAND U238 ( .A(n1496), .B(n1495), .Z(n120) );
  NANDN U239 ( .A(n1494), .B(n1493), .Z(n121) );
  NAND U240 ( .A(n120), .B(n121), .Z(n1596) );
  NAND U241 ( .A(n4025), .B(n4024), .Z(n122) );
  NAND U242 ( .A(n4022), .B(n4023), .Z(n123) );
  NAND U243 ( .A(n122), .B(n123), .Z(n4170) );
  NAND U244 ( .A(n4466), .B(n4465), .Z(n124) );
  NAND U245 ( .A(n4463), .B(n4464), .Z(n125) );
  NAND U246 ( .A(n124), .B(n125), .Z(n4614) );
  NAND U247 ( .A(n6242), .B(n6241), .Z(n126) );
  NAND U248 ( .A(n6239), .B(n6240), .Z(n127) );
  NAND U249 ( .A(n126), .B(n127), .Z(n6387) );
  NAND U250 ( .A(n8114), .B(n8113), .Z(n128) );
  NANDN U251 ( .A(n8112), .B(n8111), .Z(n129) );
  NAND U252 ( .A(n128), .B(n129), .Z(n8229) );
  NAND U253 ( .A(n9604), .B(n9603), .Z(n130) );
  NANDN U254 ( .A(n9602), .B(n9601), .Z(n131) );
  NAND U255 ( .A(n130), .B(n131), .Z(n9649) );
  XOR U256 ( .A(n8102), .B(n8103), .Z(n132) );
  NANDN U257 ( .A(n8104), .B(n132), .Z(n133) );
  NAND U258 ( .A(n8102), .B(n8103), .Z(n134) );
  AND U259 ( .A(n133), .B(n134), .Z(n8226) );
  NAND U260 ( .A(n8580), .B(n8579), .Z(n135) );
  XOR U261 ( .A(n8579), .B(n8580), .Z(n136) );
  NAND U262 ( .A(n136), .B(n8578), .Z(n137) );
  NAND U263 ( .A(n135), .B(n137), .Z(n8687) );
  XOR U264 ( .A(n9159), .B(n9158), .Z(n138) );
  NANDN U265 ( .A(n9157), .B(n138), .Z(n139) );
  NAND U266 ( .A(n9159), .B(n9158), .Z(n140) );
  AND U267 ( .A(n139), .B(n140), .Z(n9246) );
  NAND U268 ( .A(n9744), .B(n9743), .Z(n141) );
  XOR U269 ( .A(n9743), .B(n9744), .Z(n142) );
  NAND U270 ( .A(n142), .B(n9742), .Z(n143) );
  NAND U271 ( .A(n141), .B(n143), .Z(n9785) );
  NANDN U272 ( .A(n2616), .B(b[29]), .Z(n144) );
  ANDN U273 ( .B(n144), .A(n323), .Z(n145) );
  XNOR U274 ( .A(b[29]), .B(n2616), .Z(n146) );
  NANDN U275 ( .A(n2512), .B(n146), .Z(n147) );
  NAND U276 ( .A(n145), .B(n147), .Z(n2599) );
  NANDN U277 ( .A(n2520), .B(n2519), .Z(n148) );
  NANDN U278 ( .A(n2518), .B(n2517), .Z(n149) );
  NAND U279 ( .A(n148), .B(n149), .Z(n2645) );
  NAND U280 ( .A(n2972), .B(n2971), .Z(n150) );
  NANDN U281 ( .A(n2970), .B(n2969), .Z(n151) );
  NAND U282 ( .A(n150), .B(n151), .Z(n3062) );
  XNOR U283 ( .A(n3171), .B(n3170), .Z(n3172) );
  XOR U284 ( .A(n3164), .B(n3165), .Z(n3166) );
  XOR U285 ( .A(n3158), .B(n3159), .Z(n3160) );
  XOR U286 ( .A(n3447), .B(n3448), .Z(n3449) );
  XNOR U287 ( .A(n3456), .B(n3455), .Z(n3502) );
  XOR U288 ( .A(n3441), .B(n3442), .Z(n3443) );
  XOR U289 ( .A(n3891), .B(n3892), .Z(n3893) );
  XNOR U290 ( .A(n3900), .B(n3899), .Z(n3946) );
  XOR U291 ( .A(n3885), .B(n3886), .Z(n3887) );
  XOR U292 ( .A(n4185), .B(n4186), .Z(n4187) );
  XNOR U293 ( .A(n4194), .B(n4193), .Z(n4240) );
  XNOR U294 ( .A(n4180), .B(n4179), .Z(n4181) );
  XOR U295 ( .A(n4332), .B(n4333), .Z(n4334) );
  XNOR U296 ( .A(n4341), .B(n4340), .Z(n4387) );
  XNOR U297 ( .A(n4327), .B(n4326), .Z(n4328) );
  XOR U298 ( .A(n4629), .B(n4630), .Z(n4631) );
  XNOR U299 ( .A(n4638), .B(n4637), .Z(n4684) );
  XOR U300 ( .A(n4623), .B(n4624), .Z(n4625) );
  XOR U301 ( .A(n5228), .B(n5229), .Z(n5230) );
  XNOR U302 ( .A(n5237), .B(n5236), .Z(n5283) );
  XOR U303 ( .A(n5222), .B(n5223), .Z(n5224) );
  XOR U304 ( .A(n5810), .B(n5811), .Z(n5812) );
  XNOR U305 ( .A(n5819), .B(n5818), .Z(n5865) );
  XNOR U306 ( .A(n5805), .B(n5804), .Z(n5806) );
  XNOR U307 ( .A(n6116), .B(n6115), .Z(n6163) );
  XOR U308 ( .A(n6255), .B(n6256), .Z(n6257) );
  XNOR U309 ( .A(n6250), .B(n6249), .Z(n6251) );
  XOR U310 ( .A(n6576), .B(n6577), .Z(n6578) );
  NOR U311 ( .A(n1260), .B(n1261), .Z(n1357) );
  NOR U312 ( .A(b[26]), .B(n321), .Z(n152) );
  NANDN U313 ( .A(n320), .B(n9837), .Z(n153) );
  NAND U314 ( .A(n152), .B(n153), .Z(n154) );
  NANDN U315 ( .A(a[0]), .B(n9804), .Z(n155) );
  NAND U316 ( .A(n154), .B(n155), .Z(n2137) );
  NAND U317 ( .A(n2404), .B(n2403), .Z(n156) );
  NANDN U318 ( .A(n2402), .B(n2401), .Z(n157) );
  NAND U319 ( .A(n156), .B(n157), .Z(n2473) );
  XOR U320 ( .A(n2745), .B(n2746), .Z(n2747) );
  XOR U321 ( .A(n3489), .B(n3490), .Z(n3491) );
  XOR U322 ( .A(n3933), .B(n3934), .Z(n3935) );
  XOR U323 ( .A(n4227), .B(n4228), .Z(n4229) );
  XNOR U324 ( .A(n4374), .B(n4375), .Z(n4377) );
  XOR U325 ( .A(n4671), .B(n4672), .Z(n4673) );
  XOR U326 ( .A(n4975), .B(n4976), .Z(n4977) );
  XOR U327 ( .A(n5270), .B(n5271), .Z(n5272) );
  XOR U328 ( .A(n5852), .B(n5853), .Z(n5854) );
  XOR U329 ( .A(n6150), .B(n6151), .Z(n6152) );
  XNOR U330 ( .A(n6452), .B(n6453), .Z(n6455) );
  XOR U331 ( .A(n6693), .B(n6694), .Z(n6695) );
  XNOR U332 ( .A(n6702), .B(n6701), .Z(n6746) );
  XNOR U333 ( .A(n6688), .B(n6687), .Z(n6689) );
  NAND U334 ( .A(a[63]), .B(n315), .Z(n158) );
  AND U335 ( .A(b[1]), .B(n158), .Z(n7463) );
  ANDN U336 ( .B(n2616), .A(n9562), .Z(n159) );
  AND U337 ( .A(n9378), .B(n159), .Z(n160) );
  NOR U338 ( .A(n9562), .B(b[18]), .Z(n161) );
  NAND U339 ( .A(n161), .B(n9455), .Z(n162) );
  NANDN U340 ( .A(n160), .B(n162), .Z(n1249) );
  NAND U341 ( .A(n1660), .B(n1659), .Z(n163) );
  NANDN U342 ( .A(n1658), .B(n1657), .Z(n164) );
  AND U343 ( .A(n163), .B(n164), .Z(n1800) );
  NAND U344 ( .A(n1904), .B(n1903), .Z(n165) );
  NANDN U345 ( .A(n1902), .B(n1901), .Z(n166) );
  AND U346 ( .A(n165), .B(n166), .Z(n1948) );
  NAND U347 ( .A(n2244), .B(n2243), .Z(n167) );
  NANDN U348 ( .A(n2242), .B(n2241), .Z(n168) );
  NAND U349 ( .A(n167), .B(n168), .Z(n2417) );
  NAND U350 ( .A(n2263), .B(n2262), .Z(n169) );
  NANDN U351 ( .A(n2261), .B(n2260), .Z(n170) );
  NAND U352 ( .A(n169), .B(n170), .Z(n2328) );
  NAND U353 ( .A(n2472), .B(n2471), .Z(n171) );
  NANDN U354 ( .A(n2470), .B(n2469), .Z(n172) );
  AND U355 ( .A(n171), .B(n172), .Z(n2581) );
  NANDN U356 ( .A(n2742), .B(n2741), .Z(n173) );
  NANDN U357 ( .A(n2744), .B(n2743), .Z(n174) );
  NAND U358 ( .A(n173), .B(n174), .Z(n2869) );
  XOR U359 ( .A(n3126), .B(n3127), .Z(n3128) );
  NAND U360 ( .A(n3013), .B(n3012), .Z(n175) );
  NAND U361 ( .A(n3010), .B(n3011), .Z(n176) );
  NAND U362 ( .A(n175), .B(n176), .Z(n3265) );
  NAND U363 ( .A(n3151), .B(n3150), .Z(n177) );
  XOR U364 ( .A(n3150), .B(n3151), .Z(n178) );
  NAND U365 ( .A(n178), .B(n3149), .Z(n179) );
  NAND U366 ( .A(n177), .B(n179), .Z(n3412) );
  XNOR U367 ( .A(n3569), .B(n3570), .Z(n3564) );
  XNOR U368 ( .A(n3864), .B(n3865), .Z(n3859) );
  XNOR U369 ( .A(n4013), .B(n4014), .Z(n4008) );
  XNOR U370 ( .A(n4307), .B(n4308), .Z(n4302) );
  XNOR U371 ( .A(n4751), .B(n4752), .Z(n4746) );
  XNOR U372 ( .A(n4925), .B(n4926), .Z(n4920) );
  NAND U373 ( .A(n5071), .B(n5070), .Z(n180) );
  NANDN U374 ( .A(n5073), .B(n5072), .Z(n181) );
  NAND U375 ( .A(n180), .B(n181), .Z(n5211) );
  XNOR U376 ( .A(n5514), .B(n5515), .Z(n5509) );
  XNOR U377 ( .A(n5783), .B(n5784), .Z(n5778) );
  XNOR U378 ( .A(n5932), .B(n5933), .Z(n5927) );
  XNOR U379 ( .A(n6230), .B(n6231), .Z(n6225) );
  NAND U380 ( .A(n6360), .B(n6359), .Z(n182) );
  NAND U381 ( .A(n6357), .B(n6358), .Z(n183) );
  NAND U382 ( .A(n182), .B(n183), .Z(n6395) );
  NAND U383 ( .A(n6549), .B(n6548), .Z(n184) );
  NANDN U384 ( .A(n6551), .B(n6550), .Z(n185) );
  NAND U385 ( .A(n184), .B(n185), .Z(n6806) );
  XNOR U386 ( .A(n6880), .B(n6881), .Z(n6883) );
  XNOR U387 ( .A(n7571), .B(n7570), .Z(n7572) );
  XOR U388 ( .A(n7564), .B(n7565), .Z(n7567) );
  NAND U389 ( .A(n7892), .B(n7891), .Z(n186) );
  NANDN U390 ( .A(n7890), .B(n7889), .Z(n187) );
  NAND U391 ( .A(n186), .B(n187), .Z(n8084) );
  NAND U392 ( .A(n8203), .B(n8202), .Z(n188) );
  NANDN U393 ( .A(n8201), .B(n8200), .Z(n189) );
  NAND U394 ( .A(n188), .B(n189), .Z(n8249) );
  NAND U395 ( .A(n8276), .B(n8275), .Z(n190) );
  NANDN U396 ( .A(n8274), .B(n8273), .Z(n191) );
  NAND U397 ( .A(n190), .B(n191), .Z(n8377) );
  NAND U398 ( .A(n8433), .B(n8432), .Z(n192) );
  NANDN U399 ( .A(n8431), .B(n8430), .Z(n193) );
  NAND U400 ( .A(n192), .B(n193), .Z(n8550) );
  NAND U401 ( .A(n912), .B(n911), .Z(n194) );
  NANDN U402 ( .A(n910), .B(n909), .Z(n195) );
  NAND U403 ( .A(n194), .B(n195), .Z(n972) );
  NAND U404 ( .A(n836), .B(n835), .Z(n196) );
  NANDN U405 ( .A(n834), .B(n833), .Z(n197) );
  NAND U406 ( .A(n196), .B(n197), .Z(n903) );
  NAND U407 ( .A(n1110), .B(n1109), .Z(n198) );
  NANDN U408 ( .A(n1108), .B(n1107), .Z(n199) );
  AND U409 ( .A(n198), .B(n199), .Z(n1123) );
  NAND U410 ( .A(n1188), .B(n1187), .Z(n200) );
  NANDN U411 ( .A(n1186), .B(n1185), .Z(n201) );
  AND U412 ( .A(n200), .B(n201), .Z(n1224) );
  XNOR U413 ( .A(n1402), .B(n1403), .Z(n1478) );
  NANDN U414 ( .A(n1572), .B(n1571), .Z(n202) );
  NANDN U415 ( .A(n1570), .B(n1569), .Z(n203) );
  NAND U416 ( .A(n202), .B(n203), .Z(n1684) );
  NAND U417 ( .A(n1837), .B(n1836), .Z(n204) );
  NANDN U418 ( .A(n1835), .B(n1834), .Z(n205) );
  AND U419 ( .A(n204), .B(n205), .Z(n1941) );
  NANDN U420 ( .A(n2158), .B(n2157), .Z(n206) );
  NANDN U421 ( .A(n2160), .B(n2159), .Z(n207) );
  AND U422 ( .A(n206), .B(n207), .Z(n2179) );
  NAND U423 ( .A(n6987), .B(n6986), .Z(n208) );
  NANDN U424 ( .A(n6985), .B(n6984), .Z(n209) );
  NAND U425 ( .A(n208), .B(n209), .Z(n7132) );
  NAND U426 ( .A(n7713), .B(n7712), .Z(n210) );
  NANDN U427 ( .A(n7711), .B(n7710), .Z(n211) );
  NAND U428 ( .A(n210), .B(n211), .Z(n7853) );
  XNOR U429 ( .A(n8059), .B(n8060), .Z(n8062) );
  NANDN U430 ( .A(n8124), .B(n8123), .Z(n212) );
  NANDN U431 ( .A(n8122), .B(n8121), .Z(n213) );
  NAND U432 ( .A(n212), .B(n213), .Z(n8234) );
  NAND U433 ( .A(n8370), .B(n8369), .Z(n214) );
  NANDN U434 ( .A(n8368), .B(n8367), .Z(n215) );
  NAND U435 ( .A(n214), .B(n215), .Z(n8478) );
  XOR U436 ( .A(n8595), .B(n8594), .Z(n216) );
  NANDN U437 ( .A(n8593), .B(n216), .Z(n217) );
  NAND U438 ( .A(n8595), .B(n8594), .Z(n218) );
  AND U439 ( .A(n217), .B(n218), .Z(n8688) );
  NAND U440 ( .A(n8762), .B(n8761), .Z(n219) );
  NANDN U441 ( .A(n8760), .B(n8759), .Z(n220) );
  NAND U442 ( .A(n219), .B(n220), .Z(n8867) );
  NANDN U443 ( .A(n8597), .B(n8596), .Z(n221) );
  NANDN U444 ( .A(n8599), .B(n8598), .Z(n222) );
  NAND U445 ( .A(n221), .B(n222), .Z(n8707) );
  NAND U446 ( .A(n8946), .B(n8945), .Z(n223) );
  NANDN U447 ( .A(n8948), .B(n8947), .Z(n224) );
  NAND U448 ( .A(n223), .B(n224), .Z(n9001) );
  NAND U449 ( .A(n9008), .B(n9007), .Z(n225) );
  NANDN U450 ( .A(n9006), .B(n9005), .Z(n226) );
  NAND U451 ( .A(n225), .B(n226), .Z(n9142) );
  NAND U452 ( .A(n9098), .B(n9097), .Z(n227) );
  NANDN U453 ( .A(n9096), .B(n9095), .Z(n228) );
  NAND U454 ( .A(n227), .B(n228), .Z(n9229) );
  XOR U455 ( .A(n9348), .B(n9347), .Z(n229) );
  NANDN U456 ( .A(n9346), .B(n229), .Z(n230) );
  NAND U457 ( .A(n9348), .B(n9347), .Z(n231) );
  AND U458 ( .A(n230), .B(n231), .Z(n9408) );
  ANDN U459 ( .B(n2616), .A(n317), .Z(n232) );
  AND U460 ( .A(n7905), .B(n232), .Z(n233) );
  NOR U461 ( .A(n317), .B(b[4]), .Z(n234) );
  NAND U462 ( .A(n234), .B(n316), .Z(n235) );
  NANDN U463 ( .A(n233), .B(n235), .Z(n414) );
  NAND U464 ( .A(n950), .B(n949), .Z(n236) );
  NANDN U465 ( .A(n948), .B(n947), .Z(n237) );
  AND U466 ( .A(n236), .B(n237), .Z(n1025) );
  NANDN U467 ( .A(n1053), .B(n1052), .Z(n238) );
  NANDN U468 ( .A(n1055), .B(n1054), .Z(n239) );
  NAND U469 ( .A(n238), .B(n239), .Z(n1117) );
  NAND U470 ( .A(n2291), .B(n2290), .Z(n240) );
  NANDN U471 ( .A(n2289), .B(n2288), .Z(n241) );
  NAND U472 ( .A(n240), .B(n241), .Z(n2422) );
  NAND U473 ( .A(n6977), .B(n6976), .Z(n242) );
  NANDN U474 ( .A(n6975), .B(n6974), .Z(n243) );
  NAND U475 ( .A(n242), .B(n243), .Z(n7113) );
  NAND U476 ( .A(n7431), .B(n7432), .Z(n244) );
  NANDN U477 ( .A(n7430), .B(n7429), .Z(n245) );
  NAND U478 ( .A(n244), .B(n245), .Z(n7559) );
  NAND U479 ( .A(n7646), .B(n7645), .Z(n246) );
  NANDN U480 ( .A(n7644), .B(n7643), .Z(n247) );
  NAND U481 ( .A(n246), .B(n247), .Z(n7819) );
  NAND U482 ( .A(n8242), .B(n8241), .Z(n248) );
  NANDN U483 ( .A(n8240), .B(n8239), .Z(n249) );
  NAND U484 ( .A(n248), .B(n249), .Z(n8349) );
  NANDN U485 ( .A(n8701), .B(n8700), .Z(n250) );
  NANDN U486 ( .A(n8703), .B(n8702), .Z(n251) );
  NAND U487 ( .A(n250), .B(n251), .Z(n8876) );
  NAND U488 ( .A(n9094), .B(n9093), .Z(n252) );
  NANDN U489 ( .A(n9092), .B(n9091), .Z(n253) );
  AND U490 ( .A(n252), .B(n253), .Z(n9161) );
  OR U491 ( .A(n9512), .B(n9513), .Z(n254) );
  NANDN U492 ( .A(n9511), .B(n9510), .Z(n255) );
  NAND U493 ( .A(n254), .B(n255), .Z(n9580) );
  NAND U494 ( .A(n9629), .B(n9628), .Z(n256) );
  NANDN U495 ( .A(n9627), .B(n9626), .Z(n257) );
  NAND U496 ( .A(n256), .B(n257), .Z(n9681) );
  NAND U497 ( .A(n9701), .B(n9700), .Z(n258) );
  XOR U498 ( .A(n9700), .B(n9701), .Z(n259) );
  NANDN U499 ( .A(n9702), .B(n259), .Z(n260) );
  NAND U500 ( .A(n258), .B(n260), .Z(n9767) );
  OR U501 ( .A(n451), .B(n452), .Z(n261) );
  NAND U502 ( .A(n454), .B(n453), .Z(n262) );
  NAND U503 ( .A(n261), .B(n262), .Z(n466) );
  NAND U504 ( .A(n596), .B(n595), .Z(n263) );
  NANDN U505 ( .A(n594), .B(n593), .Z(n264) );
  NAND U506 ( .A(n263), .B(n264), .Z(n645) );
  NAND U507 ( .A(n2704), .B(n2703), .Z(n265) );
  NANDN U508 ( .A(n2702), .B(n2701), .Z(n266) );
  AND U509 ( .A(n265), .B(n266), .Z(n2706) );
  NAND U510 ( .A(n2997), .B(n2996), .Z(n267) );
  NANDN U511 ( .A(n2995), .B(n2994), .Z(n268) );
  NAND U512 ( .A(n267), .B(n268), .Z(n3140) );
  NAND U513 ( .A(n3581), .B(n3580), .Z(n269) );
  NAND U514 ( .A(n3578), .B(n3579), .Z(n270) );
  NAND U515 ( .A(n269), .B(n270), .Z(n3726) );
  NAND U516 ( .A(n4319), .B(n4318), .Z(n271) );
  NAND U517 ( .A(n4316), .B(n4317), .Z(n272) );
  NAND U518 ( .A(n271), .B(n272), .Z(n4466) );
  NAND U519 ( .A(n4763), .B(n4762), .Z(n273) );
  NAND U520 ( .A(n4760), .B(n4761), .Z(n274) );
  NAND U521 ( .A(n273), .B(n274), .Z(n4908) );
  NAND U522 ( .A(n5944), .B(n5943), .Z(n275) );
  NAND U523 ( .A(n5941), .B(n5942), .Z(n276) );
  NAND U524 ( .A(n275), .B(n276), .Z(n6092) );
  NAND U525 ( .A(n6387), .B(n6386), .Z(n277) );
  NAND U526 ( .A(n6384), .B(n6385), .Z(n278) );
  NAND U527 ( .A(n277), .B(n278), .Z(n6533) );
  NAND U528 ( .A(n6825), .B(n6824), .Z(n279) );
  NAND U529 ( .A(n6822), .B(n6823), .Z(n280) );
  NAND U530 ( .A(n279), .B(n280), .Z(n6971) );
  XOR U531 ( .A(n8093), .B(n8094), .Z(n8095) );
  NAND U532 ( .A(n9401), .B(n9400), .Z(n281) );
  NAND U533 ( .A(n9398), .B(n9399), .Z(n282) );
  NAND U534 ( .A(n281), .B(n282), .Z(n9461) );
  XOR U535 ( .A(n361), .B(n360), .Z(n283) );
  NANDN U536 ( .A(n359), .B(n283), .Z(n284) );
  NAND U537 ( .A(n361), .B(n360), .Z(n285) );
  AND U538 ( .A(n284), .B(n285), .Z(n373) );
  NAND U539 ( .A(n551), .B(n550), .Z(n286) );
  NANDN U540 ( .A(n549), .B(n548), .Z(n287) );
  NAND U541 ( .A(n286), .B(n287), .Z(n590) );
  NAND U542 ( .A(n767), .B(n766), .Z(n288) );
  NAND U543 ( .A(n764), .B(n765), .Z(n289) );
  NAND U544 ( .A(n288), .B(n289), .Z(n824) );
  NAND U545 ( .A(n1598), .B(n1597), .Z(n290) );
  NANDN U546 ( .A(n1596), .B(n1595), .Z(n291) );
  NAND U547 ( .A(n290), .B(n291), .Z(n1696) );
  NAND U548 ( .A(n7836), .B(n7835), .Z(n292) );
  XOR U549 ( .A(n7835), .B(n7836), .Z(n293) );
  NANDN U550 ( .A(n7837), .B(n293), .Z(n294) );
  NAND U551 ( .A(n292), .B(n294), .Z(n7976) );
  XOR U552 ( .A(n8226), .B(n8225), .Z(n295) );
  NANDN U553 ( .A(n8224), .B(n295), .Z(n296) );
  NAND U554 ( .A(n8226), .B(n8225), .Z(n297) );
  AND U555 ( .A(n296), .B(n297), .Z(n8345) );
  NAND U556 ( .A(n8686), .B(n8685), .Z(n298) );
  XOR U557 ( .A(n8685), .B(n8686), .Z(n299) );
  NANDN U558 ( .A(n8687), .B(n299), .Z(n300) );
  NAND U559 ( .A(n298), .B(n300), .Z(n8785) );
  NAND U560 ( .A(n8986), .B(n8984), .Z(n301) );
  XOR U561 ( .A(n8984), .B(n8986), .Z(n302) );
  NANDN U562 ( .A(n8985), .B(n302), .Z(n303) );
  NAND U563 ( .A(n301), .B(n303), .Z(n9077) );
  NAND U564 ( .A(n9084), .B(n9083), .Z(n304) );
  NANDN U565 ( .A(n9082), .B(n9081), .Z(n305) );
  AND U566 ( .A(n304), .B(n305), .Z(n9158) );
  NAND U567 ( .A(n9320), .B(n9319), .Z(n306) );
  XOR U568 ( .A(n9319), .B(n9320), .Z(n307) );
  NANDN U569 ( .A(n9321), .B(n307), .Z(n308) );
  NAND U570 ( .A(n306), .B(n308), .Z(n9394) );
  XOR U571 ( .A(n9645), .B(n9643), .Z(n309) );
  NANDN U572 ( .A(n9644), .B(n309), .Z(n310) );
  NAND U573 ( .A(n9645), .B(n9643), .Z(n311) );
  AND U574 ( .A(n310), .B(n311), .Z(n9697) );
  NAND U575 ( .A(n9830), .B(n9828), .Z(n312) );
  XOR U576 ( .A(n9828), .B(n9830), .Z(n313) );
  NANDN U577 ( .A(n9829), .B(n313), .Z(n314) );
  NAND U578 ( .A(n312), .B(n314), .Z(n9858) );
  IV U579 ( .A(b[0]), .Z(n315) );
  IV U580 ( .A(b[3]), .Z(n316) );
  IV U581 ( .A(b[5]), .Z(n317) );
  IV U582 ( .A(b[21]), .Z(n318) );
  IV U583 ( .A(b[23]), .Z(n319) );
  IV U584 ( .A(b[25]), .Z(n320) );
  IV U585 ( .A(b[27]), .Z(n321) );
  IV U586 ( .A(b[29]), .Z(n322) );
  IV U587 ( .A(b[31]), .Z(n323) );
  NANDN U588 ( .A(n315), .B(a[0]), .Z(n325) );
  XNOR U589 ( .A(n325), .B(sreg[32]), .Z(c[32]) );
  IV U590 ( .A(a[0]), .Z(n2616) );
  ANDN U591 ( .B(b[1]), .A(n2616), .Z(n324) );
  NANDN U592 ( .A(n315), .B(a[1]), .Z(n330) );
  XNOR U593 ( .A(n324), .B(n330), .Z(n333) );
  XNOR U594 ( .A(sreg[33]), .B(n333), .Z(n335) );
  NANDN U595 ( .A(n325), .B(sreg[32]), .Z(n334) );
  XOR U596 ( .A(n335), .B(n334), .Z(c[33]) );
  NANDN U597 ( .A(n315), .B(a[2]), .Z(n326) );
  XNOR U598 ( .A(b[1]), .B(n326), .Z(n328) );
  NANDN U599 ( .A(b[0]), .B(a[1]), .Z(n327) );
  AND U600 ( .A(n328), .B(n327), .Z(n338) );
  NANDN U601 ( .A(n2616), .B(b[2]), .Z(n329) );
  XNOR U602 ( .A(b[1]), .B(n329), .Z(n332) );
  OR U603 ( .A(n330), .B(a[0]), .Z(n331) );
  AND U604 ( .A(n332), .B(n331), .Z(n339) );
  XOR U605 ( .A(n338), .B(n339), .Z(n350) );
  NAND U606 ( .A(sreg[33]), .B(n333), .Z(n337) );
  OR U607 ( .A(n335), .B(n334), .Z(n336) );
  NAND U608 ( .A(n337), .B(n336), .Z(n349) );
  XNOR U609 ( .A(n349), .B(sreg[34]), .Z(n351) );
  XNOR U610 ( .A(n350), .B(n351), .Z(c[34]) );
  NAND U611 ( .A(n339), .B(n338), .Z(n361) );
  IV U612 ( .A(b[2]), .Z(n7756) );
  XNOR U613 ( .A(n7756), .B(b[1]), .Z(n7620) );
  XNOR U614 ( .A(n316), .B(a[0]), .Z(n342) );
  XNOR U615 ( .A(n316), .B(b[2]), .Z(n341) );
  XNOR U616 ( .A(n316), .B(b[1]), .Z(n340) );
  AND U617 ( .A(n341), .B(n340), .Z(n7622) );
  NAND U618 ( .A(n342), .B(n7622), .Z(n344) );
  XNOR U619 ( .A(n316), .B(a[1]), .Z(n362) );
  NAND U620 ( .A(n362), .B(n7620), .Z(n343) );
  NAND U621 ( .A(n344), .B(n343), .Z(n368) );
  NANDN U622 ( .A(n315), .B(a[3]), .Z(n345) );
  XNOR U623 ( .A(b[1]), .B(n345), .Z(n347) );
  IV U624 ( .A(a[2]), .Z(n2950) );
  NANDN U625 ( .A(n2950), .B(n315), .Z(n346) );
  AND U626 ( .A(n347), .B(n346), .Z(n369) );
  XOR U627 ( .A(n368), .B(n369), .Z(n359) );
  XNOR U628 ( .A(n360), .B(n359), .Z(n348) );
  XNOR U629 ( .A(n361), .B(n348), .Z(n354) );
  XNOR U630 ( .A(sreg[35]), .B(n354), .Z(n356) );
  NAND U631 ( .A(n349), .B(sreg[34]), .Z(n353) );
  NANDN U632 ( .A(n351), .B(n350), .Z(n352) );
  AND U633 ( .A(n353), .B(n352), .Z(n355) );
  XOR U634 ( .A(n356), .B(n355), .Z(c[35]) );
  NAND U635 ( .A(sreg[35]), .B(n354), .Z(n358) );
  OR U636 ( .A(n356), .B(n355), .Z(n357) );
  NAND U637 ( .A(n358), .B(n357), .Z(n391) );
  XNOR U638 ( .A(n391), .B(sreg[36]), .Z(n393) );
  NAND U639 ( .A(n362), .B(n7622), .Z(n364) );
  XNOR U640 ( .A(n316), .B(a[2]), .Z(n382) );
  NAND U641 ( .A(n382), .B(n7620), .Z(n363) );
  NAND U642 ( .A(n364), .B(n363), .Z(n385) );
  NANDN U643 ( .A(n315), .B(a[4]), .Z(n365) );
  XNOR U644 ( .A(b[1]), .B(n365), .Z(n367) );
  IV U645 ( .A(a[3]), .Z(n3094) );
  NANDN U646 ( .A(n3094), .B(n315), .Z(n366) );
  AND U647 ( .A(n367), .B(n366), .Z(n386) );
  XOR U648 ( .A(n385), .B(n386), .Z(n387) );
  XOR U649 ( .A(b[4]), .B(b[3]), .Z(n7905) );
  NANDN U650 ( .A(n2616), .B(n7905), .Z(n388) );
  XOR U651 ( .A(n387), .B(n388), .Z(n371) );
  NAND U652 ( .A(n369), .B(n368), .Z(n372) );
  XOR U653 ( .A(n371), .B(n372), .Z(n370) );
  XOR U654 ( .A(n373), .B(n370), .Z(n392) );
  XNOR U655 ( .A(n393), .B(n392), .Z(c[36]) );
  NANDN U656 ( .A(n315), .B(a[5]), .Z(n374) );
  XNOR U657 ( .A(b[1]), .B(n374), .Z(n376) );
  NANDN U658 ( .A(b[0]), .B(a[4]), .Z(n375) );
  AND U659 ( .A(n376), .B(n375), .Z(n402) );
  XNOR U660 ( .A(n317), .B(a[1]), .Z(n410) );
  AND U661 ( .A(n7905), .B(n410), .Z(n381) );
  XNOR U662 ( .A(n317), .B(a[0]), .Z(n379) );
  XNOR U663 ( .A(n317), .B(b[4]), .Z(n378) );
  XNOR U664 ( .A(n317), .B(b[3]), .Z(n377) );
  AND U665 ( .A(n378), .B(n377), .Z(n7906) );
  NAND U666 ( .A(n379), .B(n7906), .Z(n380) );
  NANDN U667 ( .A(n381), .B(n380), .Z(n403) );
  XNOR U668 ( .A(n402), .B(n403), .Z(n416) );
  XOR U669 ( .A(b[3]), .B(n3094), .Z(n404) );
  NANDN U670 ( .A(n404), .B(n7620), .Z(n384) );
  NAND U671 ( .A(n382), .B(n7622), .Z(n383) );
  AND U672 ( .A(n384), .B(n383), .Z(n413) );
  XNOR U673 ( .A(n414), .B(n413), .Z(n415) );
  XOR U674 ( .A(n416), .B(n415), .Z(n397) );
  NAND U675 ( .A(n386), .B(n385), .Z(n390) );
  NANDN U676 ( .A(n388), .B(n387), .Z(n389) );
  AND U677 ( .A(n390), .B(n389), .Z(n396) );
  XOR U678 ( .A(n397), .B(n396), .Z(n399) );
  XOR U679 ( .A(n398), .B(n399), .Z(n419) );
  XOR U680 ( .A(sreg[37]), .B(n419), .Z(n420) );
  NAND U681 ( .A(n391), .B(sreg[36]), .Z(n395) );
  NANDN U682 ( .A(n393), .B(n392), .Z(n394) );
  NAND U683 ( .A(n395), .B(n394), .Z(n421) );
  XOR U684 ( .A(n420), .B(n421), .Z(c[37]) );
  OR U685 ( .A(n397), .B(n396), .Z(n401) );
  NAND U686 ( .A(n399), .B(n398), .Z(n400) );
  NAND U687 ( .A(n401), .B(n400), .Z(n427) );
  NAND U688 ( .A(n403), .B(n402), .Z(n453) );
  NANDN U689 ( .A(n404), .B(n7622), .Z(n406) );
  XNOR U690 ( .A(n316), .B(a[4]), .Z(n435) );
  NAND U691 ( .A(n435), .B(n7620), .Z(n405) );
  NAND U692 ( .A(n406), .B(n405), .Z(n431) );
  XOR U693 ( .A(b[5]), .B(b[6]), .Z(n441) );
  AND U694 ( .A(a[0]), .B(n441), .Z(n447) );
  NANDN U695 ( .A(n315), .B(a[6]), .Z(n407) );
  XNOR U696 ( .A(b[1]), .B(n407), .Z(n409) );
  IV U697 ( .A(a[5]), .Z(n3389) );
  NANDN U698 ( .A(n3389), .B(n315), .Z(n408) );
  AND U699 ( .A(n409), .B(n408), .Z(n430) );
  XOR U700 ( .A(n447), .B(n430), .Z(n432) );
  XOR U701 ( .A(n431), .B(n432), .Z(n451) );
  XOR U702 ( .A(b[5]), .B(n2950), .Z(n438) );
  NANDN U703 ( .A(n438), .B(n7905), .Z(n412) );
  NAND U704 ( .A(n7906), .B(n410), .Z(n411) );
  NAND U705 ( .A(n412), .B(n411), .Z(n452) );
  XOR U706 ( .A(n451), .B(n452), .Z(n454) );
  XNOR U707 ( .A(n453), .B(n454), .Z(n424) );
  NANDN U708 ( .A(n414), .B(n413), .Z(n418) );
  NAND U709 ( .A(n416), .B(n415), .Z(n417) );
  NAND U710 ( .A(n418), .B(n417), .Z(n425) );
  XNOR U711 ( .A(n424), .B(n425), .Z(n426) );
  XNOR U712 ( .A(n427), .B(n426), .Z(n457) );
  OR U713 ( .A(n419), .B(sreg[37]), .Z(n423) );
  NANDN U714 ( .A(n421), .B(n420), .Z(n422) );
  AND U715 ( .A(n423), .B(n422), .Z(n455) );
  XNOR U716 ( .A(sreg[38]), .B(n455), .Z(n456) );
  XOR U717 ( .A(n457), .B(n456), .Z(c[38]) );
  NANDN U718 ( .A(n425), .B(n424), .Z(n429) );
  NAND U719 ( .A(n427), .B(n426), .Z(n428) );
  NAND U720 ( .A(n429), .B(n428), .Z(n468) );
  NAND U721 ( .A(n447), .B(n430), .Z(n434) );
  NAND U722 ( .A(n432), .B(n431), .Z(n433) );
  NAND U723 ( .A(n434), .B(n433), .Z(n473) );
  NAND U724 ( .A(n435), .B(n7622), .Z(n437) );
  XNOR U725 ( .A(n316), .B(a[5]), .Z(n486) );
  NAND U726 ( .A(n486), .B(n7620), .Z(n436) );
  NAND U727 ( .A(n437), .B(n436), .Z(n472) );
  XOR U728 ( .A(n317), .B(n3094), .Z(n494) );
  NAND U729 ( .A(n494), .B(n7905), .Z(n440) );
  NANDN U730 ( .A(n438), .B(n7906), .Z(n439) );
  NAND U731 ( .A(n440), .B(n439), .Z(n490) );
  XOR U732 ( .A(b[7]), .B(a[1]), .Z(n483) );
  IV U733 ( .A(n441), .Z(n8013) );
  ANDN U734 ( .B(n483), .A(n8013), .Z(n446) );
  XNOR U735 ( .A(b[7]), .B(n2616), .Z(n444) );
  XNOR U736 ( .A(b[7]), .B(n317), .Z(n443) );
  XOR U737 ( .A(b[7]), .B(b[6]), .Z(n442) );
  AND U738 ( .A(n443), .B(n442), .Z(n8014) );
  NAND U739 ( .A(n444), .B(n8014), .Z(n445) );
  NANDN U740 ( .A(n446), .B(n445), .Z(n489) );
  XNOR U741 ( .A(n490), .B(n489), .Z(n480) );
  NANDN U742 ( .A(n317), .B(b[6]), .Z(n8177) );
  NAND U743 ( .A(n8177), .B(b[7]), .Z(n8294) );
  NOR U744 ( .A(n8294), .B(n447), .Z(n477) );
  NANDN U745 ( .A(n315), .B(a[7]), .Z(n448) );
  XNOR U746 ( .A(b[1]), .B(n448), .Z(n450) );
  NANDN U747 ( .A(b[0]), .B(a[6]), .Z(n449) );
  AND U748 ( .A(n450), .B(n449), .Z(n478) );
  XOR U749 ( .A(n477), .B(n478), .Z(n479) );
  XOR U750 ( .A(n480), .B(n479), .Z(n471) );
  XOR U751 ( .A(n472), .B(n471), .Z(n474) );
  XNOR U752 ( .A(n473), .B(n474), .Z(n465) );
  XNOR U753 ( .A(n465), .B(n466), .Z(n467) );
  XOR U754 ( .A(n468), .B(n467), .Z(n460) );
  XNOR U755 ( .A(sreg[39]), .B(n460), .Z(n462) );
  NAND U756 ( .A(n455), .B(sreg[38]), .Z(n459) );
  OR U757 ( .A(n457), .B(n456), .Z(n458) );
  AND U758 ( .A(n459), .B(n458), .Z(n461) );
  XOR U759 ( .A(n462), .B(n461), .Z(c[39]) );
  NAND U760 ( .A(sreg[39]), .B(n460), .Z(n464) );
  OR U761 ( .A(n462), .B(n461), .Z(n463) );
  NAND U762 ( .A(n464), .B(n463), .Z(n538) );
  XNOR U763 ( .A(n538), .B(sreg[40]), .Z(n540) );
  NANDN U764 ( .A(n466), .B(n465), .Z(n470) );
  NAND U765 ( .A(n468), .B(n467), .Z(n469) );
  NAND U766 ( .A(n470), .B(n469), .Z(n500) );
  NANDN U767 ( .A(n472), .B(n471), .Z(n476) );
  OR U768 ( .A(n474), .B(n473), .Z(n475) );
  NAND U769 ( .A(n476), .B(n475), .Z(n498) );
  OR U770 ( .A(n478), .B(n477), .Z(n482) );
  NAND U771 ( .A(n480), .B(n479), .Z(n481) );
  NAND U772 ( .A(n482), .B(n481), .Z(n534) );
  XNOR U773 ( .A(b[7]), .B(a[2]), .Z(n514) );
  OR U774 ( .A(n514), .B(n8013), .Z(n485) );
  NAND U775 ( .A(n483), .B(n8014), .Z(n484) );
  NAND U776 ( .A(n485), .B(n484), .Z(n503) );
  XNOR U777 ( .A(b[3]), .B(a[6]), .Z(n523) );
  NANDN U778 ( .A(n523), .B(n7620), .Z(n488) );
  NAND U779 ( .A(n486), .B(n7622), .Z(n487) );
  AND U780 ( .A(n488), .B(n487), .Z(n504) );
  XNOR U781 ( .A(n503), .B(n504), .Z(n505) );
  NAND U782 ( .A(n490), .B(n489), .Z(n506) );
  XOR U783 ( .A(n505), .B(n506), .Z(n533) );
  XOR U784 ( .A(b[7]), .B(b[8]), .Z(n8288) );
  AND U785 ( .A(n8288), .B(a[0]), .Z(n529) );
  NANDN U786 ( .A(n315), .B(a[8]), .Z(n491) );
  XNOR U787 ( .A(b[1]), .B(n491), .Z(n493) );
  NANDN U788 ( .A(b[0]), .B(a[7]), .Z(n492) );
  AND U789 ( .A(n493), .B(n492), .Z(n527) );
  XNOR U790 ( .A(b[5]), .B(a[4]), .Z(n517) );
  NANDN U791 ( .A(n517), .B(n7905), .Z(n496) );
  NAND U792 ( .A(n7906), .B(n494), .Z(n495) );
  AND U793 ( .A(n496), .B(n495), .Z(n526) );
  XNOR U794 ( .A(n527), .B(n526), .Z(n528) );
  XNOR U795 ( .A(n529), .B(n528), .Z(n532) );
  XNOR U796 ( .A(n533), .B(n532), .Z(n535) );
  XNOR U797 ( .A(n534), .B(n535), .Z(n497) );
  XNOR U798 ( .A(n498), .B(n497), .Z(n499) );
  XOR U799 ( .A(n500), .B(n499), .Z(n539) );
  XOR U800 ( .A(n540), .B(n539), .Z(c[40]) );
  NAND U801 ( .A(n498), .B(n497), .Z(n502) );
  OR U802 ( .A(n500), .B(n499), .Z(n501) );
  NAND U803 ( .A(n502), .B(n501), .Z(n551) );
  NANDN U804 ( .A(n504), .B(n503), .Z(n508) );
  NANDN U805 ( .A(n506), .B(n505), .Z(n507) );
  NAND U806 ( .A(n508), .B(n507), .Z(n555) );
  XNOR U807 ( .A(b[9]), .B(n2616), .Z(n511) );
  XOR U808 ( .A(b[9]), .B(b[7]), .Z(n510) );
  XOR U809 ( .A(b[9]), .B(b[8]), .Z(n509) );
  AND U810 ( .A(n510), .B(n509), .Z(n8286) );
  NAND U811 ( .A(n511), .B(n8286), .Z(n513) );
  XOR U812 ( .A(b[9]), .B(a[1]), .Z(n570) );
  NAND U813 ( .A(n570), .B(n8288), .Z(n512) );
  NAND U814 ( .A(n513), .B(n512), .Z(n576) );
  XNOR U815 ( .A(b[7]), .B(a[3]), .Z(n584) );
  OR U816 ( .A(n584), .B(n8013), .Z(n516) );
  NANDN U817 ( .A(n514), .B(n8014), .Z(n515) );
  AND U818 ( .A(n516), .B(n515), .Z(n577) );
  XNOR U819 ( .A(n576), .B(n577), .Z(n561) );
  NAND U820 ( .A(b[7]), .B(b[8]), .Z(n8416) );
  NAND U821 ( .A(n8416), .B(b[9]), .Z(n8596) );
  OR U822 ( .A(n529), .B(n8596), .Z(n558) );
  XOR U823 ( .A(b[5]), .B(n3389), .Z(n573) );
  NANDN U824 ( .A(n573), .B(n7905), .Z(n519) );
  NANDN U825 ( .A(n517), .B(n7906), .Z(n518) );
  NAND U826 ( .A(n519), .B(n518), .Z(n559) );
  XOR U827 ( .A(n558), .B(n559), .Z(n560) );
  XOR U828 ( .A(n561), .B(n560), .Z(n566) );
  NANDN U829 ( .A(n315), .B(a[9]), .Z(n520) );
  XNOR U830 ( .A(b[1]), .B(n520), .Z(n522) );
  IV U831 ( .A(a[8]), .Z(n3831) );
  NANDN U832 ( .A(n3831), .B(n315), .Z(n521) );
  AND U833 ( .A(n522), .B(n521), .Z(n564) );
  XNOR U834 ( .A(b[3]), .B(a[7]), .Z(n578) );
  NANDN U835 ( .A(n578), .B(n7620), .Z(n525) );
  NANDN U836 ( .A(n523), .B(n7622), .Z(n524) );
  AND U837 ( .A(n525), .B(n524), .Z(n565) );
  XOR U838 ( .A(n564), .B(n565), .Z(n567) );
  XOR U839 ( .A(n566), .B(n567), .Z(n552) );
  NANDN U840 ( .A(n527), .B(n526), .Z(n531) );
  NANDN U841 ( .A(n529), .B(n528), .Z(n530) );
  AND U842 ( .A(n531), .B(n530), .Z(n553) );
  XOR U843 ( .A(n552), .B(n553), .Z(n554) );
  XNOR U844 ( .A(n555), .B(n554), .Z(n548) );
  NAND U845 ( .A(n533), .B(n532), .Z(n537) );
  NANDN U846 ( .A(n535), .B(n534), .Z(n536) );
  AND U847 ( .A(n537), .B(n536), .Z(n549) );
  XNOR U848 ( .A(n548), .B(n549), .Z(n550) );
  XNOR U849 ( .A(n551), .B(n550), .Z(n543) );
  XNOR U850 ( .A(n543), .B(sreg[41]), .Z(n545) );
  NAND U851 ( .A(n538), .B(sreg[40]), .Z(n542) );
  OR U852 ( .A(n540), .B(n539), .Z(n541) );
  AND U853 ( .A(n542), .B(n541), .Z(n544) );
  XOR U854 ( .A(n545), .B(n544), .Z(c[41]) );
  NAND U855 ( .A(n543), .B(sreg[41]), .Z(n547) );
  OR U856 ( .A(n545), .B(n544), .Z(n546) );
  NAND U857 ( .A(n547), .B(n546), .Z(n635) );
  XNOR U858 ( .A(n635), .B(sreg[42]), .Z(n637) );
  NAND U859 ( .A(n553), .B(n552), .Z(n557) );
  NAND U860 ( .A(n555), .B(n554), .Z(n556) );
  NAND U861 ( .A(n557), .B(n556), .Z(n587) );
  NANDN U862 ( .A(n559), .B(n558), .Z(n563) );
  OR U863 ( .A(n561), .B(n560), .Z(n562) );
  NAND U864 ( .A(n563), .B(n562), .Z(n596) );
  NANDN U865 ( .A(n565), .B(n564), .Z(n569) );
  OR U866 ( .A(n567), .B(n566), .Z(n568) );
  NAND U867 ( .A(n569), .B(n568), .Z(n594) );
  NAND U868 ( .A(n570), .B(n8286), .Z(n572) );
  XNOR U869 ( .A(b[9]), .B(n2950), .Z(n621) );
  NAND U870 ( .A(n621), .B(n8288), .Z(n571) );
  NAND U871 ( .A(n572), .B(n571), .Z(n608) );
  XNOR U872 ( .A(n317), .B(a[6]), .Z(n632) );
  NAND U873 ( .A(n632), .B(n7905), .Z(n575) );
  NANDN U874 ( .A(n573), .B(n7906), .Z(n574) );
  AND U875 ( .A(n575), .B(n574), .Z(n609) );
  XOR U876 ( .A(n608), .B(n609), .Z(n611) );
  NANDN U877 ( .A(n577), .B(n576), .Z(n610) );
  XNOR U878 ( .A(n611), .B(n610), .Z(n597) );
  NANDN U879 ( .A(n578), .B(n7622), .Z(n580) );
  XNOR U880 ( .A(n316), .B(a[8]), .Z(n618) );
  NAND U881 ( .A(n618), .B(n7620), .Z(n579) );
  NAND U882 ( .A(n580), .B(n579), .Z(n598) );
  XNOR U883 ( .A(n597), .B(n598), .Z(n599) );
  XOR U884 ( .A(b[9]), .B(b[10]), .Z(n8541) );
  AND U885 ( .A(n8541), .B(a[0]), .Z(n617) );
  NANDN U886 ( .A(n315), .B(a[10]), .Z(n581) );
  XNOR U887 ( .A(b[1]), .B(n581), .Z(n583) );
  NANDN U888 ( .A(b[0]), .B(a[9]), .Z(n582) );
  AND U889 ( .A(n583), .B(n582), .Z(n604) );
  XNOR U890 ( .A(b[7]), .B(a[4]), .Z(n614) );
  OR U891 ( .A(n614), .B(n8013), .Z(n586) );
  NANDN U892 ( .A(n584), .B(n8014), .Z(n585) );
  AND U893 ( .A(n586), .B(n585), .Z(n603) );
  XNOR U894 ( .A(n604), .B(n603), .Z(n605) );
  XNOR U895 ( .A(n617), .B(n605), .Z(n600) );
  XOR U896 ( .A(n599), .B(n600), .Z(n593) );
  XNOR U897 ( .A(n594), .B(n593), .Z(n595) );
  XNOR U898 ( .A(n596), .B(n595), .Z(n588) );
  XOR U899 ( .A(n587), .B(n588), .Z(n589) );
  XOR U900 ( .A(n590), .B(n589), .Z(n636) );
  XOR U901 ( .A(n637), .B(n636), .Z(c[42]) );
  OR U902 ( .A(n588), .B(n587), .Z(n592) );
  NAND U903 ( .A(n590), .B(n589), .Z(n591) );
  NAND U904 ( .A(n592), .B(n591), .Z(n648) );
  NANDN U905 ( .A(n598), .B(n597), .Z(n602) );
  NAND U906 ( .A(n600), .B(n599), .Z(n601) );
  NAND U907 ( .A(n602), .B(n601), .Z(n654) );
  NANDN U908 ( .A(n604), .B(n603), .Z(n607) );
  NANDN U909 ( .A(n617), .B(n605), .Z(n606) );
  NAND U910 ( .A(n607), .B(n606), .Z(n651) );
  NANDN U911 ( .A(n609), .B(n608), .Z(n613) );
  OR U912 ( .A(n611), .B(n610), .Z(n612) );
  NAND U913 ( .A(n613), .B(n612), .Z(n692) );
  XOR U914 ( .A(b[7]), .B(n3389), .Z(n674) );
  OR U915 ( .A(n674), .B(n8013), .Z(n616) );
  NANDN U916 ( .A(n614), .B(n8014), .Z(n615) );
  NAND U917 ( .A(n616), .B(n615), .Z(n660) );
  NAND U918 ( .A(b[9]), .B(b[10]), .Z(n8642) );
  NAND U919 ( .A(n8642), .B(b[11]), .Z(n8852) );
  NOR U920 ( .A(n617), .B(n8852), .Z(n658) );
  XNOR U921 ( .A(b[3]), .B(a[9]), .Z(n671) );
  NANDN U922 ( .A(n671), .B(n7620), .Z(n620) );
  NAND U923 ( .A(n618), .B(n7622), .Z(n619) );
  AND U924 ( .A(n620), .B(n619), .Z(n657) );
  XOR U925 ( .A(n658), .B(n657), .Z(n659) );
  XNOR U926 ( .A(n660), .B(n659), .Z(n689) );
  XNOR U927 ( .A(b[9]), .B(n3094), .Z(n677) );
  NAND U928 ( .A(n677), .B(n8288), .Z(n623) );
  NAND U929 ( .A(n621), .B(n8286), .Z(n622) );
  AND U930 ( .A(n623), .B(n622), .Z(n670) );
  XNOR U931 ( .A(b[11]), .B(n2616), .Z(n626) );
  XOR U932 ( .A(b[11]), .B(b[9]), .Z(n625) );
  XOR U933 ( .A(b[11]), .B(b[10]), .Z(n624) );
  AND U934 ( .A(n625), .B(n624), .Z(n8542) );
  NAND U935 ( .A(n626), .B(n8542), .Z(n628) );
  XOR U936 ( .A(b[11]), .B(a[1]), .Z(n666) );
  AND U937 ( .A(n8541), .B(n666), .Z(n627) );
  ANDN U938 ( .B(n628), .A(n627), .Z(n669) );
  XNOR U939 ( .A(n670), .B(n669), .Z(n686) );
  NANDN U940 ( .A(n315), .B(a[11]), .Z(n629) );
  XNOR U941 ( .A(b[1]), .B(n629), .Z(n631) );
  NANDN U942 ( .A(b[0]), .B(a[10]), .Z(n630) );
  AND U943 ( .A(n631), .B(n630), .Z(n684) );
  XOR U944 ( .A(n317), .B(a[7]), .Z(n663) );
  NANDN U945 ( .A(n663), .B(n7905), .Z(n634) );
  NAND U946 ( .A(n7906), .B(n632), .Z(n633) );
  AND U947 ( .A(n634), .B(n633), .Z(n683) );
  XNOR U948 ( .A(n684), .B(n683), .Z(n685) );
  XOR U949 ( .A(n686), .B(n685), .Z(n690) );
  XNOR U950 ( .A(n689), .B(n690), .Z(n691) );
  XOR U951 ( .A(n692), .B(n691), .Z(n652) );
  XNOR U952 ( .A(n651), .B(n652), .Z(n653) );
  XNOR U953 ( .A(n654), .B(n653), .Z(n646) );
  XNOR U954 ( .A(n645), .B(n646), .Z(n647) );
  XNOR U955 ( .A(n648), .B(n647), .Z(n640) );
  XNOR U956 ( .A(n640), .B(sreg[43]), .Z(n642) );
  NAND U957 ( .A(n635), .B(sreg[42]), .Z(n639) );
  OR U958 ( .A(n637), .B(n636), .Z(n638) );
  AND U959 ( .A(n639), .B(n638), .Z(n641) );
  XOR U960 ( .A(n642), .B(n641), .Z(c[43]) );
  NAND U961 ( .A(n640), .B(sreg[43]), .Z(n644) );
  OR U962 ( .A(n642), .B(n641), .Z(n643) );
  NAND U963 ( .A(n644), .B(n643), .Z(n754) );
  XNOR U964 ( .A(n754), .B(sreg[44]), .Z(n756) );
  NANDN U965 ( .A(n646), .B(n645), .Z(n650) );
  NAND U966 ( .A(n648), .B(n647), .Z(n649) );
  NAND U967 ( .A(n650), .B(n649), .Z(n698) );
  NANDN U968 ( .A(n652), .B(n651), .Z(n656) );
  NAND U969 ( .A(n654), .B(n653), .Z(n655) );
  NAND U970 ( .A(n656), .B(n655), .Z(n695) );
  NANDN U971 ( .A(n658), .B(n657), .Z(n662) );
  OR U972 ( .A(n660), .B(n659), .Z(n661) );
  NAND U973 ( .A(n662), .B(n661), .Z(n704) );
  XOR U974 ( .A(n317), .B(a[8]), .Z(n737) );
  NANDN U975 ( .A(n737), .B(n7905), .Z(n665) );
  NANDN U976 ( .A(n663), .B(n7906), .Z(n664) );
  NAND U977 ( .A(n665), .B(n664), .Z(n714) );
  XNOR U978 ( .A(b[11]), .B(a[2]), .Z(n740) );
  NANDN U979 ( .A(n740), .B(n8541), .Z(n668) );
  NAND U980 ( .A(n8542), .B(n666), .Z(n667) );
  AND U981 ( .A(n668), .B(n667), .Z(n713) );
  XNOR U982 ( .A(n714), .B(n713), .Z(n715) );
  OR U983 ( .A(n670), .B(n669), .Z(n722) );
  NANDN U984 ( .A(n671), .B(n7622), .Z(n673) );
  XNOR U985 ( .A(n316), .B(a[10]), .Z(n731) );
  NAND U986 ( .A(n731), .B(n7620), .Z(n672) );
  NAND U987 ( .A(n673), .B(n672), .Z(n720) );
  XNOR U988 ( .A(b[7]), .B(a[6]), .Z(n751) );
  OR U989 ( .A(n751), .B(n8013), .Z(n676) );
  NANDN U990 ( .A(n674), .B(n8014), .Z(n675) );
  AND U991 ( .A(n676), .B(n675), .Z(n719) );
  XNOR U992 ( .A(n720), .B(n719), .Z(n721) );
  XNOR U993 ( .A(n722), .B(n721), .Z(n716) );
  XOR U994 ( .A(n715), .B(n716), .Z(n710) );
  XOR U995 ( .A(b[11]), .B(b[12]), .Z(n8730) );
  AND U996 ( .A(n8730), .B(a[0]), .Z(n730) );
  XOR U997 ( .A(b[9]), .B(a[4]), .Z(n734) );
  NAND U998 ( .A(n734), .B(n8288), .Z(n679) );
  NAND U999 ( .A(n677), .B(n8286), .Z(n678) );
  AND U1000 ( .A(n679), .B(n678), .Z(n726) );
  NANDN U1001 ( .A(n315), .B(a[12]), .Z(n680) );
  XNOR U1002 ( .A(b[1]), .B(n680), .Z(n682) );
  NANDN U1003 ( .A(b[0]), .B(a[11]), .Z(n681) );
  AND U1004 ( .A(n682), .B(n681), .Z(n725) );
  XOR U1005 ( .A(n726), .B(n725), .Z(n727) );
  XOR U1006 ( .A(n730), .B(n727), .Z(n708) );
  NANDN U1007 ( .A(n684), .B(n683), .Z(n688) );
  NAND U1008 ( .A(n686), .B(n685), .Z(n687) );
  AND U1009 ( .A(n688), .B(n687), .Z(n707) );
  XNOR U1010 ( .A(n708), .B(n707), .Z(n709) );
  XNOR U1011 ( .A(n710), .B(n709), .Z(n701) );
  NANDN U1012 ( .A(n690), .B(n689), .Z(n694) );
  NAND U1013 ( .A(n692), .B(n691), .Z(n693) );
  NAND U1014 ( .A(n694), .B(n693), .Z(n702) );
  XNOR U1015 ( .A(n701), .B(n702), .Z(n703) );
  XNOR U1016 ( .A(n704), .B(n703), .Z(n696) );
  XNOR U1017 ( .A(n695), .B(n696), .Z(n697) );
  XOR U1018 ( .A(n698), .B(n697), .Z(n755) );
  XOR U1019 ( .A(n756), .B(n755), .Z(c[44]) );
  NANDN U1020 ( .A(n696), .B(n695), .Z(n700) );
  NAND U1021 ( .A(n698), .B(n697), .Z(n699) );
  NAND U1022 ( .A(n700), .B(n699), .Z(n767) );
  NANDN U1023 ( .A(n702), .B(n701), .Z(n706) );
  NAND U1024 ( .A(n704), .B(n703), .Z(n705) );
  NAND U1025 ( .A(n706), .B(n705), .Z(n765) );
  NANDN U1026 ( .A(n708), .B(n707), .Z(n712) );
  NAND U1027 ( .A(n710), .B(n709), .Z(n711) );
  NAND U1028 ( .A(n712), .B(n711), .Z(n771) );
  NANDN U1029 ( .A(n714), .B(n713), .Z(n718) );
  NANDN U1030 ( .A(n716), .B(n715), .Z(n717) );
  NAND U1031 ( .A(n718), .B(n717), .Z(n769) );
  NANDN U1032 ( .A(n720), .B(n719), .Z(n724) );
  NAND U1033 ( .A(n722), .B(n721), .Z(n723) );
  NAND U1034 ( .A(n724), .B(n723), .Z(n815) );
  NANDN U1035 ( .A(n726), .B(n725), .Z(n729) );
  NANDN U1036 ( .A(n727), .B(n730), .Z(n728) );
  NAND U1037 ( .A(n729), .B(n728), .Z(n816) );
  XNOR U1038 ( .A(n815), .B(n816), .Z(n817) );
  NAND U1039 ( .A(b[11]), .B(b[12]), .Z(n8795) );
  NAND U1040 ( .A(n8795), .B(b[13]), .Z(n8960) );
  IV U1041 ( .A(n8960), .Z(n9009) );
  NANDN U1042 ( .A(n730), .B(n9009), .Z(n791) );
  NAND U1043 ( .A(n731), .B(n7622), .Z(n733) );
  XNOR U1044 ( .A(n316), .B(a[11]), .Z(n806) );
  NAND U1045 ( .A(n806), .B(n7620), .Z(n732) );
  NAND U1046 ( .A(n733), .B(n732), .Z(n788) );
  NAND U1047 ( .A(n734), .B(n8286), .Z(n736) );
  XNOR U1048 ( .A(b[9]), .B(n3389), .Z(n776) );
  NAND U1049 ( .A(n776), .B(n8288), .Z(n735) );
  NAND U1050 ( .A(n736), .B(n735), .Z(n789) );
  XOR U1051 ( .A(n788), .B(n789), .Z(n790) );
  XOR U1052 ( .A(n791), .B(n790), .Z(n809) );
  XNOR U1053 ( .A(b[5]), .B(a[9]), .Z(n800) );
  NANDN U1054 ( .A(n800), .B(n7905), .Z(n739) );
  NANDN U1055 ( .A(n737), .B(n7906), .Z(n738) );
  NAND U1056 ( .A(n739), .B(n738), .Z(n810) );
  XNOR U1057 ( .A(n809), .B(n810), .Z(n811) );
  XNOR U1058 ( .A(b[11]), .B(a[3]), .Z(n797) );
  NANDN U1059 ( .A(n797), .B(n8541), .Z(n742) );
  NANDN U1060 ( .A(n740), .B(n8542), .Z(n741) );
  NAND U1061 ( .A(n742), .B(n741), .Z(n775) );
  XOR U1062 ( .A(b[13]), .B(a[1]), .Z(n779) );
  AND U1063 ( .A(n8730), .B(n779), .Z(n747) );
  XNOR U1064 ( .A(b[13]), .B(n2616), .Z(n745) );
  XOR U1065 ( .A(b[13]), .B(b[11]), .Z(n744) );
  XOR U1066 ( .A(b[13]), .B(b[12]), .Z(n743) );
  AND U1067 ( .A(n744), .B(n743), .Z(n8731) );
  NAND U1068 ( .A(n745), .B(n8731), .Z(n746) );
  NANDN U1069 ( .A(n747), .B(n746), .Z(n774) );
  XNOR U1070 ( .A(n775), .B(n774), .Z(n785) );
  NANDN U1071 ( .A(n315), .B(a[13]), .Z(n748) );
  XNOR U1072 ( .A(b[1]), .B(n748), .Z(n750) );
  NANDN U1073 ( .A(b[0]), .B(a[12]), .Z(n749) );
  AND U1074 ( .A(n750), .B(n749), .Z(n783) );
  XOR U1075 ( .A(b[7]), .B(a[7]), .Z(n803) );
  NANDN U1076 ( .A(n8013), .B(n803), .Z(n753) );
  NANDN U1077 ( .A(n751), .B(n8014), .Z(n752) );
  AND U1078 ( .A(n753), .B(n752), .Z(n782) );
  XNOR U1079 ( .A(n783), .B(n782), .Z(n784) );
  XOR U1080 ( .A(n785), .B(n784), .Z(n812) );
  XOR U1081 ( .A(n811), .B(n812), .Z(n818) );
  XOR U1082 ( .A(n817), .B(n818), .Z(n768) );
  XOR U1083 ( .A(n769), .B(n768), .Z(n770) );
  XNOR U1084 ( .A(n771), .B(n770), .Z(n764) );
  XOR U1085 ( .A(n765), .B(n764), .Z(n766) );
  XNOR U1086 ( .A(n767), .B(n766), .Z(n759) );
  XNOR U1087 ( .A(n759), .B(sreg[45]), .Z(n761) );
  NAND U1088 ( .A(n754), .B(sreg[44]), .Z(n758) );
  OR U1089 ( .A(n756), .B(n755), .Z(n757) );
  AND U1090 ( .A(n758), .B(n757), .Z(n760) );
  XOR U1091 ( .A(n761), .B(n760), .Z(c[45]) );
  NAND U1092 ( .A(n759), .B(sreg[45]), .Z(n763) );
  OR U1093 ( .A(n761), .B(n760), .Z(n762) );
  NAND U1094 ( .A(n763), .B(n762), .Z(n887) );
  XNOR U1095 ( .A(n887), .B(sreg[46]), .Z(n889) );
  NAND U1096 ( .A(n769), .B(n768), .Z(n773) );
  NANDN U1097 ( .A(n771), .B(n770), .Z(n772) );
  NAND U1098 ( .A(n773), .B(n772), .Z(n821) );
  NAND U1099 ( .A(n775), .B(n774), .Z(n835) );
  NAND U1100 ( .A(n776), .B(n8286), .Z(n778) );
  XOR U1101 ( .A(b[9]), .B(a[6]), .Z(n857) );
  NAND U1102 ( .A(n857), .B(n8288), .Z(n777) );
  NAND U1103 ( .A(n778), .B(n777), .Z(n834) );
  XNOR U1104 ( .A(b[13]), .B(a[2]), .Z(n865) );
  NANDN U1105 ( .A(n865), .B(n8730), .Z(n781) );
  NAND U1106 ( .A(n8731), .B(n779), .Z(n780) );
  AND U1107 ( .A(n781), .B(n780), .Z(n833) );
  XNOR U1108 ( .A(n834), .B(n833), .Z(n836) );
  XNOR U1109 ( .A(n835), .B(n836), .Z(n848) );
  NANDN U1110 ( .A(n783), .B(n782), .Z(n787) );
  NAND U1111 ( .A(n785), .B(n784), .Z(n786) );
  NAND U1112 ( .A(n787), .B(n786), .Z(n849) );
  XOR U1113 ( .A(n848), .B(n849), .Z(n851) );
  NAND U1114 ( .A(n789), .B(n788), .Z(n793) );
  NANDN U1115 ( .A(n791), .B(n790), .Z(n792) );
  NAND U1116 ( .A(n793), .B(n792), .Z(n845) );
  XOR U1117 ( .A(b[13]), .B(b[14]), .Z(n8963) );
  AND U1118 ( .A(n8963), .B(a[0]), .Z(n883) );
  NANDN U1119 ( .A(n315), .B(a[14]), .Z(n794) );
  XNOR U1120 ( .A(b[1]), .B(n794), .Z(n796) );
  IV U1121 ( .A(a[13]), .Z(n4578) );
  NANDN U1122 ( .A(n4578), .B(n315), .Z(n795) );
  AND U1123 ( .A(n796), .B(n795), .Z(n838) );
  XOR U1124 ( .A(b[11]), .B(a[4]), .Z(n874) );
  NAND U1125 ( .A(n8541), .B(n874), .Z(n799) );
  NANDN U1126 ( .A(n797), .B(n8542), .Z(n798) );
  AND U1127 ( .A(n799), .B(n798), .Z(n837) );
  XNOR U1128 ( .A(n838), .B(n837), .Z(n839) );
  XNOR U1129 ( .A(n883), .B(n839), .Z(n842) );
  XNOR U1130 ( .A(b[5]), .B(a[10]), .Z(n880) );
  NANDN U1131 ( .A(n880), .B(n7905), .Z(n802) );
  NANDN U1132 ( .A(n800), .B(n7906), .Z(n801) );
  NAND U1133 ( .A(n802), .B(n801), .Z(n871) );
  XNOR U1134 ( .A(b[7]), .B(n3831), .Z(n884) );
  NANDN U1135 ( .A(n8013), .B(n884), .Z(n805) );
  NAND U1136 ( .A(n803), .B(n8014), .Z(n804) );
  NAND U1137 ( .A(n805), .B(n804), .Z(n868) );
  XNOR U1138 ( .A(b[3]), .B(a[12]), .Z(n877) );
  NANDN U1139 ( .A(n877), .B(n7620), .Z(n808) );
  NAND U1140 ( .A(n806), .B(n7622), .Z(n807) );
  AND U1141 ( .A(n808), .B(n807), .Z(n869) );
  XNOR U1142 ( .A(n868), .B(n869), .Z(n870) );
  XNOR U1143 ( .A(n871), .B(n870), .Z(n843) );
  XOR U1144 ( .A(n842), .B(n843), .Z(n844) );
  XNOR U1145 ( .A(n845), .B(n844), .Z(n850) );
  XNOR U1146 ( .A(n851), .B(n850), .Z(n830) );
  NANDN U1147 ( .A(n810), .B(n809), .Z(n814) );
  NAND U1148 ( .A(n812), .B(n811), .Z(n813) );
  NAND U1149 ( .A(n814), .B(n813), .Z(n827) );
  NANDN U1150 ( .A(n816), .B(n815), .Z(n820) );
  NAND U1151 ( .A(n818), .B(n817), .Z(n819) );
  AND U1152 ( .A(n820), .B(n819), .Z(n828) );
  XNOR U1153 ( .A(n827), .B(n828), .Z(n829) );
  XNOR U1154 ( .A(n830), .B(n829), .Z(n822) );
  XNOR U1155 ( .A(n821), .B(n822), .Z(n823) );
  XOR U1156 ( .A(n824), .B(n823), .Z(n888) );
  XOR U1157 ( .A(n889), .B(n888), .Z(c[46]) );
  NANDN U1158 ( .A(n822), .B(n821), .Z(n826) );
  NAND U1159 ( .A(n824), .B(n823), .Z(n825) );
  NAND U1160 ( .A(n826), .B(n825), .Z(n900) );
  NANDN U1161 ( .A(n828), .B(n827), .Z(n832) );
  NAND U1162 ( .A(n830), .B(n829), .Z(n831) );
  NAND U1163 ( .A(n832), .B(n831), .Z(n897) );
  NANDN U1164 ( .A(n838), .B(n837), .Z(n841) );
  NANDN U1165 ( .A(n883), .B(n839), .Z(n840) );
  AND U1166 ( .A(n841), .B(n840), .Z(n904) );
  XNOR U1167 ( .A(n903), .B(n904), .Z(n905) );
  OR U1168 ( .A(n843), .B(n842), .Z(n847) );
  NAND U1169 ( .A(n845), .B(n844), .Z(n846) );
  NAND U1170 ( .A(n847), .B(n846), .Z(n906) );
  XOR U1171 ( .A(n905), .B(n906), .Z(n954) );
  NANDN U1172 ( .A(n849), .B(n848), .Z(n853) );
  OR U1173 ( .A(n851), .B(n850), .Z(n852) );
  NAND U1174 ( .A(n853), .B(n852), .Z(n951) );
  NANDN U1175 ( .A(n315), .B(a[15]), .Z(n854) );
  XNOR U1176 ( .A(b[1]), .B(n854), .Z(n856) );
  NANDN U1177 ( .A(b[0]), .B(a[14]), .Z(n855) );
  AND U1178 ( .A(n856), .B(n855), .Z(n919) );
  XOR U1179 ( .A(b[9]), .B(a[7]), .Z(n932) );
  NAND U1180 ( .A(n932), .B(n8288), .Z(n859) );
  NAND U1181 ( .A(n857), .B(n8286), .Z(n858) );
  AND U1182 ( .A(n859), .B(n858), .Z(n920) );
  XNOR U1183 ( .A(n919), .B(n920), .Z(n921) );
  XNOR U1184 ( .A(b[15]), .B(n2616), .Z(n862) );
  XOR U1185 ( .A(b[15]), .B(b[13]), .Z(n861) );
  XOR U1186 ( .A(b[15]), .B(b[14]), .Z(n860) );
  AND U1187 ( .A(n861), .B(n860), .Z(n8961) );
  NAND U1188 ( .A(n862), .B(n8961), .Z(n864) );
  XOR U1189 ( .A(b[15]), .B(a[1]), .Z(n944) );
  NAND U1190 ( .A(n944), .B(n8963), .Z(n863) );
  NAND U1191 ( .A(n864), .B(n863), .Z(n927) );
  XNOR U1192 ( .A(b[13]), .B(a[3]), .Z(n916) );
  NANDN U1193 ( .A(n916), .B(n8730), .Z(n867) );
  NANDN U1194 ( .A(n865), .B(n8731), .Z(n866) );
  AND U1195 ( .A(n867), .B(n866), .Z(n928) );
  XOR U1196 ( .A(n927), .B(n928), .Z(n922) );
  XOR U1197 ( .A(n921), .B(n922), .Z(n947) );
  NANDN U1198 ( .A(n869), .B(n868), .Z(n873) );
  NAND U1199 ( .A(n871), .B(n870), .Z(n872) );
  NAND U1200 ( .A(n873), .B(n872), .Z(n948) );
  XNOR U1201 ( .A(n947), .B(n948), .Z(n949) );
  XNOR U1202 ( .A(b[11]), .B(n3389), .Z(n938) );
  NAND U1203 ( .A(n938), .B(n8541), .Z(n876) );
  NAND U1204 ( .A(n874), .B(n8542), .Z(n875) );
  NAND U1205 ( .A(n876), .B(n875), .Z(n912) );
  NANDN U1206 ( .A(n877), .B(n7622), .Z(n879) );
  XNOR U1207 ( .A(n316), .B(a[13]), .Z(n929) );
  NAND U1208 ( .A(n929), .B(n7620), .Z(n878) );
  NAND U1209 ( .A(n879), .B(n878), .Z(n909) );
  XNOR U1210 ( .A(n317), .B(a[11]), .Z(n941) );
  NAND U1211 ( .A(n941), .B(n7905), .Z(n882) );
  NANDN U1212 ( .A(n880), .B(n7906), .Z(n881) );
  AND U1213 ( .A(n882), .B(n881), .Z(n910) );
  XNOR U1214 ( .A(n909), .B(n910), .Z(n911) );
  XNOR U1215 ( .A(n912), .B(n911), .Z(n926) );
  NAND U1216 ( .A(b[13]), .B(b[14]), .Z(n9021) );
  NAND U1217 ( .A(n9021), .B(b[15]), .Z(n9207) );
  OR U1218 ( .A(n883), .B(n9207), .Z(n923) );
  XOR U1219 ( .A(b[7]), .B(a[9]), .Z(n935) );
  NANDN U1220 ( .A(n8013), .B(n935), .Z(n886) );
  NAND U1221 ( .A(n8014), .B(n884), .Z(n885) );
  NAND U1222 ( .A(n886), .B(n885), .Z(n924) );
  XNOR U1223 ( .A(n923), .B(n924), .Z(n925) );
  XOR U1224 ( .A(n926), .B(n925), .Z(n950) );
  XOR U1225 ( .A(n949), .B(n950), .Z(n952) );
  XNOR U1226 ( .A(n951), .B(n952), .Z(n953) );
  XOR U1227 ( .A(n954), .B(n953), .Z(n898) );
  XNOR U1228 ( .A(n897), .B(n898), .Z(n899) );
  XNOR U1229 ( .A(n900), .B(n899), .Z(n892) );
  XNOR U1230 ( .A(n892), .B(sreg[47]), .Z(n894) );
  NAND U1231 ( .A(n887), .B(sreg[46]), .Z(n891) );
  OR U1232 ( .A(n889), .B(n888), .Z(n890) );
  AND U1233 ( .A(n891), .B(n890), .Z(n893) );
  XOR U1234 ( .A(n894), .B(n893), .Z(c[47]) );
  NAND U1235 ( .A(n892), .B(sreg[47]), .Z(n896) );
  OR U1236 ( .A(n894), .B(n893), .Z(n895) );
  NAND U1237 ( .A(n896), .B(n895), .Z(n1030) );
  XNOR U1238 ( .A(n1030), .B(sreg[48]), .Z(n1032) );
  NANDN U1239 ( .A(n898), .B(n897), .Z(n902) );
  NAND U1240 ( .A(n900), .B(n899), .Z(n901) );
  NAND U1241 ( .A(n902), .B(n901), .Z(n960) );
  NANDN U1242 ( .A(n904), .B(n903), .Z(n908) );
  NANDN U1243 ( .A(n906), .B(n905), .Z(n907) );
  NAND U1244 ( .A(n908), .B(n907), .Z(n1027) );
  NANDN U1245 ( .A(n315), .B(a[16]), .Z(n913) );
  XNOR U1246 ( .A(b[1]), .B(n913), .Z(n915) );
  NANDN U1247 ( .A(b[0]), .B(a[15]), .Z(n914) );
  AND U1248 ( .A(n915), .B(n914), .Z(n999) );
  XOR U1249 ( .A(b[15]), .B(b[16]), .Z(n9107) );
  AND U1250 ( .A(n9107), .B(a[0]), .Z(n1011) );
  XOR U1251 ( .A(b[13]), .B(a[4]), .Z(n985) );
  NAND U1252 ( .A(n985), .B(n8730), .Z(n918) );
  NANDN U1253 ( .A(n916), .B(n8731), .Z(n917) );
  NAND U1254 ( .A(n918), .B(n917), .Z(n998) );
  XNOR U1255 ( .A(n1011), .B(n998), .Z(n1000) );
  XNOR U1256 ( .A(n999), .B(n1000), .Z(n969) );
  XOR U1257 ( .A(n969), .B(n970), .Z(n971) );
  XOR U1258 ( .A(n972), .B(n971), .Z(n963) );
  XNOR U1259 ( .A(n963), .B(n964), .Z(n965) );
  NANDN U1260 ( .A(n928), .B(n927), .Z(n978) );
  NAND U1261 ( .A(n929), .B(n7622), .Z(n931) );
  XNOR U1262 ( .A(n316), .B(a[14]), .Z(n1018) );
  NAND U1263 ( .A(n1018), .B(n7620), .Z(n930) );
  NAND U1264 ( .A(n931), .B(n930), .Z(n976) );
  XNOR U1265 ( .A(b[9]), .B(a[8]), .Z(n1012) );
  NANDN U1266 ( .A(n1012), .B(n8288), .Z(n934) );
  NAND U1267 ( .A(n932), .B(n8286), .Z(n933) );
  AND U1268 ( .A(n934), .B(n933), .Z(n975) );
  XNOR U1269 ( .A(n976), .B(n975), .Z(n977) );
  XNOR U1270 ( .A(n978), .B(n977), .Z(n994) );
  XOR U1271 ( .A(b[7]), .B(a[10]), .Z(n979) );
  NANDN U1272 ( .A(n8013), .B(n979), .Z(n937) );
  NAND U1273 ( .A(n935), .B(n8014), .Z(n936) );
  NAND U1274 ( .A(n937), .B(n936), .Z(n993) );
  XOR U1275 ( .A(b[11]), .B(a[6]), .Z(n982) );
  NAND U1276 ( .A(n8541), .B(n982), .Z(n940) );
  NAND U1277 ( .A(n8542), .B(n938), .Z(n939) );
  AND U1278 ( .A(n940), .B(n939), .Z(n991) );
  XOR U1279 ( .A(n317), .B(a[12]), .Z(n1015) );
  NANDN U1280 ( .A(n1015), .B(n7905), .Z(n943) );
  NAND U1281 ( .A(n7906), .B(n941), .Z(n942) );
  NAND U1282 ( .A(n943), .B(n942), .Z(n988) );
  XNOR U1283 ( .A(b[15]), .B(a[2]), .Z(n1008) );
  NANDN U1284 ( .A(n1008), .B(n8963), .Z(n946) );
  NAND U1285 ( .A(n944), .B(n8961), .Z(n945) );
  AND U1286 ( .A(n946), .B(n945), .Z(n989) );
  XNOR U1287 ( .A(n988), .B(n989), .Z(n990) );
  XNOR U1288 ( .A(n991), .B(n990), .Z(n992) );
  XNOR U1289 ( .A(n993), .B(n992), .Z(n995) );
  XOR U1290 ( .A(n994), .B(n995), .Z(n966) );
  XOR U1291 ( .A(n965), .B(n966), .Z(n1024) );
  XNOR U1292 ( .A(n1024), .B(n1025), .Z(n1026) );
  XNOR U1293 ( .A(n1027), .B(n1026), .Z(n958) );
  NANDN U1294 ( .A(n952), .B(n951), .Z(n956) );
  NAND U1295 ( .A(n954), .B(n953), .Z(n955) );
  AND U1296 ( .A(n956), .B(n955), .Z(n957) );
  XNOR U1297 ( .A(n958), .B(n957), .Z(n959) );
  XOR U1298 ( .A(n960), .B(n959), .Z(n1031) );
  XOR U1299 ( .A(n1032), .B(n1031), .Z(c[48]) );
  NANDN U1300 ( .A(n958), .B(n957), .Z(n962) );
  NAND U1301 ( .A(n960), .B(n959), .Z(n961) );
  NAND U1302 ( .A(n962), .B(n961), .Z(n1043) );
  NANDN U1303 ( .A(n964), .B(n963), .Z(n968) );
  NANDN U1304 ( .A(n966), .B(n965), .Z(n967) );
  NAND U1305 ( .A(n968), .B(n967), .Z(n1046) );
  OR U1306 ( .A(n970), .B(n969), .Z(n974) );
  NANDN U1307 ( .A(n972), .B(n971), .Z(n973) );
  NAND U1308 ( .A(n974), .B(n973), .Z(n1047) );
  XNOR U1309 ( .A(n1046), .B(n1047), .Z(n1048) );
  XOR U1310 ( .A(b[7]), .B(a[11]), .Z(n1092) );
  NANDN U1311 ( .A(n8013), .B(n1092), .Z(n981) );
  NAND U1312 ( .A(n979), .B(n8014), .Z(n980) );
  NAND U1313 ( .A(n981), .B(n980), .Z(n1098) );
  XOR U1314 ( .A(b[11]), .B(a[7]), .Z(n1077) );
  NAND U1315 ( .A(n1077), .B(n8541), .Z(n984) );
  NAND U1316 ( .A(n982), .B(n8542), .Z(n983) );
  NAND U1317 ( .A(n984), .B(n983), .Z(n1095) );
  XNOR U1318 ( .A(b[13]), .B(a[5]), .Z(n1083) );
  NANDN U1319 ( .A(n1083), .B(n8730), .Z(n987) );
  NAND U1320 ( .A(n985), .B(n8731), .Z(n986) );
  AND U1321 ( .A(n987), .B(n986), .Z(n1096) );
  XNOR U1322 ( .A(n1095), .B(n1096), .Z(n1097) );
  XOR U1323 ( .A(n1098), .B(n1097), .Z(n1053) );
  XNOR U1324 ( .A(n1052), .B(n1053), .Z(n1054) );
  XNOR U1325 ( .A(n1054), .B(n1055), .Z(n1059) );
  NAND U1326 ( .A(n993), .B(n992), .Z(n997) );
  NANDN U1327 ( .A(n995), .B(n994), .Z(n996) );
  NAND U1328 ( .A(n997), .B(n996), .Z(n1056) );
  NAND U1329 ( .A(n998), .B(n1011), .Z(n1002) );
  NANDN U1330 ( .A(n1000), .B(n999), .Z(n1001) );
  NAND U1331 ( .A(n1002), .B(n1001), .Z(n1104) );
  IV U1332 ( .A(b[17]), .Z(n9455) );
  XNOR U1333 ( .A(n9455), .B(a[0]), .Z(n1005) );
  XNOR U1334 ( .A(n9455), .B(b[15]), .Z(n1004) );
  XNOR U1335 ( .A(n9455), .B(b[16]), .Z(n1003) );
  AND U1336 ( .A(n1004), .B(n1003), .Z(n9105) );
  NAND U1337 ( .A(n1005), .B(n9105), .Z(n1007) );
  XNOR U1338 ( .A(n9455), .B(a[1]), .Z(n1074) );
  NAND U1339 ( .A(n1074), .B(n9107), .Z(n1006) );
  AND U1340 ( .A(n1007), .B(n1006), .Z(n1072) );
  XNOR U1341 ( .A(b[15]), .B(a[3]), .Z(n1069) );
  NANDN U1342 ( .A(n1069), .B(n8963), .Z(n1010) );
  NANDN U1343 ( .A(n1008), .B(n8961), .Z(n1009) );
  AND U1344 ( .A(n1010), .B(n1009), .Z(n1073) );
  XNOR U1345 ( .A(n1072), .B(n1073), .Z(n1065) );
  NAND U1346 ( .A(b[15]), .B(b[16]), .Z(n9187) );
  ANDN U1347 ( .B(n9187), .A(n9455), .Z(n9372) );
  NANDN U1348 ( .A(n1011), .B(n9372), .Z(n1062) );
  NANDN U1349 ( .A(n1012), .B(n8286), .Z(n1014) );
  XOR U1350 ( .A(b[9]), .B(a[9]), .Z(n1086) );
  NAND U1351 ( .A(n1086), .B(n8288), .Z(n1013) );
  NAND U1352 ( .A(n1014), .B(n1013), .Z(n1063) );
  XNOR U1353 ( .A(n1062), .B(n1063), .Z(n1064) );
  XNOR U1354 ( .A(n1065), .B(n1064), .Z(n1101) );
  XOR U1355 ( .A(n317), .B(a[13]), .Z(n1089) );
  NANDN U1356 ( .A(n1089), .B(n7905), .Z(n1017) );
  NANDN U1357 ( .A(n1015), .B(n7906), .Z(n1016) );
  NAND U1358 ( .A(n1017), .B(n1016), .Z(n1107) );
  XNOR U1359 ( .A(b[3]), .B(a[15]), .Z(n1080) );
  NANDN U1360 ( .A(n1080), .B(n7620), .Z(n1020) );
  NAND U1361 ( .A(n1018), .B(n7622), .Z(n1019) );
  AND U1362 ( .A(n1020), .B(n1019), .Z(n1108) );
  XNOR U1363 ( .A(n1107), .B(n1108), .Z(n1110) );
  NANDN U1364 ( .A(n315), .B(a[17]), .Z(n1021) );
  XNOR U1365 ( .A(b[1]), .B(n1021), .Z(n1023) );
  NANDN U1366 ( .A(b[0]), .B(a[16]), .Z(n1022) );
  AND U1367 ( .A(n1023), .B(n1022), .Z(n1109) );
  XNOR U1368 ( .A(n1110), .B(n1109), .Z(n1102) );
  XNOR U1369 ( .A(n1101), .B(n1102), .Z(n1103) );
  XNOR U1370 ( .A(n1104), .B(n1103), .Z(n1057) );
  XNOR U1371 ( .A(n1056), .B(n1057), .Z(n1058) );
  XOR U1372 ( .A(n1059), .B(n1058), .Z(n1049) );
  XOR U1373 ( .A(n1048), .B(n1049), .Z(n1040) );
  NANDN U1374 ( .A(n1025), .B(n1024), .Z(n1029) );
  NAND U1375 ( .A(n1027), .B(n1026), .Z(n1028) );
  AND U1376 ( .A(n1029), .B(n1028), .Z(n1041) );
  XNOR U1377 ( .A(n1040), .B(n1041), .Z(n1042) );
  XNOR U1378 ( .A(n1043), .B(n1042), .Z(n1035) );
  XNOR U1379 ( .A(n1035), .B(sreg[49]), .Z(n1037) );
  NAND U1380 ( .A(n1030), .B(sreg[48]), .Z(n1034) );
  OR U1381 ( .A(n1032), .B(n1031), .Z(n1033) );
  AND U1382 ( .A(n1034), .B(n1033), .Z(n1036) );
  XOR U1383 ( .A(n1037), .B(n1036), .Z(c[49]) );
  NAND U1384 ( .A(n1035), .B(sreg[49]), .Z(n1039) );
  OR U1385 ( .A(n1037), .B(n1036), .Z(n1038) );
  NAND U1386 ( .A(n1039), .B(n1038), .Z(n1195) );
  XNOR U1387 ( .A(n1195), .B(sreg[50]), .Z(n1197) );
  NANDN U1388 ( .A(n1041), .B(n1040), .Z(n1045) );
  NAND U1389 ( .A(n1043), .B(n1042), .Z(n1044) );
  NAND U1390 ( .A(n1045), .B(n1044), .Z(n1114) );
  NANDN U1391 ( .A(n1047), .B(n1046), .Z(n1051) );
  NANDN U1392 ( .A(n1049), .B(n1048), .Z(n1050) );
  NAND U1393 ( .A(n1051), .B(n1050), .Z(n1112) );
  NANDN U1394 ( .A(n1057), .B(n1056), .Z(n1061) );
  NANDN U1395 ( .A(n1059), .B(n1058), .Z(n1060) );
  NAND U1396 ( .A(n1061), .B(n1060), .Z(n1118) );
  XNOR U1397 ( .A(n1117), .B(n1118), .Z(n1119) );
  NANDN U1398 ( .A(n315), .B(a[18]), .Z(n1066) );
  XNOR U1399 ( .A(b[1]), .B(n1066), .Z(n1068) );
  IV U1400 ( .A(a[17]), .Z(n5168) );
  NANDN U1401 ( .A(n5168), .B(n315), .Z(n1067) );
  AND U1402 ( .A(n1068), .B(n1067), .Z(n1156) );
  NANDN U1403 ( .A(n1069), .B(n8961), .Z(n1071) );
  XOR U1404 ( .A(b[15]), .B(a[4]), .Z(n1138) );
  NAND U1405 ( .A(n1138), .B(n8963), .Z(n1070) );
  NAND U1406 ( .A(n1071), .B(n1070), .Z(n1157) );
  XNOR U1407 ( .A(n1156), .B(n1157), .Z(n1159) );
  XOR U1408 ( .A(b[18]), .B(b[17]), .Z(n9378) );
  NANDN U1409 ( .A(n2616), .B(n9378), .Z(n1158) );
  XNOR U1410 ( .A(n1159), .B(n1158), .Z(n1185) );
  NAND U1411 ( .A(n1074), .B(n9105), .Z(n1076) );
  XNOR U1412 ( .A(n9455), .B(a[2]), .Z(n1167) );
  NAND U1413 ( .A(n1167), .B(n9107), .Z(n1075) );
  NAND U1414 ( .A(n1076), .B(n1075), .Z(n1180) );
  XNOR U1415 ( .A(b[11]), .B(a[8]), .Z(n1147) );
  NANDN U1416 ( .A(n1147), .B(n8541), .Z(n1079) );
  NAND U1417 ( .A(n8542), .B(n1077), .Z(n1078) );
  AND U1418 ( .A(n1079), .B(n1078), .Z(n1179) );
  XNOR U1419 ( .A(n1180), .B(n1179), .Z(n1181) );
  XNOR U1420 ( .A(n1182), .B(n1181), .Z(n1186) );
  XNOR U1421 ( .A(n1185), .B(n1186), .Z(n1187) );
  XNOR U1422 ( .A(n1188), .B(n1187), .Z(n1192) );
  NANDN U1423 ( .A(n1080), .B(n7622), .Z(n1082) );
  XNOR U1424 ( .A(n316), .B(a[16]), .Z(n1150) );
  NAND U1425 ( .A(n1150), .B(n7620), .Z(n1081) );
  NAND U1426 ( .A(n1082), .B(n1081), .Z(n1175) );
  XOR U1427 ( .A(b[13]), .B(a[6]), .Z(n1135) );
  NAND U1428 ( .A(n1135), .B(n8730), .Z(n1085) );
  NANDN U1429 ( .A(n1083), .B(n8731), .Z(n1084) );
  NAND U1430 ( .A(n1085), .B(n1084), .Z(n1173) );
  XOR U1431 ( .A(b[9]), .B(a[10]), .Z(n1170) );
  NAND U1432 ( .A(n1170), .B(n8288), .Z(n1088) );
  NAND U1433 ( .A(n1086), .B(n8286), .Z(n1087) );
  AND U1434 ( .A(n1088), .B(n1087), .Z(n1174) );
  XNOR U1435 ( .A(n1173), .B(n1174), .Z(n1176) );
  XOR U1436 ( .A(n1175), .B(n1176), .Z(n1132) );
  XNOR U1437 ( .A(b[5]), .B(a[14]), .Z(n1141) );
  NANDN U1438 ( .A(n1141), .B(n7905), .Z(n1091) );
  NANDN U1439 ( .A(n1089), .B(n7906), .Z(n1090) );
  NAND U1440 ( .A(n1091), .B(n1090), .Z(n1130) );
  XNOR U1441 ( .A(b[7]), .B(a[12]), .Z(n1153) );
  OR U1442 ( .A(n1153), .B(n8013), .Z(n1094) );
  NAND U1443 ( .A(n8014), .B(n1092), .Z(n1093) );
  AND U1444 ( .A(n1094), .B(n1093), .Z(n1129) );
  XNOR U1445 ( .A(n1130), .B(n1129), .Z(n1131) );
  XNOR U1446 ( .A(n1132), .B(n1131), .Z(n1190) );
  NANDN U1447 ( .A(n1096), .B(n1095), .Z(n1100) );
  NAND U1448 ( .A(n1098), .B(n1097), .Z(n1099) );
  AND U1449 ( .A(n1100), .B(n1099), .Z(n1189) );
  XOR U1450 ( .A(n1190), .B(n1189), .Z(n1191) );
  XOR U1451 ( .A(n1192), .B(n1191), .Z(n1126) );
  NANDN U1452 ( .A(n1102), .B(n1101), .Z(n1106) );
  NAND U1453 ( .A(n1104), .B(n1103), .Z(n1105) );
  NAND U1454 ( .A(n1106), .B(n1105), .Z(n1124) );
  XNOR U1455 ( .A(n1124), .B(n1123), .Z(n1125) );
  XOR U1456 ( .A(n1126), .B(n1125), .Z(n1120) );
  XNOR U1457 ( .A(n1119), .B(n1120), .Z(n1111) );
  XNOR U1458 ( .A(n1112), .B(n1111), .Z(n1113) );
  XOR U1459 ( .A(n1114), .B(n1113), .Z(n1196) );
  XOR U1460 ( .A(n1197), .B(n1196), .Z(c[50]) );
  NANDN U1461 ( .A(n1112), .B(n1111), .Z(n1116) );
  NAND U1462 ( .A(n1114), .B(n1113), .Z(n1115) );
  NAND U1463 ( .A(n1116), .B(n1115), .Z(n1208) );
  NANDN U1464 ( .A(n1118), .B(n1117), .Z(n1122) );
  NANDN U1465 ( .A(n1120), .B(n1119), .Z(n1121) );
  NAND U1466 ( .A(n1122), .B(n1121), .Z(n1206) );
  NANDN U1467 ( .A(n1124), .B(n1123), .Z(n1128) );
  NANDN U1468 ( .A(n1126), .B(n1125), .Z(n1127) );
  NAND U1469 ( .A(n1128), .B(n1127), .Z(n1213) );
  NANDN U1470 ( .A(n1130), .B(n1129), .Z(n1134) );
  NANDN U1471 ( .A(n1132), .B(n1131), .Z(n1133) );
  NAND U1472 ( .A(n1134), .B(n1133), .Z(n1218) );
  XOR U1473 ( .A(b[13]), .B(a[7]), .Z(n1271) );
  NAND U1474 ( .A(n1271), .B(n8730), .Z(n1137) );
  NAND U1475 ( .A(n1135), .B(n8731), .Z(n1136) );
  NAND U1476 ( .A(n1137), .B(n1136), .Z(n1232) );
  NAND U1477 ( .A(n1138), .B(n8961), .Z(n1140) );
  XNOR U1478 ( .A(b[15]), .B(n3389), .Z(n1268) );
  NAND U1479 ( .A(n1268), .B(n8963), .Z(n1139) );
  NAND U1480 ( .A(n1140), .B(n1139), .Z(n1229) );
  XNOR U1481 ( .A(b[5]), .B(a[15]), .Z(n1242) );
  NANDN U1482 ( .A(n1242), .B(n7905), .Z(n1143) );
  NANDN U1483 ( .A(n1141), .B(n7906), .Z(n1142) );
  AND U1484 ( .A(n1143), .B(n1142), .Z(n1230) );
  XNOR U1485 ( .A(n1229), .B(n1230), .Z(n1231) );
  XNOR U1486 ( .A(n1232), .B(n1231), .Z(n1280) );
  NANDN U1487 ( .A(n315), .B(a[19]), .Z(n1144) );
  XNOR U1488 ( .A(b[1]), .B(n1144), .Z(n1146) );
  NANDN U1489 ( .A(b[0]), .B(a[18]), .Z(n1145) );
  AND U1490 ( .A(n1146), .B(n1145), .Z(n1254) );
  XOR U1491 ( .A(b[11]), .B(a[9]), .Z(n1262) );
  NAND U1492 ( .A(n1262), .B(n8541), .Z(n1149) );
  NANDN U1493 ( .A(n1147), .B(n8542), .Z(n1148) );
  AND U1494 ( .A(n1149), .B(n1148), .Z(n1255) );
  XOR U1495 ( .A(n1254), .B(n1255), .Z(n1257) );
  XOR U1496 ( .A(b[3]), .B(n5168), .Z(n1239) );
  NANDN U1497 ( .A(n1239), .B(n7620), .Z(n1152) );
  NAND U1498 ( .A(n1150), .B(n7622), .Z(n1151) );
  AND U1499 ( .A(n1152), .B(n1151), .Z(n1256) );
  XNOR U1500 ( .A(n1257), .B(n1256), .Z(n1277) );
  XNOR U1501 ( .A(b[7]), .B(a[13]), .Z(n1245) );
  OR U1502 ( .A(n1245), .B(n8013), .Z(n1155) );
  NANDN U1503 ( .A(n1153), .B(n8014), .Z(n1154) );
  NAND U1504 ( .A(n1155), .B(n1154), .Z(n1278) );
  XNOR U1505 ( .A(n1277), .B(n1278), .Z(n1279) );
  XOR U1506 ( .A(n1280), .B(n1279), .Z(n1217) );
  XNOR U1507 ( .A(n1218), .B(n1217), .Z(n1220) );
  NAND U1508 ( .A(n1157), .B(n1156), .Z(n1161) );
  OR U1509 ( .A(n1159), .B(n1158), .Z(n1160) );
  AND U1510 ( .A(n1161), .B(n1160), .Z(n1219) );
  XNOR U1511 ( .A(n1220), .B(n1219), .Z(n1226) );
  IV U1512 ( .A(b[19]), .Z(n9562) );
  XNOR U1513 ( .A(n9562), .B(a[0]), .Z(n1164) );
  XNOR U1514 ( .A(n9562), .B(b[18]), .Z(n1163) );
  XNOR U1515 ( .A(n9562), .B(b[17]), .Z(n1162) );
  AND U1516 ( .A(n1163), .B(n1162), .Z(n9379) );
  NAND U1517 ( .A(n1164), .B(n9379), .Z(n1166) );
  XNOR U1518 ( .A(n9562), .B(a[1]), .Z(n1265) );
  NAND U1519 ( .A(n1265), .B(n9378), .Z(n1165) );
  AND U1520 ( .A(n1166), .B(n1165), .Z(n1260) );
  XOR U1521 ( .A(b[17]), .B(n3094), .Z(n1236) );
  NANDN U1522 ( .A(n1236), .B(n9107), .Z(n1169) );
  NAND U1523 ( .A(n1167), .B(n9105), .Z(n1168) );
  AND U1524 ( .A(n1169), .B(n1168), .Z(n1261) );
  XNOR U1525 ( .A(n1260), .B(n1261), .Z(n1250) );
  NAND U1526 ( .A(n1170), .B(n8286), .Z(n1172) );
  XOR U1527 ( .A(b[9]), .B(a[11]), .Z(n1274) );
  NAND U1528 ( .A(n1274), .B(n8288), .Z(n1171) );
  NAND U1529 ( .A(n1172), .B(n1171), .Z(n1248) );
  XOR U1530 ( .A(n1249), .B(n1248), .Z(n1251) );
  XNOR U1531 ( .A(n1250), .B(n1251), .Z(n1283) );
  NANDN U1532 ( .A(n1174), .B(n1173), .Z(n1178) );
  NAND U1533 ( .A(n1176), .B(n1175), .Z(n1177) );
  AND U1534 ( .A(n1178), .B(n1177), .Z(n1284) );
  XOR U1535 ( .A(n1283), .B(n1284), .Z(n1286) );
  NANDN U1536 ( .A(n1180), .B(n1179), .Z(n1184) );
  NAND U1537 ( .A(n1182), .B(n1181), .Z(n1183) );
  NAND U1538 ( .A(n1184), .B(n1183), .Z(n1285) );
  XNOR U1539 ( .A(n1286), .B(n1285), .Z(n1223) );
  XNOR U1540 ( .A(n1223), .B(n1224), .Z(n1225) );
  XOR U1541 ( .A(n1226), .B(n1225), .Z(n1211) );
  OR U1542 ( .A(n1190), .B(n1189), .Z(n1194) );
  NAND U1543 ( .A(n1192), .B(n1191), .Z(n1193) );
  AND U1544 ( .A(n1194), .B(n1193), .Z(n1212) );
  XNOR U1545 ( .A(n1211), .B(n1212), .Z(n1214) );
  XNOR U1546 ( .A(n1213), .B(n1214), .Z(n1205) );
  XOR U1547 ( .A(n1206), .B(n1205), .Z(n1207) );
  XNOR U1548 ( .A(n1208), .B(n1207), .Z(n1200) );
  XNOR U1549 ( .A(n1200), .B(sreg[51]), .Z(n1202) );
  NAND U1550 ( .A(n1195), .B(sreg[50]), .Z(n1199) );
  OR U1551 ( .A(n1197), .B(n1196), .Z(n1198) );
  AND U1552 ( .A(n1199), .B(n1198), .Z(n1201) );
  XOR U1553 ( .A(n1202), .B(n1201), .Z(c[51]) );
  NAND U1554 ( .A(n1200), .B(sreg[51]), .Z(n1204) );
  OR U1555 ( .A(n1202), .B(n1201), .Z(n1203) );
  NAND U1556 ( .A(n1204), .B(n1203), .Z(n1384) );
  XNOR U1557 ( .A(n1384), .B(sreg[52]), .Z(n1386) );
  NAND U1558 ( .A(n1206), .B(n1205), .Z(n1210) );
  NAND U1559 ( .A(n1208), .B(n1207), .Z(n1209) );
  NAND U1560 ( .A(n1210), .B(n1209), .Z(n1292) );
  NAND U1561 ( .A(n1212), .B(n1211), .Z(n1216) );
  NANDN U1562 ( .A(n1214), .B(n1213), .Z(n1215) );
  NAND U1563 ( .A(n1216), .B(n1215), .Z(n1289) );
  OR U1564 ( .A(n1218), .B(n1217), .Z(n1222) );
  OR U1565 ( .A(n1220), .B(n1219), .Z(n1221) );
  NAND U1566 ( .A(n1222), .B(n1221), .Z(n1298) );
  NANDN U1567 ( .A(n1224), .B(n1223), .Z(n1228) );
  NAND U1568 ( .A(n1226), .B(n1225), .Z(n1227) );
  NAND U1569 ( .A(n1228), .B(n1227), .Z(n1295) );
  NANDN U1570 ( .A(n315), .B(a[20]), .Z(n1233) );
  XNOR U1571 ( .A(b[1]), .B(n1233), .Z(n1235) );
  NANDN U1572 ( .A(b[0]), .B(a[19]), .Z(n1234) );
  AND U1573 ( .A(n1235), .B(n1234), .Z(n1324) );
  XNOR U1574 ( .A(b[17]), .B(a[4]), .Z(n1348) );
  NANDN U1575 ( .A(n1348), .B(n9107), .Z(n1238) );
  NANDN U1576 ( .A(n1236), .B(n9105), .Z(n1237) );
  AND U1577 ( .A(n1238), .B(n1237), .Z(n1325) );
  XOR U1578 ( .A(n1324), .B(n1325), .Z(n1327) );
  XOR U1579 ( .A(b[20]), .B(b[19]), .Z(n9493) );
  NANDN U1580 ( .A(n2616), .B(n9493), .Z(n1326) );
  XOR U1581 ( .A(n1327), .B(n1326), .Z(n1372) );
  XNOR U1582 ( .A(b[3]), .B(a[18]), .Z(n1333) );
  NANDN U1583 ( .A(n1333), .B(n7620), .Z(n1241) );
  NANDN U1584 ( .A(n1239), .B(n7622), .Z(n1240) );
  AND U1585 ( .A(n1241), .B(n1240), .Z(n1363) );
  XNOR U1586 ( .A(b[5]), .B(a[16]), .Z(n1342) );
  NANDN U1587 ( .A(n1342), .B(n7905), .Z(n1244) );
  NANDN U1588 ( .A(n1242), .B(n7906), .Z(n1243) );
  NAND U1589 ( .A(n1244), .B(n1243), .Z(n1360) );
  XOR U1590 ( .A(b[7]), .B(a[14]), .Z(n1339) );
  NANDN U1591 ( .A(n8013), .B(n1339), .Z(n1247) );
  NANDN U1592 ( .A(n1245), .B(n8014), .Z(n1246) );
  AND U1593 ( .A(n1247), .B(n1246), .Z(n1361) );
  XNOR U1594 ( .A(n1360), .B(n1361), .Z(n1362) );
  XOR U1595 ( .A(n1363), .B(n1362), .Z(n1373) );
  XNOR U1596 ( .A(n1372), .B(n1373), .Z(n1374) );
  XNOR U1597 ( .A(n1375), .B(n1374), .Z(n1379) );
  OR U1598 ( .A(n1249), .B(n1248), .Z(n1253) );
  NAND U1599 ( .A(n1251), .B(n1250), .Z(n1252) );
  AND U1600 ( .A(n1253), .B(n1252), .Z(n1378) );
  XNOR U1601 ( .A(n1379), .B(n1378), .Z(n1380) );
  NANDN U1602 ( .A(n1255), .B(n1254), .Z(n1259) );
  OR U1603 ( .A(n1257), .B(n1256), .Z(n1258) );
  NAND U1604 ( .A(n1259), .B(n1258), .Z(n1310) );
  XNOR U1605 ( .A(b[11]), .B(a[10]), .Z(n1321) );
  NANDN U1606 ( .A(n1321), .B(n8541), .Z(n1264) );
  NAND U1607 ( .A(n8542), .B(n1262), .Z(n1263) );
  NAND U1608 ( .A(n1264), .B(n1263), .Z(n1355) );
  NAND U1609 ( .A(n1265), .B(n9379), .Z(n1267) );
  XOR U1610 ( .A(b[19]), .B(n2950), .Z(n1313) );
  NANDN U1611 ( .A(n1313), .B(n9378), .Z(n1266) );
  AND U1612 ( .A(n1267), .B(n1266), .Z(n1354) );
  XNOR U1613 ( .A(n1355), .B(n1354), .Z(n1356) );
  XOR U1614 ( .A(n1357), .B(n1356), .Z(n1307) );
  NAND U1615 ( .A(n1268), .B(n8961), .Z(n1270) );
  XOR U1616 ( .A(b[15]), .B(a[6]), .Z(n1351) );
  NAND U1617 ( .A(n1351), .B(n8963), .Z(n1269) );
  NAND U1618 ( .A(n1270), .B(n1269), .Z(n1366) );
  XNOR U1619 ( .A(b[13]), .B(a[8]), .Z(n1345) );
  NANDN U1620 ( .A(n1345), .B(n8730), .Z(n1273) );
  NAND U1621 ( .A(n8731), .B(n1271), .Z(n1272) );
  AND U1622 ( .A(n1273), .B(n1272), .Z(n1367) );
  XOR U1623 ( .A(n1366), .B(n1367), .Z(n1368) );
  XOR U1624 ( .A(b[9]), .B(a[12]), .Z(n1336) );
  NAND U1625 ( .A(n1336), .B(n8288), .Z(n1276) );
  NAND U1626 ( .A(n1274), .B(n8286), .Z(n1275) );
  AND U1627 ( .A(n1276), .B(n1275), .Z(n1369) );
  XNOR U1628 ( .A(n1368), .B(n1369), .Z(n1308) );
  XNOR U1629 ( .A(n1307), .B(n1308), .Z(n1309) );
  XNOR U1630 ( .A(n1310), .B(n1309), .Z(n1381) );
  XOR U1631 ( .A(n1380), .B(n1381), .Z(n1304) );
  NANDN U1632 ( .A(n1278), .B(n1277), .Z(n1282) );
  NAND U1633 ( .A(n1280), .B(n1279), .Z(n1281) );
  NAND U1634 ( .A(n1282), .B(n1281), .Z(n1301) );
  NANDN U1635 ( .A(n1284), .B(n1283), .Z(n1288) );
  OR U1636 ( .A(n1286), .B(n1285), .Z(n1287) );
  NAND U1637 ( .A(n1288), .B(n1287), .Z(n1302) );
  XNOR U1638 ( .A(n1301), .B(n1302), .Z(n1303) );
  XNOR U1639 ( .A(n1304), .B(n1303), .Z(n1296) );
  XNOR U1640 ( .A(n1295), .B(n1296), .Z(n1297) );
  XOR U1641 ( .A(n1298), .B(n1297), .Z(n1290) );
  XNOR U1642 ( .A(n1289), .B(n1290), .Z(n1291) );
  XOR U1643 ( .A(n1292), .B(n1291), .Z(n1385) );
  XOR U1644 ( .A(n1386), .B(n1385), .Z(c[52]) );
  NANDN U1645 ( .A(n1290), .B(n1289), .Z(n1294) );
  NAND U1646 ( .A(n1292), .B(n1291), .Z(n1293) );
  NAND U1647 ( .A(n1294), .B(n1293), .Z(n1397) );
  NANDN U1648 ( .A(n1296), .B(n1295), .Z(n1300) );
  NANDN U1649 ( .A(n1298), .B(n1297), .Z(n1299) );
  NAND U1650 ( .A(n1300), .B(n1299), .Z(n1394) );
  NANDN U1651 ( .A(n1302), .B(n1301), .Z(n1306) );
  NAND U1652 ( .A(n1304), .B(n1303), .Z(n1305) );
  NAND U1653 ( .A(n1306), .B(n1305), .Z(n1484) );
  NANDN U1654 ( .A(n1308), .B(n1307), .Z(n1312) );
  NAND U1655 ( .A(n1310), .B(n1309), .Z(n1311) );
  NAND U1656 ( .A(n1312), .B(n1311), .Z(n1476) );
  NANDN U1657 ( .A(n1313), .B(n9379), .Z(n1315) );
  XOR U1658 ( .A(b[19]), .B(n3094), .Z(n1426) );
  NANDN U1659 ( .A(n1426), .B(n9378), .Z(n1314) );
  NAND U1660 ( .A(n1315), .B(n1314), .Z(n1425) );
  XNOR U1661 ( .A(b[21]), .B(a[1]), .Z(n1450) );
  ANDN U1662 ( .B(n9493), .A(n1450), .Z(n1320) );
  XNOR U1663 ( .A(n318), .B(a[0]), .Z(n1318) );
  XNOR U1664 ( .A(n318), .B(b[20]), .Z(n1317) );
  XNOR U1665 ( .A(n318), .B(b[19]), .Z(n1316) );
  AND U1666 ( .A(n1317), .B(n1316), .Z(n9495) );
  NAND U1667 ( .A(n1318), .B(n9495), .Z(n1319) );
  NANDN U1668 ( .A(n1320), .B(n1319), .Z(n1424) );
  XNOR U1669 ( .A(n1425), .B(n1424), .Z(n1415) );
  XOR U1670 ( .A(b[11]), .B(a[11]), .Z(n1456) );
  NAND U1671 ( .A(n8541), .B(n1456), .Z(n1323) );
  NANDN U1672 ( .A(n1321), .B(n8542), .Z(n1322) );
  AND U1673 ( .A(n1323), .B(n1322), .Z(n1412) );
  XNOR U1674 ( .A(n1413), .B(n1412), .Z(n1414) );
  XOR U1675 ( .A(n1415), .B(n1414), .Z(n1408) );
  NANDN U1676 ( .A(n1325), .B(n1324), .Z(n1329) );
  OR U1677 ( .A(n1327), .B(n1326), .Z(n1328) );
  NAND U1678 ( .A(n1329), .B(n1328), .Z(n1407) );
  NANDN U1679 ( .A(n315), .B(a[21]), .Z(n1330) );
  XNOR U1680 ( .A(b[1]), .B(n1330), .Z(n1332) );
  NANDN U1681 ( .A(b[0]), .B(a[20]), .Z(n1331) );
  AND U1682 ( .A(n1332), .B(n1331), .Z(n1464) );
  XNOR U1683 ( .A(b[3]), .B(a[19]), .Z(n1418) );
  NANDN U1684 ( .A(n1418), .B(n7620), .Z(n1335) );
  NANDN U1685 ( .A(n1333), .B(n7622), .Z(n1334) );
  AND U1686 ( .A(n1335), .B(n1334), .Z(n1463) );
  XOR U1687 ( .A(n1464), .B(n1463), .Z(n1466) );
  XNOR U1688 ( .A(b[9]), .B(a[13]), .Z(n1447) );
  NANDN U1689 ( .A(n1447), .B(n8288), .Z(n1338) );
  NAND U1690 ( .A(n1336), .B(n8286), .Z(n1337) );
  AND U1691 ( .A(n1338), .B(n1337), .Z(n1465) );
  XNOR U1692 ( .A(n1466), .B(n1465), .Z(n1406) );
  XOR U1693 ( .A(n1407), .B(n1406), .Z(n1409) );
  XNOR U1694 ( .A(n1408), .B(n1409), .Z(n1471) );
  XOR U1695 ( .A(b[7]), .B(a[15]), .Z(n1438) );
  NANDN U1696 ( .A(n8013), .B(n1438), .Z(n1341) );
  NAND U1697 ( .A(n1339), .B(n8014), .Z(n1340) );
  NAND U1698 ( .A(n1341), .B(n1340), .Z(n1432) );
  XOR U1699 ( .A(b[5]), .B(n5168), .Z(n1441) );
  NANDN U1700 ( .A(n1441), .B(n7905), .Z(n1344) );
  NANDN U1701 ( .A(n1342), .B(n7906), .Z(n1343) );
  AND U1702 ( .A(n1344), .B(n1343), .Z(n1433) );
  XNOR U1703 ( .A(n1432), .B(n1433), .Z(n1434) );
  XOR U1704 ( .A(b[13]), .B(a[9]), .Z(n1421) );
  NAND U1705 ( .A(n1421), .B(n8730), .Z(n1347) );
  NANDN U1706 ( .A(n1345), .B(n8731), .Z(n1346) );
  NAND U1707 ( .A(n1347), .B(n1346), .Z(n1462) );
  NANDN U1708 ( .A(n1348), .B(n9105), .Z(n1350) );
  XNOR U1709 ( .A(n9455), .B(a[5]), .Z(n1453) );
  NAND U1710 ( .A(n1453), .B(n9107), .Z(n1349) );
  NAND U1711 ( .A(n1350), .B(n1349), .Z(n1459) );
  XOR U1712 ( .A(b[15]), .B(a[7]), .Z(n1444) );
  NAND U1713 ( .A(n1444), .B(n8963), .Z(n1353) );
  NAND U1714 ( .A(n1351), .B(n8961), .Z(n1352) );
  AND U1715 ( .A(n1353), .B(n1352), .Z(n1460) );
  XNOR U1716 ( .A(n1459), .B(n1460), .Z(n1461) );
  XNOR U1717 ( .A(n1462), .B(n1461), .Z(n1435) );
  XNOR U1718 ( .A(n1434), .B(n1435), .Z(n1469) );
  NANDN U1719 ( .A(n1355), .B(n1354), .Z(n1359) );
  NANDN U1720 ( .A(n1357), .B(n1356), .Z(n1358) );
  AND U1721 ( .A(n1359), .B(n1358), .Z(n1470) );
  XNOR U1722 ( .A(n1469), .B(n1470), .Z(n1472) );
  XOR U1723 ( .A(n1471), .B(n1472), .Z(n1475) );
  XNOR U1724 ( .A(n1476), .B(n1475), .Z(n1477) );
  NANDN U1725 ( .A(n1361), .B(n1360), .Z(n1365) );
  NANDN U1726 ( .A(n1363), .B(n1362), .Z(n1364) );
  AND U1727 ( .A(n1365), .B(n1364), .Z(n1400) );
  NANDN U1728 ( .A(n1367), .B(n1366), .Z(n1371) );
  OR U1729 ( .A(n1369), .B(n1368), .Z(n1370) );
  AND U1730 ( .A(n1371), .B(n1370), .Z(n1401) );
  XNOR U1731 ( .A(n1400), .B(n1401), .Z(n1402) );
  NANDN U1732 ( .A(n1373), .B(n1372), .Z(n1377) );
  NAND U1733 ( .A(n1375), .B(n1374), .Z(n1376) );
  AND U1734 ( .A(n1377), .B(n1376), .Z(n1403) );
  XNOR U1735 ( .A(n1477), .B(n1478), .Z(n1481) );
  NANDN U1736 ( .A(n1379), .B(n1378), .Z(n1383) );
  NANDN U1737 ( .A(n1381), .B(n1380), .Z(n1382) );
  NAND U1738 ( .A(n1383), .B(n1382), .Z(n1482) );
  XNOR U1739 ( .A(n1481), .B(n1482), .Z(n1483) );
  XNOR U1740 ( .A(n1484), .B(n1483), .Z(n1395) );
  XNOR U1741 ( .A(n1394), .B(n1395), .Z(n1396) );
  XNOR U1742 ( .A(n1397), .B(n1396), .Z(n1389) );
  XNOR U1743 ( .A(n1389), .B(sreg[53]), .Z(n1391) );
  NAND U1744 ( .A(n1384), .B(sreg[52]), .Z(n1388) );
  OR U1745 ( .A(n1386), .B(n1385), .Z(n1387) );
  AND U1746 ( .A(n1388), .B(n1387), .Z(n1390) );
  XOR U1747 ( .A(n1391), .B(n1390), .Z(c[53]) );
  NAND U1748 ( .A(n1389), .B(sreg[53]), .Z(n1393) );
  OR U1749 ( .A(n1391), .B(n1390), .Z(n1392) );
  NAND U1750 ( .A(n1393), .B(n1392), .Z(n1585) );
  XNOR U1751 ( .A(n1585), .B(sreg[54]), .Z(n1587) );
  NANDN U1752 ( .A(n1395), .B(n1394), .Z(n1399) );
  NAND U1753 ( .A(n1397), .B(n1396), .Z(n1398) );
  NAND U1754 ( .A(n1399), .B(n1398), .Z(n1490) );
  OR U1755 ( .A(n1401), .B(n1400), .Z(n1405) );
  OR U1756 ( .A(n1403), .B(n1402), .Z(n1404) );
  NAND U1757 ( .A(n1405), .B(n1404), .Z(n1496) );
  NANDN U1758 ( .A(n1407), .B(n1406), .Z(n1411) );
  NANDN U1759 ( .A(n1409), .B(n1408), .Z(n1410) );
  NAND U1760 ( .A(n1411), .B(n1410), .Z(n1500) );
  NANDN U1761 ( .A(n1413), .B(n1412), .Z(n1417) );
  NAND U1762 ( .A(n1415), .B(n1414), .Z(n1416) );
  NAND U1763 ( .A(n1417), .B(n1416), .Z(n1576) );
  NANDN U1764 ( .A(n1418), .B(n7622), .Z(n1420) );
  XNOR U1765 ( .A(n316), .B(a[20]), .Z(n1525) );
  NAND U1766 ( .A(n1525), .B(n7620), .Z(n1419) );
  NAND U1767 ( .A(n1420), .B(n1419), .Z(n1528) );
  XOR U1768 ( .A(b[13]), .B(a[10]), .Z(n1519) );
  NAND U1769 ( .A(n1519), .B(n8730), .Z(n1423) );
  NAND U1770 ( .A(n1421), .B(n8731), .Z(n1422) );
  AND U1771 ( .A(n1423), .B(n1422), .Z(n1529) );
  XOR U1772 ( .A(n1528), .B(n1529), .Z(n1531) );
  NAND U1773 ( .A(n1425), .B(n1424), .Z(n1530) );
  XNOR U1774 ( .A(n1531), .B(n1530), .Z(n1573) );
  XNOR U1775 ( .A(b[22]), .B(b[21]), .Z(n9621) );
  NANDN U1776 ( .A(n9621), .B(a[0]), .Z(n1510) );
  NANDN U1777 ( .A(n1426), .B(n9379), .Z(n1428) );
  XNOR U1778 ( .A(n9562), .B(a[4]), .Z(n1516) );
  NAND U1779 ( .A(n1516), .B(n9378), .Z(n1427) );
  NAND U1780 ( .A(n1428), .B(n1427), .Z(n1508) );
  NANDN U1781 ( .A(n315), .B(a[22]), .Z(n1429) );
  XNOR U1782 ( .A(b[1]), .B(n1429), .Z(n1431) );
  NANDN U1783 ( .A(b[0]), .B(a[21]), .Z(n1430) );
  AND U1784 ( .A(n1431), .B(n1430), .Z(n1507) );
  XOR U1785 ( .A(n1508), .B(n1507), .Z(n1509) );
  XNOR U1786 ( .A(n1510), .B(n1509), .Z(n1574) );
  XNOR U1787 ( .A(n1573), .B(n1574), .Z(n1575) );
  XNOR U1788 ( .A(n1576), .B(n1575), .Z(n1569) );
  NANDN U1789 ( .A(n1433), .B(n1432), .Z(n1437) );
  NANDN U1790 ( .A(n1435), .B(n1434), .Z(n1436) );
  AND U1791 ( .A(n1437), .B(n1436), .Z(n1570) );
  XNOR U1792 ( .A(n1569), .B(n1570), .Z(n1571) );
  XOR U1793 ( .A(b[7]), .B(a[16]), .Z(n1548) );
  NANDN U1794 ( .A(n8013), .B(n1548), .Z(n1440) );
  NAND U1795 ( .A(n1438), .B(n8014), .Z(n1439) );
  NAND U1796 ( .A(n1440), .B(n1439), .Z(n1560) );
  XNOR U1797 ( .A(b[5]), .B(a[18]), .Z(n1554) );
  NANDN U1798 ( .A(n1554), .B(n7905), .Z(n1443) );
  NANDN U1799 ( .A(n1441), .B(n7906), .Z(n1442) );
  NAND U1800 ( .A(n1443), .B(n1442), .Z(n1557) );
  XNOR U1801 ( .A(b[15]), .B(a[8]), .Z(n1522) );
  NANDN U1802 ( .A(n1522), .B(n8963), .Z(n1446) );
  NAND U1803 ( .A(n1444), .B(n8961), .Z(n1445) );
  AND U1804 ( .A(n1446), .B(n1445), .Z(n1558) );
  XNOR U1805 ( .A(n1557), .B(n1558), .Z(n1559) );
  XOR U1806 ( .A(n1560), .B(n1559), .Z(n1504) );
  XOR U1807 ( .A(b[9]), .B(a[14]), .Z(n1551) );
  NAND U1808 ( .A(n1551), .B(n8288), .Z(n1449) );
  NANDN U1809 ( .A(n1447), .B(n8286), .Z(n1448) );
  AND U1810 ( .A(n1449), .B(n1448), .Z(n1566) );
  XOR U1811 ( .A(b[21]), .B(n2950), .Z(n1540) );
  NANDN U1812 ( .A(n1540), .B(n9493), .Z(n1452) );
  NANDN U1813 ( .A(n1450), .B(n9495), .Z(n1451) );
  NAND U1814 ( .A(n1452), .B(n1451), .Z(n1563) );
  XNOR U1815 ( .A(b[17]), .B(a[6]), .Z(n1513) );
  NANDN U1816 ( .A(n1513), .B(n9107), .Z(n1455) );
  NAND U1817 ( .A(n1453), .B(n9105), .Z(n1454) );
  AND U1818 ( .A(n1455), .B(n1454), .Z(n1564) );
  XNOR U1819 ( .A(n1563), .B(n1564), .Z(n1565) );
  XOR U1820 ( .A(n1566), .B(n1565), .Z(n1501) );
  XOR U1821 ( .A(b[11]), .B(a[12]), .Z(n1534) );
  NAND U1822 ( .A(n1534), .B(n8541), .Z(n1458) );
  NAND U1823 ( .A(n1456), .B(n8542), .Z(n1457) );
  NAND U1824 ( .A(n1458), .B(n1457), .Z(n1502) );
  XOR U1825 ( .A(n1501), .B(n1502), .Z(n1503) );
  XOR U1826 ( .A(n1504), .B(n1503), .Z(n1582) );
  NANDN U1827 ( .A(n1464), .B(n1463), .Z(n1468) );
  NANDN U1828 ( .A(n1466), .B(n1465), .Z(n1467) );
  NAND U1829 ( .A(n1468), .B(n1467), .Z(n1580) );
  XNOR U1830 ( .A(n1579), .B(n1580), .Z(n1581) );
  XOR U1831 ( .A(n1582), .B(n1581), .Z(n1572) );
  XOR U1832 ( .A(n1571), .B(n1572), .Z(n1497) );
  NAND U1833 ( .A(n1470), .B(n1469), .Z(n1474) );
  OR U1834 ( .A(n1472), .B(n1471), .Z(n1473) );
  NAND U1835 ( .A(n1474), .B(n1473), .Z(n1498) );
  XNOR U1836 ( .A(n1497), .B(n1498), .Z(n1499) );
  XNOR U1837 ( .A(n1500), .B(n1499), .Z(n1493) );
  NAND U1838 ( .A(n1476), .B(n1475), .Z(n1480) );
  OR U1839 ( .A(n1478), .B(n1477), .Z(n1479) );
  AND U1840 ( .A(n1480), .B(n1479), .Z(n1494) );
  XNOR U1841 ( .A(n1493), .B(n1494), .Z(n1495) );
  XNOR U1842 ( .A(n1496), .B(n1495), .Z(n1487) );
  NANDN U1843 ( .A(n1482), .B(n1481), .Z(n1486) );
  NAND U1844 ( .A(n1484), .B(n1483), .Z(n1485) );
  AND U1845 ( .A(n1486), .B(n1485), .Z(n1488) );
  XNOR U1846 ( .A(n1487), .B(n1488), .Z(n1489) );
  XOR U1847 ( .A(n1490), .B(n1489), .Z(n1586) );
  XOR U1848 ( .A(n1587), .B(n1586), .Z(c[54]) );
  NANDN U1849 ( .A(n1488), .B(n1487), .Z(n1492) );
  NAND U1850 ( .A(n1490), .B(n1489), .Z(n1491) );
  NAND U1851 ( .A(n1492), .B(n1491), .Z(n1598) );
  NANDN U1852 ( .A(n1502), .B(n1501), .Z(n1506) );
  OR U1853 ( .A(n1504), .B(n1503), .Z(n1505) );
  NAND U1854 ( .A(n1506), .B(n1505), .Z(n1688) );
  OR U1855 ( .A(n1508), .B(n1507), .Z(n1512) );
  NAND U1856 ( .A(n1510), .B(n1509), .Z(n1511) );
  NAND U1857 ( .A(n1512), .B(n1511), .Z(n1675) );
  NANDN U1858 ( .A(n1513), .B(n9105), .Z(n1515) );
  XNOR U1859 ( .A(n9455), .B(a[7]), .Z(n1636) );
  NAND U1860 ( .A(n1636), .B(n9107), .Z(n1514) );
  NAND U1861 ( .A(n1515), .B(n1514), .Z(n1653) );
  NAND U1862 ( .A(n1516), .B(n9379), .Z(n1518) );
  XNOR U1863 ( .A(n9562), .B(a[5]), .Z(n1624) );
  NAND U1864 ( .A(n1624), .B(n9378), .Z(n1517) );
  NAND U1865 ( .A(n1518), .B(n1517), .Z(n1651) );
  XOR U1866 ( .A(b[13]), .B(a[11]), .Z(n1663) );
  NAND U1867 ( .A(n1663), .B(n8730), .Z(n1521) );
  NAND U1868 ( .A(n1519), .B(n8731), .Z(n1520) );
  AND U1869 ( .A(n1521), .B(n1520), .Z(n1652) );
  XOR U1870 ( .A(n1651), .B(n1652), .Z(n1654) );
  XNOR U1871 ( .A(n1653), .B(n1654), .Z(n1676) );
  XNOR U1872 ( .A(n1675), .B(n1676), .Z(n1677) );
  NANDN U1873 ( .A(n1522), .B(n8961), .Z(n1524) );
  XOR U1874 ( .A(b[15]), .B(a[9]), .Z(n1618) );
  NAND U1875 ( .A(n1618), .B(n8963), .Z(n1523) );
  NAND U1876 ( .A(n1524), .B(n1523), .Z(n1642) );
  IV U1877 ( .A(b[22]), .Z(n9669) );
  NAND U1878 ( .A(n1525), .B(n7622), .Z(n1527) );
  XNOR U1879 ( .A(n316), .B(a[21]), .Z(n1666) );
  NAND U1880 ( .A(n1666), .B(n7620), .Z(n1526) );
  NAND U1881 ( .A(n1527), .B(n1526), .Z(n1639) );
  XOR U1882 ( .A(n1640), .B(n1639), .Z(n1641) );
  XNOR U1883 ( .A(n1642), .B(n1641), .Z(n1678) );
  XOR U1884 ( .A(n1677), .B(n1678), .Z(n1687) );
  XNOR U1885 ( .A(n1688), .B(n1687), .Z(n1690) );
  NANDN U1886 ( .A(n1529), .B(n1528), .Z(n1533) );
  OR U1887 ( .A(n1531), .B(n1530), .Z(n1532) );
  AND U1888 ( .A(n1533), .B(n1532), .Z(n1606) );
  XNOR U1889 ( .A(b[11]), .B(a[13]), .Z(n1615) );
  NANDN U1890 ( .A(n1615), .B(n8541), .Z(n1536) );
  NAND U1891 ( .A(n1534), .B(n8542), .Z(n1535) );
  AND U1892 ( .A(n1536), .B(n1535), .Z(n1658) );
  NANDN U1893 ( .A(n315), .B(a[23]), .Z(n1537) );
  XNOR U1894 ( .A(b[1]), .B(n1537), .Z(n1539) );
  NANDN U1895 ( .A(b[0]), .B(a[22]), .Z(n1538) );
  AND U1896 ( .A(n1539), .B(n1538), .Z(n1657) );
  XNOR U1897 ( .A(n1658), .B(n1657), .Z(n1659) );
  XOR U1898 ( .A(b[21]), .B(n3094), .Z(n1612) );
  NANDN U1899 ( .A(n1612), .B(n9493), .Z(n1542) );
  NANDN U1900 ( .A(n1540), .B(n9495), .Z(n1541) );
  NAND U1901 ( .A(n1542), .B(n1541), .Z(n1661) );
  XNOR U1902 ( .A(n319), .B(a[0]), .Z(n1545) );
  XNOR U1903 ( .A(n319), .B(b[22]), .Z(n1544) );
  XNOR U1904 ( .A(n319), .B(b[21]), .Z(n1543) );
  AND U1905 ( .A(n1544), .B(n1543), .Z(n9622) );
  NAND U1906 ( .A(n1545), .B(n9622), .Z(n1547) );
  XNOR U1907 ( .A(n319), .B(a[1]), .Z(n1627) );
  ANDN U1908 ( .B(n1627), .A(n9621), .Z(n1546) );
  ANDN U1909 ( .B(n1547), .A(n1546), .Z(n1662) );
  XNOR U1910 ( .A(n1661), .B(n1662), .Z(n1660) );
  XOR U1911 ( .A(n1659), .B(n1660), .Z(n1603) );
  XNOR U1912 ( .A(b[7]), .B(a[17]), .Z(n1630) );
  OR U1913 ( .A(n1630), .B(n8013), .Z(n1550) );
  NAND U1914 ( .A(n1548), .B(n8014), .Z(n1549) );
  NAND U1915 ( .A(n1550), .B(n1549), .Z(n1648) );
  NAND U1916 ( .A(n1551), .B(n8286), .Z(n1553) );
  XOR U1917 ( .A(b[9]), .B(a[15]), .Z(n1621) );
  NAND U1918 ( .A(n1621), .B(n8288), .Z(n1552) );
  NAND U1919 ( .A(n1553), .B(n1552), .Z(n1645) );
  XNOR U1920 ( .A(b[5]), .B(a[19]), .Z(n1633) );
  NANDN U1921 ( .A(n1633), .B(n7905), .Z(n1556) );
  NANDN U1922 ( .A(n1554), .B(n7906), .Z(n1555) );
  AND U1923 ( .A(n1556), .B(n1555), .Z(n1646) );
  XNOR U1924 ( .A(n1645), .B(n1646), .Z(n1647) );
  XNOR U1925 ( .A(n1648), .B(n1647), .Z(n1604) );
  XNOR U1926 ( .A(n1603), .B(n1604), .Z(n1605) );
  XOR U1927 ( .A(n1606), .B(n1605), .Z(n1672) );
  NANDN U1928 ( .A(n1558), .B(n1557), .Z(n1562) );
  NAND U1929 ( .A(n1560), .B(n1559), .Z(n1561) );
  NAND U1930 ( .A(n1562), .B(n1561), .Z(n1670) );
  NANDN U1931 ( .A(n1564), .B(n1563), .Z(n1568) );
  NANDN U1932 ( .A(n1566), .B(n1565), .Z(n1567) );
  AND U1933 ( .A(n1568), .B(n1567), .Z(n1669) );
  XNOR U1934 ( .A(n1670), .B(n1669), .Z(n1671) );
  XOR U1935 ( .A(n1672), .B(n1671), .Z(n1689) );
  XNOR U1936 ( .A(n1690), .B(n1689), .Z(n1599) );
  NANDN U1937 ( .A(n1574), .B(n1573), .Z(n1578) );
  NAND U1938 ( .A(n1576), .B(n1575), .Z(n1577) );
  NAND U1939 ( .A(n1578), .B(n1577), .Z(n1681) );
  NANDN U1940 ( .A(n1580), .B(n1579), .Z(n1584) );
  NANDN U1941 ( .A(n1582), .B(n1581), .Z(n1583) );
  NAND U1942 ( .A(n1584), .B(n1583), .Z(n1682) );
  XNOR U1943 ( .A(n1681), .B(n1682), .Z(n1683) );
  XOR U1944 ( .A(n1684), .B(n1683), .Z(n1600) );
  XNOR U1945 ( .A(n1599), .B(n1600), .Z(n1601) );
  XOR U1946 ( .A(n1602), .B(n1601), .Z(n1595) );
  XNOR U1947 ( .A(n1596), .B(n1595), .Z(n1597) );
  XNOR U1948 ( .A(n1598), .B(n1597), .Z(n1590) );
  XNOR U1949 ( .A(n1590), .B(sreg[55]), .Z(n1592) );
  NAND U1950 ( .A(n1585), .B(sreg[54]), .Z(n1589) );
  OR U1951 ( .A(n1587), .B(n1586), .Z(n1588) );
  AND U1952 ( .A(n1589), .B(n1588), .Z(n1591) );
  XOR U1953 ( .A(n1592), .B(n1591), .Z(c[55]) );
  NAND U1954 ( .A(n1590), .B(sreg[55]), .Z(n1594) );
  OR U1955 ( .A(n1592), .B(n1591), .Z(n1593) );
  NAND U1956 ( .A(n1594), .B(n1593), .Z(n1806) );
  XNOR U1957 ( .A(n1806), .B(sreg[56]), .Z(n1808) );
  NANDN U1958 ( .A(n1604), .B(n1603), .Z(n1608) );
  NANDN U1959 ( .A(n1606), .B(n1605), .Z(n1607) );
  NAND U1960 ( .A(n1608), .B(n1607), .Z(n1708) );
  NANDN U1961 ( .A(n315), .B(a[24]), .Z(n1609) );
  XNOR U1962 ( .A(b[1]), .B(n1609), .Z(n1611) );
  IV U1963 ( .A(a[23]), .Z(n6044) );
  NANDN U1964 ( .A(n6044), .B(n315), .Z(n1610) );
  AND U1965 ( .A(n1611), .B(n1610), .Z(n1719) );
  XNOR U1966 ( .A(b[21]), .B(a[4]), .Z(n1767) );
  NANDN U1967 ( .A(n1767), .B(n9493), .Z(n1614) );
  NANDN U1968 ( .A(n1612), .B(n9495), .Z(n1613) );
  NAND U1969 ( .A(n1614), .B(n1613), .Z(n1717) );
  XOR U1970 ( .A(b[24]), .B(b[23]), .Z(n9706) );
  NANDN U1971 ( .A(n2616), .B(n9706), .Z(n1718) );
  XNOR U1972 ( .A(n1717), .B(n1718), .Z(n1720) );
  XOR U1973 ( .A(n1719), .B(n1720), .Z(n1757) );
  XOR U1974 ( .A(b[11]), .B(a[14]), .Z(n1785) );
  NAND U1975 ( .A(n1785), .B(n8541), .Z(n1617) );
  NANDN U1976 ( .A(n1615), .B(n8542), .Z(n1616) );
  NAND U1977 ( .A(n1617), .B(n1616), .Z(n1761) );
  XOR U1978 ( .A(b[15]), .B(a[10]), .Z(n1726) );
  NAND U1979 ( .A(n1726), .B(n8963), .Z(n1620) );
  NAND U1980 ( .A(n1618), .B(n8961), .Z(n1619) );
  AND U1981 ( .A(n1620), .B(n1619), .Z(n1762) );
  XNOR U1982 ( .A(n1761), .B(n1762), .Z(n1763) );
  XOR U1983 ( .A(b[9]), .B(a[16]), .Z(n1770) );
  NAND U1984 ( .A(n1770), .B(n8288), .Z(n1623) );
  NAND U1985 ( .A(n1621), .B(n8286), .Z(n1622) );
  AND U1986 ( .A(n1623), .B(n1622), .Z(n1752) );
  NAND U1987 ( .A(n1624), .B(n9379), .Z(n1626) );
  XNOR U1988 ( .A(b[19]), .B(a[6]), .Z(n1773) );
  NANDN U1989 ( .A(n1773), .B(n9378), .Z(n1625) );
  AND U1990 ( .A(n1626), .B(n1625), .Z(n1750) );
  NAND U1991 ( .A(n1627), .B(n9622), .Z(n1629) );
  XOR U1992 ( .A(b[23]), .B(n2950), .Z(n1735) );
  OR U1993 ( .A(n1735), .B(n9621), .Z(n1628) );
  AND U1994 ( .A(n1629), .B(n1628), .Z(n1749) );
  XNOR U1995 ( .A(n1750), .B(n1749), .Z(n1751) );
  XNOR U1996 ( .A(n1752), .B(n1751), .Z(n1764) );
  XNOR U1997 ( .A(n1763), .B(n1764), .Z(n1755) );
  XOR U1998 ( .A(b[7]), .B(a[18]), .Z(n1776) );
  NANDN U1999 ( .A(n8013), .B(n1776), .Z(n1632) );
  NANDN U2000 ( .A(n1630), .B(n8014), .Z(n1631) );
  NAND U2001 ( .A(n1632), .B(n1631), .Z(n1791) );
  XNOR U2002 ( .A(b[5]), .B(a[20]), .Z(n1779) );
  NANDN U2003 ( .A(n1779), .B(n7905), .Z(n1635) );
  NANDN U2004 ( .A(n1633), .B(n7906), .Z(n1634) );
  NAND U2005 ( .A(n1635), .B(n1634), .Z(n1788) );
  XOR U2006 ( .A(b[17]), .B(n3831), .Z(n1782) );
  NANDN U2007 ( .A(n1782), .B(n9107), .Z(n1638) );
  NAND U2008 ( .A(n1636), .B(n9105), .Z(n1637) );
  AND U2009 ( .A(n1638), .B(n1637), .Z(n1789) );
  XNOR U2010 ( .A(n1788), .B(n1789), .Z(n1790) );
  XOR U2011 ( .A(n1791), .B(n1790), .Z(n1756) );
  XNOR U2012 ( .A(n1755), .B(n1756), .Z(n1758) );
  XNOR U2013 ( .A(n1757), .B(n1758), .Z(n1797) );
  OR U2014 ( .A(n1640), .B(n1639), .Z(n1644) );
  NANDN U2015 ( .A(n1642), .B(n1641), .Z(n1643) );
  NAND U2016 ( .A(n1644), .B(n1643), .Z(n1794) );
  NANDN U2017 ( .A(n1646), .B(n1645), .Z(n1650) );
  NAND U2018 ( .A(n1648), .B(n1647), .Z(n1649) );
  NAND U2019 ( .A(n1650), .B(n1649), .Z(n1795) );
  XNOR U2020 ( .A(n1794), .B(n1795), .Z(n1796) );
  XOR U2021 ( .A(n1797), .B(n1796), .Z(n1714) );
  NANDN U2022 ( .A(n1652), .B(n1651), .Z(n1656) );
  NANDN U2023 ( .A(n1654), .B(n1653), .Z(n1655) );
  NAND U2024 ( .A(n1656), .B(n1655), .Z(n1801) );
  XNOR U2025 ( .A(n1801), .B(n1800), .Z(n1802) );
  NANDN U2026 ( .A(n1662), .B(n1661), .Z(n1746) );
  XOR U2027 ( .A(b[13]), .B(a[12]), .Z(n1732) );
  NAND U2028 ( .A(n8730), .B(n1732), .Z(n1665) );
  NAND U2029 ( .A(n8731), .B(n1663), .Z(n1664) );
  NAND U2030 ( .A(n1665), .B(n1664), .Z(n1744) );
  XNOR U2031 ( .A(b[3]), .B(a[22]), .Z(n1723) );
  NANDN U2032 ( .A(n1723), .B(n7620), .Z(n1668) );
  NAND U2033 ( .A(n1666), .B(n7622), .Z(n1667) );
  AND U2034 ( .A(n1668), .B(n1667), .Z(n1743) );
  XNOR U2035 ( .A(n1744), .B(n1743), .Z(n1745) );
  XNOR U2036 ( .A(n1746), .B(n1745), .Z(n1803) );
  XOR U2037 ( .A(n1802), .B(n1803), .Z(n1711) );
  NANDN U2038 ( .A(n1670), .B(n1669), .Z(n1674) );
  NAND U2039 ( .A(n1672), .B(n1671), .Z(n1673) );
  NAND U2040 ( .A(n1674), .B(n1673), .Z(n1712) );
  XNOR U2041 ( .A(n1711), .B(n1712), .Z(n1713) );
  XNOR U2042 ( .A(n1714), .B(n1713), .Z(n1706) );
  NANDN U2043 ( .A(n1676), .B(n1675), .Z(n1680) );
  NAND U2044 ( .A(n1678), .B(n1677), .Z(n1679) );
  AND U2045 ( .A(n1680), .B(n1679), .Z(n1705) );
  XNOR U2046 ( .A(n1706), .B(n1705), .Z(n1707) );
  XNOR U2047 ( .A(n1708), .B(n1707), .Z(n1702) );
  NANDN U2048 ( .A(n1682), .B(n1681), .Z(n1686) );
  NANDN U2049 ( .A(n1684), .B(n1683), .Z(n1685) );
  NAND U2050 ( .A(n1686), .B(n1685), .Z(n1699) );
  NAND U2051 ( .A(n1688), .B(n1687), .Z(n1692) );
  NANDN U2052 ( .A(n1690), .B(n1689), .Z(n1691) );
  AND U2053 ( .A(n1692), .B(n1691), .Z(n1700) );
  XNOR U2054 ( .A(n1699), .B(n1700), .Z(n1701) );
  XOR U2055 ( .A(n1702), .B(n1701), .Z(n1693) );
  XOR U2056 ( .A(n1694), .B(n1693), .Z(n1695) );
  XOR U2057 ( .A(n1696), .B(n1695), .Z(n1807) );
  XOR U2058 ( .A(n1808), .B(n1807), .Z(c[56]) );
  NAND U2059 ( .A(n1694), .B(n1693), .Z(n1698) );
  NAND U2060 ( .A(n1696), .B(n1695), .Z(n1697) );
  NAND U2061 ( .A(n1698), .B(n1697), .Z(n1819) );
  NANDN U2062 ( .A(n1700), .B(n1699), .Z(n1704) );
  NAND U2063 ( .A(n1702), .B(n1701), .Z(n1703) );
  NAND U2064 ( .A(n1704), .B(n1703), .Z(n1816) );
  NANDN U2065 ( .A(n1706), .B(n1705), .Z(n1710) );
  NAND U2066 ( .A(n1708), .B(n1707), .Z(n1709) );
  NAND U2067 ( .A(n1710), .B(n1709), .Z(n1825) );
  NANDN U2068 ( .A(n1712), .B(n1711), .Z(n1716) );
  NAND U2069 ( .A(n1714), .B(n1713), .Z(n1715) );
  NAND U2070 ( .A(n1716), .B(n1715), .Z(n1822) );
  NANDN U2071 ( .A(n1718), .B(n1717), .Z(n1722) );
  NAND U2072 ( .A(n1720), .B(n1719), .Z(n1721) );
  NAND U2073 ( .A(n1722), .B(n1721), .Z(n1904) );
  XOR U2074 ( .A(b[3]), .B(n6044), .Z(n1849) );
  NANDN U2075 ( .A(n1849), .B(n7620), .Z(n1725) );
  NANDN U2076 ( .A(n1723), .B(n7622), .Z(n1724) );
  AND U2077 ( .A(n1725), .B(n1724), .Z(n1882) );
  XOR U2078 ( .A(n1883), .B(n1882), .Z(n1885) );
  XOR U2079 ( .A(b[15]), .B(a[11]), .Z(n1846) );
  NAND U2080 ( .A(n1846), .B(n8963), .Z(n1728) );
  NAND U2081 ( .A(n1726), .B(n8961), .Z(n1727) );
  AND U2082 ( .A(n1728), .B(n1727), .Z(n1884) );
  XNOR U2083 ( .A(n1885), .B(n1884), .Z(n1902) );
  NANDN U2084 ( .A(n315), .B(a[25]), .Z(n1729) );
  XNOR U2085 ( .A(b[1]), .B(n1729), .Z(n1731) );
  NANDN U2086 ( .A(b[0]), .B(a[24]), .Z(n1730) );
  AND U2087 ( .A(n1731), .B(n1730), .Z(n1897) );
  XNOR U2088 ( .A(b[13]), .B(a[13]), .Z(n1858) );
  NANDN U2089 ( .A(n1858), .B(n8730), .Z(n1734) );
  NAND U2090 ( .A(n1732), .B(n8731), .Z(n1733) );
  AND U2091 ( .A(n1734), .B(n1733), .Z(n1898) );
  XNOR U2092 ( .A(n1897), .B(n1898), .Z(n1899) );
  NANDN U2093 ( .A(n1735), .B(n9622), .Z(n1737) );
  XOR U2094 ( .A(b[23]), .B(n3094), .Z(n1879) );
  OR U2095 ( .A(n1879), .B(n9621), .Z(n1736) );
  NAND U2096 ( .A(n1737), .B(n1736), .Z(n1844) );
  XNOR U2097 ( .A(n320), .B(a[0]), .Z(n1740) );
  XNOR U2098 ( .A(n320), .B(b[24]), .Z(n1739) );
  XNOR U2099 ( .A(n320), .B(b[23]), .Z(n1738) );
  AND U2100 ( .A(n1739), .B(n1738), .Z(n9707) );
  NAND U2101 ( .A(n1740), .B(n9707), .Z(n1742) );
  XNOR U2102 ( .A(b[25]), .B(a[1]), .Z(n1891) );
  ANDN U2103 ( .B(n9706), .A(n1891), .Z(n1741) );
  ANDN U2104 ( .B(n1742), .A(n1741), .Z(n1845) );
  XNOR U2105 ( .A(n1844), .B(n1845), .Z(n1900) );
  XOR U2106 ( .A(n1899), .B(n1900), .Z(n1901) );
  XNOR U2107 ( .A(n1902), .B(n1901), .Z(n1903) );
  XNOR U2108 ( .A(n1904), .B(n1903), .Z(n1908) );
  NANDN U2109 ( .A(n1744), .B(n1743), .Z(n1748) );
  NAND U2110 ( .A(n1746), .B(n1745), .Z(n1747) );
  NAND U2111 ( .A(n1748), .B(n1747), .Z(n1905) );
  OR U2112 ( .A(n1750), .B(n1749), .Z(n1754) );
  OR U2113 ( .A(n1752), .B(n1751), .Z(n1753) );
  NAND U2114 ( .A(n1754), .B(n1753), .Z(n1906) );
  XNOR U2115 ( .A(n1905), .B(n1906), .Z(n1907) );
  XOR U2116 ( .A(n1908), .B(n1907), .Z(n1831) );
  OR U2117 ( .A(n1756), .B(n1755), .Z(n1760) );
  OR U2118 ( .A(n1758), .B(n1757), .Z(n1759) );
  AND U2119 ( .A(n1760), .B(n1759), .Z(n1828) );
  NANDN U2120 ( .A(n1762), .B(n1761), .Z(n1766) );
  NANDN U2121 ( .A(n1764), .B(n1763), .Z(n1765) );
  NAND U2122 ( .A(n1766), .B(n1765), .Z(n1914) );
  XOR U2123 ( .A(b[21]), .B(n3389), .Z(n1888) );
  NANDN U2124 ( .A(n1888), .B(n9493), .Z(n1769) );
  NANDN U2125 ( .A(n1767), .B(n9495), .Z(n1768) );
  NAND U2126 ( .A(n1769), .B(n1768), .Z(n1861) );
  XNOR U2127 ( .A(b[9]), .B(a[17]), .Z(n1870) );
  NANDN U2128 ( .A(n1870), .B(n8288), .Z(n1772) );
  NAND U2129 ( .A(n1770), .B(n8286), .Z(n1771) );
  AND U2130 ( .A(n1772), .B(n1771), .Z(n1862) );
  XNOR U2131 ( .A(n1861), .B(n1862), .Z(n1863) );
  NANDN U2132 ( .A(n1773), .B(n9379), .Z(n1775) );
  XNOR U2133 ( .A(b[19]), .B(a[7]), .Z(n1855) );
  NANDN U2134 ( .A(n1855), .B(n9378), .Z(n1774) );
  AND U2135 ( .A(n1775), .B(n1774), .Z(n1864) );
  XOR U2136 ( .A(n1863), .B(n1864), .Z(n1837) );
  XOR U2137 ( .A(b[7]), .B(a[19]), .Z(n1867) );
  NANDN U2138 ( .A(n8013), .B(n1867), .Z(n1778) );
  NAND U2139 ( .A(n1776), .B(n8014), .Z(n1777) );
  NAND U2140 ( .A(n1778), .B(n1777), .Z(n1841) );
  XNOR U2141 ( .A(b[5]), .B(a[21]), .Z(n1852) );
  NANDN U2142 ( .A(n1852), .B(n7905), .Z(n1781) );
  NANDN U2143 ( .A(n1779), .B(n7906), .Z(n1780) );
  NAND U2144 ( .A(n1781), .B(n1780), .Z(n1838) );
  XNOR U2145 ( .A(b[17]), .B(a[9]), .Z(n1894) );
  NANDN U2146 ( .A(n1894), .B(n9107), .Z(n1784) );
  NANDN U2147 ( .A(n1782), .B(n9105), .Z(n1783) );
  AND U2148 ( .A(n1784), .B(n1783), .Z(n1839) );
  XNOR U2149 ( .A(n1838), .B(n1839), .Z(n1840) );
  XNOR U2150 ( .A(n1841), .B(n1840), .Z(n1834) );
  XOR U2151 ( .A(b[11]), .B(a[15]), .Z(n1873) );
  NAND U2152 ( .A(n8541), .B(n1873), .Z(n1787) );
  NAND U2153 ( .A(n8542), .B(n1785), .Z(n1786) );
  NAND U2154 ( .A(n1787), .B(n1786), .Z(n1835) );
  XNOR U2155 ( .A(n1834), .B(n1835), .Z(n1836) );
  XNOR U2156 ( .A(n1837), .B(n1836), .Z(n1911) );
  NANDN U2157 ( .A(n1789), .B(n1788), .Z(n1793) );
  NAND U2158 ( .A(n1791), .B(n1790), .Z(n1792) );
  AND U2159 ( .A(n1793), .B(n1792), .Z(n1912) );
  XNOR U2160 ( .A(n1911), .B(n1912), .Z(n1913) );
  XOR U2161 ( .A(n1914), .B(n1913), .Z(n1829) );
  XOR U2162 ( .A(n1828), .B(n1829), .Z(n1830) );
  XOR U2163 ( .A(n1831), .B(n1830), .Z(n1920) );
  NANDN U2164 ( .A(n1795), .B(n1794), .Z(n1799) );
  NANDN U2165 ( .A(n1797), .B(n1796), .Z(n1798) );
  NAND U2166 ( .A(n1799), .B(n1798), .Z(n1918) );
  NANDN U2167 ( .A(n1801), .B(n1800), .Z(n1805) );
  NANDN U2168 ( .A(n1803), .B(n1802), .Z(n1804) );
  AND U2169 ( .A(n1805), .B(n1804), .Z(n1917) );
  XNOR U2170 ( .A(n1918), .B(n1917), .Z(n1919) );
  XOR U2171 ( .A(n1920), .B(n1919), .Z(n1823) );
  XNOR U2172 ( .A(n1822), .B(n1823), .Z(n1824) );
  XOR U2173 ( .A(n1825), .B(n1824), .Z(n1817) );
  XNOR U2174 ( .A(n1816), .B(n1817), .Z(n1818) );
  XNOR U2175 ( .A(n1819), .B(n1818), .Z(n1811) );
  XNOR U2176 ( .A(n1811), .B(sreg[57]), .Z(n1813) );
  NAND U2177 ( .A(n1806), .B(sreg[56]), .Z(n1810) );
  OR U2178 ( .A(n1808), .B(n1807), .Z(n1809) );
  AND U2179 ( .A(n1810), .B(n1809), .Z(n1812) );
  XOR U2180 ( .A(n1813), .B(n1812), .Z(c[57]) );
  NAND U2181 ( .A(n1811), .B(sreg[57]), .Z(n1815) );
  OR U2182 ( .A(n1813), .B(n1812), .Z(n1814) );
  NAND U2183 ( .A(n1815), .B(n1814), .Z(n2041) );
  XNOR U2184 ( .A(n2041), .B(sreg[58]), .Z(n2043) );
  NANDN U2185 ( .A(n1817), .B(n1816), .Z(n1821) );
  NAND U2186 ( .A(n1819), .B(n1818), .Z(n1820) );
  NAND U2187 ( .A(n1821), .B(n1820), .Z(n1926) );
  NANDN U2188 ( .A(n1823), .B(n1822), .Z(n1827) );
  NAND U2189 ( .A(n1825), .B(n1824), .Z(n1826) );
  NAND U2190 ( .A(n1827), .B(n1826), .Z(n1924) );
  OR U2191 ( .A(n1829), .B(n1828), .Z(n1833) );
  NAND U2192 ( .A(n1831), .B(n1830), .Z(n1832) );
  NAND U2193 ( .A(n1833), .B(n1832), .Z(n1931) );
  NANDN U2194 ( .A(n1839), .B(n1838), .Z(n1843) );
  NAND U2195 ( .A(n1841), .B(n1840), .Z(n1842) );
  NAND U2196 ( .A(n1843), .B(n1842), .Z(n1968) );
  NANDN U2197 ( .A(n1845), .B(n1844), .Z(n2027) );
  NAND U2198 ( .A(n1846), .B(n8961), .Z(n1848) );
  XOR U2199 ( .A(b[15]), .B(a[12]), .Z(n2001) );
  NAND U2200 ( .A(n2001), .B(n8963), .Z(n1847) );
  NAND U2201 ( .A(n1848), .B(n1847), .Z(n2029) );
  XNOR U2202 ( .A(b[3]), .B(a[24]), .Z(n1998) );
  NANDN U2203 ( .A(n1998), .B(n7620), .Z(n1851) );
  NANDN U2204 ( .A(n1849), .B(n7622), .Z(n1850) );
  AND U2205 ( .A(n1851), .B(n1850), .Z(n2030) );
  XNOR U2206 ( .A(n2029), .B(n2030), .Z(n2028) );
  XNOR U2207 ( .A(n2027), .B(n2028), .Z(n1965) );
  XNOR U2208 ( .A(b[5]), .B(a[22]), .Z(n2024) );
  NANDN U2209 ( .A(n2024), .B(n7905), .Z(n1854) );
  NANDN U2210 ( .A(n1852), .B(n7906), .Z(n1853) );
  NAND U2211 ( .A(n1854), .B(n1853), .Z(n1974) );
  NANDN U2212 ( .A(n1855), .B(n9379), .Z(n1857) );
  XNOR U2213 ( .A(n9562), .B(a[8]), .Z(n2021) );
  NAND U2214 ( .A(n2021), .B(n9378), .Z(n1856) );
  NAND U2215 ( .A(n1857), .B(n1856), .Z(n1971) );
  XOR U2216 ( .A(b[13]), .B(a[14]), .Z(n2015) );
  NAND U2217 ( .A(n2015), .B(n8730), .Z(n1860) );
  NANDN U2218 ( .A(n1858), .B(n8731), .Z(n1859) );
  AND U2219 ( .A(n1860), .B(n1859), .Z(n1972) );
  XNOR U2220 ( .A(n1971), .B(n1972), .Z(n1973) );
  XNOR U2221 ( .A(n1974), .B(n1973), .Z(n1966) );
  XNOR U2222 ( .A(n1965), .B(n1966), .Z(n1967) );
  XOR U2223 ( .A(n1968), .B(n1967), .Z(n1942) );
  XOR U2224 ( .A(n1941), .B(n1942), .Z(n1944) );
  NANDN U2225 ( .A(n1862), .B(n1861), .Z(n1866) );
  NANDN U2226 ( .A(n1864), .B(n1863), .Z(n1865) );
  NAND U2227 ( .A(n1866), .B(n1865), .Z(n1961) );
  XOR U2228 ( .A(b[7]), .B(a[20]), .Z(n2018) );
  NANDN U2229 ( .A(n8013), .B(n2018), .Z(n1869) );
  NAND U2230 ( .A(n1867), .B(n8014), .Z(n1868) );
  NAND U2231 ( .A(n1869), .B(n1868), .Z(n2034) );
  NANDN U2232 ( .A(n1870), .B(n8286), .Z(n1872) );
  XOR U2233 ( .A(b[9]), .B(a[18]), .Z(n1983) );
  NAND U2234 ( .A(n1983), .B(n8288), .Z(n1871) );
  NAND U2235 ( .A(n1872), .B(n1871), .Z(n2031) );
  XOR U2236 ( .A(b[11]), .B(a[16]), .Z(n1980) );
  NAND U2237 ( .A(n1980), .B(n8541), .Z(n1875) );
  NAND U2238 ( .A(n1873), .B(n8542), .Z(n1874) );
  AND U2239 ( .A(n1875), .B(n1874), .Z(n2032) );
  XNOR U2240 ( .A(n2031), .B(n2032), .Z(n2033) );
  XNOR U2241 ( .A(n2034), .B(n2033), .Z(n1959) );
  XNOR U2242 ( .A(b[26]), .B(b[25]), .Z(n9751) );
  NANDN U2243 ( .A(n9751), .B(a[0]), .Z(n1995) );
  NANDN U2244 ( .A(n315), .B(a[26]), .Z(n1876) );
  XNOR U2245 ( .A(b[1]), .B(n1876), .Z(n1878) );
  NANDN U2246 ( .A(b[0]), .B(a[25]), .Z(n1877) );
  AND U2247 ( .A(n1878), .B(n1877), .Z(n1993) );
  XNOR U2248 ( .A(b[23]), .B(a[4]), .Z(n1989) );
  OR U2249 ( .A(n1989), .B(n9621), .Z(n1881) );
  NANDN U2250 ( .A(n1879), .B(n9622), .Z(n1880) );
  AND U2251 ( .A(n1881), .B(n1880), .Z(n1992) );
  XNOR U2252 ( .A(n1993), .B(n1992), .Z(n1994) );
  XNOR U2253 ( .A(n1995), .B(n1994), .Z(n1960) );
  XOR U2254 ( .A(n1959), .B(n1960), .Z(n1962) );
  XOR U2255 ( .A(n1961), .B(n1962), .Z(n1943) );
  XOR U2256 ( .A(n1944), .B(n1943), .Z(n1949) );
  NANDN U2257 ( .A(n1883), .B(n1882), .Z(n1887) );
  NANDN U2258 ( .A(n1885), .B(n1884), .Z(n1886) );
  NAND U2259 ( .A(n1887), .B(n1886), .Z(n1956) );
  XNOR U2260 ( .A(b[21]), .B(a[6]), .Z(n1986) );
  NANDN U2261 ( .A(n1986), .B(n9493), .Z(n1890) );
  NANDN U2262 ( .A(n1888), .B(n9495), .Z(n1889) );
  NAND U2263 ( .A(n1890), .B(n1889), .Z(n2035) );
  XOR U2264 ( .A(b[25]), .B(n2950), .Z(n2004) );
  NANDN U2265 ( .A(n2004), .B(n9706), .Z(n1893) );
  NANDN U2266 ( .A(n1891), .B(n9707), .Z(n1892) );
  AND U2267 ( .A(n1893), .B(n1892), .Z(n2036) );
  XNOR U2268 ( .A(n2035), .B(n2036), .Z(n2037) );
  XNOR U2269 ( .A(b[17]), .B(a[10]), .Z(n1977) );
  NANDN U2270 ( .A(n1977), .B(n9107), .Z(n1896) );
  NANDN U2271 ( .A(n1894), .B(n9105), .Z(n1895) );
  AND U2272 ( .A(n1896), .B(n1895), .Z(n2038) );
  XOR U2273 ( .A(n2037), .B(n2038), .Z(n1953) );
  XNOR U2274 ( .A(n1953), .B(n1954), .Z(n1955) );
  XNOR U2275 ( .A(n1956), .B(n1955), .Z(n1947) );
  XOR U2276 ( .A(n1947), .B(n1948), .Z(n1950) );
  XOR U2277 ( .A(n1949), .B(n1950), .Z(n1938) );
  NANDN U2278 ( .A(n1906), .B(n1905), .Z(n1910) );
  NAND U2279 ( .A(n1908), .B(n1907), .Z(n1909) );
  NAND U2280 ( .A(n1910), .B(n1909), .Z(n1935) );
  NANDN U2281 ( .A(n1912), .B(n1911), .Z(n1916) );
  NAND U2282 ( .A(n1914), .B(n1913), .Z(n1915) );
  NAND U2283 ( .A(n1916), .B(n1915), .Z(n1936) );
  XNOR U2284 ( .A(n1935), .B(n1936), .Z(n1937) );
  XNOR U2285 ( .A(n1938), .B(n1937), .Z(n1929) );
  NANDN U2286 ( .A(n1918), .B(n1917), .Z(n1922) );
  NANDN U2287 ( .A(n1920), .B(n1919), .Z(n1921) );
  AND U2288 ( .A(n1922), .B(n1921), .Z(n1930) );
  XNOR U2289 ( .A(n1929), .B(n1930), .Z(n1932) );
  XNOR U2290 ( .A(n1931), .B(n1932), .Z(n1923) );
  XNOR U2291 ( .A(n1924), .B(n1923), .Z(n1925) );
  XOR U2292 ( .A(n1926), .B(n1925), .Z(n2042) );
  XOR U2293 ( .A(n2043), .B(n2042), .Z(c[58]) );
  NANDN U2294 ( .A(n1924), .B(n1923), .Z(n1928) );
  NAND U2295 ( .A(n1926), .B(n1925), .Z(n1927) );
  NAND U2296 ( .A(n1928), .B(n1927), .Z(n2054) );
  NAND U2297 ( .A(n1930), .B(n1929), .Z(n1934) );
  NANDN U2298 ( .A(n1932), .B(n1931), .Z(n1933) );
  NAND U2299 ( .A(n1934), .B(n1933), .Z(n2051) );
  NANDN U2300 ( .A(n1936), .B(n1935), .Z(n1940) );
  NANDN U2301 ( .A(n1938), .B(n1937), .Z(n1939) );
  NAND U2302 ( .A(n1940), .B(n1939), .Z(n2060) );
  OR U2303 ( .A(n1942), .B(n1941), .Z(n1946) );
  NAND U2304 ( .A(n1944), .B(n1943), .Z(n1945) );
  NAND U2305 ( .A(n1946), .B(n1945), .Z(n2057) );
  NANDN U2306 ( .A(n1948), .B(n1947), .Z(n1952) );
  OR U2307 ( .A(n1950), .B(n1949), .Z(n1951) );
  NAND U2308 ( .A(n1952), .B(n1951), .Z(n2164) );
  NANDN U2309 ( .A(n1954), .B(n1953), .Z(n1958) );
  NAND U2310 ( .A(n1956), .B(n1955), .Z(n1957) );
  NAND U2311 ( .A(n1958), .B(n1957), .Z(n2148) );
  NANDN U2312 ( .A(n1960), .B(n1959), .Z(n1964) );
  OR U2313 ( .A(n1962), .B(n1961), .Z(n1963) );
  NAND U2314 ( .A(n1964), .B(n1963), .Z(n2145) );
  NANDN U2315 ( .A(n1966), .B(n1965), .Z(n1970) );
  NAND U2316 ( .A(n1968), .B(n1967), .Z(n1969) );
  NAND U2317 ( .A(n1970), .B(n1969), .Z(n2146) );
  XNOR U2318 ( .A(n2145), .B(n2146), .Z(n2147) );
  XNOR U2319 ( .A(n2148), .B(n2147), .Z(n2161) );
  NANDN U2320 ( .A(n1972), .B(n1971), .Z(n1976) );
  NAND U2321 ( .A(n1974), .B(n1973), .Z(n1975) );
  NAND U2322 ( .A(n1976), .B(n1975), .Z(n2151) );
  NANDN U2323 ( .A(n1977), .B(n9105), .Z(n1979) );
  XNOR U2324 ( .A(n9455), .B(a[11]), .Z(n2093) );
  NAND U2325 ( .A(n2093), .B(n9107), .Z(n1978) );
  NAND U2326 ( .A(n1979), .B(n1978), .Z(n2111) );
  XNOR U2327 ( .A(b[11]), .B(a[17]), .Z(n2096) );
  NANDN U2328 ( .A(n2096), .B(n8541), .Z(n1982) );
  NAND U2329 ( .A(n1980), .B(n8542), .Z(n1981) );
  AND U2330 ( .A(n1982), .B(n1981), .Z(n2112) );
  XNOR U2331 ( .A(n2111), .B(n2112), .Z(n2113) );
  XOR U2332 ( .A(b[9]), .B(a[19]), .Z(n2108) );
  NAND U2333 ( .A(n2108), .B(n8288), .Z(n1985) );
  NAND U2334 ( .A(n1983), .B(n8286), .Z(n1984) );
  AND U2335 ( .A(n1985), .B(n1984), .Z(n2072) );
  XNOR U2336 ( .A(b[21]), .B(a[7]), .Z(n2105) );
  NANDN U2337 ( .A(n2105), .B(n9493), .Z(n1988) );
  NANDN U2338 ( .A(n1986), .B(n9495), .Z(n1987) );
  NAND U2339 ( .A(n1988), .B(n1987), .Z(n2069) );
  NANDN U2340 ( .A(n1989), .B(n9622), .Z(n1991) );
  XOR U2341 ( .A(b[23]), .B(n3389), .Z(n2084) );
  OR U2342 ( .A(n2084), .B(n9621), .Z(n1990) );
  AND U2343 ( .A(n1991), .B(n1990), .Z(n2070) );
  XNOR U2344 ( .A(n2069), .B(n2070), .Z(n2071) );
  XOR U2345 ( .A(n2072), .B(n2071), .Z(n2114) );
  XOR U2346 ( .A(n2113), .B(n2114), .Z(n2143) );
  NANDN U2347 ( .A(n1993), .B(n1992), .Z(n1997) );
  NAND U2348 ( .A(n1995), .B(n1994), .Z(n1996) );
  NAND U2349 ( .A(n1997), .B(n1996), .Z(n2141) );
  IV U2350 ( .A(b[26]), .Z(n9837) );
  ANDN U2351 ( .B(b[27]), .A(n9751), .Z(n9804) );
  NANDN U2352 ( .A(n1998), .B(n7622), .Z(n2000) );
  XNOR U2353 ( .A(n316), .B(a[25]), .Z(n2087) );
  NAND U2354 ( .A(n2087), .B(n7620), .Z(n1999) );
  NAND U2355 ( .A(n2000), .B(n1999), .Z(n2135) );
  XNOR U2356 ( .A(b[15]), .B(a[13]), .Z(n2127) );
  NANDN U2357 ( .A(n2127), .B(n8963), .Z(n2003) );
  NAND U2358 ( .A(n2001), .B(n8961), .Z(n2002) );
  AND U2359 ( .A(n2003), .B(n2002), .Z(n2136) );
  XOR U2360 ( .A(n2135), .B(n2136), .Z(n2138) );
  XNOR U2361 ( .A(n2137), .B(n2138), .Z(n2142) );
  XNOR U2362 ( .A(n2141), .B(n2142), .Z(n2144) );
  XNOR U2363 ( .A(n2143), .B(n2144), .Z(n2152) );
  XOR U2364 ( .A(n2151), .B(n2152), .Z(n2153) );
  XOR U2365 ( .A(b[25]), .B(n3094), .Z(n2124) );
  NANDN U2366 ( .A(n2124), .B(n9706), .Z(n2006) );
  NANDN U2367 ( .A(n2004), .B(n9707), .Z(n2005) );
  NAND U2368 ( .A(n2006), .B(n2005), .Z(n2134) );
  XNOR U2369 ( .A(b[27]), .B(a[1]), .Z(n2130) );
  NOR U2370 ( .A(n9751), .B(n2130), .Z(n2011) );
  XNOR U2371 ( .A(n321), .B(a[0]), .Z(n2009) );
  XNOR U2372 ( .A(n321), .B(b[26]), .Z(n2008) );
  XNOR U2373 ( .A(n321), .B(b[25]), .Z(n2007) );
  AND U2374 ( .A(n2008), .B(n2007), .Z(n9801) );
  NAND U2375 ( .A(n2009), .B(n9801), .Z(n2010) );
  NANDN U2376 ( .A(n2011), .B(n2010), .Z(n2133) );
  XNOR U2377 ( .A(n2134), .B(n2133), .Z(n2078) );
  NANDN U2378 ( .A(n315), .B(a[27]), .Z(n2012) );
  XNOR U2379 ( .A(b[1]), .B(n2012), .Z(n2014) );
  IV U2380 ( .A(a[26]), .Z(n6500) );
  NANDN U2381 ( .A(n6500), .B(n315), .Z(n2013) );
  AND U2382 ( .A(n2014), .B(n2013), .Z(n2076) );
  XOR U2383 ( .A(b[13]), .B(a[15]), .Z(n2081) );
  NAND U2384 ( .A(n8730), .B(n2081), .Z(n2017) );
  NAND U2385 ( .A(n8731), .B(n2015), .Z(n2016) );
  AND U2386 ( .A(n2017), .B(n2016), .Z(n2075) );
  XNOR U2387 ( .A(n2076), .B(n2075), .Z(n2077) );
  XOR U2388 ( .A(n2078), .B(n2077), .Z(n2063) );
  XOR U2389 ( .A(b[7]), .B(a[21]), .Z(n2090) );
  NANDN U2390 ( .A(n8013), .B(n2090), .Z(n2020) );
  NAND U2391 ( .A(n2018), .B(n8014), .Z(n2019) );
  NAND U2392 ( .A(n2020), .B(n2019), .Z(n2118) );
  NAND U2393 ( .A(n2021), .B(n9379), .Z(n2023) );
  XNOR U2394 ( .A(n9562), .B(a[9]), .Z(n2102) );
  NAND U2395 ( .A(n2102), .B(n9378), .Z(n2022) );
  NAND U2396 ( .A(n2023), .B(n2022), .Z(n2115) );
  XOR U2397 ( .A(b[5]), .B(n6044), .Z(n2099) );
  NANDN U2398 ( .A(n2099), .B(n7905), .Z(n2026) );
  NANDN U2399 ( .A(n2024), .B(n7906), .Z(n2025) );
  AND U2400 ( .A(n2026), .B(n2025), .Z(n2116) );
  XNOR U2401 ( .A(n2115), .B(n2116), .Z(n2117) );
  XNOR U2402 ( .A(n2118), .B(n2117), .Z(n2064) );
  XOR U2403 ( .A(n2063), .B(n2064), .Z(n2065) );
  XOR U2404 ( .A(n2065), .B(n2066), .Z(n2160) );
  NANDN U2405 ( .A(n2036), .B(n2035), .Z(n2040) );
  NANDN U2406 ( .A(n2038), .B(n2037), .Z(n2039) );
  AND U2407 ( .A(n2040), .B(n2039), .Z(n2157) );
  XNOR U2408 ( .A(n2158), .B(n2157), .Z(n2159) );
  XOR U2409 ( .A(n2160), .B(n2159), .Z(n2154) );
  XNOR U2410 ( .A(n2153), .B(n2154), .Z(n2162) );
  XNOR U2411 ( .A(n2161), .B(n2162), .Z(n2163) );
  XOR U2412 ( .A(n2164), .B(n2163), .Z(n2058) );
  XNOR U2413 ( .A(n2057), .B(n2058), .Z(n2059) );
  XNOR U2414 ( .A(n2060), .B(n2059), .Z(n2052) );
  XNOR U2415 ( .A(n2051), .B(n2052), .Z(n2053) );
  XNOR U2416 ( .A(n2054), .B(n2053), .Z(n2046) );
  XNOR U2417 ( .A(n2046), .B(sreg[59]), .Z(n2048) );
  NAND U2418 ( .A(n2041), .B(sreg[58]), .Z(n2045) );
  OR U2419 ( .A(n2043), .B(n2042), .Z(n2044) );
  AND U2420 ( .A(n2045), .B(n2044), .Z(n2047) );
  XOR U2421 ( .A(n2048), .B(n2047), .Z(c[59]) );
  NAND U2422 ( .A(n2046), .B(sreg[59]), .Z(n2050) );
  OR U2423 ( .A(n2048), .B(n2047), .Z(n2049) );
  NAND U2424 ( .A(n2050), .B(n2049), .Z(n2292) );
  XNOR U2425 ( .A(n2292), .B(sreg[60]), .Z(n2294) );
  NANDN U2426 ( .A(n2052), .B(n2051), .Z(n2056) );
  NAND U2427 ( .A(n2054), .B(n2053), .Z(n2055) );
  NAND U2428 ( .A(n2056), .B(n2055), .Z(n2170) );
  NANDN U2429 ( .A(n2058), .B(n2057), .Z(n2062) );
  NAND U2430 ( .A(n2060), .B(n2059), .Z(n2061) );
  NAND U2431 ( .A(n2062), .B(n2061), .Z(n2168) );
  OR U2432 ( .A(n2064), .B(n2063), .Z(n2068) );
  NAND U2433 ( .A(n2066), .B(n2065), .Z(n2067) );
  NAND U2434 ( .A(n2068), .B(n2067), .Z(n2267) );
  NANDN U2435 ( .A(n2070), .B(n2069), .Z(n2074) );
  NANDN U2436 ( .A(n2072), .B(n2071), .Z(n2073) );
  NAND U2437 ( .A(n2074), .B(n2073), .Z(n2279) );
  NANDN U2438 ( .A(n2076), .B(n2075), .Z(n2080) );
  NAND U2439 ( .A(n2078), .B(n2077), .Z(n2079) );
  NAND U2440 ( .A(n2080), .B(n2079), .Z(n2276) );
  XOR U2441 ( .A(b[13]), .B(a[16]), .Z(n2210) );
  NAND U2442 ( .A(n2210), .B(n8730), .Z(n2083) );
  NAND U2443 ( .A(n2081), .B(n8731), .Z(n2082) );
  NAND U2444 ( .A(n2083), .B(n2082), .Z(n2222) );
  NANDN U2445 ( .A(n2084), .B(n9622), .Z(n2086) );
  XNOR U2446 ( .A(b[23]), .B(a[6]), .Z(n2245) );
  OR U2447 ( .A(n2245), .B(n9621), .Z(n2085) );
  NAND U2448 ( .A(n2086), .B(n2085), .Z(n2219) );
  XOR U2449 ( .A(b[3]), .B(n6500), .Z(n2228) );
  NANDN U2450 ( .A(n2228), .B(n7620), .Z(n2089) );
  NAND U2451 ( .A(n2087), .B(n7622), .Z(n2088) );
  AND U2452 ( .A(n2089), .B(n2088), .Z(n2220) );
  XNOR U2453 ( .A(n2219), .B(n2220), .Z(n2221) );
  XOR U2454 ( .A(n2222), .B(n2221), .Z(n2277) );
  XNOR U2455 ( .A(n2276), .B(n2277), .Z(n2278) );
  XOR U2456 ( .A(n2279), .B(n2278), .Z(n2264) );
  XOR U2457 ( .A(b[7]), .B(a[22]), .Z(n2235) );
  NANDN U2458 ( .A(n8013), .B(n2235), .Z(n2092) );
  NAND U2459 ( .A(n2090), .B(n8014), .Z(n2091) );
  NAND U2460 ( .A(n2092), .B(n2091), .Z(n2263) );
  NAND U2461 ( .A(n2093), .B(n9105), .Z(n2095) );
  XNOR U2462 ( .A(n9455), .B(a[12]), .Z(n2231) );
  NAND U2463 ( .A(n2231), .B(n9107), .Z(n2094) );
  NAND U2464 ( .A(n2095), .B(n2094), .Z(n2260) );
  XOR U2465 ( .A(b[11]), .B(a[18]), .Z(n2216) );
  NAND U2466 ( .A(n2216), .B(n8541), .Z(n2098) );
  NANDN U2467 ( .A(n2096), .B(n8542), .Z(n2097) );
  AND U2468 ( .A(n2098), .B(n2097), .Z(n2261) );
  XNOR U2469 ( .A(n2260), .B(n2261), .Z(n2262) );
  XNOR U2470 ( .A(n2263), .B(n2262), .Z(n2273) );
  XNOR U2471 ( .A(b[5]), .B(a[24]), .Z(n2225) );
  NANDN U2472 ( .A(n2225), .B(n7905), .Z(n2101) );
  NANDN U2473 ( .A(n2099), .B(n7906), .Z(n2100) );
  NAND U2474 ( .A(n2101), .B(n2100), .Z(n2244) );
  NAND U2475 ( .A(n2102), .B(n9379), .Z(n2104) );
  XNOR U2476 ( .A(n9562), .B(a[10]), .Z(n2213) );
  NAND U2477 ( .A(n2213), .B(n9378), .Z(n2103) );
  NAND U2478 ( .A(n2104), .B(n2103), .Z(n2241) );
  XOR U2479 ( .A(n318), .B(n3831), .Z(n2238) );
  NAND U2480 ( .A(n2238), .B(n9493), .Z(n2107) );
  NANDN U2481 ( .A(n2105), .B(n9495), .Z(n2106) );
  AND U2482 ( .A(n2107), .B(n2106), .Z(n2242) );
  XNOR U2483 ( .A(n2241), .B(n2242), .Z(n2243) );
  XNOR U2484 ( .A(n2244), .B(n2243), .Z(n2270) );
  NAND U2485 ( .A(n2108), .B(n8286), .Z(n2110) );
  XOR U2486 ( .A(b[9]), .B(a[20]), .Z(n2248) );
  NAND U2487 ( .A(n2248), .B(n8288), .Z(n2109) );
  NAND U2488 ( .A(n2110), .B(n2109), .Z(n2271) );
  XNOR U2489 ( .A(n2270), .B(n2271), .Z(n2272) );
  XOR U2490 ( .A(n2273), .B(n2272), .Z(n2265) );
  XNOR U2491 ( .A(n2264), .B(n2265), .Z(n2266) );
  XNOR U2492 ( .A(n2267), .B(n2266), .Z(n2291) );
  NANDN U2493 ( .A(n2116), .B(n2115), .Z(n2120) );
  NAND U2494 ( .A(n2118), .B(n2117), .Z(n2119) );
  NAND U2495 ( .A(n2120), .B(n2119), .Z(n2285) );
  NANDN U2496 ( .A(n315), .B(a[28]), .Z(n2121) );
  XNOR U2497 ( .A(b[1]), .B(n2121), .Z(n2123) );
  NANDN U2498 ( .A(b[0]), .B(a[27]), .Z(n2122) );
  AND U2499 ( .A(n2123), .B(n2122), .Z(n2256) );
  XNOR U2500 ( .A(b[28]), .B(b[27]), .Z(n9874) );
  ANDN U2501 ( .B(a[0]), .A(n9874), .Z(n2254) );
  XNOR U2502 ( .A(b[25]), .B(a[4]), .Z(n2251) );
  NANDN U2503 ( .A(n2251), .B(n9706), .Z(n2126) );
  NANDN U2504 ( .A(n2124), .B(n9707), .Z(n2125) );
  NAND U2505 ( .A(n2126), .B(n2125), .Z(n2255) );
  XNOR U2506 ( .A(n2254), .B(n2255), .Z(n2257) );
  XNOR U2507 ( .A(n2256), .B(n2257), .Z(n2283) );
  NANDN U2508 ( .A(n2127), .B(n8961), .Z(n2129) );
  XOR U2509 ( .A(b[15]), .B(a[14]), .Z(n2197) );
  NAND U2510 ( .A(n2197), .B(n8963), .Z(n2128) );
  NAND U2511 ( .A(n2129), .B(n2128), .Z(n2191) );
  NANDN U2512 ( .A(n2130), .B(n9801), .Z(n2132) );
  XOR U2513 ( .A(b[27]), .B(n2950), .Z(n2203) );
  OR U2514 ( .A(n2203), .B(n9751), .Z(n2131) );
  AND U2515 ( .A(n2132), .B(n2131), .Z(n2192) );
  XOR U2516 ( .A(n2191), .B(n2192), .Z(n2194) );
  NAND U2517 ( .A(n2134), .B(n2133), .Z(n2193) );
  XOR U2518 ( .A(n2194), .B(n2193), .Z(n2282) );
  XOR U2519 ( .A(n2283), .B(n2282), .Z(n2284) );
  XOR U2520 ( .A(n2285), .B(n2284), .Z(n2185) );
  NANDN U2521 ( .A(n2136), .B(n2135), .Z(n2140) );
  NANDN U2522 ( .A(n2138), .B(n2137), .Z(n2139) );
  AND U2523 ( .A(n2140), .B(n2139), .Z(n2186) );
  XNOR U2524 ( .A(n2185), .B(n2186), .Z(n2187) );
  XNOR U2525 ( .A(n2188), .B(n2187), .Z(n2288) );
  XNOR U2526 ( .A(n2288), .B(n2289), .Z(n2290) );
  XOR U2527 ( .A(n2291), .B(n2290), .Z(n2175) );
  NANDN U2528 ( .A(n2146), .B(n2145), .Z(n2150) );
  NAND U2529 ( .A(n2148), .B(n2147), .Z(n2149) );
  NAND U2530 ( .A(n2150), .B(n2149), .Z(n2182) );
  OR U2531 ( .A(n2152), .B(n2151), .Z(n2156) );
  NANDN U2532 ( .A(n2154), .B(n2153), .Z(n2155) );
  NAND U2533 ( .A(n2156), .B(n2155), .Z(n2180) );
  XNOR U2534 ( .A(n2180), .B(n2179), .Z(n2181) );
  XOR U2535 ( .A(n2182), .B(n2181), .Z(n2173) );
  NANDN U2536 ( .A(n2162), .B(n2161), .Z(n2166) );
  NAND U2537 ( .A(n2164), .B(n2163), .Z(n2165) );
  NAND U2538 ( .A(n2166), .B(n2165), .Z(n2174) );
  XNOR U2539 ( .A(n2173), .B(n2174), .Z(n2176) );
  XOR U2540 ( .A(n2175), .B(n2176), .Z(n2167) );
  XOR U2541 ( .A(n2168), .B(n2167), .Z(n2169) );
  XOR U2542 ( .A(n2170), .B(n2169), .Z(n2293) );
  XOR U2543 ( .A(n2294), .B(n2293), .Z(c[60]) );
  NAND U2544 ( .A(n2168), .B(n2167), .Z(n2172) );
  NAND U2545 ( .A(n2170), .B(n2169), .Z(n2171) );
  NAND U2546 ( .A(n2172), .B(n2171), .Z(n2305) );
  NANDN U2547 ( .A(n2174), .B(n2173), .Z(n2178) );
  NAND U2548 ( .A(n2176), .B(n2175), .Z(n2177) );
  NAND U2549 ( .A(n2178), .B(n2177), .Z(n2302) );
  NANDN U2550 ( .A(n2180), .B(n2179), .Z(n2184) );
  NANDN U2551 ( .A(n2182), .B(n2181), .Z(n2183) );
  NAND U2552 ( .A(n2184), .B(n2183), .Z(n2424) );
  NANDN U2553 ( .A(n2186), .B(n2185), .Z(n2190) );
  NAND U2554 ( .A(n2188), .B(n2187), .Z(n2189) );
  NAND U2555 ( .A(n2190), .B(n2189), .Z(n2317) );
  NANDN U2556 ( .A(n2192), .B(n2191), .Z(n2196) );
  OR U2557 ( .A(n2194), .B(n2193), .Z(n2195) );
  NAND U2558 ( .A(n2196), .B(n2195), .Z(n2377) );
  NAND U2559 ( .A(n2197), .B(n8961), .Z(n2199) );
  XOR U2560 ( .A(b[15]), .B(a[15]), .Z(n2340) );
  NAND U2561 ( .A(n2340), .B(n8963), .Z(n2198) );
  NAND U2562 ( .A(n2199), .B(n2198), .Z(n2366) );
  NANDN U2563 ( .A(n315), .B(a[29]), .Z(n2200) );
  XNOR U2564 ( .A(b[1]), .B(n2200), .Z(n2202) );
  NANDN U2565 ( .A(b[0]), .B(a[28]), .Z(n2201) );
  AND U2566 ( .A(n2202), .B(n2201), .Z(n2364) );
  NANDN U2567 ( .A(n2203), .B(n9801), .Z(n2205) );
  XOR U2568 ( .A(b[27]), .B(n3094), .Z(n2383) );
  OR U2569 ( .A(n2383), .B(n9751), .Z(n2204) );
  NAND U2570 ( .A(n2205), .B(n2204), .Z(n2332) );
  XNOR U2571 ( .A(n2616), .B(b[29]), .Z(n2207) );
  XOR U2572 ( .A(b[28]), .B(b[29]), .Z(n2206) );
  AND U2573 ( .A(n2206), .B(n9874), .Z(n9875) );
  NAND U2574 ( .A(n2207), .B(n9875), .Z(n2209) );
  XNOR U2575 ( .A(b[29]), .B(a[1]), .Z(n2337) );
  NOR U2576 ( .A(n9874), .B(n2337), .Z(n2208) );
  ANDN U2577 ( .B(n2209), .A(n2208), .Z(n2333) );
  XNOR U2578 ( .A(n2332), .B(n2333), .Z(n2365) );
  XOR U2579 ( .A(n2364), .B(n2365), .Z(n2367) );
  XOR U2580 ( .A(n2366), .B(n2367), .Z(n2374) );
  XNOR U2581 ( .A(b[13]), .B(a[17]), .Z(n2355) );
  NANDN U2582 ( .A(n2355), .B(n8730), .Z(n2212) );
  NAND U2583 ( .A(n2210), .B(n8731), .Z(n2211) );
  NAND U2584 ( .A(n2212), .B(n2211), .Z(n2373) );
  NAND U2585 ( .A(n2213), .B(n9379), .Z(n2215) );
  XNOR U2586 ( .A(n9562), .B(a[11]), .Z(n2358) );
  NAND U2587 ( .A(n2358), .B(n9378), .Z(n2214) );
  NAND U2588 ( .A(n2215), .B(n2214), .Z(n2370) );
  XOR U2589 ( .A(b[11]), .B(a[19]), .Z(n2352) );
  NAND U2590 ( .A(n2352), .B(n8541), .Z(n2218) );
  NAND U2591 ( .A(n2216), .B(n8542), .Z(n2217) );
  AND U2592 ( .A(n2218), .B(n2217), .Z(n2371) );
  XNOR U2593 ( .A(n2370), .B(n2371), .Z(n2372) );
  XNOR U2594 ( .A(n2373), .B(n2372), .Z(n2375) );
  XNOR U2595 ( .A(n2374), .B(n2375), .Z(n2376) );
  XNOR U2596 ( .A(n2377), .B(n2376), .Z(n2412) );
  NANDN U2597 ( .A(n2220), .B(n2219), .Z(n2224) );
  NAND U2598 ( .A(n2222), .B(n2221), .Z(n2223) );
  NAND U2599 ( .A(n2224), .B(n2223), .Z(n2410) );
  XNOR U2600 ( .A(b[5]), .B(a[25]), .Z(n2346) );
  NANDN U2601 ( .A(n2346), .B(n7905), .Z(n2227) );
  NANDN U2602 ( .A(n2225), .B(n7906), .Z(n2226) );
  NAND U2603 ( .A(n2227), .B(n2226), .Z(n2398) );
  NANDN U2604 ( .A(n2228), .B(n7622), .Z(n2230) );
  XNOR U2605 ( .A(n316), .B(a[27]), .Z(n2343) );
  NAND U2606 ( .A(n2343), .B(n7620), .Z(n2229) );
  NAND U2607 ( .A(n2230), .B(n2229), .Z(n2395) );
  NAND U2608 ( .A(n2231), .B(n9105), .Z(n2233) );
  XNOR U2609 ( .A(n9455), .B(a[13]), .Z(n2334) );
  NAND U2610 ( .A(n2334), .B(n9107), .Z(n2232) );
  NAND U2611 ( .A(n2233), .B(n2232), .Z(n2396) );
  XOR U2612 ( .A(n2395), .B(n2396), .Z(n2397) );
  XOR U2613 ( .A(n2398), .B(n2397), .Z(n2415) );
  NANDN U2614 ( .A(n321), .B(b[28]), .Z(n2234) );
  ANDN U2615 ( .B(n2234), .A(n322), .Z(n9917) );
  NANDN U2616 ( .A(n2254), .B(n9917), .Z(n2405) );
  XNOR U2617 ( .A(b[7]), .B(a[23]), .Z(n2361) );
  OR U2618 ( .A(n2361), .B(n8013), .Z(n2237) );
  NAND U2619 ( .A(n8014), .B(n2235), .Z(n2236) );
  NAND U2620 ( .A(n2237), .B(n2236), .Z(n2406) );
  XNOR U2621 ( .A(n2405), .B(n2406), .Z(n2407) );
  XNOR U2622 ( .A(b[21]), .B(a[9]), .Z(n2392) );
  NANDN U2623 ( .A(n2392), .B(n9493), .Z(n2240) );
  NAND U2624 ( .A(n9495), .B(n2238), .Z(n2239) );
  AND U2625 ( .A(n2240), .B(n2239), .Z(n2408) );
  XNOR U2626 ( .A(n2407), .B(n2408), .Z(n2416) );
  XNOR U2627 ( .A(n2415), .B(n2416), .Z(n2418) );
  XOR U2628 ( .A(n2418), .B(n2417), .Z(n2409) );
  XNOR U2629 ( .A(n2410), .B(n2409), .Z(n2411) );
  XOR U2630 ( .A(n2412), .B(n2411), .Z(n2315) );
  NANDN U2631 ( .A(n2245), .B(n9622), .Z(n2247) );
  XNOR U2632 ( .A(b[23]), .B(a[7]), .Z(n2386) );
  OR U2633 ( .A(n2386), .B(n9621), .Z(n2246) );
  NAND U2634 ( .A(n2247), .B(n2246), .Z(n2404) );
  NAND U2635 ( .A(n2248), .B(n8286), .Z(n2250) );
  XOR U2636 ( .A(b[9]), .B(a[21]), .Z(n2349) );
  NAND U2637 ( .A(n2349), .B(n8288), .Z(n2249) );
  NAND U2638 ( .A(n2250), .B(n2249), .Z(n2401) );
  XOR U2639 ( .A(b[25]), .B(n3389), .Z(n2389) );
  NANDN U2640 ( .A(n2389), .B(n9706), .Z(n2253) );
  NANDN U2641 ( .A(n2251), .B(n9707), .Z(n2252) );
  AND U2642 ( .A(n2253), .B(n2252), .Z(n2402) );
  XNOR U2643 ( .A(n2401), .B(n2402), .Z(n2403) );
  XNOR U2644 ( .A(n2404), .B(n2403), .Z(n2326) );
  NAND U2645 ( .A(n2255), .B(n2254), .Z(n2259) );
  NANDN U2646 ( .A(n2257), .B(n2256), .Z(n2258) );
  NAND U2647 ( .A(n2259), .B(n2258), .Z(n2327) );
  XOR U2648 ( .A(n2326), .B(n2327), .Z(n2329) );
  XOR U2649 ( .A(n2329), .B(n2328), .Z(n2314) );
  XOR U2650 ( .A(n2315), .B(n2314), .Z(n2316) );
  XNOR U2651 ( .A(n2317), .B(n2316), .Z(n2311) );
  NANDN U2652 ( .A(n2265), .B(n2264), .Z(n2269) );
  NAND U2653 ( .A(n2267), .B(n2266), .Z(n2268) );
  NAND U2654 ( .A(n2269), .B(n2268), .Z(n2309) );
  NANDN U2655 ( .A(n2271), .B(n2270), .Z(n2275) );
  NAND U2656 ( .A(n2273), .B(n2272), .Z(n2274) );
  NAND U2657 ( .A(n2275), .B(n2274), .Z(n2323) );
  NANDN U2658 ( .A(n2277), .B(n2276), .Z(n2281) );
  NANDN U2659 ( .A(n2279), .B(n2278), .Z(n2280) );
  NAND U2660 ( .A(n2281), .B(n2280), .Z(n2320) );
  OR U2661 ( .A(n2283), .B(n2282), .Z(n2287) );
  NANDN U2662 ( .A(n2285), .B(n2284), .Z(n2286) );
  AND U2663 ( .A(n2287), .B(n2286), .Z(n2321) );
  XNOR U2664 ( .A(n2320), .B(n2321), .Z(n2322) );
  XOR U2665 ( .A(n2323), .B(n2322), .Z(n2308) );
  XNOR U2666 ( .A(n2309), .B(n2308), .Z(n2310) );
  XOR U2667 ( .A(n2311), .B(n2310), .Z(n2421) );
  XOR U2668 ( .A(n2421), .B(n2422), .Z(n2423) );
  XOR U2669 ( .A(n2424), .B(n2423), .Z(n2303) );
  XNOR U2670 ( .A(n2302), .B(n2303), .Z(n2304) );
  XNOR U2671 ( .A(n2305), .B(n2304), .Z(n2297) );
  XNOR U2672 ( .A(n2297), .B(sreg[61]), .Z(n2299) );
  NAND U2673 ( .A(n2292), .B(sreg[60]), .Z(n2296) );
  OR U2674 ( .A(n2294), .B(n2293), .Z(n2295) );
  AND U2675 ( .A(n2296), .B(n2295), .Z(n2298) );
  XOR U2676 ( .A(n2299), .B(n2298), .Z(c[61]) );
  NAND U2677 ( .A(n2297), .B(sreg[61]), .Z(n2301) );
  OR U2678 ( .A(n2299), .B(n2298), .Z(n2300) );
  NAND U2679 ( .A(n2301), .B(n2300), .Z(n2560) );
  XNOR U2680 ( .A(n2560), .B(sreg[62]), .Z(n2562) );
  NANDN U2681 ( .A(n2303), .B(n2302), .Z(n2307) );
  NAND U2682 ( .A(n2305), .B(n2304), .Z(n2306) );
  NAND U2683 ( .A(n2307), .B(n2306), .Z(n2430) );
  NANDN U2684 ( .A(n2309), .B(n2308), .Z(n2313) );
  NAND U2685 ( .A(n2311), .B(n2310), .Z(n2312) );
  NAND U2686 ( .A(n2313), .B(n2312), .Z(n2436) );
  OR U2687 ( .A(n2315), .B(n2314), .Z(n2319) );
  NAND U2688 ( .A(n2317), .B(n2316), .Z(n2318) );
  NAND U2689 ( .A(n2319), .B(n2318), .Z(n2433) );
  NANDN U2690 ( .A(n2321), .B(n2320), .Z(n2325) );
  NAND U2691 ( .A(n2323), .B(n2322), .Z(n2324) );
  NAND U2692 ( .A(n2325), .B(n2324), .Z(n2439) );
  NANDN U2693 ( .A(n2327), .B(n2326), .Z(n2331) );
  OR U2694 ( .A(n2329), .B(n2328), .Z(n2330) );
  NAND U2695 ( .A(n2331), .B(n2330), .Z(n2481) );
  NANDN U2696 ( .A(n2333), .B(n2332), .Z(n2515) );
  NAND U2697 ( .A(n2334), .B(n9105), .Z(n2336) );
  XNOR U2698 ( .A(n9455), .B(a[14]), .Z(n2509) );
  NAND U2699 ( .A(n2509), .B(n9107), .Z(n2335) );
  NAND U2700 ( .A(n2336), .B(n2335), .Z(n2514) );
  NANDN U2701 ( .A(n2337), .B(n9875), .Z(n2339) );
  XNOR U2702 ( .A(n322), .B(a[2]), .Z(n2449) );
  NANDN U2703 ( .A(n9874), .B(n2449), .Z(n2338) );
  AND U2704 ( .A(n2339), .B(n2338), .Z(n2513) );
  XNOR U2705 ( .A(n2514), .B(n2513), .Z(n2516) );
  XNOR U2706 ( .A(n2515), .B(n2516), .Z(n2486) );
  NAND U2707 ( .A(n2340), .B(n8961), .Z(n2342) );
  XOR U2708 ( .A(b[15]), .B(a[16]), .Z(n2460) );
  NAND U2709 ( .A(n2460), .B(n8963), .Z(n2341) );
  NAND U2710 ( .A(n2342), .B(n2341), .Z(n2529) );
  NAND U2711 ( .A(n2343), .B(n7622), .Z(n2345) );
  XNOR U2712 ( .A(n316), .B(a[28]), .Z(n2506) );
  NAND U2713 ( .A(n2506), .B(n7620), .Z(n2344) );
  NAND U2714 ( .A(n2345), .B(n2344), .Z(n2527) );
  XOR U2715 ( .A(b[5]), .B(n6500), .Z(n2503) );
  NANDN U2716 ( .A(n2503), .B(n7905), .Z(n2348) );
  NANDN U2717 ( .A(n2346), .B(n7906), .Z(n2347) );
  AND U2718 ( .A(n2348), .B(n2347), .Z(n2528) );
  XOR U2719 ( .A(n2527), .B(n2528), .Z(n2530) );
  XNOR U2720 ( .A(n2529), .B(n2530), .Z(n2485) );
  XOR U2721 ( .A(n2486), .B(n2485), .Z(n2487) );
  NAND U2722 ( .A(n2349), .B(n8286), .Z(n2351) );
  XOR U2723 ( .A(b[9]), .B(a[22]), .Z(n2533) );
  NAND U2724 ( .A(n2533), .B(n8288), .Z(n2350) );
  NAND U2725 ( .A(n2351), .B(n2350), .Z(n2517) );
  XOR U2726 ( .A(b[11]), .B(a[20]), .Z(n2551) );
  NAND U2727 ( .A(n2551), .B(n8541), .Z(n2354) );
  NAND U2728 ( .A(n2352), .B(n8542), .Z(n2353) );
  AND U2729 ( .A(n2354), .B(n2353), .Z(n2518) );
  XNOR U2730 ( .A(n2517), .B(n2518), .Z(n2519) );
  XOR U2731 ( .A(b[13]), .B(a[18]), .Z(n2536) );
  NAND U2732 ( .A(n2536), .B(n8730), .Z(n2357) );
  NANDN U2733 ( .A(n2355), .B(n8731), .Z(n2356) );
  NAND U2734 ( .A(n2357), .B(n2356), .Z(n2448) );
  NAND U2735 ( .A(n2358), .B(n9379), .Z(n2360) );
  XNOR U2736 ( .A(n9562), .B(a[12]), .Z(n2500) );
  NAND U2737 ( .A(n2500), .B(n9378), .Z(n2359) );
  NAND U2738 ( .A(n2360), .B(n2359), .Z(n2445) );
  XOR U2739 ( .A(b[7]), .B(a[24]), .Z(n2497) );
  NANDN U2740 ( .A(n8013), .B(n2497), .Z(n2363) );
  NANDN U2741 ( .A(n2361), .B(n8014), .Z(n2362) );
  AND U2742 ( .A(n2363), .B(n2362), .Z(n2446) );
  XNOR U2743 ( .A(n2445), .B(n2446), .Z(n2447) );
  XNOR U2744 ( .A(n2448), .B(n2447), .Z(n2520) );
  XNOR U2745 ( .A(n2519), .B(n2520), .Z(n2488) );
  XNOR U2746 ( .A(n2487), .B(n2488), .Z(n2471) );
  NAND U2747 ( .A(n2365), .B(n2364), .Z(n2369) );
  NAND U2748 ( .A(n2367), .B(n2366), .Z(n2368) );
  NAND U2749 ( .A(n2369), .B(n2368), .Z(n2470) );
  XNOR U2750 ( .A(n2470), .B(n2469), .Z(n2472) );
  XNOR U2751 ( .A(n2471), .B(n2472), .Z(n2479) );
  NANDN U2752 ( .A(n2375), .B(n2374), .Z(n2379) );
  NAND U2753 ( .A(n2377), .B(n2376), .Z(n2378) );
  AND U2754 ( .A(n2379), .B(n2378), .Z(n2480) );
  XOR U2755 ( .A(n2479), .B(n2480), .Z(n2482) );
  XOR U2756 ( .A(n2481), .B(n2482), .Z(n2440) );
  XNOR U2757 ( .A(n2439), .B(n2440), .Z(n2441) );
  NANDN U2758 ( .A(n315), .B(a[30]), .Z(n2380) );
  XNOR U2759 ( .A(b[1]), .B(n2380), .Z(n2382) );
  NANDN U2760 ( .A(b[0]), .B(a[29]), .Z(n2381) );
  AND U2761 ( .A(n2382), .B(n2381), .Z(n2465) );
  NANDN U2762 ( .A(n2383), .B(n9801), .Z(n2385) );
  XNOR U2763 ( .A(b[27]), .B(a[4]), .Z(n2548) );
  OR U2764 ( .A(n2548), .B(n9751), .Z(n2384) );
  NAND U2765 ( .A(n2385), .B(n2384), .Z(n2463) );
  IV U2766 ( .A(b[30]), .Z(n2512) );
  XOR U2767 ( .A(b[29]), .B(n2512), .Z(n9913) );
  OR U2768 ( .A(n9913), .B(n2616), .Z(n2464) );
  XNOR U2769 ( .A(n2463), .B(n2464), .Z(n2466) );
  XOR U2770 ( .A(n2465), .B(n2466), .Z(n2493) );
  NANDN U2771 ( .A(n2386), .B(n9622), .Z(n2388) );
  XOR U2772 ( .A(b[23]), .B(n3831), .Z(n2542) );
  OR U2773 ( .A(n2542), .B(n9621), .Z(n2387) );
  NAND U2774 ( .A(n2388), .B(n2387), .Z(n2524) );
  XNOR U2775 ( .A(b[25]), .B(a[6]), .Z(n2545) );
  NANDN U2776 ( .A(n2545), .B(n9706), .Z(n2391) );
  NANDN U2777 ( .A(n2389), .B(n9707), .Z(n2390) );
  NAND U2778 ( .A(n2391), .B(n2390), .Z(n2521) );
  XNOR U2779 ( .A(b[21]), .B(a[10]), .Z(n2539) );
  NANDN U2780 ( .A(n2539), .B(n9493), .Z(n2394) );
  NANDN U2781 ( .A(n2392), .B(n9495), .Z(n2393) );
  AND U2782 ( .A(n2394), .B(n2393), .Z(n2522) );
  XNOR U2783 ( .A(n2521), .B(n2522), .Z(n2523) );
  XNOR U2784 ( .A(n2524), .B(n2523), .Z(n2491) );
  NAND U2785 ( .A(n2396), .B(n2395), .Z(n2400) );
  NAND U2786 ( .A(n2398), .B(n2397), .Z(n2399) );
  NAND U2787 ( .A(n2400), .B(n2399), .Z(n2492) );
  XOR U2788 ( .A(n2491), .B(n2492), .Z(n2494) );
  XOR U2789 ( .A(n2493), .B(n2494), .Z(n2476) );
  XNOR U2790 ( .A(n2473), .B(n2474), .Z(n2475) );
  XNOR U2791 ( .A(n2476), .B(n2475), .Z(n2557) );
  NANDN U2792 ( .A(n2410), .B(n2409), .Z(n2414) );
  NAND U2793 ( .A(n2412), .B(n2411), .Z(n2413) );
  NAND U2794 ( .A(n2414), .B(n2413), .Z(n2554) );
  OR U2795 ( .A(n2416), .B(n2415), .Z(n2420) );
  OR U2796 ( .A(n2418), .B(n2417), .Z(n2419) );
  AND U2797 ( .A(n2420), .B(n2419), .Z(n2555) );
  XNOR U2798 ( .A(n2554), .B(n2555), .Z(n2556) );
  XOR U2799 ( .A(n2557), .B(n2556), .Z(n2442) );
  XNOR U2800 ( .A(n2441), .B(n2442), .Z(n2434) );
  XNOR U2801 ( .A(n2433), .B(n2434), .Z(n2435) );
  XOR U2802 ( .A(n2436), .B(n2435), .Z(n2427) );
  OR U2803 ( .A(n2422), .B(n2421), .Z(n2426) );
  NAND U2804 ( .A(n2424), .B(n2423), .Z(n2425) );
  NAND U2805 ( .A(n2426), .B(n2425), .Z(n2428) );
  XNOR U2806 ( .A(n2427), .B(n2428), .Z(n2429) );
  XOR U2807 ( .A(n2430), .B(n2429), .Z(n2561) );
  XOR U2808 ( .A(n2562), .B(n2561), .Z(c[62]) );
  NANDN U2809 ( .A(n2428), .B(n2427), .Z(n2432) );
  NAND U2810 ( .A(n2430), .B(n2429), .Z(n2431) );
  NAND U2811 ( .A(n2432), .B(n2431), .Z(n2573) );
  NANDN U2812 ( .A(n2434), .B(n2433), .Z(n2438) );
  NANDN U2813 ( .A(n2436), .B(n2435), .Z(n2437) );
  NAND U2814 ( .A(n2438), .B(n2437), .Z(n2570) );
  NANDN U2815 ( .A(n2440), .B(n2439), .Z(n2444) );
  NANDN U2816 ( .A(n2442), .B(n2441), .Z(n2443) );
  NAND U2817 ( .A(n2444), .B(n2443), .Z(n2704) );
  NAND U2818 ( .A(n2449), .B(n9875), .Z(n2451) );
  XOR U2819 ( .A(n322), .B(n3094), .Z(n2613) );
  NANDN U2820 ( .A(n9874), .B(n2613), .Z(n2450) );
  NAND U2821 ( .A(n2451), .B(n2450), .Z(n2685) );
  XNOR U2822 ( .A(n323), .B(a[0]), .Z(n2454) );
  XNOR U2823 ( .A(n323), .B(b[29]), .Z(n2453) );
  XNOR U2824 ( .A(n323), .B(b[30]), .Z(n2452) );
  AND U2825 ( .A(n2453), .B(n2452), .Z(n9914) );
  NAND U2826 ( .A(n2454), .B(n9914), .Z(n2456) );
  XNOR U2827 ( .A(n323), .B(a[1]), .Z(n2695) );
  NANDN U2828 ( .A(n9913), .B(n2695), .Z(n2455) );
  NAND U2829 ( .A(n2456), .B(n2455), .Z(n2684) );
  XNOR U2830 ( .A(n2685), .B(n2684), .Z(n2606) );
  NANDN U2831 ( .A(n315), .B(a[31]), .Z(n2457) );
  XNOR U2832 ( .A(b[1]), .B(n2457), .Z(n2459) );
  IV U2833 ( .A(a[30]), .Z(n6135) );
  NANDN U2834 ( .A(n6135), .B(n315), .Z(n2458) );
  AND U2835 ( .A(n2459), .B(n2458), .Z(n2605) );
  NAND U2836 ( .A(n2460), .B(n8961), .Z(n2462) );
  XNOR U2837 ( .A(b[15]), .B(n5168), .Z(n2620) );
  NAND U2838 ( .A(n2620), .B(n8963), .Z(n2461) );
  NAND U2839 ( .A(n2462), .B(n2461), .Z(n2604) );
  XOR U2840 ( .A(n2605), .B(n2604), .Z(n2607) );
  XNOR U2841 ( .A(n2606), .B(n2607), .Z(n2638) );
  NANDN U2842 ( .A(n2464), .B(n2463), .Z(n2468) );
  NAND U2843 ( .A(n2466), .B(n2465), .Z(n2467) );
  AND U2844 ( .A(n2468), .B(n2467), .Z(n2639) );
  XNOR U2845 ( .A(n2638), .B(n2639), .Z(n2640) );
  XNOR U2846 ( .A(n2641), .B(n2640), .Z(n2580) );
  XOR U2847 ( .A(n2580), .B(n2581), .Z(n2583) );
  NANDN U2848 ( .A(n2474), .B(n2473), .Z(n2478) );
  NANDN U2849 ( .A(n2476), .B(n2475), .Z(n2477) );
  NAND U2850 ( .A(n2478), .B(n2477), .Z(n2582) );
  XNOR U2851 ( .A(n2583), .B(n2582), .Z(n2579) );
  NANDN U2852 ( .A(n2480), .B(n2479), .Z(n2484) );
  OR U2853 ( .A(n2482), .B(n2481), .Z(n2483) );
  NAND U2854 ( .A(n2484), .B(n2483), .Z(n2577) );
  NAND U2855 ( .A(n2486), .B(n2485), .Z(n2490) );
  NAND U2856 ( .A(n2488), .B(n2487), .Z(n2489) );
  NAND U2857 ( .A(n2490), .B(n2489), .Z(n2586) );
  NANDN U2858 ( .A(n2492), .B(n2491), .Z(n2496) );
  OR U2859 ( .A(n2494), .B(n2493), .Z(n2495) );
  NAND U2860 ( .A(n2496), .B(n2495), .Z(n2587) );
  XNOR U2861 ( .A(n2586), .B(n2587), .Z(n2588) );
  XOR U2862 ( .A(b[7]), .B(a[25]), .Z(n2663) );
  NANDN U2863 ( .A(n8013), .B(n2663), .Z(n2499) );
  NAND U2864 ( .A(n2497), .B(n8014), .Z(n2498) );
  NAND U2865 ( .A(n2499), .B(n2498), .Z(n2681) );
  NAND U2866 ( .A(n2500), .B(n9379), .Z(n2502) );
  XNOR U2867 ( .A(n9562), .B(a[13]), .Z(n2666) );
  NAND U2868 ( .A(n2666), .B(n9378), .Z(n2501) );
  NAND U2869 ( .A(n2502), .B(n2501), .Z(n2678) );
  XNOR U2870 ( .A(b[5]), .B(a[27]), .Z(n2669) );
  NANDN U2871 ( .A(n2669), .B(n7905), .Z(n2505) );
  NANDN U2872 ( .A(n2503), .B(n7906), .Z(n2504) );
  AND U2873 ( .A(n2505), .B(n2504), .Z(n2679) );
  XNOR U2874 ( .A(n2678), .B(n2679), .Z(n2680) );
  XNOR U2875 ( .A(n2681), .B(n2680), .Z(n2633) );
  NAND U2876 ( .A(n2506), .B(n7622), .Z(n2508) );
  XNOR U2877 ( .A(n316), .B(a[29]), .Z(n2686) );
  NAND U2878 ( .A(n2686), .B(n7620), .Z(n2507) );
  NAND U2879 ( .A(n2508), .B(n2507), .Z(n2600) );
  NAND U2880 ( .A(n2509), .B(n9105), .Z(n2511) );
  XNOR U2881 ( .A(n9455), .B(a[15]), .Z(n2689) );
  NAND U2882 ( .A(n2689), .B(n9107), .Z(n2510) );
  NAND U2883 ( .A(n2511), .B(n2510), .Z(n2598) );
  XOR U2884 ( .A(n2598), .B(n2599), .Z(n2601) );
  XNOR U2885 ( .A(n2600), .B(n2601), .Z(n2632) );
  XNOR U2886 ( .A(n2633), .B(n2632), .Z(n2634) );
  XNOR U2887 ( .A(n2634), .B(n2635), .Z(n2593) );
  NANDN U2888 ( .A(n2522), .B(n2521), .Z(n2526) );
  NAND U2889 ( .A(n2524), .B(n2523), .Z(n2525) );
  NAND U2890 ( .A(n2526), .B(n2525), .Z(n2642) );
  NANDN U2891 ( .A(n2528), .B(n2527), .Z(n2532) );
  NANDN U2892 ( .A(n2530), .B(n2529), .Z(n2531) );
  AND U2893 ( .A(n2532), .B(n2531), .Z(n2643) );
  XNOR U2894 ( .A(n2642), .B(n2643), .Z(n2644) );
  XNOR U2895 ( .A(n2645), .B(n2644), .Z(n2592) );
  XNOR U2896 ( .A(n2593), .B(n2592), .Z(n2595) );
  NAND U2897 ( .A(n2533), .B(n8286), .Z(n2535) );
  XNOR U2898 ( .A(b[9]), .B(n6044), .Z(n2692) );
  NAND U2899 ( .A(n2692), .B(n8288), .Z(n2534) );
  NAND U2900 ( .A(n2535), .B(n2534), .Z(n2628) );
  XOR U2901 ( .A(b[13]), .B(a[19]), .Z(n2617) );
  NAND U2902 ( .A(n2617), .B(n8730), .Z(n2538) );
  NAND U2903 ( .A(n2536), .B(n8731), .Z(n2537) );
  NAND U2904 ( .A(n2538), .B(n2537), .Z(n2626) );
  XNOR U2905 ( .A(b[21]), .B(a[11]), .Z(n2623) );
  NANDN U2906 ( .A(n2623), .B(n9493), .Z(n2541) );
  NANDN U2907 ( .A(n2539), .B(n9495), .Z(n2540) );
  AND U2908 ( .A(n2541), .B(n2540), .Z(n2627) );
  XNOR U2909 ( .A(n2626), .B(n2627), .Z(n2629) );
  XOR U2910 ( .A(n2628), .B(n2629), .Z(n2650) );
  NANDN U2911 ( .A(n2542), .B(n9622), .Z(n2544) );
  XNOR U2912 ( .A(b[23]), .B(a[9]), .Z(n2698) );
  OR U2913 ( .A(n2698), .B(n9621), .Z(n2543) );
  NAND U2914 ( .A(n2544), .B(n2543), .Z(n2675) );
  XNOR U2915 ( .A(b[25]), .B(a[7]), .Z(n2657) );
  NANDN U2916 ( .A(n2657), .B(n9706), .Z(n2547) );
  NANDN U2917 ( .A(n2545), .B(n9707), .Z(n2546) );
  NAND U2918 ( .A(n2547), .B(n2546), .Z(n2672) );
  NANDN U2919 ( .A(n2548), .B(n9801), .Z(n2550) );
  XOR U2920 ( .A(b[27]), .B(n3389), .Z(n2660) );
  OR U2921 ( .A(n2660), .B(n9751), .Z(n2549) );
  AND U2922 ( .A(n2550), .B(n2549), .Z(n2673) );
  XNOR U2923 ( .A(n2672), .B(n2673), .Z(n2674) );
  XNOR U2924 ( .A(n2675), .B(n2674), .Z(n2648) );
  XOR U2925 ( .A(b[11]), .B(a[21]), .Z(n2654) );
  NAND U2926 ( .A(n8541), .B(n2654), .Z(n2553) );
  NAND U2927 ( .A(n8542), .B(n2551), .Z(n2552) );
  NAND U2928 ( .A(n2553), .B(n2552), .Z(n2649) );
  XOR U2929 ( .A(n2648), .B(n2649), .Z(n2651) );
  XOR U2930 ( .A(n2650), .B(n2651), .Z(n2594) );
  XNOR U2931 ( .A(n2595), .B(n2594), .Z(n2589) );
  XNOR U2932 ( .A(n2588), .B(n2589), .Z(n2576) );
  XOR U2933 ( .A(n2577), .B(n2576), .Z(n2578) );
  XNOR U2934 ( .A(n2579), .B(n2578), .Z(n2701) );
  NANDN U2935 ( .A(n2555), .B(n2554), .Z(n2559) );
  NANDN U2936 ( .A(n2557), .B(n2556), .Z(n2558) );
  AND U2937 ( .A(n2559), .B(n2558), .Z(n2702) );
  XNOR U2938 ( .A(n2701), .B(n2702), .Z(n2703) );
  XNOR U2939 ( .A(n2704), .B(n2703), .Z(n2571) );
  XOR U2940 ( .A(n2570), .B(n2571), .Z(n2572) );
  XNOR U2941 ( .A(n2573), .B(n2572), .Z(n2565) );
  XNOR U2942 ( .A(n2565), .B(sreg[63]), .Z(n2567) );
  NAND U2943 ( .A(n2560), .B(sreg[62]), .Z(n2564) );
  OR U2944 ( .A(n2562), .B(n2561), .Z(n2563) );
  AND U2945 ( .A(n2564), .B(n2563), .Z(n2566) );
  XOR U2946 ( .A(n2567), .B(n2566), .Z(c[63]) );
  NAND U2947 ( .A(n2565), .B(sreg[63]), .Z(n2569) );
  OR U2948 ( .A(n2567), .B(n2566), .Z(n2568) );
  NAND U2949 ( .A(n2569), .B(n2568), .Z(n2845) );
  XNOR U2950 ( .A(n2845), .B(sreg[64]), .Z(n2847) );
  OR U2951 ( .A(n2571), .B(n2570), .Z(n2575) );
  NAND U2952 ( .A(n2573), .B(n2572), .Z(n2574) );
  NAND U2953 ( .A(n2575), .B(n2574), .Z(n2708) );
  NANDN U2954 ( .A(n2581), .B(n2580), .Z(n2585) );
  OR U2955 ( .A(n2583), .B(n2582), .Z(n2584) );
  NAND U2956 ( .A(n2585), .B(n2584), .Z(n2842) );
  NANDN U2957 ( .A(n2587), .B(n2586), .Z(n2591) );
  NANDN U2958 ( .A(n2589), .B(n2588), .Z(n2590) );
  NAND U2959 ( .A(n2591), .B(n2590), .Z(n2711) );
  OR U2960 ( .A(n2593), .B(n2592), .Z(n2597) );
  OR U2961 ( .A(n2595), .B(n2594), .Z(n2596) );
  AND U2962 ( .A(n2597), .B(n2596), .Z(n2712) );
  XNOR U2963 ( .A(n2711), .B(n2712), .Z(n2713) );
  NANDN U2964 ( .A(n2599), .B(n2598), .Z(n2603) );
  NANDN U2965 ( .A(n2601), .B(n2600), .Z(n2602) );
  NAND U2966 ( .A(n2603), .B(n2602), .Z(n2723) );
  OR U2967 ( .A(n2605), .B(n2604), .Z(n2609) );
  NAND U2968 ( .A(n2607), .B(n2606), .Z(n2608) );
  NAND U2969 ( .A(n2609), .B(n2608), .Z(n2724) );
  XNOR U2970 ( .A(n2723), .B(n2724), .Z(n2725) );
  NANDN U2971 ( .A(n315), .B(a[32]), .Z(n2610) );
  XNOR U2972 ( .A(b[1]), .B(n2610), .Z(n2612) );
  NANDN U2973 ( .A(b[0]), .B(a[31]), .Z(n2611) );
  AND U2974 ( .A(n2612), .B(n2611), .Z(n2778) );
  NAND U2975 ( .A(n9875), .B(n2613), .Z(n2615) );
  XNOR U2976 ( .A(n322), .B(a[4]), .Z(n2763) );
  NANDN U2977 ( .A(n9874), .B(n2763), .Z(n2614) );
  AND U2978 ( .A(n2615), .B(n2614), .Z(n2779) );
  XOR U2979 ( .A(n2778), .B(n2779), .Z(n2781) );
  NANDN U2980 ( .A(n2616), .B(b[31]), .Z(n2780) );
  XOR U2981 ( .A(n2781), .B(n2780), .Z(n2835) );
  XOR U2982 ( .A(b[13]), .B(a[20]), .Z(n2826) );
  NAND U2983 ( .A(n2826), .B(n8730), .Z(n2619) );
  NAND U2984 ( .A(n2617), .B(n8731), .Z(n2618) );
  NAND U2985 ( .A(n2619), .B(n2618), .Z(n2793) );
  NAND U2986 ( .A(n2620), .B(n8961), .Z(n2622) );
  XOR U2987 ( .A(b[15]), .B(a[18]), .Z(n2760) );
  NAND U2988 ( .A(n2760), .B(n8963), .Z(n2621) );
  NAND U2989 ( .A(n2622), .B(n2621), .Z(n2790) );
  XNOR U2990 ( .A(b[21]), .B(a[12]), .Z(n2751) );
  NANDN U2991 ( .A(n2751), .B(n9493), .Z(n2625) );
  NANDN U2992 ( .A(n2623), .B(n9495), .Z(n2624) );
  AND U2993 ( .A(n2625), .B(n2624), .Z(n2791) );
  XNOR U2994 ( .A(n2790), .B(n2791), .Z(n2792) );
  XNOR U2995 ( .A(n2793), .B(n2792), .Z(n2836) );
  XOR U2996 ( .A(n2835), .B(n2836), .Z(n2838) );
  NANDN U2997 ( .A(n2627), .B(n2626), .Z(n2631) );
  NAND U2998 ( .A(n2629), .B(n2628), .Z(n2630) );
  AND U2999 ( .A(n2631), .B(n2630), .Z(n2837) );
  XOR U3000 ( .A(n2838), .B(n2837), .Z(n2726) );
  XNOR U3001 ( .A(n2725), .B(n2726), .Z(n2741) );
  NANDN U3002 ( .A(n2633), .B(n2632), .Z(n2637) );
  NAND U3003 ( .A(n2635), .B(n2634), .Z(n2636) );
  NAND U3004 ( .A(n2637), .B(n2636), .Z(n2742) );
  XNOR U3005 ( .A(n2741), .B(n2742), .Z(n2743) );
  XOR U3006 ( .A(n2743), .B(n2744), .Z(n2719) );
  NANDN U3007 ( .A(n2643), .B(n2642), .Z(n2647) );
  NAND U3008 ( .A(n2645), .B(n2644), .Z(n2646) );
  NAND U3009 ( .A(n2647), .B(n2646), .Z(n2718) );
  NANDN U3010 ( .A(n2649), .B(n2648), .Z(n2653) );
  OR U3011 ( .A(n2651), .B(n2650), .Z(n2652) );
  NAND U3012 ( .A(n2653), .B(n2652), .Z(n2748) );
  XOR U3013 ( .A(b[11]), .B(a[22]), .Z(n2802) );
  NAND U3014 ( .A(n2802), .B(n8541), .Z(n2656) );
  NAND U3015 ( .A(n2654), .B(n8542), .Z(n2655) );
  NAND U3016 ( .A(n2656), .B(n2655), .Z(n2832) );
  XOR U3017 ( .A(n320), .B(n3831), .Z(n2823) );
  NAND U3018 ( .A(n2823), .B(n9706), .Z(n2659) );
  NANDN U3019 ( .A(n2657), .B(n9707), .Z(n2658) );
  NAND U3020 ( .A(n2659), .B(n2658), .Z(n2829) );
  NANDN U3021 ( .A(n2660), .B(n9801), .Z(n2662) );
  XNOR U3022 ( .A(b[27]), .B(a[6]), .Z(n2817) );
  OR U3023 ( .A(n2817), .B(n9751), .Z(n2661) );
  AND U3024 ( .A(n2662), .B(n2661), .Z(n2830) );
  XNOR U3025 ( .A(n2829), .B(n2830), .Z(n2831) );
  XNOR U3026 ( .A(n2832), .B(n2831), .Z(n2729) );
  XNOR U3027 ( .A(b[7]), .B(n6500), .Z(n2805) );
  NANDN U3028 ( .A(n8013), .B(n2805), .Z(n2665) );
  NAND U3029 ( .A(n2663), .B(n8014), .Z(n2664) );
  NAND U3030 ( .A(n2665), .B(n2664), .Z(n2769) );
  NAND U3031 ( .A(n2666), .B(n9379), .Z(n2668) );
  XNOR U3032 ( .A(n9562), .B(a[14]), .Z(n2754) );
  NAND U3033 ( .A(n2754), .B(n9378), .Z(n2667) );
  NAND U3034 ( .A(n2668), .B(n2667), .Z(n2766) );
  XNOR U3035 ( .A(n317), .B(a[28]), .Z(n2808) );
  NAND U3036 ( .A(n2808), .B(n7905), .Z(n2671) );
  NANDN U3037 ( .A(n2669), .B(n7906), .Z(n2670) );
  AND U3038 ( .A(n2671), .B(n2670), .Z(n2767) );
  XNOR U3039 ( .A(n2766), .B(n2767), .Z(n2768) );
  XOR U3040 ( .A(n2769), .B(n2768), .Z(n2730) );
  XOR U3041 ( .A(n2729), .B(n2730), .Z(n2732) );
  NANDN U3042 ( .A(n2673), .B(n2672), .Z(n2677) );
  NAND U3043 ( .A(n2675), .B(n2674), .Z(n2676) );
  NAND U3044 ( .A(n2677), .B(n2676), .Z(n2731) );
  XOR U3045 ( .A(n2732), .B(n2731), .Z(n2745) );
  NANDN U3046 ( .A(n2679), .B(n2678), .Z(n2683) );
  NAND U3047 ( .A(n2681), .B(n2680), .Z(n2682) );
  NAND U3048 ( .A(n2683), .B(n2682), .Z(n2738) );
  AND U3049 ( .A(n2685), .B(n2684), .Z(n2787) );
  NAND U3050 ( .A(n2686), .B(n7622), .Z(n2688) );
  XNOR U3051 ( .A(n316), .B(a[30]), .Z(n2796) );
  NAND U3052 ( .A(n2796), .B(n7620), .Z(n2687) );
  NAND U3053 ( .A(n2688), .B(n2687), .Z(n2785) );
  XNOR U3054 ( .A(b[17]), .B(a[16]), .Z(n2811) );
  NANDN U3055 ( .A(n2811), .B(n9107), .Z(n2691) );
  NAND U3056 ( .A(n2689), .B(n9105), .Z(n2690) );
  AND U3057 ( .A(n2691), .B(n2690), .Z(n2784) );
  XNOR U3058 ( .A(n2785), .B(n2784), .Z(n2786) );
  XOR U3059 ( .A(n2787), .B(n2786), .Z(n2736) );
  NAND U3060 ( .A(n2692), .B(n8286), .Z(n2694) );
  XOR U3061 ( .A(b[9]), .B(a[24]), .Z(n2799) );
  NAND U3062 ( .A(n2799), .B(n8288), .Z(n2693) );
  NAND U3063 ( .A(n2694), .B(n2693), .Z(n2774) );
  NAND U3064 ( .A(n2695), .B(n9914), .Z(n2697) );
  XNOR U3065 ( .A(n323), .B(a[2]), .Z(n2814) );
  NANDN U3066 ( .A(n9913), .B(n2814), .Z(n2696) );
  NAND U3067 ( .A(n2697), .B(n2696), .Z(n2772) );
  NANDN U3068 ( .A(n2698), .B(n9622), .Z(n2700) );
  XNOR U3069 ( .A(b[23]), .B(a[10]), .Z(n2757) );
  OR U3070 ( .A(n2757), .B(n9621), .Z(n2699) );
  AND U3071 ( .A(n2700), .B(n2699), .Z(n2773) );
  XOR U3072 ( .A(n2772), .B(n2773), .Z(n2775) );
  XNOR U3073 ( .A(n2774), .B(n2775), .Z(n2735) );
  XOR U3074 ( .A(n2736), .B(n2735), .Z(n2737) );
  XNOR U3075 ( .A(n2738), .B(n2737), .Z(n2746) );
  XNOR U3076 ( .A(n2748), .B(n2747), .Z(n2717) );
  XNOR U3077 ( .A(n2718), .B(n2717), .Z(n2720) );
  XNOR U3078 ( .A(n2719), .B(n2720), .Z(n2714) );
  XOR U3079 ( .A(n2713), .B(n2714), .Z(n2841) );
  XNOR U3080 ( .A(n2842), .B(n2841), .Z(n2843) );
  XNOR U3081 ( .A(n2844), .B(n2843), .Z(n2705) );
  XNOR U3082 ( .A(n2705), .B(n2706), .Z(n2707) );
  XOR U3083 ( .A(n2708), .B(n2707), .Z(n2846) );
  XOR U3084 ( .A(n2847), .B(n2846), .Z(c[64]) );
  NANDN U3085 ( .A(n2706), .B(n2705), .Z(n2710) );
  NAND U3086 ( .A(n2708), .B(n2707), .Z(n2709) );
  NAND U3087 ( .A(n2710), .B(n2709), .Z(n2853) );
  NANDN U3088 ( .A(n2712), .B(n2711), .Z(n2716) );
  NAND U3089 ( .A(n2714), .B(n2713), .Z(n2715) );
  NAND U3090 ( .A(n2716), .B(n2715), .Z(n2856) );
  NAND U3091 ( .A(n2718), .B(n2717), .Z(n2722) );
  NANDN U3092 ( .A(n2720), .B(n2719), .Z(n2721) );
  NAND U3093 ( .A(n2722), .B(n2721), .Z(n2871) );
  NANDN U3094 ( .A(n2724), .B(n2723), .Z(n2728) );
  NAND U3095 ( .A(n2726), .B(n2725), .Z(n2727) );
  NAND U3096 ( .A(n2728), .B(n2727), .Z(n2986) );
  NANDN U3097 ( .A(n2730), .B(n2729), .Z(n2734) );
  OR U3098 ( .A(n2732), .B(n2731), .Z(n2733) );
  NAND U3099 ( .A(n2734), .B(n2733), .Z(n2983) );
  NAND U3100 ( .A(n2736), .B(n2735), .Z(n2740) );
  NAND U3101 ( .A(n2738), .B(n2737), .Z(n2739) );
  NAND U3102 ( .A(n2740), .B(n2739), .Z(n2984) );
  XNOR U3103 ( .A(n2983), .B(n2984), .Z(n2985) );
  XOR U3104 ( .A(n2986), .B(n2985), .Z(n2868) );
  XNOR U3105 ( .A(n2868), .B(n2869), .Z(n2870) );
  XNOR U3106 ( .A(n2871), .B(n2870), .Z(n2857) );
  XNOR U3107 ( .A(n2856), .B(n2857), .Z(n2858) );
  OR U3108 ( .A(n2746), .B(n2745), .Z(n2750) );
  NANDN U3109 ( .A(n2748), .B(n2747), .Z(n2749) );
  NAND U3110 ( .A(n2750), .B(n2749), .Z(n2865) );
  XOR U3111 ( .A(n318), .B(n4578), .Z(n2938) );
  NAND U3112 ( .A(n2938), .B(n9493), .Z(n2753) );
  NANDN U3113 ( .A(n2751), .B(n9495), .Z(n2752) );
  NAND U3114 ( .A(n2753), .B(n2752), .Z(n2972) );
  NAND U3115 ( .A(n2754), .B(n9379), .Z(n2756) );
  XNOR U3116 ( .A(n9562), .B(a[15]), .Z(n2911) );
  NAND U3117 ( .A(n2911), .B(n9378), .Z(n2755) );
  NAND U3118 ( .A(n2756), .B(n2755), .Z(n2969) );
  NANDN U3119 ( .A(n2757), .B(n9622), .Z(n2759) );
  XNOR U3120 ( .A(b[23]), .B(a[11]), .Z(n2954) );
  OR U3121 ( .A(n2954), .B(n9621), .Z(n2758) );
  AND U3122 ( .A(n2759), .B(n2758), .Z(n2970) );
  XNOR U3123 ( .A(n2969), .B(n2970), .Z(n2971) );
  XNOR U3124 ( .A(n2972), .B(n2971), .Z(n2874) );
  NAND U3125 ( .A(n2760), .B(n8961), .Z(n2762) );
  XOR U3126 ( .A(b[15]), .B(a[19]), .Z(n2935) );
  NAND U3127 ( .A(n2935), .B(n8963), .Z(n2761) );
  NAND U3128 ( .A(n2762), .B(n2761), .Z(n2898) );
  NAND U3129 ( .A(n9875), .B(n2763), .Z(n2765) );
  XOR U3130 ( .A(b[29]), .B(n3389), .Z(n2951) );
  OR U3131 ( .A(n2951), .B(n9874), .Z(n2764) );
  NAND U3132 ( .A(n2765), .B(n2764), .Z(n2896) );
  NANDN U3133 ( .A(n323), .B(a[1]), .Z(n2897) );
  XNOR U3134 ( .A(n2896), .B(n2897), .Z(n2899) );
  XOR U3135 ( .A(n2898), .B(n2899), .Z(n2875) );
  XNOR U3136 ( .A(n2874), .B(n2875), .Z(n2876) );
  NANDN U3137 ( .A(n2767), .B(n2766), .Z(n2771) );
  NAND U3138 ( .A(n2769), .B(n2768), .Z(n2770) );
  NAND U3139 ( .A(n2771), .B(n2770), .Z(n2877) );
  XOR U3140 ( .A(n2876), .B(n2877), .Z(n2929) );
  NANDN U3141 ( .A(n2773), .B(n2772), .Z(n2777) );
  NANDN U3142 ( .A(n2775), .B(n2774), .Z(n2776) );
  NAND U3143 ( .A(n2777), .B(n2776), .Z(n2926) );
  NANDN U3144 ( .A(n2779), .B(n2778), .Z(n2783) );
  OR U3145 ( .A(n2781), .B(n2780), .Z(n2782) );
  AND U3146 ( .A(n2783), .B(n2782), .Z(n2927) );
  XNOR U3147 ( .A(n2926), .B(n2927), .Z(n2928) );
  XNOR U3148 ( .A(n2929), .B(n2928), .Z(n2980) );
  NANDN U3149 ( .A(n2785), .B(n2784), .Z(n2789) );
  NANDN U3150 ( .A(n2787), .B(n2786), .Z(n2788) );
  NAND U3151 ( .A(n2789), .B(n2788), .Z(n2977) );
  NANDN U3152 ( .A(n2791), .B(n2790), .Z(n2795) );
  NAND U3153 ( .A(n2793), .B(n2792), .Z(n2794) );
  NAND U3154 ( .A(n2795), .B(n2794), .Z(n2923) );
  NAND U3155 ( .A(n2796), .B(n7622), .Z(n2798) );
  XNOR U3156 ( .A(n316), .B(a[31]), .Z(n2908) );
  NAND U3157 ( .A(n2908), .B(n7620), .Z(n2797) );
  NAND U3158 ( .A(n2798), .B(n2797), .Z(n2894) );
  NAND U3159 ( .A(n2799), .B(n8286), .Z(n2801) );
  XOR U3160 ( .A(b[9]), .B(a[25]), .Z(n2932) );
  NAND U3161 ( .A(n2932), .B(n8288), .Z(n2800) );
  NAND U3162 ( .A(n2801), .B(n2800), .Z(n2893) );
  XOR U3163 ( .A(b[11]), .B(n6044), .Z(n2941) );
  NANDN U3164 ( .A(n2941), .B(n8541), .Z(n2804) );
  NAND U3165 ( .A(n8542), .B(n2802), .Z(n2803) );
  NAND U3166 ( .A(n2804), .B(n2803), .Z(n2892) );
  XNOR U3167 ( .A(n2893), .B(n2892), .Z(n2895) );
  XNOR U3168 ( .A(n2894), .B(n2895), .Z(n2883) );
  XOR U3169 ( .A(b[7]), .B(a[27]), .Z(n2957) );
  NANDN U3170 ( .A(n8013), .B(n2957), .Z(n2807) );
  NAND U3171 ( .A(n8014), .B(n2805), .Z(n2806) );
  NAND U3172 ( .A(n2807), .B(n2806), .Z(n2881) );
  XNOR U3173 ( .A(b[5]), .B(a[29]), .Z(n2917) );
  NANDN U3174 ( .A(n2917), .B(n7905), .Z(n2810) );
  NAND U3175 ( .A(n7906), .B(n2808), .Z(n2809) );
  AND U3176 ( .A(n2810), .B(n2809), .Z(n2880) );
  XNOR U3177 ( .A(n2881), .B(n2880), .Z(n2882) );
  XNOR U3178 ( .A(n2883), .B(n2882), .Z(n2975) );
  NANDN U3179 ( .A(n2811), .B(n9105), .Z(n2813) );
  XNOR U3180 ( .A(n9455), .B(a[17]), .Z(n2902) );
  NAND U3181 ( .A(n2902), .B(n9107), .Z(n2812) );
  NAND U3182 ( .A(n2813), .B(n2812), .Z(n2888) );
  NAND U3183 ( .A(n2814), .B(n9914), .Z(n2816) );
  XNOR U3184 ( .A(n323), .B(a[3]), .Z(n2905) );
  NANDN U3185 ( .A(n9913), .B(n2905), .Z(n2815) );
  NAND U3186 ( .A(n2816), .B(n2815), .Z(n2886) );
  NANDN U3187 ( .A(n2817), .B(n9801), .Z(n2819) );
  XNOR U3188 ( .A(b[27]), .B(a[7]), .Z(n2914) );
  OR U3189 ( .A(n2914), .B(n9751), .Z(n2818) );
  AND U3190 ( .A(n2819), .B(n2818), .Z(n2887) );
  XOR U3191 ( .A(n2886), .B(n2887), .Z(n2889) );
  XNOR U3192 ( .A(n2888), .B(n2889), .Z(n2973) );
  NANDN U3193 ( .A(n315), .B(a[33]), .Z(n2820) );
  XNOR U3194 ( .A(b[1]), .B(n2820), .Z(n2822) );
  NANDN U3195 ( .A(b[0]), .B(a[32]), .Z(n2821) );
  AND U3196 ( .A(n2822), .B(n2821), .Z(n2964) );
  XNOR U3197 ( .A(b[25]), .B(a[9]), .Z(n2960) );
  NANDN U3198 ( .A(n2960), .B(n9706), .Z(n2825) );
  NAND U3199 ( .A(n9707), .B(n2823), .Z(n2824) );
  AND U3200 ( .A(n2825), .B(n2824), .Z(n2963) );
  XNOR U3201 ( .A(n2964), .B(n2963), .Z(n2965) );
  XNOR U3202 ( .A(b[13]), .B(a[21]), .Z(n2944) );
  NANDN U3203 ( .A(n2944), .B(n8730), .Z(n2828) );
  NAND U3204 ( .A(n8731), .B(n2826), .Z(n2827) );
  AND U3205 ( .A(n2828), .B(n2827), .Z(n2966) );
  XNOR U3206 ( .A(n2965), .B(n2966), .Z(n2974) );
  XOR U3207 ( .A(n2973), .B(n2974), .Z(n2976) );
  XOR U3208 ( .A(n2975), .B(n2976), .Z(n2921) );
  NANDN U3209 ( .A(n2830), .B(n2829), .Z(n2834) );
  NAND U3210 ( .A(n2832), .B(n2831), .Z(n2833) );
  AND U3211 ( .A(n2834), .B(n2833), .Z(n2920) );
  XOR U3212 ( .A(n2921), .B(n2920), .Z(n2922) );
  XOR U3213 ( .A(n2923), .B(n2922), .Z(n2978) );
  XNOR U3214 ( .A(n2977), .B(n2978), .Z(n2979) );
  XOR U3215 ( .A(n2980), .B(n2979), .Z(n2863) );
  NANDN U3216 ( .A(n2836), .B(n2835), .Z(n2840) );
  OR U3217 ( .A(n2838), .B(n2837), .Z(n2839) );
  AND U3218 ( .A(n2840), .B(n2839), .Z(n2862) );
  XOR U3219 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3220 ( .A(n2865), .B(n2864), .Z(n2859) );
  XOR U3221 ( .A(n2858), .B(n2859), .Z(n2850) );
  XNOR U3222 ( .A(n2850), .B(n2851), .Z(n2852) );
  XNOR U3223 ( .A(n2853), .B(n2852), .Z(n2989) );
  XNOR U3224 ( .A(n2989), .B(sreg[65]), .Z(n2991) );
  NAND U3225 ( .A(n2845), .B(sreg[64]), .Z(n2849) );
  OR U3226 ( .A(n2847), .B(n2846), .Z(n2848) );
  AND U3227 ( .A(n2849), .B(n2848), .Z(n2990) );
  XOR U3228 ( .A(n2991), .B(n2990), .Z(c[65]) );
  NANDN U3229 ( .A(n2851), .B(n2850), .Z(n2855) );
  NAND U3230 ( .A(n2853), .B(n2852), .Z(n2854) );
  NAND U3231 ( .A(n2855), .B(n2854), .Z(n2997) );
  NANDN U3232 ( .A(n2857), .B(n2856), .Z(n2861) );
  NANDN U3233 ( .A(n2859), .B(n2858), .Z(n2860) );
  NAND U3234 ( .A(n2861), .B(n2860), .Z(n2995) );
  OR U3235 ( .A(n2863), .B(n2862), .Z(n2867) );
  NAND U3236 ( .A(n2865), .B(n2864), .Z(n2866) );
  NAND U3237 ( .A(n2867), .B(n2866), .Z(n2999) );
  NANDN U3238 ( .A(n2869), .B(n2868), .Z(n2873) );
  NAND U3239 ( .A(n2871), .B(n2870), .Z(n2872) );
  AND U3240 ( .A(n2873), .B(n2872), .Z(n2998) );
  XNOR U3241 ( .A(n2999), .B(n2998), .Z(n3000) );
  NANDN U3242 ( .A(n2875), .B(n2874), .Z(n2879) );
  NANDN U3243 ( .A(n2877), .B(n2876), .Z(n2878) );
  NAND U3244 ( .A(n2879), .B(n2878), .Z(n3013) );
  NANDN U3245 ( .A(n2881), .B(n2880), .Z(n2885) );
  NANDN U3246 ( .A(n2883), .B(n2882), .Z(n2884) );
  NAND U3247 ( .A(n2885), .B(n2884), .Z(n3118) );
  NANDN U3248 ( .A(n2887), .B(n2886), .Z(n2891) );
  NANDN U3249 ( .A(n2889), .B(n2888), .Z(n2890) );
  NAND U3250 ( .A(n2891), .B(n2890), .Z(n3117) );
  XNOR U3251 ( .A(n3117), .B(n3116), .Z(n3119) );
  XOR U3252 ( .A(n3118), .B(n3119), .Z(n3010) );
  NANDN U3253 ( .A(n2897), .B(n2896), .Z(n2901) );
  NAND U3254 ( .A(n2899), .B(n2898), .Z(n2900) );
  NAND U3255 ( .A(n2901), .B(n2900), .Z(n3112) );
  NAND U3256 ( .A(n2902), .B(n9105), .Z(n2904) );
  XNOR U3257 ( .A(n9455), .B(a[18]), .Z(n3051) );
  NAND U3258 ( .A(n3051), .B(n9107), .Z(n2903) );
  NAND U3259 ( .A(n2904), .B(n2903), .Z(n3028) );
  NAND U3260 ( .A(n2905), .B(n9914), .Z(n2907) );
  XNOR U3261 ( .A(n323), .B(a[4]), .Z(n3054) );
  NANDN U3262 ( .A(n9913), .B(n3054), .Z(n2906) );
  NAND U3263 ( .A(n2907), .B(n2906), .Z(n3026) );
  NAND U3264 ( .A(n2908), .B(n7622), .Z(n2910) );
  XNOR U3265 ( .A(n316), .B(a[32]), .Z(n3057) );
  NAND U3266 ( .A(n3057), .B(n7620), .Z(n2909) );
  NAND U3267 ( .A(n2910), .B(n2909), .Z(n3027) );
  XOR U3268 ( .A(n3026), .B(n3027), .Z(n3029) );
  XNOR U3269 ( .A(n3028), .B(n3029), .Z(n3110) );
  NAND U3270 ( .A(n2911), .B(n9379), .Z(n2913) );
  XNOR U3271 ( .A(n9562), .B(a[16]), .Z(n3042) );
  NAND U3272 ( .A(n3042), .B(n9378), .Z(n2912) );
  NAND U3273 ( .A(n2913), .B(n2912), .Z(n3075) );
  NANDN U3274 ( .A(n2914), .B(n9801), .Z(n2916) );
  XOR U3275 ( .A(b[27]), .B(n3831), .Z(n3045) );
  OR U3276 ( .A(n3045), .B(n9751), .Z(n2915) );
  NAND U3277 ( .A(n2916), .B(n2915), .Z(n3073) );
  XOR U3278 ( .A(b[5]), .B(n6135), .Z(n3048) );
  NANDN U3279 ( .A(n3048), .B(n7905), .Z(n2919) );
  NANDN U3280 ( .A(n2917), .B(n7906), .Z(n2918) );
  AND U3281 ( .A(n2919), .B(n2918), .Z(n3074) );
  XNOR U3282 ( .A(n3073), .B(n3074), .Z(n3076) );
  XOR U3283 ( .A(n3075), .B(n3076), .Z(n3111) );
  XOR U3284 ( .A(n3110), .B(n3111), .Z(n3113) );
  XOR U3285 ( .A(n3112), .B(n3113), .Z(n3011) );
  XOR U3286 ( .A(n3010), .B(n3011), .Z(n3012) );
  XNOR U3287 ( .A(n3013), .B(n3012), .Z(n3129) );
  OR U3288 ( .A(n2921), .B(n2920), .Z(n2925) );
  NAND U3289 ( .A(n2923), .B(n2922), .Z(n2924) );
  AND U3290 ( .A(n2925), .B(n2924), .Z(n3126) );
  NANDN U3291 ( .A(n2927), .B(n2926), .Z(n2931) );
  NAND U3292 ( .A(n2929), .B(n2928), .Z(n2930) );
  NAND U3293 ( .A(n2931), .B(n2930), .Z(n3007) );
  NAND U3294 ( .A(n2932), .B(n8286), .Z(n2934) );
  XNOR U3295 ( .A(b[9]), .B(n6500), .Z(n3079) );
  NAND U3296 ( .A(n3079), .B(n8288), .Z(n2933) );
  NAND U3297 ( .A(n2934), .B(n2933), .Z(n3034) );
  NAND U3298 ( .A(n2935), .B(n8961), .Z(n2937) );
  XOR U3299 ( .A(b[15]), .B(a[20]), .Z(n3082) );
  NAND U3300 ( .A(n3082), .B(n8963), .Z(n2936) );
  NAND U3301 ( .A(n2937), .B(n2936), .Z(n3033) );
  XNOR U3302 ( .A(b[21]), .B(a[14]), .Z(n3085) );
  NANDN U3303 ( .A(n3085), .B(n9493), .Z(n2940) );
  NAND U3304 ( .A(n9495), .B(n2938), .Z(n2939) );
  NAND U3305 ( .A(n2940), .B(n2939), .Z(n3032) );
  XNOR U3306 ( .A(n3033), .B(n3032), .Z(n3035) );
  XNOR U3307 ( .A(n3034), .B(n3035), .Z(n3023) );
  XNOR U3308 ( .A(b[11]), .B(a[24]), .Z(n3088) );
  NANDN U3309 ( .A(n3088), .B(n8541), .Z(n2943) );
  NANDN U3310 ( .A(n2941), .B(n8542), .Z(n2942) );
  NAND U3311 ( .A(n2943), .B(n2942), .Z(n3021) );
  XNOR U3312 ( .A(b[13]), .B(a[22]), .Z(n3091) );
  NANDN U3313 ( .A(n3091), .B(n8730), .Z(n2946) );
  NANDN U3314 ( .A(n2944), .B(n8731), .Z(n2945) );
  AND U3315 ( .A(n2946), .B(n2945), .Z(n3020) );
  XNOR U3316 ( .A(n3021), .B(n3020), .Z(n3022) );
  XNOR U3317 ( .A(n3023), .B(n3022), .Z(n3017) );
  NANDN U3318 ( .A(n315), .B(a[34]), .Z(n2947) );
  XNOR U3319 ( .A(b[1]), .B(n2947), .Z(n2949) );
  IV U3320 ( .A(a[33]), .Z(n6914) );
  NANDN U3321 ( .A(n6914), .B(n315), .Z(n2948) );
  AND U3322 ( .A(n2949), .B(n2948), .Z(n3039) );
  ANDN U3323 ( .B(b[31]), .A(n2950), .Z(n3036) );
  NANDN U3324 ( .A(n2951), .B(n9875), .Z(n2953) );
  XNOR U3325 ( .A(b[29]), .B(a[6]), .Z(n3095) );
  OR U3326 ( .A(n3095), .B(n9874), .Z(n2952) );
  NAND U3327 ( .A(n2953), .B(n2952), .Z(n3037) );
  XOR U3328 ( .A(n3036), .B(n3037), .Z(n3038) );
  XOR U3329 ( .A(n3039), .B(n3038), .Z(n3014) );
  NANDN U3330 ( .A(n2954), .B(n9622), .Z(n2956) );
  XNOR U3331 ( .A(b[23]), .B(a[12]), .Z(n3101) );
  OR U3332 ( .A(n3101), .B(n9621), .Z(n2955) );
  NAND U3333 ( .A(n2956), .B(n2955), .Z(n3070) );
  XOR U3334 ( .A(b[7]), .B(a[28]), .Z(n3104) );
  NANDN U3335 ( .A(n8013), .B(n3104), .Z(n2959) );
  NAND U3336 ( .A(n2957), .B(n8014), .Z(n2958) );
  NAND U3337 ( .A(n2959), .B(n2958), .Z(n3067) );
  XNOR U3338 ( .A(b[25]), .B(a[10]), .Z(n3107) );
  NANDN U3339 ( .A(n3107), .B(n9706), .Z(n2962) );
  NANDN U3340 ( .A(n2960), .B(n9707), .Z(n2961) );
  AND U3341 ( .A(n2962), .B(n2961), .Z(n3068) );
  XNOR U3342 ( .A(n3067), .B(n3068), .Z(n3069) );
  XNOR U3343 ( .A(n3070), .B(n3069), .Z(n3015) );
  XNOR U3344 ( .A(n3014), .B(n3015), .Z(n3016) );
  XNOR U3345 ( .A(n3017), .B(n3016), .Z(n3064) );
  NANDN U3346 ( .A(n2964), .B(n2963), .Z(n2968) );
  NAND U3347 ( .A(n2966), .B(n2965), .Z(n2967) );
  NAND U3348 ( .A(n2968), .B(n2967), .Z(n3061) );
  XNOR U3349 ( .A(n3061), .B(n3062), .Z(n3063) );
  XNOR U3350 ( .A(n3064), .B(n3063), .Z(n3004) );
  XOR U3351 ( .A(n3004), .B(n3005), .Z(n3006) );
  XNOR U3352 ( .A(n3007), .B(n3006), .Z(n3127) );
  XOR U3353 ( .A(n3129), .B(n3128), .Z(n3123) );
  NANDN U3354 ( .A(n2978), .B(n2977), .Z(n2982) );
  NAND U3355 ( .A(n2980), .B(n2979), .Z(n2981) );
  NAND U3356 ( .A(n2982), .B(n2981), .Z(n3120) );
  NANDN U3357 ( .A(n2984), .B(n2983), .Z(n2988) );
  NANDN U3358 ( .A(n2986), .B(n2985), .Z(n2987) );
  AND U3359 ( .A(n2988), .B(n2987), .Z(n3121) );
  XNOR U3360 ( .A(n3120), .B(n3121), .Z(n3122) );
  XOR U3361 ( .A(n3123), .B(n3122), .Z(n3001) );
  XNOR U3362 ( .A(n3000), .B(n3001), .Z(n2994) );
  XNOR U3363 ( .A(n2995), .B(n2994), .Z(n2996) );
  XNOR U3364 ( .A(n2997), .B(n2996), .Z(n3132) );
  XNOR U3365 ( .A(n3132), .B(sreg[66]), .Z(n3134) );
  NAND U3366 ( .A(n2989), .B(sreg[65]), .Z(n2993) );
  OR U3367 ( .A(n2991), .B(n2990), .Z(n2992) );
  AND U3368 ( .A(n2993), .B(n2992), .Z(n3133) );
  XOR U3369 ( .A(n3134), .B(n3133), .Z(c[66]) );
  NANDN U3370 ( .A(n2999), .B(n2998), .Z(n3003) );
  NANDN U3371 ( .A(n3001), .B(n3000), .Z(n3002) );
  NAND U3372 ( .A(n3003), .B(n3002), .Z(n3137) );
  OR U3373 ( .A(n3005), .B(n3004), .Z(n3009) );
  NAND U3374 ( .A(n3007), .B(n3006), .Z(n3008) );
  NAND U3375 ( .A(n3009), .B(n3008), .Z(n3264) );
  XNOR U3376 ( .A(n3264), .B(n3265), .Z(n3266) );
  NANDN U3377 ( .A(n3015), .B(n3014), .Z(n3019) );
  NANDN U3378 ( .A(n3017), .B(n3016), .Z(n3018) );
  NAND U3379 ( .A(n3019), .B(n3018), .Z(n3151) );
  NANDN U3380 ( .A(n3021), .B(n3020), .Z(n3025) );
  NANDN U3381 ( .A(n3023), .B(n3022), .Z(n3024) );
  NAND U3382 ( .A(n3025), .B(n3024), .Z(n3208) );
  NAND U3383 ( .A(n3027), .B(n3026), .Z(n3031) );
  NAND U3384 ( .A(n3029), .B(n3028), .Z(n3030) );
  NAND U3385 ( .A(n3031), .B(n3030), .Z(n3207) );
  XNOR U3386 ( .A(n3207), .B(n3206), .Z(n3209) );
  XNOR U3387 ( .A(n3208), .B(n3209), .Z(n3149) );
  OR U3388 ( .A(n3037), .B(n3036), .Z(n3041) );
  NANDN U3389 ( .A(n3039), .B(n3038), .Z(n3040) );
  NAND U3390 ( .A(n3041), .B(n3040), .Z(n3219) );
  NAND U3391 ( .A(n3042), .B(n9379), .Z(n3044) );
  XNOR U3392 ( .A(n9562), .B(a[17]), .Z(n3188) );
  NAND U3393 ( .A(n3188), .B(n9378), .Z(n3043) );
  NAND U3394 ( .A(n3044), .B(n3043), .Z(n3230) );
  NANDN U3395 ( .A(n3045), .B(n9801), .Z(n3047) );
  XNOR U3396 ( .A(b[27]), .B(a[9]), .Z(n3191) );
  OR U3397 ( .A(n3191), .B(n9751), .Z(n3046) );
  NAND U3398 ( .A(n3047), .B(n3046), .Z(n3228) );
  XNOR U3399 ( .A(b[5]), .B(a[31]), .Z(n3194) );
  NANDN U3400 ( .A(n3194), .B(n7905), .Z(n3050) );
  NANDN U3401 ( .A(n3048), .B(n7906), .Z(n3049) );
  AND U3402 ( .A(n3050), .B(n3049), .Z(n3229) );
  XNOR U3403 ( .A(n3228), .B(n3229), .Z(n3231) );
  XOR U3404 ( .A(n3230), .B(n3231), .Z(n3216) );
  NAND U3405 ( .A(n3051), .B(n9105), .Z(n3053) );
  XNOR U3406 ( .A(n9455), .B(a[19]), .Z(n3197) );
  NAND U3407 ( .A(n3197), .B(n9107), .Z(n3052) );
  AND U3408 ( .A(n3053), .B(n3052), .Z(n3173) );
  NAND U3409 ( .A(n3054), .B(n9914), .Z(n3056) );
  XNOR U3410 ( .A(n323), .B(a[5]), .Z(n3200) );
  NANDN U3411 ( .A(n9913), .B(n3200), .Z(n3055) );
  AND U3412 ( .A(n3056), .B(n3055), .Z(n3171) );
  NAND U3413 ( .A(n3057), .B(n7622), .Z(n3059) );
  XNOR U3414 ( .A(n316), .B(a[33]), .Z(n3203) );
  NAND U3415 ( .A(n3203), .B(n7620), .Z(n3058) );
  NAND U3416 ( .A(n3059), .B(n3058), .Z(n3170) );
  XOR U3417 ( .A(n3216), .B(n3217), .Z(n3218) );
  XNOR U3418 ( .A(n3219), .B(n3218), .Z(n3150) );
  XNOR U3419 ( .A(n3149), .B(n3150), .Z(n3060) );
  XOR U3420 ( .A(n3151), .B(n3060), .Z(n3272) );
  NANDN U3421 ( .A(n3062), .B(n3061), .Z(n3066) );
  NANDN U3422 ( .A(n3064), .B(n3063), .Z(n3065) );
  NAND U3423 ( .A(n3066), .B(n3065), .Z(n3155) );
  NANDN U3424 ( .A(n3068), .B(n3067), .Z(n3072) );
  NAND U3425 ( .A(n3070), .B(n3069), .Z(n3071) );
  NAND U3426 ( .A(n3072), .B(n3071), .Z(n3210) );
  NANDN U3427 ( .A(n3074), .B(n3073), .Z(n3078) );
  NAND U3428 ( .A(n3076), .B(n3075), .Z(n3077) );
  AND U3429 ( .A(n3078), .B(n3077), .Z(n3211) );
  XNOR U3430 ( .A(n3210), .B(n3211), .Z(n3212) );
  NAND U3431 ( .A(n3079), .B(n8286), .Z(n3081) );
  XOR U3432 ( .A(b[9]), .B(a[27]), .Z(n3234) );
  NAND U3433 ( .A(n3234), .B(n8288), .Z(n3080) );
  NAND U3434 ( .A(n3081), .B(n3080), .Z(n3178) );
  NAND U3435 ( .A(n3082), .B(n8961), .Z(n3084) );
  XOR U3436 ( .A(b[15]), .B(a[21]), .Z(n3237) );
  NAND U3437 ( .A(n3237), .B(n8963), .Z(n3083) );
  NAND U3438 ( .A(n3084), .B(n3083), .Z(n3176) );
  XNOR U3439 ( .A(b[21]), .B(a[15]), .Z(n3240) );
  NANDN U3440 ( .A(n3240), .B(n9493), .Z(n3087) );
  NANDN U3441 ( .A(n3085), .B(n9495), .Z(n3086) );
  AND U3442 ( .A(n3087), .B(n3086), .Z(n3177) );
  XOR U3443 ( .A(n3176), .B(n3177), .Z(n3179) );
  XNOR U3444 ( .A(n3178), .B(n3179), .Z(n3167) );
  XNOR U3445 ( .A(b[11]), .B(a[25]), .Z(n3243) );
  NANDN U3446 ( .A(n3243), .B(n8541), .Z(n3090) );
  NANDN U3447 ( .A(n3088), .B(n8542), .Z(n3089) );
  NAND U3448 ( .A(n3090), .B(n3089), .Z(n3165) );
  XOR U3449 ( .A(b[13]), .B(n6044), .Z(n3246) );
  NANDN U3450 ( .A(n3246), .B(n8730), .Z(n3093) );
  NANDN U3451 ( .A(n3091), .B(n8731), .Z(n3092) );
  NAND U3452 ( .A(n3093), .B(n3092), .Z(n3164) );
  XNOR U3453 ( .A(n3167), .B(n3166), .Z(n3161) );
  ANDN U3454 ( .B(b[31]), .A(n3094), .Z(n3182) );
  NANDN U3455 ( .A(n3095), .B(n9875), .Z(n3097) );
  XNOR U3456 ( .A(n322), .B(a[7]), .Z(n3252) );
  NANDN U3457 ( .A(n9874), .B(n3252), .Z(n3096) );
  NAND U3458 ( .A(n3097), .B(n3096), .Z(n3183) );
  XOR U3459 ( .A(n3182), .B(n3183), .Z(n3184) );
  NANDN U3460 ( .A(n315), .B(a[35]), .Z(n3098) );
  XNOR U3461 ( .A(b[1]), .B(n3098), .Z(n3100) );
  NANDN U3462 ( .A(b[0]), .B(a[34]), .Z(n3099) );
  AND U3463 ( .A(n3100), .B(n3099), .Z(n3185) );
  XNOR U3464 ( .A(n3184), .B(n3185), .Z(n3158) );
  NANDN U3465 ( .A(n3101), .B(n9622), .Z(n3103) );
  XOR U3466 ( .A(b[23]), .B(n4578), .Z(n3255) );
  OR U3467 ( .A(n3255), .B(n9621), .Z(n3102) );
  NAND U3468 ( .A(n3103), .B(n3102), .Z(n3225) );
  XOR U3469 ( .A(b[7]), .B(a[29]), .Z(n3258) );
  NANDN U3470 ( .A(n8013), .B(n3258), .Z(n3106) );
  NAND U3471 ( .A(n3104), .B(n8014), .Z(n3105) );
  NAND U3472 ( .A(n3106), .B(n3105), .Z(n3222) );
  XNOR U3473 ( .A(b[25]), .B(a[11]), .Z(n3261) );
  NANDN U3474 ( .A(n3261), .B(n9706), .Z(n3109) );
  NANDN U3475 ( .A(n3107), .B(n9707), .Z(n3108) );
  AND U3476 ( .A(n3109), .B(n3108), .Z(n3223) );
  XNOR U3477 ( .A(n3222), .B(n3223), .Z(n3224) );
  XNOR U3478 ( .A(n3225), .B(n3224), .Z(n3159) );
  XOR U3479 ( .A(n3161), .B(n3160), .Z(n3213) );
  XOR U3480 ( .A(n3212), .B(n3213), .Z(n3152) );
  NANDN U3481 ( .A(n3111), .B(n3110), .Z(n3115) );
  OR U3482 ( .A(n3113), .B(n3112), .Z(n3114) );
  AND U3483 ( .A(n3115), .B(n3114), .Z(n3153) );
  XNOR U3484 ( .A(n3152), .B(n3153), .Z(n3154) );
  XOR U3485 ( .A(n3155), .B(n3154), .Z(n3270) );
  XNOR U3486 ( .A(n3270), .B(n3271), .Z(n3273) );
  XNOR U3487 ( .A(n3272), .B(n3273), .Z(n3267) );
  XOR U3488 ( .A(n3266), .B(n3267), .Z(n3146) );
  NANDN U3489 ( .A(n3121), .B(n3120), .Z(n3125) );
  NANDN U3490 ( .A(n3123), .B(n3122), .Z(n3124) );
  NAND U3491 ( .A(n3125), .B(n3124), .Z(n3143) );
  OR U3492 ( .A(n3127), .B(n3126), .Z(n3131) );
  NAND U3493 ( .A(n3129), .B(n3128), .Z(n3130) );
  NAND U3494 ( .A(n3131), .B(n3130), .Z(n3144) );
  XNOR U3495 ( .A(n3143), .B(n3144), .Z(n3145) );
  XNOR U3496 ( .A(n3146), .B(n3145), .Z(n3138) );
  XNOR U3497 ( .A(n3137), .B(n3138), .Z(n3139) );
  XNOR U3498 ( .A(n3140), .B(n3139), .Z(n3276) );
  XNOR U3499 ( .A(n3276), .B(sreg[67]), .Z(n3278) );
  NAND U3500 ( .A(n3132), .B(sreg[66]), .Z(n3136) );
  OR U3501 ( .A(n3134), .B(n3133), .Z(n3135) );
  AND U3502 ( .A(n3136), .B(n3135), .Z(n3277) );
  XOR U3503 ( .A(n3278), .B(n3277), .Z(c[67]) );
  NANDN U3504 ( .A(n3138), .B(n3137), .Z(n3142) );
  NAND U3505 ( .A(n3140), .B(n3139), .Z(n3141) );
  NAND U3506 ( .A(n3142), .B(n3141), .Z(n3284) );
  NANDN U3507 ( .A(n3144), .B(n3143), .Z(n3148) );
  NAND U3508 ( .A(n3146), .B(n3145), .Z(n3147) );
  NAND U3509 ( .A(n3148), .B(n3147), .Z(n3281) );
  NANDN U3510 ( .A(n3153), .B(n3152), .Z(n3157) );
  NAND U3511 ( .A(n3155), .B(n3154), .Z(n3156) );
  NAND U3512 ( .A(n3157), .B(n3156), .Z(n3413) );
  XOR U3513 ( .A(n3412), .B(n3413), .Z(n3415) );
  OR U3514 ( .A(n3159), .B(n3158), .Z(n3163) );
  NANDN U3515 ( .A(n3161), .B(n3160), .Z(n3162) );
  NAND U3516 ( .A(n3163), .B(n3162), .Z(n3405) );
  OR U3517 ( .A(n3165), .B(n3164), .Z(n3169) );
  NANDN U3518 ( .A(n3167), .B(n3166), .Z(n3168) );
  NAND U3519 ( .A(n3169), .B(n3168), .Z(n3343) );
  NANDN U3520 ( .A(n3171), .B(n3170), .Z(n3175) );
  NANDN U3521 ( .A(n3173), .B(n3172), .Z(n3174) );
  NAND U3522 ( .A(n3175), .B(n3174), .Z(n3342) );
  NANDN U3523 ( .A(n3177), .B(n3176), .Z(n3181) );
  NANDN U3524 ( .A(n3179), .B(n3178), .Z(n3180) );
  NAND U3525 ( .A(n3181), .B(n3180), .Z(n3341) );
  XOR U3526 ( .A(n3343), .B(n3344), .Z(n3403) );
  OR U3527 ( .A(n3183), .B(n3182), .Z(n3187) );
  NANDN U3528 ( .A(n3185), .B(n3184), .Z(n3186) );
  NAND U3529 ( .A(n3187), .B(n3186), .Z(n3356) );
  NAND U3530 ( .A(n3188), .B(n9379), .Z(n3190) );
  XNOR U3531 ( .A(n9562), .B(a[18]), .Z(n3299) );
  NAND U3532 ( .A(n3299), .B(n9378), .Z(n3189) );
  NAND U3533 ( .A(n3190), .B(n3189), .Z(n3367) );
  NANDN U3534 ( .A(n3191), .B(n9801), .Z(n3193) );
  XNOR U3535 ( .A(b[27]), .B(a[10]), .Z(n3302) );
  OR U3536 ( .A(n3302), .B(n9751), .Z(n3192) );
  NAND U3537 ( .A(n3193), .B(n3192), .Z(n3365) );
  XNOR U3538 ( .A(b[5]), .B(a[32]), .Z(n3305) );
  NANDN U3539 ( .A(n3305), .B(n7905), .Z(n3196) );
  NANDN U3540 ( .A(n3194), .B(n7906), .Z(n3195) );
  AND U3541 ( .A(n3196), .B(n3195), .Z(n3366) );
  XNOR U3542 ( .A(n3365), .B(n3366), .Z(n3368) );
  XOR U3543 ( .A(n3367), .B(n3368), .Z(n3353) );
  NAND U3544 ( .A(n3197), .B(n9105), .Z(n3199) );
  XNOR U3545 ( .A(n9455), .B(a[20]), .Z(n3308) );
  NAND U3546 ( .A(n3308), .B(n9107), .Z(n3198) );
  NAND U3547 ( .A(n3199), .B(n3198), .Z(n3325) );
  NAND U3548 ( .A(n3200), .B(n9914), .Z(n3202) );
  XNOR U3549 ( .A(n323), .B(a[6]), .Z(n3311) );
  NANDN U3550 ( .A(n9913), .B(n3311), .Z(n3201) );
  NAND U3551 ( .A(n3202), .B(n3201), .Z(n3323) );
  NAND U3552 ( .A(n3203), .B(n7622), .Z(n3205) );
  XNOR U3553 ( .A(n316), .B(a[34]), .Z(n3314) );
  NAND U3554 ( .A(n3314), .B(n7620), .Z(n3204) );
  NAND U3555 ( .A(n3205), .B(n3204), .Z(n3324) );
  XOR U3556 ( .A(n3323), .B(n3324), .Z(n3326) );
  XOR U3557 ( .A(n3325), .B(n3326), .Z(n3354) );
  XOR U3558 ( .A(n3353), .B(n3354), .Z(n3355) );
  XNOR U3559 ( .A(n3356), .B(n3355), .Z(n3402) );
  XOR U3560 ( .A(n3403), .B(n3402), .Z(n3404) );
  XNOR U3561 ( .A(n3405), .B(n3404), .Z(n3421) );
  NANDN U3562 ( .A(n3211), .B(n3210), .Z(n3215) );
  NANDN U3563 ( .A(n3213), .B(n3212), .Z(n3214) );
  NAND U3564 ( .A(n3215), .B(n3214), .Z(n3408) );
  NAND U3565 ( .A(n3217), .B(n3216), .Z(n3221) );
  NANDN U3566 ( .A(n3219), .B(n3218), .Z(n3220) );
  NAND U3567 ( .A(n3221), .B(n3220), .Z(n3407) );
  NANDN U3568 ( .A(n3223), .B(n3222), .Z(n3227) );
  NAND U3569 ( .A(n3225), .B(n3224), .Z(n3226) );
  NAND U3570 ( .A(n3227), .B(n3226), .Z(n3347) );
  NANDN U3571 ( .A(n3229), .B(n3228), .Z(n3233) );
  NAND U3572 ( .A(n3231), .B(n3230), .Z(n3232) );
  AND U3573 ( .A(n3233), .B(n3232), .Z(n3348) );
  XNOR U3574 ( .A(n3347), .B(n3348), .Z(n3349) );
  NAND U3575 ( .A(n3234), .B(n8286), .Z(n3236) );
  XOR U3576 ( .A(b[9]), .B(a[28]), .Z(n3371) );
  NAND U3577 ( .A(n3371), .B(n8288), .Z(n3235) );
  NAND U3578 ( .A(n3236), .B(n3235), .Z(n3331) );
  NAND U3579 ( .A(n3237), .B(n8961), .Z(n3239) );
  XOR U3580 ( .A(b[15]), .B(a[22]), .Z(n3374) );
  NAND U3581 ( .A(n3374), .B(n8963), .Z(n3238) );
  NAND U3582 ( .A(n3239), .B(n3238), .Z(n3329) );
  XNOR U3583 ( .A(b[21]), .B(a[16]), .Z(n3377) );
  NANDN U3584 ( .A(n3377), .B(n9493), .Z(n3242) );
  NANDN U3585 ( .A(n3240), .B(n9495), .Z(n3241) );
  AND U3586 ( .A(n3242), .B(n3241), .Z(n3330) );
  XOR U3587 ( .A(n3329), .B(n3330), .Z(n3332) );
  XNOR U3588 ( .A(n3331), .B(n3332), .Z(n3320) );
  XOR U3589 ( .A(b[11]), .B(n6500), .Z(n3380) );
  NANDN U3590 ( .A(n3380), .B(n8541), .Z(n3245) );
  NANDN U3591 ( .A(n3243), .B(n8542), .Z(n3244) );
  NAND U3592 ( .A(n3245), .B(n3244), .Z(n3318) );
  XNOR U3593 ( .A(b[13]), .B(a[24]), .Z(n3383) );
  NANDN U3594 ( .A(n3383), .B(n8730), .Z(n3248) );
  NANDN U3595 ( .A(n3246), .B(n8731), .Z(n3247) );
  AND U3596 ( .A(n3248), .B(n3247), .Z(n3317) );
  XNOR U3597 ( .A(n3318), .B(n3317), .Z(n3319) );
  XNOR U3598 ( .A(n3320), .B(n3319), .Z(n3337) );
  NANDN U3599 ( .A(n315), .B(a[36]), .Z(n3249) );
  XNOR U3600 ( .A(b[1]), .B(n3249), .Z(n3251) );
  NANDN U3601 ( .A(b[0]), .B(a[35]), .Z(n3250) );
  AND U3602 ( .A(n3251), .B(n3250), .Z(n3295) );
  NAND U3603 ( .A(n3252), .B(n9875), .Z(n3254) );
  XOR U3604 ( .A(b[29]), .B(n3831), .Z(n3390) );
  OR U3605 ( .A(n3390), .B(n9874), .Z(n3253) );
  NAND U3606 ( .A(n3254), .B(n3253), .Z(n3293) );
  NANDN U3607 ( .A(n323), .B(a[4]), .Z(n3294) );
  XNOR U3608 ( .A(n3293), .B(n3294), .Z(n3296) );
  XOR U3609 ( .A(n3295), .B(n3296), .Z(n3335) );
  NANDN U3610 ( .A(n3255), .B(n9622), .Z(n3257) );
  XNOR U3611 ( .A(b[23]), .B(a[14]), .Z(n3393) );
  OR U3612 ( .A(n3393), .B(n9621), .Z(n3256) );
  NAND U3613 ( .A(n3257), .B(n3256), .Z(n3362) );
  XNOR U3614 ( .A(b[7]), .B(a[30]), .Z(n3396) );
  OR U3615 ( .A(n3396), .B(n8013), .Z(n3260) );
  NAND U3616 ( .A(n3258), .B(n8014), .Z(n3259) );
  NAND U3617 ( .A(n3260), .B(n3259), .Z(n3359) );
  XNOR U3618 ( .A(b[25]), .B(a[12]), .Z(n3399) );
  NANDN U3619 ( .A(n3399), .B(n9706), .Z(n3263) );
  NANDN U3620 ( .A(n3261), .B(n9707), .Z(n3262) );
  AND U3621 ( .A(n3263), .B(n3262), .Z(n3360) );
  XNOR U3622 ( .A(n3359), .B(n3360), .Z(n3361) );
  XNOR U3623 ( .A(n3362), .B(n3361), .Z(n3336) );
  XOR U3624 ( .A(n3335), .B(n3336), .Z(n3338) );
  XNOR U3625 ( .A(n3337), .B(n3338), .Z(n3350) );
  XNOR U3626 ( .A(n3349), .B(n3350), .Z(n3406) );
  XNOR U3627 ( .A(n3407), .B(n3406), .Z(n3409) );
  XNOR U3628 ( .A(n3408), .B(n3409), .Z(n3418) );
  XNOR U3629 ( .A(n3419), .B(n3418), .Z(n3420) );
  XOR U3630 ( .A(n3421), .B(n3420), .Z(n3414) );
  XNOR U3631 ( .A(n3415), .B(n3414), .Z(n3290) );
  NANDN U3632 ( .A(n3265), .B(n3264), .Z(n3269) );
  NANDN U3633 ( .A(n3267), .B(n3266), .Z(n3268) );
  NAND U3634 ( .A(n3269), .B(n3268), .Z(n3288) );
  OR U3635 ( .A(n3271), .B(n3270), .Z(n3275) );
  OR U3636 ( .A(n3273), .B(n3272), .Z(n3274) );
  AND U3637 ( .A(n3275), .B(n3274), .Z(n3287) );
  XNOR U3638 ( .A(n3288), .B(n3287), .Z(n3289) );
  XNOR U3639 ( .A(n3290), .B(n3289), .Z(n3282) );
  XNOR U3640 ( .A(n3281), .B(n3282), .Z(n3283) );
  XNOR U3641 ( .A(n3284), .B(n3283), .Z(n3424) );
  XNOR U3642 ( .A(n3424), .B(sreg[68]), .Z(n3426) );
  NAND U3643 ( .A(n3276), .B(sreg[67]), .Z(n3280) );
  OR U3644 ( .A(n3278), .B(n3277), .Z(n3279) );
  AND U3645 ( .A(n3280), .B(n3279), .Z(n3425) );
  XOR U3646 ( .A(n3426), .B(n3425), .Z(c[68]) );
  NANDN U3647 ( .A(n3282), .B(n3281), .Z(n3286) );
  NAND U3648 ( .A(n3284), .B(n3283), .Z(n3285) );
  NAND U3649 ( .A(n3286), .B(n3285), .Z(n3432) );
  NANDN U3650 ( .A(n3288), .B(n3287), .Z(n3292) );
  NAND U3651 ( .A(n3290), .B(n3289), .Z(n3291) );
  NAND U3652 ( .A(n3292), .B(n3291), .Z(n3430) );
  NANDN U3653 ( .A(n3294), .B(n3293), .Z(n3298) );
  NAND U3654 ( .A(n3296), .B(n3295), .Z(n3297) );
  NAND U3655 ( .A(n3298), .B(n3297), .Z(n3504) );
  NAND U3656 ( .A(n3299), .B(n9379), .Z(n3301) );
  XNOR U3657 ( .A(n9562), .B(a[19]), .Z(n3471) );
  NAND U3658 ( .A(n3471), .B(n9378), .Z(n3300) );
  NAND U3659 ( .A(n3301), .B(n3300), .Z(n3515) );
  NANDN U3660 ( .A(n3302), .B(n9801), .Z(n3304) );
  XNOR U3661 ( .A(b[27]), .B(a[11]), .Z(n3474) );
  OR U3662 ( .A(n3474), .B(n9751), .Z(n3303) );
  NAND U3663 ( .A(n3304), .B(n3303), .Z(n3513) );
  XOR U3664 ( .A(b[5]), .B(n6914), .Z(n3477) );
  NANDN U3665 ( .A(n3477), .B(n7905), .Z(n3307) );
  NANDN U3666 ( .A(n3305), .B(n7906), .Z(n3306) );
  AND U3667 ( .A(n3307), .B(n3306), .Z(n3514) );
  XNOR U3668 ( .A(n3513), .B(n3514), .Z(n3516) );
  XOR U3669 ( .A(n3515), .B(n3516), .Z(n3501) );
  NAND U3670 ( .A(n3308), .B(n9105), .Z(n3310) );
  XNOR U3671 ( .A(n9455), .B(a[21]), .Z(n3480) );
  NAND U3672 ( .A(n3480), .B(n9107), .Z(n3309) );
  AND U3673 ( .A(n3310), .B(n3309), .Z(n3456) );
  NAND U3674 ( .A(n3311), .B(n9914), .Z(n3313) );
  XNOR U3675 ( .A(n323), .B(a[7]), .Z(n3483) );
  NANDN U3676 ( .A(n9913), .B(n3483), .Z(n3312) );
  AND U3677 ( .A(n3313), .B(n3312), .Z(n3454) );
  NAND U3678 ( .A(n3314), .B(n7622), .Z(n3316) );
  XNOR U3679 ( .A(n316), .B(a[35]), .Z(n3486) );
  NAND U3680 ( .A(n3486), .B(n7620), .Z(n3315) );
  NAND U3681 ( .A(n3316), .B(n3315), .Z(n3453) );
  XOR U3682 ( .A(n3501), .B(n3502), .Z(n3503) );
  XNOR U3683 ( .A(n3504), .B(n3503), .Z(n3549) );
  NANDN U3684 ( .A(n3318), .B(n3317), .Z(n3322) );
  NANDN U3685 ( .A(n3320), .B(n3319), .Z(n3321) );
  NAND U3686 ( .A(n3322), .B(n3321), .Z(n3492) );
  NAND U3687 ( .A(n3324), .B(n3323), .Z(n3328) );
  NAND U3688 ( .A(n3326), .B(n3325), .Z(n3327) );
  NAND U3689 ( .A(n3328), .B(n3327), .Z(n3490) );
  NANDN U3690 ( .A(n3330), .B(n3329), .Z(n3334) );
  NANDN U3691 ( .A(n3332), .B(n3331), .Z(n3333) );
  NAND U3692 ( .A(n3334), .B(n3333), .Z(n3489) );
  XNOR U3693 ( .A(n3492), .B(n3491), .Z(n3550) );
  XOR U3694 ( .A(n3549), .B(n3550), .Z(n3552) );
  NANDN U3695 ( .A(n3336), .B(n3335), .Z(n3340) );
  OR U3696 ( .A(n3338), .B(n3337), .Z(n3339) );
  NAND U3697 ( .A(n3340), .B(n3339), .Z(n3551) );
  XOR U3698 ( .A(n3552), .B(n3551), .Z(n3569) );
  OR U3699 ( .A(n3342), .B(n3341), .Z(n3346) );
  NANDN U3700 ( .A(n3344), .B(n3343), .Z(n3345) );
  NAND U3701 ( .A(n3346), .B(n3345), .Z(n3568) );
  NANDN U3702 ( .A(n3348), .B(n3347), .Z(n3352) );
  NANDN U3703 ( .A(n3350), .B(n3349), .Z(n3351) );
  NAND U3704 ( .A(n3352), .B(n3351), .Z(n3557) );
  NAND U3705 ( .A(n3354), .B(n3353), .Z(n3358) );
  NANDN U3706 ( .A(n3356), .B(n3355), .Z(n3357) );
  NAND U3707 ( .A(n3358), .B(n3357), .Z(n3556) );
  NANDN U3708 ( .A(n3360), .B(n3359), .Z(n3364) );
  NAND U3709 ( .A(n3362), .B(n3361), .Z(n3363) );
  NAND U3710 ( .A(n3364), .B(n3363), .Z(n3495) );
  NANDN U3711 ( .A(n3366), .B(n3365), .Z(n3370) );
  NAND U3712 ( .A(n3368), .B(n3367), .Z(n3369) );
  AND U3713 ( .A(n3370), .B(n3369), .Z(n3496) );
  XNOR U3714 ( .A(n3495), .B(n3496), .Z(n3497) );
  NAND U3715 ( .A(n3371), .B(n8286), .Z(n3373) );
  XOR U3716 ( .A(b[9]), .B(a[29]), .Z(n3519) );
  NAND U3717 ( .A(n3519), .B(n8288), .Z(n3372) );
  NAND U3718 ( .A(n3373), .B(n3372), .Z(n3461) );
  NAND U3719 ( .A(n3374), .B(n8961), .Z(n3376) );
  XNOR U3720 ( .A(b[15]), .B(n6044), .Z(n3522) );
  NAND U3721 ( .A(n3522), .B(n8963), .Z(n3375) );
  NAND U3722 ( .A(n3376), .B(n3375), .Z(n3459) );
  XOR U3723 ( .A(b[21]), .B(n5168), .Z(n3525) );
  NANDN U3724 ( .A(n3525), .B(n9493), .Z(n3379) );
  NANDN U3725 ( .A(n3377), .B(n9495), .Z(n3378) );
  AND U3726 ( .A(n3379), .B(n3378), .Z(n3460) );
  XOR U3727 ( .A(n3459), .B(n3460), .Z(n3462) );
  XNOR U3728 ( .A(n3461), .B(n3462), .Z(n3450) );
  XNOR U3729 ( .A(b[11]), .B(a[27]), .Z(n3528) );
  NANDN U3730 ( .A(n3528), .B(n8541), .Z(n3382) );
  NANDN U3731 ( .A(n3380), .B(n8542), .Z(n3381) );
  NAND U3732 ( .A(n3382), .B(n3381), .Z(n3448) );
  XNOR U3733 ( .A(b[13]), .B(a[25]), .Z(n3531) );
  NANDN U3734 ( .A(n3531), .B(n8730), .Z(n3385) );
  NANDN U3735 ( .A(n3383), .B(n8731), .Z(n3384) );
  NAND U3736 ( .A(n3385), .B(n3384), .Z(n3447) );
  XNOR U3737 ( .A(n3450), .B(n3449), .Z(n3444) );
  NANDN U3738 ( .A(n315), .B(a[37]), .Z(n3386) );
  XNOR U3739 ( .A(b[1]), .B(n3386), .Z(n3388) );
  IV U3740 ( .A(a[36]), .Z(n7293) );
  NANDN U3741 ( .A(n7293), .B(n315), .Z(n3387) );
  AND U3742 ( .A(n3388), .B(n3387), .Z(n3468) );
  ANDN U3743 ( .B(b[31]), .A(n3389), .Z(n3465) );
  NANDN U3744 ( .A(n3390), .B(n9875), .Z(n3392) );
  XNOR U3745 ( .A(n322), .B(a[9]), .Z(n3537) );
  NANDN U3746 ( .A(n9874), .B(n3537), .Z(n3391) );
  NAND U3747 ( .A(n3392), .B(n3391), .Z(n3466) );
  XOR U3748 ( .A(n3465), .B(n3466), .Z(n3467) );
  XNOR U3749 ( .A(n3468), .B(n3467), .Z(n3441) );
  NANDN U3750 ( .A(n3393), .B(n9622), .Z(n3395) );
  XNOR U3751 ( .A(b[23]), .B(a[15]), .Z(n3540) );
  OR U3752 ( .A(n3540), .B(n9621), .Z(n3394) );
  NAND U3753 ( .A(n3395), .B(n3394), .Z(n3510) );
  XOR U3754 ( .A(b[7]), .B(a[31]), .Z(n3543) );
  NANDN U3755 ( .A(n8013), .B(n3543), .Z(n3398) );
  NANDN U3756 ( .A(n3396), .B(n8014), .Z(n3397) );
  NAND U3757 ( .A(n3398), .B(n3397), .Z(n3507) );
  XOR U3758 ( .A(b[25]), .B(n4578), .Z(n3546) );
  NANDN U3759 ( .A(n3546), .B(n9706), .Z(n3401) );
  NANDN U3760 ( .A(n3399), .B(n9707), .Z(n3400) );
  AND U3761 ( .A(n3401), .B(n3400), .Z(n3508) );
  XNOR U3762 ( .A(n3507), .B(n3508), .Z(n3509) );
  XNOR U3763 ( .A(n3510), .B(n3509), .Z(n3442) );
  XOR U3764 ( .A(n3444), .B(n3443), .Z(n3498) );
  XNOR U3765 ( .A(n3497), .B(n3498), .Z(n3555) );
  XNOR U3766 ( .A(n3556), .B(n3555), .Z(n3558) );
  XNOR U3767 ( .A(n3557), .B(n3558), .Z(n3567) );
  XOR U3768 ( .A(n3568), .B(n3567), .Z(n3570) );
  NAND U3769 ( .A(n3407), .B(n3406), .Z(n3411) );
  NANDN U3770 ( .A(n3409), .B(n3408), .Z(n3410) );
  AND U3771 ( .A(n3411), .B(n3410), .Z(n3561) );
  XNOR U3772 ( .A(n3562), .B(n3561), .Z(n3563) );
  XOR U3773 ( .A(n3564), .B(n3563), .Z(n3437) );
  NANDN U3774 ( .A(n3413), .B(n3412), .Z(n3417) );
  OR U3775 ( .A(n3415), .B(n3414), .Z(n3416) );
  NAND U3776 ( .A(n3417), .B(n3416), .Z(n3436) );
  NANDN U3777 ( .A(n3419), .B(n3418), .Z(n3423) );
  NANDN U3778 ( .A(n3421), .B(n3420), .Z(n3422) );
  AND U3779 ( .A(n3423), .B(n3422), .Z(n3435) );
  XNOR U3780 ( .A(n3436), .B(n3435), .Z(n3438) );
  XOR U3781 ( .A(n3437), .B(n3438), .Z(n3429) );
  XOR U3782 ( .A(n3430), .B(n3429), .Z(n3431) );
  XNOR U3783 ( .A(n3432), .B(n3431), .Z(n3573) );
  XNOR U3784 ( .A(n3573), .B(sreg[69]), .Z(n3575) );
  NAND U3785 ( .A(n3424), .B(sreg[68]), .Z(n3428) );
  OR U3786 ( .A(n3426), .B(n3425), .Z(n3427) );
  AND U3787 ( .A(n3428), .B(n3427), .Z(n3574) );
  XOR U3788 ( .A(n3575), .B(n3574), .Z(c[69]) );
  NAND U3789 ( .A(n3430), .B(n3429), .Z(n3434) );
  NAND U3790 ( .A(n3432), .B(n3431), .Z(n3433) );
  NAND U3791 ( .A(n3434), .B(n3433), .Z(n3581) );
  NANDN U3792 ( .A(n3436), .B(n3435), .Z(n3440) );
  NAND U3793 ( .A(n3438), .B(n3437), .Z(n3439) );
  NAND U3794 ( .A(n3440), .B(n3439), .Z(n3579) );
  OR U3795 ( .A(n3442), .B(n3441), .Z(n3446) );
  NANDN U3796 ( .A(n3444), .B(n3443), .Z(n3445) );
  NAND U3797 ( .A(n3446), .B(n3445), .Z(n3699) );
  OR U3798 ( .A(n3448), .B(n3447), .Z(n3452) );
  NANDN U3799 ( .A(n3450), .B(n3449), .Z(n3451) );
  NAND U3800 ( .A(n3452), .B(n3451), .Z(n3638) );
  NANDN U3801 ( .A(n3454), .B(n3453), .Z(n3458) );
  NANDN U3802 ( .A(n3456), .B(n3455), .Z(n3457) );
  NAND U3803 ( .A(n3458), .B(n3457), .Z(n3637) );
  NANDN U3804 ( .A(n3460), .B(n3459), .Z(n3464) );
  NANDN U3805 ( .A(n3462), .B(n3461), .Z(n3463) );
  NAND U3806 ( .A(n3464), .B(n3463), .Z(n3636) );
  XOR U3807 ( .A(n3638), .B(n3639), .Z(n3697) );
  OR U3808 ( .A(n3466), .B(n3465), .Z(n3470) );
  NANDN U3809 ( .A(n3468), .B(n3467), .Z(n3469) );
  NAND U3810 ( .A(n3470), .B(n3469), .Z(n3651) );
  NAND U3811 ( .A(n3471), .B(n9379), .Z(n3473) );
  XNOR U3812 ( .A(n9562), .B(a[20]), .Z(n3594) );
  NAND U3813 ( .A(n3594), .B(n9378), .Z(n3472) );
  NAND U3814 ( .A(n3473), .B(n3472), .Z(n3662) );
  NANDN U3815 ( .A(n3474), .B(n9801), .Z(n3476) );
  XNOR U3816 ( .A(b[27]), .B(a[12]), .Z(n3597) );
  OR U3817 ( .A(n3597), .B(n9751), .Z(n3475) );
  NAND U3818 ( .A(n3476), .B(n3475), .Z(n3660) );
  XNOR U3819 ( .A(b[5]), .B(a[34]), .Z(n3600) );
  NANDN U3820 ( .A(n3600), .B(n7905), .Z(n3479) );
  NANDN U3821 ( .A(n3477), .B(n7906), .Z(n3478) );
  AND U3822 ( .A(n3479), .B(n3478), .Z(n3661) );
  XNOR U3823 ( .A(n3660), .B(n3661), .Z(n3663) );
  XOR U3824 ( .A(n3662), .B(n3663), .Z(n3648) );
  NAND U3825 ( .A(n3480), .B(n9105), .Z(n3482) );
  XNOR U3826 ( .A(n9455), .B(a[22]), .Z(n3603) );
  NAND U3827 ( .A(n3603), .B(n9107), .Z(n3481) );
  NAND U3828 ( .A(n3482), .B(n3481), .Z(n3620) );
  NAND U3829 ( .A(n3483), .B(n9914), .Z(n3485) );
  XNOR U3830 ( .A(n323), .B(a[8]), .Z(n3606) );
  NANDN U3831 ( .A(n9913), .B(n3606), .Z(n3484) );
  NAND U3832 ( .A(n3485), .B(n3484), .Z(n3618) );
  NAND U3833 ( .A(n3486), .B(n7622), .Z(n3488) );
  XNOR U3834 ( .A(n316), .B(a[36]), .Z(n3609) );
  NAND U3835 ( .A(n3609), .B(n7620), .Z(n3487) );
  NAND U3836 ( .A(n3488), .B(n3487), .Z(n3619) );
  XOR U3837 ( .A(n3618), .B(n3619), .Z(n3621) );
  XOR U3838 ( .A(n3620), .B(n3621), .Z(n3649) );
  XOR U3839 ( .A(n3648), .B(n3649), .Z(n3650) );
  XNOR U3840 ( .A(n3651), .B(n3650), .Z(n3696) );
  XOR U3841 ( .A(n3697), .B(n3696), .Z(n3698) );
  XNOR U3842 ( .A(n3699), .B(n3698), .Z(n3715) );
  OR U3843 ( .A(n3490), .B(n3489), .Z(n3494) );
  NAND U3844 ( .A(n3492), .B(n3491), .Z(n3493) );
  NAND U3845 ( .A(n3494), .B(n3493), .Z(n3713) );
  NANDN U3846 ( .A(n3496), .B(n3495), .Z(n3500) );
  NANDN U3847 ( .A(n3498), .B(n3497), .Z(n3499) );
  NAND U3848 ( .A(n3500), .B(n3499), .Z(n3702) );
  NAND U3849 ( .A(n3502), .B(n3501), .Z(n3506) );
  NAND U3850 ( .A(n3504), .B(n3503), .Z(n3505) );
  NAND U3851 ( .A(n3506), .B(n3505), .Z(n3701) );
  NANDN U3852 ( .A(n3508), .B(n3507), .Z(n3512) );
  NAND U3853 ( .A(n3510), .B(n3509), .Z(n3511) );
  NAND U3854 ( .A(n3512), .B(n3511), .Z(n3642) );
  NANDN U3855 ( .A(n3514), .B(n3513), .Z(n3518) );
  NAND U3856 ( .A(n3516), .B(n3515), .Z(n3517) );
  AND U3857 ( .A(n3518), .B(n3517), .Z(n3643) );
  XNOR U3858 ( .A(n3642), .B(n3643), .Z(n3644) );
  NAND U3859 ( .A(n3519), .B(n8286), .Z(n3521) );
  XNOR U3860 ( .A(b[9]), .B(n6135), .Z(n3666) );
  NAND U3861 ( .A(n3666), .B(n8288), .Z(n3520) );
  NAND U3862 ( .A(n3521), .B(n3520), .Z(n3626) );
  NAND U3863 ( .A(n3522), .B(n8961), .Z(n3524) );
  XOR U3864 ( .A(b[15]), .B(a[24]), .Z(n3669) );
  NAND U3865 ( .A(n3669), .B(n8963), .Z(n3523) );
  NAND U3866 ( .A(n3524), .B(n3523), .Z(n3624) );
  XNOR U3867 ( .A(b[21]), .B(a[18]), .Z(n3672) );
  NANDN U3868 ( .A(n3672), .B(n9493), .Z(n3527) );
  NANDN U3869 ( .A(n3525), .B(n9495), .Z(n3526) );
  AND U3870 ( .A(n3527), .B(n3526), .Z(n3625) );
  XOR U3871 ( .A(n3624), .B(n3625), .Z(n3627) );
  XNOR U3872 ( .A(n3626), .B(n3627), .Z(n3615) );
  XNOR U3873 ( .A(b[11]), .B(a[28]), .Z(n3675) );
  NANDN U3874 ( .A(n3675), .B(n8541), .Z(n3530) );
  NANDN U3875 ( .A(n3528), .B(n8542), .Z(n3529) );
  NAND U3876 ( .A(n3530), .B(n3529), .Z(n3613) );
  XOR U3877 ( .A(b[13]), .B(n6500), .Z(n3678) );
  NANDN U3878 ( .A(n3678), .B(n8730), .Z(n3533) );
  NANDN U3879 ( .A(n3531), .B(n8731), .Z(n3532) );
  AND U3880 ( .A(n3533), .B(n3532), .Z(n3612) );
  XNOR U3881 ( .A(n3613), .B(n3612), .Z(n3614) );
  XNOR U3882 ( .A(n3615), .B(n3614), .Z(n3632) );
  NANDN U3883 ( .A(n315), .B(a[38]), .Z(n3534) );
  XNOR U3884 ( .A(b[1]), .B(n3534), .Z(n3536) );
  NANDN U3885 ( .A(b[0]), .B(a[37]), .Z(n3535) );
  AND U3886 ( .A(n3536), .B(n3535), .Z(n3590) );
  NAND U3887 ( .A(n3537), .B(n9875), .Z(n3539) );
  XNOR U3888 ( .A(n322), .B(a[10]), .Z(n3684) );
  NANDN U3889 ( .A(n9874), .B(n3684), .Z(n3538) );
  NAND U3890 ( .A(n3539), .B(n3538), .Z(n3588) );
  NANDN U3891 ( .A(n323), .B(a[6]), .Z(n3589) );
  XNOR U3892 ( .A(n3588), .B(n3589), .Z(n3591) );
  XOR U3893 ( .A(n3590), .B(n3591), .Z(n3630) );
  NANDN U3894 ( .A(n3540), .B(n9622), .Z(n3542) );
  XNOR U3895 ( .A(b[23]), .B(a[16]), .Z(n3687) );
  OR U3896 ( .A(n3687), .B(n9621), .Z(n3541) );
  NAND U3897 ( .A(n3542), .B(n3541), .Z(n3657) );
  XOR U3898 ( .A(b[7]), .B(a[32]), .Z(n3690) );
  NANDN U3899 ( .A(n8013), .B(n3690), .Z(n3545) );
  NAND U3900 ( .A(n3543), .B(n8014), .Z(n3544) );
  NAND U3901 ( .A(n3545), .B(n3544), .Z(n3654) );
  XNOR U3902 ( .A(b[25]), .B(a[14]), .Z(n3693) );
  NANDN U3903 ( .A(n3693), .B(n9706), .Z(n3548) );
  NANDN U3904 ( .A(n3546), .B(n9707), .Z(n3547) );
  AND U3905 ( .A(n3548), .B(n3547), .Z(n3655) );
  XNOR U3906 ( .A(n3654), .B(n3655), .Z(n3656) );
  XNOR U3907 ( .A(n3657), .B(n3656), .Z(n3631) );
  XOR U3908 ( .A(n3630), .B(n3631), .Z(n3633) );
  XNOR U3909 ( .A(n3632), .B(n3633), .Z(n3645) );
  XNOR U3910 ( .A(n3644), .B(n3645), .Z(n3700) );
  XNOR U3911 ( .A(n3701), .B(n3700), .Z(n3703) );
  XNOR U3912 ( .A(n3702), .B(n3703), .Z(n3712) );
  XNOR U3913 ( .A(n3713), .B(n3712), .Z(n3714) );
  XOR U3914 ( .A(n3715), .B(n3714), .Z(n3709) );
  NANDN U3915 ( .A(n3550), .B(n3549), .Z(n3554) );
  OR U3916 ( .A(n3552), .B(n3551), .Z(n3553) );
  NAND U3917 ( .A(n3554), .B(n3553), .Z(n3706) );
  NAND U3918 ( .A(n3556), .B(n3555), .Z(n3560) );
  NANDN U3919 ( .A(n3558), .B(n3557), .Z(n3559) );
  NAND U3920 ( .A(n3560), .B(n3559), .Z(n3707) );
  XNOR U3921 ( .A(n3706), .B(n3707), .Z(n3708) );
  XNOR U3922 ( .A(n3709), .B(n3708), .Z(n3585) );
  NANDN U3923 ( .A(n3562), .B(n3561), .Z(n3566) );
  NAND U3924 ( .A(n3564), .B(n3563), .Z(n3565) );
  NAND U3925 ( .A(n3566), .B(n3565), .Z(n3582) );
  NANDN U3926 ( .A(n3568), .B(n3567), .Z(n3572) );
  OR U3927 ( .A(n3570), .B(n3569), .Z(n3571) );
  NAND U3928 ( .A(n3572), .B(n3571), .Z(n3583) );
  XNOR U3929 ( .A(n3582), .B(n3583), .Z(n3584) );
  XNOR U3930 ( .A(n3585), .B(n3584), .Z(n3578) );
  XOR U3931 ( .A(n3579), .B(n3578), .Z(n3580) );
  XNOR U3932 ( .A(n3581), .B(n3580), .Z(n3718) );
  XNOR U3933 ( .A(n3718), .B(sreg[70]), .Z(n3720) );
  NAND U3934 ( .A(n3573), .B(sreg[69]), .Z(n3577) );
  OR U3935 ( .A(n3575), .B(n3574), .Z(n3576) );
  AND U3936 ( .A(n3577), .B(n3576), .Z(n3719) );
  XOR U3937 ( .A(n3720), .B(n3719), .Z(c[70]) );
  NANDN U3938 ( .A(n3583), .B(n3582), .Z(n3587) );
  NANDN U3939 ( .A(n3585), .B(n3584), .Z(n3586) );
  NAND U3940 ( .A(n3587), .B(n3586), .Z(n3724) );
  NANDN U3941 ( .A(n3589), .B(n3588), .Z(n3593) );
  NAND U3942 ( .A(n3591), .B(n3590), .Z(n3592) );
  NAND U3943 ( .A(n3593), .B(n3592), .Z(n3798) );
  NAND U3944 ( .A(n3594), .B(n9379), .Z(n3596) );
  XNOR U3945 ( .A(n9562), .B(a[21]), .Z(n3741) );
  NAND U3946 ( .A(n3741), .B(n9378), .Z(n3595) );
  NAND U3947 ( .A(n3596), .B(n3595), .Z(n3809) );
  NANDN U3948 ( .A(n3597), .B(n9801), .Z(n3599) );
  XOR U3949 ( .A(b[27]), .B(n4578), .Z(n3744) );
  OR U3950 ( .A(n3744), .B(n9751), .Z(n3598) );
  NAND U3951 ( .A(n3599), .B(n3598), .Z(n3807) );
  XNOR U3952 ( .A(b[5]), .B(a[35]), .Z(n3747) );
  NANDN U3953 ( .A(n3747), .B(n7905), .Z(n3602) );
  NANDN U3954 ( .A(n3600), .B(n7906), .Z(n3601) );
  AND U3955 ( .A(n3602), .B(n3601), .Z(n3808) );
  XNOR U3956 ( .A(n3807), .B(n3808), .Z(n3810) );
  XOR U3957 ( .A(n3809), .B(n3810), .Z(n3795) );
  NAND U3958 ( .A(n3603), .B(n9105), .Z(n3605) );
  XNOR U3959 ( .A(n9455), .B(a[23]), .Z(n3750) );
  NAND U3960 ( .A(n3750), .B(n9107), .Z(n3604) );
  NAND U3961 ( .A(n3605), .B(n3604), .Z(n3767) );
  NAND U3962 ( .A(n3606), .B(n9914), .Z(n3608) );
  XNOR U3963 ( .A(n323), .B(a[9]), .Z(n3753) );
  NANDN U3964 ( .A(n9913), .B(n3753), .Z(n3607) );
  NAND U3965 ( .A(n3608), .B(n3607), .Z(n3765) );
  NAND U3966 ( .A(n3609), .B(n7622), .Z(n3611) );
  XNOR U3967 ( .A(n316), .B(a[37]), .Z(n3756) );
  NAND U3968 ( .A(n3756), .B(n7620), .Z(n3610) );
  NAND U3969 ( .A(n3611), .B(n3610), .Z(n3766) );
  XOR U3970 ( .A(n3765), .B(n3766), .Z(n3768) );
  XOR U3971 ( .A(n3767), .B(n3768), .Z(n3796) );
  XOR U3972 ( .A(n3795), .B(n3796), .Z(n3797) );
  XNOR U3973 ( .A(n3798), .B(n3797), .Z(n3844) );
  NANDN U3974 ( .A(n3613), .B(n3612), .Z(n3617) );
  NANDN U3975 ( .A(n3615), .B(n3614), .Z(n3616) );
  NAND U3976 ( .A(n3617), .B(n3616), .Z(n3786) );
  NAND U3977 ( .A(n3619), .B(n3618), .Z(n3623) );
  NAND U3978 ( .A(n3621), .B(n3620), .Z(n3622) );
  NAND U3979 ( .A(n3623), .B(n3622), .Z(n3784) );
  NANDN U3980 ( .A(n3625), .B(n3624), .Z(n3629) );
  NANDN U3981 ( .A(n3627), .B(n3626), .Z(n3628) );
  NAND U3982 ( .A(n3629), .B(n3628), .Z(n3783) );
  XNOR U3983 ( .A(n3786), .B(n3785), .Z(n3845) );
  XOR U3984 ( .A(n3844), .B(n3845), .Z(n3847) );
  NANDN U3985 ( .A(n3631), .B(n3630), .Z(n3635) );
  OR U3986 ( .A(n3633), .B(n3632), .Z(n3634) );
  NAND U3987 ( .A(n3635), .B(n3634), .Z(n3846) );
  XOR U3988 ( .A(n3847), .B(n3846), .Z(n3864) );
  OR U3989 ( .A(n3637), .B(n3636), .Z(n3641) );
  NANDN U3990 ( .A(n3639), .B(n3638), .Z(n3640) );
  NAND U3991 ( .A(n3641), .B(n3640), .Z(n3863) );
  NANDN U3992 ( .A(n3643), .B(n3642), .Z(n3647) );
  NANDN U3993 ( .A(n3645), .B(n3644), .Z(n3646) );
  NAND U3994 ( .A(n3647), .B(n3646), .Z(n3852) );
  NAND U3995 ( .A(n3649), .B(n3648), .Z(n3653) );
  NANDN U3996 ( .A(n3651), .B(n3650), .Z(n3652) );
  NAND U3997 ( .A(n3653), .B(n3652), .Z(n3851) );
  NANDN U3998 ( .A(n3655), .B(n3654), .Z(n3659) );
  NAND U3999 ( .A(n3657), .B(n3656), .Z(n3658) );
  NAND U4000 ( .A(n3659), .B(n3658), .Z(n3789) );
  NANDN U4001 ( .A(n3661), .B(n3660), .Z(n3665) );
  NAND U4002 ( .A(n3663), .B(n3662), .Z(n3664) );
  AND U4003 ( .A(n3665), .B(n3664), .Z(n3790) );
  XNOR U4004 ( .A(n3789), .B(n3790), .Z(n3791) );
  NAND U4005 ( .A(n3666), .B(n8286), .Z(n3668) );
  XOR U4006 ( .A(b[9]), .B(a[31]), .Z(n3813) );
  NAND U4007 ( .A(n3813), .B(n8288), .Z(n3667) );
  NAND U4008 ( .A(n3668), .B(n3667), .Z(n3773) );
  NAND U4009 ( .A(n3669), .B(n8961), .Z(n3671) );
  XOR U4010 ( .A(b[15]), .B(a[25]), .Z(n3816) );
  NAND U4011 ( .A(n3816), .B(n8963), .Z(n3670) );
  NAND U4012 ( .A(n3671), .B(n3670), .Z(n3771) );
  XNOR U4013 ( .A(b[21]), .B(a[19]), .Z(n3819) );
  NANDN U4014 ( .A(n3819), .B(n9493), .Z(n3674) );
  NANDN U4015 ( .A(n3672), .B(n9495), .Z(n3673) );
  AND U4016 ( .A(n3674), .B(n3673), .Z(n3772) );
  XOR U4017 ( .A(n3771), .B(n3772), .Z(n3774) );
  XNOR U4018 ( .A(n3773), .B(n3774), .Z(n3762) );
  XNOR U4019 ( .A(b[11]), .B(a[29]), .Z(n3822) );
  NANDN U4020 ( .A(n3822), .B(n8541), .Z(n3677) );
  NANDN U4021 ( .A(n3675), .B(n8542), .Z(n3676) );
  NAND U4022 ( .A(n3677), .B(n3676), .Z(n3760) );
  XNOR U4023 ( .A(b[13]), .B(a[27]), .Z(n3825) );
  NANDN U4024 ( .A(n3825), .B(n8730), .Z(n3680) );
  NANDN U4025 ( .A(n3678), .B(n8731), .Z(n3679) );
  AND U4026 ( .A(n3680), .B(n3679), .Z(n3759) );
  XNOR U4027 ( .A(n3760), .B(n3759), .Z(n3761) );
  XNOR U4028 ( .A(n3762), .B(n3761), .Z(n3779) );
  NANDN U4029 ( .A(n315), .B(a[39]), .Z(n3681) );
  XNOR U4030 ( .A(b[1]), .B(n3681), .Z(n3683) );
  IV U4031 ( .A(a[38]), .Z(n7672) );
  NANDN U4032 ( .A(n7672), .B(n315), .Z(n3682) );
  AND U4033 ( .A(n3683), .B(n3682), .Z(n3737) );
  NAND U4034 ( .A(n9875), .B(n3684), .Z(n3686) );
  XNOR U4035 ( .A(b[29]), .B(a[11]), .Z(n3832) );
  OR U4036 ( .A(n3832), .B(n9874), .Z(n3685) );
  NAND U4037 ( .A(n3686), .B(n3685), .Z(n3735) );
  NANDN U4038 ( .A(n323), .B(a[7]), .Z(n3736) );
  XNOR U4039 ( .A(n3735), .B(n3736), .Z(n3738) );
  XOR U4040 ( .A(n3737), .B(n3738), .Z(n3777) );
  NANDN U4041 ( .A(n3687), .B(n9622), .Z(n3689) );
  XOR U4042 ( .A(b[23]), .B(n5168), .Z(n3835) );
  OR U4043 ( .A(n3835), .B(n9621), .Z(n3688) );
  NAND U4044 ( .A(n3689), .B(n3688), .Z(n3804) );
  XNOR U4045 ( .A(b[7]), .B(a[33]), .Z(n3838) );
  OR U4046 ( .A(n3838), .B(n8013), .Z(n3692) );
  NAND U4047 ( .A(n3690), .B(n8014), .Z(n3691) );
  NAND U4048 ( .A(n3692), .B(n3691), .Z(n3801) );
  XNOR U4049 ( .A(b[25]), .B(a[15]), .Z(n3841) );
  NANDN U4050 ( .A(n3841), .B(n9706), .Z(n3695) );
  NANDN U4051 ( .A(n3693), .B(n9707), .Z(n3694) );
  AND U4052 ( .A(n3695), .B(n3694), .Z(n3802) );
  XNOR U4053 ( .A(n3801), .B(n3802), .Z(n3803) );
  XNOR U4054 ( .A(n3804), .B(n3803), .Z(n3778) );
  XOR U4055 ( .A(n3777), .B(n3778), .Z(n3780) );
  XNOR U4056 ( .A(n3779), .B(n3780), .Z(n3792) );
  XNOR U4057 ( .A(n3791), .B(n3792), .Z(n3850) );
  XNOR U4058 ( .A(n3851), .B(n3850), .Z(n3853) );
  XNOR U4059 ( .A(n3852), .B(n3853), .Z(n3862) );
  XOR U4060 ( .A(n3863), .B(n3862), .Z(n3865) );
  NAND U4061 ( .A(n3701), .B(n3700), .Z(n3705) );
  NANDN U4062 ( .A(n3703), .B(n3702), .Z(n3704) );
  AND U4063 ( .A(n3705), .B(n3704), .Z(n3856) );
  XNOR U4064 ( .A(n3857), .B(n3856), .Z(n3858) );
  XOR U4065 ( .A(n3859), .B(n3858), .Z(n3731) );
  NANDN U4066 ( .A(n3707), .B(n3706), .Z(n3711) );
  NAND U4067 ( .A(n3709), .B(n3708), .Z(n3710) );
  NAND U4068 ( .A(n3711), .B(n3710), .Z(n3729) );
  NANDN U4069 ( .A(n3713), .B(n3712), .Z(n3717) );
  NANDN U4070 ( .A(n3715), .B(n3714), .Z(n3716) );
  NAND U4071 ( .A(n3717), .B(n3716), .Z(n3730) );
  XNOR U4072 ( .A(n3729), .B(n3730), .Z(n3732) );
  XOR U4073 ( .A(n3731), .B(n3732), .Z(n3723) );
  XOR U4074 ( .A(n3724), .B(n3723), .Z(n3725) );
  XNOR U4075 ( .A(n3726), .B(n3725), .Z(n3868) );
  XNOR U4076 ( .A(n3868), .B(sreg[71]), .Z(n3870) );
  NAND U4077 ( .A(n3718), .B(sreg[70]), .Z(n3722) );
  OR U4078 ( .A(n3720), .B(n3719), .Z(n3721) );
  AND U4079 ( .A(n3722), .B(n3721), .Z(n3869) );
  XOR U4080 ( .A(n3870), .B(n3869), .Z(c[71]) );
  NAND U4081 ( .A(n3724), .B(n3723), .Z(n3728) );
  NAND U4082 ( .A(n3726), .B(n3725), .Z(n3727) );
  NAND U4083 ( .A(n3728), .B(n3727), .Z(n3876) );
  NANDN U4084 ( .A(n3730), .B(n3729), .Z(n3734) );
  NAND U4085 ( .A(n3732), .B(n3731), .Z(n3733) );
  NAND U4086 ( .A(n3734), .B(n3733), .Z(n3874) );
  NANDN U4087 ( .A(n3736), .B(n3735), .Z(n3740) );
  NAND U4088 ( .A(n3738), .B(n3737), .Z(n3739) );
  NAND U4089 ( .A(n3740), .B(n3739), .Z(n3948) );
  NAND U4090 ( .A(n3741), .B(n9379), .Z(n3743) );
  XNOR U4091 ( .A(n9562), .B(a[22]), .Z(n3915) );
  NAND U4092 ( .A(n3915), .B(n9378), .Z(n3742) );
  NAND U4093 ( .A(n3743), .B(n3742), .Z(n3959) );
  NANDN U4094 ( .A(n3744), .B(n9801), .Z(n3746) );
  XNOR U4095 ( .A(b[27]), .B(a[14]), .Z(n3918) );
  OR U4096 ( .A(n3918), .B(n9751), .Z(n3745) );
  NAND U4097 ( .A(n3746), .B(n3745), .Z(n3957) );
  XOR U4098 ( .A(b[5]), .B(n7293), .Z(n3921) );
  NANDN U4099 ( .A(n3921), .B(n7905), .Z(n3749) );
  NANDN U4100 ( .A(n3747), .B(n7906), .Z(n3748) );
  AND U4101 ( .A(n3749), .B(n3748), .Z(n3958) );
  XNOR U4102 ( .A(n3957), .B(n3958), .Z(n3960) );
  XOR U4103 ( .A(n3959), .B(n3960), .Z(n3945) );
  NAND U4104 ( .A(n3750), .B(n9105), .Z(n3752) );
  XNOR U4105 ( .A(n9455), .B(a[24]), .Z(n3924) );
  NAND U4106 ( .A(n3924), .B(n9107), .Z(n3751) );
  AND U4107 ( .A(n3752), .B(n3751), .Z(n3900) );
  NAND U4108 ( .A(n3753), .B(n9914), .Z(n3755) );
  XNOR U4109 ( .A(n323), .B(a[10]), .Z(n3927) );
  NANDN U4110 ( .A(n9913), .B(n3927), .Z(n3754) );
  AND U4111 ( .A(n3755), .B(n3754), .Z(n3898) );
  NAND U4112 ( .A(n3756), .B(n7622), .Z(n3758) );
  XNOR U4113 ( .A(n7672), .B(b[3]), .Z(n3930) );
  NAND U4114 ( .A(n3930), .B(n7620), .Z(n3757) );
  NAND U4115 ( .A(n3758), .B(n3757), .Z(n3897) );
  XOR U4116 ( .A(n3945), .B(n3946), .Z(n3947) );
  XNOR U4117 ( .A(n3948), .B(n3947), .Z(n3993) );
  NANDN U4118 ( .A(n3760), .B(n3759), .Z(n3764) );
  NANDN U4119 ( .A(n3762), .B(n3761), .Z(n3763) );
  NAND U4120 ( .A(n3764), .B(n3763), .Z(n3936) );
  NAND U4121 ( .A(n3766), .B(n3765), .Z(n3770) );
  NAND U4122 ( .A(n3768), .B(n3767), .Z(n3769) );
  NAND U4123 ( .A(n3770), .B(n3769), .Z(n3934) );
  NANDN U4124 ( .A(n3772), .B(n3771), .Z(n3776) );
  NANDN U4125 ( .A(n3774), .B(n3773), .Z(n3775) );
  NAND U4126 ( .A(n3776), .B(n3775), .Z(n3933) );
  XNOR U4127 ( .A(n3936), .B(n3935), .Z(n3994) );
  XOR U4128 ( .A(n3993), .B(n3994), .Z(n3996) );
  NANDN U4129 ( .A(n3778), .B(n3777), .Z(n3782) );
  OR U4130 ( .A(n3780), .B(n3779), .Z(n3781) );
  NAND U4131 ( .A(n3782), .B(n3781), .Z(n3995) );
  XOR U4132 ( .A(n3996), .B(n3995), .Z(n4013) );
  OR U4133 ( .A(n3784), .B(n3783), .Z(n3788) );
  NAND U4134 ( .A(n3786), .B(n3785), .Z(n3787) );
  NAND U4135 ( .A(n3788), .B(n3787), .Z(n4012) );
  NANDN U4136 ( .A(n3790), .B(n3789), .Z(n3794) );
  NANDN U4137 ( .A(n3792), .B(n3791), .Z(n3793) );
  NAND U4138 ( .A(n3794), .B(n3793), .Z(n4001) );
  NAND U4139 ( .A(n3796), .B(n3795), .Z(n3800) );
  NAND U4140 ( .A(n3798), .B(n3797), .Z(n3799) );
  NAND U4141 ( .A(n3800), .B(n3799), .Z(n4000) );
  NANDN U4142 ( .A(n3802), .B(n3801), .Z(n3806) );
  NAND U4143 ( .A(n3804), .B(n3803), .Z(n3805) );
  NAND U4144 ( .A(n3806), .B(n3805), .Z(n3939) );
  NANDN U4145 ( .A(n3808), .B(n3807), .Z(n3812) );
  NAND U4146 ( .A(n3810), .B(n3809), .Z(n3811) );
  AND U4147 ( .A(n3812), .B(n3811), .Z(n3940) );
  XNOR U4148 ( .A(n3939), .B(n3940), .Z(n3941) );
  NAND U4149 ( .A(n3813), .B(n8286), .Z(n3815) );
  XOR U4150 ( .A(b[9]), .B(a[32]), .Z(n3963) );
  NAND U4151 ( .A(n3963), .B(n8288), .Z(n3814) );
  NAND U4152 ( .A(n3815), .B(n3814), .Z(n3905) );
  NAND U4153 ( .A(n3816), .B(n8961), .Z(n3818) );
  XNOR U4154 ( .A(b[15]), .B(n6500), .Z(n3966) );
  NAND U4155 ( .A(n3966), .B(n8963), .Z(n3817) );
  NAND U4156 ( .A(n3818), .B(n3817), .Z(n3903) );
  XNOR U4157 ( .A(b[21]), .B(a[20]), .Z(n3969) );
  NANDN U4158 ( .A(n3969), .B(n9493), .Z(n3821) );
  NANDN U4159 ( .A(n3819), .B(n9495), .Z(n3820) );
  AND U4160 ( .A(n3821), .B(n3820), .Z(n3904) );
  XOR U4161 ( .A(n3903), .B(n3904), .Z(n3906) );
  XNOR U4162 ( .A(n3905), .B(n3906), .Z(n3894) );
  XOR U4163 ( .A(b[11]), .B(n6135), .Z(n3972) );
  NANDN U4164 ( .A(n3972), .B(n8541), .Z(n3824) );
  NANDN U4165 ( .A(n3822), .B(n8542), .Z(n3823) );
  NAND U4166 ( .A(n3824), .B(n3823), .Z(n3892) );
  XNOR U4167 ( .A(b[13]), .B(a[28]), .Z(n3975) );
  NANDN U4168 ( .A(n3975), .B(n8730), .Z(n3827) );
  NANDN U4169 ( .A(n3825), .B(n8731), .Z(n3826) );
  NAND U4170 ( .A(n3827), .B(n3826), .Z(n3891) );
  XNOR U4171 ( .A(n3894), .B(n3893), .Z(n3888) );
  NANDN U4172 ( .A(n315), .B(a[40]), .Z(n3828) );
  XNOR U4173 ( .A(b[1]), .B(n3828), .Z(n3830) );
  NANDN U4174 ( .A(b[0]), .B(a[39]), .Z(n3829) );
  AND U4175 ( .A(n3830), .B(n3829), .Z(n3912) );
  ANDN U4176 ( .B(b[31]), .A(n3831), .Z(n3909) );
  NANDN U4177 ( .A(n3832), .B(n9875), .Z(n3834) );
  XNOR U4178 ( .A(n322), .B(a[12]), .Z(n3981) );
  NANDN U4179 ( .A(n9874), .B(n3981), .Z(n3833) );
  NAND U4180 ( .A(n3834), .B(n3833), .Z(n3910) );
  XOR U4181 ( .A(n3909), .B(n3910), .Z(n3911) );
  XNOR U4182 ( .A(n3912), .B(n3911), .Z(n3885) );
  NANDN U4183 ( .A(n3835), .B(n9622), .Z(n3837) );
  XNOR U4184 ( .A(b[23]), .B(a[18]), .Z(n3984) );
  OR U4185 ( .A(n3984), .B(n9621), .Z(n3836) );
  NAND U4186 ( .A(n3837), .B(n3836), .Z(n3954) );
  XOR U4187 ( .A(b[7]), .B(a[34]), .Z(n3987) );
  NANDN U4188 ( .A(n8013), .B(n3987), .Z(n3840) );
  NANDN U4189 ( .A(n3838), .B(n8014), .Z(n3839) );
  NAND U4190 ( .A(n3840), .B(n3839), .Z(n3951) );
  XNOR U4191 ( .A(b[25]), .B(a[16]), .Z(n3990) );
  NANDN U4192 ( .A(n3990), .B(n9706), .Z(n3843) );
  NANDN U4193 ( .A(n3841), .B(n9707), .Z(n3842) );
  AND U4194 ( .A(n3843), .B(n3842), .Z(n3952) );
  XNOR U4195 ( .A(n3951), .B(n3952), .Z(n3953) );
  XNOR U4196 ( .A(n3954), .B(n3953), .Z(n3886) );
  XOR U4197 ( .A(n3888), .B(n3887), .Z(n3942) );
  XNOR U4198 ( .A(n3941), .B(n3942), .Z(n3999) );
  XNOR U4199 ( .A(n4000), .B(n3999), .Z(n4002) );
  XNOR U4200 ( .A(n4001), .B(n4002), .Z(n4011) );
  XOR U4201 ( .A(n4012), .B(n4011), .Z(n4014) );
  NANDN U4202 ( .A(n3845), .B(n3844), .Z(n3849) );
  OR U4203 ( .A(n3847), .B(n3846), .Z(n3848) );
  NAND U4204 ( .A(n3849), .B(n3848), .Z(n4005) );
  NAND U4205 ( .A(n3851), .B(n3850), .Z(n3855) );
  NANDN U4206 ( .A(n3853), .B(n3852), .Z(n3854) );
  NAND U4207 ( .A(n3855), .B(n3854), .Z(n4006) );
  XNOR U4208 ( .A(n4005), .B(n4006), .Z(n4007) );
  XOR U4209 ( .A(n4008), .B(n4007), .Z(n3881) );
  NANDN U4210 ( .A(n3857), .B(n3856), .Z(n3861) );
  NAND U4211 ( .A(n3859), .B(n3858), .Z(n3860) );
  NAND U4212 ( .A(n3861), .B(n3860), .Z(n3879) );
  NANDN U4213 ( .A(n3863), .B(n3862), .Z(n3867) );
  OR U4214 ( .A(n3865), .B(n3864), .Z(n3866) );
  NAND U4215 ( .A(n3867), .B(n3866), .Z(n3880) );
  XNOR U4216 ( .A(n3879), .B(n3880), .Z(n3882) );
  XOR U4217 ( .A(n3881), .B(n3882), .Z(n3873) );
  XOR U4218 ( .A(n3874), .B(n3873), .Z(n3875) );
  XNOR U4219 ( .A(n3876), .B(n3875), .Z(n4017) );
  XNOR U4220 ( .A(n4017), .B(sreg[72]), .Z(n4019) );
  NAND U4221 ( .A(n3868), .B(sreg[71]), .Z(n3872) );
  OR U4222 ( .A(n3870), .B(n3869), .Z(n3871) );
  AND U4223 ( .A(n3872), .B(n3871), .Z(n4018) );
  XOR U4224 ( .A(n4019), .B(n4018), .Z(c[72]) );
  NAND U4225 ( .A(n3874), .B(n3873), .Z(n3878) );
  NAND U4226 ( .A(n3876), .B(n3875), .Z(n3877) );
  NAND U4227 ( .A(n3878), .B(n3877), .Z(n4025) );
  NANDN U4228 ( .A(n3880), .B(n3879), .Z(n3884) );
  NAND U4229 ( .A(n3882), .B(n3881), .Z(n3883) );
  NAND U4230 ( .A(n3884), .B(n3883), .Z(n4023) );
  OR U4231 ( .A(n3886), .B(n3885), .Z(n3890) );
  NANDN U4232 ( .A(n3888), .B(n3887), .Z(n3889) );
  NAND U4233 ( .A(n3890), .B(n3889), .Z(n4155) );
  OR U4234 ( .A(n3892), .B(n3891), .Z(n3896) );
  NANDN U4235 ( .A(n3894), .B(n3893), .Z(n3895) );
  NAND U4236 ( .A(n3896), .B(n3895), .Z(n4094) );
  NANDN U4237 ( .A(n3898), .B(n3897), .Z(n3902) );
  NANDN U4238 ( .A(n3900), .B(n3899), .Z(n3901) );
  NAND U4239 ( .A(n3902), .B(n3901), .Z(n4093) );
  NANDN U4240 ( .A(n3904), .B(n3903), .Z(n3908) );
  NANDN U4241 ( .A(n3906), .B(n3905), .Z(n3907) );
  NAND U4242 ( .A(n3908), .B(n3907), .Z(n4092) );
  XOR U4243 ( .A(n4094), .B(n4095), .Z(n4153) );
  OR U4244 ( .A(n3910), .B(n3909), .Z(n3914) );
  NANDN U4245 ( .A(n3912), .B(n3911), .Z(n3913) );
  NAND U4246 ( .A(n3914), .B(n3913), .Z(n4107) );
  NAND U4247 ( .A(n3915), .B(n9379), .Z(n3917) );
  XNOR U4248 ( .A(n9562), .B(a[23]), .Z(n4050) );
  NAND U4249 ( .A(n4050), .B(n9378), .Z(n3916) );
  NAND U4250 ( .A(n3917), .B(n3916), .Z(n4118) );
  NANDN U4251 ( .A(n3918), .B(n9801), .Z(n3920) );
  XNOR U4252 ( .A(b[27]), .B(a[15]), .Z(n4053) );
  OR U4253 ( .A(n4053), .B(n9751), .Z(n3919) );
  NAND U4254 ( .A(n3920), .B(n3919), .Z(n4116) );
  XNOR U4255 ( .A(b[5]), .B(a[37]), .Z(n4056) );
  NANDN U4256 ( .A(n4056), .B(n7905), .Z(n3923) );
  NANDN U4257 ( .A(n3921), .B(n7906), .Z(n3922) );
  AND U4258 ( .A(n3923), .B(n3922), .Z(n4117) );
  XNOR U4259 ( .A(n4116), .B(n4117), .Z(n4119) );
  XOR U4260 ( .A(n4118), .B(n4119), .Z(n4104) );
  NAND U4261 ( .A(n3924), .B(n9105), .Z(n3926) );
  XNOR U4262 ( .A(n9455), .B(a[25]), .Z(n4059) );
  NAND U4263 ( .A(n4059), .B(n9107), .Z(n3925) );
  NAND U4264 ( .A(n3926), .B(n3925), .Z(n4076) );
  NAND U4265 ( .A(n3927), .B(n9914), .Z(n3929) );
  XNOR U4266 ( .A(n323), .B(a[11]), .Z(n4062) );
  NANDN U4267 ( .A(n9913), .B(n4062), .Z(n3928) );
  NAND U4268 ( .A(n3929), .B(n3928), .Z(n4074) );
  NAND U4269 ( .A(n3930), .B(n7622), .Z(n3932) );
  XNOR U4270 ( .A(a[39]), .B(n316), .Z(n4065) );
  NAND U4271 ( .A(n4065), .B(n7620), .Z(n3931) );
  NAND U4272 ( .A(n3932), .B(n3931), .Z(n4075) );
  XOR U4273 ( .A(n4074), .B(n4075), .Z(n4077) );
  XOR U4274 ( .A(n4076), .B(n4077), .Z(n4105) );
  XOR U4275 ( .A(n4104), .B(n4105), .Z(n4106) );
  XNOR U4276 ( .A(n4107), .B(n4106), .Z(n4152) );
  XOR U4277 ( .A(n4153), .B(n4152), .Z(n4154) );
  XNOR U4278 ( .A(n4155), .B(n4154), .Z(n4041) );
  OR U4279 ( .A(n3934), .B(n3933), .Z(n3938) );
  NAND U4280 ( .A(n3936), .B(n3935), .Z(n3937) );
  NAND U4281 ( .A(n3938), .B(n3937), .Z(n4039) );
  NANDN U4282 ( .A(n3940), .B(n3939), .Z(n3944) );
  NANDN U4283 ( .A(n3942), .B(n3941), .Z(n3943) );
  NAND U4284 ( .A(n3944), .B(n3943), .Z(n4158) );
  NAND U4285 ( .A(n3946), .B(n3945), .Z(n3950) );
  NAND U4286 ( .A(n3948), .B(n3947), .Z(n3949) );
  NAND U4287 ( .A(n3950), .B(n3949), .Z(n4157) );
  NANDN U4288 ( .A(n3952), .B(n3951), .Z(n3956) );
  NAND U4289 ( .A(n3954), .B(n3953), .Z(n3955) );
  NAND U4290 ( .A(n3956), .B(n3955), .Z(n4098) );
  NANDN U4291 ( .A(n3958), .B(n3957), .Z(n3962) );
  NAND U4292 ( .A(n3960), .B(n3959), .Z(n3961) );
  AND U4293 ( .A(n3962), .B(n3961), .Z(n4099) );
  XNOR U4294 ( .A(n4098), .B(n4099), .Z(n4100) );
  NAND U4295 ( .A(n3963), .B(n8286), .Z(n3965) );
  XNOR U4296 ( .A(b[9]), .B(n6914), .Z(n4122) );
  NAND U4297 ( .A(n4122), .B(n8288), .Z(n3964) );
  NAND U4298 ( .A(n3965), .B(n3964), .Z(n4082) );
  NAND U4299 ( .A(n3966), .B(n8961), .Z(n3968) );
  XOR U4300 ( .A(b[15]), .B(a[27]), .Z(n4125) );
  NAND U4301 ( .A(n4125), .B(n8963), .Z(n3967) );
  NAND U4302 ( .A(n3968), .B(n3967), .Z(n4080) );
  XNOR U4303 ( .A(b[21]), .B(a[21]), .Z(n4128) );
  NANDN U4304 ( .A(n4128), .B(n9493), .Z(n3971) );
  NANDN U4305 ( .A(n3969), .B(n9495), .Z(n3970) );
  AND U4306 ( .A(n3971), .B(n3970), .Z(n4081) );
  XOR U4307 ( .A(n4080), .B(n4081), .Z(n4083) );
  XNOR U4308 ( .A(n4082), .B(n4083), .Z(n4071) );
  XNOR U4309 ( .A(b[11]), .B(a[31]), .Z(n4131) );
  NANDN U4310 ( .A(n4131), .B(n8541), .Z(n3974) );
  NANDN U4311 ( .A(n3972), .B(n8542), .Z(n3973) );
  NAND U4312 ( .A(n3974), .B(n3973), .Z(n4069) );
  XNOR U4313 ( .A(b[13]), .B(a[29]), .Z(n4134) );
  NANDN U4314 ( .A(n4134), .B(n8730), .Z(n3977) );
  NANDN U4315 ( .A(n3975), .B(n8731), .Z(n3976) );
  AND U4316 ( .A(n3977), .B(n3976), .Z(n4068) );
  XNOR U4317 ( .A(n4069), .B(n4068), .Z(n4070) );
  XNOR U4318 ( .A(n4071), .B(n4070), .Z(n4088) );
  NANDN U4319 ( .A(n315), .B(a[41]), .Z(n3978) );
  XNOR U4320 ( .A(b[1]), .B(n3978), .Z(n3980) );
  IV U4321 ( .A(a[40]), .Z(n7932) );
  NANDN U4322 ( .A(n7932), .B(n315), .Z(n3979) );
  AND U4323 ( .A(n3980), .B(n3979), .Z(n4046) );
  NAND U4324 ( .A(n3981), .B(n9875), .Z(n3983) );
  XOR U4325 ( .A(n322), .B(n4578), .Z(n4140) );
  NANDN U4326 ( .A(n9874), .B(n4140), .Z(n3982) );
  NAND U4327 ( .A(n3983), .B(n3982), .Z(n4044) );
  NANDN U4328 ( .A(n323), .B(a[9]), .Z(n4045) );
  XNOR U4329 ( .A(n4044), .B(n4045), .Z(n4047) );
  XOR U4330 ( .A(n4046), .B(n4047), .Z(n4086) );
  NANDN U4331 ( .A(n3984), .B(n9622), .Z(n3986) );
  XNOR U4332 ( .A(b[23]), .B(a[19]), .Z(n4143) );
  OR U4333 ( .A(n4143), .B(n9621), .Z(n3985) );
  NAND U4334 ( .A(n3986), .B(n3985), .Z(n4113) );
  XOR U4335 ( .A(b[7]), .B(a[35]), .Z(n4146) );
  NANDN U4336 ( .A(n8013), .B(n4146), .Z(n3989) );
  NAND U4337 ( .A(n3987), .B(n8014), .Z(n3988) );
  NAND U4338 ( .A(n3989), .B(n3988), .Z(n4110) );
  XOR U4339 ( .A(b[25]), .B(n5168), .Z(n4149) );
  NANDN U4340 ( .A(n4149), .B(n9706), .Z(n3992) );
  NANDN U4341 ( .A(n3990), .B(n9707), .Z(n3991) );
  AND U4342 ( .A(n3992), .B(n3991), .Z(n4111) );
  XNOR U4343 ( .A(n4110), .B(n4111), .Z(n4112) );
  XNOR U4344 ( .A(n4113), .B(n4112), .Z(n4087) );
  XOR U4345 ( .A(n4086), .B(n4087), .Z(n4089) );
  XNOR U4346 ( .A(n4088), .B(n4089), .Z(n4101) );
  XNOR U4347 ( .A(n4100), .B(n4101), .Z(n4156) );
  XNOR U4348 ( .A(n4157), .B(n4156), .Z(n4159) );
  XNOR U4349 ( .A(n4158), .B(n4159), .Z(n4038) );
  XNOR U4350 ( .A(n4039), .B(n4038), .Z(n4040) );
  XOR U4351 ( .A(n4041), .B(n4040), .Z(n4035) );
  NANDN U4352 ( .A(n3994), .B(n3993), .Z(n3998) );
  OR U4353 ( .A(n3996), .B(n3995), .Z(n3997) );
  NAND U4354 ( .A(n3998), .B(n3997), .Z(n4032) );
  NAND U4355 ( .A(n4000), .B(n3999), .Z(n4004) );
  NANDN U4356 ( .A(n4002), .B(n4001), .Z(n4003) );
  NAND U4357 ( .A(n4004), .B(n4003), .Z(n4033) );
  XNOR U4358 ( .A(n4032), .B(n4033), .Z(n4034) );
  XNOR U4359 ( .A(n4035), .B(n4034), .Z(n4029) );
  NANDN U4360 ( .A(n4006), .B(n4005), .Z(n4010) );
  NAND U4361 ( .A(n4008), .B(n4007), .Z(n4009) );
  NAND U4362 ( .A(n4010), .B(n4009), .Z(n4026) );
  NANDN U4363 ( .A(n4012), .B(n4011), .Z(n4016) );
  OR U4364 ( .A(n4014), .B(n4013), .Z(n4015) );
  NAND U4365 ( .A(n4016), .B(n4015), .Z(n4027) );
  XNOR U4366 ( .A(n4026), .B(n4027), .Z(n4028) );
  XNOR U4367 ( .A(n4029), .B(n4028), .Z(n4022) );
  XOR U4368 ( .A(n4023), .B(n4022), .Z(n4024) );
  XNOR U4369 ( .A(n4025), .B(n4024), .Z(n4162) );
  XNOR U4370 ( .A(n4162), .B(sreg[73]), .Z(n4164) );
  NAND U4371 ( .A(n4017), .B(sreg[72]), .Z(n4021) );
  OR U4372 ( .A(n4019), .B(n4018), .Z(n4020) );
  AND U4373 ( .A(n4021), .B(n4020), .Z(n4163) );
  XOR U4374 ( .A(n4164), .B(n4163), .Z(c[73]) );
  NANDN U4375 ( .A(n4027), .B(n4026), .Z(n4031) );
  NANDN U4376 ( .A(n4029), .B(n4028), .Z(n4030) );
  NAND U4377 ( .A(n4031), .B(n4030), .Z(n4168) );
  NANDN U4378 ( .A(n4033), .B(n4032), .Z(n4037) );
  NAND U4379 ( .A(n4035), .B(n4034), .Z(n4036) );
  NAND U4380 ( .A(n4037), .B(n4036), .Z(n4173) );
  NANDN U4381 ( .A(n4039), .B(n4038), .Z(n4043) );
  NANDN U4382 ( .A(n4041), .B(n4040), .Z(n4042) );
  NAND U4383 ( .A(n4043), .B(n4042), .Z(n4174) );
  XNOR U4384 ( .A(n4173), .B(n4174), .Z(n4175) );
  NANDN U4385 ( .A(n4045), .B(n4044), .Z(n4049) );
  NAND U4386 ( .A(n4047), .B(n4046), .Z(n4048) );
  NAND U4387 ( .A(n4049), .B(n4048), .Z(n4242) );
  NAND U4388 ( .A(n4050), .B(n9379), .Z(n4052) );
  XNOR U4389 ( .A(n9562), .B(a[24]), .Z(n4209) );
  NAND U4390 ( .A(n4209), .B(n9378), .Z(n4051) );
  NAND U4391 ( .A(n4052), .B(n4051), .Z(n4253) );
  NANDN U4392 ( .A(n4053), .B(n9801), .Z(n4055) );
  XNOR U4393 ( .A(b[27]), .B(a[16]), .Z(n4212) );
  OR U4394 ( .A(n4212), .B(n9751), .Z(n4054) );
  NAND U4395 ( .A(n4055), .B(n4054), .Z(n4251) );
  XOR U4396 ( .A(b[5]), .B(n7672), .Z(n4215) );
  NANDN U4397 ( .A(n4215), .B(n7905), .Z(n4058) );
  NANDN U4398 ( .A(n4056), .B(n7906), .Z(n4057) );
  AND U4399 ( .A(n4058), .B(n4057), .Z(n4252) );
  XNOR U4400 ( .A(n4251), .B(n4252), .Z(n4254) );
  XOR U4401 ( .A(n4253), .B(n4254), .Z(n4239) );
  NAND U4402 ( .A(n4059), .B(n9105), .Z(n4061) );
  XNOR U4403 ( .A(n9455), .B(a[26]), .Z(n4218) );
  NAND U4404 ( .A(n4218), .B(n9107), .Z(n4060) );
  AND U4405 ( .A(n4061), .B(n4060), .Z(n4194) );
  NAND U4406 ( .A(n4062), .B(n9914), .Z(n4064) );
  XNOR U4407 ( .A(n323), .B(a[12]), .Z(n4221) );
  NANDN U4408 ( .A(n9913), .B(n4221), .Z(n4063) );
  AND U4409 ( .A(n4064), .B(n4063), .Z(n4192) );
  NAND U4410 ( .A(n4065), .B(n7622), .Z(n4067) );
  XNOR U4411 ( .A(n7932), .B(b[3]), .Z(n4224) );
  NAND U4412 ( .A(n4224), .B(n7620), .Z(n4066) );
  NAND U4413 ( .A(n4067), .B(n4066), .Z(n4191) );
  XOR U4414 ( .A(n4239), .B(n4240), .Z(n4241) );
  XNOR U4415 ( .A(n4242), .B(n4241), .Z(n4287) );
  NANDN U4416 ( .A(n4069), .B(n4068), .Z(n4073) );
  NANDN U4417 ( .A(n4071), .B(n4070), .Z(n4072) );
  NAND U4418 ( .A(n4073), .B(n4072), .Z(n4230) );
  NAND U4419 ( .A(n4075), .B(n4074), .Z(n4079) );
  NAND U4420 ( .A(n4077), .B(n4076), .Z(n4078) );
  NAND U4421 ( .A(n4079), .B(n4078), .Z(n4228) );
  NANDN U4422 ( .A(n4081), .B(n4080), .Z(n4085) );
  NANDN U4423 ( .A(n4083), .B(n4082), .Z(n4084) );
  NAND U4424 ( .A(n4085), .B(n4084), .Z(n4227) );
  XNOR U4425 ( .A(n4230), .B(n4229), .Z(n4288) );
  XOR U4426 ( .A(n4287), .B(n4288), .Z(n4290) );
  NANDN U4427 ( .A(n4087), .B(n4086), .Z(n4091) );
  OR U4428 ( .A(n4089), .B(n4088), .Z(n4090) );
  NAND U4429 ( .A(n4091), .B(n4090), .Z(n4289) );
  XOR U4430 ( .A(n4290), .B(n4289), .Z(n4307) );
  OR U4431 ( .A(n4093), .B(n4092), .Z(n4097) );
  NANDN U4432 ( .A(n4095), .B(n4094), .Z(n4096) );
  NAND U4433 ( .A(n4097), .B(n4096), .Z(n4306) );
  NANDN U4434 ( .A(n4099), .B(n4098), .Z(n4103) );
  NANDN U4435 ( .A(n4101), .B(n4100), .Z(n4102) );
  NAND U4436 ( .A(n4103), .B(n4102), .Z(n4295) );
  NAND U4437 ( .A(n4105), .B(n4104), .Z(n4109) );
  NANDN U4438 ( .A(n4107), .B(n4106), .Z(n4108) );
  NAND U4439 ( .A(n4109), .B(n4108), .Z(n4294) );
  NANDN U4440 ( .A(n4111), .B(n4110), .Z(n4115) );
  NAND U4441 ( .A(n4113), .B(n4112), .Z(n4114) );
  NAND U4442 ( .A(n4115), .B(n4114), .Z(n4233) );
  NANDN U4443 ( .A(n4117), .B(n4116), .Z(n4121) );
  NAND U4444 ( .A(n4119), .B(n4118), .Z(n4120) );
  AND U4445 ( .A(n4121), .B(n4120), .Z(n4234) );
  XNOR U4446 ( .A(n4233), .B(n4234), .Z(n4235) );
  NAND U4447 ( .A(n4122), .B(n8286), .Z(n4124) );
  XOR U4448 ( .A(b[9]), .B(a[34]), .Z(n4257) );
  NAND U4449 ( .A(n4257), .B(n8288), .Z(n4123) );
  NAND U4450 ( .A(n4124), .B(n4123), .Z(n4199) );
  NAND U4451 ( .A(n4125), .B(n8961), .Z(n4127) );
  XOR U4452 ( .A(b[15]), .B(a[28]), .Z(n4260) );
  NAND U4453 ( .A(n4260), .B(n8963), .Z(n4126) );
  NAND U4454 ( .A(n4127), .B(n4126), .Z(n4197) );
  XNOR U4455 ( .A(b[21]), .B(a[22]), .Z(n4263) );
  NANDN U4456 ( .A(n4263), .B(n9493), .Z(n4130) );
  NANDN U4457 ( .A(n4128), .B(n9495), .Z(n4129) );
  AND U4458 ( .A(n4130), .B(n4129), .Z(n4198) );
  XOR U4459 ( .A(n4197), .B(n4198), .Z(n4200) );
  XNOR U4460 ( .A(n4199), .B(n4200), .Z(n4188) );
  XNOR U4461 ( .A(b[11]), .B(a[32]), .Z(n4266) );
  NANDN U4462 ( .A(n4266), .B(n8541), .Z(n4133) );
  NANDN U4463 ( .A(n4131), .B(n8542), .Z(n4132) );
  NAND U4464 ( .A(n4133), .B(n4132), .Z(n4186) );
  XOR U4465 ( .A(b[13]), .B(n6135), .Z(n4269) );
  NANDN U4466 ( .A(n4269), .B(n8730), .Z(n4136) );
  NANDN U4467 ( .A(n4134), .B(n8731), .Z(n4135) );
  NAND U4468 ( .A(n4136), .B(n4135), .Z(n4185) );
  XNOR U4469 ( .A(n4188), .B(n4187), .Z(n4182) );
  NANDN U4470 ( .A(n315), .B(a[42]), .Z(n4137) );
  XNOR U4471 ( .A(b[1]), .B(n4137), .Z(n4139) );
  NANDN U4472 ( .A(b[0]), .B(a[41]), .Z(n4138) );
  AND U4473 ( .A(n4139), .B(n4138), .Z(n4205) );
  NAND U4474 ( .A(n9875), .B(n4140), .Z(n4142) );
  XNOR U4475 ( .A(n322), .B(a[14]), .Z(n4275) );
  NANDN U4476 ( .A(n9874), .B(n4275), .Z(n4141) );
  NAND U4477 ( .A(n4142), .B(n4141), .Z(n4203) );
  NANDN U4478 ( .A(n323), .B(a[10]), .Z(n4204) );
  XNOR U4479 ( .A(n4203), .B(n4204), .Z(n4206) );
  XNOR U4480 ( .A(n4205), .B(n4206), .Z(n4180) );
  NANDN U4481 ( .A(n4143), .B(n9622), .Z(n4145) );
  XNOR U4482 ( .A(b[23]), .B(a[20]), .Z(n4278) );
  OR U4483 ( .A(n4278), .B(n9621), .Z(n4144) );
  NAND U4484 ( .A(n4145), .B(n4144), .Z(n4248) );
  XNOR U4485 ( .A(b[7]), .B(a[36]), .Z(n4281) );
  OR U4486 ( .A(n4281), .B(n8013), .Z(n4148) );
  NAND U4487 ( .A(n4146), .B(n8014), .Z(n4147) );
  NAND U4488 ( .A(n4148), .B(n4147), .Z(n4245) );
  XNOR U4489 ( .A(b[25]), .B(a[18]), .Z(n4284) );
  NANDN U4490 ( .A(n4284), .B(n9706), .Z(n4151) );
  NANDN U4491 ( .A(n4149), .B(n9707), .Z(n4150) );
  AND U4492 ( .A(n4151), .B(n4150), .Z(n4246) );
  XNOR U4493 ( .A(n4245), .B(n4246), .Z(n4247) );
  XOR U4494 ( .A(n4248), .B(n4247), .Z(n4179) );
  XOR U4495 ( .A(n4182), .B(n4181), .Z(n4236) );
  XNOR U4496 ( .A(n4235), .B(n4236), .Z(n4293) );
  XNOR U4497 ( .A(n4294), .B(n4293), .Z(n4296) );
  XNOR U4498 ( .A(n4295), .B(n4296), .Z(n4305) );
  XOR U4499 ( .A(n4306), .B(n4305), .Z(n4308) );
  NAND U4500 ( .A(n4157), .B(n4156), .Z(n4161) );
  NANDN U4501 ( .A(n4159), .B(n4158), .Z(n4160) );
  AND U4502 ( .A(n4161), .B(n4160), .Z(n4299) );
  XNOR U4503 ( .A(n4300), .B(n4299), .Z(n4301) );
  XOR U4504 ( .A(n4302), .B(n4301), .Z(n4176) );
  XOR U4505 ( .A(n4175), .B(n4176), .Z(n4167) );
  XOR U4506 ( .A(n4168), .B(n4167), .Z(n4169) );
  XNOR U4507 ( .A(n4170), .B(n4169), .Z(n4311) );
  XNOR U4508 ( .A(n4311), .B(sreg[74]), .Z(n4313) );
  NAND U4509 ( .A(n4162), .B(sreg[73]), .Z(n4166) );
  OR U4510 ( .A(n4164), .B(n4163), .Z(n4165) );
  AND U4511 ( .A(n4166), .B(n4165), .Z(n4312) );
  XOR U4512 ( .A(n4313), .B(n4312), .Z(c[74]) );
  NAND U4513 ( .A(n4168), .B(n4167), .Z(n4172) );
  NAND U4514 ( .A(n4170), .B(n4169), .Z(n4171) );
  NAND U4515 ( .A(n4172), .B(n4171), .Z(n4319) );
  NANDN U4516 ( .A(n4174), .B(n4173), .Z(n4178) );
  NAND U4517 ( .A(n4176), .B(n4175), .Z(n4177) );
  NAND U4518 ( .A(n4178), .B(n4177), .Z(n4317) );
  NANDN U4519 ( .A(n4180), .B(n4179), .Z(n4184) );
  NANDN U4520 ( .A(n4182), .B(n4181), .Z(n4183) );
  NAND U4521 ( .A(n4184), .B(n4183), .Z(n4437) );
  OR U4522 ( .A(n4186), .B(n4185), .Z(n4190) );
  NANDN U4523 ( .A(n4188), .B(n4187), .Z(n4189) );
  NAND U4524 ( .A(n4190), .B(n4189), .Z(n4376) );
  NANDN U4525 ( .A(n4192), .B(n4191), .Z(n4196) );
  NANDN U4526 ( .A(n4194), .B(n4193), .Z(n4195) );
  NAND U4527 ( .A(n4196), .B(n4195), .Z(n4375) );
  NANDN U4528 ( .A(n4198), .B(n4197), .Z(n4202) );
  NANDN U4529 ( .A(n4200), .B(n4199), .Z(n4201) );
  NAND U4530 ( .A(n4202), .B(n4201), .Z(n4374) );
  XOR U4531 ( .A(n4376), .B(n4377), .Z(n4434) );
  NANDN U4532 ( .A(n4204), .B(n4203), .Z(n4208) );
  NAND U4533 ( .A(n4206), .B(n4205), .Z(n4207) );
  NAND U4534 ( .A(n4208), .B(n4207), .Z(n4389) );
  NAND U4535 ( .A(n4209), .B(n9379), .Z(n4211) );
  XNOR U4536 ( .A(n9562), .B(a[25]), .Z(n4356) );
  NAND U4537 ( .A(n4356), .B(n9378), .Z(n4210) );
  NAND U4538 ( .A(n4211), .B(n4210), .Z(n4400) );
  NANDN U4539 ( .A(n4212), .B(n9801), .Z(n4214) );
  XOR U4540 ( .A(b[27]), .B(n5168), .Z(n4359) );
  OR U4541 ( .A(n4359), .B(n9751), .Z(n4213) );
  NAND U4542 ( .A(n4214), .B(n4213), .Z(n4398) );
  XNOR U4543 ( .A(b[5]), .B(a[39]), .Z(n4362) );
  NANDN U4544 ( .A(n4362), .B(n7905), .Z(n4217) );
  NANDN U4545 ( .A(n4215), .B(n7906), .Z(n4216) );
  AND U4546 ( .A(n4217), .B(n4216), .Z(n4399) );
  XNOR U4547 ( .A(n4398), .B(n4399), .Z(n4401) );
  XOR U4548 ( .A(n4400), .B(n4401), .Z(n4386) );
  NAND U4549 ( .A(n4218), .B(n9105), .Z(n4220) );
  XNOR U4550 ( .A(n9455), .B(a[27]), .Z(n4365) );
  NAND U4551 ( .A(n4365), .B(n9107), .Z(n4219) );
  AND U4552 ( .A(n4220), .B(n4219), .Z(n4341) );
  NAND U4553 ( .A(n4221), .B(n9914), .Z(n4223) );
  XNOR U4554 ( .A(n323), .B(a[13]), .Z(n4368) );
  NANDN U4555 ( .A(n9913), .B(n4368), .Z(n4222) );
  AND U4556 ( .A(n4223), .B(n4222), .Z(n4339) );
  NAND U4557 ( .A(n4224), .B(n7622), .Z(n4226) );
  XNOR U4558 ( .A(a[41]), .B(n316), .Z(n4371) );
  NAND U4559 ( .A(n4371), .B(n7620), .Z(n4225) );
  NAND U4560 ( .A(n4226), .B(n4225), .Z(n4338) );
  XOR U4561 ( .A(n4386), .B(n4387), .Z(n4388) );
  XNOR U4562 ( .A(n4389), .B(n4388), .Z(n4435) );
  XNOR U4563 ( .A(n4434), .B(n4435), .Z(n4436) );
  XNOR U4564 ( .A(n4437), .B(n4436), .Z(n4455) );
  OR U4565 ( .A(n4228), .B(n4227), .Z(n4232) );
  NAND U4566 ( .A(n4230), .B(n4229), .Z(n4231) );
  NAND U4567 ( .A(n4232), .B(n4231), .Z(n4453) );
  NANDN U4568 ( .A(n4234), .B(n4233), .Z(n4238) );
  NANDN U4569 ( .A(n4236), .B(n4235), .Z(n4237) );
  NAND U4570 ( .A(n4238), .B(n4237), .Z(n4442) );
  NAND U4571 ( .A(n4240), .B(n4239), .Z(n4244) );
  NAND U4572 ( .A(n4242), .B(n4241), .Z(n4243) );
  NAND U4573 ( .A(n4244), .B(n4243), .Z(n4441) );
  NANDN U4574 ( .A(n4246), .B(n4245), .Z(n4250) );
  NAND U4575 ( .A(n4248), .B(n4247), .Z(n4249) );
  NAND U4576 ( .A(n4250), .B(n4249), .Z(n4380) );
  NANDN U4577 ( .A(n4252), .B(n4251), .Z(n4256) );
  NAND U4578 ( .A(n4254), .B(n4253), .Z(n4255) );
  AND U4579 ( .A(n4256), .B(n4255), .Z(n4381) );
  XNOR U4580 ( .A(n4380), .B(n4381), .Z(n4382) );
  NAND U4581 ( .A(n4257), .B(n8286), .Z(n4259) );
  XOR U4582 ( .A(b[9]), .B(a[35]), .Z(n4404) );
  NAND U4583 ( .A(n4404), .B(n8288), .Z(n4258) );
  NAND U4584 ( .A(n4259), .B(n4258), .Z(n4346) );
  NAND U4585 ( .A(n4260), .B(n8961), .Z(n4262) );
  XOR U4586 ( .A(b[15]), .B(a[29]), .Z(n4407) );
  NAND U4587 ( .A(n4407), .B(n8963), .Z(n4261) );
  NAND U4588 ( .A(n4262), .B(n4261), .Z(n4344) );
  XOR U4589 ( .A(b[21]), .B(n6044), .Z(n4410) );
  NANDN U4590 ( .A(n4410), .B(n9493), .Z(n4265) );
  NANDN U4591 ( .A(n4263), .B(n9495), .Z(n4264) );
  AND U4592 ( .A(n4265), .B(n4264), .Z(n4345) );
  XOR U4593 ( .A(n4344), .B(n4345), .Z(n4347) );
  XNOR U4594 ( .A(n4346), .B(n4347), .Z(n4335) );
  XOR U4595 ( .A(b[11]), .B(n6914), .Z(n4413) );
  NANDN U4596 ( .A(n4413), .B(n8541), .Z(n4268) );
  NANDN U4597 ( .A(n4266), .B(n8542), .Z(n4267) );
  NAND U4598 ( .A(n4268), .B(n4267), .Z(n4333) );
  XNOR U4599 ( .A(b[13]), .B(a[31]), .Z(n4416) );
  NANDN U4600 ( .A(n4416), .B(n8730), .Z(n4271) );
  NANDN U4601 ( .A(n4269), .B(n8731), .Z(n4270) );
  NAND U4602 ( .A(n4271), .B(n4270), .Z(n4332) );
  XNOR U4603 ( .A(n4335), .B(n4334), .Z(n4329) );
  NANDN U4604 ( .A(n315), .B(a[43]), .Z(n4272) );
  XNOR U4605 ( .A(b[1]), .B(n4272), .Z(n4274) );
  IV U4606 ( .A(a[42]), .Z(n8156) );
  NANDN U4607 ( .A(n8156), .B(n315), .Z(n4273) );
  AND U4608 ( .A(n4274), .B(n4273), .Z(n4352) );
  NAND U4609 ( .A(n9875), .B(n4275), .Z(n4277) );
  XNOR U4610 ( .A(n322), .B(a[15]), .Z(n4419) );
  NANDN U4611 ( .A(n9874), .B(n4419), .Z(n4276) );
  NAND U4612 ( .A(n4277), .B(n4276), .Z(n4350) );
  NANDN U4613 ( .A(n323), .B(a[11]), .Z(n4351) );
  XNOR U4614 ( .A(n4350), .B(n4351), .Z(n4353) );
  XNOR U4615 ( .A(n4352), .B(n4353), .Z(n4327) );
  NANDN U4616 ( .A(n4278), .B(n9622), .Z(n4280) );
  XNOR U4617 ( .A(b[23]), .B(a[21]), .Z(n4425) );
  OR U4618 ( .A(n4425), .B(n9621), .Z(n4279) );
  NAND U4619 ( .A(n4280), .B(n4279), .Z(n4395) );
  XOR U4620 ( .A(b[7]), .B(a[37]), .Z(n4428) );
  NANDN U4621 ( .A(n8013), .B(n4428), .Z(n4283) );
  NANDN U4622 ( .A(n4281), .B(n8014), .Z(n4282) );
  NAND U4623 ( .A(n4283), .B(n4282), .Z(n4392) );
  XNOR U4624 ( .A(b[25]), .B(a[19]), .Z(n4431) );
  NANDN U4625 ( .A(n4431), .B(n9706), .Z(n4286) );
  NANDN U4626 ( .A(n4284), .B(n9707), .Z(n4285) );
  AND U4627 ( .A(n4286), .B(n4285), .Z(n4393) );
  XNOR U4628 ( .A(n4392), .B(n4393), .Z(n4394) );
  XOR U4629 ( .A(n4395), .B(n4394), .Z(n4326) );
  XOR U4630 ( .A(n4329), .B(n4328), .Z(n4383) );
  XNOR U4631 ( .A(n4382), .B(n4383), .Z(n4440) );
  XNOR U4632 ( .A(n4441), .B(n4440), .Z(n4443) );
  XNOR U4633 ( .A(n4442), .B(n4443), .Z(n4452) );
  XNOR U4634 ( .A(n4453), .B(n4452), .Z(n4454) );
  XOR U4635 ( .A(n4455), .B(n4454), .Z(n4449) );
  NANDN U4636 ( .A(n4288), .B(n4287), .Z(n4292) );
  OR U4637 ( .A(n4290), .B(n4289), .Z(n4291) );
  NAND U4638 ( .A(n4292), .B(n4291), .Z(n4446) );
  NAND U4639 ( .A(n4294), .B(n4293), .Z(n4298) );
  NANDN U4640 ( .A(n4296), .B(n4295), .Z(n4297) );
  NAND U4641 ( .A(n4298), .B(n4297), .Z(n4447) );
  XNOR U4642 ( .A(n4446), .B(n4447), .Z(n4448) );
  XNOR U4643 ( .A(n4449), .B(n4448), .Z(n4323) );
  NANDN U4644 ( .A(n4300), .B(n4299), .Z(n4304) );
  NAND U4645 ( .A(n4302), .B(n4301), .Z(n4303) );
  NAND U4646 ( .A(n4304), .B(n4303), .Z(n4320) );
  NANDN U4647 ( .A(n4306), .B(n4305), .Z(n4310) );
  OR U4648 ( .A(n4308), .B(n4307), .Z(n4309) );
  NAND U4649 ( .A(n4310), .B(n4309), .Z(n4321) );
  XNOR U4650 ( .A(n4320), .B(n4321), .Z(n4322) );
  XNOR U4651 ( .A(n4323), .B(n4322), .Z(n4316) );
  XOR U4652 ( .A(n4317), .B(n4316), .Z(n4318) );
  XNOR U4653 ( .A(n4319), .B(n4318), .Z(n4458) );
  XNOR U4654 ( .A(n4458), .B(sreg[75]), .Z(n4460) );
  NAND U4655 ( .A(n4311), .B(sreg[74]), .Z(n4315) );
  OR U4656 ( .A(n4313), .B(n4312), .Z(n4314) );
  AND U4657 ( .A(n4315), .B(n4314), .Z(n4459) );
  XOR U4658 ( .A(n4460), .B(n4459), .Z(c[75]) );
  NANDN U4659 ( .A(n4321), .B(n4320), .Z(n4325) );
  NANDN U4660 ( .A(n4323), .B(n4322), .Z(n4324) );
  NAND U4661 ( .A(n4325), .B(n4324), .Z(n4464) );
  NANDN U4662 ( .A(n4327), .B(n4326), .Z(n4331) );
  NANDN U4663 ( .A(n4329), .B(n4328), .Z(n4330) );
  NAND U4664 ( .A(n4331), .B(n4330), .Z(n4597) );
  OR U4665 ( .A(n4333), .B(n4332), .Z(n4337) );
  NANDN U4666 ( .A(n4335), .B(n4334), .Z(n4336) );
  NAND U4667 ( .A(n4337), .B(n4336), .Z(n4535) );
  NANDN U4668 ( .A(n4339), .B(n4338), .Z(n4343) );
  NANDN U4669 ( .A(n4341), .B(n4340), .Z(n4342) );
  NAND U4670 ( .A(n4343), .B(n4342), .Z(n4534) );
  NANDN U4671 ( .A(n4345), .B(n4344), .Z(n4349) );
  NANDN U4672 ( .A(n4347), .B(n4346), .Z(n4348) );
  NAND U4673 ( .A(n4349), .B(n4348), .Z(n4533) );
  XOR U4674 ( .A(n4535), .B(n4536), .Z(n4594) );
  NANDN U4675 ( .A(n4351), .B(n4350), .Z(n4355) );
  NAND U4676 ( .A(n4353), .B(n4352), .Z(n4354) );
  NAND U4677 ( .A(n4355), .B(n4354), .Z(n4548) );
  NAND U4678 ( .A(n4356), .B(n9379), .Z(n4358) );
  XNOR U4679 ( .A(n9562), .B(a[26]), .Z(n4491) );
  NAND U4680 ( .A(n4491), .B(n9378), .Z(n4357) );
  NAND U4681 ( .A(n4358), .B(n4357), .Z(n4559) );
  NANDN U4682 ( .A(n4359), .B(n9801), .Z(n4361) );
  XNOR U4683 ( .A(b[27]), .B(a[18]), .Z(n4494) );
  OR U4684 ( .A(n4494), .B(n9751), .Z(n4360) );
  NAND U4685 ( .A(n4361), .B(n4360), .Z(n4557) );
  XOR U4686 ( .A(a[40]), .B(n317), .Z(n4497) );
  NANDN U4687 ( .A(n4497), .B(n7905), .Z(n4364) );
  NANDN U4688 ( .A(n4362), .B(n7906), .Z(n4363) );
  AND U4689 ( .A(n4364), .B(n4363), .Z(n4558) );
  XNOR U4690 ( .A(n4557), .B(n4558), .Z(n4560) );
  XOR U4691 ( .A(n4559), .B(n4560), .Z(n4545) );
  NAND U4692 ( .A(n4365), .B(n9105), .Z(n4367) );
  XNOR U4693 ( .A(n9455), .B(a[28]), .Z(n4500) );
  NAND U4694 ( .A(n4500), .B(n9107), .Z(n4366) );
  NAND U4695 ( .A(n4367), .B(n4366), .Z(n4517) );
  NAND U4696 ( .A(n4368), .B(n9914), .Z(n4370) );
  XNOR U4697 ( .A(n323), .B(a[14]), .Z(n4503) );
  NANDN U4698 ( .A(n9913), .B(n4503), .Z(n4369) );
  NAND U4699 ( .A(n4370), .B(n4369), .Z(n4515) );
  NAND U4700 ( .A(n4371), .B(n7622), .Z(n4373) );
  XNOR U4701 ( .A(n8156), .B(b[3]), .Z(n4506) );
  NAND U4702 ( .A(n4506), .B(n7620), .Z(n4372) );
  NAND U4703 ( .A(n4373), .B(n4372), .Z(n4516) );
  XOR U4704 ( .A(n4515), .B(n4516), .Z(n4518) );
  XOR U4705 ( .A(n4517), .B(n4518), .Z(n4546) );
  XOR U4706 ( .A(n4545), .B(n4546), .Z(n4547) );
  XNOR U4707 ( .A(n4548), .B(n4547), .Z(n4595) );
  XNOR U4708 ( .A(n4594), .B(n4595), .Z(n4596) );
  XNOR U4709 ( .A(n4597), .B(n4596), .Z(n4482) );
  OR U4710 ( .A(n4375), .B(n4374), .Z(n4379) );
  NANDN U4711 ( .A(n4377), .B(n4376), .Z(n4378) );
  NAND U4712 ( .A(n4379), .B(n4378), .Z(n4480) );
  NANDN U4713 ( .A(n4381), .B(n4380), .Z(n4385) );
  NANDN U4714 ( .A(n4383), .B(n4382), .Z(n4384) );
  NAND U4715 ( .A(n4385), .B(n4384), .Z(n4602) );
  NAND U4716 ( .A(n4387), .B(n4386), .Z(n4391) );
  NAND U4717 ( .A(n4389), .B(n4388), .Z(n4390) );
  NAND U4718 ( .A(n4391), .B(n4390), .Z(n4601) );
  NANDN U4719 ( .A(n4393), .B(n4392), .Z(n4397) );
  NAND U4720 ( .A(n4395), .B(n4394), .Z(n4396) );
  NAND U4721 ( .A(n4397), .B(n4396), .Z(n4539) );
  NANDN U4722 ( .A(n4399), .B(n4398), .Z(n4403) );
  NAND U4723 ( .A(n4401), .B(n4400), .Z(n4402) );
  AND U4724 ( .A(n4403), .B(n4402), .Z(n4540) );
  XNOR U4725 ( .A(n4539), .B(n4540), .Z(n4541) );
  NAND U4726 ( .A(n4404), .B(n8286), .Z(n4406) );
  XNOR U4727 ( .A(b[9]), .B(n7293), .Z(n4563) );
  NAND U4728 ( .A(n4563), .B(n8288), .Z(n4405) );
  NAND U4729 ( .A(n4406), .B(n4405), .Z(n4523) );
  NAND U4730 ( .A(n4407), .B(n8961), .Z(n4409) );
  XNOR U4731 ( .A(b[15]), .B(n6135), .Z(n4566) );
  NAND U4732 ( .A(n4566), .B(n8963), .Z(n4408) );
  NAND U4733 ( .A(n4409), .B(n4408), .Z(n4521) );
  XNOR U4734 ( .A(b[21]), .B(a[24]), .Z(n4569) );
  NANDN U4735 ( .A(n4569), .B(n9493), .Z(n4412) );
  NANDN U4736 ( .A(n4410), .B(n9495), .Z(n4411) );
  AND U4737 ( .A(n4412), .B(n4411), .Z(n4522) );
  XOR U4738 ( .A(n4521), .B(n4522), .Z(n4524) );
  XNOR U4739 ( .A(n4523), .B(n4524), .Z(n4512) );
  XNOR U4740 ( .A(b[11]), .B(a[34]), .Z(n4572) );
  NANDN U4741 ( .A(n4572), .B(n8541), .Z(n4415) );
  NANDN U4742 ( .A(n4413), .B(n8542), .Z(n4414) );
  NAND U4743 ( .A(n4415), .B(n4414), .Z(n4510) );
  XNOR U4744 ( .A(b[13]), .B(a[32]), .Z(n4575) );
  NANDN U4745 ( .A(n4575), .B(n8730), .Z(n4418) );
  NANDN U4746 ( .A(n4416), .B(n8731), .Z(n4417) );
  AND U4747 ( .A(n4418), .B(n4417), .Z(n4509) );
  XNOR U4748 ( .A(n4510), .B(n4509), .Z(n4511) );
  XNOR U4749 ( .A(n4512), .B(n4511), .Z(n4529) );
  NAND U4750 ( .A(n9875), .B(n4419), .Z(n4421) );
  XNOR U4751 ( .A(b[29]), .B(a[16]), .Z(n4579) );
  OR U4752 ( .A(n4579), .B(n9874), .Z(n4420) );
  NAND U4753 ( .A(n4421), .B(n4420), .Z(n4485) );
  NANDN U4754 ( .A(n323), .B(a[12]), .Z(n4486) );
  XNOR U4755 ( .A(n4485), .B(n4486), .Z(n4488) );
  NANDN U4756 ( .A(n315), .B(a[44]), .Z(n4422) );
  XNOR U4757 ( .A(b[1]), .B(n4422), .Z(n4424) );
  NANDN U4758 ( .A(b[0]), .B(a[43]), .Z(n4423) );
  AND U4759 ( .A(n4424), .B(n4423), .Z(n4487) );
  XOR U4760 ( .A(n4488), .B(n4487), .Z(n4527) );
  NANDN U4761 ( .A(n4425), .B(n9622), .Z(n4427) );
  XNOR U4762 ( .A(b[23]), .B(a[22]), .Z(n4585) );
  OR U4763 ( .A(n4585), .B(n9621), .Z(n4426) );
  NAND U4764 ( .A(n4427), .B(n4426), .Z(n4554) );
  XNOR U4765 ( .A(b[7]), .B(a[38]), .Z(n4588) );
  OR U4766 ( .A(n4588), .B(n8013), .Z(n4430) );
  NAND U4767 ( .A(n4428), .B(n8014), .Z(n4429) );
  NAND U4768 ( .A(n4430), .B(n4429), .Z(n4551) );
  XNOR U4769 ( .A(b[25]), .B(a[20]), .Z(n4591) );
  NANDN U4770 ( .A(n4591), .B(n9706), .Z(n4433) );
  NANDN U4771 ( .A(n4431), .B(n9707), .Z(n4432) );
  AND U4772 ( .A(n4433), .B(n4432), .Z(n4552) );
  XNOR U4773 ( .A(n4551), .B(n4552), .Z(n4553) );
  XNOR U4774 ( .A(n4554), .B(n4553), .Z(n4528) );
  XOR U4775 ( .A(n4527), .B(n4528), .Z(n4530) );
  XNOR U4776 ( .A(n4529), .B(n4530), .Z(n4542) );
  XNOR U4777 ( .A(n4541), .B(n4542), .Z(n4600) );
  XNOR U4778 ( .A(n4601), .B(n4600), .Z(n4603) );
  XNOR U4779 ( .A(n4602), .B(n4603), .Z(n4479) );
  XNOR U4780 ( .A(n4480), .B(n4479), .Z(n4481) );
  XOR U4781 ( .A(n4482), .B(n4481), .Z(n4476) );
  NANDN U4782 ( .A(n4435), .B(n4434), .Z(n4439) );
  NAND U4783 ( .A(n4437), .B(n4436), .Z(n4438) );
  NAND U4784 ( .A(n4439), .B(n4438), .Z(n4474) );
  NAND U4785 ( .A(n4441), .B(n4440), .Z(n4445) );
  NANDN U4786 ( .A(n4443), .B(n4442), .Z(n4444) );
  AND U4787 ( .A(n4445), .B(n4444), .Z(n4473) );
  XNOR U4788 ( .A(n4474), .B(n4473), .Z(n4475) );
  XNOR U4789 ( .A(n4476), .B(n4475), .Z(n4470) );
  NANDN U4790 ( .A(n4447), .B(n4446), .Z(n4451) );
  NAND U4791 ( .A(n4449), .B(n4448), .Z(n4450) );
  NAND U4792 ( .A(n4451), .B(n4450), .Z(n4467) );
  NANDN U4793 ( .A(n4453), .B(n4452), .Z(n4457) );
  NANDN U4794 ( .A(n4455), .B(n4454), .Z(n4456) );
  NAND U4795 ( .A(n4457), .B(n4456), .Z(n4468) );
  XNOR U4796 ( .A(n4467), .B(n4468), .Z(n4469) );
  XNOR U4797 ( .A(n4470), .B(n4469), .Z(n4463) );
  XOR U4798 ( .A(n4464), .B(n4463), .Z(n4465) );
  XNOR U4799 ( .A(n4466), .B(n4465), .Z(n4606) );
  XNOR U4800 ( .A(n4606), .B(sreg[76]), .Z(n4608) );
  NAND U4801 ( .A(n4458), .B(sreg[75]), .Z(n4462) );
  OR U4802 ( .A(n4460), .B(n4459), .Z(n4461) );
  AND U4803 ( .A(n4462), .B(n4461), .Z(n4607) );
  XOR U4804 ( .A(n4608), .B(n4607), .Z(c[76]) );
  NANDN U4805 ( .A(n4468), .B(n4467), .Z(n4472) );
  NANDN U4806 ( .A(n4470), .B(n4469), .Z(n4471) );
  NAND U4807 ( .A(n4472), .B(n4471), .Z(n4612) );
  NANDN U4808 ( .A(n4474), .B(n4473), .Z(n4478) );
  NAND U4809 ( .A(n4476), .B(n4475), .Z(n4477) );
  NAND U4810 ( .A(n4478), .B(n4477), .Z(n4617) );
  NANDN U4811 ( .A(n4480), .B(n4479), .Z(n4484) );
  NANDN U4812 ( .A(n4482), .B(n4481), .Z(n4483) );
  NAND U4813 ( .A(n4484), .B(n4483), .Z(n4618) );
  XNOR U4814 ( .A(n4617), .B(n4618), .Z(n4619) );
  NANDN U4815 ( .A(n4486), .B(n4485), .Z(n4490) );
  NAND U4816 ( .A(n4488), .B(n4487), .Z(n4489) );
  NAND U4817 ( .A(n4490), .B(n4489), .Z(n4686) );
  NAND U4818 ( .A(n4491), .B(n9379), .Z(n4493) );
  XNOR U4819 ( .A(n9562), .B(a[27]), .Z(n4653) );
  NAND U4820 ( .A(n4653), .B(n9378), .Z(n4492) );
  NAND U4821 ( .A(n4493), .B(n4492), .Z(n4697) );
  NANDN U4822 ( .A(n4494), .B(n9801), .Z(n4496) );
  XNOR U4823 ( .A(b[27]), .B(a[19]), .Z(n4656) );
  OR U4824 ( .A(n4656), .B(n9751), .Z(n4495) );
  NAND U4825 ( .A(n4496), .B(n4495), .Z(n4695) );
  XNOR U4826 ( .A(a[41]), .B(b[5]), .Z(n4659) );
  NANDN U4827 ( .A(n4659), .B(n7905), .Z(n4499) );
  NANDN U4828 ( .A(n4497), .B(n7906), .Z(n4498) );
  AND U4829 ( .A(n4499), .B(n4498), .Z(n4696) );
  XNOR U4830 ( .A(n4695), .B(n4696), .Z(n4698) );
  XOR U4831 ( .A(n4697), .B(n4698), .Z(n4683) );
  NAND U4832 ( .A(n4500), .B(n9105), .Z(n4502) );
  XNOR U4833 ( .A(n9455), .B(a[29]), .Z(n4662) );
  NAND U4834 ( .A(n4662), .B(n9107), .Z(n4501) );
  AND U4835 ( .A(n4502), .B(n4501), .Z(n4638) );
  NAND U4836 ( .A(n4503), .B(n9914), .Z(n4505) );
  XNOR U4837 ( .A(n323), .B(a[15]), .Z(n4665) );
  NANDN U4838 ( .A(n9913), .B(n4665), .Z(n4504) );
  AND U4839 ( .A(n4505), .B(n4504), .Z(n4636) );
  NAND U4840 ( .A(n4506), .B(n7622), .Z(n4508) );
  XNOR U4841 ( .A(a[43]), .B(n316), .Z(n4668) );
  NAND U4842 ( .A(n4668), .B(n7620), .Z(n4507) );
  NAND U4843 ( .A(n4508), .B(n4507), .Z(n4635) );
  XOR U4844 ( .A(n4683), .B(n4684), .Z(n4685) );
  XNOR U4845 ( .A(n4686), .B(n4685), .Z(n4731) );
  NANDN U4846 ( .A(n4510), .B(n4509), .Z(n4514) );
  NANDN U4847 ( .A(n4512), .B(n4511), .Z(n4513) );
  NAND U4848 ( .A(n4514), .B(n4513), .Z(n4674) );
  NAND U4849 ( .A(n4516), .B(n4515), .Z(n4520) );
  NAND U4850 ( .A(n4518), .B(n4517), .Z(n4519) );
  NAND U4851 ( .A(n4520), .B(n4519), .Z(n4672) );
  NANDN U4852 ( .A(n4522), .B(n4521), .Z(n4526) );
  NANDN U4853 ( .A(n4524), .B(n4523), .Z(n4525) );
  NAND U4854 ( .A(n4526), .B(n4525), .Z(n4671) );
  XNOR U4855 ( .A(n4674), .B(n4673), .Z(n4732) );
  XOR U4856 ( .A(n4731), .B(n4732), .Z(n4734) );
  NANDN U4857 ( .A(n4528), .B(n4527), .Z(n4532) );
  OR U4858 ( .A(n4530), .B(n4529), .Z(n4531) );
  NAND U4859 ( .A(n4532), .B(n4531), .Z(n4733) );
  XOR U4860 ( .A(n4734), .B(n4733), .Z(n4751) );
  OR U4861 ( .A(n4534), .B(n4533), .Z(n4538) );
  NANDN U4862 ( .A(n4536), .B(n4535), .Z(n4537) );
  NAND U4863 ( .A(n4538), .B(n4537), .Z(n4750) );
  NANDN U4864 ( .A(n4540), .B(n4539), .Z(n4544) );
  NANDN U4865 ( .A(n4542), .B(n4541), .Z(n4543) );
  NAND U4866 ( .A(n4544), .B(n4543), .Z(n4739) );
  NAND U4867 ( .A(n4546), .B(n4545), .Z(n4550) );
  NAND U4868 ( .A(n4548), .B(n4547), .Z(n4549) );
  NAND U4869 ( .A(n4550), .B(n4549), .Z(n4738) );
  NANDN U4870 ( .A(n4552), .B(n4551), .Z(n4556) );
  NAND U4871 ( .A(n4554), .B(n4553), .Z(n4555) );
  NAND U4872 ( .A(n4556), .B(n4555), .Z(n4677) );
  NANDN U4873 ( .A(n4558), .B(n4557), .Z(n4562) );
  NAND U4874 ( .A(n4560), .B(n4559), .Z(n4561) );
  AND U4875 ( .A(n4562), .B(n4561), .Z(n4678) );
  XNOR U4876 ( .A(n4677), .B(n4678), .Z(n4679) );
  NAND U4877 ( .A(n4563), .B(n8286), .Z(n4565) );
  XOR U4878 ( .A(b[9]), .B(a[37]), .Z(n4701) );
  NAND U4879 ( .A(n4701), .B(n8288), .Z(n4564) );
  NAND U4880 ( .A(n4565), .B(n4564), .Z(n4643) );
  NAND U4881 ( .A(n4566), .B(n8961), .Z(n4568) );
  XOR U4882 ( .A(b[15]), .B(a[31]), .Z(n4704) );
  NAND U4883 ( .A(n4704), .B(n8963), .Z(n4567) );
  NAND U4884 ( .A(n4568), .B(n4567), .Z(n4641) );
  XNOR U4885 ( .A(b[21]), .B(a[25]), .Z(n4707) );
  NANDN U4886 ( .A(n4707), .B(n9493), .Z(n4571) );
  NANDN U4887 ( .A(n4569), .B(n9495), .Z(n4570) );
  AND U4888 ( .A(n4571), .B(n4570), .Z(n4642) );
  XOR U4889 ( .A(n4641), .B(n4642), .Z(n4644) );
  XNOR U4890 ( .A(n4643), .B(n4644), .Z(n4632) );
  XNOR U4891 ( .A(b[11]), .B(a[35]), .Z(n4710) );
  NANDN U4892 ( .A(n4710), .B(n8541), .Z(n4574) );
  NANDN U4893 ( .A(n4572), .B(n8542), .Z(n4573) );
  NAND U4894 ( .A(n4574), .B(n4573), .Z(n4630) );
  XOR U4895 ( .A(b[13]), .B(n6914), .Z(n4713) );
  NANDN U4896 ( .A(n4713), .B(n8730), .Z(n4577) );
  NANDN U4897 ( .A(n4575), .B(n8731), .Z(n4576) );
  NAND U4898 ( .A(n4577), .B(n4576), .Z(n4629) );
  XNOR U4899 ( .A(n4632), .B(n4631), .Z(n4626) );
  ANDN U4900 ( .B(b[31]), .A(n4578), .Z(n4647) );
  NANDN U4901 ( .A(n4579), .B(n9875), .Z(n4581) );
  XNOR U4902 ( .A(n322), .B(a[17]), .Z(n4719) );
  NANDN U4903 ( .A(n9874), .B(n4719), .Z(n4580) );
  NAND U4904 ( .A(n4581), .B(n4580), .Z(n4648) );
  XOR U4905 ( .A(n4647), .B(n4648), .Z(n4649) );
  NANDN U4906 ( .A(n315), .B(a[45]), .Z(n4582) );
  XNOR U4907 ( .A(b[1]), .B(n4582), .Z(n4584) );
  IV U4908 ( .A(a[44]), .Z(n8444) );
  NANDN U4909 ( .A(n8444), .B(n315), .Z(n4583) );
  AND U4910 ( .A(n4584), .B(n4583), .Z(n4650) );
  XNOR U4911 ( .A(n4649), .B(n4650), .Z(n4623) );
  NANDN U4912 ( .A(n4585), .B(n9622), .Z(n4587) );
  XOR U4913 ( .A(b[23]), .B(n6044), .Z(n4722) );
  OR U4914 ( .A(n4722), .B(n9621), .Z(n4586) );
  NAND U4915 ( .A(n4587), .B(n4586), .Z(n4692) );
  XOR U4916 ( .A(b[7]), .B(a[39]), .Z(n4725) );
  NANDN U4917 ( .A(n8013), .B(n4725), .Z(n4590) );
  NANDN U4918 ( .A(n4588), .B(n8014), .Z(n4589) );
  NAND U4919 ( .A(n4590), .B(n4589), .Z(n4689) );
  XNOR U4920 ( .A(b[25]), .B(a[21]), .Z(n4728) );
  NANDN U4921 ( .A(n4728), .B(n9706), .Z(n4593) );
  NANDN U4922 ( .A(n4591), .B(n9707), .Z(n4592) );
  AND U4923 ( .A(n4593), .B(n4592), .Z(n4690) );
  XNOR U4924 ( .A(n4689), .B(n4690), .Z(n4691) );
  XNOR U4925 ( .A(n4692), .B(n4691), .Z(n4624) );
  XOR U4926 ( .A(n4626), .B(n4625), .Z(n4680) );
  XNOR U4927 ( .A(n4679), .B(n4680), .Z(n4737) );
  XNOR U4928 ( .A(n4738), .B(n4737), .Z(n4740) );
  XNOR U4929 ( .A(n4739), .B(n4740), .Z(n4749) );
  XOR U4930 ( .A(n4750), .B(n4749), .Z(n4752) );
  NANDN U4931 ( .A(n4595), .B(n4594), .Z(n4599) );
  NAND U4932 ( .A(n4597), .B(n4596), .Z(n4598) );
  NAND U4933 ( .A(n4599), .B(n4598), .Z(n4744) );
  NAND U4934 ( .A(n4601), .B(n4600), .Z(n4605) );
  NANDN U4935 ( .A(n4603), .B(n4602), .Z(n4604) );
  AND U4936 ( .A(n4605), .B(n4604), .Z(n4743) );
  XNOR U4937 ( .A(n4744), .B(n4743), .Z(n4745) );
  XOR U4938 ( .A(n4746), .B(n4745), .Z(n4620) );
  XOR U4939 ( .A(n4619), .B(n4620), .Z(n4611) );
  XOR U4940 ( .A(n4612), .B(n4611), .Z(n4613) );
  XNOR U4941 ( .A(n4614), .B(n4613), .Z(n4755) );
  XNOR U4942 ( .A(n4755), .B(sreg[77]), .Z(n4757) );
  NAND U4943 ( .A(n4606), .B(sreg[76]), .Z(n4610) );
  OR U4944 ( .A(n4608), .B(n4607), .Z(n4609) );
  AND U4945 ( .A(n4610), .B(n4609), .Z(n4756) );
  XOR U4946 ( .A(n4757), .B(n4756), .Z(c[77]) );
  NAND U4947 ( .A(n4612), .B(n4611), .Z(n4616) );
  NAND U4948 ( .A(n4614), .B(n4613), .Z(n4615) );
  NAND U4949 ( .A(n4616), .B(n4615), .Z(n4763) );
  NANDN U4950 ( .A(n4618), .B(n4617), .Z(n4622) );
  NAND U4951 ( .A(n4620), .B(n4619), .Z(n4621) );
  NAND U4952 ( .A(n4622), .B(n4621), .Z(n4761) );
  OR U4953 ( .A(n4624), .B(n4623), .Z(n4628) );
  NANDN U4954 ( .A(n4626), .B(n4625), .Z(n4627) );
  NAND U4955 ( .A(n4628), .B(n4627), .Z(n4893) );
  OR U4956 ( .A(n4630), .B(n4629), .Z(n4634) );
  NANDN U4957 ( .A(n4632), .B(n4631), .Z(n4633) );
  NAND U4958 ( .A(n4634), .B(n4633), .Z(n4832) );
  NANDN U4959 ( .A(n4636), .B(n4635), .Z(n4640) );
  NANDN U4960 ( .A(n4638), .B(n4637), .Z(n4639) );
  NAND U4961 ( .A(n4640), .B(n4639), .Z(n4831) );
  NANDN U4962 ( .A(n4642), .B(n4641), .Z(n4646) );
  NANDN U4963 ( .A(n4644), .B(n4643), .Z(n4645) );
  NAND U4964 ( .A(n4646), .B(n4645), .Z(n4830) );
  XOR U4965 ( .A(n4832), .B(n4833), .Z(n4891) );
  OR U4966 ( .A(n4648), .B(n4647), .Z(n4652) );
  NANDN U4967 ( .A(n4650), .B(n4649), .Z(n4651) );
  NAND U4968 ( .A(n4652), .B(n4651), .Z(n4845) );
  NAND U4969 ( .A(n4653), .B(n9379), .Z(n4655) );
  XNOR U4970 ( .A(n9562), .B(a[28]), .Z(n4788) );
  NAND U4971 ( .A(n4788), .B(n9378), .Z(n4654) );
  NAND U4972 ( .A(n4655), .B(n4654), .Z(n4856) );
  NANDN U4973 ( .A(n4656), .B(n9801), .Z(n4658) );
  XNOR U4974 ( .A(b[27]), .B(a[20]), .Z(n4791) );
  OR U4975 ( .A(n4791), .B(n9751), .Z(n4657) );
  NAND U4976 ( .A(n4658), .B(n4657), .Z(n4854) );
  XOR U4977 ( .A(a[42]), .B(n317), .Z(n4794) );
  NANDN U4978 ( .A(n4794), .B(n7905), .Z(n4661) );
  NANDN U4979 ( .A(n4659), .B(n7906), .Z(n4660) );
  AND U4980 ( .A(n4661), .B(n4660), .Z(n4855) );
  XNOR U4981 ( .A(n4854), .B(n4855), .Z(n4857) );
  XOR U4982 ( .A(n4856), .B(n4857), .Z(n4842) );
  NAND U4983 ( .A(n4662), .B(n9105), .Z(n4664) );
  XNOR U4984 ( .A(n9455), .B(a[30]), .Z(n4797) );
  NAND U4985 ( .A(n4797), .B(n9107), .Z(n4663) );
  NAND U4986 ( .A(n4664), .B(n4663), .Z(n4814) );
  NAND U4987 ( .A(n4665), .B(n9914), .Z(n4667) );
  XNOR U4988 ( .A(n323), .B(a[16]), .Z(n4800) );
  NANDN U4989 ( .A(n9913), .B(n4800), .Z(n4666) );
  NAND U4990 ( .A(n4667), .B(n4666), .Z(n4812) );
  NAND U4991 ( .A(n4668), .B(n7622), .Z(n4670) );
  XNOR U4992 ( .A(n8444), .B(b[3]), .Z(n4803) );
  NAND U4993 ( .A(n4803), .B(n7620), .Z(n4669) );
  NAND U4994 ( .A(n4670), .B(n4669), .Z(n4813) );
  XOR U4995 ( .A(n4812), .B(n4813), .Z(n4815) );
  XOR U4996 ( .A(n4814), .B(n4815), .Z(n4843) );
  XOR U4997 ( .A(n4842), .B(n4843), .Z(n4844) );
  XNOR U4998 ( .A(n4845), .B(n4844), .Z(n4890) );
  XOR U4999 ( .A(n4891), .B(n4890), .Z(n4892) );
  XNOR U5000 ( .A(n4893), .B(n4892), .Z(n4779) );
  OR U5001 ( .A(n4672), .B(n4671), .Z(n4676) );
  NAND U5002 ( .A(n4674), .B(n4673), .Z(n4675) );
  NAND U5003 ( .A(n4676), .B(n4675), .Z(n4777) );
  NANDN U5004 ( .A(n4678), .B(n4677), .Z(n4682) );
  NANDN U5005 ( .A(n4680), .B(n4679), .Z(n4681) );
  NAND U5006 ( .A(n4682), .B(n4681), .Z(n4896) );
  NAND U5007 ( .A(n4684), .B(n4683), .Z(n4688) );
  NAND U5008 ( .A(n4686), .B(n4685), .Z(n4687) );
  NAND U5009 ( .A(n4688), .B(n4687), .Z(n4895) );
  NANDN U5010 ( .A(n4690), .B(n4689), .Z(n4694) );
  NAND U5011 ( .A(n4692), .B(n4691), .Z(n4693) );
  NAND U5012 ( .A(n4694), .B(n4693), .Z(n4836) );
  NANDN U5013 ( .A(n4696), .B(n4695), .Z(n4700) );
  NAND U5014 ( .A(n4698), .B(n4697), .Z(n4699) );
  AND U5015 ( .A(n4700), .B(n4699), .Z(n4837) );
  XNOR U5016 ( .A(n4836), .B(n4837), .Z(n4838) );
  NAND U5017 ( .A(n4701), .B(n8286), .Z(n4703) );
  XNOR U5018 ( .A(b[9]), .B(n7672), .Z(n4860) );
  NAND U5019 ( .A(n4860), .B(n8288), .Z(n4702) );
  NAND U5020 ( .A(n4703), .B(n4702), .Z(n4820) );
  NAND U5021 ( .A(n4704), .B(n8961), .Z(n4706) );
  XOR U5022 ( .A(b[15]), .B(a[32]), .Z(n4863) );
  NAND U5023 ( .A(n4863), .B(n8963), .Z(n4705) );
  NAND U5024 ( .A(n4706), .B(n4705), .Z(n4818) );
  XOR U5025 ( .A(n318), .B(n6500), .Z(n4866) );
  NAND U5026 ( .A(n4866), .B(n9493), .Z(n4709) );
  NANDN U5027 ( .A(n4707), .B(n9495), .Z(n4708) );
  AND U5028 ( .A(n4709), .B(n4708), .Z(n4819) );
  XOR U5029 ( .A(n4818), .B(n4819), .Z(n4821) );
  XNOR U5030 ( .A(n4820), .B(n4821), .Z(n4809) );
  XOR U5031 ( .A(b[11]), .B(n7293), .Z(n4869) );
  NANDN U5032 ( .A(n4869), .B(n8541), .Z(n4712) );
  NANDN U5033 ( .A(n4710), .B(n8542), .Z(n4711) );
  NAND U5034 ( .A(n4712), .B(n4711), .Z(n4807) );
  XNOR U5035 ( .A(b[13]), .B(a[34]), .Z(n4872) );
  NANDN U5036 ( .A(n4872), .B(n8730), .Z(n4715) );
  NANDN U5037 ( .A(n4713), .B(n8731), .Z(n4714) );
  AND U5038 ( .A(n4715), .B(n4714), .Z(n4806) );
  XNOR U5039 ( .A(n4807), .B(n4806), .Z(n4808) );
  XNOR U5040 ( .A(n4809), .B(n4808), .Z(n4826) );
  NANDN U5041 ( .A(n315), .B(a[46]), .Z(n4716) );
  XNOR U5042 ( .A(b[1]), .B(n4716), .Z(n4718) );
  NANDN U5043 ( .A(b[0]), .B(a[45]), .Z(n4717) );
  AND U5044 ( .A(n4718), .B(n4717), .Z(n4784) );
  NAND U5045 ( .A(n4719), .B(n9875), .Z(n4721) );
  XNOR U5046 ( .A(n322), .B(a[18]), .Z(n4878) );
  NANDN U5047 ( .A(n9874), .B(n4878), .Z(n4720) );
  NAND U5048 ( .A(n4721), .B(n4720), .Z(n4782) );
  NANDN U5049 ( .A(n323), .B(a[14]), .Z(n4783) );
  XNOR U5050 ( .A(n4782), .B(n4783), .Z(n4785) );
  XOR U5051 ( .A(n4784), .B(n4785), .Z(n4824) );
  NANDN U5052 ( .A(n4722), .B(n9622), .Z(n4724) );
  XNOR U5053 ( .A(b[23]), .B(a[24]), .Z(n4881) );
  OR U5054 ( .A(n4881), .B(n9621), .Z(n4723) );
  NAND U5055 ( .A(n4724), .B(n4723), .Z(n4851) );
  XNOR U5056 ( .A(a[40]), .B(b[7]), .Z(n4884) );
  OR U5057 ( .A(n4884), .B(n8013), .Z(n4727) );
  NAND U5058 ( .A(n4725), .B(n8014), .Z(n4726) );
  NAND U5059 ( .A(n4727), .B(n4726), .Z(n4848) );
  XNOR U5060 ( .A(b[25]), .B(a[22]), .Z(n4887) );
  NANDN U5061 ( .A(n4887), .B(n9706), .Z(n4730) );
  NANDN U5062 ( .A(n4728), .B(n9707), .Z(n4729) );
  AND U5063 ( .A(n4730), .B(n4729), .Z(n4849) );
  XNOR U5064 ( .A(n4848), .B(n4849), .Z(n4850) );
  XNOR U5065 ( .A(n4851), .B(n4850), .Z(n4825) );
  XOR U5066 ( .A(n4824), .B(n4825), .Z(n4827) );
  XNOR U5067 ( .A(n4826), .B(n4827), .Z(n4839) );
  XNOR U5068 ( .A(n4838), .B(n4839), .Z(n4894) );
  XNOR U5069 ( .A(n4895), .B(n4894), .Z(n4897) );
  XNOR U5070 ( .A(n4896), .B(n4897), .Z(n4776) );
  XNOR U5071 ( .A(n4777), .B(n4776), .Z(n4778) );
  XOR U5072 ( .A(n4779), .B(n4778), .Z(n4773) );
  NANDN U5073 ( .A(n4732), .B(n4731), .Z(n4736) );
  OR U5074 ( .A(n4734), .B(n4733), .Z(n4735) );
  NAND U5075 ( .A(n4736), .B(n4735), .Z(n4770) );
  NAND U5076 ( .A(n4738), .B(n4737), .Z(n4742) );
  NANDN U5077 ( .A(n4740), .B(n4739), .Z(n4741) );
  NAND U5078 ( .A(n4742), .B(n4741), .Z(n4771) );
  XNOR U5079 ( .A(n4770), .B(n4771), .Z(n4772) );
  XNOR U5080 ( .A(n4773), .B(n4772), .Z(n4767) );
  NANDN U5081 ( .A(n4744), .B(n4743), .Z(n4748) );
  NAND U5082 ( .A(n4746), .B(n4745), .Z(n4747) );
  NAND U5083 ( .A(n4748), .B(n4747), .Z(n4764) );
  NANDN U5084 ( .A(n4750), .B(n4749), .Z(n4754) );
  OR U5085 ( .A(n4752), .B(n4751), .Z(n4753) );
  NAND U5086 ( .A(n4754), .B(n4753), .Z(n4765) );
  XNOR U5087 ( .A(n4764), .B(n4765), .Z(n4766) );
  XNOR U5088 ( .A(n4767), .B(n4766), .Z(n4760) );
  XOR U5089 ( .A(n4761), .B(n4760), .Z(n4762) );
  XNOR U5090 ( .A(n4763), .B(n4762), .Z(n4900) );
  XNOR U5091 ( .A(n4900), .B(sreg[78]), .Z(n4902) );
  NAND U5092 ( .A(n4755), .B(sreg[77]), .Z(n4759) );
  OR U5093 ( .A(n4757), .B(n4756), .Z(n4758) );
  AND U5094 ( .A(n4759), .B(n4758), .Z(n4901) );
  XOR U5095 ( .A(n4902), .B(n4901), .Z(c[78]) );
  NANDN U5096 ( .A(n4765), .B(n4764), .Z(n4769) );
  NANDN U5097 ( .A(n4767), .B(n4766), .Z(n4768) );
  NAND U5098 ( .A(n4769), .B(n4768), .Z(n4906) );
  NANDN U5099 ( .A(n4771), .B(n4770), .Z(n4775) );
  NAND U5100 ( .A(n4773), .B(n4772), .Z(n4774) );
  NAND U5101 ( .A(n4775), .B(n4774), .Z(n4911) );
  NANDN U5102 ( .A(n4777), .B(n4776), .Z(n4781) );
  NANDN U5103 ( .A(n4779), .B(n4778), .Z(n4780) );
  NAND U5104 ( .A(n4781), .B(n4780), .Z(n4912) );
  XNOR U5105 ( .A(n4911), .B(n4912), .Z(n4913) );
  NANDN U5106 ( .A(n4783), .B(n4782), .Z(n4787) );
  NAND U5107 ( .A(n4785), .B(n4784), .Z(n4786) );
  NAND U5108 ( .A(n4787), .B(n4786), .Z(n4990) );
  NAND U5109 ( .A(n4788), .B(n9379), .Z(n4790) );
  XNOR U5110 ( .A(n9562), .B(a[29]), .Z(n4935) );
  NAND U5111 ( .A(n4935), .B(n9378), .Z(n4789) );
  NAND U5112 ( .A(n4790), .B(n4789), .Z(n5001) );
  NANDN U5113 ( .A(n4791), .B(n9801), .Z(n4793) );
  XNOR U5114 ( .A(b[27]), .B(a[21]), .Z(n4938) );
  OR U5115 ( .A(n4938), .B(n9751), .Z(n4792) );
  NAND U5116 ( .A(n4793), .B(n4792), .Z(n4999) );
  XNOR U5117 ( .A(a[43]), .B(b[5]), .Z(n4941) );
  NANDN U5118 ( .A(n4941), .B(n7905), .Z(n4796) );
  NANDN U5119 ( .A(n4794), .B(n7906), .Z(n4795) );
  AND U5120 ( .A(n4796), .B(n4795), .Z(n5000) );
  XNOR U5121 ( .A(n4999), .B(n5000), .Z(n5002) );
  XOR U5122 ( .A(n5001), .B(n5002), .Z(n4987) );
  NAND U5123 ( .A(n4797), .B(n9105), .Z(n4799) );
  XNOR U5124 ( .A(n9455), .B(a[31]), .Z(n4944) );
  NAND U5125 ( .A(n4944), .B(n9107), .Z(n4798) );
  NAND U5126 ( .A(n4799), .B(n4798), .Z(n4961) );
  NAND U5127 ( .A(n4800), .B(n9914), .Z(n4802) );
  XNOR U5128 ( .A(n323), .B(a[17]), .Z(n4947) );
  NANDN U5129 ( .A(n9913), .B(n4947), .Z(n4801) );
  NAND U5130 ( .A(n4802), .B(n4801), .Z(n4959) );
  NAND U5131 ( .A(n4803), .B(n7622), .Z(n4805) );
  XNOR U5132 ( .A(a[45]), .B(n316), .Z(n4950) );
  NAND U5133 ( .A(n4950), .B(n7620), .Z(n4804) );
  NAND U5134 ( .A(n4805), .B(n4804), .Z(n4960) );
  XOR U5135 ( .A(n4959), .B(n4960), .Z(n4962) );
  XOR U5136 ( .A(n4961), .B(n4962), .Z(n4988) );
  XOR U5137 ( .A(n4987), .B(n4988), .Z(n4989) );
  XNOR U5138 ( .A(n4990), .B(n4989), .Z(n5035) );
  NANDN U5139 ( .A(n4807), .B(n4806), .Z(n4811) );
  NANDN U5140 ( .A(n4809), .B(n4808), .Z(n4810) );
  NAND U5141 ( .A(n4811), .B(n4810), .Z(n4978) );
  NAND U5142 ( .A(n4813), .B(n4812), .Z(n4817) );
  NAND U5143 ( .A(n4815), .B(n4814), .Z(n4816) );
  NAND U5144 ( .A(n4817), .B(n4816), .Z(n4976) );
  NANDN U5145 ( .A(n4819), .B(n4818), .Z(n4823) );
  NANDN U5146 ( .A(n4821), .B(n4820), .Z(n4822) );
  NAND U5147 ( .A(n4823), .B(n4822), .Z(n4975) );
  XNOR U5148 ( .A(n4978), .B(n4977), .Z(n5036) );
  XOR U5149 ( .A(n5035), .B(n5036), .Z(n5038) );
  NANDN U5150 ( .A(n4825), .B(n4824), .Z(n4829) );
  OR U5151 ( .A(n4827), .B(n4826), .Z(n4828) );
  NAND U5152 ( .A(n4829), .B(n4828), .Z(n5037) );
  XOR U5153 ( .A(n5038), .B(n5037), .Z(n4925) );
  OR U5154 ( .A(n4831), .B(n4830), .Z(n4835) );
  NANDN U5155 ( .A(n4833), .B(n4832), .Z(n4834) );
  NAND U5156 ( .A(n4835), .B(n4834), .Z(n4924) );
  NANDN U5157 ( .A(n4837), .B(n4836), .Z(n4841) );
  NANDN U5158 ( .A(n4839), .B(n4838), .Z(n4840) );
  NAND U5159 ( .A(n4841), .B(n4840), .Z(n5043) );
  NAND U5160 ( .A(n4843), .B(n4842), .Z(n4847) );
  NANDN U5161 ( .A(n4845), .B(n4844), .Z(n4846) );
  NAND U5162 ( .A(n4847), .B(n4846), .Z(n5042) );
  NANDN U5163 ( .A(n4849), .B(n4848), .Z(n4853) );
  NAND U5164 ( .A(n4851), .B(n4850), .Z(n4852) );
  NAND U5165 ( .A(n4853), .B(n4852), .Z(n4981) );
  NANDN U5166 ( .A(n4855), .B(n4854), .Z(n4859) );
  NAND U5167 ( .A(n4857), .B(n4856), .Z(n4858) );
  AND U5168 ( .A(n4859), .B(n4858), .Z(n4982) );
  XNOR U5169 ( .A(n4981), .B(n4982), .Z(n4983) );
  NAND U5170 ( .A(n4860), .B(n8286), .Z(n4862) );
  XOR U5171 ( .A(b[9]), .B(a[39]), .Z(n5005) );
  NAND U5172 ( .A(n5005), .B(n8288), .Z(n4861) );
  NAND U5173 ( .A(n4862), .B(n4861), .Z(n4967) );
  NAND U5174 ( .A(n4863), .B(n8961), .Z(n4865) );
  XNOR U5175 ( .A(b[15]), .B(n6914), .Z(n5008) );
  NAND U5176 ( .A(n5008), .B(n8963), .Z(n4864) );
  NAND U5177 ( .A(n4865), .B(n4864), .Z(n4966) );
  XNOR U5178 ( .A(b[21]), .B(a[27]), .Z(n5011) );
  NANDN U5179 ( .A(n5011), .B(n9493), .Z(n4868) );
  NAND U5180 ( .A(n9495), .B(n4866), .Z(n4867) );
  NAND U5181 ( .A(n4868), .B(n4867), .Z(n4965) );
  XNOR U5182 ( .A(n4966), .B(n4965), .Z(n4968) );
  XNOR U5183 ( .A(n4967), .B(n4968), .Z(n4956) );
  XNOR U5184 ( .A(b[11]), .B(a[37]), .Z(n5014) );
  NANDN U5185 ( .A(n5014), .B(n8541), .Z(n4871) );
  NANDN U5186 ( .A(n4869), .B(n8542), .Z(n4870) );
  NAND U5187 ( .A(n4871), .B(n4870), .Z(n4954) );
  XNOR U5188 ( .A(b[13]), .B(a[35]), .Z(n5017) );
  NANDN U5189 ( .A(n5017), .B(n8730), .Z(n4874) );
  NANDN U5190 ( .A(n4872), .B(n8731), .Z(n4873) );
  AND U5191 ( .A(n4874), .B(n4873), .Z(n4953) );
  XNOR U5192 ( .A(n4954), .B(n4953), .Z(n4955) );
  XNOR U5193 ( .A(n4956), .B(n4955), .Z(n4972) );
  NANDN U5194 ( .A(n315), .B(a[47]), .Z(n4875) );
  XNOR U5195 ( .A(b[1]), .B(n4875), .Z(n4877) );
  IV U5196 ( .A(a[46]), .Z(n8654) );
  NANDN U5197 ( .A(n8654), .B(n315), .Z(n4876) );
  AND U5198 ( .A(n4877), .B(n4876), .Z(n4931) );
  NAND U5199 ( .A(n9875), .B(n4878), .Z(n4880) );
  XNOR U5200 ( .A(n322), .B(a[19]), .Z(n5023) );
  NANDN U5201 ( .A(n9874), .B(n5023), .Z(n4879) );
  NAND U5202 ( .A(n4880), .B(n4879), .Z(n4929) );
  NANDN U5203 ( .A(n323), .B(a[15]), .Z(n4930) );
  XNOR U5204 ( .A(n4929), .B(n4930), .Z(n4932) );
  XNOR U5205 ( .A(n4931), .B(n4932), .Z(n4970) );
  NANDN U5206 ( .A(n4881), .B(n9622), .Z(n4883) );
  XNOR U5207 ( .A(b[23]), .B(a[25]), .Z(n5026) );
  OR U5208 ( .A(n5026), .B(n9621), .Z(n4882) );
  NAND U5209 ( .A(n4883), .B(n4882), .Z(n4996) );
  XOR U5210 ( .A(b[7]), .B(a[41]), .Z(n5029) );
  NANDN U5211 ( .A(n8013), .B(n5029), .Z(n4886) );
  NANDN U5212 ( .A(n4884), .B(n8014), .Z(n4885) );
  NAND U5213 ( .A(n4886), .B(n4885), .Z(n4993) );
  XOR U5214 ( .A(b[25]), .B(n6044), .Z(n5032) );
  NANDN U5215 ( .A(n5032), .B(n9706), .Z(n4889) );
  NANDN U5216 ( .A(n4887), .B(n9707), .Z(n4888) );
  AND U5217 ( .A(n4889), .B(n4888), .Z(n4994) );
  XNOR U5218 ( .A(n4993), .B(n4994), .Z(n4995) );
  XOR U5219 ( .A(n4996), .B(n4995), .Z(n4969) );
  XOR U5220 ( .A(n4972), .B(n4971), .Z(n4984) );
  XNOR U5221 ( .A(n4983), .B(n4984), .Z(n5041) );
  XNOR U5222 ( .A(n5042), .B(n5041), .Z(n5044) );
  XNOR U5223 ( .A(n5043), .B(n5044), .Z(n4923) );
  XOR U5224 ( .A(n4924), .B(n4923), .Z(n4926) );
  NAND U5225 ( .A(n4895), .B(n4894), .Z(n4899) );
  NANDN U5226 ( .A(n4897), .B(n4896), .Z(n4898) );
  AND U5227 ( .A(n4899), .B(n4898), .Z(n4917) );
  XNOR U5228 ( .A(n4918), .B(n4917), .Z(n4919) );
  XOR U5229 ( .A(n4920), .B(n4919), .Z(n4914) );
  XOR U5230 ( .A(n4913), .B(n4914), .Z(n4905) );
  XOR U5231 ( .A(n4906), .B(n4905), .Z(n4907) );
  XNOR U5232 ( .A(n4908), .B(n4907), .Z(n5047) );
  XNOR U5233 ( .A(n5047), .B(sreg[79]), .Z(n5049) );
  NAND U5234 ( .A(n4900), .B(sreg[78]), .Z(n4904) );
  OR U5235 ( .A(n4902), .B(n4901), .Z(n4903) );
  AND U5236 ( .A(n4904), .B(n4903), .Z(n5048) );
  XOR U5237 ( .A(n5049), .B(n5048), .Z(c[79]) );
  NAND U5238 ( .A(n4906), .B(n4905), .Z(n4910) );
  NAND U5239 ( .A(n4908), .B(n4907), .Z(n4909) );
  NAND U5240 ( .A(n4910), .B(n4909), .Z(n5055) );
  NANDN U5241 ( .A(n4912), .B(n4911), .Z(n4916) );
  NAND U5242 ( .A(n4914), .B(n4913), .Z(n4915) );
  NAND U5243 ( .A(n4916), .B(n4915), .Z(n5053) );
  NANDN U5244 ( .A(n4918), .B(n4917), .Z(n4922) );
  NAND U5245 ( .A(n4920), .B(n4919), .Z(n4921) );
  NAND U5246 ( .A(n4922), .B(n4921), .Z(n5058) );
  NANDN U5247 ( .A(n4924), .B(n4923), .Z(n4928) );
  OR U5248 ( .A(n4926), .B(n4925), .Z(n4927) );
  NAND U5249 ( .A(n4928), .B(n4927), .Z(n5059) );
  XNOR U5250 ( .A(n5058), .B(n5059), .Z(n5060) );
  NANDN U5251 ( .A(n4930), .B(n4929), .Z(n4934) );
  NAND U5252 ( .A(n4932), .B(n4931), .Z(n4933) );
  NAND U5253 ( .A(n4934), .B(n4933), .Z(n5135) );
  NAND U5254 ( .A(n4935), .B(n9379), .Z(n4937) );
  XNOR U5255 ( .A(n9562), .B(a[30]), .Z(n5080) );
  NAND U5256 ( .A(n5080), .B(n9378), .Z(n4936) );
  NAND U5257 ( .A(n4937), .B(n4936), .Z(n5146) );
  NANDN U5258 ( .A(n4938), .B(n9801), .Z(n4940) );
  XNOR U5259 ( .A(b[27]), .B(a[22]), .Z(n5083) );
  OR U5260 ( .A(n5083), .B(n9751), .Z(n4939) );
  NAND U5261 ( .A(n4940), .B(n4939), .Z(n5144) );
  XOR U5262 ( .A(a[44]), .B(n317), .Z(n5086) );
  NANDN U5263 ( .A(n5086), .B(n7905), .Z(n4943) );
  NANDN U5264 ( .A(n4941), .B(n7906), .Z(n4942) );
  AND U5265 ( .A(n4943), .B(n4942), .Z(n5145) );
  XNOR U5266 ( .A(n5144), .B(n5145), .Z(n5147) );
  XOR U5267 ( .A(n5146), .B(n5147), .Z(n5132) );
  NAND U5268 ( .A(n4944), .B(n9105), .Z(n4946) );
  XNOR U5269 ( .A(n9455), .B(a[32]), .Z(n5089) );
  NAND U5270 ( .A(n5089), .B(n9107), .Z(n4945) );
  NAND U5271 ( .A(n4946), .B(n4945), .Z(n5106) );
  NAND U5272 ( .A(n4947), .B(n9914), .Z(n4949) );
  XNOR U5273 ( .A(n323), .B(a[18]), .Z(n5092) );
  NANDN U5274 ( .A(n9913), .B(n5092), .Z(n4948) );
  NAND U5275 ( .A(n4949), .B(n4948), .Z(n5104) );
  NAND U5276 ( .A(n4950), .B(n7622), .Z(n4952) );
  XNOR U5277 ( .A(n8654), .B(b[3]), .Z(n5095) );
  NAND U5278 ( .A(n5095), .B(n7620), .Z(n4951) );
  NAND U5279 ( .A(n4952), .B(n4951), .Z(n5105) );
  XOR U5280 ( .A(n5104), .B(n5105), .Z(n5107) );
  XOR U5281 ( .A(n5106), .B(n5107), .Z(n5133) );
  XOR U5282 ( .A(n5132), .B(n5133), .Z(n5134) );
  XNOR U5283 ( .A(n5135), .B(n5134), .Z(n5071) );
  NANDN U5284 ( .A(n4954), .B(n4953), .Z(n4958) );
  NANDN U5285 ( .A(n4956), .B(n4955), .Z(n4957) );
  NAND U5286 ( .A(n4958), .B(n4957), .Z(n5124) );
  NAND U5287 ( .A(n4960), .B(n4959), .Z(n4964) );
  NAND U5288 ( .A(n4962), .B(n4961), .Z(n4963) );
  NAND U5289 ( .A(n4964), .B(n4963), .Z(n5123) );
  XNOR U5290 ( .A(n5123), .B(n5122), .Z(n5125) );
  XOR U5291 ( .A(n5124), .B(n5125), .Z(n5070) );
  XOR U5292 ( .A(n5071), .B(n5070), .Z(n5072) );
  NANDN U5293 ( .A(n4970), .B(n4969), .Z(n4974) );
  NANDN U5294 ( .A(n4972), .B(n4971), .Z(n4973) );
  NAND U5295 ( .A(n4974), .B(n4973), .Z(n5073) );
  XNOR U5296 ( .A(n5072), .B(n5073), .Z(n5189) );
  OR U5297 ( .A(n4976), .B(n4975), .Z(n4980) );
  NAND U5298 ( .A(n4978), .B(n4977), .Z(n4979) );
  NAND U5299 ( .A(n4980), .B(n4979), .Z(n5188) );
  NANDN U5300 ( .A(n4982), .B(n4981), .Z(n4986) );
  NANDN U5301 ( .A(n4984), .B(n4983), .Z(n4985) );
  NAND U5302 ( .A(n4986), .B(n4985), .Z(n5066) );
  NAND U5303 ( .A(n4988), .B(n4987), .Z(n4992) );
  NAND U5304 ( .A(n4990), .B(n4989), .Z(n4991) );
  NAND U5305 ( .A(n4992), .B(n4991), .Z(n5065) );
  NANDN U5306 ( .A(n4994), .B(n4993), .Z(n4998) );
  NAND U5307 ( .A(n4996), .B(n4995), .Z(n4997) );
  NAND U5308 ( .A(n4998), .B(n4997), .Z(n5126) );
  NANDN U5309 ( .A(n5000), .B(n4999), .Z(n5004) );
  NAND U5310 ( .A(n5002), .B(n5001), .Z(n5003) );
  AND U5311 ( .A(n5004), .B(n5003), .Z(n5127) );
  XNOR U5312 ( .A(n5126), .B(n5127), .Z(n5128) );
  NAND U5313 ( .A(n5005), .B(n8286), .Z(n5007) );
  XNOR U5314 ( .A(b[9]), .B(n7932), .Z(n5150) );
  NAND U5315 ( .A(n5150), .B(n8288), .Z(n5006) );
  NAND U5316 ( .A(n5007), .B(n5006), .Z(n5112) );
  NAND U5317 ( .A(n5008), .B(n8961), .Z(n5010) );
  XOR U5318 ( .A(b[15]), .B(a[34]), .Z(n5153) );
  NAND U5319 ( .A(n5153), .B(n8963), .Z(n5009) );
  NAND U5320 ( .A(n5010), .B(n5009), .Z(n5110) );
  XNOR U5321 ( .A(b[21]), .B(a[28]), .Z(n5156) );
  NANDN U5322 ( .A(n5156), .B(n9493), .Z(n5013) );
  NANDN U5323 ( .A(n5011), .B(n9495), .Z(n5012) );
  AND U5324 ( .A(n5013), .B(n5012), .Z(n5111) );
  XOR U5325 ( .A(n5110), .B(n5111), .Z(n5113) );
  XNOR U5326 ( .A(n5112), .B(n5113), .Z(n5101) );
  XOR U5327 ( .A(b[11]), .B(n7672), .Z(n5159) );
  NANDN U5328 ( .A(n5159), .B(n8541), .Z(n5016) );
  NANDN U5329 ( .A(n5014), .B(n8542), .Z(n5015) );
  NAND U5330 ( .A(n5016), .B(n5015), .Z(n5099) );
  XOR U5331 ( .A(b[13]), .B(n7293), .Z(n5162) );
  NANDN U5332 ( .A(n5162), .B(n8730), .Z(n5019) );
  NANDN U5333 ( .A(n5017), .B(n8731), .Z(n5018) );
  AND U5334 ( .A(n5019), .B(n5018), .Z(n5098) );
  XNOR U5335 ( .A(n5099), .B(n5098), .Z(n5100) );
  XNOR U5336 ( .A(n5101), .B(n5100), .Z(n5118) );
  NANDN U5337 ( .A(n315), .B(a[48]), .Z(n5020) );
  XNOR U5338 ( .A(b[1]), .B(n5020), .Z(n5022) );
  NANDN U5339 ( .A(b[0]), .B(a[47]), .Z(n5021) );
  AND U5340 ( .A(n5022), .B(n5021), .Z(n5076) );
  NAND U5341 ( .A(n9875), .B(n5023), .Z(n5025) );
  XNOR U5342 ( .A(b[29]), .B(a[20]), .Z(n5169) );
  OR U5343 ( .A(n5169), .B(n9874), .Z(n5024) );
  NAND U5344 ( .A(n5025), .B(n5024), .Z(n5074) );
  NANDN U5345 ( .A(n323), .B(a[16]), .Z(n5075) );
  XNOR U5346 ( .A(n5074), .B(n5075), .Z(n5077) );
  XOR U5347 ( .A(n5076), .B(n5077), .Z(n5116) );
  NANDN U5348 ( .A(n5026), .B(n9622), .Z(n5028) );
  XOR U5349 ( .A(b[23]), .B(n6500), .Z(n5172) );
  OR U5350 ( .A(n5172), .B(n9621), .Z(n5027) );
  NAND U5351 ( .A(n5028), .B(n5027), .Z(n5141) );
  XNOR U5352 ( .A(a[42]), .B(b[7]), .Z(n5175) );
  OR U5353 ( .A(n5175), .B(n8013), .Z(n5031) );
  NAND U5354 ( .A(n5029), .B(n8014), .Z(n5030) );
  NAND U5355 ( .A(n5031), .B(n5030), .Z(n5138) );
  XNOR U5356 ( .A(b[25]), .B(a[24]), .Z(n5178) );
  NANDN U5357 ( .A(n5178), .B(n9706), .Z(n5034) );
  NANDN U5358 ( .A(n5032), .B(n9707), .Z(n5033) );
  AND U5359 ( .A(n5034), .B(n5033), .Z(n5139) );
  XNOR U5360 ( .A(n5138), .B(n5139), .Z(n5140) );
  XNOR U5361 ( .A(n5141), .B(n5140), .Z(n5117) );
  XOR U5362 ( .A(n5116), .B(n5117), .Z(n5119) );
  XNOR U5363 ( .A(n5118), .B(n5119), .Z(n5129) );
  XNOR U5364 ( .A(n5128), .B(n5129), .Z(n5064) );
  XNOR U5365 ( .A(n5065), .B(n5064), .Z(n5067) );
  XNOR U5366 ( .A(n5066), .B(n5067), .Z(n5187) );
  XOR U5367 ( .A(n5188), .B(n5187), .Z(n5190) );
  NANDN U5368 ( .A(n5036), .B(n5035), .Z(n5040) );
  OR U5369 ( .A(n5038), .B(n5037), .Z(n5039) );
  NAND U5370 ( .A(n5040), .B(n5039), .Z(n5181) );
  NAND U5371 ( .A(n5042), .B(n5041), .Z(n5046) );
  NANDN U5372 ( .A(n5044), .B(n5043), .Z(n5045) );
  NAND U5373 ( .A(n5046), .B(n5045), .Z(n5182) );
  XNOR U5374 ( .A(n5181), .B(n5182), .Z(n5183) );
  XOR U5375 ( .A(n5184), .B(n5183), .Z(n5061) );
  XOR U5376 ( .A(n5060), .B(n5061), .Z(n5052) );
  XOR U5377 ( .A(n5053), .B(n5052), .Z(n5054) );
  XNOR U5378 ( .A(n5055), .B(n5054), .Z(n5193) );
  XNOR U5379 ( .A(n5193), .B(sreg[80]), .Z(n5195) );
  NAND U5380 ( .A(n5047), .B(sreg[79]), .Z(n5051) );
  OR U5381 ( .A(n5049), .B(n5048), .Z(n5050) );
  AND U5382 ( .A(n5051), .B(n5050), .Z(n5194) );
  XOR U5383 ( .A(n5195), .B(n5194), .Z(c[80]) );
  NAND U5384 ( .A(n5053), .B(n5052), .Z(n5057) );
  NAND U5385 ( .A(n5055), .B(n5054), .Z(n5056) );
  NAND U5386 ( .A(n5057), .B(n5056), .Z(n5201) );
  NANDN U5387 ( .A(n5059), .B(n5058), .Z(n5063) );
  NAND U5388 ( .A(n5061), .B(n5060), .Z(n5062) );
  NAND U5389 ( .A(n5063), .B(n5062), .Z(n5198) );
  NAND U5390 ( .A(n5065), .B(n5064), .Z(n5069) );
  NANDN U5391 ( .A(n5067), .B(n5066), .Z(n5068) );
  NAND U5392 ( .A(n5069), .B(n5068), .Z(n5210) );
  XNOR U5393 ( .A(n5210), .B(n5211), .Z(n5212) );
  NANDN U5394 ( .A(n5075), .B(n5074), .Z(n5079) );
  NAND U5395 ( .A(n5077), .B(n5076), .Z(n5078) );
  NAND U5396 ( .A(n5079), .B(n5078), .Z(n5285) );
  NAND U5397 ( .A(n5080), .B(n9379), .Z(n5082) );
  XNOR U5398 ( .A(n9562), .B(a[31]), .Z(n5252) );
  NAND U5399 ( .A(n5252), .B(n9378), .Z(n5081) );
  NAND U5400 ( .A(n5082), .B(n5081), .Z(n5296) );
  NANDN U5401 ( .A(n5083), .B(n9801), .Z(n5085) );
  XOR U5402 ( .A(b[27]), .B(n6044), .Z(n5255) );
  OR U5403 ( .A(n5255), .B(n9751), .Z(n5084) );
  NAND U5404 ( .A(n5085), .B(n5084), .Z(n5294) );
  XNOR U5405 ( .A(a[45]), .B(b[5]), .Z(n5258) );
  NANDN U5406 ( .A(n5258), .B(n7905), .Z(n5088) );
  NANDN U5407 ( .A(n5086), .B(n7906), .Z(n5087) );
  AND U5408 ( .A(n5088), .B(n5087), .Z(n5295) );
  XNOR U5409 ( .A(n5294), .B(n5295), .Z(n5297) );
  XOR U5410 ( .A(n5296), .B(n5297), .Z(n5282) );
  NAND U5411 ( .A(n5089), .B(n9105), .Z(n5091) );
  XNOR U5412 ( .A(n9455), .B(a[33]), .Z(n5261) );
  NAND U5413 ( .A(n5261), .B(n9107), .Z(n5090) );
  AND U5414 ( .A(n5091), .B(n5090), .Z(n5237) );
  NAND U5415 ( .A(n5092), .B(n9914), .Z(n5094) );
  XNOR U5416 ( .A(n323), .B(a[19]), .Z(n5264) );
  NANDN U5417 ( .A(n9913), .B(n5264), .Z(n5093) );
  AND U5418 ( .A(n5094), .B(n5093), .Z(n5235) );
  NAND U5419 ( .A(n5095), .B(n7622), .Z(n5097) );
  XNOR U5420 ( .A(a[47]), .B(n316), .Z(n5267) );
  NAND U5421 ( .A(n5267), .B(n7620), .Z(n5096) );
  NAND U5422 ( .A(n5097), .B(n5096), .Z(n5234) );
  XOR U5423 ( .A(n5282), .B(n5283), .Z(n5284) );
  XNOR U5424 ( .A(n5285), .B(n5284), .Z(n5330) );
  NANDN U5425 ( .A(n5099), .B(n5098), .Z(n5103) );
  NANDN U5426 ( .A(n5101), .B(n5100), .Z(n5102) );
  NAND U5427 ( .A(n5103), .B(n5102), .Z(n5273) );
  NAND U5428 ( .A(n5105), .B(n5104), .Z(n5109) );
  NAND U5429 ( .A(n5107), .B(n5106), .Z(n5108) );
  NAND U5430 ( .A(n5109), .B(n5108), .Z(n5271) );
  NANDN U5431 ( .A(n5111), .B(n5110), .Z(n5115) );
  NANDN U5432 ( .A(n5113), .B(n5112), .Z(n5114) );
  NAND U5433 ( .A(n5115), .B(n5114), .Z(n5270) );
  XNOR U5434 ( .A(n5273), .B(n5272), .Z(n5331) );
  XNOR U5435 ( .A(n5330), .B(n5331), .Z(n5332) );
  NANDN U5436 ( .A(n5117), .B(n5116), .Z(n5121) );
  OR U5437 ( .A(n5119), .B(n5118), .Z(n5120) );
  AND U5438 ( .A(n5121), .B(n5120), .Z(n5333) );
  XOR U5439 ( .A(n5332), .B(n5333), .Z(n5218) );
  NANDN U5440 ( .A(n5127), .B(n5126), .Z(n5131) );
  NANDN U5441 ( .A(n5129), .B(n5128), .Z(n5130) );
  NAND U5442 ( .A(n5131), .B(n5130), .Z(n5339) );
  NAND U5443 ( .A(n5133), .B(n5132), .Z(n5137) );
  NAND U5444 ( .A(n5135), .B(n5134), .Z(n5136) );
  NAND U5445 ( .A(n5137), .B(n5136), .Z(n5337) );
  NANDN U5446 ( .A(n5139), .B(n5138), .Z(n5143) );
  NAND U5447 ( .A(n5141), .B(n5140), .Z(n5142) );
  NAND U5448 ( .A(n5143), .B(n5142), .Z(n5276) );
  NANDN U5449 ( .A(n5145), .B(n5144), .Z(n5149) );
  NAND U5450 ( .A(n5147), .B(n5146), .Z(n5148) );
  AND U5451 ( .A(n5149), .B(n5148), .Z(n5277) );
  XNOR U5452 ( .A(n5276), .B(n5277), .Z(n5278) );
  NAND U5453 ( .A(n5150), .B(n8286), .Z(n5152) );
  XOR U5454 ( .A(b[9]), .B(a[41]), .Z(n5300) );
  NAND U5455 ( .A(n5300), .B(n8288), .Z(n5151) );
  NAND U5456 ( .A(n5152), .B(n5151), .Z(n5242) );
  NAND U5457 ( .A(n5153), .B(n8961), .Z(n5155) );
  XOR U5458 ( .A(b[15]), .B(a[35]), .Z(n5303) );
  NAND U5459 ( .A(n5303), .B(n8963), .Z(n5154) );
  NAND U5460 ( .A(n5155), .B(n5154), .Z(n5240) );
  XNOR U5461 ( .A(b[21]), .B(a[29]), .Z(n5306) );
  NANDN U5462 ( .A(n5306), .B(n9493), .Z(n5158) );
  NANDN U5463 ( .A(n5156), .B(n9495), .Z(n5157) );
  AND U5464 ( .A(n5158), .B(n5157), .Z(n5241) );
  XOR U5465 ( .A(n5240), .B(n5241), .Z(n5243) );
  XNOR U5466 ( .A(n5242), .B(n5243), .Z(n5231) );
  XNOR U5467 ( .A(b[11]), .B(a[39]), .Z(n5309) );
  NANDN U5468 ( .A(n5309), .B(n8541), .Z(n5161) );
  NANDN U5469 ( .A(n5159), .B(n8542), .Z(n5160) );
  NAND U5470 ( .A(n5161), .B(n5160), .Z(n5229) );
  XNOR U5471 ( .A(b[13]), .B(a[37]), .Z(n5312) );
  NANDN U5472 ( .A(n5312), .B(n8730), .Z(n5164) );
  NANDN U5473 ( .A(n5162), .B(n8731), .Z(n5163) );
  NAND U5474 ( .A(n5164), .B(n5163), .Z(n5228) );
  XNOR U5475 ( .A(n5231), .B(n5230), .Z(n5225) );
  NANDN U5476 ( .A(n315), .B(a[49]), .Z(n5165) );
  XNOR U5477 ( .A(b[1]), .B(n5165), .Z(n5167) );
  IV U5478 ( .A(a[48]), .Z(n8837) );
  NANDN U5479 ( .A(n8837), .B(n315), .Z(n5166) );
  AND U5480 ( .A(n5167), .B(n5166), .Z(n5249) );
  ANDN U5481 ( .B(b[31]), .A(n5168), .Z(n5246) );
  NANDN U5482 ( .A(n5169), .B(n9875), .Z(n5171) );
  XNOR U5483 ( .A(n322), .B(a[21]), .Z(n5318) );
  NANDN U5484 ( .A(n9874), .B(n5318), .Z(n5170) );
  NAND U5485 ( .A(n5171), .B(n5170), .Z(n5247) );
  XOR U5486 ( .A(n5246), .B(n5247), .Z(n5248) );
  XNOR U5487 ( .A(n5249), .B(n5248), .Z(n5222) );
  NANDN U5488 ( .A(n5172), .B(n9622), .Z(n5174) );
  XNOR U5489 ( .A(b[23]), .B(a[27]), .Z(n5321) );
  OR U5490 ( .A(n5321), .B(n9621), .Z(n5173) );
  NAND U5491 ( .A(n5174), .B(n5173), .Z(n5291) );
  XOR U5492 ( .A(a[43]), .B(b[7]), .Z(n5324) );
  NANDN U5493 ( .A(n8013), .B(n5324), .Z(n5177) );
  NANDN U5494 ( .A(n5175), .B(n8014), .Z(n5176) );
  NAND U5495 ( .A(n5177), .B(n5176), .Z(n5288) );
  XNOR U5496 ( .A(b[25]), .B(a[25]), .Z(n5327) );
  NANDN U5497 ( .A(n5327), .B(n9706), .Z(n5180) );
  NANDN U5498 ( .A(n5178), .B(n9707), .Z(n5179) );
  AND U5499 ( .A(n5180), .B(n5179), .Z(n5289) );
  XNOR U5500 ( .A(n5288), .B(n5289), .Z(n5290) );
  XNOR U5501 ( .A(n5291), .B(n5290), .Z(n5223) );
  XOR U5502 ( .A(n5225), .B(n5224), .Z(n5279) );
  XNOR U5503 ( .A(n5278), .B(n5279), .Z(n5336) );
  XOR U5504 ( .A(n5337), .B(n5336), .Z(n5338) );
  XNOR U5505 ( .A(n5339), .B(n5338), .Z(n5216) );
  XNOR U5506 ( .A(n5217), .B(n5216), .Z(n5219) );
  XNOR U5507 ( .A(n5218), .B(n5219), .Z(n5213) );
  XOR U5508 ( .A(n5212), .B(n5213), .Z(n5207) );
  NANDN U5509 ( .A(n5182), .B(n5181), .Z(n5186) );
  NAND U5510 ( .A(n5184), .B(n5183), .Z(n5185) );
  NAND U5511 ( .A(n5186), .B(n5185), .Z(n5204) );
  NANDN U5512 ( .A(n5188), .B(n5187), .Z(n5192) );
  OR U5513 ( .A(n5190), .B(n5189), .Z(n5191) );
  NAND U5514 ( .A(n5192), .B(n5191), .Z(n5205) );
  XNOR U5515 ( .A(n5204), .B(n5205), .Z(n5206) );
  XNOR U5516 ( .A(n5207), .B(n5206), .Z(n5199) );
  XNOR U5517 ( .A(n5198), .B(n5199), .Z(n5200) );
  XNOR U5518 ( .A(n5201), .B(n5200), .Z(n5342) );
  XNOR U5519 ( .A(n5342), .B(sreg[81]), .Z(n5344) );
  NAND U5520 ( .A(n5193), .B(sreg[80]), .Z(n5197) );
  OR U5521 ( .A(n5195), .B(n5194), .Z(n5196) );
  AND U5522 ( .A(n5197), .B(n5196), .Z(n5343) );
  XOR U5523 ( .A(n5344), .B(n5343), .Z(c[81]) );
  NANDN U5524 ( .A(n5199), .B(n5198), .Z(n5203) );
  NAND U5525 ( .A(n5201), .B(n5200), .Z(n5202) );
  NAND U5526 ( .A(n5203), .B(n5202), .Z(n5350) );
  NANDN U5527 ( .A(n5205), .B(n5204), .Z(n5209) );
  NAND U5528 ( .A(n5207), .B(n5206), .Z(n5208) );
  NAND U5529 ( .A(n5209), .B(n5208), .Z(n5348) );
  NANDN U5530 ( .A(n5211), .B(n5210), .Z(n5215) );
  NANDN U5531 ( .A(n5213), .B(n5212), .Z(n5214) );
  NAND U5532 ( .A(n5215), .B(n5214), .Z(n5354) );
  OR U5533 ( .A(n5217), .B(n5216), .Z(n5221) );
  OR U5534 ( .A(n5219), .B(n5218), .Z(n5220) );
  AND U5535 ( .A(n5221), .B(n5220), .Z(n5353) );
  XNOR U5536 ( .A(n5354), .B(n5353), .Z(n5355) );
  OR U5537 ( .A(n5223), .B(n5222), .Z(n5227) );
  NANDN U5538 ( .A(n5225), .B(n5224), .Z(n5226) );
  NAND U5539 ( .A(n5227), .B(n5226), .Z(n5482) );
  OR U5540 ( .A(n5229), .B(n5228), .Z(n5233) );
  NANDN U5541 ( .A(n5231), .B(n5230), .Z(n5232) );
  NAND U5542 ( .A(n5233), .B(n5232), .Z(n5421) );
  NANDN U5543 ( .A(n5235), .B(n5234), .Z(n5239) );
  NANDN U5544 ( .A(n5237), .B(n5236), .Z(n5238) );
  NAND U5545 ( .A(n5239), .B(n5238), .Z(n5420) );
  NANDN U5546 ( .A(n5241), .B(n5240), .Z(n5245) );
  NANDN U5547 ( .A(n5243), .B(n5242), .Z(n5244) );
  NAND U5548 ( .A(n5245), .B(n5244), .Z(n5419) );
  XOR U5549 ( .A(n5421), .B(n5422), .Z(n5480) );
  OR U5550 ( .A(n5247), .B(n5246), .Z(n5251) );
  NANDN U5551 ( .A(n5249), .B(n5248), .Z(n5250) );
  NAND U5552 ( .A(n5251), .B(n5250), .Z(n5434) );
  NAND U5553 ( .A(n5252), .B(n9379), .Z(n5254) );
  XNOR U5554 ( .A(n9562), .B(a[32]), .Z(n5377) );
  NAND U5555 ( .A(n5377), .B(n9378), .Z(n5253) );
  NAND U5556 ( .A(n5254), .B(n5253), .Z(n5445) );
  NANDN U5557 ( .A(n5255), .B(n9801), .Z(n5257) );
  XNOR U5558 ( .A(b[27]), .B(a[24]), .Z(n5380) );
  OR U5559 ( .A(n5380), .B(n9751), .Z(n5256) );
  NAND U5560 ( .A(n5257), .B(n5256), .Z(n5443) );
  XOR U5561 ( .A(a[46]), .B(n317), .Z(n5383) );
  NANDN U5562 ( .A(n5383), .B(n7905), .Z(n5260) );
  NANDN U5563 ( .A(n5258), .B(n7906), .Z(n5259) );
  AND U5564 ( .A(n5260), .B(n5259), .Z(n5444) );
  XNOR U5565 ( .A(n5443), .B(n5444), .Z(n5446) );
  XOR U5566 ( .A(n5445), .B(n5446), .Z(n5431) );
  NAND U5567 ( .A(n5261), .B(n9105), .Z(n5263) );
  XNOR U5568 ( .A(n9455), .B(a[34]), .Z(n5386) );
  NAND U5569 ( .A(n5386), .B(n9107), .Z(n5262) );
  NAND U5570 ( .A(n5263), .B(n5262), .Z(n5403) );
  NAND U5571 ( .A(n5264), .B(n9914), .Z(n5266) );
  XNOR U5572 ( .A(n323), .B(a[20]), .Z(n5389) );
  NANDN U5573 ( .A(n9913), .B(n5389), .Z(n5265) );
  NAND U5574 ( .A(n5266), .B(n5265), .Z(n5401) );
  NAND U5575 ( .A(n5267), .B(n7622), .Z(n5269) );
  XNOR U5576 ( .A(n8837), .B(b[3]), .Z(n5392) );
  NAND U5577 ( .A(n5392), .B(n7620), .Z(n5268) );
  NAND U5578 ( .A(n5269), .B(n5268), .Z(n5402) );
  XOR U5579 ( .A(n5401), .B(n5402), .Z(n5404) );
  XOR U5580 ( .A(n5403), .B(n5404), .Z(n5432) );
  XOR U5581 ( .A(n5431), .B(n5432), .Z(n5433) );
  XNOR U5582 ( .A(n5434), .B(n5433), .Z(n5479) );
  XOR U5583 ( .A(n5480), .B(n5479), .Z(n5481) );
  XNOR U5584 ( .A(n5482), .B(n5481), .Z(n5368) );
  OR U5585 ( .A(n5271), .B(n5270), .Z(n5275) );
  NAND U5586 ( .A(n5273), .B(n5272), .Z(n5274) );
  NAND U5587 ( .A(n5275), .B(n5274), .Z(n5366) );
  NANDN U5588 ( .A(n5277), .B(n5276), .Z(n5281) );
  NANDN U5589 ( .A(n5279), .B(n5278), .Z(n5280) );
  NAND U5590 ( .A(n5281), .B(n5280), .Z(n5485) );
  NAND U5591 ( .A(n5283), .B(n5282), .Z(n5287) );
  NAND U5592 ( .A(n5285), .B(n5284), .Z(n5286) );
  NAND U5593 ( .A(n5287), .B(n5286), .Z(n5484) );
  NANDN U5594 ( .A(n5289), .B(n5288), .Z(n5293) );
  NAND U5595 ( .A(n5291), .B(n5290), .Z(n5292) );
  NAND U5596 ( .A(n5293), .B(n5292), .Z(n5425) );
  NANDN U5597 ( .A(n5295), .B(n5294), .Z(n5299) );
  NAND U5598 ( .A(n5297), .B(n5296), .Z(n5298) );
  AND U5599 ( .A(n5299), .B(n5298), .Z(n5426) );
  XNOR U5600 ( .A(n5425), .B(n5426), .Z(n5427) );
  NAND U5601 ( .A(n5300), .B(n8286), .Z(n5302) );
  XNOR U5602 ( .A(b[9]), .B(n8156), .Z(n5449) );
  NAND U5603 ( .A(n5449), .B(n8288), .Z(n5301) );
  NAND U5604 ( .A(n5302), .B(n5301), .Z(n5409) );
  NAND U5605 ( .A(n5303), .B(n8961), .Z(n5305) );
  XNOR U5606 ( .A(b[15]), .B(n7293), .Z(n5452) );
  NAND U5607 ( .A(n5452), .B(n8963), .Z(n5304) );
  NAND U5608 ( .A(n5305), .B(n5304), .Z(n5407) );
  XOR U5609 ( .A(b[21]), .B(n6135), .Z(n5455) );
  NANDN U5610 ( .A(n5455), .B(n9493), .Z(n5308) );
  NANDN U5611 ( .A(n5306), .B(n9495), .Z(n5307) );
  AND U5612 ( .A(n5308), .B(n5307), .Z(n5408) );
  XOR U5613 ( .A(n5407), .B(n5408), .Z(n5410) );
  XNOR U5614 ( .A(n5409), .B(n5410), .Z(n5398) );
  XOR U5615 ( .A(b[11]), .B(n7932), .Z(n5458) );
  NANDN U5616 ( .A(n5458), .B(n8541), .Z(n5311) );
  NANDN U5617 ( .A(n5309), .B(n8542), .Z(n5310) );
  NAND U5618 ( .A(n5311), .B(n5310), .Z(n5396) );
  XOR U5619 ( .A(b[13]), .B(n7672), .Z(n5461) );
  NANDN U5620 ( .A(n5461), .B(n8730), .Z(n5314) );
  NANDN U5621 ( .A(n5312), .B(n8731), .Z(n5313) );
  AND U5622 ( .A(n5314), .B(n5313), .Z(n5395) );
  XNOR U5623 ( .A(n5396), .B(n5395), .Z(n5397) );
  XNOR U5624 ( .A(n5398), .B(n5397), .Z(n5415) );
  NANDN U5625 ( .A(n315), .B(a[50]), .Z(n5315) );
  XNOR U5626 ( .A(b[1]), .B(n5315), .Z(n5317) );
  NANDN U5627 ( .A(b[0]), .B(a[49]), .Z(n5316) );
  AND U5628 ( .A(n5317), .B(n5316), .Z(n5373) );
  NAND U5629 ( .A(n5318), .B(n9875), .Z(n5320) );
  XNOR U5630 ( .A(n322), .B(a[22]), .Z(n5467) );
  NANDN U5631 ( .A(n9874), .B(n5467), .Z(n5319) );
  NAND U5632 ( .A(n5320), .B(n5319), .Z(n5371) );
  NANDN U5633 ( .A(n323), .B(a[18]), .Z(n5372) );
  XNOR U5634 ( .A(n5371), .B(n5372), .Z(n5374) );
  XOR U5635 ( .A(n5373), .B(n5374), .Z(n5413) );
  NANDN U5636 ( .A(n5321), .B(n9622), .Z(n5323) );
  XNOR U5637 ( .A(b[23]), .B(a[28]), .Z(n5470) );
  OR U5638 ( .A(n5470), .B(n9621), .Z(n5322) );
  NAND U5639 ( .A(n5323), .B(n5322), .Z(n5440) );
  XNOR U5640 ( .A(a[44]), .B(b[7]), .Z(n5473) );
  OR U5641 ( .A(n5473), .B(n8013), .Z(n5326) );
  NAND U5642 ( .A(n5324), .B(n8014), .Z(n5325) );
  NAND U5643 ( .A(n5326), .B(n5325), .Z(n5437) );
  XOR U5644 ( .A(b[25]), .B(n6500), .Z(n5476) );
  NANDN U5645 ( .A(n5476), .B(n9706), .Z(n5329) );
  NANDN U5646 ( .A(n5327), .B(n9707), .Z(n5328) );
  AND U5647 ( .A(n5329), .B(n5328), .Z(n5438) );
  XNOR U5648 ( .A(n5437), .B(n5438), .Z(n5439) );
  XNOR U5649 ( .A(n5440), .B(n5439), .Z(n5414) );
  XOR U5650 ( .A(n5413), .B(n5414), .Z(n5416) );
  XNOR U5651 ( .A(n5415), .B(n5416), .Z(n5428) );
  XNOR U5652 ( .A(n5427), .B(n5428), .Z(n5483) );
  XNOR U5653 ( .A(n5484), .B(n5483), .Z(n5486) );
  XNOR U5654 ( .A(n5485), .B(n5486), .Z(n5365) );
  XNOR U5655 ( .A(n5366), .B(n5365), .Z(n5367) );
  XOR U5656 ( .A(n5368), .B(n5367), .Z(n5362) );
  NANDN U5657 ( .A(n5331), .B(n5330), .Z(n5335) );
  NAND U5658 ( .A(n5333), .B(n5332), .Z(n5334) );
  NAND U5659 ( .A(n5335), .B(n5334), .Z(n5359) );
  NAND U5660 ( .A(n5337), .B(n5336), .Z(n5341) );
  NAND U5661 ( .A(n5339), .B(n5338), .Z(n5340) );
  NAND U5662 ( .A(n5341), .B(n5340), .Z(n5360) );
  XNOR U5663 ( .A(n5359), .B(n5360), .Z(n5361) );
  XOR U5664 ( .A(n5362), .B(n5361), .Z(n5356) );
  XOR U5665 ( .A(n5355), .B(n5356), .Z(n5347) );
  XOR U5666 ( .A(n5348), .B(n5347), .Z(n5349) );
  XNOR U5667 ( .A(n5350), .B(n5349), .Z(n5489) );
  XNOR U5668 ( .A(n5489), .B(sreg[82]), .Z(n5491) );
  NAND U5669 ( .A(n5342), .B(sreg[81]), .Z(n5346) );
  OR U5670 ( .A(n5344), .B(n5343), .Z(n5345) );
  AND U5671 ( .A(n5346), .B(n5345), .Z(n5490) );
  XOR U5672 ( .A(n5491), .B(n5490), .Z(c[82]) );
  NAND U5673 ( .A(n5348), .B(n5347), .Z(n5352) );
  NAND U5674 ( .A(n5350), .B(n5349), .Z(n5351) );
  NAND U5675 ( .A(n5352), .B(n5351), .Z(n5497) );
  NANDN U5676 ( .A(n5354), .B(n5353), .Z(n5358) );
  NAND U5677 ( .A(n5356), .B(n5355), .Z(n5357) );
  NAND U5678 ( .A(n5358), .B(n5357), .Z(n5495) );
  NANDN U5679 ( .A(n5360), .B(n5359), .Z(n5364) );
  NAND U5680 ( .A(n5362), .B(n5361), .Z(n5363) );
  NAND U5681 ( .A(n5364), .B(n5363), .Z(n5500) );
  NANDN U5682 ( .A(n5366), .B(n5365), .Z(n5370) );
  NANDN U5683 ( .A(n5368), .B(n5367), .Z(n5369) );
  NAND U5684 ( .A(n5370), .B(n5369), .Z(n5501) );
  XNOR U5685 ( .A(n5500), .B(n5501), .Z(n5502) );
  NANDN U5686 ( .A(n5372), .B(n5371), .Z(n5376) );
  NAND U5687 ( .A(n5374), .B(n5373), .Z(n5375) );
  NAND U5688 ( .A(n5376), .B(n5375), .Z(n5581) );
  NAND U5689 ( .A(n5377), .B(n9379), .Z(n5379) );
  XNOR U5690 ( .A(n9562), .B(a[33]), .Z(n5524) );
  NAND U5691 ( .A(n5524), .B(n9378), .Z(n5378) );
  NAND U5692 ( .A(n5379), .B(n5378), .Z(n5592) );
  NANDN U5693 ( .A(n5380), .B(n9801), .Z(n5382) );
  XNOR U5694 ( .A(b[27]), .B(a[25]), .Z(n5527) );
  OR U5695 ( .A(n5527), .B(n9751), .Z(n5381) );
  NAND U5696 ( .A(n5382), .B(n5381), .Z(n5590) );
  XNOR U5697 ( .A(a[47]), .B(b[5]), .Z(n5530) );
  NANDN U5698 ( .A(n5530), .B(n7905), .Z(n5385) );
  NANDN U5699 ( .A(n5383), .B(n7906), .Z(n5384) );
  AND U5700 ( .A(n5385), .B(n5384), .Z(n5591) );
  XNOR U5701 ( .A(n5590), .B(n5591), .Z(n5593) );
  XOR U5702 ( .A(n5592), .B(n5593), .Z(n5578) );
  NAND U5703 ( .A(n5386), .B(n9105), .Z(n5388) );
  XNOR U5704 ( .A(n9455), .B(a[35]), .Z(n5533) );
  NAND U5705 ( .A(n5533), .B(n9107), .Z(n5387) );
  NAND U5706 ( .A(n5388), .B(n5387), .Z(n5550) );
  NAND U5707 ( .A(n5389), .B(n9914), .Z(n5391) );
  XNOR U5708 ( .A(n323), .B(a[21]), .Z(n5536) );
  NANDN U5709 ( .A(n9913), .B(n5536), .Z(n5390) );
  NAND U5710 ( .A(n5391), .B(n5390), .Z(n5548) );
  NAND U5711 ( .A(n5392), .B(n7622), .Z(n5394) );
  XNOR U5712 ( .A(a[49]), .B(n316), .Z(n5539) );
  NAND U5713 ( .A(n5539), .B(n7620), .Z(n5393) );
  NAND U5714 ( .A(n5394), .B(n5393), .Z(n5549) );
  XOR U5715 ( .A(n5548), .B(n5549), .Z(n5551) );
  XOR U5716 ( .A(n5550), .B(n5551), .Z(n5579) );
  XOR U5717 ( .A(n5578), .B(n5579), .Z(n5580) );
  XNOR U5718 ( .A(n5581), .B(n5580), .Z(n5626) );
  NANDN U5719 ( .A(n5396), .B(n5395), .Z(n5400) );
  NANDN U5720 ( .A(n5398), .B(n5397), .Z(n5399) );
  NAND U5721 ( .A(n5400), .B(n5399), .Z(n5569) );
  NAND U5722 ( .A(n5402), .B(n5401), .Z(n5406) );
  NAND U5723 ( .A(n5404), .B(n5403), .Z(n5405) );
  NAND U5724 ( .A(n5406), .B(n5405), .Z(n5567) );
  NANDN U5725 ( .A(n5408), .B(n5407), .Z(n5412) );
  NANDN U5726 ( .A(n5410), .B(n5409), .Z(n5411) );
  NAND U5727 ( .A(n5412), .B(n5411), .Z(n5566) );
  XNOR U5728 ( .A(n5569), .B(n5568), .Z(n5627) );
  XOR U5729 ( .A(n5626), .B(n5627), .Z(n5629) );
  NANDN U5730 ( .A(n5414), .B(n5413), .Z(n5418) );
  OR U5731 ( .A(n5416), .B(n5415), .Z(n5417) );
  NAND U5732 ( .A(n5418), .B(n5417), .Z(n5628) );
  XOR U5733 ( .A(n5629), .B(n5628), .Z(n5514) );
  OR U5734 ( .A(n5420), .B(n5419), .Z(n5424) );
  NANDN U5735 ( .A(n5422), .B(n5421), .Z(n5423) );
  NAND U5736 ( .A(n5424), .B(n5423), .Z(n5513) );
  NANDN U5737 ( .A(n5426), .B(n5425), .Z(n5430) );
  NANDN U5738 ( .A(n5428), .B(n5427), .Z(n5429) );
  NAND U5739 ( .A(n5430), .B(n5429), .Z(n5634) );
  NAND U5740 ( .A(n5432), .B(n5431), .Z(n5436) );
  NANDN U5741 ( .A(n5434), .B(n5433), .Z(n5435) );
  NAND U5742 ( .A(n5436), .B(n5435), .Z(n5633) );
  NANDN U5743 ( .A(n5438), .B(n5437), .Z(n5442) );
  NAND U5744 ( .A(n5440), .B(n5439), .Z(n5441) );
  NAND U5745 ( .A(n5442), .B(n5441), .Z(n5572) );
  NANDN U5746 ( .A(n5444), .B(n5443), .Z(n5448) );
  NAND U5747 ( .A(n5446), .B(n5445), .Z(n5447) );
  AND U5748 ( .A(n5448), .B(n5447), .Z(n5573) );
  XNOR U5749 ( .A(n5572), .B(n5573), .Z(n5574) );
  NAND U5750 ( .A(n5449), .B(n8286), .Z(n5451) );
  XOR U5751 ( .A(b[9]), .B(a[43]), .Z(n5596) );
  NAND U5752 ( .A(n5596), .B(n8288), .Z(n5450) );
  NAND U5753 ( .A(n5451), .B(n5450), .Z(n5556) );
  NAND U5754 ( .A(n5452), .B(n8961), .Z(n5454) );
  XOR U5755 ( .A(b[15]), .B(a[37]), .Z(n5599) );
  NAND U5756 ( .A(n5599), .B(n8963), .Z(n5453) );
  NAND U5757 ( .A(n5454), .B(n5453), .Z(n5554) );
  XNOR U5758 ( .A(b[21]), .B(a[31]), .Z(n5602) );
  NANDN U5759 ( .A(n5602), .B(n9493), .Z(n5457) );
  NANDN U5760 ( .A(n5455), .B(n9495), .Z(n5456) );
  AND U5761 ( .A(n5457), .B(n5456), .Z(n5555) );
  XOR U5762 ( .A(n5554), .B(n5555), .Z(n5557) );
  XNOR U5763 ( .A(n5556), .B(n5557), .Z(n5545) );
  XNOR U5764 ( .A(b[11]), .B(a[41]), .Z(n5605) );
  NANDN U5765 ( .A(n5605), .B(n8541), .Z(n5460) );
  NANDN U5766 ( .A(n5458), .B(n8542), .Z(n5459) );
  NAND U5767 ( .A(n5460), .B(n5459), .Z(n5543) );
  XNOR U5768 ( .A(b[13]), .B(a[39]), .Z(n5608) );
  NANDN U5769 ( .A(n5608), .B(n8730), .Z(n5463) );
  NANDN U5770 ( .A(n5461), .B(n8731), .Z(n5462) );
  AND U5771 ( .A(n5463), .B(n5462), .Z(n5542) );
  XNOR U5772 ( .A(n5543), .B(n5542), .Z(n5544) );
  XNOR U5773 ( .A(n5545), .B(n5544), .Z(n5562) );
  NANDN U5774 ( .A(n315), .B(a[51]), .Z(n5464) );
  XNOR U5775 ( .A(b[1]), .B(n5464), .Z(n5466) );
  IV U5776 ( .A(a[50]), .Z(n9033) );
  NANDN U5777 ( .A(n9033), .B(n315), .Z(n5465) );
  AND U5778 ( .A(n5466), .B(n5465), .Z(n5520) );
  NAND U5779 ( .A(n9875), .B(n5467), .Z(n5469) );
  XOR U5780 ( .A(n322), .B(n6044), .Z(n5614) );
  NANDN U5781 ( .A(n9874), .B(n5614), .Z(n5468) );
  NAND U5782 ( .A(n5469), .B(n5468), .Z(n5518) );
  NANDN U5783 ( .A(n323), .B(a[19]), .Z(n5519) );
  XNOR U5784 ( .A(n5518), .B(n5519), .Z(n5521) );
  XOR U5785 ( .A(n5520), .B(n5521), .Z(n5560) );
  NANDN U5786 ( .A(n5470), .B(n9622), .Z(n5472) );
  XNOR U5787 ( .A(b[23]), .B(a[29]), .Z(n5617) );
  OR U5788 ( .A(n5617), .B(n9621), .Z(n5471) );
  NAND U5789 ( .A(n5472), .B(n5471), .Z(n5587) );
  XOR U5790 ( .A(a[45]), .B(b[7]), .Z(n5620) );
  NANDN U5791 ( .A(n8013), .B(n5620), .Z(n5475) );
  NANDN U5792 ( .A(n5473), .B(n8014), .Z(n5474) );
  NAND U5793 ( .A(n5475), .B(n5474), .Z(n5584) );
  XNOR U5794 ( .A(b[25]), .B(a[27]), .Z(n5623) );
  NANDN U5795 ( .A(n5623), .B(n9706), .Z(n5478) );
  NANDN U5796 ( .A(n5476), .B(n9707), .Z(n5477) );
  AND U5797 ( .A(n5478), .B(n5477), .Z(n5585) );
  XNOR U5798 ( .A(n5584), .B(n5585), .Z(n5586) );
  XNOR U5799 ( .A(n5587), .B(n5586), .Z(n5561) );
  XOR U5800 ( .A(n5560), .B(n5561), .Z(n5563) );
  XNOR U5801 ( .A(n5562), .B(n5563), .Z(n5575) );
  XNOR U5802 ( .A(n5574), .B(n5575), .Z(n5632) );
  XNOR U5803 ( .A(n5633), .B(n5632), .Z(n5635) );
  XNOR U5804 ( .A(n5634), .B(n5635), .Z(n5512) );
  XOR U5805 ( .A(n5513), .B(n5512), .Z(n5515) );
  NAND U5806 ( .A(n5484), .B(n5483), .Z(n5488) );
  NANDN U5807 ( .A(n5486), .B(n5485), .Z(n5487) );
  AND U5808 ( .A(n5488), .B(n5487), .Z(n5506) );
  XNOR U5809 ( .A(n5507), .B(n5506), .Z(n5508) );
  XOR U5810 ( .A(n5509), .B(n5508), .Z(n5503) );
  XOR U5811 ( .A(n5502), .B(n5503), .Z(n5494) );
  XOR U5812 ( .A(n5495), .B(n5494), .Z(n5496) );
  XNOR U5813 ( .A(n5497), .B(n5496), .Z(n5638) );
  XNOR U5814 ( .A(n5638), .B(sreg[83]), .Z(n5640) );
  NAND U5815 ( .A(n5489), .B(sreg[82]), .Z(n5493) );
  OR U5816 ( .A(n5491), .B(n5490), .Z(n5492) );
  AND U5817 ( .A(n5493), .B(n5492), .Z(n5639) );
  XOR U5818 ( .A(n5640), .B(n5639), .Z(c[83]) );
  NAND U5819 ( .A(n5495), .B(n5494), .Z(n5499) );
  NAND U5820 ( .A(n5497), .B(n5496), .Z(n5498) );
  NAND U5821 ( .A(n5499), .B(n5498), .Z(n5646) );
  NANDN U5822 ( .A(n5501), .B(n5500), .Z(n5505) );
  NAND U5823 ( .A(n5503), .B(n5502), .Z(n5504) );
  NAND U5824 ( .A(n5505), .B(n5504), .Z(n5644) );
  NANDN U5825 ( .A(n5507), .B(n5506), .Z(n5511) );
  NAND U5826 ( .A(n5509), .B(n5508), .Z(n5510) );
  NAND U5827 ( .A(n5511), .B(n5510), .Z(n5649) );
  NANDN U5828 ( .A(n5513), .B(n5512), .Z(n5517) );
  OR U5829 ( .A(n5515), .B(n5514), .Z(n5516) );
  NAND U5830 ( .A(n5517), .B(n5516), .Z(n5650) );
  XNOR U5831 ( .A(n5649), .B(n5650), .Z(n5651) );
  NANDN U5832 ( .A(n5519), .B(n5518), .Z(n5523) );
  NAND U5833 ( .A(n5521), .B(n5520), .Z(n5522) );
  NAND U5834 ( .A(n5523), .B(n5522), .Z(n5718) );
  NAND U5835 ( .A(n5524), .B(n9379), .Z(n5526) );
  XNOR U5836 ( .A(n9562), .B(a[34]), .Z(n5661) );
  NAND U5837 ( .A(n5661), .B(n9378), .Z(n5525) );
  NAND U5838 ( .A(n5526), .B(n5525), .Z(n5729) );
  NANDN U5839 ( .A(n5527), .B(n9801), .Z(n5529) );
  XOR U5840 ( .A(b[27]), .B(n6500), .Z(n5664) );
  OR U5841 ( .A(n5664), .B(n9751), .Z(n5528) );
  NAND U5842 ( .A(n5529), .B(n5528), .Z(n5727) );
  XOR U5843 ( .A(a[48]), .B(n317), .Z(n5667) );
  NANDN U5844 ( .A(n5667), .B(n7905), .Z(n5532) );
  NANDN U5845 ( .A(n5530), .B(n7906), .Z(n5531) );
  AND U5846 ( .A(n5532), .B(n5531), .Z(n5728) );
  XNOR U5847 ( .A(n5727), .B(n5728), .Z(n5730) );
  XOR U5848 ( .A(n5729), .B(n5730), .Z(n5715) );
  NAND U5849 ( .A(n5533), .B(n9105), .Z(n5535) );
  XNOR U5850 ( .A(n9455), .B(a[36]), .Z(n5670) );
  NAND U5851 ( .A(n5670), .B(n9107), .Z(n5534) );
  NAND U5852 ( .A(n5535), .B(n5534), .Z(n5687) );
  NAND U5853 ( .A(n5536), .B(n9914), .Z(n5538) );
  XNOR U5854 ( .A(n323), .B(a[22]), .Z(n5673) );
  NANDN U5855 ( .A(n9913), .B(n5673), .Z(n5537) );
  NAND U5856 ( .A(n5538), .B(n5537), .Z(n5685) );
  NAND U5857 ( .A(n5539), .B(n7622), .Z(n5541) );
  XNOR U5858 ( .A(n9033), .B(b[3]), .Z(n5676) );
  NAND U5859 ( .A(n5676), .B(n7620), .Z(n5540) );
  NAND U5860 ( .A(n5541), .B(n5540), .Z(n5686) );
  XOR U5861 ( .A(n5685), .B(n5686), .Z(n5688) );
  XOR U5862 ( .A(n5687), .B(n5688), .Z(n5716) );
  XOR U5863 ( .A(n5715), .B(n5716), .Z(n5717) );
  XNOR U5864 ( .A(n5718), .B(n5717), .Z(n5763) );
  NANDN U5865 ( .A(n5543), .B(n5542), .Z(n5547) );
  NANDN U5866 ( .A(n5545), .B(n5544), .Z(n5546) );
  NAND U5867 ( .A(n5547), .B(n5546), .Z(n5706) );
  NAND U5868 ( .A(n5549), .B(n5548), .Z(n5553) );
  NAND U5869 ( .A(n5551), .B(n5550), .Z(n5552) );
  NAND U5870 ( .A(n5553), .B(n5552), .Z(n5704) );
  NANDN U5871 ( .A(n5555), .B(n5554), .Z(n5559) );
  NANDN U5872 ( .A(n5557), .B(n5556), .Z(n5558) );
  NAND U5873 ( .A(n5559), .B(n5558), .Z(n5703) );
  XNOR U5874 ( .A(n5706), .B(n5705), .Z(n5764) );
  XOR U5875 ( .A(n5763), .B(n5764), .Z(n5766) );
  NANDN U5876 ( .A(n5561), .B(n5560), .Z(n5565) );
  OR U5877 ( .A(n5563), .B(n5562), .Z(n5564) );
  NAND U5878 ( .A(n5565), .B(n5564), .Z(n5765) );
  XOR U5879 ( .A(n5766), .B(n5765), .Z(n5783) );
  OR U5880 ( .A(n5567), .B(n5566), .Z(n5571) );
  NAND U5881 ( .A(n5569), .B(n5568), .Z(n5570) );
  NAND U5882 ( .A(n5571), .B(n5570), .Z(n5782) );
  NANDN U5883 ( .A(n5573), .B(n5572), .Z(n5577) );
  NANDN U5884 ( .A(n5575), .B(n5574), .Z(n5576) );
  NAND U5885 ( .A(n5577), .B(n5576), .Z(n5771) );
  NAND U5886 ( .A(n5579), .B(n5578), .Z(n5583) );
  NAND U5887 ( .A(n5581), .B(n5580), .Z(n5582) );
  NAND U5888 ( .A(n5583), .B(n5582), .Z(n5770) );
  NANDN U5889 ( .A(n5585), .B(n5584), .Z(n5589) );
  NAND U5890 ( .A(n5587), .B(n5586), .Z(n5588) );
  NAND U5891 ( .A(n5589), .B(n5588), .Z(n5709) );
  NANDN U5892 ( .A(n5591), .B(n5590), .Z(n5595) );
  NAND U5893 ( .A(n5593), .B(n5592), .Z(n5594) );
  AND U5894 ( .A(n5595), .B(n5594), .Z(n5710) );
  XNOR U5895 ( .A(n5709), .B(n5710), .Z(n5711) );
  NAND U5896 ( .A(n5596), .B(n8286), .Z(n5598) );
  XNOR U5897 ( .A(n8444), .B(b[9]), .Z(n5733) );
  NAND U5898 ( .A(n5733), .B(n8288), .Z(n5597) );
  NAND U5899 ( .A(n5598), .B(n5597), .Z(n5693) );
  NAND U5900 ( .A(n5599), .B(n8961), .Z(n5601) );
  XNOR U5901 ( .A(b[15]), .B(n7672), .Z(n5736) );
  NAND U5902 ( .A(n5736), .B(n8963), .Z(n5600) );
  NAND U5903 ( .A(n5601), .B(n5600), .Z(n5691) );
  XNOR U5904 ( .A(b[21]), .B(a[32]), .Z(n5739) );
  NANDN U5905 ( .A(n5739), .B(n9493), .Z(n5604) );
  NANDN U5906 ( .A(n5602), .B(n9495), .Z(n5603) );
  AND U5907 ( .A(n5604), .B(n5603), .Z(n5692) );
  XOR U5908 ( .A(n5691), .B(n5692), .Z(n5694) );
  XNOR U5909 ( .A(n5693), .B(n5694), .Z(n5682) );
  XOR U5910 ( .A(b[11]), .B(n8156), .Z(n5742) );
  NANDN U5911 ( .A(n5742), .B(n8541), .Z(n5607) );
  NANDN U5912 ( .A(n5605), .B(n8542), .Z(n5606) );
  NAND U5913 ( .A(n5607), .B(n5606), .Z(n5680) );
  XOR U5914 ( .A(b[13]), .B(n7932), .Z(n5745) );
  NANDN U5915 ( .A(n5745), .B(n8730), .Z(n5610) );
  NANDN U5916 ( .A(n5608), .B(n8731), .Z(n5609) );
  AND U5917 ( .A(n5610), .B(n5609), .Z(n5679) );
  XNOR U5918 ( .A(n5680), .B(n5679), .Z(n5681) );
  XNOR U5919 ( .A(n5682), .B(n5681), .Z(n5699) );
  NANDN U5920 ( .A(n315), .B(a[52]), .Z(n5611) );
  XNOR U5921 ( .A(b[1]), .B(n5611), .Z(n5613) );
  IV U5922 ( .A(a[51]), .Z(n9457) );
  NANDN U5923 ( .A(n9457), .B(n315), .Z(n5612) );
  AND U5924 ( .A(n5613), .B(n5612), .Z(n5657) );
  NAND U5925 ( .A(n9875), .B(n5614), .Z(n5616) );
  XNOR U5926 ( .A(n322), .B(a[24]), .Z(n5751) );
  NANDN U5927 ( .A(n9874), .B(n5751), .Z(n5615) );
  NAND U5928 ( .A(n5616), .B(n5615), .Z(n5655) );
  NANDN U5929 ( .A(n323), .B(a[20]), .Z(n5656) );
  XNOR U5930 ( .A(n5655), .B(n5656), .Z(n5658) );
  XOR U5931 ( .A(n5657), .B(n5658), .Z(n5697) );
  NANDN U5932 ( .A(n5617), .B(n9622), .Z(n5619) );
  XOR U5933 ( .A(b[23]), .B(n6135), .Z(n5754) );
  OR U5934 ( .A(n5754), .B(n9621), .Z(n5618) );
  NAND U5935 ( .A(n5619), .B(n5618), .Z(n5724) );
  XNOR U5936 ( .A(a[46]), .B(b[7]), .Z(n5757) );
  OR U5937 ( .A(n5757), .B(n8013), .Z(n5622) );
  NAND U5938 ( .A(n5620), .B(n8014), .Z(n5621) );
  NAND U5939 ( .A(n5622), .B(n5621), .Z(n5721) );
  XNOR U5940 ( .A(b[25]), .B(a[28]), .Z(n5760) );
  NANDN U5941 ( .A(n5760), .B(n9706), .Z(n5625) );
  NANDN U5942 ( .A(n5623), .B(n9707), .Z(n5624) );
  AND U5943 ( .A(n5625), .B(n5624), .Z(n5722) );
  XNOR U5944 ( .A(n5721), .B(n5722), .Z(n5723) );
  XNOR U5945 ( .A(n5724), .B(n5723), .Z(n5698) );
  XOR U5946 ( .A(n5697), .B(n5698), .Z(n5700) );
  XNOR U5947 ( .A(n5699), .B(n5700), .Z(n5712) );
  XNOR U5948 ( .A(n5711), .B(n5712), .Z(n5769) );
  XNOR U5949 ( .A(n5770), .B(n5769), .Z(n5772) );
  XNOR U5950 ( .A(n5771), .B(n5772), .Z(n5781) );
  XOR U5951 ( .A(n5782), .B(n5781), .Z(n5784) );
  NANDN U5952 ( .A(n5627), .B(n5626), .Z(n5631) );
  OR U5953 ( .A(n5629), .B(n5628), .Z(n5630) );
  NAND U5954 ( .A(n5631), .B(n5630), .Z(n5775) );
  NAND U5955 ( .A(n5633), .B(n5632), .Z(n5637) );
  NANDN U5956 ( .A(n5635), .B(n5634), .Z(n5636) );
  NAND U5957 ( .A(n5637), .B(n5636), .Z(n5776) );
  XNOR U5958 ( .A(n5775), .B(n5776), .Z(n5777) );
  XOR U5959 ( .A(n5778), .B(n5777), .Z(n5652) );
  XOR U5960 ( .A(n5651), .B(n5652), .Z(n5643) );
  XOR U5961 ( .A(n5644), .B(n5643), .Z(n5645) );
  XNOR U5962 ( .A(n5646), .B(n5645), .Z(n5787) );
  XNOR U5963 ( .A(n5787), .B(sreg[84]), .Z(n5789) );
  NAND U5964 ( .A(n5638), .B(sreg[83]), .Z(n5642) );
  OR U5965 ( .A(n5640), .B(n5639), .Z(n5641) );
  AND U5966 ( .A(n5642), .B(n5641), .Z(n5788) );
  XOR U5967 ( .A(n5789), .B(n5788), .Z(c[84]) );
  NAND U5968 ( .A(n5644), .B(n5643), .Z(n5648) );
  NAND U5969 ( .A(n5646), .B(n5645), .Z(n5647) );
  NAND U5970 ( .A(n5648), .B(n5647), .Z(n5795) );
  NANDN U5971 ( .A(n5650), .B(n5649), .Z(n5654) );
  NAND U5972 ( .A(n5652), .B(n5651), .Z(n5653) );
  NAND U5973 ( .A(n5654), .B(n5653), .Z(n5793) );
  NANDN U5974 ( .A(n5656), .B(n5655), .Z(n5660) );
  NAND U5975 ( .A(n5658), .B(n5657), .Z(n5659) );
  NAND U5976 ( .A(n5660), .B(n5659), .Z(n5867) );
  NAND U5977 ( .A(n5661), .B(n9379), .Z(n5663) );
  XNOR U5978 ( .A(n9562), .B(a[35]), .Z(n5834) );
  NAND U5979 ( .A(n5834), .B(n9378), .Z(n5662) );
  NAND U5980 ( .A(n5663), .B(n5662), .Z(n5878) );
  NANDN U5981 ( .A(n5664), .B(n9801), .Z(n5666) );
  XNOR U5982 ( .A(b[27]), .B(a[27]), .Z(n5837) );
  OR U5983 ( .A(n5837), .B(n9751), .Z(n5665) );
  NAND U5984 ( .A(n5666), .B(n5665), .Z(n5876) );
  XNOR U5985 ( .A(a[49]), .B(b[5]), .Z(n5840) );
  NANDN U5986 ( .A(n5840), .B(n7905), .Z(n5669) );
  NANDN U5987 ( .A(n5667), .B(n7906), .Z(n5668) );
  AND U5988 ( .A(n5669), .B(n5668), .Z(n5877) );
  XNOR U5989 ( .A(n5876), .B(n5877), .Z(n5879) );
  XOR U5990 ( .A(n5878), .B(n5879), .Z(n5864) );
  NAND U5991 ( .A(n5670), .B(n9105), .Z(n5672) );
  XNOR U5992 ( .A(n9455), .B(a[37]), .Z(n5843) );
  NAND U5993 ( .A(n5843), .B(n9107), .Z(n5671) );
  AND U5994 ( .A(n5672), .B(n5671), .Z(n5819) );
  NAND U5995 ( .A(n5673), .B(n9914), .Z(n5675) );
  XNOR U5996 ( .A(n323), .B(a[23]), .Z(n5846) );
  NANDN U5997 ( .A(n9913), .B(n5846), .Z(n5674) );
  AND U5998 ( .A(n5675), .B(n5674), .Z(n5817) );
  NAND U5999 ( .A(n5676), .B(n7622), .Z(n5678) );
  XNOR U6000 ( .A(n9457), .B(b[3]), .Z(n5849) );
  NAND U6001 ( .A(n5849), .B(n7620), .Z(n5677) );
  NAND U6002 ( .A(n5678), .B(n5677), .Z(n5816) );
  XOR U6003 ( .A(n5864), .B(n5865), .Z(n5866) );
  XNOR U6004 ( .A(n5867), .B(n5866), .Z(n5912) );
  NANDN U6005 ( .A(n5680), .B(n5679), .Z(n5684) );
  NANDN U6006 ( .A(n5682), .B(n5681), .Z(n5683) );
  NAND U6007 ( .A(n5684), .B(n5683), .Z(n5855) );
  NAND U6008 ( .A(n5686), .B(n5685), .Z(n5690) );
  NAND U6009 ( .A(n5688), .B(n5687), .Z(n5689) );
  NAND U6010 ( .A(n5690), .B(n5689), .Z(n5853) );
  NANDN U6011 ( .A(n5692), .B(n5691), .Z(n5696) );
  NANDN U6012 ( .A(n5694), .B(n5693), .Z(n5695) );
  NAND U6013 ( .A(n5696), .B(n5695), .Z(n5852) );
  XNOR U6014 ( .A(n5855), .B(n5854), .Z(n5913) );
  XOR U6015 ( .A(n5912), .B(n5913), .Z(n5915) );
  NANDN U6016 ( .A(n5698), .B(n5697), .Z(n5702) );
  OR U6017 ( .A(n5700), .B(n5699), .Z(n5701) );
  NAND U6018 ( .A(n5702), .B(n5701), .Z(n5914) );
  XOR U6019 ( .A(n5915), .B(n5914), .Z(n5932) );
  OR U6020 ( .A(n5704), .B(n5703), .Z(n5708) );
  NAND U6021 ( .A(n5706), .B(n5705), .Z(n5707) );
  NAND U6022 ( .A(n5708), .B(n5707), .Z(n5931) );
  NANDN U6023 ( .A(n5710), .B(n5709), .Z(n5714) );
  NANDN U6024 ( .A(n5712), .B(n5711), .Z(n5713) );
  NAND U6025 ( .A(n5714), .B(n5713), .Z(n5920) );
  NAND U6026 ( .A(n5716), .B(n5715), .Z(n5720) );
  NAND U6027 ( .A(n5718), .B(n5717), .Z(n5719) );
  NAND U6028 ( .A(n5720), .B(n5719), .Z(n5919) );
  NANDN U6029 ( .A(n5722), .B(n5721), .Z(n5726) );
  NAND U6030 ( .A(n5724), .B(n5723), .Z(n5725) );
  NAND U6031 ( .A(n5726), .B(n5725), .Z(n5858) );
  NANDN U6032 ( .A(n5728), .B(n5727), .Z(n5732) );
  NAND U6033 ( .A(n5730), .B(n5729), .Z(n5731) );
  AND U6034 ( .A(n5732), .B(n5731), .Z(n5859) );
  XNOR U6035 ( .A(n5858), .B(n5859), .Z(n5860) );
  NAND U6036 ( .A(n5733), .B(n8286), .Z(n5735) );
  XOR U6037 ( .A(a[45]), .B(b[9]), .Z(n5882) );
  NAND U6038 ( .A(n5882), .B(n8288), .Z(n5734) );
  NAND U6039 ( .A(n5735), .B(n5734), .Z(n5824) );
  NAND U6040 ( .A(n5736), .B(n8961), .Z(n5738) );
  XOR U6041 ( .A(b[15]), .B(a[39]), .Z(n5885) );
  NAND U6042 ( .A(n5885), .B(n8963), .Z(n5737) );
  NAND U6043 ( .A(n5738), .B(n5737), .Z(n5822) );
  XOR U6044 ( .A(b[21]), .B(n6914), .Z(n5888) );
  NANDN U6045 ( .A(n5888), .B(n9493), .Z(n5741) );
  NANDN U6046 ( .A(n5739), .B(n9495), .Z(n5740) );
  AND U6047 ( .A(n5741), .B(n5740), .Z(n5823) );
  XOR U6048 ( .A(n5822), .B(n5823), .Z(n5825) );
  XNOR U6049 ( .A(n5824), .B(n5825), .Z(n5813) );
  XNOR U6050 ( .A(b[11]), .B(a[43]), .Z(n5891) );
  NANDN U6051 ( .A(n5891), .B(n8541), .Z(n5744) );
  NANDN U6052 ( .A(n5742), .B(n8542), .Z(n5743) );
  NAND U6053 ( .A(n5744), .B(n5743), .Z(n5811) );
  XNOR U6054 ( .A(b[13]), .B(a[41]), .Z(n5894) );
  NANDN U6055 ( .A(n5894), .B(n8730), .Z(n5747) );
  NANDN U6056 ( .A(n5745), .B(n8731), .Z(n5746) );
  NAND U6057 ( .A(n5747), .B(n5746), .Z(n5810) );
  XNOR U6058 ( .A(n5813), .B(n5812), .Z(n5807) );
  NANDN U6059 ( .A(n315), .B(a[53]), .Z(n5748) );
  XNOR U6060 ( .A(b[1]), .B(n5748), .Z(n5750) );
  IV U6061 ( .A(a[52]), .Z(n9217) );
  NANDN U6062 ( .A(n9217), .B(n315), .Z(n5749) );
  AND U6063 ( .A(n5750), .B(n5749), .Z(n5830) );
  NAND U6064 ( .A(n9875), .B(n5751), .Z(n5753) );
  XNOR U6065 ( .A(n322), .B(a[25]), .Z(n5900) );
  NANDN U6066 ( .A(n9874), .B(n5900), .Z(n5752) );
  NAND U6067 ( .A(n5753), .B(n5752), .Z(n5828) );
  NANDN U6068 ( .A(n323), .B(a[21]), .Z(n5829) );
  XNOR U6069 ( .A(n5828), .B(n5829), .Z(n5831) );
  XNOR U6070 ( .A(n5830), .B(n5831), .Z(n5805) );
  NANDN U6071 ( .A(n5754), .B(n9622), .Z(n5756) );
  XNOR U6072 ( .A(b[23]), .B(a[31]), .Z(n5903) );
  OR U6073 ( .A(n5903), .B(n9621), .Z(n5755) );
  NAND U6074 ( .A(n5756), .B(n5755), .Z(n5873) );
  XOR U6075 ( .A(a[47]), .B(b[7]), .Z(n5906) );
  NANDN U6076 ( .A(n8013), .B(n5906), .Z(n5759) );
  NANDN U6077 ( .A(n5757), .B(n8014), .Z(n5758) );
  NAND U6078 ( .A(n5759), .B(n5758), .Z(n5870) );
  XNOR U6079 ( .A(b[25]), .B(a[29]), .Z(n5909) );
  NANDN U6080 ( .A(n5909), .B(n9706), .Z(n5762) );
  NANDN U6081 ( .A(n5760), .B(n9707), .Z(n5761) );
  AND U6082 ( .A(n5762), .B(n5761), .Z(n5871) );
  XNOR U6083 ( .A(n5870), .B(n5871), .Z(n5872) );
  XOR U6084 ( .A(n5873), .B(n5872), .Z(n5804) );
  XOR U6085 ( .A(n5807), .B(n5806), .Z(n5861) );
  XNOR U6086 ( .A(n5860), .B(n5861), .Z(n5918) );
  XNOR U6087 ( .A(n5919), .B(n5918), .Z(n5921) );
  XNOR U6088 ( .A(n5920), .B(n5921), .Z(n5930) );
  XOR U6089 ( .A(n5931), .B(n5930), .Z(n5933) );
  NANDN U6090 ( .A(n5764), .B(n5763), .Z(n5768) );
  OR U6091 ( .A(n5766), .B(n5765), .Z(n5767) );
  NAND U6092 ( .A(n5768), .B(n5767), .Z(n5924) );
  NAND U6093 ( .A(n5770), .B(n5769), .Z(n5774) );
  NANDN U6094 ( .A(n5772), .B(n5771), .Z(n5773) );
  NAND U6095 ( .A(n5774), .B(n5773), .Z(n5925) );
  XNOR U6096 ( .A(n5924), .B(n5925), .Z(n5926) );
  XOR U6097 ( .A(n5927), .B(n5926), .Z(n5800) );
  NANDN U6098 ( .A(n5776), .B(n5775), .Z(n5780) );
  NAND U6099 ( .A(n5778), .B(n5777), .Z(n5779) );
  NAND U6100 ( .A(n5780), .B(n5779), .Z(n5798) );
  NANDN U6101 ( .A(n5782), .B(n5781), .Z(n5786) );
  OR U6102 ( .A(n5784), .B(n5783), .Z(n5785) );
  NAND U6103 ( .A(n5786), .B(n5785), .Z(n5799) );
  XNOR U6104 ( .A(n5798), .B(n5799), .Z(n5801) );
  XOR U6105 ( .A(n5800), .B(n5801), .Z(n5792) );
  XOR U6106 ( .A(n5793), .B(n5792), .Z(n5794) );
  XNOR U6107 ( .A(n5795), .B(n5794), .Z(n5936) );
  XNOR U6108 ( .A(n5936), .B(sreg[85]), .Z(n5938) );
  NAND U6109 ( .A(n5787), .B(sreg[84]), .Z(n5791) );
  OR U6110 ( .A(n5789), .B(n5788), .Z(n5790) );
  AND U6111 ( .A(n5791), .B(n5790), .Z(n5937) );
  XOR U6112 ( .A(n5938), .B(n5937), .Z(c[85]) );
  NAND U6113 ( .A(n5793), .B(n5792), .Z(n5797) );
  NAND U6114 ( .A(n5795), .B(n5794), .Z(n5796) );
  NAND U6115 ( .A(n5797), .B(n5796), .Z(n5944) );
  NANDN U6116 ( .A(n5799), .B(n5798), .Z(n5803) );
  NAND U6117 ( .A(n5801), .B(n5800), .Z(n5802) );
  NAND U6118 ( .A(n5803), .B(n5802), .Z(n5942) );
  NANDN U6119 ( .A(n5805), .B(n5804), .Z(n5809) );
  NANDN U6120 ( .A(n5807), .B(n5806), .Z(n5808) );
  NAND U6121 ( .A(n5809), .B(n5808), .Z(n6063) );
  OR U6122 ( .A(n5811), .B(n5810), .Z(n5815) );
  NANDN U6123 ( .A(n5813), .B(n5812), .Z(n5814) );
  NAND U6124 ( .A(n5815), .B(n5814), .Z(n6001) );
  NANDN U6125 ( .A(n5817), .B(n5816), .Z(n5821) );
  NANDN U6126 ( .A(n5819), .B(n5818), .Z(n5820) );
  NAND U6127 ( .A(n5821), .B(n5820), .Z(n6000) );
  NANDN U6128 ( .A(n5823), .B(n5822), .Z(n5827) );
  NANDN U6129 ( .A(n5825), .B(n5824), .Z(n5826) );
  NAND U6130 ( .A(n5827), .B(n5826), .Z(n5999) );
  XOR U6131 ( .A(n6001), .B(n6002), .Z(n6060) );
  NANDN U6132 ( .A(n5829), .B(n5828), .Z(n5833) );
  NAND U6133 ( .A(n5831), .B(n5830), .Z(n5832) );
  NAND U6134 ( .A(n5833), .B(n5832), .Z(n6014) );
  NAND U6135 ( .A(n5834), .B(n9379), .Z(n5836) );
  XNOR U6136 ( .A(n9562), .B(a[36]), .Z(n5957) );
  NAND U6137 ( .A(n5957), .B(n9378), .Z(n5835) );
  NAND U6138 ( .A(n5836), .B(n5835), .Z(n6025) );
  NANDN U6139 ( .A(n5837), .B(n9801), .Z(n5839) );
  XNOR U6140 ( .A(b[27]), .B(a[28]), .Z(n5960) );
  OR U6141 ( .A(n5960), .B(n9751), .Z(n5838) );
  NAND U6142 ( .A(n5839), .B(n5838), .Z(n6023) );
  XOR U6143 ( .A(a[50]), .B(n317), .Z(n5963) );
  NANDN U6144 ( .A(n5963), .B(n7905), .Z(n5842) );
  NANDN U6145 ( .A(n5840), .B(n7906), .Z(n5841) );
  AND U6146 ( .A(n5842), .B(n5841), .Z(n6024) );
  XNOR U6147 ( .A(n6023), .B(n6024), .Z(n6026) );
  XOR U6148 ( .A(n6025), .B(n6026), .Z(n6011) );
  NAND U6149 ( .A(n5843), .B(n9105), .Z(n5845) );
  XNOR U6150 ( .A(n9455), .B(a[38]), .Z(n5966) );
  NAND U6151 ( .A(n5966), .B(n9107), .Z(n5844) );
  NAND U6152 ( .A(n5845), .B(n5844), .Z(n5983) );
  NAND U6153 ( .A(n5846), .B(n9914), .Z(n5848) );
  XNOR U6154 ( .A(n323), .B(a[24]), .Z(n5969) );
  NANDN U6155 ( .A(n9913), .B(n5969), .Z(n5847) );
  NAND U6156 ( .A(n5848), .B(n5847), .Z(n5981) );
  NAND U6157 ( .A(n5849), .B(n7622), .Z(n5851) );
  XNOR U6158 ( .A(n9217), .B(b[3]), .Z(n5972) );
  NAND U6159 ( .A(n5972), .B(n7620), .Z(n5850) );
  NAND U6160 ( .A(n5851), .B(n5850), .Z(n5982) );
  XOR U6161 ( .A(n5981), .B(n5982), .Z(n5984) );
  XOR U6162 ( .A(n5983), .B(n5984), .Z(n6012) );
  XOR U6163 ( .A(n6011), .B(n6012), .Z(n6013) );
  XNOR U6164 ( .A(n6014), .B(n6013), .Z(n6061) );
  XNOR U6165 ( .A(n6060), .B(n6061), .Z(n6062) );
  XNOR U6166 ( .A(n6063), .B(n6062), .Z(n6081) );
  OR U6167 ( .A(n5853), .B(n5852), .Z(n5857) );
  NAND U6168 ( .A(n5855), .B(n5854), .Z(n5856) );
  NAND U6169 ( .A(n5857), .B(n5856), .Z(n6079) );
  NANDN U6170 ( .A(n5859), .B(n5858), .Z(n5863) );
  NANDN U6171 ( .A(n5861), .B(n5860), .Z(n5862) );
  NAND U6172 ( .A(n5863), .B(n5862), .Z(n6068) );
  NAND U6173 ( .A(n5865), .B(n5864), .Z(n5869) );
  NAND U6174 ( .A(n5867), .B(n5866), .Z(n5868) );
  NAND U6175 ( .A(n5869), .B(n5868), .Z(n6067) );
  NANDN U6176 ( .A(n5871), .B(n5870), .Z(n5875) );
  NAND U6177 ( .A(n5873), .B(n5872), .Z(n5874) );
  NAND U6178 ( .A(n5875), .B(n5874), .Z(n6005) );
  NANDN U6179 ( .A(n5877), .B(n5876), .Z(n5881) );
  NAND U6180 ( .A(n5879), .B(n5878), .Z(n5880) );
  AND U6181 ( .A(n5881), .B(n5880), .Z(n6006) );
  XNOR U6182 ( .A(n6005), .B(n6006), .Z(n6007) );
  NAND U6183 ( .A(n5882), .B(n8286), .Z(n5884) );
  XNOR U6184 ( .A(n8654), .B(b[9]), .Z(n6029) );
  NAND U6185 ( .A(n6029), .B(n8288), .Z(n5883) );
  NAND U6186 ( .A(n5884), .B(n5883), .Z(n5989) );
  NAND U6187 ( .A(n5885), .B(n8961), .Z(n5887) );
  XNOR U6188 ( .A(b[15]), .B(n7932), .Z(n6032) );
  NAND U6189 ( .A(n6032), .B(n8963), .Z(n5886) );
  NAND U6190 ( .A(n5887), .B(n5886), .Z(n5987) );
  XNOR U6191 ( .A(b[21]), .B(a[34]), .Z(n6035) );
  NANDN U6192 ( .A(n6035), .B(n9493), .Z(n5890) );
  NANDN U6193 ( .A(n5888), .B(n9495), .Z(n5889) );
  AND U6194 ( .A(n5890), .B(n5889), .Z(n5988) );
  XOR U6195 ( .A(n5987), .B(n5988), .Z(n5990) );
  XNOR U6196 ( .A(n5989), .B(n5990), .Z(n5978) );
  XOR U6197 ( .A(b[11]), .B(n8444), .Z(n6038) );
  NANDN U6198 ( .A(n6038), .B(n8541), .Z(n5893) );
  NANDN U6199 ( .A(n5891), .B(n8542), .Z(n5892) );
  NAND U6200 ( .A(n5893), .B(n5892), .Z(n5976) );
  XOR U6201 ( .A(b[13]), .B(n8156), .Z(n6041) );
  NANDN U6202 ( .A(n6041), .B(n8730), .Z(n5896) );
  NANDN U6203 ( .A(n5894), .B(n8731), .Z(n5895) );
  AND U6204 ( .A(n5896), .B(n5895), .Z(n5975) );
  XNOR U6205 ( .A(n5976), .B(n5975), .Z(n5977) );
  XNOR U6206 ( .A(n5978), .B(n5977), .Z(n5995) );
  NANDN U6207 ( .A(n315), .B(a[54]), .Z(n5897) );
  XNOR U6208 ( .A(b[1]), .B(n5897), .Z(n5899) );
  IV U6209 ( .A(a[53]), .Z(n9564) );
  NANDN U6210 ( .A(n9564), .B(n315), .Z(n5898) );
  AND U6211 ( .A(n5899), .B(n5898), .Z(n5953) );
  NAND U6212 ( .A(n9875), .B(n5900), .Z(n5902) );
  XOR U6213 ( .A(b[29]), .B(n6500), .Z(n6045) );
  OR U6214 ( .A(n6045), .B(n9874), .Z(n5901) );
  NAND U6215 ( .A(n5902), .B(n5901), .Z(n5951) );
  NANDN U6216 ( .A(n323), .B(a[22]), .Z(n5952) );
  XNOR U6217 ( .A(n5951), .B(n5952), .Z(n5954) );
  XOR U6218 ( .A(n5953), .B(n5954), .Z(n5993) );
  NANDN U6219 ( .A(n5903), .B(n9622), .Z(n5905) );
  XNOR U6220 ( .A(b[23]), .B(a[32]), .Z(n6051) );
  OR U6221 ( .A(n6051), .B(n9621), .Z(n5904) );
  NAND U6222 ( .A(n5905), .B(n5904), .Z(n6020) );
  XNOR U6223 ( .A(a[48]), .B(b[7]), .Z(n6054) );
  OR U6224 ( .A(n6054), .B(n8013), .Z(n5908) );
  NAND U6225 ( .A(n5906), .B(n8014), .Z(n5907) );
  NAND U6226 ( .A(n5908), .B(n5907), .Z(n6017) );
  XOR U6227 ( .A(b[25]), .B(n6135), .Z(n6057) );
  NANDN U6228 ( .A(n6057), .B(n9706), .Z(n5911) );
  NANDN U6229 ( .A(n5909), .B(n9707), .Z(n5910) );
  AND U6230 ( .A(n5911), .B(n5910), .Z(n6018) );
  XNOR U6231 ( .A(n6017), .B(n6018), .Z(n6019) );
  XNOR U6232 ( .A(n6020), .B(n6019), .Z(n5994) );
  XOR U6233 ( .A(n5993), .B(n5994), .Z(n5996) );
  XNOR U6234 ( .A(n5995), .B(n5996), .Z(n6008) );
  XNOR U6235 ( .A(n6007), .B(n6008), .Z(n6066) );
  XNOR U6236 ( .A(n6067), .B(n6066), .Z(n6069) );
  XNOR U6237 ( .A(n6068), .B(n6069), .Z(n6078) );
  XNOR U6238 ( .A(n6079), .B(n6078), .Z(n6080) );
  XOR U6239 ( .A(n6081), .B(n6080), .Z(n6075) );
  NANDN U6240 ( .A(n5913), .B(n5912), .Z(n5917) );
  OR U6241 ( .A(n5915), .B(n5914), .Z(n5916) );
  NAND U6242 ( .A(n5917), .B(n5916), .Z(n6072) );
  NAND U6243 ( .A(n5919), .B(n5918), .Z(n5923) );
  NANDN U6244 ( .A(n5921), .B(n5920), .Z(n5922) );
  NAND U6245 ( .A(n5923), .B(n5922), .Z(n6073) );
  XNOR U6246 ( .A(n6072), .B(n6073), .Z(n6074) );
  XNOR U6247 ( .A(n6075), .B(n6074), .Z(n5948) );
  NANDN U6248 ( .A(n5925), .B(n5924), .Z(n5929) );
  NAND U6249 ( .A(n5927), .B(n5926), .Z(n5928) );
  NAND U6250 ( .A(n5929), .B(n5928), .Z(n5945) );
  NANDN U6251 ( .A(n5931), .B(n5930), .Z(n5935) );
  OR U6252 ( .A(n5933), .B(n5932), .Z(n5934) );
  NAND U6253 ( .A(n5935), .B(n5934), .Z(n5946) );
  XNOR U6254 ( .A(n5945), .B(n5946), .Z(n5947) );
  XNOR U6255 ( .A(n5948), .B(n5947), .Z(n5941) );
  XOR U6256 ( .A(n5942), .B(n5941), .Z(n5943) );
  XNOR U6257 ( .A(n5944), .B(n5943), .Z(n6084) );
  XNOR U6258 ( .A(n6084), .B(sreg[86]), .Z(n6086) );
  NAND U6259 ( .A(n5936), .B(sreg[85]), .Z(n5940) );
  OR U6260 ( .A(n5938), .B(n5937), .Z(n5939) );
  AND U6261 ( .A(n5940), .B(n5939), .Z(n6085) );
  XOR U6262 ( .A(n6086), .B(n6085), .Z(c[86]) );
  NANDN U6263 ( .A(n5946), .B(n5945), .Z(n5950) );
  NANDN U6264 ( .A(n5948), .B(n5947), .Z(n5949) );
  NAND U6265 ( .A(n5950), .B(n5949), .Z(n6090) );
  NANDN U6266 ( .A(n5952), .B(n5951), .Z(n5956) );
  NAND U6267 ( .A(n5954), .B(n5953), .Z(n5955) );
  NAND U6268 ( .A(n5956), .B(n5955), .Z(n6165) );
  NAND U6269 ( .A(n5957), .B(n9379), .Z(n5959) );
  XNOR U6270 ( .A(n9562), .B(a[37]), .Z(n6131) );
  NAND U6271 ( .A(n6131), .B(n9378), .Z(n5958) );
  NAND U6272 ( .A(n5959), .B(n5958), .Z(n6176) );
  NANDN U6273 ( .A(n5960), .B(n9801), .Z(n5962) );
  XNOR U6274 ( .A(b[27]), .B(a[29]), .Z(n6134) );
  OR U6275 ( .A(n6134), .B(n9751), .Z(n5961) );
  NAND U6276 ( .A(n5962), .B(n5961), .Z(n6174) );
  XOR U6277 ( .A(a[51]), .B(n317), .Z(n6138) );
  NANDN U6278 ( .A(n6138), .B(n7905), .Z(n5965) );
  NANDN U6279 ( .A(n5963), .B(n7906), .Z(n5964) );
  AND U6280 ( .A(n5965), .B(n5964), .Z(n6175) );
  XNOR U6281 ( .A(n6174), .B(n6175), .Z(n6177) );
  XOR U6282 ( .A(n6176), .B(n6177), .Z(n6162) );
  NAND U6283 ( .A(n5966), .B(n9105), .Z(n5968) );
  XNOR U6284 ( .A(n9455), .B(a[39]), .Z(n6141) );
  NAND U6285 ( .A(n6141), .B(n9107), .Z(n5967) );
  AND U6286 ( .A(n5968), .B(n5967), .Z(n6116) );
  NAND U6287 ( .A(n5969), .B(n9914), .Z(n5971) );
  XNOR U6288 ( .A(n323), .B(a[25]), .Z(n6144) );
  NANDN U6289 ( .A(n9913), .B(n6144), .Z(n5970) );
  AND U6290 ( .A(n5971), .B(n5970), .Z(n6114) );
  NAND U6291 ( .A(n5972), .B(n7622), .Z(n5974) );
  XNOR U6292 ( .A(n9564), .B(b[3]), .Z(n6147) );
  NAND U6293 ( .A(n6147), .B(n7620), .Z(n5973) );
  NAND U6294 ( .A(n5974), .B(n5973), .Z(n6113) );
  XOR U6295 ( .A(n6162), .B(n6163), .Z(n6164) );
  XNOR U6296 ( .A(n6165), .B(n6164), .Z(n6210) );
  NANDN U6297 ( .A(n5976), .B(n5975), .Z(n5980) );
  NANDN U6298 ( .A(n5978), .B(n5977), .Z(n5979) );
  NAND U6299 ( .A(n5980), .B(n5979), .Z(n6153) );
  NAND U6300 ( .A(n5982), .B(n5981), .Z(n5986) );
  NAND U6301 ( .A(n5984), .B(n5983), .Z(n5985) );
  NAND U6302 ( .A(n5986), .B(n5985), .Z(n6151) );
  NANDN U6303 ( .A(n5988), .B(n5987), .Z(n5992) );
  NANDN U6304 ( .A(n5990), .B(n5989), .Z(n5991) );
  NAND U6305 ( .A(n5992), .B(n5991), .Z(n6150) );
  XNOR U6306 ( .A(n6153), .B(n6152), .Z(n6211) );
  XOR U6307 ( .A(n6210), .B(n6211), .Z(n6213) );
  NANDN U6308 ( .A(n5994), .B(n5993), .Z(n5998) );
  OR U6309 ( .A(n5996), .B(n5995), .Z(n5997) );
  NAND U6310 ( .A(n5998), .B(n5997), .Z(n6212) );
  XOR U6311 ( .A(n6213), .B(n6212), .Z(n6230) );
  OR U6312 ( .A(n6000), .B(n5999), .Z(n6004) );
  NANDN U6313 ( .A(n6002), .B(n6001), .Z(n6003) );
  NAND U6314 ( .A(n6004), .B(n6003), .Z(n6229) );
  NANDN U6315 ( .A(n6006), .B(n6005), .Z(n6010) );
  NANDN U6316 ( .A(n6008), .B(n6007), .Z(n6009) );
  NAND U6317 ( .A(n6010), .B(n6009), .Z(n6218) );
  NAND U6318 ( .A(n6012), .B(n6011), .Z(n6016) );
  NAND U6319 ( .A(n6014), .B(n6013), .Z(n6015) );
  NAND U6320 ( .A(n6016), .B(n6015), .Z(n6217) );
  NANDN U6321 ( .A(n6018), .B(n6017), .Z(n6022) );
  NAND U6322 ( .A(n6020), .B(n6019), .Z(n6021) );
  NAND U6323 ( .A(n6022), .B(n6021), .Z(n6156) );
  NANDN U6324 ( .A(n6024), .B(n6023), .Z(n6028) );
  NAND U6325 ( .A(n6026), .B(n6025), .Z(n6027) );
  AND U6326 ( .A(n6028), .B(n6027), .Z(n6157) );
  XNOR U6327 ( .A(n6156), .B(n6157), .Z(n6158) );
  NAND U6328 ( .A(n6029), .B(n8286), .Z(n6031) );
  XOR U6329 ( .A(a[47]), .B(b[9]), .Z(n6180) );
  NAND U6330 ( .A(n6180), .B(n8288), .Z(n6030) );
  NAND U6331 ( .A(n6031), .B(n6030), .Z(n6121) );
  NAND U6332 ( .A(n6032), .B(n8961), .Z(n6034) );
  XOR U6333 ( .A(b[15]), .B(a[41]), .Z(n6183) );
  NAND U6334 ( .A(n6183), .B(n8963), .Z(n6033) );
  NAND U6335 ( .A(n6034), .B(n6033), .Z(n6119) );
  XNOR U6336 ( .A(b[21]), .B(a[35]), .Z(n6186) );
  NANDN U6337 ( .A(n6186), .B(n9493), .Z(n6037) );
  NANDN U6338 ( .A(n6035), .B(n9495), .Z(n6036) );
  AND U6339 ( .A(n6037), .B(n6036), .Z(n6120) );
  XOR U6340 ( .A(n6119), .B(n6120), .Z(n6122) );
  XNOR U6341 ( .A(n6121), .B(n6122), .Z(n6110) );
  XNOR U6342 ( .A(b[11]), .B(a[45]), .Z(n6189) );
  NANDN U6343 ( .A(n6189), .B(n8541), .Z(n6040) );
  NANDN U6344 ( .A(n6038), .B(n8542), .Z(n6039) );
  NAND U6345 ( .A(n6040), .B(n6039), .Z(n6108) );
  XNOR U6346 ( .A(b[13]), .B(a[43]), .Z(n6192) );
  NANDN U6347 ( .A(n6192), .B(n8730), .Z(n6043) );
  NANDN U6348 ( .A(n6041), .B(n8731), .Z(n6042) );
  NAND U6349 ( .A(n6043), .B(n6042), .Z(n6107) );
  XNOR U6350 ( .A(n6110), .B(n6109), .Z(n6104) );
  ANDN U6351 ( .B(b[31]), .A(n6044), .Z(n6125) );
  NANDN U6352 ( .A(n6045), .B(n9875), .Z(n6047) );
  XNOR U6353 ( .A(n322), .B(a[27]), .Z(n6198) );
  NANDN U6354 ( .A(n9874), .B(n6198), .Z(n6046) );
  NAND U6355 ( .A(n6047), .B(n6046), .Z(n6126) );
  XOR U6356 ( .A(n6125), .B(n6126), .Z(n6127) );
  NANDN U6357 ( .A(n315), .B(a[55]), .Z(n6048) );
  XNOR U6358 ( .A(b[1]), .B(n6048), .Z(n6050) );
  IV U6359 ( .A(a[54]), .Z(n9353) );
  NANDN U6360 ( .A(n9353), .B(n315), .Z(n6049) );
  AND U6361 ( .A(n6050), .B(n6049), .Z(n6128) );
  XNOR U6362 ( .A(n6127), .B(n6128), .Z(n6101) );
  NANDN U6363 ( .A(n6051), .B(n9622), .Z(n6053) );
  XOR U6364 ( .A(b[23]), .B(n6914), .Z(n6201) );
  OR U6365 ( .A(n6201), .B(n9621), .Z(n6052) );
  NAND U6366 ( .A(n6053), .B(n6052), .Z(n6171) );
  XOR U6367 ( .A(a[49]), .B(b[7]), .Z(n6204) );
  NANDN U6368 ( .A(n8013), .B(n6204), .Z(n6056) );
  NANDN U6369 ( .A(n6054), .B(n8014), .Z(n6055) );
  NAND U6370 ( .A(n6056), .B(n6055), .Z(n6168) );
  XNOR U6371 ( .A(b[25]), .B(a[31]), .Z(n6207) );
  NANDN U6372 ( .A(n6207), .B(n9706), .Z(n6059) );
  NANDN U6373 ( .A(n6057), .B(n9707), .Z(n6058) );
  AND U6374 ( .A(n6059), .B(n6058), .Z(n6169) );
  XNOR U6375 ( .A(n6168), .B(n6169), .Z(n6170) );
  XNOR U6376 ( .A(n6171), .B(n6170), .Z(n6102) );
  XOR U6377 ( .A(n6104), .B(n6103), .Z(n6159) );
  XNOR U6378 ( .A(n6158), .B(n6159), .Z(n6216) );
  XNOR U6379 ( .A(n6217), .B(n6216), .Z(n6219) );
  XNOR U6380 ( .A(n6218), .B(n6219), .Z(n6228) );
  XOR U6381 ( .A(n6229), .B(n6228), .Z(n6231) );
  NANDN U6382 ( .A(n6061), .B(n6060), .Z(n6065) );
  NAND U6383 ( .A(n6063), .B(n6062), .Z(n6064) );
  NAND U6384 ( .A(n6065), .B(n6064), .Z(n6223) );
  NAND U6385 ( .A(n6067), .B(n6066), .Z(n6071) );
  NANDN U6386 ( .A(n6069), .B(n6068), .Z(n6070) );
  AND U6387 ( .A(n6071), .B(n6070), .Z(n6222) );
  XNOR U6388 ( .A(n6223), .B(n6222), .Z(n6224) );
  XOR U6389 ( .A(n6225), .B(n6224), .Z(n6097) );
  NANDN U6390 ( .A(n6073), .B(n6072), .Z(n6077) );
  NAND U6391 ( .A(n6075), .B(n6074), .Z(n6076) );
  NAND U6392 ( .A(n6077), .B(n6076), .Z(n6095) );
  NANDN U6393 ( .A(n6079), .B(n6078), .Z(n6083) );
  NANDN U6394 ( .A(n6081), .B(n6080), .Z(n6082) );
  NAND U6395 ( .A(n6083), .B(n6082), .Z(n6096) );
  XNOR U6396 ( .A(n6095), .B(n6096), .Z(n6098) );
  XOR U6397 ( .A(n6097), .B(n6098), .Z(n6089) );
  XOR U6398 ( .A(n6090), .B(n6089), .Z(n6091) );
  XNOR U6399 ( .A(n6092), .B(n6091), .Z(n6234) );
  XNOR U6400 ( .A(n6234), .B(sreg[87]), .Z(n6236) );
  NAND U6401 ( .A(n6084), .B(sreg[86]), .Z(n6088) );
  OR U6402 ( .A(n6086), .B(n6085), .Z(n6087) );
  AND U6403 ( .A(n6088), .B(n6087), .Z(n6235) );
  XOR U6404 ( .A(n6236), .B(n6235), .Z(c[87]) );
  NAND U6405 ( .A(n6090), .B(n6089), .Z(n6094) );
  NAND U6406 ( .A(n6092), .B(n6091), .Z(n6093) );
  NAND U6407 ( .A(n6094), .B(n6093), .Z(n6242) );
  NANDN U6408 ( .A(n6096), .B(n6095), .Z(n6100) );
  NAND U6409 ( .A(n6098), .B(n6097), .Z(n6099) );
  NAND U6410 ( .A(n6100), .B(n6099), .Z(n6240) );
  OR U6411 ( .A(n6102), .B(n6101), .Z(n6106) );
  NANDN U6412 ( .A(n6104), .B(n6103), .Z(n6105) );
  NAND U6413 ( .A(n6106), .B(n6105), .Z(n6360) );
  OR U6414 ( .A(n6108), .B(n6107), .Z(n6112) );
  NANDN U6415 ( .A(n6110), .B(n6109), .Z(n6111) );
  NAND U6416 ( .A(n6112), .B(n6111), .Z(n6299) );
  NANDN U6417 ( .A(n6114), .B(n6113), .Z(n6118) );
  NANDN U6418 ( .A(n6116), .B(n6115), .Z(n6117) );
  NAND U6419 ( .A(n6118), .B(n6117), .Z(n6298) );
  NANDN U6420 ( .A(n6120), .B(n6119), .Z(n6124) );
  NANDN U6421 ( .A(n6122), .B(n6121), .Z(n6123) );
  NAND U6422 ( .A(n6124), .B(n6123), .Z(n6297) );
  XOR U6423 ( .A(n6299), .B(n6300), .Z(n6358) );
  OR U6424 ( .A(n6126), .B(n6125), .Z(n6130) );
  NANDN U6425 ( .A(n6128), .B(n6127), .Z(n6129) );
  NAND U6426 ( .A(n6130), .B(n6129), .Z(n6312) );
  NAND U6427 ( .A(n6131), .B(n9379), .Z(n6133) );
  XNOR U6428 ( .A(n9562), .B(a[38]), .Z(n6279) );
  NAND U6429 ( .A(n6279), .B(n9378), .Z(n6132) );
  NAND U6430 ( .A(n6133), .B(n6132), .Z(n6323) );
  NANDN U6431 ( .A(n6134), .B(n9801), .Z(n6137) );
  XOR U6432 ( .A(b[27]), .B(n6135), .Z(n6282) );
  OR U6433 ( .A(n6282), .B(n9751), .Z(n6136) );
  NAND U6434 ( .A(n6137), .B(n6136), .Z(n6321) );
  XOR U6435 ( .A(a[52]), .B(n317), .Z(n6285) );
  NANDN U6436 ( .A(n6285), .B(n7905), .Z(n6140) );
  NANDN U6437 ( .A(n6138), .B(n7906), .Z(n6139) );
  AND U6438 ( .A(n6140), .B(n6139), .Z(n6322) );
  XNOR U6439 ( .A(n6321), .B(n6322), .Z(n6324) );
  XOR U6440 ( .A(n6323), .B(n6324), .Z(n6309) );
  NAND U6441 ( .A(n6141), .B(n9105), .Z(n6143) );
  XNOR U6442 ( .A(n9455), .B(a[40]), .Z(n6288) );
  NAND U6443 ( .A(n6288), .B(n9107), .Z(n6142) );
  AND U6444 ( .A(n6143), .B(n6142), .Z(n6264) );
  NAND U6445 ( .A(n6144), .B(n9914), .Z(n6146) );
  XNOR U6446 ( .A(n323), .B(a[26]), .Z(n6291) );
  NANDN U6447 ( .A(n9913), .B(n6291), .Z(n6145) );
  AND U6448 ( .A(n6146), .B(n6145), .Z(n6262) );
  NAND U6449 ( .A(n6147), .B(n7622), .Z(n6149) );
  XNOR U6450 ( .A(n9353), .B(b[3]), .Z(n6294) );
  NAND U6451 ( .A(n6294), .B(n7620), .Z(n6148) );
  NAND U6452 ( .A(n6149), .B(n6148), .Z(n6261) );
  XOR U6453 ( .A(n6309), .B(n6310), .Z(n6311) );
  XNOR U6454 ( .A(n6312), .B(n6311), .Z(n6357) );
  XOR U6455 ( .A(n6358), .B(n6357), .Z(n6359) );
  XNOR U6456 ( .A(n6360), .B(n6359), .Z(n6376) );
  OR U6457 ( .A(n6151), .B(n6150), .Z(n6155) );
  NAND U6458 ( .A(n6153), .B(n6152), .Z(n6154) );
  NAND U6459 ( .A(n6155), .B(n6154), .Z(n6374) );
  NANDN U6460 ( .A(n6157), .B(n6156), .Z(n6161) );
  NANDN U6461 ( .A(n6159), .B(n6158), .Z(n6160) );
  NAND U6462 ( .A(n6161), .B(n6160), .Z(n6363) );
  NAND U6463 ( .A(n6163), .B(n6162), .Z(n6167) );
  NAND U6464 ( .A(n6165), .B(n6164), .Z(n6166) );
  NAND U6465 ( .A(n6167), .B(n6166), .Z(n6362) );
  NANDN U6466 ( .A(n6169), .B(n6168), .Z(n6173) );
  NAND U6467 ( .A(n6171), .B(n6170), .Z(n6172) );
  NAND U6468 ( .A(n6173), .B(n6172), .Z(n6303) );
  NANDN U6469 ( .A(n6175), .B(n6174), .Z(n6179) );
  NAND U6470 ( .A(n6177), .B(n6176), .Z(n6178) );
  AND U6471 ( .A(n6179), .B(n6178), .Z(n6304) );
  XNOR U6472 ( .A(n6303), .B(n6304), .Z(n6305) );
  NAND U6473 ( .A(n6180), .B(n8286), .Z(n6182) );
  XNOR U6474 ( .A(n8837), .B(b[9]), .Z(n6327) );
  NAND U6475 ( .A(n6327), .B(n8288), .Z(n6181) );
  NAND U6476 ( .A(n6182), .B(n6181), .Z(n6269) );
  NAND U6477 ( .A(n6183), .B(n8961), .Z(n6185) );
  XNOR U6478 ( .A(b[15]), .B(n8156), .Z(n6330) );
  NAND U6479 ( .A(n6330), .B(n8963), .Z(n6184) );
  NAND U6480 ( .A(n6185), .B(n6184), .Z(n6267) );
  XOR U6481 ( .A(n318), .B(n7293), .Z(n6333) );
  NAND U6482 ( .A(n6333), .B(n9493), .Z(n6188) );
  NANDN U6483 ( .A(n6186), .B(n9495), .Z(n6187) );
  AND U6484 ( .A(n6188), .B(n6187), .Z(n6268) );
  XOR U6485 ( .A(n6267), .B(n6268), .Z(n6270) );
  XNOR U6486 ( .A(n6269), .B(n6270), .Z(n6258) );
  XOR U6487 ( .A(n8654), .B(b[11]), .Z(n6336) );
  NANDN U6488 ( .A(n6336), .B(n8541), .Z(n6191) );
  NANDN U6489 ( .A(n6189), .B(n8542), .Z(n6190) );
  NAND U6490 ( .A(n6191), .B(n6190), .Z(n6256) );
  XOR U6491 ( .A(b[13]), .B(n8444), .Z(n6339) );
  NANDN U6492 ( .A(n6339), .B(n8730), .Z(n6194) );
  NANDN U6493 ( .A(n6192), .B(n8731), .Z(n6193) );
  NAND U6494 ( .A(n6194), .B(n6193), .Z(n6255) );
  XNOR U6495 ( .A(n6258), .B(n6257), .Z(n6252) );
  NANDN U6496 ( .A(n315), .B(a[56]), .Z(n6195) );
  XNOR U6497 ( .A(b[1]), .B(n6195), .Z(n6197) );
  NANDN U6498 ( .A(b[0]), .B(a[55]), .Z(n6196) );
  AND U6499 ( .A(n6197), .B(n6196), .Z(n6275) );
  NAND U6500 ( .A(n6198), .B(n9875), .Z(n6200) );
  XNOR U6501 ( .A(n322), .B(a[28]), .Z(n6342) );
  NANDN U6502 ( .A(n9874), .B(n6342), .Z(n6199) );
  NAND U6503 ( .A(n6200), .B(n6199), .Z(n6273) );
  NANDN U6504 ( .A(n323), .B(a[24]), .Z(n6274) );
  XNOR U6505 ( .A(n6273), .B(n6274), .Z(n6276) );
  XNOR U6506 ( .A(n6275), .B(n6276), .Z(n6250) );
  NANDN U6507 ( .A(n6201), .B(n9622), .Z(n6203) );
  XNOR U6508 ( .A(b[23]), .B(a[34]), .Z(n6348) );
  OR U6509 ( .A(n6348), .B(n9621), .Z(n6202) );
  NAND U6510 ( .A(n6203), .B(n6202), .Z(n6318) );
  XNOR U6511 ( .A(a[50]), .B(b[7]), .Z(n6351) );
  OR U6512 ( .A(n6351), .B(n8013), .Z(n6206) );
  NAND U6513 ( .A(n6204), .B(n8014), .Z(n6205) );
  NAND U6514 ( .A(n6206), .B(n6205), .Z(n6315) );
  XNOR U6515 ( .A(b[25]), .B(a[32]), .Z(n6354) );
  NANDN U6516 ( .A(n6354), .B(n9706), .Z(n6209) );
  NANDN U6517 ( .A(n6207), .B(n9707), .Z(n6208) );
  AND U6518 ( .A(n6209), .B(n6208), .Z(n6316) );
  XNOR U6519 ( .A(n6315), .B(n6316), .Z(n6317) );
  XOR U6520 ( .A(n6318), .B(n6317), .Z(n6249) );
  XOR U6521 ( .A(n6252), .B(n6251), .Z(n6306) );
  XNOR U6522 ( .A(n6305), .B(n6306), .Z(n6361) );
  XNOR U6523 ( .A(n6362), .B(n6361), .Z(n6364) );
  XNOR U6524 ( .A(n6363), .B(n6364), .Z(n6373) );
  XNOR U6525 ( .A(n6374), .B(n6373), .Z(n6375) );
  XOR U6526 ( .A(n6376), .B(n6375), .Z(n6370) );
  NANDN U6527 ( .A(n6211), .B(n6210), .Z(n6215) );
  OR U6528 ( .A(n6213), .B(n6212), .Z(n6214) );
  NAND U6529 ( .A(n6215), .B(n6214), .Z(n6367) );
  NAND U6530 ( .A(n6217), .B(n6216), .Z(n6221) );
  NANDN U6531 ( .A(n6219), .B(n6218), .Z(n6220) );
  NAND U6532 ( .A(n6221), .B(n6220), .Z(n6368) );
  XNOR U6533 ( .A(n6367), .B(n6368), .Z(n6369) );
  XNOR U6534 ( .A(n6370), .B(n6369), .Z(n6246) );
  NANDN U6535 ( .A(n6223), .B(n6222), .Z(n6227) );
  NAND U6536 ( .A(n6225), .B(n6224), .Z(n6226) );
  NAND U6537 ( .A(n6227), .B(n6226), .Z(n6243) );
  NANDN U6538 ( .A(n6229), .B(n6228), .Z(n6233) );
  OR U6539 ( .A(n6231), .B(n6230), .Z(n6232) );
  NAND U6540 ( .A(n6233), .B(n6232), .Z(n6244) );
  XNOR U6541 ( .A(n6243), .B(n6244), .Z(n6245) );
  XNOR U6542 ( .A(n6246), .B(n6245), .Z(n6239) );
  XOR U6543 ( .A(n6240), .B(n6239), .Z(n6241) );
  XNOR U6544 ( .A(n6242), .B(n6241), .Z(n6379) );
  XNOR U6545 ( .A(n6379), .B(sreg[88]), .Z(n6381) );
  NAND U6546 ( .A(n6234), .B(sreg[87]), .Z(n6238) );
  OR U6547 ( .A(n6236), .B(n6235), .Z(n6237) );
  AND U6548 ( .A(n6238), .B(n6237), .Z(n6380) );
  XOR U6549 ( .A(n6381), .B(n6380), .Z(c[88]) );
  NANDN U6550 ( .A(n6244), .B(n6243), .Z(n6248) );
  NANDN U6551 ( .A(n6246), .B(n6245), .Z(n6247) );
  NAND U6552 ( .A(n6248), .B(n6247), .Z(n6385) );
  NANDN U6553 ( .A(n6250), .B(n6249), .Z(n6254) );
  NANDN U6554 ( .A(n6252), .B(n6251), .Z(n6253) );
  NAND U6555 ( .A(n6254), .B(n6253), .Z(n6516) );
  OR U6556 ( .A(n6256), .B(n6255), .Z(n6260) );
  NANDN U6557 ( .A(n6258), .B(n6257), .Z(n6259) );
  NAND U6558 ( .A(n6260), .B(n6259), .Z(n6454) );
  NANDN U6559 ( .A(n6262), .B(n6261), .Z(n6266) );
  NANDN U6560 ( .A(n6264), .B(n6263), .Z(n6265) );
  NAND U6561 ( .A(n6266), .B(n6265), .Z(n6453) );
  NANDN U6562 ( .A(n6268), .B(n6267), .Z(n6272) );
  NANDN U6563 ( .A(n6270), .B(n6269), .Z(n6271) );
  NAND U6564 ( .A(n6272), .B(n6271), .Z(n6452) );
  XOR U6565 ( .A(n6454), .B(n6455), .Z(n6513) );
  NANDN U6566 ( .A(n6274), .B(n6273), .Z(n6278) );
  NAND U6567 ( .A(n6276), .B(n6275), .Z(n6277) );
  NAND U6568 ( .A(n6278), .B(n6277), .Z(n6467) );
  NAND U6569 ( .A(n6279), .B(n9379), .Z(n6281) );
  XNOR U6570 ( .A(n9562), .B(a[39]), .Z(n6412) );
  NAND U6571 ( .A(n6412), .B(n9378), .Z(n6280) );
  NAND U6572 ( .A(n6281), .B(n6280), .Z(n6478) );
  NANDN U6573 ( .A(n6282), .B(n9801), .Z(n6284) );
  XNOR U6574 ( .A(b[27]), .B(a[31]), .Z(n6415) );
  OR U6575 ( .A(n6415), .B(n9751), .Z(n6283) );
  NAND U6576 ( .A(n6284), .B(n6283), .Z(n6476) );
  XOR U6577 ( .A(a[53]), .B(n317), .Z(n6418) );
  NANDN U6578 ( .A(n6418), .B(n7905), .Z(n6287) );
  NANDN U6579 ( .A(n6285), .B(n7906), .Z(n6286) );
  AND U6580 ( .A(n6287), .B(n6286), .Z(n6477) );
  XNOR U6581 ( .A(n6476), .B(n6477), .Z(n6479) );
  XOR U6582 ( .A(n6478), .B(n6479), .Z(n6464) );
  NAND U6583 ( .A(n6288), .B(n9105), .Z(n6290) );
  XNOR U6584 ( .A(n9455), .B(a[41]), .Z(n6421) );
  NAND U6585 ( .A(n6421), .B(n9107), .Z(n6289) );
  NAND U6586 ( .A(n6290), .B(n6289), .Z(n6438) );
  NAND U6587 ( .A(n6291), .B(n9914), .Z(n6293) );
  XNOR U6588 ( .A(n323), .B(a[27]), .Z(n6424) );
  NANDN U6589 ( .A(n9913), .B(n6424), .Z(n6292) );
  NAND U6590 ( .A(n6293), .B(n6292), .Z(n6436) );
  NAND U6591 ( .A(n6294), .B(n7622), .Z(n6296) );
  XNOR U6592 ( .A(a[55]), .B(n316), .Z(n6427) );
  NAND U6593 ( .A(n6427), .B(n7620), .Z(n6295) );
  NAND U6594 ( .A(n6296), .B(n6295), .Z(n6437) );
  XOR U6595 ( .A(n6436), .B(n6437), .Z(n6439) );
  XOR U6596 ( .A(n6438), .B(n6439), .Z(n6465) );
  XOR U6597 ( .A(n6464), .B(n6465), .Z(n6466) );
  XNOR U6598 ( .A(n6467), .B(n6466), .Z(n6514) );
  XNOR U6599 ( .A(n6513), .B(n6514), .Z(n6515) );
  XNOR U6600 ( .A(n6516), .B(n6515), .Z(n6403) );
  OR U6601 ( .A(n6298), .B(n6297), .Z(n6302) );
  NANDN U6602 ( .A(n6300), .B(n6299), .Z(n6301) );
  NAND U6603 ( .A(n6302), .B(n6301), .Z(n6401) );
  NANDN U6604 ( .A(n6304), .B(n6303), .Z(n6308) );
  NANDN U6605 ( .A(n6306), .B(n6305), .Z(n6307) );
  NAND U6606 ( .A(n6308), .B(n6307), .Z(n6521) );
  NAND U6607 ( .A(n6310), .B(n6309), .Z(n6314) );
  NANDN U6608 ( .A(n6312), .B(n6311), .Z(n6313) );
  NAND U6609 ( .A(n6314), .B(n6313), .Z(n6520) );
  NANDN U6610 ( .A(n6316), .B(n6315), .Z(n6320) );
  NAND U6611 ( .A(n6318), .B(n6317), .Z(n6319) );
  NAND U6612 ( .A(n6320), .B(n6319), .Z(n6458) );
  NANDN U6613 ( .A(n6322), .B(n6321), .Z(n6326) );
  NAND U6614 ( .A(n6324), .B(n6323), .Z(n6325) );
  AND U6615 ( .A(n6326), .B(n6325), .Z(n6459) );
  XNOR U6616 ( .A(n6458), .B(n6459), .Z(n6460) );
  NAND U6617 ( .A(n6327), .B(n8286), .Z(n6329) );
  XOR U6618 ( .A(a[49]), .B(b[9]), .Z(n6488) );
  NAND U6619 ( .A(n6488), .B(n8288), .Z(n6328) );
  NAND U6620 ( .A(n6329), .B(n6328), .Z(n6444) );
  NAND U6621 ( .A(n6330), .B(n8961), .Z(n6332) );
  XOR U6622 ( .A(b[15]), .B(a[43]), .Z(n6482) );
  NAND U6623 ( .A(n6482), .B(n8963), .Z(n6331) );
  NAND U6624 ( .A(n6332), .B(n6331), .Z(n6443) );
  XNOR U6625 ( .A(b[21]), .B(a[37]), .Z(n6485) );
  NANDN U6626 ( .A(n6485), .B(n9493), .Z(n6335) );
  NAND U6627 ( .A(n9495), .B(n6333), .Z(n6334) );
  NAND U6628 ( .A(n6335), .B(n6334), .Z(n6442) );
  XNOR U6629 ( .A(n6443), .B(n6442), .Z(n6445) );
  XNOR U6630 ( .A(n6444), .B(n6445), .Z(n6433) );
  XNOR U6631 ( .A(a[47]), .B(b[11]), .Z(n6491) );
  NANDN U6632 ( .A(n6491), .B(n8541), .Z(n6338) );
  NANDN U6633 ( .A(n6336), .B(n8542), .Z(n6337) );
  NAND U6634 ( .A(n6338), .B(n6337), .Z(n6431) );
  XNOR U6635 ( .A(b[13]), .B(a[45]), .Z(n6494) );
  NANDN U6636 ( .A(n6494), .B(n8730), .Z(n6341) );
  NANDN U6637 ( .A(n6339), .B(n8731), .Z(n6340) );
  AND U6638 ( .A(n6341), .B(n6340), .Z(n6430) );
  XNOR U6639 ( .A(n6431), .B(n6430), .Z(n6432) );
  XNOR U6640 ( .A(n6433), .B(n6432), .Z(n6449) );
  NAND U6641 ( .A(n9875), .B(n6342), .Z(n6344) );
  XNOR U6642 ( .A(b[29]), .B(a[29]), .Z(n6501) );
  OR U6643 ( .A(n6501), .B(n9874), .Z(n6343) );
  NAND U6644 ( .A(n6344), .B(n6343), .Z(n6406) );
  NANDN U6645 ( .A(n323), .B(a[25]), .Z(n6407) );
  XNOR U6646 ( .A(n6406), .B(n6407), .Z(n6409) );
  NANDN U6647 ( .A(n315), .B(a[57]), .Z(n6345) );
  XNOR U6648 ( .A(b[1]), .B(n6345), .Z(n6347) );
  IV U6649 ( .A(a[56]), .Z(n9357) );
  NANDN U6650 ( .A(n9357), .B(n315), .Z(n6346) );
  AND U6651 ( .A(n6347), .B(n6346), .Z(n6408) );
  XNOR U6652 ( .A(n6409), .B(n6408), .Z(n6447) );
  NANDN U6653 ( .A(n6348), .B(n9622), .Z(n6350) );
  XNOR U6654 ( .A(b[23]), .B(a[35]), .Z(n6504) );
  OR U6655 ( .A(n6504), .B(n9621), .Z(n6349) );
  NAND U6656 ( .A(n6350), .B(n6349), .Z(n6473) );
  XNOR U6657 ( .A(a[51]), .B(b[7]), .Z(n6507) );
  OR U6658 ( .A(n6507), .B(n8013), .Z(n6353) );
  NANDN U6659 ( .A(n6351), .B(n8014), .Z(n6352) );
  NAND U6660 ( .A(n6353), .B(n6352), .Z(n6470) );
  XOR U6661 ( .A(b[25]), .B(n6914), .Z(n6510) );
  NANDN U6662 ( .A(n6510), .B(n9706), .Z(n6356) );
  NANDN U6663 ( .A(n6354), .B(n9707), .Z(n6355) );
  AND U6664 ( .A(n6356), .B(n6355), .Z(n6471) );
  XNOR U6665 ( .A(n6470), .B(n6471), .Z(n6472) );
  XOR U6666 ( .A(n6473), .B(n6472), .Z(n6446) );
  XOR U6667 ( .A(n6449), .B(n6448), .Z(n6461) );
  XNOR U6668 ( .A(n6460), .B(n6461), .Z(n6519) );
  XNOR U6669 ( .A(n6520), .B(n6519), .Z(n6522) );
  XNOR U6670 ( .A(n6521), .B(n6522), .Z(n6400) );
  XNOR U6671 ( .A(n6401), .B(n6400), .Z(n6402) );
  XOR U6672 ( .A(n6403), .B(n6402), .Z(n6397) );
  NAND U6673 ( .A(n6362), .B(n6361), .Z(n6366) );
  NANDN U6674 ( .A(n6364), .B(n6363), .Z(n6365) );
  AND U6675 ( .A(n6366), .B(n6365), .Z(n6394) );
  XNOR U6676 ( .A(n6395), .B(n6394), .Z(n6396) );
  XNOR U6677 ( .A(n6397), .B(n6396), .Z(n6391) );
  NANDN U6678 ( .A(n6368), .B(n6367), .Z(n6372) );
  NAND U6679 ( .A(n6370), .B(n6369), .Z(n6371) );
  NAND U6680 ( .A(n6372), .B(n6371), .Z(n6388) );
  NANDN U6681 ( .A(n6374), .B(n6373), .Z(n6378) );
  NANDN U6682 ( .A(n6376), .B(n6375), .Z(n6377) );
  NAND U6683 ( .A(n6378), .B(n6377), .Z(n6389) );
  XNOR U6684 ( .A(n6388), .B(n6389), .Z(n6390) );
  XNOR U6685 ( .A(n6391), .B(n6390), .Z(n6384) );
  XOR U6686 ( .A(n6385), .B(n6384), .Z(n6386) );
  XNOR U6687 ( .A(n6387), .B(n6386), .Z(n6525) );
  XNOR U6688 ( .A(n6525), .B(sreg[89]), .Z(n6527) );
  NAND U6689 ( .A(n6379), .B(sreg[88]), .Z(n6383) );
  OR U6690 ( .A(n6381), .B(n6380), .Z(n6382) );
  AND U6691 ( .A(n6383), .B(n6382), .Z(n6526) );
  XOR U6692 ( .A(n6527), .B(n6526), .Z(c[89]) );
  NANDN U6693 ( .A(n6389), .B(n6388), .Z(n6393) );
  NANDN U6694 ( .A(n6391), .B(n6390), .Z(n6392) );
  NAND U6695 ( .A(n6393), .B(n6392), .Z(n6531) );
  NANDN U6696 ( .A(n6395), .B(n6394), .Z(n6399) );
  NAND U6697 ( .A(n6397), .B(n6396), .Z(n6398) );
  NAND U6698 ( .A(n6399), .B(n6398), .Z(n6536) );
  NANDN U6699 ( .A(n6401), .B(n6400), .Z(n6405) );
  NANDN U6700 ( .A(n6403), .B(n6402), .Z(n6404) );
  NAND U6701 ( .A(n6405), .B(n6404), .Z(n6537) );
  XNOR U6702 ( .A(n6536), .B(n6537), .Z(n6538) );
  NANDN U6703 ( .A(n6407), .B(n6406), .Z(n6411) );
  NAND U6704 ( .A(n6409), .B(n6408), .Z(n6410) );
  NAND U6705 ( .A(n6411), .B(n6410), .Z(n6613) );
  NAND U6706 ( .A(n6412), .B(n9379), .Z(n6414) );
  XNOR U6707 ( .A(n9562), .B(a[40]), .Z(n6558) );
  NAND U6708 ( .A(n6558), .B(n9378), .Z(n6413) );
  NAND U6709 ( .A(n6414), .B(n6413), .Z(n6624) );
  NANDN U6710 ( .A(n6415), .B(n9801), .Z(n6417) );
  XNOR U6711 ( .A(b[27]), .B(a[32]), .Z(n6561) );
  OR U6712 ( .A(n6561), .B(n9751), .Z(n6416) );
  NAND U6713 ( .A(n6417), .B(n6416), .Z(n6622) );
  XOR U6714 ( .A(a[54]), .B(n317), .Z(n6564) );
  NANDN U6715 ( .A(n6564), .B(n7905), .Z(n6420) );
  NANDN U6716 ( .A(n6418), .B(n7906), .Z(n6419) );
  AND U6717 ( .A(n6420), .B(n6419), .Z(n6623) );
  XNOR U6718 ( .A(n6622), .B(n6623), .Z(n6625) );
  XOR U6719 ( .A(n6624), .B(n6625), .Z(n6610) );
  NAND U6720 ( .A(n6421), .B(n9105), .Z(n6423) );
  XNOR U6721 ( .A(n9455), .B(a[42]), .Z(n6567) );
  NAND U6722 ( .A(n6567), .B(n9107), .Z(n6422) );
  NAND U6723 ( .A(n6423), .B(n6422), .Z(n6584) );
  NAND U6724 ( .A(n6424), .B(n9914), .Z(n6426) );
  XNOR U6725 ( .A(n323), .B(a[28]), .Z(n6570) );
  NANDN U6726 ( .A(n9913), .B(n6570), .Z(n6425) );
  NAND U6727 ( .A(n6426), .B(n6425), .Z(n6582) );
  NAND U6728 ( .A(n6427), .B(n7622), .Z(n6429) );
  XNOR U6729 ( .A(n9357), .B(b[3]), .Z(n6573) );
  NAND U6730 ( .A(n6573), .B(n7620), .Z(n6428) );
  NAND U6731 ( .A(n6429), .B(n6428), .Z(n6583) );
  XOR U6732 ( .A(n6582), .B(n6583), .Z(n6585) );
  XOR U6733 ( .A(n6584), .B(n6585), .Z(n6611) );
  XOR U6734 ( .A(n6610), .B(n6611), .Z(n6612) );
  XNOR U6735 ( .A(n6613), .B(n6612), .Z(n6549) );
  NANDN U6736 ( .A(n6431), .B(n6430), .Z(n6435) );
  NANDN U6737 ( .A(n6433), .B(n6432), .Z(n6434) );
  NAND U6738 ( .A(n6435), .B(n6434), .Z(n6602) );
  NAND U6739 ( .A(n6437), .B(n6436), .Z(n6441) );
  NAND U6740 ( .A(n6439), .B(n6438), .Z(n6440) );
  NAND U6741 ( .A(n6441), .B(n6440), .Z(n6601) );
  XNOR U6742 ( .A(n6601), .B(n6600), .Z(n6603) );
  XOR U6743 ( .A(n6602), .B(n6603), .Z(n6548) );
  XOR U6744 ( .A(n6549), .B(n6548), .Z(n6550) );
  NANDN U6745 ( .A(n6447), .B(n6446), .Z(n6451) );
  NANDN U6746 ( .A(n6449), .B(n6448), .Z(n6450) );
  NAND U6747 ( .A(n6451), .B(n6450), .Z(n6551) );
  XNOR U6748 ( .A(n6550), .B(n6551), .Z(n6666) );
  OR U6749 ( .A(n6453), .B(n6452), .Z(n6457) );
  NANDN U6750 ( .A(n6455), .B(n6454), .Z(n6456) );
  NAND U6751 ( .A(n6457), .B(n6456), .Z(n6665) );
  NANDN U6752 ( .A(n6459), .B(n6458), .Z(n6463) );
  NANDN U6753 ( .A(n6461), .B(n6460), .Z(n6462) );
  NAND U6754 ( .A(n6463), .B(n6462), .Z(n6544) );
  NAND U6755 ( .A(n6465), .B(n6464), .Z(n6469) );
  NAND U6756 ( .A(n6467), .B(n6466), .Z(n6468) );
  NAND U6757 ( .A(n6469), .B(n6468), .Z(n6543) );
  NANDN U6758 ( .A(n6471), .B(n6470), .Z(n6475) );
  NAND U6759 ( .A(n6473), .B(n6472), .Z(n6474) );
  NAND U6760 ( .A(n6475), .B(n6474), .Z(n6604) );
  NANDN U6761 ( .A(n6477), .B(n6476), .Z(n6481) );
  NAND U6762 ( .A(n6479), .B(n6478), .Z(n6480) );
  AND U6763 ( .A(n6481), .B(n6480), .Z(n6605) );
  XNOR U6764 ( .A(n6604), .B(n6605), .Z(n6606) );
  NAND U6765 ( .A(n6482), .B(n8961), .Z(n6484) );
  XNOR U6766 ( .A(b[15]), .B(n8444), .Z(n6631) );
  NAND U6767 ( .A(n6631), .B(n8963), .Z(n6483) );
  NAND U6768 ( .A(n6484), .B(n6483), .Z(n6594) );
  XOR U6769 ( .A(b[21]), .B(n7672), .Z(n6634) );
  NANDN U6770 ( .A(n6634), .B(n9493), .Z(n6487) );
  NANDN U6771 ( .A(n6485), .B(n9495), .Z(n6486) );
  AND U6772 ( .A(n6487), .B(n6486), .Z(n6595) );
  XOR U6773 ( .A(n6594), .B(n6595), .Z(n6597) );
  NAND U6774 ( .A(n6488), .B(n8286), .Z(n6490) );
  XNOR U6775 ( .A(n9033), .B(b[9]), .Z(n6628) );
  NAND U6776 ( .A(n6628), .B(n8288), .Z(n6489) );
  NAND U6777 ( .A(n6490), .B(n6489), .Z(n6596) );
  XNOR U6778 ( .A(n6597), .B(n6596), .Z(n6591) );
  XOR U6779 ( .A(n8837), .B(b[11]), .Z(n6637) );
  NANDN U6780 ( .A(n6637), .B(n8541), .Z(n6493) );
  NANDN U6781 ( .A(n6491), .B(n8542), .Z(n6492) );
  NAND U6782 ( .A(n6493), .B(n6492), .Z(n6589) );
  XOR U6783 ( .A(b[13]), .B(n8654), .Z(n6640) );
  NANDN U6784 ( .A(n6640), .B(n8730), .Z(n6496) );
  NANDN U6785 ( .A(n6494), .B(n8731), .Z(n6495) );
  NAND U6786 ( .A(n6496), .B(n6495), .Z(n6588) );
  XNOR U6787 ( .A(n6589), .B(n6588), .Z(n6590) );
  XOR U6788 ( .A(n6591), .B(n6590), .Z(n6579) );
  NANDN U6789 ( .A(n315), .B(a[58]), .Z(n6497) );
  XNOR U6790 ( .A(b[1]), .B(n6497), .Z(n6499) );
  NANDN U6791 ( .A(b[0]), .B(a[57]), .Z(n6498) );
  AND U6792 ( .A(n6499), .B(n6498), .Z(n6555) );
  ANDN U6793 ( .B(b[31]), .A(n6500), .Z(n6552) );
  NANDN U6794 ( .A(n6501), .B(n9875), .Z(n6503) );
  XNOR U6795 ( .A(n322), .B(a[30]), .Z(n6643) );
  NANDN U6796 ( .A(n9874), .B(n6643), .Z(n6502) );
  NAND U6797 ( .A(n6503), .B(n6502), .Z(n6553) );
  XOR U6798 ( .A(n6552), .B(n6553), .Z(n6554) );
  XNOR U6799 ( .A(n6555), .B(n6554), .Z(n6576) );
  NANDN U6800 ( .A(n6504), .B(n9622), .Z(n6506) );
  XOR U6801 ( .A(b[23]), .B(n7293), .Z(n6649) );
  OR U6802 ( .A(n6649), .B(n9621), .Z(n6505) );
  NAND U6803 ( .A(n6506), .B(n6505), .Z(n6619) );
  XNOR U6804 ( .A(a[52]), .B(b[7]), .Z(n6652) );
  OR U6805 ( .A(n6652), .B(n8013), .Z(n6509) );
  NANDN U6806 ( .A(n6507), .B(n8014), .Z(n6508) );
  NAND U6807 ( .A(n6509), .B(n6508), .Z(n6616) );
  XNOR U6808 ( .A(b[25]), .B(a[34]), .Z(n6655) );
  NANDN U6809 ( .A(n6655), .B(n9706), .Z(n6512) );
  NANDN U6810 ( .A(n6510), .B(n9707), .Z(n6511) );
  AND U6811 ( .A(n6512), .B(n6511), .Z(n6617) );
  XNOR U6812 ( .A(n6616), .B(n6617), .Z(n6618) );
  XNOR U6813 ( .A(n6619), .B(n6618), .Z(n6577) );
  XOR U6814 ( .A(n6579), .B(n6578), .Z(n6607) );
  XNOR U6815 ( .A(n6606), .B(n6607), .Z(n6542) );
  XNOR U6816 ( .A(n6543), .B(n6542), .Z(n6545) );
  XNOR U6817 ( .A(n6544), .B(n6545), .Z(n6664) );
  XOR U6818 ( .A(n6665), .B(n6664), .Z(n6667) );
  NANDN U6819 ( .A(n6514), .B(n6513), .Z(n6518) );
  NAND U6820 ( .A(n6516), .B(n6515), .Z(n6517) );
  NAND U6821 ( .A(n6518), .B(n6517), .Z(n6659) );
  NAND U6822 ( .A(n6520), .B(n6519), .Z(n6524) );
  NANDN U6823 ( .A(n6522), .B(n6521), .Z(n6523) );
  AND U6824 ( .A(n6524), .B(n6523), .Z(n6658) );
  XNOR U6825 ( .A(n6659), .B(n6658), .Z(n6660) );
  XOR U6826 ( .A(n6661), .B(n6660), .Z(n6539) );
  XOR U6827 ( .A(n6538), .B(n6539), .Z(n6530) );
  XOR U6828 ( .A(n6531), .B(n6530), .Z(n6532) );
  XNOR U6829 ( .A(n6533), .B(n6532), .Z(n6670) );
  XNOR U6830 ( .A(n6670), .B(sreg[90]), .Z(n6672) );
  NAND U6831 ( .A(n6525), .B(sreg[89]), .Z(n6529) );
  OR U6832 ( .A(n6527), .B(n6526), .Z(n6528) );
  AND U6833 ( .A(n6529), .B(n6528), .Z(n6671) );
  XOR U6834 ( .A(n6672), .B(n6671), .Z(c[90]) );
  NAND U6835 ( .A(n6531), .B(n6530), .Z(n6535) );
  NAND U6836 ( .A(n6533), .B(n6532), .Z(n6534) );
  NAND U6837 ( .A(n6535), .B(n6534), .Z(n6678) );
  NANDN U6838 ( .A(n6537), .B(n6536), .Z(n6541) );
  NAND U6839 ( .A(n6539), .B(n6538), .Z(n6540) );
  NAND U6840 ( .A(n6541), .B(n6540), .Z(n6675) );
  NAND U6841 ( .A(n6543), .B(n6542), .Z(n6547) );
  NANDN U6842 ( .A(n6545), .B(n6544), .Z(n6546) );
  NAND U6843 ( .A(n6547), .B(n6546), .Z(n6805) );
  XNOR U6844 ( .A(n6805), .B(n6806), .Z(n6807) );
  OR U6845 ( .A(n6553), .B(n6552), .Z(n6557) );
  NANDN U6846 ( .A(n6555), .B(n6554), .Z(n6556) );
  NAND U6847 ( .A(n6557), .B(n6556), .Z(n6748) );
  NAND U6848 ( .A(n6558), .B(n9379), .Z(n6560) );
  XNOR U6849 ( .A(n9562), .B(a[41]), .Z(n6720) );
  NAND U6850 ( .A(n6720), .B(n9378), .Z(n6559) );
  NAND U6851 ( .A(n6560), .B(n6559), .Z(n6789) );
  NANDN U6852 ( .A(n6561), .B(n9801), .Z(n6563) );
  XOR U6853 ( .A(b[27]), .B(n6914), .Z(n6717) );
  OR U6854 ( .A(n6717), .B(n9751), .Z(n6562) );
  NAND U6855 ( .A(n6563), .B(n6562), .Z(n6787) );
  XNOR U6856 ( .A(a[55]), .B(b[5]), .Z(n6723) );
  NANDN U6857 ( .A(n6723), .B(n7905), .Z(n6566) );
  NANDN U6858 ( .A(n6564), .B(n7906), .Z(n6565) );
  AND U6859 ( .A(n6566), .B(n6565), .Z(n6788) );
  XNOR U6860 ( .A(n6787), .B(n6788), .Z(n6790) );
  XOR U6861 ( .A(n6789), .B(n6790), .Z(n6745) );
  NAND U6862 ( .A(n6567), .B(n9105), .Z(n6569) );
  XNOR U6863 ( .A(n9455), .B(a[43]), .Z(n6726) );
  NAND U6864 ( .A(n6726), .B(n9107), .Z(n6568) );
  AND U6865 ( .A(n6569), .B(n6568), .Z(n6702) );
  NAND U6866 ( .A(n6570), .B(n9914), .Z(n6572) );
  XNOR U6867 ( .A(n323), .B(a[29]), .Z(n6729) );
  NANDN U6868 ( .A(n9913), .B(n6729), .Z(n6571) );
  AND U6869 ( .A(n6572), .B(n6571), .Z(n6700) );
  NAND U6870 ( .A(n6573), .B(n7622), .Z(n6575) );
  XNOR U6871 ( .A(a[57]), .B(n316), .Z(n6732) );
  NAND U6872 ( .A(n6732), .B(n7620), .Z(n6574) );
  NAND U6873 ( .A(n6575), .B(n6574), .Z(n6699) );
  XOR U6874 ( .A(n6745), .B(n6746), .Z(n6747) );
  XOR U6875 ( .A(n6748), .B(n6747), .Z(n6799) );
  OR U6876 ( .A(n6577), .B(n6576), .Z(n6581) );
  NANDN U6877 ( .A(n6579), .B(n6578), .Z(n6580) );
  NAND U6878 ( .A(n6581), .B(n6580), .Z(n6800) );
  XNOR U6879 ( .A(n6799), .B(n6800), .Z(n6801) );
  NAND U6880 ( .A(n6583), .B(n6582), .Z(n6587) );
  NAND U6881 ( .A(n6585), .B(n6584), .Z(n6586) );
  NAND U6882 ( .A(n6587), .B(n6586), .Z(n6738) );
  OR U6883 ( .A(n6589), .B(n6588), .Z(n6593) );
  OR U6884 ( .A(n6591), .B(n6590), .Z(n6592) );
  NAND U6885 ( .A(n6593), .B(n6592), .Z(n6736) );
  NANDN U6886 ( .A(n6595), .B(n6594), .Z(n6599) );
  NANDN U6887 ( .A(n6597), .B(n6596), .Z(n6598) );
  AND U6888 ( .A(n6599), .B(n6598), .Z(n6735) );
  XNOR U6889 ( .A(n6736), .B(n6735), .Z(n6737) );
  XOR U6890 ( .A(n6738), .B(n6737), .Z(n6802) );
  XOR U6891 ( .A(n6801), .B(n6802), .Z(n6813) );
  NANDN U6892 ( .A(n6605), .B(n6604), .Z(n6609) );
  NANDN U6893 ( .A(n6607), .B(n6606), .Z(n6608) );
  NAND U6894 ( .A(n6609), .B(n6608), .Z(n6796) );
  NAND U6895 ( .A(n6611), .B(n6610), .Z(n6615) );
  NAND U6896 ( .A(n6613), .B(n6612), .Z(n6614) );
  NAND U6897 ( .A(n6615), .B(n6614), .Z(n6794) );
  NANDN U6898 ( .A(n6617), .B(n6616), .Z(n6621) );
  NAND U6899 ( .A(n6619), .B(n6618), .Z(n6620) );
  NAND U6900 ( .A(n6621), .B(n6620), .Z(n6739) );
  NANDN U6901 ( .A(n6623), .B(n6622), .Z(n6627) );
  NAND U6902 ( .A(n6625), .B(n6624), .Z(n6626) );
  AND U6903 ( .A(n6627), .B(n6626), .Z(n6740) );
  XNOR U6904 ( .A(n6739), .B(n6740), .Z(n6741) );
  NAND U6905 ( .A(n6628), .B(n8286), .Z(n6630) );
  XNOR U6906 ( .A(n9457), .B(b[9]), .Z(n6757) );
  NAND U6907 ( .A(n6757), .B(n8288), .Z(n6629) );
  NAND U6908 ( .A(n6630), .B(n6629), .Z(n6707) );
  NAND U6909 ( .A(n6631), .B(n8961), .Z(n6633) );
  XOR U6910 ( .A(b[15]), .B(a[45]), .Z(n6751) );
  NAND U6911 ( .A(n6751), .B(n8963), .Z(n6632) );
  NAND U6912 ( .A(n6633), .B(n6632), .Z(n6705) );
  XNOR U6913 ( .A(b[21]), .B(a[39]), .Z(n6754) );
  NANDN U6914 ( .A(n6754), .B(n9493), .Z(n6636) );
  NANDN U6915 ( .A(n6634), .B(n9495), .Z(n6635) );
  AND U6916 ( .A(n6636), .B(n6635), .Z(n6706) );
  XOR U6917 ( .A(n6705), .B(n6706), .Z(n6708) );
  XNOR U6918 ( .A(n6707), .B(n6708), .Z(n6696) );
  XNOR U6919 ( .A(a[49]), .B(b[11]), .Z(n6760) );
  NANDN U6920 ( .A(n6760), .B(n8541), .Z(n6639) );
  NANDN U6921 ( .A(n6637), .B(n8542), .Z(n6638) );
  NAND U6922 ( .A(n6639), .B(n6638), .Z(n6694) );
  XNOR U6923 ( .A(b[13]), .B(a[47]), .Z(n6763) );
  NANDN U6924 ( .A(n6763), .B(n8730), .Z(n6642) );
  NANDN U6925 ( .A(n6640), .B(n8731), .Z(n6641) );
  NAND U6926 ( .A(n6642), .B(n6641), .Z(n6693) );
  XNOR U6927 ( .A(n6696), .B(n6695), .Z(n6690) );
  NAND U6928 ( .A(n6643), .B(n9875), .Z(n6645) );
  XNOR U6929 ( .A(n322), .B(a[31]), .Z(n6778) );
  NANDN U6930 ( .A(n9874), .B(n6778), .Z(n6644) );
  NAND U6931 ( .A(n6645), .B(n6644), .Z(n6711) );
  NANDN U6932 ( .A(n323), .B(a[27]), .Z(n6712) );
  XNOR U6933 ( .A(n6711), .B(n6712), .Z(n6714) );
  NANDN U6934 ( .A(n315), .B(a[59]), .Z(n6646) );
  XNOR U6935 ( .A(b[1]), .B(n6646), .Z(n6648) );
  NANDN U6936 ( .A(b[0]), .B(a[58]), .Z(n6647) );
  AND U6937 ( .A(n6648), .B(n6647), .Z(n6713) );
  XNOR U6938 ( .A(n6714), .B(n6713), .Z(n6688) );
  NANDN U6939 ( .A(n6649), .B(n9622), .Z(n6651) );
  XNOR U6940 ( .A(b[23]), .B(a[37]), .Z(n6769) );
  OR U6941 ( .A(n6769), .B(n9621), .Z(n6650) );
  NAND U6942 ( .A(n6651), .B(n6650), .Z(n6784) );
  XNOR U6943 ( .A(a[53]), .B(b[7]), .Z(n6772) );
  OR U6944 ( .A(n6772), .B(n8013), .Z(n6654) );
  NANDN U6945 ( .A(n6652), .B(n8014), .Z(n6653) );
  NAND U6946 ( .A(n6654), .B(n6653), .Z(n6781) );
  XNOR U6947 ( .A(b[25]), .B(a[35]), .Z(n6766) );
  NANDN U6948 ( .A(n6766), .B(n9706), .Z(n6657) );
  NANDN U6949 ( .A(n6655), .B(n9707), .Z(n6656) );
  AND U6950 ( .A(n6657), .B(n6656), .Z(n6782) );
  XNOR U6951 ( .A(n6781), .B(n6782), .Z(n6783) );
  XOR U6952 ( .A(n6784), .B(n6783), .Z(n6687) );
  XOR U6953 ( .A(n6690), .B(n6689), .Z(n6742) );
  XNOR U6954 ( .A(n6741), .B(n6742), .Z(n6793) );
  XOR U6955 ( .A(n6794), .B(n6793), .Z(n6795) );
  XNOR U6956 ( .A(n6796), .B(n6795), .Z(n6811) );
  XNOR U6957 ( .A(n6812), .B(n6811), .Z(n6814) );
  XNOR U6958 ( .A(n6813), .B(n6814), .Z(n6808) );
  XOR U6959 ( .A(n6807), .B(n6808), .Z(n6684) );
  NANDN U6960 ( .A(n6659), .B(n6658), .Z(n6663) );
  NAND U6961 ( .A(n6661), .B(n6660), .Z(n6662) );
  NAND U6962 ( .A(n6663), .B(n6662), .Z(n6681) );
  NANDN U6963 ( .A(n6665), .B(n6664), .Z(n6669) );
  OR U6964 ( .A(n6667), .B(n6666), .Z(n6668) );
  NAND U6965 ( .A(n6669), .B(n6668), .Z(n6682) );
  XNOR U6966 ( .A(n6681), .B(n6682), .Z(n6683) );
  XNOR U6967 ( .A(n6684), .B(n6683), .Z(n6676) );
  XNOR U6968 ( .A(n6675), .B(n6676), .Z(n6677) );
  XNOR U6969 ( .A(n6678), .B(n6677), .Z(n6817) );
  XNOR U6970 ( .A(n6817), .B(sreg[91]), .Z(n6819) );
  NAND U6971 ( .A(n6670), .B(sreg[90]), .Z(n6674) );
  OR U6972 ( .A(n6672), .B(n6671), .Z(n6673) );
  AND U6973 ( .A(n6674), .B(n6673), .Z(n6818) );
  XOR U6974 ( .A(n6819), .B(n6818), .Z(c[91]) );
  NANDN U6975 ( .A(n6676), .B(n6675), .Z(n6680) );
  NAND U6976 ( .A(n6678), .B(n6677), .Z(n6679) );
  NAND U6977 ( .A(n6680), .B(n6679), .Z(n6825) );
  NANDN U6978 ( .A(n6682), .B(n6681), .Z(n6686) );
  NAND U6979 ( .A(n6684), .B(n6683), .Z(n6685) );
  NAND U6980 ( .A(n6686), .B(n6685), .Z(n6823) );
  NANDN U6981 ( .A(n6688), .B(n6687), .Z(n6692) );
  NANDN U6982 ( .A(n6690), .B(n6689), .Z(n6691) );
  NAND U6983 ( .A(n6692), .B(n6691), .Z(n6944) );
  OR U6984 ( .A(n6694), .B(n6693), .Z(n6698) );
  NANDN U6985 ( .A(n6696), .B(n6695), .Z(n6697) );
  NAND U6986 ( .A(n6698), .B(n6697), .Z(n6882) );
  NANDN U6987 ( .A(n6700), .B(n6699), .Z(n6704) );
  NANDN U6988 ( .A(n6702), .B(n6701), .Z(n6703) );
  NAND U6989 ( .A(n6704), .B(n6703), .Z(n6881) );
  NANDN U6990 ( .A(n6706), .B(n6705), .Z(n6710) );
  NANDN U6991 ( .A(n6708), .B(n6707), .Z(n6709) );
  NAND U6992 ( .A(n6710), .B(n6709), .Z(n6880) );
  XOR U6993 ( .A(n6882), .B(n6883), .Z(n6941) );
  NANDN U6994 ( .A(n6712), .B(n6711), .Z(n6716) );
  NAND U6995 ( .A(n6714), .B(n6713), .Z(n6715) );
  NAND U6996 ( .A(n6716), .B(n6715), .Z(n6895) );
  NANDN U6997 ( .A(n6717), .B(n9801), .Z(n6719) );
  XNOR U6998 ( .A(b[27]), .B(a[34]), .Z(n6865) );
  OR U6999 ( .A(n6865), .B(n9751), .Z(n6718) );
  NAND U7000 ( .A(n6719), .B(n6718), .Z(n6901) );
  NAND U7001 ( .A(n6720), .B(n9379), .Z(n6722) );
  XNOR U7002 ( .A(n9562), .B(a[42]), .Z(n6871) );
  NAND U7003 ( .A(n6871), .B(n9378), .Z(n6721) );
  NAND U7004 ( .A(n6722), .B(n6721), .Z(n6898) );
  XOR U7005 ( .A(a[56]), .B(n317), .Z(n6868) );
  NANDN U7006 ( .A(n6868), .B(n7905), .Z(n6725) );
  NANDN U7007 ( .A(n6723), .B(n7906), .Z(n6724) );
  AND U7008 ( .A(n6725), .B(n6724), .Z(n6899) );
  XNOR U7009 ( .A(n6898), .B(n6899), .Z(n6900) );
  XNOR U7010 ( .A(n6901), .B(n6900), .Z(n6893) );
  XOR U7011 ( .A(b[17]), .B(n8444), .Z(n6862) );
  NANDN U7012 ( .A(n6862), .B(n9107), .Z(n6728) );
  NAND U7013 ( .A(n6726), .B(n9105), .Z(n6727) );
  AND U7014 ( .A(n6728), .B(n6727), .Z(n6847) );
  NAND U7015 ( .A(n6729), .B(n9914), .Z(n6731) );
  XNOR U7016 ( .A(n323), .B(a[30]), .Z(n6856) );
  NANDN U7017 ( .A(n9913), .B(n6856), .Z(n6730) );
  NAND U7018 ( .A(n6731), .B(n6730), .Z(n6844) );
  NAND U7019 ( .A(n6732), .B(n7622), .Z(n6734) );
  XNOR U7020 ( .A(a[58]), .B(n316), .Z(n6859) );
  NAND U7021 ( .A(n6859), .B(n7620), .Z(n6733) );
  NAND U7022 ( .A(n6734), .B(n6733), .Z(n6845) );
  XOR U7023 ( .A(n6844), .B(n6845), .Z(n6846) );
  XNOR U7024 ( .A(n6847), .B(n6846), .Z(n6892) );
  XNOR U7025 ( .A(n6893), .B(n6892), .Z(n6894) );
  XNOR U7026 ( .A(n6895), .B(n6894), .Z(n6942) );
  XNOR U7027 ( .A(n6941), .B(n6942), .Z(n6943) );
  XNOR U7028 ( .A(n6944), .B(n6943), .Z(n6953) );
  NANDN U7029 ( .A(n6740), .B(n6739), .Z(n6744) );
  NANDN U7030 ( .A(n6742), .B(n6741), .Z(n6743) );
  NAND U7031 ( .A(n6744), .B(n6743), .Z(n6948) );
  NAND U7032 ( .A(n6746), .B(n6745), .Z(n6750) );
  NANDN U7033 ( .A(n6748), .B(n6747), .Z(n6749) );
  NAND U7034 ( .A(n6750), .B(n6749), .Z(n6945) );
  NAND U7035 ( .A(n6751), .B(n8961), .Z(n6753) );
  XNOR U7036 ( .A(b[15]), .B(n8654), .Z(n6929) );
  NAND U7037 ( .A(n6929), .B(n8963), .Z(n6752) );
  NAND U7038 ( .A(n6753), .B(n6752), .Z(n6850) );
  XOR U7039 ( .A(b[21]), .B(n7932), .Z(n6932) );
  NANDN U7040 ( .A(n6932), .B(n9493), .Z(n6756) );
  NANDN U7041 ( .A(n6754), .B(n9495), .Z(n6755) );
  AND U7042 ( .A(n6756), .B(n6755), .Z(n6851) );
  XOR U7043 ( .A(n6850), .B(n6851), .Z(n6853) );
  XNOR U7044 ( .A(a[52]), .B(b[9]), .Z(n6926) );
  NANDN U7045 ( .A(n6926), .B(n8288), .Z(n6759) );
  NAND U7046 ( .A(n6757), .B(n8286), .Z(n6758) );
  AND U7047 ( .A(n6759), .B(n6758), .Z(n6852) );
  XNOR U7048 ( .A(n6853), .B(n6852), .Z(n6841) );
  XOR U7049 ( .A(n9033), .B(b[11]), .Z(n6938) );
  NANDN U7050 ( .A(n6938), .B(n8541), .Z(n6762) );
  NANDN U7051 ( .A(n6760), .B(n8542), .Z(n6761) );
  NAND U7052 ( .A(n6762), .B(n6761), .Z(n6839) );
  XOR U7053 ( .A(n8837), .B(b[13]), .Z(n6935) );
  NANDN U7054 ( .A(n6935), .B(n8730), .Z(n6765) );
  NANDN U7055 ( .A(n6763), .B(n8731), .Z(n6764) );
  AND U7056 ( .A(n6765), .B(n6764), .Z(n6838) );
  XNOR U7057 ( .A(n6839), .B(n6838), .Z(n6840) );
  XNOR U7058 ( .A(n6841), .B(n6840), .Z(n6835) );
  XOR U7059 ( .A(b[25]), .B(n7293), .Z(n6923) );
  NANDN U7060 ( .A(n6923), .B(n9706), .Z(n6768) );
  NANDN U7061 ( .A(n6766), .B(n9707), .Z(n6767) );
  NAND U7062 ( .A(n6768), .B(n6767), .Z(n6907) );
  NANDN U7063 ( .A(n6769), .B(n9622), .Z(n6771) );
  XOR U7064 ( .A(b[23]), .B(n7672), .Z(n6917) );
  OR U7065 ( .A(n6917), .B(n9621), .Z(n6770) );
  NAND U7066 ( .A(n6771), .B(n6770), .Z(n6904) );
  XNOR U7067 ( .A(a[54]), .B(b[7]), .Z(n6920) );
  OR U7068 ( .A(n6920), .B(n8013), .Z(n6774) );
  NANDN U7069 ( .A(n6772), .B(n8014), .Z(n6773) );
  AND U7070 ( .A(n6774), .B(n6773), .Z(n6905) );
  XNOR U7071 ( .A(n6904), .B(n6905), .Z(n6906) );
  XNOR U7072 ( .A(n6907), .B(n6906), .Z(n6832) );
  NANDN U7073 ( .A(n315), .B(a[60]), .Z(n6775) );
  XNOR U7074 ( .A(b[1]), .B(n6775), .Z(n6777) );
  NANDN U7075 ( .A(b[0]), .B(a[59]), .Z(n6776) );
  AND U7076 ( .A(n6777), .B(n6776), .Z(n6876) );
  NAND U7077 ( .A(n9875), .B(n6778), .Z(n6780) );
  XNOR U7078 ( .A(n322), .B(a[32]), .Z(n6913) );
  NANDN U7079 ( .A(n9874), .B(n6913), .Z(n6779) );
  NAND U7080 ( .A(n6780), .B(n6779), .Z(n6874) );
  NANDN U7081 ( .A(n323), .B(a[28]), .Z(n6875) );
  XNOR U7082 ( .A(n6874), .B(n6875), .Z(n6877) );
  XOR U7083 ( .A(n6876), .B(n6877), .Z(n6833) );
  XNOR U7084 ( .A(n6832), .B(n6833), .Z(n6834) );
  XOR U7085 ( .A(n6835), .B(n6834), .Z(n6889) );
  NANDN U7086 ( .A(n6782), .B(n6781), .Z(n6786) );
  NAND U7087 ( .A(n6784), .B(n6783), .Z(n6785) );
  NAND U7088 ( .A(n6786), .B(n6785), .Z(n6886) );
  NANDN U7089 ( .A(n6788), .B(n6787), .Z(n6792) );
  NAND U7090 ( .A(n6790), .B(n6789), .Z(n6791) );
  AND U7091 ( .A(n6792), .B(n6791), .Z(n6887) );
  XNOR U7092 ( .A(n6886), .B(n6887), .Z(n6888) );
  XNOR U7093 ( .A(n6889), .B(n6888), .Z(n6946) );
  XNOR U7094 ( .A(n6945), .B(n6946), .Z(n6947) );
  XOR U7095 ( .A(n6948), .B(n6947), .Z(n6952) );
  XOR U7096 ( .A(n6951), .B(n6952), .Z(n6954) );
  XNOR U7097 ( .A(n6953), .B(n6954), .Z(n6960) );
  NAND U7098 ( .A(n6794), .B(n6793), .Z(n6798) );
  NAND U7099 ( .A(n6796), .B(n6795), .Z(n6797) );
  NAND U7100 ( .A(n6798), .B(n6797), .Z(n6957) );
  NANDN U7101 ( .A(n6800), .B(n6799), .Z(n6804) );
  NAND U7102 ( .A(n6802), .B(n6801), .Z(n6803) );
  NAND U7103 ( .A(n6804), .B(n6803), .Z(n6958) );
  XNOR U7104 ( .A(n6957), .B(n6958), .Z(n6959) );
  XNOR U7105 ( .A(n6960), .B(n6959), .Z(n6829) );
  NANDN U7106 ( .A(n6806), .B(n6805), .Z(n6810) );
  NANDN U7107 ( .A(n6808), .B(n6807), .Z(n6809) );
  NAND U7108 ( .A(n6810), .B(n6809), .Z(n6827) );
  OR U7109 ( .A(n6812), .B(n6811), .Z(n6816) );
  OR U7110 ( .A(n6814), .B(n6813), .Z(n6815) );
  AND U7111 ( .A(n6816), .B(n6815), .Z(n6826) );
  XNOR U7112 ( .A(n6827), .B(n6826), .Z(n6828) );
  XNOR U7113 ( .A(n6829), .B(n6828), .Z(n6822) );
  XOR U7114 ( .A(n6823), .B(n6822), .Z(n6824) );
  XNOR U7115 ( .A(n6825), .B(n6824), .Z(n6963) );
  XNOR U7116 ( .A(n6963), .B(sreg[92]), .Z(n6965) );
  NAND U7117 ( .A(n6817), .B(sreg[91]), .Z(n6821) );
  OR U7118 ( .A(n6819), .B(n6818), .Z(n6820) );
  AND U7119 ( .A(n6821), .B(n6820), .Z(n6964) );
  XOR U7120 ( .A(n6965), .B(n6964), .Z(c[92]) );
  NANDN U7121 ( .A(n6827), .B(n6826), .Z(n6831) );
  NANDN U7122 ( .A(n6829), .B(n6828), .Z(n6830) );
  NAND U7123 ( .A(n6831), .B(n6830), .Z(n6969) );
  NANDN U7124 ( .A(n6833), .B(n6832), .Z(n6837) );
  NANDN U7125 ( .A(n6835), .B(n6834), .Z(n6836) );
  NAND U7126 ( .A(n6837), .B(n6836), .Z(n6987) );
  NANDN U7127 ( .A(n6839), .B(n6838), .Z(n6843) );
  NAND U7128 ( .A(n6841), .B(n6840), .Z(n6842) );
  NAND U7129 ( .A(n6843), .B(n6842), .Z(n7039) );
  NAND U7130 ( .A(n6845), .B(n6844), .Z(n6849) );
  NANDN U7131 ( .A(n6847), .B(n6846), .Z(n6848) );
  NAND U7132 ( .A(n6849), .B(n6848), .Z(n7037) );
  NANDN U7133 ( .A(n6851), .B(n6850), .Z(n6855) );
  OR U7134 ( .A(n6853), .B(n6852), .Z(n6854) );
  AND U7135 ( .A(n6855), .B(n6854), .Z(n7036) );
  XNOR U7136 ( .A(n7037), .B(n7036), .Z(n7038) );
  XNOR U7137 ( .A(n7039), .B(n7038), .Z(n6985) );
  NAND U7138 ( .A(n6856), .B(n9914), .Z(n6858) );
  XNOR U7139 ( .A(n323), .B(a[31]), .Z(n7006) );
  NANDN U7140 ( .A(n9913), .B(n7006), .Z(n6857) );
  NAND U7141 ( .A(n6858), .B(n6857), .Z(n6994) );
  NAND U7142 ( .A(n6859), .B(n7622), .Z(n6861) );
  XNOR U7143 ( .A(a[59]), .B(n316), .Z(n7009) );
  NAND U7144 ( .A(n7009), .B(n7620), .Z(n6860) );
  NAND U7145 ( .A(n6861), .B(n6860), .Z(n6995) );
  XOR U7146 ( .A(n6994), .B(n6995), .Z(n6996) );
  XNOR U7147 ( .A(b[17]), .B(a[45]), .Z(n7012) );
  NANDN U7148 ( .A(n7012), .B(n9107), .Z(n6864) );
  NANDN U7149 ( .A(n6862), .B(n9105), .Z(n6863) );
  AND U7150 ( .A(n6864), .B(n6863), .Z(n6997) );
  XOR U7151 ( .A(n6996), .B(n6997), .Z(n7042) );
  NANDN U7152 ( .A(n6865), .B(n9801), .Z(n6867) );
  XNOR U7153 ( .A(b[27]), .B(a[35]), .Z(n7015) );
  OR U7154 ( .A(n7015), .B(n9751), .Z(n6866) );
  NAND U7155 ( .A(n6867), .B(n6866), .Z(n7093) );
  XNOR U7156 ( .A(a[57]), .B(b[5]), .Z(n7021) );
  NANDN U7157 ( .A(n7021), .B(n7905), .Z(n6870) );
  NANDN U7158 ( .A(n6868), .B(n7906), .Z(n6869) );
  NAND U7159 ( .A(n6870), .B(n6869), .Z(n7090) );
  NAND U7160 ( .A(n6871), .B(n9379), .Z(n6873) );
  XNOR U7161 ( .A(b[19]), .B(a[43]), .Z(n7018) );
  NANDN U7162 ( .A(n7018), .B(n9378), .Z(n6872) );
  AND U7163 ( .A(n6873), .B(n6872), .Z(n7091) );
  XNOR U7164 ( .A(n7090), .B(n7091), .Z(n7092) );
  XOR U7165 ( .A(n7093), .B(n7092), .Z(n7043) );
  XNOR U7166 ( .A(n7042), .B(n7043), .Z(n7044) );
  NANDN U7167 ( .A(n6875), .B(n6874), .Z(n6879) );
  NAND U7168 ( .A(n6877), .B(n6876), .Z(n6878) );
  AND U7169 ( .A(n6879), .B(n6878), .Z(n7045) );
  XOR U7170 ( .A(n7044), .B(n7045), .Z(n6984) );
  XNOR U7171 ( .A(n6985), .B(n6984), .Z(n6986) );
  XNOR U7172 ( .A(n6987), .B(n6986), .Z(n7104) );
  OR U7173 ( .A(n6881), .B(n6880), .Z(n6885) );
  NANDN U7174 ( .A(n6883), .B(n6882), .Z(n6884) );
  NAND U7175 ( .A(n6885), .B(n6884), .Z(n7103) );
  NANDN U7176 ( .A(n6887), .B(n6886), .Z(n6891) );
  NAND U7177 ( .A(n6889), .B(n6888), .Z(n6890) );
  NAND U7178 ( .A(n6891), .B(n6890), .Z(n6981) );
  NANDN U7179 ( .A(n6893), .B(n6892), .Z(n6897) );
  NAND U7180 ( .A(n6895), .B(n6894), .Z(n6896) );
  NAND U7181 ( .A(n6897), .B(n6896), .Z(n6978) );
  NANDN U7182 ( .A(n6899), .B(n6898), .Z(n6903) );
  NAND U7183 ( .A(n6901), .B(n6900), .Z(n6902) );
  NAND U7184 ( .A(n6903), .B(n6902), .Z(n7049) );
  NANDN U7185 ( .A(n6905), .B(n6904), .Z(n6909) );
  NAND U7186 ( .A(n6907), .B(n6906), .Z(n6908) );
  AND U7187 ( .A(n6909), .B(n6908), .Z(n7048) );
  XNOR U7188 ( .A(n7049), .B(n7048), .Z(n7050) );
  NANDN U7189 ( .A(n315), .B(a[61]), .Z(n6910) );
  XNOR U7190 ( .A(b[1]), .B(n6910), .Z(n6912) );
  IV U7191 ( .A(a[60]), .Z(n9805) );
  NANDN U7192 ( .A(n9805), .B(n315), .Z(n6911) );
  AND U7193 ( .A(n6912), .B(n6911), .Z(n7026) );
  NAND U7194 ( .A(n9875), .B(n6913), .Z(n6916) );
  XOR U7195 ( .A(b[29]), .B(n6914), .Z(n7081) );
  OR U7196 ( .A(n7081), .B(n9874), .Z(n6915) );
  NAND U7197 ( .A(n6916), .B(n6915), .Z(n7024) );
  NANDN U7198 ( .A(n323), .B(a[29]), .Z(n7025) );
  XNOR U7199 ( .A(n7024), .B(n7025), .Z(n7027) );
  XOR U7200 ( .A(n7026), .B(n7027), .Z(n7032) );
  NANDN U7201 ( .A(n6917), .B(n9622), .Z(n6919) );
  XNOR U7202 ( .A(b[23]), .B(a[39]), .Z(n7072) );
  OR U7203 ( .A(n7072), .B(n9621), .Z(n6918) );
  NAND U7204 ( .A(n6919), .B(n6918), .Z(n7087) );
  XOR U7205 ( .A(a[55]), .B(b[7]), .Z(n7075) );
  NANDN U7206 ( .A(n8013), .B(n7075), .Z(n6922) );
  NANDN U7207 ( .A(n6920), .B(n8014), .Z(n6921) );
  NAND U7208 ( .A(n6922), .B(n6921), .Z(n7084) );
  XNOR U7209 ( .A(b[25]), .B(a[37]), .Z(n7069) );
  NANDN U7210 ( .A(n7069), .B(n9706), .Z(n6925) );
  NANDN U7211 ( .A(n6923), .B(n9707), .Z(n6924) );
  AND U7212 ( .A(n6925), .B(n6924), .Z(n7085) );
  XNOR U7213 ( .A(n7084), .B(n7085), .Z(n7086) );
  XOR U7214 ( .A(n7087), .B(n7086), .Z(n7030) );
  NANDN U7215 ( .A(n6926), .B(n8286), .Z(n6928) );
  XNOR U7216 ( .A(n9564), .B(b[9]), .Z(n7063) );
  NAND U7217 ( .A(n7063), .B(n8288), .Z(n6927) );
  NAND U7218 ( .A(n6928), .B(n6927), .Z(n7002) );
  NAND U7219 ( .A(n6929), .B(n8961), .Z(n6931) );
  XOR U7220 ( .A(b[15]), .B(a[47]), .Z(n7060) );
  NAND U7221 ( .A(n7060), .B(n8963), .Z(n6930) );
  NAND U7222 ( .A(n6931), .B(n6930), .Z(n7000) );
  XNOR U7223 ( .A(b[21]), .B(a[41]), .Z(n7066) );
  NANDN U7224 ( .A(n7066), .B(n9493), .Z(n6934) );
  NANDN U7225 ( .A(n6932), .B(n9495), .Z(n6933) );
  AND U7226 ( .A(n6934), .B(n6933), .Z(n7001) );
  XOR U7227 ( .A(n7000), .B(n7001), .Z(n7003) );
  XNOR U7228 ( .A(n7002), .B(n7003), .Z(n6991) );
  XOR U7229 ( .A(a[49]), .B(b[13]), .Z(n7057) );
  NAND U7230 ( .A(n8730), .B(n7057), .Z(n6937) );
  NANDN U7231 ( .A(n6935), .B(n8731), .Z(n6936) );
  NAND U7232 ( .A(n6937), .B(n6936), .Z(n6989) );
  XNOR U7233 ( .A(a[51]), .B(b[11]), .Z(n7054) );
  NANDN U7234 ( .A(n7054), .B(n8541), .Z(n6940) );
  NANDN U7235 ( .A(n6938), .B(n8542), .Z(n6939) );
  AND U7236 ( .A(n6940), .B(n6939), .Z(n6988) );
  XNOR U7237 ( .A(n6989), .B(n6988), .Z(n6990) );
  XOR U7238 ( .A(n6991), .B(n6990), .Z(n7031) );
  XNOR U7239 ( .A(n7030), .B(n7031), .Z(n7033) );
  XNOR U7240 ( .A(n7032), .B(n7033), .Z(n7051) );
  XNOR U7241 ( .A(n7050), .B(n7051), .Z(n6979) );
  XNOR U7242 ( .A(n6978), .B(n6979), .Z(n6980) );
  XOR U7243 ( .A(n6981), .B(n6980), .Z(n7102) );
  XOR U7244 ( .A(n7103), .B(n7102), .Z(n7105) );
  XNOR U7245 ( .A(n7104), .B(n7105), .Z(n7099) );
  NANDN U7246 ( .A(n6946), .B(n6945), .Z(n6950) );
  NAND U7247 ( .A(n6948), .B(n6947), .Z(n6949) );
  AND U7248 ( .A(n6950), .B(n6949), .Z(n7096) );
  XNOR U7249 ( .A(n7097), .B(n7096), .Z(n7098) );
  XNOR U7250 ( .A(n7099), .B(n7098), .Z(n6976) );
  NANDN U7251 ( .A(n6952), .B(n6951), .Z(n6956) );
  NANDN U7252 ( .A(n6954), .B(n6953), .Z(n6955) );
  NAND U7253 ( .A(n6956), .B(n6955), .Z(n6974) );
  NANDN U7254 ( .A(n6958), .B(n6957), .Z(n6962) );
  NANDN U7255 ( .A(n6960), .B(n6959), .Z(n6961) );
  NAND U7256 ( .A(n6962), .B(n6961), .Z(n6975) );
  XNOR U7257 ( .A(n6974), .B(n6975), .Z(n6977) );
  XOR U7258 ( .A(n6976), .B(n6977), .Z(n6968) );
  XOR U7259 ( .A(n6969), .B(n6968), .Z(n6970) );
  XNOR U7260 ( .A(n6971), .B(n6970), .Z(n7108) );
  XNOR U7261 ( .A(n7108), .B(sreg[93]), .Z(n7110) );
  NAND U7262 ( .A(n6963), .B(sreg[92]), .Z(n6967) );
  OR U7263 ( .A(n6965), .B(n6964), .Z(n6966) );
  AND U7264 ( .A(n6967), .B(n6966), .Z(n7109) );
  XOR U7265 ( .A(n7110), .B(n7109), .Z(c[93]) );
  NAND U7266 ( .A(n6969), .B(n6968), .Z(n6973) );
  NAND U7267 ( .A(n6971), .B(n6970), .Z(n6972) );
  NAND U7268 ( .A(n6973), .B(n6972), .Z(n7116) );
  NANDN U7269 ( .A(n6979), .B(n6978), .Z(n6983) );
  NAND U7270 ( .A(n6981), .B(n6980), .Z(n6982) );
  NAND U7271 ( .A(n6983), .B(n6982), .Z(n7131) );
  XNOR U7272 ( .A(n7131), .B(n7132), .Z(n7133) );
  NANDN U7273 ( .A(n6989), .B(n6988), .Z(n6993) );
  NANDN U7274 ( .A(n6991), .B(n6990), .Z(n6992) );
  NAND U7275 ( .A(n6993), .B(n6992), .Z(n7194) );
  NAND U7276 ( .A(n6995), .B(n6994), .Z(n6999) );
  NANDN U7277 ( .A(n6997), .B(n6996), .Z(n6998) );
  NAND U7278 ( .A(n6999), .B(n6998), .Z(n7192) );
  NANDN U7279 ( .A(n7001), .B(n7000), .Z(n7005) );
  NANDN U7280 ( .A(n7003), .B(n7002), .Z(n7004) );
  AND U7281 ( .A(n7005), .B(n7004), .Z(n7191) );
  XNOR U7282 ( .A(n7192), .B(n7191), .Z(n7193) );
  XNOR U7283 ( .A(n7194), .B(n7193), .Z(n7251) );
  NAND U7284 ( .A(n7006), .B(n9914), .Z(n7008) );
  XNOR U7285 ( .A(n323), .B(a[32]), .Z(n7215) );
  NANDN U7286 ( .A(n9913), .B(n7215), .Z(n7007) );
  NAND U7287 ( .A(n7008), .B(n7007), .Z(n7233) );
  NAND U7288 ( .A(n7009), .B(n7622), .Z(n7011) );
  XNOR U7289 ( .A(n9805), .B(b[3]), .Z(n7218) );
  NAND U7290 ( .A(n7218), .B(n7620), .Z(n7010) );
  NAND U7291 ( .A(n7011), .B(n7010), .Z(n7234) );
  XOR U7292 ( .A(n7233), .B(n7234), .Z(n7235) );
  XOR U7293 ( .A(b[17]), .B(n8654), .Z(n7212) );
  NANDN U7294 ( .A(n7212), .B(n9107), .Z(n7014) );
  NANDN U7295 ( .A(n7012), .B(n9105), .Z(n7013) );
  AND U7296 ( .A(n7014), .B(n7013), .Z(n7236) );
  XOR U7297 ( .A(n7235), .B(n7236), .Z(n7143) );
  NANDN U7298 ( .A(n7015), .B(n9801), .Z(n7017) );
  XOR U7299 ( .A(b[27]), .B(n7293), .Z(n7203) );
  OR U7300 ( .A(n7203), .B(n9751), .Z(n7016) );
  NAND U7301 ( .A(n7017), .B(n7016), .Z(n7188) );
  NANDN U7302 ( .A(n7018), .B(n9379), .Z(n7020) );
  XNOR U7303 ( .A(n9562), .B(a[44]), .Z(n7209) );
  NAND U7304 ( .A(n7209), .B(n9378), .Z(n7019) );
  NAND U7305 ( .A(n7020), .B(n7019), .Z(n7185) );
  XNOR U7306 ( .A(a[58]), .B(b[5]), .Z(n7206) );
  NANDN U7307 ( .A(n7206), .B(n7905), .Z(n7023) );
  NANDN U7308 ( .A(n7021), .B(n7906), .Z(n7022) );
  AND U7309 ( .A(n7023), .B(n7022), .Z(n7186) );
  XNOR U7310 ( .A(n7185), .B(n7186), .Z(n7187) );
  XOR U7311 ( .A(n7188), .B(n7187), .Z(n7144) );
  XNOR U7312 ( .A(n7143), .B(n7144), .Z(n7145) );
  NANDN U7313 ( .A(n7025), .B(n7024), .Z(n7029) );
  NAND U7314 ( .A(n7027), .B(n7026), .Z(n7028) );
  NAND U7315 ( .A(n7029), .B(n7028), .Z(n7146) );
  XNOR U7316 ( .A(n7145), .B(n7146), .Z(n7252) );
  XNOR U7317 ( .A(n7251), .B(n7252), .Z(n7253) );
  OR U7318 ( .A(n7031), .B(n7030), .Z(n7035) );
  OR U7319 ( .A(n7033), .B(n7032), .Z(n7034) );
  AND U7320 ( .A(n7035), .B(n7034), .Z(n7254) );
  XNOR U7321 ( .A(n7253), .B(n7254), .Z(n7127) );
  NANDN U7322 ( .A(n7037), .B(n7036), .Z(n7041) );
  NAND U7323 ( .A(n7039), .B(n7038), .Z(n7040) );
  NAND U7324 ( .A(n7041), .B(n7040), .Z(n7126) );
  NANDN U7325 ( .A(n7043), .B(n7042), .Z(n7047) );
  NAND U7326 ( .A(n7045), .B(n7044), .Z(n7046) );
  NAND U7327 ( .A(n7047), .B(n7046), .Z(n7246) );
  NANDN U7328 ( .A(n7049), .B(n7048), .Z(n7053) );
  NANDN U7329 ( .A(n7051), .B(n7050), .Z(n7052) );
  AND U7330 ( .A(n7053), .B(n7052), .Z(n7245) );
  XNOR U7331 ( .A(n7246), .B(n7245), .Z(n7247) );
  XNOR U7332 ( .A(n9217), .B(b[11]), .Z(n7176) );
  NAND U7333 ( .A(n7176), .B(n8541), .Z(n7056) );
  NANDN U7334 ( .A(n7054), .B(n8542), .Z(n7055) );
  NAND U7335 ( .A(n7056), .B(n7055), .Z(n7242) );
  XNOR U7336 ( .A(n9033), .B(b[13]), .Z(n7173) );
  NAND U7337 ( .A(n7173), .B(n8730), .Z(n7059) );
  NAND U7338 ( .A(n7057), .B(n8731), .Z(n7058) );
  NAND U7339 ( .A(n7059), .B(n7058), .Z(n7240) );
  NAND U7340 ( .A(n7060), .B(n8961), .Z(n7062) );
  XNOR U7341 ( .A(b[15]), .B(n8837), .Z(n7164) );
  NAND U7342 ( .A(n7164), .B(n8963), .Z(n7061) );
  NAND U7343 ( .A(n7062), .B(n7061), .Z(n7229) );
  NAND U7344 ( .A(n7063), .B(n8286), .Z(n7065) );
  XNOR U7345 ( .A(n9353), .B(b[9]), .Z(n7167) );
  NAND U7346 ( .A(n7167), .B(n8288), .Z(n7064) );
  NAND U7347 ( .A(n7065), .B(n7064), .Z(n7227) );
  XOR U7348 ( .A(b[21]), .B(n8156), .Z(n7170) );
  NANDN U7349 ( .A(n7170), .B(n9493), .Z(n7068) );
  NANDN U7350 ( .A(n7066), .B(n9495), .Z(n7067) );
  AND U7351 ( .A(n7068), .B(n7067), .Z(n7228) );
  XOR U7352 ( .A(n7227), .B(n7228), .Z(n7230) );
  XNOR U7353 ( .A(n7229), .B(n7230), .Z(n7239) );
  XOR U7354 ( .A(n7240), .B(n7239), .Z(n7241) );
  XNOR U7355 ( .A(n7242), .B(n7241), .Z(n7199) );
  XOR U7356 ( .A(b[25]), .B(n7672), .Z(n7149) );
  NANDN U7357 ( .A(n7149), .B(n9706), .Z(n7071) );
  NANDN U7358 ( .A(n7069), .B(n9707), .Z(n7070) );
  NAND U7359 ( .A(n7071), .B(n7070), .Z(n7182) );
  NANDN U7360 ( .A(n7072), .B(n9622), .Z(n7074) );
  XOR U7361 ( .A(b[23]), .B(n7932), .Z(n7152) );
  OR U7362 ( .A(n7152), .B(n9621), .Z(n7073) );
  NAND U7363 ( .A(n7074), .B(n7073), .Z(n7179) );
  XNOR U7364 ( .A(a[56]), .B(b[7]), .Z(n7155) );
  OR U7365 ( .A(n7155), .B(n8013), .Z(n7077) );
  NAND U7366 ( .A(n7075), .B(n8014), .Z(n7076) );
  AND U7367 ( .A(n7077), .B(n7076), .Z(n7180) );
  XNOR U7368 ( .A(n7179), .B(n7180), .Z(n7181) );
  XNOR U7369 ( .A(n7182), .B(n7181), .Z(n7197) );
  NAND U7370 ( .A(a[30]), .B(b[31]), .Z(n7224) );
  NANDN U7371 ( .A(n315), .B(a[62]), .Z(n7078) );
  XNOR U7372 ( .A(b[1]), .B(n7078), .Z(n7080) );
  NANDN U7373 ( .A(b[0]), .B(a[61]), .Z(n7079) );
  AND U7374 ( .A(n7080), .B(n7079), .Z(n7222) );
  NANDN U7375 ( .A(n7081), .B(n9875), .Z(n7083) );
  XNOR U7376 ( .A(n322), .B(a[34]), .Z(n7161) );
  NANDN U7377 ( .A(n9874), .B(n7161), .Z(n7082) );
  AND U7378 ( .A(n7083), .B(n7082), .Z(n7221) );
  XNOR U7379 ( .A(n7222), .B(n7221), .Z(n7223) );
  XNOR U7380 ( .A(n7224), .B(n7223), .Z(n7198) );
  XOR U7381 ( .A(n7197), .B(n7198), .Z(n7200) );
  XNOR U7382 ( .A(n7199), .B(n7200), .Z(n7140) );
  NANDN U7383 ( .A(n7085), .B(n7084), .Z(n7089) );
  NAND U7384 ( .A(n7087), .B(n7086), .Z(n7088) );
  NAND U7385 ( .A(n7089), .B(n7088), .Z(n7137) );
  NANDN U7386 ( .A(n7091), .B(n7090), .Z(n7095) );
  NAND U7387 ( .A(n7093), .B(n7092), .Z(n7094) );
  AND U7388 ( .A(n7095), .B(n7094), .Z(n7138) );
  XNOR U7389 ( .A(n7137), .B(n7138), .Z(n7139) );
  XOR U7390 ( .A(n7140), .B(n7139), .Z(n7248) );
  XNOR U7391 ( .A(n7247), .B(n7248), .Z(n7125) );
  XOR U7392 ( .A(n7126), .B(n7125), .Z(n7128) );
  XOR U7393 ( .A(n7127), .B(n7128), .Z(n7134) );
  XNOR U7394 ( .A(n7133), .B(n7134), .Z(n7122) );
  NANDN U7395 ( .A(n7097), .B(n7096), .Z(n7101) );
  NANDN U7396 ( .A(n7099), .B(n7098), .Z(n7100) );
  NAND U7397 ( .A(n7101), .B(n7100), .Z(n7119) );
  NANDN U7398 ( .A(n7103), .B(n7102), .Z(n7107) );
  NANDN U7399 ( .A(n7105), .B(n7104), .Z(n7106) );
  NAND U7400 ( .A(n7107), .B(n7106), .Z(n7120) );
  XNOR U7401 ( .A(n7119), .B(n7120), .Z(n7121) );
  XNOR U7402 ( .A(n7122), .B(n7121), .Z(n7114) );
  XNOR U7403 ( .A(n7113), .B(n7114), .Z(n7115) );
  XNOR U7404 ( .A(n7116), .B(n7115), .Z(n7257) );
  XNOR U7405 ( .A(n7257), .B(sreg[94]), .Z(n7259) );
  NAND U7406 ( .A(n7108), .B(sreg[93]), .Z(n7112) );
  OR U7407 ( .A(n7110), .B(n7109), .Z(n7111) );
  AND U7408 ( .A(n7112), .B(n7111), .Z(n7258) );
  XOR U7409 ( .A(n7259), .B(n7258), .Z(c[94]) );
  NANDN U7410 ( .A(n7114), .B(n7113), .Z(n7118) );
  NAND U7411 ( .A(n7116), .B(n7115), .Z(n7117) );
  NAND U7412 ( .A(n7118), .B(n7117), .Z(n7265) );
  NANDN U7413 ( .A(n7120), .B(n7119), .Z(n7124) );
  NAND U7414 ( .A(n7122), .B(n7121), .Z(n7123) );
  NAND U7415 ( .A(n7124), .B(n7123), .Z(n7262) );
  NANDN U7416 ( .A(n7126), .B(n7125), .Z(n7130) );
  OR U7417 ( .A(n7128), .B(n7127), .Z(n7129) );
  NAND U7418 ( .A(n7130), .B(n7129), .Z(n7398) );
  NANDN U7419 ( .A(n7132), .B(n7131), .Z(n7136) );
  NAND U7420 ( .A(n7134), .B(n7133), .Z(n7135) );
  AND U7421 ( .A(n7136), .B(n7135), .Z(n7399) );
  XNOR U7422 ( .A(n7398), .B(n7399), .Z(n7400) );
  NANDN U7423 ( .A(n7138), .B(n7137), .Z(n7142) );
  NANDN U7424 ( .A(n7140), .B(n7139), .Z(n7141) );
  NAND U7425 ( .A(n7142), .B(n7141), .Z(n7383) );
  NANDN U7426 ( .A(n7144), .B(n7143), .Z(n7148) );
  NANDN U7427 ( .A(n7146), .B(n7145), .Z(n7147) );
  NAND U7428 ( .A(n7148), .B(n7147), .Z(n7380) );
  XNOR U7429 ( .A(b[25]), .B(a[39]), .Z(n7302) );
  NANDN U7430 ( .A(n7302), .B(n9706), .Z(n7151) );
  NANDN U7431 ( .A(n7149), .B(n9707), .Z(n7150) );
  NAND U7432 ( .A(n7151), .B(n7150), .Z(n7289) );
  NANDN U7433 ( .A(n7152), .B(n9622), .Z(n7154) );
  XNOR U7434 ( .A(b[23]), .B(a[41]), .Z(n7296) );
  OR U7435 ( .A(n7296), .B(n9621), .Z(n7153) );
  NAND U7436 ( .A(n7154), .B(n7153), .Z(n7286) );
  XOR U7437 ( .A(a[57]), .B(b[7]), .Z(n7299) );
  NANDN U7438 ( .A(n8013), .B(n7299), .Z(n7157) );
  NANDN U7439 ( .A(n7155), .B(n8014), .Z(n7156) );
  AND U7440 ( .A(n7157), .B(n7156), .Z(n7287) );
  XNOR U7441 ( .A(n7286), .B(n7287), .Z(n7288) );
  XOR U7442 ( .A(n7289), .B(n7288), .Z(n7332) );
  IV U7443 ( .A(a[63]), .Z(n9946) );
  NANDN U7444 ( .A(n9946), .B(b[0]), .Z(n7158) );
  XNOR U7445 ( .A(b[1]), .B(n7158), .Z(n7160) );
  IV U7446 ( .A(a[62]), .Z(n9810) );
  NANDN U7447 ( .A(n9810), .B(n315), .Z(n7159) );
  AND U7448 ( .A(n7160), .B(n7159), .Z(n7358) );
  NAND U7449 ( .A(n7161), .B(n9875), .Z(n7163) );
  XNOR U7450 ( .A(n322), .B(a[35]), .Z(n7292) );
  NANDN U7451 ( .A(n9874), .B(n7292), .Z(n7162) );
  NAND U7452 ( .A(n7163), .B(n7162), .Z(n7356) );
  NANDN U7453 ( .A(n323), .B(a[31]), .Z(n7357) );
  XNOR U7454 ( .A(n7356), .B(n7357), .Z(n7359) );
  XOR U7455 ( .A(n7358), .B(n7359), .Z(n7333) );
  XNOR U7456 ( .A(n7332), .B(n7333), .Z(n7335) );
  NAND U7457 ( .A(n7164), .B(n8961), .Z(n7166) );
  XOR U7458 ( .A(b[15]), .B(a[49]), .Z(n7305) );
  NAND U7459 ( .A(n7305), .B(n8963), .Z(n7165) );
  NAND U7460 ( .A(n7166), .B(n7165), .Z(n7376) );
  NAND U7461 ( .A(n7167), .B(n8286), .Z(n7169) );
  XOR U7462 ( .A(a[55]), .B(b[9]), .Z(n7308) );
  NAND U7463 ( .A(n7308), .B(n8288), .Z(n7168) );
  NAND U7464 ( .A(n7169), .B(n7168), .Z(n7374) );
  XNOR U7465 ( .A(b[21]), .B(a[43]), .Z(n7311) );
  NANDN U7466 ( .A(n7311), .B(n9493), .Z(n7172) );
  NANDN U7467 ( .A(n7170), .B(n9495), .Z(n7171) );
  AND U7468 ( .A(n7172), .B(n7171), .Z(n7375) );
  XOR U7469 ( .A(n7374), .B(n7375), .Z(n7377) );
  XNOR U7470 ( .A(n7376), .B(n7377), .Z(n7365) );
  XOR U7471 ( .A(n9457), .B(b[13]), .Z(n7314) );
  NANDN U7472 ( .A(n7314), .B(n8730), .Z(n7175) );
  NAND U7473 ( .A(n8731), .B(n7173), .Z(n7174) );
  NAND U7474 ( .A(n7175), .B(n7174), .Z(n7363) );
  XOR U7475 ( .A(n9564), .B(b[11]), .Z(n7317) );
  NANDN U7476 ( .A(n7317), .B(n8541), .Z(n7178) );
  NAND U7477 ( .A(n8542), .B(n7176), .Z(n7177) );
  AND U7478 ( .A(n7178), .B(n7177), .Z(n7362) );
  XNOR U7479 ( .A(n7363), .B(n7362), .Z(n7364) );
  XNOR U7480 ( .A(n7365), .B(n7364), .Z(n7334) );
  XNOR U7481 ( .A(n7335), .B(n7334), .Z(n7277) );
  NANDN U7482 ( .A(n7180), .B(n7179), .Z(n7184) );
  NAND U7483 ( .A(n7182), .B(n7181), .Z(n7183) );
  NAND U7484 ( .A(n7184), .B(n7183), .Z(n7274) );
  NANDN U7485 ( .A(n7186), .B(n7185), .Z(n7190) );
  NAND U7486 ( .A(n7188), .B(n7187), .Z(n7189) );
  AND U7487 ( .A(n7190), .B(n7189), .Z(n7275) );
  XNOR U7488 ( .A(n7274), .B(n7275), .Z(n7276) );
  XOR U7489 ( .A(n7277), .B(n7276), .Z(n7381) );
  XOR U7490 ( .A(n7380), .B(n7381), .Z(n7382) );
  XNOR U7491 ( .A(n7383), .B(n7382), .Z(n7395) );
  NANDN U7492 ( .A(n7192), .B(n7191), .Z(n7196) );
  NAND U7493 ( .A(n7194), .B(n7193), .Z(n7195) );
  NAND U7494 ( .A(n7196), .B(n7195), .Z(n7392) );
  NANDN U7495 ( .A(n7198), .B(n7197), .Z(n7202) );
  NANDN U7496 ( .A(n7200), .B(n7199), .Z(n7201) );
  NAND U7497 ( .A(n7202), .B(n7201), .Z(n7389) );
  NANDN U7498 ( .A(n7203), .B(n9801), .Z(n7205) );
  XNOR U7499 ( .A(b[27]), .B(a[37]), .Z(n7350) );
  OR U7500 ( .A(n7350), .B(n9751), .Z(n7204) );
  NAND U7501 ( .A(n7205), .B(n7204), .Z(n7283) );
  XNOR U7502 ( .A(a[59]), .B(b[5]), .Z(n7353) );
  NANDN U7503 ( .A(n7353), .B(n7905), .Z(n7208) );
  NANDN U7504 ( .A(n7206), .B(n7906), .Z(n7207) );
  NAND U7505 ( .A(n7208), .B(n7207), .Z(n7280) );
  NAND U7506 ( .A(n7209), .B(n9379), .Z(n7211) );
  XNOR U7507 ( .A(b[19]), .B(a[45]), .Z(n7347) );
  NANDN U7508 ( .A(n7347), .B(n9378), .Z(n7210) );
  AND U7509 ( .A(n7211), .B(n7210), .Z(n7281) );
  XNOR U7510 ( .A(n7280), .B(n7281), .Z(n7282) );
  XNOR U7511 ( .A(n7283), .B(n7282), .Z(n7321) );
  XNOR U7512 ( .A(b[17]), .B(a[47]), .Z(n7338) );
  NANDN U7513 ( .A(n7338), .B(n9107), .Z(n7214) );
  NANDN U7514 ( .A(n7212), .B(n9105), .Z(n7213) );
  AND U7515 ( .A(n7214), .B(n7213), .Z(n7371) );
  NAND U7516 ( .A(n7215), .B(n9914), .Z(n7217) );
  XNOR U7517 ( .A(n323), .B(a[33]), .Z(n7341) );
  NANDN U7518 ( .A(n9913), .B(n7341), .Z(n7216) );
  NAND U7519 ( .A(n7217), .B(n7216), .Z(n7368) );
  NAND U7520 ( .A(n7218), .B(n7622), .Z(n7220) );
  XNOR U7521 ( .A(a[61]), .B(n316), .Z(n7344) );
  NAND U7522 ( .A(n7344), .B(n7620), .Z(n7219) );
  NAND U7523 ( .A(n7220), .B(n7219), .Z(n7369) );
  XOR U7524 ( .A(n7368), .B(n7369), .Z(n7370) );
  XNOR U7525 ( .A(n7371), .B(n7370), .Z(n7320) );
  XOR U7526 ( .A(n7321), .B(n7320), .Z(n7323) );
  NANDN U7527 ( .A(n7222), .B(n7221), .Z(n7226) );
  NAND U7528 ( .A(n7224), .B(n7223), .Z(n7225) );
  NAND U7529 ( .A(n7226), .B(n7225), .Z(n7322) );
  XNOR U7530 ( .A(n7323), .B(n7322), .Z(n7386) );
  NANDN U7531 ( .A(n7228), .B(n7227), .Z(n7232) );
  NANDN U7532 ( .A(n7230), .B(n7229), .Z(n7231) );
  NAND U7533 ( .A(n7232), .B(n7231), .Z(n7327) );
  NAND U7534 ( .A(n7234), .B(n7233), .Z(n7238) );
  NANDN U7535 ( .A(n7236), .B(n7235), .Z(n7237) );
  AND U7536 ( .A(n7238), .B(n7237), .Z(n7326) );
  XNOR U7537 ( .A(n7327), .B(n7326), .Z(n7328) );
  NAND U7538 ( .A(n7240), .B(n7239), .Z(n7244) );
  NAND U7539 ( .A(n7242), .B(n7241), .Z(n7243) );
  AND U7540 ( .A(n7244), .B(n7243), .Z(n7329) );
  XNOR U7541 ( .A(n7328), .B(n7329), .Z(n7387) );
  XNOR U7542 ( .A(n7386), .B(n7387), .Z(n7388) );
  XNOR U7543 ( .A(n7389), .B(n7388), .Z(n7393) );
  XNOR U7544 ( .A(n7392), .B(n7393), .Z(n7394) );
  XOR U7545 ( .A(n7395), .B(n7394), .Z(n7271) );
  NANDN U7546 ( .A(n7246), .B(n7245), .Z(n7250) );
  NANDN U7547 ( .A(n7248), .B(n7247), .Z(n7249) );
  NAND U7548 ( .A(n7250), .B(n7249), .Z(n7268) );
  NANDN U7549 ( .A(n7252), .B(n7251), .Z(n7256) );
  NAND U7550 ( .A(n7254), .B(n7253), .Z(n7255) );
  AND U7551 ( .A(n7256), .B(n7255), .Z(n7269) );
  XNOR U7552 ( .A(n7268), .B(n7269), .Z(n7270) );
  XOR U7553 ( .A(n7271), .B(n7270), .Z(n7401) );
  XNOR U7554 ( .A(n7400), .B(n7401), .Z(n7263) );
  XNOR U7555 ( .A(n7262), .B(n7263), .Z(n7264) );
  XNOR U7556 ( .A(n7265), .B(n7264), .Z(n7404) );
  XNOR U7557 ( .A(n7404), .B(sreg[95]), .Z(n7406) );
  NAND U7558 ( .A(n7257), .B(sreg[94]), .Z(n7261) );
  OR U7559 ( .A(n7259), .B(n7258), .Z(n7260) );
  AND U7560 ( .A(n7261), .B(n7260), .Z(n7405) );
  XOR U7561 ( .A(n7406), .B(n7405), .Z(c[95]) );
  NANDN U7562 ( .A(n7263), .B(n7262), .Z(n7267) );
  NAND U7563 ( .A(n7265), .B(n7264), .Z(n7266) );
  NAND U7564 ( .A(n7267), .B(n7266), .Z(n7414) );
  NANDN U7565 ( .A(n7269), .B(n7268), .Z(n7273) );
  NANDN U7566 ( .A(n7271), .B(n7270), .Z(n7272) );
  NAND U7567 ( .A(n7273), .B(n7272), .Z(n7547) );
  NANDN U7568 ( .A(n7275), .B(n7274), .Z(n7279) );
  NANDN U7569 ( .A(n7277), .B(n7276), .Z(n7278) );
  NAND U7570 ( .A(n7279), .B(n7278), .Z(n7432) );
  NANDN U7571 ( .A(n7281), .B(n7280), .Z(n7285) );
  NAND U7572 ( .A(n7283), .B(n7282), .Z(n7284) );
  NAND U7573 ( .A(n7285), .B(n7284), .Z(n7527) );
  NANDN U7574 ( .A(n7287), .B(n7286), .Z(n7291) );
  NAND U7575 ( .A(n7289), .B(n7288), .Z(n7290) );
  AND U7576 ( .A(n7291), .B(n7290), .Z(n7526) );
  XNOR U7577 ( .A(n7527), .B(n7526), .Z(n7528) );
  NAND U7578 ( .A(n9875), .B(n7292), .Z(n7295) );
  XOR U7579 ( .A(b[29]), .B(n7293), .Z(n7511) );
  OR U7580 ( .A(n7511), .B(n9874), .Z(n7294) );
  NAND U7581 ( .A(n7295), .B(n7294), .Z(n7460) );
  NANDN U7582 ( .A(n323), .B(a[32]), .Z(n7461) );
  XNOR U7583 ( .A(n7460), .B(n7461), .Z(n7462) );
  XNOR U7584 ( .A(n7463), .B(n7462), .Z(n7439) );
  NANDN U7585 ( .A(n7296), .B(n9622), .Z(n7298) );
  XOR U7586 ( .A(b[23]), .B(n8156), .Z(n7499) );
  OR U7587 ( .A(n7499), .B(n9621), .Z(n7297) );
  NAND U7588 ( .A(n7298), .B(n7297), .Z(n7517) );
  XOR U7589 ( .A(a[58]), .B(b[7]), .Z(n7490) );
  NANDN U7590 ( .A(n8013), .B(n7490), .Z(n7301) );
  NAND U7591 ( .A(n7299), .B(n8014), .Z(n7300) );
  NAND U7592 ( .A(n7301), .B(n7300), .Z(n7514) );
  XOR U7593 ( .A(b[25]), .B(n7932), .Z(n7445) );
  NANDN U7594 ( .A(n7445), .B(n9706), .Z(n7304) );
  NANDN U7595 ( .A(n7302), .B(n9707), .Z(n7303) );
  AND U7596 ( .A(n7304), .B(n7303), .Z(n7515) );
  XNOR U7597 ( .A(n7514), .B(n7515), .Z(n7516) );
  XOR U7598 ( .A(n7517), .B(n7516), .Z(n7440) );
  XOR U7599 ( .A(n7439), .B(n7440), .Z(n7442) );
  NAND U7600 ( .A(n7305), .B(n8961), .Z(n7307) );
  XNOR U7601 ( .A(n9033), .B(b[15]), .Z(n7454) );
  NAND U7602 ( .A(n7454), .B(n8963), .Z(n7306) );
  NAND U7603 ( .A(n7307), .B(n7306), .Z(n7480) );
  NAND U7604 ( .A(n7308), .B(n8286), .Z(n7310) );
  XNOR U7605 ( .A(n9357), .B(b[9]), .Z(n7484) );
  NAND U7606 ( .A(n7484), .B(n8288), .Z(n7309) );
  NAND U7607 ( .A(n7310), .B(n7309), .Z(n7478) );
  XOR U7608 ( .A(b[21]), .B(n8444), .Z(n7502) );
  NANDN U7609 ( .A(n7502), .B(n9493), .Z(n7313) );
  NANDN U7610 ( .A(n7311), .B(n9495), .Z(n7312) );
  AND U7611 ( .A(n7313), .B(n7312), .Z(n7479) );
  XOR U7612 ( .A(n7478), .B(n7479), .Z(n7481) );
  XNOR U7613 ( .A(n7480), .B(n7481), .Z(n7469) );
  XNOR U7614 ( .A(a[52]), .B(b[13]), .Z(n7496) );
  NANDN U7615 ( .A(n7496), .B(n8730), .Z(n7316) );
  NANDN U7616 ( .A(n7314), .B(n8731), .Z(n7315) );
  NAND U7617 ( .A(n7316), .B(n7315), .Z(n7467) );
  XNOR U7618 ( .A(a[54]), .B(b[11]), .Z(n7487) );
  NANDN U7619 ( .A(n7487), .B(n8541), .Z(n7319) );
  NANDN U7620 ( .A(n7317), .B(n8542), .Z(n7318) );
  AND U7621 ( .A(n7319), .B(n7318), .Z(n7466) );
  XNOR U7622 ( .A(n7467), .B(n7466), .Z(n7468) );
  XNOR U7623 ( .A(n7469), .B(n7468), .Z(n7441) );
  XNOR U7624 ( .A(n7442), .B(n7441), .Z(n7529) );
  XNOR U7625 ( .A(n7528), .B(n7529), .Z(n7429) );
  NANDN U7626 ( .A(n7321), .B(n7320), .Z(n7325) );
  OR U7627 ( .A(n7323), .B(n7322), .Z(n7324) );
  AND U7628 ( .A(n7325), .B(n7324), .Z(n7430) );
  XNOR U7629 ( .A(n7429), .B(n7430), .Z(n7431) );
  XNOR U7630 ( .A(n7432), .B(n7431), .Z(n7538) );
  NANDN U7631 ( .A(n7327), .B(n7326), .Z(n7331) );
  NAND U7632 ( .A(n7329), .B(n7328), .Z(n7330) );
  AND U7633 ( .A(n7331), .B(n7330), .Z(n7539) );
  XOR U7634 ( .A(n7538), .B(n7539), .Z(n7541) );
  OR U7635 ( .A(n7333), .B(n7332), .Z(n7337) );
  NANDN U7636 ( .A(n7335), .B(n7334), .Z(n7336) );
  NAND U7637 ( .A(n7337), .B(n7336), .Z(n7423) );
  NANDN U7638 ( .A(n7338), .B(n9105), .Z(n7340) );
  XNOR U7639 ( .A(n9455), .B(a[48]), .Z(n7451) );
  NAND U7640 ( .A(n7451), .B(n9107), .Z(n7339) );
  NAND U7641 ( .A(n7340), .B(n7339), .Z(n7474) );
  NAND U7642 ( .A(n7341), .B(n9914), .Z(n7343) );
  XNOR U7643 ( .A(n323), .B(a[34]), .Z(n7508) );
  NANDN U7644 ( .A(n9913), .B(n7508), .Z(n7342) );
  NAND U7645 ( .A(n7343), .B(n7342), .Z(n7472) );
  NAND U7646 ( .A(n7344), .B(n7622), .Z(n7346) );
  XNOR U7647 ( .A(n9810), .B(b[3]), .Z(n7448) );
  NAND U7648 ( .A(n7448), .B(n7620), .Z(n7345) );
  NAND U7649 ( .A(n7346), .B(n7345), .Z(n7473) );
  XOR U7650 ( .A(n7472), .B(n7473), .Z(n7475) );
  XNOR U7651 ( .A(n7474), .B(n7475), .Z(n7532) );
  NANDN U7652 ( .A(n7347), .B(n9379), .Z(n7349) );
  XNOR U7653 ( .A(n9562), .B(a[46]), .Z(n7493) );
  NAND U7654 ( .A(n7493), .B(n9378), .Z(n7348) );
  NAND U7655 ( .A(n7349), .B(n7348), .Z(n7522) );
  NANDN U7656 ( .A(n7350), .B(n9801), .Z(n7352) );
  XOR U7657 ( .A(n321), .B(n7672), .Z(n7457) );
  NANDN U7658 ( .A(n9751), .B(n7457), .Z(n7351) );
  NAND U7659 ( .A(n7352), .B(n7351), .Z(n7520) );
  XOR U7660 ( .A(a[60]), .B(n317), .Z(n7505) );
  NANDN U7661 ( .A(n7505), .B(n7905), .Z(n7355) );
  NANDN U7662 ( .A(n7353), .B(n7906), .Z(n7354) );
  AND U7663 ( .A(n7355), .B(n7354), .Z(n7521) );
  XNOR U7664 ( .A(n7520), .B(n7521), .Z(n7523) );
  XOR U7665 ( .A(n7522), .B(n7523), .Z(n7533) );
  XNOR U7666 ( .A(n7532), .B(n7533), .Z(n7534) );
  NANDN U7667 ( .A(n7357), .B(n7356), .Z(n7361) );
  NAND U7668 ( .A(n7359), .B(n7358), .Z(n7360) );
  AND U7669 ( .A(n7361), .B(n7360), .Z(n7535) );
  XNOR U7670 ( .A(n7534), .B(n7535), .Z(n7424) );
  XNOR U7671 ( .A(n7423), .B(n7424), .Z(n7425) );
  NANDN U7672 ( .A(n7363), .B(n7362), .Z(n7367) );
  NANDN U7673 ( .A(n7365), .B(n7364), .Z(n7366) );
  NAND U7674 ( .A(n7367), .B(n7366), .Z(n7436) );
  NAND U7675 ( .A(n7369), .B(n7368), .Z(n7373) );
  NANDN U7676 ( .A(n7371), .B(n7370), .Z(n7372) );
  NAND U7677 ( .A(n7373), .B(n7372), .Z(n7434) );
  NANDN U7678 ( .A(n7375), .B(n7374), .Z(n7379) );
  NANDN U7679 ( .A(n7377), .B(n7376), .Z(n7378) );
  AND U7680 ( .A(n7379), .B(n7378), .Z(n7433) );
  XNOR U7681 ( .A(n7434), .B(n7433), .Z(n7435) );
  XOR U7682 ( .A(n7436), .B(n7435), .Z(n7426) );
  XOR U7683 ( .A(n7425), .B(n7426), .Z(n7540) );
  XOR U7684 ( .A(n7541), .B(n7540), .Z(n7420) );
  OR U7685 ( .A(n7381), .B(n7380), .Z(n7385) );
  NAND U7686 ( .A(n7383), .B(n7382), .Z(n7384) );
  NAND U7687 ( .A(n7385), .B(n7384), .Z(n7417) );
  NANDN U7688 ( .A(n7387), .B(n7386), .Z(n7391) );
  NAND U7689 ( .A(n7389), .B(n7388), .Z(n7390) );
  NAND U7690 ( .A(n7391), .B(n7390), .Z(n7418) );
  XNOR U7691 ( .A(n7417), .B(n7418), .Z(n7419) );
  XNOR U7692 ( .A(n7420), .B(n7419), .Z(n7545) );
  NANDN U7693 ( .A(n7393), .B(n7392), .Z(n7397) );
  NAND U7694 ( .A(n7395), .B(n7394), .Z(n7396) );
  AND U7695 ( .A(n7397), .B(n7396), .Z(n7544) );
  XNOR U7696 ( .A(n7545), .B(n7544), .Z(n7546) );
  XNOR U7697 ( .A(n7547), .B(n7546), .Z(n7411) );
  NANDN U7698 ( .A(n7399), .B(n7398), .Z(n7403) );
  NANDN U7699 ( .A(n7401), .B(n7400), .Z(n7402) );
  NAND U7700 ( .A(n7403), .B(n7402), .Z(n7412) );
  XNOR U7701 ( .A(n7411), .B(n7412), .Z(n7413) );
  XOR U7702 ( .A(n7414), .B(n7413), .Z(n7410) );
  NAND U7703 ( .A(n7404), .B(sreg[95]), .Z(n7408) );
  OR U7704 ( .A(n7406), .B(n7405), .Z(n7407) );
  AND U7705 ( .A(n7408), .B(n7407), .Z(n7409) );
  XOR U7706 ( .A(n7410), .B(n7409), .Z(c[96]) );
  OR U7707 ( .A(n7410), .B(n7409), .Z(n7551) );
  NANDN U7708 ( .A(n7412), .B(n7411), .Z(n7416) );
  NAND U7709 ( .A(n7414), .B(n7413), .Z(n7415) );
  NAND U7710 ( .A(n7416), .B(n7415), .Z(n7555) );
  NANDN U7711 ( .A(n7418), .B(n7417), .Z(n7422) );
  NAND U7712 ( .A(n7420), .B(n7419), .Z(n7421) );
  NAND U7713 ( .A(n7422), .B(n7421), .Z(n7689) );
  NANDN U7714 ( .A(n7424), .B(n7423), .Z(n7428) );
  NAND U7715 ( .A(n7426), .B(n7425), .Z(n7427) );
  NAND U7716 ( .A(n7428), .B(n7427), .Z(n7558) );
  XNOR U7717 ( .A(n7558), .B(n7559), .Z(n7560) );
  NANDN U7718 ( .A(n7434), .B(n7433), .Z(n7438) );
  NAND U7719 ( .A(n7436), .B(n7435), .Z(n7437) );
  NAND U7720 ( .A(n7438), .B(n7437), .Z(n7681) );
  NANDN U7721 ( .A(n7440), .B(n7439), .Z(n7444) );
  NANDN U7722 ( .A(n7442), .B(n7441), .Z(n7443) );
  NAND U7723 ( .A(n7444), .B(n7443), .Z(n7637) );
  XNOR U7724 ( .A(b[25]), .B(a[41]), .Z(n7597) );
  NANDN U7725 ( .A(n7597), .B(n9706), .Z(n7447) );
  NANDN U7726 ( .A(n7445), .B(n9707), .Z(n7446) );
  AND U7727 ( .A(n7447), .B(n7446), .Z(n7573) );
  NAND U7728 ( .A(n7448), .B(n7622), .Z(n7450) );
  XOR U7729 ( .A(n9946), .B(n316), .Z(n7621) );
  NAND U7730 ( .A(n7621), .B(n7620), .Z(n7449) );
  AND U7731 ( .A(n7450), .B(n7449), .Z(n7571) );
  NAND U7732 ( .A(n7451), .B(n9105), .Z(n7453) );
  XNOR U7733 ( .A(n9455), .B(a[49]), .Z(n7617) );
  NAND U7734 ( .A(n7617), .B(n9107), .Z(n7452) );
  NAND U7735 ( .A(n7453), .B(n7452), .Z(n7570) );
  XOR U7736 ( .A(n7573), .B(n7572), .Z(n7601) );
  NAND U7737 ( .A(n7454), .B(n8961), .Z(n7456) );
  XNOR U7738 ( .A(n9457), .B(b[15]), .Z(n7665) );
  NAND U7739 ( .A(n7665), .B(n8963), .Z(n7455) );
  NAND U7740 ( .A(n7456), .B(n7455), .Z(n7606) );
  XOR U7741 ( .A(b[1]), .B(n7606), .Z(n7608) );
  XOR U7742 ( .A(n321), .B(a[39]), .Z(n7614) );
  OR U7743 ( .A(n7614), .B(n9751), .Z(n7459) );
  NAND U7744 ( .A(n9801), .B(n7457), .Z(n7458) );
  AND U7745 ( .A(n7459), .B(n7458), .Z(n7607) );
  XNOR U7746 ( .A(n7608), .B(n7607), .Z(n7600) );
  XOR U7747 ( .A(n7601), .B(n7600), .Z(n7602) );
  NANDN U7748 ( .A(n7461), .B(n7460), .Z(n7465) );
  NAND U7749 ( .A(n7463), .B(n7462), .Z(n7464) );
  AND U7750 ( .A(n7465), .B(n7464), .Z(n7603) );
  XNOR U7751 ( .A(n7602), .B(n7603), .Z(n7638) );
  XNOR U7752 ( .A(n7637), .B(n7638), .Z(n7639) );
  NANDN U7753 ( .A(n7467), .B(n7466), .Z(n7471) );
  NANDN U7754 ( .A(n7469), .B(n7468), .Z(n7470) );
  NAND U7755 ( .A(n7471), .B(n7470), .Z(n7656) );
  NAND U7756 ( .A(n7473), .B(n7472), .Z(n7477) );
  NAND U7757 ( .A(n7475), .B(n7474), .Z(n7476) );
  NAND U7758 ( .A(n7477), .B(n7476), .Z(n7654) );
  NANDN U7759 ( .A(n7479), .B(n7478), .Z(n7483) );
  NANDN U7760 ( .A(n7481), .B(n7480), .Z(n7482) );
  AND U7761 ( .A(n7483), .B(n7482), .Z(n7653) );
  XNOR U7762 ( .A(n7654), .B(n7653), .Z(n7655) );
  XOR U7763 ( .A(n7656), .B(n7655), .Z(n7640) );
  XOR U7764 ( .A(n7639), .B(n7640), .Z(n7680) );
  XNOR U7765 ( .A(n7681), .B(n7680), .Z(n7683) );
  NAND U7766 ( .A(n7484), .B(n8286), .Z(n7486) );
  XOR U7767 ( .A(a[57]), .B(b[9]), .Z(n7582) );
  NAND U7768 ( .A(n7582), .B(n8288), .Z(n7485) );
  NAND U7769 ( .A(n7486), .B(n7485), .Z(n7566) );
  XOR U7770 ( .A(a[55]), .B(b[11]), .Z(n7594) );
  NAND U7771 ( .A(n7594), .B(n8541), .Z(n7489) );
  NANDN U7772 ( .A(n7487), .B(n8542), .Z(n7488) );
  AND U7773 ( .A(n7489), .B(n7488), .Z(n7564) );
  XOR U7774 ( .A(a[59]), .B(b[7]), .Z(n7585) );
  NANDN U7775 ( .A(n8013), .B(n7585), .Z(n7492) );
  NAND U7776 ( .A(n7490), .B(n8014), .Z(n7491) );
  NAND U7777 ( .A(n7492), .B(n7491), .Z(n7579) );
  NAND U7778 ( .A(n7493), .B(n9379), .Z(n7495) );
  XNOR U7779 ( .A(n9562), .B(a[47]), .Z(n7625) );
  NAND U7780 ( .A(n7625), .B(n9378), .Z(n7494) );
  NAND U7781 ( .A(n7495), .B(n7494), .Z(n7576) );
  XNOR U7782 ( .A(a[53]), .B(b[13]), .Z(n7591) );
  NANDN U7783 ( .A(n7591), .B(n8730), .Z(n7498) );
  NANDN U7784 ( .A(n7496), .B(n8731), .Z(n7497) );
  AND U7785 ( .A(n7498), .B(n7497), .Z(n7577) );
  XNOR U7786 ( .A(n7576), .B(n7577), .Z(n7578) );
  XNOR U7787 ( .A(n7579), .B(n7578), .Z(n7565) );
  XOR U7788 ( .A(n7566), .B(n7567), .Z(n7633) );
  NANDN U7789 ( .A(n7499), .B(n9622), .Z(n7501) );
  XNOR U7790 ( .A(n319), .B(a[43]), .Z(n7611) );
  NANDN U7791 ( .A(n9621), .B(n7611), .Z(n7500) );
  NAND U7792 ( .A(n7501), .B(n7500), .Z(n7662) );
  XNOR U7793 ( .A(b[21]), .B(a[45]), .Z(n7588) );
  NANDN U7794 ( .A(n7588), .B(n9493), .Z(n7504) );
  NANDN U7795 ( .A(n7502), .B(n9495), .Z(n7503) );
  NAND U7796 ( .A(n7504), .B(n7503), .Z(n7659) );
  XNOR U7797 ( .A(a[61]), .B(b[5]), .Z(n7628) );
  NANDN U7798 ( .A(n7628), .B(n7905), .Z(n7507) );
  NANDN U7799 ( .A(n7505), .B(n7906), .Z(n7506) );
  AND U7800 ( .A(n7507), .B(n7506), .Z(n7660) );
  XNOR U7801 ( .A(n7659), .B(n7660), .Z(n7661) );
  XOR U7802 ( .A(n7662), .B(n7661), .Z(n7632) );
  NAND U7803 ( .A(n7508), .B(n9914), .Z(n7510) );
  XNOR U7804 ( .A(n323), .B(a[35]), .Z(n7668) );
  NANDN U7805 ( .A(n9913), .B(n7668), .Z(n7509) );
  NAND U7806 ( .A(n7510), .B(n7509), .Z(n7676) );
  ANDN U7807 ( .B(a[33]), .A(n323), .Z(n7785) );
  IV U7808 ( .A(n7785), .Z(n7868) );
  NANDN U7809 ( .A(n7511), .B(n9875), .Z(n7513) );
  XNOR U7810 ( .A(n322), .B(a[37]), .Z(n7671) );
  NANDN U7811 ( .A(n9874), .B(n7671), .Z(n7512) );
  AND U7812 ( .A(n7513), .B(n7512), .Z(n7675) );
  XOR U7813 ( .A(n7868), .B(n7675), .Z(n7677) );
  XOR U7814 ( .A(n7676), .B(n7677), .Z(n7631) );
  XOR U7815 ( .A(n7632), .B(n7631), .Z(n7634) );
  XNOR U7816 ( .A(n7633), .B(n7634), .Z(n7650) );
  NANDN U7817 ( .A(n7515), .B(n7514), .Z(n7519) );
  NAND U7818 ( .A(n7517), .B(n7516), .Z(n7518) );
  NAND U7819 ( .A(n7519), .B(n7518), .Z(n7648) );
  NANDN U7820 ( .A(n7521), .B(n7520), .Z(n7525) );
  NAND U7821 ( .A(n7523), .B(n7522), .Z(n7524) );
  AND U7822 ( .A(n7525), .B(n7524), .Z(n7647) );
  XNOR U7823 ( .A(n7648), .B(n7647), .Z(n7649) );
  XNOR U7824 ( .A(n7650), .B(n7649), .Z(n7645) );
  NANDN U7825 ( .A(n7527), .B(n7526), .Z(n7531) );
  NAND U7826 ( .A(n7529), .B(n7528), .Z(n7530) );
  NAND U7827 ( .A(n7531), .B(n7530), .Z(n7643) );
  NANDN U7828 ( .A(n7533), .B(n7532), .Z(n7537) );
  NAND U7829 ( .A(n7535), .B(n7534), .Z(n7536) );
  AND U7830 ( .A(n7537), .B(n7536), .Z(n7644) );
  XNOR U7831 ( .A(n7643), .B(n7644), .Z(n7646) );
  XOR U7832 ( .A(n7645), .B(n7646), .Z(n7682) );
  XOR U7833 ( .A(n7683), .B(n7682), .Z(n7561) );
  XOR U7834 ( .A(n7560), .B(n7561), .Z(n7686) );
  NANDN U7835 ( .A(n7539), .B(n7538), .Z(n7543) );
  NANDN U7836 ( .A(n7541), .B(n7540), .Z(n7542) );
  NAND U7837 ( .A(n7543), .B(n7542), .Z(n7687) );
  XNOR U7838 ( .A(n7686), .B(n7687), .Z(n7688) );
  XNOR U7839 ( .A(n7689), .B(n7688), .Z(n7552) );
  NANDN U7840 ( .A(n7545), .B(n7544), .Z(n7549) );
  NAND U7841 ( .A(n7547), .B(n7546), .Z(n7548) );
  NAND U7842 ( .A(n7549), .B(n7548), .Z(n7553) );
  XNOR U7843 ( .A(n7552), .B(n7553), .Z(n7554) );
  XOR U7844 ( .A(n7555), .B(n7554), .Z(n7550) );
  XOR U7845 ( .A(n7551), .B(n7550), .Z(c[97]) );
  OR U7846 ( .A(n7551), .B(n7550), .Z(n7832) );
  NANDN U7847 ( .A(n7553), .B(n7552), .Z(n7557) );
  NAND U7848 ( .A(n7555), .B(n7554), .Z(n7556) );
  NAND U7849 ( .A(n7557), .B(n7556), .Z(n7695) );
  NANDN U7850 ( .A(n7559), .B(n7558), .Z(n7563) );
  NANDN U7851 ( .A(n7561), .B(n7560), .Z(n7562) );
  NAND U7852 ( .A(n7563), .B(n7562), .Z(n7700) );
  OR U7853 ( .A(n7565), .B(n7564), .Z(n7569) );
  NAND U7854 ( .A(n7567), .B(n7566), .Z(n7568) );
  NAND U7855 ( .A(n7569), .B(n7568), .Z(n7706) );
  NANDN U7856 ( .A(n7571), .B(n7570), .Z(n7575) );
  NANDN U7857 ( .A(n7573), .B(n7572), .Z(n7574) );
  NAND U7858 ( .A(n7575), .B(n7574), .Z(n7705) );
  NANDN U7859 ( .A(n7577), .B(n7576), .Z(n7581) );
  NAND U7860 ( .A(n7579), .B(n7578), .Z(n7580) );
  NAND U7861 ( .A(n7581), .B(n7580), .Z(n7770) );
  NAND U7862 ( .A(n7582), .B(n8286), .Z(n7584) );
  XOR U7863 ( .A(a[58]), .B(b[9]), .Z(n7747) );
  NAND U7864 ( .A(n7747), .B(n8288), .Z(n7583) );
  NAND U7865 ( .A(n7584), .B(n7583), .Z(n7802) );
  XNOR U7866 ( .A(a[60]), .B(b[7]), .Z(n7723) );
  OR U7867 ( .A(n7723), .B(n8013), .Z(n7587) );
  NAND U7868 ( .A(n8014), .B(n7585), .Z(n7586) );
  NAND U7869 ( .A(n7587), .B(n7586), .Z(n7800) );
  XOR U7870 ( .A(b[21]), .B(n8654), .Z(n7729) );
  NANDN U7871 ( .A(n7729), .B(n9493), .Z(n7590) );
  NANDN U7872 ( .A(n7588), .B(n9495), .Z(n7589) );
  AND U7873 ( .A(n7590), .B(n7589), .Z(n7801) );
  XOR U7874 ( .A(n7800), .B(n7801), .Z(n7803) );
  XOR U7875 ( .A(n7802), .B(n7803), .Z(n7768) );
  XNOR U7876 ( .A(a[54]), .B(b[13]), .Z(n7773) );
  NANDN U7877 ( .A(n7773), .B(n8730), .Z(n7593) );
  NANDN U7878 ( .A(n7591), .B(n8731), .Z(n7592) );
  NAND U7879 ( .A(n7593), .B(n7592), .Z(n7741) );
  XNOR U7880 ( .A(a[56]), .B(b[11]), .Z(n7714) );
  NANDN U7881 ( .A(n7714), .B(n8541), .Z(n7596) );
  NAND U7882 ( .A(n7594), .B(n8542), .Z(n7595) );
  NAND U7883 ( .A(n7596), .B(n7595), .Z(n7738) );
  XOR U7884 ( .A(b[25]), .B(n8156), .Z(n7717) );
  NANDN U7885 ( .A(n7717), .B(n9706), .Z(n7599) );
  NANDN U7886 ( .A(n7597), .B(n9707), .Z(n7598) );
  AND U7887 ( .A(n7599), .B(n7598), .Z(n7739) );
  XNOR U7888 ( .A(n7738), .B(n7739), .Z(n7740) );
  XNOR U7889 ( .A(n7741), .B(n7740), .Z(n7767) );
  XOR U7890 ( .A(n7768), .B(n7767), .Z(n7769) );
  XNOR U7891 ( .A(n7770), .B(n7769), .Z(n7704) );
  XOR U7892 ( .A(n7705), .B(n7704), .Z(n7707) );
  XNOR U7893 ( .A(n7706), .B(n7707), .Z(n7825) );
  NAND U7894 ( .A(n7601), .B(n7600), .Z(n7605) );
  NAND U7895 ( .A(n7603), .B(n7602), .Z(n7604) );
  NAND U7896 ( .A(n7605), .B(n7604), .Z(n7808) );
  NANDN U7897 ( .A(n7606), .B(b[1]), .Z(n7610) );
  NANDN U7898 ( .A(n7608), .B(n7607), .Z(n7609) );
  NAND U7899 ( .A(n7610), .B(n7609), .Z(n7713) );
  XOR U7900 ( .A(b[23]), .B(n8444), .Z(n7744) );
  OR U7901 ( .A(n7744), .B(n9621), .Z(n7613) );
  NAND U7902 ( .A(n9622), .B(n7611), .Z(n7612) );
  NAND U7903 ( .A(n7613), .B(n7612), .Z(n7790) );
  XOR U7904 ( .A(b[27]), .B(n7932), .Z(n7720) );
  OR U7905 ( .A(n7720), .B(n9751), .Z(n7616) );
  NANDN U7906 ( .A(n7614), .B(n9801), .Z(n7615) );
  NAND U7907 ( .A(n7616), .B(n7615), .Z(n7789) );
  NAND U7908 ( .A(n7617), .B(n9105), .Z(n7619) );
  XNOR U7909 ( .A(n9033), .B(b[17]), .Z(n7779) );
  NAND U7910 ( .A(n7779), .B(n9107), .Z(n7618) );
  NAND U7911 ( .A(n7619), .B(n7618), .Z(n7788) );
  XOR U7912 ( .A(n7789), .B(n7788), .Z(n7791) );
  XNOR U7913 ( .A(n7790), .B(n7791), .Z(n7710) );
  NANDN U7914 ( .A(n316), .B(n7620), .Z(n7624) );
  NAND U7915 ( .A(n7622), .B(n7621), .Z(n7623) );
  NAND U7916 ( .A(n7624), .B(n7623), .Z(n7782) );
  NANDN U7917 ( .A(n323), .B(a[34]), .Z(n7783) );
  XNOR U7918 ( .A(n7782), .B(n7783), .Z(n7784) );
  XNOR U7919 ( .A(n7868), .B(n7784), .Z(n7797) );
  NAND U7920 ( .A(n7625), .B(n9379), .Z(n7627) );
  XNOR U7921 ( .A(n9562), .B(a[48]), .Z(n7753) );
  NAND U7922 ( .A(n7753), .B(n9378), .Z(n7626) );
  NAND U7923 ( .A(n7627), .B(n7626), .Z(n7795) );
  XOR U7924 ( .A(n9810), .B(n317), .Z(n7758) );
  NAND U7925 ( .A(n7758), .B(n7905), .Z(n7630) );
  NANDN U7926 ( .A(n7628), .B(n7906), .Z(n7629) );
  AND U7927 ( .A(n7630), .B(n7629), .Z(n7794) );
  XNOR U7928 ( .A(n7795), .B(n7794), .Z(n7796) );
  XNOR U7929 ( .A(n7797), .B(n7796), .Z(n7711) );
  XNOR U7930 ( .A(n7710), .B(n7711), .Z(n7712) );
  XNOR U7931 ( .A(n7713), .B(n7712), .Z(n7806) );
  NANDN U7932 ( .A(n7632), .B(n7631), .Z(n7636) );
  OR U7933 ( .A(n7634), .B(n7633), .Z(n7635) );
  NAND U7934 ( .A(n7636), .B(n7635), .Z(n7807) );
  XOR U7935 ( .A(n7806), .B(n7807), .Z(n7809) );
  XOR U7936 ( .A(n7808), .B(n7809), .Z(n7824) );
  XNOR U7937 ( .A(n7825), .B(n7824), .Z(n7827) );
  NANDN U7938 ( .A(n7638), .B(n7637), .Z(n7642) );
  NAND U7939 ( .A(n7640), .B(n7639), .Z(n7641) );
  NAND U7940 ( .A(n7642), .B(n7641), .Z(n7826) );
  XNOR U7941 ( .A(n7827), .B(n7826), .Z(n7821) );
  NANDN U7942 ( .A(n7648), .B(n7647), .Z(n7652) );
  NANDN U7943 ( .A(n7650), .B(n7649), .Z(n7651) );
  NAND U7944 ( .A(n7652), .B(n7651), .Z(n7814) );
  NANDN U7945 ( .A(n7654), .B(n7653), .Z(n7658) );
  NAND U7946 ( .A(n7656), .B(n7655), .Z(n7657) );
  NAND U7947 ( .A(n7658), .B(n7657), .Z(n7813) );
  NANDN U7948 ( .A(n7660), .B(n7659), .Z(n7664) );
  NAND U7949 ( .A(n7662), .B(n7661), .Z(n7663) );
  NAND U7950 ( .A(n7664), .B(n7663), .Z(n7764) );
  NAND U7951 ( .A(n7665), .B(n8961), .Z(n7667) );
  XNOR U7952 ( .A(n9217), .B(b[15]), .Z(n7776) );
  NAND U7953 ( .A(n7776), .B(n8963), .Z(n7666) );
  NAND U7954 ( .A(n7667), .B(n7666), .Z(n7734) );
  NAND U7955 ( .A(n7668), .B(n9914), .Z(n7670) );
  XNOR U7956 ( .A(n323), .B(a[36]), .Z(n7726) );
  NANDN U7957 ( .A(n9913), .B(n7726), .Z(n7669) );
  NAND U7958 ( .A(n7670), .B(n7669), .Z(n7732) );
  NAND U7959 ( .A(n7671), .B(n9875), .Z(n7674) );
  XOR U7960 ( .A(n322), .B(n7672), .Z(n7750) );
  NANDN U7961 ( .A(n9874), .B(n7750), .Z(n7673) );
  AND U7962 ( .A(n7674), .B(n7673), .Z(n7733) );
  XOR U7963 ( .A(n7732), .B(n7733), .Z(n7735) );
  XNOR U7964 ( .A(n7734), .B(n7735), .Z(n7762) );
  NANDN U7965 ( .A(n7868), .B(n7675), .Z(n7679) );
  OR U7966 ( .A(n7677), .B(n7676), .Z(n7678) );
  AND U7967 ( .A(n7679), .B(n7678), .Z(n7761) );
  XOR U7968 ( .A(n7762), .B(n7761), .Z(n7763) );
  XNOR U7969 ( .A(n7764), .B(n7763), .Z(n7812) );
  XNOR U7970 ( .A(n7813), .B(n7812), .Z(n7815) );
  XNOR U7971 ( .A(n7814), .B(n7815), .Z(n7818) );
  XOR U7972 ( .A(n7819), .B(n7818), .Z(n7820) );
  XNOR U7973 ( .A(n7821), .B(n7820), .Z(n7698) );
  NAND U7974 ( .A(n7681), .B(n7680), .Z(n7685) );
  NANDN U7975 ( .A(n7683), .B(n7682), .Z(n7684) );
  NAND U7976 ( .A(n7685), .B(n7684), .Z(n7699) );
  XOR U7977 ( .A(n7698), .B(n7699), .Z(n7701) );
  XNOR U7978 ( .A(n7700), .B(n7701), .Z(n7692) );
  NANDN U7979 ( .A(n7687), .B(n7686), .Z(n7691) );
  NAND U7980 ( .A(n7689), .B(n7688), .Z(n7690) );
  NAND U7981 ( .A(n7691), .B(n7690), .Z(n7693) );
  XNOR U7982 ( .A(n7692), .B(n7693), .Z(n7694) );
  XOR U7983 ( .A(n7695), .B(n7694), .Z(n7831) );
  XOR U7984 ( .A(n7832), .B(n7831), .Z(c[98]) );
  NANDN U7985 ( .A(n7693), .B(n7692), .Z(n7697) );
  NAND U7986 ( .A(n7695), .B(n7694), .Z(n7696) );
  NAND U7987 ( .A(n7697), .B(n7696), .Z(n7837) );
  NANDN U7988 ( .A(n7699), .B(n7698), .Z(n7703) );
  OR U7989 ( .A(n7701), .B(n7700), .Z(n7702) );
  NAND U7990 ( .A(n7703), .B(n7702), .Z(n7835) );
  NANDN U7991 ( .A(n7705), .B(n7704), .Z(n7709) );
  OR U7992 ( .A(n7707), .B(n7706), .Z(n7708) );
  NAND U7993 ( .A(n7709), .B(n7708), .Z(n7845) );
  XOR U7994 ( .A(a[57]), .B(b[11]), .Z(n7922) );
  NAND U7995 ( .A(n7922), .B(n8541), .Z(n7716) );
  NANDN U7996 ( .A(n7714), .B(n8542), .Z(n7715) );
  NAND U7997 ( .A(n7716), .B(n7715), .Z(n7913) );
  XNOR U7998 ( .A(b[25]), .B(a[43]), .Z(n7919) );
  NANDN U7999 ( .A(n7919), .B(n9706), .Z(n7719) );
  NANDN U8000 ( .A(n7717), .B(n9707), .Z(n7718) );
  NAND U8001 ( .A(n7719), .B(n7718), .Z(n7910) );
  NANDN U8002 ( .A(n7720), .B(n9801), .Z(n7722) );
  XNOR U8003 ( .A(b[27]), .B(a[41]), .Z(n7899) );
  OR U8004 ( .A(n7899), .B(n9751), .Z(n7721) );
  AND U8005 ( .A(n7722), .B(n7721), .Z(n7911) );
  XNOR U8006 ( .A(n7910), .B(n7911), .Z(n7912) );
  XNOR U8007 ( .A(n7913), .B(n7912), .Z(n7953) );
  XOR U8008 ( .A(a[61]), .B(b[7]), .Z(n7925) );
  NANDN U8009 ( .A(n8013), .B(n7925), .Z(n7725) );
  NANDN U8010 ( .A(n7723), .B(n8014), .Z(n7724) );
  NAND U8011 ( .A(n7725), .B(n7724), .Z(n7859) );
  NAND U8012 ( .A(n7726), .B(n9914), .Z(n7728) );
  XNOR U8013 ( .A(n323), .B(a[37]), .Z(n7902) );
  NANDN U8014 ( .A(n9913), .B(n7902), .Z(n7727) );
  NAND U8015 ( .A(n7728), .B(n7727), .Z(n7856) );
  XNOR U8016 ( .A(b[21]), .B(a[47]), .Z(n7893) );
  NANDN U8017 ( .A(n7893), .B(n9493), .Z(n7731) );
  NANDN U8018 ( .A(n7729), .B(n9495), .Z(n7730) );
  AND U8019 ( .A(n7731), .B(n7730), .Z(n7857) );
  XNOR U8020 ( .A(n7856), .B(n7857), .Z(n7858) );
  XOR U8021 ( .A(n7859), .B(n7858), .Z(n7954) );
  XNOR U8022 ( .A(n7953), .B(n7954), .Z(n7955) );
  NANDN U8023 ( .A(n7733), .B(n7732), .Z(n7737) );
  NANDN U8024 ( .A(n7735), .B(n7734), .Z(n7736) );
  AND U8025 ( .A(n7737), .B(n7736), .Z(n7956) );
  XOR U8026 ( .A(n7955), .B(n7956), .Z(n7850) );
  NANDN U8027 ( .A(n7739), .B(n7738), .Z(n7743) );
  NAND U8028 ( .A(n7741), .B(n7740), .Z(n7742) );
  NAND U8029 ( .A(n7743), .B(n7742), .Z(n7950) );
  NANDN U8030 ( .A(n7744), .B(n9622), .Z(n7746) );
  XNOR U8031 ( .A(b[23]), .B(a[45]), .Z(n7916) );
  OR U8032 ( .A(n7916), .B(n9621), .Z(n7745) );
  NAND U8033 ( .A(n7746), .B(n7745), .Z(n7892) );
  NAND U8034 ( .A(n7747), .B(n8286), .Z(n7749) );
  XOR U8035 ( .A(a[59]), .B(b[9]), .Z(n7896) );
  NAND U8036 ( .A(n7896), .B(n8288), .Z(n7748) );
  NAND U8037 ( .A(n7749), .B(n7748), .Z(n7889) );
  NAND U8038 ( .A(n9875), .B(n7750), .Z(n7752) );
  XNOR U8039 ( .A(n322), .B(a[39]), .Z(n7931) );
  NANDN U8040 ( .A(n9874), .B(n7931), .Z(n7751) );
  AND U8041 ( .A(n7752), .B(n7751), .Z(n7890) );
  XNOR U8042 ( .A(n7889), .B(n7890), .Z(n7891) );
  XNOR U8043 ( .A(n7892), .B(n7891), .Z(n7948) );
  NAND U8044 ( .A(n7753), .B(n9379), .Z(n7755) );
  XNOR U8045 ( .A(n9562), .B(a[49]), .Z(n7928) );
  NAND U8046 ( .A(n7928), .B(n9378), .Z(n7754) );
  NAND U8047 ( .A(n7755), .B(n7754), .Z(n7864) );
  NANDN U8048 ( .A(n323), .B(a[35]), .Z(n7871) );
  NANDN U8049 ( .A(n7756), .B(b[1]), .Z(n7757) );
  ANDN U8050 ( .B(n7757), .A(n316), .Z(n7869) );
  XNOR U8051 ( .A(n7868), .B(n7869), .Z(n7870) );
  XNOR U8052 ( .A(n7871), .B(n7870), .Z(n7862) );
  XOR U8053 ( .A(n9946), .B(b[5]), .Z(n7907) );
  NANDN U8054 ( .A(n7907), .B(n7905), .Z(n7760) );
  NAND U8055 ( .A(n7906), .B(n7758), .Z(n7759) );
  NAND U8056 ( .A(n7760), .B(n7759), .Z(n7863) );
  XOR U8057 ( .A(n7862), .B(n7863), .Z(n7865) );
  XOR U8058 ( .A(n7864), .B(n7865), .Z(n7947) );
  XNOR U8059 ( .A(n7948), .B(n7947), .Z(n7949) );
  XOR U8060 ( .A(n7950), .B(n7949), .Z(n7851) );
  XOR U8061 ( .A(n7850), .B(n7851), .Z(n7852) );
  XOR U8062 ( .A(n7853), .B(n7852), .Z(n7844) );
  XNOR U8063 ( .A(n7845), .B(n7844), .Z(n7847) );
  OR U8064 ( .A(n7762), .B(n7761), .Z(n7766) );
  NANDN U8065 ( .A(n7764), .B(n7763), .Z(n7765) );
  NAND U8066 ( .A(n7766), .B(n7765), .Z(n7962) );
  NAND U8067 ( .A(n7768), .B(n7767), .Z(n7772) );
  NANDN U8068 ( .A(n7770), .B(n7769), .Z(n7771) );
  NAND U8069 ( .A(n7772), .B(n7771), .Z(n7960) );
  XOR U8070 ( .A(a[55]), .B(b[13]), .Z(n7880) );
  NAND U8071 ( .A(n7880), .B(n8730), .Z(n7775) );
  NANDN U8072 ( .A(n7773), .B(n8731), .Z(n7774) );
  NAND U8073 ( .A(n7775), .B(n7774), .Z(n7886) );
  NAND U8074 ( .A(n7776), .B(n8961), .Z(n7778) );
  XNOR U8075 ( .A(n9564), .B(b[15]), .Z(n7874) );
  NAND U8076 ( .A(n7874), .B(n8963), .Z(n7777) );
  NAND U8077 ( .A(n7778), .B(n7777), .Z(n7883) );
  NAND U8078 ( .A(n7779), .B(n9105), .Z(n7781) );
  XNOR U8079 ( .A(n9455), .B(a[51]), .Z(n7877) );
  NAND U8080 ( .A(n7877), .B(n9107), .Z(n7780) );
  NAND U8081 ( .A(n7781), .B(n7780), .Z(n7884) );
  XOR U8082 ( .A(n7883), .B(n7884), .Z(n7885) );
  XNOR U8083 ( .A(n7886), .B(n7885), .Z(n7938) );
  NANDN U8084 ( .A(n7783), .B(n7782), .Z(n7787) );
  NANDN U8085 ( .A(n7785), .B(n7784), .Z(n7786) );
  NAND U8086 ( .A(n7787), .B(n7786), .Z(n7936) );
  NAND U8087 ( .A(n7789), .B(n7788), .Z(n7793) );
  NAND U8088 ( .A(n7791), .B(n7790), .Z(n7792) );
  AND U8089 ( .A(n7793), .B(n7792), .Z(n7935) );
  XNOR U8090 ( .A(n7936), .B(n7935), .Z(n7937) );
  XNOR U8091 ( .A(n7938), .B(n7937), .Z(n7944) );
  NANDN U8092 ( .A(n7795), .B(n7794), .Z(n7799) );
  NAND U8093 ( .A(n7797), .B(n7796), .Z(n7798) );
  NAND U8094 ( .A(n7799), .B(n7798), .Z(n7942) );
  NANDN U8095 ( .A(n7801), .B(n7800), .Z(n7805) );
  NANDN U8096 ( .A(n7803), .B(n7802), .Z(n7804) );
  AND U8097 ( .A(n7805), .B(n7804), .Z(n7941) );
  XOR U8098 ( .A(n7942), .B(n7941), .Z(n7943) );
  XNOR U8099 ( .A(n7944), .B(n7943), .Z(n7959) );
  XOR U8100 ( .A(n7960), .B(n7959), .Z(n7961) );
  XOR U8101 ( .A(n7962), .B(n7961), .Z(n7846) );
  XOR U8102 ( .A(n7847), .B(n7846), .Z(n7841) );
  NANDN U8103 ( .A(n7807), .B(n7806), .Z(n7811) );
  OR U8104 ( .A(n7809), .B(n7808), .Z(n7810) );
  NAND U8105 ( .A(n7811), .B(n7810), .Z(n7838) );
  NAND U8106 ( .A(n7813), .B(n7812), .Z(n7817) );
  NANDN U8107 ( .A(n7815), .B(n7814), .Z(n7816) );
  NAND U8108 ( .A(n7817), .B(n7816), .Z(n7839) );
  XNOR U8109 ( .A(n7838), .B(n7839), .Z(n7840) );
  XNOR U8110 ( .A(n7841), .B(n7840), .Z(n7968) );
  NAND U8111 ( .A(n7819), .B(n7818), .Z(n7823) );
  NAND U8112 ( .A(n7821), .B(n7820), .Z(n7822) );
  NAND U8113 ( .A(n7823), .B(n7822), .Z(n7965) );
  NAND U8114 ( .A(n7825), .B(n7824), .Z(n7829) );
  OR U8115 ( .A(n7827), .B(n7826), .Z(n7828) );
  NAND U8116 ( .A(n7829), .B(n7828), .Z(n7966) );
  XNOR U8117 ( .A(n7965), .B(n7966), .Z(n7967) );
  XNOR U8118 ( .A(n7968), .B(n7967), .Z(n7836) );
  XNOR U8119 ( .A(n7835), .B(n7836), .Z(n7830) );
  XNOR U8120 ( .A(n7837), .B(n7830), .Z(n7834) );
  OR U8121 ( .A(n7832), .B(n7831), .Z(n7833) );
  XOR U8122 ( .A(n7834), .B(n7833), .Z(c[99]) );
  OR U8123 ( .A(n7834), .B(n7833), .Z(n7973) );
  NANDN U8124 ( .A(n7839), .B(n7838), .Z(n7843) );
  NAND U8125 ( .A(n7841), .B(n7840), .Z(n7842) );
  NAND U8126 ( .A(n7843), .B(n7842), .Z(n8096) );
  NAND U8127 ( .A(n7845), .B(n7844), .Z(n7849) );
  NANDN U8128 ( .A(n7847), .B(n7846), .Z(n7848) );
  AND U8129 ( .A(n7849), .B(n7848), .Z(n8093) );
  NAND U8130 ( .A(n7851), .B(n7850), .Z(n7855) );
  NAND U8131 ( .A(n7853), .B(n7852), .Z(n7854) );
  NAND U8132 ( .A(n7855), .B(n7854), .Z(n8068) );
  NANDN U8133 ( .A(n7857), .B(n7856), .Z(n7861) );
  NAND U8134 ( .A(n7859), .B(n7858), .Z(n7860) );
  NAND U8135 ( .A(n7861), .B(n7860), .Z(n8087) );
  NANDN U8136 ( .A(n7863), .B(n7862), .Z(n7867) );
  OR U8137 ( .A(n7865), .B(n7864), .Z(n7866) );
  NAND U8138 ( .A(n7867), .B(n7866), .Z(n8088) );
  XNOR U8139 ( .A(n8087), .B(n8088), .Z(n8089) );
  OR U8140 ( .A(n7869), .B(n7868), .Z(n7873) );
  OR U8141 ( .A(n7871), .B(n7870), .Z(n7872) );
  AND U8142 ( .A(n7873), .B(n7872), .Z(n8060) );
  NAND U8143 ( .A(n7874), .B(n8961), .Z(n7876) );
  XNOR U8144 ( .A(n9353), .B(b[15]), .Z(n7995) );
  NAND U8145 ( .A(n7995), .B(n8963), .Z(n7875) );
  NAND U8146 ( .A(n7876), .B(n7875), .Z(n8051) );
  NAND U8147 ( .A(n7877), .B(n9105), .Z(n7879) );
  XNOR U8148 ( .A(n9217), .B(b[17]), .Z(n8001) );
  NAND U8149 ( .A(n8001), .B(n9107), .Z(n7878) );
  NAND U8150 ( .A(n7879), .B(n7878), .Z(n8049) );
  XNOR U8151 ( .A(a[56]), .B(b[13]), .Z(n7998) );
  NANDN U8152 ( .A(n7998), .B(n8730), .Z(n7882) );
  NAND U8153 ( .A(n7880), .B(n8731), .Z(n7881) );
  AND U8154 ( .A(n7882), .B(n7881), .Z(n8050) );
  XOR U8155 ( .A(n8049), .B(n8050), .Z(n8052) );
  XOR U8156 ( .A(n8051), .B(n8052), .Z(n8059) );
  NAND U8157 ( .A(n7884), .B(n7883), .Z(n7888) );
  NAND U8158 ( .A(n7886), .B(n7885), .Z(n7887) );
  AND U8159 ( .A(n7888), .B(n7887), .Z(n8061) );
  XNOR U8160 ( .A(n8062), .B(n8061), .Z(n8090) );
  XOR U8161 ( .A(n8089), .B(n8090), .Z(n8065) );
  XOR U8162 ( .A(b[21]), .B(n8837), .Z(n8018) );
  NANDN U8163 ( .A(n8018), .B(n9493), .Z(n7895) );
  NANDN U8164 ( .A(n7893), .B(n9495), .Z(n7894) );
  NAND U8165 ( .A(n7895), .B(n7894), .Z(n8058) );
  NAND U8166 ( .A(n7896), .B(n8286), .Z(n7898) );
  XNOR U8167 ( .A(n9805), .B(b[9]), .Z(n8035) );
  NAND U8168 ( .A(n8035), .B(n8288), .Z(n7897) );
  NAND U8169 ( .A(n7898), .B(n7897), .Z(n8055) );
  NANDN U8170 ( .A(n7899), .B(n9801), .Z(n7901) );
  XOR U8171 ( .A(b[27]), .B(n8156), .Z(n8038) );
  OR U8172 ( .A(n8038), .B(n9751), .Z(n7900) );
  AND U8173 ( .A(n7901), .B(n7900), .Z(n8056) );
  XNOR U8174 ( .A(n8055), .B(n8056), .Z(n8057) );
  XNOR U8175 ( .A(n8058), .B(n8057), .Z(n8082) );
  NAND U8176 ( .A(n7902), .B(n9914), .Z(n7904) );
  XNOR U8177 ( .A(n323), .B(a[38]), .Z(n8041) );
  NANDN U8178 ( .A(n9913), .B(n8041), .Z(n7903) );
  NAND U8179 ( .A(n7904), .B(n7903), .Z(n8028) );
  NANDN U8180 ( .A(n317), .B(n7905), .Z(n7909) );
  NANDN U8181 ( .A(n7907), .B(n7906), .Z(n7908) );
  NAND U8182 ( .A(n7909), .B(n7908), .Z(n8027) );
  ANDN U8183 ( .B(a[36]), .A(n323), .Z(n8045) );
  IV U8184 ( .A(n8045), .Z(n8207) );
  XNOR U8185 ( .A(n8027), .B(n8207), .Z(n8029) );
  XOR U8186 ( .A(n8028), .B(n8029), .Z(n8081) );
  XOR U8187 ( .A(n8082), .B(n8081), .Z(n8083) );
  XOR U8188 ( .A(n8084), .B(n8083), .Z(n7983) );
  NANDN U8189 ( .A(n7911), .B(n7910), .Z(n7915) );
  NAND U8190 ( .A(n7913), .B(n7912), .Z(n7914) );
  NAND U8191 ( .A(n7915), .B(n7914), .Z(n8077) );
  NANDN U8192 ( .A(n7916), .B(n9622), .Z(n7918) );
  XOR U8193 ( .A(b[23]), .B(n8654), .Z(n8032) );
  OR U8194 ( .A(n8032), .B(n9621), .Z(n7917) );
  NAND U8195 ( .A(n7918), .B(n7917), .Z(n7992) );
  XOR U8196 ( .A(b[25]), .B(n8444), .Z(n8004) );
  NANDN U8197 ( .A(n8004), .B(n9706), .Z(n7921) );
  NANDN U8198 ( .A(n7919), .B(n9707), .Z(n7920) );
  NAND U8199 ( .A(n7921), .B(n7920), .Z(n7989) );
  XOR U8200 ( .A(a[58]), .B(b[11]), .Z(n8007) );
  NAND U8201 ( .A(n8007), .B(n8541), .Z(n7924) );
  NAND U8202 ( .A(n7922), .B(n8542), .Z(n7923) );
  AND U8203 ( .A(n7924), .B(n7923), .Z(n7990) );
  XNOR U8204 ( .A(n7989), .B(n7990), .Z(n7991) );
  XNOR U8205 ( .A(n7992), .B(n7991), .Z(n8075) );
  XNOR U8206 ( .A(a[62]), .B(b[7]), .Z(n8015) );
  OR U8207 ( .A(n8015), .B(n8013), .Z(n7927) );
  NAND U8208 ( .A(n7925), .B(n8014), .Z(n7926) );
  NAND U8209 ( .A(n7927), .B(n7926), .Z(n8024) );
  NAND U8210 ( .A(n7928), .B(n9379), .Z(n7930) );
  XNOR U8211 ( .A(n9562), .B(a[50]), .Z(n8046) );
  NAND U8212 ( .A(n8046), .B(n9378), .Z(n7929) );
  NAND U8213 ( .A(n7930), .B(n7929), .Z(n8021) );
  NAND U8214 ( .A(n9875), .B(n7931), .Z(n7934) );
  XOR U8215 ( .A(n322), .B(n7932), .Z(n8010) );
  NANDN U8216 ( .A(n9874), .B(n8010), .Z(n7933) );
  AND U8217 ( .A(n7934), .B(n7933), .Z(n8022) );
  XNOR U8218 ( .A(n8021), .B(n8022), .Z(n8023) );
  XOR U8219 ( .A(n8024), .B(n8023), .Z(n8076) );
  XOR U8220 ( .A(n8075), .B(n8076), .Z(n8078) );
  XOR U8221 ( .A(n8077), .B(n8078), .Z(n7984) );
  XNOR U8222 ( .A(n7983), .B(n7984), .Z(n7985) );
  NANDN U8223 ( .A(n7936), .B(n7935), .Z(n7940) );
  NAND U8224 ( .A(n7938), .B(n7937), .Z(n7939) );
  NAND U8225 ( .A(n7940), .B(n7939), .Z(n7986) );
  XNOR U8226 ( .A(n7985), .B(n7986), .Z(n8066) );
  XNOR U8227 ( .A(n8065), .B(n8066), .Z(n8067) );
  XNOR U8228 ( .A(n8068), .B(n8067), .Z(n7979) );
  NAND U8229 ( .A(n7942), .B(n7941), .Z(n7946) );
  NANDN U8230 ( .A(n7944), .B(n7943), .Z(n7945) );
  NAND U8231 ( .A(n7946), .B(n7945), .Z(n8074) );
  NAND U8232 ( .A(n7948), .B(n7947), .Z(n7952) );
  OR U8233 ( .A(n7950), .B(n7949), .Z(n7951) );
  NAND U8234 ( .A(n7952), .B(n7951), .Z(n8071) );
  NANDN U8235 ( .A(n7954), .B(n7953), .Z(n7958) );
  NAND U8236 ( .A(n7956), .B(n7955), .Z(n7957) );
  AND U8237 ( .A(n7958), .B(n7957), .Z(n8072) );
  XNOR U8238 ( .A(n8071), .B(n8072), .Z(n8073) );
  XOR U8239 ( .A(n8074), .B(n8073), .Z(n7978) );
  NAND U8240 ( .A(n7960), .B(n7959), .Z(n7964) );
  NAND U8241 ( .A(n7962), .B(n7961), .Z(n7963) );
  AND U8242 ( .A(n7964), .B(n7963), .Z(n7977) );
  XNOR U8243 ( .A(n7978), .B(n7977), .Z(n7980) );
  XOR U8244 ( .A(n7979), .B(n7980), .Z(n8094) );
  XOR U8245 ( .A(n8096), .B(n8095), .Z(n7974) );
  NANDN U8246 ( .A(n7966), .B(n7965), .Z(n7970) );
  NAND U8247 ( .A(n7968), .B(n7967), .Z(n7969) );
  AND U8248 ( .A(n7970), .B(n7969), .Z(n7975) );
  XOR U8249 ( .A(n7974), .B(n7975), .Z(n7971) );
  XOR U8250 ( .A(n7976), .B(n7971), .Z(n7972) );
  XNOR U8251 ( .A(n7973), .B(n7972), .Z(c[100]) );
  NANDN U8252 ( .A(n7973), .B(n7972), .Z(n8101) );
  NANDN U8253 ( .A(n7978), .B(n7977), .Z(n7982) );
  NAND U8254 ( .A(n7980), .B(n7979), .Z(n7981) );
  NAND U8255 ( .A(n7982), .B(n7981), .Z(n8108) );
  NANDN U8256 ( .A(n7984), .B(n7983), .Z(n7988) );
  NANDN U8257 ( .A(n7986), .B(n7985), .Z(n7987) );
  NAND U8258 ( .A(n7988), .B(n7987), .Z(n8222) );
  NANDN U8259 ( .A(n7990), .B(n7989), .Z(n7994) );
  NAND U8260 ( .A(n7992), .B(n7991), .Z(n7993) );
  NAND U8261 ( .A(n7994), .B(n7993), .Z(n8122) );
  NAND U8262 ( .A(n7995), .B(n8961), .Z(n7997) );
  XOR U8263 ( .A(a[55]), .B(b[15]), .Z(n8210) );
  NAND U8264 ( .A(n8210), .B(n8963), .Z(n7996) );
  NAND U8265 ( .A(n7997), .B(n7996), .Z(n8190) );
  XOR U8266 ( .A(a[57]), .B(b[13]), .Z(n8213) );
  NAND U8267 ( .A(n8213), .B(n8730), .Z(n8000) );
  NANDN U8268 ( .A(n7998), .B(n8731), .Z(n7999) );
  NAND U8269 ( .A(n8000), .B(n7999), .Z(n8189) );
  NAND U8270 ( .A(n8001), .B(n9105), .Z(n8003) );
  XNOR U8271 ( .A(n9564), .B(b[17]), .Z(n8152) );
  NAND U8272 ( .A(n8152), .B(n9107), .Z(n8002) );
  NAND U8273 ( .A(n8003), .B(n8002), .Z(n8145) );
  XNOR U8274 ( .A(b[25]), .B(a[45]), .Z(n8216) );
  NANDN U8275 ( .A(n8216), .B(n9706), .Z(n8006) );
  NANDN U8276 ( .A(n8004), .B(n9707), .Z(n8005) );
  NAND U8277 ( .A(n8006), .B(n8005), .Z(n8143) );
  XOR U8278 ( .A(a[59]), .B(b[11]), .Z(n8171) );
  NAND U8279 ( .A(n8171), .B(n8541), .Z(n8009) );
  NAND U8280 ( .A(n8007), .B(n8542), .Z(n8008) );
  AND U8281 ( .A(n8009), .B(n8008), .Z(n8144) );
  XNOR U8282 ( .A(n8143), .B(n8144), .Z(n8146) );
  XOR U8283 ( .A(n8145), .B(n8146), .Z(n8188) );
  XOR U8284 ( .A(n8189), .B(n8188), .Z(n8191) );
  XOR U8285 ( .A(n8190), .B(n8191), .Z(n8127) );
  NAND U8286 ( .A(n9875), .B(n8010), .Z(n8012) );
  XNOR U8287 ( .A(n322), .B(a[41]), .Z(n8155) );
  NANDN U8288 ( .A(n9874), .B(n8155), .Z(n8011) );
  NAND U8289 ( .A(n8012), .B(n8011), .Z(n8197) );
  XNOR U8290 ( .A(n9946), .B(b[7]), .Z(n8179) );
  NANDN U8291 ( .A(n8013), .B(n8179), .Z(n8017) );
  NANDN U8292 ( .A(n8015), .B(n8014), .Z(n8016) );
  NAND U8293 ( .A(n8017), .B(n8016), .Z(n8194) );
  XNOR U8294 ( .A(b[21]), .B(a[49]), .Z(n8165) );
  NANDN U8295 ( .A(n8165), .B(n9493), .Z(n8020) );
  NANDN U8296 ( .A(n8018), .B(n9495), .Z(n8019) );
  AND U8297 ( .A(n8020), .B(n8019), .Z(n8195) );
  XNOR U8298 ( .A(n8194), .B(n8195), .Z(n8196) );
  XNOR U8299 ( .A(n8197), .B(n8196), .Z(n8125) );
  NANDN U8300 ( .A(n8022), .B(n8021), .Z(n8026) );
  NAND U8301 ( .A(n8024), .B(n8023), .Z(n8025) );
  NAND U8302 ( .A(n8026), .B(n8025), .Z(n8126) );
  XOR U8303 ( .A(n8125), .B(n8126), .Z(n8128) );
  XOR U8304 ( .A(n8127), .B(n8128), .Z(n8121) );
  XNOR U8305 ( .A(n8122), .B(n8121), .Z(n8123) );
  OR U8306 ( .A(n8027), .B(n8207), .Z(n8031) );
  OR U8307 ( .A(n8029), .B(n8028), .Z(n8030) );
  NAND U8308 ( .A(n8031), .B(n8030), .Z(n8134) );
  NANDN U8309 ( .A(n8032), .B(n9622), .Z(n8034) );
  XNOR U8310 ( .A(b[23]), .B(a[47]), .Z(n8162) );
  OR U8311 ( .A(n8162), .B(n9621), .Z(n8033) );
  NAND U8312 ( .A(n8034), .B(n8033), .Z(n8203) );
  NAND U8313 ( .A(n8035), .B(n8286), .Z(n8037) );
  XOR U8314 ( .A(a[61]), .B(b[9]), .Z(n8168) );
  NAND U8315 ( .A(n8168), .B(n8288), .Z(n8036) );
  NAND U8316 ( .A(n8037), .B(n8036), .Z(n8200) );
  NANDN U8317 ( .A(n8038), .B(n9801), .Z(n8040) );
  XNOR U8318 ( .A(b[27]), .B(a[43]), .Z(n8149) );
  OR U8319 ( .A(n8149), .B(n9751), .Z(n8039) );
  AND U8320 ( .A(n8040), .B(n8039), .Z(n8201) );
  XNOR U8321 ( .A(n8200), .B(n8201), .Z(n8202) );
  XNOR U8322 ( .A(n8203), .B(n8202), .Z(n8131) );
  NAND U8323 ( .A(n8041), .B(n9914), .Z(n8043) );
  XNOR U8324 ( .A(n323), .B(a[39]), .Z(n8174) );
  NANDN U8325 ( .A(n9913), .B(n8174), .Z(n8042) );
  NAND U8326 ( .A(n8043), .B(n8042), .Z(n8137) );
  NANDN U8327 ( .A(n323), .B(a[37]), .Z(n8204) );
  NANDN U8328 ( .A(n316), .B(b[4]), .Z(n8044) );
  ANDN U8329 ( .B(n8044), .A(n317), .Z(n8205) );
  XOR U8330 ( .A(n8204), .B(n8205), .Z(n8206) );
  XOR U8331 ( .A(n8045), .B(n8206), .Z(n8138) );
  XOR U8332 ( .A(n8137), .B(n8138), .Z(n8139) );
  NAND U8333 ( .A(n8046), .B(n9379), .Z(n8048) );
  XOR U8334 ( .A(b[19]), .B(n9457), .Z(n8159) );
  NANDN U8335 ( .A(n8159), .B(n9378), .Z(n8047) );
  AND U8336 ( .A(n8048), .B(n8047), .Z(n8140) );
  XNOR U8337 ( .A(n8139), .B(n8140), .Z(n8132) );
  XNOR U8338 ( .A(n8131), .B(n8132), .Z(n8133) );
  XNOR U8339 ( .A(n8134), .B(n8133), .Z(n8185) );
  NANDN U8340 ( .A(n8050), .B(n8049), .Z(n8054) );
  NANDN U8341 ( .A(n8052), .B(n8051), .Z(n8053) );
  NAND U8342 ( .A(n8054), .B(n8053), .Z(n8183) );
  XNOR U8343 ( .A(n8183), .B(n8182), .Z(n8184) );
  XOR U8344 ( .A(n8185), .B(n8184), .Z(n8124) );
  XOR U8345 ( .A(n8123), .B(n8124), .Z(n8219) );
  OR U8346 ( .A(n8060), .B(n8059), .Z(n8064) );
  OR U8347 ( .A(n8062), .B(n8061), .Z(n8063) );
  AND U8348 ( .A(n8064), .B(n8063), .Z(n8220) );
  XNOR U8349 ( .A(n8219), .B(n8220), .Z(n8221) );
  XNOR U8350 ( .A(n8222), .B(n8221), .Z(n8106) );
  NANDN U8351 ( .A(n8066), .B(n8065), .Z(n8070) );
  NAND U8352 ( .A(n8068), .B(n8067), .Z(n8069) );
  NAND U8353 ( .A(n8070), .B(n8069), .Z(n8114) );
  NANDN U8354 ( .A(n8076), .B(n8075), .Z(n8080) );
  OR U8355 ( .A(n8078), .B(n8077), .Z(n8079) );
  NAND U8356 ( .A(n8080), .B(n8079), .Z(n8115) );
  NAND U8357 ( .A(n8082), .B(n8081), .Z(n8086) );
  NANDN U8358 ( .A(n8084), .B(n8083), .Z(n8085) );
  AND U8359 ( .A(n8086), .B(n8085), .Z(n8116) );
  XNOR U8360 ( .A(n8115), .B(n8116), .Z(n8117) );
  NANDN U8361 ( .A(n8088), .B(n8087), .Z(n8092) );
  NANDN U8362 ( .A(n8090), .B(n8089), .Z(n8091) );
  AND U8363 ( .A(n8092), .B(n8091), .Z(n8118) );
  XNOR U8364 ( .A(n8117), .B(n8118), .Z(n8112) );
  XNOR U8365 ( .A(n8111), .B(n8112), .Z(n8113) );
  XOR U8366 ( .A(n8114), .B(n8113), .Z(n8105) );
  XNOR U8367 ( .A(n8106), .B(n8105), .Z(n8107) );
  XOR U8368 ( .A(n8108), .B(n8107), .Z(n8102) );
  OR U8369 ( .A(n8094), .B(n8093), .Z(n8098) );
  NANDN U8370 ( .A(n8096), .B(n8095), .Z(n8097) );
  NAND U8371 ( .A(n8098), .B(n8097), .Z(n8103) );
  XOR U8372 ( .A(n8102), .B(n8103), .Z(n8099) );
  XOR U8373 ( .A(n8104), .B(n8099), .Z(n8100) );
  XNOR U8374 ( .A(n8101), .B(n8100), .Z(c[101]) );
  NANDN U8375 ( .A(n8101), .B(n8100), .Z(n8339) );
  NAND U8376 ( .A(n8106), .B(n8105), .Z(n8110) );
  OR U8377 ( .A(n8108), .B(n8107), .Z(n8109) );
  AND U8378 ( .A(n8110), .B(n8109), .Z(n8225) );
  NANDN U8379 ( .A(n8116), .B(n8115), .Z(n8120) );
  NAND U8380 ( .A(n8118), .B(n8117), .Z(n8119) );
  NAND U8381 ( .A(n8120), .B(n8119), .Z(n8235) );
  NANDN U8382 ( .A(n8126), .B(n8125), .Z(n8130) );
  OR U8383 ( .A(n8128), .B(n8127), .Z(n8129) );
  NAND U8384 ( .A(n8130), .B(n8129), .Z(n8264) );
  NANDN U8385 ( .A(n8132), .B(n8131), .Z(n8136) );
  NAND U8386 ( .A(n8134), .B(n8133), .Z(n8135) );
  NAND U8387 ( .A(n8136), .B(n8135), .Z(n8262) );
  OR U8388 ( .A(n8138), .B(n8137), .Z(n8142) );
  NAND U8389 ( .A(n8140), .B(n8139), .Z(n8141) );
  NAND U8390 ( .A(n8142), .B(n8141), .Z(n8243) );
  NANDN U8391 ( .A(n8144), .B(n8143), .Z(n8148) );
  NAND U8392 ( .A(n8146), .B(n8145), .Z(n8147) );
  NAND U8393 ( .A(n8148), .B(n8147), .Z(n8244) );
  XNOR U8394 ( .A(n8243), .B(n8244), .Z(n8245) );
  NANDN U8395 ( .A(n8149), .B(n9801), .Z(n8151) );
  XOR U8396 ( .A(b[27]), .B(n8444), .Z(n8316) );
  OR U8397 ( .A(n8316), .B(n9751), .Z(n8150) );
  NAND U8398 ( .A(n8151), .B(n8150), .Z(n8276) );
  NAND U8399 ( .A(n8152), .B(n9105), .Z(n8154) );
  XNOR U8400 ( .A(n9353), .B(b[17]), .Z(n8310) );
  NAND U8401 ( .A(n8310), .B(n9107), .Z(n8153) );
  NAND U8402 ( .A(n8154), .B(n8153), .Z(n8273) );
  NAND U8403 ( .A(n9875), .B(n8155), .Z(n8158) );
  XOR U8404 ( .A(n322), .B(n8156), .Z(n8295) );
  NANDN U8405 ( .A(n9874), .B(n8295), .Z(n8157) );
  AND U8406 ( .A(n8158), .B(n8157), .Z(n8274) );
  XNOR U8407 ( .A(n8273), .B(n8274), .Z(n8275) );
  XNOR U8408 ( .A(n8276), .B(n8275), .Z(n8334) );
  NANDN U8409 ( .A(n8159), .B(n9379), .Z(n8161) );
  XNOR U8410 ( .A(n9217), .B(b[19]), .Z(n8307) );
  NAND U8411 ( .A(n8307), .B(n9378), .Z(n8160) );
  NAND U8412 ( .A(n8161), .B(n8160), .Z(n8332) );
  NANDN U8413 ( .A(n8162), .B(n9622), .Z(n8164) );
  XOR U8414 ( .A(b[23]), .B(n8837), .Z(n8301) );
  OR U8415 ( .A(n8301), .B(n9621), .Z(n8163) );
  AND U8416 ( .A(n8164), .B(n8163), .Z(n8331) );
  XNOR U8417 ( .A(n8332), .B(n8331), .Z(n8333) );
  XNOR U8418 ( .A(n8334), .B(n8333), .Z(n8258) );
  XOR U8419 ( .A(b[21]), .B(n9033), .Z(n8291) );
  NANDN U8420 ( .A(n8291), .B(n9493), .Z(n8167) );
  NANDN U8421 ( .A(n8165), .B(n9495), .Z(n8166) );
  NAND U8422 ( .A(n8167), .B(n8166), .Z(n8280) );
  NAND U8423 ( .A(n8168), .B(n8286), .Z(n8170) );
  XNOR U8424 ( .A(n9810), .B(b[9]), .Z(n8287) );
  NAND U8425 ( .A(n8287), .B(n8288), .Z(n8169) );
  NAND U8426 ( .A(n8170), .B(n8169), .Z(n8277) );
  XNOR U8427 ( .A(a[60]), .B(b[11]), .Z(n8319) );
  NANDN U8428 ( .A(n8319), .B(n8541), .Z(n8173) );
  NAND U8429 ( .A(n8171), .B(n8542), .Z(n8172) );
  AND U8430 ( .A(n8173), .B(n8172), .Z(n8278) );
  XNOR U8431 ( .A(n8277), .B(n8278), .Z(n8279) );
  XNOR U8432 ( .A(n8280), .B(n8279), .Z(n8256) );
  NAND U8433 ( .A(n8174), .B(n9914), .Z(n8176) );
  XNOR U8434 ( .A(n323), .B(a[40]), .Z(n8298) );
  NANDN U8435 ( .A(n9913), .B(n8298), .Z(n8175) );
  NAND U8436 ( .A(n8176), .B(n8175), .Z(n8282) );
  XNOR U8437 ( .A(b[7]), .B(n8177), .Z(n8181) );
  XOR U8438 ( .A(b[6]), .B(n317), .Z(n8178) );
  NANDN U8439 ( .A(n8179), .B(n8178), .Z(n8180) );
  AND U8440 ( .A(n8181), .B(n8180), .Z(n8281) );
  AND U8441 ( .A(a[38]), .B(b[31]), .Z(n8426) );
  XOR U8442 ( .A(n8281), .B(n8426), .Z(n8283) );
  XOR U8443 ( .A(n8282), .B(n8283), .Z(n8255) );
  XOR U8444 ( .A(n8256), .B(n8255), .Z(n8257) );
  XOR U8445 ( .A(n8258), .B(n8257), .Z(n8246) );
  XNOR U8446 ( .A(n8245), .B(n8246), .Z(n8261) );
  XOR U8447 ( .A(n8262), .B(n8261), .Z(n8263) );
  XNOR U8448 ( .A(n8264), .B(n8263), .Z(n8242) );
  NANDN U8449 ( .A(n8183), .B(n8182), .Z(n8187) );
  NANDN U8450 ( .A(n8185), .B(n8184), .Z(n8186) );
  NAND U8451 ( .A(n8187), .B(n8186), .Z(n8240) );
  NAND U8452 ( .A(n8189), .B(n8188), .Z(n8193) );
  NAND U8453 ( .A(n8191), .B(n8190), .Z(n8192) );
  NAND U8454 ( .A(n8193), .B(n8192), .Z(n8269) );
  NANDN U8455 ( .A(n8195), .B(n8194), .Z(n8199) );
  NAND U8456 ( .A(n8197), .B(n8196), .Z(n8198) );
  NAND U8457 ( .A(n8199), .B(n8198), .Z(n8268) );
  OR U8458 ( .A(n8205), .B(n8204), .Z(n8209) );
  NANDN U8459 ( .A(n8207), .B(n8206), .Z(n8208) );
  AND U8460 ( .A(n8209), .B(n8208), .Z(n8250) );
  XNOR U8461 ( .A(n8249), .B(n8250), .Z(n8251) );
  NAND U8462 ( .A(n8210), .B(n8961), .Z(n8212) );
  XNOR U8463 ( .A(n9357), .B(b[15]), .Z(n8322) );
  NAND U8464 ( .A(n8322), .B(n8963), .Z(n8211) );
  NAND U8465 ( .A(n8212), .B(n8211), .Z(n8327) );
  XOR U8466 ( .A(a[58]), .B(b[13]), .Z(n8304) );
  NAND U8467 ( .A(n8730), .B(n8304), .Z(n8215) );
  NAND U8468 ( .A(n8731), .B(n8213), .Z(n8214) );
  NAND U8469 ( .A(n8215), .B(n8214), .Z(n8325) );
  XOR U8470 ( .A(b[25]), .B(n8654), .Z(n8313) );
  NANDN U8471 ( .A(n8313), .B(n9706), .Z(n8218) );
  NANDN U8472 ( .A(n8216), .B(n9707), .Z(n8217) );
  AND U8473 ( .A(n8218), .B(n8217), .Z(n8326) );
  XOR U8474 ( .A(n8325), .B(n8326), .Z(n8328) );
  XNOR U8475 ( .A(n8327), .B(n8328), .Z(n8252) );
  XOR U8476 ( .A(n8251), .B(n8252), .Z(n8267) );
  XNOR U8477 ( .A(n8268), .B(n8267), .Z(n8270) );
  XNOR U8478 ( .A(n8269), .B(n8270), .Z(n8239) );
  XNOR U8479 ( .A(n8240), .B(n8239), .Z(n8241) );
  XOR U8480 ( .A(n8242), .B(n8241), .Z(n8233) );
  XOR U8481 ( .A(n8234), .B(n8233), .Z(n8236) );
  XNOR U8482 ( .A(n8235), .B(n8236), .Z(n8228) );
  XOR U8483 ( .A(n8228), .B(n8227), .Z(n8230) );
  XOR U8484 ( .A(n8229), .B(n8230), .Z(n8224) );
  XNOR U8485 ( .A(n8225), .B(n8224), .Z(n8223) );
  XNOR U8486 ( .A(n8226), .B(n8223), .Z(n8338) );
  XOR U8487 ( .A(n8339), .B(n8338), .Z(c[102]) );
  NAND U8488 ( .A(n8228), .B(n8227), .Z(n8232) );
  NAND U8489 ( .A(n8230), .B(n8229), .Z(n8231) );
  AND U8490 ( .A(n8232), .B(n8231), .Z(n8343) );
  NANDN U8491 ( .A(n8234), .B(n8233), .Z(n8238) );
  OR U8492 ( .A(n8236), .B(n8235), .Z(n8237) );
  NAND U8493 ( .A(n8238), .B(n8237), .Z(n8352) );
  NANDN U8494 ( .A(n8244), .B(n8243), .Z(n8248) );
  NANDN U8495 ( .A(n8246), .B(n8245), .Z(n8247) );
  NAND U8496 ( .A(n8248), .B(n8247), .Z(n8364) );
  NANDN U8497 ( .A(n8250), .B(n8249), .Z(n8254) );
  NAND U8498 ( .A(n8252), .B(n8251), .Z(n8253) );
  NAND U8499 ( .A(n8254), .B(n8253), .Z(n8361) );
  NAND U8500 ( .A(n8256), .B(n8255), .Z(n8260) );
  NANDN U8501 ( .A(n8258), .B(n8257), .Z(n8259) );
  NAND U8502 ( .A(n8260), .B(n8259), .Z(n8362) );
  XNOR U8503 ( .A(n8361), .B(n8362), .Z(n8363) );
  XOR U8504 ( .A(n8364), .B(n8363), .Z(n8355) );
  NAND U8505 ( .A(n8262), .B(n8261), .Z(n8266) );
  NAND U8506 ( .A(n8264), .B(n8263), .Z(n8265) );
  AND U8507 ( .A(n8266), .B(n8265), .Z(n8356) );
  XNOR U8508 ( .A(n8355), .B(n8356), .Z(n8357) );
  NAND U8509 ( .A(n8268), .B(n8267), .Z(n8272) );
  NANDN U8510 ( .A(n8270), .B(n8269), .Z(n8271) );
  NAND U8511 ( .A(n8272), .B(n8271), .Z(n8459) );
  XNOR U8512 ( .A(n8377), .B(n8378), .Z(n8379) );
  NANDN U8513 ( .A(n8281), .B(n8426), .Z(n8285) );
  OR U8514 ( .A(n8283), .B(n8282), .Z(n8284) );
  NAND U8515 ( .A(n8285), .B(n8284), .Z(n8374) );
  NAND U8516 ( .A(n8287), .B(n8286), .Z(n8290) );
  XNOR U8517 ( .A(n9946), .B(b[9]), .Z(n8418) );
  NAND U8518 ( .A(n8418), .B(n8288), .Z(n8289) );
  NAND U8519 ( .A(n8290), .B(n8289), .Z(n8450) );
  XOR U8520 ( .A(b[21]), .B(n9457), .Z(n8447) );
  NANDN U8521 ( .A(n8447), .B(n9493), .Z(n8293) );
  NANDN U8522 ( .A(n8291), .B(n9495), .Z(n8292) );
  AND U8523 ( .A(n8293), .B(n8292), .Z(n8451) );
  XOR U8524 ( .A(n8450), .B(n8451), .Z(n8453) );
  IV U8525 ( .A(n8294), .Z(n8424) );
  NANDN U8526 ( .A(n323), .B(a[39]), .Z(n8425) );
  XNOR U8527 ( .A(n8424), .B(n8425), .Z(n8427) );
  XOR U8528 ( .A(n8426), .B(n8427), .Z(n8452) );
  XOR U8529 ( .A(n8453), .B(n8452), .Z(n8371) );
  NAND U8530 ( .A(n9875), .B(n8295), .Z(n8297) );
  XNOR U8531 ( .A(n322), .B(a[43]), .Z(n8443) );
  NANDN U8532 ( .A(n9874), .B(n8443), .Z(n8296) );
  NAND U8533 ( .A(n8297), .B(n8296), .Z(n8433) );
  NAND U8534 ( .A(n8298), .B(n9914), .Z(n8300) );
  XNOR U8535 ( .A(n323), .B(a[41]), .Z(n8421) );
  NANDN U8536 ( .A(n9913), .B(n8421), .Z(n8299) );
  NAND U8537 ( .A(n8300), .B(n8299), .Z(n8430) );
  NANDN U8538 ( .A(n8301), .B(n9622), .Z(n8303) );
  XNOR U8539 ( .A(b[23]), .B(a[49]), .Z(n8395) );
  OR U8540 ( .A(n8395), .B(n9621), .Z(n8302) );
  AND U8541 ( .A(n8303), .B(n8302), .Z(n8431) );
  XNOR U8542 ( .A(n8430), .B(n8431), .Z(n8432) );
  XNOR U8543 ( .A(n8433), .B(n8432), .Z(n8372) );
  XNOR U8544 ( .A(n8371), .B(n8372), .Z(n8373) );
  XOR U8545 ( .A(n8374), .B(n8373), .Z(n8380) );
  XOR U8546 ( .A(n8379), .B(n8380), .Z(n8456) );
  XOR U8547 ( .A(a[59]), .B(b[13]), .Z(n8404) );
  NAND U8548 ( .A(n8404), .B(n8730), .Z(n8306) );
  NAND U8549 ( .A(n8304), .B(n8731), .Z(n8305) );
  NAND U8550 ( .A(n8306), .B(n8305), .Z(n8434) );
  NAND U8551 ( .A(n8307), .B(n9379), .Z(n8309) );
  XOR U8552 ( .A(b[19]), .B(n9564), .Z(n8401) );
  NANDN U8553 ( .A(n8401), .B(n9378), .Z(n8308) );
  AND U8554 ( .A(n8309), .B(n8308), .Z(n8435) );
  XNOR U8555 ( .A(n8434), .B(n8435), .Z(n8436) );
  XNOR U8556 ( .A(a[55]), .B(b[17]), .Z(n8407) );
  NANDN U8557 ( .A(n8407), .B(n9107), .Z(n8312) );
  NAND U8558 ( .A(n8310), .B(n9105), .Z(n8311) );
  AND U8559 ( .A(n8312), .B(n8311), .Z(n8437) );
  XOR U8560 ( .A(n8436), .B(n8437), .Z(n8370) );
  XNOR U8561 ( .A(b[25]), .B(a[47]), .Z(n8389) );
  NANDN U8562 ( .A(n8389), .B(n9706), .Z(n8315) );
  NANDN U8563 ( .A(n8313), .B(n9707), .Z(n8314) );
  NAND U8564 ( .A(n8315), .B(n8314), .Z(n8413) );
  NANDN U8565 ( .A(n8316), .B(n9801), .Z(n8318) );
  XNOR U8566 ( .A(b[27]), .B(a[45]), .Z(n8392) );
  OR U8567 ( .A(n8392), .B(n9751), .Z(n8317) );
  NAND U8568 ( .A(n8318), .B(n8317), .Z(n8410) );
  XOR U8569 ( .A(a[61]), .B(b[11]), .Z(n8440) );
  NAND U8570 ( .A(n8440), .B(n8541), .Z(n8321) );
  NANDN U8571 ( .A(n8319), .B(n8542), .Z(n8320) );
  AND U8572 ( .A(n8321), .B(n8320), .Z(n8411) );
  XNOR U8573 ( .A(n8410), .B(n8411), .Z(n8412) );
  XNOR U8574 ( .A(n8413), .B(n8412), .Z(n8367) );
  NAND U8575 ( .A(n8322), .B(n8961), .Z(n8324) );
  XOR U8576 ( .A(a[57]), .B(b[15]), .Z(n8398) );
  NAND U8577 ( .A(n8398), .B(n8963), .Z(n8323) );
  NAND U8578 ( .A(n8324), .B(n8323), .Z(n8368) );
  XNOR U8579 ( .A(n8367), .B(n8368), .Z(n8369) );
  XNOR U8580 ( .A(n8370), .B(n8369), .Z(n8383) );
  NANDN U8581 ( .A(n8326), .B(n8325), .Z(n8330) );
  NANDN U8582 ( .A(n8328), .B(n8327), .Z(n8329) );
  AND U8583 ( .A(n8330), .B(n8329), .Z(n8384) );
  XOR U8584 ( .A(n8383), .B(n8384), .Z(n8386) );
  NANDN U8585 ( .A(n8332), .B(n8331), .Z(n8336) );
  NAND U8586 ( .A(n8334), .B(n8333), .Z(n8335) );
  NAND U8587 ( .A(n8336), .B(n8335), .Z(n8385) );
  XOR U8588 ( .A(n8386), .B(n8385), .Z(n8457) );
  XNOR U8589 ( .A(n8456), .B(n8457), .Z(n8458) );
  XOR U8590 ( .A(n8459), .B(n8458), .Z(n8358) );
  XNOR U8591 ( .A(n8357), .B(n8358), .Z(n8350) );
  XNOR U8592 ( .A(n8349), .B(n8350), .Z(n8351) );
  XOR U8593 ( .A(n8352), .B(n8351), .Z(n8344) );
  IV U8594 ( .A(n8344), .Z(n8342) );
  XOR U8595 ( .A(n8343), .B(n8342), .Z(n8337) );
  XNOR U8596 ( .A(n8345), .B(n8337), .Z(n8341) );
  OR U8597 ( .A(n8339), .B(n8338), .Z(n8340) );
  XOR U8598 ( .A(n8341), .B(n8340), .Z(c[103]) );
  OR U8599 ( .A(n8341), .B(n8340), .Z(n8575) );
  NANDN U8600 ( .A(n8342), .B(n8343), .Z(n8348) );
  NOR U8601 ( .A(n8344), .B(n8343), .Z(n8346) );
  OR U8602 ( .A(n8346), .B(n8345), .Z(n8347) );
  NAND U8603 ( .A(n8348), .B(n8347), .Z(n8464) );
  NANDN U8604 ( .A(n8350), .B(n8349), .Z(n8354) );
  NAND U8605 ( .A(n8352), .B(n8351), .Z(n8353) );
  NAND U8606 ( .A(n8354), .B(n8353), .Z(n8463) );
  NANDN U8607 ( .A(n8356), .B(n8355), .Z(n8360) );
  NANDN U8608 ( .A(n8358), .B(n8357), .Z(n8359) );
  NAND U8609 ( .A(n8360), .B(n8359), .Z(n8471) );
  NANDN U8610 ( .A(n8362), .B(n8361), .Z(n8366) );
  NANDN U8611 ( .A(n8364), .B(n8363), .Z(n8365) );
  NAND U8612 ( .A(n8366), .B(n8365), .Z(n8472) );
  NANDN U8613 ( .A(n8372), .B(n8371), .Z(n8376) );
  NANDN U8614 ( .A(n8374), .B(n8373), .Z(n8375) );
  NAND U8615 ( .A(n8376), .B(n8375), .Z(n8479) );
  XNOR U8616 ( .A(n8478), .B(n8479), .Z(n8480) );
  NANDN U8617 ( .A(n8378), .B(n8377), .Z(n8382) );
  NANDN U8618 ( .A(n8380), .B(n8379), .Z(n8381) );
  NAND U8619 ( .A(n8382), .B(n8381), .Z(n8481) );
  XNOR U8620 ( .A(n8480), .B(n8481), .Z(n8473) );
  XNOR U8621 ( .A(n8472), .B(n8473), .Z(n8474) );
  NANDN U8622 ( .A(n8384), .B(n8383), .Z(n8388) );
  OR U8623 ( .A(n8386), .B(n8385), .Z(n8387) );
  NAND U8624 ( .A(n8388), .B(n8387), .Z(n8570) );
  XOR U8625 ( .A(b[25]), .B(n8837), .Z(n8496) );
  NANDN U8626 ( .A(n8496), .B(n9706), .Z(n8391) );
  NANDN U8627 ( .A(n8389), .B(n9707), .Z(n8390) );
  NAND U8628 ( .A(n8391), .B(n8390), .Z(n8514) );
  NANDN U8629 ( .A(n8392), .B(n9801), .Z(n8394) );
  XOR U8630 ( .A(b[27]), .B(n8654), .Z(n8502) );
  OR U8631 ( .A(n8502), .B(n9751), .Z(n8393) );
  NAND U8632 ( .A(n8394), .B(n8393), .Z(n8511) );
  NANDN U8633 ( .A(n8395), .B(n9622), .Z(n8397) );
  XOR U8634 ( .A(b[23]), .B(n9033), .Z(n8546) );
  OR U8635 ( .A(n8546), .B(n9621), .Z(n8396) );
  AND U8636 ( .A(n8397), .B(n8396), .Z(n8512) );
  XNOR U8637 ( .A(n8511), .B(n8512), .Z(n8513) );
  XNOR U8638 ( .A(n8514), .B(n8513), .Z(n8564) );
  NAND U8639 ( .A(n8398), .B(n8961), .Z(n8400) );
  XOR U8640 ( .A(a[58]), .B(b[15]), .Z(n8535) );
  NAND U8641 ( .A(n8535), .B(n8963), .Z(n8399) );
  NAND U8642 ( .A(n8400), .B(n8399), .Z(n8525) );
  NANDN U8643 ( .A(n8401), .B(n9379), .Z(n8403) );
  XNOR U8644 ( .A(n9353), .B(b[19]), .Z(n8499) );
  NAND U8645 ( .A(n8499), .B(n9378), .Z(n8402) );
  NAND U8646 ( .A(n8403), .B(n8402), .Z(n8523) );
  XNOR U8647 ( .A(a[60]), .B(b[13]), .Z(n8538) );
  NANDN U8648 ( .A(n8538), .B(n8730), .Z(n8406) );
  NAND U8649 ( .A(n8404), .B(n8731), .Z(n8405) );
  AND U8650 ( .A(n8406), .B(n8405), .Z(n8524) );
  XOR U8651 ( .A(n8523), .B(n8524), .Z(n8526) );
  XNOR U8652 ( .A(n8525), .B(n8526), .Z(n8561) );
  NANDN U8653 ( .A(n8407), .B(n9105), .Z(n8409) );
  XNOR U8654 ( .A(n9357), .B(b[17]), .Z(n8532) );
  NAND U8655 ( .A(n8532), .B(n9107), .Z(n8408) );
  NAND U8656 ( .A(n8409), .B(n8408), .Z(n8562) );
  XOR U8657 ( .A(n8561), .B(n8562), .Z(n8563) );
  XOR U8658 ( .A(n8564), .B(n8563), .Z(n8551) );
  NANDN U8659 ( .A(n8411), .B(n8410), .Z(n8415) );
  NAND U8660 ( .A(n8413), .B(n8412), .Z(n8414) );
  NAND U8661 ( .A(n8415), .B(n8414), .Z(n8487) );
  XNOR U8662 ( .A(b[9]), .B(n8416), .Z(n8420) );
  XNOR U8663 ( .A(b[8]), .B(b[7]), .Z(n8417) );
  NANDN U8664 ( .A(n8418), .B(n8417), .Z(n8419) );
  AND U8665 ( .A(n8420), .B(n8419), .Z(n8517) );
  AND U8666 ( .A(a[40]), .B(b[31]), .Z(n8598) );
  XOR U8667 ( .A(n8517), .B(n8598), .Z(n8519) );
  NAND U8668 ( .A(n8421), .B(n9914), .Z(n8423) );
  XNOR U8669 ( .A(n323), .B(a[42]), .Z(n8505) );
  NANDN U8670 ( .A(n9913), .B(n8505), .Z(n8422) );
  NAND U8671 ( .A(n8423), .B(n8422), .Z(n8518) );
  XNOR U8672 ( .A(n8519), .B(n8518), .Z(n8484) );
  OR U8673 ( .A(n8425), .B(n8424), .Z(n8429) );
  NANDN U8674 ( .A(n8427), .B(n8426), .Z(n8428) );
  AND U8675 ( .A(n8429), .B(n8428), .Z(n8485) );
  XNOR U8676 ( .A(n8484), .B(n8485), .Z(n8486) );
  XNOR U8677 ( .A(n8487), .B(n8486), .Z(n8549) );
  XOR U8678 ( .A(n8549), .B(n8550), .Z(n8552) );
  XOR U8679 ( .A(n8551), .B(n8552), .Z(n8567) );
  NANDN U8680 ( .A(n8435), .B(n8434), .Z(n8439) );
  NANDN U8681 ( .A(n8437), .B(n8436), .Z(n8438) );
  NAND U8682 ( .A(n8439), .B(n8438), .Z(n8557) );
  XNOR U8683 ( .A(n9810), .B(b[11]), .Z(n8543) );
  NAND U8684 ( .A(n8543), .B(n8541), .Z(n8442) );
  NAND U8685 ( .A(n8440), .B(n8542), .Z(n8441) );
  NAND U8686 ( .A(n8442), .B(n8441), .Z(n8493) );
  NAND U8687 ( .A(n9875), .B(n8443), .Z(n8446) );
  XOR U8688 ( .A(b[29]), .B(n8444), .Z(n8529) );
  OR U8689 ( .A(n8529), .B(n9874), .Z(n8445) );
  NAND U8690 ( .A(n8446), .B(n8445), .Z(n8490) );
  XOR U8691 ( .A(n318), .B(n9217), .Z(n8508) );
  NAND U8692 ( .A(n8508), .B(n9493), .Z(n8449) );
  NANDN U8693 ( .A(n8447), .B(n9495), .Z(n8448) );
  AND U8694 ( .A(n8449), .B(n8448), .Z(n8491) );
  XNOR U8695 ( .A(n8490), .B(n8491), .Z(n8492) );
  XNOR U8696 ( .A(n8493), .B(n8492), .Z(n8555) );
  NANDN U8697 ( .A(n8451), .B(n8450), .Z(n8455) );
  OR U8698 ( .A(n8453), .B(n8452), .Z(n8454) );
  NAND U8699 ( .A(n8455), .B(n8454), .Z(n8556) );
  XOR U8700 ( .A(n8555), .B(n8556), .Z(n8558) );
  XOR U8701 ( .A(n8557), .B(n8558), .Z(n8568) );
  XNOR U8702 ( .A(n8567), .B(n8568), .Z(n8569) );
  XOR U8703 ( .A(n8570), .B(n8569), .Z(n8475) );
  XNOR U8704 ( .A(n8474), .B(n8475), .Z(n8468) );
  NANDN U8705 ( .A(n8457), .B(n8456), .Z(n8461) );
  NANDN U8706 ( .A(n8459), .B(n8458), .Z(n8460) );
  AND U8707 ( .A(n8461), .B(n8460), .Z(n8469) );
  XNOR U8708 ( .A(n8468), .B(n8469), .Z(n8470) );
  XOR U8709 ( .A(n8471), .B(n8470), .Z(n8462) );
  XOR U8710 ( .A(n8463), .B(n8462), .Z(n8465) );
  XOR U8711 ( .A(n8464), .B(n8465), .Z(n8574) );
  XOR U8712 ( .A(n8575), .B(n8574), .Z(c[104]) );
  NANDN U8713 ( .A(n8463), .B(n8462), .Z(n8467) );
  OR U8714 ( .A(n8465), .B(n8464), .Z(n8466) );
  AND U8715 ( .A(n8467), .B(n8466), .Z(n8580) );
  NANDN U8716 ( .A(n8473), .B(n8472), .Z(n8477) );
  NAND U8717 ( .A(n8475), .B(n8474), .Z(n8476) );
  NAND U8718 ( .A(n8477), .B(n8476), .Z(n8678) );
  NANDN U8719 ( .A(n8479), .B(n8478), .Z(n8483) );
  NANDN U8720 ( .A(n8481), .B(n8480), .Z(n8482) );
  NAND U8721 ( .A(n8483), .B(n8482), .Z(n8671) );
  NANDN U8722 ( .A(n8485), .B(n8484), .Z(n8489) );
  NAND U8723 ( .A(n8487), .B(n8486), .Z(n8488) );
  NAND U8724 ( .A(n8489), .B(n8488), .Z(n8589) );
  NANDN U8725 ( .A(n8491), .B(n8490), .Z(n8495) );
  NAND U8726 ( .A(n8493), .B(n8492), .Z(n8494) );
  NAND U8727 ( .A(n8495), .B(n8494), .Z(n8620) );
  XNOR U8728 ( .A(b[25]), .B(a[49]), .Z(n8630) );
  NANDN U8729 ( .A(n8630), .B(n9706), .Z(n8498) );
  NANDN U8730 ( .A(n8496), .B(n9707), .Z(n8497) );
  NAND U8731 ( .A(n8498), .B(n8497), .Z(n8669) );
  NAND U8732 ( .A(n8499), .B(n9379), .Z(n8501) );
  XNOR U8733 ( .A(a[55]), .B(n9562), .Z(n8633) );
  NAND U8734 ( .A(n8633), .B(n9378), .Z(n8500) );
  NAND U8735 ( .A(n8501), .B(n8500), .Z(n8666) );
  NANDN U8736 ( .A(n8502), .B(n9801), .Z(n8504) );
  XNOR U8737 ( .A(b[27]), .B(a[47]), .Z(n8647) );
  OR U8738 ( .A(n8647), .B(n9751), .Z(n8503) );
  AND U8739 ( .A(n8504), .B(n8503), .Z(n8667) );
  XNOR U8740 ( .A(n8666), .B(n8667), .Z(n8668) );
  XNOR U8741 ( .A(n8669), .B(n8668), .Z(n8618) );
  NANDN U8742 ( .A(n323), .B(a[41]), .Z(n8597) );
  XOR U8743 ( .A(n8596), .B(n8597), .Z(n8599) );
  XNOR U8744 ( .A(n8598), .B(n8599), .Z(n8624) );
  NAND U8745 ( .A(n8505), .B(n9914), .Z(n8507) );
  XNOR U8746 ( .A(n323), .B(a[43]), .Z(n8639) );
  NANDN U8747 ( .A(n9913), .B(n8639), .Z(n8506) );
  NAND U8748 ( .A(n8507), .B(n8506), .Z(n8625) );
  XOR U8749 ( .A(n8624), .B(n8625), .Z(n8626) );
  XOR U8750 ( .A(b[21]), .B(n9564), .Z(n8636) );
  NANDN U8751 ( .A(n8636), .B(n9493), .Z(n8510) );
  NAND U8752 ( .A(n9495), .B(n8508), .Z(n8509) );
  AND U8753 ( .A(n8510), .B(n8509), .Z(n8627) );
  XNOR U8754 ( .A(n8626), .B(n8627), .Z(n8619) );
  XOR U8755 ( .A(n8618), .B(n8619), .Z(n8621) );
  XOR U8756 ( .A(n8620), .B(n8621), .Z(n8595) );
  NANDN U8757 ( .A(n8512), .B(n8511), .Z(n8516) );
  NAND U8758 ( .A(n8514), .B(n8513), .Z(n8515) );
  AND U8759 ( .A(n8516), .B(n8515), .Z(n8594) );
  NANDN U8760 ( .A(n8517), .B(n8598), .Z(n8521) );
  OR U8761 ( .A(n8519), .B(n8518), .Z(n8520) );
  AND U8762 ( .A(n8521), .B(n8520), .Z(n8593) );
  XNOR U8763 ( .A(n8594), .B(n8593), .Z(n8522) );
  XNOR U8764 ( .A(n8595), .B(n8522), .Z(n8588) );
  NANDN U8765 ( .A(n8524), .B(n8523), .Z(n8528) );
  NANDN U8766 ( .A(n8526), .B(n8525), .Z(n8527) );
  NAND U8767 ( .A(n8528), .B(n8527), .Z(n8614) );
  NANDN U8768 ( .A(n8529), .B(n9875), .Z(n8531) );
  XNOR U8769 ( .A(n322), .B(a[45]), .Z(n8653) );
  NANDN U8770 ( .A(n9874), .B(n8653), .Z(n8530) );
  NAND U8771 ( .A(n8531), .B(n8530), .Z(n8608) );
  NAND U8772 ( .A(n8532), .B(n9105), .Z(n8534) );
  XNOR U8773 ( .A(a[57]), .B(n9455), .Z(n8650) );
  NAND U8774 ( .A(n8650), .B(n9107), .Z(n8533) );
  NAND U8775 ( .A(n8534), .B(n8533), .Z(n8606) );
  NAND U8776 ( .A(n8535), .B(n8961), .Z(n8537) );
  XOR U8777 ( .A(a[59]), .B(b[15]), .Z(n8663) );
  NAND U8778 ( .A(n8663), .B(n8963), .Z(n8536) );
  NAND U8779 ( .A(n8537), .B(n8536), .Z(n8607) );
  XOR U8780 ( .A(n8606), .B(n8607), .Z(n8609) );
  XNOR U8781 ( .A(n8608), .B(n8609), .Z(n8612) );
  XOR U8782 ( .A(a[61]), .B(b[13]), .Z(n8660) );
  NAND U8783 ( .A(n8660), .B(n8730), .Z(n8540) );
  NANDN U8784 ( .A(n8538), .B(n8731), .Z(n8539) );
  NAND U8785 ( .A(n8540), .B(n8539), .Z(n8603) );
  XNOR U8786 ( .A(n9946), .B(b[11]), .Z(n8644) );
  NAND U8787 ( .A(n8644), .B(n8541), .Z(n8545) );
  NAND U8788 ( .A(n8543), .B(n8542), .Z(n8544) );
  NAND U8789 ( .A(n8545), .B(n8544), .Z(n8600) );
  NANDN U8790 ( .A(n8546), .B(n9622), .Z(n8548) );
  XOR U8791 ( .A(b[23]), .B(n9457), .Z(n8657) );
  OR U8792 ( .A(n8657), .B(n9621), .Z(n8547) );
  AND U8793 ( .A(n8548), .B(n8547), .Z(n8601) );
  XNOR U8794 ( .A(n8600), .B(n8601), .Z(n8602) );
  XOR U8795 ( .A(n8603), .B(n8602), .Z(n8613) );
  XOR U8796 ( .A(n8612), .B(n8613), .Z(n8615) );
  XOR U8797 ( .A(n8614), .B(n8615), .Z(n8587) );
  XOR U8798 ( .A(n8588), .B(n8587), .Z(n8590) );
  XOR U8799 ( .A(n8589), .B(n8590), .Z(n8670) );
  XNOR U8800 ( .A(n8671), .B(n8670), .Z(n8673) );
  NANDN U8801 ( .A(n8550), .B(n8549), .Z(n8554) );
  NANDN U8802 ( .A(n8552), .B(n8551), .Z(n8553) );
  NAND U8803 ( .A(n8554), .B(n8553), .Z(n8584) );
  NANDN U8804 ( .A(n8556), .B(n8555), .Z(n8560) );
  OR U8805 ( .A(n8558), .B(n8557), .Z(n8559) );
  NAND U8806 ( .A(n8560), .B(n8559), .Z(n8581) );
  OR U8807 ( .A(n8562), .B(n8561), .Z(n8566) );
  NAND U8808 ( .A(n8564), .B(n8563), .Z(n8565) );
  AND U8809 ( .A(n8566), .B(n8565), .Z(n8582) );
  XNOR U8810 ( .A(n8581), .B(n8582), .Z(n8583) );
  XOR U8811 ( .A(n8584), .B(n8583), .Z(n8672) );
  XOR U8812 ( .A(n8673), .B(n8672), .Z(n8677) );
  NANDN U8813 ( .A(n8568), .B(n8567), .Z(n8572) );
  NAND U8814 ( .A(n8570), .B(n8569), .Z(n8571) );
  NAND U8815 ( .A(n8572), .B(n8571), .Z(n8676) );
  XOR U8816 ( .A(n8677), .B(n8676), .Z(n8679) );
  XOR U8817 ( .A(n8678), .B(n8679), .Z(n8578) );
  XOR U8818 ( .A(n8579), .B(n8578), .Z(n8573) );
  XOR U8819 ( .A(n8580), .B(n8573), .Z(n8576) );
  OR U8820 ( .A(n8575), .B(n8574), .Z(n8577) );
  XNOR U8821 ( .A(n8576), .B(n8577), .Z(c[105]) );
  NANDN U8822 ( .A(n8577), .B(n8576), .Z(n8684) );
  NANDN U8823 ( .A(n8582), .B(n8581), .Z(n8586) );
  NAND U8824 ( .A(n8584), .B(n8583), .Z(n8585) );
  NAND U8825 ( .A(n8586), .B(n8585), .Z(n8775) );
  NANDN U8826 ( .A(n8588), .B(n8587), .Z(n8592) );
  OR U8827 ( .A(n8590), .B(n8589), .Z(n8591) );
  NAND U8828 ( .A(n8592), .B(n8591), .Z(n8691) );
  NANDN U8829 ( .A(n8601), .B(n8600), .Z(n8605) );
  NAND U8830 ( .A(n8603), .B(n8602), .Z(n8604) );
  NAND U8831 ( .A(n8605), .B(n8604), .Z(n8705) );
  NAND U8832 ( .A(n8607), .B(n8606), .Z(n8611) );
  NAND U8833 ( .A(n8609), .B(n8608), .Z(n8610) );
  AND U8834 ( .A(n8611), .B(n8610), .Z(n8704) );
  XNOR U8835 ( .A(n8705), .B(n8704), .Z(n8706) );
  XOR U8836 ( .A(n8707), .B(n8706), .Z(n8694) );
  NANDN U8837 ( .A(n8613), .B(n8612), .Z(n8617) );
  OR U8838 ( .A(n8615), .B(n8614), .Z(n8616) );
  NAND U8839 ( .A(n8617), .B(n8616), .Z(n8695) );
  XNOR U8840 ( .A(n8694), .B(n8695), .Z(n8696) );
  NANDN U8841 ( .A(n8619), .B(n8618), .Z(n8623) );
  OR U8842 ( .A(n8621), .B(n8620), .Z(n8622) );
  NAND U8843 ( .A(n8623), .B(n8622), .Z(n8703) );
  OR U8844 ( .A(n8625), .B(n8624), .Z(n8629) );
  NAND U8845 ( .A(n8627), .B(n8626), .Z(n8628) );
  NAND U8846 ( .A(n8629), .B(n8628), .Z(n8769) );
  XOR U8847 ( .A(b[25]), .B(n9033), .Z(n8744) );
  NANDN U8848 ( .A(n8744), .B(n9706), .Z(n8632) );
  NANDN U8849 ( .A(n8630), .B(n9707), .Z(n8631) );
  NAND U8850 ( .A(n8632), .B(n8631), .Z(n8756) );
  NAND U8851 ( .A(n8633), .B(n9379), .Z(n8635) );
  XNOR U8852 ( .A(n9357), .B(b[19]), .Z(n8747) );
  NAND U8853 ( .A(n8747), .B(n9378), .Z(n8634) );
  NAND U8854 ( .A(n8635), .B(n8634), .Z(n8753) );
  XOR U8855 ( .A(b[21]), .B(n9353), .Z(n8735) );
  NANDN U8856 ( .A(n8735), .B(n9493), .Z(n8638) );
  NANDN U8857 ( .A(n8636), .B(n9495), .Z(n8637) );
  AND U8858 ( .A(n8638), .B(n8637), .Z(n8754) );
  XNOR U8859 ( .A(n8753), .B(n8754), .Z(n8755) );
  XOR U8860 ( .A(n8756), .B(n8755), .Z(n8770) );
  XNOR U8861 ( .A(n8769), .B(n8770), .Z(n8771) );
  NAND U8862 ( .A(n8639), .B(n9914), .Z(n8641) );
  XNOR U8863 ( .A(n323), .B(a[44]), .Z(n8724) );
  NANDN U8864 ( .A(n9913), .B(n8724), .Z(n8640) );
  NAND U8865 ( .A(n8641), .B(n8640), .Z(n8717) );
  XNOR U8866 ( .A(b[11]), .B(n8642), .Z(n8646) );
  XNOR U8867 ( .A(b[10]), .B(b[9]), .Z(n8643) );
  NANDN U8868 ( .A(n8644), .B(n8643), .Z(n8645) );
  AND U8869 ( .A(n8646), .B(n8645), .Z(n8716) );
  AND U8870 ( .A(a[42]), .B(b[31]), .Z(n8854) );
  XOR U8871 ( .A(n8716), .B(n8854), .Z(n8718) );
  XOR U8872 ( .A(n8717), .B(n8718), .Z(n8772) );
  XNOR U8873 ( .A(n8771), .B(n8772), .Z(n8700) );
  NANDN U8874 ( .A(n8647), .B(n9801), .Z(n8649) );
  XOR U8875 ( .A(b[27]), .B(n8837), .Z(n8750) );
  OR U8876 ( .A(n8750), .B(n9751), .Z(n8648) );
  NAND U8877 ( .A(n8649), .B(n8648), .Z(n8762) );
  NAND U8878 ( .A(n8650), .B(n9105), .Z(n8652) );
  XNOR U8879 ( .A(a[58]), .B(n9455), .Z(n8738) );
  NAND U8880 ( .A(n8738), .B(n9107), .Z(n8651) );
  NAND U8881 ( .A(n8652), .B(n8651), .Z(n8759) );
  NAND U8882 ( .A(n9875), .B(n8653), .Z(n8656) );
  XOR U8883 ( .A(n322), .B(n8654), .Z(n8727) );
  NANDN U8884 ( .A(n9874), .B(n8727), .Z(n8655) );
  AND U8885 ( .A(n8656), .B(n8655), .Z(n8760) );
  XNOR U8886 ( .A(n8759), .B(n8760), .Z(n8761) );
  XNOR U8887 ( .A(n8762), .B(n8761), .Z(n8763) );
  NANDN U8888 ( .A(n8657), .B(n9622), .Z(n8659) );
  XOR U8889 ( .A(b[23]), .B(n9217), .Z(n8721) );
  OR U8890 ( .A(n8721), .B(n9621), .Z(n8658) );
  NAND U8891 ( .A(n8659), .B(n8658), .Z(n8713) );
  XNOR U8892 ( .A(a[62]), .B(b[13]), .Z(n8732) );
  NANDN U8893 ( .A(n8732), .B(n8730), .Z(n8662) );
  NAND U8894 ( .A(n8660), .B(n8731), .Z(n8661) );
  NAND U8895 ( .A(n8662), .B(n8661), .Z(n8710) );
  XNOR U8896 ( .A(a[60]), .B(b[15]), .Z(n8741) );
  NANDN U8897 ( .A(n8741), .B(n8963), .Z(n8665) );
  NAND U8898 ( .A(n8663), .B(n8961), .Z(n8664) );
  AND U8899 ( .A(n8665), .B(n8664), .Z(n8711) );
  XNOR U8900 ( .A(n8710), .B(n8711), .Z(n8712) );
  XOR U8901 ( .A(n8713), .B(n8712), .Z(n8764) );
  XOR U8902 ( .A(n8763), .B(n8764), .Z(n8766) );
  XOR U8903 ( .A(n8766), .B(n8765), .Z(n8701) );
  XNOR U8904 ( .A(n8700), .B(n8701), .Z(n8702) );
  XOR U8905 ( .A(n8703), .B(n8702), .Z(n8697) );
  XNOR U8906 ( .A(n8696), .B(n8697), .Z(n8689) );
  XOR U8907 ( .A(n8688), .B(n8689), .Z(n8690) );
  XOR U8908 ( .A(n8691), .B(n8690), .Z(n8776) );
  XOR U8909 ( .A(n8775), .B(n8776), .Z(n8777) );
  NAND U8910 ( .A(n8671), .B(n8670), .Z(n8675) );
  NANDN U8911 ( .A(n8673), .B(n8672), .Z(n8674) );
  AND U8912 ( .A(n8675), .B(n8674), .Z(n8778) );
  XNOR U8913 ( .A(n8777), .B(n8778), .Z(n8685) );
  NAND U8914 ( .A(n8677), .B(n8676), .Z(n8681) );
  NAND U8915 ( .A(n8679), .B(n8678), .Z(n8680) );
  AND U8916 ( .A(n8681), .B(n8680), .Z(n8686) );
  XOR U8917 ( .A(n8685), .B(n8686), .Z(n8682) );
  XNOR U8918 ( .A(n8687), .B(n8682), .Z(n8683) );
  XOR U8919 ( .A(n8684), .B(n8683), .Z(c[106]) );
  OR U8920 ( .A(n8684), .B(n8683), .Z(n8782) );
  NAND U8921 ( .A(n8689), .B(n8688), .Z(n8693) );
  NANDN U8922 ( .A(n8691), .B(n8690), .Z(n8692) );
  NAND U8923 ( .A(n8693), .B(n8692), .Z(n8885) );
  NANDN U8924 ( .A(n8695), .B(n8694), .Z(n8699) );
  NANDN U8925 ( .A(n8697), .B(n8696), .Z(n8698) );
  NAND U8926 ( .A(n8699), .B(n8698), .Z(n8883) );
  NANDN U8927 ( .A(n8705), .B(n8704), .Z(n8709) );
  NANDN U8928 ( .A(n8707), .B(n8706), .Z(n8708) );
  NAND U8929 ( .A(n8709), .B(n8708), .Z(n8877) );
  XNOR U8930 ( .A(n8876), .B(n8877), .Z(n8878) );
  NANDN U8931 ( .A(n8711), .B(n8710), .Z(n8715) );
  NAND U8932 ( .A(n8713), .B(n8712), .Z(n8714) );
  AND U8933 ( .A(n8715), .B(n8714), .Z(n8859) );
  NANDN U8934 ( .A(n8716), .B(n8854), .Z(n8720) );
  OR U8935 ( .A(n8718), .B(n8717), .Z(n8719) );
  NAND U8936 ( .A(n8720), .B(n8719), .Z(n8811) );
  NANDN U8937 ( .A(n8721), .B(n9622), .Z(n8723) );
  XOR U8938 ( .A(b[23]), .B(n9564), .Z(n8840) );
  OR U8939 ( .A(n8840), .B(n9621), .Z(n8722) );
  NAND U8940 ( .A(n8723), .B(n8722), .Z(n8792) );
  NAND U8941 ( .A(n8724), .B(n9914), .Z(n8726) );
  XNOR U8942 ( .A(n323), .B(a[45]), .Z(n8800) );
  NANDN U8943 ( .A(n9913), .B(n8800), .Z(n8725) );
  NAND U8944 ( .A(n8726), .B(n8725), .Z(n8789) );
  NANDN U8945 ( .A(n323), .B(a[43]), .Z(n8853) );
  XOR U8946 ( .A(n8852), .B(n8853), .Z(n8855) );
  XOR U8947 ( .A(n8854), .B(n8855), .Z(n8790) );
  XNOR U8948 ( .A(n8789), .B(n8790), .Z(n8791) );
  XNOR U8949 ( .A(n8792), .B(n8791), .Z(n8810) );
  NAND U8950 ( .A(n9875), .B(n8727), .Z(n8729) );
  XNOR U8951 ( .A(b[29]), .B(a[47]), .Z(n8836) );
  OR U8952 ( .A(n8836), .B(n9874), .Z(n8728) );
  NAND U8953 ( .A(n8729), .B(n8728), .Z(n8824) );
  XNOR U8954 ( .A(n9946), .B(b[13]), .Z(n8797) );
  NAND U8955 ( .A(n8797), .B(n8730), .Z(n8734) );
  NANDN U8956 ( .A(n8732), .B(n8731), .Z(n8733) );
  NAND U8957 ( .A(n8734), .B(n8733), .Z(n8821) );
  XNOR U8958 ( .A(b[21]), .B(a[55]), .Z(n8830) );
  NANDN U8959 ( .A(n8830), .B(n9493), .Z(n8737) );
  NANDN U8960 ( .A(n8735), .B(n9495), .Z(n8736) );
  AND U8961 ( .A(n8737), .B(n8736), .Z(n8822) );
  XNOR U8962 ( .A(n8821), .B(n8822), .Z(n8823) );
  XOR U8963 ( .A(n8824), .B(n8823), .Z(n8809) );
  XOR U8964 ( .A(n8810), .B(n8809), .Z(n8812) );
  XOR U8965 ( .A(n8811), .B(n8812), .Z(n8858) );
  XNOR U8966 ( .A(n8859), .B(n8858), .Z(n8861) );
  NAND U8967 ( .A(n8738), .B(n9105), .Z(n8740) );
  XNOR U8968 ( .A(a[59]), .B(n9455), .Z(n8843) );
  NAND U8969 ( .A(n8843), .B(n9107), .Z(n8739) );
  NAND U8970 ( .A(n8740), .B(n8739), .Z(n8817) );
  NANDN U8971 ( .A(n8741), .B(n8961), .Z(n8743) );
  XOR U8972 ( .A(a[61]), .B(b[15]), .Z(n8849) );
  NAND U8973 ( .A(n8849), .B(n8963), .Z(n8742) );
  NAND U8974 ( .A(n8743), .B(n8742), .Z(n8815) );
  XOR U8975 ( .A(b[25]), .B(n9457), .Z(n8846) );
  NANDN U8976 ( .A(n8846), .B(n9706), .Z(n8746) );
  NANDN U8977 ( .A(n8744), .B(n9707), .Z(n8745) );
  NAND U8978 ( .A(n8746), .B(n8745), .Z(n8805) );
  NAND U8979 ( .A(n8747), .B(n9379), .Z(n8749) );
  XNOR U8980 ( .A(a[57]), .B(n9562), .Z(n8827) );
  NAND U8981 ( .A(n8827), .B(n9378), .Z(n8748) );
  NAND U8982 ( .A(n8749), .B(n8748), .Z(n8803) );
  NANDN U8983 ( .A(n8750), .B(n9801), .Z(n8752) );
  XNOR U8984 ( .A(n321), .B(a[49]), .Z(n8833) );
  NANDN U8985 ( .A(n9751), .B(n8833), .Z(n8751) );
  AND U8986 ( .A(n8752), .B(n8751), .Z(n8804) );
  XOR U8987 ( .A(n8803), .B(n8804), .Z(n8806) );
  XOR U8988 ( .A(n8805), .B(n8806), .Z(n8816) );
  XOR U8989 ( .A(n8815), .B(n8816), .Z(n8818) );
  XNOR U8990 ( .A(n8817), .B(n8818), .Z(n8860) );
  XOR U8991 ( .A(n8861), .B(n8860), .Z(n8864) );
  NANDN U8992 ( .A(n8754), .B(n8753), .Z(n8758) );
  NAND U8993 ( .A(n8756), .B(n8755), .Z(n8757) );
  NAND U8994 ( .A(n8758), .B(n8757), .Z(n8865) );
  XOR U8995 ( .A(n8864), .B(n8865), .Z(n8866) );
  XOR U8996 ( .A(n8866), .B(n8867), .Z(n8873) );
  NANDN U8997 ( .A(n8764), .B(n8763), .Z(n8768) );
  OR U8998 ( .A(n8766), .B(n8765), .Z(n8767) );
  NAND U8999 ( .A(n8768), .B(n8767), .Z(n8871) );
  NANDN U9000 ( .A(n8770), .B(n8769), .Z(n8774) );
  NAND U9001 ( .A(n8772), .B(n8771), .Z(n8773) );
  AND U9002 ( .A(n8774), .B(n8773), .Z(n8870) );
  XNOR U9003 ( .A(n8871), .B(n8870), .Z(n8872) );
  XOR U9004 ( .A(n8873), .B(n8872), .Z(n8879) );
  XOR U9005 ( .A(n8878), .B(n8879), .Z(n8882) );
  XOR U9006 ( .A(n8883), .B(n8882), .Z(n8884) );
  XNOR U9007 ( .A(n8885), .B(n8884), .Z(n8783) );
  OR U9008 ( .A(n8776), .B(n8775), .Z(n8780) );
  NAND U9009 ( .A(n8778), .B(n8777), .Z(n8779) );
  NAND U9010 ( .A(n8780), .B(n8779), .Z(n8784) );
  XOR U9011 ( .A(n8783), .B(n8784), .Z(n8786) );
  XNOR U9012 ( .A(n8785), .B(n8786), .Z(n8781) );
  XOR U9013 ( .A(n8782), .B(n8781), .Z(c[107]) );
  OR U9014 ( .A(n8782), .B(n8781), .Z(n8981) );
  NANDN U9015 ( .A(n8784), .B(n8783), .Z(n8788) );
  NANDN U9016 ( .A(n8786), .B(n8785), .Z(n8787) );
  NAND U9017 ( .A(n8788), .B(n8787), .Z(n8891) );
  NANDN U9018 ( .A(n8790), .B(n8789), .Z(n8794) );
  NAND U9019 ( .A(n8792), .B(n8791), .Z(n8793) );
  NAND U9020 ( .A(n8794), .B(n8793), .Z(n8909) );
  XNOR U9021 ( .A(b[13]), .B(n8795), .Z(n8799) );
  XNOR U9022 ( .A(b[12]), .B(b[11]), .Z(n8796) );
  NANDN U9023 ( .A(n8797), .B(n8796), .Z(n8798) );
  AND U9024 ( .A(n8799), .B(n8798), .Z(n8956) );
  NAND U9025 ( .A(n8800), .B(n9914), .Z(n8802) );
  XNOR U9026 ( .A(n323), .B(a[46]), .Z(n8930) );
  NANDN U9027 ( .A(n9913), .B(n8930), .Z(n8801) );
  NAND U9028 ( .A(n8802), .B(n8801), .Z(n8955) );
  AND U9029 ( .A(b[31]), .B(a[44]), .Z(n9011) );
  XOR U9030 ( .A(n8955), .B(n9011), .Z(n8957) );
  XNOR U9031 ( .A(n8956), .B(n8957), .Z(n8906) );
  NANDN U9032 ( .A(n8804), .B(n8803), .Z(n8808) );
  NANDN U9033 ( .A(n8806), .B(n8805), .Z(n8807) );
  NAND U9034 ( .A(n8808), .B(n8807), .Z(n8907) );
  XOR U9035 ( .A(n8906), .B(n8907), .Z(n8908) );
  XNOR U9036 ( .A(n8909), .B(n8908), .Z(n8973) );
  NANDN U9037 ( .A(n8810), .B(n8809), .Z(n8814) );
  OR U9038 ( .A(n8812), .B(n8811), .Z(n8813) );
  AND U9039 ( .A(n8814), .B(n8813), .Z(n8974) );
  XNOR U9040 ( .A(n8973), .B(n8974), .Z(n8975) );
  NANDN U9041 ( .A(n8816), .B(n8815), .Z(n8820) );
  NANDN U9042 ( .A(n8818), .B(n8817), .Z(n8819) );
  NAND U9043 ( .A(n8820), .B(n8819), .Z(n8915) );
  NANDN U9044 ( .A(n8822), .B(n8821), .Z(n8826) );
  NAND U9045 ( .A(n8824), .B(n8823), .Z(n8825) );
  NAND U9046 ( .A(n8826), .B(n8825), .Z(n8912) );
  NAND U9047 ( .A(n8827), .B(n9379), .Z(n8829) );
  XNOR U9048 ( .A(a[58]), .B(n9562), .Z(n8939) );
  NAND U9049 ( .A(n8939), .B(n9378), .Z(n8828) );
  NAND U9050 ( .A(n8829), .B(n8828), .Z(n8947) );
  XOR U9051 ( .A(n9357), .B(n318), .Z(n8942) );
  NAND U9052 ( .A(n8942), .B(n9493), .Z(n8832) );
  NANDN U9053 ( .A(n8830), .B(n9495), .Z(n8831) );
  NAND U9054 ( .A(n8832), .B(n8831), .Z(n8946) );
  XOR U9055 ( .A(n321), .B(a[50]), .Z(n8933) );
  OR U9056 ( .A(n8933), .B(n9751), .Z(n8835) );
  NAND U9057 ( .A(n9801), .B(n8833), .Z(n8834) );
  NAND U9058 ( .A(n8835), .B(n8834), .Z(n8971) );
  NANDN U9059 ( .A(n8836), .B(n9875), .Z(n8839) );
  XOR U9060 ( .A(b[29]), .B(n8837), .Z(n8936) );
  OR U9061 ( .A(n8936), .B(n9874), .Z(n8838) );
  NAND U9062 ( .A(n8839), .B(n8838), .Z(n8969) );
  NANDN U9063 ( .A(n8840), .B(n9622), .Z(n8842) );
  XOR U9064 ( .A(n319), .B(n9353), .Z(n8924) );
  NANDN U9065 ( .A(n9621), .B(n8924), .Z(n8841) );
  AND U9066 ( .A(n8842), .B(n8841), .Z(n8970) );
  XNOR U9067 ( .A(n8969), .B(n8970), .Z(n8972) );
  XOR U9068 ( .A(n8971), .B(n8972), .Z(n8945) );
  XNOR U9069 ( .A(n8946), .B(n8945), .Z(n8948) );
  XNOR U9070 ( .A(n8947), .B(n8948), .Z(n8952) );
  NAND U9071 ( .A(n8843), .B(n9105), .Z(n8845) );
  XNOR U9072 ( .A(n9805), .B(b[17]), .Z(n8927) );
  NAND U9073 ( .A(n8927), .B(n9107), .Z(n8844) );
  NAND U9074 ( .A(n8845), .B(n8844), .Z(n8920) );
  XOR U9075 ( .A(n320), .B(n9217), .Z(n8966) );
  NAND U9076 ( .A(n8966), .B(n9706), .Z(n8848) );
  NANDN U9077 ( .A(n8846), .B(n9707), .Z(n8847) );
  NAND U9078 ( .A(n8848), .B(n8847), .Z(n8918) );
  XNOR U9079 ( .A(a[62]), .B(b[15]), .Z(n8962) );
  NANDN U9080 ( .A(n8962), .B(n8963), .Z(n8851) );
  NAND U9081 ( .A(n8849), .B(n8961), .Z(n8850) );
  AND U9082 ( .A(n8851), .B(n8850), .Z(n8919) );
  XNOR U9083 ( .A(n8918), .B(n8919), .Z(n8921) );
  XOR U9084 ( .A(n8920), .B(n8921), .Z(n8949) );
  NANDN U9085 ( .A(n8853), .B(n8852), .Z(n8857) );
  NANDN U9086 ( .A(n8855), .B(n8854), .Z(n8856) );
  NAND U9087 ( .A(n8857), .B(n8856), .Z(n8950) );
  XOR U9088 ( .A(n8949), .B(n8950), .Z(n8951) );
  XOR U9089 ( .A(n8952), .B(n8951), .Z(n8913) );
  XOR U9090 ( .A(n8912), .B(n8913), .Z(n8914) );
  XOR U9091 ( .A(n8915), .B(n8914), .Z(n8976) );
  XNOR U9092 ( .A(n8975), .B(n8976), .Z(n8903) );
  NANDN U9093 ( .A(n8859), .B(n8858), .Z(n8863) );
  NAND U9094 ( .A(n8861), .B(n8860), .Z(n8862) );
  NAND U9095 ( .A(n8863), .B(n8862), .Z(n8900) );
  OR U9096 ( .A(n8865), .B(n8864), .Z(n8869) );
  NANDN U9097 ( .A(n8867), .B(n8866), .Z(n8868) );
  NAND U9098 ( .A(n8869), .B(n8868), .Z(n8901) );
  XNOR U9099 ( .A(n8900), .B(n8901), .Z(n8902) );
  XNOR U9100 ( .A(n8903), .B(n8902), .Z(n8894) );
  NANDN U9101 ( .A(n8871), .B(n8870), .Z(n8875) );
  NAND U9102 ( .A(n8873), .B(n8872), .Z(n8874) );
  NAND U9103 ( .A(n8875), .B(n8874), .Z(n8895) );
  XNOR U9104 ( .A(n8894), .B(n8895), .Z(n8896) );
  NANDN U9105 ( .A(n8877), .B(n8876), .Z(n8881) );
  NAND U9106 ( .A(n8879), .B(n8878), .Z(n8880) );
  AND U9107 ( .A(n8881), .B(n8880), .Z(n8897) );
  XNOR U9108 ( .A(n8896), .B(n8897), .Z(n8889) );
  NAND U9109 ( .A(n8883), .B(n8882), .Z(n8887) );
  NAND U9110 ( .A(n8885), .B(n8884), .Z(n8886) );
  AND U9111 ( .A(n8887), .B(n8886), .Z(n8888) );
  XNOR U9112 ( .A(n8889), .B(n8888), .Z(n8890) );
  XOR U9113 ( .A(n8891), .B(n8890), .Z(n8980) );
  XOR U9114 ( .A(n8981), .B(n8980), .Z(c[108]) );
  NANDN U9115 ( .A(n8889), .B(n8888), .Z(n8893) );
  NAND U9116 ( .A(n8891), .B(n8890), .Z(n8892) );
  NAND U9117 ( .A(n8893), .B(n8892), .Z(n8986) );
  NANDN U9118 ( .A(n8895), .B(n8894), .Z(n8899) );
  NAND U9119 ( .A(n8897), .B(n8896), .Z(n8898) );
  AND U9120 ( .A(n8899), .B(n8898), .Z(n8985) );
  NANDN U9121 ( .A(n8901), .B(n8900), .Z(n8905) );
  NAND U9122 ( .A(n8903), .B(n8902), .Z(n8904) );
  NAND U9123 ( .A(n8905), .B(n8904), .Z(n8990) );
  OR U9124 ( .A(n8907), .B(n8906), .Z(n8911) );
  NANDN U9125 ( .A(n8909), .B(n8908), .Z(n8910) );
  NAND U9126 ( .A(n8911), .B(n8910), .Z(n9070) );
  OR U9127 ( .A(n8913), .B(n8912), .Z(n8917) );
  NANDN U9128 ( .A(n8915), .B(n8914), .Z(n8916) );
  AND U9129 ( .A(n8917), .B(n8916), .Z(n9069) );
  XNOR U9130 ( .A(n9070), .B(n9069), .Z(n9071) );
  NANDN U9131 ( .A(n8919), .B(n8918), .Z(n8923) );
  NAND U9132 ( .A(n8921), .B(n8920), .Z(n8922) );
  NAND U9133 ( .A(n8923), .B(n8922), .Z(n9000) );
  XNOR U9134 ( .A(b[23]), .B(a[55]), .Z(n9045) );
  OR U9135 ( .A(n9045), .B(n9621), .Z(n8926) );
  NAND U9136 ( .A(n9622), .B(n8924), .Z(n8925) );
  NAND U9137 ( .A(n8926), .B(n8925), .Z(n9053) );
  NAND U9138 ( .A(n8927), .B(n9105), .Z(n8929) );
  XNOR U9139 ( .A(a[61]), .B(n9455), .Z(n9042) );
  NAND U9140 ( .A(n9042), .B(n9107), .Z(n8928) );
  NAND U9141 ( .A(n8929), .B(n8928), .Z(n9051) );
  NAND U9142 ( .A(n8930), .B(n9914), .Z(n8932) );
  XNOR U9143 ( .A(n323), .B(a[47]), .Z(n9026) );
  NANDN U9144 ( .A(n9913), .B(n9026), .Z(n8931) );
  NAND U9145 ( .A(n8932), .B(n8931), .Z(n9052) );
  XOR U9146 ( .A(n9051), .B(n9052), .Z(n9054) );
  XNOR U9147 ( .A(n9053), .B(n9054), .Z(n9008) );
  XOR U9148 ( .A(b[27]), .B(n9457), .Z(n9029) );
  OR U9149 ( .A(n9029), .B(n9751), .Z(n8935) );
  NANDN U9150 ( .A(n8933), .B(n9801), .Z(n8934) );
  NAND U9151 ( .A(n8935), .B(n8934), .Z(n9059) );
  NANDN U9152 ( .A(n8936), .B(n9875), .Z(n8938) );
  XNOR U9153 ( .A(n322), .B(a[49]), .Z(n9032) );
  NANDN U9154 ( .A(n9874), .B(n9032), .Z(n8937) );
  NAND U9155 ( .A(n8938), .B(n8937), .Z(n9058) );
  NAND U9156 ( .A(n8939), .B(n9379), .Z(n8941) );
  XNOR U9157 ( .A(a[59]), .B(n9562), .Z(n9048) );
  NAND U9158 ( .A(n9048), .B(n9378), .Z(n8940) );
  NAND U9159 ( .A(n8941), .B(n8940), .Z(n9057) );
  XOR U9160 ( .A(n9058), .B(n9057), .Z(n9060) );
  XNOR U9161 ( .A(n9059), .B(n9060), .Z(n9005) );
  XNOR U9162 ( .A(a[57]), .B(b[21]), .Z(n9039) );
  NANDN U9163 ( .A(n9039), .B(n9493), .Z(n8944) );
  NAND U9164 ( .A(n9495), .B(n8942), .Z(n8943) );
  NAND U9165 ( .A(n8944), .B(n8943), .Z(n9006) );
  XNOR U9166 ( .A(n9005), .B(n9006), .Z(n9007) );
  XOR U9167 ( .A(n9008), .B(n9007), .Z(n8999) );
  XOR U9168 ( .A(n9000), .B(n8999), .Z(n9002) );
  XNOR U9169 ( .A(n9002), .B(n9001), .Z(n9066) );
  OR U9170 ( .A(n8950), .B(n8949), .Z(n8954) );
  NANDN U9171 ( .A(n8952), .B(n8951), .Z(n8953) );
  NAND U9172 ( .A(n8954), .B(n8953), .Z(n9064) );
  NANDN U9173 ( .A(n9011), .B(n8955), .Z(n8959) );
  NANDN U9174 ( .A(n8957), .B(n8956), .Z(n8958) );
  NAND U9175 ( .A(n8959), .B(n8958), .Z(n8996) );
  NANDN U9176 ( .A(n323), .B(a[45]), .Z(n9010) );
  XOR U9177 ( .A(n8960), .B(n9010), .Z(n9012) );
  XNOR U9178 ( .A(n9011), .B(n9012), .Z(n9015) );
  NANDN U9179 ( .A(n8962), .B(n8961), .Z(n8965) );
  XNOR U9180 ( .A(n9946), .B(b[15]), .Z(n9023) );
  NAND U9181 ( .A(n9023), .B(n8963), .Z(n8964) );
  NAND U9182 ( .A(n8965), .B(n8964), .Z(n9016) );
  XOR U9183 ( .A(n9015), .B(n9016), .Z(n9017) );
  XOR U9184 ( .A(b[25]), .B(n9564), .Z(n9036) );
  NANDN U9185 ( .A(n9036), .B(n9706), .Z(n8968) );
  NAND U9186 ( .A(n9707), .B(n8966), .Z(n8967) );
  NAND U9187 ( .A(n8968), .B(n8967), .Z(n9018) );
  XOR U9188 ( .A(n9017), .B(n9018), .Z(n8993) );
  XNOR U9189 ( .A(n8993), .B(n8994), .Z(n8995) );
  XOR U9190 ( .A(n8996), .B(n8995), .Z(n9063) );
  XNOR U9191 ( .A(n9064), .B(n9063), .Z(n9065) );
  XNOR U9192 ( .A(n9066), .B(n9065), .Z(n9072) );
  XOR U9193 ( .A(n9071), .B(n9072), .Z(n8987) );
  NAND U9194 ( .A(n8974), .B(n8973), .Z(n8978) );
  OR U9195 ( .A(n8976), .B(n8975), .Z(n8977) );
  AND U9196 ( .A(n8978), .B(n8977), .Z(n8988) );
  XNOR U9197 ( .A(n8987), .B(n8988), .Z(n8989) );
  XNOR U9198 ( .A(n8990), .B(n8989), .Z(n8984) );
  XOR U9199 ( .A(n8985), .B(n8984), .Z(n8979) );
  XOR U9200 ( .A(n8986), .B(n8979), .Z(n8982) );
  OR U9201 ( .A(n8981), .B(n8980), .Z(n8983) );
  XNOR U9202 ( .A(n8982), .B(n8983), .Z(c[109]) );
  NANDN U9203 ( .A(n8983), .B(n8982), .Z(n9156) );
  NANDN U9204 ( .A(n8988), .B(n8987), .Z(n8992) );
  NANDN U9205 ( .A(n8990), .B(n8989), .Z(n8991) );
  NAND U9206 ( .A(n8992), .B(n8991), .Z(n9076) );
  NANDN U9207 ( .A(n8994), .B(n8993), .Z(n8998) );
  NAND U9208 ( .A(n8996), .B(n8995), .Z(n8997) );
  NAND U9209 ( .A(n8998), .B(n8997), .Z(n9148) );
  NANDN U9210 ( .A(n9000), .B(n8999), .Z(n9004) );
  OR U9211 ( .A(n9002), .B(n9001), .Z(n9003) );
  NAND U9212 ( .A(n9004), .B(n9003), .Z(n9149) );
  XNOR U9213 ( .A(n9148), .B(n9149), .Z(n9150) );
  OR U9214 ( .A(n9010), .B(n9009), .Z(n9014) );
  NANDN U9215 ( .A(n9012), .B(n9011), .Z(n9013) );
  NAND U9216 ( .A(n9014), .B(n9013), .Z(n9085) );
  OR U9217 ( .A(n9016), .B(n9015), .Z(n9020) );
  NANDN U9218 ( .A(n9018), .B(n9017), .Z(n9019) );
  NAND U9219 ( .A(n9020), .B(n9019), .Z(n9086) );
  XNOR U9220 ( .A(n9085), .B(n9086), .Z(n9087) );
  XNOR U9221 ( .A(b[15]), .B(n9021), .Z(n9025) );
  XNOR U9222 ( .A(b[14]), .B(b[13]), .Z(n9022) );
  NANDN U9223 ( .A(n9023), .B(n9022), .Z(n9024) );
  AND U9224 ( .A(n9025), .B(n9024), .Z(n9132) );
  NAND U9225 ( .A(n9026), .B(n9914), .Z(n9028) );
  XNOR U9226 ( .A(n323), .B(a[48]), .Z(n9116) );
  NANDN U9227 ( .A(n9913), .B(n9116), .Z(n9027) );
  NAND U9228 ( .A(n9028), .B(n9027), .Z(n9131) );
  AND U9229 ( .A(b[31]), .B(a[46]), .Z(n9209) );
  XOR U9230 ( .A(n9131), .B(n9209), .Z(n9133) );
  XOR U9231 ( .A(n9132), .B(n9133), .Z(n9088) );
  XOR U9232 ( .A(n9087), .B(n9088), .Z(n9143) );
  XOR U9233 ( .A(n9142), .B(n9143), .Z(n9144) );
  NANDN U9234 ( .A(n9029), .B(n9801), .Z(n9031) );
  XOR U9235 ( .A(b[27]), .B(n9217), .Z(n9122) );
  OR U9236 ( .A(n9122), .B(n9751), .Z(n9030) );
  NAND U9237 ( .A(n9031), .B(n9030), .Z(n9113) );
  NAND U9238 ( .A(n9032), .B(n9875), .Z(n9035) );
  XOR U9239 ( .A(n322), .B(n9033), .Z(n9125) );
  NANDN U9240 ( .A(n9874), .B(n9125), .Z(n9034) );
  NAND U9241 ( .A(n9035), .B(n9034), .Z(n9110) );
  XOR U9242 ( .A(b[25]), .B(n9353), .Z(n9119) );
  NANDN U9243 ( .A(n9119), .B(n9706), .Z(n9038) );
  NANDN U9244 ( .A(n9036), .B(n9707), .Z(n9037) );
  AND U9245 ( .A(n9038), .B(n9037), .Z(n9111) );
  XNOR U9246 ( .A(n9110), .B(n9111), .Z(n9112) );
  XNOR U9247 ( .A(n9113), .B(n9112), .Z(n9139) );
  XNOR U9248 ( .A(a[58]), .B(b[21]), .Z(n9128) );
  NANDN U9249 ( .A(n9128), .B(n9493), .Z(n9041) );
  NANDN U9250 ( .A(n9039), .B(n9495), .Z(n9040) );
  NAND U9251 ( .A(n9041), .B(n9040), .Z(n9098) );
  NAND U9252 ( .A(n9042), .B(n9105), .Z(n9044) );
  XNOR U9253 ( .A(n9810), .B(b[17]), .Z(n9106) );
  NAND U9254 ( .A(n9106), .B(n9107), .Z(n9043) );
  NAND U9255 ( .A(n9044), .B(n9043), .Z(n9095) );
  NANDN U9256 ( .A(n9045), .B(n9622), .Z(n9047) );
  XOR U9257 ( .A(b[23]), .B(n9357), .Z(n9099) );
  OR U9258 ( .A(n9099), .B(n9621), .Z(n9046) );
  AND U9259 ( .A(n9047), .B(n9046), .Z(n9096) );
  XNOR U9260 ( .A(n9095), .B(n9096), .Z(n9097) );
  XNOR U9261 ( .A(n9098), .B(n9097), .Z(n9136) );
  NAND U9262 ( .A(n9048), .B(n9379), .Z(n9050) );
  XNOR U9263 ( .A(n9805), .B(b[19]), .Z(n9102) );
  NAND U9264 ( .A(n9102), .B(n9378), .Z(n9049) );
  NAND U9265 ( .A(n9050), .B(n9049), .Z(n9137) );
  XNOR U9266 ( .A(n9136), .B(n9137), .Z(n9138) );
  XNOR U9267 ( .A(n9139), .B(n9138), .Z(n9094) );
  NAND U9268 ( .A(n9052), .B(n9051), .Z(n9056) );
  NAND U9269 ( .A(n9054), .B(n9053), .Z(n9055) );
  NAND U9270 ( .A(n9056), .B(n9055), .Z(n9091) );
  NAND U9271 ( .A(n9058), .B(n9057), .Z(n9062) );
  NAND U9272 ( .A(n9060), .B(n9059), .Z(n9061) );
  AND U9273 ( .A(n9062), .B(n9061), .Z(n9092) );
  XNOR U9274 ( .A(n9091), .B(n9092), .Z(n9093) );
  XNOR U9275 ( .A(n9094), .B(n9093), .Z(n9145) );
  XNOR U9276 ( .A(n9144), .B(n9145), .Z(n9151) );
  XNOR U9277 ( .A(n9150), .B(n9151), .Z(n9081) );
  NANDN U9278 ( .A(n9064), .B(n9063), .Z(n9068) );
  NAND U9279 ( .A(n9066), .B(n9065), .Z(n9067) );
  NAND U9280 ( .A(n9068), .B(n9067), .Z(n9082) );
  XNOR U9281 ( .A(n9081), .B(n9082), .Z(n9083) );
  NANDN U9282 ( .A(n9070), .B(n9069), .Z(n9074) );
  NANDN U9283 ( .A(n9072), .B(n9071), .Z(n9073) );
  AND U9284 ( .A(n9074), .B(n9073), .Z(n9084) );
  XOR U9285 ( .A(n9083), .B(n9084), .Z(n9075) );
  XOR U9286 ( .A(n9076), .B(n9075), .Z(n9078) );
  XOR U9287 ( .A(n9077), .B(n9078), .Z(n9155) );
  XOR U9288 ( .A(n9156), .B(n9155), .Z(c[110]) );
  NAND U9289 ( .A(n9076), .B(n9075), .Z(n9080) );
  NAND U9290 ( .A(n9078), .B(n9077), .Z(n9079) );
  AND U9291 ( .A(n9080), .B(n9079), .Z(n9159) );
  NANDN U9292 ( .A(n9086), .B(n9085), .Z(n9090) );
  NANDN U9293 ( .A(n9088), .B(n9087), .Z(n9089) );
  NAND U9294 ( .A(n9090), .B(n9089), .Z(n9160) );
  XOR U9295 ( .A(n9160), .B(n9161), .Z(n9163) );
  NANDN U9296 ( .A(n9099), .B(n9622), .Z(n9101) );
  XNOR U9297 ( .A(b[23]), .B(a[57]), .Z(n9220) );
  OR U9298 ( .A(n9220), .B(n9621), .Z(n9100) );
  NAND U9299 ( .A(n9101), .B(n9100), .Z(n9174) );
  NAND U9300 ( .A(n9102), .B(n9379), .Z(n9104) );
  XNOR U9301 ( .A(a[61]), .B(n9562), .Z(n9181) );
  NAND U9302 ( .A(n9181), .B(n9378), .Z(n9103) );
  NAND U9303 ( .A(n9104), .B(n9103), .Z(n9172) );
  NAND U9304 ( .A(n9106), .B(n9105), .Z(n9109) );
  XNOR U9305 ( .A(n9946), .B(b[17]), .Z(n9189) );
  NAND U9306 ( .A(n9189), .B(n9107), .Z(n9108) );
  NAND U9307 ( .A(n9109), .B(n9108), .Z(n9173) );
  XOR U9308 ( .A(n9172), .B(n9173), .Z(n9175) );
  XNOR U9309 ( .A(n9174), .B(n9175), .Z(n9227) );
  NANDN U9310 ( .A(n9111), .B(n9110), .Z(n9115) );
  NAND U9311 ( .A(n9113), .B(n9112), .Z(n9114) );
  NAND U9312 ( .A(n9115), .B(n9114), .Z(n9228) );
  XOR U9313 ( .A(n9227), .B(n9228), .Z(n9230) );
  XNOR U9314 ( .A(n9229), .B(n9230), .Z(n9169) );
  NAND U9315 ( .A(n9116), .B(n9914), .Z(n9118) );
  XNOR U9316 ( .A(n323), .B(a[49]), .Z(n9192) );
  NANDN U9317 ( .A(n9913), .B(n9192), .Z(n9117) );
  NAND U9318 ( .A(n9118), .B(n9117), .Z(n9195) );
  XNOR U9319 ( .A(b[25]), .B(a[55]), .Z(n9213) );
  NANDN U9320 ( .A(n9213), .B(n9706), .Z(n9121) );
  NANDN U9321 ( .A(n9119), .B(n9707), .Z(n9120) );
  AND U9322 ( .A(n9121), .B(n9120), .Z(n9196) );
  XOR U9323 ( .A(n9195), .B(n9196), .Z(n9198) );
  NANDN U9324 ( .A(n323), .B(a[47]), .Z(n9208) );
  XOR U9325 ( .A(n9207), .B(n9208), .Z(n9210) );
  XOR U9326 ( .A(n9209), .B(n9210), .Z(n9197) );
  XNOR U9327 ( .A(n9198), .B(n9197), .Z(n9226) );
  NANDN U9328 ( .A(n9122), .B(n9801), .Z(n9124) );
  XOR U9329 ( .A(b[27]), .B(n9564), .Z(n9184) );
  OR U9330 ( .A(n9184), .B(n9751), .Z(n9123) );
  NAND U9331 ( .A(n9124), .B(n9123), .Z(n9204) );
  NAND U9332 ( .A(n9875), .B(n9125), .Z(n9127) );
  XOR U9333 ( .A(n322), .B(n9457), .Z(n9216) );
  NANDN U9334 ( .A(n9874), .B(n9216), .Z(n9126) );
  NAND U9335 ( .A(n9127), .B(n9126), .Z(n9201) );
  XNOR U9336 ( .A(a[59]), .B(b[21]), .Z(n9178) );
  NANDN U9337 ( .A(n9178), .B(n9493), .Z(n9130) );
  NANDN U9338 ( .A(n9128), .B(n9495), .Z(n9129) );
  AND U9339 ( .A(n9130), .B(n9129), .Z(n9202) );
  XNOR U9340 ( .A(n9201), .B(n9202), .Z(n9203) );
  XNOR U9341 ( .A(n9204), .B(n9203), .Z(n9223) );
  NANDN U9342 ( .A(n9209), .B(n9131), .Z(n9135) );
  NANDN U9343 ( .A(n9133), .B(n9132), .Z(n9134) );
  NAND U9344 ( .A(n9135), .B(n9134), .Z(n9224) );
  XNOR U9345 ( .A(n9223), .B(n9224), .Z(n9225) );
  XNOR U9346 ( .A(n9226), .B(n9225), .Z(n9166) );
  NANDN U9347 ( .A(n9137), .B(n9136), .Z(n9141) );
  NAND U9348 ( .A(n9139), .B(n9138), .Z(n9140) );
  NAND U9349 ( .A(n9141), .B(n9140), .Z(n9167) );
  XNOR U9350 ( .A(n9166), .B(n9167), .Z(n9168) );
  XNOR U9351 ( .A(n9169), .B(n9168), .Z(n9162) );
  XNOR U9352 ( .A(n9163), .B(n9162), .Z(n9233) );
  OR U9353 ( .A(n9143), .B(n9142), .Z(n9147) );
  NANDN U9354 ( .A(n9145), .B(n9144), .Z(n9146) );
  NAND U9355 ( .A(n9147), .B(n9146), .Z(n9234) );
  XNOR U9356 ( .A(n9233), .B(n9234), .Z(n9235) );
  NANDN U9357 ( .A(n9149), .B(n9148), .Z(n9153) );
  NAND U9358 ( .A(n9151), .B(n9150), .Z(n9152) );
  NAND U9359 ( .A(n9153), .B(n9152), .Z(n9236) );
  XNOR U9360 ( .A(n9235), .B(n9236), .Z(n9157) );
  XNOR U9361 ( .A(n9158), .B(n9157), .Z(n9154) );
  XNOR U9362 ( .A(n9159), .B(n9154), .Z(n9240) );
  OR U9363 ( .A(n9156), .B(n9155), .Z(n9239) );
  XOR U9364 ( .A(n9240), .B(n9239), .Z(c[111]) );
  NANDN U9365 ( .A(n9161), .B(n9160), .Z(n9165) );
  OR U9366 ( .A(n9163), .B(n9162), .Z(n9164) );
  NAND U9367 ( .A(n9165), .B(n9164), .Z(n9252) );
  NANDN U9368 ( .A(n9167), .B(n9166), .Z(n9171) );
  NAND U9369 ( .A(n9169), .B(n9168), .Z(n9170) );
  NAND U9370 ( .A(n9171), .B(n9170), .Z(n9250) );
  NAND U9371 ( .A(n9173), .B(n9172), .Z(n9177) );
  NAND U9372 ( .A(n9175), .B(n9174), .Z(n9176) );
  NAND U9373 ( .A(n9177), .B(n9176), .Z(n9297) );
  XOR U9374 ( .A(n9805), .B(n318), .Z(n9285) );
  NAND U9375 ( .A(n9285), .B(n9493), .Z(n9180) );
  NANDN U9376 ( .A(n9178), .B(n9495), .Z(n9179) );
  NAND U9377 ( .A(n9180), .B(n9179), .Z(n9310) );
  NAND U9378 ( .A(n9181), .B(n9379), .Z(n9183) );
  XNOR U9379 ( .A(n9810), .B(b[19]), .Z(n9273) );
  NAND U9380 ( .A(n9273), .B(n9378), .Z(n9182) );
  NAND U9381 ( .A(n9183), .B(n9182), .Z(n9307) );
  NANDN U9382 ( .A(n9184), .B(n9801), .Z(n9186) );
  XOR U9383 ( .A(b[27]), .B(n9353), .Z(n9276) );
  OR U9384 ( .A(n9276), .B(n9751), .Z(n9185) );
  AND U9385 ( .A(n9186), .B(n9185), .Z(n9308) );
  XNOR U9386 ( .A(n9307), .B(n9308), .Z(n9309) );
  XNOR U9387 ( .A(n9310), .B(n9309), .Z(n9295) );
  XOR U9388 ( .A(n9455), .B(n9187), .Z(n9191) );
  XNOR U9389 ( .A(b[16]), .B(b[15]), .Z(n9188) );
  NANDN U9390 ( .A(n9189), .B(n9188), .Z(n9190) );
  AND U9391 ( .A(n9191), .B(n9190), .Z(n9312) );
  NAND U9392 ( .A(n9192), .B(n9914), .Z(n9194) );
  XNOR U9393 ( .A(n323), .B(a[50]), .Z(n9288) );
  NANDN U9394 ( .A(n9913), .B(n9288), .Z(n9193) );
  NAND U9395 ( .A(n9194), .B(n9193), .Z(n9311) );
  AND U9396 ( .A(b[31]), .B(a[48]), .Z(n9374) );
  XOR U9397 ( .A(n9311), .B(n9374), .Z(n9313) );
  XNOR U9398 ( .A(n9312), .B(n9313), .Z(n9296) );
  XOR U9399 ( .A(n9295), .B(n9296), .Z(n9298) );
  XNOR U9400 ( .A(n9297), .B(n9298), .Z(n9261) );
  NANDN U9401 ( .A(n9196), .B(n9195), .Z(n9200) );
  OR U9402 ( .A(n9198), .B(n9197), .Z(n9199) );
  AND U9403 ( .A(n9200), .B(n9199), .Z(n9262) );
  XNOR U9404 ( .A(n9261), .B(n9262), .Z(n9263) );
  NANDN U9405 ( .A(n9202), .B(n9201), .Z(n9206) );
  NAND U9406 ( .A(n9204), .B(n9203), .Z(n9205) );
  NAND U9407 ( .A(n9206), .B(n9205), .Z(n9304) );
  NANDN U9408 ( .A(n9208), .B(n9207), .Z(n9212) );
  NANDN U9409 ( .A(n9210), .B(n9209), .Z(n9211) );
  NAND U9410 ( .A(n9212), .B(n9211), .Z(n9301) );
  XOR U9411 ( .A(n320), .B(n9357), .Z(n9291) );
  NAND U9412 ( .A(n9291), .B(n9706), .Z(n9215) );
  NANDN U9413 ( .A(n9213), .B(n9707), .Z(n9214) );
  NAND U9414 ( .A(n9215), .B(n9214), .Z(n9270) );
  NAND U9415 ( .A(n9875), .B(n9216), .Z(n9219) );
  XOR U9416 ( .A(n322), .B(n9217), .Z(n9279) );
  NANDN U9417 ( .A(n9874), .B(n9279), .Z(n9218) );
  NAND U9418 ( .A(n9219), .B(n9218), .Z(n9267) );
  NANDN U9419 ( .A(n9220), .B(n9622), .Z(n9222) );
  XNOR U9420 ( .A(a[58]), .B(b[23]), .Z(n9282) );
  OR U9421 ( .A(n9282), .B(n9621), .Z(n9221) );
  AND U9422 ( .A(n9222), .B(n9221), .Z(n9268) );
  XNOR U9423 ( .A(n9267), .B(n9268), .Z(n9269) );
  XNOR U9424 ( .A(n9270), .B(n9269), .Z(n9302) );
  XNOR U9425 ( .A(n9301), .B(n9302), .Z(n9303) );
  XNOR U9426 ( .A(n9304), .B(n9303), .Z(n9264) );
  XOR U9427 ( .A(n9263), .B(n9264), .Z(n9258) );
  NANDN U9428 ( .A(n9228), .B(n9227), .Z(n9232) );
  OR U9429 ( .A(n9230), .B(n9229), .Z(n9231) );
  AND U9430 ( .A(n9232), .B(n9231), .Z(n9256) );
  XNOR U9431 ( .A(n9255), .B(n9256), .Z(n9257) );
  XOR U9432 ( .A(n9258), .B(n9257), .Z(n9249) );
  XNOR U9433 ( .A(n9250), .B(n9249), .Z(n9251) );
  XOR U9434 ( .A(n9252), .B(n9251), .Z(n9243) );
  NANDN U9435 ( .A(n9234), .B(n9233), .Z(n9238) );
  NANDN U9436 ( .A(n9236), .B(n9235), .Z(n9237) );
  NAND U9437 ( .A(n9238), .B(n9237), .Z(n9244) );
  XNOR U9438 ( .A(n9243), .B(n9244), .Z(n9245) );
  XNOR U9439 ( .A(n9246), .B(n9245), .Z(n9241) );
  OR U9440 ( .A(n9240), .B(n9239), .Z(n9242) );
  XNOR U9441 ( .A(n9241), .B(n9242), .Z(c[112]) );
  NANDN U9442 ( .A(n9242), .B(n9241), .Z(n9318) );
  NANDN U9443 ( .A(n9244), .B(n9243), .Z(n9248) );
  NANDN U9444 ( .A(n9246), .B(n9245), .Z(n9247) );
  AND U9445 ( .A(n9248), .B(n9247), .Z(n9321) );
  NANDN U9446 ( .A(n9250), .B(n9249), .Z(n9254) );
  NANDN U9447 ( .A(n9252), .B(n9251), .Z(n9253) );
  AND U9448 ( .A(n9254), .B(n9253), .Z(n9320) );
  NANDN U9449 ( .A(n9256), .B(n9255), .Z(n9260) );
  NAND U9450 ( .A(n9258), .B(n9257), .Z(n9259) );
  NAND U9451 ( .A(n9260), .B(n9259), .Z(n9389) );
  NANDN U9452 ( .A(n9262), .B(n9261), .Z(n9266) );
  NANDN U9453 ( .A(n9264), .B(n9263), .Z(n9265) );
  NAND U9454 ( .A(n9266), .B(n9265), .Z(n9387) );
  NANDN U9455 ( .A(n9268), .B(n9267), .Z(n9272) );
  NAND U9456 ( .A(n9270), .B(n9269), .Z(n9271) );
  NAND U9457 ( .A(n9272), .B(n9271), .Z(n9337) );
  NAND U9458 ( .A(n9273), .B(n9379), .Z(n9275) );
  XOR U9459 ( .A(a[63]), .B(n9562), .Z(n9380) );
  NANDN U9460 ( .A(n9380), .B(n9378), .Z(n9274) );
  NAND U9461 ( .A(n9275), .B(n9274), .Z(n9366) );
  NANDN U9462 ( .A(n9276), .B(n9801), .Z(n9278) );
  XNOR U9463 ( .A(b[27]), .B(a[55]), .Z(n9356) );
  OR U9464 ( .A(n9356), .B(n9751), .Z(n9277) );
  AND U9465 ( .A(n9278), .B(n9277), .Z(n9367) );
  XOR U9466 ( .A(n9366), .B(n9367), .Z(n9369) );
  NANDN U9467 ( .A(n323), .B(a[49]), .Z(n9373) );
  XNOR U9468 ( .A(n9372), .B(n9373), .Z(n9375) );
  XOR U9469 ( .A(n9374), .B(n9375), .Z(n9368) );
  XNOR U9470 ( .A(n9369), .B(n9368), .Z(n9334) );
  NAND U9471 ( .A(n9875), .B(n9279), .Z(n9281) );
  XOR U9472 ( .A(n322), .B(n9564), .Z(n9352) );
  NANDN U9473 ( .A(n9874), .B(n9352), .Z(n9280) );
  NAND U9474 ( .A(n9281), .B(n9280), .Z(n9343) );
  NANDN U9475 ( .A(n9282), .B(n9622), .Z(n9284) );
  XNOR U9476 ( .A(a[59]), .B(b[23]), .Z(n9363) );
  OR U9477 ( .A(n9363), .B(n9621), .Z(n9283) );
  NAND U9478 ( .A(n9284), .B(n9283), .Z(n9340) );
  XNOR U9479 ( .A(a[61]), .B(b[21]), .Z(n9360) );
  NANDN U9480 ( .A(n9360), .B(n9493), .Z(n9287) );
  NAND U9481 ( .A(n9495), .B(n9285), .Z(n9286) );
  AND U9482 ( .A(n9287), .B(n9286), .Z(n9348) );
  NAND U9483 ( .A(n9288), .B(n9914), .Z(n9290) );
  XNOR U9484 ( .A(n323), .B(a[51]), .Z(n9383) );
  NANDN U9485 ( .A(n9913), .B(n9383), .Z(n9289) );
  NAND U9486 ( .A(n9290), .B(n9289), .Z(n9346) );
  XNOR U9487 ( .A(b[25]), .B(a[57]), .Z(n9349) );
  NANDN U9488 ( .A(n9349), .B(n9706), .Z(n9293) );
  NAND U9489 ( .A(n9707), .B(n9291), .Z(n9292) );
  AND U9490 ( .A(n9293), .B(n9292), .Z(n9347) );
  XOR U9491 ( .A(n9346), .B(n9347), .Z(n9294) );
  XNOR U9492 ( .A(n9348), .B(n9294), .Z(n9341) );
  XNOR U9493 ( .A(n9340), .B(n9341), .Z(n9342) );
  XOR U9494 ( .A(n9343), .B(n9342), .Z(n9335) );
  XNOR U9495 ( .A(n9334), .B(n9335), .Z(n9336) );
  XOR U9496 ( .A(n9337), .B(n9336), .Z(n9322) );
  NANDN U9497 ( .A(n9296), .B(n9295), .Z(n9300) );
  OR U9498 ( .A(n9298), .B(n9297), .Z(n9299) );
  NAND U9499 ( .A(n9300), .B(n9299), .Z(n9323) );
  XNOR U9500 ( .A(n9322), .B(n9323), .Z(n9324) );
  NANDN U9501 ( .A(n9302), .B(n9301), .Z(n9306) );
  NAND U9502 ( .A(n9304), .B(n9303), .Z(n9305) );
  NAND U9503 ( .A(n9306), .B(n9305), .Z(n9331) );
  NANDN U9504 ( .A(n9374), .B(n9311), .Z(n9315) );
  NANDN U9505 ( .A(n9313), .B(n9312), .Z(n9314) );
  AND U9506 ( .A(n9315), .B(n9314), .Z(n9329) );
  XNOR U9507 ( .A(n9328), .B(n9329), .Z(n9330) );
  XOR U9508 ( .A(n9331), .B(n9330), .Z(n9325) );
  XOR U9509 ( .A(n9324), .B(n9325), .Z(n9386) );
  XNOR U9510 ( .A(n9387), .B(n9386), .Z(n9388) );
  XOR U9511 ( .A(n9389), .B(n9388), .Z(n9319) );
  XNOR U9512 ( .A(n9320), .B(n9319), .Z(n9316) );
  XNOR U9513 ( .A(n9321), .B(n9316), .Z(n9317) );
  XOR U9514 ( .A(n9318), .B(n9317), .Z(c[113]) );
  OR U9515 ( .A(n9318), .B(n9317), .Z(n9459) );
  NANDN U9516 ( .A(n9323), .B(n9322), .Z(n9327) );
  NAND U9517 ( .A(n9325), .B(n9324), .Z(n9326) );
  NAND U9518 ( .A(n9327), .B(n9326), .Z(n9401) );
  NANDN U9519 ( .A(n9329), .B(n9328), .Z(n9333) );
  NAND U9520 ( .A(n9331), .B(n9330), .Z(n9332) );
  NAND U9521 ( .A(n9333), .B(n9332), .Z(n9399) );
  NANDN U9522 ( .A(n9335), .B(n9334), .Z(n9339) );
  NANDN U9523 ( .A(n9337), .B(n9336), .Z(n9338) );
  NAND U9524 ( .A(n9339), .B(n9338), .Z(n9405) );
  NANDN U9525 ( .A(n9341), .B(n9340), .Z(n9345) );
  NAND U9526 ( .A(n9343), .B(n9342), .Z(n9344) );
  NAND U9527 ( .A(n9345), .B(n9344), .Z(n9403) );
  XNOR U9528 ( .A(b[25]), .B(a[58]), .Z(n9440) );
  NANDN U9529 ( .A(n9440), .B(n9706), .Z(n9351) );
  NANDN U9530 ( .A(n9349), .B(n9707), .Z(n9350) );
  NAND U9531 ( .A(n9351), .B(n9350), .Z(n9434) );
  NAND U9532 ( .A(n9875), .B(n9352), .Z(n9355) );
  XOR U9533 ( .A(n322), .B(n9353), .Z(n9437) );
  NANDN U9534 ( .A(n9874), .B(n9437), .Z(n9354) );
  NAND U9535 ( .A(n9355), .B(n9354), .Z(n9431) );
  NANDN U9536 ( .A(n9356), .B(n9801), .Z(n9359) );
  XOR U9537 ( .A(b[27]), .B(n9357), .Z(n9452) );
  OR U9538 ( .A(n9452), .B(n9751), .Z(n9358) );
  AND U9539 ( .A(n9359), .B(n9358), .Z(n9432) );
  XNOR U9540 ( .A(n9431), .B(n9432), .Z(n9433) );
  XNOR U9541 ( .A(n9434), .B(n9433), .Z(n9417) );
  XOR U9542 ( .A(a[62]), .B(n318), .Z(n9449) );
  NANDN U9543 ( .A(n9449), .B(n9493), .Z(n9362) );
  NANDN U9544 ( .A(n9360), .B(n9495), .Z(n9361) );
  NAND U9545 ( .A(n9362), .B(n9361), .Z(n9414) );
  NANDN U9546 ( .A(n9363), .B(n9622), .Z(n9365) );
  XOR U9547 ( .A(a[60]), .B(n319), .Z(n9446) );
  OR U9548 ( .A(n9446), .B(n9621), .Z(n9364) );
  AND U9549 ( .A(n9365), .B(n9364), .Z(n9415) );
  XNOR U9550 ( .A(n9414), .B(n9415), .Z(n9416) );
  XOR U9551 ( .A(n9417), .B(n9416), .Z(n9409) );
  XNOR U9552 ( .A(n9408), .B(n9409), .Z(n9410) );
  NANDN U9553 ( .A(n9367), .B(n9366), .Z(n9371) );
  OR U9554 ( .A(n9369), .B(n9368), .Z(n9370) );
  NAND U9555 ( .A(n9371), .B(n9370), .Z(n9422) );
  OR U9556 ( .A(n9373), .B(n9372), .Z(n9377) );
  NANDN U9557 ( .A(n9375), .B(n9374), .Z(n9376) );
  NAND U9558 ( .A(n9377), .B(n9376), .Z(n9421) );
  NANDN U9559 ( .A(n9562), .B(n9378), .Z(n9382) );
  NANDN U9560 ( .A(n9380), .B(n9379), .Z(n9381) );
  NAND U9561 ( .A(n9382), .B(n9381), .Z(n9427) );
  NAND U9562 ( .A(n9383), .B(n9914), .Z(n9385) );
  XNOR U9563 ( .A(n323), .B(a[52]), .Z(n9443) );
  NANDN U9564 ( .A(n9913), .B(n9443), .Z(n9384) );
  NAND U9565 ( .A(n9385), .B(n9384), .Z(n9426) );
  ANDN U9566 ( .B(a[50]), .A(n323), .Z(n9510) );
  XOR U9567 ( .A(n9426), .B(n9510), .Z(n9428) );
  XNOR U9568 ( .A(n9427), .B(n9428), .Z(n9420) );
  XNOR U9569 ( .A(n9421), .B(n9420), .Z(n9423) );
  XNOR U9570 ( .A(n9422), .B(n9423), .Z(n9411) );
  XOR U9571 ( .A(n9410), .B(n9411), .Z(n9402) );
  XOR U9572 ( .A(n9403), .B(n9402), .Z(n9404) );
  XNOR U9573 ( .A(n9405), .B(n9404), .Z(n9398) );
  XOR U9574 ( .A(n9399), .B(n9398), .Z(n9400) );
  XNOR U9575 ( .A(n9401), .B(n9400), .Z(n9392) );
  NAND U9576 ( .A(n9387), .B(n9386), .Z(n9391) );
  OR U9577 ( .A(n9389), .B(n9388), .Z(n9390) );
  NAND U9578 ( .A(n9391), .B(n9390), .Z(n9393) );
  XOR U9579 ( .A(n9392), .B(n9393), .Z(n9395) );
  XOR U9580 ( .A(n9394), .B(n9395), .Z(n9458) );
  XOR U9581 ( .A(n9459), .B(n9458), .Z(c[114]) );
  NANDN U9582 ( .A(n9393), .B(n9392), .Z(n9397) );
  OR U9583 ( .A(n9395), .B(n9394), .Z(n9396) );
  NAND U9584 ( .A(n9397), .B(n9396), .Z(n9463) );
  NAND U9585 ( .A(n9403), .B(n9402), .Z(n9407) );
  NANDN U9586 ( .A(n9405), .B(n9404), .Z(n9406) );
  NAND U9587 ( .A(n9407), .B(n9406), .Z(n9468) );
  NANDN U9588 ( .A(n9409), .B(n9408), .Z(n9413) );
  NAND U9589 ( .A(n9411), .B(n9410), .Z(n9412) );
  NAND U9590 ( .A(n9413), .B(n9412), .Z(n9467) );
  NANDN U9591 ( .A(n9415), .B(n9414), .Z(n9419) );
  NANDN U9592 ( .A(n9417), .B(n9416), .Z(n9418) );
  NAND U9593 ( .A(n9419), .B(n9418), .Z(n9472) );
  NAND U9594 ( .A(n9421), .B(n9420), .Z(n9425) );
  NANDN U9595 ( .A(n9423), .B(n9422), .Z(n9424) );
  AND U9596 ( .A(n9425), .B(n9424), .Z(n9473) );
  XNOR U9597 ( .A(n9472), .B(n9473), .Z(n9474) );
  NANDN U9598 ( .A(n9510), .B(n9426), .Z(n9430) );
  NANDN U9599 ( .A(n9428), .B(n9427), .Z(n9429) );
  NAND U9600 ( .A(n9430), .B(n9429), .Z(n9520) );
  NANDN U9601 ( .A(n9432), .B(n9431), .Z(n9436) );
  NAND U9602 ( .A(n9434), .B(n9433), .Z(n9435) );
  AND U9603 ( .A(n9436), .B(n9435), .Z(n9521) );
  XNOR U9604 ( .A(n9520), .B(n9521), .Z(n9522) );
  NAND U9605 ( .A(n9875), .B(n9437), .Z(n9439) );
  XNOR U9606 ( .A(b[29]), .B(a[55]), .Z(n9487) );
  OR U9607 ( .A(n9487), .B(n9874), .Z(n9438) );
  NAND U9608 ( .A(n9439), .B(n9438), .Z(n9498) );
  XNOR U9609 ( .A(a[59]), .B(b[25]), .Z(n9478) );
  NANDN U9610 ( .A(n9478), .B(n9706), .Z(n9442) );
  NANDN U9611 ( .A(n9440), .B(n9707), .Z(n9441) );
  NAND U9612 ( .A(n9442), .B(n9441), .Z(n9507) );
  NAND U9613 ( .A(n9443), .B(n9914), .Z(n9445) );
  XNOR U9614 ( .A(n323), .B(a[53]), .Z(n9490) );
  NANDN U9615 ( .A(n9913), .B(n9490), .Z(n9444) );
  NAND U9616 ( .A(n9445), .B(n9444), .Z(n9504) );
  NANDN U9617 ( .A(n9446), .B(n9622), .Z(n9448) );
  XNOR U9618 ( .A(a[61]), .B(b[23]), .Z(n9481) );
  OR U9619 ( .A(n9481), .B(n9621), .Z(n9447) );
  AND U9620 ( .A(n9448), .B(n9447), .Z(n9505) );
  XNOR U9621 ( .A(n9504), .B(n9505), .Z(n9506) );
  XNOR U9622 ( .A(n9507), .B(n9506), .Z(n9499) );
  XNOR U9623 ( .A(n9498), .B(n9499), .Z(n9500) );
  XOR U9624 ( .A(n9946), .B(n318), .Z(n9494) );
  NAND U9625 ( .A(n9494), .B(n9493), .Z(n9451) );
  NANDN U9626 ( .A(n9449), .B(n9495), .Z(n9450) );
  NAND U9627 ( .A(n9451), .B(n9450), .Z(n9514) );
  NANDN U9628 ( .A(n9452), .B(n9801), .Z(n9454) );
  XNOR U9629 ( .A(b[27]), .B(a[57]), .Z(n9484) );
  OR U9630 ( .A(n9484), .B(n9751), .Z(n9453) );
  AND U9631 ( .A(n9454), .B(n9453), .Z(n9515) );
  XNOR U9632 ( .A(n9514), .B(n9515), .Z(n9516) );
  NANDN U9633 ( .A(n9455), .B(b[18]), .Z(n9456) );
  ANDN U9634 ( .B(n9456), .A(n9562), .Z(n9511) );
  XOR U9635 ( .A(n9510), .B(n9511), .Z(n9513) );
  NANDN U9636 ( .A(n9457), .B(b[31]), .Z(n9512) );
  XOR U9637 ( .A(n9513), .B(n9512), .Z(n9517) );
  XOR U9638 ( .A(n9516), .B(n9517), .Z(n9501) );
  XOR U9639 ( .A(n9500), .B(n9501), .Z(n9523) );
  XOR U9640 ( .A(n9522), .B(n9523), .Z(n9475) );
  XOR U9641 ( .A(n9474), .B(n9475), .Z(n9466) );
  XNOR U9642 ( .A(n9467), .B(n9466), .Z(n9469) );
  XNOR U9643 ( .A(n9468), .B(n9469), .Z(n9460) );
  XOR U9644 ( .A(n9461), .B(n9460), .Z(n9462) );
  XNOR U9645 ( .A(n9463), .B(n9462), .Z(n9526) );
  OR U9646 ( .A(n9459), .B(n9458), .Z(n9527) );
  XNOR U9647 ( .A(n9526), .B(n9527), .Z(c[115]) );
  NAND U9648 ( .A(n9461), .B(n9460), .Z(n9465) );
  NANDN U9649 ( .A(n9463), .B(n9462), .Z(n9464) );
  NAND U9650 ( .A(n9465), .B(n9464), .Z(n9531) );
  NAND U9651 ( .A(n9467), .B(n9466), .Z(n9471) );
  NANDN U9652 ( .A(n9469), .B(n9468), .Z(n9470) );
  NAND U9653 ( .A(n9471), .B(n9470), .Z(n9528) );
  NANDN U9654 ( .A(n9473), .B(n9472), .Z(n9477) );
  NAND U9655 ( .A(n9475), .B(n9474), .Z(n9476) );
  NAND U9656 ( .A(n9477), .B(n9476), .Z(n9537) );
  XOR U9657 ( .A(a[60]), .B(n320), .Z(n9565) );
  NANDN U9658 ( .A(n9565), .B(n9706), .Z(n9480) );
  NANDN U9659 ( .A(n9478), .B(n9707), .Z(n9479) );
  NAND U9660 ( .A(n9480), .B(n9479), .Z(n9553) );
  NANDN U9661 ( .A(n9481), .B(n9622), .Z(n9483) );
  XOR U9662 ( .A(a[62]), .B(n319), .Z(n9556) );
  OR U9663 ( .A(n9556), .B(n9621), .Z(n9482) );
  NAND U9664 ( .A(n9483), .B(n9482), .Z(n9550) );
  NANDN U9665 ( .A(n9484), .B(n9801), .Z(n9486) );
  XNOR U9666 ( .A(b[27]), .B(a[58]), .Z(n9559) );
  OR U9667 ( .A(n9559), .B(n9751), .Z(n9485) );
  AND U9668 ( .A(n9486), .B(n9485), .Z(n9551) );
  XNOR U9669 ( .A(n9550), .B(n9551), .Z(n9552) );
  XNOR U9670 ( .A(n9553), .B(n9552), .Z(n9546) );
  NANDN U9671 ( .A(n9487), .B(n9875), .Z(n9489) );
  XNOR U9672 ( .A(n322), .B(a[56]), .Z(n9571) );
  NANDN U9673 ( .A(n9874), .B(n9571), .Z(n9488) );
  NAND U9674 ( .A(n9489), .B(n9488), .Z(n9547) );
  XNOR U9675 ( .A(n9546), .B(n9547), .Z(n9548) );
  NAND U9676 ( .A(n9490), .B(n9914), .Z(n9492) );
  XNOR U9677 ( .A(n323), .B(a[54]), .Z(n9568) );
  NANDN U9678 ( .A(n9913), .B(n9568), .Z(n9491) );
  NAND U9679 ( .A(n9492), .B(n9491), .Z(n9575) );
  NANDN U9680 ( .A(n318), .B(n9493), .Z(n9497) );
  NAND U9681 ( .A(n9495), .B(n9494), .Z(n9496) );
  NAND U9682 ( .A(n9497), .B(n9496), .Z(n9574) );
  AND U9683 ( .A(a[52]), .B(b[31]), .Z(n9638) );
  XOR U9684 ( .A(n9574), .B(n9638), .Z(n9576) );
  XOR U9685 ( .A(n9575), .B(n9576), .Z(n9549) );
  XOR U9686 ( .A(n9548), .B(n9549), .Z(n9540) );
  NANDN U9687 ( .A(n9499), .B(n9498), .Z(n9503) );
  NAND U9688 ( .A(n9501), .B(n9500), .Z(n9502) );
  AND U9689 ( .A(n9503), .B(n9502), .Z(n9541) );
  XNOR U9690 ( .A(n9540), .B(n9541), .Z(n9542) );
  NANDN U9691 ( .A(n9505), .B(n9504), .Z(n9509) );
  NAND U9692 ( .A(n9507), .B(n9506), .Z(n9508) );
  NAND U9693 ( .A(n9509), .B(n9508), .Z(n9582) );
  NANDN U9694 ( .A(n9515), .B(n9514), .Z(n9519) );
  NAND U9695 ( .A(n9517), .B(n9516), .Z(n9518) );
  AND U9696 ( .A(n9519), .B(n9518), .Z(n9579) );
  XNOR U9697 ( .A(n9580), .B(n9579), .Z(n9581) );
  XOR U9698 ( .A(n9582), .B(n9581), .Z(n9543) );
  XNOR U9699 ( .A(n9542), .B(n9543), .Z(n9534) );
  NANDN U9700 ( .A(n9521), .B(n9520), .Z(n9525) );
  NAND U9701 ( .A(n9523), .B(n9522), .Z(n9524) );
  AND U9702 ( .A(n9525), .B(n9524), .Z(n9535) );
  XNOR U9703 ( .A(n9534), .B(n9535), .Z(n9536) );
  XNOR U9704 ( .A(n9537), .B(n9536), .Z(n9529) );
  XNOR U9705 ( .A(n9528), .B(n9529), .Z(n9530) );
  XNOR U9706 ( .A(n9531), .B(n9530), .Z(n9586) );
  NANDN U9707 ( .A(n9527), .B(n9526), .Z(n9585) );
  XOR U9708 ( .A(n9586), .B(n9585), .Z(c[116]) );
  NANDN U9709 ( .A(n9529), .B(n9528), .Z(n9533) );
  NAND U9710 ( .A(n9531), .B(n9530), .Z(n9532) );
  NAND U9711 ( .A(n9533), .B(n9532), .Z(n9597) );
  NANDN U9712 ( .A(n9535), .B(n9534), .Z(n9539) );
  NAND U9713 ( .A(n9537), .B(n9536), .Z(n9538) );
  NAND U9714 ( .A(n9539), .B(n9538), .Z(n9596) );
  NAND U9715 ( .A(n9541), .B(n9540), .Z(n9545) );
  OR U9716 ( .A(n9543), .B(n9542), .Z(n9544) );
  NAND U9717 ( .A(n9545), .B(n9544), .Z(n9591) );
  NANDN U9718 ( .A(n9551), .B(n9550), .Z(n9555) );
  NAND U9719 ( .A(n9553), .B(n9552), .Z(n9554) );
  NAND U9720 ( .A(n9555), .B(n9554), .Z(n9608) );
  NANDN U9721 ( .A(n9556), .B(n9622), .Z(n9558) );
  XOR U9722 ( .A(a[63]), .B(n319), .Z(n9623) );
  OR U9723 ( .A(n9623), .B(n9621), .Z(n9557) );
  NAND U9724 ( .A(n9558), .B(n9557), .Z(n9630) );
  NANDN U9725 ( .A(n9559), .B(n9801), .Z(n9561) );
  XNOR U9726 ( .A(b[27]), .B(a[59]), .Z(n9609) );
  OR U9727 ( .A(n9609), .B(n9751), .Z(n9560) );
  AND U9728 ( .A(n9561), .B(n9560), .Z(n9631) );
  XNOR U9729 ( .A(n9630), .B(n9631), .Z(n9632) );
  NANDN U9730 ( .A(n9562), .B(b[20]), .Z(n9563) );
  NANDN U9731 ( .A(n318), .B(n9563), .Z(n9637) );
  ANDN U9732 ( .B(b[31]), .A(n9564), .Z(n9636) );
  XNOR U9733 ( .A(n9637), .B(n9636), .Z(n9639) );
  XOR U9734 ( .A(n9638), .B(n9639), .Z(n9633) );
  XNOR U9735 ( .A(n9632), .B(n9633), .Z(n9605) );
  XNOR U9736 ( .A(a[61]), .B(b[25]), .Z(n9612) );
  NANDN U9737 ( .A(n9612), .B(n9706), .Z(n9567) );
  NANDN U9738 ( .A(n9565), .B(n9707), .Z(n9566) );
  NAND U9739 ( .A(n9567), .B(n9566), .Z(n9629) );
  NAND U9740 ( .A(n9568), .B(n9914), .Z(n9570) );
  XNOR U9741 ( .A(n323), .B(a[55]), .Z(n9618) );
  NANDN U9742 ( .A(n9913), .B(n9618), .Z(n9569) );
  NAND U9743 ( .A(n9570), .B(n9569), .Z(n9626) );
  NAND U9744 ( .A(n9571), .B(n9875), .Z(n9573) );
  XNOR U9745 ( .A(n322), .B(a[57]), .Z(n9615) );
  NANDN U9746 ( .A(n9874), .B(n9615), .Z(n9572) );
  AND U9747 ( .A(n9573), .B(n9572), .Z(n9627) );
  XNOR U9748 ( .A(n9626), .B(n9627), .Z(n9628) );
  XNOR U9749 ( .A(n9629), .B(n9628), .Z(n9606) );
  XNOR U9750 ( .A(n9605), .B(n9606), .Z(n9607) );
  XNOR U9751 ( .A(n9608), .B(n9607), .Z(n9601) );
  NANDN U9752 ( .A(n9574), .B(n9638), .Z(n9578) );
  OR U9753 ( .A(n9576), .B(n9575), .Z(n9577) );
  AND U9754 ( .A(n9578), .B(n9577), .Z(n9602) );
  XNOR U9755 ( .A(n9601), .B(n9602), .Z(n9603) );
  XNOR U9756 ( .A(n9604), .B(n9603), .Z(n9589) );
  NANDN U9757 ( .A(n9580), .B(n9579), .Z(n9584) );
  NANDN U9758 ( .A(n9582), .B(n9581), .Z(n9583) );
  NAND U9759 ( .A(n9584), .B(n9583), .Z(n9590) );
  XOR U9760 ( .A(n9589), .B(n9590), .Z(n9592) );
  XOR U9761 ( .A(n9591), .B(n9592), .Z(n9595) );
  XNOR U9762 ( .A(n9596), .B(n9595), .Z(n9598) );
  XNOR U9763 ( .A(n9597), .B(n9598), .Z(n9587) );
  OR U9764 ( .A(n9586), .B(n9585), .Z(n9588) );
  XNOR U9765 ( .A(n9587), .B(n9588), .Z(c[117]) );
  NANDN U9766 ( .A(n9588), .B(n9587), .Z(n9691) );
  NANDN U9767 ( .A(n9590), .B(n9589), .Z(n9594) );
  OR U9768 ( .A(n9592), .B(n9591), .Z(n9593) );
  NAND U9769 ( .A(n9594), .B(n9593), .Z(n9643) );
  NAND U9770 ( .A(n9596), .B(n9595), .Z(n9600) );
  NANDN U9771 ( .A(n9598), .B(n9597), .Z(n9599) );
  NAND U9772 ( .A(n9600), .B(n9599), .Z(n9645) );
  NANDN U9773 ( .A(n9609), .B(n9801), .Z(n9611) );
  XOR U9774 ( .A(b[27]), .B(n9805), .Z(n9675) );
  OR U9775 ( .A(n9675), .B(n9751), .Z(n9610) );
  NAND U9776 ( .A(n9611), .B(n9610), .Z(n9655) );
  XOR U9777 ( .A(n9810), .B(n320), .Z(n9671) );
  NAND U9778 ( .A(n9671), .B(n9706), .Z(n9614) );
  NANDN U9779 ( .A(n9612), .B(n9707), .Z(n9613) );
  NAND U9780 ( .A(n9614), .B(n9613), .Z(n9652) );
  NAND U9781 ( .A(n9875), .B(n9615), .Z(n9617) );
  XNOR U9782 ( .A(b[29]), .B(a[58]), .Z(n9666) );
  OR U9783 ( .A(n9666), .B(n9874), .Z(n9616) );
  AND U9784 ( .A(n9617), .B(n9616), .Z(n9653) );
  XNOR U9785 ( .A(n9652), .B(n9653), .Z(n9654) );
  XNOR U9786 ( .A(n9655), .B(n9654), .Z(n9679) );
  NAND U9787 ( .A(n9618), .B(n9914), .Z(n9620) );
  XNOR U9788 ( .A(n323), .B(a[56]), .Z(n9663) );
  NANDN U9789 ( .A(n9913), .B(n9663), .Z(n9619) );
  NAND U9790 ( .A(n9620), .B(n9619), .Z(n9659) );
  NANDN U9791 ( .A(n9621), .B(b[23]), .Z(n9625) );
  NANDN U9792 ( .A(n9623), .B(n9622), .Z(n9624) );
  NAND U9793 ( .A(n9625), .B(n9624), .Z(n9658) );
  AND U9794 ( .A(a[54]), .B(b[31]), .Z(n9713) );
  XOR U9795 ( .A(n9658), .B(n9713), .Z(n9660) );
  XOR U9796 ( .A(n9659), .B(n9660), .Z(n9678) );
  XOR U9797 ( .A(n9679), .B(n9678), .Z(n9680) );
  XOR U9798 ( .A(n9680), .B(n9681), .Z(n9687) );
  NANDN U9799 ( .A(n9631), .B(n9630), .Z(n9635) );
  NANDN U9800 ( .A(n9633), .B(n9632), .Z(n9634) );
  NAND U9801 ( .A(n9635), .B(n9634), .Z(n9684) );
  NAND U9802 ( .A(n9637), .B(n9636), .Z(n9641) );
  NANDN U9803 ( .A(n9639), .B(n9638), .Z(n9640) );
  AND U9804 ( .A(n9641), .B(n9640), .Z(n9685) );
  XNOR U9805 ( .A(n9684), .B(n9685), .Z(n9686) );
  XNOR U9806 ( .A(n9687), .B(n9686), .Z(n9647) );
  XNOR U9807 ( .A(n9646), .B(n9647), .Z(n9648) );
  XOR U9808 ( .A(n9649), .B(n9648), .Z(n9644) );
  XOR U9809 ( .A(n9645), .B(n9644), .Z(n9642) );
  XNOR U9810 ( .A(n9643), .B(n9642), .Z(n9690) );
  XNOR U9811 ( .A(n9691), .B(n9690), .Z(c[118]) );
  NANDN U9812 ( .A(n9647), .B(n9646), .Z(n9651) );
  NANDN U9813 ( .A(n9649), .B(n9648), .Z(n9650) );
  NAND U9814 ( .A(n9651), .B(n9650), .Z(n9694) );
  NANDN U9815 ( .A(n9653), .B(n9652), .Z(n9657) );
  NAND U9816 ( .A(n9655), .B(n9654), .Z(n9656) );
  NAND U9817 ( .A(n9657), .B(n9656), .Z(n9732) );
  NANDN U9818 ( .A(n9658), .B(n9713), .Z(n9662) );
  OR U9819 ( .A(n9660), .B(n9659), .Z(n9661) );
  NAND U9820 ( .A(n9662), .B(n9661), .Z(n9729) );
  NAND U9821 ( .A(n9663), .B(n9914), .Z(n9665) );
  XNOR U9822 ( .A(n323), .B(a[57]), .Z(n9703) );
  NANDN U9823 ( .A(n9913), .B(n9703), .Z(n9664) );
  NAND U9824 ( .A(n9665), .B(n9664), .Z(n9725) );
  NANDN U9825 ( .A(n9666), .B(n9875), .Z(n9668) );
  XNOR U9826 ( .A(n322), .B(a[59]), .Z(n9717) );
  NANDN U9827 ( .A(n9874), .B(n9717), .Z(n9667) );
  NAND U9828 ( .A(n9668), .B(n9667), .Z(n9700) );
  NANDN U9829 ( .A(n323), .B(a[55]), .Z(n9711) );
  NANDN U9830 ( .A(n9669), .B(b[21]), .Z(n9670) );
  ANDN U9831 ( .B(n9670), .A(n319), .Z(n9712) );
  XOR U9832 ( .A(n9711), .B(n9712), .Z(n9714) );
  XNOR U9833 ( .A(n9713), .B(n9714), .Z(n9702) );
  XOR U9834 ( .A(n9946), .B(b[25]), .Z(n9708) );
  NANDN U9835 ( .A(n9708), .B(n9706), .Z(n9673) );
  NAND U9836 ( .A(n9707), .B(n9671), .Z(n9672) );
  NAND U9837 ( .A(n9673), .B(n9672), .Z(n9701) );
  XOR U9838 ( .A(n9702), .B(n9701), .Z(n9674) );
  XNOR U9839 ( .A(n9700), .B(n9674), .Z(n9723) );
  NANDN U9840 ( .A(n9675), .B(n9801), .Z(n9677) );
  XNOR U9841 ( .A(a[61]), .B(b[27]), .Z(n9720) );
  OR U9842 ( .A(n9720), .B(n9751), .Z(n9676) );
  NAND U9843 ( .A(n9677), .B(n9676), .Z(n9724) );
  XNOR U9844 ( .A(n9723), .B(n9724), .Z(n9726) );
  XOR U9845 ( .A(n9725), .B(n9726), .Z(n9730) );
  XOR U9846 ( .A(n9729), .B(n9730), .Z(n9731) );
  XNOR U9847 ( .A(n9732), .B(n9731), .Z(n9735) );
  NAND U9848 ( .A(n9679), .B(n9678), .Z(n9683) );
  NANDN U9849 ( .A(n9681), .B(n9680), .Z(n9682) );
  AND U9850 ( .A(n9683), .B(n9682), .Z(n9736) );
  XOR U9851 ( .A(n9735), .B(n9736), .Z(n9738) );
  NANDN U9852 ( .A(n9685), .B(n9684), .Z(n9689) );
  NAND U9853 ( .A(n9687), .B(n9686), .Z(n9688) );
  NAND U9854 ( .A(n9689), .B(n9688), .Z(n9737) );
  XOR U9855 ( .A(n9738), .B(n9737), .Z(n9695) );
  XNOR U9856 ( .A(n9694), .B(n9695), .Z(n9696) );
  XNOR U9857 ( .A(n9697), .B(n9696), .Z(n9692) );
  NANDN U9858 ( .A(n9691), .B(n9690), .Z(n9693) );
  XNOR U9859 ( .A(n9692), .B(n9693), .Z(c[119]) );
  NANDN U9860 ( .A(n9693), .B(n9692), .Z(n9780) );
  NANDN U9861 ( .A(n9695), .B(n9694), .Z(n9699) );
  NANDN U9862 ( .A(n9697), .B(n9696), .Z(n9698) );
  NAND U9863 ( .A(n9699), .B(n9698), .Z(n9744) );
  XNOR U9864 ( .A(b[31]), .B(a[58]), .Z(n9754) );
  OR U9865 ( .A(n9754), .B(n9913), .Z(n9705) );
  NAND U9866 ( .A(n9703), .B(n9914), .Z(n9704) );
  AND U9867 ( .A(n9705), .B(n9704), .Z(n9746) );
  NANDN U9868 ( .A(n320), .B(n9706), .Z(n9710) );
  NANDN U9869 ( .A(n9708), .B(n9707), .Z(n9709) );
  NAND U9870 ( .A(n9710), .B(n9709), .Z(n9745) );
  AND U9871 ( .A(b[31]), .B(a[56]), .Z(n9816) );
  XOR U9872 ( .A(n9745), .B(n9816), .Z(n9747) );
  XOR U9873 ( .A(n9746), .B(n9747), .Z(n9768) );
  XOR U9874 ( .A(n9767), .B(n9768), .Z(n9769) );
  OR U9875 ( .A(n9712), .B(n9711), .Z(n9716) );
  NAND U9876 ( .A(n9714), .B(n9713), .Z(n9715) );
  NAND U9877 ( .A(n9716), .B(n9715), .Z(n9764) );
  NAND U9878 ( .A(n9717), .B(n9875), .Z(n9719) );
  XOR U9879 ( .A(n322), .B(n9805), .Z(n9757) );
  NANDN U9880 ( .A(n9874), .B(n9757), .Z(n9718) );
  NAND U9881 ( .A(n9719), .B(n9718), .Z(n9761) );
  NANDN U9882 ( .A(n9720), .B(n9801), .Z(n9722) );
  XOR U9883 ( .A(b[27]), .B(n9810), .Z(n9750) );
  OR U9884 ( .A(n9750), .B(n9751), .Z(n9721) );
  AND U9885 ( .A(n9722), .B(n9721), .Z(n9762) );
  XNOR U9886 ( .A(n9761), .B(n9762), .Z(n9763) );
  XNOR U9887 ( .A(n9764), .B(n9763), .Z(n9770) );
  XOR U9888 ( .A(n9769), .B(n9770), .Z(n9773) );
  NAND U9889 ( .A(n9724), .B(n9723), .Z(n9728) );
  NANDN U9890 ( .A(n9726), .B(n9725), .Z(n9727) );
  NAND U9891 ( .A(n9728), .B(n9727), .Z(n9774) );
  XNOR U9892 ( .A(n9773), .B(n9774), .Z(n9775) );
  OR U9893 ( .A(n9730), .B(n9729), .Z(n9734) );
  NAND U9894 ( .A(n9732), .B(n9731), .Z(n9733) );
  AND U9895 ( .A(n9734), .B(n9733), .Z(n9776) );
  XNOR U9896 ( .A(n9775), .B(n9776), .Z(n9742) );
  NANDN U9897 ( .A(n9736), .B(n9735), .Z(n9740) );
  OR U9898 ( .A(n9738), .B(n9737), .Z(n9739) );
  AND U9899 ( .A(n9740), .B(n9739), .Z(n9743) );
  XOR U9900 ( .A(n9742), .B(n9743), .Z(n9741) );
  XOR U9901 ( .A(n9744), .B(n9741), .Z(n9779) );
  XNOR U9902 ( .A(n9780), .B(n9779), .Z(c[120]) );
  NANDN U9903 ( .A(n9816), .B(n9745), .Z(n9749) );
  OR U9904 ( .A(n9747), .B(n9746), .Z(n9748) );
  NAND U9905 ( .A(n9749), .B(n9748), .Z(n9792) );
  NANDN U9906 ( .A(n9750), .B(n9801), .Z(n9753) );
  XOR U9907 ( .A(a[63]), .B(n321), .Z(n9802) );
  OR U9908 ( .A(n9802), .B(n9751), .Z(n9752) );
  NAND U9909 ( .A(n9753), .B(n9752), .Z(n9790) );
  NANDN U9910 ( .A(n9754), .B(n9914), .Z(n9756) );
  XNOR U9911 ( .A(n323), .B(a[59]), .Z(n9806) );
  NANDN U9912 ( .A(n9913), .B(n9806), .Z(n9755) );
  NAND U9913 ( .A(n9756), .B(n9755), .Z(n9795) );
  NAND U9914 ( .A(n9875), .B(n9757), .Z(n9759) );
  XNOR U9915 ( .A(n322), .B(a[61]), .Z(n9809) );
  NANDN U9916 ( .A(n9874), .B(n9809), .Z(n9758) );
  AND U9917 ( .A(n9759), .B(n9758), .Z(n9796) );
  XOR U9918 ( .A(n9795), .B(n9796), .Z(n9798) );
  NANDN U9919 ( .A(n323), .B(a[57]), .Z(n9813) );
  NANDN U9920 ( .A(n319), .B(b[24]), .Z(n9760) );
  ANDN U9921 ( .B(n9760), .A(n320), .Z(n9814) );
  XOR U9922 ( .A(n9813), .B(n9814), .Z(n9815) );
  XNOR U9923 ( .A(n9816), .B(n9815), .Z(n9797) );
  XOR U9924 ( .A(n9798), .B(n9797), .Z(n9789) );
  XOR U9925 ( .A(n9790), .B(n9789), .Z(n9791) );
  XNOR U9926 ( .A(n9792), .B(n9791), .Z(n9819) );
  NANDN U9927 ( .A(n9762), .B(n9761), .Z(n9766) );
  NAND U9928 ( .A(n9764), .B(n9763), .Z(n9765) );
  NAND U9929 ( .A(n9766), .B(n9765), .Z(n9820) );
  XOR U9930 ( .A(n9819), .B(n9820), .Z(n9822) );
  NAND U9931 ( .A(n9768), .B(n9767), .Z(n9772) );
  NANDN U9932 ( .A(n9770), .B(n9769), .Z(n9771) );
  NAND U9933 ( .A(n9772), .B(n9771), .Z(n9821) );
  XNOR U9934 ( .A(n9822), .B(n9821), .Z(n9783) );
  NANDN U9935 ( .A(n9774), .B(n9773), .Z(n9778) );
  NAND U9936 ( .A(n9776), .B(n9775), .Z(n9777) );
  NAND U9937 ( .A(n9778), .B(n9777), .Z(n9784) );
  XNOR U9938 ( .A(n9783), .B(n9784), .Z(n9786) );
  XOR U9939 ( .A(n9785), .B(n9786), .Z(n9781) );
  NANDN U9940 ( .A(n9780), .B(n9779), .Z(n9782) );
  XNOR U9941 ( .A(n9781), .B(n9782), .Z(c[121]) );
  NANDN U9942 ( .A(n9782), .B(n9781), .Z(n9827) );
  NANDN U9943 ( .A(n9784), .B(n9783), .Z(n9788) );
  NAND U9944 ( .A(n9786), .B(n9785), .Z(n9787) );
  AND U9945 ( .A(n9788), .B(n9787), .Z(n9830) );
  NAND U9946 ( .A(n9790), .B(n9789), .Z(n9794) );
  NAND U9947 ( .A(n9792), .B(n9791), .Z(n9793) );
  NAND U9948 ( .A(n9794), .B(n9793), .Z(n9852) );
  NANDN U9949 ( .A(n9796), .B(n9795), .Z(n9800) );
  OR U9950 ( .A(n9798), .B(n9797), .Z(n9799) );
  NAND U9951 ( .A(n9800), .B(n9799), .Z(n9851) );
  AND U9952 ( .A(a[58]), .B(b[31]), .Z(n9884) );
  NANDN U9953 ( .A(n9802), .B(n9801), .Z(n9803) );
  NANDN U9954 ( .A(n9804), .B(n9803), .Z(n9839) );
  XNOR U9955 ( .A(n9884), .B(n9839), .Z(n9840) );
  XOR U9956 ( .A(b[31]), .B(n9805), .Z(n9831) );
  OR U9957 ( .A(n9831), .B(n9913), .Z(n9808) );
  NAND U9958 ( .A(n9806), .B(n9914), .Z(n9807) );
  AND U9959 ( .A(n9808), .B(n9807), .Z(n9841) );
  XOR U9960 ( .A(n9840), .B(n9841), .Z(n9847) );
  NAND U9961 ( .A(n9875), .B(n9809), .Z(n9812) );
  XOR U9962 ( .A(n322), .B(n9810), .Z(n9834) );
  NANDN U9963 ( .A(n9874), .B(n9834), .Z(n9811) );
  NAND U9964 ( .A(n9812), .B(n9811), .Z(n9844) );
  OR U9965 ( .A(n9814), .B(n9813), .Z(n9818) );
  NAND U9966 ( .A(n9816), .B(n9815), .Z(n9817) );
  AND U9967 ( .A(n9818), .B(n9817), .Z(n9845) );
  XNOR U9968 ( .A(n9844), .B(n9845), .Z(n9846) );
  XNOR U9969 ( .A(n9847), .B(n9846), .Z(n9850) );
  XNOR U9970 ( .A(n9851), .B(n9850), .Z(n9853) );
  XOR U9971 ( .A(n9852), .B(n9853), .Z(n9828) );
  NANDN U9972 ( .A(n9820), .B(n9819), .Z(n9824) );
  OR U9973 ( .A(n9822), .B(n9821), .Z(n9823) );
  AND U9974 ( .A(n9824), .B(n9823), .Z(n9829) );
  XOR U9975 ( .A(n9828), .B(n9829), .Z(n9825) );
  XOR U9976 ( .A(n9830), .B(n9825), .Z(n9826) );
  XNOR U9977 ( .A(n9827), .B(n9826), .Z(c[122]) );
  NANDN U9978 ( .A(n9827), .B(n9826), .Z(n9889) );
  NANDN U9979 ( .A(n9831), .B(n9914), .Z(n9833) );
  XNOR U9980 ( .A(n323), .B(a[61]), .Z(n9879) );
  NANDN U9981 ( .A(n9913), .B(n9879), .Z(n9832) );
  NAND U9982 ( .A(n9833), .B(n9832), .Z(n9868) );
  NAND U9983 ( .A(n9875), .B(n9834), .Z(n9836) );
  XOR U9984 ( .A(b[29]), .B(n9946), .Z(n9876) );
  OR U9985 ( .A(n9876), .B(n9874), .Z(n9835) );
  AND U9986 ( .A(n9836), .B(n9835), .Z(n9869) );
  XOR U9987 ( .A(n9868), .B(n9869), .Z(n9871) );
  NANDN U9988 ( .A(n323), .B(a[59]), .Z(n9882) );
  NANDN U9989 ( .A(n9837), .B(b[25]), .Z(n9838) );
  ANDN U9990 ( .B(n9838), .A(n321), .Z(n9883) );
  XOR U9991 ( .A(n9882), .B(n9883), .Z(n9885) );
  XNOR U9992 ( .A(n9884), .B(n9885), .Z(n9870) );
  XNOR U9993 ( .A(n9871), .B(n9870), .Z(n9862) );
  NANDN U9994 ( .A(n9839), .B(n9884), .Z(n9843) );
  NAND U9995 ( .A(n9841), .B(n9840), .Z(n9842) );
  AND U9996 ( .A(n9843), .B(n9842), .Z(n9863) );
  XNOR U9997 ( .A(n9862), .B(n9863), .Z(n9864) );
  NANDN U9998 ( .A(n9845), .B(n9844), .Z(n9849) );
  NANDN U9999 ( .A(n9847), .B(n9846), .Z(n9848) );
  AND U10000 ( .A(n9849), .B(n9848), .Z(n9865) );
  XNOR U10001 ( .A(n9864), .B(n9865), .Z(n9857) );
  NAND U10002 ( .A(n9851), .B(n9850), .Z(n9855) );
  NANDN U10003 ( .A(n9853), .B(n9852), .Z(n9854) );
  AND U10004 ( .A(n9855), .B(n9854), .Z(n9856) );
  XNOR U10005 ( .A(n9857), .B(n9856), .Z(n9859) );
  XOR U10006 ( .A(n9858), .B(n9859), .Z(n9888) );
  XOR U10007 ( .A(n9889), .B(n9888), .Z(c[123]) );
  NANDN U10008 ( .A(n9857), .B(n9856), .Z(n9861) );
  NAND U10009 ( .A(n9859), .B(n9858), .Z(n9860) );
  NAND U10010 ( .A(n9861), .B(n9860), .Z(n9894) );
  NANDN U10011 ( .A(n9863), .B(n9862), .Z(n9867) );
  NAND U10012 ( .A(n9865), .B(n9864), .Z(n9866) );
  NAND U10013 ( .A(n9867), .B(n9866), .Z(n9893) );
  NANDN U10014 ( .A(n9869), .B(n9868), .Z(n9873) );
  OR U10015 ( .A(n9871), .B(n9870), .Z(n9872) );
  NAND U10016 ( .A(n9873), .B(n9872), .Z(n9909) );
  NANDN U10017 ( .A(n9874), .B(b[29]), .Z(n9878) );
  NANDN U10018 ( .A(n9876), .B(n9875), .Z(n9877) );
  NAND U10019 ( .A(n9878), .B(n9877), .Z(n9898) );
  AND U10020 ( .A(a[60]), .B(b[31]), .Z(n9919) );
  XOR U10021 ( .A(n9898), .B(n9919), .Z(n9900) );
  NAND U10022 ( .A(n9879), .B(n9914), .Z(n9881) );
  XNOR U10023 ( .A(n323), .B(a[62]), .Z(n9903) );
  NANDN U10024 ( .A(n9913), .B(n9903), .Z(n9880) );
  NAND U10025 ( .A(n9881), .B(n9880), .Z(n9899) );
  XNOR U10026 ( .A(n9900), .B(n9899), .Z(n9906) );
  OR U10027 ( .A(n9883), .B(n9882), .Z(n9887) );
  NAND U10028 ( .A(n9885), .B(n9884), .Z(n9886) );
  AND U10029 ( .A(n9887), .B(n9886), .Z(n9907) );
  XNOR U10030 ( .A(n9906), .B(n9907), .Z(n9908) );
  XOR U10031 ( .A(n9909), .B(n9908), .Z(n9892) );
  XOR U10032 ( .A(n9893), .B(n9892), .Z(n9895) );
  XOR U10033 ( .A(n9894), .B(n9895), .Z(n9890) );
  OR U10034 ( .A(n9889), .B(n9888), .Z(n9891) );
  XNOR U10035 ( .A(n9890), .B(n9891), .Z(c[124]) );
  NANDN U10036 ( .A(n9891), .B(n9890), .Z(n9939) );
  NANDN U10037 ( .A(n9893), .B(n9892), .Z(n9897) );
  OR U10038 ( .A(n9895), .B(n9894), .Z(n9896) );
  AND U10039 ( .A(n9897), .B(n9896), .Z(n9927) );
  NANDN U10040 ( .A(n323), .B(a[61]), .Z(n9918) );
  XNOR U10041 ( .A(n9918), .B(n9917), .Z(n9920) );
  XOR U10042 ( .A(n9919), .B(n9920), .Z(n9933) );
  NANDN U10043 ( .A(n9898), .B(n9919), .Z(n9902) );
  OR U10044 ( .A(n9900), .B(n9899), .Z(n9901) );
  NAND U10045 ( .A(n9902), .B(n9901), .Z(n9932) );
  XOR U10046 ( .A(b[31]), .B(n9946), .Z(n9915) );
  OR U10047 ( .A(n9915), .B(n9913), .Z(n9905) );
  NAND U10048 ( .A(n9903), .B(n9914), .Z(n9904) );
  AND U10049 ( .A(n9905), .B(n9904), .Z(n9931) );
  XOR U10050 ( .A(n9932), .B(n9931), .Z(n9934) );
  XOR U10051 ( .A(n9933), .B(n9934), .Z(n9926) );
  IV U10052 ( .A(n9926), .Z(n9924) );
  NANDN U10053 ( .A(n9907), .B(n9906), .Z(n9911) );
  NAND U10054 ( .A(n9909), .B(n9908), .Z(n9910) );
  AND U10055 ( .A(n9911), .B(n9910), .Z(n9925) );
  XOR U10056 ( .A(n9924), .B(n9925), .Z(n9912) );
  XOR U10057 ( .A(n9927), .B(n9912), .Z(n9938) );
  XNOR U10058 ( .A(n9939), .B(n9938), .Z(c[125]) );
  ANDN U10059 ( .B(b[31]), .A(n9913), .Z(n9948) );
  NANDN U10060 ( .A(n9915), .B(n9914), .Z(n9916) );
  NANDN U10061 ( .A(n9948), .B(n9916), .Z(n9954) );
  OR U10062 ( .A(n9918), .B(n9917), .Z(n9922) );
  NANDN U10063 ( .A(n9920), .B(n9919), .Z(n9921) );
  NAND U10064 ( .A(n9922), .B(n9921), .Z(n9956) );
  AND U10065 ( .A(a[62]), .B(b[31]), .Z(n9953) );
  XNOR U10066 ( .A(n9956), .B(n9953), .Z(n9923) );
  XNOR U10067 ( .A(n9954), .B(n9923), .Z(n9943) );
  NANDN U10068 ( .A(n9924), .B(n9925), .Z(n9930) );
  NOR U10069 ( .A(n9926), .B(n9925), .Z(n9928) );
  NANDN U10070 ( .A(n9928), .B(n9927), .Z(n9929) );
  NAND U10071 ( .A(n9930), .B(n9929), .Z(n9941) );
  NAND U10072 ( .A(n9932), .B(n9931), .Z(n9936) );
  NAND U10073 ( .A(n9934), .B(n9933), .Z(n9935) );
  AND U10074 ( .A(n9936), .B(n9935), .Z(n9942) );
  XNOR U10075 ( .A(n9941), .B(n9942), .Z(n9937) );
  XNOR U10076 ( .A(n9943), .B(n9937), .Z(n9961) );
  NANDN U10077 ( .A(n9939), .B(n9938), .Z(n9962) );
  XNOR U10078 ( .A(n9961), .B(n9962), .Z(c[126]) );
  XNOR U10079 ( .A(n9943), .B(n9942), .Z(n9940) );
  NANDN U10080 ( .A(n9941), .B(n9940), .Z(n9945) );
  NANDN U10081 ( .A(n9943), .B(n9942), .Z(n9944) );
  AND U10082 ( .A(n9945), .B(n9944), .Z(n9952) );
  NANDN U10083 ( .A(b[29]), .B(n323), .Z(n9947) );
  ANDN U10084 ( .B(n9947), .A(n9946), .Z(n9950) );
  OR U10085 ( .A(n9948), .B(b[30]), .Z(n9949) );
  AND U10086 ( .A(n9950), .B(n9949), .Z(n9951) );
  XNOR U10087 ( .A(n9952), .B(n9951), .Z(n9960) );
  NANDN U10088 ( .A(n9953), .B(n9954), .Z(n9958) );
  XNOR U10089 ( .A(n9954), .B(n9953), .Z(n9955) );
  NANDN U10090 ( .A(n9956), .B(n9955), .Z(n9957) );
  AND U10091 ( .A(n9958), .B(n9957), .Z(n9959) );
  XNOR U10092 ( .A(n9960), .B(n9959), .Z(n9964) );
  NANDN U10093 ( .A(n9962), .B(n9961), .Z(n9963) );
  XNOR U10094 ( .A(n9964), .B(n9963), .Z(c[127]) );
endmodule

