
module sum_N1024_CC16 ( clk, rst, a, b, c );
  input [63:0] a;
  input [63:0] b;
  output [63:0] c;
  input clk, rst;
  wire   N130, N131, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952;
  wire   [1:0] carry_on;

  DFF \carry_on_reg[1]  ( .D(N131), .CLK(clk), .RST(rst), .Q(carry_on[1]) );
  DFF \carry_on_reg[0]  ( .D(N130), .CLK(clk), .RST(rst), .Q(carry_on[0]) );
  DFF \rc_reg[63]  ( .D(n256), .CLK(clk), .RST(1'b0), .Q(c[63]) );
  DFF \rc_reg[62]  ( .D(n255), .CLK(clk), .RST(1'b0), .Q(c[62]) );
  DFF \rc_reg[61]  ( .D(n254), .CLK(clk), .RST(1'b0), .Q(c[61]) );
  DFF \rc_reg[60]  ( .D(n253), .CLK(clk), .RST(1'b0), .Q(c[60]) );
  DFF \rc_reg[59]  ( .D(n252), .CLK(clk), .RST(1'b0), .Q(c[59]) );
  DFF \rc_reg[58]  ( .D(n251), .CLK(clk), .RST(1'b0), .Q(c[58]) );
  DFF \rc_reg[57]  ( .D(n250), .CLK(clk), .RST(1'b0), .Q(c[57]) );
  DFF \rc_reg[56]  ( .D(n249), .CLK(clk), .RST(1'b0), .Q(c[56]) );
  DFF \rc_reg[55]  ( .D(n248), .CLK(clk), .RST(1'b0), .Q(c[55]) );
  DFF \rc_reg[54]  ( .D(n247), .CLK(clk), .RST(1'b0), .Q(c[54]) );
  DFF \rc_reg[53]  ( .D(n246), .CLK(clk), .RST(1'b0), .Q(c[53]) );
  DFF \rc_reg[52]  ( .D(n245), .CLK(clk), .RST(1'b0), .Q(c[52]) );
  DFF \rc_reg[51]  ( .D(n244), .CLK(clk), .RST(1'b0), .Q(c[51]) );
  DFF \rc_reg[50]  ( .D(n243), .CLK(clk), .RST(1'b0), .Q(c[50]) );
  DFF \rc_reg[49]  ( .D(n242), .CLK(clk), .RST(1'b0), .Q(c[49]) );
  DFF \rc_reg[48]  ( .D(n241), .CLK(clk), .RST(1'b0), .Q(c[48]) );
  DFF \rc_reg[47]  ( .D(n240), .CLK(clk), .RST(1'b0), .Q(c[47]) );
  DFF \rc_reg[46]  ( .D(n239), .CLK(clk), .RST(1'b0), .Q(c[46]) );
  DFF \rc_reg[45]  ( .D(n238), .CLK(clk), .RST(1'b0), .Q(c[45]) );
  DFF \rc_reg[44]  ( .D(n237), .CLK(clk), .RST(1'b0), .Q(c[44]) );
  DFF \rc_reg[43]  ( .D(n236), .CLK(clk), .RST(1'b0), .Q(c[43]) );
  DFF \rc_reg[42]  ( .D(n235), .CLK(clk), .RST(1'b0), .Q(c[42]) );
  DFF \rc_reg[41]  ( .D(n234), .CLK(clk), .RST(1'b0), .Q(c[41]) );
  DFF \rc_reg[40]  ( .D(n233), .CLK(clk), .RST(1'b0), .Q(c[40]) );
  DFF \rc_reg[39]  ( .D(n232), .CLK(clk), .RST(1'b0), .Q(c[39]) );
  DFF \rc_reg[38]  ( .D(n231), .CLK(clk), .RST(1'b0), .Q(c[38]) );
  DFF \rc_reg[37]  ( .D(n230), .CLK(clk), .RST(1'b0), .Q(c[37]) );
  DFF \rc_reg[36]  ( .D(n229), .CLK(clk), .RST(1'b0), .Q(c[36]) );
  DFF \rc_reg[35]  ( .D(n228), .CLK(clk), .RST(1'b0), .Q(c[35]) );
  DFF \rc_reg[34]  ( .D(n227), .CLK(clk), .RST(1'b0), .Q(c[34]) );
  DFF \rc_reg[33]  ( .D(n226), .CLK(clk), .RST(1'b0), .Q(c[33]) );
  DFF \rc_reg[32]  ( .D(n225), .CLK(clk), .RST(1'b0), .Q(c[32]) );
  DFF \rc_reg[31]  ( .D(n224), .CLK(clk), .RST(1'b0), .Q(c[31]) );
  DFF \rc_reg[30]  ( .D(n223), .CLK(clk), .RST(1'b0), .Q(c[30]) );
  DFF \rc_reg[29]  ( .D(n222), .CLK(clk), .RST(1'b0), .Q(c[29]) );
  DFF \rc_reg[28]  ( .D(n221), .CLK(clk), .RST(1'b0), .Q(c[28]) );
  DFF \rc_reg[27]  ( .D(n220), .CLK(clk), .RST(1'b0), .Q(c[27]) );
  DFF \rc_reg[26]  ( .D(n219), .CLK(clk), .RST(1'b0), .Q(c[26]) );
  DFF \rc_reg[25]  ( .D(n218), .CLK(clk), .RST(1'b0), .Q(c[25]) );
  DFF \rc_reg[24]  ( .D(n217), .CLK(clk), .RST(1'b0), .Q(c[24]) );
  DFF \rc_reg[23]  ( .D(n216), .CLK(clk), .RST(1'b0), .Q(c[23]) );
  DFF \rc_reg[22]  ( .D(n215), .CLK(clk), .RST(1'b0), .Q(c[22]) );
  DFF \rc_reg[21]  ( .D(n214), .CLK(clk), .RST(1'b0), .Q(c[21]) );
  DFF \rc_reg[20]  ( .D(n213), .CLK(clk), .RST(1'b0), .Q(c[20]) );
  DFF \rc_reg[19]  ( .D(n212), .CLK(clk), .RST(1'b0), .Q(c[19]) );
  DFF \rc_reg[18]  ( .D(n211), .CLK(clk), .RST(1'b0), .Q(c[18]) );
  DFF \rc_reg[17]  ( .D(n210), .CLK(clk), .RST(1'b0), .Q(c[17]) );
  DFF \rc_reg[16]  ( .D(n209), .CLK(clk), .RST(1'b0), .Q(c[16]) );
  DFF \rc_reg[15]  ( .D(n208), .CLK(clk), .RST(1'b0), .Q(c[15]) );
  DFF \rc_reg[14]  ( .D(n207), .CLK(clk), .RST(1'b0), .Q(c[14]) );
  DFF \rc_reg[13]  ( .D(n206), .CLK(clk), .RST(1'b0), .Q(c[13]) );
  DFF \rc_reg[12]  ( .D(n205), .CLK(clk), .RST(1'b0), .Q(c[12]) );
  DFF \rc_reg[11]  ( .D(n204), .CLK(clk), .RST(1'b0), .Q(c[11]) );
  DFF \rc_reg[10]  ( .D(n203), .CLK(clk), .RST(1'b0), .Q(c[10]) );
  DFF \rc_reg[9]  ( .D(n202), .CLK(clk), .RST(1'b0), .Q(c[9]) );
  DFF \rc_reg[8]  ( .D(n201), .CLK(clk), .RST(1'b0), .Q(c[8]) );
  DFF \rc_reg[7]  ( .D(n200), .CLK(clk), .RST(1'b0), .Q(c[7]) );
  DFF \rc_reg[6]  ( .D(n199), .CLK(clk), .RST(1'b0), .Q(c[6]) );
  DFF \rc_reg[5]  ( .D(n198), .CLK(clk), .RST(1'b0), .Q(c[5]) );
  DFF \rc_reg[4]  ( .D(n197), .CLK(clk), .RST(1'b0), .Q(c[4]) );
  DFF \rc_reg[3]  ( .D(n196), .CLK(clk), .RST(1'b0), .Q(c[3]) );
  DFF \rc_reg[2]  ( .D(n195), .CLK(clk), .RST(1'b0), .Q(c[2]) );
  DFF \rc_reg[1]  ( .D(n194), .CLK(clk), .RST(1'b0), .Q(c[1]) );
  DFF \rc_reg[0]  ( .D(n193), .CLK(clk), .RST(1'b0), .Q(c[0]) );
  NANDN U259 ( .A(n625), .B(n626), .Z(n257) );
  NANDN U260 ( .A(n939), .B(n938), .Z(n258) );
  AND U261 ( .A(n257), .B(n258), .Z(n259) );
  NAND U262 ( .A(n944), .B(n943), .Z(n260) );
  NANDN U263 ( .A(n259), .B(n627), .Z(n261) );
  AND U264 ( .A(n260), .B(n261), .Z(n628) );
  XOR U265 ( .A(n316), .B(n315), .Z(n678) );
  XOR U266 ( .A(n340), .B(n339), .Z(n698) );
  XOR U267 ( .A(n364), .B(n363), .Z(n718) );
  XOR U268 ( .A(n388), .B(n387), .Z(n738) );
  XOR U269 ( .A(n412), .B(n411), .Z(n758) );
  XOR U270 ( .A(n436), .B(n435), .Z(n778) );
  XOR U271 ( .A(n460), .B(n459), .Z(n798) );
  XOR U272 ( .A(n484), .B(n483), .Z(n818) );
  XOR U273 ( .A(n508), .B(n507), .Z(n838) );
  XOR U274 ( .A(n532), .B(n531), .Z(n858) );
  XOR U275 ( .A(n556), .B(n555), .Z(n878) );
  XOR U276 ( .A(n580), .B(n579), .Z(n898) );
  XOR U277 ( .A(n604), .B(n603), .Z(n918) );
  XOR U278 ( .A(n279), .B(n278), .Z(n648) );
  XOR U279 ( .A(n304), .B(n303), .Z(n668) );
  XOR U280 ( .A(n328), .B(n327), .Z(n688) );
  XOR U281 ( .A(n352), .B(n351), .Z(n708) );
  XOR U282 ( .A(n376), .B(n375), .Z(n728) );
  XOR U283 ( .A(n400), .B(n399), .Z(n748) );
  XOR U284 ( .A(n424), .B(n423), .Z(n768) );
  XOR U285 ( .A(n448), .B(n447), .Z(n788) );
  XOR U286 ( .A(n472), .B(n471), .Z(n808) );
  XOR U287 ( .A(n496), .B(n495), .Z(n828) );
  XOR U288 ( .A(n520), .B(n519), .Z(n848) );
  XOR U289 ( .A(n544), .B(n543), .Z(n868) );
  XOR U290 ( .A(n568), .B(n567), .Z(n888) );
  XOR U291 ( .A(n592), .B(n591), .Z(n908) );
  XOR U292 ( .A(n616), .B(n615), .Z(n928) );
  AND U293 ( .A(b[63]), .B(a[63]), .Z(n633) );
  NAND U294 ( .A(a[61]), .B(b[61]), .Z(n627) );
  AND U295 ( .A(a[60]), .B(b[60]), .Z(n625) );
  XNOR U296 ( .A(a[1]), .B(b[1]), .Z(n264) );
  XNOR U297 ( .A(carry_on[1]), .B(n264), .Z(n639) );
  NAND U298 ( .A(a[0]), .B(b[0]), .Z(n263) );
  XOR U299 ( .A(a[0]), .B(b[0]), .Z(n634) );
  NAND U300 ( .A(n634), .B(carry_on[0]), .Z(n262) );
  NAND U301 ( .A(n263), .B(n262), .Z(n638) );
  NAND U302 ( .A(n639), .B(n638), .Z(n266) );
  ANDN U303 ( .B(carry_on[1]), .A(n264), .Z(n267) );
  ANDN U304 ( .B(n266), .A(n267), .Z(n265) );
  NAND U305 ( .A(a[1]), .B(b[1]), .Z(n268) );
  NAND U306 ( .A(n265), .B(n268), .Z(n272) );
  XNOR U307 ( .A(n268), .B(n266), .Z(n270) );
  NAND U308 ( .A(n268), .B(n267), .Z(n269) );
  NAND U309 ( .A(n270), .B(n269), .Z(n644) );
  XNOR U310 ( .A(a[2]), .B(b[2]), .Z(n643) );
  NAND U311 ( .A(n644), .B(n643), .Z(n271) );
  NAND U312 ( .A(n272), .B(n271), .Z(n278) );
  NAND U313 ( .A(a[2]), .B(b[2]), .Z(n279) );
  AND U314 ( .A(n278), .B(n279), .Z(n274) );
  XOR U315 ( .A(a[3]), .B(b[3]), .Z(n649) );
  ANDN U316 ( .B(n648), .A(n649), .Z(n273) );
  OR U317 ( .A(n274), .B(n273), .Z(n275) );
  AND U318 ( .A(a[3]), .B(b[3]), .Z(n277) );
  ANDN U319 ( .B(n275), .A(n277), .Z(n284) );
  NOR U320 ( .A(n279), .B(n278), .Z(n276) );
  XNOR U321 ( .A(n277), .B(n276), .Z(n282) );
  XOR U322 ( .A(n279), .B(n278), .Z(n280) );
  NAND U323 ( .A(n280), .B(n649), .Z(n281) );
  NAND U324 ( .A(n282), .B(n281), .Z(n654) );
  XNOR U325 ( .A(a[4]), .B(b[4]), .Z(n653) );
  NAND U326 ( .A(n654), .B(n653), .Z(n283) );
  NANDN U327 ( .A(n284), .B(n283), .Z(n291) );
  AND U328 ( .A(a[4]), .B(b[4]), .Z(n285) );
  IV U329 ( .A(n285), .Z(n292) );
  AND U330 ( .A(n291), .B(n292), .Z(n287) );
  XOR U331 ( .A(a[5]), .B(b[5]), .Z(n659) );
  XNOR U332 ( .A(n285), .B(n291), .Z(n658) );
  NANDN U333 ( .A(n659), .B(n658), .Z(n286) );
  NANDN U334 ( .A(n287), .B(n286), .Z(n288) );
  AND U335 ( .A(a[5]), .B(b[5]), .Z(n290) );
  ANDN U336 ( .B(n288), .A(n290), .Z(n297) );
  NOR U337 ( .A(n292), .B(n291), .Z(n289) );
  XNOR U338 ( .A(n290), .B(n289), .Z(n295) );
  XOR U339 ( .A(n292), .B(n291), .Z(n293) );
  NAND U340 ( .A(n293), .B(n659), .Z(n294) );
  NAND U341 ( .A(n295), .B(n294), .Z(n664) );
  XNOR U342 ( .A(a[6]), .B(b[6]), .Z(n663) );
  NAND U343 ( .A(n664), .B(n663), .Z(n296) );
  NANDN U344 ( .A(n297), .B(n296), .Z(n303) );
  NAND U345 ( .A(a[6]), .B(b[6]), .Z(n304) );
  AND U346 ( .A(n303), .B(n304), .Z(n299) );
  XOR U347 ( .A(a[7]), .B(b[7]), .Z(n669) );
  ANDN U348 ( .B(n668), .A(n669), .Z(n298) );
  OR U349 ( .A(n299), .B(n298), .Z(n300) );
  AND U350 ( .A(a[7]), .B(b[7]), .Z(n302) );
  ANDN U351 ( .B(n300), .A(n302), .Z(n309) );
  NOR U352 ( .A(n304), .B(n303), .Z(n301) );
  XNOR U353 ( .A(n302), .B(n301), .Z(n307) );
  XOR U354 ( .A(n304), .B(n303), .Z(n305) );
  NAND U355 ( .A(n305), .B(n669), .Z(n306) );
  NAND U356 ( .A(n307), .B(n306), .Z(n674) );
  XNOR U357 ( .A(a[8]), .B(b[8]), .Z(n673) );
  NAND U358 ( .A(n674), .B(n673), .Z(n308) );
  NANDN U359 ( .A(n309), .B(n308), .Z(n315) );
  NAND U360 ( .A(a[8]), .B(b[8]), .Z(n316) );
  AND U361 ( .A(n315), .B(n316), .Z(n311) );
  XOR U362 ( .A(a[9]), .B(b[9]), .Z(n679) );
  ANDN U363 ( .B(n678), .A(n679), .Z(n310) );
  OR U364 ( .A(n311), .B(n310), .Z(n312) );
  AND U365 ( .A(a[9]), .B(b[9]), .Z(n314) );
  ANDN U366 ( .B(n312), .A(n314), .Z(n321) );
  NOR U367 ( .A(n316), .B(n315), .Z(n313) );
  XNOR U368 ( .A(n314), .B(n313), .Z(n319) );
  XOR U369 ( .A(n316), .B(n315), .Z(n317) );
  NAND U370 ( .A(n317), .B(n679), .Z(n318) );
  NAND U371 ( .A(n319), .B(n318), .Z(n684) );
  XNOR U372 ( .A(a[10]), .B(b[10]), .Z(n683) );
  NAND U373 ( .A(n684), .B(n683), .Z(n320) );
  NANDN U374 ( .A(n321), .B(n320), .Z(n327) );
  NAND U375 ( .A(a[10]), .B(b[10]), .Z(n328) );
  AND U376 ( .A(n327), .B(n328), .Z(n323) );
  XOR U377 ( .A(a[11]), .B(b[11]), .Z(n689) );
  ANDN U378 ( .B(n688), .A(n689), .Z(n322) );
  OR U379 ( .A(n323), .B(n322), .Z(n324) );
  AND U380 ( .A(a[11]), .B(b[11]), .Z(n326) );
  ANDN U381 ( .B(n324), .A(n326), .Z(n333) );
  NOR U382 ( .A(n328), .B(n327), .Z(n325) );
  XNOR U383 ( .A(n326), .B(n325), .Z(n331) );
  XOR U384 ( .A(n328), .B(n327), .Z(n329) );
  NAND U385 ( .A(n329), .B(n689), .Z(n330) );
  NAND U386 ( .A(n331), .B(n330), .Z(n694) );
  XNOR U387 ( .A(a[12]), .B(b[12]), .Z(n693) );
  NAND U388 ( .A(n694), .B(n693), .Z(n332) );
  NANDN U389 ( .A(n333), .B(n332), .Z(n339) );
  NAND U390 ( .A(a[12]), .B(b[12]), .Z(n340) );
  AND U391 ( .A(n339), .B(n340), .Z(n335) );
  XOR U392 ( .A(a[13]), .B(b[13]), .Z(n699) );
  ANDN U393 ( .B(n698), .A(n699), .Z(n334) );
  OR U394 ( .A(n335), .B(n334), .Z(n336) );
  AND U395 ( .A(a[13]), .B(b[13]), .Z(n338) );
  ANDN U396 ( .B(n336), .A(n338), .Z(n345) );
  NOR U397 ( .A(n340), .B(n339), .Z(n337) );
  XNOR U398 ( .A(n338), .B(n337), .Z(n343) );
  XOR U399 ( .A(n340), .B(n339), .Z(n341) );
  NAND U400 ( .A(n341), .B(n699), .Z(n342) );
  NAND U401 ( .A(n343), .B(n342), .Z(n704) );
  XNOR U402 ( .A(a[14]), .B(b[14]), .Z(n703) );
  NAND U403 ( .A(n704), .B(n703), .Z(n344) );
  NANDN U404 ( .A(n345), .B(n344), .Z(n351) );
  NAND U405 ( .A(a[14]), .B(b[14]), .Z(n352) );
  AND U406 ( .A(n351), .B(n352), .Z(n347) );
  XOR U407 ( .A(a[15]), .B(b[15]), .Z(n709) );
  ANDN U408 ( .B(n708), .A(n709), .Z(n346) );
  OR U409 ( .A(n347), .B(n346), .Z(n348) );
  AND U410 ( .A(a[15]), .B(b[15]), .Z(n350) );
  ANDN U411 ( .B(n348), .A(n350), .Z(n357) );
  NOR U412 ( .A(n352), .B(n351), .Z(n349) );
  XNOR U413 ( .A(n350), .B(n349), .Z(n355) );
  XOR U414 ( .A(n352), .B(n351), .Z(n353) );
  NAND U415 ( .A(n353), .B(n709), .Z(n354) );
  NAND U416 ( .A(n355), .B(n354), .Z(n714) );
  XNOR U417 ( .A(a[16]), .B(b[16]), .Z(n713) );
  NAND U418 ( .A(n714), .B(n713), .Z(n356) );
  NANDN U419 ( .A(n357), .B(n356), .Z(n363) );
  NAND U420 ( .A(a[16]), .B(b[16]), .Z(n364) );
  AND U421 ( .A(n363), .B(n364), .Z(n359) );
  XOR U422 ( .A(a[17]), .B(b[17]), .Z(n719) );
  ANDN U423 ( .B(n718), .A(n719), .Z(n358) );
  OR U424 ( .A(n359), .B(n358), .Z(n360) );
  AND U425 ( .A(a[17]), .B(b[17]), .Z(n362) );
  ANDN U426 ( .B(n360), .A(n362), .Z(n369) );
  NOR U427 ( .A(n364), .B(n363), .Z(n361) );
  XNOR U428 ( .A(n362), .B(n361), .Z(n367) );
  XOR U429 ( .A(n364), .B(n363), .Z(n365) );
  NAND U430 ( .A(n365), .B(n719), .Z(n366) );
  NAND U431 ( .A(n367), .B(n366), .Z(n724) );
  XNOR U432 ( .A(a[18]), .B(b[18]), .Z(n723) );
  NAND U433 ( .A(n724), .B(n723), .Z(n368) );
  NANDN U434 ( .A(n369), .B(n368), .Z(n375) );
  NAND U435 ( .A(a[18]), .B(b[18]), .Z(n376) );
  AND U436 ( .A(n375), .B(n376), .Z(n371) );
  XOR U437 ( .A(a[19]), .B(b[19]), .Z(n729) );
  ANDN U438 ( .B(n728), .A(n729), .Z(n370) );
  OR U439 ( .A(n371), .B(n370), .Z(n372) );
  AND U440 ( .A(a[19]), .B(b[19]), .Z(n374) );
  ANDN U441 ( .B(n372), .A(n374), .Z(n381) );
  NOR U442 ( .A(n376), .B(n375), .Z(n373) );
  XNOR U443 ( .A(n374), .B(n373), .Z(n379) );
  XOR U444 ( .A(n376), .B(n375), .Z(n377) );
  NAND U445 ( .A(n377), .B(n729), .Z(n378) );
  NAND U446 ( .A(n379), .B(n378), .Z(n734) );
  XNOR U447 ( .A(a[20]), .B(b[20]), .Z(n733) );
  NAND U448 ( .A(n734), .B(n733), .Z(n380) );
  NANDN U449 ( .A(n381), .B(n380), .Z(n387) );
  NAND U450 ( .A(a[20]), .B(b[20]), .Z(n388) );
  AND U451 ( .A(n387), .B(n388), .Z(n383) );
  XOR U452 ( .A(a[21]), .B(b[21]), .Z(n739) );
  ANDN U453 ( .B(n738), .A(n739), .Z(n382) );
  OR U454 ( .A(n383), .B(n382), .Z(n384) );
  AND U455 ( .A(a[21]), .B(b[21]), .Z(n386) );
  ANDN U456 ( .B(n384), .A(n386), .Z(n393) );
  NOR U457 ( .A(n388), .B(n387), .Z(n385) );
  XNOR U458 ( .A(n386), .B(n385), .Z(n391) );
  XOR U459 ( .A(n388), .B(n387), .Z(n389) );
  NAND U460 ( .A(n389), .B(n739), .Z(n390) );
  NAND U461 ( .A(n391), .B(n390), .Z(n744) );
  XNOR U462 ( .A(a[22]), .B(b[22]), .Z(n743) );
  NAND U463 ( .A(n744), .B(n743), .Z(n392) );
  NANDN U464 ( .A(n393), .B(n392), .Z(n399) );
  NAND U465 ( .A(a[22]), .B(b[22]), .Z(n400) );
  AND U466 ( .A(n399), .B(n400), .Z(n395) );
  XOR U467 ( .A(a[23]), .B(b[23]), .Z(n749) );
  ANDN U468 ( .B(n748), .A(n749), .Z(n394) );
  OR U469 ( .A(n395), .B(n394), .Z(n396) );
  AND U470 ( .A(a[23]), .B(b[23]), .Z(n398) );
  ANDN U471 ( .B(n396), .A(n398), .Z(n405) );
  NOR U472 ( .A(n400), .B(n399), .Z(n397) );
  XNOR U473 ( .A(n398), .B(n397), .Z(n403) );
  XOR U474 ( .A(n400), .B(n399), .Z(n401) );
  NAND U475 ( .A(n401), .B(n749), .Z(n402) );
  NAND U476 ( .A(n403), .B(n402), .Z(n754) );
  XNOR U477 ( .A(a[24]), .B(b[24]), .Z(n753) );
  NAND U478 ( .A(n754), .B(n753), .Z(n404) );
  NANDN U479 ( .A(n405), .B(n404), .Z(n411) );
  NAND U480 ( .A(a[24]), .B(b[24]), .Z(n412) );
  AND U481 ( .A(n411), .B(n412), .Z(n407) );
  XOR U482 ( .A(a[25]), .B(b[25]), .Z(n759) );
  ANDN U483 ( .B(n758), .A(n759), .Z(n406) );
  OR U484 ( .A(n407), .B(n406), .Z(n408) );
  AND U485 ( .A(a[25]), .B(b[25]), .Z(n410) );
  ANDN U486 ( .B(n408), .A(n410), .Z(n417) );
  NOR U487 ( .A(n412), .B(n411), .Z(n409) );
  XNOR U488 ( .A(n410), .B(n409), .Z(n415) );
  XOR U489 ( .A(n412), .B(n411), .Z(n413) );
  NAND U490 ( .A(n413), .B(n759), .Z(n414) );
  NAND U491 ( .A(n415), .B(n414), .Z(n764) );
  XNOR U492 ( .A(a[26]), .B(b[26]), .Z(n763) );
  NAND U493 ( .A(n764), .B(n763), .Z(n416) );
  NANDN U494 ( .A(n417), .B(n416), .Z(n423) );
  NAND U495 ( .A(a[26]), .B(b[26]), .Z(n424) );
  AND U496 ( .A(n423), .B(n424), .Z(n419) );
  XOR U497 ( .A(a[27]), .B(b[27]), .Z(n769) );
  ANDN U498 ( .B(n768), .A(n769), .Z(n418) );
  OR U499 ( .A(n419), .B(n418), .Z(n420) );
  AND U500 ( .A(a[27]), .B(b[27]), .Z(n422) );
  ANDN U501 ( .B(n420), .A(n422), .Z(n429) );
  NOR U502 ( .A(n424), .B(n423), .Z(n421) );
  XNOR U503 ( .A(n422), .B(n421), .Z(n427) );
  XOR U504 ( .A(n424), .B(n423), .Z(n425) );
  NAND U505 ( .A(n425), .B(n769), .Z(n426) );
  NAND U506 ( .A(n427), .B(n426), .Z(n774) );
  XNOR U507 ( .A(a[28]), .B(b[28]), .Z(n773) );
  NAND U508 ( .A(n774), .B(n773), .Z(n428) );
  NANDN U509 ( .A(n429), .B(n428), .Z(n435) );
  NAND U510 ( .A(a[28]), .B(b[28]), .Z(n436) );
  AND U511 ( .A(n435), .B(n436), .Z(n431) );
  XOR U512 ( .A(a[29]), .B(b[29]), .Z(n779) );
  ANDN U513 ( .B(n778), .A(n779), .Z(n430) );
  OR U514 ( .A(n431), .B(n430), .Z(n432) );
  AND U515 ( .A(a[29]), .B(b[29]), .Z(n434) );
  ANDN U516 ( .B(n432), .A(n434), .Z(n441) );
  NOR U517 ( .A(n436), .B(n435), .Z(n433) );
  XNOR U518 ( .A(n434), .B(n433), .Z(n439) );
  XOR U519 ( .A(n436), .B(n435), .Z(n437) );
  NAND U520 ( .A(n437), .B(n779), .Z(n438) );
  NAND U521 ( .A(n439), .B(n438), .Z(n784) );
  XNOR U522 ( .A(a[30]), .B(b[30]), .Z(n783) );
  NAND U523 ( .A(n784), .B(n783), .Z(n440) );
  NANDN U524 ( .A(n441), .B(n440), .Z(n447) );
  NAND U525 ( .A(a[30]), .B(b[30]), .Z(n448) );
  AND U526 ( .A(n447), .B(n448), .Z(n443) );
  XOR U527 ( .A(a[31]), .B(b[31]), .Z(n789) );
  ANDN U528 ( .B(n788), .A(n789), .Z(n442) );
  OR U529 ( .A(n443), .B(n442), .Z(n444) );
  AND U530 ( .A(a[31]), .B(b[31]), .Z(n446) );
  ANDN U531 ( .B(n444), .A(n446), .Z(n453) );
  NOR U532 ( .A(n448), .B(n447), .Z(n445) );
  XNOR U533 ( .A(n446), .B(n445), .Z(n451) );
  XOR U534 ( .A(n448), .B(n447), .Z(n449) );
  NAND U535 ( .A(n449), .B(n789), .Z(n450) );
  NAND U536 ( .A(n451), .B(n450), .Z(n794) );
  XNOR U537 ( .A(a[32]), .B(b[32]), .Z(n793) );
  NAND U538 ( .A(n794), .B(n793), .Z(n452) );
  NANDN U539 ( .A(n453), .B(n452), .Z(n459) );
  NAND U540 ( .A(a[32]), .B(b[32]), .Z(n460) );
  AND U541 ( .A(n459), .B(n460), .Z(n455) );
  XOR U542 ( .A(a[33]), .B(b[33]), .Z(n799) );
  ANDN U543 ( .B(n798), .A(n799), .Z(n454) );
  OR U544 ( .A(n455), .B(n454), .Z(n456) );
  AND U545 ( .A(a[33]), .B(b[33]), .Z(n458) );
  ANDN U546 ( .B(n456), .A(n458), .Z(n465) );
  NOR U547 ( .A(n460), .B(n459), .Z(n457) );
  XNOR U548 ( .A(n458), .B(n457), .Z(n463) );
  XOR U549 ( .A(n460), .B(n459), .Z(n461) );
  NAND U550 ( .A(n461), .B(n799), .Z(n462) );
  NAND U551 ( .A(n463), .B(n462), .Z(n804) );
  XNOR U552 ( .A(a[34]), .B(b[34]), .Z(n803) );
  NAND U553 ( .A(n804), .B(n803), .Z(n464) );
  NANDN U554 ( .A(n465), .B(n464), .Z(n471) );
  NAND U555 ( .A(a[34]), .B(b[34]), .Z(n472) );
  AND U556 ( .A(n471), .B(n472), .Z(n467) );
  XOR U557 ( .A(a[35]), .B(b[35]), .Z(n809) );
  ANDN U558 ( .B(n808), .A(n809), .Z(n466) );
  OR U559 ( .A(n467), .B(n466), .Z(n468) );
  AND U560 ( .A(a[35]), .B(b[35]), .Z(n470) );
  ANDN U561 ( .B(n468), .A(n470), .Z(n477) );
  NOR U562 ( .A(n472), .B(n471), .Z(n469) );
  XNOR U563 ( .A(n470), .B(n469), .Z(n475) );
  XOR U564 ( .A(n472), .B(n471), .Z(n473) );
  NAND U565 ( .A(n473), .B(n809), .Z(n474) );
  NAND U566 ( .A(n475), .B(n474), .Z(n814) );
  XNOR U567 ( .A(a[36]), .B(b[36]), .Z(n813) );
  NAND U568 ( .A(n814), .B(n813), .Z(n476) );
  NANDN U569 ( .A(n477), .B(n476), .Z(n483) );
  NAND U570 ( .A(a[36]), .B(b[36]), .Z(n484) );
  AND U571 ( .A(n483), .B(n484), .Z(n479) );
  XOR U572 ( .A(a[37]), .B(b[37]), .Z(n819) );
  ANDN U573 ( .B(n818), .A(n819), .Z(n478) );
  OR U574 ( .A(n479), .B(n478), .Z(n480) );
  AND U575 ( .A(a[37]), .B(b[37]), .Z(n482) );
  ANDN U576 ( .B(n480), .A(n482), .Z(n489) );
  NOR U577 ( .A(n484), .B(n483), .Z(n481) );
  XNOR U578 ( .A(n482), .B(n481), .Z(n487) );
  XOR U579 ( .A(n484), .B(n483), .Z(n485) );
  NAND U580 ( .A(n485), .B(n819), .Z(n486) );
  NAND U581 ( .A(n487), .B(n486), .Z(n824) );
  XNOR U582 ( .A(a[38]), .B(b[38]), .Z(n823) );
  NAND U583 ( .A(n824), .B(n823), .Z(n488) );
  NANDN U584 ( .A(n489), .B(n488), .Z(n495) );
  NAND U585 ( .A(a[38]), .B(b[38]), .Z(n496) );
  AND U586 ( .A(n495), .B(n496), .Z(n491) );
  XOR U587 ( .A(a[39]), .B(b[39]), .Z(n829) );
  ANDN U588 ( .B(n828), .A(n829), .Z(n490) );
  OR U589 ( .A(n491), .B(n490), .Z(n492) );
  AND U590 ( .A(a[39]), .B(b[39]), .Z(n494) );
  ANDN U591 ( .B(n492), .A(n494), .Z(n501) );
  NOR U592 ( .A(n496), .B(n495), .Z(n493) );
  XNOR U593 ( .A(n494), .B(n493), .Z(n499) );
  XOR U594 ( .A(n496), .B(n495), .Z(n497) );
  NAND U595 ( .A(n497), .B(n829), .Z(n498) );
  NAND U596 ( .A(n499), .B(n498), .Z(n834) );
  XNOR U597 ( .A(a[40]), .B(b[40]), .Z(n833) );
  NAND U598 ( .A(n834), .B(n833), .Z(n500) );
  NANDN U599 ( .A(n501), .B(n500), .Z(n507) );
  NAND U600 ( .A(a[40]), .B(b[40]), .Z(n508) );
  AND U601 ( .A(n507), .B(n508), .Z(n503) );
  XOR U602 ( .A(a[41]), .B(b[41]), .Z(n839) );
  ANDN U603 ( .B(n838), .A(n839), .Z(n502) );
  OR U604 ( .A(n503), .B(n502), .Z(n504) );
  AND U605 ( .A(a[41]), .B(b[41]), .Z(n506) );
  ANDN U606 ( .B(n504), .A(n506), .Z(n513) );
  NOR U607 ( .A(n508), .B(n507), .Z(n505) );
  XNOR U608 ( .A(n506), .B(n505), .Z(n511) );
  XOR U609 ( .A(n508), .B(n507), .Z(n509) );
  NAND U610 ( .A(n509), .B(n839), .Z(n510) );
  NAND U611 ( .A(n511), .B(n510), .Z(n844) );
  XNOR U612 ( .A(a[42]), .B(b[42]), .Z(n843) );
  NAND U613 ( .A(n844), .B(n843), .Z(n512) );
  NANDN U614 ( .A(n513), .B(n512), .Z(n519) );
  NAND U615 ( .A(a[42]), .B(b[42]), .Z(n520) );
  AND U616 ( .A(n519), .B(n520), .Z(n515) );
  XOR U617 ( .A(a[43]), .B(b[43]), .Z(n849) );
  ANDN U618 ( .B(n848), .A(n849), .Z(n514) );
  OR U619 ( .A(n515), .B(n514), .Z(n516) );
  AND U620 ( .A(a[43]), .B(b[43]), .Z(n518) );
  ANDN U621 ( .B(n516), .A(n518), .Z(n525) );
  NOR U622 ( .A(n520), .B(n519), .Z(n517) );
  XNOR U623 ( .A(n518), .B(n517), .Z(n523) );
  XOR U624 ( .A(n520), .B(n519), .Z(n521) );
  NAND U625 ( .A(n521), .B(n849), .Z(n522) );
  NAND U626 ( .A(n523), .B(n522), .Z(n854) );
  XNOR U627 ( .A(a[44]), .B(b[44]), .Z(n853) );
  NAND U628 ( .A(n854), .B(n853), .Z(n524) );
  NANDN U629 ( .A(n525), .B(n524), .Z(n531) );
  NAND U630 ( .A(a[44]), .B(b[44]), .Z(n532) );
  AND U631 ( .A(n531), .B(n532), .Z(n527) );
  XOR U632 ( .A(a[45]), .B(b[45]), .Z(n859) );
  ANDN U633 ( .B(n858), .A(n859), .Z(n526) );
  OR U634 ( .A(n527), .B(n526), .Z(n528) );
  AND U635 ( .A(a[45]), .B(b[45]), .Z(n530) );
  ANDN U636 ( .B(n528), .A(n530), .Z(n537) );
  NOR U637 ( .A(n532), .B(n531), .Z(n529) );
  XNOR U638 ( .A(n530), .B(n529), .Z(n535) );
  XOR U639 ( .A(n532), .B(n531), .Z(n533) );
  NAND U640 ( .A(n533), .B(n859), .Z(n534) );
  NAND U641 ( .A(n535), .B(n534), .Z(n864) );
  XNOR U642 ( .A(a[46]), .B(b[46]), .Z(n863) );
  NAND U643 ( .A(n864), .B(n863), .Z(n536) );
  NANDN U644 ( .A(n537), .B(n536), .Z(n543) );
  NAND U645 ( .A(a[46]), .B(b[46]), .Z(n544) );
  AND U646 ( .A(n543), .B(n544), .Z(n539) );
  XOR U647 ( .A(a[47]), .B(b[47]), .Z(n869) );
  ANDN U648 ( .B(n868), .A(n869), .Z(n538) );
  OR U649 ( .A(n539), .B(n538), .Z(n540) );
  AND U650 ( .A(a[47]), .B(b[47]), .Z(n542) );
  ANDN U651 ( .B(n540), .A(n542), .Z(n549) );
  NOR U652 ( .A(n544), .B(n543), .Z(n541) );
  XNOR U653 ( .A(n542), .B(n541), .Z(n547) );
  XOR U654 ( .A(n544), .B(n543), .Z(n545) );
  NAND U655 ( .A(n545), .B(n869), .Z(n546) );
  NAND U656 ( .A(n547), .B(n546), .Z(n874) );
  XNOR U657 ( .A(a[48]), .B(b[48]), .Z(n873) );
  NAND U658 ( .A(n874), .B(n873), .Z(n548) );
  NANDN U659 ( .A(n549), .B(n548), .Z(n555) );
  NAND U660 ( .A(a[48]), .B(b[48]), .Z(n556) );
  AND U661 ( .A(n555), .B(n556), .Z(n551) );
  XOR U662 ( .A(a[49]), .B(b[49]), .Z(n879) );
  ANDN U663 ( .B(n878), .A(n879), .Z(n550) );
  OR U664 ( .A(n551), .B(n550), .Z(n552) );
  AND U665 ( .A(a[49]), .B(b[49]), .Z(n554) );
  ANDN U666 ( .B(n552), .A(n554), .Z(n561) );
  NOR U667 ( .A(n556), .B(n555), .Z(n553) );
  XNOR U668 ( .A(n554), .B(n553), .Z(n559) );
  XOR U669 ( .A(n556), .B(n555), .Z(n557) );
  NAND U670 ( .A(n557), .B(n879), .Z(n558) );
  NAND U671 ( .A(n559), .B(n558), .Z(n884) );
  XNOR U672 ( .A(a[50]), .B(b[50]), .Z(n883) );
  NAND U673 ( .A(n884), .B(n883), .Z(n560) );
  NANDN U674 ( .A(n561), .B(n560), .Z(n567) );
  NAND U675 ( .A(a[50]), .B(b[50]), .Z(n568) );
  AND U676 ( .A(n567), .B(n568), .Z(n563) );
  XOR U677 ( .A(a[51]), .B(b[51]), .Z(n889) );
  ANDN U678 ( .B(n888), .A(n889), .Z(n562) );
  OR U679 ( .A(n563), .B(n562), .Z(n564) );
  AND U680 ( .A(a[51]), .B(b[51]), .Z(n566) );
  ANDN U681 ( .B(n564), .A(n566), .Z(n573) );
  NOR U682 ( .A(n568), .B(n567), .Z(n565) );
  XNOR U683 ( .A(n566), .B(n565), .Z(n571) );
  XOR U684 ( .A(n568), .B(n567), .Z(n569) );
  NAND U685 ( .A(n569), .B(n889), .Z(n570) );
  NAND U686 ( .A(n571), .B(n570), .Z(n894) );
  XNOR U687 ( .A(a[52]), .B(b[52]), .Z(n893) );
  NAND U688 ( .A(n894), .B(n893), .Z(n572) );
  NANDN U689 ( .A(n573), .B(n572), .Z(n579) );
  NAND U690 ( .A(a[52]), .B(b[52]), .Z(n580) );
  AND U691 ( .A(n579), .B(n580), .Z(n575) );
  XOR U692 ( .A(a[53]), .B(b[53]), .Z(n899) );
  ANDN U693 ( .B(n898), .A(n899), .Z(n574) );
  OR U694 ( .A(n575), .B(n574), .Z(n576) );
  AND U695 ( .A(a[53]), .B(b[53]), .Z(n578) );
  ANDN U696 ( .B(n576), .A(n578), .Z(n585) );
  NOR U697 ( .A(n580), .B(n579), .Z(n577) );
  XNOR U698 ( .A(n578), .B(n577), .Z(n583) );
  XOR U699 ( .A(n580), .B(n579), .Z(n581) );
  NAND U700 ( .A(n581), .B(n899), .Z(n582) );
  NAND U701 ( .A(n583), .B(n582), .Z(n904) );
  XNOR U702 ( .A(a[54]), .B(b[54]), .Z(n903) );
  NAND U703 ( .A(n904), .B(n903), .Z(n584) );
  NANDN U704 ( .A(n585), .B(n584), .Z(n591) );
  NAND U705 ( .A(a[54]), .B(b[54]), .Z(n592) );
  AND U706 ( .A(n591), .B(n592), .Z(n587) );
  XOR U707 ( .A(a[55]), .B(b[55]), .Z(n909) );
  ANDN U708 ( .B(n908), .A(n909), .Z(n586) );
  OR U709 ( .A(n587), .B(n586), .Z(n588) );
  AND U710 ( .A(a[55]), .B(b[55]), .Z(n590) );
  ANDN U711 ( .B(n588), .A(n590), .Z(n597) );
  NOR U712 ( .A(n592), .B(n591), .Z(n589) );
  XNOR U713 ( .A(n590), .B(n589), .Z(n595) );
  XOR U714 ( .A(n592), .B(n591), .Z(n593) );
  NAND U715 ( .A(n593), .B(n909), .Z(n594) );
  NAND U716 ( .A(n595), .B(n594), .Z(n914) );
  XNOR U717 ( .A(a[56]), .B(b[56]), .Z(n913) );
  NAND U718 ( .A(n914), .B(n913), .Z(n596) );
  NANDN U719 ( .A(n597), .B(n596), .Z(n603) );
  NAND U720 ( .A(a[56]), .B(b[56]), .Z(n604) );
  AND U721 ( .A(n603), .B(n604), .Z(n599) );
  XOR U722 ( .A(a[57]), .B(b[57]), .Z(n919) );
  ANDN U723 ( .B(n918), .A(n919), .Z(n598) );
  OR U724 ( .A(n599), .B(n598), .Z(n600) );
  AND U725 ( .A(a[57]), .B(b[57]), .Z(n602) );
  ANDN U726 ( .B(n600), .A(n602), .Z(n609) );
  NOR U727 ( .A(n604), .B(n603), .Z(n601) );
  XNOR U728 ( .A(n602), .B(n601), .Z(n607) );
  XOR U729 ( .A(n604), .B(n603), .Z(n605) );
  NAND U730 ( .A(n605), .B(n919), .Z(n606) );
  NAND U731 ( .A(n607), .B(n606), .Z(n924) );
  XNOR U732 ( .A(a[58]), .B(b[58]), .Z(n923) );
  NAND U733 ( .A(n924), .B(n923), .Z(n608) );
  NANDN U734 ( .A(n609), .B(n608), .Z(n615) );
  NAND U735 ( .A(a[58]), .B(b[58]), .Z(n616) );
  AND U736 ( .A(n615), .B(n616), .Z(n611) );
  XOR U737 ( .A(a[59]), .B(b[59]), .Z(n929) );
  ANDN U738 ( .B(n928), .A(n929), .Z(n610) );
  OR U739 ( .A(n611), .B(n610), .Z(n612) );
  AND U740 ( .A(a[59]), .B(b[59]), .Z(n614) );
  ANDN U741 ( .B(n612), .A(n614), .Z(n621) );
  NOR U742 ( .A(n616), .B(n615), .Z(n613) );
  XNOR U743 ( .A(n614), .B(n613), .Z(n619) );
  XOR U744 ( .A(n616), .B(n615), .Z(n617) );
  NAND U745 ( .A(n617), .B(n929), .Z(n618) );
  NAND U746 ( .A(n619), .B(n618), .Z(n934) );
  XNOR U747 ( .A(a[60]), .B(b[60]), .Z(n933) );
  NAND U748 ( .A(n934), .B(n933), .Z(n620) );
  NANDN U749 ( .A(n621), .B(n620), .Z(n626) );
  ANDN U750 ( .B(n625), .A(n626), .Z(n622) );
  XOR U751 ( .A(n627), .B(n622), .Z(n624) );
  XOR U752 ( .A(a[61]), .B(b[61]), .Z(n939) );
  XNOR U753 ( .A(n625), .B(n626), .Z(n938) );
  NAND U754 ( .A(n939), .B(n938), .Z(n623) );
  NAND U755 ( .A(n624), .B(n623), .Z(n944) );
  XNOR U756 ( .A(a[62]), .B(b[62]), .Z(n943) );
  NAND U757 ( .A(a[62]), .B(b[62]), .Z(n629) );
  ANDN U758 ( .B(n628), .A(n629), .Z(n632) );
  XNOR U759 ( .A(n633), .B(n632), .Z(n631) );
  XNOR U760 ( .A(n629), .B(n628), .Z(n948) );
  XOR U761 ( .A(b[63]), .B(a[63]), .Z(n949) );
  NAND U762 ( .A(n948), .B(n949), .Z(n630) );
  NAND U763 ( .A(n631), .B(n630), .Z(N130) );
  AND U764 ( .A(n633), .B(n632), .Z(N131) );
  NAND U766 ( .A(c[0]), .B(rst), .Z(n637) );
  XOR U767 ( .A(n634), .B(carry_on[0]), .Z(n635) );
  NANDN U768 ( .A(rst), .B(n635), .Z(n636) );
  NAND U769 ( .A(n637), .B(n636), .Z(n193) );
  NAND U770 ( .A(c[1]), .B(rst), .Z(n642) );
  XOR U771 ( .A(n639), .B(n638), .Z(n640) );
  NANDN U772 ( .A(rst), .B(n640), .Z(n641) );
  NAND U773 ( .A(n642), .B(n641), .Z(n194) );
  NAND U774 ( .A(c[2]), .B(rst), .Z(n647) );
  XNOR U775 ( .A(n644), .B(n643), .Z(n645) );
  NANDN U776 ( .A(rst), .B(n645), .Z(n646) );
  NAND U777 ( .A(n647), .B(n646), .Z(n195) );
  NAND U778 ( .A(c[3]), .B(rst), .Z(n652) );
  XOR U779 ( .A(n649), .B(n648), .Z(n650) );
  NANDN U780 ( .A(rst), .B(n650), .Z(n651) );
  NAND U781 ( .A(n652), .B(n651), .Z(n196) );
  NAND U782 ( .A(c[4]), .B(rst), .Z(n657) );
  XNOR U783 ( .A(n654), .B(n653), .Z(n655) );
  NANDN U784 ( .A(rst), .B(n655), .Z(n656) );
  NAND U785 ( .A(n657), .B(n656), .Z(n197) );
  NAND U786 ( .A(c[5]), .B(rst), .Z(n662) );
  XOR U787 ( .A(n659), .B(n658), .Z(n660) );
  NANDN U788 ( .A(rst), .B(n660), .Z(n661) );
  NAND U789 ( .A(n662), .B(n661), .Z(n198) );
  NAND U790 ( .A(c[6]), .B(rst), .Z(n667) );
  XNOR U791 ( .A(n664), .B(n663), .Z(n665) );
  NANDN U792 ( .A(rst), .B(n665), .Z(n666) );
  NAND U793 ( .A(n667), .B(n666), .Z(n199) );
  NAND U794 ( .A(c[7]), .B(rst), .Z(n672) );
  XOR U795 ( .A(n669), .B(n668), .Z(n670) );
  NANDN U796 ( .A(rst), .B(n670), .Z(n671) );
  NAND U797 ( .A(n672), .B(n671), .Z(n200) );
  NAND U798 ( .A(c[8]), .B(rst), .Z(n677) );
  XNOR U799 ( .A(n674), .B(n673), .Z(n675) );
  NANDN U800 ( .A(rst), .B(n675), .Z(n676) );
  NAND U801 ( .A(n677), .B(n676), .Z(n201) );
  NAND U802 ( .A(c[9]), .B(rst), .Z(n682) );
  XOR U803 ( .A(n679), .B(n678), .Z(n680) );
  NANDN U804 ( .A(rst), .B(n680), .Z(n681) );
  NAND U805 ( .A(n682), .B(n681), .Z(n202) );
  NAND U806 ( .A(c[10]), .B(rst), .Z(n687) );
  XNOR U807 ( .A(n684), .B(n683), .Z(n685) );
  NANDN U808 ( .A(rst), .B(n685), .Z(n686) );
  NAND U809 ( .A(n687), .B(n686), .Z(n203) );
  NAND U810 ( .A(c[11]), .B(rst), .Z(n692) );
  XOR U811 ( .A(n689), .B(n688), .Z(n690) );
  NANDN U812 ( .A(rst), .B(n690), .Z(n691) );
  NAND U813 ( .A(n692), .B(n691), .Z(n204) );
  NAND U814 ( .A(c[12]), .B(rst), .Z(n697) );
  XNOR U815 ( .A(n694), .B(n693), .Z(n695) );
  NANDN U816 ( .A(rst), .B(n695), .Z(n696) );
  NAND U817 ( .A(n697), .B(n696), .Z(n205) );
  NAND U818 ( .A(c[13]), .B(rst), .Z(n702) );
  XOR U819 ( .A(n699), .B(n698), .Z(n700) );
  NANDN U820 ( .A(rst), .B(n700), .Z(n701) );
  NAND U821 ( .A(n702), .B(n701), .Z(n206) );
  NAND U822 ( .A(c[14]), .B(rst), .Z(n707) );
  XNOR U823 ( .A(n704), .B(n703), .Z(n705) );
  NANDN U824 ( .A(rst), .B(n705), .Z(n706) );
  NAND U825 ( .A(n707), .B(n706), .Z(n207) );
  NAND U826 ( .A(c[15]), .B(rst), .Z(n712) );
  XOR U827 ( .A(n709), .B(n708), .Z(n710) );
  NANDN U828 ( .A(rst), .B(n710), .Z(n711) );
  NAND U829 ( .A(n712), .B(n711), .Z(n208) );
  NAND U830 ( .A(c[16]), .B(rst), .Z(n717) );
  XNOR U831 ( .A(n714), .B(n713), .Z(n715) );
  NANDN U832 ( .A(rst), .B(n715), .Z(n716) );
  NAND U833 ( .A(n717), .B(n716), .Z(n209) );
  NAND U834 ( .A(c[17]), .B(rst), .Z(n722) );
  XOR U835 ( .A(n719), .B(n718), .Z(n720) );
  NANDN U836 ( .A(rst), .B(n720), .Z(n721) );
  NAND U837 ( .A(n722), .B(n721), .Z(n210) );
  NAND U838 ( .A(c[18]), .B(rst), .Z(n727) );
  XNOR U839 ( .A(n724), .B(n723), .Z(n725) );
  NANDN U840 ( .A(rst), .B(n725), .Z(n726) );
  NAND U841 ( .A(n727), .B(n726), .Z(n211) );
  NAND U842 ( .A(c[19]), .B(rst), .Z(n732) );
  XOR U843 ( .A(n729), .B(n728), .Z(n730) );
  NANDN U844 ( .A(rst), .B(n730), .Z(n731) );
  NAND U845 ( .A(n732), .B(n731), .Z(n212) );
  NAND U846 ( .A(c[20]), .B(rst), .Z(n737) );
  XNOR U847 ( .A(n734), .B(n733), .Z(n735) );
  NANDN U848 ( .A(rst), .B(n735), .Z(n736) );
  NAND U849 ( .A(n737), .B(n736), .Z(n213) );
  NAND U850 ( .A(c[21]), .B(rst), .Z(n742) );
  XOR U851 ( .A(n739), .B(n738), .Z(n740) );
  NANDN U852 ( .A(rst), .B(n740), .Z(n741) );
  NAND U853 ( .A(n742), .B(n741), .Z(n214) );
  NAND U854 ( .A(c[22]), .B(rst), .Z(n747) );
  XNOR U855 ( .A(n744), .B(n743), .Z(n745) );
  NANDN U856 ( .A(rst), .B(n745), .Z(n746) );
  NAND U857 ( .A(n747), .B(n746), .Z(n215) );
  NAND U858 ( .A(c[23]), .B(rst), .Z(n752) );
  XOR U859 ( .A(n749), .B(n748), .Z(n750) );
  NANDN U860 ( .A(rst), .B(n750), .Z(n751) );
  NAND U861 ( .A(n752), .B(n751), .Z(n216) );
  NAND U862 ( .A(c[24]), .B(rst), .Z(n757) );
  XNOR U863 ( .A(n754), .B(n753), .Z(n755) );
  NANDN U864 ( .A(rst), .B(n755), .Z(n756) );
  NAND U865 ( .A(n757), .B(n756), .Z(n217) );
  NAND U866 ( .A(c[25]), .B(rst), .Z(n762) );
  XOR U867 ( .A(n759), .B(n758), .Z(n760) );
  NANDN U868 ( .A(rst), .B(n760), .Z(n761) );
  NAND U869 ( .A(n762), .B(n761), .Z(n218) );
  NAND U870 ( .A(c[26]), .B(rst), .Z(n767) );
  XNOR U871 ( .A(n764), .B(n763), .Z(n765) );
  NANDN U872 ( .A(rst), .B(n765), .Z(n766) );
  NAND U873 ( .A(n767), .B(n766), .Z(n219) );
  NAND U874 ( .A(c[27]), .B(rst), .Z(n772) );
  XOR U875 ( .A(n769), .B(n768), .Z(n770) );
  NANDN U876 ( .A(rst), .B(n770), .Z(n771) );
  NAND U877 ( .A(n772), .B(n771), .Z(n220) );
  NAND U878 ( .A(c[28]), .B(rst), .Z(n777) );
  XNOR U879 ( .A(n774), .B(n773), .Z(n775) );
  NANDN U880 ( .A(rst), .B(n775), .Z(n776) );
  NAND U881 ( .A(n777), .B(n776), .Z(n221) );
  NAND U882 ( .A(c[29]), .B(rst), .Z(n782) );
  XOR U883 ( .A(n779), .B(n778), .Z(n780) );
  NANDN U884 ( .A(rst), .B(n780), .Z(n781) );
  NAND U885 ( .A(n782), .B(n781), .Z(n222) );
  NAND U886 ( .A(c[30]), .B(rst), .Z(n787) );
  XNOR U887 ( .A(n784), .B(n783), .Z(n785) );
  NANDN U888 ( .A(rst), .B(n785), .Z(n786) );
  NAND U889 ( .A(n787), .B(n786), .Z(n223) );
  NAND U890 ( .A(c[31]), .B(rst), .Z(n792) );
  XOR U891 ( .A(n789), .B(n788), .Z(n790) );
  NANDN U892 ( .A(rst), .B(n790), .Z(n791) );
  NAND U893 ( .A(n792), .B(n791), .Z(n224) );
  NAND U894 ( .A(c[32]), .B(rst), .Z(n797) );
  XNOR U895 ( .A(n794), .B(n793), .Z(n795) );
  NANDN U896 ( .A(rst), .B(n795), .Z(n796) );
  NAND U897 ( .A(n797), .B(n796), .Z(n225) );
  NAND U898 ( .A(c[33]), .B(rst), .Z(n802) );
  XOR U899 ( .A(n799), .B(n798), .Z(n800) );
  NANDN U900 ( .A(rst), .B(n800), .Z(n801) );
  NAND U901 ( .A(n802), .B(n801), .Z(n226) );
  NAND U902 ( .A(c[34]), .B(rst), .Z(n807) );
  XNOR U903 ( .A(n804), .B(n803), .Z(n805) );
  NANDN U904 ( .A(rst), .B(n805), .Z(n806) );
  NAND U905 ( .A(n807), .B(n806), .Z(n227) );
  NAND U906 ( .A(c[35]), .B(rst), .Z(n812) );
  XOR U907 ( .A(n809), .B(n808), .Z(n810) );
  NANDN U908 ( .A(rst), .B(n810), .Z(n811) );
  NAND U909 ( .A(n812), .B(n811), .Z(n228) );
  NAND U910 ( .A(c[36]), .B(rst), .Z(n817) );
  XNOR U911 ( .A(n814), .B(n813), .Z(n815) );
  NANDN U912 ( .A(rst), .B(n815), .Z(n816) );
  NAND U913 ( .A(n817), .B(n816), .Z(n229) );
  NAND U914 ( .A(c[37]), .B(rst), .Z(n822) );
  XOR U915 ( .A(n819), .B(n818), .Z(n820) );
  NANDN U916 ( .A(rst), .B(n820), .Z(n821) );
  NAND U917 ( .A(n822), .B(n821), .Z(n230) );
  NAND U918 ( .A(c[38]), .B(rst), .Z(n827) );
  XNOR U919 ( .A(n824), .B(n823), .Z(n825) );
  NANDN U920 ( .A(rst), .B(n825), .Z(n826) );
  NAND U921 ( .A(n827), .B(n826), .Z(n231) );
  NAND U922 ( .A(c[39]), .B(rst), .Z(n832) );
  XOR U923 ( .A(n829), .B(n828), .Z(n830) );
  NANDN U924 ( .A(rst), .B(n830), .Z(n831) );
  NAND U925 ( .A(n832), .B(n831), .Z(n232) );
  NAND U926 ( .A(c[40]), .B(rst), .Z(n837) );
  XNOR U927 ( .A(n834), .B(n833), .Z(n835) );
  NANDN U928 ( .A(rst), .B(n835), .Z(n836) );
  NAND U929 ( .A(n837), .B(n836), .Z(n233) );
  NAND U930 ( .A(c[41]), .B(rst), .Z(n842) );
  XOR U931 ( .A(n839), .B(n838), .Z(n840) );
  NANDN U932 ( .A(rst), .B(n840), .Z(n841) );
  NAND U933 ( .A(n842), .B(n841), .Z(n234) );
  NAND U934 ( .A(c[42]), .B(rst), .Z(n847) );
  XNOR U935 ( .A(n844), .B(n843), .Z(n845) );
  NANDN U936 ( .A(rst), .B(n845), .Z(n846) );
  NAND U937 ( .A(n847), .B(n846), .Z(n235) );
  NAND U938 ( .A(c[43]), .B(rst), .Z(n852) );
  XOR U939 ( .A(n849), .B(n848), .Z(n850) );
  NANDN U940 ( .A(rst), .B(n850), .Z(n851) );
  NAND U941 ( .A(n852), .B(n851), .Z(n236) );
  NAND U942 ( .A(c[44]), .B(rst), .Z(n857) );
  XNOR U943 ( .A(n854), .B(n853), .Z(n855) );
  NANDN U944 ( .A(rst), .B(n855), .Z(n856) );
  NAND U945 ( .A(n857), .B(n856), .Z(n237) );
  NAND U946 ( .A(c[45]), .B(rst), .Z(n862) );
  XOR U947 ( .A(n859), .B(n858), .Z(n860) );
  NANDN U948 ( .A(rst), .B(n860), .Z(n861) );
  NAND U949 ( .A(n862), .B(n861), .Z(n238) );
  NAND U950 ( .A(c[46]), .B(rst), .Z(n867) );
  XNOR U951 ( .A(n864), .B(n863), .Z(n865) );
  NANDN U952 ( .A(rst), .B(n865), .Z(n866) );
  NAND U953 ( .A(n867), .B(n866), .Z(n239) );
  NAND U954 ( .A(c[47]), .B(rst), .Z(n872) );
  XOR U955 ( .A(n869), .B(n868), .Z(n870) );
  NANDN U956 ( .A(rst), .B(n870), .Z(n871) );
  NAND U957 ( .A(n872), .B(n871), .Z(n240) );
  NAND U958 ( .A(c[48]), .B(rst), .Z(n877) );
  XNOR U959 ( .A(n874), .B(n873), .Z(n875) );
  NANDN U960 ( .A(rst), .B(n875), .Z(n876) );
  NAND U961 ( .A(n877), .B(n876), .Z(n241) );
  NAND U962 ( .A(c[49]), .B(rst), .Z(n882) );
  XOR U963 ( .A(n879), .B(n878), .Z(n880) );
  NANDN U964 ( .A(rst), .B(n880), .Z(n881) );
  NAND U965 ( .A(n882), .B(n881), .Z(n242) );
  NAND U966 ( .A(c[50]), .B(rst), .Z(n887) );
  XNOR U967 ( .A(n884), .B(n883), .Z(n885) );
  NANDN U968 ( .A(rst), .B(n885), .Z(n886) );
  NAND U969 ( .A(n887), .B(n886), .Z(n243) );
  NAND U970 ( .A(c[51]), .B(rst), .Z(n892) );
  XOR U971 ( .A(n889), .B(n888), .Z(n890) );
  NANDN U972 ( .A(rst), .B(n890), .Z(n891) );
  NAND U973 ( .A(n892), .B(n891), .Z(n244) );
  NAND U974 ( .A(c[52]), .B(rst), .Z(n897) );
  XNOR U975 ( .A(n894), .B(n893), .Z(n895) );
  NANDN U976 ( .A(rst), .B(n895), .Z(n896) );
  NAND U977 ( .A(n897), .B(n896), .Z(n245) );
  NAND U978 ( .A(c[53]), .B(rst), .Z(n902) );
  XOR U979 ( .A(n899), .B(n898), .Z(n900) );
  NANDN U980 ( .A(rst), .B(n900), .Z(n901) );
  NAND U981 ( .A(n902), .B(n901), .Z(n246) );
  NAND U982 ( .A(c[54]), .B(rst), .Z(n907) );
  XNOR U983 ( .A(n904), .B(n903), .Z(n905) );
  NANDN U984 ( .A(rst), .B(n905), .Z(n906) );
  NAND U985 ( .A(n907), .B(n906), .Z(n247) );
  NAND U986 ( .A(c[55]), .B(rst), .Z(n912) );
  XOR U987 ( .A(n909), .B(n908), .Z(n910) );
  NANDN U988 ( .A(rst), .B(n910), .Z(n911) );
  NAND U989 ( .A(n912), .B(n911), .Z(n248) );
  NAND U990 ( .A(c[56]), .B(rst), .Z(n917) );
  XNOR U991 ( .A(n914), .B(n913), .Z(n915) );
  NANDN U992 ( .A(rst), .B(n915), .Z(n916) );
  NAND U993 ( .A(n917), .B(n916), .Z(n249) );
  NAND U994 ( .A(c[57]), .B(rst), .Z(n922) );
  XOR U995 ( .A(n919), .B(n918), .Z(n920) );
  NANDN U996 ( .A(rst), .B(n920), .Z(n921) );
  NAND U997 ( .A(n922), .B(n921), .Z(n250) );
  NAND U998 ( .A(c[58]), .B(rst), .Z(n927) );
  XNOR U999 ( .A(n924), .B(n923), .Z(n925) );
  NANDN U1000 ( .A(rst), .B(n925), .Z(n926) );
  NAND U1001 ( .A(n927), .B(n926), .Z(n251) );
  NAND U1002 ( .A(c[59]), .B(rst), .Z(n932) );
  XOR U1003 ( .A(n929), .B(n928), .Z(n930) );
  NANDN U1004 ( .A(rst), .B(n930), .Z(n931) );
  NAND U1005 ( .A(n932), .B(n931), .Z(n252) );
  NAND U1006 ( .A(c[60]), .B(rst), .Z(n937) );
  XNOR U1007 ( .A(n934), .B(n933), .Z(n935) );
  NANDN U1008 ( .A(rst), .B(n935), .Z(n936) );
  NAND U1009 ( .A(n937), .B(n936), .Z(n253) );
  NAND U1010 ( .A(c[61]), .B(rst), .Z(n942) );
  XOR U1011 ( .A(n939), .B(n938), .Z(n940) );
  NANDN U1012 ( .A(rst), .B(n940), .Z(n941) );
  NAND U1013 ( .A(n942), .B(n941), .Z(n254) );
  NAND U1014 ( .A(c[62]), .B(rst), .Z(n947) );
  XNOR U1015 ( .A(n944), .B(n943), .Z(n945) );
  NANDN U1016 ( .A(rst), .B(n945), .Z(n946) );
  NAND U1017 ( .A(n947), .B(n946), .Z(n255) );
  NAND U1018 ( .A(c[63]), .B(rst), .Z(n952) );
  XOR U1019 ( .A(n949), .B(n948), .Z(n950) );
  NANDN U1020 ( .A(rst), .B(n950), .Z(n951) );
  NAND U1021 ( .A(n952), .B(n951), .Z(n256) );
endmodule

