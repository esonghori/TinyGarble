
module sum_N1024_CC1 ( clk, rst, a, b, c );
  input [1023:0] a;
  input [1023:0] b;
  output [1023:0] c;
  input clk, rst;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092;

  XOR U2 ( .A(a[1]), .B(b[1]), .Z(n2) );
  NANDN U3 ( .A(n2316), .B(n2), .Z(n3) );
  NAND U4 ( .A(a[1]), .B(b[1]), .Z(n4) );
  AND U5 ( .A(n3), .B(n4), .Z(n2538) );
  XOR U6 ( .A(a[0]), .B(b[0]), .Z(c[0]) );
  XOR U7 ( .A(b[1000]), .B(a[1000]), .Z(n2002) );
  OR U8 ( .A(a[999]), .B(b[999]), .Z(n2000) );
  XOR U9 ( .A(a[999]), .B(b[999]), .Z(n4088) );
  OR U10 ( .A(a[998]), .B(b[998]), .Z(n1998) );
  XOR U11 ( .A(a[998]), .B(b[998]), .Z(n4086) );
  OR U12 ( .A(a[997]), .B(b[997]), .Z(n1996) );
  XOR U13 ( .A(a[997]), .B(b[997]), .Z(n4084) );
  OR U14 ( .A(a[996]), .B(b[996]), .Z(n1994) );
  XOR U15 ( .A(a[996]), .B(b[996]), .Z(n4082) );
  OR U16 ( .A(a[995]), .B(b[995]), .Z(n1992) );
  XOR U17 ( .A(a[995]), .B(b[995]), .Z(n4080) );
  OR U18 ( .A(a[994]), .B(b[994]), .Z(n1990) );
  XOR U19 ( .A(a[994]), .B(b[994]), .Z(n4078) );
  OR U20 ( .A(a[993]), .B(b[993]), .Z(n1988) );
  XOR U21 ( .A(a[993]), .B(b[993]), .Z(n4076) );
  OR U22 ( .A(a[992]), .B(b[992]), .Z(n1986) );
  XOR U23 ( .A(a[992]), .B(b[992]), .Z(n4074) );
  OR U24 ( .A(a[991]), .B(b[991]), .Z(n1984) );
  XOR U25 ( .A(a[991]), .B(b[991]), .Z(n4072) );
  OR U26 ( .A(a[990]), .B(b[990]), .Z(n1982) );
  XOR U27 ( .A(a[990]), .B(b[990]), .Z(n4070) );
  OR U28 ( .A(a[989]), .B(b[989]), .Z(n1980) );
  XOR U29 ( .A(a[989]), .B(b[989]), .Z(n4066) );
  OR U30 ( .A(a[988]), .B(b[988]), .Z(n1978) );
  XOR U31 ( .A(a[988]), .B(b[988]), .Z(n4064) );
  OR U32 ( .A(a[987]), .B(b[987]), .Z(n1976) );
  XOR U33 ( .A(a[987]), .B(b[987]), .Z(n4062) );
  OR U34 ( .A(a[986]), .B(b[986]), .Z(n1974) );
  XOR U35 ( .A(a[986]), .B(b[986]), .Z(n4060) );
  OR U36 ( .A(a[985]), .B(b[985]), .Z(n1972) );
  XOR U37 ( .A(a[985]), .B(b[985]), .Z(n4058) );
  OR U38 ( .A(a[984]), .B(b[984]), .Z(n1970) );
  XOR U39 ( .A(a[984]), .B(b[984]), .Z(n4056) );
  OR U40 ( .A(a[983]), .B(b[983]), .Z(n1968) );
  XOR U41 ( .A(a[983]), .B(b[983]), .Z(n4054) );
  OR U42 ( .A(a[982]), .B(b[982]), .Z(n1966) );
  XOR U43 ( .A(a[982]), .B(b[982]), .Z(n4052) );
  OR U44 ( .A(a[981]), .B(b[981]), .Z(n1964) );
  XOR U45 ( .A(a[981]), .B(b[981]), .Z(n4050) );
  OR U46 ( .A(a[980]), .B(b[980]), .Z(n1962) );
  XOR U47 ( .A(a[980]), .B(b[980]), .Z(n4048) );
  OR U48 ( .A(a[979]), .B(b[979]), .Z(n1960) );
  XOR U49 ( .A(a[979]), .B(b[979]), .Z(n4044) );
  OR U50 ( .A(a[978]), .B(b[978]), .Z(n1958) );
  XOR U51 ( .A(a[978]), .B(b[978]), .Z(n4042) );
  OR U52 ( .A(a[977]), .B(b[977]), .Z(n1956) );
  XOR U53 ( .A(a[977]), .B(b[977]), .Z(n4040) );
  OR U54 ( .A(a[976]), .B(b[976]), .Z(n1954) );
  XOR U55 ( .A(a[976]), .B(b[976]), .Z(n4038) );
  OR U56 ( .A(a[975]), .B(b[975]), .Z(n1952) );
  XOR U57 ( .A(a[975]), .B(b[975]), .Z(n4036) );
  OR U58 ( .A(a[974]), .B(b[974]), .Z(n1950) );
  XOR U59 ( .A(a[974]), .B(b[974]), .Z(n4034) );
  OR U60 ( .A(a[973]), .B(b[973]), .Z(n1948) );
  XOR U61 ( .A(a[973]), .B(b[973]), .Z(n4032) );
  OR U62 ( .A(a[972]), .B(b[972]), .Z(n1946) );
  XOR U63 ( .A(a[972]), .B(b[972]), .Z(n4030) );
  OR U64 ( .A(a[971]), .B(b[971]), .Z(n1944) );
  XOR U65 ( .A(a[971]), .B(b[971]), .Z(n4028) );
  OR U66 ( .A(a[970]), .B(b[970]), .Z(n1942) );
  XOR U67 ( .A(a[970]), .B(b[970]), .Z(n4026) );
  OR U68 ( .A(a[969]), .B(b[969]), .Z(n1940) );
  XOR U69 ( .A(a[969]), .B(b[969]), .Z(n4022) );
  OR U70 ( .A(a[968]), .B(b[968]), .Z(n1938) );
  XOR U71 ( .A(a[968]), .B(b[968]), .Z(n4020) );
  OR U72 ( .A(a[967]), .B(b[967]), .Z(n1936) );
  XOR U73 ( .A(a[967]), .B(b[967]), .Z(n4018) );
  OR U74 ( .A(a[966]), .B(b[966]), .Z(n1934) );
  XOR U75 ( .A(a[966]), .B(b[966]), .Z(n4016) );
  OR U76 ( .A(a[965]), .B(b[965]), .Z(n1932) );
  XOR U77 ( .A(a[965]), .B(b[965]), .Z(n4014) );
  OR U78 ( .A(a[964]), .B(b[964]), .Z(n1930) );
  XOR U79 ( .A(a[964]), .B(b[964]), .Z(n4012) );
  OR U80 ( .A(a[963]), .B(b[963]), .Z(n1928) );
  XOR U81 ( .A(a[963]), .B(b[963]), .Z(n4010) );
  OR U82 ( .A(a[962]), .B(b[962]), .Z(n1926) );
  XOR U83 ( .A(a[962]), .B(b[962]), .Z(n4008) );
  OR U84 ( .A(a[961]), .B(b[961]), .Z(n1924) );
  XOR U85 ( .A(a[961]), .B(b[961]), .Z(n4006) );
  OR U86 ( .A(a[960]), .B(b[960]), .Z(n1922) );
  XOR U87 ( .A(a[960]), .B(b[960]), .Z(n4004) );
  OR U88 ( .A(a[959]), .B(b[959]), .Z(n1920) );
  XOR U89 ( .A(a[959]), .B(b[959]), .Z(n4000) );
  OR U90 ( .A(a[958]), .B(b[958]), .Z(n1918) );
  XOR U91 ( .A(a[958]), .B(b[958]), .Z(n3998) );
  OR U92 ( .A(a[957]), .B(b[957]), .Z(n1916) );
  XOR U93 ( .A(a[957]), .B(b[957]), .Z(n3996) );
  OR U94 ( .A(a[956]), .B(b[956]), .Z(n1914) );
  XOR U95 ( .A(a[956]), .B(b[956]), .Z(n3994) );
  OR U96 ( .A(a[955]), .B(b[955]), .Z(n1912) );
  XOR U97 ( .A(a[955]), .B(b[955]), .Z(n3992) );
  OR U98 ( .A(a[954]), .B(b[954]), .Z(n1910) );
  XOR U99 ( .A(a[954]), .B(b[954]), .Z(n3990) );
  OR U100 ( .A(a[953]), .B(b[953]), .Z(n1908) );
  XOR U101 ( .A(a[953]), .B(b[953]), .Z(n3988) );
  OR U102 ( .A(a[952]), .B(b[952]), .Z(n1906) );
  XOR U103 ( .A(a[952]), .B(b[952]), .Z(n3986) );
  OR U104 ( .A(a[951]), .B(b[951]), .Z(n1904) );
  XOR U105 ( .A(a[951]), .B(b[951]), .Z(n3984) );
  OR U106 ( .A(a[950]), .B(b[950]), .Z(n1902) );
  XOR U107 ( .A(a[950]), .B(b[950]), .Z(n3982) );
  OR U108 ( .A(a[949]), .B(b[949]), .Z(n1900) );
  XOR U109 ( .A(a[949]), .B(b[949]), .Z(n3978) );
  OR U110 ( .A(a[948]), .B(b[948]), .Z(n1898) );
  XOR U111 ( .A(a[948]), .B(b[948]), .Z(n3976) );
  OR U112 ( .A(a[947]), .B(b[947]), .Z(n1896) );
  XOR U113 ( .A(a[947]), .B(b[947]), .Z(n3974) );
  OR U114 ( .A(a[946]), .B(b[946]), .Z(n1894) );
  XOR U115 ( .A(a[946]), .B(b[946]), .Z(n3972) );
  OR U116 ( .A(a[945]), .B(b[945]), .Z(n1892) );
  XOR U117 ( .A(a[945]), .B(b[945]), .Z(n3970) );
  OR U118 ( .A(a[944]), .B(b[944]), .Z(n1890) );
  XOR U119 ( .A(a[944]), .B(b[944]), .Z(n3968) );
  OR U120 ( .A(a[943]), .B(b[943]), .Z(n1888) );
  XOR U121 ( .A(a[943]), .B(b[943]), .Z(n3966) );
  OR U122 ( .A(a[942]), .B(b[942]), .Z(n1886) );
  XOR U123 ( .A(a[942]), .B(b[942]), .Z(n3964) );
  OR U124 ( .A(a[941]), .B(b[941]), .Z(n1884) );
  XOR U125 ( .A(a[941]), .B(b[941]), .Z(n3962) );
  OR U126 ( .A(a[940]), .B(b[940]), .Z(n1882) );
  XOR U127 ( .A(a[940]), .B(b[940]), .Z(n3960) );
  OR U128 ( .A(a[939]), .B(b[939]), .Z(n1880) );
  XOR U129 ( .A(a[939]), .B(b[939]), .Z(n3956) );
  OR U130 ( .A(a[938]), .B(b[938]), .Z(n1878) );
  XOR U131 ( .A(a[938]), .B(b[938]), .Z(n3954) );
  OR U132 ( .A(a[937]), .B(b[937]), .Z(n1876) );
  XOR U133 ( .A(a[937]), .B(b[937]), .Z(n3952) );
  OR U134 ( .A(a[936]), .B(b[936]), .Z(n1874) );
  XOR U135 ( .A(a[936]), .B(b[936]), .Z(n3950) );
  OR U136 ( .A(a[935]), .B(b[935]), .Z(n1872) );
  XOR U137 ( .A(a[935]), .B(b[935]), .Z(n3948) );
  OR U138 ( .A(a[934]), .B(b[934]), .Z(n1870) );
  XOR U139 ( .A(a[934]), .B(b[934]), .Z(n3946) );
  OR U140 ( .A(a[933]), .B(b[933]), .Z(n1868) );
  XOR U141 ( .A(a[933]), .B(b[933]), .Z(n3944) );
  OR U142 ( .A(a[932]), .B(b[932]), .Z(n1866) );
  XOR U143 ( .A(a[932]), .B(b[932]), .Z(n3942) );
  OR U144 ( .A(a[931]), .B(b[931]), .Z(n1864) );
  XOR U145 ( .A(a[931]), .B(b[931]), .Z(n3940) );
  OR U146 ( .A(a[930]), .B(b[930]), .Z(n1862) );
  XOR U147 ( .A(a[930]), .B(b[930]), .Z(n3938) );
  OR U148 ( .A(a[929]), .B(b[929]), .Z(n1860) );
  XOR U149 ( .A(a[929]), .B(b[929]), .Z(n3934) );
  OR U150 ( .A(a[928]), .B(b[928]), .Z(n1858) );
  XOR U151 ( .A(a[928]), .B(b[928]), .Z(n3932) );
  OR U152 ( .A(a[927]), .B(b[927]), .Z(n1856) );
  XOR U153 ( .A(a[927]), .B(b[927]), .Z(n3930) );
  OR U154 ( .A(a[926]), .B(b[926]), .Z(n1854) );
  XOR U155 ( .A(a[926]), .B(b[926]), .Z(n3928) );
  OR U156 ( .A(a[925]), .B(b[925]), .Z(n1852) );
  XOR U157 ( .A(a[925]), .B(b[925]), .Z(n3926) );
  OR U158 ( .A(a[924]), .B(b[924]), .Z(n1850) );
  XOR U159 ( .A(a[924]), .B(b[924]), .Z(n3924) );
  OR U160 ( .A(a[923]), .B(b[923]), .Z(n1848) );
  XOR U161 ( .A(a[923]), .B(b[923]), .Z(n3922) );
  OR U162 ( .A(a[922]), .B(b[922]), .Z(n1846) );
  XOR U163 ( .A(a[922]), .B(b[922]), .Z(n3920) );
  OR U164 ( .A(a[921]), .B(b[921]), .Z(n1844) );
  XOR U165 ( .A(a[921]), .B(b[921]), .Z(n3918) );
  OR U166 ( .A(a[920]), .B(b[920]), .Z(n1842) );
  XOR U167 ( .A(a[920]), .B(b[920]), .Z(n3916) );
  OR U168 ( .A(a[919]), .B(b[919]), .Z(n1840) );
  XOR U169 ( .A(a[919]), .B(b[919]), .Z(n3912) );
  OR U170 ( .A(a[918]), .B(b[918]), .Z(n1838) );
  XOR U171 ( .A(a[918]), .B(b[918]), .Z(n3910) );
  OR U172 ( .A(a[917]), .B(b[917]), .Z(n1836) );
  XOR U173 ( .A(a[917]), .B(b[917]), .Z(n3908) );
  OR U174 ( .A(a[916]), .B(b[916]), .Z(n1834) );
  XOR U175 ( .A(a[916]), .B(b[916]), .Z(n3906) );
  OR U176 ( .A(a[915]), .B(b[915]), .Z(n1832) );
  XOR U177 ( .A(a[915]), .B(b[915]), .Z(n3904) );
  OR U178 ( .A(a[914]), .B(b[914]), .Z(n1830) );
  XOR U179 ( .A(a[914]), .B(b[914]), .Z(n3902) );
  OR U180 ( .A(a[913]), .B(b[913]), .Z(n1828) );
  XOR U181 ( .A(a[913]), .B(b[913]), .Z(n3900) );
  OR U182 ( .A(a[912]), .B(b[912]), .Z(n1826) );
  XOR U183 ( .A(a[912]), .B(b[912]), .Z(n3898) );
  OR U184 ( .A(a[911]), .B(b[911]), .Z(n1824) );
  XOR U185 ( .A(a[911]), .B(b[911]), .Z(n3896) );
  OR U186 ( .A(a[910]), .B(b[910]), .Z(n1822) );
  XOR U187 ( .A(a[910]), .B(b[910]), .Z(n3894) );
  OR U188 ( .A(a[909]), .B(b[909]), .Z(n1820) );
  XOR U189 ( .A(a[909]), .B(b[909]), .Z(n3890) );
  OR U190 ( .A(a[908]), .B(b[908]), .Z(n1818) );
  XOR U191 ( .A(a[908]), .B(b[908]), .Z(n3888) );
  OR U192 ( .A(a[907]), .B(b[907]), .Z(n1816) );
  XOR U193 ( .A(a[907]), .B(b[907]), .Z(n3886) );
  OR U194 ( .A(a[906]), .B(b[906]), .Z(n1814) );
  XOR U195 ( .A(a[906]), .B(b[906]), .Z(n3884) );
  OR U196 ( .A(a[905]), .B(b[905]), .Z(n1812) );
  XOR U197 ( .A(a[905]), .B(b[905]), .Z(n3882) );
  OR U198 ( .A(a[904]), .B(b[904]), .Z(n1810) );
  XOR U199 ( .A(a[904]), .B(b[904]), .Z(n3880) );
  OR U200 ( .A(a[903]), .B(b[903]), .Z(n1808) );
  XOR U201 ( .A(a[903]), .B(b[903]), .Z(n3878) );
  OR U202 ( .A(a[902]), .B(b[902]), .Z(n1806) );
  XOR U203 ( .A(a[902]), .B(b[902]), .Z(n3876) );
  OR U204 ( .A(a[901]), .B(b[901]), .Z(n1804) );
  XOR U205 ( .A(a[901]), .B(b[901]), .Z(n3874) );
  OR U206 ( .A(a[900]), .B(b[900]), .Z(n1802) );
  XOR U207 ( .A(a[900]), .B(b[900]), .Z(n3872) );
  OR U208 ( .A(a[899]), .B(b[899]), .Z(n1800) );
  XOR U209 ( .A(a[899]), .B(b[899]), .Z(n3866) );
  OR U210 ( .A(a[898]), .B(b[898]), .Z(n1798) );
  XOR U211 ( .A(a[898]), .B(b[898]), .Z(n3864) );
  OR U212 ( .A(a[897]), .B(b[897]), .Z(n1796) );
  XOR U213 ( .A(a[897]), .B(b[897]), .Z(n3862) );
  OR U214 ( .A(a[896]), .B(b[896]), .Z(n1794) );
  XOR U215 ( .A(a[896]), .B(b[896]), .Z(n3860) );
  OR U216 ( .A(a[895]), .B(b[895]), .Z(n1792) );
  XOR U217 ( .A(a[895]), .B(b[895]), .Z(n3858) );
  OR U218 ( .A(a[894]), .B(b[894]), .Z(n1790) );
  XOR U219 ( .A(a[894]), .B(b[894]), .Z(n3856) );
  OR U220 ( .A(a[893]), .B(b[893]), .Z(n1788) );
  XOR U221 ( .A(a[893]), .B(b[893]), .Z(n3854) );
  OR U222 ( .A(a[892]), .B(b[892]), .Z(n1786) );
  XOR U223 ( .A(a[892]), .B(b[892]), .Z(n3852) );
  OR U224 ( .A(a[891]), .B(b[891]), .Z(n1784) );
  XOR U225 ( .A(a[891]), .B(b[891]), .Z(n3850) );
  OR U226 ( .A(a[890]), .B(b[890]), .Z(n1782) );
  XOR U227 ( .A(a[890]), .B(b[890]), .Z(n3848) );
  OR U228 ( .A(a[889]), .B(b[889]), .Z(n1780) );
  XOR U229 ( .A(a[889]), .B(b[889]), .Z(n3844) );
  OR U230 ( .A(a[888]), .B(b[888]), .Z(n1778) );
  XOR U231 ( .A(a[888]), .B(b[888]), .Z(n3842) );
  OR U232 ( .A(a[887]), .B(b[887]), .Z(n1776) );
  XOR U233 ( .A(a[887]), .B(b[887]), .Z(n3840) );
  OR U234 ( .A(a[886]), .B(b[886]), .Z(n1774) );
  XOR U235 ( .A(a[886]), .B(b[886]), .Z(n3838) );
  OR U236 ( .A(a[885]), .B(b[885]), .Z(n1772) );
  XOR U237 ( .A(a[885]), .B(b[885]), .Z(n3836) );
  OR U238 ( .A(a[884]), .B(b[884]), .Z(n1770) );
  XOR U239 ( .A(a[884]), .B(b[884]), .Z(n3834) );
  OR U240 ( .A(a[883]), .B(b[883]), .Z(n1768) );
  XOR U241 ( .A(a[883]), .B(b[883]), .Z(n3832) );
  OR U242 ( .A(a[882]), .B(b[882]), .Z(n1766) );
  XOR U243 ( .A(a[882]), .B(b[882]), .Z(n3830) );
  OR U244 ( .A(a[881]), .B(b[881]), .Z(n1764) );
  XOR U245 ( .A(a[881]), .B(b[881]), .Z(n3828) );
  OR U246 ( .A(a[880]), .B(b[880]), .Z(n1762) );
  XOR U247 ( .A(a[880]), .B(b[880]), .Z(n3826) );
  OR U248 ( .A(a[879]), .B(b[879]), .Z(n1760) );
  XOR U249 ( .A(a[879]), .B(b[879]), .Z(n3822) );
  OR U250 ( .A(a[878]), .B(b[878]), .Z(n1758) );
  XOR U251 ( .A(a[878]), .B(b[878]), .Z(n3820) );
  OR U252 ( .A(a[877]), .B(b[877]), .Z(n1756) );
  XOR U253 ( .A(a[877]), .B(b[877]), .Z(n3818) );
  OR U254 ( .A(a[876]), .B(b[876]), .Z(n1754) );
  XOR U255 ( .A(a[876]), .B(b[876]), .Z(n3816) );
  OR U256 ( .A(a[875]), .B(b[875]), .Z(n1752) );
  XOR U257 ( .A(a[875]), .B(b[875]), .Z(n3814) );
  OR U258 ( .A(a[874]), .B(b[874]), .Z(n1750) );
  XOR U259 ( .A(a[874]), .B(b[874]), .Z(n3812) );
  OR U260 ( .A(a[873]), .B(b[873]), .Z(n1748) );
  XOR U261 ( .A(a[873]), .B(b[873]), .Z(n3810) );
  OR U262 ( .A(a[872]), .B(b[872]), .Z(n1746) );
  XOR U263 ( .A(a[872]), .B(b[872]), .Z(n3808) );
  OR U264 ( .A(a[871]), .B(b[871]), .Z(n1744) );
  XOR U265 ( .A(a[871]), .B(b[871]), .Z(n3806) );
  OR U266 ( .A(a[870]), .B(b[870]), .Z(n1742) );
  XOR U267 ( .A(a[870]), .B(b[870]), .Z(n3804) );
  OR U268 ( .A(a[869]), .B(b[869]), .Z(n1740) );
  XOR U269 ( .A(a[869]), .B(b[869]), .Z(n3800) );
  OR U270 ( .A(a[868]), .B(b[868]), .Z(n1738) );
  XOR U271 ( .A(a[868]), .B(b[868]), .Z(n3798) );
  OR U272 ( .A(a[867]), .B(b[867]), .Z(n1736) );
  XOR U273 ( .A(a[867]), .B(b[867]), .Z(n3796) );
  OR U274 ( .A(a[866]), .B(b[866]), .Z(n1734) );
  XOR U275 ( .A(a[866]), .B(b[866]), .Z(n3794) );
  OR U276 ( .A(a[865]), .B(b[865]), .Z(n1732) );
  XOR U277 ( .A(a[865]), .B(b[865]), .Z(n3792) );
  OR U278 ( .A(a[864]), .B(b[864]), .Z(n1730) );
  XOR U279 ( .A(a[864]), .B(b[864]), .Z(n3790) );
  OR U280 ( .A(a[863]), .B(b[863]), .Z(n1728) );
  XOR U281 ( .A(a[863]), .B(b[863]), .Z(n3788) );
  OR U282 ( .A(a[862]), .B(b[862]), .Z(n1726) );
  XOR U283 ( .A(a[862]), .B(b[862]), .Z(n3786) );
  OR U284 ( .A(a[861]), .B(b[861]), .Z(n1724) );
  XOR U285 ( .A(a[861]), .B(b[861]), .Z(n3784) );
  OR U286 ( .A(a[860]), .B(b[860]), .Z(n1722) );
  XOR U287 ( .A(a[860]), .B(b[860]), .Z(n3782) );
  OR U288 ( .A(a[859]), .B(b[859]), .Z(n1720) );
  XOR U289 ( .A(a[859]), .B(b[859]), .Z(n3778) );
  OR U290 ( .A(a[858]), .B(b[858]), .Z(n1718) );
  XOR U291 ( .A(a[858]), .B(b[858]), .Z(n3776) );
  OR U292 ( .A(a[857]), .B(b[857]), .Z(n1716) );
  XOR U293 ( .A(a[857]), .B(b[857]), .Z(n3774) );
  OR U294 ( .A(a[856]), .B(b[856]), .Z(n1714) );
  XOR U295 ( .A(a[856]), .B(b[856]), .Z(n3772) );
  OR U296 ( .A(a[855]), .B(b[855]), .Z(n1712) );
  XOR U297 ( .A(a[855]), .B(b[855]), .Z(n3770) );
  OR U298 ( .A(a[854]), .B(b[854]), .Z(n1710) );
  XOR U299 ( .A(a[854]), .B(b[854]), .Z(n3768) );
  OR U300 ( .A(a[853]), .B(b[853]), .Z(n1708) );
  XOR U301 ( .A(a[853]), .B(b[853]), .Z(n3766) );
  OR U302 ( .A(a[852]), .B(b[852]), .Z(n1706) );
  XOR U303 ( .A(a[852]), .B(b[852]), .Z(n3764) );
  OR U304 ( .A(a[851]), .B(b[851]), .Z(n1704) );
  XOR U305 ( .A(a[851]), .B(b[851]), .Z(n3762) );
  OR U306 ( .A(a[850]), .B(b[850]), .Z(n1702) );
  XOR U307 ( .A(a[850]), .B(b[850]), .Z(n3760) );
  OR U308 ( .A(a[849]), .B(b[849]), .Z(n1700) );
  XOR U309 ( .A(a[849]), .B(b[849]), .Z(n3756) );
  OR U310 ( .A(a[848]), .B(b[848]), .Z(n1698) );
  XOR U311 ( .A(a[848]), .B(b[848]), .Z(n3754) );
  OR U312 ( .A(a[847]), .B(b[847]), .Z(n1696) );
  XOR U313 ( .A(a[847]), .B(b[847]), .Z(n3752) );
  OR U314 ( .A(a[846]), .B(b[846]), .Z(n1694) );
  XOR U315 ( .A(a[846]), .B(b[846]), .Z(n3750) );
  OR U316 ( .A(a[845]), .B(b[845]), .Z(n1692) );
  XOR U317 ( .A(a[845]), .B(b[845]), .Z(n3748) );
  OR U318 ( .A(a[844]), .B(b[844]), .Z(n1690) );
  XOR U319 ( .A(a[844]), .B(b[844]), .Z(n3746) );
  OR U320 ( .A(a[843]), .B(b[843]), .Z(n1688) );
  XOR U321 ( .A(a[843]), .B(b[843]), .Z(n3744) );
  OR U322 ( .A(a[842]), .B(b[842]), .Z(n1686) );
  XOR U323 ( .A(a[842]), .B(b[842]), .Z(n3742) );
  OR U324 ( .A(a[841]), .B(b[841]), .Z(n1684) );
  XOR U325 ( .A(a[841]), .B(b[841]), .Z(n3740) );
  OR U326 ( .A(a[840]), .B(b[840]), .Z(n1682) );
  XOR U327 ( .A(a[840]), .B(b[840]), .Z(n3738) );
  OR U328 ( .A(a[839]), .B(b[839]), .Z(n1680) );
  XOR U329 ( .A(a[839]), .B(b[839]), .Z(n3734) );
  OR U330 ( .A(a[838]), .B(b[838]), .Z(n1678) );
  XOR U331 ( .A(a[838]), .B(b[838]), .Z(n3732) );
  OR U332 ( .A(a[837]), .B(b[837]), .Z(n1676) );
  XOR U333 ( .A(a[837]), .B(b[837]), .Z(n3730) );
  OR U334 ( .A(a[836]), .B(b[836]), .Z(n1674) );
  XOR U335 ( .A(a[836]), .B(b[836]), .Z(n3728) );
  OR U336 ( .A(a[835]), .B(b[835]), .Z(n1672) );
  XOR U337 ( .A(a[835]), .B(b[835]), .Z(n3726) );
  OR U338 ( .A(a[834]), .B(b[834]), .Z(n1670) );
  XOR U339 ( .A(a[834]), .B(b[834]), .Z(n3724) );
  OR U340 ( .A(a[833]), .B(b[833]), .Z(n1668) );
  XOR U341 ( .A(a[833]), .B(b[833]), .Z(n3722) );
  OR U342 ( .A(a[832]), .B(b[832]), .Z(n1666) );
  XOR U343 ( .A(a[832]), .B(b[832]), .Z(n3720) );
  OR U344 ( .A(a[831]), .B(b[831]), .Z(n1664) );
  XOR U345 ( .A(a[831]), .B(b[831]), .Z(n3718) );
  OR U346 ( .A(a[830]), .B(b[830]), .Z(n1662) );
  XOR U347 ( .A(a[830]), .B(b[830]), .Z(n3716) );
  OR U348 ( .A(a[829]), .B(b[829]), .Z(n1660) );
  XOR U349 ( .A(a[829]), .B(b[829]), .Z(n3712) );
  OR U350 ( .A(a[828]), .B(b[828]), .Z(n1658) );
  XOR U351 ( .A(a[828]), .B(b[828]), .Z(n3710) );
  OR U352 ( .A(a[827]), .B(b[827]), .Z(n1656) );
  XOR U353 ( .A(a[827]), .B(b[827]), .Z(n3708) );
  OR U354 ( .A(a[826]), .B(b[826]), .Z(n1654) );
  XOR U355 ( .A(a[826]), .B(b[826]), .Z(n3706) );
  OR U356 ( .A(a[825]), .B(b[825]), .Z(n1652) );
  XOR U357 ( .A(a[825]), .B(b[825]), .Z(n3704) );
  OR U358 ( .A(a[824]), .B(b[824]), .Z(n1650) );
  XOR U359 ( .A(a[824]), .B(b[824]), .Z(n3702) );
  OR U360 ( .A(a[823]), .B(b[823]), .Z(n1648) );
  XOR U361 ( .A(a[823]), .B(b[823]), .Z(n3700) );
  OR U362 ( .A(a[822]), .B(b[822]), .Z(n1646) );
  XOR U363 ( .A(a[822]), .B(b[822]), .Z(n3698) );
  OR U364 ( .A(a[821]), .B(b[821]), .Z(n1644) );
  XOR U365 ( .A(a[821]), .B(b[821]), .Z(n3696) );
  OR U366 ( .A(a[820]), .B(b[820]), .Z(n1642) );
  XOR U367 ( .A(a[820]), .B(b[820]), .Z(n3694) );
  OR U368 ( .A(a[819]), .B(b[819]), .Z(n1640) );
  XOR U369 ( .A(a[819]), .B(b[819]), .Z(n3690) );
  OR U370 ( .A(a[818]), .B(b[818]), .Z(n1638) );
  XOR U371 ( .A(a[818]), .B(b[818]), .Z(n3688) );
  OR U372 ( .A(a[817]), .B(b[817]), .Z(n1636) );
  XOR U373 ( .A(a[817]), .B(b[817]), .Z(n3686) );
  OR U374 ( .A(a[816]), .B(b[816]), .Z(n1634) );
  XOR U375 ( .A(a[816]), .B(b[816]), .Z(n3684) );
  OR U376 ( .A(a[815]), .B(b[815]), .Z(n1632) );
  XOR U377 ( .A(a[815]), .B(b[815]), .Z(n3682) );
  OR U378 ( .A(a[814]), .B(b[814]), .Z(n1630) );
  XOR U379 ( .A(a[814]), .B(b[814]), .Z(n3680) );
  OR U380 ( .A(a[813]), .B(b[813]), .Z(n1628) );
  XOR U381 ( .A(a[813]), .B(b[813]), .Z(n3678) );
  OR U382 ( .A(a[812]), .B(b[812]), .Z(n1626) );
  XOR U383 ( .A(a[812]), .B(b[812]), .Z(n3676) );
  OR U384 ( .A(a[811]), .B(b[811]), .Z(n1624) );
  XOR U385 ( .A(a[811]), .B(b[811]), .Z(n3674) );
  OR U386 ( .A(a[810]), .B(b[810]), .Z(n1622) );
  XOR U387 ( .A(a[810]), .B(b[810]), .Z(n3672) );
  OR U388 ( .A(a[809]), .B(b[809]), .Z(n1620) );
  XOR U389 ( .A(a[809]), .B(b[809]), .Z(n3668) );
  OR U390 ( .A(a[808]), .B(b[808]), .Z(n1618) );
  XOR U391 ( .A(a[808]), .B(b[808]), .Z(n3666) );
  OR U392 ( .A(a[807]), .B(b[807]), .Z(n1616) );
  XOR U393 ( .A(a[807]), .B(b[807]), .Z(n3664) );
  OR U394 ( .A(a[806]), .B(b[806]), .Z(n1614) );
  XOR U395 ( .A(a[806]), .B(b[806]), .Z(n3662) );
  OR U396 ( .A(a[805]), .B(b[805]), .Z(n1612) );
  XOR U397 ( .A(a[805]), .B(b[805]), .Z(n3660) );
  OR U398 ( .A(a[804]), .B(b[804]), .Z(n1610) );
  XOR U399 ( .A(a[804]), .B(b[804]), .Z(n3658) );
  OR U400 ( .A(a[803]), .B(b[803]), .Z(n1608) );
  XOR U401 ( .A(a[803]), .B(b[803]), .Z(n3656) );
  OR U402 ( .A(a[802]), .B(b[802]), .Z(n1606) );
  XOR U403 ( .A(a[802]), .B(b[802]), .Z(n3654) );
  OR U404 ( .A(a[801]), .B(b[801]), .Z(n1604) );
  XOR U405 ( .A(a[801]), .B(b[801]), .Z(n3652) );
  OR U406 ( .A(a[800]), .B(b[800]), .Z(n1602) );
  XOR U407 ( .A(a[800]), .B(b[800]), .Z(n3650) );
  OR U408 ( .A(a[799]), .B(b[799]), .Z(n1600) );
  XOR U409 ( .A(a[799]), .B(b[799]), .Z(n3644) );
  OR U410 ( .A(a[798]), .B(b[798]), .Z(n1598) );
  XOR U411 ( .A(a[798]), .B(b[798]), .Z(n3642) );
  OR U412 ( .A(a[797]), .B(b[797]), .Z(n1596) );
  XOR U413 ( .A(a[797]), .B(b[797]), .Z(n3640) );
  OR U414 ( .A(a[796]), .B(b[796]), .Z(n1594) );
  XOR U415 ( .A(a[796]), .B(b[796]), .Z(n3638) );
  OR U416 ( .A(a[795]), .B(b[795]), .Z(n1592) );
  XOR U417 ( .A(a[795]), .B(b[795]), .Z(n3636) );
  OR U418 ( .A(a[794]), .B(b[794]), .Z(n1590) );
  XOR U419 ( .A(a[794]), .B(b[794]), .Z(n3634) );
  OR U420 ( .A(a[793]), .B(b[793]), .Z(n1588) );
  XOR U421 ( .A(a[793]), .B(b[793]), .Z(n3632) );
  OR U422 ( .A(a[792]), .B(b[792]), .Z(n1586) );
  XOR U423 ( .A(a[792]), .B(b[792]), .Z(n3630) );
  OR U424 ( .A(a[791]), .B(b[791]), .Z(n1584) );
  XOR U425 ( .A(a[791]), .B(b[791]), .Z(n3628) );
  OR U426 ( .A(a[790]), .B(b[790]), .Z(n1582) );
  XOR U427 ( .A(a[790]), .B(b[790]), .Z(n3626) );
  OR U428 ( .A(a[789]), .B(b[789]), .Z(n1580) );
  XOR U429 ( .A(a[789]), .B(b[789]), .Z(n3622) );
  OR U430 ( .A(a[788]), .B(b[788]), .Z(n1578) );
  XOR U431 ( .A(a[788]), .B(b[788]), .Z(n3620) );
  OR U432 ( .A(a[787]), .B(b[787]), .Z(n1576) );
  XOR U433 ( .A(a[787]), .B(b[787]), .Z(n3618) );
  OR U434 ( .A(a[786]), .B(b[786]), .Z(n1574) );
  XOR U435 ( .A(a[786]), .B(b[786]), .Z(n3616) );
  OR U436 ( .A(a[785]), .B(b[785]), .Z(n1572) );
  XOR U437 ( .A(a[785]), .B(b[785]), .Z(n3614) );
  OR U438 ( .A(a[784]), .B(b[784]), .Z(n1570) );
  XOR U439 ( .A(a[784]), .B(b[784]), .Z(n3612) );
  OR U440 ( .A(a[783]), .B(b[783]), .Z(n1568) );
  XOR U441 ( .A(a[783]), .B(b[783]), .Z(n3610) );
  OR U442 ( .A(a[782]), .B(b[782]), .Z(n1566) );
  XOR U443 ( .A(a[782]), .B(b[782]), .Z(n3608) );
  OR U444 ( .A(a[781]), .B(b[781]), .Z(n1564) );
  XOR U445 ( .A(a[781]), .B(b[781]), .Z(n3606) );
  OR U446 ( .A(a[780]), .B(b[780]), .Z(n1562) );
  XOR U447 ( .A(a[780]), .B(b[780]), .Z(n3604) );
  OR U448 ( .A(a[779]), .B(b[779]), .Z(n1560) );
  XOR U449 ( .A(a[779]), .B(b[779]), .Z(n3600) );
  OR U450 ( .A(a[778]), .B(b[778]), .Z(n1558) );
  XOR U451 ( .A(a[778]), .B(b[778]), .Z(n3598) );
  OR U452 ( .A(a[777]), .B(b[777]), .Z(n1556) );
  XOR U453 ( .A(a[777]), .B(b[777]), .Z(n3596) );
  OR U454 ( .A(a[776]), .B(b[776]), .Z(n1554) );
  XOR U455 ( .A(a[776]), .B(b[776]), .Z(n3594) );
  OR U456 ( .A(a[775]), .B(b[775]), .Z(n1552) );
  XOR U457 ( .A(a[775]), .B(b[775]), .Z(n3592) );
  OR U458 ( .A(a[774]), .B(b[774]), .Z(n1550) );
  XOR U459 ( .A(a[774]), .B(b[774]), .Z(n3590) );
  OR U460 ( .A(a[773]), .B(b[773]), .Z(n1548) );
  XOR U461 ( .A(a[773]), .B(b[773]), .Z(n3588) );
  OR U462 ( .A(a[772]), .B(b[772]), .Z(n1546) );
  XOR U463 ( .A(a[772]), .B(b[772]), .Z(n3586) );
  OR U464 ( .A(a[771]), .B(b[771]), .Z(n1544) );
  XOR U465 ( .A(a[771]), .B(b[771]), .Z(n3584) );
  OR U466 ( .A(a[770]), .B(b[770]), .Z(n1542) );
  XOR U467 ( .A(a[770]), .B(b[770]), .Z(n3582) );
  OR U468 ( .A(a[769]), .B(b[769]), .Z(n1540) );
  XOR U469 ( .A(a[769]), .B(b[769]), .Z(n3578) );
  OR U470 ( .A(a[768]), .B(b[768]), .Z(n1538) );
  XOR U471 ( .A(a[768]), .B(b[768]), .Z(n3576) );
  OR U472 ( .A(a[767]), .B(b[767]), .Z(n1536) );
  XOR U473 ( .A(a[767]), .B(b[767]), .Z(n3574) );
  OR U474 ( .A(a[766]), .B(b[766]), .Z(n1534) );
  XOR U475 ( .A(a[766]), .B(b[766]), .Z(n3572) );
  OR U476 ( .A(a[765]), .B(b[765]), .Z(n1532) );
  XOR U477 ( .A(a[765]), .B(b[765]), .Z(n3570) );
  OR U478 ( .A(a[764]), .B(b[764]), .Z(n1530) );
  XOR U479 ( .A(a[764]), .B(b[764]), .Z(n3568) );
  OR U480 ( .A(a[763]), .B(b[763]), .Z(n1528) );
  XOR U481 ( .A(a[763]), .B(b[763]), .Z(n3566) );
  OR U482 ( .A(a[762]), .B(b[762]), .Z(n1526) );
  XOR U483 ( .A(a[762]), .B(b[762]), .Z(n3564) );
  OR U484 ( .A(a[761]), .B(b[761]), .Z(n1524) );
  XOR U485 ( .A(a[761]), .B(b[761]), .Z(n3562) );
  OR U486 ( .A(a[760]), .B(b[760]), .Z(n1522) );
  XOR U487 ( .A(a[760]), .B(b[760]), .Z(n3560) );
  OR U488 ( .A(a[759]), .B(b[759]), .Z(n1520) );
  XOR U489 ( .A(a[759]), .B(b[759]), .Z(n3556) );
  OR U490 ( .A(a[758]), .B(b[758]), .Z(n1518) );
  XOR U491 ( .A(a[758]), .B(b[758]), .Z(n3554) );
  OR U492 ( .A(a[757]), .B(b[757]), .Z(n1516) );
  XOR U493 ( .A(a[757]), .B(b[757]), .Z(n3552) );
  OR U494 ( .A(a[756]), .B(b[756]), .Z(n1514) );
  XOR U495 ( .A(a[756]), .B(b[756]), .Z(n3550) );
  OR U496 ( .A(a[755]), .B(b[755]), .Z(n1512) );
  XOR U497 ( .A(a[755]), .B(b[755]), .Z(n3548) );
  OR U498 ( .A(a[754]), .B(b[754]), .Z(n1510) );
  XOR U499 ( .A(a[754]), .B(b[754]), .Z(n3546) );
  OR U500 ( .A(a[753]), .B(b[753]), .Z(n1508) );
  XOR U501 ( .A(a[753]), .B(b[753]), .Z(n3544) );
  OR U502 ( .A(a[752]), .B(b[752]), .Z(n1506) );
  XOR U503 ( .A(a[752]), .B(b[752]), .Z(n3542) );
  OR U504 ( .A(a[751]), .B(b[751]), .Z(n1504) );
  XOR U505 ( .A(a[751]), .B(b[751]), .Z(n3540) );
  OR U506 ( .A(a[750]), .B(b[750]), .Z(n1502) );
  XOR U507 ( .A(a[750]), .B(b[750]), .Z(n3538) );
  OR U508 ( .A(a[749]), .B(b[749]), .Z(n1500) );
  XOR U509 ( .A(a[749]), .B(b[749]), .Z(n3534) );
  OR U510 ( .A(a[748]), .B(b[748]), .Z(n1498) );
  XOR U511 ( .A(a[748]), .B(b[748]), .Z(n3532) );
  OR U512 ( .A(a[747]), .B(b[747]), .Z(n1496) );
  XOR U513 ( .A(a[747]), .B(b[747]), .Z(n3530) );
  OR U514 ( .A(a[746]), .B(b[746]), .Z(n1494) );
  XOR U515 ( .A(a[746]), .B(b[746]), .Z(n3528) );
  OR U516 ( .A(a[745]), .B(b[745]), .Z(n1492) );
  XOR U517 ( .A(a[745]), .B(b[745]), .Z(n3526) );
  OR U518 ( .A(a[744]), .B(b[744]), .Z(n1490) );
  XOR U519 ( .A(a[744]), .B(b[744]), .Z(n3524) );
  OR U520 ( .A(a[743]), .B(b[743]), .Z(n1488) );
  XOR U521 ( .A(a[743]), .B(b[743]), .Z(n3522) );
  OR U522 ( .A(a[742]), .B(b[742]), .Z(n1486) );
  XOR U523 ( .A(a[742]), .B(b[742]), .Z(n3520) );
  OR U524 ( .A(a[741]), .B(b[741]), .Z(n1484) );
  XOR U525 ( .A(a[741]), .B(b[741]), .Z(n3518) );
  OR U526 ( .A(a[740]), .B(b[740]), .Z(n1482) );
  XOR U527 ( .A(a[740]), .B(b[740]), .Z(n3516) );
  OR U528 ( .A(a[739]), .B(b[739]), .Z(n1480) );
  XOR U529 ( .A(a[739]), .B(b[739]), .Z(n3512) );
  OR U530 ( .A(a[738]), .B(b[738]), .Z(n1478) );
  XOR U531 ( .A(a[738]), .B(b[738]), .Z(n3510) );
  OR U532 ( .A(a[737]), .B(b[737]), .Z(n1476) );
  XOR U533 ( .A(a[737]), .B(b[737]), .Z(n3508) );
  OR U534 ( .A(a[736]), .B(b[736]), .Z(n1474) );
  XOR U535 ( .A(a[736]), .B(b[736]), .Z(n3506) );
  OR U536 ( .A(a[735]), .B(b[735]), .Z(n1472) );
  XOR U537 ( .A(a[735]), .B(b[735]), .Z(n3504) );
  OR U538 ( .A(a[734]), .B(b[734]), .Z(n1470) );
  XOR U539 ( .A(a[734]), .B(b[734]), .Z(n3502) );
  OR U540 ( .A(a[733]), .B(b[733]), .Z(n1468) );
  XOR U541 ( .A(a[733]), .B(b[733]), .Z(n3500) );
  OR U542 ( .A(a[732]), .B(b[732]), .Z(n1466) );
  XOR U543 ( .A(a[732]), .B(b[732]), .Z(n3498) );
  OR U544 ( .A(a[731]), .B(b[731]), .Z(n1464) );
  XOR U545 ( .A(a[731]), .B(b[731]), .Z(n3496) );
  OR U546 ( .A(a[730]), .B(b[730]), .Z(n1462) );
  XOR U547 ( .A(a[730]), .B(b[730]), .Z(n3494) );
  OR U548 ( .A(a[729]), .B(b[729]), .Z(n1460) );
  XOR U549 ( .A(a[729]), .B(b[729]), .Z(n3490) );
  OR U550 ( .A(a[728]), .B(b[728]), .Z(n1458) );
  XOR U551 ( .A(a[728]), .B(b[728]), .Z(n3488) );
  OR U552 ( .A(a[727]), .B(b[727]), .Z(n1456) );
  XOR U553 ( .A(a[727]), .B(b[727]), .Z(n3486) );
  OR U554 ( .A(a[726]), .B(b[726]), .Z(n1454) );
  XOR U555 ( .A(a[726]), .B(b[726]), .Z(n3484) );
  OR U556 ( .A(a[725]), .B(b[725]), .Z(n1452) );
  XOR U557 ( .A(a[725]), .B(b[725]), .Z(n3482) );
  OR U558 ( .A(a[724]), .B(b[724]), .Z(n1450) );
  XOR U559 ( .A(a[724]), .B(b[724]), .Z(n3480) );
  OR U560 ( .A(a[723]), .B(b[723]), .Z(n1448) );
  XOR U561 ( .A(a[723]), .B(b[723]), .Z(n3478) );
  OR U562 ( .A(a[722]), .B(b[722]), .Z(n1446) );
  XOR U563 ( .A(a[722]), .B(b[722]), .Z(n3476) );
  OR U564 ( .A(a[721]), .B(b[721]), .Z(n1444) );
  XOR U565 ( .A(a[721]), .B(b[721]), .Z(n3474) );
  OR U566 ( .A(a[720]), .B(b[720]), .Z(n1442) );
  XOR U567 ( .A(a[720]), .B(b[720]), .Z(n3472) );
  OR U568 ( .A(a[719]), .B(b[719]), .Z(n1440) );
  XOR U569 ( .A(a[719]), .B(b[719]), .Z(n3468) );
  OR U570 ( .A(a[718]), .B(b[718]), .Z(n1438) );
  XOR U571 ( .A(a[718]), .B(b[718]), .Z(n3466) );
  OR U572 ( .A(a[717]), .B(b[717]), .Z(n1436) );
  XOR U573 ( .A(a[717]), .B(b[717]), .Z(n3464) );
  OR U574 ( .A(a[716]), .B(b[716]), .Z(n1434) );
  XOR U575 ( .A(a[716]), .B(b[716]), .Z(n3462) );
  OR U576 ( .A(a[715]), .B(b[715]), .Z(n1432) );
  XOR U577 ( .A(a[715]), .B(b[715]), .Z(n3460) );
  OR U578 ( .A(a[714]), .B(b[714]), .Z(n1430) );
  XOR U579 ( .A(a[714]), .B(b[714]), .Z(n3458) );
  OR U580 ( .A(a[713]), .B(b[713]), .Z(n1428) );
  XOR U581 ( .A(a[713]), .B(b[713]), .Z(n3456) );
  OR U582 ( .A(a[712]), .B(b[712]), .Z(n1426) );
  XOR U583 ( .A(a[712]), .B(b[712]), .Z(n3454) );
  OR U584 ( .A(a[711]), .B(b[711]), .Z(n1424) );
  XOR U585 ( .A(a[711]), .B(b[711]), .Z(n3452) );
  OR U586 ( .A(a[710]), .B(b[710]), .Z(n1422) );
  XOR U587 ( .A(a[710]), .B(b[710]), .Z(n3450) );
  OR U588 ( .A(a[709]), .B(b[709]), .Z(n1420) );
  XOR U589 ( .A(a[709]), .B(b[709]), .Z(n3446) );
  OR U590 ( .A(a[708]), .B(b[708]), .Z(n1418) );
  XOR U591 ( .A(a[708]), .B(b[708]), .Z(n3444) );
  OR U592 ( .A(a[707]), .B(b[707]), .Z(n1416) );
  XOR U593 ( .A(a[707]), .B(b[707]), .Z(n3442) );
  OR U594 ( .A(a[706]), .B(b[706]), .Z(n1414) );
  XOR U595 ( .A(a[706]), .B(b[706]), .Z(n3440) );
  OR U596 ( .A(a[705]), .B(b[705]), .Z(n1412) );
  XOR U597 ( .A(a[705]), .B(b[705]), .Z(n3438) );
  OR U598 ( .A(a[704]), .B(b[704]), .Z(n1410) );
  XOR U599 ( .A(a[704]), .B(b[704]), .Z(n3436) );
  OR U600 ( .A(a[703]), .B(b[703]), .Z(n1408) );
  XOR U601 ( .A(a[703]), .B(b[703]), .Z(n3434) );
  OR U602 ( .A(a[702]), .B(b[702]), .Z(n1406) );
  XOR U603 ( .A(a[702]), .B(b[702]), .Z(n3432) );
  OR U604 ( .A(a[701]), .B(b[701]), .Z(n1404) );
  XOR U605 ( .A(a[701]), .B(b[701]), .Z(n3430) );
  OR U606 ( .A(a[700]), .B(b[700]), .Z(n1402) );
  XOR U607 ( .A(a[700]), .B(b[700]), .Z(n3428) );
  OR U608 ( .A(a[699]), .B(b[699]), .Z(n1400) );
  XOR U609 ( .A(a[699]), .B(b[699]), .Z(n3422) );
  OR U610 ( .A(a[698]), .B(b[698]), .Z(n1398) );
  XOR U611 ( .A(a[698]), .B(b[698]), .Z(n3420) );
  OR U612 ( .A(a[697]), .B(b[697]), .Z(n1396) );
  XOR U613 ( .A(a[697]), .B(b[697]), .Z(n3418) );
  OR U614 ( .A(a[696]), .B(b[696]), .Z(n1394) );
  XOR U615 ( .A(a[696]), .B(b[696]), .Z(n3416) );
  OR U616 ( .A(a[695]), .B(b[695]), .Z(n1392) );
  XOR U617 ( .A(a[695]), .B(b[695]), .Z(n3414) );
  OR U618 ( .A(a[694]), .B(b[694]), .Z(n1390) );
  XOR U619 ( .A(a[694]), .B(b[694]), .Z(n3412) );
  OR U620 ( .A(a[693]), .B(b[693]), .Z(n1388) );
  XOR U621 ( .A(a[693]), .B(b[693]), .Z(n3410) );
  OR U622 ( .A(a[692]), .B(b[692]), .Z(n1386) );
  XOR U623 ( .A(a[692]), .B(b[692]), .Z(n3408) );
  OR U624 ( .A(a[691]), .B(b[691]), .Z(n1384) );
  XOR U625 ( .A(a[691]), .B(b[691]), .Z(n3406) );
  OR U626 ( .A(a[690]), .B(b[690]), .Z(n1382) );
  XOR U627 ( .A(a[690]), .B(b[690]), .Z(n3404) );
  OR U628 ( .A(a[689]), .B(b[689]), .Z(n1380) );
  XOR U629 ( .A(a[689]), .B(b[689]), .Z(n3400) );
  OR U630 ( .A(a[688]), .B(b[688]), .Z(n1378) );
  XOR U631 ( .A(a[688]), .B(b[688]), .Z(n3398) );
  OR U632 ( .A(a[687]), .B(b[687]), .Z(n1376) );
  XOR U633 ( .A(a[687]), .B(b[687]), .Z(n3396) );
  OR U634 ( .A(a[686]), .B(b[686]), .Z(n1374) );
  XOR U635 ( .A(a[686]), .B(b[686]), .Z(n3394) );
  OR U636 ( .A(a[685]), .B(b[685]), .Z(n1372) );
  XOR U637 ( .A(a[685]), .B(b[685]), .Z(n3392) );
  OR U638 ( .A(a[684]), .B(b[684]), .Z(n1370) );
  XOR U639 ( .A(a[684]), .B(b[684]), .Z(n3390) );
  OR U640 ( .A(a[683]), .B(b[683]), .Z(n1368) );
  XOR U641 ( .A(a[683]), .B(b[683]), .Z(n3388) );
  OR U642 ( .A(a[682]), .B(b[682]), .Z(n1366) );
  XOR U643 ( .A(a[682]), .B(b[682]), .Z(n3386) );
  OR U644 ( .A(a[681]), .B(b[681]), .Z(n1364) );
  XOR U645 ( .A(a[681]), .B(b[681]), .Z(n3384) );
  OR U646 ( .A(a[680]), .B(b[680]), .Z(n1362) );
  XOR U647 ( .A(a[680]), .B(b[680]), .Z(n3382) );
  OR U648 ( .A(a[679]), .B(b[679]), .Z(n1360) );
  XOR U649 ( .A(a[679]), .B(b[679]), .Z(n3378) );
  OR U650 ( .A(a[678]), .B(b[678]), .Z(n1358) );
  XOR U651 ( .A(a[678]), .B(b[678]), .Z(n3376) );
  OR U652 ( .A(a[677]), .B(b[677]), .Z(n1356) );
  XOR U653 ( .A(a[677]), .B(b[677]), .Z(n3374) );
  OR U654 ( .A(a[676]), .B(b[676]), .Z(n1354) );
  XOR U655 ( .A(a[676]), .B(b[676]), .Z(n3372) );
  OR U656 ( .A(a[675]), .B(b[675]), .Z(n1352) );
  XOR U657 ( .A(a[675]), .B(b[675]), .Z(n3370) );
  OR U658 ( .A(a[674]), .B(b[674]), .Z(n1350) );
  XOR U659 ( .A(a[674]), .B(b[674]), .Z(n3368) );
  OR U660 ( .A(a[673]), .B(b[673]), .Z(n1348) );
  XOR U661 ( .A(a[673]), .B(b[673]), .Z(n3366) );
  OR U662 ( .A(a[672]), .B(b[672]), .Z(n1346) );
  XOR U663 ( .A(a[672]), .B(b[672]), .Z(n3364) );
  OR U664 ( .A(a[671]), .B(b[671]), .Z(n1344) );
  XOR U665 ( .A(a[671]), .B(b[671]), .Z(n3362) );
  OR U666 ( .A(a[670]), .B(b[670]), .Z(n1342) );
  XOR U667 ( .A(a[670]), .B(b[670]), .Z(n3360) );
  OR U668 ( .A(a[669]), .B(b[669]), .Z(n1340) );
  XOR U669 ( .A(a[669]), .B(b[669]), .Z(n3356) );
  OR U670 ( .A(a[668]), .B(b[668]), .Z(n1338) );
  XOR U671 ( .A(a[668]), .B(b[668]), .Z(n3354) );
  OR U672 ( .A(a[667]), .B(b[667]), .Z(n1336) );
  XOR U673 ( .A(a[667]), .B(b[667]), .Z(n3352) );
  OR U674 ( .A(a[666]), .B(b[666]), .Z(n1334) );
  XOR U675 ( .A(a[666]), .B(b[666]), .Z(n3350) );
  OR U676 ( .A(a[665]), .B(b[665]), .Z(n1332) );
  XOR U677 ( .A(a[665]), .B(b[665]), .Z(n3348) );
  OR U678 ( .A(a[664]), .B(b[664]), .Z(n1330) );
  XOR U679 ( .A(a[664]), .B(b[664]), .Z(n3346) );
  OR U680 ( .A(a[663]), .B(b[663]), .Z(n1328) );
  XOR U681 ( .A(a[663]), .B(b[663]), .Z(n3344) );
  OR U682 ( .A(a[662]), .B(b[662]), .Z(n1326) );
  XOR U683 ( .A(a[662]), .B(b[662]), .Z(n3342) );
  OR U684 ( .A(a[661]), .B(b[661]), .Z(n1324) );
  XOR U685 ( .A(a[661]), .B(b[661]), .Z(n3340) );
  OR U686 ( .A(a[660]), .B(b[660]), .Z(n1322) );
  XOR U687 ( .A(a[660]), .B(b[660]), .Z(n3338) );
  OR U688 ( .A(a[659]), .B(b[659]), .Z(n1320) );
  XOR U689 ( .A(a[659]), .B(b[659]), .Z(n3334) );
  OR U690 ( .A(a[658]), .B(b[658]), .Z(n1318) );
  XOR U691 ( .A(a[658]), .B(b[658]), .Z(n3332) );
  OR U692 ( .A(a[657]), .B(b[657]), .Z(n1316) );
  XOR U693 ( .A(a[657]), .B(b[657]), .Z(n3330) );
  OR U694 ( .A(a[656]), .B(b[656]), .Z(n1314) );
  XOR U695 ( .A(a[656]), .B(b[656]), .Z(n3328) );
  OR U696 ( .A(a[655]), .B(b[655]), .Z(n1312) );
  XOR U697 ( .A(a[655]), .B(b[655]), .Z(n3326) );
  OR U698 ( .A(a[654]), .B(b[654]), .Z(n1310) );
  XOR U699 ( .A(a[654]), .B(b[654]), .Z(n3324) );
  OR U700 ( .A(a[653]), .B(b[653]), .Z(n1308) );
  XOR U701 ( .A(a[653]), .B(b[653]), .Z(n3322) );
  OR U702 ( .A(a[652]), .B(b[652]), .Z(n1306) );
  XOR U703 ( .A(a[652]), .B(b[652]), .Z(n3320) );
  OR U704 ( .A(a[651]), .B(b[651]), .Z(n1304) );
  XOR U705 ( .A(a[651]), .B(b[651]), .Z(n3318) );
  OR U706 ( .A(a[650]), .B(b[650]), .Z(n1302) );
  XOR U707 ( .A(a[650]), .B(b[650]), .Z(n3316) );
  OR U708 ( .A(a[649]), .B(b[649]), .Z(n1300) );
  XOR U709 ( .A(a[649]), .B(b[649]), .Z(n3312) );
  OR U710 ( .A(a[648]), .B(b[648]), .Z(n1298) );
  XOR U711 ( .A(a[648]), .B(b[648]), .Z(n3310) );
  OR U712 ( .A(a[647]), .B(b[647]), .Z(n1296) );
  XOR U713 ( .A(a[647]), .B(b[647]), .Z(n3308) );
  OR U714 ( .A(a[646]), .B(b[646]), .Z(n1294) );
  XOR U715 ( .A(a[646]), .B(b[646]), .Z(n3306) );
  OR U716 ( .A(a[645]), .B(b[645]), .Z(n1292) );
  XOR U717 ( .A(a[645]), .B(b[645]), .Z(n3304) );
  OR U718 ( .A(a[644]), .B(b[644]), .Z(n1290) );
  XOR U719 ( .A(a[644]), .B(b[644]), .Z(n3302) );
  OR U720 ( .A(a[643]), .B(b[643]), .Z(n1288) );
  XOR U721 ( .A(a[643]), .B(b[643]), .Z(n3300) );
  OR U722 ( .A(a[642]), .B(b[642]), .Z(n1286) );
  XOR U723 ( .A(a[642]), .B(b[642]), .Z(n3298) );
  OR U724 ( .A(a[641]), .B(b[641]), .Z(n1284) );
  XOR U725 ( .A(a[641]), .B(b[641]), .Z(n3296) );
  OR U726 ( .A(a[640]), .B(b[640]), .Z(n1282) );
  XOR U727 ( .A(a[640]), .B(b[640]), .Z(n3294) );
  OR U728 ( .A(a[639]), .B(b[639]), .Z(n1280) );
  XOR U729 ( .A(a[639]), .B(b[639]), .Z(n3290) );
  OR U730 ( .A(a[638]), .B(b[638]), .Z(n1278) );
  XOR U731 ( .A(a[638]), .B(b[638]), .Z(n3288) );
  OR U732 ( .A(a[637]), .B(b[637]), .Z(n1276) );
  XOR U733 ( .A(a[637]), .B(b[637]), .Z(n3286) );
  OR U734 ( .A(a[636]), .B(b[636]), .Z(n1274) );
  XOR U735 ( .A(a[636]), .B(b[636]), .Z(n3284) );
  OR U736 ( .A(a[635]), .B(b[635]), .Z(n1272) );
  XOR U737 ( .A(a[635]), .B(b[635]), .Z(n3282) );
  OR U738 ( .A(a[634]), .B(b[634]), .Z(n1270) );
  XOR U739 ( .A(a[634]), .B(b[634]), .Z(n3280) );
  OR U740 ( .A(a[633]), .B(b[633]), .Z(n1268) );
  XOR U741 ( .A(a[633]), .B(b[633]), .Z(n3278) );
  OR U742 ( .A(a[632]), .B(b[632]), .Z(n1266) );
  XOR U743 ( .A(a[632]), .B(b[632]), .Z(n3276) );
  OR U744 ( .A(a[631]), .B(b[631]), .Z(n1264) );
  XOR U745 ( .A(a[631]), .B(b[631]), .Z(n3274) );
  OR U746 ( .A(a[630]), .B(b[630]), .Z(n1262) );
  XOR U747 ( .A(a[630]), .B(b[630]), .Z(n3272) );
  OR U748 ( .A(a[629]), .B(b[629]), .Z(n1260) );
  XOR U749 ( .A(a[629]), .B(b[629]), .Z(n3268) );
  OR U750 ( .A(a[628]), .B(b[628]), .Z(n1258) );
  XOR U751 ( .A(a[628]), .B(b[628]), .Z(n3266) );
  OR U752 ( .A(a[627]), .B(b[627]), .Z(n1256) );
  XOR U753 ( .A(a[627]), .B(b[627]), .Z(n3264) );
  OR U754 ( .A(a[626]), .B(b[626]), .Z(n1254) );
  XOR U755 ( .A(a[626]), .B(b[626]), .Z(n3262) );
  OR U756 ( .A(a[625]), .B(b[625]), .Z(n1252) );
  XOR U757 ( .A(a[625]), .B(b[625]), .Z(n3260) );
  OR U758 ( .A(a[624]), .B(b[624]), .Z(n1250) );
  XOR U759 ( .A(a[624]), .B(b[624]), .Z(n3258) );
  OR U760 ( .A(a[623]), .B(b[623]), .Z(n1248) );
  XOR U761 ( .A(a[623]), .B(b[623]), .Z(n3256) );
  OR U762 ( .A(a[622]), .B(b[622]), .Z(n1246) );
  XOR U763 ( .A(a[622]), .B(b[622]), .Z(n3254) );
  OR U764 ( .A(a[621]), .B(b[621]), .Z(n1244) );
  XOR U765 ( .A(a[621]), .B(b[621]), .Z(n3252) );
  OR U766 ( .A(a[620]), .B(b[620]), .Z(n1242) );
  XOR U767 ( .A(a[620]), .B(b[620]), .Z(n3250) );
  OR U768 ( .A(a[619]), .B(b[619]), .Z(n1240) );
  XOR U769 ( .A(a[619]), .B(b[619]), .Z(n3246) );
  OR U770 ( .A(a[618]), .B(b[618]), .Z(n1238) );
  XOR U771 ( .A(a[618]), .B(b[618]), .Z(n3244) );
  OR U772 ( .A(a[617]), .B(b[617]), .Z(n1236) );
  XOR U773 ( .A(a[617]), .B(b[617]), .Z(n3242) );
  OR U774 ( .A(a[616]), .B(b[616]), .Z(n1234) );
  XOR U775 ( .A(a[616]), .B(b[616]), .Z(n3240) );
  OR U776 ( .A(a[615]), .B(b[615]), .Z(n1232) );
  XOR U777 ( .A(a[615]), .B(b[615]), .Z(n3238) );
  OR U778 ( .A(a[614]), .B(b[614]), .Z(n1230) );
  XOR U779 ( .A(a[614]), .B(b[614]), .Z(n3236) );
  OR U780 ( .A(a[613]), .B(b[613]), .Z(n1228) );
  XOR U781 ( .A(a[613]), .B(b[613]), .Z(n3234) );
  OR U782 ( .A(a[612]), .B(b[612]), .Z(n1226) );
  XOR U783 ( .A(a[612]), .B(b[612]), .Z(n3232) );
  OR U784 ( .A(a[611]), .B(b[611]), .Z(n1224) );
  XOR U785 ( .A(a[611]), .B(b[611]), .Z(n3230) );
  OR U786 ( .A(a[610]), .B(b[610]), .Z(n1222) );
  XOR U787 ( .A(a[610]), .B(b[610]), .Z(n3228) );
  OR U788 ( .A(a[609]), .B(b[609]), .Z(n1220) );
  XOR U789 ( .A(a[609]), .B(b[609]), .Z(n3224) );
  OR U790 ( .A(a[608]), .B(b[608]), .Z(n1218) );
  XOR U791 ( .A(a[608]), .B(b[608]), .Z(n3222) );
  OR U792 ( .A(a[607]), .B(b[607]), .Z(n1216) );
  XOR U793 ( .A(a[607]), .B(b[607]), .Z(n3220) );
  OR U794 ( .A(a[606]), .B(b[606]), .Z(n1214) );
  XOR U795 ( .A(a[606]), .B(b[606]), .Z(n3218) );
  OR U796 ( .A(a[605]), .B(b[605]), .Z(n1212) );
  XOR U797 ( .A(a[605]), .B(b[605]), .Z(n3216) );
  OR U798 ( .A(a[604]), .B(b[604]), .Z(n1210) );
  XOR U799 ( .A(a[604]), .B(b[604]), .Z(n3214) );
  OR U800 ( .A(a[603]), .B(b[603]), .Z(n1208) );
  XOR U801 ( .A(a[603]), .B(b[603]), .Z(n3212) );
  OR U802 ( .A(a[602]), .B(b[602]), .Z(n1206) );
  XOR U803 ( .A(a[602]), .B(b[602]), .Z(n3210) );
  OR U804 ( .A(a[601]), .B(b[601]), .Z(n1204) );
  XOR U805 ( .A(a[601]), .B(b[601]), .Z(n3208) );
  OR U806 ( .A(a[600]), .B(b[600]), .Z(n1202) );
  XOR U807 ( .A(a[600]), .B(b[600]), .Z(n3206) );
  OR U808 ( .A(a[599]), .B(b[599]), .Z(n1200) );
  XOR U809 ( .A(a[599]), .B(b[599]), .Z(n3200) );
  OR U810 ( .A(a[598]), .B(b[598]), .Z(n1198) );
  XOR U811 ( .A(a[598]), .B(b[598]), .Z(n3198) );
  OR U812 ( .A(a[597]), .B(b[597]), .Z(n1196) );
  XOR U813 ( .A(a[597]), .B(b[597]), .Z(n3196) );
  OR U814 ( .A(a[596]), .B(b[596]), .Z(n1194) );
  XOR U815 ( .A(a[596]), .B(b[596]), .Z(n3194) );
  OR U816 ( .A(a[595]), .B(b[595]), .Z(n1192) );
  XOR U817 ( .A(a[595]), .B(b[595]), .Z(n3192) );
  OR U818 ( .A(a[594]), .B(b[594]), .Z(n1190) );
  XOR U819 ( .A(a[594]), .B(b[594]), .Z(n3190) );
  OR U820 ( .A(a[593]), .B(b[593]), .Z(n1188) );
  XOR U821 ( .A(a[593]), .B(b[593]), .Z(n3188) );
  OR U822 ( .A(a[592]), .B(b[592]), .Z(n1186) );
  XOR U823 ( .A(a[592]), .B(b[592]), .Z(n3186) );
  OR U824 ( .A(a[591]), .B(b[591]), .Z(n1184) );
  XOR U825 ( .A(a[591]), .B(b[591]), .Z(n3184) );
  OR U826 ( .A(a[590]), .B(b[590]), .Z(n1182) );
  XOR U827 ( .A(a[590]), .B(b[590]), .Z(n3182) );
  OR U828 ( .A(a[589]), .B(b[589]), .Z(n1180) );
  XOR U829 ( .A(a[589]), .B(b[589]), .Z(n3178) );
  OR U830 ( .A(a[588]), .B(b[588]), .Z(n1178) );
  XOR U831 ( .A(a[588]), .B(b[588]), .Z(n3176) );
  OR U832 ( .A(a[587]), .B(b[587]), .Z(n1176) );
  XOR U833 ( .A(a[587]), .B(b[587]), .Z(n3174) );
  OR U834 ( .A(a[586]), .B(b[586]), .Z(n1174) );
  XOR U835 ( .A(a[586]), .B(b[586]), .Z(n3172) );
  OR U836 ( .A(a[585]), .B(b[585]), .Z(n1172) );
  XOR U837 ( .A(a[585]), .B(b[585]), .Z(n3170) );
  OR U838 ( .A(a[584]), .B(b[584]), .Z(n1170) );
  XOR U839 ( .A(a[584]), .B(b[584]), .Z(n3168) );
  OR U840 ( .A(a[583]), .B(b[583]), .Z(n1168) );
  XOR U841 ( .A(a[583]), .B(b[583]), .Z(n3166) );
  OR U842 ( .A(a[582]), .B(b[582]), .Z(n1166) );
  XOR U843 ( .A(a[582]), .B(b[582]), .Z(n3164) );
  OR U844 ( .A(a[581]), .B(b[581]), .Z(n1164) );
  XOR U845 ( .A(a[581]), .B(b[581]), .Z(n3162) );
  OR U846 ( .A(a[580]), .B(b[580]), .Z(n1162) );
  XOR U847 ( .A(a[580]), .B(b[580]), .Z(n3160) );
  OR U848 ( .A(a[579]), .B(b[579]), .Z(n1160) );
  XOR U849 ( .A(a[579]), .B(b[579]), .Z(n3156) );
  OR U850 ( .A(a[578]), .B(b[578]), .Z(n1158) );
  XOR U851 ( .A(a[578]), .B(b[578]), .Z(n3154) );
  OR U852 ( .A(a[577]), .B(b[577]), .Z(n1156) );
  XOR U853 ( .A(a[577]), .B(b[577]), .Z(n3152) );
  OR U854 ( .A(a[576]), .B(b[576]), .Z(n1154) );
  XOR U855 ( .A(a[576]), .B(b[576]), .Z(n3150) );
  OR U856 ( .A(a[575]), .B(b[575]), .Z(n1152) );
  XOR U857 ( .A(a[575]), .B(b[575]), .Z(n3148) );
  OR U858 ( .A(a[574]), .B(b[574]), .Z(n1150) );
  XOR U859 ( .A(a[574]), .B(b[574]), .Z(n3146) );
  OR U860 ( .A(a[573]), .B(b[573]), .Z(n1148) );
  XOR U861 ( .A(a[573]), .B(b[573]), .Z(n3144) );
  OR U862 ( .A(a[572]), .B(b[572]), .Z(n1146) );
  XOR U863 ( .A(a[572]), .B(b[572]), .Z(n3142) );
  OR U864 ( .A(a[571]), .B(b[571]), .Z(n1144) );
  XOR U865 ( .A(a[571]), .B(b[571]), .Z(n3140) );
  OR U866 ( .A(a[570]), .B(b[570]), .Z(n1142) );
  XOR U867 ( .A(a[570]), .B(b[570]), .Z(n3138) );
  OR U868 ( .A(a[569]), .B(b[569]), .Z(n1140) );
  XOR U869 ( .A(a[569]), .B(b[569]), .Z(n3134) );
  OR U870 ( .A(a[568]), .B(b[568]), .Z(n1138) );
  XOR U871 ( .A(a[568]), .B(b[568]), .Z(n3132) );
  OR U872 ( .A(a[567]), .B(b[567]), .Z(n1136) );
  XOR U873 ( .A(a[567]), .B(b[567]), .Z(n3130) );
  OR U874 ( .A(a[566]), .B(b[566]), .Z(n1134) );
  XOR U875 ( .A(a[566]), .B(b[566]), .Z(n3128) );
  OR U876 ( .A(a[565]), .B(b[565]), .Z(n1132) );
  XOR U877 ( .A(a[565]), .B(b[565]), .Z(n3126) );
  OR U878 ( .A(a[564]), .B(b[564]), .Z(n1130) );
  XOR U879 ( .A(a[564]), .B(b[564]), .Z(n3124) );
  OR U880 ( .A(a[563]), .B(b[563]), .Z(n1128) );
  XOR U881 ( .A(a[563]), .B(b[563]), .Z(n3122) );
  OR U882 ( .A(a[562]), .B(b[562]), .Z(n1126) );
  XOR U883 ( .A(a[562]), .B(b[562]), .Z(n3120) );
  OR U884 ( .A(a[561]), .B(b[561]), .Z(n1124) );
  XOR U885 ( .A(a[561]), .B(b[561]), .Z(n3118) );
  OR U886 ( .A(a[560]), .B(b[560]), .Z(n1122) );
  XOR U887 ( .A(a[560]), .B(b[560]), .Z(n3116) );
  OR U888 ( .A(a[559]), .B(b[559]), .Z(n1120) );
  XOR U889 ( .A(a[559]), .B(b[559]), .Z(n3112) );
  OR U890 ( .A(a[558]), .B(b[558]), .Z(n1118) );
  XOR U891 ( .A(a[558]), .B(b[558]), .Z(n3110) );
  OR U892 ( .A(a[557]), .B(b[557]), .Z(n1116) );
  XOR U893 ( .A(a[557]), .B(b[557]), .Z(n3108) );
  OR U894 ( .A(a[556]), .B(b[556]), .Z(n1114) );
  XOR U895 ( .A(a[556]), .B(b[556]), .Z(n3106) );
  OR U896 ( .A(a[555]), .B(b[555]), .Z(n1112) );
  XOR U897 ( .A(a[555]), .B(b[555]), .Z(n3104) );
  OR U898 ( .A(a[554]), .B(b[554]), .Z(n1110) );
  XOR U899 ( .A(a[554]), .B(b[554]), .Z(n3102) );
  OR U900 ( .A(a[553]), .B(b[553]), .Z(n1108) );
  XOR U901 ( .A(a[553]), .B(b[553]), .Z(n3100) );
  OR U902 ( .A(a[552]), .B(b[552]), .Z(n1106) );
  XOR U903 ( .A(a[552]), .B(b[552]), .Z(n3098) );
  OR U904 ( .A(a[551]), .B(b[551]), .Z(n1104) );
  XOR U905 ( .A(a[551]), .B(b[551]), .Z(n3096) );
  OR U906 ( .A(a[550]), .B(b[550]), .Z(n1102) );
  XOR U907 ( .A(a[550]), .B(b[550]), .Z(n3094) );
  OR U908 ( .A(a[549]), .B(b[549]), .Z(n1100) );
  XOR U909 ( .A(a[549]), .B(b[549]), .Z(n3090) );
  OR U910 ( .A(a[548]), .B(b[548]), .Z(n1098) );
  XOR U911 ( .A(a[548]), .B(b[548]), .Z(n3088) );
  OR U912 ( .A(a[547]), .B(b[547]), .Z(n1096) );
  XOR U913 ( .A(a[547]), .B(b[547]), .Z(n3086) );
  OR U914 ( .A(a[546]), .B(b[546]), .Z(n1094) );
  XOR U915 ( .A(a[546]), .B(b[546]), .Z(n3084) );
  OR U916 ( .A(a[545]), .B(b[545]), .Z(n1092) );
  XOR U917 ( .A(a[545]), .B(b[545]), .Z(n3082) );
  OR U918 ( .A(a[544]), .B(b[544]), .Z(n1090) );
  XOR U919 ( .A(a[544]), .B(b[544]), .Z(n3080) );
  OR U920 ( .A(a[543]), .B(b[543]), .Z(n1088) );
  XOR U921 ( .A(a[543]), .B(b[543]), .Z(n3078) );
  OR U922 ( .A(a[542]), .B(b[542]), .Z(n1086) );
  XOR U923 ( .A(a[542]), .B(b[542]), .Z(n3076) );
  OR U924 ( .A(a[541]), .B(b[541]), .Z(n1084) );
  XOR U925 ( .A(a[541]), .B(b[541]), .Z(n3074) );
  OR U926 ( .A(a[540]), .B(b[540]), .Z(n1082) );
  XOR U927 ( .A(a[540]), .B(b[540]), .Z(n3072) );
  OR U928 ( .A(a[539]), .B(b[539]), .Z(n1080) );
  XOR U929 ( .A(a[539]), .B(b[539]), .Z(n3068) );
  OR U930 ( .A(a[538]), .B(b[538]), .Z(n1078) );
  XOR U931 ( .A(a[538]), .B(b[538]), .Z(n3066) );
  OR U932 ( .A(a[537]), .B(b[537]), .Z(n1076) );
  XOR U933 ( .A(a[537]), .B(b[537]), .Z(n3064) );
  OR U934 ( .A(a[536]), .B(b[536]), .Z(n1074) );
  XOR U935 ( .A(a[536]), .B(b[536]), .Z(n3062) );
  OR U936 ( .A(a[535]), .B(b[535]), .Z(n1072) );
  XOR U937 ( .A(a[535]), .B(b[535]), .Z(n3060) );
  OR U938 ( .A(a[534]), .B(b[534]), .Z(n1070) );
  XOR U939 ( .A(a[534]), .B(b[534]), .Z(n3058) );
  OR U940 ( .A(a[533]), .B(b[533]), .Z(n1068) );
  XOR U941 ( .A(a[533]), .B(b[533]), .Z(n3056) );
  OR U942 ( .A(a[532]), .B(b[532]), .Z(n1066) );
  XOR U943 ( .A(a[532]), .B(b[532]), .Z(n3054) );
  OR U944 ( .A(a[531]), .B(b[531]), .Z(n1064) );
  XOR U945 ( .A(a[531]), .B(b[531]), .Z(n3052) );
  OR U946 ( .A(a[530]), .B(b[530]), .Z(n1062) );
  XOR U947 ( .A(a[530]), .B(b[530]), .Z(n3050) );
  OR U948 ( .A(a[529]), .B(b[529]), .Z(n1060) );
  XOR U949 ( .A(a[529]), .B(b[529]), .Z(n3046) );
  OR U950 ( .A(a[528]), .B(b[528]), .Z(n1058) );
  XOR U951 ( .A(a[528]), .B(b[528]), .Z(n3044) );
  OR U952 ( .A(a[527]), .B(b[527]), .Z(n1056) );
  XOR U953 ( .A(a[527]), .B(b[527]), .Z(n3042) );
  OR U954 ( .A(a[526]), .B(b[526]), .Z(n1054) );
  XOR U955 ( .A(a[526]), .B(b[526]), .Z(n3040) );
  OR U956 ( .A(a[525]), .B(b[525]), .Z(n1052) );
  XOR U957 ( .A(a[525]), .B(b[525]), .Z(n3038) );
  OR U958 ( .A(a[524]), .B(b[524]), .Z(n1050) );
  XOR U959 ( .A(a[524]), .B(b[524]), .Z(n3036) );
  OR U960 ( .A(a[523]), .B(b[523]), .Z(n1048) );
  XOR U961 ( .A(a[523]), .B(b[523]), .Z(n3034) );
  OR U962 ( .A(a[522]), .B(b[522]), .Z(n1046) );
  XOR U963 ( .A(a[522]), .B(b[522]), .Z(n3032) );
  OR U964 ( .A(a[521]), .B(b[521]), .Z(n1044) );
  XOR U965 ( .A(a[521]), .B(b[521]), .Z(n3030) );
  OR U966 ( .A(a[520]), .B(b[520]), .Z(n1042) );
  XOR U967 ( .A(a[520]), .B(b[520]), .Z(n3028) );
  OR U968 ( .A(a[519]), .B(b[519]), .Z(n1040) );
  XOR U969 ( .A(a[519]), .B(b[519]), .Z(n3024) );
  OR U970 ( .A(a[518]), .B(b[518]), .Z(n1038) );
  XOR U971 ( .A(a[518]), .B(b[518]), .Z(n3022) );
  OR U972 ( .A(a[517]), .B(b[517]), .Z(n1036) );
  XOR U973 ( .A(a[517]), .B(b[517]), .Z(n3020) );
  OR U974 ( .A(a[516]), .B(b[516]), .Z(n1034) );
  XOR U975 ( .A(a[516]), .B(b[516]), .Z(n3018) );
  OR U976 ( .A(a[515]), .B(b[515]), .Z(n1032) );
  XOR U977 ( .A(a[515]), .B(b[515]), .Z(n3016) );
  OR U978 ( .A(a[514]), .B(b[514]), .Z(n1030) );
  XOR U979 ( .A(a[514]), .B(b[514]), .Z(n3014) );
  OR U980 ( .A(a[513]), .B(b[513]), .Z(n1028) );
  XOR U981 ( .A(a[513]), .B(b[513]), .Z(n3012) );
  OR U982 ( .A(a[512]), .B(b[512]), .Z(n1026) );
  XOR U983 ( .A(a[512]), .B(b[512]), .Z(n3010) );
  OR U984 ( .A(a[511]), .B(b[511]), .Z(n1024) );
  XOR U985 ( .A(a[511]), .B(b[511]), .Z(n3008) );
  OR U986 ( .A(a[510]), .B(b[510]), .Z(n1022) );
  XOR U987 ( .A(a[510]), .B(b[510]), .Z(n3006) );
  OR U988 ( .A(a[509]), .B(b[509]), .Z(n1020) );
  XOR U989 ( .A(a[509]), .B(b[509]), .Z(n3002) );
  OR U990 ( .A(a[508]), .B(b[508]), .Z(n1018) );
  XOR U991 ( .A(a[508]), .B(b[508]), .Z(n3000) );
  OR U992 ( .A(a[507]), .B(b[507]), .Z(n1016) );
  XOR U993 ( .A(a[507]), .B(b[507]), .Z(n2998) );
  OR U994 ( .A(a[506]), .B(b[506]), .Z(n1014) );
  XOR U995 ( .A(a[506]), .B(b[506]), .Z(n2996) );
  OR U996 ( .A(a[505]), .B(b[505]), .Z(n1012) );
  XOR U997 ( .A(a[505]), .B(b[505]), .Z(n2994) );
  OR U998 ( .A(a[504]), .B(b[504]), .Z(n1010) );
  XOR U999 ( .A(a[504]), .B(b[504]), .Z(n2992) );
  OR U1000 ( .A(a[503]), .B(b[503]), .Z(n1008) );
  XOR U1001 ( .A(a[503]), .B(b[503]), .Z(n2990) );
  OR U1002 ( .A(a[502]), .B(b[502]), .Z(n1006) );
  XOR U1003 ( .A(a[502]), .B(b[502]), .Z(n2988) );
  OR U1004 ( .A(a[501]), .B(b[501]), .Z(n1004) );
  XOR U1005 ( .A(a[501]), .B(b[501]), .Z(n2986) );
  OR U1006 ( .A(a[500]), .B(b[500]), .Z(n1002) );
  XOR U1007 ( .A(a[500]), .B(b[500]), .Z(n2984) );
  OR U1008 ( .A(a[499]), .B(b[499]), .Z(n1000) );
  XOR U1009 ( .A(a[499]), .B(b[499]), .Z(n2978) );
  OR U1010 ( .A(a[498]), .B(b[498]), .Z(n998) );
  XOR U1011 ( .A(a[498]), .B(b[498]), .Z(n2976) );
  OR U1012 ( .A(a[497]), .B(b[497]), .Z(n996) );
  XOR U1013 ( .A(a[497]), .B(b[497]), .Z(n2974) );
  OR U1014 ( .A(a[496]), .B(b[496]), .Z(n994) );
  XOR U1015 ( .A(a[496]), .B(b[496]), .Z(n2972) );
  OR U1016 ( .A(a[495]), .B(b[495]), .Z(n992) );
  XOR U1017 ( .A(a[495]), .B(b[495]), .Z(n2970) );
  OR U1018 ( .A(a[494]), .B(b[494]), .Z(n990) );
  XOR U1019 ( .A(a[494]), .B(b[494]), .Z(n2968) );
  OR U1020 ( .A(a[493]), .B(b[493]), .Z(n988) );
  XOR U1021 ( .A(a[493]), .B(b[493]), .Z(n2966) );
  OR U1022 ( .A(a[492]), .B(b[492]), .Z(n986) );
  XOR U1023 ( .A(a[492]), .B(b[492]), .Z(n2964) );
  OR U1024 ( .A(a[491]), .B(b[491]), .Z(n984) );
  XOR U1025 ( .A(a[491]), .B(b[491]), .Z(n2962) );
  OR U1026 ( .A(a[490]), .B(b[490]), .Z(n982) );
  XOR U1027 ( .A(a[490]), .B(b[490]), .Z(n2960) );
  OR U1028 ( .A(a[489]), .B(b[489]), .Z(n980) );
  XOR U1029 ( .A(a[489]), .B(b[489]), .Z(n2956) );
  OR U1030 ( .A(a[488]), .B(b[488]), .Z(n978) );
  XOR U1031 ( .A(a[488]), .B(b[488]), .Z(n2954) );
  OR U1032 ( .A(a[487]), .B(b[487]), .Z(n976) );
  XOR U1033 ( .A(a[487]), .B(b[487]), .Z(n2952) );
  OR U1034 ( .A(a[486]), .B(b[486]), .Z(n974) );
  XOR U1035 ( .A(a[486]), .B(b[486]), .Z(n2950) );
  OR U1036 ( .A(a[485]), .B(b[485]), .Z(n972) );
  XOR U1037 ( .A(a[485]), .B(b[485]), .Z(n2948) );
  OR U1038 ( .A(a[484]), .B(b[484]), .Z(n970) );
  XOR U1039 ( .A(a[484]), .B(b[484]), .Z(n2946) );
  OR U1040 ( .A(a[483]), .B(b[483]), .Z(n968) );
  XOR U1041 ( .A(a[483]), .B(b[483]), .Z(n2944) );
  OR U1042 ( .A(a[482]), .B(b[482]), .Z(n966) );
  XOR U1043 ( .A(a[482]), .B(b[482]), .Z(n2942) );
  OR U1044 ( .A(a[481]), .B(b[481]), .Z(n964) );
  XOR U1045 ( .A(a[481]), .B(b[481]), .Z(n2940) );
  OR U1046 ( .A(a[480]), .B(b[480]), .Z(n962) );
  XOR U1047 ( .A(a[480]), .B(b[480]), .Z(n2938) );
  OR U1048 ( .A(a[479]), .B(b[479]), .Z(n960) );
  XOR U1049 ( .A(a[479]), .B(b[479]), .Z(n2934) );
  OR U1050 ( .A(a[478]), .B(b[478]), .Z(n958) );
  XOR U1051 ( .A(a[478]), .B(b[478]), .Z(n2932) );
  OR U1052 ( .A(a[477]), .B(b[477]), .Z(n956) );
  XOR U1053 ( .A(a[477]), .B(b[477]), .Z(n2930) );
  OR U1054 ( .A(a[476]), .B(b[476]), .Z(n954) );
  XOR U1055 ( .A(a[476]), .B(b[476]), .Z(n2928) );
  OR U1056 ( .A(a[475]), .B(b[475]), .Z(n952) );
  XOR U1057 ( .A(a[475]), .B(b[475]), .Z(n2926) );
  OR U1058 ( .A(a[474]), .B(b[474]), .Z(n950) );
  XOR U1059 ( .A(a[474]), .B(b[474]), .Z(n2924) );
  OR U1060 ( .A(a[473]), .B(b[473]), .Z(n948) );
  XOR U1061 ( .A(a[473]), .B(b[473]), .Z(n2922) );
  OR U1062 ( .A(a[472]), .B(b[472]), .Z(n946) );
  XOR U1063 ( .A(a[472]), .B(b[472]), .Z(n2920) );
  OR U1064 ( .A(a[471]), .B(b[471]), .Z(n944) );
  XOR U1065 ( .A(a[471]), .B(b[471]), .Z(n2918) );
  OR U1066 ( .A(a[470]), .B(b[470]), .Z(n942) );
  XOR U1067 ( .A(a[470]), .B(b[470]), .Z(n2916) );
  OR U1068 ( .A(a[469]), .B(b[469]), .Z(n940) );
  XOR U1069 ( .A(a[469]), .B(b[469]), .Z(n2912) );
  OR U1070 ( .A(a[468]), .B(b[468]), .Z(n938) );
  XOR U1071 ( .A(a[468]), .B(b[468]), .Z(n2910) );
  OR U1072 ( .A(a[467]), .B(b[467]), .Z(n936) );
  XOR U1073 ( .A(a[467]), .B(b[467]), .Z(n2908) );
  OR U1074 ( .A(a[466]), .B(b[466]), .Z(n934) );
  XOR U1075 ( .A(a[466]), .B(b[466]), .Z(n2906) );
  OR U1076 ( .A(a[465]), .B(b[465]), .Z(n932) );
  XOR U1077 ( .A(a[465]), .B(b[465]), .Z(n2904) );
  OR U1078 ( .A(a[464]), .B(b[464]), .Z(n930) );
  XOR U1079 ( .A(a[464]), .B(b[464]), .Z(n2902) );
  OR U1080 ( .A(a[463]), .B(b[463]), .Z(n928) );
  XOR U1081 ( .A(a[463]), .B(b[463]), .Z(n2900) );
  OR U1082 ( .A(a[462]), .B(b[462]), .Z(n926) );
  XOR U1083 ( .A(a[462]), .B(b[462]), .Z(n2898) );
  OR U1084 ( .A(a[461]), .B(b[461]), .Z(n924) );
  XOR U1085 ( .A(a[461]), .B(b[461]), .Z(n2896) );
  OR U1086 ( .A(a[460]), .B(b[460]), .Z(n922) );
  XOR U1087 ( .A(a[460]), .B(b[460]), .Z(n2894) );
  OR U1088 ( .A(a[459]), .B(b[459]), .Z(n920) );
  XOR U1089 ( .A(a[459]), .B(b[459]), .Z(n2890) );
  OR U1090 ( .A(a[458]), .B(b[458]), .Z(n918) );
  XOR U1091 ( .A(a[458]), .B(b[458]), .Z(n2888) );
  OR U1092 ( .A(a[457]), .B(b[457]), .Z(n916) );
  XOR U1093 ( .A(a[457]), .B(b[457]), .Z(n2886) );
  OR U1094 ( .A(a[456]), .B(b[456]), .Z(n914) );
  XOR U1095 ( .A(a[456]), .B(b[456]), .Z(n2884) );
  OR U1096 ( .A(a[455]), .B(b[455]), .Z(n912) );
  XOR U1097 ( .A(a[455]), .B(b[455]), .Z(n2882) );
  OR U1098 ( .A(a[454]), .B(b[454]), .Z(n910) );
  XOR U1099 ( .A(a[454]), .B(b[454]), .Z(n2880) );
  OR U1100 ( .A(a[453]), .B(b[453]), .Z(n908) );
  XOR U1101 ( .A(a[453]), .B(b[453]), .Z(n2878) );
  OR U1102 ( .A(a[452]), .B(b[452]), .Z(n906) );
  XOR U1103 ( .A(a[452]), .B(b[452]), .Z(n2876) );
  OR U1104 ( .A(a[451]), .B(b[451]), .Z(n904) );
  XOR U1105 ( .A(a[451]), .B(b[451]), .Z(n2874) );
  OR U1106 ( .A(a[450]), .B(b[450]), .Z(n902) );
  XOR U1107 ( .A(a[450]), .B(b[450]), .Z(n2872) );
  OR U1108 ( .A(a[449]), .B(b[449]), .Z(n900) );
  XOR U1109 ( .A(a[449]), .B(b[449]), .Z(n2868) );
  OR U1110 ( .A(a[448]), .B(b[448]), .Z(n898) );
  XOR U1111 ( .A(a[448]), .B(b[448]), .Z(n2866) );
  OR U1112 ( .A(a[447]), .B(b[447]), .Z(n896) );
  XOR U1113 ( .A(a[447]), .B(b[447]), .Z(n2864) );
  OR U1114 ( .A(a[446]), .B(b[446]), .Z(n894) );
  XOR U1115 ( .A(a[446]), .B(b[446]), .Z(n2862) );
  OR U1116 ( .A(a[445]), .B(b[445]), .Z(n892) );
  XOR U1117 ( .A(a[445]), .B(b[445]), .Z(n2860) );
  OR U1118 ( .A(a[444]), .B(b[444]), .Z(n890) );
  XOR U1119 ( .A(a[444]), .B(b[444]), .Z(n2858) );
  OR U1120 ( .A(a[443]), .B(b[443]), .Z(n888) );
  XOR U1121 ( .A(a[443]), .B(b[443]), .Z(n2856) );
  OR U1122 ( .A(a[442]), .B(b[442]), .Z(n886) );
  XOR U1123 ( .A(a[442]), .B(b[442]), .Z(n2854) );
  OR U1124 ( .A(a[441]), .B(b[441]), .Z(n884) );
  XOR U1125 ( .A(a[441]), .B(b[441]), .Z(n2852) );
  OR U1126 ( .A(a[440]), .B(b[440]), .Z(n882) );
  XOR U1127 ( .A(a[440]), .B(b[440]), .Z(n2850) );
  OR U1128 ( .A(a[439]), .B(b[439]), .Z(n880) );
  XOR U1129 ( .A(a[439]), .B(b[439]), .Z(n2846) );
  OR U1130 ( .A(a[438]), .B(b[438]), .Z(n878) );
  XOR U1131 ( .A(a[438]), .B(b[438]), .Z(n2844) );
  OR U1132 ( .A(a[437]), .B(b[437]), .Z(n876) );
  XOR U1133 ( .A(a[437]), .B(b[437]), .Z(n2842) );
  OR U1134 ( .A(a[436]), .B(b[436]), .Z(n874) );
  XOR U1135 ( .A(a[436]), .B(b[436]), .Z(n2840) );
  OR U1136 ( .A(a[435]), .B(b[435]), .Z(n872) );
  XOR U1137 ( .A(a[435]), .B(b[435]), .Z(n2838) );
  OR U1138 ( .A(a[434]), .B(b[434]), .Z(n870) );
  XOR U1139 ( .A(a[434]), .B(b[434]), .Z(n2836) );
  OR U1140 ( .A(a[433]), .B(b[433]), .Z(n868) );
  XOR U1141 ( .A(a[433]), .B(b[433]), .Z(n2834) );
  OR U1142 ( .A(a[432]), .B(b[432]), .Z(n866) );
  XOR U1143 ( .A(a[432]), .B(b[432]), .Z(n2832) );
  OR U1144 ( .A(a[431]), .B(b[431]), .Z(n864) );
  XOR U1145 ( .A(a[431]), .B(b[431]), .Z(n2830) );
  OR U1146 ( .A(a[430]), .B(b[430]), .Z(n862) );
  XOR U1147 ( .A(a[430]), .B(b[430]), .Z(n2828) );
  OR U1148 ( .A(a[429]), .B(b[429]), .Z(n860) );
  XOR U1149 ( .A(a[429]), .B(b[429]), .Z(n2824) );
  OR U1150 ( .A(a[428]), .B(b[428]), .Z(n858) );
  XOR U1151 ( .A(a[428]), .B(b[428]), .Z(n2822) );
  OR U1152 ( .A(a[427]), .B(b[427]), .Z(n856) );
  XOR U1153 ( .A(a[427]), .B(b[427]), .Z(n2820) );
  OR U1154 ( .A(a[426]), .B(b[426]), .Z(n854) );
  XOR U1155 ( .A(a[426]), .B(b[426]), .Z(n2818) );
  OR U1156 ( .A(a[425]), .B(b[425]), .Z(n852) );
  XOR U1157 ( .A(a[425]), .B(b[425]), .Z(n2816) );
  OR U1158 ( .A(a[424]), .B(b[424]), .Z(n850) );
  XOR U1159 ( .A(a[424]), .B(b[424]), .Z(n2814) );
  OR U1160 ( .A(a[423]), .B(b[423]), .Z(n848) );
  XOR U1161 ( .A(a[423]), .B(b[423]), .Z(n2812) );
  OR U1162 ( .A(a[422]), .B(b[422]), .Z(n846) );
  XOR U1163 ( .A(a[422]), .B(b[422]), .Z(n2810) );
  OR U1164 ( .A(a[421]), .B(b[421]), .Z(n844) );
  XOR U1165 ( .A(a[421]), .B(b[421]), .Z(n2808) );
  OR U1166 ( .A(a[420]), .B(b[420]), .Z(n842) );
  XOR U1167 ( .A(a[420]), .B(b[420]), .Z(n2806) );
  OR U1168 ( .A(a[419]), .B(b[419]), .Z(n840) );
  XOR U1169 ( .A(a[419]), .B(b[419]), .Z(n2802) );
  OR U1170 ( .A(a[418]), .B(b[418]), .Z(n838) );
  XOR U1171 ( .A(a[418]), .B(b[418]), .Z(n2800) );
  OR U1172 ( .A(a[417]), .B(b[417]), .Z(n836) );
  XOR U1173 ( .A(a[417]), .B(b[417]), .Z(n2798) );
  OR U1174 ( .A(a[416]), .B(b[416]), .Z(n834) );
  XOR U1175 ( .A(a[416]), .B(b[416]), .Z(n2796) );
  OR U1176 ( .A(a[415]), .B(b[415]), .Z(n832) );
  XOR U1177 ( .A(a[415]), .B(b[415]), .Z(n2794) );
  OR U1178 ( .A(a[414]), .B(b[414]), .Z(n830) );
  XOR U1179 ( .A(a[414]), .B(b[414]), .Z(n2792) );
  OR U1180 ( .A(a[413]), .B(b[413]), .Z(n828) );
  XOR U1181 ( .A(a[413]), .B(b[413]), .Z(n2790) );
  OR U1182 ( .A(a[412]), .B(b[412]), .Z(n826) );
  XOR U1183 ( .A(a[412]), .B(b[412]), .Z(n2788) );
  OR U1184 ( .A(a[411]), .B(b[411]), .Z(n824) );
  XOR U1185 ( .A(a[411]), .B(b[411]), .Z(n2786) );
  OR U1186 ( .A(a[410]), .B(b[410]), .Z(n822) );
  XOR U1187 ( .A(a[410]), .B(b[410]), .Z(n2784) );
  OR U1188 ( .A(a[409]), .B(b[409]), .Z(n820) );
  XOR U1189 ( .A(a[409]), .B(b[409]), .Z(n2780) );
  OR U1190 ( .A(a[408]), .B(b[408]), .Z(n818) );
  XOR U1191 ( .A(a[408]), .B(b[408]), .Z(n2778) );
  OR U1192 ( .A(a[407]), .B(b[407]), .Z(n816) );
  XOR U1193 ( .A(a[407]), .B(b[407]), .Z(n2776) );
  OR U1194 ( .A(a[406]), .B(b[406]), .Z(n814) );
  XOR U1195 ( .A(a[406]), .B(b[406]), .Z(n2774) );
  OR U1196 ( .A(a[405]), .B(b[405]), .Z(n812) );
  XOR U1197 ( .A(a[405]), .B(b[405]), .Z(n2772) );
  OR U1198 ( .A(a[404]), .B(b[404]), .Z(n810) );
  XOR U1199 ( .A(a[404]), .B(b[404]), .Z(n2770) );
  OR U1200 ( .A(a[403]), .B(b[403]), .Z(n808) );
  XOR U1201 ( .A(a[403]), .B(b[403]), .Z(n2768) );
  OR U1202 ( .A(a[402]), .B(b[402]), .Z(n806) );
  XOR U1203 ( .A(a[402]), .B(b[402]), .Z(n2766) );
  OR U1204 ( .A(a[401]), .B(b[401]), .Z(n804) );
  XOR U1205 ( .A(a[401]), .B(b[401]), .Z(n2764) );
  OR U1206 ( .A(a[400]), .B(b[400]), .Z(n802) );
  XOR U1207 ( .A(a[400]), .B(b[400]), .Z(n2762) );
  OR U1208 ( .A(a[399]), .B(b[399]), .Z(n800) );
  XOR U1209 ( .A(a[399]), .B(b[399]), .Z(n2756) );
  OR U1210 ( .A(a[398]), .B(b[398]), .Z(n798) );
  XOR U1211 ( .A(a[398]), .B(b[398]), .Z(n2754) );
  OR U1212 ( .A(a[397]), .B(b[397]), .Z(n796) );
  XOR U1213 ( .A(a[397]), .B(b[397]), .Z(n2752) );
  OR U1214 ( .A(a[396]), .B(b[396]), .Z(n794) );
  XOR U1215 ( .A(a[396]), .B(b[396]), .Z(n2750) );
  OR U1216 ( .A(a[395]), .B(b[395]), .Z(n792) );
  XOR U1217 ( .A(a[395]), .B(b[395]), .Z(n2748) );
  OR U1218 ( .A(a[394]), .B(b[394]), .Z(n790) );
  XOR U1219 ( .A(a[394]), .B(b[394]), .Z(n2746) );
  OR U1220 ( .A(a[393]), .B(b[393]), .Z(n788) );
  XOR U1221 ( .A(a[393]), .B(b[393]), .Z(n2744) );
  OR U1222 ( .A(a[392]), .B(b[392]), .Z(n786) );
  XOR U1223 ( .A(a[392]), .B(b[392]), .Z(n2742) );
  OR U1224 ( .A(a[391]), .B(b[391]), .Z(n784) );
  XOR U1225 ( .A(a[391]), .B(b[391]), .Z(n2740) );
  OR U1226 ( .A(a[390]), .B(b[390]), .Z(n782) );
  XOR U1227 ( .A(a[390]), .B(b[390]), .Z(n2738) );
  OR U1228 ( .A(a[389]), .B(b[389]), .Z(n780) );
  XOR U1229 ( .A(a[389]), .B(b[389]), .Z(n2734) );
  OR U1230 ( .A(a[388]), .B(b[388]), .Z(n778) );
  XOR U1231 ( .A(a[388]), .B(b[388]), .Z(n2732) );
  OR U1232 ( .A(a[387]), .B(b[387]), .Z(n776) );
  XOR U1233 ( .A(a[387]), .B(b[387]), .Z(n2730) );
  OR U1234 ( .A(a[386]), .B(b[386]), .Z(n774) );
  XOR U1235 ( .A(a[386]), .B(b[386]), .Z(n2728) );
  OR U1236 ( .A(a[385]), .B(b[385]), .Z(n772) );
  XOR U1237 ( .A(a[385]), .B(b[385]), .Z(n2726) );
  OR U1238 ( .A(a[384]), .B(b[384]), .Z(n770) );
  XOR U1239 ( .A(a[384]), .B(b[384]), .Z(n2724) );
  OR U1240 ( .A(a[383]), .B(b[383]), .Z(n768) );
  XOR U1241 ( .A(a[383]), .B(b[383]), .Z(n2722) );
  OR U1242 ( .A(a[382]), .B(b[382]), .Z(n766) );
  XOR U1243 ( .A(a[382]), .B(b[382]), .Z(n2720) );
  OR U1244 ( .A(a[381]), .B(b[381]), .Z(n764) );
  XOR U1245 ( .A(a[381]), .B(b[381]), .Z(n2718) );
  OR U1246 ( .A(a[380]), .B(b[380]), .Z(n762) );
  XOR U1247 ( .A(a[380]), .B(b[380]), .Z(n2716) );
  OR U1248 ( .A(a[379]), .B(b[379]), .Z(n760) );
  XOR U1249 ( .A(a[379]), .B(b[379]), .Z(n2712) );
  OR U1250 ( .A(a[378]), .B(b[378]), .Z(n758) );
  XOR U1251 ( .A(a[378]), .B(b[378]), .Z(n2710) );
  OR U1252 ( .A(a[377]), .B(b[377]), .Z(n756) );
  XOR U1253 ( .A(a[377]), .B(b[377]), .Z(n2708) );
  OR U1254 ( .A(a[376]), .B(b[376]), .Z(n754) );
  XOR U1255 ( .A(a[376]), .B(b[376]), .Z(n2706) );
  OR U1256 ( .A(a[375]), .B(b[375]), .Z(n752) );
  XOR U1257 ( .A(a[375]), .B(b[375]), .Z(n2704) );
  OR U1258 ( .A(a[374]), .B(b[374]), .Z(n750) );
  XOR U1259 ( .A(a[374]), .B(b[374]), .Z(n2702) );
  OR U1260 ( .A(a[373]), .B(b[373]), .Z(n748) );
  XOR U1261 ( .A(a[373]), .B(b[373]), .Z(n2700) );
  OR U1262 ( .A(a[372]), .B(b[372]), .Z(n746) );
  XOR U1263 ( .A(a[372]), .B(b[372]), .Z(n2698) );
  OR U1264 ( .A(a[371]), .B(b[371]), .Z(n744) );
  XOR U1265 ( .A(a[371]), .B(b[371]), .Z(n2696) );
  OR U1266 ( .A(a[370]), .B(b[370]), .Z(n742) );
  XOR U1267 ( .A(a[370]), .B(b[370]), .Z(n2694) );
  OR U1268 ( .A(a[369]), .B(b[369]), .Z(n740) );
  XOR U1269 ( .A(a[369]), .B(b[369]), .Z(n2690) );
  OR U1270 ( .A(a[368]), .B(b[368]), .Z(n738) );
  XOR U1271 ( .A(a[368]), .B(b[368]), .Z(n2688) );
  OR U1272 ( .A(a[367]), .B(b[367]), .Z(n736) );
  XOR U1273 ( .A(a[367]), .B(b[367]), .Z(n2686) );
  OR U1274 ( .A(a[366]), .B(b[366]), .Z(n734) );
  XOR U1275 ( .A(a[366]), .B(b[366]), .Z(n2684) );
  OR U1276 ( .A(a[365]), .B(b[365]), .Z(n732) );
  XOR U1277 ( .A(a[365]), .B(b[365]), .Z(n2682) );
  OR U1278 ( .A(a[364]), .B(b[364]), .Z(n730) );
  XOR U1279 ( .A(a[364]), .B(b[364]), .Z(n2680) );
  OR U1280 ( .A(a[363]), .B(b[363]), .Z(n728) );
  XOR U1281 ( .A(a[363]), .B(b[363]), .Z(n2678) );
  OR U1282 ( .A(a[362]), .B(b[362]), .Z(n726) );
  XOR U1283 ( .A(a[362]), .B(b[362]), .Z(n2676) );
  OR U1284 ( .A(a[361]), .B(b[361]), .Z(n724) );
  XOR U1285 ( .A(a[361]), .B(b[361]), .Z(n2674) );
  OR U1286 ( .A(a[360]), .B(b[360]), .Z(n722) );
  XOR U1287 ( .A(a[360]), .B(b[360]), .Z(n2672) );
  OR U1288 ( .A(a[359]), .B(b[359]), .Z(n720) );
  XOR U1289 ( .A(a[359]), .B(b[359]), .Z(n2668) );
  OR U1290 ( .A(a[358]), .B(b[358]), .Z(n718) );
  XOR U1291 ( .A(a[358]), .B(b[358]), .Z(n2666) );
  OR U1292 ( .A(a[357]), .B(b[357]), .Z(n716) );
  XOR U1293 ( .A(a[357]), .B(b[357]), .Z(n2664) );
  OR U1294 ( .A(a[356]), .B(b[356]), .Z(n714) );
  XOR U1295 ( .A(a[356]), .B(b[356]), .Z(n2662) );
  OR U1296 ( .A(a[355]), .B(b[355]), .Z(n712) );
  XOR U1297 ( .A(a[355]), .B(b[355]), .Z(n2660) );
  OR U1298 ( .A(a[354]), .B(b[354]), .Z(n710) );
  XOR U1299 ( .A(a[354]), .B(b[354]), .Z(n2658) );
  OR U1300 ( .A(a[353]), .B(b[353]), .Z(n708) );
  XOR U1301 ( .A(a[353]), .B(b[353]), .Z(n2656) );
  OR U1302 ( .A(a[352]), .B(b[352]), .Z(n706) );
  XOR U1303 ( .A(a[352]), .B(b[352]), .Z(n2654) );
  OR U1304 ( .A(a[351]), .B(b[351]), .Z(n704) );
  XOR U1305 ( .A(a[351]), .B(b[351]), .Z(n2652) );
  OR U1306 ( .A(a[350]), .B(b[350]), .Z(n702) );
  XOR U1307 ( .A(a[350]), .B(b[350]), .Z(n2650) );
  OR U1308 ( .A(a[349]), .B(b[349]), .Z(n700) );
  XOR U1309 ( .A(a[349]), .B(b[349]), .Z(n2646) );
  OR U1310 ( .A(a[348]), .B(b[348]), .Z(n698) );
  XOR U1311 ( .A(a[348]), .B(b[348]), .Z(n2644) );
  OR U1312 ( .A(a[347]), .B(b[347]), .Z(n696) );
  XOR U1313 ( .A(a[347]), .B(b[347]), .Z(n2642) );
  OR U1314 ( .A(a[346]), .B(b[346]), .Z(n694) );
  XOR U1315 ( .A(a[346]), .B(b[346]), .Z(n2640) );
  OR U1316 ( .A(a[345]), .B(b[345]), .Z(n692) );
  XOR U1317 ( .A(a[345]), .B(b[345]), .Z(n2638) );
  OR U1318 ( .A(a[344]), .B(b[344]), .Z(n690) );
  XOR U1319 ( .A(a[344]), .B(b[344]), .Z(n2636) );
  OR U1320 ( .A(a[343]), .B(b[343]), .Z(n688) );
  XOR U1321 ( .A(a[343]), .B(b[343]), .Z(n2634) );
  OR U1322 ( .A(a[342]), .B(b[342]), .Z(n686) );
  XOR U1323 ( .A(a[342]), .B(b[342]), .Z(n2632) );
  OR U1324 ( .A(a[341]), .B(b[341]), .Z(n684) );
  XOR U1325 ( .A(a[341]), .B(b[341]), .Z(n2630) );
  OR U1326 ( .A(a[340]), .B(b[340]), .Z(n682) );
  XOR U1327 ( .A(a[340]), .B(b[340]), .Z(n2628) );
  OR U1328 ( .A(a[339]), .B(b[339]), .Z(n680) );
  XOR U1329 ( .A(a[339]), .B(b[339]), .Z(n2624) );
  OR U1330 ( .A(a[338]), .B(b[338]), .Z(n678) );
  XOR U1331 ( .A(a[338]), .B(b[338]), .Z(n2622) );
  OR U1332 ( .A(a[337]), .B(b[337]), .Z(n676) );
  XOR U1333 ( .A(a[337]), .B(b[337]), .Z(n2620) );
  OR U1334 ( .A(a[336]), .B(b[336]), .Z(n674) );
  XOR U1335 ( .A(a[336]), .B(b[336]), .Z(n2618) );
  OR U1336 ( .A(a[335]), .B(b[335]), .Z(n672) );
  XOR U1337 ( .A(a[335]), .B(b[335]), .Z(n2616) );
  OR U1338 ( .A(a[334]), .B(b[334]), .Z(n670) );
  XOR U1339 ( .A(a[334]), .B(b[334]), .Z(n2614) );
  OR U1340 ( .A(a[333]), .B(b[333]), .Z(n668) );
  XOR U1341 ( .A(a[333]), .B(b[333]), .Z(n2612) );
  OR U1342 ( .A(a[332]), .B(b[332]), .Z(n666) );
  XOR U1343 ( .A(a[332]), .B(b[332]), .Z(n2610) );
  OR U1344 ( .A(a[331]), .B(b[331]), .Z(n664) );
  XOR U1345 ( .A(a[331]), .B(b[331]), .Z(n2608) );
  OR U1346 ( .A(a[330]), .B(b[330]), .Z(n662) );
  XOR U1347 ( .A(a[330]), .B(b[330]), .Z(n2606) );
  OR U1348 ( .A(a[329]), .B(b[329]), .Z(n660) );
  XOR U1349 ( .A(a[329]), .B(b[329]), .Z(n2602) );
  OR U1350 ( .A(a[328]), .B(b[328]), .Z(n658) );
  XOR U1351 ( .A(a[328]), .B(b[328]), .Z(n2600) );
  OR U1352 ( .A(a[327]), .B(b[327]), .Z(n656) );
  XOR U1353 ( .A(a[327]), .B(b[327]), .Z(n2598) );
  OR U1354 ( .A(a[326]), .B(b[326]), .Z(n654) );
  XOR U1355 ( .A(a[326]), .B(b[326]), .Z(n2596) );
  OR U1356 ( .A(a[325]), .B(b[325]), .Z(n652) );
  XOR U1357 ( .A(a[325]), .B(b[325]), .Z(n2594) );
  OR U1358 ( .A(a[324]), .B(b[324]), .Z(n650) );
  XOR U1359 ( .A(a[324]), .B(b[324]), .Z(n2592) );
  OR U1360 ( .A(a[323]), .B(b[323]), .Z(n648) );
  XOR U1361 ( .A(a[323]), .B(b[323]), .Z(n2590) );
  OR U1362 ( .A(a[322]), .B(b[322]), .Z(n646) );
  XOR U1363 ( .A(a[322]), .B(b[322]), .Z(n2588) );
  OR U1364 ( .A(a[321]), .B(b[321]), .Z(n644) );
  XOR U1365 ( .A(a[321]), .B(b[321]), .Z(n2586) );
  OR U1366 ( .A(a[320]), .B(b[320]), .Z(n642) );
  XOR U1367 ( .A(a[320]), .B(b[320]), .Z(n2584) );
  OR U1368 ( .A(a[319]), .B(b[319]), .Z(n640) );
  XOR U1369 ( .A(a[319]), .B(b[319]), .Z(n2580) );
  OR U1370 ( .A(a[318]), .B(b[318]), .Z(n638) );
  XOR U1371 ( .A(a[318]), .B(b[318]), .Z(n2578) );
  OR U1372 ( .A(a[317]), .B(b[317]), .Z(n636) );
  XOR U1373 ( .A(a[317]), .B(b[317]), .Z(n2576) );
  OR U1374 ( .A(a[316]), .B(b[316]), .Z(n634) );
  XOR U1375 ( .A(a[316]), .B(b[316]), .Z(n2574) );
  OR U1376 ( .A(a[315]), .B(b[315]), .Z(n632) );
  XOR U1377 ( .A(a[315]), .B(b[315]), .Z(n2572) );
  OR U1378 ( .A(a[314]), .B(b[314]), .Z(n630) );
  XOR U1379 ( .A(a[314]), .B(b[314]), .Z(n2570) );
  OR U1380 ( .A(a[313]), .B(b[313]), .Z(n628) );
  XOR U1381 ( .A(a[313]), .B(b[313]), .Z(n2568) );
  OR U1382 ( .A(a[312]), .B(b[312]), .Z(n626) );
  XOR U1383 ( .A(a[312]), .B(b[312]), .Z(n2566) );
  OR U1384 ( .A(a[311]), .B(b[311]), .Z(n624) );
  XOR U1385 ( .A(a[311]), .B(b[311]), .Z(n2564) );
  OR U1386 ( .A(a[310]), .B(b[310]), .Z(n622) );
  XOR U1387 ( .A(a[310]), .B(b[310]), .Z(n2562) );
  OR U1388 ( .A(a[309]), .B(b[309]), .Z(n620) );
  XOR U1389 ( .A(a[309]), .B(b[309]), .Z(n2558) );
  OR U1390 ( .A(a[308]), .B(b[308]), .Z(n618) );
  XOR U1391 ( .A(a[308]), .B(b[308]), .Z(n2556) );
  OR U1392 ( .A(a[307]), .B(b[307]), .Z(n616) );
  XOR U1393 ( .A(a[307]), .B(b[307]), .Z(n2554) );
  OR U1394 ( .A(a[306]), .B(b[306]), .Z(n614) );
  XOR U1395 ( .A(a[306]), .B(b[306]), .Z(n2552) );
  OR U1396 ( .A(a[305]), .B(b[305]), .Z(n612) );
  XOR U1397 ( .A(a[305]), .B(b[305]), .Z(n2550) );
  OR U1398 ( .A(a[304]), .B(b[304]), .Z(n610) );
  XOR U1399 ( .A(a[304]), .B(b[304]), .Z(n2548) );
  OR U1400 ( .A(a[303]), .B(b[303]), .Z(n608) );
  XOR U1401 ( .A(a[303]), .B(b[303]), .Z(n2546) );
  OR U1402 ( .A(a[302]), .B(b[302]), .Z(n606) );
  XOR U1403 ( .A(a[302]), .B(b[302]), .Z(n2544) );
  OR U1404 ( .A(a[301]), .B(b[301]), .Z(n604) );
  XOR U1405 ( .A(a[301]), .B(b[301]), .Z(n2542) );
  OR U1406 ( .A(a[300]), .B(b[300]), .Z(n602) );
  XOR U1407 ( .A(a[300]), .B(b[300]), .Z(n2540) );
  OR U1408 ( .A(a[299]), .B(b[299]), .Z(n600) );
  XOR U1409 ( .A(a[299]), .B(b[299]), .Z(n2534) );
  OR U1410 ( .A(a[298]), .B(b[298]), .Z(n598) );
  XOR U1411 ( .A(a[298]), .B(b[298]), .Z(n2532) );
  OR U1412 ( .A(a[297]), .B(b[297]), .Z(n596) );
  XOR U1413 ( .A(a[297]), .B(b[297]), .Z(n2530) );
  OR U1414 ( .A(a[296]), .B(b[296]), .Z(n594) );
  XOR U1415 ( .A(a[296]), .B(b[296]), .Z(n2528) );
  OR U1416 ( .A(a[295]), .B(b[295]), .Z(n592) );
  XOR U1417 ( .A(a[295]), .B(b[295]), .Z(n2526) );
  OR U1418 ( .A(a[294]), .B(b[294]), .Z(n590) );
  XOR U1419 ( .A(a[294]), .B(b[294]), .Z(n2524) );
  OR U1420 ( .A(a[293]), .B(b[293]), .Z(n588) );
  XOR U1421 ( .A(a[293]), .B(b[293]), .Z(n2522) );
  OR U1422 ( .A(a[292]), .B(b[292]), .Z(n586) );
  XOR U1423 ( .A(a[292]), .B(b[292]), .Z(n2520) );
  OR U1424 ( .A(a[291]), .B(b[291]), .Z(n584) );
  XOR U1425 ( .A(a[291]), .B(b[291]), .Z(n2518) );
  OR U1426 ( .A(a[290]), .B(b[290]), .Z(n582) );
  XOR U1427 ( .A(a[290]), .B(b[290]), .Z(n2516) );
  OR U1428 ( .A(a[289]), .B(b[289]), .Z(n580) );
  XOR U1429 ( .A(a[289]), .B(b[289]), .Z(n2512) );
  OR U1430 ( .A(a[288]), .B(b[288]), .Z(n578) );
  XOR U1431 ( .A(a[288]), .B(b[288]), .Z(n2510) );
  OR U1432 ( .A(a[287]), .B(b[287]), .Z(n576) );
  XOR U1433 ( .A(a[287]), .B(b[287]), .Z(n2508) );
  OR U1434 ( .A(a[286]), .B(b[286]), .Z(n574) );
  XOR U1435 ( .A(a[286]), .B(b[286]), .Z(n2506) );
  OR U1436 ( .A(a[285]), .B(b[285]), .Z(n572) );
  XOR U1437 ( .A(a[285]), .B(b[285]), .Z(n2504) );
  OR U1438 ( .A(a[284]), .B(b[284]), .Z(n570) );
  XOR U1439 ( .A(a[284]), .B(b[284]), .Z(n2502) );
  OR U1440 ( .A(a[283]), .B(b[283]), .Z(n568) );
  XOR U1441 ( .A(a[283]), .B(b[283]), .Z(n2500) );
  OR U1442 ( .A(a[282]), .B(b[282]), .Z(n566) );
  XOR U1443 ( .A(a[282]), .B(b[282]), .Z(n2498) );
  OR U1444 ( .A(a[281]), .B(b[281]), .Z(n564) );
  XOR U1445 ( .A(a[281]), .B(b[281]), .Z(n2496) );
  OR U1446 ( .A(a[280]), .B(b[280]), .Z(n562) );
  XOR U1447 ( .A(a[280]), .B(b[280]), .Z(n2494) );
  OR U1448 ( .A(a[279]), .B(b[279]), .Z(n560) );
  XOR U1449 ( .A(a[279]), .B(b[279]), .Z(n2490) );
  OR U1450 ( .A(a[278]), .B(b[278]), .Z(n558) );
  XOR U1451 ( .A(a[278]), .B(b[278]), .Z(n2488) );
  OR U1452 ( .A(a[277]), .B(b[277]), .Z(n556) );
  XOR U1453 ( .A(a[277]), .B(b[277]), .Z(n2486) );
  OR U1454 ( .A(a[276]), .B(b[276]), .Z(n554) );
  XOR U1455 ( .A(a[276]), .B(b[276]), .Z(n2484) );
  OR U1456 ( .A(a[275]), .B(b[275]), .Z(n552) );
  XOR U1457 ( .A(a[275]), .B(b[275]), .Z(n2482) );
  OR U1458 ( .A(a[274]), .B(b[274]), .Z(n550) );
  XOR U1459 ( .A(a[274]), .B(b[274]), .Z(n2480) );
  OR U1460 ( .A(a[273]), .B(b[273]), .Z(n548) );
  XOR U1461 ( .A(a[273]), .B(b[273]), .Z(n2478) );
  OR U1462 ( .A(a[272]), .B(b[272]), .Z(n546) );
  XOR U1463 ( .A(a[272]), .B(b[272]), .Z(n2476) );
  OR U1464 ( .A(a[271]), .B(b[271]), .Z(n544) );
  XOR U1465 ( .A(a[271]), .B(b[271]), .Z(n2474) );
  OR U1466 ( .A(a[270]), .B(b[270]), .Z(n542) );
  XOR U1467 ( .A(a[270]), .B(b[270]), .Z(n2472) );
  OR U1468 ( .A(a[269]), .B(b[269]), .Z(n540) );
  XOR U1469 ( .A(a[269]), .B(b[269]), .Z(n2468) );
  OR U1470 ( .A(a[268]), .B(b[268]), .Z(n538) );
  XOR U1471 ( .A(a[268]), .B(b[268]), .Z(n2466) );
  OR U1472 ( .A(a[267]), .B(b[267]), .Z(n536) );
  XOR U1473 ( .A(a[267]), .B(b[267]), .Z(n2464) );
  OR U1474 ( .A(a[266]), .B(b[266]), .Z(n534) );
  XOR U1475 ( .A(a[266]), .B(b[266]), .Z(n2462) );
  OR U1476 ( .A(a[265]), .B(b[265]), .Z(n532) );
  XOR U1477 ( .A(a[265]), .B(b[265]), .Z(n2460) );
  OR U1478 ( .A(a[264]), .B(b[264]), .Z(n530) );
  XOR U1479 ( .A(a[264]), .B(b[264]), .Z(n2458) );
  OR U1480 ( .A(a[263]), .B(b[263]), .Z(n528) );
  XOR U1481 ( .A(a[263]), .B(b[263]), .Z(n2456) );
  OR U1482 ( .A(a[262]), .B(b[262]), .Z(n526) );
  XOR U1483 ( .A(a[262]), .B(b[262]), .Z(n2454) );
  OR U1484 ( .A(a[261]), .B(b[261]), .Z(n524) );
  XOR U1485 ( .A(a[261]), .B(b[261]), .Z(n2452) );
  OR U1486 ( .A(a[260]), .B(b[260]), .Z(n522) );
  XOR U1487 ( .A(a[260]), .B(b[260]), .Z(n2450) );
  OR U1488 ( .A(a[259]), .B(b[259]), .Z(n520) );
  XOR U1489 ( .A(a[259]), .B(b[259]), .Z(n2446) );
  OR U1490 ( .A(a[258]), .B(b[258]), .Z(n518) );
  XOR U1491 ( .A(a[258]), .B(b[258]), .Z(n2444) );
  OR U1492 ( .A(a[257]), .B(b[257]), .Z(n516) );
  XOR U1493 ( .A(a[257]), .B(b[257]), .Z(n2442) );
  OR U1494 ( .A(a[256]), .B(b[256]), .Z(n514) );
  XOR U1495 ( .A(a[256]), .B(b[256]), .Z(n2440) );
  OR U1496 ( .A(a[255]), .B(b[255]), .Z(n512) );
  XOR U1497 ( .A(a[255]), .B(b[255]), .Z(n2438) );
  OR U1498 ( .A(a[254]), .B(b[254]), .Z(n510) );
  XOR U1499 ( .A(a[254]), .B(b[254]), .Z(n2436) );
  OR U1500 ( .A(a[253]), .B(b[253]), .Z(n508) );
  XOR U1501 ( .A(a[253]), .B(b[253]), .Z(n2434) );
  OR U1502 ( .A(a[252]), .B(b[252]), .Z(n506) );
  XOR U1503 ( .A(a[252]), .B(b[252]), .Z(n2432) );
  OR U1504 ( .A(a[251]), .B(b[251]), .Z(n504) );
  XOR U1505 ( .A(a[251]), .B(b[251]), .Z(n2430) );
  OR U1506 ( .A(a[250]), .B(b[250]), .Z(n502) );
  XOR U1507 ( .A(a[250]), .B(b[250]), .Z(n2428) );
  OR U1508 ( .A(a[249]), .B(b[249]), .Z(n500) );
  XOR U1509 ( .A(a[249]), .B(b[249]), .Z(n2424) );
  OR U1510 ( .A(a[248]), .B(b[248]), .Z(n498) );
  XOR U1511 ( .A(a[248]), .B(b[248]), .Z(n2422) );
  OR U1512 ( .A(a[247]), .B(b[247]), .Z(n496) );
  XOR U1513 ( .A(a[247]), .B(b[247]), .Z(n2420) );
  OR U1514 ( .A(a[246]), .B(b[246]), .Z(n494) );
  XOR U1515 ( .A(a[246]), .B(b[246]), .Z(n2418) );
  OR U1516 ( .A(a[245]), .B(b[245]), .Z(n492) );
  XOR U1517 ( .A(a[245]), .B(b[245]), .Z(n2416) );
  OR U1518 ( .A(a[244]), .B(b[244]), .Z(n490) );
  XOR U1519 ( .A(a[244]), .B(b[244]), .Z(n2414) );
  OR U1520 ( .A(a[243]), .B(b[243]), .Z(n488) );
  XOR U1521 ( .A(a[243]), .B(b[243]), .Z(n2412) );
  OR U1522 ( .A(a[242]), .B(b[242]), .Z(n486) );
  XOR U1523 ( .A(a[242]), .B(b[242]), .Z(n2410) );
  OR U1524 ( .A(a[241]), .B(b[241]), .Z(n484) );
  XOR U1525 ( .A(a[241]), .B(b[241]), .Z(n2408) );
  OR U1526 ( .A(a[240]), .B(b[240]), .Z(n482) );
  XOR U1527 ( .A(a[240]), .B(b[240]), .Z(n2406) );
  OR U1528 ( .A(a[239]), .B(b[239]), .Z(n480) );
  XOR U1529 ( .A(a[239]), .B(b[239]), .Z(n2402) );
  OR U1530 ( .A(a[238]), .B(b[238]), .Z(n478) );
  XOR U1531 ( .A(a[238]), .B(b[238]), .Z(n2400) );
  OR U1532 ( .A(a[237]), .B(b[237]), .Z(n476) );
  XOR U1533 ( .A(a[237]), .B(b[237]), .Z(n2398) );
  OR U1534 ( .A(a[236]), .B(b[236]), .Z(n474) );
  XOR U1535 ( .A(a[236]), .B(b[236]), .Z(n2396) );
  OR U1536 ( .A(a[235]), .B(b[235]), .Z(n472) );
  XOR U1537 ( .A(a[235]), .B(b[235]), .Z(n2394) );
  OR U1538 ( .A(a[234]), .B(b[234]), .Z(n470) );
  XOR U1539 ( .A(a[234]), .B(b[234]), .Z(n2392) );
  OR U1540 ( .A(a[233]), .B(b[233]), .Z(n468) );
  XOR U1541 ( .A(a[233]), .B(b[233]), .Z(n2390) );
  OR U1542 ( .A(a[232]), .B(b[232]), .Z(n466) );
  XOR U1543 ( .A(a[232]), .B(b[232]), .Z(n2388) );
  OR U1544 ( .A(a[231]), .B(b[231]), .Z(n464) );
  XOR U1545 ( .A(a[231]), .B(b[231]), .Z(n2386) );
  OR U1546 ( .A(a[230]), .B(b[230]), .Z(n462) );
  XOR U1547 ( .A(a[230]), .B(b[230]), .Z(n2384) );
  OR U1548 ( .A(a[229]), .B(b[229]), .Z(n460) );
  XOR U1549 ( .A(a[229]), .B(b[229]), .Z(n2380) );
  OR U1550 ( .A(a[228]), .B(b[228]), .Z(n458) );
  XOR U1551 ( .A(a[228]), .B(b[228]), .Z(n2378) );
  OR U1552 ( .A(a[227]), .B(b[227]), .Z(n456) );
  XOR U1553 ( .A(a[227]), .B(b[227]), .Z(n2376) );
  OR U1554 ( .A(a[226]), .B(b[226]), .Z(n454) );
  XOR U1555 ( .A(a[226]), .B(b[226]), .Z(n2374) );
  OR U1556 ( .A(a[225]), .B(b[225]), .Z(n452) );
  XOR U1557 ( .A(a[225]), .B(b[225]), .Z(n2372) );
  OR U1558 ( .A(a[224]), .B(b[224]), .Z(n450) );
  XOR U1559 ( .A(a[224]), .B(b[224]), .Z(n2370) );
  OR U1560 ( .A(a[223]), .B(b[223]), .Z(n448) );
  XOR U1561 ( .A(a[223]), .B(b[223]), .Z(n2368) );
  OR U1562 ( .A(a[222]), .B(b[222]), .Z(n446) );
  XOR U1563 ( .A(a[222]), .B(b[222]), .Z(n2366) );
  OR U1564 ( .A(a[221]), .B(b[221]), .Z(n444) );
  XOR U1565 ( .A(a[221]), .B(b[221]), .Z(n2364) );
  OR U1566 ( .A(a[220]), .B(b[220]), .Z(n442) );
  XOR U1567 ( .A(a[220]), .B(b[220]), .Z(n2362) );
  OR U1568 ( .A(a[219]), .B(b[219]), .Z(n440) );
  XOR U1569 ( .A(a[219]), .B(b[219]), .Z(n2358) );
  OR U1570 ( .A(a[218]), .B(b[218]), .Z(n438) );
  XOR U1571 ( .A(a[218]), .B(b[218]), .Z(n2356) );
  OR U1572 ( .A(a[217]), .B(b[217]), .Z(n436) );
  XOR U1573 ( .A(a[217]), .B(b[217]), .Z(n2354) );
  OR U1574 ( .A(a[216]), .B(b[216]), .Z(n434) );
  XOR U1575 ( .A(a[216]), .B(b[216]), .Z(n2352) );
  OR U1576 ( .A(a[215]), .B(b[215]), .Z(n432) );
  XOR U1577 ( .A(a[215]), .B(b[215]), .Z(n2350) );
  OR U1578 ( .A(a[214]), .B(b[214]), .Z(n430) );
  XOR U1579 ( .A(a[214]), .B(b[214]), .Z(n2348) );
  OR U1580 ( .A(a[213]), .B(b[213]), .Z(n428) );
  XOR U1581 ( .A(a[213]), .B(b[213]), .Z(n2346) );
  OR U1582 ( .A(a[212]), .B(b[212]), .Z(n426) );
  XOR U1583 ( .A(a[212]), .B(b[212]), .Z(n2344) );
  OR U1584 ( .A(a[211]), .B(b[211]), .Z(n424) );
  XOR U1585 ( .A(a[211]), .B(b[211]), .Z(n2342) );
  OR U1586 ( .A(a[210]), .B(b[210]), .Z(n422) );
  XOR U1587 ( .A(a[210]), .B(b[210]), .Z(n2340) );
  OR U1588 ( .A(a[209]), .B(b[209]), .Z(n420) );
  XOR U1589 ( .A(a[209]), .B(b[209]), .Z(n2336) );
  OR U1590 ( .A(a[208]), .B(b[208]), .Z(n418) );
  XOR U1591 ( .A(a[208]), .B(b[208]), .Z(n2334) );
  OR U1592 ( .A(a[207]), .B(b[207]), .Z(n416) );
  XOR U1593 ( .A(a[207]), .B(b[207]), .Z(n2332) );
  OR U1594 ( .A(a[206]), .B(b[206]), .Z(n414) );
  XOR U1595 ( .A(a[206]), .B(b[206]), .Z(n2330) );
  OR U1596 ( .A(a[205]), .B(b[205]), .Z(n412) );
  XOR U1597 ( .A(a[205]), .B(b[205]), .Z(n2328) );
  OR U1598 ( .A(a[204]), .B(b[204]), .Z(n410) );
  XOR U1599 ( .A(a[204]), .B(b[204]), .Z(n2326) );
  OR U1600 ( .A(a[203]), .B(b[203]), .Z(n408) );
  XOR U1601 ( .A(a[203]), .B(b[203]), .Z(n2324) );
  OR U1602 ( .A(a[202]), .B(b[202]), .Z(n406) );
  XOR U1603 ( .A(a[202]), .B(b[202]), .Z(n2322) );
  OR U1604 ( .A(a[201]), .B(b[201]), .Z(n404) );
  XOR U1605 ( .A(a[201]), .B(b[201]), .Z(n2320) );
  OR U1606 ( .A(a[200]), .B(b[200]), .Z(n402) );
  XOR U1607 ( .A(a[200]), .B(b[200]), .Z(n2318) );
  OR U1608 ( .A(a[199]), .B(b[199]), .Z(n400) );
  XOR U1609 ( .A(a[199]), .B(b[199]), .Z(n2312) );
  OR U1610 ( .A(a[198]), .B(b[198]), .Z(n398) );
  XOR U1611 ( .A(a[198]), .B(b[198]), .Z(n2310) );
  OR U1612 ( .A(a[197]), .B(b[197]), .Z(n396) );
  XOR U1613 ( .A(a[197]), .B(b[197]), .Z(n2308) );
  OR U1614 ( .A(a[196]), .B(b[196]), .Z(n394) );
  XOR U1615 ( .A(a[196]), .B(b[196]), .Z(n2306) );
  OR U1616 ( .A(a[195]), .B(b[195]), .Z(n392) );
  XOR U1617 ( .A(a[195]), .B(b[195]), .Z(n2304) );
  OR U1618 ( .A(a[194]), .B(b[194]), .Z(n390) );
  XOR U1619 ( .A(a[194]), .B(b[194]), .Z(n2302) );
  OR U1620 ( .A(a[193]), .B(b[193]), .Z(n388) );
  XOR U1621 ( .A(a[193]), .B(b[193]), .Z(n2300) );
  OR U1622 ( .A(a[192]), .B(b[192]), .Z(n386) );
  XOR U1623 ( .A(a[192]), .B(b[192]), .Z(n2298) );
  OR U1624 ( .A(a[191]), .B(b[191]), .Z(n384) );
  XOR U1625 ( .A(a[191]), .B(b[191]), .Z(n2296) );
  OR U1626 ( .A(a[190]), .B(b[190]), .Z(n382) );
  XOR U1627 ( .A(a[190]), .B(b[190]), .Z(n2294) );
  OR U1628 ( .A(a[189]), .B(b[189]), .Z(n380) );
  XOR U1629 ( .A(a[189]), .B(b[189]), .Z(n2290) );
  OR U1630 ( .A(a[188]), .B(b[188]), .Z(n378) );
  XOR U1631 ( .A(a[188]), .B(b[188]), .Z(n2288) );
  OR U1632 ( .A(a[187]), .B(b[187]), .Z(n376) );
  XOR U1633 ( .A(a[187]), .B(b[187]), .Z(n2286) );
  OR U1634 ( .A(a[186]), .B(b[186]), .Z(n374) );
  XOR U1635 ( .A(a[186]), .B(b[186]), .Z(n2284) );
  OR U1636 ( .A(a[185]), .B(b[185]), .Z(n372) );
  XOR U1637 ( .A(a[185]), .B(b[185]), .Z(n2282) );
  OR U1638 ( .A(a[184]), .B(b[184]), .Z(n370) );
  XOR U1639 ( .A(a[184]), .B(b[184]), .Z(n2280) );
  OR U1640 ( .A(a[183]), .B(b[183]), .Z(n368) );
  XOR U1641 ( .A(a[183]), .B(b[183]), .Z(n2278) );
  OR U1642 ( .A(a[182]), .B(b[182]), .Z(n366) );
  XOR U1643 ( .A(a[182]), .B(b[182]), .Z(n2276) );
  OR U1644 ( .A(a[181]), .B(b[181]), .Z(n364) );
  XOR U1645 ( .A(a[181]), .B(b[181]), .Z(n2274) );
  OR U1646 ( .A(a[180]), .B(b[180]), .Z(n362) );
  XOR U1647 ( .A(a[180]), .B(b[180]), .Z(n2272) );
  OR U1648 ( .A(a[179]), .B(b[179]), .Z(n360) );
  XOR U1649 ( .A(a[179]), .B(b[179]), .Z(n2268) );
  OR U1650 ( .A(a[178]), .B(b[178]), .Z(n358) );
  XOR U1651 ( .A(a[178]), .B(b[178]), .Z(n2266) );
  OR U1652 ( .A(a[177]), .B(b[177]), .Z(n356) );
  XOR U1653 ( .A(a[177]), .B(b[177]), .Z(n2264) );
  OR U1654 ( .A(a[176]), .B(b[176]), .Z(n354) );
  XOR U1655 ( .A(a[176]), .B(b[176]), .Z(n2262) );
  OR U1656 ( .A(a[175]), .B(b[175]), .Z(n352) );
  XOR U1657 ( .A(a[175]), .B(b[175]), .Z(n2260) );
  OR U1658 ( .A(a[174]), .B(b[174]), .Z(n350) );
  XOR U1659 ( .A(a[174]), .B(b[174]), .Z(n2258) );
  OR U1660 ( .A(a[173]), .B(b[173]), .Z(n348) );
  XOR U1661 ( .A(a[173]), .B(b[173]), .Z(n2256) );
  OR U1662 ( .A(a[172]), .B(b[172]), .Z(n346) );
  XOR U1663 ( .A(a[172]), .B(b[172]), .Z(n2254) );
  OR U1664 ( .A(a[171]), .B(b[171]), .Z(n344) );
  XOR U1665 ( .A(a[171]), .B(b[171]), .Z(n2252) );
  OR U1666 ( .A(a[170]), .B(b[170]), .Z(n342) );
  XOR U1667 ( .A(a[170]), .B(b[170]), .Z(n2250) );
  OR U1668 ( .A(a[169]), .B(b[169]), .Z(n340) );
  XOR U1669 ( .A(a[169]), .B(b[169]), .Z(n2246) );
  OR U1670 ( .A(a[168]), .B(b[168]), .Z(n338) );
  XOR U1671 ( .A(a[168]), .B(b[168]), .Z(n2244) );
  OR U1672 ( .A(a[167]), .B(b[167]), .Z(n336) );
  XOR U1673 ( .A(a[167]), .B(b[167]), .Z(n2242) );
  OR U1674 ( .A(a[166]), .B(b[166]), .Z(n334) );
  XOR U1675 ( .A(a[166]), .B(b[166]), .Z(n2240) );
  OR U1676 ( .A(a[165]), .B(b[165]), .Z(n332) );
  XOR U1677 ( .A(a[165]), .B(b[165]), .Z(n2238) );
  OR U1678 ( .A(a[164]), .B(b[164]), .Z(n330) );
  XOR U1679 ( .A(a[164]), .B(b[164]), .Z(n2236) );
  OR U1680 ( .A(a[163]), .B(b[163]), .Z(n328) );
  XOR U1681 ( .A(a[163]), .B(b[163]), .Z(n2234) );
  OR U1682 ( .A(a[162]), .B(b[162]), .Z(n326) );
  XOR U1683 ( .A(a[162]), .B(b[162]), .Z(n2232) );
  OR U1684 ( .A(a[161]), .B(b[161]), .Z(n324) );
  XOR U1685 ( .A(a[161]), .B(b[161]), .Z(n2230) );
  OR U1686 ( .A(a[160]), .B(b[160]), .Z(n322) );
  XOR U1687 ( .A(a[160]), .B(b[160]), .Z(n2228) );
  OR U1688 ( .A(a[159]), .B(b[159]), .Z(n320) );
  XOR U1689 ( .A(a[159]), .B(b[159]), .Z(n2224) );
  OR U1690 ( .A(a[158]), .B(b[158]), .Z(n318) );
  XOR U1691 ( .A(a[158]), .B(b[158]), .Z(n2222) );
  OR U1692 ( .A(a[157]), .B(b[157]), .Z(n316) );
  XOR U1693 ( .A(a[157]), .B(b[157]), .Z(n2220) );
  OR U1694 ( .A(a[156]), .B(b[156]), .Z(n314) );
  XOR U1695 ( .A(a[156]), .B(b[156]), .Z(n2218) );
  OR U1696 ( .A(a[155]), .B(b[155]), .Z(n312) );
  XOR U1697 ( .A(a[155]), .B(b[155]), .Z(n2216) );
  OR U1698 ( .A(a[154]), .B(b[154]), .Z(n310) );
  XOR U1699 ( .A(a[154]), .B(b[154]), .Z(n2214) );
  OR U1700 ( .A(a[153]), .B(b[153]), .Z(n308) );
  XOR U1701 ( .A(a[153]), .B(b[153]), .Z(n2212) );
  OR U1702 ( .A(a[152]), .B(b[152]), .Z(n306) );
  XOR U1703 ( .A(a[152]), .B(b[152]), .Z(n2210) );
  OR U1704 ( .A(a[151]), .B(b[151]), .Z(n304) );
  XOR U1705 ( .A(a[151]), .B(b[151]), .Z(n2208) );
  OR U1706 ( .A(a[150]), .B(b[150]), .Z(n302) );
  XOR U1707 ( .A(a[150]), .B(b[150]), .Z(n2206) );
  OR U1708 ( .A(a[149]), .B(b[149]), .Z(n300) );
  XOR U1709 ( .A(a[149]), .B(b[149]), .Z(n2202) );
  OR U1710 ( .A(a[148]), .B(b[148]), .Z(n298) );
  XOR U1711 ( .A(a[148]), .B(b[148]), .Z(n2200) );
  OR U1712 ( .A(a[147]), .B(b[147]), .Z(n296) );
  XOR U1713 ( .A(a[147]), .B(b[147]), .Z(n2198) );
  OR U1714 ( .A(a[146]), .B(b[146]), .Z(n294) );
  XOR U1715 ( .A(a[146]), .B(b[146]), .Z(n2196) );
  OR U1716 ( .A(a[145]), .B(b[145]), .Z(n292) );
  XOR U1717 ( .A(a[145]), .B(b[145]), .Z(n2194) );
  OR U1718 ( .A(a[144]), .B(b[144]), .Z(n290) );
  XOR U1719 ( .A(a[144]), .B(b[144]), .Z(n2192) );
  OR U1720 ( .A(a[143]), .B(b[143]), .Z(n288) );
  XOR U1721 ( .A(a[143]), .B(b[143]), .Z(n2190) );
  OR U1722 ( .A(a[142]), .B(b[142]), .Z(n286) );
  XOR U1723 ( .A(a[142]), .B(b[142]), .Z(n2188) );
  OR U1724 ( .A(a[141]), .B(b[141]), .Z(n284) );
  XOR U1725 ( .A(a[141]), .B(b[141]), .Z(n2186) );
  OR U1726 ( .A(a[140]), .B(b[140]), .Z(n282) );
  XOR U1727 ( .A(a[140]), .B(b[140]), .Z(n2184) );
  OR U1728 ( .A(a[139]), .B(b[139]), .Z(n280) );
  XOR U1729 ( .A(a[139]), .B(b[139]), .Z(n2180) );
  OR U1730 ( .A(a[138]), .B(b[138]), .Z(n278) );
  XOR U1731 ( .A(a[138]), .B(b[138]), .Z(n2178) );
  OR U1732 ( .A(a[137]), .B(b[137]), .Z(n276) );
  XOR U1733 ( .A(a[137]), .B(b[137]), .Z(n2176) );
  OR U1734 ( .A(a[136]), .B(b[136]), .Z(n274) );
  XOR U1735 ( .A(a[136]), .B(b[136]), .Z(n2174) );
  OR U1736 ( .A(a[135]), .B(b[135]), .Z(n272) );
  XOR U1737 ( .A(a[135]), .B(b[135]), .Z(n2172) );
  OR U1738 ( .A(a[134]), .B(b[134]), .Z(n270) );
  XOR U1739 ( .A(a[134]), .B(b[134]), .Z(n2170) );
  OR U1740 ( .A(a[133]), .B(b[133]), .Z(n268) );
  XOR U1741 ( .A(a[133]), .B(b[133]), .Z(n2168) );
  OR U1742 ( .A(a[132]), .B(b[132]), .Z(n266) );
  XOR U1743 ( .A(a[132]), .B(b[132]), .Z(n2166) );
  OR U1744 ( .A(a[131]), .B(b[131]), .Z(n264) );
  XOR U1745 ( .A(a[131]), .B(b[131]), .Z(n2164) );
  OR U1746 ( .A(a[130]), .B(b[130]), .Z(n262) );
  XOR U1747 ( .A(a[130]), .B(b[130]), .Z(n2162) );
  OR U1748 ( .A(a[129]), .B(b[129]), .Z(n260) );
  XOR U1749 ( .A(a[129]), .B(b[129]), .Z(n2158) );
  OR U1750 ( .A(a[128]), .B(b[128]), .Z(n258) );
  XOR U1751 ( .A(a[128]), .B(b[128]), .Z(n2156) );
  OR U1752 ( .A(a[127]), .B(b[127]), .Z(n256) );
  XOR U1753 ( .A(a[127]), .B(b[127]), .Z(n2154) );
  OR U1754 ( .A(a[126]), .B(b[126]), .Z(n254) );
  XOR U1755 ( .A(a[126]), .B(b[126]), .Z(n2152) );
  OR U1756 ( .A(a[125]), .B(b[125]), .Z(n252) );
  XOR U1757 ( .A(a[125]), .B(b[125]), .Z(n2150) );
  OR U1758 ( .A(a[124]), .B(b[124]), .Z(n250) );
  XOR U1759 ( .A(a[124]), .B(b[124]), .Z(n2148) );
  OR U1760 ( .A(a[123]), .B(b[123]), .Z(n248) );
  XOR U1761 ( .A(a[123]), .B(b[123]), .Z(n2146) );
  OR U1762 ( .A(a[122]), .B(b[122]), .Z(n246) );
  XOR U1763 ( .A(a[122]), .B(b[122]), .Z(n2144) );
  OR U1764 ( .A(a[121]), .B(b[121]), .Z(n244) );
  XOR U1765 ( .A(a[121]), .B(b[121]), .Z(n2142) );
  OR U1766 ( .A(a[120]), .B(b[120]), .Z(n242) );
  XOR U1767 ( .A(a[120]), .B(b[120]), .Z(n2140) );
  OR U1768 ( .A(a[119]), .B(b[119]), .Z(n240) );
  XOR U1769 ( .A(a[119]), .B(b[119]), .Z(n2136) );
  OR U1770 ( .A(a[118]), .B(b[118]), .Z(n238) );
  XOR U1771 ( .A(a[118]), .B(b[118]), .Z(n2134) );
  OR U1772 ( .A(a[117]), .B(b[117]), .Z(n236) );
  XOR U1773 ( .A(a[117]), .B(b[117]), .Z(n2132) );
  OR U1774 ( .A(a[116]), .B(b[116]), .Z(n234) );
  XOR U1775 ( .A(a[116]), .B(b[116]), .Z(n2130) );
  OR U1776 ( .A(a[115]), .B(b[115]), .Z(n232) );
  XOR U1777 ( .A(a[115]), .B(b[115]), .Z(n2128) );
  OR U1778 ( .A(a[114]), .B(b[114]), .Z(n230) );
  XOR U1779 ( .A(a[114]), .B(b[114]), .Z(n2126) );
  OR U1780 ( .A(a[113]), .B(b[113]), .Z(n228) );
  XOR U1781 ( .A(a[113]), .B(b[113]), .Z(n2124) );
  OR U1782 ( .A(a[112]), .B(b[112]), .Z(n226) );
  XOR U1783 ( .A(a[112]), .B(b[112]), .Z(n2122) );
  OR U1784 ( .A(a[111]), .B(b[111]), .Z(n224) );
  XOR U1785 ( .A(a[111]), .B(b[111]), .Z(n2120) );
  OR U1786 ( .A(a[110]), .B(b[110]), .Z(n222) );
  XOR U1787 ( .A(a[110]), .B(b[110]), .Z(n2118) );
  OR U1788 ( .A(a[109]), .B(b[109]), .Z(n220) );
  XOR U1789 ( .A(a[109]), .B(b[109]), .Z(n2114) );
  OR U1790 ( .A(a[108]), .B(b[108]), .Z(n218) );
  XOR U1791 ( .A(a[108]), .B(b[108]), .Z(n2112) );
  OR U1792 ( .A(a[107]), .B(b[107]), .Z(n216) );
  XOR U1793 ( .A(a[107]), .B(b[107]), .Z(n2110) );
  OR U1794 ( .A(a[106]), .B(b[106]), .Z(n214) );
  XOR U1795 ( .A(a[106]), .B(b[106]), .Z(n2108) );
  OR U1796 ( .A(a[105]), .B(b[105]), .Z(n212) );
  XOR U1797 ( .A(a[105]), .B(b[105]), .Z(n2106) );
  OR U1798 ( .A(a[104]), .B(b[104]), .Z(n210) );
  XOR U1799 ( .A(a[104]), .B(b[104]), .Z(n2104) );
  OR U1800 ( .A(a[103]), .B(b[103]), .Z(n208) );
  XOR U1801 ( .A(a[103]), .B(b[103]), .Z(n2102) );
  OR U1802 ( .A(a[102]), .B(b[102]), .Z(n206) );
  XOR U1803 ( .A(a[102]), .B(b[102]), .Z(n2100) );
  OR U1804 ( .A(a[101]), .B(b[101]), .Z(n204) );
  XOR U1805 ( .A(a[101]), .B(b[101]), .Z(n2080) );
  OR U1806 ( .A(a[100]), .B(b[100]), .Z(n202) );
  XOR U1807 ( .A(a[100]), .B(b[100]), .Z(n2038) );
  OR U1808 ( .A(a[99]), .B(b[99]), .Z(n200) );
  XOR U1809 ( .A(a[99]), .B(b[99]), .Z(n4090) );
  OR U1810 ( .A(a[98]), .B(b[98]), .Z(n198) );
  XOR U1811 ( .A(a[98]), .B(b[98]), .Z(n4068) );
  OR U1812 ( .A(a[97]), .B(b[97]), .Z(n196) );
  XOR U1813 ( .A(a[97]), .B(b[97]), .Z(n4046) );
  OR U1814 ( .A(a[96]), .B(b[96]), .Z(n194) );
  XOR U1815 ( .A(a[96]), .B(b[96]), .Z(n4024) );
  OR U1816 ( .A(a[95]), .B(b[95]), .Z(n192) );
  XOR U1817 ( .A(a[95]), .B(b[95]), .Z(n4002) );
  OR U1818 ( .A(a[94]), .B(b[94]), .Z(n190) );
  XOR U1819 ( .A(a[94]), .B(b[94]), .Z(n3980) );
  OR U1820 ( .A(a[93]), .B(b[93]), .Z(n188) );
  XOR U1821 ( .A(a[93]), .B(b[93]), .Z(n3958) );
  OR U1822 ( .A(a[92]), .B(b[92]), .Z(n186) );
  XOR U1823 ( .A(a[92]), .B(b[92]), .Z(n3936) );
  OR U1824 ( .A(a[91]), .B(b[91]), .Z(n184) );
  XOR U1825 ( .A(a[91]), .B(b[91]), .Z(n3914) );
  OR U1826 ( .A(a[90]), .B(b[90]), .Z(n182) );
  XOR U1827 ( .A(a[90]), .B(b[90]), .Z(n3892) );
  OR U1828 ( .A(a[89]), .B(b[89]), .Z(n180) );
  XOR U1829 ( .A(a[89]), .B(b[89]), .Z(n3868) );
  OR U1830 ( .A(a[88]), .B(b[88]), .Z(n178) );
  XOR U1831 ( .A(a[88]), .B(b[88]), .Z(n3846) );
  OR U1832 ( .A(a[87]), .B(b[87]), .Z(n176) );
  XOR U1833 ( .A(a[87]), .B(b[87]), .Z(n3824) );
  OR U1834 ( .A(a[86]), .B(b[86]), .Z(n174) );
  XOR U1835 ( .A(a[86]), .B(b[86]), .Z(n3802) );
  OR U1836 ( .A(a[85]), .B(b[85]), .Z(n172) );
  XOR U1837 ( .A(a[85]), .B(b[85]), .Z(n3780) );
  OR U1838 ( .A(a[84]), .B(b[84]), .Z(n170) );
  XOR U1839 ( .A(a[84]), .B(b[84]), .Z(n3758) );
  OR U1840 ( .A(a[83]), .B(b[83]), .Z(n168) );
  XOR U1841 ( .A(a[83]), .B(b[83]), .Z(n3736) );
  OR U1842 ( .A(a[82]), .B(b[82]), .Z(n166) );
  XOR U1843 ( .A(a[82]), .B(b[82]), .Z(n3714) );
  OR U1844 ( .A(a[81]), .B(b[81]), .Z(n164) );
  XOR U1845 ( .A(a[81]), .B(b[81]), .Z(n3692) );
  OR U1846 ( .A(a[80]), .B(b[80]), .Z(n162) );
  XOR U1847 ( .A(a[80]), .B(b[80]), .Z(n3670) );
  OR U1848 ( .A(a[79]), .B(b[79]), .Z(n160) );
  XOR U1849 ( .A(a[79]), .B(b[79]), .Z(n3646) );
  OR U1850 ( .A(a[78]), .B(b[78]), .Z(n158) );
  XOR U1851 ( .A(a[78]), .B(b[78]), .Z(n3624) );
  OR U1852 ( .A(a[77]), .B(b[77]), .Z(n156) );
  XOR U1853 ( .A(a[77]), .B(b[77]), .Z(n3602) );
  OR U1854 ( .A(a[76]), .B(b[76]), .Z(n154) );
  XOR U1855 ( .A(a[76]), .B(b[76]), .Z(n3580) );
  OR U1856 ( .A(a[75]), .B(b[75]), .Z(n152) );
  XOR U1857 ( .A(a[75]), .B(b[75]), .Z(n3558) );
  OR U1858 ( .A(a[74]), .B(b[74]), .Z(n150) );
  XOR U1859 ( .A(a[74]), .B(b[74]), .Z(n3536) );
  OR U1860 ( .A(a[73]), .B(b[73]), .Z(n148) );
  XOR U1861 ( .A(a[73]), .B(b[73]), .Z(n3514) );
  OR U1862 ( .A(a[72]), .B(b[72]), .Z(n146) );
  XOR U1863 ( .A(a[72]), .B(b[72]), .Z(n3492) );
  OR U1864 ( .A(a[71]), .B(b[71]), .Z(n144) );
  XOR U1865 ( .A(a[71]), .B(b[71]), .Z(n3470) );
  OR U1866 ( .A(a[70]), .B(b[70]), .Z(n142) );
  XOR U1867 ( .A(a[70]), .B(b[70]), .Z(n3448) );
  OR U1868 ( .A(a[69]), .B(b[69]), .Z(n140) );
  XOR U1869 ( .A(a[69]), .B(b[69]), .Z(n3424) );
  OR U1870 ( .A(a[68]), .B(b[68]), .Z(n138) );
  XOR U1871 ( .A(a[68]), .B(b[68]), .Z(n3402) );
  OR U1872 ( .A(a[67]), .B(b[67]), .Z(n136) );
  XOR U1873 ( .A(a[67]), .B(b[67]), .Z(n3380) );
  OR U1874 ( .A(a[66]), .B(b[66]), .Z(n134) );
  XOR U1875 ( .A(a[66]), .B(b[66]), .Z(n3358) );
  OR U1876 ( .A(a[65]), .B(b[65]), .Z(n132) );
  XOR U1877 ( .A(a[65]), .B(b[65]), .Z(n3336) );
  OR U1878 ( .A(a[64]), .B(b[64]), .Z(n130) );
  XOR U1879 ( .A(a[64]), .B(b[64]), .Z(n3314) );
  OR U1880 ( .A(a[63]), .B(b[63]), .Z(n128) );
  XOR U1881 ( .A(a[63]), .B(b[63]), .Z(n3292) );
  OR U1882 ( .A(a[62]), .B(b[62]), .Z(n126) );
  XOR U1883 ( .A(a[62]), .B(b[62]), .Z(n3270) );
  OR U1884 ( .A(a[61]), .B(b[61]), .Z(n124) );
  XOR U1885 ( .A(a[61]), .B(b[61]), .Z(n3248) );
  OR U1886 ( .A(a[60]), .B(b[60]), .Z(n122) );
  XOR U1887 ( .A(a[60]), .B(b[60]), .Z(n3226) );
  OR U1888 ( .A(a[59]), .B(b[59]), .Z(n120) );
  XOR U1889 ( .A(a[59]), .B(b[59]), .Z(n3202) );
  OR U1890 ( .A(a[58]), .B(b[58]), .Z(n118) );
  XOR U1891 ( .A(a[58]), .B(b[58]), .Z(n3180) );
  OR U1892 ( .A(a[57]), .B(b[57]), .Z(n116) );
  XOR U1893 ( .A(a[57]), .B(b[57]), .Z(n3158) );
  OR U1894 ( .A(a[56]), .B(b[56]), .Z(n114) );
  XOR U1895 ( .A(a[56]), .B(b[56]), .Z(n3136) );
  OR U1896 ( .A(a[55]), .B(b[55]), .Z(n112) );
  XOR U1897 ( .A(a[55]), .B(b[55]), .Z(n3114) );
  OR U1898 ( .A(a[54]), .B(b[54]), .Z(n110) );
  XOR U1899 ( .A(a[54]), .B(b[54]), .Z(n3092) );
  OR U1900 ( .A(a[53]), .B(b[53]), .Z(n108) );
  XOR U1901 ( .A(a[53]), .B(b[53]), .Z(n3070) );
  OR U1902 ( .A(a[52]), .B(b[52]), .Z(n106) );
  XOR U1903 ( .A(a[52]), .B(b[52]), .Z(n3048) );
  OR U1904 ( .A(a[51]), .B(b[51]), .Z(n104) );
  XOR U1905 ( .A(a[51]), .B(b[51]), .Z(n3026) );
  OR U1906 ( .A(a[50]), .B(b[50]), .Z(n102) );
  XOR U1907 ( .A(a[50]), .B(b[50]), .Z(n3004) );
  OR U1908 ( .A(a[49]), .B(b[49]), .Z(n100) );
  XOR U1909 ( .A(a[49]), .B(b[49]), .Z(n2980) );
  OR U1910 ( .A(a[48]), .B(b[48]), .Z(n98) );
  XOR U1911 ( .A(a[48]), .B(b[48]), .Z(n2958) );
  OR U1912 ( .A(a[47]), .B(b[47]), .Z(n96) );
  XOR U1913 ( .A(a[47]), .B(b[47]), .Z(n2936) );
  OR U1914 ( .A(a[46]), .B(b[46]), .Z(n94) );
  XOR U1915 ( .A(a[46]), .B(b[46]), .Z(n2914) );
  OR U1916 ( .A(a[45]), .B(b[45]), .Z(n92) );
  XOR U1917 ( .A(a[45]), .B(b[45]), .Z(n2892) );
  OR U1918 ( .A(a[44]), .B(b[44]), .Z(n90) );
  XOR U1919 ( .A(a[44]), .B(b[44]), .Z(n2870) );
  OR U1920 ( .A(a[43]), .B(b[43]), .Z(n88) );
  XOR U1921 ( .A(a[43]), .B(b[43]), .Z(n2848) );
  OR U1922 ( .A(a[42]), .B(b[42]), .Z(n86) );
  XOR U1923 ( .A(a[42]), .B(b[42]), .Z(n2826) );
  OR U1924 ( .A(a[41]), .B(b[41]), .Z(n84) );
  XOR U1925 ( .A(a[41]), .B(b[41]), .Z(n2804) );
  OR U1926 ( .A(a[40]), .B(b[40]), .Z(n82) );
  XOR U1927 ( .A(a[40]), .B(b[40]), .Z(n2782) );
  OR U1928 ( .A(a[39]), .B(b[39]), .Z(n80) );
  XOR U1929 ( .A(a[39]), .B(b[39]), .Z(n2758) );
  OR U1930 ( .A(a[38]), .B(b[38]), .Z(n78) );
  XOR U1931 ( .A(a[38]), .B(b[38]), .Z(n2736) );
  OR U1932 ( .A(a[37]), .B(b[37]), .Z(n76) );
  XOR U1933 ( .A(a[37]), .B(b[37]), .Z(n2714) );
  OR U1934 ( .A(a[36]), .B(b[36]), .Z(n74) );
  XOR U1935 ( .A(a[36]), .B(b[36]), .Z(n2692) );
  OR U1936 ( .A(a[35]), .B(b[35]), .Z(n72) );
  XOR U1937 ( .A(a[35]), .B(b[35]), .Z(n2670) );
  OR U1938 ( .A(a[34]), .B(b[34]), .Z(n70) );
  XOR U1939 ( .A(a[34]), .B(b[34]), .Z(n2648) );
  OR U1940 ( .A(a[33]), .B(b[33]), .Z(n68) );
  XOR U1941 ( .A(a[33]), .B(b[33]), .Z(n2626) );
  OR U1942 ( .A(a[32]), .B(b[32]), .Z(n66) );
  XOR U1943 ( .A(a[32]), .B(b[32]), .Z(n2604) );
  OR U1944 ( .A(a[31]), .B(b[31]), .Z(n64) );
  XOR U1945 ( .A(a[31]), .B(b[31]), .Z(n2582) );
  OR U1946 ( .A(a[30]), .B(b[30]), .Z(n62) );
  XOR U1947 ( .A(a[30]), .B(b[30]), .Z(n2560) );
  OR U1948 ( .A(a[29]), .B(b[29]), .Z(n60) );
  XOR U1949 ( .A(a[29]), .B(b[29]), .Z(n2536) );
  OR U1950 ( .A(a[28]), .B(b[28]), .Z(n58) );
  XOR U1951 ( .A(a[28]), .B(b[28]), .Z(n2514) );
  OR U1952 ( .A(a[27]), .B(b[27]), .Z(n56) );
  XOR U1953 ( .A(a[27]), .B(b[27]), .Z(n2492) );
  OR U1954 ( .A(a[26]), .B(b[26]), .Z(n54) );
  XOR U1955 ( .A(a[26]), .B(b[26]), .Z(n2470) );
  OR U1956 ( .A(a[25]), .B(b[25]), .Z(n52) );
  XOR U1957 ( .A(a[25]), .B(b[25]), .Z(n2448) );
  OR U1958 ( .A(a[24]), .B(b[24]), .Z(n50) );
  XOR U1959 ( .A(a[24]), .B(b[24]), .Z(n2426) );
  OR U1960 ( .A(a[23]), .B(b[23]), .Z(n48) );
  XOR U1961 ( .A(a[23]), .B(b[23]), .Z(n2404) );
  OR U1962 ( .A(a[22]), .B(b[22]), .Z(n46) );
  XOR U1963 ( .A(a[22]), .B(b[22]), .Z(n2382) );
  OR U1964 ( .A(a[21]), .B(b[21]), .Z(n44) );
  XOR U1965 ( .A(a[21]), .B(b[21]), .Z(n2360) );
  OR U1966 ( .A(a[20]), .B(b[20]), .Z(n42) );
  XOR U1967 ( .A(a[20]), .B(b[20]), .Z(n2338) );
  OR U1968 ( .A(a[19]), .B(b[19]), .Z(n40) );
  XOR U1969 ( .A(a[19]), .B(b[19]), .Z(n2314) );
  OR U1970 ( .A(a[18]), .B(b[18]), .Z(n38) );
  XOR U1971 ( .A(a[18]), .B(b[18]), .Z(n2292) );
  OR U1972 ( .A(a[17]), .B(b[17]), .Z(n36) );
  XOR U1973 ( .A(a[17]), .B(b[17]), .Z(n2270) );
  OR U1974 ( .A(a[16]), .B(b[16]), .Z(n34) );
  XOR U1975 ( .A(a[16]), .B(b[16]), .Z(n2248) );
  OR U1976 ( .A(a[15]), .B(b[15]), .Z(n32) );
  XOR U1977 ( .A(a[15]), .B(b[15]), .Z(n2226) );
  OR U1978 ( .A(a[14]), .B(b[14]), .Z(n30) );
  XOR U1979 ( .A(a[14]), .B(b[14]), .Z(n2204) );
  OR U1980 ( .A(a[13]), .B(b[13]), .Z(n28) );
  XOR U1981 ( .A(a[13]), .B(b[13]), .Z(n2182) );
  OR U1982 ( .A(a[12]), .B(b[12]), .Z(n26) );
  XOR U1983 ( .A(a[12]), .B(b[12]), .Z(n2160) );
  OR U1984 ( .A(a[11]), .B(b[11]), .Z(n24) );
  XOR U1985 ( .A(a[11]), .B(b[11]), .Z(n2138) );
  OR U1986 ( .A(a[10]), .B(b[10]), .Z(n22) );
  XOR U1987 ( .A(a[10]), .B(b[10]), .Z(n2116) );
  OR U1988 ( .A(a[9]), .B(b[9]), .Z(n20) );
  XOR U1989 ( .A(a[9]), .B(b[9]), .Z(n4092) );
  OR U1990 ( .A(a[8]), .B(b[8]), .Z(n18) );
  XOR U1991 ( .A(a[8]), .B(b[8]), .Z(n3870) );
  OR U1992 ( .A(a[7]), .B(b[7]), .Z(n16) );
  XOR U1993 ( .A(a[7]), .B(b[7]), .Z(n3648) );
  OR U1994 ( .A(a[6]), .B(b[6]), .Z(n14) );
  XOR U1995 ( .A(a[6]), .B(b[6]), .Z(n3426) );
  OR U1996 ( .A(a[5]), .B(b[5]), .Z(n12) );
  XOR U1997 ( .A(a[5]), .B(b[5]), .Z(n3204) );
  OR U1998 ( .A(a[4]), .B(b[4]), .Z(n10) );
  NAND U1999 ( .A(b[3]), .B(a[3]), .Z(n8) );
  XOR U2000 ( .A(b[3]), .B(a[3]), .Z(n2760) );
  NAND U2001 ( .A(b[2]), .B(a[2]), .Z(n6) );
  NAND U2002 ( .A(a[0]), .B(b[0]), .Z(n2316) );
  XOR U2003 ( .A(b[2]), .B(a[2]), .Z(n2537) );
  NANDN U2004 ( .A(n2538), .B(n2537), .Z(n5) );
  NAND U2005 ( .A(n6), .B(n5), .Z(n2759) );
  NAND U2006 ( .A(n2760), .B(n2759), .Z(n7) );
  AND U2007 ( .A(n8), .B(n7), .Z(n2982) );
  XOR U2008 ( .A(a[4]), .B(b[4]), .Z(n2981) );
  NAND U2009 ( .A(n2982), .B(n2981), .Z(n9) );
  NAND U2010 ( .A(n10), .B(n9), .Z(n3203) );
  NAND U2011 ( .A(n3204), .B(n3203), .Z(n11) );
  NAND U2012 ( .A(n12), .B(n11), .Z(n3425) );
  NAND U2013 ( .A(n3426), .B(n3425), .Z(n13) );
  NAND U2014 ( .A(n14), .B(n13), .Z(n3647) );
  NAND U2015 ( .A(n3648), .B(n3647), .Z(n15) );
  NAND U2016 ( .A(n16), .B(n15), .Z(n3869) );
  NAND U2017 ( .A(n3870), .B(n3869), .Z(n17) );
  NAND U2018 ( .A(n18), .B(n17), .Z(n4091) );
  NAND U2019 ( .A(n4092), .B(n4091), .Z(n19) );
  NAND U2020 ( .A(n20), .B(n19), .Z(n2115) );
  NAND U2021 ( .A(n2116), .B(n2115), .Z(n21) );
  NAND U2022 ( .A(n22), .B(n21), .Z(n2137) );
  NAND U2023 ( .A(n2138), .B(n2137), .Z(n23) );
  NAND U2024 ( .A(n24), .B(n23), .Z(n2159) );
  NAND U2025 ( .A(n2160), .B(n2159), .Z(n25) );
  NAND U2026 ( .A(n26), .B(n25), .Z(n2181) );
  NAND U2027 ( .A(n2182), .B(n2181), .Z(n27) );
  NAND U2028 ( .A(n28), .B(n27), .Z(n2203) );
  NAND U2029 ( .A(n2204), .B(n2203), .Z(n29) );
  NAND U2030 ( .A(n30), .B(n29), .Z(n2225) );
  NAND U2031 ( .A(n2226), .B(n2225), .Z(n31) );
  NAND U2032 ( .A(n32), .B(n31), .Z(n2247) );
  NAND U2033 ( .A(n2248), .B(n2247), .Z(n33) );
  NAND U2034 ( .A(n34), .B(n33), .Z(n2269) );
  NAND U2035 ( .A(n2270), .B(n2269), .Z(n35) );
  NAND U2036 ( .A(n36), .B(n35), .Z(n2291) );
  NAND U2037 ( .A(n2292), .B(n2291), .Z(n37) );
  NAND U2038 ( .A(n38), .B(n37), .Z(n2313) );
  NAND U2039 ( .A(n2314), .B(n2313), .Z(n39) );
  NAND U2040 ( .A(n40), .B(n39), .Z(n2337) );
  NAND U2041 ( .A(n2338), .B(n2337), .Z(n41) );
  NAND U2042 ( .A(n42), .B(n41), .Z(n2359) );
  NAND U2043 ( .A(n2360), .B(n2359), .Z(n43) );
  NAND U2044 ( .A(n44), .B(n43), .Z(n2381) );
  NAND U2045 ( .A(n2382), .B(n2381), .Z(n45) );
  NAND U2046 ( .A(n46), .B(n45), .Z(n2403) );
  NAND U2047 ( .A(n2404), .B(n2403), .Z(n47) );
  NAND U2048 ( .A(n48), .B(n47), .Z(n2425) );
  NAND U2049 ( .A(n2426), .B(n2425), .Z(n49) );
  NAND U2050 ( .A(n50), .B(n49), .Z(n2447) );
  NAND U2051 ( .A(n2448), .B(n2447), .Z(n51) );
  NAND U2052 ( .A(n52), .B(n51), .Z(n2469) );
  NAND U2053 ( .A(n2470), .B(n2469), .Z(n53) );
  NAND U2054 ( .A(n54), .B(n53), .Z(n2491) );
  NAND U2055 ( .A(n2492), .B(n2491), .Z(n55) );
  NAND U2056 ( .A(n56), .B(n55), .Z(n2513) );
  NAND U2057 ( .A(n2514), .B(n2513), .Z(n57) );
  NAND U2058 ( .A(n58), .B(n57), .Z(n2535) );
  NAND U2059 ( .A(n2536), .B(n2535), .Z(n59) );
  NAND U2060 ( .A(n60), .B(n59), .Z(n2559) );
  NAND U2061 ( .A(n2560), .B(n2559), .Z(n61) );
  NAND U2062 ( .A(n62), .B(n61), .Z(n2581) );
  NAND U2063 ( .A(n2582), .B(n2581), .Z(n63) );
  NAND U2064 ( .A(n64), .B(n63), .Z(n2603) );
  NAND U2065 ( .A(n2604), .B(n2603), .Z(n65) );
  NAND U2066 ( .A(n66), .B(n65), .Z(n2625) );
  NAND U2067 ( .A(n2626), .B(n2625), .Z(n67) );
  NAND U2068 ( .A(n68), .B(n67), .Z(n2647) );
  NAND U2069 ( .A(n2648), .B(n2647), .Z(n69) );
  NAND U2070 ( .A(n70), .B(n69), .Z(n2669) );
  NAND U2071 ( .A(n2670), .B(n2669), .Z(n71) );
  NAND U2072 ( .A(n72), .B(n71), .Z(n2691) );
  NAND U2073 ( .A(n2692), .B(n2691), .Z(n73) );
  NAND U2074 ( .A(n74), .B(n73), .Z(n2713) );
  NAND U2075 ( .A(n2714), .B(n2713), .Z(n75) );
  NAND U2076 ( .A(n76), .B(n75), .Z(n2735) );
  NAND U2077 ( .A(n2736), .B(n2735), .Z(n77) );
  NAND U2078 ( .A(n78), .B(n77), .Z(n2757) );
  NAND U2079 ( .A(n2758), .B(n2757), .Z(n79) );
  NAND U2080 ( .A(n80), .B(n79), .Z(n2781) );
  NAND U2081 ( .A(n2782), .B(n2781), .Z(n81) );
  NAND U2082 ( .A(n82), .B(n81), .Z(n2803) );
  NAND U2083 ( .A(n2804), .B(n2803), .Z(n83) );
  NAND U2084 ( .A(n84), .B(n83), .Z(n2825) );
  NAND U2085 ( .A(n2826), .B(n2825), .Z(n85) );
  NAND U2086 ( .A(n86), .B(n85), .Z(n2847) );
  NAND U2087 ( .A(n2848), .B(n2847), .Z(n87) );
  NAND U2088 ( .A(n88), .B(n87), .Z(n2869) );
  NAND U2089 ( .A(n2870), .B(n2869), .Z(n89) );
  NAND U2090 ( .A(n90), .B(n89), .Z(n2891) );
  NAND U2091 ( .A(n2892), .B(n2891), .Z(n91) );
  NAND U2092 ( .A(n92), .B(n91), .Z(n2913) );
  NAND U2093 ( .A(n2914), .B(n2913), .Z(n93) );
  NAND U2094 ( .A(n94), .B(n93), .Z(n2935) );
  NAND U2095 ( .A(n2936), .B(n2935), .Z(n95) );
  NAND U2096 ( .A(n96), .B(n95), .Z(n2957) );
  NAND U2097 ( .A(n2958), .B(n2957), .Z(n97) );
  NAND U2098 ( .A(n98), .B(n97), .Z(n2979) );
  NAND U2099 ( .A(n2980), .B(n2979), .Z(n99) );
  NAND U2100 ( .A(n100), .B(n99), .Z(n3003) );
  NAND U2101 ( .A(n3004), .B(n3003), .Z(n101) );
  NAND U2102 ( .A(n102), .B(n101), .Z(n3025) );
  NAND U2103 ( .A(n3026), .B(n3025), .Z(n103) );
  NAND U2104 ( .A(n104), .B(n103), .Z(n3047) );
  NAND U2105 ( .A(n3048), .B(n3047), .Z(n105) );
  NAND U2106 ( .A(n106), .B(n105), .Z(n3069) );
  NAND U2107 ( .A(n3070), .B(n3069), .Z(n107) );
  NAND U2108 ( .A(n108), .B(n107), .Z(n3091) );
  NAND U2109 ( .A(n3092), .B(n3091), .Z(n109) );
  NAND U2110 ( .A(n110), .B(n109), .Z(n3113) );
  NAND U2111 ( .A(n3114), .B(n3113), .Z(n111) );
  NAND U2112 ( .A(n112), .B(n111), .Z(n3135) );
  NAND U2113 ( .A(n3136), .B(n3135), .Z(n113) );
  NAND U2114 ( .A(n114), .B(n113), .Z(n3157) );
  NAND U2115 ( .A(n3158), .B(n3157), .Z(n115) );
  NAND U2116 ( .A(n116), .B(n115), .Z(n3179) );
  NAND U2117 ( .A(n3180), .B(n3179), .Z(n117) );
  NAND U2118 ( .A(n118), .B(n117), .Z(n3201) );
  NAND U2119 ( .A(n3202), .B(n3201), .Z(n119) );
  NAND U2120 ( .A(n120), .B(n119), .Z(n3225) );
  NAND U2121 ( .A(n3226), .B(n3225), .Z(n121) );
  NAND U2122 ( .A(n122), .B(n121), .Z(n3247) );
  NAND U2123 ( .A(n3248), .B(n3247), .Z(n123) );
  NAND U2124 ( .A(n124), .B(n123), .Z(n3269) );
  NAND U2125 ( .A(n3270), .B(n3269), .Z(n125) );
  NAND U2126 ( .A(n126), .B(n125), .Z(n3291) );
  NAND U2127 ( .A(n3292), .B(n3291), .Z(n127) );
  NAND U2128 ( .A(n128), .B(n127), .Z(n3313) );
  NAND U2129 ( .A(n3314), .B(n3313), .Z(n129) );
  NAND U2130 ( .A(n130), .B(n129), .Z(n3335) );
  NAND U2131 ( .A(n3336), .B(n3335), .Z(n131) );
  NAND U2132 ( .A(n132), .B(n131), .Z(n3357) );
  NAND U2133 ( .A(n3358), .B(n3357), .Z(n133) );
  NAND U2134 ( .A(n134), .B(n133), .Z(n3379) );
  NAND U2135 ( .A(n3380), .B(n3379), .Z(n135) );
  NAND U2136 ( .A(n136), .B(n135), .Z(n3401) );
  NAND U2137 ( .A(n3402), .B(n3401), .Z(n137) );
  NAND U2138 ( .A(n138), .B(n137), .Z(n3423) );
  NAND U2139 ( .A(n3424), .B(n3423), .Z(n139) );
  NAND U2140 ( .A(n140), .B(n139), .Z(n3447) );
  NAND U2141 ( .A(n3448), .B(n3447), .Z(n141) );
  NAND U2142 ( .A(n142), .B(n141), .Z(n3469) );
  NAND U2143 ( .A(n3470), .B(n3469), .Z(n143) );
  NAND U2144 ( .A(n144), .B(n143), .Z(n3491) );
  NAND U2145 ( .A(n3492), .B(n3491), .Z(n145) );
  NAND U2146 ( .A(n146), .B(n145), .Z(n3513) );
  NAND U2147 ( .A(n3514), .B(n3513), .Z(n147) );
  NAND U2148 ( .A(n148), .B(n147), .Z(n3535) );
  NAND U2149 ( .A(n3536), .B(n3535), .Z(n149) );
  NAND U2150 ( .A(n150), .B(n149), .Z(n3557) );
  NAND U2151 ( .A(n3558), .B(n3557), .Z(n151) );
  NAND U2152 ( .A(n152), .B(n151), .Z(n3579) );
  NAND U2153 ( .A(n3580), .B(n3579), .Z(n153) );
  NAND U2154 ( .A(n154), .B(n153), .Z(n3601) );
  NAND U2155 ( .A(n3602), .B(n3601), .Z(n155) );
  NAND U2156 ( .A(n156), .B(n155), .Z(n3623) );
  NAND U2157 ( .A(n3624), .B(n3623), .Z(n157) );
  NAND U2158 ( .A(n158), .B(n157), .Z(n3645) );
  NAND U2159 ( .A(n3646), .B(n3645), .Z(n159) );
  NAND U2160 ( .A(n160), .B(n159), .Z(n3669) );
  NAND U2161 ( .A(n3670), .B(n3669), .Z(n161) );
  NAND U2162 ( .A(n162), .B(n161), .Z(n3691) );
  NAND U2163 ( .A(n3692), .B(n3691), .Z(n163) );
  NAND U2164 ( .A(n164), .B(n163), .Z(n3713) );
  NAND U2165 ( .A(n3714), .B(n3713), .Z(n165) );
  NAND U2166 ( .A(n166), .B(n165), .Z(n3735) );
  NAND U2167 ( .A(n3736), .B(n3735), .Z(n167) );
  NAND U2168 ( .A(n168), .B(n167), .Z(n3757) );
  NAND U2169 ( .A(n3758), .B(n3757), .Z(n169) );
  NAND U2170 ( .A(n170), .B(n169), .Z(n3779) );
  NAND U2171 ( .A(n3780), .B(n3779), .Z(n171) );
  NAND U2172 ( .A(n172), .B(n171), .Z(n3801) );
  NAND U2173 ( .A(n3802), .B(n3801), .Z(n173) );
  NAND U2174 ( .A(n174), .B(n173), .Z(n3823) );
  NAND U2175 ( .A(n3824), .B(n3823), .Z(n175) );
  NAND U2176 ( .A(n176), .B(n175), .Z(n3845) );
  NAND U2177 ( .A(n3846), .B(n3845), .Z(n177) );
  NAND U2178 ( .A(n178), .B(n177), .Z(n3867) );
  NAND U2179 ( .A(n3868), .B(n3867), .Z(n179) );
  NAND U2180 ( .A(n180), .B(n179), .Z(n3891) );
  NAND U2181 ( .A(n3892), .B(n3891), .Z(n181) );
  NAND U2182 ( .A(n182), .B(n181), .Z(n3913) );
  NAND U2183 ( .A(n3914), .B(n3913), .Z(n183) );
  NAND U2184 ( .A(n184), .B(n183), .Z(n3935) );
  NAND U2185 ( .A(n3936), .B(n3935), .Z(n185) );
  NAND U2186 ( .A(n186), .B(n185), .Z(n3957) );
  NAND U2187 ( .A(n3958), .B(n3957), .Z(n187) );
  NAND U2188 ( .A(n188), .B(n187), .Z(n3979) );
  NAND U2189 ( .A(n3980), .B(n3979), .Z(n189) );
  NAND U2190 ( .A(n190), .B(n189), .Z(n4001) );
  NAND U2191 ( .A(n4002), .B(n4001), .Z(n191) );
  NAND U2192 ( .A(n192), .B(n191), .Z(n4023) );
  NAND U2193 ( .A(n4024), .B(n4023), .Z(n193) );
  NAND U2194 ( .A(n194), .B(n193), .Z(n4045) );
  NAND U2195 ( .A(n4046), .B(n4045), .Z(n195) );
  NAND U2196 ( .A(n196), .B(n195), .Z(n4067) );
  NAND U2197 ( .A(n4068), .B(n4067), .Z(n197) );
  NAND U2198 ( .A(n198), .B(n197), .Z(n4089) );
  NAND U2199 ( .A(n4090), .B(n4089), .Z(n199) );
  NAND U2200 ( .A(n200), .B(n199), .Z(n2037) );
  NAND U2201 ( .A(n2038), .B(n2037), .Z(n201) );
  NAND U2202 ( .A(n202), .B(n201), .Z(n2079) );
  NAND U2203 ( .A(n2080), .B(n2079), .Z(n203) );
  NAND U2204 ( .A(n204), .B(n203), .Z(n2099) );
  NAND U2205 ( .A(n2100), .B(n2099), .Z(n205) );
  NAND U2206 ( .A(n206), .B(n205), .Z(n2101) );
  NAND U2207 ( .A(n2102), .B(n2101), .Z(n207) );
  NAND U2208 ( .A(n208), .B(n207), .Z(n2103) );
  NAND U2209 ( .A(n2104), .B(n2103), .Z(n209) );
  NAND U2210 ( .A(n210), .B(n209), .Z(n2105) );
  NAND U2211 ( .A(n2106), .B(n2105), .Z(n211) );
  NAND U2212 ( .A(n212), .B(n211), .Z(n2107) );
  NAND U2213 ( .A(n2108), .B(n2107), .Z(n213) );
  NAND U2214 ( .A(n214), .B(n213), .Z(n2109) );
  NAND U2215 ( .A(n2110), .B(n2109), .Z(n215) );
  NAND U2216 ( .A(n216), .B(n215), .Z(n2111) );
  NAND U2217 ( .A(n2112), .B(n2111), .Z(n217) );
  NAND U2218 ( .A(n218), .B(n217), .Z(n2113) );
  NAND U2219 ( .A(n2114), .B(n2113), .Z(n219) );
  NAND U2220 ( .A(n220), .B(n219), .Z(n2117) );
  NAND U2221 ( .A(n2118), .B(n2117), .Z(n221) );
  NAND U2222 ( .A(n222), .B(n221), .Z(n2119) );
  NAND U2223 ( .A(n2120), .B(n2119), .Z(n223) );
  NAND U2224 ( .A(n224), .B(n223), .Z(n2121) );
  NAND U2225 ( .A(n2122), .B(n2121), .Z(n225) );
  NAND U2226 ( .A(n226), .B(n225), .Z(n2123) );
  NAND U2227 ( .A(n2124), .B(n2123), .Z(n227) );
  NAND U2228 ( .A(n228), .B(n227), .Z(n2125) );
  NAND U2229 ( .A(n2126), .B(n2125), .Z(n229) );
  NAND U2230 ( .A(n230), .B(n229), .Z(n2127) );
  NAND U2231 ( .A(n2128), .B(n2127), .Z(n231) );
  NAND U2232 ( .A(n232), .B(n231), .Z(n2129) );
  NAND U2233 ( .A(n2130), .B(n2129), .Z(n233) );
  NAND U2234 ( .A(n234), .B(n233), .Z(n2131) );
  NAND U2235 ( .A(n2132), .B(n2131), .Z(n235) );
  NAND U2236 ( .A(n236), .B(n235), .Z(n2133) );
  NAND U2237 ( .A(n2134), .B(n2133), .Z(n237) );
  NAND U2238 ( .A(n238), .B(n237), .Z(n2135) );
  NAND U2239 ( .A(n2136), .B(n2135), .Z(n239) );
  NAND U2240 ( .A(n240), .B(n239), .Z(n2139) );
  NAND U2241 ( .A(n2140), .B(n2139), .Z(n241) );
  NAND U2242 ( .A(n242), .B(n241), .Z(n2141) );
  NAND U2243 ( .A(n2142), .B(n2141), .Z(n243) );
  NAND U2244 ( .A(n244), .B(n243), .Z(n2143) );
  NAND U2245 ( .A(n2144), .B(n2143), .Z(n245) );
  NAND U2246 ( .A(n246), .B(n245), .Z(n2145) );
  NAND U2247 ( .A(n2146), .B(n2145), .Z(n247) );
  NAND U2248 ( .A(n248), .B(n247), .Z(n2147) );
  NAND U2249 ( .A(n2148), .B(n2147), .Z(n249) );
  NAND U2250 ( .A(n250), .B(n249), .Z(n2149) );
  NAND U2251 ( .A(n2150), .B(n2149), .Z(n251) );
  NAND U2252 ( .A(n252), .B(n251), .Z(n2151) );
  NAND U2253 ( .A(n2152), .B(n2151), .Z(n253) );
  NAND U2254 ( .A(n254), .B(n253), .Z(n2153) );
  NAND U2255 ( .A(n2154), .B(n2153), .Z(n255) );
  NAND U2256 ( .A(n256), .B(n255), .Z(n2155) );
  NAND U2257 ( .A(n2156), .B(n2155), .Z(n257) );
  NAND U2258 ( .A(n258), .B(n257), .Z(n2157) );
  NAND U2259 ( .A(n2158), .B(n2157), .Z(n259) );
  NAND U2260 ( .A(n260), .B(n259), .Z(n2161) );
  NAND U2261 ( .A(n2162), .B(n2161), .Z(n261) );
  NAND U2262 ( .A(n262), .B(n261), .Z(n2163) );
  NAND U2263 ( .A(n2164), .B(n2163), .Z(n263) );
  NAND U2264 ( .A(n264), .B(n263), .Z(n2165) );
  NAND U2265 ( .A(n2166), .B(n2165), .Z(n265) );
  NAND U2266 ( .A(n266), .B(n265), .Z(n2167) );
  NAND U2267 ( .A(n2168), .B(n2167), .Z(n267) );
  NAND U2268 ( .A(n268), .B(n267), .Z(n2169) );
  NAND U2269 ( .A(n2170), .B(n2169), .Z(n269) );
  NAND U2270 ( .A(n270), .B(n269), .Z(n2171) );
  NAND U2271 ( .A(n2172), .B(n2171), .Z(n271) );
  NAND U2272 ( .A(n272), .B(n271), .Z(n2173) );
  NAND U2273 ( .A(n2174), .B(n2173), .Z(n273) );
  NAND U2274 ( .A(n274), .B(n273), .Z(n2175) );
  NAND U2275 ( .A(n2176), .B(n2175), .Z(n275) );
  NAND U2276 ( .A(n276), .B(n275), .Z(n2177) );
  NAND U2277 ( .A(n2178), .B(n2177), .Z(n277) );
  NAND U2278 ( .A(n278), .B(n277), .Z(n2179) );
  NAND U2279 ( .A(n2180), .B(n2179), .Z(n279) );
  NAND U2280 ( .A(n280), .B(n279), .Z(n2183) );
  NAND U2281 ( .A(n2184), .B(n2183), .Z(n281) );
  NAND U2282 ( .A(n282), .B(n281), .Z(n2185) );
  NAND U2283 ( .A(n2186), .B(n2185), .Z(n283) );
  NAND U2284 ( .A(n284), .B(n283), .Z(n2187) );
  NAND U2285 ( .A(n2188), .B(n2187), .Z(n285) );
  NAND U2286 ( .A(n286), .B(n285), .Z(n2189) );
  NAND U2287 ( .A(n2190), .B(n2189), .Z(n287) );
  NAND U2288 ( .A(n288), .B(n287), .Z(n2191) );
  NAND U2289 ( .A(n2192), .B(n2191), .Z(n289) );
  NAND U2290 ( .A(n290), .B(n289), .Z(n2193) );
  NAND U2291 ( .A(n2194), .B(n2193), .Z(n291) );
  NAND U2292 ( .A(n292), .B(n291), .Z(n2195) );
  NAND U2293 ( .A(n2196), .B(n2195), .Z(n293) );
  NAND U2294 ( .A(n294), .B(n293), .Z(n2197) );
  NAND U2295 ( .A(n2198), .B(n2197), .Z(n295) );
  NAND U2296 ( .A(n296), .B(n295), .Z(n2199) );
  NAND U2297 ( .A(n2200), .B(n2199), .Z(n297) );
  NAND U2298 ( .A(n298), .B(n297), .Z(n2201) );
  NAND U2299 ( .A(n2202), .B(n2201), .Z(n299) );
  NAND U2300 ( .A(n300), .B(n299), .Z(n2205) );
  NAND U2301 ( .A(n2206), .B(n2205), .Z(n301) );
  NAND U2302 ( .A(n302), .B(n301), .Z(n2207) );
  NAND U2303 ( .A(n2208), .B(n2207), .Z(n303) );
  NAND U2304 ( .A(n304), .B(n303), .Z(n2209) );
  NAND U2305 ( .A(n2210), .B(n2209), .Z(n305) );
  NAND U2306 ( .A(n306), .B(n305), .Z(n2211) );
  NAND U2307 ( .A(n2212), .B(n2211), .Z(n307) );
  NAND U2308 ( .A(n308), .B(n307), .Z(n2213) );
  NAND U2309 ( .A(n2214), .B(n2213), .Z(n309) );
  NAND U2310 ( .A(n310), .B(n309), .Z(n2215) );
  NAND U2311 ( .A(n2216), .B(n2215), .Z(n311) );
  NAND U2312 ( .A(n312), .B(n311), .Z(n2217) );
  NAND U2313 ( .A(n2218), .B(n2217), .Z(n313) );
  NAND U2314 ( .A(n314), .B(n313), .Z(n2219) );
  NAND U2315 ( .A(n2220), .B(n2219), .Z(n315) );
  NAND U2316 ( .A(n316), .B(n315), .Z(n2221) );
  NAND U2317 ( .A(n2222), .B(n2221), .Z(n317) );
  NAND U2318 ( .A(n318), .B(n317), .Z(n2223) );
  NAND U2319 ( .A(n2224), .B(n2223), .Z(n319) );
  NAND U2320 ( .A(n320), .B(n319), .Z(n2227) );
  NAND U2321 ( .A(n2228), .B(n2227), .Z(n321) );
  NAND U2322 ( .A(n322), .B(n321), .Z(n2229) );
  NAND U2323 ( .A(n2230), .B(n2229), .Z(n323) );
  NAND U2324 ( .A(n324), .B(n323), .Z(n2231) );
  NAND U2325 ( .A(n2232), .B(n2231), .Z(n325) );
  NAND U2326 ( .A(n326), .B(n325), .Z(n2233) );
  NAND U2327 ( .A(n2234), .B(n2233), .Z(n327) );
  NAND U2328 ( .A(n328), .B(n327), .Z(n2235) );
  NAND U2329 ( .A(n2236), .B(n2235), .Z(n329) );
  NAND U2330 ( .A(n330), .B(n329), .Z(n2237) );
  NAND U2331 ( .A(n2238), .B(n2237), .Z(n331) );
  NAND U2332 ( .A(n332), .B(n331), .Z(n2239) );
  NAND U2333 ( .A(n2240), .B(n2239), .Z(n333) );
  NAND U2334 ( .A(n334), .B(n333), .Z(n2241) );
  NAND U2335 ( .A(n2242), .B(n2241), .Z(n335) );
  NAND U2336 ( .A(n336), .B(n335), .Z(n2243) );
  NAND U2337 ( .A(n2244), .B(n2243), .Z(n337) );
  NAND U2338 ( .A(n338), .B(n337), .Z(n2245) );
  NAND U2339 ( .A(n2246), .B(n2245), .Z(n339) );
  NAND U2340 ( .A(n340), .B(n339), .Z(n2249) );
  NAND U2341 ( .A(n2250), .B(n2249), .Z(n341) );
  NAND U2342 ( .A(n342), .B(n341), .Z(n2251) );
  NAND U2343 ( .A(n2252), .B(n2251), .Z(n343) );
  NAND U2344 ( .A(n344), .B(n343), .Z(n2253) );
  NAND U2345 ( .A(n2254), .B(n2253), .Z(n345) );
  NAND U2346 ( .A(n346), .B(n345), .Z(n2255) );
  NAND U2347 ( .A(n2256), .B(n2255), .Z(n347) );
  NAND U2348 ( .A(n348), .B(n347), .Z(n2257) );
  NAND U2349 ( .A(n2258), .B(n2257), .Z(n349) );
  NAND U2350 ( .A(n350), .B(n349), .Z(n2259) );
  NAND U2351 ( .A(n2260), .B(n2259), .Z(n351) );
  NAND U2352 ( .A(n352), .B(n351), .Z(n2261) );
  NAND U2353 ( .A(n2262), .B(n2261), .Z(n353) );
  NAND U2354 ( .A(n354), .B(n353), .Z(n2263) );
  NAND U2355 ( .A(n2264), .B(n2263), .Z(n355) );
  NAND U2356 ( .A(n356), .B(n355), .Z(n2265) );
  NAND U2357 ( .A(n2266), .B(n2265), .Z(n357) );
  NAND U2358 ( .A(n358), .B(n357), .Z(n2267) );
  NAND U2359 ( .A(n2268), .B(n2267), .Z(n359) );
  NAND U2360 ( .A(n360), .B(n359), .Z(n2271) );
  NAND U2361 ( .A(n2272), .B(n2271), .Z(n361) );
  NAND U2362 ( .A(n362), .B(n361), .Z(n2273) );
  NAND U2363 ( .A(n2274), .B(n2273), .Z(n363) );
  NAND U2364 ( .A(n364), .B(n363), .Z(n2275) );
  NAND U2365 ( .A(n2276), .B(n2275), .Z(n365) );
  NAND U2366 ( .A(n366), .B(n365), .Z(n2277) );
  NAND U2367 ( .A(n2278), .B(n2277), .Z(n367) );
  NAND U2368 ( .A(n368), .B(n367), .Z(n2279) );
  NAND U2369 ( .A(n2280), .B(n2279), .Z(n369) );
  NAND U2370 ( .A(n370), .B(n369), .Z(n2281) );
  NAND U2371 ( .A(n2282), .B(n2281), .Z(n371) );
  NAND U2372 ( .A(n372), .B(n371), .Z(n2283) );
  NAND U2373 ( .A(n2284), .B(n2283), .Z(n373) );
  NAND U2374 ( .A(n374), .B(n373), .Z(n2285) );
  NAND U2375 ( .A(n2286), .B(n2285), .Z(n375) );
  NAND U2376 ( .A(n376), .B(n375), .Z(n2287) );
  NAND U2377 ( .A(n2288), .B(n2287), .Z(n377) );
  NAND U2378 ( .A(n378), .B(n377), .Z(n2289) );
  NAND U2379 ( .A(n2290), .B(n2289), .Z(n379) );
  NAND U2380 ( .A(n380), .B(n379), .Z(n2293) );
  NAND U2381 ( .A(n2294), .B(n2293), .Z(n381) );
  NAND U2382 ( .A(n382), .B(n381), .Z(n2295) );
  NAND U2383 ( .A(n2296), .B(n2295), .Z(n383) );
  NAND U2384 ( .A(n384), .B(n383), .Z(n2297) );
  NAND U2385 ( .A(n2298), .B(n2297), .Z(n385) );
  NAND U2386 ( .A(n386), .B(n385), .Z(n2299) );
  NAND U2387 ( .A(n2300), .B(n2299), .Z(n387) );
  NAND U2388 ( .A(n388), .B(n387), .Z(n2301) );
  NAND U2389 ( .A(n2302), .B(n2301), .Z(n389) );
  NAND U2390 ( .A(n390), .B(n389), .Z(n2303) );
  NAND U2391 ( .A(n2304), .B(n2303), .Z(n391) );
  NAND U2392 ( .A(n392), .B(n391), .Z(n2305) );
  NAND U2393 ( .A(n2306), .B(n2305), .Z(n393) );
  NAND U2394 ( .A(n394), .B(n393), .Z(n2307) );
  NAND U2395 ( .A(n2308), .B(n2307), .Z(n395) );
  NAND U2396 ( .A(n396), .B(n395), .Z(n2309) );
  NAND U2397 ( .A(n2310), .B(n2309), .Z(n397) );
  NAND U2398 ( .A(n398), .B(n397), .Z(n2311) );
  NAND U2399 ( .A(n2312), .B(n2311), .Z(n399) );
  NAND U2400 ( .A(n400), .B(n399), .Z(n2317) );
  NAND U2401 ( .A(n2318), .B(n2317), .Z(n401) );
  NAND U2402 ( .A(n402), .B(n401), .Z(n2319) );
  NAND U2403 ( .A(n2320), .B(n2319), .Z(n403) );
  NAND U2404 ( .A(n404), .B(n403), .Z(n2321) );
  NAND U2405 ( .A(n2322), .B(n2321), .Z(n405) );
  NAND U2406 ( .A(n406), .B(n405), .Z(n2323) );
  NAND U2407 ( .A(n2324), .B(n2323), .Z(n407) );
  NAND U2408 ( .A(n408), .B(n407), .Z(n2325) );
  NAND U2409 ( .A(n2326), .B(n2325), .Z(n409) );
  NAND U2410 ( .A(n410), .B(n409), .Z(n2327) );
  NAND U2411 ( .A(n2328), .B(n2327), .Z(n411) );
  NAND U2412 ( .A(n412), .B(n411), .Z(n2329) );
  NAND U2413 ( .A(n2330), .B(n2329), .Z(n413) );
  NAND U2414 ( .A(n414), .B(n413), .Z(n2331) );
  NAND U2415 ( .A(n2332), .B(n2331), .Z(n415) );
  NAND U2416 ( .A(n416), .B(n415), .Z(n2333) );
  NAND U2417 ( .A(n2334), .B(n2333), .Z(n417) );
  NAND U2418 ( .A(n418), .B(n417), .Z(n2335) );
  NAND U2419 ( .A(n2336), .B(n2335), .Z(n419) );
  NAND U2420 ( .A(n420), .B(n419), .Z(n2339) );
  NAND U2421 ( .A(n2340), .B(n2339), .Z(n421) );
  NAND U2422 ( .A(n422), .B(n421), .Z(n2341) );
  NAND U2423 ( .A(n2342), .B(n2341), .Z(n423) );
  NAND U2424 ( .A(n424), .B(n423), .Z(n2343) );
  NAND U2425 ( .A(n2344), .B(n2343), .Z(n425) );
  NAND U2426 ( .A(n426), .B(n425), .Z(n2345) );
  NAND U2427 ( .A(n2346), .B(n2345), .Z(n427) );
  NAND U2428 ( .A(n428), .B(n427), .Z(n2347) );
  NAND U2429 ( .A(n2348), .B(n2347), .Z(n429) );
  NAND U2430 ( .A(n430), .B(n429), .Z(n2349) );
  NAND U2431 ( .A(n2350), .B(n2349), .Z(n431) );
  NAND U2432 ( .A(n432), .B(n431), .Z(n2351) );
  NAND U2433 ( .A(n2352), .B(n2351), .Z(n433) );
  NAND U2434 ( .A(n434), .B(n433), .Z(n2353) );
  NAND U2435 ( .A(n2354), .B(n2353), .Z(n435) );
  NAND U2436 ( .A(n436), .B(n435), .Z(n2355) );
  NAND U2437 ( .A(n2356), .B(n2355), .Z(n437) );
  NAND U2438 ( .A(n438), .B(n437), .Z(n2357) );
  NAND U2439 ( .A(n2358), .B(n2357), .Z(n439) );
  NAND U2440 ( .A(n440), .B(n439), .Z(n2361) );
  NAND U2441 ( .A(n2362), .B(n2361), .Z(n441) );
  NAND U2442 ( .A(n442), .B(n441), .Z(n2363) );
  NAND U2443 ( .A(n2364), .B(n2363), .Z(n443) );
  NAND U2444 ( .A(n444), .B(n443), .Z(n2365) );
  NAND U2445 ( .A(n2366), .B(n2365), .Z(n445) );
  NAND U2446 ( .A(n446), .B(n445), .Z(n2367) );
  NAND U2447 ( .A(n2368), .B(n2367), .Z(n447) );
  NAND U2448 ( .A(n448), .B(n447), .Z(n2369) );
  NAND U2449 ( .A(n2370), .B(n2369), .Z(n449) );
  NAND U2450 ( .A(n450), .B(n449), .Z(n2371) );
  NAND U2451 ( .A(n2372), .B(n2371), .Z(n451) );
  NAND U2452 ( .A(n452), .B(n451), .Z(n2373) );
  NAND U2453 ( .A(n2374), .B(n2373), .Z(n453) );
  NAND U2454 ( .A(n454), .B(n453), .Z(n2375) );
  NAND U2455 ( .A(n2376), .B(n2375), .Z(n455) );
  NAND U2456 ( .A(n456), .B(n455), .Z(n2377) );
  NAND U2457 ( .A(n2378), .B(n2377), .Z(n457) );
  NAND U2458 ( .A(n458), .B(n457), .Z(n2379) );
  NAND U2459 ( .A(n2380), .B(n2379), .Z(n459) );
  NAND U2460 ( .A(n460), .B(n459), .Z(n2383) );
  NAND U2461 ( .A(n2384), .B(n2383), .Z(n461) );
  NAND U2462 ( .A(n462), .B(n461), .Z(n2385) );
  NAND U2463 ( .A(n2386), .B(n2385), .Z(n463) );
  NAND U2464 ( .A(n464), .B(n463), .Z(n2387) );
  NAND U2465 ( .A(n2388), .B(n2387), .Z(n465) );
  NAND U2466 ( .A(n466), .B(n465), .Z(n2389) );
  NAND U2467 ( .A(n2390), .B(n2389), .Z(n467) );
  NAND U2468 ( .A(n468), .B(n467), .Z(n2391) );
  NAND U2469 ( .A(n2392), .B(n2391), .Z(n469) );
  NAND U2470 ( .A(n470), .B(n469), .Z(n2393) );
  NAND U2471 ( .A(n2394), .B(n2393), .Z(n471) );
  NAND U2472 ( .A(n472), .B(n471), .Z(n2395) );
  NAND U2473 ( .A(n2396), .B(n2395), .Z(n473) );
  NAND U2474 ( .A(n474), .B(n473), .Z(n2397) );
  NAND U2475 ( .A(n2398), .B(n2397), .Z(n475) );
  NAND U2476 ( .A(n476), .B(n475), .Z(n2399) );
  NAND U2477 ( .A(n2400), .B(n2399), .Z(n477) );
  NAND U2478 ( .A(n478), .B(n477), .Z(n2401) );
  NAND U2479 ( .A(n2402), .B(n2401), .Z(n479) );
  NAND U2480 ( .A(n480), .B(n479), .Z(n2405) );
  NAND U2481 ( .A(n2406), .B(n2405), .Z(n481) );
  NAND U2482 ( .A(n482), .B(n481), .Z(n2407) );
  NAND U2483 ( .A(n2408), .B(n2407), .Z(n483) );
  NAND U2484 ( .A(n484), .B(n483), .Z(n2409) );
  NAND U2485 ( .A(n2410), .B(n2409), .Z(n485) );
  NAND U2486 ( .A(n486), .B(n485), .Z(n2411) );
  NAND U2487 ( .A(n2412), .B(n2411), .Z(n487) );
  NAND U2488 ( .A(n488), .B(n487), .Z(n2413) );
  NAND U2489 ( .A(n2414), .B(n2413), .Z(n489) );
  NAND U2490 ( .A(n490), .B(n489), .Z(n2415) );
  NAND U2491 ( .A(n2416), .B(n2415), .Z(n491) );
  NAND U2492 ( .A(n492), .B(n491), .Z(n2417) );
  NAND U2493 ( .A(n2418), .B(n2417), .Z(n493) );
  NAND U2494 ( .A(n494), .B(n493), .Z(n2419) );
  NAND U2495 ( .A(n2420), .B(n2419), .Z(n495) );
  NAND U2496 ( .A(n496), .B(n495), .Z(n2421) );
  NAND U2497 ( .A(n2422), .B(n2421), .Z(n497) );
  NAND U2498 ( .A(n498), .B(n497), .Z(n2423) );
  NAND U2499 ( .A(n2424), .B(n2423), .Z(n499) );
  NAND U2500 ( .A(n500), .B(n499), .Z(n2427) );
  NAND U2501 ( .A(n2428), .B(n2427), .Z(n501) );
  NAND U2502 ( .A(n502), .B(n501), .Z(n2429) );
  NAND U2503 ( .A(n2430), .B(n2429), .Z(n503) );
  NAND U2504 ( .A(n504), .B(n503), .Z(n2431) );
  NAND U2505 ( .A(n2432), .B(n2431), .Z(n505) );
  NAND U2506 ( .A(n506), .B(n505), .Z(n2433) );
  NAND U2507 ( .A(n2434), .B(n2433), .Z(n507) );
  NAND U2508 ( .A(n508), .B(n507), .Z(n2435) );
  NAND U2509 ( .A(n2436), .B(n2435), .Z(n509) );
  NAND U2510 ( .A(n510), .B(n509), .Z(n2437) );
  NAND U2511 ( .A(n2438), .B(n2437), .Z(n511) );
  NAND U2512 ( .A(n512), .B(n511), .Z(n2439) );
  NAND U2513 ( .A(n2440), .B(n2439), .Z(n513) );
  NAND U2514 ( .A(n514), .B(n513), .Z(n2441) );
  NAND U2515 ( .A(n2442), .B(n2441), .Z(n515) );
  NAND U2516 ( .A(n516), .B(n515), .Z(n2443) );
  NAND U2517 ( .A(n2444), .B(n2443), .Z(n517) );
  NAND U2518 ( .A(n518), .B(n517), .Z(n2445) );
  NAND U2519 ( .A(n2446), .B(n2445), .Z(n519) );
  NAND U2520 ( .A(n520), .B(n519), .Z(n2449) );
  NAND U2521 ( .A(n2450), .B(n2449), .Z(n521) );
  NAND U2522 ( .A(n522), .B(n521), .Z(n2451) );
  NAND U2523 ( .A(n2452), .B(n2451), .Z(n523) );
  NAND U2524 ( .A(n524), .B(n523), .Z(n2453) );
  NAND U2525 ( .A(n2454), .B(n2453), .Z(n525) );
  NAND U2526 ( .A(n526), .B(n525), .Z(n2455) );
  NAND U2527 ( .A(n2456), .B(n2455), .Z(n527) );
  NAND U2528 ( .A(n528), .B(n527), .Z(n2457) );
  NAND U2529 ( .A(n2458), .B(n2457), .Z(n529) );
  NAND U2530 ( .A(n530), .B(n529), .Z(n2459) );
  NAND U2531 ( .A(n2460), .B(n2459), .Z(n531) );
  NAND U2532 ( .A(n532), .B(n531), .Z(n2461) );
  NAND U2533 ( .A(n2462), .B(n2461), .Z(n533) );
  NAND U2534 ( .A(n534), .B(n533), .Z(n2463) );
  NAND U2535 ( .A(n2464), .B(n2463), .Z(n535) );
  NAND U2536 ( .A(n536), .B(n535), .Z(n2465) );
  NAND U2537 ( .A(n2466), .B(n2465), .Z(n537) );
  NAND U2538 ( .A(n538), .B(n537), .Z(n2467) );
  NAND U2539 ( .A(n2468), .B(n2467), .Z(n539) );
  NAND U2540 ( .A(n540), .B(n539), .Z(n2471) );
  NAND U2541 ( .A(n2472), .B(n2471), .Z(n541) );
  NAND U2542 ( .A(n542), .B(n541), .Z(n2473) );
  NAND U2543 ( .A(n2474), .B(n2473), .Z(n543) );
  NAND U2544 ( .A(n544), .B(n543), .Z(n2475) );
  NAND U2545 ( .A(n2476), .B(n2475), .Z(n545) );
  NAND U2546 ( .A(n546), .B(n545), .Z(n2477) );
  NAND U2547 ( .A(n2478), .B(n2477), .Z(n547) );
  NAND U2548 ( .A(n548), .B(n547), .Z(n2479) );
  NAND U2549 ( .A(n2480), .B(n2479), .Z(n549) );
  NAND U2550 ( .A(n550), .B(n549), .Z(n2481) );
  NAND U2551 ( .A(n2482), .B(n2481), .Z(n551) );
  NAND U2552 ( .A(n552), .B(n551), .Z(n2483) );
  NAND U2553 ( .A(n2484), .B(n2483), .Z(n553) );
  NAND U2554 ( .A(n554), .B(n553), .Z(n2485) );
  NAND U2555 ( .A(n2486), .B(n2485), .Z(n555) );
  NAND U2556 ( .A(n556), .B(n555), .Z(n2487) );
  NAND U2557 ( .A(n2488), .B(n2487), .Z(n557) );
  NAND U2558 ( .A(n558), .B(n557), .Z(n2489) );
  NAND U2559 ( .A(n2490), .B(n2489), .Z(n559) );
  NAND U2560 ( .A(n560), .B(n559), .Z(n2493) );
  NAND U2561 ( .A(n2494), .B(n2493), .Z(n561) );
  NAND U2562 ( .A(n562), .B(n561), .Z(n2495) );
  NAND U2563 ( .A(n2496), .B(n2495), .Z(n563) );
  NAND U2564 ( .A(n564), .B(n563), .Z(n2497) );
  NAND U2565 ( .A(n2498), .B(n2497), .Z(n565) );
  NAND U2566 ( .A(n566), .B(n565), .Z(n2499) );
  NAND U2567 ( .A(n2500), .B(n2499), .Z(n567) );
  NAND U2568 ( .A(n568), .B(n567), .Z(n2501) );
  NAND U2569 ( .A(n2502), .B(n2501), .Z(n569) );
  NAND U2570 ( .A(n570), .B(n569), .Z(n2503) );
  NAND U2571 ( .A(n2504), .B(n2503), .Z(n571) );
  NAND U2572 ( .A(n572), .B(n571), .Z(n2505) );
  NAND U2573 ( .A(n2506), .B(n2505), .Z(n573) );
  NAND U2574 ( .A(n574), .B(n573), .Z(n2507) );
  NAND U2575 ( .A(n2508), .B(n2507), .Z(n575) );
  NAND U2576 ( .A(n576), .B(n575), .Z(n2509) );
  NAND U2577 ( .A(n2510), .B(n2509), .Z(n577) );
  NAND U2578 ( .A(n578), .B(n577), .Z(n2511) );
  NAND U2579 ( .A(n2512), .B(n2511), .Z(n579) );
  NAND U2580 ( .A(n580), .B(n579), .Z(n2515) );
  NAND U2581 ( .A(n2516), .B(n2515), .Z(n581) );
  NAND U2582 ( .A(n582), .B(n581), .Z(n2517) );
  NAND U2583 ( .A(n2518), .B(n2517), .Z(n583) );
  NAND U2584 ( .A(n584), .B(n583), .Z(n2519) );
  NAND U2585 ( .A(n2520), .B(n2519), .Z(n585) );
  NAND U2586 ( .A(n586), .B(n585), .Z(n2521) );
  NAND U2587 ( .A(n2522), .B(n2521), .Z(n587) );
  NAND U2588 ( .A(n588), .B(n587), .Z(n2523) );
  NAND U2589 ( .A(n2524), .B(n2523), .Z(n589) );
  NAND U2590 ( .A(n590), .B(n589), .Z(n2525) );
  NAND U2591 ( .A(n2526), .B(n2525), .Z(n591) );
  NAND U2592 ( .A(n592), .B(n591), .Z(n2527) );
  NAND U2593 ( .A(n2528), .B(n2527), .Z(n593) );
  NAND U2594 ( .A(n594), .B(n593), .Z(n2529) );
  NAND U2595 ( .A(n2530), .B(n2529), .Z(n595) );
  NAND U2596 ( .A(n596), .B(n595), .Z(n2531) );
  NAND U2597 ( .A(n2532), .B(n2531), .Z(n597) );
  NAND U2598 ( .A(n598), .B(n597), .Z(n2533) );
  NAND U2599 ( .A(n2534), .B(n2533), .Z(n599) );
  NAND U2600 ( .A(n600), .B(n599), .Z(n2539) );
  NAND U2601 ( .A(n2540), .B(n2539), .Z(n601) );
  NAND U2602 ( .A(n602), .B(n601), .Z(n2541) );
  NAND U2603 ( .A(n2542), .B(n2541), .Z(n603) );
  NAND U2604 ( .A(n604), .B(n603), .Z(n2543) );
  NAND U2605 ( .A(n2544), .B(n2543), .Z(n605) );
  NAND U2606 ( .A(n606), .B(n605), .Z(n2545) );
  NAND U2607 ( .A(n2546), .B(n2545), .Z(n607) );
  NAND U2608 ( .A(n608), .B(n607), .Z(n2547) );
  NAND U2609 ( .A(n2548), .B(n2547), .Z(n609) );
  NAND U2610 ( .A(n610), .B(n609), .Z(n2549) );
  NAND U2611 ( .A(n2550), .B(n2549), .Z(n611) );
  NAND U2612 ( .A(n612), .B(n611), .Z(n2551) );
  NAND U2613 ( .A(n2552), .B(n2551), .Z(n613) );
  NAND U2614 ( .A(n614), .B(n613), .Z(n2553) );
  NAND U2615 ( .A(n2554), .B(n2553), .Z(n615) );
  NAND U2616 ( .A(n616), .B(n615), .Z(n2555) );
  NAND U2617 ( .A(n2556), .B(n2555), .Z(n617) );
  NAND U2618 ( .A(n618), .B(n617), .Z(n2557) );
  NAND U2619 ( .A(n2558), .B(n2557), .Z(n619) );
  NAND U2620 ( .A(n620), .B(n619), .Z(n2561) );
  NAND U2621 ( .A(n2562), .B(n2561), .Z(n621) );
  NAND U2622 ( .A(n622), .B(n621), .Z(n2563) );
  NAND U2623 ( .A(n2564), .B(n2563), .Z(n623) );
  NAND U2624 ( .A(n624), .B(n623), .Z(n2565) );
  NAND U2625 ( .A(n2566), .B(n2565), .Z(n625) );
  NAND U2626 ( .A(n626), .B(n625), .Z(n2567) );
  NAND U2627 ( .A(n2568), .B(n2567), .Z(n627) );
  NAND U2628 ( .A(n628), .B(n627), .Z(n2569) );
  NAND U2629 ( .A(n2570), .B(n2569), .Z(n629) );
  NAND U2630 ( .A(n630), .B(n629), .Z(n2571) );
  NAND U2631 ( .A(n2572), .B(n2571), .Z(n631) );
  NAND U2632 ( .A(n632), .B(n631), .Z(n2573) );
  NAND U2633 ( .A(n2574), .B(n2573), .Z(n633) );
  NAND U2634 ( .A(n634), .B(n633), .Z(n2575) );
  NAND U2635 ( .A(n2576), .B(n2575), .Z(n635) );
  NAND U2636 ( .A(n636), .B(n635), .Z(n2577) );
  NAND U2637 ( .A(n2578), .B(n2577), .Z(n637) );
  NAND U2638 ( .A(n638), .B(n637), .Z(n2579) );
  NAND U2639 ( .A(n2580), .B(n2579), .Z(n639) );
  NAND U2640 ( .A(n640), .B(n639), .Z(n2583) );
  NAND U2641 ( .A(n2584), .B(n2583), .Z(n641) );
  NAND U2642 ( .A(n642), .B(n641), .Z(n2585) );
  NAND U2643 ( .A(n2586), .B(n2585), .Z(n643) );
  NAND U2644 ( .A(n644), .B(n643), .Z(n2587) );
  NAND U2645 ( .A(n2588), .B(n2587), .Z(n645) );
  NAND U2646 ( .A(n646), .B(n645), .Z(n2589) );
  NAND U2647 ( .A(n2590), .B(n2589), .Z(n647) );
  NAND U2648 ( .A(n648), .B(n647), .Z(n2591) );
  NAND U2649 ( .A(n2592), .B(n2591), .Z(n649) );
  NAND U2650 ( .A(n650), .B(n649), .Z(n2593) );
  NAND U2651 ( .A(n2594), .B(n2593), .Z(n651) );
  NAND U2652 ( .A(n652), .B(n651), .Z(n2595) );
  NAND U2653 ( .A(n2596), .B(n2595), .Z(n653) );
  NAND U2654 ( .A(n654), .B(n653), .Z(n2597) );
  NAND U2655 ( .A(n2598), .B(n2597), .Z(n655) );
  NAND U2656 ( .A(n656), .B(n655), .Z(n2599) );
  NAND U2657 ( .A(n2600), .B(n2599), .Z(n657) );
  NAND U2658 ( .A(n658), .B(n657), .Z(n2601) );
  NAND U2659 ( .A(n2602), .B(n2601), .Z(n659) );
  NAND U2660 ( .A(n660), .B(n659), .Z(n2605) );
  NAND U2661 ( .A(n2606), .B(n2605), .Z(n661) );
  NAND U2662 ( .A(n662), .B(n661), .Z(n2607) );
  NAND U2663 ( .A(n2608), .B(n2607), .Z(n663) );
  NAND U2664 ( .A(n664), .B(n663), .Z(n2609) );
  NAND U2665 ( .A(n2610), .B(n2609), .Z(n665) );
  NAND U2666 ( .A(n666), .B(n665), .Z(n2611) );
  NAND U2667 ( .A(n2612), .B(n2611), .Z(n667) );
  NAND U2668 ( .A(n668), .B(n667), .Z(n2613) );
  NAND U2669 ( .A(n2614), .B(n2613), .Z(n669) );
  NAND U2670 ( .A(n670), .B(n669), .Z(n2615) );
  NAND U2671 ( .A(n2616), .B(n2615), .Z(n671) );
  NAND U2672 ( .A(n672), .B(n671), .Z(n2617) );
  NAND U2673 ( .A(n2618), .B(n2617), .Z(n673) );
  NAND U2674 ( .A(n674), .B(n673), .Z(n2619) );
  NAND U2675 ( .A(n2620), .B(n2619), .Z(n675) );
  NAND U2676 ( .A(n676), .B(n675), .Z(n2621) );
  NAND U2677 ( .A(n2622), .B(n2621), .Z(n677) );
  NAND U2678 ( .A(n678), .B(n677), .Z(n2623) );
  NAND U2679 ( .A(n2624), .B(n2623), .Z(n679) );
  NAND U2680 ( .A(n680), .B(n679), .Z(n2627) );
  NAND U2681 ( .A(n2628), .B(n2627), .Z(n681) );
  NAND U2682 ( .A(n682), .B(n681), .Z(n2629) );
  NAND U2683 ( .A(n2630), .B(n2629), .Z(n683) );
  NAND U2684 ( .A(n684), .B(n683), .Z(n2631) );
  NAND U2685 ( .A(n2632), .B(n2631), .Z(n685) );
  NAND U2686 ( .A(n686), .B(n685), .Z(n2633) );
  NAND U2687 ( .A(n2634), .B(n2633), .Z(n687) );
  NAND U2688 ( .A(n688), .B(n687), .Z(n2635) );
  NAND U2689 ( .A(n2636), .B(n2635), .Z(n689) );
  NAND U2690 ( .A(n690), .B(n689), .Z(n2637) );
  NAND U2691 ( .A(n2638), .B(n2637), .Z(n691) );
  NAND U2692 ( .A(n692), .B(n691), .Z(n2639) );
  NAND U2693 ( .A(n2640), .B(n2639), .Z(n693) );
  NAND U2694 ( .A(n694), .B(n693), .Z(n2641) );
  NAND U2695 ( .A(n2642), .B(n2641), .Z(n695) );
  NAND U2696 ( .A(n696), .B(n695), .Z(n2643) );
  NAND U2697 ( .A(n2644), .B(n2643), .Z(n697) );
  NAND U2698 ( .A(n698), .B(n697), .Z(n2645) );
  NAND U2699 ( .A(n2646), .B(n2645), .Z(n699) );
  NAND U2700 ( .A(n700), .B(n699), .Z(n2649) );
  NAND U2701 ( .A(n2650), .B(n2649), .Z(n701) );
  NAND U2702 ( .A(n702), .B(n701), .Z(n2651) );
  NAND U2703 ( .A(n2652), .B(n2651), .Z(n703) );
  NAND U2704 ( .A(n704), .B(n703), .Z(n2653) );
  NAND U2705 ( .A(n2654), .B(n2653), .Z(n705) );
  NAND U2706 ( .A(n706), .B(n705), .Z(n2655) );
  NAND U2707 ( .A(n2656), .B(n2655), .Z(n707) );
  NAND U2708 ( .A(n708), .B(n707), .Z(n2657) );
  NAND U2709 ( .A(n2658), .B(n2657), .Z(n709) );
  NAND U2710 ( .A(n710), .B(n709), .Z(n2659) );
  NAND U2711 ( .A(n2660), .B(n2659), .Z(n711) );
  NAND U2712 ( .A(n712), .B(n711), .Z(n2661) );
  NAND U2713 ( .A(n2662), .B(n2661), .Z(n713) );
  NAND U2714 ( .A(n714), .B(n713), .Z(n2663) );
  NAND U2715 ( .A(n2664), .B(n2663), .Z(n715) );
  NAND U2716 ( .A(n716), .B(n715), .Z(n2665) );
  NAND U2717 ( .A(n2666), .B(n2665), .Z(n717) );
  NAND U2718 ( .A(n718), .B(n717), .Z(n2667) );
  NAND U2719 ( .A(n2668), .B(n2667), .Z(n719) );
  NAND U2720 ( .A(n720), .B(n719), .Z(n2671) );
  NAND U2721 ( .A(n2672), .B(n2671), .Z(n721) );
  NAND U2722 ( .A(n722), .B(n721), .Z(n2673) );
  NAND U2723 ( .A(n2674), .B(n2673), .Z(n723) );
  NAND U2724 ( .A(n724), .B(n723), .Z(n2675) );
  NAND U2725 ( .A(n2676), .B(n2675), .Z(n725) );
  NAND U2726 ( .A(n726), .B(n725), .Z(n2677) );
  NAND U2727 ( .A(n2678), .B(n2677), .Z(n727) );
  NAND U2728 ( .A(n728), .B(n727), .Z(n2679) );
  NAND U2729 ( .A(n2680), .B(n2679), .Z(n729) );
  NAND U2730 ( .A(n730), .B(n729), .Z(n2681) );
  NAND U2731 ( .A(n2682), .B(n2681), .Z(n731) );
  NAND U2732 ( .A(n732), .B(n731), .Z(n2683) );
  NAND U2733 ( .A(n2684), .B(n2683), .Z(n733) );
  NAND U2734 ( .A(n734), .B(n733), .Z(n2685) );
  NAND U2735 ( .A(n2686), .B(n2685), .Z(n735) );
  NAND U2736 ( .A(n736), .B(n735), .Z(n2687) );
  NAND U2737 ( .A(n2688), .B(n2687), .Z(n737) );
  NAND U2738 ( .A(n738), .B(n737), .Z(n2689) );
  NAND U2739 ( .A(n2690), .B(n2689), .Z(n739) );
  NAND U2740 ( .A(n740), .B(n739), .Z(n2693) );
  NAND U2741 ( .A(n2694), .B(n2693), .Z(n741) );
  NAND U2742 ( .A(n742), .B(n741), .Z(n2695) );
  NAND U2743 ( .A(n2696), .B(n2695), .Z(n743) );
  NAND U2744 ( .A(n744), .B(n743), .Z(n2697) );
  NAND U2745 ( .A(n2698), .B(n2697), .Z(n745) );
  NAND U2746 ( .A(n746), .B(n745), .Z(n2699) );
  NAND U2747 ( .A(n2700), .B(n2699), .Z(n747) );
  NAND U2748 ( .A(n748), .B(n747), .Z(n2701) );
  NAND U2749 ( .A(n2702), .B(n2701), .Z(n749) );
  NAND U2750 ( .A(n750), .B(n749), .Z(n2703) );
  NAND U2751 ( .A(n2704), .B(n2703), .Z(n751) );
  NAND U2752 ( .A(n752), .B(n751), .Z(n2705) );
  NAND U2753 ( .A(n2706), .B(n2705), .Z(n753) );
  NAND U2754 ( .A(n754), .B(n753), .Z(n2707) );
  NAND U2755 ( .A(n2708), .B(n2707), .Z(n755) );
  NAND U2756 ( .A(n756), .B(n755), .Z(n2709) );
  NAND U2757 ( .A(n2710), .B(n2709), .Z(n757) );
  NAND U2758 ( .A(n758), .B(n757), .Z(n2711) );
  NAND U2759 ( .A(n2712), .B(n2711), .Z(n759) );
  NAND U2760 ( .A(n760), .B(n759), .Z(n2715) );
  NAND U2761 ( .A(n2716), .B(n2715), .Z(n761) );
  NAND U2762 ( .A(n762), .B(n761), .Z(n2717) );
  NAND U2763 ( .A(n2718), .B(n2717), .Z(n763) );
  NAND U2764 ( .A(n764), .B(n763), .Z(n2719) );
  NAND U2765 ( .A(n2720), .B(n2719), .Z(n765) );
  NAND U2766 ( .A(n766), .B(n765), .Z(n2721) );
  NAND U2767 ( .A(n2722), .B(n2721), .Z(n767) );
  NAND U2768 ( .A(n768), .B(n767), .Z(n2723) );
  NAND U2769 ( .A(n2724), .B(n2723), .Z(n769) );
  NAND U2770 ( .A(n770), .B(n769), .Z(n2725) );
  NAND U2771 ( .A(n2726), .B(n2725), .Z(n771) );
  NAND U2772 ( .A(n772), .B(n771), .Z(n2727) );
  NAND U2773 ( .A(n2728), .B(n2727), .Z(n773) );
  NAND U2774 ( .A(n774), .B(n773), .Z(n2729) );
  NAND U2775 ( .A(n2730), .B(n2729), .Z(n775) );
  NAND U2776 ( .A(n776), .B(n775), .Z(n2731) );
  NAND U2777 ( .A(n2732), .B(n2731), .Z(n777) );
  NAND U2778 ( .A(n778), .B(n777), .Z(n2733) );
  NAND U2779 ( .A(n2734), .B(n2733), .Z(n779) );
  NAND U2780 ( .A(n780), .B(n779), .Z(n2737) );
  NAND U2781 ( .A(n2738), .B(n2737), .Z(n781) );
  NAND U2782 ( .A(n782), .B(n781), .Z(n2739) );
  NAND U2783 ( .A(n2740), .B(n2739), .Z(n783) );
  NAND U2784 ( .A(n784), .B(n783), .Z(n2741) );
  NAND U2785 ( .A(n2742), .B(n2741), .Z(n785) );
  NAND U2786 ( .A(n786), .B(n785), .Z(n2743) );
  NAND U2787 ( .A(n2744), .B(n2743), .Z(n787) );
  NAND U2788 ( .A(n788), .B(n787), .Z(n2745) );
  NAND U2789 ( .A(n2746), .B(n2745), .Z(n789) );
  NAND U2790 ( .A(n790), .B(n789), .Z(n2747) );
  NAND U2791 ( .A(n2748), .B(n2747), .Z(n791) );
  NAND U2792 ( .A(n792), .B(n791), .Z(n2749) );
  NAND U2793 ( .A(n2750), .B(n2749), .Z(n793) );
  NAND U2794 ( .A(n794), .B(n793), .Z(n2751) );
  NAND U2795 ( .A(n2752), .B(n2751), .Z(n795) );
  NAND U2796 ( .A(n796), .B(n795), .Z(n2753) );
  NAND U2797 ( .A(n2754), .B(n2753), .Z(n797) );
  NAND U2798 ( .A(n798), .B(n797), .Z(n2755) );
  NAND U2799 ( .A(n2756), .B(n2755), .Z(n799) );
  NAND U2800 ( .A(n800), .B(n799), .Z(n2761) );
  NAND U2801 ( .A(n2762), .B(n2761), .Z(n801) );
  NAND U2802 ( .A(n802), .B(n801), .Z(n2763) );
  NAND U2803 ( .A(n2764), .B(n2763), .Z(n803) );
  NAND U2804 ( .A(n804), .B(n803), .Z(n2765) );
  NAND U2805 ( .A(n2766), .B(n2765), .Z(n805) );
  NAND U2806 ( .A(n806), .B(n805), .Z(n2767) );
  NAND U2807 ( .A(n2768), .B(n2767), .Z(n807) );
  NAND U2808 ( .A(n808), .B(n807), .Z(n2769) );
  NAND U2809 ( .A(n2770), .B(n2769), .Z(n809) );
  NAND U2810 ( .A(n810), .B(n809), .Z(n2771) );
  NAND U2811 ( .A(n2772), .B(n2771), .Z(n811) );
  NAND U2812 ( .A(n812), .B(n811), .Z(n2773) );
  NAND U2813 ( .A(n2774), .B(n2773), .Z(n813) );
  NAND U2814 ( .A(n814), .B(n813), .Z(n2775) );
  NAND U2815 ( .A(n2776), .B(n2775), .Z(n815) );
  NAND U2816 ( .A(n816), .B(n815), .Z(n2777) );
  NAND U2817 ( .A(n2778), .B(n2777), .Z(n817) );
  NAND U2818 ( .A(n818), .B(n817), .Z(n2779) );
  NAND U2819 ( .A(n2780), .B(n2779), .Z(n819) );
  NAND U2820 ( .A(n820), .B(n819), .Z(n2783) );
  NAND U2821 ( .A(n2784), .B(n2783), .Z(n821) );
  NAND U2822 ( .A(n822), .B(n821), .Z(n2785) );
  NAND U2823 ( .A(n2786), .B(n2785), .Z(n823) );
  NAND U2824 ( .A(n824), .B(n823), .Z(n2787) );
  NAND U2825 ( .A(n2788), .B(n2787), .Z(n825) );
  NAND U2826 ( .A(n826), .B(n825), .Z(n2789) );
  NAND U2827 ( .A(n2790), .B(n2789), .Z(n827) );
  NAND U2828 ( .A(n828), .B(n827), .Z(n2791) );
  NAND U2829 ( .A(n2792), .B(n2791), .Z(n829) );
  NAND U2830 ( .A(n830), .B(n829), .Z(n2793) );
  NAND U2831 ( .A(n2794), .B(n2793), .Z(n831) );
  NAND U2832 ( .A(n832), .B(n831), .Z(n2795) );
  NAND U2833 ( .A(n2796), .B(n2795), .Z(n833) );
  NAND U2834 ( .A(n834), .B(n833), .Z(n2797) );
  NAND U2835 ( .A(n2798), .B(n2797), .Z(n835) );
  NAND U2836 ( .A(n836), .B(n835), .Z(n2799) );
  NAND U2837 ( .A(n2800), .B(n2799), .Z(n837) );
  NAND U2838 ( .A(n838), .B(n837), .Z(n2801) );
  NAND U2839 ( .A(n2802), .B(n2801), .Z(n839) );
  NAND U2840 ( .A(n840), .B(n839), .Z(n2805) );
  NAND U2841 ( .A(n2806), .B(n2805), .Z(n841) );
  NAND U2842 ( .A(n842), .B(n841), .Z(n2807) );
  NAND U2843 ( .A(n2808), .B(n2807), .Z(n843) );
  NAND U2844 ( .A(n844), .B(n843), .Z(n2809) );
  NAND U2845 ( .A(n2810), .B(n2809), .Z(n845) );
  NAND U2846 ( .A(n846), .B(n845), .Z(n2811) );
  NAND U2847 ( .A(n2812), .B(n2811), .Z(n847) );
  NAND U2848 ( .A(n848), .B(n847), .Z(n2813) );
  NAND U2849 ( .A(n2814), .B(n2813), .Z(n849) );
  NAND U2850 ( .A(n850), .B(n849), .Z(n2815) );
  NAND U2851 ( .A(n2816), .B(n2815), .Z(n851) );
  NAND U2852 ( .A(n852), .B(n851), .Z(n2817) );
  NAND U2853 ( .A(n2818), .B(n2817), .Z(n853) );
  NAND U2854 ( .A(n854), .B(n853), .Z(n2819) );
  NAND U2855 ( .A(n2820), .B(n2819), .Z(n855) );
  NAND U2856 ( .A(n856), .B(n855), .Z(n2821) );
  NAND U2857 ( .A(n2822), .B(n2821), .Z(n857) );
  NAND U2858 ( .A(n858), .B(n857), .Z(n2823) );
  NAND U2859 ( .A(n2824), .B(n2823), .Z(n859) );
  NAND U2860 ( .A(n860), .B(n859), .Z(n2827) );
  NAND U2861 ( .A(n2828), .B(n2827), .Z(n861) );
  NAND U2862 ( .A(n862), .B(n861), .Z(n2829) );
  NAND U2863 ( .A(n2830), .B(n2829), .Z(n863) );
  NAND U2864 ( .A(n864), .B(n863), .Z(n2831) );
  NAND U2865 ( .A(n2832), .B(n2831), .Z(n865) );
  NAND U2866 ( .A(n866), .B(n865), .Z(n2833) );
  NAND U2867 ( .A(n2834), .B(n2833), .Z(n867) );
  NAND U2868 ( .A(n868), .B(n867), .Z(n2835) );
  NAND U2869 ( .A(n2836), .B(n2835), .Z(n869) );
  NAND U2870 ( .A(n870), .B(n869), .Z(n2837) );
  NAND U2871 ( .A(n2838), .B(n2837), .Z(n871) );
  NAND U2872 ( .A(n872), .B(n871), .Z(n2839) );
  NAND U2873 ( .A(n2840), .B(n2839), .Z(n873) );
  NAND U2874 ( .A(n874), .B(n873), .Z(n2841) );
  NAND U2875 ( .A(n2842), .B(n2841), .Z(n875) );
  NAND U2876 ( .A(n876), .B(n875), .Z(n2843) );
  NAND U2877 ( .A(n2844), .B(n2843), .Z(n877) );
  NAND U2878 ( .A(n878), .B(n877), .Z(n2845) );
  NAND U2879 ( .A(n2846), .B(n2845), .Z(n879) );
  NAND U2880 ( .A(n880), .B(n879), .Z(n2849) );
  NAND U2881 ( .A(n2850), .B(n2849), .Z(n881) );
  NAND U2882 ( .A(n882), .B(n881), .Z(n2851) );
  NAND U2883 ( .A(n2852), .B(n2851), .Z(n883) );
  NAND U2884 ( .A(n884), .B(n883), .Z(n2853) );
  NAND U2885 ( .A(n2854), .B(n2853), .Z(n885) );
  NAND U2886 ( .A(n886), .B(n885), .Z(n2855) );
  NAND U2887 ( .A(n2856), .B(n2855), .Z(n887) );
  NAND U2888 ( .A(n888), .B(n887), .Z(n2857) );
  NAND U2889 ( .A(n2858), .B(n2857), .Z(n889) );
  NAND U2890 ( .A(n890), .B(n889), .Z(n2859) );
  NAND U2891 ( .A(n2860), .B(n2859), .Z(n891) );
  NAND U2892 ( .A(n892), .B(n891), .Z(n2861) );
  NAND U2893 ( .A(n2862), .B(n2861), .Z(n893) );
  NAND U2894 ( .A(n894), .B(n893), .Z(n2863) );
  NAND U2895 ( .A(n2864), .B(n2863), .Z(n895) );
  NAND U2896 ( .A(n896), .B(n895), .Z(n2865) );
  NAND U2897 ( .A(n2866), .B(n2865), .Z(n897) );
  NAND U2898 ( .A(n898), .B(n897), .Z(n2867) );
  NAND U2899 ( .A(n2868), .B(n2867), .Z(n899) );
  NAND U2900 ( .A(n900), .B(n899), .Z(n2871) );
  NAND U2901 ( .A(n2872), .B(n2871), .Z(n901) );
  NAND U2902 ( .A(n902), .B(n901), .Z(n2873) );
  NAND U2903 ( .A(n2874), .B(n2873), .Z(n903) );
  NAND U2904 ( .A(n904), .B(n903), .Z(n2875) );
  NAND U2905 ( .A(n2876), .B(n2875), .Z(n905) );
  NAND U2906 ( .A(n906), .B(n905), .Z(n2877) );
  NAND U2907 ( .A(n2878), .B(n2877), .Z(n907) );
  NAND U2908 ( .A(n908), .B(n907), .Z(n2879) );
  NAND U2909 ( .A(n2880), .B(n2879), .Z(n909) );
  NAND U2910 ( .A(n910), .B(n909), .Z(n2881) );
  NAND U2911 ( .A(n2882), .B(n2881), .Z(n911) );
  NAND U2912 ( .A(n912), .B(n911), .Z(n2883) );
  NAND U2913 ( .A(n2884), .B(n2883), .Z(n913) );
  NAND U2914 ( .A(n914), .B(n913), .Z(n2885) );
  NAND U2915 ( .A(n2886), .B(n2885), .Z(n915) );
  NAND U2916 ( .A(n916), .B(n915), .Z(n2887) );
  NAND U2917 ( .A(n2888), .B(n2887), .Z(n917) );
  NAND U2918 ( .A(n918), .B(n917), .Z(n2889) );
  NAND U2919 ( .A(n2890), .B(n2889), .Z(n919) );
  NAND U2920 ( .A(n920), .B(n919), .Z(n2893) );
  NAND U2921 ( .A(n2894), .B(n2893), .Z(n921) );
  NAND U2922 ( .A(n922), .B(n921), .Z(n2895) );
  NAND U2923 ( .A(n2896), .B(n2895), .Z(n923) );
  NAND U2924 ( .A(n924), .B(n923), .Z(n2897) );
  NAND U2925 ( .A(n2898), .B(n2897), .Z(n925) );
  NAND U2926 ( .A(n926), .B(n925), .Z(n2899) );
  NAND U2927 ( .A(n2900), .B(n2899), .Z(n927) );
  NAND U2928 ( .A(n928), .B(n927), .Z(n2901) );
  NAND U2929 ( .A(n2902), .B(n2901), .Z(n929) );
  NAND U2930 ( .A(n930), .B(n929), .Z(n2903) );
  NAND U2931 ( .A(n2904), .B(n2903), .Z(n931) );
  NAND U2932 ( .A(n932), .B(n931), .Z(n2905) );
  NAND U2933 ( .A(n2906), .B(n2905), .Z(n933) );
  NAND U2934 ( .A(n934), .B(n933), .Z(n2907) );
  NAND U2935 ( .A(n2908), .B(n2907), .Z(n935) );
  NAND U2936 ( .A(n936), .B(n935), .Z(n2909) );
  NAND U2937 ( .A(n2910), .B(n2909), .Z(n937) );
  NAND U2938 ( .A(n938), .B(n937), .Z(n2911) );
  NAND U2939 ( .A(n2912), .B(n2911), .Z(n939) );
  NAND U2940 ( .A(n940), .B(n939), .Z(n2915) );
  NAND U2941 ( .A(n2916), .B(n2915), .Z(n941) );
  NAND U2942 ( .A(n942), .B(n941), .Z(n2917) );
  NAND U2943 ( .A(n2918), .B(n2917), .Z(n943) );
  NAND U2944 ( .A(n944), .B(n943), .Z(n2919) );
  NAND U2945 ( .A(n2920), .B(n2919), .Z(n945) );
  NAND U2946 ( .A(n946), .B(n945), .Z(n2921) );
  NAND U2947 ( .A(n2922), .B(n2921), .Z(n947) );
  NAND U2948 ( .A(n948), .B(n947), .Z(n2923) );
  NAND U2949 ( .A(n2924), .B(n2923), .Z(n949) );
  NAND U2950 ( .A(n950), .B(n949), .Z(n2925) );
  NAND U2951 ( .A(n2926), .B(n2925), .Z(n951) );
  NAND U2952 ( .A(n952), .B(n951), .Z(n2927) );
  NAND U2953 ( .A(n2928), .B(n2927), .Z(n953) );
  NAND U2954 ( .A(n954), .B(n953), .Z(n2929) );
  NAND U2955 ( .A(n2930), .B(n2929), .Z(n955) );
  NAND U2956 ( .A(n956), .B(n955), .Z(n2931) );
  NAND U2957 ( .A(n2932), .B(n2931), .Z(n957) );
  NAND U2958 ( .A(n958), .B(n957), .Z(n2933) );
  NAND U2959 ( .A(n2934), .B(n2933), .Z(n959) );
  NAND U2960 ( .A(n960), .B(n959), .Z(n2937) );
  NAND U2961 ( .A(n2938), .B(n2937), .Z(n961) );
  NAND U2962 ( .A(n962), .B(n961), .Z(n2939) );
  NAND U2963 ( .A(n2940), .B(n2939), .Z(n963) );
  NAND U2964 ( .A(n964), .B(n963), .Z(n2941) );
  NAND U2965 ( .A(n2942), .B(n2941), .Z(n965) );
  NAND U2966 ( .A(n966), .B(n965), .Z(n2943) );
  NAND U2967 ( .A(n2944), .B(n2943), .Z(n967) );
  NAND U2968 ( .A(n968), .B(n967), .Z(n2945) );
  NAND U2969 ( .A(n2946), .B(n2945), .Z(n969) );
  NAND U2970 ( .A(n970), .B(n969), .Z(n2947) );
  NAND U2971 ( .A(n2948), .B(n2947), .Z(n971) );
  NAND U2972 ( .A(n972), .B(n971), .Z(n2949) );
  NAND U2973 ( .A(n2950), .B(n2949), .Z(n973) );
  NAND U2974 ( .A(n974), .B(n973), .Z(n2951) );
  NAND U2975 ( .A(n2952), .B(n2951), .Z(n975) );
  NAND U2976 ( .A(n976), .B(n975), .Z(n2953) );
  NAND U2977 ( .A(n2954), .B(n2953), .Z(n977) );
  NAND U2978 ( .A(n978), .B(n977), .Z(n2955) );
  NAND U2979 ( .A(n2956), .B(n2955), .Z(n979) );
  NAND U2980 ( .A(n980), .B(n979), .Z(n2959) );
  NAND U2981 ( .A(n2960), .B(n2959), .Z(n981) );
  NAND U2982 ( .A(n982), .B(n981), .Z(n2961) );
  NAND U2983 ( .A(n2962), .B(n2961), .Z(n983) );
  NAND U2984 ( .A(n984), .B(n983), .Z(n2963) );
  NAND U2985 ( .A(n2964), .B(n2963), .Z(n985) );
  NAND U2986 ( .A(n986), .B(n985), .Z(n2965) );
  NAND U2987 ( .A(n2966), .B(n2965), .Z(n987) );
  NAND U2988 ( .A(n988), .B(n987), .Z(n2967) );
  NAND U2989 ( .A(n2968), .B(n2967), .Z(n989) );
  NAND U2990 ( .A(n990), .B(n989), .Z(n2969) );
  NAND U2991 ( .A(n2970), .B(n2969), .Z(n991) );
  NAND U2992 ( .A(n992), .B(n991), .Z(n2971) );
  NAND U2993 ( .A(n2972), .B(n2971), .Z(n993) );
  NAND U2994 ( .A(n994), .B(n993), .Z(n2973) );
  NAND U2995 ( .A(n2974), .B(n2973), .Z(n995) );
  NAND U2996 ( .A(n996), .B(n995), .Z(n2975) );
  NAND U2997 ( .A(n2976), .B(n2975), .Z(n997) );
  NAND U2998 ( .A(n998), .B(n997), .Z(n2977) );
  NAND U2999 ( .A(n2978), .B(n2977), .Z(n999) );
  NAND U3000 ( .A(n1000), .B(n999), .Z(n2983) );
  NAND U3001 ( .A(n2984), .B(n2983), .Z(n1001) );
  NAND U3002 ( .A(n1002), .B(n1001), .Z(n2985) );
  NAND U3003 ( .A(n2986), .B(n2985), .Z(n1003) );
  NAND U3004 ( .A(n1004), .B(n1003), .Z(n2987) );
  NAND U3005 ( .A(n2988), .B(n2987), .Z(n1005) );
  NAND U3006 ( .A(n1006), .B(n1005), .Z(n2989) );
  NAND U3007 ( .A(n2990), .B(n2989), .Z(n1007) );
  NAND U3008 ( .A(n1008), .B(n1007), .Z(n2991) );
  NAND U3009 ( .A(n2992), .B(n2991), .Z(n1009) );
  NAND U3010 ( .A(n1010), .B(n1009), .Z(n2993) );
  NAND U3011 ( .A(n2994), .B(n2993), .Z(n1011) );
  NAND U3012 ( .A(n1012), .B(n1011), .Z(n2995) );
  NAND U3013 ( .A(n2996), .B(n2995), .Z(n1013) );
  NAND U3014 ( .A(n1014), .B(n1013), .Z(n2997) );
  NAND U3015 ( .A(n2998), .B(n2997), .Z(n1015) );
  NAND U3016 ( .A(n1016), .B(n1015), .Z(n2999) );
  NAND U3017 ( .A(n3000), .B(n2999), .Z(n1017) );
  NAND U3018 ( .A(n1018), .B(n1017), .Z(n3001) );
  NAND U3019 ( .A(n3002), .B(n3001), .Z(n1019) );
  NAND U3020 ( .A(n1020), .B(n1019), .Z(n3005) );
  NAND U3021 ( .A(n3006), .B(n3005), .Z(n1021) );
  NAND U3022 ( .A(n1022), .B(n1021), .Z(n3007) );
  NAND U3023 ( .A(n3008), .B(n3007), .Z(n1023) );
  NAND U3024 ( .A(n1024), .B(n1023), .Z(n3009) );
  NAND U3025 ( .A(n3010), .B(n3009), .Z(n1025) );
  NAND U3026 ( .A(n1026), .B(n1025), .Z(n3011) );
  NAND U3027 ( .A(n3012), .B(n3011), .Z(n1027) );
  NAND U3028 ( .A(n1028), .B(n1027), .Z(n3013) );
  NAND U3029 ( .A(n3014), .B(n3013), .Z(n1029) );
  NAND U3030 ( .A(n1030), .B(n1029), .Z(n3015) );
  NAND U3031 ( .A(n3016), .B(n3015), .Z(n1031) );
  NAND U3032 ( .A(n1032), .B(n1031), .Z(n3017) );
  NAND U3033 ( .A(n3018), .B(n3017), .Z(n1033) );
  NAND U3034 ( .A(n1034), .B(n1033), .Z(n3019) );
  NAND U3035 ( .A(n3020), .B(n3019), .Z(n1035) );
  NAND U3036 ( .A(n1036), .B(n1035), .Z(n3021) );
  NAND U3037 ( .A(n3022), .B(n3021), .Z(n1037) );
  NAND U3038 ( .A(n1038), .B(n1037), .Z(n3023) );
  NAND U3039 ( .A(n3024), .B(n3023), .Z(n1039) );
  NAND U3040 ( .A(n1040), .B(n1039), .Z(n3027) );
  NAND U3041 ( .A(n3028), .B(n3027), .Z(n1041) );
  NAND U3042 ( .A(n1042), .B(n1041), .Z(n3029) );
  NAND U3043 ( .A(n3030), .B(n3029), .Z(n1043) );
  NAND U3044 ( .A(n1044), .B(n1043), .Z(n3031) );
  NAND U3045 ( .A(n3032), .B(n3031), .Z(n1045) );
  NAND U3046 ( .A(n1046), .B(n1045), .Z(n3033) );
  NAND U3047 ( .A(n3034), .B(n3033), .Z(n1047) );
  NAND U3048 ( .A(n1048), .B(n1047), .Z(n3035) );
  NAND U3049 ( .A(n3036), .B(n3035), .Z(n1049) );
  NAND U3050 ( .A(n1050), .B(n1049), .Z(n3037) );
  NAND U3051 ( .A(n3038), .B(n3037), .Z(n1051) );
  NAND U3052 ( .A(n1052), .B(n1051), .Z(n3039) );
  NAND U3053 ( .A(n3040), .B(n3039), .Z(n1053) );
  NAND U3054 ( .A(n1054), .B(n1053), .Z(n3041) );
  NAND U3055 ( .A(n3042), .B(n3041), .Z(n1055) );
  NAND U3056 ( .A(n1056), .B(n1055), .Z(n3043) );
  NAND U3057 ( .A(n3044), .B(n3043), .Z(n1057) );
  NAND U3058 ( .A(n1058), .B(n1057), .Z(n3045) );
  NAND U3059 ( .A(n3046), .B(n3045), .Z(n1059) );
  NAND U3060 ( .A(n1060), .B(n1059), .Z(n3049) );
  NAND U3061 ( .A(n3050), .B(n3049), .Z(n1061) );
  NAND U3062 ( .A(n1062), .B(n1061), .Z(n3051) );
  NAND U3063 ( .A(n3052), .B(n3051), .Z(n1063) );
  NAND U3064 ( .A(n1064), .B(n1063), .Z(n3053) );
  NAND U3065 ( .A(n3054), .B(n3053), .Z(n1065) );
  NAND U3066 ( .A(n1066), .B(n1065), .Z(n3055) );
  NAND U3067 ( .A(n3056), .B(n3055), .Z(n1067) );
  NAND U3068 ( .A(n1068), .B(n1067), .Z(n3057) );
  NAND U3069 ( .A(n3058), .B(n3057), .Z(n1069) );
  NAND U3070 ( .A(n1070), .B(n1069), .Z(n3059) );
  NAND U3071 ( .A(n3060), .B(n3059), .Z(n1071) );
  NAND U3072 ( .A(n1072), .B(n1071), .Z(n3061) );
  NAND U3073 ( .A(n3062), .B(n3061), .Z(n1073) );
  NAND U3074 ( .A(n1074), .B(n1073), .Z(n3063) );
  NAND U3075 ( .A(n3064), .B(n3063), .Z(n1075) );
  NAND U3076 ( .A(n1076), .B(n1075), .Z(n3065) );
  NAND U3077 ( .A(n3066), .B(n3065), .Z(n1077) );
  NAND U3078 ( .A(n1078), .B(n1077), .Z(n3067) );
  NAND U3079 ( .A(n3068), .B(n3067), .Z(n1079) );
  NAND U3080 ( .A(n1080), .B(n1079), .Z(n3071) );
  NAND U3081 ( .A(n3072), .B(n3071), .Z(n1081) );
  NAND U3082 ( .A(n1082), .B(n1081), .Z(n3073) );
  NAND U3083 ( .A(n3074), .B(n3073), .Z(n1083) );
  NAND U3084 ( .A(n1084), .B(n1083), .Z(n3075) );
  NAND U3085 ( .A(n3076), .B(n3075), .Z(n1085) );
  NAND U3086 ( .A(n1086), .B(n1085), .Z(n3077) );
  NAND U3087 ( .A(n3078), .B(n3077), .Z(n1087) );
  NAND U3088 ( .A(n1088), .B(n1087), .Z(n3079) );
  NAND U3089 ( .A(n3080), .B(n3079), .Z(n1089) );
  NAND U3090 ( .A(n1090), .B(n1089), .Z(n3081) );
  NAND U3091 ( .A(n3082), .B(n3081), .Z(n1091) );
  NAND U3092 ( .A(n1092), .B(n1091), .Z(n3083) );
  NAND U3093 ( .A(n3084), .B(n3083), .Z(n1093) );
  NAND U3094 ( .A(n1094), .B(n1093), .Z(n3085) );
  NAND U3095 ( .A(n3086), .B(n3085), .Z(n1095) );
  NAND U3096 ( .A(n1096), .B(n1095), .Z(n3087) );
  NAND U3097 ( .A(n3088), .B(n3087), .Z(n1097) );
  NAND U3098 ( .A(n1098), .B(n1097), .Z(n3089) );
  NAND U3099 ( .A(n3090), .B(n3089), .Z(n1099) );
  NAND U3100 ( .A(n1100), .B(n1099), .Z(n3093) );
  NAND U3101 ( .A(n3094), .B(n3093), .Z(n1101) );
  NAND U3102 ( .A(n1102), .B(n1101), .Z(n3095) );
  NAND U3103 ( .A(n3096), .B(n3095), .Z(n1103) );
  NAND U3104 ( .A(n1104), .B(n1103), .Z(n3097) );
  NAND U3105 ( .A(n3098), .B(n3097), .Z(n1105) );
  NAND U3106 ( .A(n1106), .B(n1105), .Z(n3099) );
  NAND U3107 ( .A(n3100), .B(n3099), .Z(n1107) );
  NAND U3108 ( .A(n1108), .B(n1107), .Z(n3101) );
  NAND U3109 ( .A(n3102), .B(n3101), .Z(n1109) );
  NAND U3110 ( .A(n1110), .B(n1109), .Z(n3103) );
  NAND U3111 ( .A(n3104), .B(n3103), .Z(n1111) );
  NAND U3112 ( .A(n1112), .B(n1111), .Z(n3105) );
  NAND U3113 ( .A(n3106), .B(n3105), .Z(n1113) );
  NAND U3114 ( .A(n1114), .B(n1113), .Z(n3107) );
  NAND U3115 ( .A(n3108), .B(n3107), .Z(n1115) );
  NAND U3116 ( .A(n1116), .B(n1115), .Z(n3109) );
  NAND U3117 ( .A(n3110), .B(n3109), .Z(n1117) );
  NAND U3118 ( .A(n1118), .B(n1117), .Z(n3111) );
  NAND U3119 ( .A(n3112), .B(n3111), .Z(n1119) );
  NAND U3120 ( .A(n1120), .B(n1119), .Z(n3115) );
  NAND U3121 ( .A(n3116), .B(n3115), .Z(n1121) );
  NAND U3122 ( .A(n1122), .B(n1121), .Z(n3117) );
  NAND U3123 ( .A(n3118), .B(n3117), .Z(n1123) );
  NAND U3124 ( .A(n1124), .B(n1123), .Z(n3119) );
  NAND U3125 ( .A(n3120), .B(n3119), .Z(n1125) );
  NAND U3126 ( .A(n1126), .B(n1125), .Z(n3121) );
  NAND U3127 ( .A(n3122), .B(n3121), .Z(n1127) );
  NAND U3128 ( .A(n1128), .B(n1127), .Z(n3123) );
  NAND U3129 ( .A(n3124), .B(n3123), .Z(n1129) );
  NAND U3130 ( .A(n1130), .B(n1129), .Z(n3125) );
  NAND U3131 ( .A(n3126), .B(n3125), .Z(n1131) );
  NAND U3132 ( .A(n1132), .B(n1131), .Z(n3127) );
  NAND U3133 ( .A(n3128), .B(n3127), .Z(n1133) );
  NAND U3134 ( .A(n1134), .B(n1133), .Z(n3129) );
  NAND U3135 ( .A(n3130), .B(n3129), .Z(n1135) );
  NAND U3136 ( .A(n1136), .B(n1135), .Z(n3131) );
  NAND U3137 ( .A(n3132), .B(n3131), .Z(n1137) );
  NAND U3138 ( .A(n1138), .B(n1137), .Z(n3133) );
  NAND U3139 ( .A(n3134), .B(n3133), .Z(n1139) );
  NAND U3140 ( .A(n1140), .B(n1139), .Z(n3137) );
  NAND U3141 ( .A(n3138), .B(n3137), .Z(n1141) );
  NAND U3142 ( .A(n1142), .B(n1141), .Z(n3139) );
  NAND U3143 ( .A(n3140), .B(n3139), .Z(n1143) );
  NAND U3144 ( .A(n1144), .B(n1143), .Z(n3141) );
  NAND U3145 ( .A(n3142), .B(n3141), .Z(n1145) );
  NAND U3146 ( .A(n1146), .B(n1145), .Z(n3143) );
  NAND U3147 ( .A(n3144), .B(n3143), .Z(n1147) );
  NAND U3148 ( .A(n1148), .B(n1147), .Z(n3145) );
  NAND U3149 ( .A(n3146), .B(n3145), .Z(n1149) );
  NAND U3150 ( .A(n1150), .B(n1149), .Z(n3147) );
  NAND U3151 ( .A(n3148), .B(n3147), .Z(n1151) );
  NAND U3152 ( .A(n1152), .B(n1151), .Z(n3149) );
  NAND U3153 ( .A(n3150), .B(n3149), .Z(n1153) );
  NAND U3154 ( .A(n1154), .B(n1153), .Z(n3151) );
  NAND U3155 ( .A(n3152), .B(n3151), .Z(n1155) );
  NAND U3156 ( .A(n1156), .B(n1155), .Z(n3153) );
  NAND U3157 ( .A(n3154), .B(n3153), .Z(n1157) );
  NAND U3158 ( .A(n1158), .B(n1157), .Z(n3155) );
  NAND U3159 ( .A(n3156), .B(n3155), .Z(n1159) );
  NAND U3160 ( .A(n1160), .B(n1159), .Z(n3159) );
  NAND U3161 ( .A(n3160), .B(n3159), .Z(n1161) );
  NAND U3162 ( .A(n1162), .B(n1161), .Z(n3161) );
  NAND U3163 ( .A(n3162), .B(n3161), .Z(n1163) );
  NAND U3164 ( .A(n1164), .B(n1163), .Z(n3163) );
  NAND U3165 ( .A(n3164), .B(n3163), .Z(n1165) );
  NAND U3166 ( .A(n1166), .B(n1165), .Z(n3165) );
  NAND U3167 ( .A(n3166), .B(n3165), .Z(n1167) );
  NAND U3168 ( .A(n1168), .B(n1167), .Z(n3167) );
  NAND U3169 ( .A(n3168), .B(n3167), .Z(n1169) );
  NAND U3170 ( .A(n1170), .B(n1169), .Z(n3169) );
  NAND U3171 ( .A(n3170), .B(n3169), .Z(n1171) );
  NAND U3172 ( .A(n1172), .B(n1171), .Z(n3171) );
  NAND U3173 ( .A(n3172), .B(n3171), .Z(n1173) );
  NAND U3174 ( .A(n1174), .B(n1173), .Z(n3173) );
  NAND U3175 ( .A(n3174), .B(n3173), .Z(n1175) );
  NAND U3176 ( .A(n1176), .B(n1175), .Z(n3175) );
  NAND U3177 ( .A(n3176), .B(n3175), .Z(n1177) );
  NAND U3178 ( .A(n1178), .B(n1177), .Z(n3177) );
  NAND U3179 ( .A(n3178), .B(n3177), .Z(n1179) );
  NAND U3180 ( .A(n1180), .B(n1179), .Z(n3181) );
  NAND U3181 ( .A(n3182), .B(n3181), .Z(n1181) );
  NAND U3182 ( .A(n1182), .B(n1181), .Z(n3183) );
  NAND U3183 ( .A(n3184), .B(n3183), .Z(n1183) );
  NAND U3184 ( .A(n1184), .B(n1183), .Z(n3185) );
  NAND U3185 ( .A(n3186), .B(n3185), .Z(n1185) );
  NAND U3186 ( .A(n1186), .B(n1185), .Z(n3187) );
  NAND U3187 ( .A(n3188), .B(n3187), .Z(n1187) );
  NAND U3188 ( .A(n1188), .B(n1187), .Z(n3189) );
  NAND U3189 ( .A(n3190), .B(n3189), .Z(n1189) );
  NAND U3190 ( .A(n1190), .B(n1189), .Z(n3191) );
  NAND U3191 ( .A(n3192), .B(n3191), .Z(n1191) );
  NAND U3192 ( .A(n1192), .B(n1191), .Z(n3193) );
  NAND U3193 ( .A(n3194), .B(n3193), .Z(n1193) );
  NAND U3194 ( .A(n1194), .B(n1193), .Z(n3195) );
  NAND U3195 ( .A(n3196), .B(n3195), .Z(n1195) );
  NAND U3196 ( .A(n1196), .B(n1195), .Z(n3197) );
  NAND U3197 ( .A(n3198), .B(n3197), .Z(n1197) );
  NAND U3198 ( .A(n1198), .B(n1197), .Z(n3199) );
  NAND U3199 ( .A(n3200), .B(n3199), .Z(n1199) );
  NAND U3200 ( .A(n1200), .B(n1199), .Z(n3205) );
  NAND U3201 ( .A(n3206), .B(n3205), .Z(n1201) );
  NAND U3202 ( .A(n1202), .B(n1201), .Z(n3207) );
  NAND U3203 ( .A(n3208), .B(n3207), .Z(n1203) );
  NAND U3204 ( .A(n1204), .B(n1203), .Z(n3209) );
  NAND U3205 ( .A(n3210), .B(n3209), .Z(n1205) );
  NAND U3206 ( .A(n1206), .B(n1205), .Z(n3211) );
  NAND U3207 ( .A(n3212), .B(n3211), .Z(n1207) );
  NAND U3208 ( .A(n1208), .B(n1207), .Z(n3213) );
  NAND U3209 ( .A(n3214), .B(n3213), .Z(n1209) );
  NAND U3210 ( .A(n1210), .B(n1209), .Z(n3215) );
  NAND U3211 ( .A(n3216), .B(n3215), .Z(n1211) );
  NAND U3212 ( .A(n1212), .B(n1211), .Z(n3217) );
  NAND U3213 ( .A(n3218), .B(n3217), .Z(n1213) );
  NAND U3214 ( .A(n1214), .B(n1213), .Z(n3219) );
  NAND U3215 ( .A(n3220), .B(n3219), .Z(n1215) );
  NAND U3216 ( .A(n1216), .B(n1215), .Z(n3221) );
  NAND U3217 ( .A(n3222), .B(n3221), .Z(n1217) );
  NAND U3218 ( .A(n1218), .B(n1217), .Z(n3223) );
  NAND U3219 ( .A(n3224), .B(n3223), .Z(n1219) );
  NAND U3220 ( .A(n1220), .B(n1219), .Z(n3227) );
  NAND U3221 ( .A(n3228), .B(n3227), .Z(n1221) );
  NAND U3222 ( .A(n1222), .B(n1221), .Z(n3229) );
  NAND U3223 ( .A(n3230), .B(n3229), .Z(n1223) );
  NAND U3224 ( .A(n1224), .B(n1223), .Z(n3231) );
  NAND U3225 ( .A(n3232), .B(n3231), .Z(n1225) );
  NAND U3226 ( .A(n1226), .B(n1225), .Z(n3233) );
  NAND U3227 ( .A(n3234), .B(n3233), .Z(n1227) );
  NAND U3228 ( .A(n1228), .B(n1227), .Z(n3235) );
  NAND U3229 ( .A(n3236), .B(n3235), .Z(n1229) );
  NAND U3230 ( .A(n1230), .B(n1229), .Z(n3237) );
  NAND U3231 ( .A(n3238), .B(n3237), .Z(n1231) );
  NAND U3232 ( .A(n1232), .B(n1231), .Z(n3239) );
  NAND U3233 ( .A(n3240), .B(n3239), .Z(n1233) );
  NAND U3234 ( .A(n1234), .B(n1233), .Z(n3241) );
  NAND U3235 ( .A(n3242), .B(n3241), .Z(n1235) );
  NAND U3236 ( .A(n1236), .B(n1235), .Z(n3243) );
  NAND U3237 ( .A(n3244), .B(n3243), .Z(n1237) );
  NAND U3238 ( .A(n1238), .B(n1237), .Z(n3245) );
  NAND U3239 ( .A(n3246), .B(n3245), .Z(n1239) );
  NAND U3240 ( .A(n1240), .B(n1239), .Z(n3249) );
  NAND U3241 ( .A(n3250), .B(n3249), .Z(n1241) );
  NAND U3242 ( .A(n1242), .B(n1241), .Z(n3251) );
  NAND U3243 ( .A(n3252), .B(n3251), .Z(n1243) );
  NAND U3244 ( .A(n1244), .B(n1243), .Z(n3253) );
  NAND U3245 ( .A(n3254), .B(n3253), .Z(n1245) );
  NAND U3246 ( .A(n1246), .B(n1245), .Z(n3255) );
  NAND U3247 ( .A(n3256), .B(n3255), .Z(n1247) );
  NAND U3248 ( .A(n1248), .B(n1247), .Z(n3257) );
  NAND U3249 ( .A(n3258), .B(n3257), .Z(n1249) );
  NAND U3250 ( .A(n1250), .B(n1249), .Z(n3259) );
  NAND U3251 ( .A(n3260), .B(n3259), .Z(n1251) );
  NAND U3252 ( .A(n1252), .B(n1251), .Z(n3261) );
  NAND U3253 ( .A(n3262), .B(n3261), .Z(n1253) );
  NAND U3254 ( .A(n1254), .B(n1253), .Z(n3263) );
  NAND U3255 ( .A(n3264), .B(n3263), .Z(n1255) );
  NAND U3256 ( .A(n1256), .B(n1255), .Z(n3265) );
  NAND U3257 ( .A(n3266), .B(n3265), .Z(n1257) );
  NAND U3258 ( .A(n1258), .B(n1257), .Z(n3267) );
  NAND U3259 ( .A(n3268), .B(n3267), .Z(n1259) );
  NAND U3260 ( .A(n1260), .B(n1259), .Z(n3271) );
  NAND U3261 ( .A(n3272), .B(n3271), .Z(n1261) );
  NAND U3262 ( .A(n1262), .B(n1261), .Z(n3273) );
  NAND U3263 ( .A(n3274), .B(n3273), .Z(n1263) );
  NAND U3264 ( .A(n1264), .B(n1263), .Z(n3275) );
  NAND U3265 ( .A(n3276), .B(n3275), .Z(n1265) );
  NAND U3266 ( .A(n1266), .B(n1265), .Z(n3277) );
  NAND U3267 ( .A(n3278), .B(n3277), .Z(n1267) );
  NAND U3268 ( .A(n1268), .B(n1267), .Z(n3279) );
  NAND U3269 ( .A(n3280), .B(n3279), .Z(n1269) );
  NAND U3270 ( .A(n1270), .B(n1269), .Z(n3281) );
  NAND U3271 ( .A(n3282), .B(n3281), .Z(n1271) );
  NAND U3272 ( .A(n1272), .B(n1271), .Z(n3283) );
  NAND U3273 ( .A(n3284), .B(n3283), .Z(n1273) );
  NAND U3274 ( .A(n1274), .B(n1273), .Z(n3285) );
  NAND U3275 ( .A(n3286), .B(n3285), .Z(n1275) );
  NAND U3276 ( .A(n1276), .B(n1275), .Z(n3287) );
  NAND U3277 ( .A(n3288), .B(n3287), .Z(n1277) );
  NAND U3278 ( .A(n1278), .B(n1277), .Z(n3289) );
  NAND U3279 ( .A(n3290), .B(n3289), .Z(n1279) );
  NAND U3280 ( .A(n1280), .B(n1279), .Z(n3293) );
  NAND U3281 ( .A(n3294), .B(n3293), .Z(n1281) );
  NAND U3282 ( .A(n1282), .B(n1281), .Z(n3295) );
  NAND U3283 ( .A(n3296), .B(n3295), .Z(n1283) );
  NAND U3284 ( .A(n1284), .B(n1283), .Z(n3297) );
  NAND U3285 ( .A(n3298), .B(n3297), .Z(n1285) );
  NAND U3286 ( .A(n1286), .B(n1285), .Z(n3299) );
  NAND U3287 ( .A(n3300), .B(n3299), .Z(n1287) );
  NAND U3288 ( .A(n1288), .B(n1287), .Z(n3301) );
  NAND U3289 ( .A(n3302), .B(n3301), .Z(n1289) );
  NAND U3290 ( .A(n1290), .B(n1289), .Z(n3303) );
  NAND U3291 ( .A(n3304), .B(n3303), .Z(n1291) );
  NAND U3292 ( .A(n1292), .B(n1291), .Z(n3305) );
  NAND U3293 ( .A(n3306), .B(n3305), .Z(n1293) );
  NAND U3294 ( .A(n1294), .B(n1293), .Z(n3307) );
  NAND U3295 ( .A(n3308), .B(n3307), .Z(n1295) );
  NAND U3296 ( .A(n1296), .B(n1295), .Z(n3309) );
  NAND U3297 ( .A(n3310), .B(n3309), .Z(n1297) );
  NAND U3298 ( .A(n1298), .B(n1297), .Z(n3311) );
  NAND U3299 ( .A(n3312), .B(n3311), .Z(n1299) );
  NAND U3300 ( .A(n1300), .B(n1299), .Z(n3315) );
  NAND U3301 ( .A(n3316), .B(n3315), .Z(n1301) );
  NAND U3302 ( .A(n1302), .B(n1301), .Z(n3317) );
  NAND U3303 ( .A(n3318), .B(n3317), .Z(n1303) );
  NAND U3304 ( .A(n1304), .B(n1303), .Z(n3319) );
  NAND U3305 ( .A(n3320), .B(n3319), .Z(n1305) );
  NAND U3306 ( .A(n1306), .B(n1305), .Z(n3321) );
  NAND U3307 ( .A(n3322), .B(n3321), .Z(n1307) );
  NAND U3308 ( .A(n1308), .B(n1307), .Z(n3323) );
  NAND U3309 ( .A(n3324), .B(n3323), .Z(n1309) );
  NAND U3310 ( .A(n1310), .B(n1309), .Z(n3325) );
  NAND U3311 ( .A(n3326), .B(n3325), .Z(n1311) );
  NAND U3312 ( .A(n1312), .B(n1311), .Z(n3327) );
  NAND U3313 ( .A(n3328), .B(n3327), .Z(n1313) );
  NAND U3314 ( .A(n1314), .B(n1313), .Z(n3329) );
  NAND U3315 ( .A(n3330), .B(n3329), .Z(n1315) );
  NAND U3316 ( .A(n1316), .B(n1315), .Z(n3331) );
  NAND U3317 ( .A(n3332), .B(n3331), .Z(n1317) );
  NAND U3318 ( .A(n1318), .B(n1317), .Z(n3333) );
  NAND U3319 ( .A(n3334), .B(n3333), .Z(n1319) );
  NAND U3320 ( .A(n1320), .B(n1319), .Z(n3337) );
  NAND U3321 ( .A(n3338), .B(n3337), .Z(n1321) );
  NAND U3322 ( .A(n1322), .B(n1321), .Z(n3339) );
  NAND U3323 ( .A(n3340), .B(n3339), .Z(n1323) );
  NAND U3324 ( .A(n1324), .B(n1323), .Z(n3341) );
  NAND U3325 ( .A(n3342), .B(n3341), .Z(n1325) );
  NAND U3326 ( .A(n1326), .B(n1325), .Z(n3343) );
  NAND U3327 ( .A(n3344), .B(n3343), .Z(n1327) );
  NAND U3328 ( .A(n1328), .B(n1327), .Z(n3345) );
  NAND U3329 ( .A(n3346), .B(n3345), .Z(n1329) );
  NAND U3330 ( .A(n1330), .B(n1329), .Z(n3347) );
  NAND U3331 ( .A(n3348), .B(n3347), .Z(n1331) );
  NAND U3332 ( .A(n1332), .B(n1331), .Z(n3349) );
  NAND U3333 ( .A(n3350), .B(n3349), .Z(n1333) );
  NAND U3334 ( .A(n1334), .B(n1333), .Z(n3351) );
  NAND U3335 ( .A(n3352), .B(n3351), .Z(n1335) );
  NAND U3336 ( .A(n1336), .B(n1335), .Z(n3353) );
  NAND U3337 ( .A(n3354), .B(n3353), .Z(n1337) );
  NAND U3338 ( .A(n1338), .B(n1337), .Z(n3355) );
  NAND U3339 ( .A(n3356), .B(n3355), .Z(n1339) );
  NAND U3340 ( .A(n1340), .B(n1339), .Z(n3359) );
  NAND U3341 ( .A(n3360), .B(n3359), .Z(n1341) );
  NAND U3342 ( .A(n1342), .B(n1341), .Z(n3361) );
  NAND U3343 ( .A(n3362), .B(n3361), .Z(n1343) );
  NAND U3344 ( .A(n1344), .B(n1343), .Z(n3363) );
  NAND U3345 ( .A(n3364), .B(n3363), .Z(n1345) );
  NAND U3346 ( .A(n1346), .B(n1345), .Z(n3365) );
  NAND U3347 ( .A(n3366), .B(n3365), .Z(n1347) );
  NAND U3348 ( .A(n1348), .B(n1347), .Z(n3367) );
  NAND U3349 ( .A(n3368), .B(n3367), .Z(n1349) );
  NAND U3350 ( .A(n1350), .B(n1349), .Z(n3369) );
  NAND U3351 ( .A(n3370), .B(n3369), .Z(n1351) );
  NAND U3352 ( .A(n1352), .B(n1351), .Z(n3371) );
  NAND U3353 ( .A(n3372), .B(n3371), .Z(n1353) );
  NAND U3354 ( .A(n1354), .B(n1353), .Z(n3373) );
  NAND U3355 ( .A(n3374), .B(n3373), .Z(n1355) );
  NAND U3356 ( .A(n1356), .B(n1355), .Z(n3375) );
  NAND U3357 ( .A(n3376), .B(n3375), .Z(n1357) );
  NAND U3358 ( .A(n1358), .B(n1357), .Z(n3377) );
  NAND U3359 ( .A(n3378), .B(n3377), .Z(n1359) );
  NAND U3360 ( .A(n1360), .B(n1359), .Z(n3381) );
  NAND U3361 ( .A(n3382), .B(n3381), .Z(n1361) );
  NAND U3362 ( .A(n1362), .B(n1361), .Z(n3383) );
  NAND U3363 ( .A(n3384), .B(n3383), .Z(n1363) );
  NAND U3364 ( .A(n1364), .B(n1363), .Z(n3385) );
  NAND U3365 ( .A(n3386), .B(n3385), .Z(n1365) );
  NAND U3366 ( .A(n1366), .B(n1365), .Z(n3387) );
  NAND U3367 ( .A(n3388), .B(n3387), .Z(n1367) );
  NAND U3368 ( .A(n1368), .B(n1367), .Z(n3389) );
  NAND U3369 ( .A(n3390), .B(n3389), .Z(n1369) );
  NAND U3370 ( .A(n1370), .B(n1369), .Z(n3391) );
  NAND U3371 ( .A(n3392), .B(n3391), .Z(n1371) );
  NAND U3372 ( .A(n1372), .B(n1371), .Z(n3393) );
  NAND U3373 ( .A(n3394), .B(n3393), .Z(n1373) );
  NAND U3374 ( .A(n1374), .B(n1373), .Z(n3395) );
  NAND U3375 ( .A(n3396), .B(n3395), .Z(n1375) );
  NAND U3376 ( .A(n1376), .B(n1375), .Z(n3397) );
  NAND U3377 ( .A(n3398), .B(n3397), .Z(n1377) );
  NAND U3378 ( .A(n1378), .B(n1377), .Z(n3399) );
  NAND U3379 ( .A(n3400), .B(n3399), .Z(n1379) );
  NAND U3380 ( .A(n1380), .B(n1379), .Z(n3403) );
  NAND U3381 ( .A(n3404), .B(n3403), .Z(n1381) );
  NAND U3382 ( .A(n1382), .B(n1381), .Z(n3405) );
  NAND U3383 ( .A(n3406), .B(n3405), .Z(n1383) );
  NAND U3384 ( .A(n1384), .B(n1383), .Z(n3407) );
  NAND U3385 ( .A(n3408), .B(n3407), .Z(n1385) );
  NAND U3386 ( .A(n1386), .B(n1385), .Z(n3409) );
  NAND U3387 ( .A(n3410), .B(n3409), .Z(n1387) );
  NAND U3388 ( .A(n1388), .B(n1387), .Z(n3411) );
  NAND U3389 ( .A(n3412), .B(n3411), .Z(n1389) );
  NAND U3390 ( .A(n1390), .B(n1389), .Z(n3413) );
  NAND U3391 ( .A(n3414), .B(n3413), .Z(n1391) );
  NAND U3392 ( .A(n1392), .B(n1391), .Z(n3415) );
  NAND U3393 ( .A(n3416), .B(n3415), .Z(n1393) );
  NAND U3394 ( .A(n1394), .B(n1393), .Z(n3417) );
  NAND U3395 ( .A(n3418), .B(n3417), .Z(n1395) );
  NAND U3396 ( .A(n1396), .B(n1395), .Z(n3419) );
  NAND U3397 ( .A(n3420), .B(n3419), .Z(n1397) );
  NAND U3398 ( .A(n1398), .B(n1397), .Z(n3421) );
  NAND U3399 ( .A(n3422), .B(n3421), .Z(n1399) );
  NAND U3400 ( .A(n1400), .B(n1399), .Z(n3427) );
  NAND U3401 ( .A(n3428), .B(n3427), .Z(n1401) );
  NAND U3402 ( .A(n1402), .B(n1401), .Z(n3429) );
  NAND U3403 ( .A(n3430), .B(n3429), .Z(n1403) );
  NAND U3404 ( .A(n1404), .B(n1403), .Z(n3431) );
  NAND U3405 ( .A(n3432), .B(n3431), .Z(n1405) );
  NAND U3406 ( .A(n1406), .B(n1405), .Z(n3433) );
  NAND U3407 ( .A(n3434), .B(n3433), .Z(n1407) );
  NAND U3408 ( .A(n1408), .B(n1407), .Z(n3435) );
  NAND U3409 ( .A(n3436), .B(n3435), .Z(n1409) );
  NAND U3410 ( .A(n1410), .B(n1409), .Z(n3437) );
  NAND U3411 ( .A(n3438), .B(n3437), .Z(n1411) );
  NAND U3412 ( .A(n1412), .B(n1411), .Z(n3439) );
  NAND U3413 ( .A(n3440), .B(n3439), .Z(n1413) );
  NAND U3414 ( .A(n1414), .B(n1413), .Z(n3441) );
  NAND U3415 ( .A(n3442), .B(n3441), .Z(n1415) );
  NAND U3416 ( .A(n1416), .B(n1415), .Z(n3443) );
  NAND U3417 ( .A(n3444), .B(n3443), .Z(n1417) );
  NAND U3418 ( .A(n1418), .B(n1417), .Z(n3445) );
  NAND U3419 ( .A(n3446), .B(n3445), .Z(n1419) );
  NAND U3420 ( .A(n1420), .B(n1419), .Z(n3449) );
  NAND U3421 ( .A(n3450), .B(n3449), .Z(n1421) );
  NAND U3422 ( .A(n1422), .B(n1421), .Z(n3451) );
  NAND U3423 ( .A(n3452), .B(n3451), .Z(n1423) );
  NAND U3424 ( .A(n1424), .B(n1423), .Z(n3453) );
  NAND U3425 ( .A(n3454), .B(n3453), .Z(n1425) );
  NAND U3426 ( .A(n1426), .B(n1425), .Z(n3455) );
  NAND U3427 ( .A(n3456), .B(n3455), .Z(n1427) );
  NAND U3428 ( .A(n1428), .B(n1427), .Z(n3457) );
  NAND U3429 ( .A(n3458), .B(n3457), .Z(n1429) );
  NAND U3430 ( .A(n1430), .B(n1429), .Z(n3459) );
  NAND U3431 ( .A(n3460), .B(n3459), .Z(n1431) );
  NAND U3432 ( .A(n1432), .B(n1431), .Z(n3461) );
  NAND U3433 ( .A(n3462), .B(n3461), .Z(n1433) );
  NAND U3434 ( .A(n1434), .B(n1433), .Z(n3463) );
  NAND U3435 ( .A(n3464), .B(n3463), .Z(n1435) );
  NAND U3436 ( .A(n1436), .B(n1435), .Z(n3465) );
  NAND U3437 ( .A(n3466), .B(n3465), .Z(n1437) );
  NAND U3438 ( .A(n1438), .B(n1437), .Z(n3467) );
  NAND U3439 ( .A(n3468), .B(n3467), .Z(n1439) );
  NAND U3440 ( .A(n1440), .B(n1439), .Z(n3471) );
  NAND U3441 ( .A(n3472), .B(n3471), .Z(n1441) );
  NAND U3442 ( .A(n1442), .B(n1441), .Z(n3473) );
  NAND U3443 ( .A(n3474), .B(n3473), .Z(n1443) );
  NAND U3444 ( .A(n1444), .B(n1443), .Z(n3475) );
  NAND U3445 ( .A(n3476), .B(n3475), .Z(n1445) );
  NAND U3446 ( .A(n1446), .B(n1445), .Z(n3477) );
  NAND U3447 ( .A(n3478), .B(n3477), .Z(n1447) );
  NAND U3448 ( .A(n1448), .B(n1447), .Z(n3479) );
  NAND U3449 ( .A(n3480), .B(n3479), .Z(n1449) );
  NAND U3450 ( .A(n1450), .B(n1449), .Z(n3481) );
  NAND U3451 ( .A(n3482), .B(n3481), .Z(n1451) );
  NAND U3452 ( .A(n1452), .B(n1451), .Z(n3483) );
  NAND U3453 ( .A(n3484), .B(n3483), .Z(n1453) );
  NAND U3454 ( .A(n1454), .B(n1453), .Z(n3485) );
  NAND U3455 ( .A(n3486), .B(n3485), .Z(n1455) );
  NAND U3456 ( .A(n1456), .B(n1455), .Z(n3487) );
  NAND U3457 ( .A(n3488), .B(n3487), .Z(n1457) );
  NAND U3458 ( .A(n1458), .B(n1457), .Z(n3489) );
  NAND U3459 ( .A(n3490), .B(n3489), .Z(n1459) );
  NAND U3460 ( .A(n1460), .B(n1459), .Z(n3493) );
  NAND U3461 ( .A(n3494), .B(n3493), .Z(n1461) );
  NAND U3462 ( .A(n1462), .B(n1461), .Z(n3495) );
  NAND U3463 ( .A(n3496), .B(n3495), .Z(n1463) );
  NAND U3464 ( .A(n1464), .B(n1463), .Z(n3497) );
  NAND U3465 ( .A(n3498), .B(n3497), .Z(n1465) );
  NAND U3466 ( .A(n1466), .B(n1465), .Z(n3499) );
  NAND U3467 ( .A(n3500), .B(n3499), .Z(n1467) );
  NAND U3468 ( .A(n1468), .B(n1467), .Z(n3501) );
  NAND U3469 ( .A(n3502), .B(n3501), .Z(n1469) );
  NAND U3470 ( .A(n1470), .B(n1469), .Z(n3503) );
  NAND U3471 ( .A(n3504), .B(n3503), .Z(n1471) );
  NAND U3472 ( .A(n1472), .B(n1471), .Z(n3505) );
  NAND U3473 ( .A(n3506), .B(n3505), .Z(n1473) );
  NAND U3474 ( .A(n1474), .B(n1473), .Z(n3507) );
  NAND U3475 ( .A(n3508), .B(n3507), .Z(n1475) );
  NAND U3476 ( .A(n1476), .B(n1475), .Z(n3509) );
  NAND U3477 ( .A(n3510), .B(n3509), .Z(n1477) );
  NAND U3478 ( .A(n1478), .B(n1477), .Z(n3511) );
  NAND U3479 ( .A(n3512), .B(n3511), .Z(n1479) );
  NAND U3480 ( .A(n1480), .B(n1479), .Z(n3515) );
  NAND U3481 ( .A(n3516), .B(n3515), .Z(n1481) );
  NAND U3482 ( .A(n1482), .B(n1481), .Z(n3517) );
  NAND U3483 ( .A(n3518), .B(n3517), .Z(n1483) );
  NAND U3484 ( .A(n1484), .B(n1483), .Z(n3519) );
  NAND U3485 ( .A(n3520), .B(n3519), .Z(n1485) );
  NAND U3486 ( .A(n1486), .B(n1485), .Z(n3521) );
  NAND U3487 ( .A(n3522), .B(n3521), .Z(n1487) );
  NAND U3488 ( .A(n1488), .B(n1487), .Z(n3523) );
  NAND U3489 ( .A(n3524), .B(n3523), .Z(n1489) );
  NAND U3490 ( .A(n1490), .B(n1489), .Z(n3525) );
  NAND U3491 ( .A(n3526), .B(n3525), .Z(n1491) );
  NAND U3492 ( .A(n1492), .B(n1491), .Z(n3527) );
  NAND U3493 ( .A(n3528), .B(n3527), .Z(n1493) );
  NAND U3494 ( .A(n1494), .B(n1493), .Z(n3529) );
  NAND U3495 ( .A(n3530), .B(n3529), .Z(n1495) );
  NAND U3496 ( .A(n1496), .B(n1495), .Z(n3531) );
  NAND U3497 ( .A(n3532), .B(n3531), .Z(n1497) );
  NAND U3498 ( .A(n1498), .B(n1497), .Z(n3533) );
  NAND U3499 ( .A(n3534), .B(n3533), .Z(n1499) );
  NAND U3500 ( .A(n1500), .B(n1499), .Z(n3537) );
  NAND U3501 ( .A(n3538), .B(n3537), .Z(n1501) );
  NAND U3502 ( .A(n1502), .B(n1501), .Z(n3539) );
  NAND U3503 ( .A(n3540), .B(n3539), .Z(n1503) );
  NAND U3504 ( .A(n1504), .B(n1503), .Z(n3541) );
  NAND U3505 ( .A(n3542), .B(n3541), .Z(n1505) );
  NAND U3506 ( .A(n1506), .B(n1505), .Z(n3543) );
  NAND U3507 ( .A(n3544), .B(n3543), .Z(n1507) );
  NAND U3508 ( .A(n1508), .B(n1507), .Z(n3545) );
  NAND U3509 ( .A(n3546), .B(n3545), .Z(n1509) );
  NAND U3510 ( .A(n1510), .B(n1509), .Z(n3547) );
  NAND U3511 ( .A(n3548), .B(n3547), .Z(n1511) );
  NAND U3512 ( .A(n1512), .B(n1511), .Z(n3549) );
  NAND U3513 ( .A(n3550), .B(n3549), .Z(n1513) );
  NAND U3514 ( .A(n1514), .B(n1513), .Z(n3551) );
  NAND U3515 ( .A(n3552), .B(n3551), .Z(n1515) );
  NAND U3516 ( .A(n1516), .B(n1515), .Z(n3553) );
  NAND U3517 ( .A(n3554), .B(n3553), .Z(n1517) );
  NAND U3518 ( .A(n1518), .B(n1517), .Z(n3555) );
  NAND U3519 ( .A(n3556), .B(n3555), .Z(n1519) );
  NAND U3520 ( .A(n1520), .B(n1519), .Z(n3559) );
  NAND U3521 ( .A(n3560), .B(n3559), .Z(n1521) );
  NAND U3522 ( .A(n1522), .B(n1521), .Z(n3561) );
  NAND U3523 ( .A(n3562), .B(n3561), .Z(n1523) );
  NAND U3524 ( .A(n1524), .B(n1523), .Z(n3563) );
  NAND U3525 ( .A(n3564), .B(n3563), .Z(n1525) );
  NAND U3526 ( .A(n1526), .B(n1525), .Z(n3565) );
  NAND U3527 ( .A(n3566), .B(n3565), .Z(n1527) );
  NAND U3528 ( .A(n1528), .B(n1527), .Z(n3567) );
  NAND U3529 ( .A(n3568), .B(n3567), .Z(n1529) );
  NAND U3530 ( .A(n1530), .B(n1529), .Z(n3569) );
  NAND U3531 ( .A(n3570), .B(n3569), .Z(n1531) );
  NAND U3532 ( .A(n1532), .B(n1531), .Z(n3571) );
  NAND U3533 ( .A(n3572), .B(n3571), .Z(n1533) );
  NAND U3534 ( .A(n1534), .B(n1533), .Z(n3573) );
  NAND U3535 ( .A(n3574), .B(n3573), .Z(n1535) );
  NAND U3536 ( .A(n1536), .B(n1535), .Z(n3575) );
  NAND U3537 ( .A(n3576), .B(n3575), .Z(n1537) );
  NAND U3538 ( .A(n1538), .B(n1537), .Z(n3577) );
  NAND U3539 ( .A(n3578), .B(n3577), .Z(n1539) );
  NAND U3540 ( .A(n1540), .B(n1539), .Z(n3581) );
  NAND U3541 ( .A(n3582), .B(n3581), .Z(n1541) );
  NAND U3542 ( .A(n1542), .B(n1541), .Z(n3583) );
  NAND U3543 ( .A(n3584), .B(n3583), .Z(n1543) );
  NAND U3544 ( .A(n1544), .B(n1543), .Z(n3585) );
  NAND U3545 ( .A(n3586), .B(n3585), .Z(n1545) );
  NAND U3546 ( .A(n1546), .B(n1545), .Z(n3587) );
  NAND U3547 ( .A(n3588), .B(n3587), .Z(n1547) );
  NAND U3548 ( .A(n1548), .B(n1547), .Z(n3589) );
  NAND U3549 ( .A(n3590), .B(n3589), .Z(n1549) );
  NAND U3550 ( .A(n1550), .B(n1549), .Z(n3591) );
  NAND U3551 ( .A(n3592), .B(n3591), .Z(n1551) );
  NAND U3552 ( .A(n1552), .B(n1551), .Z(n3593) );
  NAND U3553 ( .A(n3594), .B(n3593), .Z(n1553) );
  NAND U3554 ( .A(n1554), .B(n1553), .Z(n3595) );
  NAND U3555 ( .A(n3596), .B(n3595), .Z(n1555) );
  NAND U3556 ( .A(n1556), .B(n1555), .Z(n3597) );
  NAND U3557 ( .A(n3598), .B(n3597), .Z(n1557) );
  NAND U3558 ( .A(n1558), .B(n1557), .Z(n3599) );
  NAND U3559 ( .A(n3600), .B(n3599), .Z(n1559) );
  NAND U3560 ( .A(n1560), .B(n1559), .Z(n3603) );
  NAND U3561 ( .A(n3604), .B(n3603), .Z(n1561) );
  NAND U3562 ( .A(n1562), .B(n1561), .Z(n3605) );
  NAND U3563 ( .A(n3606), .B(n3605), .Z(n1563) );
  NAND U3564 ( .A(n1564), .B(n1563), .Z(n3607) );
  NAND U3565 ( .A(n3608), .B(n3607), .Z(n1565) );
  NAND U3566 ( .A(n1566), .B(n1565), .Z(n3609) );
  NAND U3567 ( .A(n3610), .B(n3609), .Z(n1567) );
  NAND U3568 ( .A(n1568), .B(n1567), .Z(n3611) );
  NAND U3569 ( .A(n3612), .B(n3611), .Z(n1569) );
  NAND U3570 ( .A(n1570), .B(n1569), .Z(n3613) );
  NAND U3571 ( .A(n3614), .B(n3613), .Z(n1571) );
  NAND U3572 ( .A(n1572), .B(n1571), .Z(n3615) );
  NAND U3573 ( .A(n3616), .B(n3615), .Z(n1573) );
  NAND U3574 ( .A(n1574), .B(n1573), .Z(n3617) );
  NAND U3575 ( .A(n3618), .B(n3617), .Z(n1575) );
  NAND U3576 ( .A(n1576), .B(n1575), .Z(n3619) );
  NAND U3577 ( .A(n3620), .B(n3619), .Z(n1577) );
  NAND U3578 ( .A(n1578), .B(n1577), .Z(n3621) );
  NAND U3579 ( .A(n3622), .B(n3621), .Z(n1579) );
  NAND U3580 ( .A(n1580), .B(n1579), .Z(n3625) );
  NAND U3581 ( .A(n3626), .B(n3625), .Z(n1581) );
  NAND U3582 ( .A(n1582), .B(n1581), .Z(n3627) );
  NAND U3583 ( .A(n3628), .B(n3627), .Z(n1583) );
  NAND U3584 ( .A(n1584), .B(n1583), .Z(n3629) );
  NAND U3585 ( .A(n3630), .B(n3629), .Z(n1585) );
  NAND U3586 ( .A(n1586), .B(n1585), .Z(n3631) );
  NAND U3587 ( .A(n3632), .B(n3631), .Z(n1587) );
  NAND U3588 ( .A(n1588), .B(n1587), .Z(n3633) );
  NAND U3589 ( .A(n3634), .B(n3633), .Z(n1589) );
  NAND U3590 ( .A(n1590), .B(n1589), .Z(n3635) );
  NAND U3591 ( .A(n3636), .B(n3635), .Z(n1591) );
  NAND U3592 ( .A(n1592), .B(n1591), .Z(n3637) );
  NAND U3593 ( .A(n3638), .B(n3637), .Z(n1593) );
  NAND U3594 ( .A(n1594), .B(n1593), .Z(n3639) );
  NAND U3595 ( .A(n3640), .B(n3639), .Z(n1595) );
  NAND U3596 ( .A(n1596), .B(n1595), .Z(n3641) );
  NAND U3597 ( .A(n3642), .B(n3641), .Z(n1597) );
  NAND U3598 ( .A(n1598), .B(n1597), .Z(n3643) );
  NAND U3599 ( .A(n3644), .B(n3643), .Z(n1599) );
  NAND U3600 ( .A(n1600), .B(n1599), .Z(n3649) );
  NAND U3601 ( .A(n3650), .B(n3649), .Z(n1601) );
  NAND U3602 ( .A(n1602), .B(n1601), .Z(n3651) );
  NAND U3603 ( .A(n3652), .B(n3651), .Z(n1603) );
  NAND U3604 ( .A(n1604), .B(n1603), .Z(n3653) );
  NAND U3605 ( .A(n3654), .B(n3653), .Z(n1605) );
  NAND U3606 ( .A(n1606), .B(n1605), .Z(n3655) );
  NAND U3607 ( .A(n3656), .B(n3655), .Z(n1607) );
  NAND U3608 ( .A(n1608), .B(n1607), .Z(n3657) );
  NAND U3609 ( .A(n3658), .B(n3657), .Z(n1609) );
  NAND U3610 ( .A(n1610), .B(n1609), .Z(n3659) );
  NAND U3611 ( .A(n3660), .B(n3659), .Z(n1611) );
  NAND U3612 ( .A(n1612), .B(n1611), .Z(n3661) );
  NAND U3613 ( .A(n3662), .B(n3661), .Z(n1613) );
  NAND U3614 ( .A(n1614), .B(n1613), .Z(n3663) );
  NAND U3615 ( .A(n3664), .B(n3663), .Z(n1615) );
  NAND U3616 ( .A(n1616), .B(n1615), .Z(n3665) );
  NAND U3617 ( .A(n3666), .B(n3665), .Z(n1617) );
  NAND U3618 ( .A(n1618), .B(n1617), .Z(n3667) );
  NAND U3619 ( .A(n3668), .B(n3667), .Z(n1619) );
  NAND U3620 ( .A(n1620), .B(n1619), .Z(n3671) );
  NAND U3621 ( .A(n3672), .B(n3671), .Z(n1621) );
  NAND U3622 ( .A(n1622), .B(n1621), .Z(n3673) );
  NAND U3623 ( .A(n3674), .B(n3673), .Z(n1623) );
  NAND U3624 ( .A(n1624), .B(n1623), .Z(n3675) );
  NAND U3625 ( .A(n3676), .B(n3675), .Z(n1625) );
  NAND U3626 ( .A(n1626), .B(n1625), .Z(n3677) );
  NAND U3627 ( .A(n3678), .B(n3677), .Z(n1627) );
  NAND U3628 ( .A(n1628), .B(n1627), .Z(n3679) );
  NAND U3629 ( .A(n3680), .B(n3679), .Z(n1629) );
  NAND U3630 ( .A(n1630), .B(n1629), .Z(n3681) );
  NAND U3631 ( .A(n3682), .B(n3681), .Z(n1631) );
  NAND U3632 ( .A(n1632), .B(n1631), .Z(n3683) );
  NAND U3633 ( .A(n3684), .B(n3683), .Z(n1633) );
  NAND U3634 ( .A(n1634), .B(n1633), .Z(n3685) );
  NAND U3635 ( .A(n3686), .B(n3685), .Z(n1635) );
  NAND U3636 ( .A(n1636), .B(n1635), .Z(n3687) );
  NAND U3637 ( .A(n3688), .B(n3687), .Z(n1637) );
  NAND U3638 ( .A(n1638), .B(n1637), .Z(n3689) );
  NAND U3639 ( .A(n3690), .B(n3689), .Z(n1639) );
  NAND U3640 ( .A(n1640), .B(n1639), .Z(n3693) );
  NAND U3641 ( .A(n3694), .B(n3693), .Z(n1641) );
  NAND U3642 ( .A(n1642), .B(n1641), .Z(n3695) );
  NAND U3643 ( .A(n3696), .B(n3695), .Z(n1643) );
  NAND U3644 ( .A(n1644), .B(n1643), .Z(n3697) );
  NAND U3645 ( .A(n3698), .B(n3697), .Z(n1645) );
  NAND U3646 ( .A(n1646), .B(n1645), .Z(n3699) );
  NAND U3647 ( .A(n3700), .B(n3699), .Z(n1647) );
  NAND U3648 ( .A(n1648), .B(n1647), .Z(n3701) );
  NAND U3649 ( .A(n3702), .B(n3701), .Z(n1649) );
  NAND U3650 ( .A(n1650), .B(n1649), .Z(n3703) );
  NAND U3651 ( .A(n3704), .B(n3703), .Z(n1651) );
  NAND U3652 ( .A(n1652), .B(n1651), .Z(n3705) );
  NAND U3653 ( .A(n3706), .B(n3705), .Z(n1653) );
  NAND U3654 ( .A(n1654), .B(n1653), .Z(n3707) );
  NAND U3655 ( .A(n3708), .B(n3707), .Z(n1655) );
  NAND U3656 ( .A(n1656), .B(n1655), .Z(n3709) );
  NAND U3657 ( .A(n3710), .B(n3709), .Z(n1657) );
  NAND U3658 ( .A(n1658), .B(n1657), .Z(n3711) );
  NAND U3659 ( .A(n3712), .B(n3711), .Z(n1659) );
  NAND U3660 ( .A(n1660), .B(n1659), .Z(n3715) );
  NAND U3661 ( .A(n3716), .B(n3715), .Z(n1661) );
  NAND U3662 ( .A(n1662), .B(n1661), .Z(n3717) );
  NAND U3663 ( .A(n3718), .B(n3717), .Z(n1663) );
  NAND U3664 ( .A(n1664), .B(n1663), .Z(n3719) );
  NAND U3665 ( .A(n3720), .B(n3719), .Z(n1665) );
  NAND U3666 ( .A(n1666), .B(n1665), .Z(n3721) );
  NAND U3667 ( .A(n3722), .B(n3721), .Z(n1667) );
  NAND U3668 ( .A(n1668), .B(n1667), .Z(n3723) );
  NAND U3669 ( .A(n3724), .B(n3723), .Z(n1669) );
  NAND U3670 ( .A(n1670), .B(n1669), .Z(n3725) );
  NAND U3671 ( .A(n3726), .B(n3725), .Z(n1671) );
  NAND U3672 ( .A(n1672), .B(n1671), .Z(n3727) );
  NAND U3673 ( .A(n3728), .B(n3727), .Z(n1673) );
  NAND U3674 ( .A(n1674), .B(n1673), .Z(n3729) );
  NAND U3675 ( .A(n3730), .B(n3729), .Z(n1675) );
  NAND U3676 ( .A(n1676), .B(n1675), .Z(n3731) );
  NAND U3677 ( .A(n3732), .B(n3731), .Z(n1677) );
  NAND U3678 ( .A(n1678), .B(n1677), .Z(n3733) );
  NAND U3679 ( .A(n3734), .B(n3733), .Z(n1679) );
  NAND U3680 ( .A(n1680), .B(n1679), .Z(n3737) );
  NAND U3681 ( .A(n3738), .B(n3737), .Z(n1681) );
  NAND U3682 ( .A(n1682), .B(n1681), .Z(n3739) );
  NAND U3683 ( .A(n3740), .B(n3739), .Z(n1683) );
  NAND U3684 ( .A(n1684), .B(n1683), .Z(n3741) );
  NAND U3685 ( .A(n3742), .B(n3741), .Z(n1685) );
  NAND U3686 ( .A(n1686), .B(n1685), .Z(n3743) );
  NAND U3687 ( .A(n3744), .B(n3743), .Z(n1687) );
  NAND U3688 ( .A(n1688), .B(n1687), .Z(n3745) );
  NAND U3689 ( .A(n3746), .B(n3745), .Z(n1689) );
  NAND U3690 ( .A(n1690), .B(n1689), .Z(n3747) );
  NAND U3691 ( .A(n3748), .B(n3747), .Z(n1691) );
  NAND U3692 ( .A(n1692), .B(n1691), .Z(n3749) );
  NAND U3693 ( .A(n3750), .B(n3749), .Z(n1693) );
  NAND U3694 ( .A(n1694), .B(n1693), .Z(n3751) );
  NAND U3695 ( .A(n3752), .B(n3751), .Z(n1695) );
  NAND U3696 ( .A(n1696), .B(n1695), .Z(n3753) );
  NAND U3697 ( .A(n3754), .B(n3753), .Z(n1697) );
  NAND U3698 ( .A(n1698), .B(n1697), .Z(n3755) );
  NAND U3699 ( .A(n3756), .B(n3755), .Z(n1699) );
  NAND U3700 ( .A(n1700), .B(n1699), .Z(n3759) );
  NAND U3701 ( .A(n3760), .B(n3759), .Z(n1701) );
  NAND U3702 ( .A(n1702), .B(n1701), .Z(n3761) );
  NAND U3703 ( .A(n3762), .B(n3761), .Z(n1703) );
  NAND U3704 ( .A(n1704), .B(n1703), .Z(n3763) );
  NAND U3705 ( .A(n3764), .B(n3763), .Z(n1705) );
  NAND U3706 ( .A(n1706), .B(n1705), .Z(n3765) );
  NAND U3707 ( .A(n3766), .B(n3765), .Z(n1707) );
  NAND U3708 ( .A(n1708), .B(n1707), .Z(n3767) );
  NAND U3709 ( .A(n3768), .B(n3767), .Z(n1709) );
  NAND U3710 ( .A(n1710), .B(n1709), .Z(n3769) );
  NAND U3711 ( .A(n3770), .B(n3769), .Z(n1711) );
  NAND U3712 ( .A(n1712), .B(n1711), .Z(n3771) );
  NAND U3713 ( .A(n3772), .B(n3771), .Z(n1713) );
  NAND U3714 ( .A(n1714), .B(n1713), .Z(n3773) );
  NAND U3715 ( .A(n3774), .B(n3773), .Z(n1715) );
  NAND U3716 ( .A(n1716), .B(n1715), .Z(n3775) );
  NAND U3717 ( .A(n3776), .B(n3775), .Z(n1717) );
  NAND U3718 ( .A(n1718), .B(n1717), .Z(n3777) );
  NAND U3719 ( .A(n3778), .B(n3777), .Z(n1719) );
  NAND U3720 ( .A(n1720), .B(n1719), .Z(n3781) );
  NAND U3721 ( .A(n3782), .B(n3781), .Z(n1721) );
  NAND U3722 ( .A(n1722), .B(n1721), .Z(n3783) );
  NAND U3723 ( .A(n3784), .B(n3783), .Z(n1723) );
  NAND U3724 ( .A(n1724), .B(n1723), .Z(n3785) );
  NAND U3725 ( .A(n3786), .B(n3785), .Z(n1725) );
  NAND U3726 ( .A(n1726), .B(n1725), .Z(n3787) );
  NAND U3727 ( .A(n3788), .B(n3787), .Z(n1727) );
  NAND U3728 ( .A(n1728), .B(n1727), .Z(n3789) );
  NAND U3729 ( .A(n3790), .B(n3789), .Z(n1729) );
  NAND U3730 ( .A(n1730), .B(n1729), .Z(n3791) );
  NAND U3731 ( .A(n3792), .B(n3791), .Z(n1731) );
  NAND U3732 ( .A(n1732), .B(n1731), .Z(n3793) );
  NAND U3733 ( .A(n3794), .B(n3793), .Z(n1733) );
  NAND U3734 ( .A(n1734), .B(n1733), .Z(n3795) );
  NAND U3735 ( .A(n3796), .B(n3795), .Z(n1735) );
  NAND U3736 ( .A(n1736), .B(n1735), .Z(n3797) );
  NAND U3737 ( .A(n3798), .B(n3797), .Z(n1737) );
  NAND U3738 ( .A(n1738), .B(n1737), .Z(n3799) );
  NAND U3739 ( .A(n3800), .B(n3799), .Z(n1739) );
  NAND U3740 ( .A(n1740), .B(n1739), .Z(n3803) );
  NAND U3741 ( .A(n3804), .B(n3803), .Z(n1741) );
  NAND U3742 ( .A(n1742), .B(n1741), .Z(n3805) );
  NAND U3743 ( .A(n3806), .B(n3805), .Z(n1743) );
  NAND U3744 ( .A(n1744), .B(n1743), .Z(n3807) );
  NAND U3745 ( .A(n3808), .B(n3807), .Z(n1745) );
  NAND U3746 ( .A(n1746), .B(n1745), .Z(n3809) );
  NAND U3747 ( .A(n3810), .B(n3809), .Z(n1747) );
  NAND U3748 ( .A(n1748), .B(n1747), .Z(n3811) );
  NAND U3749 ( .A(n3812), .B(n3811), .Z(n1749) );
  NAND U3750 ( .A(n1750), .B(n1749), .Z(n3813) );
  NAND U3751 ( .A(n3814), .B(n3813), .Z(n1751) );
  NAND U3752 ( .A(n1752), .B(n1751), .Z(n3815) );
  NAND U3753 ( .A(n3816), .B(n3815), .Z(n1753) );
  NAND U3754 ( .A(n1754), .B(n1753), .Z(n3817) );
  NAND U3755 ( .A(n3818), .B(n3817), .Z(n1755) );
  NAND U3756 ( .A(n1756), .B(n1755), .Z(n3819) );
  NAND U3757 ( .A(n3820), .B(n3819), .Z(n1757) );
  NAND U3758 ( .A(n1758), .B(n1757), .Z(n3821) );
  NAND U3759 ( .A(n3822), .B(n3821), .Z(n1759) );
  NAND U3760 ( .A(n1760), .B(n1759), .Z(n3825) );
  NAND U3761 ( .A(n3826), .B(n3825), .Z(n1761) );
  NAND U3762 ( .A(n1762), .B(n1761), .Z(n3827) );
  NAND U3763 ( .A(n3828), .B(n3827), .Z(n1763) );
  NAND U3764 ( .A(n1764), .B(n1763), .Z(n3829) );
  NAND U3765 ( .A(n3830), .B(n3829), .Z(n1765) );
  NAND U3766 ( .A(n1766), .B(n1765), .Z(n3831) );
  NAND U3767 ( .A(n3832), .B(n3831), .Z(n1767) );
  NAND U3768 ( .A(n1768), .B(n1767), .Z(n3833) );
  NAND U3769 ( .A(n3834), .B(n3833), .Z(n1769) );
  NAND U3770 ( .A(n1770), .B(n1769), .Z(n3835) );
  NAND U3771 ( .A(n3836), .B(n3835), .Z(n1771) );
  NAND U3772 ( .A(n1772), .B(n1771), .Z(n3837) );
  NAND U3773 ( .A(n3838), .B(n3837), .Z(n1773) );
  NAND U3774 ( .A(n1774), .B(n1773), .Z(n3839) );
  NAND U3775 ( .A(n3840), .B(n3839), .Z(n1775) );
  NAND U3776 ( .A(n1776), .B(n1775), .Z(n3841) );
  NAND U3777 ( .A(n3842), .B(n3841), .Z(n1777) );
  NAND U3778 ( .A(n1778), .B(n1777), .Z(n3843) );
  NAND U3779 ( .A(n3844), .B(n3843), .Z(n1779) );
  NAND U3780 ( .A(n1780), .B(n1779), .Z(n3847) );
  NAND U3781 ( .A(n3848), .B(n3847), .Z(n1781) );
  NAND U3782 ( .A(n1782), .B(n1781), .Z(n3849) );
  NAND U3783 ( .A(n3850), .B(n3849), .Z(n1783) );
  NAND U3784 ( .A(n1784), .B(n1783), .Z(n3851) );
  NAND U3785 ( .A(n3852), .B(n3851), .Z(n1785) );
  NAND U3786 ( .A(n1786), .B(n1785), .Z(n3853) );
  NAND U3787 ( .A(n3854), .B(n3853), .Z(n1787) );
  NAND U3788 ( .A(n1788), .B(n1787), .Z(n3855) );
  NAND U3789 ( .A(n3856), .B(n3855), .Z(n1789) );
  NAND U3790 ( .A(n1790), .B(n1789), .Z(n3857) );
  NAND U3791 ( .A(n3858), .B(n3857), .Z(n1791) );
  NAND U3792 ( .A(n1792), .B(n1791), .Z(n3859) );
  NAND U3793 ( .A(n3860), .B(n3859), .Z(n1793) );
  NAND U3794 ( .A(n1794), .B(n1793), .Z(n3861) );
  NAND U3795 ( .A(n3862), .B(n3861), .Z(n1795) );
  NAND U3796 ( .A(n1796), .B(n1795), .Z(n3863) );
  NAND U3797 ( .A(n3864), .B(n3863), .Z(n1797) );
  NAND U3798 ( .A(n1798), .B(n1797), .Z(n3865) );
  NAND U3799 ( .A(n3866), .B(n3865), .Z(n1799) );
  NAND U3800 ( .A(n1800), .B(n1799), .Z(n3871) );
  NAND U3801 ( .A(n3872), .B(n3871), .Z(n1801) );
  NAND U3802 ( .A(n1802), .B(n1801), .Z(n3873) );
  NAND U3803 ( .A(n3874), .B(n3873), .Z(n1803) );
  NAND U3804 ( .A(n1804), .B(n1803), .Z(n3875) );
  NAND U3805 ( .A(n3876), .B(n3875), .Z(n1805) );
  NAND U3806 ( .A(n1806), .B(n1805), .Z(n3877) );
  NAND U3807 ( .A(n3878), .B(n3877), .Z(n1807) );
  NAND U3808 ( .A(n1808), .B(n1807), .Z(n3879) );
  NAND U3809 ( .A(n3880), .B(n3879), .Z(n1809) );
  NAND U3810 ( .A(n1810), .B(n1809), .Z(n3881) );
  NAND U3811 ( .A(n3882), .B(n3881), .Z(n1811) );
  NAND U3812 ( .A(n1812), .B(n1811), .Z(n3883) );
  NAND U3813 ( .A(n3884), .B(n3883), .Z(n1813) );
  NAND U3814 ( .A(n1814), .B(n1813), .Z(n3885) );
  NAND U3815 ( .A(n3886), .B(n3885), .Z(n1815) );
  NAND U3816 ( .A(n1816), .B(n1815), .Z(n3887) );
  NAND U3817 ( .A(n3888), .B(n3887), .Z(n1817) );
  NAND U3818 ( .A(n1818), .B(n1817), .Z(n3889) );
  NAND U3819 ( .A(n3890), .B(n3889), .Z(n1819) );
  NAND U3820 ( .A(n1820), .B(n1819), .Z(n3893) );
  NAND U3821 ( .A(n3894), .B(n3893), .Z(n1821) );
  NAND U3822 ( .A(n1822), .B(n1821), .Z(n3895) );
  NAND U3823 ( .A(n3896), .B(n3895), .Z(n1823) );
  NAND U3824 ( .A(n1824), .B(n1823), .Z(n3897) );
  NAND U3825 ( .A(n3898), .B(n3897), .Z(n1825) );
  NAND U3826 ( .A(n1826), .B(n1825), .Z(n3899) );
  NAND U3827 ( .A(n3900), .B(n3899), .Z(n1827) );
  NAND U3828 ( .A(n1828), .B(n1827), .Z(n3901) );
  NAND U3829 ( .A(n3902), .B(n3901), .Z(n1829) );
  NAND U3830 ( .A(n1830), .B(n1829), .Z(n3903) );
  NAND U3831 ( .A(n3904), .B(n3903), .Z(n1831) );
  NAND U3832 ( .A(n1832), .B(n1831), .Z(n3905) );
  NAND U3833 ( .A(n3906), .B(n3905), .Z(n1833) );
  NAND U3834 ( .A(n1834), .B(n1833), .Z(n3907) );
  NAND U3835 ( .A(n3908), .B(n3907), .Z(n1835) );
  NAND U3836 ( .A(n1836), .B(n1835), .Z(n3909) );
  NAND U3837 ( .A(n3910), .B(n3909), .Z(n1837) );
  NAND U3838 ( .A(n1838), .B(n1837), .Z(n3911) );
  NAND U3839 ( .A(n3912), .B(n3911), .Z(n1839) );
  NAND U3840 ( .A(n1840), .B(n1839), .Z(n3915) );
  NAND U3841 ( .A(n3916), .B(n3915), .Z(n1841) );
  NAND U3842 ( .A(n1842), .B(n1841), .Z(n3917) );
  NAND U3843 ( .A(n3918), .B(n3917), .Z(n1843) );
  NAND U3844 ( .A(n1844), .B(n1843), .Z(n3919) );
  NAND U3845 ( .A(n3920), .B(n3919), .Z(n1845) );
  NAND U3846 ( .A(n1846), .B(n1845), .Z(n3921) );
  NAND U3847 ( .A(n3922), .B(n3921), .Z(n1847) );
  NAND U3848 ( .A(n1848), .B(n1847), .Z(n3923) );
  NAND U3849 ( .A(n3924), .B(n3923), .Z(n1849) );
  NAND U3850 ( .A(n1850), .B(n1849), .Z(n3925) );
  NAND U3851 ( .A(n3926), .B(n3925), .Z(n1851) );
  NAND U3852 ( .A(n1852), .B(n1851), .Z(n3927) );
  NAND U3853 ( .A(n3928), .B(n3927), .Z(n1853) );
  NAND U3854 ( .A(n1854), .B(n1853), .Z(n3929) );
  NAND U3855 ( .A(n3930), .B(n3929), .Z(n1855) );
  NAND U3856 ( .A(n1856), .B(n1855), .Z(n3931) );
  NAND U3857 ( .A(n3932), .B(n3931), .Z(n1857) );
  NAND U3858 ( .A(n1858), .B(n1857), .Z(n3933) );
  NAND U3859 ( .A(n3934), .B(n3933), .Z(n1859) );
  NAND U3860 ( .A(n1860), .B(n1859), .Z(n3937) );
  NAND U3861 ( .A(n3938), .B(n3937), .Z(n1861) );
  NAND U3862 ( .A(n1862), .B(n1861), .Z(n3939) );
  NAND U3863 ( .A(n3940), .B(n3939), .Z(n1863) );
  NAND U3864 ( .A(n1864), .B(n1863), .Z(n3941) );
  NAND U3865 ( .A(n3942), .B(n3941), .Z(n1865) );
  NAND U3866 ( .A(n1866), .B(n1865), .Z(n3943) );
  NAND U3867 ( .A(n3944), .B(n3943), .Z(n1867) );
  NAND U3868 ( .A(n1868), .B(n1867), .Z(n3945) );
  NAND U3869 ( .A(n3946), .B(n3945), .Z(n1869) );
  NAND U3870 ( .A(n1870), .B(n1869), .Z(n3947) );
  NAND U3871 ( .A(n3948), .B(n3947), .Z(n1871) );
  NAND U3872 ( .A(n1872), .B(n1871), .Z(n3949) );
  NAND U3873 ( .A(n3950), .B(n3949), .Z(n1873) );
  NAND U3874 ( .A(n1874), .B(n1873), .Z(n3951) );
  NAND U3875 ( .A(n3952), .B(n3951), .Z(n1875) );
  NAND U3876 ( .A(n1876), .B(n1875), .Z(n3953) );
  NAND U3877 ( .A(n3954), .B(n3953), .Z(n1877) );
  NAND U3878 ( .A(n1878), .B(n1877), .Z(n3955) );
  NAND U3879 ( .A(n3956), .B(n3955), .Z(n1879) );
  NAND U3880 ( .A(n1880), .B(n1879), .Z(n3959) );
  NAND U3881 ( .A(n3960), .B(n3959), .Z(n1881) );
  NAND U3882 ( .A(n1882), .B(n1881), .Z(n3961) );
  NAND U3883 ( .A(n3962), .B(n3961), .Z(n1883) );
  NAND U3884 ( .A(n1884), .B(n1883), .Z(n3963) );
  NAND U3885 ( .A(n3964), .B(n3963), .Z(n1885) );
  NAND U3886 ( .A(n1886), .B(n1885), .Z(n3965) );
  NAND U3887 ( .A(n3966), .B(n3965), .Z(n1887) );
  NAND U3888 ( .A(n1888), .B(n1887), .Z(n3967) );
  NAND U3889 ( .A(n3968), .B(n3967), .Z(n1889) );
  NAND U3890 ( .A(n1890), .B(n1889), .Z(n3969) );
  NAND U3891 ( .A(n3970), .B(n3969), .Z(n1891) );
  NAND U3892 ( .A(n1892), .B(n1891), .Z(n3971) );
  NAND U3893 ( .A(n3972), .B(n3971), .Z(n1893) );
  NAND U3894 ( .A(n1894), .B(n1893), .Z(n3973) );
  NAND U3895 ( .A(n3974), .B(n3973), .Z(n1895) );
  NAND U3896 ( .A(n1896), .B(n1895), .Z(n3975) );
  NAND U3897 ( .A(n3976), .B(n3975), .Z(n1897) );
  NAND U3898 ( .A(n1898), .B(n1897), .Z(n3977) );
  NAND U3899 ( .A(n3978), .B(n3977), .Z(n1899) );
  NAND U3900 ( .A(n1900), .B(n1899), .Z(n3981) );
  NAND U3901 ( .A(n3982), .B(n3981), .Z(n1901) );
  NAND U3902 ( .A(n1902), .B(n1901), .Z(n3983) );
  NAND U3903 ( .A(n3984), .B(n3983), .Z(n1903) );
  NAND U3904 ( .A(n1904), .B(n1903), .Z(n3985) );
  NAND U3905 ( .A(n3986), .B(n3985), .Z(n1905) );
  NAND U3906 ( .A(n1906), .B(n1905), .Z(n3987) );
  NAND U3907 ( .A(n3988), .B(n3987), .Z(n1907) );
  NAND U3908 ( .A(n1908), .B(n1907), .Z(n3989) );
  NAND U3909 ( .A(n3990), .B(n3989), .Z(n1909) );
  NAND U3910 ( .A(n1910), .B(n1909), .Z(n3991) );
  NAND U3911 ( .A(n3992), .B(n3991), .Z(n1911) );
  NAND U3912 ( .A(n1912), .B(n1911), .Z(n3993) );
  NAND U3913 ( .A(n3994), .B(n3993), .Z(n1913) );
  NAND U3914 ( .A(n1914), .B(n1913), .Z(n3995) );
  NAND U3915 ( .A(n3996), .B(n3995), .Z(n1915) );
  NAND U3916 ( .A(n1916), .B(n1915), .Z(n3997) );
  NAND U3917 ( .A(n3998), .B(n3997), .Z(n1917) );
  NAND U3918 ( .A(n1918), .B(n1917), .Z(n3999) );
  NAND U3919 ( .A(n4000), .B(n3999), .Z(n1919) );
  NAND U3920 ( .A(n1920), .B(n1919), .Z(n4003) );
  NAND U3921 ( .A(n4004), .B(n4003), .Z(n1921) );
  NAND U3922 ( .A(n1922), .B(n1921), .Z(n4005) );
  NAND U3923 ( .A(n4006), .B(n4005), .Z(n1923) );
  NAND U3924 ( .A(n1924), .B(n1923), .Z(n4007) );
  NAND U3925 ( .A(n4008), .B(n4007), .Z(n1925) );
  NAND U3926 ( .A(n1926), .B(n1925), .Z(n4009) );
  NAND U3927 ( .A(n4010), .B(n4009), .Z(n1927) );
  NAND U3928 ( .A(n1928), .B(n1927), .Z(n4011) );
  NAND U3929 ( .A(n4012), .B(n4011), .Z(n1929) );
  NAND U3930 ( .A(n1930), .B(n1929), .Z(n4013) );
  NAND U3931 ( .A(n4014), .B(n4013), .Z(n1931) );
  NAND U3932 ( .A(n1932), .B(n1931), .Z(n4015) );
  NAND U3933 ( .A(n4016), .B(n4015), .Z(n1933) );
  NAND U3934 ( .A(n1934), .B(n1933), .Z(n4017) );
  NAND U3935 ( .A(n4018), .B(n4017), .Z(n1935) );
  NAND U3936 ( .A(n1936), .B(n1935), .Z(n4019) );
  NAND U3937 ( .A(n4020), .B(n4019), .Z(n1937) );
  NAND U3938 ( .A(n1938), .B(n1937), .Z(n4021) );
  NAND U3939 ( .A(n4022), .B(n4021), .Z(n1939) );
  NAND U3940 ( .A(n1940), .B(n1939), .Z(n4025) );
  NAND U3941 ( .A(n4026), .B(n4025), .Z(n1941) );
  NAND U3942 ( .A(n1942), .B(n1941), .Z(n4027) );
  NAND U3943 ( .A(n4028), .B(n4027), .Z(n1943) );
  NAND U3944 ( .A(n1944), .B(n1943), .Z(n4029) );
  NAND U3945 ( .A(n4030), .B(n4029), .Z(n1945) );
  NAND U3946 ( .A(n1946), .B(n1945), .Z(n4031) );
  NAND U3947 ( .A(n4032), .B(n4031), .Z(n1947) );
  NAND U3948 ( .A(n1948), .B(n1947), .Z(n4033) );
  NAND U3949 ( .A(n4034), .B(n4033), .Z(n1949) );
  NAND U3950 ( .A(n1950), .B(n1949), .Z(n4035) );
  NAND U3951 ( .A(n4036), .B(n4035), .Z(n1951) );
  NAND U3952 ( .A(n1952), .B(n1951), .Z(n4037) );
  NAND U3953 ( .A(n4038), .B(n4037), .Z(n1953) );
  NAND U3954 ( .A(n1954), .B(n1953), .Z(n4039) );
  NAND U3955 ( .A(n4040), .B(n4039), .Z(n1955) );
  NAND U3956 ( .A(n1956), .B(n1955), .Z(n4041) );
  NAND U3957 ( .A(n4042), .B(n4041), .Z(n1957) );
  NAND U3958 ( .A(n1958), .B(n1957), .Z(n4043) );
  NAND U3959 ( .A(n4044), .B(n4043), .Z(n1959) );
  NAND U3960 ( .A(n1960), .B(n1959), .Z(n4047) );
  NAND U3961 ( .A(n4048), .B(n4047), .Z(n1961) );
  NAND U3962 ( .A(n1962), .B(n1961), .Z(n4049) );
  NAND U3963 ( .A(n4050), .B(n4049), .Z(n1963) );
  NAND U3964 ( .A(n1964), .B(n1963), .Z(n4051) );
  NAND U3965 ( .A(n4052), .B(n4051), .Z(n1965) );
  NAND U3966 ( .A(n1966), .B(n1965), .Z(n4053) );
  NAND U3967 ( .A(n4054), .B(n4053), .Z(n1967) );
  NAND U3968 ( .A(n1968), .B(n1967), .Z(n4055) );
  NAND U3969 ( .A(n4056), .B(n4055), .Z(n1969) );
  NAND U3970 ( .A(n1970), .B(n1969), .Z(n4057) );
  NAND U3971 ( .A(n4058), .B(n4057), .Z(n1971) );
  NAND U3972 ( .A(n1972), .B(n1971), .Z(n4059) );
  NAND U3973 ( .A(n4060), .B(n4059), .Z(n1973) );
  NAND U3974 ( .A(n1974), .B(n1973), .Z(n4061) );
  NAND U3975 ( .A(n4062), .B(n4061), .Z(n1975) );
  NAND U3976 ( .A(n1976), .B(n1975), .Z(n4063) );
  NAND U3977 ( .A(n4064), .B(n4063), .Z(n1977) );
  NAND U3978 ( .A(n1978), .B(n1977), .Z(n4065) );
  NAND U3979 ( .A(n4066), .B(n4065), .Z(n1979) );
  NAND U3980 ( .A(n1980), .B(n1979), .Z(n4069) );
  NAND U3981 ( .A(n4070), .B(n4069), .Z(n1981) );
  NAND U3982 ( .A(n1982), .B(n1981), .Z(n4071) );
  NAND U3983 ( .A(n4072), .B(n4071), .Z(n1983) );
  NAND U3984 ( .A(n1984), .B(n1983), .Z(n4073) );
  NAND U3985 ( .A(n4074), .B(n4073), .Z(n1985) );
  NAND U3986 ( .A(n1986), .B(n1985), .Z(n4075) );
  NAND U3987 ( .A(n4076), .B(n4075), .Z(n1987) );
  NAND U3988 ( .A(n1988), .B(n1987), .Z(n4077) );
  NAND U3989 ( .A(n4078), .B(n4077), .Z(n1989) );
  NAND U3990 ( .A(n1990), .B(n1989), .Z(n4079) );
  NAND U3991 ( .A(n4080), .B(n4079), .Z(n1991) );
  NAND U3992 ( .A(n1992), .B(n1991), .Z(n4081) );
  NAND U3993 ( .A(n4082), .B(n4081), .Z(n1993) );
  NAND U3994 ( .A(n1994), .B(n1993), .Z(n4083) );
  NAND U3995 ( .A(n4084), .B(n4083), .Z(n1995) );
  NAND U3996 ( .A(n1996), .B(n1995), .Z(n4085) );
  NAND U3997 ( .A(n4086), .B(n4085), .Z(n1997) );
  NAND U3998 ( .A(n1998), .B(n1997), .Z(n4087) );
  NAND U3999 ( .A(n4088), .B(n4087), .Z(n1999) );
  NAND U4000 ( .A(n2000), .B(n1999), .Z(n2001) );
  XNOR U4001 ( .A(n2002), .B(n2001), .Z(c[1000]) );
  XOR U4002 ( .A(b[1001]), .B(a[1001]), .Z(n2006) );
  OR U4003 ( .A(b[1000]), .B(a[1000]), .Z(n2004) );
  NAND U4004 ( .A(n2002), .B(n2001), .Z(n2003) );
  NAND U4005 ( .A(n2004), .B(n2003), .Z(n2005) );
  XNOR U4006 ( .A(n2006), .B(n2005), .Z(c[1001]) );
  XOR U4007 ( .A(b[1002]), .B(a[1002]), .Z(n2010) );
  OR U4008 ( .A(b[1001]), .B(a[1001]), .Z(n2008) );
  NAND U4009 ( .A(n2006), .B(n2005), .Z(n2007) );
  NAND U4010 ( .A(n2008), .B(n2007), .Z(n2009) );
  XNOR U4011 ( .A(n2010), .B(n2009), .Z(c[1002]) );
  XOR U4012 ( .A(b[1003]), .B(a[1003]), .Z(n2014) );
  OR U4013 ( .A(b[1002]), .B(a[1002]), .Z(n2012) );
  NAND U4014 ( .A(n2010), .B(n2009), .Z(n2011) );
  NAND U4015 ( .A(n2012), .B(n2011), .Z(n2013) );
  XNOR U4016 ( .A(n2014), .B(n2013), .Z(c[1003]) );
  XOR U4017 ( .A(b[1004]), .B(a[1004]), .Z(n2018) );
  OR U4018 ( .A(b[1003]), .B(a[1003]), .Z(n2016) );
  NAND U4019 ( .A(n2014), .B(n2013), .Z(n2015) );
  NAND U4020 ( .A(n2016), .B(n2015), .Z(n2017) );
  XNOR U4021 ( .A(n2018), .B(n2017), .Z(c[1004]) );
  XOR U4022 ( .A(b[1005]), .B(a[1005]), .Z(n2022) );
  OR U4023 ( .A(b[1004]), .B(a[1004]), .Z(n2020) );
  NAND U4024 ( .A(n2018), .B(n2017), .Z(n2019) );
  NAND U4025 ( .A(n2020), .B(n2019), .Z(n2021) );
  XNOR U4026 ( .A(n2022), .B(n2021), .Z(c[1005]) );
  XOR U4027 ( .A(b[1006]), .B(a[1006]), .Z(n2026) );
  OR U4028 ( .A(b[1005]), .B(a[1005]), .Z(n2024) );
  NAND U4029 ( .A(n2022), .B(n2021), .Z(n2023) );
  NAND U4030 ( .A(n2024), .B(n2023), .Z(n2025) );
  XNOR U4031 ( .A(n2026), .B(n2025), .Z(c[1006]) );
  XOR U4032 ( .A(b[1007]), .B(a[1007]), .Z(n2030) );
  OR U4033 ( .A(b[1006]), .B(a[1006]), .Z(n2028) );
  NAND U4034 ( .A(n2026), .B(n2025), .Z(n2027) );
  NAND U4035 ( .A(n2028), .B(n2027), .Z(n2029) );
  XNOR U4036 ( .A(n2030), .B(n2029), .Z(c[1007]) );
  XOR U4037 ( .A(b[1008]), .B(a[1008]), .Z(n2034) );
  OR U4038 ( .A(b[1007]), .B(a[1007]), .Z(n2032) );
  NAND U4039 ( .A(n2030), .B(n2029), .Z(n2031) );
  NAND U4040 ( .A(n2032), .B(n2031), .Z(n2033) );
  XNOR U4041 ( .A(n2034), .B(n2033), .Z(c[1008]) );
  XOR U4042 ( .A(b[1009]), .B(a[1009]), .Z(n2040) );
  OR U4043 ( .A(b[1008]), .B(a[1008]), .Z(n2036) );
  NAND U4044 ( .A(n2034), .B(n2033), .Z(n2035) );
  NAND U4045 ( .A(n2036), .B(n2035), .Z(n2039) );
  XNOR U4046 ( .A(n2040), .B(n2039), .Z(c[1009]) );
  XNOR U4047 ( .A(n2038), .B(n2037), .Z(c[100]) );
  XOR U4048 ( .A(b[1010]), .B(a[1010]), .Z(n2044) );
  OR U4049 ( .A(b[1009]), .B(a[1009]), .Z(n2042) );
  NAND U4050 ( .A(n2040), .B(n2039), .Z(n2041) );
  NAND U4051 ( .A(n2042), .B(n2041), .Z(n2043) );
  XNOR U4052 ( .A(n2044), .B(n2043), .Z(c[1010]) );
  XOR U4053 ( .A(b[1011]), .B(a[1011]), .Z(n2048) );
  OR U4054 ( .A(b[1010]), .B(a[1010]), .Z(n2046) );
  NAND U4055 ( .A(n2044), .B(n2043), .Z(n2045) );
  NAND U4056 ( .A(n2046), .B(n2045), .Z(n2047) );
  XNOR U4057 ( .A(n2048), .B(n2047), .Z(c[1011]) );
  XOR U4058 ( .A(b[1012]), .B(a[1012]), .Z(n2052) );
  OR U4059 ( .A(b[1011]), .B(a[1011]), .Z(n2050) );
  NAND U4060 ( .A(n2048), .B(n2047), .Z(n2049) );
  NAND U4061 ( .A(n2050), .B(n2049), .Z(n2051) );
  XNOR U4062 ( .A(n2052), .B(n2051), .Z(c[1012]) );
  XOR U4063 ( .A(b[1013]), .B(a[1013]), .Z(n2056) );
  OR U4064 ( .A(b[1012]), .B(a[1012]), .Z(n2054) );
  NAND U4065 ( .A(n2052), .B(n2051), .Z(n2053) );
  NAND U4066 ( .A(n2054), .B(n2053), .Z(n2055) );
  XNOR U4067 ( .A(n2056), .B(n2055), .Z(c[1013]) );
  XOR U4068 ( .A(b[1014]), .B(a[1014]), .Z(n2060) );
  OR U4069 ( .A(b[1013]), .B(a[1013]), .Z(n2058) );
  NAND U4070 ( .A(n2056), .B(n2055), .Z(n2057) );
  NAND U4071 ( .A(n2058), .B(n2057), .Z(n2059) );
  XNOR U4072 ( .A(n2060), .B(n2059), .Z(c[1014]) );
  XOR U4073 ( .A(b[1015]), .B(a[1015]), .Z(n2064) );
  OR U4074 ( .A(b[1014]), .B(a[1014]), .Z(n2062) );
  NAND U4075 ( .A(n2060), .B(n2059), .Z(n2061) );
  NAND U4076 ( .A(n2062), .B(n2061), .Z(n2063) );
  XNOR U4077 ( .A(n2064), .B(n2063), .Z(c[1015]) );
  XOR U4078 ( .A(b[1016]), .B(a[1016]), .Z(n2068) );
  OR U4079 ( .A(b[1015]), .B(a[1015]), .Z(n2066) );
  NAND U4080 ( .A(n2064), .B(n2063), .Z(n2065) );
  NAND U4081 ( .A(n2066), .B(n2065), .Z(n2067) );
  XNOR U4082 ( .A(n2068), .B(n2067), .Z(c[1016]) );
  XOR U4083 ( .A(b[1017]), .B(a[1017]), .Z(n2072) );
  OR U4084 ( .A(b[1016]), .B(a[1016]), .Z(n2070) );
  NAND U4085 ( .A(n2068), .B(n2067), .Z(n2069) );
  NAND U4086 ( .A(n2070), .B(n2069), .Z(n2071) );
  XNOR U4087 ( .A(n2072), .B(n2071), .Z(c[1017]) );
  XOR U4088 ( .A(b[1018]), .B(a[1018]), .Z(n2076) );
  OR U4089 ( .A(b[1017]), .B(a[1017]), .Z(n2074) );
  NAND U4090 ( .A(n2072), .B(n2071), .Z(n2073) );
  NAND U4091 ( .A(n2074), .B(n2073), .Z(n2075) );
  XNOR U4092 ( .A(n2076), .B(n2075), .Z(c[1018]) );
  XOR U4093 ( .A(b[1019]), .B(a[1019]), .Z(n2082) );
  OR U4094 ( .A(b[1018]), .B(a[1018]), .Z(n2078) );
  NAND U4095 ( .A(n2076), .B(n2075), .Z(n2077) );
  NAND U4096 ( .A(n2078), .B(n2077), .Z(n2081) );
  XNOR U4097 ( .A(n2082), .B(n2081), .Z(c[1019]) );
  XNOR U4098 ( .A(n2080), .B(n2079), .Z(c[101]) );
  XOR U4099 ( .A(b[1020]), .B(a[1020]), .Z(n2086) );
  OR U4100 ( .A(b[1019]), .B(a[1019]), .Z(n2084) );
  NAND U4101 ( .A(n2082), .B(n2081), .Z(n2083) );
  NAND U4102 ( .A(n2084), .B(n2083), .Z(n2085) );
  XNOR U4103 ( .A(n2086), .B(n2085), .Z(c[1020]) );
  XOR U4104 ( .A(b[1021]), .B(a[1021]), .Z(n2090) );
  OR U4105 ( .A(b[1020]), .B(a[1020]), .Z(n2088) );
  NAND U4106 ( .A(n2086), .B(n2085), .Z(n2087) );
  NAND U4107 ( .A(n2088), .B(n2087), .Z(n2089) );
  XNOR U4108 ( .A(n2090), .B(n2089), .Z(c[1021]) );
  XOR U4109 ( .A(b[1022]), .B(a[1022]), .Z(n2094) );
  OR U4110 ( .A(b[1021]), .B(a[1021]), .Z(n2092) );
  NAND U4111 ( .A(n2090), .B(n2089), .Z(n2091) );
  NAND U4112 ( .A(n2092), .B(n2091), .Z(n2093) );
  XNOR U4113 ( .A(n2094), .B(n2093), .Z(c[1022]) );
  NAND U4114 ( .A(n2094), .B(n2093), .Z(n2096) );
  OR U4115 ( .A(b[1022]), .B(a[1022]), .Z(n2095) );
  AND U4116 ( .A(n2096), .B(n2095), .Z(n2098) );
  XNOR U4117 ( .A(b[1023]), .B(a[1023]), .Z(n2097) );
  XNOR U4118 ( .A(n2098), .B(n2097), .Z(c[1023]) );
  XNOR U4119 ( .A(n2100), .B(n2099), .Z(c[102]) );
  XNOR U4120 ( .A(n2102), .B(n2101), .Z(c[103]) );
  XNOR U4121 ( .A(n2104), .B(n2103), .Z(c[104]) );
  XNOR U4122 ( .A(n2106), .B(n2105), .Z(c[105]) );
  XNOR U4123 ( .A(n2108), .B(n2107), .Z(c[106]) );
  XNOR U4124 ( .A(n2110), .B(n2109), .Z(c[107]) );
  XNOR U4125 ( .A(n2112), .B(n2111), .Z(c[108]) );
  XNOR U4126 ( .A(n2114), .B(n2113), .Z(c[109]) );
  XNOR U4127 ( .A(n2116), .B(n2115), .Z(c[10]) );
  XNOR U4128 ( .A(n2118), .B(n2117), .Z(c[110]) );
  XNOR U4129 ( .A(n2120), .B(n2119), .Z(c[111]) );
  XNOR U4130 ( .A(n2122), .B(n2121), .Z(c[112]) );
  XNOR U4131 ( .A(n2124), .B(n2123), .Z(c[113]) );
  XNOR U4132 ( .A(n2126), .B(n2125), .Z(c[114]) );
  XNOR U4133 ( .A(n2128), .B(n2127), .Z(c[115]) );
  XNOR U4134 ( .A(n2130), .B(n2129), .Z(c[116]) );
  XNOR U4135 ( .A(n2132), .B(n2131), .Z(c[117]) );
  XNOR U4136 ( .A(n2134), .B(n2133), .Z(c[118]) );
  XNOR U4137 ( .A(n2136), .B(n2135), .Z(c[119]) );
  XNOR U4138 ( .A(n2138), .B(n2137), .Z(c[11]) );
  XNOR U4139 ( .A(n2140), .B(n2139), .Z(c[120]) );
  XNOR U4140 ( .A(n2142), .B(n2141), .Z(c[121]) );
  XNOR U4141 ( .A(n2144), .B(n2143), .Z(c[122]) );
  XNOR U4142 ( .A(n2146), .B(n2145), .Z(c[123]) );
  XNOR U4143 ( .A(n2148), .B(n2147), .Z(c[124]) );
  XNOR U4144 ( .A(n2150), .B(n2149), .Z(c[125]) );
  XNOR U4145 ( .A(n2152), .B(n2151), .Z(c[126]) );
  XNOR U4146 ( .A(n2154), .B(n2153), .Z(c[127]) );
  XNOR U4147 ( .A(n2156), .B(n2155), .Z(c[128]) );
  XNOR U4148 ( .A(n2158), .B(n2157), .Z(c[129]) );
  XNOR U4149 ( .A(n2160), .B(n2159), .Z(c[12]) );
  XNOR U4150 ( .A(n2162), .B(n2161), .Z(c[130]) );
  XNOR U4151 ( .A(n2164), .B(n2163), .Z(c[131]) );
  XNOR U4152 ( .A(n2166), .B(n2165), .Z(c[132]) );
  XNOR U4153 ( .A(n2168), .B(n2167), .Z(c[133]) );
  XNOR U4154 ( .A(n2170), .B(n2169), .Z(c[134]) );
  XNOR U4155 ( .A(n2172), .B(n2171), .Z(c[135]) );
  XNOR U4156 ( .A(n2174), .B(n2173), .Z(c[136]) );
  XNOR U4157 ( .A(n2176), .B(n2175), .Z(c[137]) );
  XNOR U4158 ( .A(n2178), .B(n2177), .Z(c[138]) );
  XNOR U4159 ( .A(n2180), .B(n2179), .Z(c[139]) );
  XNOR U4160 ( .A(n2182), .B(n2181), .Z(c[13]) );
  XNOR U4161 ( .A(n2184), .B(n2183), .Z(c[140]) );
  XNOR U4162 ( .A(n2186), .B(n2185), .Z(c[141]) );
  XNOR U4163 ( .A(n2188), .B(n2187), .Z(c[142]) );
  XNOR U4164 ( .A(n2190), .B(n2189), .Z(c[143]) );
  XNOR U4165 ( .A(n2192), .B(n2191), .Z(c[144]) );
  XNOR U4166 ( .A(n2194), .B(n2193), .Z(c[145]) );
  XNOR U4167 ( .A(n2196), .B(n2195), .Z(c[146]) );
  XNOR U4168 ( .A(n2198), .B(n2197), .Z(c[147]) );
  XNOR U4169 ( .A(n2200), .B(n2199), .Z(c[148]) );
  XNOR U4170 ( .A(n2202), .B(n2201), .Z(c[149]) );
  XNOR U4171 ( .A(n2204), .B(n2203), .Z(c[14]) );
  XNOR U4172 ( .A(n2206), .B(n2205), .Z(c[150]) );
  XNOR U4173 ( .A(n2208), .B(n2207), .Z(c[151]) );
  XNOR U4174 ( .A(n2210), .B(n2209), .Z(c[152]) );
  XNOR U4175 ( .A(n2212), .B(n2211), .Z(c[153]) );
  XNOR U4176 ( .A(n2214), .B(n2213), .Z(c[154]) );
  XNOR U4177 ( .A(n2216), .B(n2215), .Z(c[155]) );
  XNOR U4178 ( .A(n2218), .B(n2217), .Z(c[156]) );
  XNOR U4179 ( .A(n2220), .B(n2219), .Z(c[157]) );
  XNOR U4180 ( .A(n2222), .B(n2221), .Z(c[158]) );
  XNOR U4181 ( .A(n2224), .B(n2223), .Z(c[159]) );
  XNOR U4182 ( .A(n2226), .B(n2225), .Z(c[15]) );
  XNOR U4183 ( .A(n2228), .B(n2227), .Z(c[160]) );
  XNOR U4184 ( .A(n2230), .B(n2229), .Z(c[161]) );
  XNOR U4185 ( .A(n2232), .B(n2231), .Z(c[162]) );
  XNOR U4186 ( .A(n2234), .B(n2233), .Z(c[163]) );
  XNOR U4187 ( .A(n2236), .B(n2235), .Z(c[164]) );
  XNOR U4188 ( .A(n2238), .B(n2237), .Z(c[165]) );
  XNOR U4189 ( .A(n2240), .B(n2239), .Z(c[166]) );
  XNOR U4190 ( .A(n2242), .B(n2241), .Z(c[167]) );
  XNOR U4191 ( .A(n2244), .B(n2243), .Z(c[168]) );
  XNOR U4192 ( .A(n2246), .B(n2245), .Z(c[169]) );
  XNOR U4193 ( .A(n2248), .B(n2247), .Z(c[16]) );
  XNOR U4194 ( .A(n2250), .B(n2249), .Z(c[170]) );
  XNOR U4195 ( .A(n2252), .B(n2251), .Z(c[171]) );
  XNOR U4196 ( .A(n2254), .B(n2253), .Z(c[172]) );
  XNOR U4197 ( .A(n2256), .B(n2255), .Z(c[173]) );
  XNOR U4198 ( .A(n2258), .B(n2257), .Z(c[174]) );
  XNOR U4199 ( .A(n2260), .B(n2259), .Z(c[175]) );
  XNOR U4200 ( .A(n2262), .B(n2261), .Z(c[176]) );
  XNOR U4201 ( .A(n2264), .B(n2263), .Z(c[177]) );
  XNOR U4202 ( .A(n2266), .B(n2265), .Z(c[178]) );
  XNOR U4203 ( .A(n2268), .B(n2267), .Z(c[179]) );
  XNOR U4204 ( .A(n2270), .B(n2269), .Z(c[17]) );
  XNOR U4205 ( .A(n2272), .B(n2271), .Z(c[180]) );
  XNOR U4206 ( .A(n2274), .B(n2273), .Z(c[181]) );
  XNOR U4207 ( .A(n2276), .B(n2275), .Z(c[182]) );
  XNOR U4208 ( .A(n2278), .B(n2277), .Z(c[183]) );
  XNOR U4209 ( .A(n2280), .B(n2279), .Z(c[184]) );
  XNOR U4210 ( .A(n2282), .B(n2281), .Z(c[185]) );
  XNOR U4211 ( .A(n2284), .B(n2283), .Z(c[186]) );
  XNOR U4212 ( .A(n2286), .B(n2285), .Z(c[187]) );
  XNOR U4213 ( .A(n2288), .B(n2287), .Z(c[188]) );
  XNOR U4214 ( .A(n2290), .B(n2289), .Z(c[189]) );
  XNOR U4215 ( .A(n2292), .B(n2291), .Z(c[18]) );
  XNOR U4216 ( .A(n2294), .B(n2293), .Z(c[190]) );
  XNOR U4217 ( .A(n2296), .B(n2295), .Z(c[191]) );
  XNOR U4218 ( .A(n2298), .B(n2297), .Z(c[192]) );
  XNOR U4219 ( .A(n2300), .B(n2299), .Z(c[193]) );
  XNOR U4220 ( .A(n2302), .B(n2301), .Z(c[194]) );
  XNOR U4221 ( .A(n2304), .B(n2303), .Z(c[195]) );
  XNOR U4222 ( .A(n2306), .B(n2305), .Z(c[196]) );
  XNOR U4223 ( .A(n2308), .B(n2307), .Z(c[197]) );
  XNOR U4224 ( .A(n2310), .B(n2309), .Z(c[198]) );
  XNOR U4225 ( .A(n2312), .B(n2311), .Z(c[199]) );
  XNOR U4226 ( .A(n2314), .B(n2313), .Z(c[19]) );
  XOR U4227 ( .A(b[1]), .B(a[1]), .Z(n2315) );
  XNOR U4228 ( .A(n2316), .B(n2315), .Z(c[1]) );
  XNOR U4229 ( .A(n2318), .B(n2317), .Z(c[200]) );
  XNOR U4230 ( .A(n2320), .B(n2319), .Z(c[201]) );
  XNOR U4231 ( .A(n2322), .B(n2321), .Z(c[202]) );
  XNOR U4232 ( .A(n2324), .B(n2323), .Z(c[203]) );
  XNOR U4233 ( .A(n2326), .B(n2325), .Z(c[204]) );
  XNOR U4234 ( .A(n2328), .B(n2327), .Z(c[205]) );
  XNOR U4235 ( .A(n2330), .B(n2329), .Z(c[206]) );
  XNOR U4236 ( .A(n2332), .B(n2331), .Z(c[207]) );
  XNOR U4237 ( .A(n2334), .B(n2333), .Z(c[208]) );
  XNOR U4238 ( .A(n2336), .B(n2335), .Z(c[209]) );
  XNOR U4239 ( .A(n2338), .B(n2337), .Z(c[20]) );
  XNOR U4240 ( .A(n2340), .B(n2339), .Z(c[210]) );
  XNOR U4241 ( .A(n2342), .B(n2341), .Z(c[211]) );
  XNOR U4242 ( .A(n2344), .B(n2343), .Z(c[212]) );
  XNOR U4243 ( .A(n2346), .B(n2345), .Z(c[213]) );
  XNOR U4244 ( .A(n2348), .B(n2347), .Z(c[214]) );
  XNOR U4245 ( .A(n2350), .B(n2349), .Z(c[215]) );
  XNOR U4246 ( .A(n2352), .B(n2351), .Z(c[216]) );
  XNOR U4247 ( .A(n2354), .B(n2353), .Z(c[217]) );
  XNOR U4248 ( .A(n2356), .B(n2355), .Z(c[218]) );
  XNOR U4249 ( .A(n2358), .B(n2357), .Z(c[219]) );
  XNOR U4250 ( .A(n2360), .B(n2359), .Z(c[21]) );
  XNOR U4251 ( .A(n2362), .B(n2361), .Z(c[220]) );
  XNOR U4252 ( .A(n2364), .B(n2363), .Z(c[221]) );
  XNOR U4253 ( .A(n2366), .B(n2365), .Z(c[222]) );
  XNOR U4254 ( .A(n2368), .B(n2367), .Z(c[223]) );
  XNOR U4255 ( .A(n2370), .B(n2369), .Z(c[224]) );
  XNOR U4256 ( .A(n2372), .B(n2371), .Z(c[225]) );
  XNOR U4257 ( .A(n2374), .B(n2373), .Z(c[226]) );
  XNOR U4258 ( .A(n2376), .B(n2375), .Z(c[227]) );
  XNOR U4259 ( .A(n2378), .B(n2377), .Z(c[228]) );
  XNOR U4260 ( .A(n2380), .B(n2379), .Z(c[229]) );
  XNOR U4261 ( .A(n2382), .B(n2381), .Z(c[22]) );
  XNOR U4262 ( .A(n2384), .B(n2383), .Z(c[230]) );
  XNOR U4263 ( .A(n2386), .B(n2385), .Z(c[231]) );
  XNOR U4264 ( .A(n2388), .B(n2387), .Z(c[232]) );
  XNOR U4265 ( .A(n2390), .B(n2389), .Z(c[233]) );
  XNOR U4266 ( .A(n2392), .B(n2391), .Z(c[234]) );
  XNOR U4267 ( .A(n2394), .B(n2393), .Z(c[235]) );
  XNOR U4268 ( .A(n2396), .B(n2395), .Z(c[236]) );
  XNOR U4269 ( .A(n2398), .B(n2397), .Z(c[237]) );
  XNOR U4270 ( .A(n2400), .B(n2399), .Z(c[238]) );
  XNOR U4271 ( .A(n2402), .B(n2401), .Z(c[239]) );
  XNOR U4272 ( .A(n2404), .B(n2403), .Z(c[23]) );
  XNOR U4273 ( .A(n2406), .B(n2405), .Z(c[240]) );
  XNOR U4274 ( .A(n2408), .B(n2407), .Z(c[241]) );
  XNOR U4275 ( .A(n2410), .B(n2409), .Z(c[242]) );
  XNOR U4276 ( .A(n2412), .B(n2411), .Z(c[243]) );
  XNOR U4277 ( .A(n2414), .B(n2413), .Z(c[244]) );
  XNOR U4278 ( .A(n2416), .B(n2415), .Z(c[245]) );
  XNOR U4279 ( .A(n2418), .B(n2417), .Z(c[246]) );
  XNOR U4280 ( .A(n2420), .B(n2419), .Z(c[247]) );
  XNOR U4281 ( .A(n2422), .B(n2421), .Z(c[248]) );
  XNOR U4282 ( .A(n2424), .B(n2423), .Z(c[249]) );
  XNOR U4283 ( .A(n2426), .B(n2425), .Z(c[24]) );
  XNOR U4284 ( .A(n2428), .B(n2427), .Z(c[250]) );
  XNOR U4285 ( .A(n2430), .B(n2429), .Z(c[251]) );
  XNOR U4286 ( .A(n2432), .B(n2431), .Z(c[252]) );
  XNOR U4287 ( .A(n2434), .B(n2433), .Z(c[253]) );
  XNOR U4288 ( .A(n2436), .B(n2435), .Z(c[254]) );
  XNOR U4289 ( .A(n2438), .B(n2437), .Z(c[255]) );
  XNOR U4290 ( .A(n2440), .B(n2439), .Z(c[256]) );
  XNOR U4291 ( .A(n2442), .B(n2441), .Z(c[257]) );
  XNOR U4292 ( .A(n2444), .B(n2443), .Z(c[258]) );
  XNOR U4293 ( .A(n2446), .B(n2445), .Z(c[259]) );
  XNOR U4294 ( .A(n2448), .B(n2447), .Z(c[25]) );
  XNOR U4295 ( .A(n2450), .B(n2449), .Z(c[260]) );
  XNOR U4296 ( .A(n2452), .B(n2451), .Z(c[261]) );
  XNOR U4297 ( .A(n2454), .B(n2453), .Z(c[262]) );
  XNOR U4298 ( .A(n2456), .B(n2455), .Z(c[263]) );
  XNOR U4299 ( .A(n2458), .B(n2457), .Z(c[264]) );
  XNOR U4300 ( .A(n2460), .B(n2459), .Z(c[265]) );
  XNOR U4301 ( .A(n2462), .B(n2461), .Z(c[266]) );
  XNOR U4302 ( .A(n2464), .B(n2463), .Z(c[267]) );
  XNOR U4303 ( .A(n2466), .B(n2465), .Z(c[268]) );
  XNOR U4304 ( .A(n2468), .B(n2467), .Z(c[269]) );
  XNOR U4305 ( .A(n2470), .B(n2469), .Z(c[26]) );
  XNOR U4306 ( .A(n2472), .B(n2471), .Z(c[270]) );
  XNOR U4307 ( .A(n2474), .B(n2473), .Z(c[271]) );
  XNOR U4308 ( .A(n2476), .B(n2475), .Z(c[272]) );
  XNOR U4309 ( .A(n2478), .B(n2477), .Z(c[273]) );
  XNOR U4310 ( .A(n2480), .B(n2479), .Z(c[274]) );
  XNOR U4311 ( .A(n2482), .B(n2481), .Z(c[275]) );
  XNOR U4312 ( .A(n2484), .B(n2483), .Z(c[276]) );
  XNOR U4313 ( .A(n2486), .B(n2485), .Z(c[277]) );
  XNOR U4314 ( .A(n2488), .B(n2487), .Z(c[278]) );
  XNOR U4315 ( .A(n2490), .B(n2489), .Z(c[279]) );
  XNOR U4316 ( .A(n2492), .B(n2491), .Z(c[27]) );
  XNOR U4317 ( .A(n2494), .B(n2493), .Z(c[280]) );
  XNOR U4318 ( .A(n2496), .B(n2495), .Z(c[281]) );
  XNOR U4319 ( .A(n2498), .B(n2497), .Z(c[282]) );
  XNOR U4320 ( .A(n2500), .B(n2499), .Z(c[283]) );
  XNOR U4321 ( .A(n2502), .B(n2501), .Z(c[284]) );
  XNOR U4322 ( .A(n2504), .B(n2503), .Z(c[285]) );
  XNOR U4323 ( .A(n2506), .B(n2505), .Z(c[286]) );
  XNOR U4324 ( .A(n2508), .B(n2507), .Z(c[287]) );
  XNOR U4325 ( .A(n2510), .B(n2509), .Z(c[288]) );
  XNOR U4326 ( .A(n2512), .B(n2511), .Z(c[289]) );
  XNOR U4327 ( .A(n2514), .B(n2513), .Z(c[28]) );
  XNOR U4328 ( .A(n2516), .B(n2515), .Z(c[290]) );
  XNOR U4329 ( .A(n2518), .B(n2517), .Z(c[291]) );
  XNOR U4330 ( .A(n2520), .B(n2519), .Z(c[292]) );
  XNOR U4331 ( .A(n2522), .B(n2521), .Z(c[293]) );
  XNOR U4332 ( .A(n2524), .B(n2523), .Z(c[294]) );
  XNOR U4333 ( .A(n2526), .B(n2525), .Z(c[295]) );
  XNOR U4334 ( .A(n2528), .B(n2527), .Z(c[296]) );
  XNOR U4335 ( .A(n2530), .B(n2529), .Z(c[297]) );
  XNOR U4336 ( .A(n2532), .B(n2531), .Z(c[298]) );
  XNOR U4337 ( .A(n2534), .B(n2533), .Z(c[299]) );
  XNOR U4338 ( .A(n2536), .B(n2535), .Z(c[29]) );
  XNOR U4339 ( .A(n2538), .B(n2537), .Z(c[2]) );
  XNOR U4340 ( .A(n2540), .B(n2539), .Z(c[300]) );
  XNOR U4341 ( .A(n2542), .B(n2541), .Z(c[301]) );
  XNOR U4342 ( .A(n2544), .B(n2543), .Z(c[302]) );
  XNOR U4343 ( .A(n2546), .B(n2545), .Z(c[303]) );
  XNOR U4344 ( .A(n2548), .B(n2547), .Z(c[304]) );
  XNOR U4345 ( .A(n2550), .B(n2549), .Z(c[305]) );
  XNOR U4346 ( .A(n2552), .B(n2551), .Z(c[306]) );
  XNOR U4347 ( .A(n2554), .B(n2553), .Z(c[307]) );
  XNOR U4348 ( .A(n2556), .B(n2555), .Z(c[308]) );
  XNOR U4349 ( .A(n2558), .B(n2557), .Z(c[309]) );
  XNOR U4350 ( .A(n2560), .B(n2559), .Z(c[30]) );
  XNOR U4351 ( .A(n2562), .B(n2561), .Z(c[310]) );
  XNOR U4352 ( .A(n2564), .B(n2563), .Z(c[311]) );
  XNOR U4353 ( .A(n2566), .B(n2565), .Z(c[312]) );
  XNOR U4354 ( .A(n2568), .B(n2567), .Z(c[313]) );
  XNOR U4355 ( .A(n2570), .B(n2569), .Z(c[314]) );
  XNOR U4356 ( .A(n2572), .B(n2571), .Z(c[315]) );
  XNOR U4357 ( .A(n2574), .B(n2573), .Z(c[316]) );
  XNOR U4358 ( .A(n2576), .B(n2575), .Z(c[317]) );
  XNOR U4359 ( .A(n2578), .B(n2577), .Z(c[318]) );
  XNOR U4360 ( .A(n2580), .B(n2579), .Z(c[319]) );
  XNOR U4361 ( .A(n2582), .B(n2581), .Z(c[31]) );
  XNOR U4362 ( .A(n2584), .B(n2583), .Z(c[320]) );
  XNOR U4363 ( .A(n2586), .B(n2585), .Z(c[321]) );
  XNOR U4364 ( .A(n2588), .B(n2587), .Z(c[322]) );
  XNOR U4365 ( .A(n2590), .B(n2589), .Z(c[323]) );
  XNOR U4366 ( .A(n2592), .B(n2591), .Z(c[324]) );
  XNOR U4367 ( .A(n2594), .B(n2593), .Z(c[325]) );
  XNOR U4368 ( .A(n2596), .B(n2595), .Z(c[326]) );
  XNOR U4369 ( .A(n2598), .B(n2597), .Z(c[327]) );
  XNOR U4370 ( .A(n2600), .B(n2599), .Z(c[328]) );
  XNOR U4371 ( .A(n2602), .B(n2601), .Z(c[329]) );
  XNOR U4372 ( .A(n2604), .B(n2603), .Z(c[32]) );
  XNOR U4373 ( .A(n2606), .B(n2605), .Z(c[330]) );
  XNOR U4374 ( .A(n2608), .B(n2607), .Z(c[331]) );
  XNOR U4375 ( .A(n2610), .B(n2609), .Z(c[332]) );
  XNOR U4376 ( .A(n2612), .B(n2611), .Z(c[333]) );
  XNOR U4377 ( .A(n2614), .B(n2613), .Z(c[334]) );
  XNOR U4378 ( .A(n2616), .B(n2615), .Z(c[335]) );
  XNOR U4379 ( .A(n2618), .B(n2617), .Z(c[336]) );
  XNOR U4380 ( .A(n2620), .B(n2619), .Z(c[337]) );
  XNOR U4381 ( .A(n2622), .B(n2621), .Z(c[338]) );
  XNOR U4382 ( .A(n2624), .B(n2623), .Z(c[339]) );
  XNOR U4383 ( .A(n2626), .B(n2625), .Z(c[33]) );
  XNOR U4384 ( .A(n2628), .B(n2627), .Z(c[340]) );
  XNOR U4385 ( .A(n2630), .B(n2629), .Z(c[341]) );
  XNOR U4386 ( .A(n2632), .B(n2631), .Z(c[342]) );
  XNOR U4387 ( .A(n2634), .B(n2633), .Z(c[343]) );
  XNOR U4388 ( .A(n2636), .B(n2635), .Z(c[344]) );
  XNOR U4389 ( .A(n2638), .B(n2637), .Z(c[345]) );
  XNOR U4390 ( .A(n2640), .B(n2639), .Z(c[346]) );
  XNOR U4391 ( .A(n2642), .B(n2641), .Z(c[347]) );
  XNOR U4392 ( .A(n2644), .B(n2643), .Z(c[348]) );
  XNOR U4393 ( .A(n2646), .B(n2645), .Z(c[349]) );
  XNOR U4394 ( .A(n2648), .B(n2647), .Z(c[34]) );
  XNOR U4395 ( .A(n2650), .B(n2649), .Z(c[350]) );
  XNOR U4396 ( .A(n2652), .B(n2651), .Z(c[351]) );
  XNOR U4397 ( .A(n2654), .B(n2653), .Z(c[352]) );
  XNOR U4398 ( .A(n2656), .B(n2655), .Z(c[353]) );
  XNOR U4399 ( .A(n2658), .B(n2657), .Z(c[354]) );
  XNOR U4400 ( .A(n2660), .B(n2659), .Z(c[355]) );
  XNOR U4401 ( .A(n2662), .B(n2661), .Z(c[356]) );
  XNOR U4402 ( .A(n2664), .B(n2663), .Z(c[357]) );
  XNOR U4403 ( .A(n2666), .B(n2665), .Z(c[358]) );
  XNOR U4404 ( .A(n2668), .B(n2667), .Z(c[359]) );
  XNOR U4405 ( .A(n2670), .B(n2669), .Z(c[35]) );
  XNOR U4406 ( .A(n2672), .B(n2671), .Z(c[360]) );
  XNOR U4407 ( .A(n2674), .B(n2673), .Z(c[361]) );
  XNOR U4408 ( .A(n2676), .B(n2675), .Z(c[362]) );
  XNOR U4409 ( .A(n2678), .B(n2677), .Z(c[363]) );
  XNOR U4410 ( .A(n2680), .B(n2679), .Z(c[364]) );
  XNOR U4411 ( .A(n2682), .B(n2681), .Z(c[365]) );
  XNOR U4412 ( .A(n2684), .B(n2683), .Z(c[366]) );
  XNOR U4413 ( .A(n2686), .B(n2685), .Z(c[367]) );
  XNOR U4414 ( .A(n2688), .B(n2687), .Z(c[368]) );
  XNOR U4415 ( .A(n2690), .B(n2689), .Z(c[369]) );
  XNOR U4416 ( .A(n2692), .B(n2691), .Z(c[36]) );
  XNOR U4417 ( .A(n2694), .B(n2693), .Z(c[370]) );
  XNOR U4418 ( .A(n2696), .B(n2695), .Z(c[371]) );
  XNOR U4419 ( .A(n2698), .B(n2697), .Z(c[372]) );
  XNOR U4420 ( .A(n2700), .B(n2699), .Z(c[373]) );
  XNOR U4421 ( .A(n2702), .B(n2701), .Z(c[374]) );
  XNOR U4422 ( .A(n2704), .B(n2703), .Z(c[375]) );
  XNOR U4423 ( .A(n2706), .B(n2705), .Z(c[376]) );
  XNOR U4424 ( .A(n2708), .B(n2707), .Z(c[377]) );
  XNOR U4425 ( .A(n2710), .B(n2709), .Z(c[378]) );
  XNOR U4426 ( .A(n2712), .B(n2711), .Z(c[379]) );
  XNOR U4427 ( .A(n2714), .B(n2713), .Z(c[37]) );
  XNOR U4428 ( .A(n2716), .B(n2715), .Z(c[380]) );
  XNOR U4429 ( .A(n2718), .B(n2717), .Z(c[381]) );
  XNOR U4430 ( .A(n2720), .B(n2719), .Z(c[382]) );
  XNOR U4431 ( .A(n2722), .B(n2721), .Z(c[383]) );
  XNOR U4432 ( .A(n2724), .B(n2723), .Z(c[384]) );
  XNOR U4433 ( .A(n2726), .B(n2725), .Z(c[385]) );
  XNOR U4434 ( .A(n2728), .B(n2727), .Z(c[386]) );
  XNOR U4435 ( .A(n2730), .B(n2729), .Z(c[387]) );
  XNOR U4436 ( .A(n2732), .B(n2731), .Z(c[388]) );
  XNOR U4437 ( .A(n2734), .B(n2733), .Z(c[389]) );
  XNOR U4438 ( .A(n2736), .B(n2735), .Z(c[38]) );
  XNOR U4439 ( .A(n2738), .B(n2737), .Z(c[390]) );
  XNOR U4440 ( .A(n2740), .B(n2739), .Z(c[391]) );
  XNOR U4441 ( .A(n2742), .B(n2741), .Z(c[392]) );
  XNOR U4442 ( .A(n2744), .B(n2743), .Z(c[393]) );
  XNOR U4443 ( .A(n2746), .B(n2745), .Z(c[394]) );
  XNOR U4444 ( .A(n2748), .B(n2747), .Z(c[395]) );
  XNOR U4445 ( .A(n2750), .B(n2749), .Z(c[396]) );
  XNOR U4446 ( .A(n2752), .B(n2751), .Z(c[397]) );
  XNOR U4447 ( .A(n2754), .B(n2753), .Z(c[398]) );
  XNOR U4448 ( .A(n2756), .B(n2755), .Z(c[399]) );
  XNOR U4449 ( .A(n2758), .B(n2757), .Z(c[39]) );
  XOR U4450 ( .A(n2760), .B(n2759), .Z(c[3]) );
  XNOR U4451 ( .A(n2762), .B(n2761), .Z(c[400]) );
  XNOR U4452 ( .A(n2764), .B(n2763), .Z(c[401]) );
  XNOR U4453 ( .A(n2766), .B(n2765), .Z(c[402]) );
  XNOR U4454 ( .A(n2768), .B(n2767), .Z(c[403]) );
  XNOR U4455 ( .A(n2770), .B(n2769), .Z(c[404]) );
  XNOR U4456 ( .A(n2772), .B(n2771), .Z(c[405]) );
  XNOR U4457 ( .A(n2774), .B(n2773), .Z(c[406]) );
  XNOR U4458 ( .A(n2776), .B(n2775), .Z(c[407]) );
  XNOR U4459 ( .A(n2778), .B(n2777), .Z(c[408]) );
  XNOR U4460 ( .A(n2780), .B(n2779), .Z(c[409]) );
  XNOR U4461 ( .A(n2782), .B(n2781), .Z(c[40]) );
  XNOR U4462 ( .A(n2784), .B(n2783), .Z(c[410]) );
  XNOR U4463 ( .A(n2786), .B(n2785), .Z(c[411]) );
  XNOR U4464 ( .A(n2788), .B(n2787), .Z(c[412]) );
  XNOR U4465 ( .A(n2790), .B(n2789), .Z(c[413]) );
  XNOR U4466 ( .A(n2792), .B(n2791), .Z(c[414]) );
  XNOR U4467 ( .A(n2794), .B(n2793), .Z(c[415]) );
  XNOR U4468 ( .A(n2796), .B(n2795), .Z(c[416]) );
  XNOR U4469 ( .A(n2798), .B(n2797), .Z(c[417]) );
  XNOR U4470 ( .A(n2800), .B(n2799), .Z(c[418]) );
  XNOR U4471 ( .A(n2802), .B(n2801), .Z(c[419]) );
  XNOR U4472 ( .A(n2804), .B(n2803), .Z(c[41]) );
  XNOR U4473 ( .A(n2806), .B(n2805), .Z(c[420]) );
  XNOR U4474 ( .A(n2808), .B(n2807), .Z(c[421]) );
  XNOR U4475 ( .A(n2810), .B(n2809), .Z(c[422]) );
  XNOR U4476 ( .A(n2812), .B(n2811), .Z(c[423]) );
  XNOR U4477 ( .A(n2814), .B(n2813), .Z(c[424]) );
  XNOR U4478 ( .A(n2816), .B(n2815), .Z(c[425]) );
  XNOR U4479 ( .A(n2818), .B(n2817), .Z(c[426]) );
  XNOR U4480 ( .A(n2820), .B(n2819), .Z(c[427]) );
  XNOR U4481 ( .A(n2822), .B(n2821), .Z(c[428]) );
  XNOR U4482 ( .A(n2824), .B(n2823), .Z(c[429]) );
  XNOR U4483 ( .A(n2826), .B(n2825), .Z(c[42]) );
  XNOR U4484 ( .A(n2828), .B(n2827), .Z(c[430]) );
  XNOR U4485 ( .A(n2830), .B(n2829), .Z(c[431]) );
  XNOR U4486 ( .A(n2832), .B(n2831), .Z(c[432]) );
  XNOR U4487 ( .A(n2834), .B(n2833), .Z(c[433]) );
  XNOR U4488 ( .A(n2836), .B(n2835), .Z(c[434]) );
  XNOR U4489 ( .A(n2838), .B(n2837), .Z(c[435]) );
  XNOR U4490 ( .A(n2840), .B(n2839), .Z(c[436]) );
  XNOR U4491 ( .A(n2842), .B(n2841), .Z(c[437]) );
  XNOR U4492 ( .A(n2844), .B(n2843), .Z(c[438]) );
  XNOR U4493 ( .A(n2846), .B(n2845), .Z(c[439]) );
  XNOR U4494 ( .A(n2848), .B(n2847), .Z(c[43]) );
  XNOR U4495 ( .A(n2850), .B(n2849), .Z(c[440]) );
  XNOR U4496 ( .A(n2852), .B(n2851), .Z(c[441]) );
  XNOR U4497 ( .A(n2854), .B(n2853), .Z(c[442]) );
  XNOR U4498 ( .A(n2856), .B(n2855), .Z(c[443]) );
  XNOR U4499 ( .A(n2858), .B(n2857), .Z(c[444]) );
  XNOR U4500 ( .A(n2860), .B(n2859), .Z(c[445]) );
  XNOR U4501 ( .A(n2862), .B(n2861), .Z(c[446]) );
  XNOR U4502 ( .A(n2864), .B(n2863), .Z(c[447]) );
  XNOR U4503 ( .A(n2866), .B(n2865), .Z(c[448]) );
  XNOR U4504 ( .A(n2868), .B(n2867), .Z(c[449]) );
  XNOR U4505 ( .A(n2870), .B(n2869), .Z(c[44]) );
  XNOR U4506 ( .A(n2872), .B(n2871), .Z(c[450]) );
  XNOR U4507 ( .A(n2874), .B(n2873), .Z(c[451]) );
  XNOR U4508 ( .A(n2876), .B(n2875), .Z(c[452]) );
  XNOR U4509 ( .A(n2878), .B(n2877), .Z(c[453]) );
  XNOR U4510 ( .A(n2880), .B(n2879), .Z(c[454]) );
  XNOR U4511 ( .A(n2882), .B(n2881), .Z(c[455]) );
  XNOR U4512 ( .A(n2884), .B(n2883), .Z(c[456]) );
  XNOR U4513 ( .A(n2886), .B(n2885), .Z(c[457]) );
  XNOR U4514 ( .A(n2888), .B(n2887), .Z(c[458]) );
  XNOR U4515 ( .A(n2890), .B(n2889), .Z(c[459]) );
  XNOR U4516 ( .A(n2892), .B(n2891), .Z(c[45]) );
  XNOR U4517 ( .A(n2894), .B(n2893), .Z(c[460]) );
  XNOR U4518 ( .A(n2896), .B(n2895), .Z(c[461]) );
  XNOR U4519 ( .A(n2898), .B(n2897), .Z(c[462]) );
  XNOR U4520 ( .A(n2900), .B(n2899), .Z(c[463]) );
  XNOR U4521 ( .A(n2902), .B(n2901), .Z(c[464]) );
  XNOR U4522 ( .A(n2904), .B(n2903), .Z(c[465]) );
  XNOR U4523 ( .A(n2906), .B(n2905), .Z(c[466]) );
  XNOR U4524 ( .A(n2908), .B(n2907), .Z(c[467]) );
  XNOR U4525 ( .A(n2910), .B(n2909), .Z(c[468]) );
  XNOR U4526 ( .A(n2912), .B(n2911), .Z(c[469]) );
  XNOR U4527 ( .A(n2914), .B(n2913), .Z(c[46]) );
  XNOR U4528 ( .A(n2916), .B(n2915), .Z(c[470]) );
  XNOR U4529 ( .A(n2918), .B(n2917), .Z(c[471]) );
  XNOR U4530 ( .A(n2920), .B(n2919), .Z(c[472]) );
  XNOR U4531 ( .A(n2922), .B(n2921), .Z(c[473]) );
  XNOR U4532 ( .A(n2924), .B(n2923), .Z(c[474]) );
  XNOR U4533 ( .A(n2926), .B(n2925), .Z(c[475]) );
  XNOR U4534 ( .A(n2928), .B(n2927), .Z(c[476]) );
  XNOR U4535 ( .A(n2930), .B(n2929), .Z(c[477]) );
  XNOR U4536 ( .A(n2932), .B(n2931), .Z(c[478]) );
  XNOR U4537 ( .A(n2934), .B(n2933), .Z(c[479]) );
  XNOR U4538 ( .A(n2936), .B(n2935), .Z(c[47]) );
  XNOR U4539 ( .A(n2938), .B(n2937), .Z(c[480]) );
  XNOR U4540 ( .A(n2940), .B(n2939), .Z(c[481]) );
  XNOR U4541 ( .A(n2942), .B(n2941), .Z(c[482]) );
  XNOR U4542 ( .A(n2944), .B(n2943), .Z(c[483]) );
  XNOR U4543 ( .A(n2946), .B(n2945), .Z(c[484]) );
  XNOR U4544 ( .A(n2948), .B(n2947), .Z(c[485]) );
  XNOR U4545 ( .A(n2950), .B(n2949), .Z(c[486]) );
  XNOR U4546 ( .A(n2952), .B(n2951), .Z(c[487]) );
  XNOR U4547 ( .A(n2954), .B(n2953), .Z(c[488]) );
  XNOR U4548 ( .A(n2956), .B(n2955), .Z(c[489]) );
  XNOR U4549 ( .A(n2958), .B(n2957), .Z(c[48]) );
  XNOR U4550 ( .A(n2960), .B(n2959), .Z(c[490]) );
  XNOR U4551 ( .A(n2962), .B(n2961), .Z(c[491]) );
  XNOR U4552 ( .A(n2964), .B(n2963), .Z(c[492]) );
  XNOR U4553 ( .A(n2966), .B(n2965), .Z(c[493]) );
  XNOR U4554 ( .A(n2968), .B(n2967), .Z(c[494]) );
  XNOR U4555 ( .A(n2970), .B(n2969), .Z(c[495]) );
  XNOR U4556 ( .A(n2972), .B(n2971), .Z(c[496]) );
  XNOR U4557 ( .A(n2974), .B(n2973), .Z(c[497]) );
  XNOR U4558 ( .A(n2976), .B(n2975), .Z(c[498]) );
  XNOR U4559 ( .A(n2978), .B(n2977), .Z(c[499]) );
  XNOR U4560 ( .A(n2980), .B(n2979), .Z(c[49]) );
  XNOR U4561 ( .A(n2982), .B(n2981), .Z(c[4]) );
  XNOR U4562 ( .A(n2984), .B(n2983), .Z(c[500]) );
  XNOR U4563 ( .A(n2986), .B(n2985), .Z(c[501]) );
  XNOR U4564 ( .A(n2988), .B(n2987), .Z(c[502]) );
  XNOR U4565 ( .A(n2990), .B(n2989), .Z(c[503]) );
  XNOR U4566 ( .A(n2992), .B(n2991), .Z(c[504]) );
  XNOR U4567 ( .A(n2994), .B(n2993), .Z(c[505]) );
  XNOR U4568 ( .A(n2996), .B(n2995), .Z(c[506]) );
  XNOR U4569 ( .A(n2998), .B(n2997), .Z(c[507]) );
  XNOR U4570 ( .A(n3000), .B(n2999), .Z(c[508]) );
  XNOR U4571 ( .A(n3002), .B(n3001), .Z(c[509]) );
  XNOR U4572 ( .A(n3004), .B(n3003), .Z(c[50]) );
  XNOR U4573 ( .A(n3006), .B(n3005), .Z(c[510]) );
  XNOR U4574 ( .A(n3008), .B(n3007), .Z(c[511]) );
  XNOR U4575 ( .A(n3010), .B(n3009), .Z(c[512]) );
  XNOR U4576 ( .A(n3012), .B(n3011), .Z(c[513]) );
  XNOR U4577 ( .A(n3014), .B(n3013), .Z(c[514]) );
  XNOR U4578 ( .A(n3016), .B(n3015), .Z(c[515]) );
  XNOR U4579 ( .A(n3018), .B(n3017), .Z(c[516]) );
  XNOR U4580 ( .A(n3020), .B(n3019), .Z(c[517]) );
  XNOR U4581 ( .A(n3022), .B(n3021), .Z(c[518]) );
  XNOR U4582 ( .A(n3024), .B(n3023), .Z(c[519]) );
  XNOR U4583 ( .A(n3026), .B(n3025), .Z(c[51]) );
  XNOR U4584 ( .A(n3028), .B(n3027), .Z(c[520]) );
  XNOR U4585 ( .A(n3030), .B(n3029), .Z(c[521]) );
  XNOR U4586 ( .A(n3032), .B(n3031), .Z(c[522]) );
  XNOR U4587 ( .A(n3034), .B(n3033), .Z(c[523]) );
  XNOR U4588 ( .A(n3036), .B(n3035), .Z(c[524]) );
  XNOR U4589 ( .A(n3038), .B(n3037), .Z(c[525]) );
  XNOR U4590 ( .A(n3040), .B(n3039), .Z(c[526]) );
  XNOR U4591 ( .A(n3042), .B(n3041), .Z(c[527]) );
  XNOR U4592 ( .A(n3044), .B(n3043), .Z(c[528]) );
  XNOR U4593 ( .A(n3046), .B(n3045), .Z(c[529]) );
  XNOR U4594 ( .A(n3048), .B(n3047), .Z(c[52]) );
  XNOR U4595 ( .A(n3050), .B(n3049), .Z(c[530]) );
  XNOR U4596 ( .A(n3052), .B(n3051), .Z(c[531]) );
  XNOR U4597 ( .A(n3054), .B(n3053), .Z(c[532]) );
  XNOR U4598 ( .A(n3056), .B(n3055), .Z(c[533]) );
  XNOR U4599 ( .A(n3058), .B(n3057), .Z(c[534]) );
  XNOR U4600 ( .A(n3060), .B(n3059), .Z(c[535]) );
  XNOR U4601 ( .A(n3062), .B(n3061), .Z(c[536]) );
  XNOR U4602 ( .A(n3064), .B(n3063), .Z(c[537]) );
  XNOR U4603 ( .A(n3066), .B(n3065), .Z(c[538]) );
  XNOR U4604 ( .A(n3068), .B(n3067), .Z(c[539]) );
  XNOR U4605 ( .A(n3070), .B(n3069), .Z(c[53]) );
  XNOR U4606 ( .A(n3072), .B(n3071), .Z(c[540]) );
  XNOR U4607 ( .A(n3074), .B(n3073), .Z(c[541]) );
  XNOR U4608 ( .A(n3076), .B(n3075), .Z(c[542]) );
  XNOR U4609 ( .A(n3078), .B(n3077), .Z(c[543]) );
  XNOR U4610 ( .A(n3080), .B(n3079), .Z(c[544]) );
  XNOR U4611 ( .A(n3082), .B(n3081), .Z(c[545]) );
  XNOR U4612 ( .A(n3084), .B(n3083), .Z(c[546]) );
  XNOR U4613 ( .A(n3086), .B(n3085), .Z(c[547]) );
  XNOR U4614 ( .A(n3088), .B(n3087), .Z(c[548]) );
  XNOR U4615 ( .A(n3090), .B(n3089), .Z(c[549]) );
  XNOR U4616 ( .A(n3092), .B(n3091), .Z(c[54]) );
  XNOR U4617 ( .A(n3094), .B(n3093), .Z(c[550]) );
  XNOR U4618 ( .A(n3096), .B(n3095), .Z(c[551]) );
  XNOR U4619 ( .A(n3098), .B(n3097), .Z(c[552]) );
  XNOR U4620 ( .A(n3100), .B(n3099), .Z(c[553]) );
  XNOR U4621 ( .A(n3102), .B(n3101), .Z(c[554]) );
  XNOR U4622 ( .A(n3104), .B(n3103), .Z(c[555]) );
  XNOR U4623 ( .A(n3106), .B(n3105), .Z(c[556]) );
  XNOR U4624 ( .A(n3108), .B(n3107), .Z(c[557]) );
  XNOR U4625 ( .A(n3110), .B(n3109), .Z(c[558]) );
  XNOR U4626 ( .A(n3112), .B(n3111), .Z(c[559]) );
  XNOR U4627 ( .A(n3114), .B(n3113), .Z(c[55]) );
  XNOR U4628 ( .A(n3116), .B(n3115), .Z(c[560]) );
  XNOR U4629 ( .A(n3118), .B(n3117), .Z(c[561]) );
  XNOR U4630 ( .A(n3120), .B(n3119), .Z(c[562]) );
  XNOR U4631 ( .A(n3122), .B(n3121), .Z(c[563]) );
  XNOR U4632 ( .A(n3124), .B(n3123), .Z(c[564]) );
  XNOR U4633 ( .A(n3126), .B(n3125), .Z(c[565]) );
  XNOR U4634 ( .A(n3128), .B(n3127), .Z(c[566]) );
  XNOR U4635 ( .A(n3130), .B(n3129), .Z(c[567]) );
  XNOR U4636 ( .A(n3132), .B(n3131), .Z(c[568]) );
  XNOR U4637 ( .A(n3134), .B(n3133), .Z(c[569]) );
  XNOR U4638 ( .A(n3136), .B(n3135), .Z(c[56]) );
  XNOR U4639 ( .A(n3138), .B(n3137), .Z(c[570]) );
  XNOR U4640 ( .A(n3140), .B(n3139), .Z(c[571]) );
  XNOR U4641 ( .A(n3142), .B(n3141), .Z(c[572]) );
  XNOR U4642 ( .A(n3144), .B(n3143), .Z(c[573]) );
  XNOR U4643 ( .A(n3146), .B(n3145), .Z(c[574]) );
  XNOR U4644 ( .A(n3148), .B(n3147), .Z(c[575]) );
  XNOR U4645 ( .A(n3150), .B(n3149), .Z(c[576]) );
  XNOR U4646 ( .A(n3152), .B(n3151), .Z(c[577]) );
  XNOR U4647 ( .A(n3154), .B(n3153), .Z(c[578]) );
  XNOR U4648 ( .A(n3156), .B(n3155), .Z(c[579]) );
  XNOR U4649 ( .A(n3158), .B(n3157), .Z(c[57]) );
  XNOR U4650 ( .A(n3160), .B(n3159), .Z(c[580]) );
  XNOR U4651 ( .A(n3162), .B(n3161), .Z(c[581]) );
  XNOR U4652 ( .A(n3164), .B(n3163), .Z(c[582]) );
  XNOR U4653 ( .A(n3166), .B(n3165), .Z(c[583]) );
  XNOR U4654 ( .A(n3168), .B(n3167), .Z(c[584]) );
  XNOR U4655 ( .A(n3170), .B(n3169), .Z(c[585]) );
  XNOR U4656 ( .A(n3172), .B(n3171), .Z(c[586]) );
  XNOR U4657 ( .A(n3174), .B(n3173), .Z(c[587]) );
  XNOR U4658 ( .A(n3176), .B(n3175), .Z(c[588]) );
  XNOR U4659 ( .A(n3178), .B(n3177), .Z(c[589]) );
  XNOR U4660 ( .A(n3180), .B(n3179), .Z(c[58]) );
  XNOR U4661 ( .A(n3182), .B(n3181), .Z(c[590]) );
  XNOR U4662 ( .A(n3184), .B(n3183), .Z(c[591]) );
  XNOR U4663 ( .A(n3186), .B(n3185), .Z(c[592]) );
  XNOR U4664 ( .A(n3188), .B(n3187), .Z(c[593]) );
  XNOR U4665 ( .A(n3190), .B(n3189), .Z(c[594]) );
  XNOR U4666 ( .A(n3192), .B(n3191), .Z(c[595]) );
  XNOR U4667 ( .A(n3194), .B(n3193), .Z(c[596]) );
  XNOR U4668 ( .A(n3196), .B(n3195), .Z(c[597]) );
  XNOR U4669 ( .A(n3198), .B(n3197), .Z(c[598]) );
  XNOR U4670 ( .A(n3200), .B(n3199), .Z(c[599]) );
  XNOR U4671 ( .A(n3202), .B(n3201), .Z(c[59]) );
  XNOR U4672 ( .A(n3204), .B(n3203), .Z(c[5]) );
  XNOR U4673 ( .A(n3206), .B(n3205), .Z(c[600]) );
  XNOR U4674 ( .A(n3208), .B(n3207), .Z(c[601]) );
  XNOR U4675 ( .A(n3210), .B(n3209), .Z(c[602]) );
  XNOR U4676 ( .A(n3212), .B(n3211), .Z(c[603]) );
  XNOR U4677 ( .A(n3214), .B(n3213), .Z(c[604]) );
  XNOR U4678 ( .A(n3216), .B(n3215), .Z(c[605]) );
  XNOR U4679 ( .A(n3218), .B(n3217), .Z(c[606]) );
  XNOR U4680 ( .A(n3220), .B(n3219), .Z(c[607]) );
  XNOR U4681 ( .A(n3222), .B(n3221), .Z(c[608]) );
  XNOR U4682 ( .A(n3224), .B(n3223), .Z(c[609]) );
  XNOR U4683 ( .A(n3226), .B(n3225), .Z(c[60]) );
  XNOR U4684 ( .A(n3228), .B(n3227), .Z(c[610]) );
  XNOR U4685 ( .A(n3230), .B(n3229), .Z(c[611]) );
  XNOR U4686 ( .A(n3232), .B(n3231), .Z(c[612]) );
  XNOR U4687 ( .A(n3234), .B(n3233), .Z(c[613]) );
  XNOR U4688 ( .A(n3236), .B(n3235), .Z(c[614]) );
  XNOR U4689 ( .A(n3238), .B(n3237), .Z(c[615]) );
  XNOR U4690 ( .A(n3240), .B(n3239), .Z(c[616]) );
  XNOR U4691 ( .A(n3242), .B(n3241), .Z(c[617]) );
  XNOR U4692 ( .A(n3244), .B(n3243), .Z(c[618]) );
  XNOR U4693 ( .A(n3246), .B(n3245), .Z(c[619]) );
  XNOR U4694 ( .A(n3248), .B(n3247), .Z(c[61]) );
  XNOR U4695 ( .A(n3250), .B(n3249), .Z(c[620]) );
  XNOR U4696 ( .A(n3252), .B(n3251), .Z(c[621]) );
  XNOR U4697 ( .A(n3254), .B(n3253), .Z(c[622]) );
  XNOR U4698 ( .A(n3256), .B(n3255), .Z(c[623]) );
  XNOR U4699 ( .A(n3258), .B(n3257), .Z(c[624]) );
  XNOR U4700 ( .A(n3260), .B(n3259), .Z(c[625]) );
  XNOR U4701 ( .A(n3262), .B(n3261), .Z(c[626]) );
  XNOR U4702 ( .A(n3264), .B(n3263), .Z(c[627]) );
  XNOR U4703 ( .A(n3266), .B(n3265), .Z(c[628]) );
  XNOR U4704 ( .A(n3268), .B(n3267), .Z(c[629]) );
  XNOR U4705 ( .A(n3270), .B(n3269), .Z(c[62]) );
  XNOR U4706 ( .A(n3272), .B(n3271), .Z(c[630]) );
  XNOR U4707 ( .A(n3274), .B(n3273), .Z(c[631]) );
  XNOR U4708 ( .A(n3276), .B(n3275), .Z(c[632]) );
  XNOR U4709 ( .A(n3278), .B(n3277), .Z(c[633]) );
  XNOR U4710 ( .A(n3280), .B(n3279), .Z(c[634]) );
  XNOR U4711 ( .A(n3282), .B(n3281), .Z(c[635]) );
  XNOR U4712 ( .A(n3284), .B(n3283), .Z(c[636]) );
  XNOR U4713 ( .A(n3286), .B(n3285), .Z(c[637]) );
  XNOR U4714 ( .A(n3288), .B(n3287), .Z(c[638]) );
  XNOR U4715 ( .A(n3290), .B(n3289), .Z(c[639]) );
  XNOR U4716 ( .A(n3292), .B(n3291), .Z(c[63]) );
  XNOR U4717 ( .A(n3294), .B(n3293), .Z(c[640]) );
  XNOR U4718 ( .A(n3296), .B(n3295), .Z(c[641]) );
  XNOR U4719 ( .A(n3298), .B(n3297), .Z(c[642]) );
  XNOR U4720 ( .A(n3300), .B(n3299), .Z(c[643]) );
  XNOR U4721 ( .A(n3302), .B(n3301), .Z(c[644]) );
  XNOR U4722 ( .A(n3304), .B(n3303), .Z(c[645]) );
  XNOR U4723 ( .A(n3306), .B(n3305), .Z(c[646]) );
  XNOR U4724 ( .A(n3308), .B(n3307), .Z(c[647]) );
  XNOR U4725 ( .A(n3310), .B(n3309), .Z(c[648]) );
  XNOR U4726 ( .A(n3312), .B(n3311), .Z(c[649]) );
  XNOR U4727 ( .A(n3314), .B(n3313), .Z(c[64]) );
  XNOR U4728 ( .A(n3316), .B(n3315), .Z(c[650]) );
  XNOR U4729 ( .A(n3318), .B(n3317), .Z(c[651]) );
  XNOR U4730 ( .A(n3320), .B(n3319), .Z(c[652]) );
  XNOR U4731 ( .A(n3322), .B(n3321), .Z(c[653]) );
  XNOR U4732 ( .A(n3324), .B(n3323), .Z(c[654]) );
  XNOR U4733 ( .A(n3326), .B(n3325), .Z(c[655]) );
  XNOR U4734 ( .A(n3328), .B(n3327), .Z(c[656]) );
  XNOR U4735 ( .A(n3330), .B(n3329), .Z(c[657]) );
  XNOR U4736 ( .A(n3332), .B(n3331), .Z(c[658]) );
  XNOR U4737 ( .A(n3334), .B(n3333), .Z(c[659]) );
  XNOR U4738 ( .A(n3336), .B(n3335), .Z(c[65]) );
  XNOR U4739 ( .A(n3338), .B(n3337), .Z(c[660]) );
  XNOR U4740 ( .A(n3340), .B(n3339), .Z(c[661]) );
  XNOR U4741 ( .A(n3342), .B(n3341), .Z(c[662]) );
  XNOR U4742 ( .A(n3344), .B(n3343), .Z(c[663]) );
  XNOR U4743 ( .A(n3346), .B(n3345), .Z(c[664]) );
  XNOR U4744 ( .A(n3348), .B(n3347), .Z(c[665]) );
  XNOR U4745 ( .A(n3350), .B(n3349), .Z(c[666]) );
  XNOR U4746 ( .A(n3352), .B(n3351), .Z(c[667]) );
  XNOR U4747 ( .A(n3354), .B(n3353), .Z(c[668]) );
  XNOR U4748 ( .A(n3356), .B(n3355), .Z(c[669]) );
  XNOR U4749 ( .A(n3358), .B(n3357), .Z(c[66]) );
  XNOR U4750 ( .A(n3360), .B(n3359), .Z(c[670]) );
  XNOR U4751 ( .A(n3362), .B(n3361), .Z(c[671]) );
  XNOR U4752 ( .A(n3364), .B(n3363), .Z(c[672]) );
  XNOR U4753 ( .A(n3366), .B(n3365), .Z(c[673]) );
  XNOR U4754 ( .A(n3368), .B(n3367), .Z(c[674]) );
  XNOR U4755 ( .A(n3370), .B(n3369), .Z(c[675]) );
  XNOR U4756 ( .A(n3372), .B(n3371), .Z(c[676]) );
  XNOR U4757 ( .A(n3374), .B(n3373), .Z(c[677]) );
  XNOR U4758 ( .A(n3376), .B(n3375), .Z(c[678]) );
  XNOR U4759 ( .A(n3378), .B(n3377), .Z(c[679]) );
  XNOR U4760 ( .A(n3380), .B(n3379), .Z(c[67]) );
  XNOR U4761 ( .A(n3382), .B(n3381), .Z(c[680]) );
  XNOR U4762 ( .A(n3384), .B(n3383), .Z(c[681]) );
  XNOR U4763 ( .A(n3386), .B(n3385), .Z(c[682]) );
  XNOR U4764 ( .A(n3388), .B(n3387), .Z(c[683]) );
  XNOR U4765 ( .A(n3390), .B(n3389), .Z(c[684]) );
  XNOR U4766 ( .A(n3392), .B(n3391), .Z(c[685]) );
  XNOR U4767 ( .A(n3394), .B(n3393), .Z(c[686]) );
  XNOR U4768 ( .A(n3396), .B(n3395), .Z(c[687]) );
  XNOR U4769 ( .A(n3398), .B(n3397), .Z(c[688]) );
  XNOR U4770 ( .A(n3400), .B(n3399), .Z(c[689]) );
  XNOR U4771 ( .A(n3402), .B(n3401), .Z(c[68]) );
  XNOR U4772 ( .A(n3404), .B(n3403), .Z(c[690]) );
  XNOR U4773 ( .A(n3406), .B(n3405), .Z(c[691]) );
  XNOR U4774 ( .A(n3408), .B(n3407), .Z(c[692]) );
  XNOR U4775 ( .A(n3410), .B(n3409), .Z(c[693]) );
  XNOR U4776 ( .A(n3412), .B(n3411), .Z(c[694]) );
  XNOR U4777 ( .A(n3414), .B(n3413), .Z(c[695]) );
  XNOR U4778 ( .A(n3416), .B(n3415), .Z(c[696]) );
  XNOR U4779 ( .A(n3418), .B(n3417), .Z(c[697]) );
  XNOR U4780 ( .A(n3420), .B(n3419), .Z(c[698]) );
  XNOR U4781 ( .A(n3422), .B(n3421), .Z(c[699]) );
  XNOR U4782 ( .A(n3424), .B(n3423), .Z(c[69]) );
  XNOR U4783 ( .A(n3426), .B(n3425), .Z(c[6]) );
  XNOR U4784 ( .A(n3428), .B(n3427), .Z(c[700]) );
  XNOR U4785 ( .A(n3430), .B(n3429), .Z(c[701]) );
  XNOR U4786 ( .A(n3432), .B(n3431), .Z(c[702]) );
  XNOR U4787 ( .A(n3434), .B(n3433), .Z(c[703]) );
  XNOR U4788 ( .A(n3436), .B(n3435), .Z(c[704]) );
  XNOR U4789 ( .A(n3438), .B(n3437), .Z(c[705]) );
  XNOR U4790 ( .A(n3440), .B(n3439), .Z(c[706]) );
  XNOR U4791 ( .A(n3442), .B(n3441), .Z(c[707]) );
  XNOR U4792 ( .A(n3444), .B(n3443), .Z(c[708]) );
  XNOR U4793 ( .A(n3446), .B(n3445), .Z(c[709]) );
  XNOR U4794 ( .A(n3448), .B(n3447), .Z(c[70]) );
  XNOR U4795 ( .A(n3450), .B(n3449), .Z(c[710]) );
  XNOR U4796 ( .A(n3452), .B(n3451), .Z(c[711]) );
  XNOR U4797 ( .A(n3454), .B(n3453), .Z(c[712]) );
  XNOR U4798 ( .A(n3456), .B(n3455), .Z(c[713]) );
  XNOR U4799 ( .A(n3458), .B(n3457), .Z(c[714]) );
  XNOR U4800 ( .A(n3460), .B(n3459), .Z(c[715]) );
  XNOR U4801 ( .A(n3462), .B(n3461), .Z(c[716]) );
  XNOR U4802 ( .A(n3464), .B(n3463), .Z(c[717]) );
  XNOR U4803 ( .A(n3466), .B(n3465), .Z(c[718]) );
  XNOR U4804 ( .A(n3468), .B(n3467), .Z(c[719]) );
  XNOR U4805 ( .A(n3470), .B(n3469), .Z(c[71]) );
  XNOR U4806 ( .A(n3472), .B(n3471), .Z(c[720]) );
  XNOR U4807 ( .A(n3474), .B(n3473), .Z(c[721]) );
  XNOR U4808 ( .A(n3476), .B(n3475), .Z(c[722]) );
  XNOR U4809 ( .A(n3478), .B(n3477), .Z(c[723]) );
  XNOR U4810 ( .A(n3480), .B(n3479), .Z(c[724]) );
  XNOR U4811 ( .A(n3482), .B(n3481), .Z(c[725]) );
  XNOR U4812 ( .A(n3484), .B(n3483), .Z(c[726]) );
  XNOR U4813 ( .A(n3486), .B(n3485), .Z(c[727]) );
  XNOR U4814 ( .A(n3488), .B(n3487), .Z(c[728]) );
  XNOR U4815 ( .A(n3490), .B(n3489), .Z(c[729]) );
  XNOR U4816 ( .A(n3492), .B(n3491), .Z(c[72]) );
  XNOR U4817 ( .A(n3494), .B(n3493), .Z(c[730]) );
  XNOR U4818 ( .A(n3496), .B(n3495), .Z(c[731]) );
  XNOR U4819 ( .A(n3498), .B(n3497), .Z(c[732]) );
  XNOR U4820 ( .A(n3500), .B(n3499), .Z(c[733]) );
  XNOR U4821 ( .A(n3502), .B(n3501), .Z(c[734]) );
  XNOR U4822 ( .A(n3504), .B(n3503), .Z(c[735]) );
  XNOR U4823 ( .A(n3506), .B(n3505), .Z(c[736]) );
  XNOR U4824 ( .A(n3508), .B(n3507), .Z(c[737]) );
  XNOR U4825 ( .A(n3510), .B(n3509), .Z(c[738]) );
  XNOR U4826 ( .A(n3512), .B(n3511), .Z(c[739]) );
  XNOR U4827 ( .A(n3514), .B(n3513), .Z(c[73]) );
  XNOR U4828 ( .A(n3516), .B(n3515), .Z(c[740]) );
  XNOR U4829 ( .A(n3518), .B(n3517), .Z(c[741]) );
  XNOR U4830 ( .A(n3520), .B(n3519), .Z(c[742]) );
  XNOR U4831 ( .A(n3522), .B(n3521), .Z(c[743]) );
  XNOR U4832 ( .A(n3524), .B(n3523), .Z(c[744]) );
  XNOR U4833 ( .A(n3526), .B(n3525), .Z(c[745]) );
  XNOR U4834 ( .A(n3528), .B(n3527), .Z(c[746]) );
  XNOR U4835 ( .A(n3530), .B(n3529), .Z(c[747]) );
  XNOR U4836 ( .A(n3532), .B(n3531), .Z(c[748]) );
  XNOR U4837 ( .A(n3534), .B(n3533), .Z(c[749]) );
  XNOR U4838 ( .A(n3536), .B(n3535), .Z(c[74]) );
  XNOR U4839 ( .A(n3538), .B(n3537), .Z(c[750]) );
  XNOR U4840 ( .A(n3540), .B(n3539), .Z(c[751]) );
  XNOR U4841 ( .A(n3542), .B(n3541), .Z(c[752]) );
  XNOR U4842 ( .A(n3544), .B(n3543), .Z(c[753]) );
  XNOR U4843 ( .A(n3546), .B(n3545), .Z(c[754]) );
  XNOR U4844 ( .A(n3548), .B(n3547), .Z(c[755]) );
  XNOR U4845 ( .A(n3550), .B(n3549), .Z(c[756]) );
  XNOR U4846 ( .A(n3552), .B(n3551), .Z(c[757]) );
  XNOR U4847 ( .A(n3554), .B(n3553), .Z(c[758]) );
  XNOR U4848 ( .A(n3556), .B(n3555), .Z(c[759]) );
  XNOR U4849 ( .A(n3558), .B(n3557), .Z(c[75]) );
  XNOR U4850 ( .A(n3560), .B(n3559), .Z(c[760]) );
  XNOR U4851 ( .A(n3562), .B(n3561), .Z(c[761]) );
  XNOR U4852 ( .A(n3564), .B(n3563), .Z(c[762]) );
  XNOR U4853 ( .A(n3566), .B(n3565), .Z(c[763]) );
  XNOR U4854 ( .A(n3568), .B(n3567), .Z(c[764]) );
  XNOR U4855 ( .A(n3570), .B(n3569), .Z(c[765]) );
  XNOR U4856 ( .A(n3572), .B(n3571), .Z(c[766]) );
  XNOR U4857 ( .A(n3574), .B(n3573), .Z(c[767]) );
  XNOR U4858 ( .A(n3576), .B(n3575), .Z(c[768]) );
  XNOR U4859 ( .A(n3578), .B(n3577), .Z(c[769]) );
  XNOR U4860 ( .A(n3580), .B(n3579), .Z(c[76]) );
  XNOR U4861 ( .A(n3582), .B(n3581), .Z(c[770]) );
  XNOR U4862 ( .A(n3584), .B(n3583), .Z(c[771]) );
  XNOR U4863 ( .A(n3586), .B(n3585), .Z(c[772]) );
  XNOR U4864 ( .A(n3588), .B(n3587), .Z(c[773]) );
  XNOR U4865 ( .A(n3590), .B(n3589), .Z(c[774]) );
  XNOR U4866 ( .A(n3592), .B(n3591), .Z(c[775]) );
  XNOR U4867 ( .A(n3594), .B(n3593), .Z(c[776]) );
  XNOR U4868 ( .A(n3596), .B(n3595), .Z(c[777]) );
  XNOR U4869 ( .A(n3598), .B(n3597), .Z(c[778]) );
  XNOR U4870 ( .A(n3600), .B(n3599), .Z(c[779]) );
  XNOR U4871 ( .A(n3602), .B(n3601), .Z(c[77]) );
  XNOR U4872 ( .A(n3604), .B(n3603), .Z(c[780]) );
  XNOR U4873 ( .A(n3606), .B(n3605), .Z(c[781]) );
  XNOR U4874 ( .A(n3608), .B(n3607), .Z(c[782]) );
  XNOR U4875 ( .A(n3610), .B(n3609), .Z(c[783]) );
  XNOR U4876 ( .A(n3612), .B(n3611), .Z(c[784]) );
  XNOR U4877 ( .A(n3614), .B(n3613), .Z(c[785]) );
  XNOR U4878 ( .A(n3616), .B(n3615), .Z(c[786]) );
  XNOR U4879 ( .A(n3618), .B(n3617), .Z(c[787]) );
  XNOR U4880 ( .A(n3620), .B(n3619), .Z(c[788]) );
  XNOR U4881 ( .A(n3622), .B(n3621), .Z(c[789]) );
  XNOR U4882 ( .A(n3624), .B(n3623), .Z(c[78]) );
  XNOR U4883 ( .A(n3626), .B(n3625), .Z(c[790]) );
  XNOR U4884 ( .A(n3628), .B(n3627), .Z(c[791]) );
  XNOR U4885 ( .A(n3630), .B(n3629), .Z(c[792]) );
  XNOR U4886 ( .A(n3632), .B(n3631), .Z(c[793]) );
  XNOR U4887 ( .A(n3634), .B(n3633), .Z(c[794]) );
  XNOR U4888 ( .A(n3636), .B(n3635), .Z(c[795]) );
  XNOR U4889 ( .A(n3638), .B(n3637), .Z(c[796]) );
  XNOR U4890 ( .A(n3640), .B(n3639), .Z(c[797]) );
  XNOR U4891 ( .A(n3642), .B(n3641), .Z(c[798]) );
  XNOR U4892 ( .A(n3644), .B(n3643), .Z(c[799]) );
  XNOR U4893 ( .A(n3646), .B(n3645), .Z(c[79]) );
  XNOR U4894 ( .A(n3648), .B(n3647), .Z(c[7]) );
  XNOR U4895 ( .A(n3650), .B(n3649), .Z(c[800]) );
  XNOR U4896 ( .A(n3652), .B(n3651), .Z(c[801]) );
  XNOR U4897 ( .A(n3654), .B(n3653), .Z(c[802]) );
  XNOR U4898 ( .A(n3656), .B(n3655), .Z(c[803]) );
  XNOR U4899 ( .A(n3658), .B(n3657), .Z(c[804]) );
  XNOR U4900 ( .A(n3660), .B(n3659), .Z(c[805]) );
  XNOR U4901 ( .A(n3662), .B(n3661), .Z(c[806]) );
  XNOR U4902 ( .A(n3664), .B(n3663), .Z(c[807]) );
  XNOR U4903 ( .A(n3666), .B(n3665), .Z(c[808]) );
  XNOR U4904 ( .A(n3668), .B(n3667), .Z(c[809]) );
  XNOR U4905 ( .A(n3670), .B(n3669), .Z(c[80]) );
  XNOR U4906 ( .A(n3672), .B(n3671), .Z(c[810]) );
  XNOR U4907 ( .A(n3674), .B(n3673), .Z(c[811]) );
  XNOR U4908 ( .A(n3676), .B(n3675), .Z(c[812]) );
  XNOR U4909 ( .A(n3678), .B(n3677), .Z(c[813]) );
  XNOR U4910 ( .A(n3680), .B(n3679), .Z(c[814]) );
  XNOR U4911 ( .A(n3682), .B(n3681), .Z(c[815]) );
  XNOR U4912 ( .A(n3684), .B(n3683), .Z(c[816]) );
  XNOR U4913 ( .A(n3686), .B(n3685), .Z(c[817]) );
  XNOR U4914 ( .A(n3688), .B(n3687), .Z(c[818]) );
  XNOR U4915 ( .A(n3690), .B(n3689), .Z(c[819]) );
  XNOR U4916 ( .A(n3692), .B(n3691), .Z(c[81]) );
  XNOR U4917 ( .A(n3694), .B(n3693), .Z(c[820]) );
  XNOR U4918 ( .A(n3696), .B(n3695), .Z(c[821]) );
  XNOR U4919 ( .A(n3698), .B(n3697), .Z(c[822]) );
  XNOR U4920 ( .A(n3700), .B(n3699), .Z(c[823]) );
  XNOR U4921 ( .A(n3702), .B(n3701), .Z(c[824]) );
  XNOR U4922 ( .A(n3704), .B(n3703), .Z(c[825]) );
  XNOR U4923 ( .A(n3706), .B(n3705), .Z(c[826]) );
  XNOR U4924 ( .A(n3708), .B(n3707), .Z(c[827]) );
  XNOR U4925 ( .A(n3710), .B(n3709), .Z(c[828]) );
  XNOR U4926 ( .A(n3712), .B(n3711), .Z(c[829]) );
  XNOR U4927 ( .A(n3714), .B(n3713), .Z(c[82]) );
  XNOR U4928 ( .A(n3716), .B(n3715), .Z(c[830]) );
  XNOR U4929 ( .A(n3718), .B(n3717), .Z(c[831]) );
  XNOR U4930 ( .A(n3720), .B(n3719), .Z(c[832]) );
  XNOR U4931 ( .A(n3722), .B(n3721), .Z(c[833]) );
  XNOR U4932 ( .A(n3724), .B(n3723), .Z(c[834]) );
  XNOR U4933 ( .A(n3726), .B(n3725), .Z(c[835]) );
  XNOR U4934 ( .A(n3728), .B(n3727), .Z(c[836]) );
  XNOR U4935 ( .A(n3730), .B(n3729), .Z(c[837]) );
  XNOR U4936 ( .A(n3732), .B(n3731), .Z(c[838]) );
  XNOR U4937 ( .A(n3734), .B(n3733), .Z(c[839]) );
  XNOR U4938 ( .A(n3736), .B(n3735), .Z(c[83]) );
  XNOR U4939 ( .A(n3738), .B(n3737), .Z(c[840]) );
  XNOR U4940 ( .A(n3740), .B(n3739), .Z(c[841]) );
  XNOR U4941 ( .A(n3742), .B(n3741), .Z(c[842]) );
  XNOR U4942 ( .A(n3744), .B(n3743), .Z(c[843]) );
  XNOR U4943 ( .A(n3746), .B(n3745), .Z(c[844]) );
  XNOR U4944 ( .A(n3748), .B(n3747), .Z(c[845]) );
  XNOR U4945 ( .A(n3750), .B(n3749), .Z(c[846]) );
  XNOR U4946 ( .A(n3752), .B(n3751), .Z(c[847]) );
  XNOR U4947 ( .A(n3754), .B(n3753), .Z(c[848]) );
  XNOR U4948 ( .A(n3756), .B(n3755), .Z(c[849]) );
  XNOR U4949 ( .A(n3758), .B(n3757), .Z(c[84]) );
  XNOR U4950 ( .A(n3760), .B(n3759), .Z(c[850]) );
  XNOR U4951 ( .A(n3762), .B(n3761), .Z(c[851]) );
  XNOR U4952 ( .A(n3764), .B(n3763), .Z(c[852]) );
  XNOR U4953 ( .A(n3766), .B(n3765), .Z(c[853]) );
  XNOR U4954 ( .A(n3768), .B(n3767), .Z(c[854]) );
  XNOR U4955 ( .A(n3770), .B(n3769), .Z(c[855]) );
  XNOR U4956 ( .A(n3772), .B(n3771), .Z(c[856]) );
  XNOR U4957 ( .A(n3774), .B(n3773), .Z(c[857]) );
  XNOR U4958 ( .A(n3776), .B(n3775), .Z(c[858]) );
  XNOR U4959 ( .A(n3778), .B(n3777), .Z(c[859]) );
  XNOR U4960 ( .A(n3780), .B(n3779), .Z(c[85]) );
  XNOR U4961 ( .A(n3782), .B(n3781), .Z(c[860]) );
  XNOR U4962 ( .A(n3784), .B(n3783), .Z(c[861]) );
  XNOR U4963 ( .A(n3786), .B(n3785), .Z(c[862]) );
  XNOR U4964 ( .A(n3788), .B(n3787), .Z(c[863]) );
  XNOR U4965 ( .A(n3790), .B(n3789), .Z(c[864]) );
  XNOR U4966 ( .A(n3792), .B(n3791), .Z(c[865]) );
  XNOR U4967 ( .A(n3794), .B(n3793), .Z(c[866]) );
  XNOR U4968 ( .A(n3796), .B(n3795), .Z(c[867]) );
  XNOR U4969 ( .A(n3798), .B(n3797), .Z(c[868]) );
  XNOR U4970 ( .A(n3800), .B(n3799), .Z(c[869]) );
  XNOR U4971 ( .A(n3802), .B(n3801), .Z(c[86]) );
  XNOR U4972 ( .A(n3804), .B(n3803), .Z(c[870]) );
  XNOR U4973 ( .A(n3806), .B(n3805), .Z(c[871]) );
  XNOR U4974 ( .A(n3808), .B(n3807), .Z(c[872]) );
  XNOR U4975 ( .A(n3810), .B(n3809), .Z(c[873]) );
  XNOR U4976 ( .A(n3812), .B(n3811), .Z(c[874]) );
  XNOR U4977 ( .A(n3814), .B(n3813), .Z(c[875]) );
  XNOR U4978 ( .A(n3816), .B(n3815), .Z(c[876]) );
  XNOR U4979 ( .A(n3818), .B(n3817), .Z(c[877]) );
  XNOR U4980 ( .A(n3820), .B(n3819), .Z(c[878]) );
  XNOR U4981 ( .A(n3822), .B(n3821), .Z(c[879]) );
  XNOR U4982 ( .A(n3824), .B(n3823), .Z(c[87]) );
  XNOR U4983 ( .A(n3826), .B(n3825), .Z(c[880]) );
  XNOR U4984 ( .A(n3828), .B(n3827), .Z(c[881]) );
  XNOR U4985 ( .A(n3830), .B(n3829), .Z(c[882]) );
  XNOR U4986 ( .A(n3832), .B(n3831), .Z(c[883]) );
  XNOR U4987 ( .A(n3834), .B(n3833), .Z(c[884]) );
  XNOR U4988 ( .A(n3836), .B(n3835), .Z(c[885]) );
  XNOR U4989 ( .A(n3838), .B(n3837), .Z(c[886]) );
  XNOR U4990 ( .A(n3840), .B(n3839), .Z(c[887]) );
  XNOR U4991 ( .A(n3842), .B(n3841), .Z(c[888]) );
  XNOR U4992 ( .A(n3844), .B(n3843), .Z(c[889]) );
  XNOR U4993 ( .A(n3846), .B(n3845), .Z(c[88]) );
  XNOR U4994 ( .A(n3848), .B(n3847), .Z(c[890]) );
  XNOR U4995 ( .A(n3850), .B(n3849), .Z(c[891]) );
  XNOR U4996 ( .A(n3852), .B(n3851), .Z(c[892]) );
  XNOR U4997 ( .A(n3854), .B(n3853), .Z(c[893]) );
  XNOR U4998 ( .A(n3856), .B(n3855), .Z(c[894]) );
  XNOR U4999 ( .A(n3858), .B(n3857), .Z(c[895]) );
  XNOR U5000 ( .A(n3860), .B(n3859), .Z(c[896]) );
  XNOR U5001 ( .A(n3862), .B(n3861), .Z(c[897]) );
  XNOR U5002 ( .A(n3864), .B(n3863), .Z(c[898]) );
  XNOR U5003 ( .A(n3866), .B(n3865), .Z(c[899]) );
  XNOR U5004 ( .A(n3868), .B(n3867), .Z(c[89]) );
  XNOR U5005 ( .A(n3870), .B(n3869), .Z(c[8]) );
  XNOR U5006 ( .A(n3872), .B(n3871), .Z(c[900]) );
  XNOR U5007 ( .A(n3874), .B(n3873), .Z(c[901]) );
  XNOR U5008 ( .A(n3876), .B(n3875), .Z(c[902]) );
  XNOR U5009 ( .A(n3878), .B(n3877), .Z(c[903]) );
  XNOR U5010 ( .A(n3880), .B(n3879), .Z(c[904]) );
  XNOR U5011 ( .A(n3882), .B(n3881), .Z(c[905]) );
  XNOR U5012 ( .A(n3884), .B(n3883), .Z(c[906]) );
  XNOR U5013 ( .A(n3886), .B(n3885), .Z(c[907]) );
  XNOR U5014 ( .A(n3888), .B(n3887), .Z(c[908]) );
  XNOR U5015 ( .A(n3890), .B(n3889), .Z(c[909]) );
  XNOR U5016 ( .A(n3892), .B(n3891), .Z(c[90]) );
  XNOR U5017 ( .A(n3894), .B(n3893), .Z(c[910]) );
  XNOR U5018 ( .A(n3896), .B(n3895), .Z(c[911]) );
  XNOR U5019 ( .A(n3898), .B(n3897), .Z(c[912]) );
  XNOR U5020 ( .A(n3900), .B(n3899), .Z(c[913]) );
  XNOR U5021 ( .A(n3902), .B(n3901), .Z(c[914]) );
  XNOR U5022 ( .A(n3904), .B(n3903), .Z(c[915]) );
  XNOR U5023 ( .A(n3906), .B(n3905), .Z(c[916]) );
  XNOR U5024 ( .A(n3908), .B(n3907), .Z(c[917]) );
  XNOR U5025 ( .A(n3910), .B(n3909), .Z(c[918]) );
  XNOR U5026 ( .A(n3912), .B(n3911), .Z(c[919]) );
  XNOR U5027 ( .A(n3914), .B(n3913), .Z(c[91]) );
  XNOR U5028 ( .A(n3916), .B(n3915), .Z(c[920]) );
  XNOR U5029 ( .A(n3918), .B(n3917), .Z(c[921]) );
  XNOR U5030 ( .A(n3920), .B(n3919), .Z(c[922]) );
  XNOR U5031 ( .A(n3922), .B(n3921), .Z(c[923]) );
  XNOR U5032 ( .A(n3924), .B(n3923), .Z(c[924]) );
  XNOR U5033 ( .A(n3926), .B(n3925), .Z(c[925]) );
  XNOR U5034 ( .A(n3928), .B(n3927), .Z(c[926]) );
  XNOR U5035 ( .A(n3930), .B(n3929), .Z(c[927]) );
  XNOR U5036 ( .A(n3932), .B(n3931), .Z(c[928]) );
  XNOR U5037 ( .A(n3934), .B(n3933), .Z(c[929]) );
  XNOR U5038 ( .A(n3936), .B(n3935), .Z(c[92]) );
  XNOR U5039 ( .A(n3938), .B(n3937), .Z(c[930]) );
  XNOR U5040 ( .A(n3940), .B(n3939), .Z(c[931]) );
  XNOR U5041 ( .A(n3942), .B(n3941), .Z(c[932]) );
  XNOR U5042 ( .A(n3944), .B(n3943), .Z(c[933]) );
  XNOR U5043 ( .A(n3946), .B(n3945), .Z(c[934]) );
  XNOR U5044 ( .A(n3948), .B(n3947), .Z(c[935]) );
  XNOR U5045 ( .A(n3950), .B(n3949), .Z(c[936]) );
  XNOR U5046 ( .A(n3952), .B(n3951), .Z(c[937]) );
  XNOR U5047 ( .A(n3954), .B(n3953), .Z(c[938]) );
  XNOR U5048 ( .A(n3956), .B(n3955), .Z(c[939]) );
  XNOR U5049 ( .A(n3958), .B(n3957), .Z(c[93]) );
  XNOR U5050 ( .A(n3960), .B(n3959), .Z(c[940]) );
  XNOR U5051 ( .A(n3962), .B(n3961), .Z(c[941]) );
  XNOR U5052 ( .A(n3964), .B(n3963), .Z(c[942]) );
  XNOR U5053 ( .A(n3966), .B(n3965), .Z(c[943]) );
  XNOR U5054 ( .A(n3968), .B(n3967), .Z(c[944]) );
  XNOR U5055 ( .A(n3970), .B(n3969), .Z(c[945]) );
  XNOR U5056 ( .A(n3972), .B(n3971), .Z(c[946]) );
  XNOR U5057 ( .A(n3974), .B(n3973), .Z(c[947]) );
  XNOR U5058 ( .A(n3976), .B(n3975), .Z(c[948]) );
  XNOR U5059 ( .A(n3978), .B(n3977), .Z(c[949]) );
  XNOR U5060 ( .A(n3980), .B(n3979), .Z(c[94]) );
  XNOR U5061 ( .A(n3982), .B(n3981), .Z(c[950]) );
  XNOR U5062 ( .A(n3984), .B(n3983), .Z(c[951]) );
  XNOR U5063 ( .A(n3986), .B(n3985), .Z(c[952]) );
  XNOR U5064 ( .A(n3988), .B(n3987), .Z(c[953]) );
  XNOR U5065 ( .A(n3990), .B(n3989), .Z(c[954]) );
  XNOR U5066 ( .A(n3992), .B(n3991), .Z(c[955]) );
  XNOR U5067 ( .A(n3994), .B(n3993), .Z(c[956]) );
  XNOR U5068 ( .A(n3996), .B(n3995), .Z(c[957]) );
  XNOR U5069 ( .A(n3998), .B(n3997), .Z(c[958]) );
  XNOR U5070 ( .A(n4000), .B(n3999), .Z(c[959]) );
  XNOR U5071 ( .A(n4002), .B(n4001), .Z(c[95]) );
  XNOR U5072 ( .A(n4004), .B(n4003), .Z(c[960]) );
  XNOR U5073 ( .A(n4006), .B(n4005), .Z(c[961]) );
  XNOR U5074 ( .A(n4008), .B(n4007), .Z(c[962]) );
  XNOR U5075 ( .A(n4010), .B(n4009), .Z(c[963]) );
  XNOR U5076 ( .A(n4012), .B(n4011), .Z(c[964]) );
  XNOR U5077 ( .A(n4014), .B(n4013), .Z(c[965]) );
  XNOR U5078 ( .A(n4016), .B(n4015), .Z(c[966]) );
  XNOR U5079 ( .A(n4018), .B(n4017), .Z(c[967]) );
  XNOR U5080 ( .A(n4020), .B(n4019), .Z(c[968]) );
  XNOR U5081 ( .A(n4022), .B(n4021), .Z(c[969]) );
  XNOR U5082 ( .A(n4024), .B(n4023), .Z(c[96]) );
  XNOR U5083 ( .A(n4026), .B(n4025), .Z(c[970]) );
  XNOR U5084 ( .A(n4028), .B(n4027), .Z(c[971]) );
  XNOR U5085 ( .A(n4030), .B(n4029), .Z(c[972]) );
  XNOR U5086 ( .A(n4032), .B(n4031), .Z(c[973]) );
  XNOR U5087 ( .A(n4034), .B(n4033), .Z(c[974]) );
  XNOR U5088 ( .A(n4036), .B(n4035), .Z(c[975]) );
  XNOR U5089 ( .A(n4038), .B(n4037), .Z(c[976]) );
  XNOR U5090 ( .A(n4040), .B(n4039), .Z(c[977]) );
  XNOR U5091 ( .A(n4042), .B(n4041), .Z(c[978]) );
  XNOR U5092 ( .A(n4044), .B(n4043), .Z(c[979]) );
  XNOR U5093 ( .A(n4046), .B(n4045), .Z(c[97]) );
  XNOR U5094 ( .A(n4048), .B(n4047), .Z(c[980]) );
  XNOR U5095 ( .A(n4050), .B(n4049), .Z(c[981]) );
  XNOR U5096 ( .A(n4052), .B(n4051), .Z(c[982]) );
  XNOR U5097 ( .A(n4054), .B(n4053), .Z(c[983]) );
  XNOR U5098 ( .A(n4056), .B(n4055), .Z(c[984]) );
  XNOR U5099 ( .A(n4058), .B(n4057), .Z(c[985]) );
  XNOR U5100 ( .A(n4060), .B(n4059), .Z(c[986]) );
  XNOR U5101 ( .A(n4062), .B(n4061), .Z(c[987]) );
  XNOR U5102 ( .A(n4064), .B(n4063), .Z(c[988]) );
  XNOR U5103 ( .A(n4066), .B(n4065), .Z(c[989]) );
  XNOR U5104 ( .A(n4068), .B(n4067), .Z(c[98]) );
  XNOR U5105 ( .A(n4070), .B(n4069), .Z(c[990]) );
  XNOR U5106 ( .A(n4072), .B(n4071), .Z(c[991]) );
  XNOR U5107 ( .A(n4074), .B(n4073), .Z(c[992]) );
  XNOR U5108 ( .A(n4076), .B(n4075), .Z(c[993]) );
  XNOR U5109 ( .A(n4078), .B(n4077), .Z(c[994]) );
  XNOR U5110 ( .A(n4080), .B(n4079), .Z(c[995]) );
  XNOR U5111 ( .A(n4082), .B(n4081), .Z(c[996]) );
  XNOR U5112 ( .A(n4084), .B(n4083), .Z(c[997]) );
  XNOR U5113 ( .A(n4086), .B(n4085), .Z(c[998]) );
  XNOR U5114 ( .A(n4088), .B(n4087), .Z(c[999]) );
  XNOR U5115 ( .A(n4090), .B(n4089), .Z(c[99]) );
  XNOR U5116 ( .A(n4092), .B(n4091), .Z(c[9]) );
endmodule

