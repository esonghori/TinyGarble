
module FA_0 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(A), .B(B), .Z(CO) );
  XOR U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_99 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_98 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_97 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_96 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_95 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_94 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_93 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_92 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_91 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_90 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_89 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_88 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_87 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_86 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_85 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_84 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_83 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_82 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_81 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_80 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_79 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_78 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_77 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_76 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_75 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_74 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_73 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_72 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_71 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_70 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_69 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_68 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_67 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_66 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_65 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_64 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_63 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_62 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_61 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_60 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_59 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_58 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_57 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_56 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_55 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_54 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_53 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_52 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_51 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_50 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_49 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_48 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_47 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_46 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_45 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_44 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_43 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_42 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_41 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_40 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_39 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_38 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_37 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_36 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_35 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_34 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_33 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_32 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_31 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_30 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_29 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_28 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_27 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_26 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_25 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_24 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_23 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_22 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_21 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_20 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_19 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_18 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_17 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_16 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_15 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_14 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_13 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_12 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_11 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_10 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_9 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_8 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_7 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_6 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_5 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_4 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_3 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_2 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  XOR U2 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_1 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N256 ( A, B, CI, S, CO );
  input [255:0] A;
  input [255:0] B;
  output [255:0] S;
  input CI;
  output CO;

  wire   [255:1] C;

  FA_0 \FAINST[0].FA_  ( .A(A[0]), .B(B[0]), .CI(1'b0), .S(S[0]), .CO(C[1]) );
  FA_255 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(C[1]), .S(S[1]), .CO(C[2])
         );
  FA_254 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_253 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_252 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_251 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_250 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_249 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_248 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_247 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10])
         );
  FA_246 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_245 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_244 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_243 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_242 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_241 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_240 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_239 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_238 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_237 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_236 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_235 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_234 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_233 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_232 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_231 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_230 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_229 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_228 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_227 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_226 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_225 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]), .CO(
        C[32]) );
  FA_224 \FAINST[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), .S(S[32]), .CO(
        C[33]) );
  FA_223 \FAINST[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), .S(S[33]), .CO(
        C[34]) );
  FA_222 \FAINST[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), .S(S[34]), .CO(
        C[35]) );
  FA_221 \FAINST[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), .S(S[35]), .CO(
        C[36]) );
  FA_220 \FAINST[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), .S(S[36]), .CO(
        C[37]) );
  FA_219 \FAINST[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), .S(S[37]), .CO(
        C[38]) );
  FA_218 \FAINST[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), .S(S[38]), .CO(
        C[39]) );
  FA_217 \FAINST[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), .S(S[39]), .CO(
        C[40]) );
  FA_216 \FAINST[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), .S(S[40]), .CO(
        C[41]) );
  FA_215 \FAINST[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), .S(S[41]), .CO(
        C[42]) );
  FA_214 \FAINST[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), .S(S[42]), .CO(
        C[43]) );
  FA_213 \FAINST[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), .S(S[43]), .CO(
        C[44]) );
  FA_212 \FAINST[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), .S(S[44]), .CO(
        C[45]) );
  FA_211 \FAINST[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), .S(S[45]), .CO(
        C[46]) );
  FA_210 \FAINST[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), .S(S[46]), .CO(
        C[47]) );
  FA_209 \FAINST[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), .S(S[47]), .CO(
        C[48]) );
  FA_208 \FAINST[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), .S(S[48]), .CO(
        C[49]) );
  FA_207 \FAINST[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), .S(S[49]), .CO(
        C[50]) );
  FA_206 \FAINST[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), .S(S[50]), .CO(
        C[51]) );
  FA_205 \FAINST[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), .S(S[51]), .CO(
        C[52]) );
  FA_204 \FAINST[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), .S(S[52]), .CO(
        C[53]) );
  FA_203 \FAINST[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), .S(S[53]), .CO(
        C[54]) );
  FA_202 \FAINST[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), .S(S[54]), .CO(
        C[55]) );
  FA_201 \FAINST[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), .S(S[55]), .CO(
        C[56]) );
  FA_200 \FAINST[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), .S(S[56]), .CO(
        C[57]) );
  FA_199 \FAINST[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), .S(S[57]), .CO(
        C[58]) );
  FA_198 \FAINST[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), .S(S[58]), .CO(
        C[59]) );
  FA_197 \FAINST[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), .S(S[59]), .CO(
        C[60]) );
  FA_196 \FAINST[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), .S(S[60]), .CO(
        C[61]) );
  FA_195 \FAINST[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), .S(S[61]), .CO(
        C[62]) );
  FA_194 \FAINST[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), .S(S[62]), .CO(
        C[63]) );
  FA_193 \FAINST[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), .S(S[63]), .CO(
        C[64]) );
  FA_192 \FAINST[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), .S(S[64]), .CO(
        C[65]) );
  FA_191 \FAINST[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), .S(S[65]), .CO(
        C[66]) );
  FA_190 \FAINST[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), .S(S[66]), .CO(
        C[67]) );
  FA_189 \FAINST[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), .S(S[67]), .CO(
        C[68]) );
  FA_188 \FAINST[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), .S(S[68]), .CO(
        C[69]) );
  FA_187 \FAINST[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), .S(S[69]), .CO(
        C[70]) );
  FA_186 \FAINST[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), .S(S[70]), .CO(
        C[71]) );
  FA_185 \FAINST[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), .S(S[71]), .CO(
        C[72]) );
  FA_184 \FAINST[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), .S(S[72]), .CO(
        C[73]) );
  FA_183 \FAINST[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), .S(S[73]), .CO(
        C[74]) );
  FA_182 \FAINST[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), .S(S[74]), .CO(
        C[75]) );
  FA_181 \FAINST[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), .S(S[75]), .CO(
        C[76]) );
  FA_180 \FAINST[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), .S(S[76]), .CO(
        C[77]) );
  FA_179 \FAINST[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), .S(S[77]), .CO(
        C[78]) );
  FA_178 \FAINST[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), .S(S[78]), .CO(
        C[79]) );
  FA_177 \FAINST[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), .S(S[79]), .CO(
        C[80]) );
  FA_176 \FAINST[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), .S(S[80]), .CO(
        C[81]) );
  FA_175 \FAINST[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), .S(S[81]), .CO(
        C[82]) );
  FA_174 \FAINST[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), .S(S[82]), .CO(
        C[83]) );
  FA_173 \FAINST[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), .S(S[83]), .CO(
        C[84]) );
  FA_172 \FAINST[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), .S(S[84]), .CO(
        C[85]) );
  FA_171 \FAINST[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), .S(S[85]), .CO(
        C[86]) );
  FA_170 \FAINST[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), .S(S[86]), .CO(
        C[87]) );
  FA_169 \FAINST[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), .S(S[87]), .CO(
        C[88]) );
  FA_168 \FAINST[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), .S(S[88]), .CO(
        C[89]) );
  FA_167 \FAINST[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), .S(S[89]), .CO(
        C[90]) );
  FA_166 \FAINST[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), .S(S[90]), .CO(
        C[91]) );
  FA_165 \FAINST[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), .S(S[91]), .CO(
        C[92]) );
  FA_164 \FAINST[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), .S(S[92]), .CO(
        C[93]) );
  FA_163 \FAINST[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), .S(S[93]), .CO(
        C[94]) );
  FA_162 \FAINST[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), .S(S[94]), .CO(
        C[95]) );
  FA_161 \FAINST[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), .S(S[95]), .CO(
        C[96]) );
  FA_160 \FAINST[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), .S(S[96]), .CO(
        C[97]) );
  FA_159 \FAINST[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), .S(S[97]), .CO(
        C[98]) );
  FA_158 \FAINST[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), .S(S[98]), .CO(
        C[99]) );
  FA_157 \FAINST[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), .S(S[99]), .CO(
        C[100]) );
  FA_156 \FAINST[100].FA_  ( .A(A[100]), .B(B[100]), .CI(C[100]), .S(S[100]), 
        .CO(C[101]) );
  FA_155 \FAINST[101].FA_  ( .A(A[101]), .B(B[101]), .CI(C[101]), .S(S[101]), 
        .CO(C[102]) );
  FA_154 \FAINST[102].FA_  ( .A(A[102]), .B(B[102]), .CI(C[102]), .S(S[102]), 
        .CO(C[103]) );
  FA_153 \FAINST[103].FA_  ( .A(A[103]), .B(B[103]), .CI(C[103]), .S(S[103]), 
        .CO(C[104]) );
  FA_152 \FAINST[104].FA_  ( .A(A[104]), .B(B[104]), .CI(C[104]), .S(S[104]), 
        .CO(C[105]) );
  FA_151 \FAINST[105].FA_  ( .A(A[105]), .B(B[105]), .CI(C[105]), .S(S[105]), 
        .CO(C[106]) );
  FA_150 \FAINST[106].FA_  ( .A(A[106]), .B(B[106]), .CI(C[106]), .S(S[106]), 
        .CO(C[107]) );
  FA_149 \FAINST[107].FA_  ( .A(A[107]), .B(B[107]), .CI(C[107]), .S(S[107]), 
        .CO(C[108]) );
  FA_148 \FAINST[108].FA_  ( .A(A[108]), .B(B[108]), .CI(C[108]), .S(S[108]), 
        .CO(C[109]) );
  FA_147 \FAINST[109].FA_  ( .A(A[109]), .B(B[109]), .CI(C[109]), .S(S[109]), 
        .CO(C[110]) );
  FA_146 \FAINST[110].FA_  ( .A(A[110]), .B(B[110]), .CI(C[110]), .S(S[110]), 
        .CO(C[111]) );
  FA_145 \FAINST[111].FA_  ( .A(A[111]), .B(B[111]), .CI(C[111]), .S(S[111]), 
        .CO(C[112]) );
  FA_144 \FAINST[112].FA_  ( .A(A[112]), .B(B[112]), .CI(C[112]), .S(S[112]), 
        .CO(C[113]) );
  FA_143 \FAINST[113].FA_  ( .A(A[113]), .B(B[113]), .CI(C[113]), .S(S[113]), 
        .CO(C[114]) );
  FA_142 \FAINST[114].FA_  ( .A(A[114]), .B(B[114]), .CI(C[114]), .S(S[114]), 
        .CO(C[115]) );
  FA_141 \FAINST[115].FA_  ( .A(A[115]), .B(B[115]), .CI(C[115]), .S(S[115]), 
        .CO(C[116]) );
  FA_140 \FAINST[116].FA_  ( .A(A[116]), .B(B[116]), .CI(C[116]), .S(S[116]), 
        .CO(C[117]) );
  FA_139 \FAINST[117].FA_  ( .A(A[117]), .B(B[117]), .CI(C[117]), .S(S[117]), 
        .CO(C[118]) );
  FA_138 \FAINST[118].FA_  ( .A(A[118]), .B(B[118]), .CI(C[118]), .S(S[118]), 
        .CO(C[119]) );
  FA_137 \FAINST[119].FA_  ( .A(A[119]), .B(B[119]), .CI(C[119]), .S(S[119]), 
        .CO(C[120]) );
  FA_136 \FAINST[120].FA_  ( .A(A[120]), .B(B[120]), .CI(C[120]), .S(S[120]), 
        .CO(C[121]) );
  FA_135 \FAINST[121].FA_  ( .A(A[121]), .B(B[121]), .CI(C[121]), .S(S[121]), 
        .CO(C[122]) );
  FA_134 \FAINST[122].FA_  ( .A(A[122]), .B(B[122]), .CI(C[122]), .S(S[122]), 
        .CO(C[123]) );
  FA_133 \FAINST[123].FA_  ( .A(A[123]), .B(B[123]), .CI(C[123]), .S(S[123]), 
        .CO(C[124]) );
  FA_132 \FAINST[124].FA_  ( .A(A[124]), .B(B[124]), .CI(C[124]), .S(S[124]), 
        .CO(C[125]) );
  FA_131 \FAINST[125].FA_  ( .A(A[125]), .B(B[125]), .CI(C[125]), .S(S[125]), 
        .CO(C[126]) );
  FA_130 \FAINST[126].FA_  ( .A(A[126]), .B(B[126]), .CI(C[126]), .S(S[126]), 
        .CO(C[127]) );
  FA_129 \FAINST[127].FA_  ( .A(A[127]), .B(B[127]), .CI(C[127]), .S(S[127]), 
        .CO(C[128]) );
  FA_128 \FAINST[128].FA_  ( .A(A[128]), .B(B[128]), .CI(C[128]), .S(S[128]), 
        .CO(C[129]) );
  FA_127 \FAINST[129].FA_  ( .A(A[129]), .B(B[129]), .CI(C[129]), .S(S[129]), 
        .CO(C[130]) );
  FA_126 \FAINST[130].FA_  ( .A(A[130]), .B(B[130]), .CI(C[130]), .S(S[130]), 
        .CO(C[131]) );
  FA_125 \FAINST[131].FA_  ( .A(A[131]), .B(B[131]), .CI(C[131]), .S(S[131]), 
        .CO(C[132]) );
  FA_124 \FAINST[132].FA_  ( .A(A[132]), .B(B[132]), .CI(C[132]), .S(S[132]), 
        .CO(C[133]) );
  FA_123 \FAINST[133].FA_  ( .A(A[133]), .B(B[133]), .CI(C[133]), .S(S[133]), 
        .CO(C[134]) );
  FA_122 \FAINST[134].FA_  ( .A(A[134]), .B(B[134]), .CI(C[134]), .S(S[134]), 
        .CO(C[135]) );
  FA_121 \FAINST[135].FA_  ( .A(A[135]), .B(B[135]), .CI(C[135]), .S(S[135]), 
        .CO(C[136]) );
  FA_120 \FAINST[136].FA_  ( .A(A[136]), .B(B[136]), .CI(C[136]), .S(S[136]), 
        .CO(C[137]) );
  FA_119 \FAINST[137].FA_  ( .A(A[137]), .B(B[137]), .CI(C[137]), .S(S[137]), 
        .CO(C[138]) );
  FA_118 \FAINST[138].FA_  ( .A(A[138]), .B(B[138]), .CI(C[138]), .S(S[138]), 
        .CO(C[139]) );
  FA_117 \FAINST[139].FA_  ( .A(A[139]), .B(B[139]), .CI(C[139]), .S(S[139]), 
        .CO(C[140]) );
  FA_116 \FAINST[140].FA_  ( .A(A[140]), .B(B[140]), .CI(C[140]), .S(S[140]), 
        .CO(C[141]) );
  FA_115 \FAINST[141].FA_  ( .A(A[141]), .B(B[141]), .CI(C[141]), .S(S[141]), 
        .CO(C[142]) );
  FA_114 \FAINST[142].FA_  ( .A(A[142]), .B(B[142]), .CI(C[142]), .S(S[142]), 
        .CO(C[143]) );
  FA_113 \FAINST[143].FA_  ( .A(A[143]), .B(B[143]), .CI(C[143]), .S(S[143]), 
        .CO(C[144]) );
  FA_112 \FAINST[144].FA_  ( .A(A[144]), .B(B[144]), .CI(C[144]), .S(S[144]), 
        .CO(C[145]) );
  FA_111 \FAINST[145].FA_  ( .A(A[145]), .B(B[145]), .CI(C[145]), .S(S[145]), 
        .CO(C[146]) );
  FA_110 \FAINST[146].FA_  ( .A(A[146]), .B(B[146]), .CI(C[146]), .S(S[146]), 
        .CO(C[147]) );
  FA_109 \FAINST[147].FA_  ( .A(A[147]), .B(B[147]), .CI(C[147]), .S(S[147]), 
        .CO(C[148]) );
  FA_108 \FAINST[148].FA_  ( .A(A[148]), .B(B[148]), .CI(C[148]), .S(S[148]), 
        .CO(C[149]) );
  FA_107 \FAINST[149].FA_  ( .A(A[149]), .B(B[149]), .CI(C[149]), .S(S[149]), 
        .CO(C[150]) );
  FA_106 \FAINST[150].FA_  ( .A(A[150]), .B(B[150]), .CI(C[150]), .S(S[150]), 
        .CO(C[151]) );
  FA_105 \FAINST[151].FA_  ( .A(A[151]), .B(B[151]), .CI(C[151]), .S(S[151]), 
        .CO(C[152]) );
  FA_104 \FAINST[152].FA_  ( .A(A[152]), .B(B[152]), .CI(C[152]), .S(S[152]), 
        .CO(C[153]) );
  FA_103 \FAINST[153].FA_  ( .A(A[153]), .B(B[153]), .CI(C[153]), .S(S[153]), 
        .CO(C[154]) );
  FA_102 \FAINST[154].FA_  ( .A(A[154]), .B(B[154]), .CI(C[154]), .S(S[154]), 
        .CO(C[155]) );
  FA_101 \FAINST[155].FA_  ( .A(A[155]), .B(B[155]), .CI(C[155]), .S(S[155]), 
        .CO(C[156]) );
  FA_100 \FAINST[156].FA_  ( .A(A[156]), .B(B[156]), .CI(C[156]), .S(S[156]), 
        .CO(C[157]) );
  FA_99 \FAINST[157].FA_  ( .A(A[157]), .B(B[157]), .CI(C[157]), .S(S[157]), 
        .CO(C[158]) );
  FA_98 \FAINST[158].FA_  ( .A(A[158]), .B(B[158]), .CI(C[158]), .S(S[158]), 
        .CO(C[159]) );
  FA_97 \FAINST[159].FA_  ( .A(A[159]), .B(B[159]), .CI(C[159]), .S(S[159]), 
        .CO(C[160]) );
  FA_96 \FAINST[160].FA_  ( .A(A[160]), .B(B[160]), .CI(C[160]), .S(S[160]), 
        .CO(C[161]) );
  FA_95 \FAINST[161].FA_  ( .A(A[161]), .B(B[161]), .CI(C[161]), .S(S[161]), 
        .CO(C[162]) );
  FA_94 \FAINST[162].FA_  ( .A(A[162]), .B(B[162]), .CI(C[162]), .S(S[162]), 
        .CO(C[163]) );
  FA_93 \FAINST[163].FA_  ( .A(A[163]), .B(B[163]), .CI(C[163]), .S(S[163]), 
        .CO(C[164]) );
  FA_92 \FAINST[164].FA_  ( .A(A[164]), .B(B[164]), .CI(C[164]), .S(S[164]), 
        .CO(C[165]) );
  FA_91 \FAINST[165].FA_  ( .A(A[165]), .B(B[165]), .CI(C[165]), .S(S[165]), 
        .CO(C[166]) );
  FA_90 \FAINST[166].FA_  ( .A(A[166]), .B(B[166]), .CI(C[166]), .S(S[166]), 
        .CO(C[167]) );
  FA_89 \FAINST[167].FA_  ( .A(A[167]), .B(B[167]), .CI(C[167]), .S(S[167]), 
        .CO(C[168]) );
  FA_88 \FAINST[168].FA_  ( .A(A[168]), .B(B[168]), .CI(C[168]), .S(S[168]), 
        .CO(C[169]) );
  FA_87 \FAINST[169].FA_  ( .A(A[169]), .B(B[169]), .CI(C[169]), .S(S[169]), 
        .CO(C[170]) );
  FA_86 \FAINST[170].FA_  ( .A(A[170]), .B(B[170]), .CI(C[170]), .S(S[170]), 
        .CO(C[171]) );
  FA_85 \FAINST[171].FA_  ( .A(A[171]), .B(B[171]), .CI(C[171]), .S(S[171]), 
        .CO(C[172]) );
  FA_84 \FAINST[172].FA_  ( .A(A[172]), .B(B[172]), .CI(C[172]), .S(S[172]), 
        .CO(C[173]) );
  FA_83 \FAINST[173].FA_  ( .A(A[173]), .B(B[173]), .CI(C[173]), .S(S[173]), 
        .CO(C[174]) );
  FA_82 \FAINST[174].FA_  ( .A(A[174]), .B(B[174]), .CI(C[174]), .S(S[174]), 
        .CO(C[175]) );
  FA_81 \FAINST[175].FA_  ( .A(A[175]), .B(B[175]), .CI(C[175]), .S(S[175]), 
        .CO(C[176]) );
  FA_80 \FAINST[176].FA_  ( .A(A[176]), .B(B[176]), .CI(C[176]), .S(S[176]), 
        .CO(C[177]) );
  FA_79 \FAINST[177].FA_  ( .A(A[177]), .B(B[177]), .CI(C[177]), .S(S[177]), 
        .CO(C[178]) );
  FA_78 \FAINST[178].FA_  ( .A(A[178]), .B(B[178]), .CI(C[178]), .S(S[178]), 
        .CO(C[179]) );
  FA_77 \FAINST[179].FA_  ( .A(A[179]), .B(B[179]), .CI(C[179]), .S(S[179]), 
        .CO(C[180]) );
  FA_76 \FAINST[180].FA_  ( .A(A[180]), .B(B[180]), .CI(C[180]), .S(S[180]), 
        .CO(C[181]) );
  FA_75 \FAINST[181].FA_  ( .A(A[181]), .B(B[181]), .CI(C[181]), .S(S[181]), 
        .CO(C[182]) );
  FA_74 \FAINST[182].FA_  ( .A(A[182]), .B(B[182]), .CI(C[182]), .S(S[182]), 
        .CO(C[183]) );
  FA_73 \FAINST[183].FA_  ( .A(A[183]), .B(B[183]), .CI(C[183]), .S(S[183]), 
        .CO(C[184]) );
  FA_72 \FAINST[184].FA_  ( .A(A[184]), .B(B[184]), .CI(C[184]), .S(S[184]), 
        .CO(C[185]) );
  FA_71 \FAINST[185].FA_  ( .A(A[185]), .B(B[185]), .CI(C[185]), .S(S[185]), 
        .CO(C[186]) );
  FA_70 \FAINST[186].FA_  ( .A(A[186]), .B(B[186]), .CI(C[186]), .S(S[186]), 
        .CO(C[187]) );
  FA_69 \FAINST[187].FA_  ( .A(A[187]), .B(B[187]), .CI(C[187]), .S(S[187]), 
        .CO(C[188]) );
  FA_68 \FAINST[188].FA_  ( .A(A[188]), .B(B[188]), .CI(C[188]), .S(S[188]), 
        .CO(C[189]) );
  FA_67 \FAINST[189].FA_  ( .A(A[189]), .B(B[189]), .CI(C[189]), .S(S[189]), 
        .CO(C[190]) );
  FA_66 \FAINST[190].FA_  ( .A(A[190]), .B(B[190]), .CI(C[190]), .S(S[190]), 
        .CO(C[191]) );
  FA_65 \FAINST[191].FA_  ( .A(A[191]), .B(B[191]), .CI(C[191]), .S(S[191]), 
        .CO(C[192]) );
  FA_64 \FAINST[192].FA_  ( .A(A[192]), .B(B[192]), .CI(C[192]), .S(S[192]), 
        .CO(C[193]) );
  FA_63 \FAINST[193].FA_  ( .A(A[193]), .B(B[193]), .CI(C[193]), .S(S[193]), 
        .CO(C[194]) );
  FA_62 \FAINST[194].FA_  ( .A(A[194]), .B(B[194]), .CI(C[194]), .S(S[194]), 
        .CO(C[195]) );
  FA_61 \FAINST[195].FA_  ( .A(A[195]), .B(B[195]), .CI(C[195]), .S(S[195]), 
        .CO(C[196]) );
  FA_60 \FAINST[196].FA_  ( .A(A[196]), .B(B[196]), .CI(C[196]), .S(S[196]), 
        .CO(C[197]) );
  FA_59 \FAINST[197].FA_  ( .A(A[197]), .B(B[197]), .CI(C[197]), .S(S[197]), 
        .CO(C[198]) );
  FA_58 \FAINST[198].FA_  ( .A(A[198]), .B(B[198]), .CI(C[198]), .S(S[198]), 
        .CO(C[199]) );
  FA_57 \FAINST[199].FA_  ( .A(A[199]), .B(B[199]), .CI(C[199]), .S(S[199]), 
        .CO(C[200]) );
  FA_56 \FAINST[200].FA_  ( .A(A[200]), .B(B[200]), .CI(C[200]), .S(S[200]), 
        .CO(C[201]) );
  FA_55 \FAINST[201].FA_  ( .A(A[201]), .B(B[201]), .CI(C[201]), .S(S[201]), 
        .CO(C[202]) );
  FA_54 \FAINST[202].FA_  ( .A(A[202]), .B(B[202]), .CI(C[202]), .S(S[202]), 
        .CO(C[203]) );
  FA_53 \FAINST[203].FA_  ( .A(A[203]), .B(B[203]), .CI(C[203]), .S(S[203]), 
        .CO(C[204]) );
  FA_52 \FAINST[204].FA_  ( .A(A[204]), .B(B[204]), .CI(C[204]), .S(S[204]), 
        .CO(C[205]) );
  FA_51 \FAINST[205].FA_  ( .A(A[205]), .B(B[205]), .CI(C[205]), .S(S[205]), 
        .CO(C[206]) );
  FA_50 \FAINST[206].FA_  ( .A(A[206]), .B(B[206]), .CI(C[206]), .S(S[206]), 
        .CO(C[207]) );
  FA_49 \FAINST[207].FA_  ( .A(A[207]), .B(B[207]), .CI(C[207]), .S(S[207]), 
        .CO(C[208]) );
  FA_48 \FAINST[208].FA_  ( .A(A[208]), .B(B[208]), .CI(C[208]), .S(S[208]), 
        .CO(C[209]) );
  FA_47 \FAINST[209].FA_  ( .A(A[209]), .B(B[209]), .CI(C[209]), .S(S[209]), 
        .CO(C[210]) );
  FA_46 \FAINST[210].FA_  ( .A(A[210]), .B(B[210]), .CI(C[210]), .S(S[210]), 
        .CO(C[211]) );
  FA_45 \FAINST[211].FA_  ( .A(A[211]), .B(B[211]), .CI(C[211]), .S(S[211]), 
        .CO(C[212]) );
  FA_44 \FAINST[212].FA_  ( .A(A[212]), .B(B[212]), .CI(C[212]), .S(S[212]), 
        .CO(C[213]) );
  FA_43 \FAINST[213].FA_  ( .A(A[213]), .B(B[213]), .CI(C[213]), .S(S[213]), 
        .CO(C[214]) );
  FA_42 \FAINST[214].FA_  ( .A(A[214]), .B(B[214]), .CI(C[214]), .S(S[214]), 
        .CO(C[215]) );
  FA_41 \FAINST[215].FA_  ( .A(A[215]), .B(B[215]), .CI(C[215]), .S(S[215]), 
        .CO(C[216]) );
  FA_40 \FAINST[216].FA_  ( .A(A[216]), .B(B[216]), .CI(C[216]), .S(S[216]), 
        .CO(C[217]) );
  FA_39 \FAINST[217].FA_  ( .A(A[217]), .B(B[217]), .CI(C[217]), .S(S[217]), 
        .CO(C[218]) );
  FA_38 \FAINST[218].FA_  ( .A(A[218]), .B(B[218]), .CI(C[218]), .S(S[218]), 
        .CO(C[219]) );
  FA_37 \FAINST[219].FA_  ( .A(A[219]), .B(B[219]), .CI(C[219]), .S(S[219]), 
        .CO(C[220]) );
  FA_36 \FAINST[220].FA_  ( .A(A[220]), .B(B[220]), .CI(C[220]), .S(S[220]), 
        .CO(C[221]) );
  FA_35 \FAINST[221].FA_  ( .A(A[221]), .B(B[221]), .CI(C[221]), .S(S[221]), 
        .CO(C[222]) );
  FA_34 \FAINST[222].FA_  ( .A(A[222]), .B(B[222]), .CI(C[222]), .S(S[222]), 
        .CO(C[223]) );
  FA_33 \FAINST[223].FA_  ( .A(A[223]), .B(B[223]), .CI(C[223]), .S(S[223]), 
        .CO(C[224]) );
  FA_32 \FAINST[224].FA_  ( .A(A[224]), .B(B[224]), .CI(C[224]), .S(S[224]), 
        .CO(C[225]) );
  FA_31 \FAINST[225].FA_  ( .A(A[225]), .B(B[225]), .CI(C[225]), .S(S[225]), 
        .CO(C[226]) );
  FA_30 \FAINST[226].FA_  ( .A(A[226]), .B(B[226]), .CI(C[226]), .S(S[226]), 
        .CO(C[227]) );
  FA_29 \FAINST[227].FA_  ( .A(A[227]), .B(B[227]), .CI(C[227]), .S(S[227]), 
        .CO(C[228]) );
  FA_28 \FAINST[228].FA_  ( .A(A[228]), .B(B[228]), .CI(C[228]), .S(S[228]), 
        .CO(C[229]) );
  FA_27 \FAINST[229].FA_  ( .A(A[229]), .B(B[229]), .CI(C[229]), .S(S[229]), 
        .CO(C[230]) );
  FA_26 \FAINST[230].FA_  ( .A(A[230]), .B(B[230]), .CI(C[230]), .S(S[230]), 
        .CO(C[231]) );
  FA_25 \FAINST[231].FA_  ( .A(A[231]), .B(B[231]), .CI(C[231]), .S(S[231]), 
        .CO(C[232]) );
  FA_24 \FAINST[232].FA_  ( .A(A[232]), .B(B[232]), .CI(C[232]), .S(S[232]), 
        .CO(C[233]) );
  FA_23 \FAINST[233].FA_  ( .A(A[233]), .B(B[233]), .CI(C[233]), .S(S[233]), 
        .CO(C[234]) );
  FA_22 \FAINST[234].FA_  ( .A(A[234]), .B(B[234]), .CI(C[234]), .S(S[234]), 
        .CO(C[235]) );
  FA_21 \FAINST[235].FA_  ( .A(A[235]), .B(B[235]), .CI(C[235]), .S(S[235]), 
        .CO(C[236]) );
  FA_20 \FAINST[236].FA_  ( .A(A[236]), .B(B[236]), .CI(C[236]), .S(S[236]), 
        .CO(C[237]) );
  FA_19 \FAINST[237].FA_  ( .A(A[237]), .B(B[237]), .CI(C[237]), .S(S[237]), 
        .CO(C[238]) );
  FA_18 \FAINST[238].FA_  ( .A(A[238]), .B(B[238]), .CI(C[238]), .S(S[238]), 
        .CO(C[239]) );
  FA_17 \FAINST[239].FA_  ( .A(A[239]), .B(B[239]), .CI(C[239]), .S(S[239]), 
        .CO(C[240]) );
  FA_16 \FAINST[240].FA_  ( .A(1'b0), .B(B[240]), .CI(C[240]), .S(S[240]), 
        .CO(C[241]) );
  FA_15 \FAINST[241].FA_  ( .A(1'b0), .B(B[241]), .CI(C[241]), .S(S[241]), 
        .CO(C[242]) );
  FA_14 \FAINST[242].FA_  ( .A(1'b0), .B(B[242]), .CI(C[242]), .S(S[242]), 
        .CO(C[243]) );
  FA_13 \FAINST[243].FA_  ( .A(1'b0), .B(B[243]), .CI(C[243]), .S(S[243]), 
        .CO(C[244]) );
  FA_12 \FAINST[244].FA_  ( .A(1'b0), .B(B[244]), .CI(C[244]), .S(S[244]), 
        .CO(C[245]) );
  FA_11 \FAINST[245].FA_  ( .A(1'b0), .B(B[245]), .CI(C[245]), .S(S[245]), 
        .CO(C[246]) );
  FA_10 \FAINST[246].FA_  ( .A(1'b0), .B(B[246]), .CI(C[246]), .S(S[246]), 
        .CO(C[247]) );
  FA_9 \FAINST[247].FA_  ( .A(1'b0), .B(B[247]), .CI(C[247]), .S(S[247]), .CO(
        C[248]) );
  FA_8 \FAINST[248].FA_  ( .A(1'b0), .B(B[248]), .CI(C[248]), .S(S[248]), .CO(
        C[249]) );
  FA_7 \FAINST[249].FA_  ( .A(1'b0), .B(B[249]), .CI(C[249]), .S(S[249]), .CO(
        C[250]) );
  FA_6 \FAINST[250].FA_  ( .A(1'b0), .B(B[250]), .CI(C[250]), .S(S[250]), .CO(
        C[251]) );
  FA_5 \FAINST[251].FA_  ( .A(1'b0), .B(B[251]), .CI(C[251]), .S(S[251]), .CO(
        C[252]) );
  FA_4 \FAINST[252].FA_  ( .A(1'b0), .B(B[252]), .CI(C[252]), .S(S[252]), .CO(
        C[253]) );
  FA_3 \FAINST[253].FA_  ( .A(1'b0), .B(B[253]), .CI(C[253]), .S(S[253]), .CO(
        C[254]) );
  FA_2 \FAINST[254].FA_  ( .A(1'b0), .B(B[254]), .CI(C[254]), .S(S[254]) );
  FA_1 \FAINST[255].FA_  ( .A(1'b0), .B(B[255]), .CI(1'b0), .S(S[255]) );
endmodule


module mult_N256_CC16_DW01_add_0 ( A, B, CI, SUM, CO );
  input [269:0] A;
  input [269:0] B;
  output [269:0] SUM;
  input CI;
  output CO;
  wire   \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] ,
         \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764;
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  NAND U2 ( .A(n15), .B(n18), .Z(n19) );
  XOR U3 ( .A(n1), .B(n2), .Z(SUM[99]) );
  NANDN U4 ( .A(n3), .B(n4), .Z(n2) );
  ANDN U5 ( .B(n5), .A(n6), .Z(n1) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  XNOR U7 ( .A(n7), .B(n9), .Z(SUM[98]) );
  NANDN U8 ( .A(n6), .B(n8), .Z(n9) );
  NANDN U9 ( .A(n10), .B(n11), .Z(n7) );
  NAND U10 ( .A(n12), .B(n13), .Z(n11) );
  XNOR U11 ( .A(n12), .B(n14), .Z(SUM[97]) );
  NANDN U12 ( .A(n10), .B(n13), .Z(n14) );
  NAND U13 ( .A(n15), .B(n16), .Z(n12) );
  NANDN U14 ( .A(n17), .B(n18), .Z(n16) );
  XOR U15 ( .A(n17), .B(n19), .Z(SUM[96]) );
  XOR U16 ( .A(n20), .B(n21), .Z(SUM[95]) );
  OR U17 ( .A(n22), .B(n23), .Z(n21) );
  ANDN U18 ( .B(n24), .A(n25), .Z(n20) );
  NANDN U19 ( .A(n26), .B(n27), .Z(n24) );
  XNOR U20 ( .A(n27), .B(n28), .Z(SUM[94]) );
  OR U21 ( .A(n26), .B(n25), .Z(n28) );
  NANDN U22 ( .A(n29), .B(n30), .Z(n27) );
  NANDN U23 ( .A(n31), .B(n32), .Z(n30) );
  XNOR U24 ( .A(n32), .B(n33), .Z(SUM[93]) );
  OR U25 ( .A(n31), .B(n29), .Z(n33) );
  NANDN U26 ( .A(n34), .B(n35), .Z(n32) );
  NAND U27 ( .A(n36), .B(n37), .Z(n35) );
  XNOR U28 ( .A(n36), .B(n38), .Z(SUM[92]) );
  NANDN U29 ( .A(n34), .B(n37), .Z(n38) );
  NANDN U30 ( .A(n39), .B(n40), .Z(n36) );
  NANDN U31 ( .A(n41), .B(n42), .Z(n40) );
  XOR U32 ( .A(n43), .B(n44), .Z(SUM[91]) );
  NANDN U33 ( .A(n45), .B(n46), .Z(n44) );
  ANDN U34 ( .B(n47), .A(n48), .Z(n43) );
  NAND U35 ( .A(n49), .B(n50), .Z(n47) );
  XNOR U36 ( .A(n49), .B(n51), .Z(SUM[90]) );
  NANDN U37 ( .A(n48), .B(n50), .Z(n51) );
  NANDN U38 ( .A(n52), .B(n53), .Z(n49) );
  NAND U39 ( .A(n54), .B(n55), .Z(n53) );
  XNOR U40 ( .A(n54), .B(n56), .Z(SUM[89]) );
  NANDN U41 ( .A(n52), .B(n55), .Z(n56) );
  NANDN U42 ( .A(n57), .B(n58), .Z(n54) );
  NAND U43 ( .A(n42), .B(n59), .Z(n58) );
  XNOR U44 ( .A(n42), .B(n60), .Z(SUM[88]) );
  NANDN U45 ( .A(n57), .B(n59), .Z(n60) );
  NANDN U46 ( .A(n61), .B(n62), .Z(n42) );
  NANDN U47 ( .A(n63), .B(n64), .Z(n62) );
  XOR U48 ( .A(n65), .B(n66), .Z(SUM[87]) );
  NANDN U49 ( .A(n67), .B(n68), .Z(n66) );
  ANDN U50 ( .B(n69), .A(n70), .Z(n65) );
  NAND U51 ( .A(n71), .B(n72), .Z(n69) );
  XNOR U52 ( .A(n71), .B(n73), .Z(SUM[86]) );
  NANDN U53 ( .A(n70), .B(n72), .Z(n73) );
  NANDN U54 ( .A(n74), .B(n75), .Z(n71) );
  NAND U55 ( .A(n76), .B(n77), .Z(n75) );
  XNOR U56 ( .A(n76), .B(n78), .Z(SUM[85]) );
  NANDN U57 ( .A(n74), .B(n77), .Z(n78) );
  NANDN U58 ( .A(n79), .B(n80), .Z(n76) );
  NANDN U59 ( .A(n63), .B(n81), .Z(n80) );
  XOR U60 ( .A(n63), .B(n82), .Z(SUM[84]) );
  NANDN U61 ( .A(n79), .B(n81), .Z(n82) );
  ANDN U62 ( .B(n83), .A(n84), .Z(n63) );
  OR U63 ( .A(n85), .B(n86), .Z(n83) );
  XOR U64 ( .A(n87), .B(n88), .Z(SUM[83]) );
  NANDN U65 ( .A(n89), .B(n90), .Z(n88) );
  ANDN U66 ( .B(n91), .A(n92), .Z(n87) );
  NANDN U67 ( .A(n93), .B(n94), .Z(n91) );
  XNOR U68 ( .A(n94), .B(n95), .Z(SUM[82]) );
  OR U69 ( .A(n93), .B(n92), .Z(n95) );
  NANDN U70 ( .A(n96), .B(n97), .Z(n94) );
  NAND U71 ( .A(n98), .B(n99), .Z(n97) );
  XNOR U72 ( .A(n98), .B(n100), .Z(SUM[81]) );
  NANDN U73 ( .A(n96), .B(n99), .Z(n100) );
  NANDN U74 ( .A(n101), .B(n102), .Z(n98) );
  NANDN U75 ( .A(n86), .B(n103), .Z(n102) );
  XOR U76 ( .A(n86), .B(n104), .Z(SUM[80]) );
  NANDN U77 ( .A(n101), .B(n103), .Z(n104) );
  XOR U78 ( .A(n105), .B(n106), .Z(SUM[79]) );
  OR U79 ( .A(n107), .B(n108), .Z(n106) );
  ANDN U80 ( .B(n109), .A(n110), .Z(n105) );
  NANDN U81 ( .A(n111), .B(n112), .Z(n109) );
  XNOR U82 ( .A(n112), .B(n113), .Z(SUM[78]) );
  OR U83 ( .A(n111), .B(n110), .Z(n113) );
  NANDN U84 ( .A(n114), .B(n115), .Z(n112) );
  NANDN U85 ( .A(n116), .B(n117), .Z(n115) );
  XNOR U86 ( .A(n117), .B(n118), .Z(SUM[77]) );
  OR U87 ( .A(n116), .B(n114), .Z(n118) );
  NANDN U88 ( .A(n119), .B(n120), .Z(n117) );
  NAND U89 ( .A(n121), .B(n122), .Z(n120) );
  XNOR U90 ( .A(n121), .B(n123), .Z(SUM[76]) );
  NANDN U91 ( .A(n119), .B(n122), .Z(n123) );
  NANDN U92 ( .A(n124), .B(n125), .Z(n121) );
  NANDN U93 ( .A(n126), .B(n127), .Z(n125) );
  XOR U94 ( .A(n128), .B(n129), .Z(SUM[75]) );
  NANDN U95 ( .A(n130), .B(n131), .Z(n129) );
  ANDN U96 ( .B(n132), .A(n133), .Z(n128) );
  NAND U97 ( .A(n134), .B(n135), .Z(n132) );
  XNOR U98 ( .A(n134), .B(n136), .Z(SUM[74]) );
  NANDN U99 ( .A(n133), .B(n135), .Z(n136) );
  NANDN U100 ( .A(n137), .B(n138), .Z(n134) );
  NAND U101 ( .A(n139), .B(n140), .Z(n138) );
  XNOR U102 ( .A(n139), .B(n141), .Z(SUM[73]) );
  NANDN U103 ( .A(n137), .B(n140), .Z(n141) );
  NANDN U104 ( .A(n142), .B(n143), .Z(n139) );
  NAND U105 ( .A(n127), .B(n144), .Z(n143) );
  XNOR U106 ( .A(n127), .B(n145), .Z(SUM[72]) );
  NANDN U107 ( .A(n142), .B(n144), .Z(n145) );
  NANDN U108 ( .A(n146), .B(n147), .Z(n127) );
  NANDN U109 ( .A(n148), .B(n149), .Z(n147) );
  XOR U110 ( .A(n150), .B(n151), .Z(SUM[71]) );
  NANDN U111 ( .A(n152), .B(n153), .Z(n151) );
  ANDN U112 ( .B(n154), .A(n155), .Z(n150) );
  NAND U113 ( .A(n156), .B(n157), .Z(n154) );
  XNOR U114 ( .A(n156), .B(n158), .Z(SUM[70]) );
  NANDN U115 ( .A(n155), .B(n157), .Z(n158) );
  NANDN U116 ( .A(n159), .B(n160), .Z(n156) );
  NAND U117 ( .A(n161), .B(n162), .Z(n160) );
  XNOR U118 ( .A(n161), .B(n163), .Z(SUM[69]) );
  NANDN U119 ( .A(n159), .B(n162), .Z(n163) );
  NANDN U120 ( .A(n164), .B(n165), .Z(n161) );
  NANDN U121 ( .A(n148), .B(n166), .Z(n165) );
  XOR U122 ( .A(n148), .B(n167), .Z(SUM[68]) );
  NANDN U123 ( .A(n164), .B(n166), .Z(n167) );
  ANDN U124 ( .B(n168), .A(n169), .Z(n148) );
  OR U125 ( .A(n170), .B(n171), .Z(n168) );
  XOR U126 ( .A(n172), .B(n173), .Z(SUM[67]) );
  NANDN U127 ( .A(n174), .B(n175), .Z(n173) );
  ANDN U128 ( .B(n176), .A(n177), .Z(n172) );
  NANDN U129 ( .A(n178), .B(n179), .Z(n176) );
  XNOR U130 ( .A(n179), .B(n180), .Z(SUM[66]) );
  OR U131 ( .A(n178), .B(n177), .Z(n180) );
  NANDN U132 ( .A(n181), .B(n182), .Z(n179) );
  NAND U133 ( .A(n183), .B(n184), .Z(n182) );
  XNOR U134 ( .A(n183), .B(n185), .Z(SUM[65]) );
  NANDN U135 ( .A(n181), .B(n184), .Z(n185) );
  NANDN U136 ( .A(n186), .B(n187), .Z(n183) );
  NANDN U137 ( .A(n171), .B(n188), .Z(n187) );
  XOR U138 ( .A(n171), .B(n189), .Z(SUM[64]) );
  NANDN U139 ( .A(n186), .B(n188), .Z(n189) );
  XOR U140 ( .A(n190), .B(n191), .Z(SUM[63]) );
  OR U141 ( .A(n192), .B(n193), .Z(n191) );
  ANDN U142 ( .B(n194), .A(n195), .Z(n190) );
  NANDN U143 ( .A(n196), .B(n197), .Z(n194) );
  XNOR U144 ( .A(n197), .B(n198), .Z(SUM[62]) );
  OR U145 ( .A(n196), .B(n195), .Z(n198) );
  NANDN U146 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U147 ( .A(n201), .B(n202), .Z(n200) );
  XNOR U148 ( .A(n202), .B(n203), .Z(SUM[61]) );
  OR U149 ( .A(n201), .B(n199), .Z(n203) );
  NANDN U150 ( .A(n204), .B(n205), .Z(n202) );
  NANDN U151 ( .A(n206), .B(n207), .Z(n205) );
  XNOR U152 ( .A(n207), .B(n208), .Z(SUM[60]) );
  OR U153 ( .A(n206), .B(n204), .Z(n208) );
  NANDN U154 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U155 ( .A(n211), .B(n212), .Z(n210) );
  XOR U156 ( .A(n213), .B(n214), .Z(SUM[59]) );
  NANDN U157 ( .A(n215), .B(n216), .Z(n214) );
  ANDN U158 ( .B(n217), .A(n218), .Z(n213) );
  NAND U159 ( .A(n219), .B(n220), .Z(n217) );
  XNOR U160 ( .A(n219), .B(n221), .Z(SUM[58]) );
  NANDN U161 ( .A(n218), .B(n220), .Z(n221) );
  NANDN U162 ( .A(n222), .B(n223), .Z(n219) );
  NAND U163 ( .A(n224), .B(n225), .Z(n223) );
  XNOR U164 ( .A(n224), .B(n226), .Z(SUM[57]) );
  NANDN U165 ( .A(n222), .B(n225), .Z(n226) );
  NANDN U166 ( .A(n227), .B(n228), .Z(n224) );
  NAND U167 ( .A(n212), .B(n229), .Z(n228) );
  XNOR U168 ( .A(n212), .B(n230), .Z(SUM[56]) );
  NANDN U169 ( .A(n227), .B(n229), .Z(n230) );
  NANDN U170 ( .A(n231), .B(n232), .Z(n212) );
  OR U171 ( .A(n233), .B(n234), .Z(n232) );
  XOR U172 ( .A(n235), .B(n236), .Z(SUM[55]) );
  NANDN U173 ( .A(n237), .B(n238), .Z(n236) );
  ANDN U174 ( .B(n239), .A(n240), .Z(n235) );
  NAND U175 ( .A(n241), .B(n242), .Z(n239) );
  XNOR U176 ( .A(n241), .B(n243), .Z(SUM[54]) );
  NANDN U177 ( .A(n240), .B(n242), .Z(n243) );
  NANDN U178 ( .A(n244), .B(n245), .Z(n241) );
  NAND U179 ( .A(n246), .B(n247), .Z(n245) );
  XNOR U180 ( .A(n246), .B(n248), .Z(SUM[53]) );
  NANDN U181 ( .A(n244), .B(n247), .Z(n248) );
  NANDN U182 ( .A(n249), .B(n250), .Z(n246) );
  NANDN U183 ( .A(n234), .B(n251), .Z(n250) );
  XOR U184 ( .A(n234), .B(n252), .Z(SUM[52]) );
  NANDN U185 ( .A(n249), .B(n251), .Z(n252) );
  NOR U186 ( .A(n253), .B(n254), .Z(n234) );
  XOR U187 ( .A(n255), .B(n256), .Z(SUM[51]) );
  NANDN U188 ( .A(n257), .B(n258), .Z(n256) );
  ANDN U189 ( .B(n259), .A(n260), .Z(n255) );
  NAND U190 ( .A(n261), .B(n262), .Z(n259) );
  XNOR U191 ( .A(n261), .B(n263), .Z(SUM[50]) );
  NANDN U192 ( .A(n260), .B(n262), .Z(n263) );
  NANDN U193 ( .A(n264), .B(n265), .Z(n261) );
  NAND U194 ( .A(n266), .B(n267), .Z(n265) );
  XNOR U195 ( .A(n266), .B(n268), .Z(SUM[49]) );
  NANDN U196 ( .A(n264), .B(n267), .Z(n268) );
  NANDN U197 ( .A(n269), .B(n270), .Z(n266) );
  NANDN U198 ( .A(n271), .B(n272), .Z(n270) );
  XOR U199 ( .A(n271), .B(n273), .Z(SUM[48]) );
  NANDN U200 ( .A(n269), .B(n272), .Z(n273) );
  XOR U201 ( .A(n274), .B(n275), .Z(SUM[47]) );
  OR U202 ( .A(n276), .B(n277), .Z(n275) );
  ANDN U203 ( .B(n278), .A(n279), .Z(n274) );
  NANDN U204 ( .A(n280), .B(n281), .Z(n278) );
  XNOR U205 ( .A(n281), .B(n282), .Z(SUM[46]) );
  OR U206 ( .A(n280), .B(n279), .Z(n282) );
  NANDN U207 ( .A(n283), .B(n284), .Z(n281) );
  NANDN U208 ( .A(n285), .B(n286), .Z(n284) );
  XNOR U209 ( .A(n286), .B(n287), .Z(SUM[45]) );
  OR U210 ( .A(n285), .B(n283), .Z(n287) );
  NANDN U211 ( .A(n288), .B(n289), .Z(n286) );
  NAND U212 ( .A(n290), .B(n291), .Z(n289) );
  XNOR U213 ( .A(n290), .B(n292), .Z(SUM[44]) );
  NANDN U214 ( .A(n288), .B(n291), .Z(n292) );
  NANDN U215 ( .A(n293), .B(n294), .Z(n290) );
  NANDN U216 ( .A(n295), .B(n296), .Z(n294) );
  XOR U217 ( .A(n297), .B(n298), .Z(SUM[43]) );
  NANDN U218 ( .A(n299), .B(n300), .Z(n298) );
  ANDN U219 ( .B(n301), .A(n302), .Z(n297) );
  NAND U220 ( .A(n303), .B(n304), .Z(n301) );
  XNOR U221 ( .A(n303), .B(n305), .Z(SUM[42]) );
  NANDN U222 ( .A(n302), .B(n304), .Z(n305) );
  NANDN U223 ( .A(n306), .B(n307), .Z(n303) );
  NAND U224 ( .A(n308), .B(n309), .Z(n307) );
  XNOR U225 ( .A(n308), .B(n310), .Z(SUM[41]) );
  NANDN U226 ( .A(n306), .B(n309), .Z(n310) );
  NANDN U227 ( .A(n311), .B(n312), .Z(n308) );
  NAND U228 ( .A(n296), .B(n313), .Z(n312) );
  XNOR U229 ( .A(n296), .B(n314), .Z(SUM[40]) );
  NANDN U230 ( .A(n311), .B(n313), .Z(n314) );
  NANDN U231 ( .A(n315), .B(n316), .Z(n296) );
  NANDN U232 ( .A(n317), .B(n318), .Z(n316) );
  XOR U233 ( .A(n319), .B(n320), .Z(SUM[39]) );
  NANDN U234 ( .A(n321), .B(n322), .Z(n320) );
  ANDN U235 ( .B(n323), .A(n324), .Z(n319) );
  NAND U236 ( .A(n325), .B(n326), .Z(n323) );
  XNOR U237 ( .A(n325), .B(n327), .Z(SUM[38]) );
  NANDN U238 ( .A(n324), .B(n326), .Z(n327) );
  NANDN U239 ( .A(n328), .B(n329), .Z(n325) );
  NAND U240 ( .A(n330), .B(n331), .Z(n329) );
  XNOR U241 ( .A(n330), .B(n332), .Z(SUM[37]) );
  NANDN U242 ( .A(n328), .B(n331), .Z(n332) );
  NANDN U243 ( .A(n333), .B(n334), .Z(n330) );
  NANDN U244 ( .A(n317), .B(n335), .Z(n334) );
  XOR U245 ( .A(n317), .B(n336), .Z(SUM[36]) );
  NANDN U246 ( .A(n333), .B(n335), .Z(n336) );
  ANDN U247 ( .B(n337), .A(n338), .Z(n317) );
  OR U248 ( .A(n339), .B(n340), .Z(n337) );
  XOR U249 ( .A(n341), .B(n342), .Z(SUM[35]) );
  NANDN U250 ( .A(n343), .B(n344), .Z(n342) );
  ANDN U251 ( .B(n345), .A(n346), .Z(n341) );
  NANDN U252 ( .A(n347), .B(n348), .Z(n345) );
  XNOR U253 ( .A(n348), .B(n349), .Z(SUM[34]) );
  OR U254 ( .A(n347), .B(n346), .Z(n349) );
  NANDN U255 ( .A(n350), .B(n351), .Z(n348) );
  NAND U256 ( .A(n352), .B(n353), .Z(n351) );
  XNOR U257 ( .A(n352), .B(n354), .Z(SUM[33]) );
  NANDN U258 ( .A(n350), .B(n353), .Z(n354) );
  NANDN U259 ( .A(n355), .B(n356), .Z(n352) );
  NANDN U260 ( .A(n340), .B(n357), .Z(n356) );
  XOR U261 ( .A(n340), .B(n358), .Z(SUM[32]) );
  NANDN U262 ( .A(n355), .B(n357), .Z(n358) );
  XOR U263 ( .A(n359), .B(n360), .Z(SUM[31]) );
  OR U264 ( .A(n361), .B(n362), .Z(n360) );
  ANDN U265 ( .B(n363), .A(n364), .Z(n359) );
  NANDN U266 ( .A(n365), .B(n366), .Z(n363) );
  XNOR U267 ( .A(n366), .B(n367), .Z(SUM[30]) );
  OR U268 ( .A(n365), .B(n364), .Z(n367) );
  NANDN U269 ( .A(n368), .B(n369), .Z(n366) );
  NANDN U270 ( .A(n370), .B(n371), .Z(n369) );
  XNOR U271 ( .A(n371), .B(n372), .Z(SUM[29]) );
  OR U272 ( .A(n370), .B(n368), .Z(n372) );
  NANDN U273 ( .A(n373), .B(n374), .Z(n371) );
  NAND U274 ( .A(n375), .B(n376), .Z(n374) );
  XNOR U275 ( .A(n375), .B(n377), .Z(SUM[28]) );
  NANDN U276 ( .A(n373), .B(n376), .Z(n377) );
  NANDN U277 ( .A(n378), .B(n379), .Z(n375) );
  NANDN U278 ( .A(n380), .B(n381), .Z(n379) );
  XOR U279 ( .A(n382), .B(n383), .Z(SUM[27]) );
  NANDN U280 ( .A(n384), .B(n385), .Z(n383) );
  ANDN U281 ( .B(n386), .A(n387), .Z(n382) );
  NAND U282 ( .A(n388), .B(n389), .Z(n386) );
  XNOR U283 ( .A(n388), .B(n390), .Z(SUM[26]) );
  NANDN U284 ( .A(n387), .B(n389), .Z(n390) );
  NANDN U285 ( .A(n391), .B(n392), .Z(n388) );
  NAND U286 ( .A(n393), .B(n394), .Z(n392) );
  XNOR U287 ( .A(n393), .B(n395), .Z(SUM[25]) );
  NANDN U288 ( .A(n391), .B(n394), .Z(n395) );
  NANDN U289 ( .A(n396), .B(n397), .Z(n393) );
  NAND U290 ( .A(n381), .B(n398), .Z(n397) );
  XOR U291 ( .A(n399), .B(n400), .Z(SUM[253]) );
  XNOR U292 ( .A(B[253]), .B(A[253]), .Z(n400) );
  ANDN U293 ( .B(n401), .A(n402), .Z(n399) );
  NAND U294 ( .A(n403), .B(n404), .Z(n401) );
  XNOR U295 ( .A(n403), .B(n405), .Z(SUM[252]) );
  NANDN U296 ( .A(n402), .B(n404), .Z(n405) );
  OR U297 ( .A(B[252]), .B(A[252]), .Z(n404) );
  AND U298 ( .A(B[252]), .B(A[252]), .Z(n402) );
  NANDN U299 ( .A(n406), .B(n407), .Z(n403) );
  NAND U300 ( .A(n408), .B(n409), .Z(n407) );
  XNOR U301 ( .A(n408), .B(n410), .Z(SUM[251]) );
  NANDN U302 ( .A(n406), .B(n409), .Z(n410) );
  OR U303 ( .A(B[251]), .B(A[251]), .Z(n409) );
  AND U304 ( .A(B[251]), .B(A[251]), .Z(n406) );
  NANDN U305 ( .A(n411), .B(n412), .Z(n408) );
  NAND U306 ( .A(n413), .B(n414), .Z(n412) );
  XNOR U307 ( .A(n413), .B(n415), .Z(SUM[250]) );
  NANDN U308 ( .A(n411), .B(n414), .Z(n415) );
  OR U309 ( .A(B[250]), .B(A[250]), .Z(n414) );
  AND U310 ( .A(B[250]), .B(A[250]), .Z(n411) );
  NANDN U311 ( .A(n416), .B(n417), .Z(n413) );
  NAND U312 ( .A(n418), .B(n419), .Z(n417) );
  XNOR U313 ( .A(n381), .B(n420), .Z(SUM[24]) );
  NANDN U314 ( .A(n396), .B(n398), .Z(n420) );
  NANDN U315 ( .A(n421), .B(n422), .Z(n381) );
  NANDN U316 ( .A(n423), .B(n424), .Z(n422) );
  XNOR U317 ( .A(n418), .B(n425), .Z(SUM[249]) );
  NANDN U318 ( .A(n416), .B(n419), .Z(n425) );
  OR U319 ( .A(B[249]), .B(A[249]), .Z(n419) );
  AND U320 ( .A(B[249]), .B(A[249]), .Z(n416) );
  NANDN U321 ( .A(n426), .B(n427), .Z(n418) );
  NAND U322 ( .A(n428), .B(n429), .Z(n427) );
  XNOR U323 ( .A(n428), .B(n430), .Z(SUM[248]) );
  NANDN U324 ( .A(n426), .B(n429), .Z(n430) );
  OR U325 ( .A(B[248]), .B(A[248]), .Z(n429) );
  AND U326 ( .A(B[248]), .B(A[248]), .Z(n426) );
  NANDN U327 ( .A(n431), .B(n432), .Z(n428) );
  NAND U328 ( .A(n433), .B(n434), .Z(n432) );
  XNOR U329 ( .A(n433), .B(n435), .Z(SUM[247]) );
  NANDN U330 ( .A(n431), .B(n434), .Z(n435) );
  OR U331 ( .A(B[247]), .B(A[247]), .Z(n434) );
  AND U332 ( .A(B[247]), .B(A[247]), .Z(n431) );
  NANDN U333 ( .A(n436), .B(n437), .Z(n433) );
  NAND U334 ( .A(n438), .B(n439), .Z(n437) );
  XNOR U335 ( .A(n438), .B(n440), .Z(SUM[246]) );
  NANDN U336 ( .A(n436), .B(n439), .Z(n440) );
  OR U337 ( .A(B[246]), .B(A[246]), .Z(n439) );
  AND U338 ( .A(B[246]), .B(A[246]), .Z(n436) );
  NANDN U339 ( .A(n441), .B(n442), .Z(n438) );
  NAND U340 ( .A(n443), .B(n444), .Z(n442) );
  XNOR U341 ( .A(n443), .B(n445), .Z(SUM[245]) );
  NANDN U342 ( .A(n441), .B(n444), .Z(n445) );
  OR U343 ( .A(B[245]), .B(A[245]), .Z(n444) );
  AND U344 ( .A(B[245]), .B(A[245]), .Z(n441) );
  NANDN U345 ( .A(n446), .B(n447), .Z(n443) );
  NAND U346 ( .A(n448), .B(n449), .Z(n447) );
  XNOR U347 ( .A(n448), .B(n450), .Z(SUM[244]) );
  NANDN U348 ( .A(n446), .B(n449), .Z(n450) );
  OR U349 ( .A(B[244]), .B(A[244]), .Z(n449) );
  AND U350 ( .A(B[244]), .B(A[244]), .Z(n446) );
  NANDN U351 ( .A(n451), .B(n452), .Z(n448) );
  NAND U352 ( .A(n453), .B(n454), .Z(n452) );
  XNOR U353 ( .A(n453), .B(n455), .Z(SUM[243]) );
  NANDN U354 ( .A(n451), .B(n454), .Z(n455) );
  OR U355 ( .A(B[243]), .B(A[243]), .Z(n454) );
  AND U356 ( .A(B[243]), .B(A[243]), .Z(n451) );
  NANDN U357 ( .A(n456), .B(n457), .Z(n453) );
  NAND U358 ( .A(n458), .B(n459), .Z(n457) );
  XNOR U359 ( .A(n458), .B(n460), .Z(SUM[242]) );
  NANDN U360 ( .A(n456), .B(n459), .Z(n460) );
  OR U361 ( .A(B[242]), .B(A[242]), .Z(n459) );
  AND U362 ( .A(B[242]), .B(A[242]), .Z(n456) );
  NANDN U363 ( .A(n461), .B(n462), .Z(n458) );
  NAND U364 ( .A(n463), .B(n464), .Z(n462) );
  XNOR U365 ( .A(n463), .B(n465), .Z(SUM[241]) );
  NANDN U366 ( .A(n461), .B(n464), .Z(n465) );
  OR U367 ( .A(B[241]), .B(A[241]), .Z(n464) );
  AND U368 ( .A(B[241]), .B(A[241]), .Z(n461) );
  NANDN U369 ( .A(n466), .B(n467), .Z(n463) );
  NAND U370 ( .A(n468), .B(n469), .Z(n467) );
  XNOR U371 ( .A(n468), .B(n470), .Z(SUM[240]) );
  NANDN U372 ( .A(n466), .B(n469), .Z(n470) );
  OR U373 ( .A(B[240]), .B(A[240]), .Z(n469) );
  AND U374 ( .A(B[240]), .B(A[240]), .Z(n466) );
  NANDN U375 ( .A(n471), .B(n472), .Z(n468) );
  NANDN U376 ( .A(n473), .B(n474), .Z(n472) );
  NANDN U377 ( .A(n475), .B(n476), .Z(n474) );
  NANDN U378 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U379 ( .A(n479), .B(n480), .Z(n478) );
  NANDN U380 ( .A(n481), .B(n482), .Z(n480) );
  NANDN U381 ( .A(n483), .B(n484), .Z(n482) );
  NANDN U382 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U383 ( .A(n487), .B(n488), .Z(n486) );
  NANDN U384 ( .A(n489), .B(n490), .Z(n488) );
  NANDN U385 ( .A(n491), .B(n492), .Z(n490) );
  AND U386 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U387 ( .A(n495), .B(n496), .Z(n494) );
  NANDN U388 ( .A(n495), .B(n497), .Z(n493) );
  XOR U389 ( .A(n498), .B(n499), .Z(SUM[23]) );
  NANDN U390 ( .A(n500), .B(n501), .Z(n499) );
  ANDN U391 ( .B(n502), .A(n503), .Z(n498) );
  NAND U392 ( .A(n504), .B(n505), .Z(n502) );
  XOR U393 ( .A(n506), .B(n507), .Z(SUM[239]) );
  OR U394 ( .A(n473), .B(n471), .Z(n507) );
  AND U395 ( .A(B[239]), .B(A[239]), .Z(n471) );
  NOR U396 ( .A(B[239]), .B(A[239]), .Z(n473) );
  ANDN U397 ( .B(n508), .A(n475), .Z(n506) );
  NANDN U398 ( .A(n477), .B(n509), .Z(n508) );
  XNOR U399 ( .A(n509), .B(n510), .Z(SUM[238]) );
  OR U400 ( .A(n477), .B(n475), .Z(n510) );
  AND U401 ( .A(B[238]), .B(A[238]), .Z(n475) );
  NOR U402 ( .A(B[238]), .B(A[238]), .Z(n477) );
  NANDN U403 ( .A(n479), .B(n511), .Z(n509) );
  NANDN U404 ( .A(n481), .B(n512), .Z(n511) );
  XNOR U405 ( .A(n512), .B(n513), .Z(SUM[237]) );
  OR U406 ( .A(n481), .B(n479), .Z(n513) );
  AND U407 ( .A(B[237]), .B(A[237]), .Z(n479) );
  NOR U408 ( .A(B[237]), .B(A[237]), .Z(n481) );
  NANDN U409 ( .A(n483), .B(n514), .Z(n512) );
  NANDN U410 ( .A(n485), .B(n515), .Z(n514) );
  XNOR U411 ( .A(n515), .B(n516), .Z(SUM[236]) );
  OR U412 ( .A(n485), .B(n483), .Z(n516) );
  AND U413 ( .A(B[236]), .B(A[236]), .Z(n483) );
  NOR U414 ( .A(B[236]), .B(A[236]), .Z(n485) );
  NANDN U415 ( .A(n487), .B(n517), .Z(n515) );
  NANDN U416 ( .A(n489), .B(n518), .Z(n517) );
  NAND U417 ( .A(n519), .B(n520), .Z(n489) );
  AND U418 ( .A(n521), .B(n522), .Z(n520) );
  AND U419 ( .A(n523), .B(n524), .Z(n519) );
  NANDN U420 ( .A(n525), .B(n526), .Z(n487) );
  NAND U421 ( .A(n527), .B(n524), .Z(n526) );
  NANDN U422 ( .A(n528), .B(n529), .Z(n527) );
  NAND U423 ( .A(n530), .B(n523), .Z(n529) );
  NANDN U424 ( .A(n531), .B(n532), .Z(n530) );
  NAND U425 ( .A(n522), .B(n533), .Z(n532) );
  XOR U426 ( .A(n534), .B(n535), .Z(SUM[235]) );
  NANDN U427 ( .A(n525), .B(n524), .Z(n535) );
  OR U428 ( .A(B[235]), .B(A[235]), .Z(n524) );
  AND U429 ( .A(B[235]), .B(A[235]), .Z(n525) );
  ANDN U430 ( .B(n536), .A(n528), .Z(n534) );
  NAND U431 ( .A(n537), .B(n523), .Z(n536) );
  XNOR U432 ( .A(n537), .B(n538), .Z(SUM[234]) );
  NANDN U433 ( .A(n528), .B(n523), .Z(n538) );
  OR U434 ( .A(B[234]), .B(A[234]), .Z(n523) );
  AND U435 ( .A(B[234]), .B(A[234]), .Z(n528) );
  NANDN U436 ( .A(n531), .B(n539), .Z(n537) );
  NAND U437 ( .A(n540), .B(n522), .Z(n539) );
  XNOR U438 ( .A(n540), .B(n541), .Z(SUM[233]) );
  NANDN U439 ( .A(n531), .B(n522), .Z(n541) );
  OR U440 ( .A(B[233]), .B(A[233]), .Z(n522) );
  AND U441 ( .A(B[233]), .B(A[233]), .Z(n531) );
  NANDN U442 ( .A(n533), .B(n542), .Z(n540) );
  NAND U443 ( .A(n518), .B(n521), .Z(n542) );
  XNOR U444 ( .A(n518), .B(n543), .Z(SUM[232]) );
  NANDN U445 ( .A(n533), .B(n521), .Z(n543) );
  OR U446 ( .A(B[232]), .B(A[232]), .Z(n521) );
  AND U447 ( .A(B[232]), .B(A[232]), .Z(n533) );
  NANDN U448 ( .A(n491), .B(n544), .Z(n518) );
  OR U449 ( .A(n495), .B(n545), .Z(n544) );
  NAND U450 ( .A(n546), .B(n547), .Z(n495) );
  AND U451 ( .A(n548), .B(n549), .Z(n547) );
  AND U452 ( .A(n550), .B(n551), .Z(n546) );
  NANDN U453 ( .A(n552), .B(n553), .Z(n491) );
  NAND U454 ( .A(n554), .B(n551), .Z(n553) );
  NANDN U455 ( .A(n555), .B(n556), .Z(n554) );
  NAND U456 ( .A(n557), .B(n550), .Z(n556) );
  NANDN U457 ( .A(n558), .B(n559), .Z(n557) );
  NAND U458 ( .A(n549), .B(n560), .Z(n559) );
  XOR U459 ( .A(n561), .B(n562), .Z(SUM[231]) );
  NANDN U460 ( .A(n552), .B(n551), .Z(n562) );
  OR U461 ( .A(B[231]), .B(A[231]), .Z(n551) );
  AND U462 ( .A(B[231]), .B(A[231]), .Z(n552) );
  ANDN U463 ( .B(n563), .A(n555), .Z(n561) );
  NAND U464 ( .A(n564), .B(n550), .Z(n563) );
  XNOR U465 ( .A(n564), .B(n565), .Z(SUM[230]) );
  NANDN U466 ( .A(n555), .B(n550), .Z(n565) );
  OR U467 ( .A(A[230]), .B(B[230]), .Z(n550) );
  AND U468 ( .A(A[230]), .B(B[230]), .Z(n555) );
  NANDN U469 ( .A(n558), .B(n566), .Z(n564) );
  NAND U470 ( .A(n567), .B(n549), .Z(n566) );
  XNOR U471 ( .A(n504), .B(n568), .Z(SUM[22]) );
  NANDN U472 ( .A(n503), .B(n505), .Z(n568) );
  NANDN U473 ( .A(n569), .B(n570), .Z(n504) );
  NAND U474 ( .A(n571), .B(n572), .Z(n570) );
  XNOR U475 ( .A(n567), .B(n573), .Z(SUM[229]) );
  NANDN U476 ( .A(n558), .B(n549), .Z(n573) );
  OR U477 ( .A(A[229]), .B(B[229]), .Z(n549) );
  AND U478 ( .A(A[229]), .B(B[229]), .Z(n558) );
  NANDN U479 ( .A(n560), .B(n574), .Z(n567) );
  NANDN U480 ( .A(n545), .B(n548), .Z(n574) );
  XOR U481 ( .A(n545), .B(n575), .Z(SUM[228]) );
  NANDN U482 ( .A(n560), .B(n548), .Z(n575) );
  OR U483 ( .A(A[228]), .B(B[228]), .Z(n548) );
  AND U484 ( .A(A[228]), .B(B[228]), .Z(n560) );
  NOR U485 ( .A(n496), .B(n497), .Z(n545) );
  AND U486 ( .A(n576), .B(n577), .Z(n497) );
  AND U487 ( .A(n578), .B(n579), .Z(n577) );
  NOR U488 ( .A(n580), .B(n581), .Z(n579) );
  AND U489 ( .A(n582), .B(n583), .Z(n576) );
  NANDN U490 ( .A(n584), .B(n585), .Z(n496) );
  NAND U491 ( .A(n586), .B(n583), .Z(n585) );
  NANDN U492 ( .A(n587), .B(n588), .Z(n586) );
  NAND U493 ( .A(n589), .B(n582), .Z(n588) );
  NANDN U494 ( .A(n590), .B(n591), .Z(n589) );
  NAND U495 ( .A(n578), .B(n592), .Z(n591) );
  XOR U496 ( .A(n593), .B(n594), .Z(SUM[227]) );
  NANDN U497 ( .A(n584), .B(n583), .Z(n594) );
  OR U498 ( .A(B[227]), .B(A[227]), .Z(n583) );
  AND U499 ( .A(B[227]), .B(A[227]), .Z(n584) );
  ANDN U500 ( .B(n595), .A(n587), .Z(n593) );
  NAND U501 ( .A(n596), .B(n582), .Z(n595) );
  XNOR U502 ( .A(n596), .B(n597), .Z(SUM[226]) );
  NANDN U503 ( .A(n587), .B(n582), .Z(n597) );
  OR U504 ( .A(A[226]), .B(B[226]), .Z(n582) );
  AND U505 ( .A(A[226]), .B(B[226]), .Z(n587) );
  NANDN U506 ( .A(n590), .B(n598), .Z(n596) );
  NAND U507 ( .A(n599), .B(n578), .Z(n598) );
  XNOR U508 ( .A(n599), .B(n600), .Z(SUM[225]) );
  NANDN U509 ( .A(n590), .B(n578), .Z(n600) );
  OR U510 ( .A(A[225]), .B(B[225]), .Z(n578) );
  AND U511 ( .A(A[225]), .B(B[225]), .Z(n590) );
  NANDN U512 ( .A(n592), .B(n601), .Z(n599) );
  OR U513 ( .A(n580), .B(n581), .Z(n601) );
  XOR U514 ( .A(n580), .B(n602), .Z(SUM[224]) );
  OR U515 ( .A(n581), .B(n592), .Z(n602) );
  AND U516 ( .A(A[224]), .B(B[224]), .Z(n592) );
  NOR U517 ( .A(B[224]), .B(A[224]), .Z(n581) );
  ANDN U518 ( .B(n603), .A(n604), .Z(n580) );
  NANDN U519 ( .A(n605), .B(n606), .Z(n603) );
  NANDN U520 ( .A(n607), .B(n608), .Z(n606) );
  NANDN U521 ( .A(n609), .B(n610), .Z(n608) );
  NANDN U522 ( .A(n611), .B(n612), .Z(n610) );
  NANDN U523 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U524 ( .A(n615), .B(n616), .Z(n614) );
  NANDN U525 ( .A(n617), .B(n618), .Z(n616) );
  NANDN U526 ( .A(n619), .B(n620), .Z(n618) );
  NANDN U527 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U528 ( .A(n623), .B(n624), .Z(n622) );
  AND U529 ( .A(n625), .B(n626), .Z(n624) );
  NANDN U530 ( .A(n627), .B(n628), .Z(n626) );
  NANDN U531 ( .A(n627), .B(n629), .Z(n625) );
  XOR U532 ( .A(n630), .B(n631), .Z(SUM[223]) );
  OR U533 ( .A(n605), .B(n604), .Z(n631) );
  AND U534 ( .A(B[223]), .B(A[223]), .Z(n604) );
  NOR U535 ( .A(B[223]), .B(A[223]), .Z(n605) );
  ANDN U536 ( .B(n632), .A(n607), .Z(n630) );
  NANDN U537 ( .A(n609), .B(n633), .Z(n632) );
  XNOR U538 ( .A(n633), .B(n634), .Z(SUM[222]) );
  OR U539 ( .A(n609), .B(n607), .Z(n634) );
  AND U540 ( .A(B[222]), .B(A[222]), .Z(n607) );
  NOR U541 ( .A(B[222]), .B(A[222]), .Z(n609) );
  NANDN U542 ( .A(n611), .B(n635), .Z(n633) );
  NANDN U543 ( .A(n613), .B(n636), .Z(n635) );
  XNOR U544 ( .A(n636), .B(n637), .Z(SUM[221]) );
  OR U545 ( .A(n613), .B(n611), .Z(n637) );
  AND U546 ( .A(B[221]), .B(A[221]), .Z(n611) );
  NOR U547 ( .A(B[221]), .B(A[221]), .Z(n613) );
  NANDN U548 ( .A(n615), .B(n638), .Z(n636) );
  NANDN U549 ( .A(n617), .B(n639), .Z(n638) );
  XNOR U550 ( .A(n639), .B(n640), .Z(SUM[220]) );
  OR U551 ( .A(n617), .B(n615), .Z(n640) );
  AND U552 ( .A(B[220]), .B(A[220]), .Z(n615) );
  NOR U553 ( .A(B[220]), .B(A[220]), .Z(n617) );
  NANDN U554 ( .A(n619), .B(n641), .Z(n639) );
  NANDN U555 ( .A(n621), .B(n642), .Z(n641) );
  NAND U556 ( .A(n643), .B(n644), .Z(n621) );
  AND U557 ( .A(n645), .B(n646), .Z(n644) );
  AND U558 ( .A(n647), .B(n648), .Z(n643) );
  NANDN U559 ( .A(n649), .B(n650), .Z(n619) );
  NAND U560 ( .A(n651), .B(n648), .Z(n650) );
  NANDN U561 ( .A(n652), .B(n653), .Z(n651) );
  NAND U562 ( .A(n654), .B(n647), .Z(n653) );
  NANDN U563 ( .A(n655), .B(n656), .Z(n654) );
  NAND U564 ( .A(n646), .B(n657), .Z(n656) );
  XNOR U565 ( .A(n571), .B(n658), .Z(SUM[21]) );
  NANDN U566 ( .A(n569), .B(n572), .Z(n658) );
  NANDN U567 ( .A(n659), .B(n660), .Z(n571) );
  NANDN U568 ( .A(n423), .B(n661), .Z(n660) );
  XOR U569 ( .A(n662), .B(n663), .Z(SUM[219]) );
  NANDN U570 ( .A(n649), .B(n648), .Z(n663) );
  OR U571 ( .A(B[219]), .B(A[219]), .Z(n648) );
  AND U572 ( .A(B[219]), .B(A[219]), .Z(n649) );
  ANDN U573 ( .B(n664), .A(n652), .Z(n662) );
  NAND U574 ( .A(n665), .B(n647), .Z(n664) );
  XNOR U575 ( .A(n665), .B(n666), .Z(SUM[218]) );
  NANDN U576 ( .A(n652), .B(n647), .Z(n666) );
  OR U577 ( .A(B[218]), .B(A[218]), .Z(n647) );
  AND U578 ( .A(B[218]), .B(A[218]), .Z(n652) );
  NANDN U579 ( .A(n655), .B(n667), .Z(n665) );
  NAND U580 ( .A(n668), .B(n646), .Z(n667) );
  XNOR U581 ( .A(n668), .B(n669), .Z(SUM[217]) );
  NANDN U582 ( .A(n655), .B(n646), .Z(n669) );
  OR U583 ( .A(B[217]), .B(A[217]), .Z(n646) );
  AND U584 ( .A(B[217]), .B(A[217]), .Z(n655) );
  NANDN U585 ( .A(n657), .B(n670), .Z(n668) );
  NAND U586 ( .A(n642), .B(n645), .Z(n670) );
  XNOR U587 ( .A(n642), .B(n671), .Z(SUM[216]) );
  NANDN U588 ( .A(n657), .B(n645), .Z(n671) );
  OR U589 ( .A(B[216]), .B(A[216]), .Z(n645) );
  AND U590 ( .A(B[216]), .B(A[216]), .Z(n657) );
  NANDN U591 ( .A(n623), .B(n672), .Z(n642) );
  OR U592 ( .A(n627), .B(n673), .Z(n672) );
  NAND U593 ( .A(n674), .B(n675), .Z(n627) );
  AND U594 ( .A(n676), .B(n677), .Z(n675) );
  AND U595 ( .A(n678), .B(n679), .Z(n674) );
  NANDN U596 ( .A(n680), .B(n681), .Z(n623) );
  NAND U597 ( .A(n682), .B(n679), .Z(n681) );
  NANDN U598 ( .A(n683), .B(n684), .Z(n682) );
  NAND U599 ( .A(n685), .B(n678), .Z(n684) );
  NANDN U600 ( .A(n686), .B(n687), .Z(n685) );
  NAND U601 ( .A(n677), .B(n688), .Z(n687) );
  XOR U602 ( .A(n689), .B(n690), .Z(SUM[215]) );
  NANDN U603 ( .A(n680), .B(n679), .Z(n690) );
  OR U604 ( .A(B[215]), .B(A[215]), .Z(n679) );
  AND U605 ( .A(B[215]), .B(A[215]), .Z(n680) );
  ANDN U606 ( .B(n691), .A(n683), .Z(n689) );
  NAND U607 ( .A(n692), .B(n678), .Z(n691) );
  XNOR U608 ( .A(n692), .B(n693), .Z(SUM[214]) );
  NANDN U609 ( .A(n683), .B(n678), .Z(n693) );
  OR U610 ( .A(A[214]), .B(B[214]), .Z(n678) );
  AND U611 ( .A(A[214]), .B(B[214]), .Z(n683) );
  NANDN U612 ( .A(n686), .B(n694), .Z(n692) );
  NAND U613 ( .A(n695), .B(n677), .Z(n694) );
  XNOR U614 ( .A(n695), .B(n696), .Z(SUM[213]) );
  NANDN U615 ( .A(n686), .B(n677), .Z(n696) );
  OR U616 ( .A(A[213]), .B(B[213]), .Z(n677) );
  AND U617 ( .A(A[213]), .B(B[213]), .Z(n686) );
  NANDN U618 ( .A(n688), .B(n697), .Z(n695) );
  NANDN U619 ( .A(n673), .B(n676), .Z(n697) );
  XOR U620 ( .A(n673), .B(n698), .Z(SUM[212]) );
  NANDN U621 ( .A(n688), .B(n676), .Z(n698) );
  OR U622 ( .A(A[212]), .B(B[212]), .Z(n676) );
  AND U623 ( .A(A[212]), .B(B[212]), .Z(n688) );
  NOR U624 ( .A(n628), .B(n629), .Z(n673) );
  AND U625 ( .A(n699), .B(n700), .Z(n629) );
  AND U626 ( .A(n701), .B(n702), .Z(n700) );
  NOR U627 ( .A(n703), .B(n704), .Z(n702) );
  AND U628 ( .A(n705), .B(n706), .Z(n699) );
  NANDN U629 ( .A(n707), .B(n708), .Z(n628) );
  NAND U630 ( .A(n709), .B(n706), .Z(n708) );
  NANDN U631 ( .A(n710), .B(n711), .Z(n709) );
  NAND U632 ( .A(n712), .B(n705), .Z(n711) );
  NANDN U633 ( .A(n713), .B(n714), .Z(n712) );
  NAND U634 ( .A(n701), .B(n715), .Z(n714) );
  XOR U635 ( .A(n716), .B(n717), .Z(SUM[211]) );
  NANDN U636 ( .A(n707), .B(n706), .Z(n717) );
  OR U637 ( .A(B[211]), .B(A[211]), .Z(n706) );
  AND U638 ( .A(B[211]), .B(A[211]), .Z(n707) );
  ANDN U639 ( .B(n718), .A(n710), .Z(n716) );
  NAND U640 ( .A(n719), .B(n705), .Z(n718) );
  XNOR U641 ( .A(n719), .B(n720), .Z(SUM[210]) );
  NANDN U642 ( .A(n710), .B(n705), .Z(n720) );
  OR U643 ( .A(A[210]), .B(B[210]), .Z(n705) );
  AND U644 ( .A(A[210]), .B(B[210]), .Z(n710) );
  NANDN U645 ( .A(n713), .B(n721), .Z(n719) );
  NAND U646 ( .A(n722), .B(n701), .Z(n721) );
  XOR U647 ( .A(n423), .B(n723), .Z(SUM[20]) );
  NANDN U648 ( .A(n659), .B(n661), .Z(n723) );
  ANDN U649 ( .B(n724), .A(n725), .Z(n423) );
  NANDN U650 ( .A(n726), .B(n727), .Z(n724) );
  XNOR U651 ( .A(n722), .B(n728), .Z(SUM[209]) );
  NANDN U652 ( .A(n713), .B(n701), .Z(n728) );
  OR U653 ( .A(A[209]), .B(B[209]), .Z(n701) );
  AND U654 ( .A(A[209]), .B(B[209]), .Z(n713) );
  NANDN U655 ( .A(n715), .B(n729), .Z(n722) );
  OR U656 ( .A(n703), .B(n704), .Z(n729) );
  XOR U657 ( .A(n703), .B(n730), .Z(SUM[208]) );
  OR U658 ( .A(n704), .B(n715), .Z(n730) );
  AND U659 ( .A(A[208]), .B(B[208]), .Z(n715) );
  NOR U660 ( .A(B[208]), .B(A[208]), .Z(n704) );
  ANDN U661 ( .B(n731), .A(n732), .Z(n703) );
  NANDN U662 ( .A(n733), .B(n734), .Z(n731) );
  NANDN U663 ( .A(n735), .B(n736), .Z(n734) );
  NANDN U664 ( .A(n737), .B(n738), .Z(n736) );
  NANDN U665 ( .A(n739), .B(n740), .Z(n738) );
  NANDN U666 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U667 ( .A(n743), .B(n744), .Z(n742) );
  NANDN U668 ( .A(n745), .B(n746), .Z(n744) );
  NANDN U669 ( .A(n747), .B(n748), .Z(n746) );
  NANDN U670 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U671 ( .A(n751), .B(n752), .Z(n750) );
  AND U672 ( .A(n753), .B(n754), .Z(n752) );
  NANDN U673 ( .A(n755), .B(n756), .Z(n754) );
  NANDN U674 ( .A(n755), .B(n757), .Z(n753) );
  XOR U675 ( .A(n758), .B(n759), .Z(SUM[207]) );
  OR U676 ( .A(n733), .B(n732), .Z(n759) );
  AND U677 ( .A(B[207]), .B(A[207]), .Z(n732) );
  NOR U678 ( .A(B[207]), .B(A[207]), .Z(n733) );
  ANDN U679 ( .B(n760), .A(n735), .Z(n758) );
  NANDN U680 ( .A(n737), .B(n761), .Z(n760) );
  XNOR U681 ( .A(n761), .B(n762), .Z(SUM[206]) );
  OR U682 ( .A(n737), .B(n735), .Z(n762) );
  AND U683 ( .A(B[206]), .B(A[206]), .Z(n735) );
  NOR U684 ( .A(B[206]), .B(A[206]), .Z(n737) );
  NANDN U685 ( .A(n739), .B(n763), .Z(n761) );
  NANDN U686 ( .A(n741), .B(n764), .Z(n763) );
  XNOR U687 ( .A(n764), .B(n765), .Z(SUM[205]) );
  OR U688 ( .A(n741), .B(n739), .Z(n765) );
  AND U689 ( .A(B[205]), .B(A[205]), .Z(n739) );
  NOR U690 ( .A(B[205]), .B(A[205]), .Z(n741) );
  NANDN U691 ( .A(n743), .B(n766), .Z(n764) );
  NANDN U692 ( .A(n745), .B(n767), .Z(n766) );
  XNOR U693 ( .A(n767), .B(n768), .Z(SUM[204]) );
  OR U694 ( .A(n745), .B(n743), .Z(n768) );
  AND U695 ( .A(B[204]), .B(A[204]), .Z(n743) );
  NOR U696 ( .A(B[204]), .B(A[204]), .Z(n745) );
  NANDN U697 ( .A(n747), .B(n769), .Z(n767) );
  NANDN U698 ( .A(n749), .B(n770), .Z(n769) );
  NAND U699 ( .A(n771), .B(n772), .Z(n749) );
  AND U700 ( .A(n773), .B(n774), .Z(n772) );
  AND U701 ( .A(n775), .B(n776), .Z(n771) );
  NANDN U702 ( .A(n777), .B(n778), .Z(n747) );
  NAND U703 ( .A(n779), .B(n776), .Z(n778) );
  NANDN U704 ( .A(n780), .B(n781), .Z(n779) );
  NAND U705 ( .A(n782), .B(n775), .Z(n781) );
  NANDN U706 ( .A(n783), .B(n784), .Z(n782) );
  NAND U707 ( .A(n774), .B(n785), .Z(n784) );
  XOR U708 ( .A(n786), .B(n787), .Z(SUM[203]) );
  NANDN U709 ( .A(n777), .B(n776), .Z(n787) );
  OR U710 ( .A(B[203]), .B(A[203]), .Z(n776) );
  AND U711 ( .A(B[203]), .B(A[203]), .Z(n777) );
  ANDN U712 ( .B(n788), .A(n780), .Z(n786) );
  NAND U713 ( .A(n789), .B(n775), .Z(n788) );
  XNOR U714 ( .A(n789), .B(n790), .Z(SUM[202]) );
  NANDN U715 ( .A(n780), .B(n775), .Z(n790) );
  OR U716 ( .A(B[202]), .B(A[202]), .Z(n775) );
  AND U717 ( .A(B[202]), .B(A[202]), .Z(n780) );
  NANDN U718 ( .A(n783), .B(n791), .Z(n789) );
  NAND U719 ( .A(n792), .B(n774), .Z(n791) );
  XNOR U720 ( .A(n792), .B(n793), .Z(SUM[201]) );
  NANDN U721 ( .A(n783), .B(n774), .Z(n793) );
  OR U722 ( .A(B[201]), .B(A[201]), .Z(n774) );
  AND U723 ( .A(B[201]), .B(A[201]), .Z(n783) );
  NANDN U724 ( .A(n785), .B(n794), .Z(n792) );
  NAND U725 ( .A(n770), .B(n773), .Z(n794) );
  XNOR U726 ( .A(n770), .B(n795), .Z(SUM[200]) );
  NANDN U727 ( .A(n785), .B(n773), .Z(n795) );
  OR U728 ( .A(B[200]), .B(A[200]), .Z(n773) );
  AND U729 ( .A(B[200]), .B(A[200]), .Z(n785) );
  NANDN U730 ( .A(n751), .B(n796), .Z(n770) );
  OR U731 ( .A(n755), .B(n797), .Z(n796) );
  NAND U732 ( .A(n798), .B(n799), .Z(n755) );
  AND U733 ( .A(n800), .B(n801), .Z(n799) );
  AND U734 ( .A(n802), .B(n803), .Z(n798) );
  NANDN U735 ( .A(n804), .B(n805), .Z(n751) );
  NAND U736 ( .A(n806), .B(n803), .Z(n805) );
  NANDN U737 ( .A(n807), .B(n808), .Z(n806) );
  NAND U738 ( .A(n809), .B(n802), .Z(n808) );
  NANDN U739 ( .A(n810), .B(n811), .Z(n809) );
  NAND U740 ( .A(n801), .B(n812), .Z(n811) );
  XOR U741 ( .A(n813), .B(n814), .Z(SUM[19]) );
  NANDN U742 ( .A(n815), .B(n816), .Z(n814) );
  ANDN U743 ( .B(n817), .A(n818), .Z(n813) );
  NANDN U744 ( .A(n819), .B(n820), .Z(n817) );
  XOR U745 ( .A(n821), .B(n822), .Z(SUM[199]) );
  NANDN U746 ( .A(n804), .B(n803), .Z(n822) );
  OR U747 ( .A(B[199]), .B(A[199]), .Z(n803) );
  AND U748 ( .A(B[199]), .B(A[199]), .Z(n804) );
  ANDN U749 ( .B(n823), .A(n807), .Z(n821) );
  NAND U750 ( .A(n824), .B(n802), .Z(n823) );
  XNOR U751 ( .A(n824), .B(n825), .Z(SUM[198]) );
  NANDN U752 ( .A(n807), .B(n802), .Z(n825) );
  OR U753 ( .A(A[198]), .B(B[198]), .Z(n802) );
  AND U754 ( .A(A[198]), .B(B[198]), .Z(n807) );
  NANDN U755 ( .A(n810), .B(n826), .Z(n824) );
  NAND U756 ( .A(n827), .B(n801), .Z(n826) );
  XNOR U757 ( .A(n827), .B(n828), .Z(SUM[197]) );
  NANDN U758 ( .A(n810), .B(n801), .Z(n828) );
  OR U759 ( .A(A[197]), .B(B[197]), .Z(n801) );
  AND U760 ( .A(A[197]), .B(B[197]), .Z(n810) );
  NANDN U761 ( .A(n812), .B(n829), .Z(n827) );
  NANDN U762 ( .A(n797), .B(n800), .Z(n829) );
  XOR U763 ( .A(n797), .B(n830), .Z(SUM[196]) );
  NANDN U764 ( .A(n812), .B(n800), .Z(n830) );
  OR U765 ( .A(A[196]), .B(B[196]), .Z(n800) );
  AND U766 ( .A(A[196]), .B(B[196]), .Z(n812) );
  NOR U767 ( .A(n756), .B(n757), .Z(n797) );
  AND U768 ( .A(n831), .B(n832), .Z(n757) );
  AND U769 ( .A(n833), .B(n834), .Z(n832) );
  NOR U770 ( .A(n835), .B(n836), .Z(n834) );
  AND U771 ( .A(n837), .B(n838), .Z(n831) );
  NANDN U772 ( .A(n839), .B(n840), .Z(n756) );
  NAND U773 ( .A(n841), .B(n838), .Z(n840) );
  NANDN U774 ( .A(n842), .B(n843), .Z(n841) );
  NAND U775 ( .A(n844), .B(n837), .Z(n843) );
  NANDN U776 ( .A(n845), .B(n846), .Z(n844) );
  NAND U777 ( .A(n833), .B(n847), .Z(n846) );
  XOR U778 ( .A(n848), .B(n849), .Z(SUM[195]) );
  NANDN U779 ( .A(n839), .B(n838), .Z(n849) );
  OR U780 ( .A(B[195]), .B(A[195]), .Z(n838) );
  AND U781 ( .A(B[195]), .B(A[195]), .Z(n839) );
  ANDN U782 ( .B(n850), .A(n842), .Z(n848) );
  NAND U783 ( .A(n851), .B(n837), .Z(n850) );
  XNOR U784 ( .A(n851), .B(n852), .Z(SUM[194]) );
  NANDN U785 ( .A(n842), .B(n837), .Z(n852) );
  OR U786 ( .A(A[194]), .B(B[194]), .Z(n837) );
  AND U787 ( .A(A[194]), .B(B[194]), .Z(n842) );
  NANDN U788 ( .A(n845), .B(n853), .Z(n851) );
  NAND U789 ( .A(n854), .B(n833), .Z(n853) );
  XNOR U790 ( .A(n854), .B(n855), .Z(SUM[193]) );
  NANDN U791 ( .A(n845), .B(n833), .Z(n855) );
  OR U792 ( .A(A[193]), .B(B[193]), .Z(n833) );
  AND U793 ( .A(A[193]), .B(B[193]), .Z(n845) );
  NANDN U794 ( .A(n847), .B(n856), .Z(n854) );
  OR U795 ( .A(n835), .B(n836), .Z(n856) );
  XOR U796 ( .A(n835), .B(n857), .Z(SUM[192]) );
  OR U797 ( .A(n836), .B(n847), .Z(n857) );
  AND U798 ( .A(A[192]), .B(B[192]), .Z(n847) );
  NOR U799 ( .A(B[192]), .B(A[192]), .Z(n836) );
  ANDN U800 ( .B(n858), .A(n859), .Z(n835) );
  NANDN U801 ( .A(n860), .B(n861), .Z(n858) );
  NANDN U802 ( .A(n862), .B(n863), .Z(n861) );
  NANDN U803 ( .A(n864), .B(n865), .Z(n863) );
  NANDN U804 ( .A(n866), .B(n867), .Z(n865) );
  NANDN U805 ( .A(n868), .B(n869), .Z(n867) );
  NAND U806 ( .A(n870), .B(n871), .Z(n869) );
  NAND U807 ( .A(n872), .B(n873), .Z(n871) );
  AND U808 ( .A(n874), .B(n875), .Z(n873) );
  ANDN U809 ( .B(n876), .A(n877), .Z(n875) );
  NOR U810 ( .A(n878), .B(n879), .Z(n872) );
  ANDN U811 ( .B(n880), .A(n881), .Z(n870) );
  NAND U812 ( .A(n882), .B(n876), .Z(n880) );
  NANDN U813 ( .A(n883), .B(n884), .Z(n882) );
  NANDN U814 ( .A(n879), .B(n885), .Z(n884) );
  NANDN U815 ( .A(n886), .B(n887), .Z(n885) );
  NAND U816 ( .A(n888), .B(n874), .Z(n887) );
  XOR U817 ( .A(n889), .B(n890), .Z(SUM[191]) );
  OR U818 ( .A(n860), .B(n859), .Z(n890) );
  AND U819 ( .A(B[191]), .B(A[191]), .Z(n859) );
  NOR U820 ( .A(B[191]), .B(A[191]), .Z(n860) );
  ANDN U821 ( .B(n891), .A(n862), .Z(n889) );
  NANDN U822 ( .A(n864), .B(n892), .Z(n891) );
  XNOR U823 ( .A(n892), .B(n893), .Z(SUM[190]) );
  OR U824 ( .A(n864), .B(n862), .Z(n893) );
  AND U825 ( .A(B[190]), .B(A[190]), .Z(n862) );
  NOR U826 ( .A(B[190]), .B(A[190]), .Z(n864) );
  NANDN U827 ( .A(n866), .B(n894), .Z(n892) );
  NANDN U828 ( .A(n868), .B(n895), .Z(n894) );
  XNOR U829 ( .A(n820), .B(n896), .Z(SUM[18]) );
  OR U830 ( .A(n819), .B(n818), .Z(n896) );
  NANDN U831 ( .A(n897), .B(n898), .Z(n820) );
  NAND U832 ( .A(n899), .B(n900), .Z(n898) );
  XNOR U833 ( .A(n895), .B(n901), .Z(SUM[189]) );
  OR U834 ( .A(n868), .B(n866), .Z(n901) );
  AND U835 ( .A(B[189]), .B(A[189]), .Z(n866) );
  NOR U836 ( .A(B[189]), .B(A[189]), .Z(n868) );
  NANDN U837 ( .A(n881), .B(n902), .Z(n895) );
  NAND U838 ( .A(n903), .B(n876), .Z(n902) );
  XNOR U839 ( .A(n903), .B(n904), .Z(SUM[188]) );
  NANDN U840 ( .A(n881), .B(n876), .Z(n904) );
  OR U841 ( .A(A[188]), .B(B[188]), .Z(n876) );
  AND U842 ( .A(B[188]), .B(A[188]), .Z(n881) );
  NANDN U843 ( .A(n883), .B(n905), .Z(n903) );
  NANDN U844 ( .A(n879), .B(n906), .Z(n905) );
  NAND U845 ( .A(n907), .B(n908), .Z(n879) );
  AND U846 ( .A(n909), .B(n910), .Z(n908) );
  AND U847 ( .A(n911), .B(n912), .Z(n907) );
  NANDN U848 ( .A(n913), .B(n914), .Z(n883) );
  NAND U849 ( .A(n915), .B(n912), .Z(n914) );
  NANDN U850 ( .A(n916), .B(n917), .Z(n915) );
  NAND U851 ( .A(n918), .B(n911), .Z(n917) );
  NANDN U852 ( .A(n919), .B(n920), .Z(n918) );
  NAND U853 ( .A(n910), .B(n921), .Z(n920) );
  XOR U854 ( .A(n922), .B(n923), .Z(SUM[187]) );
  NANDN U855 ( .A(n913), .B(n912), .Z(n923) );
  OR U856 ( .A(B[187]), .B(A[187]), .Z(n912) );
  AND U857 ( .A(B[187]), .B(A[187]), .Z(n913) );
  ANDN U858 ( .B(n924), .A(n916), .Z(n922) );
  NAND U859 ( .A(n925), .B(n911), .Z(n924) );
  XNOR U860 ( .A(n925), .B(n926), .Z(SUM[186]) );
  NANDN U861 ( .A(n916), .B(n911), .Z(n926) );
  OR U862 ( .A(B[186]), .B(A[186]), .Z(n911) );
  AND U863 ( .A(B[186]), .B(A[186]), .Z(n916) );
  NANDN U864 ( .A(n919), .B(n927), .Z(n925) );
  NAND U865 ( .A(n928), .B(n910), .Z(n927) );
  XNOR U866 ( .A(n928), .B(n929), .Z(SUM[185]) );
  NANDN U867 ( .A(n919), .B(n910), .Z(n929) );
  OR U868 ( .A(B[185]), .B(A[185]), .Z(n910) );
  AND U869 ( .A(B[185]), .B(A[185]), .Z(n919) );
  NANDN U870 ( .A(n921), .B(n930), .Z(n928) );
  NAND U871 ( .A(n906), .B(n909), .Z(n930) );
  XNOR U872 ( .A(n906), .B(n931), .Z(SUM[184]) );
  NANDN U873 ( .A(n921), .B(n909), .Z(n931) );
  OR U874 ( .A(B[184]), .B(A[184]), .Z(n909) );
  AND U875 ( .A(B[184]), .B(A[184]), .Z(n921) );
  NANDN U876 ( .A(n886), .B(n932), .Z(n906) );
  NANDN U877 ( .A(n933), .B(n874), .Z(n932) );
  AND U878 ( .A(n934), .B(n935), .Z(n874) );
  AND U879 ( .A(n936), .B(n937), .Z(n935) );
  AND U880 ( .A(n938), .B(n939), .Z(n934) );
  NANDN U881 ( .A(n940), .B(n941), .Z(n886) );
  NAND U882 ( .A(n942), .B(n939), .Z(n941) );
  NANDN U883 ( .A(n943), .B(n944), .Z(n942) );
  NAND U884 ( .A(n945), .B(n938), .Z(n944) );
  NANDN U885 ( .A(n946), .B(n947), .Z(n945) );
  NAND U886 ( .A(n937), .B(n948), .Z(n947) );
  XOR U887 ( .A(n949), .B(n950), .Z(SUM[183]) );
  NANDN U888 ( .A(n940), .B(n939), .Z(n950) );
  OR U889 ( .A(B[183]), .B(A[183]), .Z(n939) );
  AND U890 ( .A(B[183]), .B(A[183]), .Z(n940) );
  ANDN U891 ( .B(n951), .A(n943), .Z(n949) );
  NAND U892 ( .A(n952), .B(n938), .Z(n951) );
  XNOR U893 ( .A(n952), .B(n953), .Z(SUM[182]) );
  NANDN U894 ( .A(n943), .B(n938), .Z(n953) );
  OR U895 ( .A(B[182]), .B(A[182]), .Z(n938) );
  AND U896 ( .A(B[182]), .B(A[182]), .Z(n943) );
  NANDN U897 ( .A(n946), .B(n954), .Z(n952) );
  NAND U898 ( .A(n955), .B(n937), .Z(n954) );
  XNOR U899 ( .A(n955), .B(n956), .Z(SUM[181]) );
  NANDN U900 ( .A(n946), .B(n937), .Z(n956) );
  OR U901 ( .A(B[181]), .B(A[181]), .Z(n937) );
  AND U902 ( .A(B[181]), .B(A[181]), .Z(n946) );
  NANDN U903 ( .A(n948), .B(n957), .Z(n955) );
  NANDN U904 ( .A(n933), .B(n936), .Z(n957) );
  XOR U905 ( .A(n933), .B(n958), .Z(SUM[180]) );
  NANDN U906 ( .A(n948), .B(n936), .Z(n958) );
  OR U907 ( .A(B[180]), .B(A[180]), .Z(n936) );
  AND U908 ( .A(B[180]), .B(A[180]), .Z(n948) );
  ANDN U909 ( .B(n959), .A(n888), .Z(n933) );
  NANDN U910 ( .A(n960), .B(n961), .Z(n888) );
  NAND U911 ( .A(n962), .B(n963), .Z(n961) );
  NANDN U912 ( .A(n964), .B(n965), .Z(n962) );
  NANDN U913 ( .A(n966), .B(n967), .Z(n965) );
  NANDN U914 ( .A(n968), .B(n969), .Z(n967) );
  NAND U915 ( .A(n970), .B(n971), .Z(n969) );
  OR U916 ( .A(n878), .B(n877), .Z(n959) );
  NAND U917 ( .A(n972), .B(n973), .Z(n878) );
  AND U918 ( .A(n974), .B(n970), .Z(n973) );
  ANDN U919 ( .B(n963), .A(n966), .Z(n972) );
  XNOR U920 ( .A(n899), .B(n975), .Z(SUM[17]) );
  NANDN U921 ( .A(n897), .B(n900), .Z(n975) );
  NANDN U922 ( .A(n976), .B(n977), .Z(n899) );
  NAND U923 ( .A(n978), .B(n727), .Z(n977) );
  XOR U924 ( .A(n979), .B(n980), .Z(SUM[179]) );
  NANDN U925 ( .A(n960), .B(n963), .Z(n980) );
  OR U926 ( .A(B[179]), .B(A[179]), .Z(n963) );
  AND U927 ( .A(B[179]), .B(A[179]), .Z(n960) );
  ANDN U928 ( .B(n981), .A(n964), .Z(n979) );
  NANDN U929 ( .A(n966), .B(n982), .Z(n981) );
  XNOR U930 ( .A(n982), .B(n983), .Z(SUM[178]) );
  OR U931 ( .A(n966), .B(n964), .Z(n983) );
  AND U932 ( .A(B[178]), .B(A[178]), .Z(n964) );
  NOR U933 ( .A(B[178]), .B(A[178]), .Z(n966) );
  NANDN U934 ( .A(n968), .B(n984), .Z(n982) );
  NAND U935 ( .A(n985), .B(n970), .Z(n984) );
  XNOR U936 ( .A(n985), .B(n986), .Z(SUM[177]) );
  NANDN U937 ( .A(n968), .B(n970), .Z(n986) );
  OR U938 ( .A(B[177]), .B(A[177]), .Z(n970) );
  AND U939 ( .A(B[177]), .B(A[177]), .Z(n968) );
  NANDN U940 ( .A(n971), .B(n987), .Z(n985) );
  NANDN U941 ( .A(n877), .B(n974), .Z(n987) );
  XOR U942 ( .A(n877), .B(n988), .Z(SUM[176]) );
  NANDN U943 ( .A(n971), .B(n974), .Z(n988) );
  OR U944 ( .A(B[176]), .B(A[176]), .Z(n974) );
  AND U945 ( .A(A[176]), .B(B[176]), .Z(n971) );
  ANDN U946 ( .B(n989), .A(n990), .Z(n877) );
  NANDN U947 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U948 ( .A(n993), .B(n994), .Z(n992) );
  NANDN U949 ( .A(n995), .B(n996), .Z(n994) );
  NANDN U950 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U951 ( .A(n999), .B(n1000), .Z(n998) );
  NAND U952 ( .A(n1001), .B(n1002), .Z(n1000) );
  NAND U953 ( .A(n1003), .B(n1004), .Z(n1002) );
  AND U954 ( .A(n1005), .B(n1006), .Z(n1004) );
  ANDN U955 ( .B(n1007), .A(n1008), .Z(n1006) );
  NOR U956 ( .A(n1009), .B(n1010), .Z(n1003) );
  ANDN U957 ( .B(n1011), .A(n1012), .Z(n1001) );
  NAND U958 ( .A(n1013), .B(n1007), .Z(n1011) );
  NANDN U959 ( .A(n1014), .B(n1015), .Z(n1013) );
  NANDN U960 ( .A(n1010), .B(n1016), .Z(n1015) );
  NANDN U961 ( .A(n1017), .B(n1018), .Z(n1016) );
  NAND U962 ( .A(n1019), .B(n1005), .Z(n1018) );
  XOR U963 ( .A(n1020), .B(n1021), .Z(SUM[175]) );
  OR U964 ( .A(n991), .B(n990), .Z(n1021) );
  AND U965 ( .A(B[175]), .B(A[175]), .Z(n990) );
  NOR U966 ( .A(B[175]), .B(A[175]), .Z(n991) );
  ANDN U967 ( .B(n1022), .A(n993), .Z(n1020) );
  NANDN U968 ( .A(n995), .B(n1023), .Z(n1022) );
  XNOR U969 ( .A(n1023), .B(n1024), .Z(SUM[174]) );
  OR U970 ( .A(n995), .B(n993), .Z(n1024) );
  AND U971 ( .A(B[174]), .B(A[174]), .Z(n993) );
  NOR U972 ( .A(B[174]), .B(A[174]), .Z(n995) );
  NANDN U973 ( .A(n997), .B(n1025), .Z(n1023) );
  NANDN U974 ( .A(n999), .B(n1026), .Z(n1025) );
  XNOR U975 ( .A(n1026), .B(n1027), .Z(SUM[173]) );
  OR U976 ( .A(n999), .B(n997), .Z(n1027) );
  AND U977 ( .A(B[173]), .B(A[173]), .Z(n997) );
  NOR U978 ( .A(B[173]), .B(A[173]), .Z(n999) );
  NANDN U979 ( .A(n1012), .B(n1028), .Z(n1026) );
  NAND U980 ( .A(n1029), .B(n1007), .Z(n1028) );
  XNOR U981 ( .A(n1029), .B(n1030), .Z(SUM[172]) );
  NANDN U982 ( .A(n1012), .B(n1007), .Z(n1030) );
  OR U983 ( .A(A[172]), .B(B[172]), .Z(n1007) );
  AND U984 ( .A(B[172]), .B(A[172]), .Z(n1012) );
  NANDN U985 ( .A(n1014), .B(n1031), .Z(n1029) );
  NANDN U986 ( .A(n1010), .B(n1032), .Z(n1031) );
  NAND U987 ( .A(n1033), .B(n1034), .Z(n1010) );
  AND U988 ( .A(n1035), .B(n1036), .Z(n1034) );
  AND U989 ( .A(n1037), .B(n1038), .Z(n1033) );
  NANDN U990 ( .A(n1039), .B(n1040), .Z(n1014) );
  NAND U991 ( .A(n1041), .B(n1038), .Z(n1040) );
  NANDN U992 ( .A(n1042), .B(n1043), .Z(n1041) );
  NAND U993 ( .A(n1044), .B(n1037), .Z(n1043) );
  NANDN U994 ( .A(n1045), .B(n1046), .Z(n1044) );
  NAND U995 ( .A(n1036), .B(n1047), .Z(n1046) );
  XOR U996 ( .A(n1048), .B(n1049), .Z(SUM[171]) );
  NANDN U997 ( .A(n1039), .B(n1038), .Z(n1049) );
  OR U998 ( .A(B[171]), .B(A[171]), .Z(n1038) );
  AND U999 ( .A(B[171]), .B(A[171]), .Z(n1039) );
  ANDN U1000 ( .B(n1050), .A(n1042), .Z(n1048) );
  NAND U1001 ( .A(n1051), .B(n1037), .Z(n1050) );
  XNOR U1002 ( .A(n1051), .B(n1052), .Z(SUM[170]) );
  NANDN U1003 ( .A(n1042), .B(n1037), .Z(n1052) );
  OR U1004 ( .A(B[170]), .B(A[170]), .Z(n1037) );
  AND U1005 ( .A(B[170]), .B(A[170]), .Z(n1042) );
  NANDN U1006 ( .A(n1045), .B(n1053), .Z(n1051) );
  NAND U1007 ( .A(n1054), .B(n1036), .Z(n1053) );
  XOR U1008 ( .A(n727), .B(n1055), .Z(SUM[16]) );
  ANDN U1009 ( .B(n978), .A(n976), .Z(n1055) );
  XNOR U1010 ( .A(n1054), .B(n1056), .Z(SUM[169]) );
  NANDN U1011 ( .A(n1045), .B(n1036), .Z(n1056) );
  OR U1012 ( .A(B[169]), .B(A[169]), .Z(n1036) );
  AND U1013 ( .A(B[169]), .B(A[169]), .Z(n1045) );
  NANDN U1014 ( .A(n1047), .B(n1057), .Z(n1054) );
  NAND U1015 ( .A(n1032), .B(n1035), .Z(n1057) );
  XNOR U1016 ( .A(n1032), .B(n1058), .Z(SUM[168]) );
  NANDN U1017 ( .A(n1047), .B(n1035), .Z(n1058) );
  OR U1018 ( .A(B[168]), .B(A[168]), .Z(n1035) );
  AND U1019 ( .A(B[168]), .B(A[168]), .Z(n1047) );
  NANDN U1020 ( .A(n1017), .B(n1059), .Z(n1032) );
  NANDN U1021 ( .A(n1060), .B(n1005), .Z(n1059) );
  AND U1022 ( .A(n1061), .B(n1062), .Z(n1005) );
  AND U1023 ( .A(n1063), .B(n1064), .Z(n1062) );
  AND U1024 ( .A(n1065), .B(n1066), .Z(n1061) );
  NANDN U1025 ( .A(n1067), .B(n1068), .Z(n1017) );
  NAND U1026 ( .A(n1069), .B(n1066), .Z(n1068) );
  NANDN U1027 ( .A(n1070), .B(n1071), .Z(n1069) );
  NAND U1028 ( .A(n1072), .B(n1065), .Z(n1071) );
  NANDN U1029 ( .A(n1073), .B(n1074), .Z(n1072) );
  NAND U1030 ( .A(n1064), .B(n1075), .Z(n1074) );
  XOR U1031 ( .A(n1076), .B(n1077), .Z(SUM[167]) );
  NANDN U1032 ( .A(n1067), .B(n1066), .Z(n1077) );
  OR U1033 ( .A(B[167]), .B(A[167]), .Z(n1066) );
  AND U1034 ( .A(B[167]), .B(A[167]), .Z(n1067) );
  ANDN U1035 ( .B(n1078), .A(n1070), .Z(n1076) );
  NAND U1036 ( .A(n1079), .B(n1065), .Z(n1078) );
  XNOR U1037 ( .A(n1079), .B(n1080), .Z(SUM[166]) );
  NANDN U1038 ( .A(n1070), .B(n1065), .Z(n1080) );
  OR U1039 ( .A(B[166]), .B(A[166]), .Z(n1065) );
  AND U1040 ( .A(B[166]), .B(A[166]), .Z(n1070) );
  NANDN U1041 ( .A(n1073), .B(n1081), .Z(n1079) );
  NAND U1042 ( .A(n1082), .B(n1064), .Z(n1081) );
  XNOR U1043 ( .A(n1082), .B(n1083), .Z(SUM[165]) );
  NANDN U1044 ( .A(n1073), .B(n1064), .Z(n1083) );
  OR U1045 ( .A(B[165]), .B(A[165]), .Z(n1064) );
  AND U1046 ( .A(B[165]), .B(A[165]), .Z(n1073) );
  NANDN U1047 ( .A(n1075), .B(n1084), .Z(n1082) );
  NANDN U1048 ( .A(n1060), .B(n1063), .Z(n1084) );
  XOR U1049 ( .A(n1060), .B(n1085), .Z(SUM[164]) );
  NANDN U1050 ( .A(n1075), .B(n1063), .Z(n1085) );
  OR U1051 ( .A(B[164]), .B(A[164]), .Z(n1063) );
  AND U1052 ( .A(B[164]), .B(A[164]), .Z(n1075) );
  ANDN U1053 ( .B(n1086), .A(n1019), .Z(n1060) );
  NANDN U1054 ( .A(n1087), .B(n1088), .Z(n1019) );
  NAND U1055 ( .A(n1089), .B(n1090), .Z(n1088) );
  NANDN U1056 ( .A(n1091), .B(n1092), .Z(n1089) );
  NANDN U1057 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1058 ( .A(n1095), .B(n1096), .Z(n1094) );
  NAND U1059 ( .A(n1097), .B(n1098), .Z(n1096) );
  OR U1060 ( .A(n1009), .B(n1008), .Z(n1086) );
  NAND U1061 ( .A(n1099), .B(n1100), .Z(n1009) );
  AND U1062 ( .A(n1101), .B(n1097), .Z(n1100) );
  ANDN U1063 ( .B(n1090), .A(n1093), .Z(n1099) );
  XOR U1064 ( .A(n1102), .B(n1103), .Z(SUM[163]) );
  NANDN U1065 ( .A(n1087), .B(n1090), .Z(n1103) );
  OR U1066 ( .A(B[163]), .B(A[163]), .Z(n1090) );
  AND U1067 ( .A(B[163]), .B(A[163]), .Z(n1087) );
  ANDN U1068 ( .B(n1104), .A(n1091), .Z(n1102) );
  NANDN U1069 ( .A(n1093), .B(n1105), .Z(n1104) );
  XNOR U1070 ( .A(n1105), .B(n1106), .Z(SUM[162]) );
  OR U1071 ( .A(n1093), .B(n1091), .Z(n1106) );
  AND U1072 ( .A(B[162]), .B(A[162]), .Z(n1091) );
  NOR U1073 ( .A(B[162]), .B(A[162]), .Z(n1093) );
  NANDN U1074 ( .A(n1095), .B(n1107), .Z(n1105) );
  NAND U1075 ( .A(n1108), .B(n1097), .Z(n1107) );
  XNOR U1076 ( .A(n1108), .B(n1109), .Z(SUM[161]) );
  NANDN U1077 ( .A(n1095), .B(n1097), .Z(n1109) );
  OR U1078 ( .A(B[161]), .B(A[161]), .Z(n1097) );
  AND U1079 ( .A(B[161]), .B(A[161]), .Z(n1095) );
  NANDN U1080 ( .A(n1098), .B(n1110), .Z(n1108) );
  NANDN U1081 ( .A(n1008), .B(n1101), .Z(n1110) );
  XOR U1082 ( .A(n1008), .B(n1111), .Z(SUM[160]) );
  NANDN U1083 ( .A(n1098), .B(n1101), .Z(n1111) );
  OR U1084 ( .A(B[160]), .B(A[160]), .Z(n1101) );
  AND U1085 ( .A(A[160]), .B(B[160]), .Z(n1098) );
  ANDN U1086 ( .B(n1112), .A(n1113), .Z(n1008) );
  NANDN U1087 ( .A(n1114), .B(n1115), .Z(n1112) );
  NANDN U1088 ( .A(n1116), .B(n1117), .Z(n1115) );
  NANDN U1089 ( .A(n1118), .B(n1119), .Z(n1117) );
  NANDN U1090 ( .A(n1120), .B(n1121), .Z(n1119) );
  NANDN U1091 ( .A(n1122), .B(n1123), .Z(n1121) );
  NAND U1092 ( .A(n1124), .B(n1125), .Z(n1123) );
  NAND U1093 ( .A(n1126), .B(n1127), .Z(n1125) );
  AND U1094 ( .A(n1128), .B(n1129), .Z(n1127) );
  ANDN U1095 ( .B(n1130), .A(n1131), .Z(n1129) );
  NOR U1096 ( .A(n1132), .B(n1133), .Z(n1126) );
  ANDN U1097 ( .B(n1134), .A(n1135), .Z(n1124) );
  NAND U1098 ( .A(n1136), .B(n1130), .Z(n1134) );
  NANDN U1099 ( .A(n1137), .B(n1138), .Z(n1136) );
  NANDN U1100 ( .A(n1133), .B(n1139), .Z(n1138) );
  NANDN U1101 ( .A(n1140), .B(n1141), .Z(n1139) );
  NAND U1102 ( .A(n1142), .B(n1128), .Z(n1141) );
  ANDN U1103 ( .B(n1143), .A(n727), .Z(SUM[15]) );
  OR U1104 ( .A(A[15]), .B(B[15]), .Z(n1143) );
  XOR U1105 ( .A(n1144), .B(n1145), .Z(SUM[159]) );
  OR U1106 ( .A(n1114), .B(n1113), .Z(n1145) );
  AND U1107 ( .A(B[159]), .B(A[159]), .Z(n1113) );
  NOR U1108 ( .A(B[159]), .B(A[159]), .Z(n1114) );
  ANDN U1109 ( .B(n1146), .A(n1116), .Z(n1144) );
  NANDN U1110 ( .A(n1118), .B(n1147), .Z(n1146) );
  XNOR U1111 ( .A(n1147), .B(n1148), .Z(SUM[158]) );
  OR U1112 ( .A(n1118), .B(n1116), .Z(n1148) );
  AND U1113 ( .A(B[158]), .B(A[158]), .Z(n1116) );
  NOR U1114 ( .A(B[158]), .B(A[158]), .Z(n1118) );
  NANDN U1115 ( .A(n1120), .B(n1149), .Z(n1147) );
  NANDN U1116 ( .A(n1122), .B(n1150), .Z(n1149) );
  XNOR U1117 ( .A(n1150), .B(n1151), .Z(SUM[157]) );
  OR U1118 ( .A(n1122), .B(n1120), .Z(n1151) );
  AND U1119 ( .A(B[157]), .B(A[157]), .Z(n1120) );
  NOR U1120 ( .A(B[157]), .B(A[157]), .Z(n1122) );
  NANDN U1121 ( .A(n1135), .B(n1152), .Z(n1150) );
  NAND U1122 ( .A(n1153), .B(n1130), .Z(n1152) );
  XNOR U1123 ( .A(n1153), .B(n1154), .Z(SUM[156]) );
  NANDN U1124 ( .A(n1135), .B(n1130), .Z(n1154) );
  OR U1125 ( .A(A[156]), .B(B[156]), .Z(n1130) );
  AND U1126 ( .A(B[156]), .B(A[156]), .Z(n1135) );
  NANDN U1127 ( .A(n1137), .B(n1155), .Z(n1153) );
  NANDN U1128 ( .A(n1133), .B(n1156), .Z(n1155) );
  NAND U1129 ( .A(n1157), .B(n1158), .Z(n1133) );
  AND U1130 ( .A(n1159), .B(n1160), .Z(n1158) );
  AND U1131 ( .A(n1161), .B(n1162), .Z(n1157) );
  NANDN U1132 ( .A(n1163), .B(n1164), .Z(n1137) );
  NAND U1133 ( .A(n1165), .B(n1162), .Z(n1164) );
  NANDN U1134 ( .A(n1166), .B(n1167), .Z(n1165) );
  NAND U1135 ( .A(n1168), .B(n1161), .Z(n1167) );
  NANDN U1136 ( .A(n1169), .B(n1170), .Z(n1168) );
  NAND U1137 ( .A(n1160), .B(n1171), .Z(n1170) );
  XOR U1138 ( .A(n1172), .B(n1173), .Z(SUM[155]) );
  NANDN U1139 ( .A(n1163), .B(n1162), .Z(n1173) );
  OR U1140 ( .A(B[155]), .B(A[155]), .Z(n1162) );
  AND U1141 ( .A(B[155]), .B(A[155]), .Z(n1163) );
  ANDN U1142 ( .B(n1174), .A(n1166), .Z(n1172) );
  NAND U1143 ( .A(n1175), .B(n1161), .Z(n1174) );
  XNOR U1144 ( .A(n1175), .B(n1176), .Z(SUM[154]) );
  NANDN U1145 ( .A(n1166), .B(n1161), .Z(n1176) );
  OR U1146 ( .A(B[154]), .B(A[154]), .Z(n1161) );
  AND U1147 ( .A(B[154]), .B(A[154]), .Z(n1166) );
  NANDN U1148 ( .A(n1169), .B(n1177), .Z(n1175) );
  NAND U1149 ( .A(n1178), .B(n1160), .Z(n1177) );
  XNOR U1150 ( .A(n1178), .B(n1179), .Z(SUM[153]) );
  NANDN U1151 ( .A(n1169), .B(n1160), .Z(n1179) );
  OR U1152 ( .A(B[153]), .B(A[153]), .Z(n1160) );
  AND U1153 ( .A(B[153]), .B(A[153]), .Z(n1169) );
  NANDN U1154 ( .A(n1171), .B(n1180), .Z(n1178) );
  NAND U1155 ( .A(n1156), .B(n1159), .Z(n1180) );
  XNOR U1156 ( .A(n1156), .B(n1181), .Z(SUM[152]) );
  NANDN U1157 ( .A(n1171), .B(n1159), .Z(n1181) );
  OR U1158 ( .A(B[152]), .B(A[152]), .Z(n1159) );
  AND U1159 ( .A(B[152]), .B(A[152]), .Z(n1171) );
  NANDN U1160 ( .A(n1140), .B(n1182), .Z(n1156) );
  NANDN U1161 ( .A(n1183), .B(n1128), .Z(n1182) );
  AND U1162 ( .A(n1184), .B(n1185), .Z(n1128) );
  AND U1163 ( .A(n1186), .B(n1187), .Z(n1185) );
  AND U1164 ( .A(n1188), .B(n1189), .Z(n1184) );
  NANDN U1165 ( .A(n1190), .B(n1191), .Z(n1140) );
  NAND U1166 ( .A(n1192), .B(n1189), .Z(n1191) );
  NANDN U1167 ( .A(n1193), .B(n1194), .Z(n1192) );
  NAND U1168 ( .A(n1195), .B(n1188), .Z(n1194) );
  NANDN U1169 ( .A(n1196), .B(n1197), .Z(n1195) );
  NAND U1170 ( .A(n1187), .B(n1198), .Z(n1197) );
  XOR U1171 ( .A(n1199), .B(n1200), .Z(SUM[151]) );
  NANDN U1172 ( .A(n1190), .B(n1189), .Z(n1200) );
  OR U1173 ( .A(B[151]), .B(A[151]), .Z(n1189) );
  AND U1174 ( .A(B[151]), .B(A[151]), .Z(n1190) );
  ANDN U1175 ( .B(n1201), .A(n1193), .Z(n1199) );
  NAND U1176 ( .A(n1202), .B(n1188), .Z(n1201) );
  XNOR U1177 ( .A(n1202), .B(n1203), .Z(SUM[150]) );
  NANDN U1178 ( .A(n1193), .B(n1188), .Z(n1203) );
  OR U1179 ( .A(B[150]), .B(A[150]), .Z(n1188) );
  AND U1180 ( .A(B[150]), .B(A[150]), .Z(n1193) );
  NANDN U1181 ( .A(n1196), .B(n1204), .Z(n1202) );
  NAND U1182 ( .A(n1205), .B(n1187), .Z(n1204) );
  XNOR U1183 ( .A(n1205), .B(n1206), .Z(SUM[149]) );
  NANDN U1184 ( .A(n1196), .B(n1187), .Z(n1206) );
  OR U1185 ( .A(B[149]), .B(A[149]), .Z(n1187) );
  AND U1186 ( .A(B[149]), .B(A[149]), .Z(n1196) );
  NANDN U1187 ( .A(n1198), .B(n1207), .Z(n1205) );
  NANDN U1188 ( .A(n1183), .B(n1186), .Z(n1207) );
  XOR U1189 ( .A(n1183), .B(n1208), .Z(SUM[148]) );
  NANDN U1190 ( .A(n1198), .B(n1186), .Z(n1208) );
  OR U1191 ( .A(B[148]), .B(A[148]), .Z(n1186) );
  AND U1192 ( .A(B[148]), .B(A[148]), .Z(n1198) );
  ANDN U1193 ( .B(n1209), .A(n1142), .Z(n1183) );
  NANDN U1194 ( .A(n1210), .B(n1211), .Z(n1142) );
  NAND U1195 ( .A(n1212), .B(n1213), .Z(n1211) );
  NANDN U1196 ( .A(n1214), .B(n1215), .Z(n1212) );
  NANDN U1197 ( .A(n1216), .B(n1217), .Z(n1215) );
  NANDN U1198 ( .A(n1218), .B(n1219), .Z(n1217) );
  NAND U1199 ( .A(n1220), .B(n1221), .Z(n1219) );
  OR U1200 ( .A(n1132), .B(n1131), .Z(n1209) );
  NAND U1201 ( .A(n1222), .B(n1223), .Z(n1132) );
  AND U1202 ( .A(n1224), .B(n1220), .Z(n1223) );
  ANDN U1203 ( .B(n1213), .A(n1216), .Z(n1222) );
  XOR U1204 ( .A(n1225), .B(n1226), .Z(SUM[147]) );
  NANDN U1205 ( .A(n1210), .B(n1213), .Z(n1226) );
  OR U1206 ( .A(B[147]), .B(A[147]), .Z(n1213) );
  AND U1207 ( .A(B[147]), .B(A[147]), .Z(n1210) );
  ANDN U1208 ( .B(n1227), .A(n1214), .Z(n1225) );
  NANDN U1209 ( .A(n1216), .B(n1228), .Z(n1227) );
  XNOR U1210 ( .A(n1228), .B(n1229), .Z(SUM[146]) );
  OR U1211 ( .A(n1216), .B(n1214), .Z(n1229) );
  AND U1212 ( .A(B[146]), .B(A[146]), .Z(n1214) );
  NOR U1213 ( .A(B[146]), .B(A[146]), .Z(n1216) );
  NANDN U1214 ( .A(n1218), .B(n1230), .Z(n1228) );
  NAND U1215 ( .A(n1231), .B(n1220), .Z(n1230) );
  XNOR U1216 ( .A(n1231), .B(n1232), .Z(SUM[145]) );
  NANDN U1217 ( .A(n1218), .B(n1220), .Z(n1232) );
  OR U1218 ( .A(B[145]), .B(A[145]), .Z(n1220) );
  AND U1219 ( .A(B[145]), .B(A[145]), .Z(n1218) );
  NANDN U1220 ( .A(n1221), .B(n1233), .Z(n1231) );
  NANDN U1221 ( .A(n1131), .B(n1224), .Z(n1233) );
  XOR U1222 ( .A(n1131), .B(n1234), .Z(SUM[144]) );
  NANDN U1223 ( .A(n1221), .B(n1224), .Z(n1234) );
  OR U1224 ( .A(B[144]), .B(A[144]), .Z(n1224) );
  AND U1225 ( .A(A[144]), .B(B[144]), .Z(n1221) );
  ANDN U1226 ( .B(n1235), .A(n1236), .Z(n1131) );
  NANDN U1227 ( .A(n1237), .B(n1238), .Z(n1235) );
  NANDN U1228 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1229 ( .A(n1241), .B(n1242), .Z(n1240) );
  NANDN U1230 ( .A(n1243), .B(n1244), .Z(n1242) );
  NANDN U1231 ( .A(n1245), .B(n1246), .Z(n1244) );
  NAND U1232 ( .A(n1247), .B(n1248), .Z(n1246) );
  NAND U1233 ( .A(n1249), .B(n1250), .Z(n1248) );
  AND U1234 ( .A(n1251), .B(n1252), .Z(n1250) );
  ANDN U1235 ( .B(n1253), .A(n1254), .Z(n1252) );
  NOR U1236 ( .A(n1255), .B(n1256), .Z(n1249) );
  ANDN U1237 ( .B(n1257), .A(n1258), .Z(n1247) );
  NAND U1238 ( .A(n1259), .B(n1253), .Z(n1257) );
  NANDN U1239 ( .A(n1260), .B(n1261), .Z(n1259) );
  NANDN U1240 ( .A(n1256), .B(n1262), .Z(n1261) );
  NANDN U1241 ( .A(n1263), .B(n1264), .Z(n1262) );
  NAND U1242 ( .A(n1265), .B(n1251), .Z(n1264) );
  XOR U1243 ( .A(n1266), .B(n1267), .Z(SUM[143]) );
  OR U1244 ( .A(n1237), .B(n1236), .Z(n1267) );
  AND U1245 ( .A(B[143]), .B(A[143]), .Z(n1236) );
  NOR U1246 ( .A(B[143]), .B(A[143]), .Z(n1237) );
  ANDN U1247 ( .B(n1268), .A(n1239), .Z(n1266) );
  NANDN U1248 ( .A(n1241), .B(n1269), .Z(n1268) );
  XNOR U1249 ( .A(n1269), .B(n1270), .Z(SUM[142]) );
  OR U1250 ( .A(n1241), .B(n1239), .Z(n1270) );
  AND U1251 ( .A(B[142]), .B(A[142]), .Z(n1239) );
  NOR U1252 ( .A(B[142]), .B(A[142]), .Z(n1241) );
  NANDN U1253 ( .A(n1243), .B(n1271), .Z(n1269) );
  NANDN U1254 ( .A(n1245), .B(n1272), .Z(n1271) );
  XNOR U1255 ( .A(n1272), .B(n1273), .Z(SUM[141]) );
  OR U1256 ( .A(n1245), .B(n1243), .Z(n1273) );
  AND U1257 ( .A(B[141]), .B(A[141]), .Z(n1243) );
  NOR U1258 ( .A(B[141]), .B(A[141]), .Z(n1245) );
  NANDN U1259 ( .A(n1258), .B(n1274), .Z(n1272) );
  NAND U1260 ( .A(n1275), .B(n1253), .Z(n1274) );
  XNOR U1261 ( .A(n1275), .B(n1276), .Z(SUM[140]) );
  NANDN U1262 ( .A(n1258), .B(n1253), .Z(n1276) );
  OR U1263 ( .A(A[140]), .B(B[140]), .Z(n1253) );
  AND U1264 ( .A(B[140]), .B(A[140]), .Z(n1258) );
  NANDN U1265 ( .A(n1260), .B(n1277), .Z(n1275) );
  NANDN U1266 ( .A(n1256), .B(n1278), .Z(n1277) );
  NAND U1267 ( .A(n1279), .B(n1280), .Z(n1256) );
  AND U1268 ( .A(n1281), .B(n1282), .Z(n1280) );
  AND U1269 ( .A(n1283), .B(n1284), .Z(n1279) );
  NANDN U1270 ( .A(n1285), .B(n1286), .Z(n1260) );
  NAND U1271 ( .A(n1287), .B(n1284), .Z(n1286) );
  NANDN U1272 ( .A(n1288), .B(n1289), .Z(n1287) );
  NAND U1273 ( .A(n1290), .B(n1283), .Z(n1289) );
  NANDN U1274 ( .A(n1291), .B(n1292), .Z(n1290) );
  NAND U1275 ( .A(n1282), .B(n1293), .Z(n1292) );
  XOR U1276 ( .A(n1294), .B(n1295), .Z(SUM[139]) );
  NANDN U1277 ( .A(n1285), .B(n1284), .Z(n1295) );
  OR U1278 ( .A(B[139]), .B(A[139]), .Z(n1284) );
  AND U1279 ( .A(B[139]), .B(A[139]), .Z(n1285) );
  ANDN U1280 ( .B(n1296), .A(n1288), .Z(n1294) );
  NAND U1281 ( .A(n1297), .B(n1283), .Z(n1296) );
  XNOR U1282 ( .A(n1297), .B(n1298), .Z(SUM[138]) );
  NANDN U1283 ( .A(n1288), .B(n1283), .Z(n1298) );
  OR U1284 ( .A(B[138]), .B(A[138]), .Z(n1283) );
  AND U1285 ( .A(B[138]), .B(A[138]), .Z(n1288) );
  NANDN U1286 ( .A(n1291), .B(n1299), .Z(n1297) );
  NAND U1287 ( .A(n1300), .B(n1282), .Z(n1299) );
  XNOR U1288 ( .A(n1300), .B(n1301), .Z(SUM[137]) );
  NANDN U1289 ( .A(n1291), .B(n1282), .Z(n1301) );
  OR U1290 ( .A(B[137]), .B(A[137]), .Z(n1282) );
  AND U1291 ( .A(B[137]), .B(A[137]), .Z(n1291) );
  NANDN U1292 ( .A(n1293), .B(n1302), .Z(n1300) );
  NAND U1293 ( .A(n1278), .B(n1281), .Z(n1302) );
  XNOR U1294 ( .A(n1278), .B(n1303), .Z(SUM[136]) );
  NANDN U1295 ( .A(n1293), .B(n1281), .Z(n1303) );
  OR U1296 ( .A(B[136]), .B(A[136]), .Z(n1281) );
  AND U1297 ( .A(B[136]), .B(A[136]), .Z(n1293) );
  NANDN U1298 ( .A(n1263), .B(n1304), .Z(n1278) );
  NANDN U1299 ( .A(n1305), .B(n1251), .Z(n1304) );
  AND U1300 ( .A(n1306), .B(n1307), .Z(n1251) );
  AND U1301 ( .A(n1308), .B(n1309), .Z(n1307) );
  AND U1302 ( .A(n1310), .B(n1311), .Z(n1306) );
  NANDN U1303 ( .A(n1312), .B(n1313), .Z(n1263) );
  NAND U1304 ( .A(n1314), .B(n1311), .Z(n1313) );
  NANDN U1305 ( .A(n1315), .B(n1316), .Z(n1314) );
  NAND U1306 ( .A(n1317), .B(n1310), .Z(n1316) );
  NANDN U1307 ( .A(n1318), .B(n1319), .Z(n1317) );
  NAND U1308 ( .A(n1309), .B(n1320), .Z(n1319) );
  XOR U1309 ( .A(n1321), .B(n1322), .Z(SUM[135]) );
  NANDN U1310 ( .A(n1312), .B(n1311), .Z(n1322) );
  OR U1311 ( .A(B[135]), .B(A[135]), .Z(n1311) );
  AND U1312 ( .A(B[135]), .B(A[135]), .Z(n1312) );
  ANDN U1313 ( .B(n1323), .A(n1315), .Z(n1321) );
  NAND U1314 ( .A(n1324), .B(n1310), .Z(n1323) );
  XNOR U1315 ( .A(n1324), .B(n1325), .Z(SUM[134]) );
  NANDN U1316 ( .A(n1315), .B(n1310), .Z(n1325) );
  OR U1317 ( .A(B[134]), .B(A[134]), .Z(n1310) );
  AND U1318 ( .A(B[134]), .B(A[134]), .Z(n1315) );
  NANDN U1319 ( .A(n1318), .B(n1326), .Z(n1324) );
  NAND U1320 ( .A(n1327), .B(n1309), .Z(n1326) );
  XNOR U1321 ( .A(n1327), .B(n1328), .Z(SUM[133]) );
  NANDN U1322 ( .A(n1318), .B(n1309), .Z(n1328) );
  OR U1323 ( .A(B[133]), .B(A[133]), .Z(n1309) );
  AND U1324 ( .A(B[133]), .B(A[133]), .Z(n1318) );
  NANDN U1325 ( .A(n1320), .B(n1329), .Z(n1327) );
  NANDN U1326 ( .A(n1305), .B(n1308), .Z(n1329) );
  XOR U1327 ( .A(n1305), .B(n1330), .Z(SUM[132]) );
  NANDN U1328 ( .A(n1320), .B(n1308), .Z(n1330) );
  OR U1329 ( .A(B[132]), .B(A[132]), .Z(n1308) );
  AND U1330 ( .A(B[132]), .B(A[132]), .Z(n1320) );
  ANDN U1331 ( .B(n1331), .A(n1265), .Z(n1305) );
  NANDN U1332 ( .A(n1332), .B(n1333), .Z(n1265) );
  NAND U1333 ( .A(n1334), .B(n1335), .Z(n1333) );
  NANDN U1334 ( .A(n1336), .B(n1337), .Z(n1334) );
  NANDN U1335 ( .A(n1338), .B(n1339), .Z(n1337) );
  NANDN U1336 ( .A(n1340), .B(n1341), .Z(n1339) );
  NAND U1337 ( .A(n1342), .B(n1343), .Z(n1341) );
  OR U1338 ( .A(n1255), .B(n1254), .Z(n1331) );
  NAND U1339 ( .A(n1344), .B(n1345), .Z(n1255) );
  AND U1340 ( .A(n1346), .B(n1342), .Z(n1345) );
  ANDN U1341 ( .B(n1335), .A(n1338), .Z(n1344) );
  XOR U1342 ( .A(n1347), .B(n1348), .Z(SUM[131]) );
  NANDN U1343 ( .A(n1332), .B(n1335), .Z(n1348) );
  OR U1344 ( .A(B[131]), .B(A[131]), .Z(n1335) );
  AND U1345 ( .A(B[131]), .B(A[131]), .Z(n1332) );
  ANDN U1346 ( .B(n1349), .A(n1336), .Z(n1347) );
  NANDN U1347 ( .A(n1338), .B(n1350), .Z(n1349) );
  XNOR U1348 ( .A(n1350), .B(n1351), .Z(SUM[130]) );
  OR U1349 ( .A(n1338), .B(n1336), .Z(n1351) );
  AND U1350 ( .A(B[130]), .B(A[130]), .Z(n1336) );
  NOR U1351 ( .A(B[130]), .B(A[130]), .Z(n1338) );
  NANDN U1352 ( .A(n1340), .B(n1352), .Z(n1350) );
  NAND U1353 ( .A(n1353), .B(n1342), .Z(n1352) );
  XNOR U1354 ( .A(n1353), .B(n1354), .Z(SUM[129]) );
  NANDN U1355 ( .A(n1340), .B(n1342), .Z(n1354) );
  OR U1356 ( .A(B[129]), .B(A[129]), .Z(n1342) );
  AND U1357 ( .A(B[129]), .B(A[129]), .Z(n1340) );
  NANDN U1358 ( .A(n1343), .B(n1355), .Z(n1353) );
  NANDN U1359 ( .A(n1254), .B(n1346), .Z(n1355) );
  XOR U1360 ( .A(n1254), .B(n1356), .Z(SUM[128]) );
  NANDN U1361 ( .A(n1343), .B(n1346), .Z(n1356) );
  OR U1362 ( .A(B[128]), .B(A[128]), .Z(n1346) );
  AND U1363 ( .A(A[128]), .B(B[128]), .Z(n1343) );
  ANDN U1364 ( .B(n1357), .A(n1358), .Z(n1254) );
  NANDN U1365 ( .A(n1359), .B(n1360), .Z(n1357) );
  NANDN U1366 ( .A(n1361), .B(n1362), .Z(n1360) );
  NANDN U1367 ( .A(n1363), .B(n1364), .Z(n1362) );
  NANDN U1368 ( .A(n1365), .B(n1366), .Z(n1364) );
  NANDN U1369 ( .A(n1367), .B(n1368), .Z(n1366) );
  NAND U1370 ( .A(n1369), .B(n1370), .Z(n1368) );
  NAND U1371 ( .A(n1371), .B(n1372), .Z(n1370) );
  AND U1372 ( .A(n1373), .B(n1374), .Z(n1372) );
  ANDN U1373 ( .B(n1375), .A(n1376), .Z(n1374) );
  NOR U1374 ( .A(n1377), .B(n1378), .Z(n1371) );
  ANDN U1375 ( .B(n1379), .A(n1380), .Z(n1369) );
  NAND U1376 ( .A(n1381), .B(n1375), .Z(n1379) );
  NANDN U1377 ( .A(n1382), .B(n1383), .Z(n1381) );
  NANDN U1378 ( .A(n1378), .B(n1384), .Z(n1383) );
  NANDN U1379 ( .A(n1385), .B(n1386), .Z(n1384) );
  NAND U1380 ( .A(n1387), .B(n1373), .Z(n1386) );
  XOR U1381 ( .A(n1388), .B(n1389), .Z(SUM[127]) );
  OR U1382 ( .A(n1359), .B(n1358), .Z(n1389) );
  AND U1383 ( .A(B[127]), .B(A[127]), .Z(n1358) );
  NOR U1384 ( .A(B[127]), .B(A[127]), .Z(n1359) );
  ANDN U1385 ( .B(n1390), .A(n1361), .Z(n1388) );
  NANDN U1386 ( .A(n1363), .B(n1391), .Z(n1390) );
  XNOR U1387 ( .A(n1391), .B(n1392), .Z(SUM[126]) );
  OR U1388 ( .A(n1363), .B(n1361), .Z(n1392) );
  AND U1389 ( .A(B[126]), .B(A[126]), .Z(n1361) );
  NOR U1390 ( .A(B[126]), .B(A[126]), .Z(n1363) );
  NANDN U1391 ( .A(n1365), .B(n1393), .Z(n1391) );
  NANDN U1392 ( .A(n1367), .B(n1394), .Z(n1393) );
  XNOR U1393 ( .A(n1394), .B(n1395), .Z(SUM[125]) );
  OR U1394 ( .A(n1367), .B(n1365), .Z(n1395) );
  AND U1395 ( .A(B[125]), .B(A[125]), .Z(n1365) );
  NOR U1396 ( .A(B[125]), .B(A[125]), .Z(n1367) );
  NANDN U1397 ( .A(n1380), .B(n1396), .Z(n1394) );
  NAND U1398 ( .A(n1397), .B(n1375), .Z(n1396) );
  XNOR U1399 ( .A(n1397), .B(n1398), .Z(SUM[124]) );
  NANDN U1400 ( .A(n1380), .B(n1375), .Z(n1398) );
  OR U1401 ( .A(A[124]), .B(B[124]), .Z(n1375) );
  AND U1402 ( .A(B[124]), .B(A[124]), .Z(n1380) );
  NANDN U1403 ( .A(n1382), .B(n1399), .Z(n1397) );
  NANDN U1404 ( .A(n1378), .B(n1400), .Z(n1399) );
  NAND U1405 ( .A(n1401), .B(n1402), .Z(n1378) );
  AND U1406 ( .A(n1403), .B(n1404), .Z(n1402) );
  AND U1407 ( .A(n1405), .B(n1406), .Z(n1401) );
  NANDN U1408 ( .A(n1407), .B(n1408), .Z(n1382) );
  NAND U1409 ( .A(n1409), .B(n1406), .Z(n1408) );
  NANDN U1410 ( .A(n1410), .B(n1411), .Z(n1409) );
  NAND U1411 ( .A(n1412), .B(n1405), .Z(n1411) );
  NANDN U1412 ( .A(n1413), .B(n1414), .Z(n1412) );
  NAND U1413 ( .A(n1404), .B(n1415), .Z(n1414) );
  XOR U1414 ( .A(n1416), .B(n1417), .Z(SUM[123]) );
  NANDN U1415 ( .A(n1407), .B(n1406), .Z(n1417) );
  OR U1416 ( .A(B[123]), .B(A[123]), .Z(n1406) );
  AND U1417 ( .A(B[123]), .B(A[123]), .Z(n1407) );
  ANDN U1418 ( .B(n1418), .A(n1410), .Z(n1416) );
  NAND U1419 ( .A(n1419), .B(n1405), .Z(n1418) );
  XNOR U1420 ( .A(n1419), .B(n1420), .Z(SUM[122]) );
  NANDN U1421 ( .A(n1410), .B(n1405), .Z(n1420) );
  OR U1422 ( .A(B[122]), .B(A[122]), .Z(n1405) );
  AND U1423 ( .A(B[122]), .B(A[122]), .Z(n1410) );
  NANDN U1424 ( .A(n1413), .B(n1421), .Z(n1419) );
  NAND U1425 ( .A(n1422), .B(n1404), .Z(n1421) );
  XNOR U1426 ( .A(n1422), .B(n1423), .Z(SUM[121]) );
  NANDN U1427 ( .A(n1413), .B(n1404), .Z(n1423) );
  OR U1428 ( .A(B[121]), .B(A[121]), .Z(n1404) );
  AND U1429 ( .A(B[121]), .B(A[121]), .Z(n1413) );
  NANDN U1430 ( .A(n1415), .B(n1424), .Z(n1422) );
  NAND U1431 ( .A(n1400), .B(n1403), .Z(n1424) );
  XNOR U1432 ( .A(n1400), .B(n1425), .Z(SUM[120]) );
  NANDN U1433 ( .A(n1415), .B(n1403), .Z(n1425) );
  OR U1434 ( .A(B[120]), .B(A[120]), .Z(n1403) );
  AND U1435 ( .A(B[120]), .B(A[120]), .Z(n1415) );
  NANDN U1436 ( .A(n1385), .B(n1426), .Z(n1400) );
  NANDN U1437 ( .A(n1427), .B(n1373), .Z(n1426) );
  AND U1438 ( .A(n1428), .B(n1429), .Z(n1373) );
  AND U1439 ( .A(n1430), .B(n1431), .Z(n1429) );
  AND U1440 ( .A(n1432), .B(n1433), .Z(n1428) );
  NANDN U1441 ( .A(n1434), .B(n1435), .Z(n1385) );
  NAND U1442 ( .A(n1436), .B(n1433), .Z(n1435) );
  NANDN U1443 ( .A(n1437), .B(n1438), .Z(n1436) );
  NAND U1444 ( .A(n1439), .B(n1432), .Z(n1438) );
  NANDN U1445 ( .A(n1440), .B(n1441), .Z(n1439) );
  NAND U1446 ( .A(n1431), .B(n1442), .Z(n1441) );
  XOR U1447 ( .A(n1443), .B(n1444), .Z(SUM[119]) );
  NANDN U1448 ( .A(n1434), .B(n1433), .Z(n1444) );
  OR U1449 ( .A(B[119]), .B(A[119]), .Z(n1433) );
  AND U1450 ( .A(B[119]), .B(A[119]), .Z(n1434) );
  ANDN U1451 ( .B(n1445), .A(n1437), .Z(n1443) );
  NAND U1452 ( .A(n1446), .B(n1432), .Z(n1445) );
  XNOR U1453 ( .A(n1446), .B(n1447), .Z(SUM[118]) );
  NANDN U1454 ( .A(n1437), .B(n1432), .Z(n1447) );
  OR U1455 ( .A(B[118]), .B(A[118]), .Z(n1432) );
  AND U1456 ( .A(B[118]), .B(A[118]), .Z(n1437) );
  NANDN U1457 ( .A(n1440), .B(n1448), .Z(n1446) );
  NAND U1458 ( .A(n1449), .B(n1431), .Z(n1448) );
  XNOR U1459 ( .A(n1449), .B(n1450), .Z(SUM[117]) );
  NANDN U1460 ( .A(n1440), .B(n1431), .Z(n1450) );
  OR U1461 ( .A(B[117]), .B(A[117]), .Z(n1431) );
  AND U1462 ( .A(B[117]), .B(A[117]), .Z(n1440) );
  NANDN U1463 ( .A(n1442), .B(n1451), .Z(n1449) );
  NANDN U1464 ( .A(n1427), .B(n1430), .Z(n1451) );
  XOR U1465 ( .A(n1427), .B(n1452), .Z(SUM[116]) );
  NANDN U1466 ( .A(n1442), .B(n1430), .Z(n1452) );
  OR U1467 ( .A(B[116]), .B(A[116]), .Z(n1430) );
  AND U1468 ( .A(B[116]), .B(A[116]), .Z(n1442) );
  ANDN U1469 ( .B(n1453), .A(n1387), .Z(n1427) );
  NANDN U1470 ( .A(n1454), .B(n1455), .Z(n1387) );
  NAND U1471 ( .A(n1456), .B(n1457), .Z(n1455) );
  NANDN U1472 ( .A(n1458), .B(n1459), .Z(n1456) );
  NANDN U1473 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1474 ( .A(n1462), .B(n1463), .Z(n1461) );
  NAND U1475 ( .A(n1464), .B(n1465), .Z(n1463) );
  OR U1476 ( .A(n1377), .B(n1376), .Z(n1453) );
  NAND U1477 ( .A(n1466), .B(n1467), .Z(n1377) );
  AND U1478 ( .A(n1468), .B(n1464), .Z(n1467) );
  ANDN U1479 ( .B(n1457), .A(n1460), .Z(n1466) );
  XOR U1480 ( .A(n1469), .B(n1470), .Z(SUM[115]) );
  NANDN U1481 ( .A(n1454), .B(n1457), .Z(n1470) );
  OR U1482 ( .A(B[115]), .B(A[115]), .Z(n1457) );
  AND U1483 ( .A(B[115]), .B(A[115]), .Z(n1454) );
  ANDN U1484 ( .B(n1471), .A(n1458), .Z(n1469) );
  NANDN U1485 ( .A(n1460), .B(n1472), .Z(n1471) );
  XNOR U1486 ( .A(n1472), .B(n1473), .Z(SUM[114]) );
  OR U1487 ( .A(n1460), .B(n1458), .Z(n1473) );
  AND U1488 ( .A(B[114]), .B(A[114]), .Z(n1458) );
  NOR U1489 ( .A(B[114]), .B(A[114]), .Z(n1460) );
  NANDN U1490 ( .A(n1462), .B(n1474), .Z(n1472) );
  NAND U1491 ( .A(n1475), .B(n1464), .Z(n1474) );
  XNOR U1492 ( .A(n1475), .B(n1476), .Z(SUM[113]) );
  NANDN U1493 ( .A(n1462), .B(n1464), .Z(n1476) );
  OR U1494 ( .A(B[113]), .B(A[113]), .Z(n1464) );
  AND U1495 ( .A(B[113]), .B(A[113]), .Z(n1462) );
  NANDN U1496 ( .A(n1465), .B(n1477), .Z(n1475) );
  NANDN U1497 ( .A(n1376), .B(n1468), .Z(n1477) );
  XOR U1498 ( .A(n1376), .B(n1478), .Z(SUM[112]) );
  NANDN U1499 ( .A(n1465), .B(n1468), .Z(n1478) );
  OR U1500 ( .A(B[112]), .B(A[112]), .Z(n1468) );
  AND U1501 ( .A(A[112]), .B(B[112]), .Z(n1465) );
  ANDN U1502 ( .B(n1479), .A(n1480), .Z(n1376) );
  NANDN U1503 ( .A(n1481), .B(n1482), .Z(n1479) );
  NANDN U1504 ( .A(n1483), .B(n1484), .Z(n1482) );
  NANDN U1505 ( .A(n1485), .B(n1486), .Z(n1484) );
  NANDN U1506 ( .A(n1487), .B(n1488), .Z(n1486) );
  NANDN U1507 ( .A(n1489), .B(n1490), .Z(n1488) );
  NAND U1508 ( .A(n1491), .B(n1492), .Z(n1490) );
  NAND U1509 ( .A(n1493), .B(n1494), .Z(n1492) );
  AND U1510 ( .A(n1495), .B(n1496), .Z(n1494) );
  ANDN U1511 ( .B(n1497), .A(n17), .Z(n1496) );
  NOR U1512 ( .A(n1498), .B(n1499), .Z(n1493) );
  ANDN U1513 ( .B(n1500), .A(n1501), .Z(n1491) );
  NAND U1514 ( .A(n1502), .B(n1497), .Z(n1500) );
  NANDN U1515 ( .A(n1503), .B(n1504), .Z(n1502) );
  NANDN U1516 ( .A(n1499), .B(n1505), .Z(n1504) );
  NANDN U1517 ( .A(n1506), .B(n1507), .Z(n1505) );
  NAND U1518 ( .A(n1508), .B(n1495), .Z(n1507) );
  XOR U1519 ( .A(n1509), .B(n1510), .Z(SUM[111]) );
  OR U1520 ( .A(n1481), .B(n1480), .Z(n1510) );
  AND U1521 ( .A(B[111]), .B(A[111]), .Z(n1480) );
  NOR U1522 ( .A(B[111]), .B(A[111]), .Z(n1481) );
  ANDN U1523 ( .B(n1511), .A(n1483), .Z(n1509) );
  NANDN U1524 ( .A(n1485), .B(n1512), .Z(n1511) );
  XNOR U1525 ( .A(n1512), .B(n1513), .Z(SUM[110]) );
  OR U1526 ( .A(n1485), .B(n1483), .Z(n1513) );
  AND U1527 ( .A(B[110]), .B(A[110]), .Z(n1483) );
  NOR U1528 ( .A(B[110]), .B(A[110]), .Z(n1485) );
  NANDN U1529 ( .A(n1487), .B(n1514), .Z(n1512) );
  NANDN U1530 ( .A(n1489), .B(n1515), .Z(n1514) );
  XNOR U1531 ( .A(n1515), .B(n1516), .Z(SUM[109]) );
  OR U1532 ( .A(n1489), .B(n1487), .Z(n1516) );
  AND U1533 ( .A(B[109]), .B(A[109]), .Z(n1487) );
  NOR U1534 ( .A(B[109]), .B(A[109]), .Z(n1489) );
  NANDN U1535 ( .A(n1501), .B(n1517), .Z(n1515) );
  NAND U1536 ( .A(n1518), .B(n1497), .Z(n1517) );
  XNOR U1537 ( .A(n1518), .B(n1519), .Z(SUM[108]) );
  NANDN U1538 ( .A(n1501), .B(n1497), .Z(n1519) );
  OR U1539 ( .A(A[108]), .B(B[108]), .Z(n1497) );
  AND U1540 ( .A(B[108]), .B(A[108]), .Z(n1501) );
  NANDN U1541 ( .A(n1503), .B(n1520), .Z(n1518) );
  NANDN U1542 ( .A(n1499), .B(n1521), .Z(n1520) );
  NAND U1543 ( .A(n1522), .B(n1523), .Z(n1499) );
  AND U1544 ( .A(n1524), .B(n1525), .Z(n1523) );
  AND U1545 ( .A(n1526), .B(n1527), .Z(n1522) );
  NANDN U1546 ( .A(n1528), .B(n1529), .Z(n1503) );
  NAND U1547 ( .A(n1530), .B(n1527), .Z(n1529) );
  NANDN U1548 ( .A(n1531), .B(n1532), .Z(n1530) );
  NAND U1549 ( .A(n1533), .B(n1526), .Z(n1532) );
  NANDN U1550 ( .A(n1534), .B(n1535), .Z(n1533) );
  NAND U1551 ( .A(n1525), .B(n1536), .Z(n1535) );
  XOR U1552 ( .A(n1537), .B(n1538), .Z(SUM[107]) );
  NANDN U1553 ( .A(n1528), .B(n1527), .Z(n1538) );
  OR U1554 ( .A(B[107]), .B(A[107]), .Z(n1527) );
  AND U1555 ( .A(B[107]), .B(A[107]), .Z(n1528) );
  ANDN U1556 ( .B(n1539), .A(n1531), .Z(n1537) );
  NAND U1557 ( .A(n1540), .B(n1526), .Z(n1539) );
  XNOR U1558 ( .A(n1540), .B(n1541), .Z(SUM[106]) );
  NANDN U1559 ( .A(n1531), .B(n1526), .Z(n1541) );
  OR U1560 ( .A(B[106]), .B(A[106]), .Z(n1526) );
  AND U1561 ( .A(B[106]), .B(A[106]), .Z(n1531) );
  NANDN U1562 ( .A(n1534), .B(n1542), .Z(n1540) );
  NAND U1563 ( .A(n1543), .B(n1525), .Z(n1542) );
  XNOR U1564 ( .A(n1543), .B(n1544), .Z(SUM[105]) );
  NANDN U1565 ( .A(n1534), .B(n1525), .Z(n1544) );
  OR U1566 ( .A(B[105]), .B(A[105]), .Z(n1525) );
  AND U1567 ( .A(B[105]), .B(A[105]), .Z(n1534) );
  NANDN U1568 ( .A(n1536), .B(n1545), .Z(n1543) );
  NAND U1569 ( .A(n1521), .B(n1524), .Z(n1545) );
  XNOR U1570 ( .A(n1521), .B(n1546), .Z(SUM[104]) );
  NANDN U1571 ( .A(n1536), .B(n1524), .Z(n1546) );
  OR U1572 ( .A(B[104]), .B(A[104]), .Z(n1524) );
  AND U1573 ( .A(B[104]), .B(A[104]), .Z(n1536) );
  NANDN U1574 ( .A(n1506), .B(n1547), .Z(n1521) );
  NANDN U1575 ( .A(n1548), .B(n1495), .Z(n1547) );
  AND U1576 ( .A(n1549), .B(n1550), .Z(n1495) );
  AND U1577 ( .A(n1551), .B(n1552), .Z(n1550) );
  AND U1578 ( .A(n1553), .B(n1554), .Z(n1549) );
  NANDN U1579 ( .A(n1555), .B(n1556), .Z(n1506) );
  NAND U1580 ( .A(n1557), .B(n1554), .Z(n1556) );
  NANDN U1581 ( .A(n1558), .B(n1559), .Z(n1557) );
  NAND U1582 ( .A(n1560), .B(n1553), .Z(n1559) );
  NANDN U1583 ( .A(n1561), .B(n1562), .Z(n1560) );
  NAND U1584 ( .A(n1552), .B(n1563), .Z(n1562) );
  XOR U1585 ( .A(n1564), .B(n1565), .Z(SUM[103]) );
  NANDN U1586 ( .A(n1555), .B(n1554), .Z(n1565) );
  OR U1587 ( .A(B[103]), .B(A[103]), .Z(n1554) );
  AND U1588 ( .A(B[103]), .B(A[103]), .Z(n1555) );
  ANDN U1589 ( .B(n1566), .A(n1558), .Z(n1564) );
  NAND U1590 ( .A(n1567), .B(n1553), .Z(n1566) );
  XNOR U1591 ( .A(n1567), .B(n1568), .Z(SUM[102]) );
  NANDN U1592 ( .A(n1558), .B(n1553), .Z(n1568) );
  OR U1593 ( .A(B[102]), .B(A[102]), .Z(n1553) );
  AND U1594 ( .A(B[102]), .B(A[102]), .Z(n1558) );
  NANDN U1595 ( .A(n1561), .B(n1569), .Z(n1567) );
  NAND U1596 ( .A(n1570), .B(n1552), .Z(n1569) );
  XNOR U1597 ( .A(n1570), .B(n1571), .Z(SUM[101]) );
  NANDN U1598 ( .A(n1561), .B(n1552), .Z(n1571) );
  OR U1599 ( .A(B[101]), .B(A[101]), .Z(n1552) );
  AND U1600 ( .A(B[101]), .B(A[101]), .Z(n1561) );
  NANDN U1601 ( .A(n1563), .B(n1572), .Z(n1570) );
  NANDN U1602 ( .A(n1548), .B(n1551), .Z(n1572) );
  XOR U1603 ( .A(n1548), .B(n1573), .Z(SUM[100]) );
  NANDN U1604 ( .A(n1563), .B(n1551), .Z(n1573) );
  OR U1605 ( .A(B[100]), .B(A[100]), .Z(n1551) );
  AND U1606 ( .A(B[100]), .B(A[100]), .Z(n1563) );
  ANDN U1607 ( .B(n1574), .A(n1508), .Z(n1548) );
  NANDN U1608 ( .A(n3), .B(n1575), .Z(n1508) );
  NAND U1609 ( .A(n1576), .B(n4), .Z(n1575) );
  NANDN U1610 ( .A(n6), .B(n1577), .Z(n1576) );
  NAND U1611 ( .A(n1578), .B(n8), .Z(n1577) );
  NANDN U1612 ( .A(n10), .B(n1579), .Z(n1578) );
  NANDN U1613 ( .A(n15), .B(n13), .Z(n1579) );
  NAND U1614 ( .A(B[96]), .B(A[96]), .Z(n15) );
  AND U1615 ( .A(B[97]), .B(A[97]), .Z(n10) );
  AND U1616 ( .A(A[98]), .B(B[98]), .Z(n6) );
  AND U1617 ( .A(B[99]), .B(A[99]), .Z(n3) );
  OR U1618 ( .A(n1498), .B(n17), .Z(n1574) );
  ANDN U1619 ( .B(n1580), .A(n23), .Z(n17) );
  AND U1620 ( .A(B[95]), .B(A[95]), .Z(n23) );
  NANDN U1621 ( .A(n22), .B(n1581), .Z(n1580) );
  NANDN U1622 ( .A(n25), .B(n1582), .Z(n1581) );
  NANDN U1623 ( .A(n26), .B(n1583), .Z(n1582) );
  NANDN U1624 ( .A(n29), .B(n1584), .Z(n1583) );
  NANDN U1625 ( .A(n31), .B(n1585), .Z(n1584) );
  NAND U1626 ( .A(n1586), .B(n1587), .Z(n1585) );
  NAND U1627 ( .A(n1588), .B(n1589), .Z(n1587) );
  AND U1628 ( .A(n64), .B(n1590), .Z(n1589) );
  ANDN U1629 ( .B(n37), .A(n86), .Z(n1590) );
  ANDN U1630 ( .B(n1591), .A(n108), .Z(n86) );
  AND U1631 ( .A(B[79]), .B(A[79]), .Z(n108) );
  NANDN U1632 ( .A(n107), .B(n1592), .Z(n1591) );
  NANDN U1633 ( .A(n110), .B(n1593), .Z(n1592) );
  NANDN U1634 ( .A(n111), .B(n1594), .Z(n1593) );
  NANDN U1635 ( .A(n114), .B(n1595), .Z(n1594) );
  NANDN U1636 ( .A(n116), .B(n1596), .Z(n1595) );
  NAND U1637 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1638 ( .A(n1599), .B(n1600), .Z(n1598) );
  AND U1639 ( .A(n149), .B(n1601), .Z(n1600) );
  ANDN U1640 ( .B(n122), .A(n171), .Z(n1601) );
  ANDN U1641 ( .B(n1602), .A(n193), .Z(n171) );
  AND U1642 ( .A(B[63]), .B(A[63]), .Z(n193) );
  NANDN U1643 ( .A(n192), .B(n1603), .Z(n1602) );
  NANDN U1644 ( .A(n195), .B(n1604), .Z(n1603) );
  NANDN U1645 ( .A(n196), .B(n1605), .Z(n1604) );
  NANDN U1646 ( .A(n199), .B(n1606), .Z(n1605) );
  NANDN U1647 ( .A(n201), .B(n1607), .Z(n1606) );
  NANDN U1648 ( .A(n204), .B(n1608), .Z(n1607) );
  NANDN U1649 ( .A(n206), .B(n1609), .Z(n1608) );
  NANDN U1650 ( .A(n209), .B(n1610), .Z(n1609) );
  NANDN U1651 ( .A(n211), .B(n1611), .Z(n1610) );
  NANDN U1652 ( .A(n231), .B(n1612), .Z(n1611) );
  AND U1653 ( .A(n1613), .B(n1614), .Z(n1612) );
  NANDN U1654 ( .A(n233), .B(n253), .Z(n1614) );
  NANDN U1655 ( .A(n257), .B(n1615), .Z(n253) );
  NAND U1656 ( .A(n1616), .B(n258), .Z(n1615) );
  NANDN U1657 ( .A(n260), .B(n1617), .Z(n1616) );
  NAND U1658 ( .A(n1618), .B(n262), .Z(n1617) );
  NANDN U1659 ( .A(n264), .B(n1619), .Z(n1618) );
  NAND U1660 ( .A(n267), .B(n269), .Z(n1619) );
  AND U1661 ( .A(A[48]), .B(B[48]), .Z(n269) );
  AND U1662 ( .A(A[49]), .B(B[49]), .Z(n264) );
  AND U1663 ( .A(A[50]), .B(B[50]), .Z(n260) );
  AND U1664 ( .A(B[51]), .B(A[51]), .Z(n257) );
  NANDN U1665 ( .A(n233), .B(n254), .Z(n1613) );
  AND U1666 ( .A(n1620), .B(n1621), .Z(n254) );
  AND U1667 ( .A(n262), .B(n1622), .Z(n1621) );
  AND U1668 ( .A(n272), .B(n267), .Z(n1622) );
  OR U1669 ( .A(A[49]), .B(B[49]), .Z(n267) );
  OR U1670 ( .A(A[48]), .B(B[48]), .Z(n272) );
  OR U1671 ( .A(A[50]), .B(B[50]), .Z(n262) );
  ANDN U1672 ( .B(n258), .A(n271), .Z(n1620) );
  ANDN U1673 ( .B(n1623), .A(n277), .Z(n271) );
  AND U1674 ( .A(B[47]), .B(A[47]), .Z(n277) );
  NANDN U1675 ( .A(n276), .B(n1624), .Z(n1623) );
  NANDN U1676 ( .A(n279), .B(n1625), .Z(n1624) );
  NANDN U1677 ( .A(n280), .B(n1626), .Z(n1625) );
  NANDN U1678 ( .A(n283), .B(n1627), .Z(n1626) );
  NANDN U1679 ( .A(n285), .B(n1628), .Z(n1627) );
  NAND U1680 ( .A(n1629), .B(n1630), .Z(n1628) );
  NAND U1681 ( .A(n1631), .B(n1632), .Z(n1630) );
  AND U1682 ( .A(n318), .B(n1633), .Z(n1632) );
  ANDN U1683 ( .B(n291), .A(n340), .Z(n1633) );
  ANDN U1684 ( .B(n1634), .A(n362), .Z(n340) );
  AND U1685 ( .A(B[31]), .B(A[31]), .Z(n362) );
  NANDN U1686 ( .A(n361), .B(n1635), .Z(n1634) );
  NANDN U1687 ( .A(n364), .B(n1636), .Z(n1635) );
  NANDN U1688 ( .A(n365), .B(n1637), .Z(n1636) );
  NANDN U1689 ( .A(n368), .B(n1638), .Z(n1637) );
  NANDN U1690 ( .A(n370), .B(n1639), .Z(n1638) );
  NAND U1691 ( .A(n1640), .B(n1641), .Z(n1639) );
  NAND U1692 ( .A(n1642), .B(n1643), .Z(n1641) );
  ANDN U1693 ( .B(n1644), .A(n380), .Z(n1643) );
  AND U1694 ( .A(n376), .B(n424), .Z(n1644) );
  ANDN U1695 ( .B(n727), .A(n726), .Z(n1642) );
  NAND U1696 ( .A(n1645), .B(n1646), .Z(n726) );
  AND U1697 ( .A(n978), .B(n900), .Z(n1646) );
  OR U1698 ( .A(B[16]), .B(A[16]), .Z(n978) );
  ANDN U1699 ( .B(n816), .A(n819), .Z(n1645) );
  AND U1700 ( .A(A[15]), .B(B[15]), .Z(n727) );
  ANDN U1701 ( .B(n1647), .A(n373), .Z(n1640) );
  AND U1702 ( .A(B[28]), .B(A[28]), .Z(n373) );
  NAND U1703 ( .A(n1648), .B(n376), .Z(n1647) );
  OR U1704 ( .A(A[28]), .B(B[28]), .Z(n376) );
  NANDN U1705 ( .A(n378), .B(n1649), .Z(n1648) );
  NANDN U1706 ( .A(n380), .B(n1650), .Z(n1649) );
  NANDN U1707 ( .A(n421), .B(n1651), .Z(n1650) );
  NAND U1708 ( .A(n725), .B(n424), .Z(n1651) );
  AND U1709 ( .A(n1652), .B(n1653), .Z(n424) );
  AND U1710 ( .A(n661), .B(n572), .Z(n1653) );
  OR U1711 ( .A(B[20]), .B(A[20]), .Z(n661) );
  AND U1712 ( .A(n505), .B(n501), .Z(n1652) );
  NANDN U1713 ( .A(n815), .B(n1654), .Z(n725) );
  NAND U1714 ( .A(n1655), .B(n816), .Z(n1654) );
  OR U1715 ( .A(B[19]), .B(A[19]), .Z(n816) );
  NANDN U1716 ( .A(n818), .B(n1656), .Z(n1655) );
  NANDN U1717 ( .A(n819), .B(n1657), .Z(n1656) );
  NANDN U1718 ( .A(n897), .B(n1658), .Z(n1657) );
  NAND U1719 ( .A(n900), .B(n976), .Z(n1658) );
  AND U1720 ( .A(A[16]), .B(B[16]), .Z(n976) );
  OR U1721 ( .A(B[17]), .B(A[17]), .Z(n900) );
  AND U1722 ( .A(B[17]), .B(A[17]), .Z(n897) );
  NOR U1723 ( .A(B[18]), .B(A[18]), .Z(n819) );
  AND U1724 ( .A(B[18]), .B(A[18]), .Z(n818) );
  AND U1725 ( .A(B[19]), .B(A[19]), .Z(n815) );
  NANDN U1726 ( .A(n500), .B(n1659), .Z(n421) );
  NAND U1727 ( .A(n1660), .B(n501), .Z(n1659) );
  OR U1728 ( .A(B[23]), .B(A[23]), .Z(n501) );
  NANDN U1729 ( .A(n503), .B(n1661), .Z(n1660) );
  NAND U1730 ( .A(n1662), .B(n505), .Z(n1661) );
  OR U1731 ( .A(B[22]), .B(A[22]), .Z(n505) );
  NANDN U1732 ( .A(n569), .B(n1663), .Z(n1662) );
  NAND U1733 ( .A(n572), .B(n659), .Z(n1663) );
  AND U1734 ( .A(B[20]), .B(A[20]), .Z(n659) );
  OR U1735 ( .A(B[21]), .B(A[21]), .Z(n572) );
  AND U1736 ( .A(B[21]), .B(A[21]), .Z(n569) );
  AND U1737 ( .A(B[22]), .B(A[22]), .Z(n503) );
  AND U1738 ( .A(B[23]), .B(A[23]), .Z(n500) );
  NAND U1739 ( .A(n1664), .B(n1665), .Z(n380) );
  AND U1740 ( .A(n398), .B(n394), .Z(n1665) );
  OR U1741 ( .A(B[24]), .B(A[24]), .Z(n398) );
  AND U1742 ( .A(n389), .B(n385), .Z(n1664) );
  NANDN U1743 ( .A(n384), .B(n1666), .Z(n378) );
  NAND U1744 ( .A(n1667), .B(n385), .Z(n1666) );
  OR U1745 ( .A(B[27]), .B(A[27]), .Z(n385) );
  NANDN U1746 ( .A(n387), .B(n1668), .Z(n1667) );
  NAND U1747 ( .A(n1669), .B(n389), .Z(n1668) );
  OR U1748 ( .A(B[26]), .B(A[26]), .Z(n389) );
  NANDN U1749 ( .A(n391), .B(n1670), .Z(n1669) );
  NAND U1750 ( .A(n394), .B(n396), .Z(n1670) );
  AND U1751 ( .A(B[24]), .B(A[24]), .Z(n396) );
  OR U1752 ( .A(B[25]), .B(A[25]), .Z(n394) );
  AND U1753 ( .A(B[25]), .B(A[25]), .Z(n391) );
  AND U1754 ( .A(B[26]), .B(A[26]), .Z(n387) );
  AND U1755 ( .A(B[27]), .B(A[27]), .Z(n384) );
  NOR U1756 ( .A(B[29]), .B(A[29]), .Z(n370) );
  AND U1757 ( .A(B[29]), .B(A[29]), .Z(n368) );
  NOR U1758 ( .A(B[30]), .B(A[30]), .Z(n365) );
  AND U1759 ( .A(B[30]), .B(A[30]), .Z(n364) );
  NOR U1760 ( .A(B[31]), .B(A[31]), .Z(n361) );
  NOR U1761 ( .A(n339), .B(n295), .Z(n1631) );
  NAND U1762 ( .A(n1671), .B(n1672), .Z(n339) );
  AND U1763 ( .A(n357), .B(n353), .Z(n1672) );
  OR U1764 ( .A(B[32]), .B(A[32]), .Z(n357) );
  ANDN U1765 ( .B(n344), .A(n347), .Z(n1671) );
  ANDN U1766 ( .B(n1673), .A(n288), .Z(n1629) );
  AND U1767 ( .A(B[44]), .B(A[44]), .Z(n288) );
  NAND U1768 ( .A(n1674), .B(n291), .Z(n1673) );
  OR U1769 ( .A(A[44]), .B(B[44]), .Z(n291) );
  NANDN U1770 ( .A(n293), .B(n1675), .Z(n1674) );
  NANDN U1771 ( .A(n295), .B(n1676), .Z(n1675) );
  NANDN U1772 ( .A(n315), .B(n1677), .Z(n1676) );
  NAND U1773 ( .A(n338), .B(n318), .Z(n1677) );
  AND U1774 ( .A(n1678), .B(n1679), .Z(n318) );
  AND U1775 ( .A(n335), .B(n331), .Z(n1679) );
  OR U1776 ( .A(B[36]), .B(A[36]), .Z(n335) );
  AND U1777 ( .A(n326), .B(n322), .Z(n1678) );
  NANDN U1778 ( .A(n343), .B(n1680), .Z(n338) );
  NAND U1779 ( .A(n1681), .B(n344), .Z(n1680) );
  OR U1780 ( .A(B[35]), .B(A[35]), .Z(n344) );
  NANDN U1781 ( .A(n346), .B(n1682), .Z(n1681) );
  NANDN U1782 ( .A(n347), .B(n1683), .Z(n1682) );
  NANDN U1783 ( .A(n350), .B(n1684), .Z(n1683) );
  NAND U1784 ( .A(n353), .B(n355), .Z(n1684) );
  AND U1785 ( .A(A[32]), .B(B[32]), .Z(n355) );
  OR U1786 ( .A(B[33]), .B(A[33]), .Z(n353) );
  AND U1787 ( .A(B[33]), .B(A[33]), .Z(n350) );
  NOR U1788 ( .A(B[34]), .B(A[34]), .Z(n347) );
  AND U1789 ( .A(B[34]), .B(A[34]), .Z(n346) );
  AND U1790 ( .A(B[35]), .B(A[35]), .Z(n343) );
  NANDN U1791 ( .A(n321), .B(n1685), .Z(n315) );
  NAND U1792 ( .A(n1686), .B(n322), .Z(n1685) );
  OR U1793 ( .A(B[39]), .B(A[39]), .Z(n322) );
  NANDN U1794 ( .A(n324), .B(n1687), .Z(n1686) );
  NAND U1795 ( .A(n1688), .B(n326), .Z(n1687) );
  OR U1796 ( .A(B[38]), .B(A[38]), .Z(n326) );
  NANDN U1797 ( .A(n328), .B(n1689), .Z(n1688) );
  NAND U1798 ( .A(n331), .B(n333), .Z(n1689) );
  AND U1799 ( .A(B[36]), .B(A[36]), .Z(n333) );
  OR U1800 ( .A(B[37]), .B(A[37]), .Z(n331) );
  AND U1801 ( .A(B[37]), .B(A[37]), .Z(n328) );
  AND U1802 ( .A(B[38]), .B(A[38]), .Z(n324) );
  AND U1803 ( .A(B[39]), .B(A[39]), .Z(n321) );
  NAND U1804 ( .A(n1690), .B(n1691), .Z(n295) );
  AND U1805 ( .A(n313), .B(n309), .Z(n1691) );
  OR U1806 ( .A(B[40]), .B(A[40]), .Z(n313) );
  AND U1807 ( .A(n304), .B(n300), .Z(n1690) );
  NANDN U1808 ( .A(n299), .B(n1692), .Z(n293) );
  NAND U1809 ( .A(n1693), .B(n300), .Z(n1692) );
  OR U1810 ( .A(B[43]), .B(A[43]), .Z(n300) );
  NANDN U1811 ( .A(n302), .B(n1694), .Z(n1693) );
  NAND U1812 ( .A(n1695), .B(n304), .Z(n1694) );
  OR U1813 ( .A(B[42]), .B(A[42]), .Z(n304) );
  NANDN U1814 ( .A(n306), .B(n1696), .Z(n1695) );
  NAND U1815 ( .A(n309), .B(n311), .Z(n1696) );
  AND U1816 ( .A(B[40]), .B(A[40]), .Z(n311) );
  OR U1817 ( .A(B[41]), .B(A[41]), .Z(n309) );
  AND U1818 ( .A(B[41]), .B(A[41]), .Z(n306) );
  AND U1819 ( .A(B[42]), .B(A[42]), .Z(n302) );
  AND U1820 ( .A(B[43]), .B(A[43]), .Z(n299) );
  NOR U1821 ( .A(B[45]), .B(A[45]), .Z(n285) );
  AND U1822 ( .A(B[45]), .B(A[45]), .Z(n283) );
  NOR U1823 ( .A(B[46]), .B(A[46]), .Z(n280) );
  AND U1824 ( .A(B[46]), .B(A[46]), .Z(n279) );
  NOR U1825 ( .A(B[47]), .B(A[47]), .Z(n276) );
  OR U1826 ( .A(B[51]), .B(A[51]), .Z(n258) );
  NAND U1827 ( .A(n1697), .B(n1698), .Z(n233) );
  AND U1828 ( .A(n251), .B(n247), .Z(n1698) );
  OR U1829 ( .A(A[52]), .B(B[52]), .Z(n251) );
  AND U1830 ( .A(n242), .B(n238), .Z(n1697) );
  NANDN U1831 ( .A(n237), .B(n1699), .Z(n231) );
  NAND U1832 ( .A(n1700), .B(n238), .Z(n1699) );
  OR U1833 ( .A(B[55]), .B(A[55]), .Z(n238) );
  NANDN U1834 ( .A(n240), .B(n1701), .Z(n1700) );
  NAND U1835 ( .A(n1702), .B(n242), .Z(n1701) );
  OR U1836 ( .A(A[54]), .B(B[54]), .Z(n242) );
  NANDN U1837 ( .A(n244), .B(n1703), .Z(n1702) );
  NAND U1838 ( .A(n247), .B(n249), .Z(n1703) );
  AND U1839 ( .A(A[52]), .B(B[52]), .Z(n249) );
  OR U1840 ( .A(A[53]), .B(B[53]), .Z(n247) );
  AND U1841 ( .A(A[53]), .B(B[53]), .Z(n244) );
  AND U1842 ( .A(A[54]), .B(B[54]), .Z(n240) );
  AND U1843 ( .A(B[55]), .B(A[55]), .Z(n237) );
  NAND U1844 ( .A(n1704), .B(n1705), .Z(n211) );
  AND U1845 ( .A(n229), .B(n225), .Z(n1705) );
  OR U1846 ( .A(B[56]), .B(A[56]), .Z(n229) );
  AND U1847 ( .A(n220), .B(n216), .Z(n1704) );
  NANDN U1848 ( .A(n215), .B(n1706), .Z(n209) );
  NAND U1849 ( .A(n1707), .B(n216), .Z(n1706) );
  OR U1850 ( .A(B[59]), .B(A[59]), .Z(n216) );
  NANDN U1851 ( .A(n218), .B(n1708), .Z(n1707) );
  NAND U1852 ( .A(n1709), .B(n220), .Z(n1708) );
  OR U1853 ( .A(B[58]), .B(A[58]), .Z(n220) );
  NANDN U1854 ( .A(n222), .B(n1710), .Z(n1709) );
  NAND U1855 ( .A(n225), .B(n227), .Z(n1710) );
  AND U1856 ( .A(B[56]), .B(A[56]), .Z(n227) );
  OR U1857 ( .A(B[57]), .B(A[57]), .Z(n225) );
  AND U1858 ( .A(B[57]), .B(A[57]), .Z(n222) );
  AND U1859 ( .A(B[58]), .B(A[58]), .Z(n218) );
  AND U1860 ( .A(B[59]), .B(A[59]), .Z(n215) );
  NOR U1861 ( .A(B[60]), .B(A[60]), .Z(n206) );
  AND U1862 ( .A(B[60]), .B(A[60]), .Z(n204) );
  NOR U1863 ( .A(B[61]), .B(A[61]), .Z(n201) );
  AND U1864 ( .A(B[61]), .B(A[61]), .Z(n199) );
  NOR U1865 ( .A(B[62]), .B(A[62]), .Z(n196) );
  AND U1866 ( .A(B[62]), .B(A[62]), .Z(n195) );
  NOR U1867 ( .A(B[63]), .B(A[63]), .Z(n192) );
  NOR U1868 ( .A(n170), .B(n126), .Z(n1599) );
  NAND U1869 ( .A(n1711), .B(n1712), .Z(n170) );
  AND U1870 ( .A(n188), .B(n184), .Z(n1712) );
  OR U1871 ( .A(B[64]), .B(A[64]), .Z(n188) );
  ANDN U1872 ( .B(n175), .A(n178), .Z(n1711) );
  ANDN U1873 ( .B(n1713), .A(n119), .Z(n1597) );
  AND U1874 ( .A(B[76]), .B(A[76]), .Z(n119) );
  NAND U1875 ( .A(n1714), .B(n122), .Z(n1713) );
  OR U1876 ( .A(A[76]), .B(B[76]), .Z(n122) );
  NANDN U1877 ( .A(n124), .B(n1715), .Z(n1714) );
  NANDN U1878 ( .A(n126), .B(n1716), .Z(n1715) );
  NANDN U1879 ( .A(n146), .B(n1717), .Z(n1716) );
  NAND U1880 ( .A(n169), .B(n149), .Z(n1717) );
  AND U1881 ( .A(n1718), .B(n1719), .Z(n149) );
  AND U1882 ( .A(n166), .B(n162), .Z(n1719) );
  OR U1883 ( .A(B[68]), .B(A[68]), .Z(n166) );
  AND U1884 ( .A(n157), .B(n153), .Z(n1718) );
  NANDN U1885 ( .A(n174), .B(n1720), .Z(n169) );
  NAND U1886 ( .A(n1721), .B(n175), .Z(n1720) );
  OR U1887 ( .A(B[67]), .B(A[67]), .Z(n175) );
  NANDN U1888 ( .A(n177), .B(n1722), .Z(n1721) );
  NANDN U1889 ( .A(n178), .B(n1723), .Z(n1722) );
  NANDN U1890 ( .A(n181), .B(n1724), .Z(n1723) );
  NAND U1891 ( .A(n184), .B(n186), .Z(n1724) );
  AND U1892 ( .A(A[64]), .B(B[64]), .Z(n186) );
  OR U1893 ( .A(B[65]), .B(A[65]), .Z(n184) );
  AND U1894 ( .A(B[65]), .B(A[65]), .Z(n181) );
  NOR U1895 ( .A(B[66]), .B(A[66]), .Z(n178) );
  AND U1896 ( .A(B[66]), .B(A[66]), .Z(n177) );
  AND U1897 ( .A(B[67]), .B(A[67]), .Z(n174) );
  NANDN U1898 ( .A(n152), .B(n1725), .Z(n146) );
  NAND U1899 ( .A(n1726), .B(n153), .Z(n1725) );
  OR U1900 ( .A(B[71]), .B(A[71]), .Z(n153) );
  NANDN U1901 ( .A(n155), .B(n1727), .Z(n1726) );
  NAND U1902 ( .A(n1728), .B(n157), .Z(n1727) );
  OR U1903 ( .A(B[70]), .B(A[70]), .Z(n157) );
  NANDN U1904 ( .A(n159), .B(n1729), .Z(n1728) );
  NAND U1905 ( .A(n162), .B(n164), .Z(n1729) );
  AND U1906 ( .A(B[68]), .B(A[68]), .Z(n164) );
  OR U1907 ( .A(B[69]), .B(A[69]), .Z(n162) );
  AND U1908 ( .A(B[69]), .B(A[69]), .Z(n159) );
  AND U1909 ( .A(B[70]), .B(A[70]), .Z(n155) );
  AND U1910 ( .A(B[71]), .B(A[71]), .Z(n152) );
  NAND U1911 ( .A(n1730), .B(n1731), .Z(n126) );
  AND U1912 ( .A(n144), .B(n140), .Z(n1731) );
  OR U1913 ( .A(B[72]), .B(A[72]), .Z(n144) );
  AND U1914 ( .A(n135), .B(n131), .Z(n1730) );
  NANDN U1915 ( .A(n130), .B(n1732), .Z(n124) );
  NAND U1916 ( .A(n1733), .B(n131), .Z(n1732) );
  OR U1917 ( .A(B[75]), .B(A[75]), .Z(n131) );
  NANDN U1918 ( .A(n133), .B(n1734), .Z(n1733) );
  NAND U1919 ( .A(n1735), .B(n135), .Z(n1734) );
  OR U1920 ( .A(B[74]), .B(A[74]), .Z(n135) );
  NANDN U1921 ( .A(n137), .B(n1736), .Z(n1735) );
  NAND U1922 ( .A(n140), .B(n142), .Z(n1736) );
  AND U1923 ( .A(B[72]), .B(A[72]), .Z(n142) );
  OR U1924 ( .A(B[73]), .B(A[73]), .Z(n140) );
  AND U1925 ( .A(B[73]), .B(A[73]), .Z(n137) );
  AND U1926 ( .A(B[74]), .B(A[74]), .Z(n133) );
  AND U1927 ( .A(B[75]), .B(A[75]), .Z(n130) );
  NOR U1928 ( .A(B[77]), .B(A[77]), .Z(n116) );
  AND U1929 ( .A(B[77]), .B(A[77]), .Z(n114) );
  NOR U1930 ( .A(B[78]), .B(A[78]), .Z(n111) );
  AND U1931 ( .A(B[78]), .B(A[78]), .Z(n110) );
  NOR U1932 ( .A(B[79]), .B(A[79]), .Z(n107) );
  NOR U1933 ( .A(n85), .B(n41), .Z(n1588) );
  NAND U1934 ( .A(n1737), .B(n1738), .Z(n85) );
  AND U1935 ( .A(n103), .B(n99), .Z(n1738) );
  OR U1936 ( .A(B[80]), .B(A[80]), .Z(n103) );
  ANDN U1937 ( .B(n90), .A(n93), .Z(n1737) );
  ANDN U1938 ( .B(n1739), .A(n34), .Z(n1586) );
  AND U1939 ( .A(B[92]), .B(A[92]), .Z(n34) );
  NAND U1940 ( .A(n1740), .B(n37), .Z(n1739) );
  OR U1941 ( .A(A[92]), .B(B[92]), .Z(n37) );
  NANDN U1942 ( .A(n39), .B(n1741), .Z(n1740) );
  NANDN U1943 ( .A(n41), .B(n1742), .Z(n1741) );
  NANDN U1944 ( .A(n61), .B(n1743), .Z(n1742) );
  NAND U1945 ( .A(n84), .B(n64), .Z(n1743) );
  AND U1946 ( .A(n1744), .B(n1745), .Z(n64) );
  AND U1947 ( .A(n81), .B(n77), .Z(n1745) );
  OR U1948 ( .A(B[84]), .B(A[84]), .Z(n81) );
  AND U1949 ( .A(n72), .B(n68), .Z(n1744) );
  NANDN U1950 ( .A(n89), .B(n1746), .Z(n84) );
  NAND U1951 ( .A(n1747), .B(n90), .Z(n1746) );
  OR U1952 ( .A(B[83]), .B(A[83]), .Z(n90) );
  NANDN U1953 ( .A(n92), .B(n1748), .Z(n1747) );
  NANDN U1954 ( .A(n93), .B(n1749), .Z(n1748) );
  NANDN U1955 ( .A(n96), .B(n1750), .Z(n1749) );
  NAND U1956 ( .A(n99), .B(n101), .Z(n1750) );
  AND U1957 ( .A(A[80]), .B(B[80]), .Z(n101) );
  OR U1958 ( .A(B[81]), .B(A[81]), .Z(n99) );
  AND U1959 ( .A(B[81]), .B(A[81]), .Z(n96) );
  NOR U1960 ( .A(B[82]), .B(A[82]), .Z(n93) );
  AND U1961 ( .A(B[82]), .B(A[82]), .Z(n92) );
  AND U1962 ( .A(B[83]), .B(A[83]), .Z(n89) );
  NANDN U1963 ( .A(n67), .B(n1751), .Z(n61) );
  NAND U1964 ( .A(n1752), .B(n68), .Z(n1751) );
  OR U1965 ( .A(B[87]), .B(A[87]), .Z(n68) );
  NANDN U1966 ( .A(n70), .B(n1753), .Z(n1752) );
  NAND U1967 ( .A(n1754), .B(n72), .Z(n1753) );
  OR U1968 ( .A(B[86]), .B(A[86]), .Z(n72) );
  NANDN U1969 ( .A(n74), .B(n1755), .Z(n1754) );
  NAND U1970 ( .A(n77), .B(n79), .Z(n1755) );
  AND U1971 ( .A(B[84]), .B(A[84]), .Z(n79) );
  OR U1972 ( .A(B[85]), .B(A[85]), .Z(n77) );
  AND U1973 ( .A(B[85]), .B(A[85]), .Z(n74) );
  AND U1974 ( .A(B[86]), .B(A[86]), .Z(n70) );
  AND U1975 ( .A(B[87]), .B(A[87]), .Z(n67) );
  NAND U1976 ( .A(n1756), .B(n1757), .Z(n41) );
  AND U1977 ( .A(n59), .B(n55), .Z(n1757) );
  OR U1978 ( .A(B[88]), .B(A[88]), .Z(n59) );
  AND U1979 ( .A(n50), .B(n46), .Z(n1756) );
  NANDN U1980 ( .A(n45), .B(n1758), .Z(n39) );
  NAND U1981 ( .A(n1759), .B(n46), .Z(n1758) );
  OR U1982 ( .A(B[91]), .B(A[91]), .Z(n46) );
  NANDN U1983 ( .A(n48), .B(n1760), .Z(n1759) );
  NAND U1984 ( .A(n1761), .B(n50), .Z(n1760) );
  OR U1985 ( .A(B[90]), .B(A[90]), .Z(n50) );
  NANDN U1986 ( .A(n52), .B(n1762), .Z(n1761) );
  NAND U1987 ( .A(n55), .B(n57), .Z(n1762) );
  AND U1988 ( .A(B[88]), .B(A[88]), .Z(n57) );
  OR U1989 ( .A(B[89]), .B(A[89]), .Z(n55) );
  AND U1990 ( .A(B[89]), .B(A[89]), .Z(n52) );
  AND U1991 ( .A(B[90]), .B(A[90]), .Z(n48) );
  AND U1992 ( .A(B[91]), .B(A[91]), .Z(n45) );
  NOR U1993 ( .A(B[93]), .B(A[93]), .Z(n31) );
  AND U1994 ( .A(B[93]), .B(A[93]), .Z(n29) );
  NOR U1995 ( .A(B[94]), .B(A[94]), .Z(n26) );
  AND U1996 ( .A(B[94]), .B(A[94]), .Z(n25) );
  NOR U1997 ( .A(B[95]), .B(A[95]), .Z(n22) );
  NAND U1998 ( .A(n1763), .B(n1764), .Z(n1498) );
  AND U1999 ( .A(n13), .B(n8), .Z(n1764) );
  OR U2000 ( .A(B[98]), .B(A[98]), .Z(n8) );
  OR U2001 ( .A(B[97]), .B(A[97]), .Z(n13) );
  AND U2002 ( .A(n4), .B(n18), .Z(n1763) );
  OR U2003 ( .A(B[96]), .B(A[96]), .Z(n18) );
  OR U2004 ( .A(B[99]), .B(A[99]), .Z(n4) );
endmodule


module mult_N256_CC16_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [255:0] B;
  output [271:0] PRODUCT;
  input TC;
  wire   \A1[268] , \A1[267] , \A1[266] , \A1[265] , \A1[264] , \A1[263] ,
         \A1[262] , \A1[261] , \A1[260] , \A1[259] , \A1[258] , \A1[257] ,
         \A1[256] , \A1[255] , \A1[254] , \A1[253] , \A1[252] , \A1[251] ,
         \A1[250] , \A1[249] , \A1[248] , \A1[247] , \A1[246] , \A1[245] ,
         \A1[244] , \A1[243] , \A1[242] , \A1[241] , \A1[240] , \A1[239] ,
         \A1[238] , \A1[237] , \A1[236] , \A1[235] , \A1[234] , \A1[233] ,
         \A1[232] , \A1[231] , \A1[230] , \A1[229] , \A1[228] , \A1[227] ,
         \A1[226] , \A1[225] , \A1[224] , \A1[223] , \A1[222] , \A1[221] ,
         \A1[220] , \A1[219] , \A1[218] , \A1[217] , \A1[216] , \A1[215] ,
         \A1[214] , \A1[213] , \A1[212] , \A1[211] , \A1[210] , \A1[209] ,
         \A1[208] , \A1[207] , \A1[206] , \A1[205] , \A1[204] , \A1[203] ,
         \A1[202] , \A1[201] , \A1[200] , \A1[199] , \A1[198] , \A1[197] ,
         \A1[196] , \A1[195] , \A1[194] , \A1[193] , \A1[192] , \A1[191] ,
         \A1[190] , \A1[189] , \A1[188] , \A1[187] , \A1[186] , \A1[185] ,
         \A1[184] , \A1[183] , \A1[182] , \A1[181] , \A1[180] , \A1[179] ,
         \A1[178] , \A1[177] , \A1[176] , \A1[175] , \A1[174] , \A1[173] ,
         \A1[172] , \A1[171] , \A1[170] , \A1[169] , \A1[168] , \A1[167] ,
         \A1[166] , \A1[165] , \A1[164] , \A1[163] , \A1[162] , \A1[161] ,
         \A1[160] , \A1[159] , \A1[158] , \A1[157] , \A1[156] , \A1[155] ,
         \A1[154] , \A1[153] , \A1[152] , \A1[151] , \A1[150] , \A1[149] ,
         \A1[148] , \A1[147] , \A1[146] , \A1[145] , \A1[144] , \A1[143] ,
         \A1[142] , \A1[141] , \A1[140] , \A1[139] , \A1[138] , \A1[137] ,
         \A1[136] , \A1[135] , \A1[134] , \A1[133] , \A1[132] , \A1[131] ,
         \A1[130] , \A1[129] , \A1[128] , \A1[127] , \A1[126] , \A1[125] ,
         \A1[124] , \A1[123] , \A1[122] , \A1[121] , \A1[120] , \A1[119] ,
         \A1[118] , \A1[117] , \A1[116] , \A1[115] , \A1[114] , \A1[113] ,
         \A1[112] , \A1[111] , \A1[110] , \A1[109] , \A1[108] , \A1[107] ,
         \A1[106] , \A1[105] , \A1[104] , \A1[103] , \A1[102] , \A1[101] ,
         \A1[100] , \A1[99] , \A1[98] , \A1[97] , \A1[96] , \A1[95] , \A1[94] ,
         \A1[93] , \A1[92] , \A1[91] , \A1[90] , \A1[89] , \A1[88] , \A1[87] ,
         \A1[86] , \A1[85] , \A1[84] , \A1[83] , \A1[82] , \A1[81] , \A1[80] ,
         \A1[79] , \A1[78] , \A1[77] , \A1[76] , \A1[75] , \A1[74] , \A1[73] ,
         \A1[72] , \A1[71] , \A1[70] , \A1[69] , \A1[68] , \A1[67] , \A1[66] ,
         \A1[65] , \A1[64] , \A1[63] , \A1[62] , \A1[61] , \A1[60] , \A1[59] ,
         \A1[58] , \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] ,
         \A1[51] , \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[45] ,
         \A1[44] , \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] ,
         \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] ,
         \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] ,
         \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] ,
         \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] ,
         \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] ,
         \A1[2] , \A1[1] , \A1[0] , \A2[269] , \A2[268] , \A2[267] , \A2[266] ,
         \A2[265] , \A2[264] , \A2[263] , \A2[262] , \A2[261] , \A2[260] ,
         \A2[259] , \A2[258] , \A2[257] , \A2[256] , \A2[255] , \A2[254] ,
         \A2[253] , \A2[252] , \A2[251] , \A2[250] , \A2[249] , \A2[248] ,
         \A2[247] , \A2[246] , \A2[245] , \A2[244] , \A2[243] , \A2[242] ,
         \A2[241] , \A2[240] , \A2[239] , \A2[238] , \A2[237] , \A2[236] ,
         \A2[235] , \A2[234] , \A2[233] , \A2[232] , \A2[231] , \A2[230] ,
         \A2[229] , \A2[228] , \A2[227] , \A2[226] , \A2[225] , \A2[224] ,
         \A2[223] , \A2[222] , \A2[221] , \A2[220] , \A2[219] , \A2[218] ,
         \A2[217] , \A2[216] , \A2[215] , \A2[214] , \A2[213] , \A2[212] ,
         \A2[211] , \A2[210] , \A2[209] , \A2[208] , \A2[207] , \A2[206] ,
         \A2[205] , \A2[204] , \A2[203] , \A2[202] , \A2[201] , \A2[200] ,
         \A2[199] , \A2[198] , \A2[197] , \A2[196] , \A2[195] , \A2[194] ,
         \A2[193] , \A2[192] , \A2[191] , \A2[190] , \A2[189] , \A2[188] ,
         \A2[187] , \A2[186] , \A2[185] , \A2[184] , \A2[183] , \A2[182] ,
         \A2[181] , \A2[180] , \A2[179] , \A2[178] , \A2[177] , \A2[176] ,
         \A2[175] , \A2[174] , \A2[173] , \A2[172] , \A2[171] , \A2[170] ,
         \A2[169] , \A2[168] , \A2[167] , \A2[166] , \A2[165] , \A2[164] ,
         \A2[163] , \A2[162] , \A2[161] , \A2[160] , \A2[159] , \A2[158] ,
         \A2[157] , \A2[156] , \A2[155] , \A2[154] , \A2[153] , \A2[152] ,
         \A2[151] , \A2[150] , \A2[149] , \A2[148] , \A2[147] , \A2[146] ,
         \A2[145] , \A2[144] , \A2[143] , \A2[142] , \A2[141] , \A2[140] ,
         \A2[139] , \A2[138] , \A2[137] , \A2[136] , \A2[135] , \A2[134] ,
         \A2[133] , \A2[132] , \A2[131] , \A2[130] , \A2[129] , \A2[128] ,
         \A2[127] , \A2[126] , \A2[125] , \A2[124] , \A2[123] , \A2[122] ,
         \A2[121] , \A2[120] , \A2[119] , \A2[118] , \A2[117] , \A2[116] ,
         \A2[115] , \A2[114] , \A2[113] , \A2[112] , \A2[111] , \A2[110] ,
         \A2[109] , \A2[108] , \A2[107] , \A2[106] , \A2[105] , \A2[104] ,
         \A2[103] , \A2[102] , \A2[101] , \A2[100] , \A2[99] , \A2[98] ,
         \A2[97] , \A2[96] , \A2[95] , \A2[94] , \A2[93] , \A2[92] , \A2[91] ,
         \A2[90] , \A2[89] , \A2[88] , \A2[87] , \A2[86] , \A2[85] , \A2[84] ,
         \A2[83] , \A2[82] , \A2[81] , \A2[80] , \A2[79] , \A2[78] , \A2[77] ,
         \A2[76] , \A2[75] , \A2[74] , \A2[73] , \A2[72] , \A2[71] , \A2[70] ,
         \A2[69] , \A2[68] , \A2[67] , \A2[66] , \A2[65] , \A2[64] , \A2[63] ,
         \A2[62] , \A2[61] , \A2[60] , \A2[59] , \A2[58] , \A2[57] , \A2[56] ,
         \A2[55] , \A2[54] , \A2[53] , \A2[52] , \A2[51] , \A2[50] , \A2[49] ,
         \A2[48] , \A2[47] , \A2[46] , \A2[45] , \A2[44] , \A2[43] , \A2[42] ,
         \A2[41] , \A2[40] , \A2[39] , \A2[38] , \A2[37] , \A2[36] , \A2[35] ,
         \A2[34] , \A2[33] , \A2[32] , \A2[31] , \A2[30] , \A2[29] , \A2[28] ,
         \A2[27] , \A2[26] , \A2[25] , \A2[24] , \A2[23] , \A2[22] , \A2[21] ,
         \A2[20] , \A2[19] , \A2[18] , \A2[17] , \A2[16] , \A2[15] , n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
         n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
         n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
         n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
         n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275,
         n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
         n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
         n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
         n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
         n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
         n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331,
         n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
         n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347,
         n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
         n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
         n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
         n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
         n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
         n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395,
         n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
         n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
         n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
         n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443,
         n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451,
         n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
         n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467,
         n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
         n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
         n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
         n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
         n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
         n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
         n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539,
         n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
         n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
         n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563,
         n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
         n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
         n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
         n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
         n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
         n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
         n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
         n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
         n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
         n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
         n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707,
         n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
         n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
         n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731,
         n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
         n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
         n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755,
         n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
         n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
         n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
         n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
         n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
         n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
         n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
         n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
         n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827,
         n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
         n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
         n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
         n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
         n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
         n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875,
         n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
         n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
         n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899,
         n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
         n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
         n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
         n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
         n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
         n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947,
         n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
         n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971,
         n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
         n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
         n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
         n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
         n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
         n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
         n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
         n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
         n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
         n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115,
         n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
         n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
         n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
         n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
         n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
         n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163,
         n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
         n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
         n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
         n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
         n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211,
         n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
         n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
         n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
         n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243,
         n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
         n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
         n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355,
         n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
         n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
         n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
         n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
         n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
         n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
         n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
         n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
         n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
         n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
         n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
         n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
         n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
         n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
         n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
         n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
         n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
         n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
         n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
         n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
         n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
         n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
         n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
         n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
         n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
         n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
         n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
         n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787,
         n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
         n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
         n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
         n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
         n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
         n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
         n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003,
         n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
         n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
         n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027,
         n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035,
         n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
         n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051,
         n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
         n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
         n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075,
         n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
         n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
         n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099,
         n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
         n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
         n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
         n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
         n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147,
         n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
         n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
         n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171,
         n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
         n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
         n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195,
         n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
         n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
         n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219,
         n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
         n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
         n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243,
         n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
         n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
         n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267,
         n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275,
         n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
         n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
         n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
         n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315,
         n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
         n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
         n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
         n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
         n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363,
         n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
         n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
         n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387,
         n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419,
         n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
         n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435,
         n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
         n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
         n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459,
         n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
         n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483,
         n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491,
         n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
         n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507,
         n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
         n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
         n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531,
         n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
         n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
         n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555,
         n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
         n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
         n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579,
         n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
         n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
         n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603,
         n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
         n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
         n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627,
         n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635,
         n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
         n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651,
         n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
         n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
         n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
         n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
         n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
         n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699,
         n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707,
         n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
         n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
         n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
         n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
         n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
         n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
         n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771,
         n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779,
         n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
         n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
         n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
         n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
         n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819,
         n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827,
         n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
         n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843,
         n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851,
         n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
         n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
         n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
         n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
         n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
         n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
         n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
         n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915,
         n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
         n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
         n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
         n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
         n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987,
         n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
         n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
         n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
         n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
         n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
         n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035,
         n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
         n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
         n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059,
         n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067,
         n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
         n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
         n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
         n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
         n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107,
         n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
         n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
         n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131,
         n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139,
         n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
         n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155,
         n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
         n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
         n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179,
         n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
         n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
         n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
         n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211,
         n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
         n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227,
         n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
         n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
         n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
         n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
         n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
         n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275,
         n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283,
         n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
         n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299,
         n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
         n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
         n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323,
         n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
         n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
         n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
         n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
         n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
         n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
         n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395,
         n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403,
         n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
         n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
         n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427,
         n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
         n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443,
         n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
         n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459,
         n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467,
         n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499,
         n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
         n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
         n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539,
         n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
         n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
         n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
         n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
         n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
         n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611,
         n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
         n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
         n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659,
         n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755,
         n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
         n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
         n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
         n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803,
         n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
         n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
         n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
         n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
         n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
         n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
         n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875,
         n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
         n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
         n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
         n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
         n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
         n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947,
         n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
         n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
         n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971,
         n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
         n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003,
         n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
         n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019,
         n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
         n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
         n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043,
         n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051,
         n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
         n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
         n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075,
         n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083,
         n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091,
         n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
         n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
         n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115,
         n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123,
         n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
         n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139,
         n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147,
         n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
         n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163,
         n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
         n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179,
         n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187,
         n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195,
         n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
         n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211,
         n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219,
         n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227,
         n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235,
         n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
         n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
         n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259,
         n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267,
         n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
         n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283,
         n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291,
         n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
         n26300, n26301, n26302, n26303, n26304;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  mult_N256_CC16_DW01_add_0 FS_1 ( .A({1'b0, \A1[268] , \A1[267] , \A1[266] , 
        \A1[265] , \A1[264] , \A1[263] , \A1[262] , \A1[261] , \A1[260] , 
        \A1[259] , \A1[258] , \A1[257] , \A1[256] , \A1[255] , \A1[254] , 
        \A1[253] , \A1[252] , \A1[251] , \A1[250] , \A1[249] , \A1[248] , 
        \A1[247] , \A1[246] , \A1[245] , \A1[244] , \A1[243] , \A1[242] , 
        \A1[241] , \A1[240] , \A1[239] , \A1[238] , \A1[237] , \A1[236] , 
        \A1[235] , \A1[234] , \A1[233] , \A1[232] , \A1[231] , \A1[230] , 
        \A1[229] , \A1[228] , \A1[227] , \A1[226] , \A1[225] , \A1[224] , 
        \A1[223] , \A1[222] , \A1[221] , \A1[220] , \A1[219] , \A1[218] , 
        \A1[217] , \A1[216] , \A1[215] , \A1[214] , \A1[213] , \A1[212] , 
        \A1[211] , \A1[210] , \A1[209] , \A1[208] , \A1[207] , \A1[206] , 
        \A1[205] , \A1[204] , \A1[203] , \A1[202] , \A1[201] , \A1[200] , 
        \A1[199] , \A1[198] , \A1[197] , \A1[196] , \A1[195] , \A1[194] , 
        \A1[193] , \A1[192] , \A1[191] , \A1[190] , \A1[189] , \A1[188] , 
        \A1[187] , \A1[186] , \A1[185] , \A1[184] , \A1[183] , \A1[182] , 
        \A1[181] , \A1[180] , \A1[179] , \A1[178] , \A1[177] , \A1[176] , 
        \A1[175] , \A1[174] , \A1[173] , \A1[172] , \A1[171] , \A1[170] , 
        \A1[169] , \A1[168] , \A1[167] , \A1[166] , \A1[165] , \A1[164] , 
        \A1[163] , \A1[162] , \A1[161] , \A1[160] , \A1[159] , \A1[158] , 
        \A1[157] , \A1[156] , \A1[155] , \A1[154] , \A1[153] , \A1[152] , 
        \A1[151] , \A1[150] , \A1[149] , \A1[148] , \A1[147] , \A1[146] , 
        \A1[145] , \A1[144] , \A1[143] , \A1[142] , \A1[141] , \A1[140] , 
        \A1[139] , \A1[138] , \A1[137] , \A1[136] , \A1[135] , \A1[134] , 
        \A1[133] , \A1[132] , \A1[131] , \A1[130] , \A1[129] , \A1[128] , 
        \A1[127] , \A1[126] , \A1[125] , \A1[124] , \A1[123] , \A1[122] , 
        \A1[121] , \A1[120] , \A1[119] , \A1[118] , \A1[117] , \A1[116] , 
        \A1[115] , \A1[114] , \A1[113] , \A1[112] , \A1[111] , \A1[110] , 
        \A1[109] , \A1[108] , \A1[107] , \A1[106] , \A1[105] , \A1[104] , 
        \A1[103] , \A1[102] , \A1[101] , \A1[100] , \A1[99] , \A1[98] , 
        \A1[97] , \A1[96] , \A1[95] , \A1[94] , \A1[93] , \A1[92] , \A1[91] , 
        \A1[90] , \A1[89] , \A1[88] , \A1[87] , \A1[86] , \A1[85] , \A1[84] , 
        \A1[83] , \A1[82] , \A1[81] , \A1[80] , \A1[79] , \A1[78] , \A1[77] , 
        \A1[76] , \A1[75] , \A1[74] , \A1[73] , \A1[72] , \A1[71] , \A1[70] , 
        \A1[69] , \A1[68] , \A1[67] , \A1[66] , \A1[65] , \A1[64] , \A1[63] , 
        \A1[62] , \A1[61] , \A1[60] , \A1[59] , \A1[58] , \A1[57] , \A1[56] , 
        \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] , \A1[49] , 
        \A1[48] , \A1[47] , \A1[46] , \A1[45] , \A1[44] , \A1[43] , \A1[42] , 
        \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , 
        \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , 
        \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , 
        \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , 
        \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , 
        \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({
        \A2[269] , \A2[268] , \A2[267] , \A2[266] , \A2[265] , \A2[264] , 
        \A2[263] , \A2[262] , \A2[261] , \A2[260] , \A2[259] , \A2[258] , 
        \A2[257] , \A2[256] , \A2[255] , \A2[254] , \A2[253] , \A2[252] , 
        \A2[251] , \A2[250] , \A2[249] , \A2[248] , \A2[247] , \A2[246] , 
        \A2[245] , \A2[244] , \A2[243] , \A2[242] , \A2[241] , \A2[240] , 
        \A2[239] , \A2[238] , \A2[237] , \A2[236] , \A2[235] , \A2[234] , 
        \A2[233] , \A2[232] , \A2[231] , \A2[230] , \A2[229] , \A2[228] , 
        \A2[227] , \A2[226] , \A2[225] , \A2[224] , \A2[223] , \A2[222] , 
        \A2[221] , \A2[220] , \A2[219] , \A2[218] , \A2[217] , \A2[216] , 
        \A2[215] , \A2[214] , \A2[213] , \A2[212] , \A2[211] , \A2[210] , 
        \A2[209] , \A2[208] , \A2[207] , \A2[206] , \A2[205] , \A2[204] , 
        \A2[203] , \A2[202] , \A2[201] , \A2[200] , \A2[199] , \A2[198] , 
        \A2[197] , \A2[196] , \A2[195] , \A2[194] , \A2[193] , \A2[192] , 
        \A2[191] , \A2[190] , \A2[189] , \A2[188] , \A2[187] , \A2[186] , 
        \A2[185] , \A2[184] , \A2[183] , \A2[182] , \A2[181] , \A2[180] , 
        \A2[179] , \A2[178] , \A2[177] , \A2[176] , \A2[175] , \A2[174] , 
        \A2[173] , \A2[172] , \A2[171] , \A2[170] , \A2[169] , \A2[168] , 
        \A2[167] , \A2[166] , \A2[165] , \A2[164] , \A2[163] , \A2[162] , 
        \A2[161] , \A2[160] , \A2[159] , \A2[158] , \A2[157] , \A2[156] , 
        \A2[155] , \A2[154] , \A2[153] , \A2[152] , \A2[151] , \A2[150] , 
        \A2[149] , \A2[148] , \A2[147] , \A2[146] , \A2[145] , \A2[144] , 
        \A2[143] , \A2[142] , \A2[141] , \A2[140] , \A2[139] , \A2[138] , 
        \A2[137] , \A2[136] , \A2[135] , \A2[134] , \A2[133] , \A2[132] , 
        \A2[131] , \A2[130] , \A2[129] , \A2[128] , \A2[127] , \A2[126] , 
        \A2[125] , \A2[124] , \A2[123] , \A2[122] , \A2[121] , \A2[120] , 
        \A2[119] , \A2[118] , \A2[117] , \A2[116] , \A2[115] , \A2[114] , 
        \A2[113] , \A2[112] , \A2[111] , \A2[110] , \A2[109] , \A2[108] , 
        \A2[107] , \A2[106] , \A2[105] , \A2[104] , \A2[103] , \A2[102] , 
        \A2[101] , \A2[100] , \A2[99] , \A2[98] , \A2[97] , \A2[96] , \A2[95] , 
        \A2[94] , \A2[93] , \A2[92] , \A2[91] , \A2[90] , \A2[89] , \A2[88] , 
        \A2[87] , \A2[86] , \A2[85] , \A2[84] , \A2[83] , \A2[82] , \A2[81] , 
        \A2[80] , \A2[79] , \A2[78] , \A2[77] , \A2[76] , \A2[75] , \A2[74] , 
        \A2[73] , \A2[72] , \A2[71] , \A2[70] , \A2[69] , \A2[68] , \A2[67] , 
        \A2[66] , \A2[65] , \A2[64] , \A2[63] , \A2[62] , \A2[61] , \A2[60] , 
        \A2[59] , \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , 
        \A2[52] , \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , \A2[46] , 
        \A2[45] , \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , 
        \A2[38] , \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , 
        \A2[31] , \A2[30] , \A2[29] , \A2[28] , \A2[27] , \A2[26] , \A2[25] , 
        \A2[24] , \A2[23] , \A2[22] , \A2[21] , \A2[20] , \A2[19] , \A2[18] , 
        \A2[17] , \A2[16] , \A2[15] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, PRODUCT[255:2]})
         );
  OR U2 ( .A(n10237), .B(n10236), .Z(n10232) );
  OR U3 ( .A(n26292), .B(n26289), .Z(n26294) );
  NANDN U4 ( .A(n1122), .B(n1121), .Z(n1117) );
  NAND U5 ( .A(B[255]), .B(n8321), .Z(n8220) );
  NANDN U6 ( .A(n881), .B(n880), .Z(n876) );
  OR U7 ( .A(n25782), .B(n25780), .Z(n25852) );
  NANDN U8 ( .A(n707), .B(n706), .Z(n702) );
  OR U9 ( .A(n25750), .B(n25748), .Z(n25840) );
  NANDN U10 ( .A(n596), .B(n595), .Z(n591) );
  OR U11 ( .A(n24361), .B(n24358), .Z(n24412) );
  OR U12 ( .A(n10439), .B(n10438), .Z(n10434) );
  OR U13 ( .A(n10641), .B(n10640), .Z(n10636) );
  OR U14 ( .A(n10843), .B(n10842), .Z(n10838) );
  OR U15 ( .A(n11146), .B(n11145), .Z(n11141) );
  OR U16 ( .A(n11348), .B(n11347), .Z(n11343) );
  OR U17 ( .A(n11550), .B(n11549), .Z(n11545) );
  OR U18 ( .A(n11752), .B(n11751), .Z(n11747) );
  OR U19 ( .A(n11954), .B(n11953), .Z(n11949) );
  OR U20 ( .A(n12257), .B(n12256), .Z(n12252) );
  OR U21 ( .A(n12459), .B(n12458), .Z(n12454) );
  OR U22 ( .A(n12661), .B(n12660), .Z(n12656) );
  OR U23 ( .A(n12863), .B(n12862), .Z(n12858) );
  OR U24 ( .A(n13065), .B(n13064), .Z(n13060) );
  OR U25 ( .A(n13368), .B(n13367), .Z(n13363) );
  OR U26 ( .A(n13570), .B(n13569), .Z(n13565) );
  OR U27 ( .A(n13772), .B(n13771), .Z(n13767) );
  OR U28 ( .A(n13974), .B(n13973), .Z(n13969) );
  OR U29 ( .A(n14176), .B(n14175), .Z(n14171) );
  OR U30 ( .A(n14483), .B(n14482), .Z(n14478) );
  OR U31 ( .A(n14685), .B(n14684), .Z(n14680) );
  OR U32 ( .A(n14887), .B(n14886), .Z(n14882) );
  OR U33 ( .A(n15089), .B(n15088), .Z(n15084) );
  OR U34 ( .A(n15291), .B(n15290), .Z(n15286) );
  OR U35 ( .A(n15594), .B(n15593), .Z(n15589) );
  OR U36 ( .A(n15796), .B(n15795), .Z(n15791) );
  OR U37 ( .A(n15998), .B(n15997), .Z(n15993) );
  OR U38 ( .A(n16200), .B(n16199), .Z(n16195) );
  OR U39 ( .A(n16402), .B(n16401), .Z(n16397) );
  OR U40 ( .A(n16705), .B(n16704), .Z(n16700) );
  OR U41 ( .A(n16907), .B(n16906), .Z(n16902) );
  OR U42 ( .A(n17109), .B(n17108), .Z(n17104) );
  OR U43 ( .A(n17311), .B(n17310), .Z(n17306) );
  OR U44 ( .A(n17513), .B(n17512), .Z(n17508) );
  OR U45 ( .A(n17816), .B(n17815), .Z(n17811) );
  OR U46 ( .A(n18018), .B(n18017), .Z(n18013) );
  OR U47 ( .A(n18220), .B(n18219), .Z(n18215) );
  OR U48 ( .A(n18422), .B(n18421), .Z(n18417) );
  OR U49 ( .A(n18624), .B(n18623), .Z(n18619) );
  OR U50 ( .A(n18927), .B(n18926), .Z(n18922) );
  OR U51 ( .A(n19129), .B(n19128), .Z(n19124) );
  OR U52 ( .A(n19331), .B(n19330), .Z(n19326) );
  OR U53 ( .A(n19533), .B(n19532), .Z(n19528) );
  OR U54 ( .A(n19735), .B(n19734), .Z(n19730) );
  OR U55 ( .A(n20038), .B(n20037), .Z(n20033) );
  OR U56 ( .A(n20240), .B(n20239), .Z(n20235) );
  OR U57 ( .A(n20442), .B(n20441), .Z(n20437) );
  OR U58 ( .A(n20644), .B(n20643), .Z(n20639) );
  OR U59 ( .A(n20846), .B(n20845), .Z(n20841) );
  OR U60 ( .A(n21143), .B(n21142), .Z(n21138) );
  OR U61 ( .A(n21345), .B(n21344), .Z(n21340) );
  OR U62 ( .A(n21547), .B(n21546), .Z(n21542) );
  OR U63 ( .A(n21749), .B(n21748), .Z(n21744) );
  OR U64 ( .A(n21951), .B(n21950), .Z(n21946) );
  OR U65 ( .A(n22241), .B(n22240), .Z(n22236) );
  OR U66 ( .A(n22443), .B(n22442), .Z(n22438) );
  OR U67 ( .A(n22645), .B(n22644), .Z(n22640) );
  OR U68 ( .A(n22847), .B(n22846), .Z(n22842) );
  OR U69 ( .A(n23049), .B(n23048), .Z(n23044) );
  OR U70 ( .A(n23332), .B(n23331), .Z(n23327) );
  OR U71 ( .A(n23534), .B(n23533), .Z(n23529) );
  OR U72 ( .A(n23736), .B(n23735), .Z(n23731) );
  OR U73 ( .A(n23938), .B(n23937), .Z(n23933) );
  OR U74 ( .A(n24140), .B(n24139), .Z(n24135) );
  OR U75 ( .A(n24735), .B(n24734), .Z(n24730) );
  OR U76 ( .A(n24937), .B(n24936), .Z(n24932) );
  OR U77 ( .A(n25139), .B(n25138), .Z(n25134) );
  OR U78 ( .A(n25341), .B(n25340), .Z(n25336) );
  OR U79 ( .A(n25543), .B(n25542), .Z(n25538) );
  NANDN U80 ( .A(n1316), .B(n1319), .Z(n25828) );
  OR U81 ( .A(n26274), .B(n26271), .Z(n26283) );
  OR U82 ( .A(n26217), .B(n26214), .Z(n26240) );
  OR U83 ( .A(n26132), .B(n26129), .Z(n26169) );
  OR U84 ( .A(n26019), .B(n26016), .Z(n26070) );
  OR U85 ( .A(n25878), .B(n25875), .Z(n25943) );
  OR U86 ( .A(n1619), .B(n1618), .Z(n1614) );
  OR U87 ( .A(n1821), .B(n1820), .Z(n1816) );
  OR U88 ( .A(n2026), .B(n2025), .Z(n2021) );
  OR U89 ( .A(n2228), .B(n2227), .Z(n2223) );
  OR U90 ( .A(n2430), .B(n2429), .Z(n2425) );
  OR U91 ( .A(n2632), .B(n2631), .Z(n2627) );
  OR U92 ( .A(n2834), .B(n2833), .Z(n2829) );
  OR U93 ( .A(n3040), .B(n3039), .Z(n3035) );
  OR U94 ( .A(n3242), .B(n3241), .Z(n3237) );
  OR U95 ( .A(n3444), .B(n3443), .Z(n3439) );
  OR U96 ( .A(n3646), .B(n3645), .Z(n3641) );
  OR U97 ( .A(n3848), .B(n3847), .Z(n3843) );
  OR U98 ( .A(n4053), .B(n4052), .Z(n4048) );
  OR U99 ( .A(n4255), .B(n4254), .Z(n4250) );
  OR U100 ( .A(n4457), .B(n4456), .Z(n4452) );
  OR U101 ( .A(n4659), .B(n4658), .Z(n4654) );
  OR U102 ( .A(n4861), .B(n4860), .Z(n4856) );
  OR U103 ( .A(n5067), .B(n5066), .Z(n5062) );
  OR U104 ( .A(n5269), .B(n5268), .Z(n5264) );
  OR U105 ( .A(n5471), .B(n5470), .Z(n5466) );
  OR U106 ( .A(n5673), .B(n5672), .Z(n5668) );
  OR U107 ( .A(n5875), .B(n5874), .Z(n5870) );
  OR U108 ( .A(n6080), .B(n6079), .Z(n6075) );
  OR U109 ( .A(n6282), .B(n6281), .Z(n6277) );
  OR U110 ( .A(n6484), .B(n6483), .Z(n6479) );
  OR U111 ( .A(n6686), .B(n6685), .Z(n6681) );
  OR U112 ( .A(n6888), .B(n6887), .Z(n6883) );
  OR U113 ( .A(n7094), .B(n7093), .Z(n7089) );
  OR U114 ( .A(n7296), .B(n7295), .Z(n7291) );
  OR U115 ( .A(n7805), .B(n7804), .Z(n7800) );
  OR U116 ( .A(n9934), .B(n9933), .Z(n9929) );
  OR U117 ( .A(n12156), .B(n12155), .Z(n12151) );
  OR U118 ( .A(n14382), .B(n14381), .Z(n14377) );
  OR U119 ( .A(n16604), .B(n16603), .Z(n16599) );
  OR U120 ( .A(n10136), .B(n10135), .Z(n10131) );
  OR U121 ( .A(n18826), .B(n18825), .Z(n18821) );
  OR U122 ( .A(n21048), .B(n21047), .Z(n21043) );
  NANDN U123 ( .A(n1036), .B(n1035), .Z(n1031) );
  OR U124 ( .A(n9833), .B(n9832), .Z(n9828) );
  OR U125 ( .A(n8319), .B(n8318), .Z(n8314) );
  OR U126 ( .A(n9631), .B(n9630), .Z(n9626) );
  OR U127 ( .A(n8520), .B(n8519), .Z(n8515) );
  OR U128 ( .A(n9429), .B(n9428), .Z(n9424) );
  OR U129 ( .A(n9227), .B(n9226), .Z(n9222) );
  OR U130 ( .A(n8722), .B(n8721), .Z(n8717) );
  OR U131 ( .A(n9025), .B(n9024), .Z(n9020) );
  OR U132 ( .A(n25798), .B(n25796), .Z(n25858) );
  OR U133 ( .A(n23237), .B(n23236), .Z(n23232) );
  NANDN U134 ( .A(n816), .B(n815), .Z(n811) );
  OR U135 ( .A(n24616), .B(n24613), .Z(n24625) );
  OR U136 ( .A(n24559), .B(n24556), .Z(n24582) );
  NANDN U137 ( .A(n663), .B(n662), .Z(n658) );
  NANDN U138 ( .A(n25666), .B(n25665), .Z(n25661) );
  OR U139 ( .A(n24474), .B(n24471), .Z(n24511) );
  OR U140 ( .A(n573), .B(n576), .Z(n25741) );
  NANDN U141 ( .A(n572), .B(n571), .Z(n567) );
  OR U142 ( .A(n24304), .B(n24302), .Z(n24347) );
  OR U143 ( .A(n24274), .B(n24272), .Z(n24335) );
  OR U144 ( .A(n10338), .B(n10337), .Z(n10333) );
  OR U145 ( .A(n10540), .B(n10539), .Z(n10535) );
  OR U146 ( .A(n10742), .B(n10741), .Z(n10737) );
  OR U147 ( .A(n10944), .B(n10943), .Z(n10939) );
  OR U148 ( .A(n11247), .B(n11246), .Z(n11242) );
  OR U149 ( .A(n11449), .B(n11448), .Z(n11444) );
  OR U150 ( .A(n11651), .B(n11650), .Z(n11646) );
  OR U151 ( .A(n11853), .B(n11852), .Z(n11848) );
  OR U152 ( .A(n12055), .B(n12054), .Z(n12050) );
  OR U153 ( .A(n12358), .B(n12357), .Z(n12353) );
  OR U154 ( .A(n12560), .B(n12559), .Z(n12555) );
  OR U155 ( .A(n12762), .B(n12761), .Z(n12757) );
  OR U156 ( .A(n12964), .B(n12963), .Z(n12959) );
  OR U157 ( .A(n13166), .B(n13165), .Z(n13161) );
  OR U158 ( .A(n13469), .B(n13468), .Z(n13464) );
  OR U159 ( .A(n13671), .B(n13670), .Z(n13666) );
  OR U160 ( .A(n13873), .B(n13872), .Z(n13868) );
  OR U161 ( .A(n14075), .B(n14074), .Z(n14070) );
  OR U162 ( .A(n14277), .B(n14276), .Z(n14272) );
  OR U163 ( .A(n14584), .B(n14583), .Z(n14579) );
  OR U164 ( .A(n14786), .B(n14785), .Z(n14781) );
  OR U165 ( .A(n14988), .B(n14987), .Z(n14983) );
  OR U166 ( .A(n15190), .B(n15189), .Z(n15185) );
  OR U167 ( .A(n15392), .B(n15391), .Z(n15387) );
  OR U168 ( .A(n15695), .B(n15694), .Z(n15690) );
  OR U169 ( .A(n15897), .B(n15896), .Z(n15892) );
  OR U170 ( .A(n16099), .B(n16098), .Z(n16094) );
  OR U171 ( .A(n16301), .B(n16300), .Z(n16296) );
  OR U172 ( .A(n16503), .B(n16502), .Z(n16498) );
  OR U173 ( .A(n16806), .B(n16805), .Z(n16801) );
  OR U174 ( .A(n17008), .B(n17007), .Z(n17003) );
  OR U175 ( .A(n17210), .B(n17209), .Z(n17205) );
  OR U176 ( .A(n17412), .B(n17411), .Z(n17407) );
  OR U177 ( .A(n17614), .B(n17613), .Z(n17609) );
  OR U178 ( .A(n17917), .B(n17916), .Z(n17912) );
  OR U179 ( .A(n18119), .B(n18118), .Z(n18114) );
  OR U180 ( .A(n18321), .B(n18320), .Z(n18316) );
  OR U181 ( .A(n18523), .B(n18522), .Z(n18518) );
  OR U182 ( .A(n18725), .B(n18724), .Z(n18720) );
  OR U183 ( .A(n19028), .B(n19027), .Z(n19023) );
  OR U184 ( .A(n19230), .B(n19229), .Z(n19225) );
  OR U185 ( .A(n19432), .B(n19431), .Z(n19427) );
  OR U186 ( .A(n19634), .B(n19633), .Z(n19629) );
  OR U187 ( .A(n19836), .B(n19835), .Z(n19831) );
  OR U188 ( .A(n20139), .B(n20138), .Z(n20134) );
  OR U189 ( .A(n20341), .B(n20340), .Z(n20336) );
  OR U190 ( .A(n20543), .B(n20542), .Z(n20538) );
  OR U191 ( .A(n20745), .B(n20744), .Z(n20740) );
  OR U192 ( .A(n20947), .B(n20946), .Z(n20942) );
  OR U193 ( .A(n21244), .B(n21243), .Z(n21239) );
  OR U194 ( .A(n21446), .B(n21445), .Z(n21441) );
  OR U195 ( .A(n21648), .B(n21647), .Z(n21643) );
  OR U196 ( .A(n21850), .B(n21849), .Z(n21845) );
  OR U197 ( .A(n22052), .B(n22051), .Z(n22047) );
  OR U198 ( .A(n22342), .B(n22341), .Z(n22337) );
  OR U199 ( .A(n22544), .B(n22543), .Z(n22539) );
  OR U200 ( .A(n22746), .B(n22745), .Z(n22741) );
  OR U201 ( .A(n22948), .B(n22947), .Z(n22943) );
  OR U202 ( .A(n23150), .B(n23149), .Z(n23145) );
  OR U203 ( .A(n23433), .B(n23432), .Z(n23428) );
  OR U204 ( .A(n23635), .B(n23634), .Z(n23630) );
  OR U205 ( .A(n23837), .B(n23836), .Z(n23832) );
  OR U206 ( .A(n24039), .B(n24038), .Z(n24034) );
  OR U207 ( .A(n24241), .B(n24240), .Z(n24236) );
  OR U208 ( .A(n24836), .B(n24835), .Z(n24831) );
  OR U209 ( .A(n25038), .B(n25037), .Z(n25033) );
  OR U210 ( .A(n25240), .B(n25239), .Z(n25235) );
  OR U211 ( .A(n25442), .B(n25441), .Z(n25437) );
  OR U212 ( .A(n25644), .B(n25643), .Z(n25639) );
  OR U213 ( .A(n26249), .B(n26246), .Z(n26265) );
  OR U214 ( .A(n26178), .B(n26175), .Z(n26208) );
  OR U215 ( .A(n26079), .B(n26076), .Z(n26123) );
  OR U216 ( .A(n25952), .B(n25949), .Z(n26010) );
  OR U217 ( .A(n1416), .B(n1415), .Z(n1411) );
  OR U218 ( .A(n1518), .B(n1517), .Z(n1513) );
  OR U219 ( .A(n1720), .B(n1719), .Z(n1715) );
  OR U220 ( .A(n1922), .B(n1921), .Z(n1917) );
  OR U221 ( .A(n2127), .B(n2126), .Z(n2122) );
  OR U222 ( .A(n2329), .B(n2328), .Z(n2324) );
  OR U223 ( .A(n2531), .B(n2530), .Z(n2526) );
  OR U224 ( .A(n2733), .B(n2732), .Z(n2728) );
  OR U225 ( .A(n2935), .B(n2934), .Z(n2930) );
  OR U226 ( .A(n3141), .B(n3140), .Z(n3136) );
  OR U227 ( .A(n3343), .B(n3342), .Z(n3338) );
  OR U228 ( .A(n3545), .B(n3544), .Z(n3540) );
  OR U229 ( .A(n3747), .B(n3746), .Z(n3742) );
  OR U230 ( .A(n3949), .B(n3948), .Z(n3944) );
  OR U231 ( .A(n4154), .B(n4153), .Z(n4149) );
  OR U232 ( .A(n4356), .B(n4355), .Z(n4351) );
  OR U233 ( .A(n4558), .B(n4557), .Z(n4553) );
  OR U234 ( .A(n4760), .B(n4759), .Z(n4755) );
  OR U235 ( .A(n4962), .B(n4961), .Z(n4957) );
  OR U236 ( .A(n5168), .B(n5167), .Z(n5163) );
  OR U237 ( .A(n5370), .B(n5369), .Z(n5365) );
  OR U238 ( .A(n5572), .B(n5571), .Z(n5567) );
  OR U239 ( .A(n5774), .B(n5773), .Z(n5769) );
  OR U240 ( .A(n5976), .B(n5975), .Z(n5971) );
  OR U241 ( .A(n6181), .B(n6180), .Z(n6176) );
  OR U242 ( .A(n6383), .B(n6382), .Z(n6378) );
  OR U243 ( .A(n6585), .B(n6584), .Z(n6580) );
  OR U244 ( .A(n6787), .B(n6786), .Z(n6782) );
  OR U245 ( .A(n6989), .B(n6988), .Z(n6984) );
  OR U246 ( .A(n7195), .B(n7194), .Z(n7190) );
  OR U247 ( .A(n7397), .B(n7396), .Z(n7392) );
  OR U248 ( .A(n8823), .B(n8822), .Z(n8818) );
  OR U249 ( .A(n11045), .B(n11044), .Z(n11040) );
  OR U250 ( .A(n13267), .B(n13266), .Z(n13262) );
  OR U251 ( .A(n15493), .B(n15492), .Z(n15488) );
  OR U252 ( .A(n17715), .B(n17714), .Z(n17710) );
  NANDN U253 ( .A(n1215), .B(n1214), .Z(n1210) );
  OR U254 ( .A(n10035), .B(n10034), .Z(n10030) );
  NANDN U255 ( .A(n25722), .B(n25721), .Z(n25717) );
  OR U256 ( .A(n25814), .B(n25812), .Z(n25864) );
  OR U257 ( .A(n19937), .B(n19936), .Z(n19932) );
  OR U258 ( .A(n9732), .B(n9731), .Z(n9727) );
  OR U259 ( .A(n8419), .B(n8418), .Z(n8414) );
  OR U260 ( .A(n9530), .B(n9529), .Z(n9525) );
  OR U261 ( .A(n9328), .B(n9327), .Z(n9323) );
  OR U262 ( .A(n8621), .B(n8620), .Z(n8616) );
  OR U263 ( .A(n9126), .B(n9125), .Z(n9121) );
  OR U264 ( .A(n8924), .B(n8923), .Z(n8919) );
  OR U265 ( .A(n22146), .B(n22145), .Z(n22141) );
  NANDN U266 ( .A(n25708), .B(n25707), .Z(n25703) );
  NANDN U267 ( .A(n953), .B(n952), .Z(n948) );
  NANDN U268 ( .A(n8127), .B(n8124), .Z(n8123) );
  OR U269 ( .A(n24634), .B(n24631), .Z(n24636) );
  NANDN U270 ( .A(n25694), .B(n25693), .Z(n25689) );
  NANDN U271 ( .A(n758), .B(n757), .Z(n753) );
  OR U272 ( .A(n24591), .B(n24588), .Z(n24607) );
  NANDN U273 ( .A(n25680), .B(n25679), .Z(n25675) );
  OR U274 ( .A(n25766), .B(n25764), .Z(n25846) );
  OR U275 ( .A(n24520), .B(n24517), .Z(n24550) );
  NANDN U276 ( .A(n626), .B(n625), .Z(n621) );
  OR U277 ( .A(n24421), .B(n24418), .Z(n24465) );
  OR U278 ( .A(n25559), .B(n25560), .Z(n25558) );
  NANDN U279 ( .A(n565), .B(n564), .Z(n560) );
  OR U280 ( .A(n24325), .B(n24322), .Z(n24351) );
  OR U281 ( .A(n24289), .B(n24287), .Z(n24341) );
  OR U282 ( .A(n24259), .B(n24257), .Z(n24329) );
  OR U283 ( .A(n7426), .B(n7427), .Z(n7425) );
  OR U284 ( .A(n7473), .B(n7474), .Z(n7472) );
  OR U285 ( .A(n7548), .B(n7549), .Z(n7547) );
  OR U286 ( .A(n7651), .B(n7652), .Z(n7650) );
  OR U287 ( .A(n7883), .B(n7884), .Z(n7882) );
  OR U288 ( .A(n8042), .B(n8043), .Z(n8041) );
  IV U289 ( .A(n8217), .Z(n2) );
  IV U290 ( .A(B[100]), .Z(n3) );
  IV U291 ( .A(n25652), .Z(n4) );
  IV U292 ( .A(B[99]), .Z(n5) );
  IV U293 ( .A(n25747), .Z(n6) );
  IV U294 ( .A(n25755), .Z(n7) );
  IV U295 ( .A(B[97]), .Z(n8) );
  IV U296 ( .A(n25763), .Z(n9) );
  IV U297 ( .A(B[96]), .Z(n10) );
  IV U298 ( .A(n25771), .Z(n11) );
  IV U299 ( .A(B[95]), .Z(n12) );
  IV U300 ( .A(n25779), .Z(n13) );
  IV U301 ( .A(B[94]), .Z(n14) );
  IV U302 ( .A(n25787), .Z(n15) );
  IV U303 ( .A(B[93]), .Z(n16) );
  IV U304 ( .A(n25795), .Z(n17) );
  IV U305 ( .A(n25803), .Z(n18) );
  IV U306 ( .A(n25811), .Z(n19) );
  IV U307 ( .A(n25819), .Z(n20) );
  IV U308 ( .A(n25871), .Z(n21) );
  IV U309 ( .A(n25827), .Z(n22) );
  IV U310 ( .A(n1308), .Z(n23) );
  IV U311 ( .A(n24256), .Z(n24) );
  IV U312 ( .A(n24271), .Z(n25) );
  IV U313 ( .A(n24286), .Z(n26) );
  IV U314 ( .A(n24301), .Z(n27) );
  IV U315 ( .A(n24321), .Z(n28) );
  IV U316 ( .A(A[15]), .Z(n29) );
  IV U317 ( .A(A[14]), .Z(n30) );
  IV U318 ( .A(A[13]), .Z(n31) );
  IV U319 ( .A(A[12]), .Z(n32) );
  IV U320 ( .A(A[11]), .Z(n33) );
  IV U321 ( .A(A[10]), .Z(n34) );
  IV U322 ( .A(A[9]), .Z(n35) );
  IV U323 ( .A(A[8]), .Z(n36) );
  IV U324 ( .A(A[7]), .Z(n37) );
  IV U325 ( .A(A[6]), .Z(n38) );
  IV U326 ( .A(A[5]), .Z(n39) );
  IV U327 ( .A(A[4]), .Z(n40) );
  IV U328 ( .A(A[3]), .Z(n41) );
  XNOR U329 ( .A(n43), .B(n44), .Z(PRODUCT[1]) );
  AND U330 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  AND U331 ( .A(n45), .B(n46), .Z(\A2[99] ) );
  AND U332 ( .A(n47), .B(n48), .Z(\A2[98] ) );
  AND U333 ( .A(n49), .B(n50), .Z(\A2[97] ) );
  AND U334 ( .A(n51), .B(n52), .Z(\A2[96] ) );
  AND U335 ( .A(n53), .B(n54), .Z(\A2[95] ) );
  AND U336 ( .A(n55), .B(n56), .Z(\A2[94] ) );
  AND U337 ( .A(n57), .B(n58), .Z(\A2[93] ) );
  AND U338 ( .A(n59), .B(n60), .Z(\A2[92] ) );
  AND U339 ( .A(n61), .B(n62), .Z(\A2[91] ) );
  AND U340 ( .A(n63), .B(n64), .Z(\A2[90] ) );
  AND U341 ( .A(n65), .B(n66), .Z(\A2[89] ) );
  AND U342 ( .A(n67), .B(n68), .Z(\A2[88] ) );
  AND U343 ( .A(n69), .B(n70), .Z(\A2[87] ) );
  AND U344 ( .A(n71), .B(n72), .Z(\A2[86] ) );
  AND U345 ( .A(n73), .B(n74), .Z(\A2[85] ) );
  AND U346 ( .A(n75), .B(n76), .Z(\A2[84] ) );
  AND U347 ( .A(n77), .B(n78), .Z(\A2[83] ) );
  AND U348 ( .A(n79), .B(n80), .Z(\A2[82] ) );
  AND U349 ( .A(n81), .B(n82), .Z(\A2[81] ) );
  AND U350 ( .A(n83), .B(n84), .Z(\A2[80] ) );
  AND U351 ( .A(n85), .B(n86), .Z(\A2[79] ) );
  AND U352 ( .A(n87), .B(n88), .Z(\A2[78] ) );
  AND U353 ( .A(n89), .B(n90), .Z(\A2[77] ) );
  AND U354 ( .A(n91), .B(n92), .Z(\A2[76] ) );
  AND U355 ( .A(n93), .B(n94), .Z(\A2[75] ) );
  AND U356 ( .A(n95), .B(n96), .Z(\A2[74] ) );
  AND U357 ( .A(n97), .B(n98), .Z(\A2[73] ) );
  AND U358 ( .A(n99), .B(n100), .Z(\A2[72] ) );
  AND U359 ( .A(n101), .B(n102), .Z(\A2[71] ) );
  AND U360 ( .A(n103), .B(n104), .Z(\A2[70] ) );
  AND U361 ( .A(n105), .B(n106), .Z(\A2[69] ) );
  AND U362 ( .A(n107), .B(n108), .Z(\A2[68] ) );
  AND U363 ( .A(n109), .B(n110), .Z(\A2[67] ) );
  AND U364 ( .A(n111), .B(n112), .Z(\A2[66] ) );
  AND U365 ( .A(n113), .B(n114), .Z(\A2[65] ) );
  AND U366 ( .A(n115), .B(n116), .Z(\A2[64] ) );
  AND U367 ( .A(n117), .B(n118), .Z(\A2[63] ) );
  AND U368 ( .A(n119), .B(n120), .Z(\A2[62] ) );
  AND U369 ( .A(n121), .B(n122), .Z(\A2[61] ) );
  AND U370 ( .A(n123), .B(n124), .Z(\A2[60] ) );
  AND U371 ( .A(n125), .B(n126), .Z(\A2[59] ) );
  AND U372 ( .A(n127), .B(n128), .Z(\A2[58] ) );
  AND U373 ( .A(n129), .B(n130), .Z(\A2[57] ) );
  AND U374 ( .A(n131), .B(n132), .Z(\A2[56] ) );
  AND U375 ( .A(n133), .B(n134), .Z(\A2[55] ) );
  AND U376 ( .A(n135), .B(n136), .Z(\A2[54] ) );
  AND U377 ( .A(n137), .B(n138), .Z(\A2[53] ) );
  AND U378 ( .A(n139), .B(n140), .Z(\A2[52] ) );
  AND U379 ( .A(n141), .B(n142), .Z(\A2[51] ) );
  AND U380 ( .A(n143), .B(n144), .Z(\A2[50] ) );
  AND U381 ( .A(n145), .B(n146), .Z(\A2[49] ) );
  AND U382 ( .A(n147), .B(n148), .Z(\A2[48] ) );
  AND U383 ( .A(n149), .B(n150), .Z(\A2[47] ) );
  AND U384 ( .A(n151), .B(n152), .Z(\A2[46] ) );
  AND U385 ( .A(n153), .B(n154), .Z(\A2[45] ) );
  AND U386 ( .A(n155), .B(n156), .Z(\A2[44] ) );
  AND U387 ( .A(n157), .B(n158), .Z(\A2[43] ) );
  AND U388 ( .A(n159), .B(n160), .Z(\A2[42] ) );
  AND U389 ( .A(n161), .B(n162), .Z(\A2[41] ) );
  AND U390 ( .A(n163), .B(n164), .Z(\A2[40] ) );
  AND U391 ( .A(n165), .B(n166), .Z(\A2[39] ) );
  AND U392 ( .A(n167), .B(n168), .Z(\A2[38] ) );
  AND U393 ( .A(n169), .B(n170), .Z(\A2[37] ) );
  AND U394 ( .A(n171), .B(n172), .Z(\A2[36] ) );
  AND U395 ( .A(n173), .B(n174), .Z(\A2[35] ) );
  AND U396 ( .A(n175), .B(n176), .Z(\A2[34] ) );
  AND U397 ( .A(n177), .B(n178), .Z(\A2[33] ) );
  AND U398 ( .A(n179), .B(n180), .Z(\A2[32] ) );
  AND U399 ( .A(n181), .B(n182), .Z(\A2[31] ) );
  AND U400 ( .A(n183), .B(n184), .Z(\A2[30] ) );
  AND U401 ( .A(n185), .B(n186), .Z(\A2[29] ) );
  AND U402 ( .A(n187), .B(n188), .Z(\A2[28] ) );
  AND U403 ( .A(n189), .B(n190), .Z(\A2[27] ) );
  AND U404 ( .A(n191), .B(n192), .Z(\A2[26] ) );
  AND U405 ( .A(n193), .B(A[15]), .Z(\A2[269] ) );
  AND U406 ( .A(n194), .B(n195), .Z(\A2[268] ) );
  AND U407 ( .A(n196), .B(n197), .Z(\A2[267] ) );
  AND U408 ( .A(n198), .B(n199), .Z(\A2[266] ) );
  AND U409 ( .A(n200), .B(n201), .Z(\A2[265] ) );
  AND U410 ( .A(n202), .B(n203), .Z(\A2[264] ) );
  AND U411 ( .A(n204), .B(n205), .Z(\A2[263] ) );
  AND U412 ( .A(n206), .B(n207), .Z(\A2[262] ) );
  AND U413 ( .A(n208), .B(n209), .Z(\A2[261] ) );
  AND U414 ( .A(n210), .B(n211), .Z(\A2[260] ) );
  AND U415 ( .A(n212), .B(n213), .Z(\A2[25] ) );
  AND U416 ( .A(n214), .B(n215), .Z(\A2[259] ) );
  AND U417 ( .A(n216), .B(n217), .Z(\A2[258] ) );
  AND U418 ( .A(n218), .B(n219), .Z(\A2[257] ) );
  AND U419 ( .A(n220), .B(n221), .Z(\A2[256] ) );
  AND U420 ( .A(n222), .B(n223), .Z(\A2[255] ) );
  AND U421 ( .A(n224), .B(n225), .Z(\A2[254] ) );
  AND U422 ( .A(n226), .B(n227), .Z(\A2[253] ) );
  AND U423 ( .A(n228), .B(n229), .Z(\A2[252] ) );
  AND U424 ( .A(n230), .B(n231), .Z(\A2[251] ) );
  AND U425 ( .A(n232), .B(n233), .Z(\A2[250] ) );
  AND U426 ( .A(n234), .B(n235), .Z(\A2[24] ) );
  AND U427 ( .A(n236), .B(n237), .Z(\A2[249] ) );
  AND U428 ( .A(n238), .B(n239), .Z(\A2[248] ) );
  AND U429 ( .A(n240), .B(n241), .Z(\A2[247] ) );
  AND U430 ( .A(n242), .B(n243), .Z(\A2[246] ) );
  AND U431 ( .A(n244), .B(n245), .Z(\A2[245] ) );
  AND U432 ( .A(n246), .B(n247), .Z(\A2[244] ) );
  AND U433 ( .A(n248), .B(n249), .Z(\A2[243] ) );
  AND U434 ( .A(n250), .B(n251), .Z(\A2[242] ) );
  AND U435 ( .A(n252), .B(n253), .Z(\A2[241] ) );
  AND U436 ( .A(n254), .B(n255), .Z(\A2[240] ) );
  AND U437 ( .A(n256), .B(n257), .Z(\A2[23] ) );
  AND U438 ( .A(n258), .B(n259), .Z(\A2[239] ) );
  AND U439 ( .A(n260), .B(n261), .Z(\A2[238] ) );
  AND U440 ( .A(n262), .B(n263), .Z(\A2[237] ) );
  AND U441 ( .A(n264), .B(n265), .Z(\A2[236] ) );
  AND U442 ( .A(n266), .B(n267), .Z(\A2[235] ) );
  AND U443 ( .A(n268), .B(n269), .Z(\A2[234] ) );
  AND U444 ( .A(n270), .B(n271), .Z(\A2[233] ) );
  AND U445 ( .A(n272), .B(n273), .Z(\A2[232] ) );
  AND U446 ( .A(n274), .B(n275), .Z(\A2[231] ) );
  AND U447 ( .A(n276), .B(n277), .Z(\A2[230] ) );
  AND U448 ( .A(n278), .B(n279), .Z(\A2[22] ) );
  AND U449 ( .A(n280), .B(n281), .Z(\A2[229] ) );
  AND U450 ( .A(n282), .B(n283), .Z(\A2[228] ) );
  AND U451 ( .A(n284), .B(n285), .Z(\A2[227] ) );
  AND U452 ( .A(n286), .B(n287), .Z(\A2[226] ) );
  AND U453 ( .A(n288), .B(n289), .Z(\A2[225] ) );
  AND U454 ( .A(n290), .B(n291), .Z(\A2[224] ) );
  AND U455 ( .A(n292), .B(n293), .Z(\A2[223] ) );
  AND U456 ( .A(n294), .B(n295), .Z(\A2[222] ) );
  AND U457 ( .A(n296), .B(n297), .Z(\A2[221] ) );
  AND U458 ( .A(n298), .B(n299), .Z(\A2[220] ) );
  AND U459 ( .A(n300), .B(n301), .Z(\A2[21] ) );
  AND U460 ( .A(n302), .B(n303), .Z(\A2[219] ) );
  AND U461 ( .A(n304), .B(n305), .Z(\A2[218] ) );
  AND U462 ( .A(n306), .B(n307), .Z(\A2[217] ) );
  AND U463 ( .A(n308), .B(n309), .Z(\A2[216] ) );
  AND U464 ( .A(n310), .B(n311), .Z(\A2[215] ) );
  AND U465 ( .A(n312), .B(n313), .Z(\A2[214] ) );
  AND U466 ( .A(n314), .B(n315), .Z(\A2[213] ) );
  AND U467 ( .A(n316), .B(n317), .Z(\A2[212] ) );
  AND U468 ( .A(n318), .B(n319), .Z(\A2[211] ) );
  AND U469 ( .A(n320), .B(n321), .Z(\A2[210] ) );
  AND U470 ( .A(n322), .B(n323), .Z(\A2[20] ) );
  AND U471 ( .A(n324), .B(n325), .Z(\A2[209] ) );
  AND U472 ( .A(n326), .B(n327), .Z(\A2[208] ) );
  AND U473 ( .A(n328), .B(n329), .Z(\A2[207] ) );
  AND U474 ( .A(n330), .B(n331), .Z(\A2[206] ) );
  AND U475 ( .A(n332), .B(n333), .Z(\A2[205] ) );
  AND U476 ( .A(n334), .B(n335), .Z(\A2[204] ) );
  AND U477 ( .A(n336), .B(n337), .Z(\A2[203] ) );
  AND U478 ( .A(n338), .B(n339), .Z(\A2[202] ) );
  AND U479 ( .A(n340), .B(n341), .Z(\A2[201] ) );
  AND U480 ( .A(n342), .B(n343), .Z(\A2[200] ) );
  AND U481 ( .A(n344), .B(n345), .Z(\A2[19] ) );
  AND U482 ( .A(n346), .B(n347), .Z(\A2[199] ) );
  AND U483 ( .A(n348), .B(n349), .Z(\A2[198] ) );
  AND U484 ( .A(n350), .B(n351), .Z(\A2[197] ) );
  AND U485 ( .A(n352), .B(n353), .Z(\A2[196] ) );
  AND U486 ( .A(n354), .B(n355), .Z(\A2[195] ) );
  AND U487 ( .A(n356), .B(n357), .Z(\A2[194] ) );
  AND U488 ( .A(n358), .B(n359), .Z(\A2[193] ) );
  AND U489 ( .A(n360), .B(n361), .Z(\A2[192] ) );
  AND U490 ( .A(n362), .B(n363), .Z(\A2[191] ) );
  AND U491 ( .A(n364), .B(n365), .Z(\A2[190] ) );
  AND U492 ( .A(n366), .B(n367), .Z(\A2[18] ) );
  AND U493 ( .A(n368), .B(n369), .Z(\A2[189] ) );
  AND U494 ( .A(n370), .B(n371), .Z(\A2[188] ) );
  AND U495 ( .A(n372), .B(n373), .Z(\A2[187] ) );
  AND U496 ( .A(n374), .B(n375), .Z(\A2[186] ) );
  AND U497 ( .A(n376), .B(n377), .Z(\A2[185] ) );
  AND U498 ( .A(n378), .B(n379), .Z(\A2[184] ) );
  AND U499 ( .A(n380), .B(n381), .Z(\A2[183] ) );
  AND U500 ( .A(n382), .B(n383), .Z(\A2[182] ) );
  AND U501 ( .A(n384), .B(n385), .Z(\A2[181] ) );
  AND U502 ( .A(n386), .B(n387), .Z(\A2[180] ) );
  AND U503 ( .A(n388), .B(n389), .Z(\A2[17] ) );
  AND U504 ( .A(n390), .B(n391), .Z(\A2[179] ) );
  AND U505 ( .A(n392), .B(n393), .Z(\A2[178] ) );
  AND U506 ( .A(n394), .B(n395), .Z(\A2[177] ) );
  AND U507 ( .A(n396), .B(n397), .Z(\A2[176] ) );
  AND U508 ( .A(n398), .B(n399), .Z(\A2[175] ) );
  AND U509 ( .A(n400), .B(n401), .Z(\A2[174] ) );
  AND U510 ( .A(n402), .B(n403), .Z(\A2[173] ) );
  AND U511 ( .A(n404), .B(n405), .Z(\A2[172] ) );
  AND U512 ( .A(n406), .B(n407), .Z(\A2[171] ) );
  AND U513 ( .A(n408), .B(n409), .Z(\A2[170] ) );
  AND U514 ( .A(n410), .B(n411), .Z(\A2[16] ) );
  AND U515 ( .A(n412), .B(n413), .Z(\A2[169] ) );
  AND U516 ( .A(n414), .B(n415), .Z(\A2[168] ) );
  AND U517 ( .A(n416), .B(n417), .Z(\A2[167] ) );
  AND U518 ( .A(n418), .B(n419), .Z(\A2[166] ) );
  AND U519 ( .A(n420), .B(n421), .Z(\A2[165] ) );
  AND U520 ( .A(n422), .B(n423), .Z(\A2[164] ) );
  AND U521 ( .A(n424), .B(n425), .Z(\A2[163] ) );
  AND U522 ( .A(n426), .B(n427), .Z(\A2[162] ) );
  AND U523 ( .A(n428), .B(n429), .Z(\A2[161] ) );
  AND U524 ( .A(n430), .B(n431), .Z(\A2[160] ) );
  AND U525 ( .A(n432), .B(n433), .Z(\A2[15] ) );
  AND U526 ( .A(n434), .B(n435), .Z(\A2[159] ) );
  AND U527 ( .A(n436), .B(n437), .Z(\A2[158] ) );
  AND U528 ( .A(n438), .B(n439), .Z(\A2[157] ) );
  AND U529 ( .A(n440), .B(n441), .Z(\A2[156] ) );
  AND U530 ( .A(n442), .B(n443), .Z(\A2[155] ) );
  AND U531 ( .A(n444), .B(n445), .Z(\A2[154] ) );
  AND U532 ( .A(n446), .B(n447), .Z(\A2[153] ) );
  AND U533 ( .A(n448), .B(n449), .Z(\A2[152] ) );
  AND U534 ( .A(n450), .B(n451), .Z(\A2[151] ) );
  AND U535 ( .A(n452), .B(n453), .Z(\A2[150] ) );
  AND U536 ( .A(n454), .B(n455), .Z(\A2[149] ) );
  AND U537 ( .A(n456), .B(n457), .Z(\A2[148] ) );
  AND U538 ( .A(n458), .B(n459), .Z(\A2[147] ) );
  AND U539 ( .A(n460), .B(n461), .Z(\A2[146] ) );
  AND U540 ( .A(n462), .B(n463), .Z(\A2[145] ) );
  AND U541 ( .A(n464), .B(n465), .Z(\A2[144] ) );
  AND U542 ( .A(n466), .B(n467), .Z(\A2[143] ) );
  AND U543 ( .A(n468), .B(n469), .Z(\A2[142] ) );
  AND U544 ( .A(n470), .B(n471), .Z(\A2[141] ) );
  AND U545 ( .A(n472), .B(n473), .Z(\A2[140] ) );
  AND U546 ( .A(n474), .B(n475), .Z(\A2[139] ) );
  AND U547 ( .A(n476), .B(n477), .Z(\A2[138] ) );
  AND U548 ( .A(n478), .B(n479), .Z(\A2[137] ) );
  AND U549 ( .A(n480), .B(n481), .Z(\A2[136] ) );
  AND U550 ( .A(n482), .B(n483), .Z(\A2[135] ) );
  AND U551 ( .A(n484), .B(n485), .Z(\A2[134] ) );
  AND U552 ( .A(n486), .B(n487), .Z(\A2[133] ) );
  AND U553 ( .A(n488), .B(n489), .Z(\A2[132] ) );
  AND U554 ( .A(n490), .B(n491), .Z(\A2[131] ) );
  AND U555 ( .A(n492), .B(n493), .Z(\A2[130] ) );
  AND U556 ( .A(n494), .B(n495), .Z(\A2[129] ) );
  AND U557 ( .A(n496), .B(n497), .Z(\A2[128] ) );
  AND U558 ( .A(n498), .B(n499), .Z(\A2[127] ) );
  AND U559 ( .A(n500), .B(n501), .Z(\A2[126] ) );
  AND U560 ( .A(n502), .B(n503), .Z(\A2[125] ) );
  AND U561 ( .A(n504), .B(n505), .Z(\A2[124] ) );
  AND U562 ( .A(n506), .B(n507), .Z(\A2[123] ) );
  AND U563 ( .A(n508), .B(n509), .Z(\A2[122] ) );
  AND U564 ( .A(n510), .B(n511), .Z(\A2[121] ) );
  AND U565 ( .A(n512), .B(n513), .Z(\A2[120] ) );
  AND U566 ( .A(n514), .B(n515), .Z(\A2[119] ) );
  AND U567 ( .A(n516), .B(n517), .Z(\A2[118] ) );
  AND U568 ( .A(n518), .B(n519), .Z(\A2[117] ) );
  AND U569 ( .A(n520), .B(n521), .Z(\A2[116] ) );
  AND U570 ( .A(n522), .B(n523), .Z(\A2[115] ) );
  AND U571 ( .A(n524), .B(n525), .Z(\A2[114] ) );
  AND U572 ( .A(n526), .B(n527), .Z(\A2[113] ) );
  AND U573 ( .A(n528), .B(n529), .Z(\A2[112] ) );
  AND U574 ( .A(n530), .B(n531), .Z(\A2[111] ) );
  AND U575 ( .A(n532), .B(n533), .Z(\A2[110] ) );
  AND U576 ( .A(n534), .B(n535), .Z(\A2[109] ) );
  AND U577 ( .A(n536), .B(n537), .Z(\A2[108] ) );
  AND U578 ( .A(n538), .B(n539), .Z(\A2[107] ) );
  AND U579 ( .A(n540), .B(n541), .Z(\A2[106] ) );
  AND U580 ( .A(n542), .B(n543), .Z(\A2[105] ) );
  AND U581 ( .A(n544), .B(n545), .Z(\A2[104] ) );
  AND U582 ( .A(n546), .B(n547), .Z(\A2[103] ) );
  AND U583 ( .A(n548), .B(n549), .Z(\A2[102] ) );
  AND U584 ( .A(n550), .B(n551), .Z(\A2[101] ) );
  AND U585 ( .A(n552), .B(n553), .Z(\A2[100] ) );
  XOR U586 ( .A(n554), .B(n555), .Z(\A1[9] ) );
  XNOR U587 ( .A(n556), .B(n24), .Z(n555) );
  XOR U588 ( .A(n553), .B(n552), .Z(\A1[99] ) );
  XOR U589 ( .A(n557), .B(n558), .Z(n552) );
  XNOR U590 ( .A(n559), .B(n4), .Z(n558) );
  NAND U591 ( .A(n560), .B(n561), .Z(n553) );
  NANDN U592 ( .A(n562), .B(n563), .Z(n561) );
  NANDN U593 ( .A(n564), .B(n565), .Z(n563) );
  XOR U594 ( .A(n46), .B(n45), .Z(\A1[98] ) );
  XNOR U595 ( .A(n562), .B(n566), .Z(n45) );
  XNOR U596 ( .A(n564), .B(n565), .Z(n566) );
  AND U597 ( .A(n567), .B(n568), .Z(n565) );
  NAND U598 ( .A(n569), .B(n570), .Z(n568) );
  NANDN U599 ( .A(n571), .B(n572), .Z(n569) );
  ANDN U600 ( .B(B[85]), .A(n29), .Z(n564) );
  XOR U601 ( .A(n573), .B(n574), .Z(n562) );
  XOR U602 ( .A(n575), .B(n576), .Z(n574) );
  NAND U603 ( .A(n577), .B(n578), .Z(n46) );
  NANDN U604 ( .A(n579), .B(n580), .Z(n578) );
  OR U605 ( .A(n581), .B(n582), .Z(n580) );
  NAND U606 ( .A(n582), .B(n581), .Z(n577) );
  XOR U607 ( .A(n48), .B(n47), .Z(\A1[97] ) );
  XOR U608 ( .A(n582), .B(n583), .Z(n47) );
  XNOR U609 ( .A(n581), .B(n579), .Z(n583) );
  AND U610 ( .A(n584), .B(n585), .Z(n579) );
  NANDN U611 ( .A(n586), .B(n587), .Z(n585) );
  NANDN U612 ( .A(n588), .B(n589), .Z(n587) );
  NANDN U613 ( .A(n589), .B(n588), .Z(n584) );
  ANDN U614 ( .B(B[84]), .A(n29), .Z(n581) );
  XOR U615 ( .A(n570), .B(n590), .Z(n582) );
  XNOR U616 ( .A(n571), .B(n572), .Z(n590) );
  AND U617 ( .A(n591), .B(n592), .Z(n572) );
  NANDN U618 ( .A(n593), .B(n594), .Z(n592) );
  NANDN U619 ( .A(n595), .B(n596), .Z(n594) );
  ANDN U620 ( .B(B[85]), .A(n30), .Z(n571) );
  XOR U621 ( .A(n597), .B(n598), .Z(n570) );
  XNOR U622 ( .A(n599), .B(n6), .Z(n598) );
  NAND U623 ( .A(n600), .B(n601), .Z(n48) );
  NANDN U624 ( .A(n602), .B(n603), .Z(n601) );
  OR U625 ( .A(n604), .B(n605), .Z(n603) );
  NAND U626 ( .A(n605), .B(n604), .Z(n600) );
  XOR U627 ( .A(n50), .B(n49), .Z(\A1[96] ) );
  XOR U628 ( .A(n605), .B(n606), .Z(n49) );
  XNOR U629 ( .A(n604), .B(n602), .Z(n606) );
  AND U630 ( .A(n607), .B(n608), .Z(n602) );
  NANDN U631 ( .A(n609), .B(n610), .Z(n608) );
  NANDN U632 ( .A(n611), .B(n612), .Z(n610) );
  NANDN U633 ( .A(n612), .B(n611), .Z(n607) );
  ANDN U634 ( .B(B[83]), .A(n29), .Z(n604) );
  XNOR U635 ( .A(n589), .B(n613), .Z(n605) );
  XNOR U636 ( .A(n588), .B(n586), .Z(n613) );
  AND U637 ( .A(n614), .B(n615), .Z(n586) );
  NANDN U638 ( .A(n616), .B(n617), .Z(n615) );
  OR U639 ( .A(n618), .B(n619), .Z(n617) );
  NAND U640 ( .A(n619), .B(n618), .Z(n614) );
  ANDN U641 ( .B(B[84]), .A(n30), .Z(n588) );
  XOR U642 ( .A(n593), .B(n620), .Z(n589) );
  XNOR U643 ( .A(n595), .B(n596), .Z(n620) );
  AND U644 ( .A(n621), .B(n622), .Z(n596) );
  NAND U645 ( .A(n623), .B(n624), .Z(n622) );
  NANDN U646 ( .A(n625), .B(n626), .Z(n623) );
  ANDN U647 ( .B(B[85]), .A(n31), .Z(n595) );
  XNOR U648 ( .A(n627), .B(n628), .Z(n593) );
  XNOR U649 ( .A(n629), .B(n7), .Z(n628) );
  NAND U650 ( .A(n630), .B(n631), .Z(n50) );
  NANDN U651 ( .A(n632), .B(n633), .Z(n631) );
  OR U652 ( .A(n634), .B(n635), .Z(n633) );
  NAND U653 ( .A(n635), .B(n634), .Z(n630) );
  XOR U654 ( .A(n52), .B(n51), .Z(\A1[95] ) );
  XOR U655 ( .A(n635), .B(n636), .Z(n51) );
  XNOR U656 ( .A(n634), .B(n632), .Z(n636) );
  AND U657 ( .A(n637), .B(n638), .Z(n632) );
  NANDN U658 ( .A(n639), .B(n640), .Z(n638) );
  NANDN U659 ( .A(n641), .B(n642), .Z(n640) );
  NANDN U660 ( .A(n642), .B(n641), .Z(n637) );
  ANDN U661 ( .B(B[82]), .A(n29), .Z(n634) );
  XNOR U662 ( .A(n612), .B(n643), .Z(n635) );
  XNOR U663 ( .A(n611), .B(n609), .Z(n643) );
  AND U664 ( .A(n644), .B(n645), .Z(n609) );
  NANDN U665 ( .A(n646), .B(n647), .Z(n645) );
  OR U666 ( .A(n648), .B(n649), .Z(n647) );
  NAND U667 ( .A(n649), .B(n648), .Z(n644) );
  ANDN U668 ( .B(B[83]), .A(n30), .Z(n611) );
  XNOR U669 ( .A(n619), .B(n650), .Z(n612) );
  XNOR U670 ( .A(n618), .B(n616), .Z(n650) );
  AND U671 ( .A(n651), .B(n652), .Z(n616) );
  NANDN U672 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U673 ( .A(n655), .B(n656), .Z(n654) );
  NANDN U674 ( .A(n656), .B(n655), .Z(n651) );
  ANDN U675 ( .B(B[84]), .A(n31), .Z(n618) );
  XOR U676 ( .A(n624), .B(n657), .Z(n619) );
  XNOR U677 ( .A(n625), .B(n626), .Z(n657) );
  AND U678 ( .A(n658), .B(n659), .Z(n626) );
  NANDN U679 ( .A(n660), .B(n661), .Z(n659) );
  NANDN U680 ( .A(n662), .B(n663), .Z(n661) );
  ANDN U681 ( .B(B[85]), .A(n32), .Z(n625) );
  XOR U682 ( .A(n664), .B(n665), .Z(n624) );
  XNOR U683 ( .A(n666), .B(n9), .Z(n665) );
  NAND U684 ( .A(n667), .B(n668), .Z(n52) );
  NANDN U685 ( .A(n669), .B(n670), .Z(n668) );
  OR U686 ( .A(n671), .B(n672), .Z(n670) );
  NAND U687 ( .A(n672), .B(n671), .Z(n667) );
  XOR U688 ( .A(n54), .B(n53), .Z(\A1[94] ) );
  XOR U689 ( .A(n672), .B(n673), .Z(n53) );
  XNOR U690 ( .A(n671), .B(n669), .Z(n673) );
  AND U691 ( .A(n674), .B(n675), .Z(n669) );
  NANDN U692 ( .A(n676), .B(n677), .Z(n675) );
  NANDN U693 ( .A(n678), .B(n679), .Z(n677) );
  NANDN U694 ( .A(n679), .B(n678), .Z(n674) );
  ANDN U695 ( .B(B[81]), .A(n29), .Z(n671) );
  XNOR U696 ( .A(n642), .B(n680), .Z(n672) );
  XNOR U697 ( .A(n641), .B(n639), .Z(n680) );
  AND U698 ( .A(n681), .B(n682), .Z(n639) );
  NANDN U699 ( .A(n683), .B(n684), .Z(n682) );
  OR U700 ( .A(n685), .B(n686), .Z(n684) );
  NAND U701 ( .A(n686), .B(n685), .Z(n681) );
  ANDN U702 ( .B(B[82]), .A(n30), .Z(n641) );
  XNOR U703 ( .A(n649), .B(n687), .Z(n642) );
  XNOR U704 ( .A(n648), .B(n646), .Z(n687) );
  AND U705 ( .A(n688), .B(n689), .Z(n646) );
  NANDN U706 ( .A(n690), .B(n691), .Z(n689) );
  NANDN U707 ( .A(n692), .B(n693), .Z(n691) );
  NANDN U708 ( .A(n693), .B(n692), .Z(n688) );
  ANDN U709 ( .B(B[83]), .A(n31), .Z(n648) );
  XNOR U710 ( .A(n656), .B(n694), .Z(n649) );
  XNOR U711 ( .A(n655), .B(n653), .Z(n694) );
  AND U712 ( .A(n695), .B(n696), .Z(n653) );
  NANDN U713 ( .A(n697), .B(n698), .Z(n696) );
  OR U714 ( .A(n699), .B(n700), .Z(n698) );
  NAND U715 ( .A(n700), .B(n699), .Z(n695) );
  ANDN U716 ( .B(B[84]), .A(n32), .Z(n655) );
  XOR U717 ( .A(n660), .B(n701), .Z(n656) );
  XNOR U718 ( .A(n662), .B(n663), .Z(n701) );
  AND U719 ( .A(n702), .B(n703), .Z(n663) );
  NAND U720 ( .A(n704), .B(n705), .Z(n703) );
  NANDN U721 ( .A(n706), .B(n707), .Z(n704) );
  ANDN U722 ( .B(B[85]), .A(n33), .Z(n662) );
  XNOR U723 ( .A(n708), .B(n709), .Z(n660) );
  XNOR U724 ( .A(n710), .B(n11), .Z(n709) );
  NAND U725 ( .A(n711), .B(n712), .Z(n54) );
  NANDN U726 ( .A(n713), .B(n714), .Z(n712) );
  OR U727 ( .A(n715), .B(n716), .Z(n714) );
  NAND U728 ( .A(n716), .B(n715), .Z(n711) );
  XOR U729 ( .A(n56), .B(n55), .Z(\A1[93] ) );
  XOR U730 ( .A(n716), .B(n717), .Z(n55) );
  XNOR U731 ( .A(n715), .B(n713), .Z(n717) );
  AND U732 ( .A(n718), .B(n719), .Z(n713) );
  NANDN U733 ( .A(n720), .B(n721), .Z(n719) );
  NANDN U734 ( .A(n722), .B(n723), .Z(n721) );
  NANDN U735 ( .A(n723), .B(n722), .Z(n718) );
  ANDN U736 ( .B(B[80]), .A(n29), .Z(n715) );
  XNOR U737 ( .A(n679), .B(n724), .Z(n716) );
  XNOR U738 ( .A(n678), .B(n676), .Z(n724) );
  AND U739 ( .A(n725), .B(n726), .Z(n676) );
  NANDN U740 ( .A(n727), .B(n728), .Z(n726) );
  OR U741 ( .A(n729), .B(n730), .Z(n728) );
  NAND U742 ( .A(n730), .B(n729), .Z(n725) );
  ANDN U743 ( .B(B[81]), .A(n30), .Z(n678) );
  XNOR U744 ( .A(n686), .B(n731), .Z(n679) );
  XNOR U745 ( .A(n685), .B(n683), .Z(n731) );
  AND U746 ( .A(n732), .B(n733), .Z(n683) );
  NANDN U747 ( .A(n734), .B(n735), .Z(n733) );
  NANDN U748 ( .A(n736), .B(n737), .Z(n735) );
  NANDN U749 ( .A(n737), .B(n736), .Z(n732) );
  ANDN U750 ( .B(B[82]), .A(n31), .Z(n685) );
  XNOR U751 ( .A(n693), .B(n738), .Z(n686) );
  XNOR U752 ( .A(n692), .B(n690), .Z(n738) );
  AND U753 ( .A(n739), .B(n740), .Z(n690) );
  NANDN U754 ( .A(n741), .B(n742), .Z(n740) );
  OR U755 ( .A(n743), .B(n744), .Z(n742) );
  NAND U756 ( .A(n744), .B(n743), .Z(n739) );
  ANDN U757 ( .B(B[83]), .A(n32), .Z(n692) );
  XNOR U758 ( .A(n700), .B(n745), .Z(n693) );
  XNOR U759 ( .A(n699), .B(n697), .Z(n745) );
  AND U760 ( .A(n746), .B(n747), .Z(n697) );
  NANDN U761 ( .A(n748), .B(n749), .Z(n747) );
  NANDN U762 ( .A(n750), .B(n751), .Z(n749) );
  NANDN U763 ( .A(n751), .B(n750), .Z(n746) );
  ANDN U764 ( .B(B[84]), .A(n33), .Z(n699) );
  XOR U765 ( .A(n705), .B(n752), .Z(n700) );
  XNOR U766 ( .A(n706), .B(n707), .Z(n752) );
  AND U767 ( .A(n753), .B(n754), .Z(n707) );
  NANDN U768 ( .A(n755), .B(n756), .Z(n754) );
  NANDN U769 ( .A(n757), .B(n758), .Z(n756) );
  ANDN U770 ( .B(B[85]), .A(n34), .Z(n706) );
  XOR U771 ( .A(n759), .B(n760), .Z(n705) );
  XNOR U772 ( .A(n761), .B(n13), .Z(n760) );
  NAND U773 ( .A(n762), .B(n763), .Z(n56) );
  NANDN U774 ( .A(n764), .B(n765), .Z(n763) );
  OR U775 ( .A(n766), .B(n767), .Z(n765) );
  NAND U776 ( .A(n767), .B(n766), .Z(n762) );
  XOR U777 ( .A(n58), .B(n57), .Z(\A1[92] ) );
  XOR U778 ( .A(n767), .B(n768), .Z(n57) );
  XNOR U779 ( .A(n766), .B(n764), .Z(n768) );
  AND U780 ( .A(n769), .B(n770), .Z(n764) );
  NANDN U781 ( .A(n771), .B(n772), .Z(n770) );
  NANDN U782 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U783 ( .A(n774), .B(n773), .Z(n769) );
  ANDN U784 ( .B(B[79]), .A(n29), .Z(n766) );
  XNOR U785 ( .A(n723), .B(n775), .Z(n767) );
  XNOR U786 ( .A(n722), .B(n720), .Z(n775) );
  AND U787 ( .A(n776), .B(n777), .Z(n720) );
  NANDN U788 ( .A(n778), .B(n779), .Z(n777) );
  OR U789 ( .A(n780), .B(n781), .Z(n779) );
  NAND U790 ( .A(n781), .B(n780), .Z(n776) );
  ANDN U791 ( .B(B[80]), .A(n30), .Z(n722) );
  XNOR U792 ( .A(n730), .B(n782), .Z(n723) );
  XNOR U793 ( .A(n729), .B(n727), .Z(n782) );
  AND U794 ( .A(n783), .B(n784), .Z(n727) );
  NANDN U795 ( .A(n785), .B(n786), .Z(n784) );
  NANDN U796 ( .A(n787), .B(n788), .Z(n786) );
  NANDN U797 ( .A(n788), .B(n787), .Z(n783) );
  ANDN U798 ( .B(B[81]), .A(n31), .Z(n729) );
  XNOR U799 ( .A(n737), .B(n789), .Z(n730) );
  XNOR U800 ( .A(n736), .B(n734), .Z(n789) );
  AND U801 ( .A(n790), .B(n791), .Z(n734) );
  NANDN U802 ( .A(n792), .B(n793), .Z(n791) );
  OR U803 ( .A(n794), .B(n795), .Z(n793) );
  NAND U804 ( .A(n795), .B(n794), .Z(n790) );
  ANDN U805 ( .B(B[82]), .A(n32), .Z(n736) );
  XNOR U806 ( .A(n744), .B(n796), .Z(n737) );
  XNOR U807 ( .A(n743), .B(n741), .Z(n796) );
  AND U808 ( .A(n797), .B(n798), .Z(n741) );
  NANDN U809 ( .A(n799), .B(n800), .Z(n798) );
  NANDN U810 ( .A(n801), .B(n802), .Z(n800) );
  NANDN U811 ( .A(n802), .B(n801), .Z(n797) );
  ANDN U812 ( .B(B[83]), .A(n33), .Z(n743) );
  XNOR U813 ( .A(n751), .B(n803), .Z(n744) );
  XNOR U814 ( .A(n750), .B(n748), .Z(n803) );
  AND U815 ( .A(n804), .B(n805), .Z(n748) );
  NANDN U816 ( .A(n806), .B(n807), .Z(n805) );
  OR U817 ( .A(n808), .B(n809), .Z(n807) );
  NAND U818 ( .A(n809), .B(n808), .Z(n804) );
  ANDN U819 ( .B(B[84]), .A(n34), .Z(n750) );
  XOR U820 ( .A(n755), .B(n810), .Z(n751) );
  XNOR U821 ( .A(n757), .B(n758), .Z(n810) );
  AND U822 ( .A(n811), .B(n812), .Z(n758) );
  NAND U823 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U824 ( .A(n815), .B(n816), .Z(n813) );
  ANDN U825 ( .B(B[85]), .A(n35), .Z(n757) );
  XNOR U826 ( .A(n817), .B(n818), .Z(n755) );
  XNOR U827 ( .A(n819), .B(n15), .Z(n818) );
  NAND U828 ( .A(n820), .B(n821), .Z(n58) );
  NANDN U829 ( .A(n822), .B(n823), .Z(n821) );
  OR U830 ( .A(n824), .B(n825), .Z(n823) );
  NAND U831 ( .A(n825), .B(n824), .Z(n820) );
  XOR U832 ( .A(n60), .B(n59), .Z(\A1[91] ) );
  XOR U833 ( .A(n825), .B(n826), .Z(n59) );
  XNOR U834 ( .A(n824), .B(n822), .Z(n826) );
  AND U835 ( .A(n827), .B(n828), .Z(n822) );
  NANDN U836 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U837 ( .A(n831), .B(n832), .Z(n830) );
  NANDN U838 ( .A(n832), .B(n831), .Z(n827) );
  ANDN U839 ( .B(B[78]), .A(n29), .Z(n824) );
  XNOR U840 ( .A(n774), .B(n833), .Z(n825) );
  XNOR U841 ( .A(n773), .B(n771), .Z(n833) );
  AND U842 ( .A(n834), .B(n835), .Z(n771) );
  NANDN U843 ( .A(n836), .B(n837), .Z(n835) );
  OR U844 ( .A(n838), .B(n839), .Z(n837) );
  NAND U845 ( .A(n839), .B(n838), .Z(n834) );
  ANDN U846 ( .B(B[79]), .A(n30), .Z(n773) );
  XNOR U847 ( .A(n781), .B(n840), .Z(n774) );
  XNOR U848 ( .A(n780), .B(n778), .Z(n840) );
  AND U849 ( .A(n841), .B(n842), .Z(n778) );
  NANDN U850 ( .A(n843), .B(n844), .Z(n842) );
  NANDN U851 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U852 ( .A(n846), .B(n845), .Z(n841) );
  ANDN U853 ( .B(B[80]), .A(n31), .Z(n780) );
  XNOR U854 ( .A(n788), .B(n847), .Z(n781) );
  XNOR U855 ( .A(n787), .B(n785), .Z(n847) );
  AND U856 ( .A(n848), .B(n849), .Z(n785) );
  NANDN U857 ( .A(n850), .B(n851), .Z(n849) );
  OR U858 ( .A(n852), .B(n853), .Z(n851) );
  NAND U859 ( .A(n853), .B(n852), .Z(n848) );
  ANDN U860 ( .B(B[81]), .A(n32), .Z(n787) );
  XNOR U861 ( .A(n795), .B(n854), .Z(n788) );
  XNOR U862 ( .A(n794), .B(n792), .Z(n854) );
  AND U863 ( .A(n855), .B(n856), .Z(n792) );
  NANDN U864 ( .A(n857), .B(n858), .Z(n856) );
  NANDN U865 ( .A(n859), .B(n860), .Z(n858) );
  NANDN U866 ( .A(n860), .B(n859), .Z(n855) );
  ANDN U867 ( .B(B[82]), .A(n33), .Z(n794) );
  XNOR U868 ( .A(n802), .B(n861), .Z(n795) );
  XNOR U869 ( .A(n801), .B(n799), .Z(n861) );
  AND U870 ( .A(n862), .B(n863), .Z(n799) );
  NANDN U871 ( .A(n864), .B(n865), .Z(n863) );
  OR U872 ( .A(n866), .B(n867), .Z(n865) );
  NAND U873 ( .A(n867), .B(n866), .Z(n862) );
  ANDN U874 ( .B(B[83]), .A(n34), .Z(n801) );
  XNOR U875 ( .A(n809), .B(n868), .Z(n802) );
  XNOR U876 ( .A(n808), .B(n806), .Z(n868) );
  AND U877 ( .A(n869), .B(n870), .Z(n806) );
  NANDN U878 ( .A(n871), .B(n872), .Z(n870) );
  NANDN U879 ( .A(n873), .B(n874), .Z(n872) );
  NANDN U880 ( .A(n874), .B(n873), .Z(n869) );
  ANDN U881 ( .B(B[84]), .A(n35), .Z(n808) );
  XOR U882 ( .A(n814), .B(n875), .Z(n809) );
  XNOR U883 ( .A(n815), .B(n816), .Z(n875) );
  AND U884 ( .A(n876), .B(n877), .Z(n816) );
  NANDN U885 ( .A(n878), .B(n879), .Z(n877) );
  NANDN U886 ( .A(n880), .B(n881), .Z(n879) );
  ANDN U887 ( .B(B[85]), .A(n36), .Z(n815) );
  XOR U888 ( .A(n882), .B(n883), .Z(n814) );
  XNOR U889 ( .A(n884), .B(n17), .Z(n883) );
  NAND U890 ( .A(n885), .B(n886), .Z(n60) );
  NANDN U891 ( .A(n887), .B(n888), .Z(n886) );
  OR U892 ( .A(n889), .B(n890), .Z(n888) );
  NAND U893 ( .A(n890), .B(n889), .Z(n885) );
  XOR U894 ( .A(n62), .B(n61), .Z(\A1[90] ) );
  XOR U895 ( .A(n890), .B(n891), .Z(n61) );
  XNOR U896 ( .A(n889), .B(n887), .Z(n891) );
  AND U897 ( .A(n892), .B(n893), .Z(n887) );
  NANDN U898 ( .A(n894), .B(n895), .Z(n893) );
  NANDN U899 ( .A(n896), .B(n897), .Z(n895) );
  NANDN U900 ( .A(n897), .B(n896), .Z(n892) );
  ANDN U901 ( .B(B[77]), .A(n29), .Z(n889) );
  XNOR U902 ( .A(n832), .B(n898), .Z(n890) );
  XNOR U903 ( .A(n831), .B(n829), .Z(n898) );
  AND U904 ( .A(n899), .B(n900), .Z(n829) );
  NANDN U905 ( .A(n901), .B(n902), .Z(n900) );
  OR U906 ( .A(n903), .B(n904), .Z(n902) );
  NAND U907 ( .A(n904), .B(n903), .Z(n899) );
  ANDN U908 ( .B(B[78]), .A(n30), .Z(n831) );
  XNOR U909 ( .A(n839), .B(n905), .Z(n832) );
  XNOR U910 ( .A(n838), .B(n836), .Z(n905) );
  AND U911 ( .A(n906), .B(n907), .Z(n836) );
  NANDN U912 ( .A(n908), .B(n909), .Z(n907) );
  NANDN U913 ( .A(n910), .B(n911), .Z(n909) );
  NANDN U914 ( .A(n911), .B(n910), .Z(n906) );
  ANDN U915 ( .B(B[79]), .A(n31), .Z(n838) );
  XNOR U916 ( .A(n846), .B(n912), .Z(n839) );
  XNOR U917 ( .A(n845), .B(n843), .Z(n912) );
  AND U918 ( .A(n913), .B(n914), .Z(n843) );
  NANDN U919 ( .A(n915), .B(n916), .Z(n914) );
  OR U920 ( .A(n917), .B(n918), .Z(n916) );
  NAND U921 ( .A(n918), .B(n917), .Z(n913) );
  ANDN U922 ( .B(B[80]), .A(n32), .Z(n845) );
  XNOR U923 ( .A(n853), .B(n919), .Z(n846) );
  XNOR U924 ( .A(n852), .B(n850), .Z(n919) );
  AND U925 ( .A(n920), .B(n921), .Z(n850) );
  NANDN U926 ( .A(n922), .B(n923), .Z(n921) );
  NANDN U927 ( .A(n924), .B(n925), .Z(n923) );
  NANDN U928 ( .A(n925), .B(n924), .Z(n920) );
  ANDN U929 ( .B(B[81]), .A(n33), .Z(n852) );
  XNOR U930 ( .A(n860), .B(n926), .Z(n853) );
  XNOR U931 ( .A(n859), .B(n857), .Z(n926) );
  AND U932 ( .A(n927), .B(n928), .Z(n857) );
  NANDN U933 ( .A(n929), .B(n930), .Z(n928) );
  OR U934 ( .A(n931), .B(n932), .Z(n930) );
  NAND U935 ( .A(n932), .B(n931), .Z(n927) );
  ANDN U936 ( .B(B[82]), .A(n34), .Z(n859) );
  XNOR U937 ( .A(n867), .B(n933), .Z(n860) );
  XNOR U938 ( .A(n866), .B(n864), .Z(n933) );
  AND U939 ( .A(n934), .B(n935), .Z(n864) );
  NANDN U940 ( .A(n936), .B(n937), .Z(n935) );
  NANDN U941 ( .A(n938), .B(n939), .Z(n937) );
  NANDN U942 ( .A(n939), .B(n938), .Z(n934) );
  ANDN U943 ( .B(B[83]), .A(n35), .Z(n866) );
  XNOR U944 ( .A(n874), .B(n940), .Z(n867) );
  XNOR U945 ( .A(n873), .B(n871), .Z(n940) );
  AND U946 ( .A(n941), .B(n942), .Z(n871) );
  NANDN U947 ( .A(n943), .B(n944), .Z(n942) );
  OR U948 ( .A(n945), .B(n946), .Z(n944) );
  NAND U949 ( .A(n946), .B(n945), .Z(n941) );
  ANDN U950 ( .B(B[84]), .A(n36), .Z(n873) );
  XOR U951 ( .A(n878), .B(n947), .Z(n874) );
  XNOR U952 ( .A(n880), .B(n881), .Z(n947) );
  AND U953 ( .A(n948), .B(n949), .Z(n881) );
  NAND U954 ( .A(n950), .B(n951), .Z(n949) );
  NANDN U955 ( .A(n952), .B(n953), .Z(n950) );
  ANDN U956 ( .B(B[85]), .A(n37), .Z(n880) );
  XNOR U957 ( .A(n954), .B(n955), .Z(n878) );
  XNOR U958 ( .A(n956), .B(n18), .Z(n955) );
  NAND U959 ( .A(n957), .B(n958), .Z(n62) );
  NANDN U960 ( .A(n959), .B(n960), .Z(n958) );
  OR U961 ( .A(n961), .B(n962), .Z(n960) );
  NAND U962 ( .A(n962), .B(n961), .Z(n957) );
  XNOR U963 ( .A(n963), .B(n964), .Z(\A1[8] ) );
  XNOR U964 ( .A(n965), .B(n966), .Z(n964) );
  XOR U965 ( .A(n64), .B(n63), .Z(\A1[89] ) );
  XOR U966 ( .A(n962), .B(n967), .Z(n63) );
  XNOR U967 ( .A(n961), .B(n959), .Z(n967) );
  AND U968 ( .A(n968), .B(n969), .Z(n959) );
  NANDN U969 ( .A(n970), .B(n971), .Z(n969) );
  NANDN U970 ( .A(n972), .B(n973), .Z(n971) );
  NANDN U971 ( .A(n973), .B(n972), .Z(n968) );
  ANDN U972 ( .B(B[76]), .A(n29), .Z(n961) );
  XNOR U973 ( .A(n897), .B(n974), .Z(n962) );
  XNOR U974 ( .A(n896), .B(n894), .Z(n974) );
  AND U975 ( .A(n975), .B(n976), .Z(n894) );
  NANDN U976 ( .A(n977), .B(n978), .Z(n976) );
  OR U977 ( .A(n979), .B(n980), .Z(n978) );
  NAND U978 ( .A(n980), .B(n979), .Z(n975) );
  ANDN U979 ( .B(B[77]), .A(n30), .Z(n896) );
  XNOR U980 ( .A(n904), .B(n981), .Z(n897) );
  XNOR U981 ( .A(n903), .B(n901), .Z(n981) );
  AND U982 ( .A(n982), .B(n983), .Z(n901) );
  NANDN U983 ( .A(n984), .B(n985), .Z(n983) );
  NANDN U984 ( .A(n986), .B(n987), .Z(n985) );
  NANDN U985 ( .A(n987), .B(n986), .Z(n982) );
  ANDN U986 ( .B(B[78]), .A(n31), .Z(n903) );
  XNOR U987 ( .A(n911), .B(n988), .Z(n904) );
  XNOR U988 ( .A(n910), .B(n908), .Z(n988) );
  AND U989 ( .A(n989), .B(n990), .Z(n908) );
  NANDN U990 ( .A(n991), .B(n992), .Z(n990) );
  OR U991 ( .A(n993), .B(n994), .Z(n992) );
  NAND U992 ( .A(n994), .B(n993), .Z(n989) );
  ANDN U993 ( .B(B[79]), .A(n32), .Z(n910) );
  XNOR U994 ( .A(n918), .B(n995), .Z(n911) );
  XNOR U995 ( .A(n917), .B(n915), .Z(n995) );
  AND U996 ( .A(n996), .B(n997), .Z(n915) );
  NANDN U997 ( .A(n998), .B(n999), .Z(n997) );
  NANDN U998 ( .A(n1000), .B(n1001), .Z(n999) );
  NANDN U999 ( .A(n1001), .B(n1000), .Z(n996) );
  ANDN U1000 ( .B(B[80]), .A(n33), .Z(n917) );
  XNOR U1001 ( .A(n925), .B(n1002), .Z(n918) );
  XNOR U1002 ( .A(n924), .B(n922), .Z(n1002) );
  AND U1003 ( .A(n1003), .B(n1004), .Z(n922) );
  NANDN U1004 ( .A(n1005), .B(n1006), .Z(n1004) );
  OR U1005 ( .A(n1007), .B(n1008), .Z(n1006) );
  NAND U1006 ( .A(n1008), .B(n1007), .Z(n1003) );
  ANDN U1007 ( .B(B[81]), .A(n34), .Z(n924) );
  XNOR U1008 ( .A(n932), .B(n1009), .Z(n925) );
  XNOR U1009 ( .A(n931), .B(n929), .Z(n1009) );
  AND U1010 ( .A(n1010), .B(n1011), .Z(n929) );
  NANDN U1011 ( .A(n1012), .B(n1013), .Z(n1011) );
  NANDN U1012 ( .A(n1014), .B(n1015), .Z(n1013) );
  NANDN U1013 ( .A(n1015), .B(n1014), .Z(n1010) );
  ANDN U1014 ( .B(B[82]), .A(n35), .Z(n931) );
  XNOR U1015 ( .A(n939), .B(n1016), .Z(n932) );
  XNOR U1016 ( .A(n938), .B(n936), .Z(n1016) );
  AND U1017 ( .A(n1017), .B(n1018), .Z(n936) );
  NANDN U1018 ( .A(n1019), .B(n1020), .Z(n1018) );
  OR U1019 ( .A(n1021), .B(n1022), .Z(n1020) );
  NAND U1020 ( .A(n1022), .B(n1021), .Z(n1017) );
  ANDN U1021 ( .B(B[83]), .A(n36), .Z(n938) );
  XNOR U1022 ( .A(n946), .B(n1023), .Z(n939) );
  XNOR U1023 ( .A(n945), .B(n943), .Z(n1023) );
  AND U1024 ( .A(n1024), .B(n1025), .Z(n943) );
  NANDN U1025 ( .A(n1026), .B(n1027), .Z(n1025) );
  NANDN U1026 ( .A(n1028), .B(n1029), .Z(n1027) );
  NANDN U1027 ( .A(n1029), .B(n1028), .Z(n1024) );
  ANDN U1028 ( .B(B[84]), .A(n37), .Z(n945) );
  XOR U1029 ( .A(n951), .B(n1030), .Z(n946) );
  XNOR U1030 ( .A(n952), .B(n953), .Z(n1030) );
  AND U1031 ( .A(n1031), .B(n1032), .Z(n953) );
  NANDN U1032 ( .A(n1033), .B(n1034), .Z(n1032) );
  NANDN U1033 ( .A(n1035), .B(n1036), .Z(n1034) );
  ANDN U1034 ( .B(B[85]), .A(n38), .Z(n952) );
  XOR U1035 ( .A(n1037), .B(n1038), .Z(n951) );
  XNOR U1036 ( .A(n1039), .B(n19), .Z(n1038) );
  NAND U1037 ( .A(n1040), .B(n1041), .Z(n64) );
  NANDN U1038 ( .A(n1042), .B(n1043), .Z(n1041) );
  OR U1039 ( .A(n1044), .B(n1045), .Z(n1043) );
  NAND U1040 ( .A(n1045), .B(n1044), .Z(n1040) );
  XOR U1041 ( .A(n66), .B(n65), .Z(\A1[88] ) );
  XOR U1042 ( .A(n1045), .B(n1046), .Z(n65) );
  XNOR U1043 ( .A(n1044), .B(n1042), .Z(n1046) );
  AND U1044 ( .A(n1047), .B(n1048), .Z(n1042) );
  NANDN U1045 ( .A(n1049), .B(n1050), .Z(n1048) );
  NANDN U1046 ( .A(n1051), .B(n1052), .Z(n1050) );
  NANDN U1047 ( .A(n1052), .B(n1051), .Z(n1047) );
  ANDN U1048 ( .B(B[75]), .A(n29), .Z(n1044) );
  XNOR U1049 ( .A(n973), .B(n1053), .Z(n1045) );
  XNOR U1050 ( .A(n972), .B(n970), .Z(n1053) );
  AND U1051 ( .A(n1054), .B(n1055), .Z(n970) );
  NANDN U1052 ( .A(n1056), .B(n1057), .Z(n1055) );
  OR U1053 ( .A(n1058), .B(n1059), .Z(n1057) );
  NAND U1054 ( .A(n1059), .B(n1058), .Z(n1054) );
  ANDN U1055 ( .B(B[76]), .A(n30), .Z(n972) );
  XNOR U1056 ( .A(n980), .B(n1060), .Z(n973) );
  XNOR U1057 ( .A(n979), .B(n977), .Z(n1060) );
  AND U1058 ( .A(n1061), .B(n1062), .Z(n977) );
  NANDN U1059 ( .A(n1063), .B(n1064), .Z(n1062) );
  NANDN U1060 ( .A(n1065), .B(n1066), .Z(n1064) );
  NANDN U1061 ( .A(n1066), .B(n1065), .Z(n1061) );
  ANDN U1062 ( .B(B[77]), .A(n31), .Z(n979) );
  XNOR U1063 ( .A(n987), .B(n1067), .Z(n980) );
  XNOR U1064 ( .A(n986), .B(n984), .Z(n1067) );
  AND U1065 ( .A(n1068), .B(n1069), .Z(n984) );
  NANDN U1066 ( .A(n1070), .B(n1071), .Z(n1069) );
  OR U1067 ( .A(n1072), .B(n1073), .Z(n1071) );
  NAND U1068 ( .A(n1073), .B(n1072), .Z(n1068) );
  ANDN U1069 ( .B(B[78]), .A(n32), .Z(n986) );
  XNOR U1070 ( .A(n994), .B(n1074), .Z(n987) );
  XNOR U1071 ( .A(n993), .B(n991), .Z(n1074) );
  AND U1072 ( .A(n1075), .B(n1076), .Z(n991) );
  NANDN U1073 ( .A(n1077), .B(n1078), .Z(n1076) );
  NANDN U1074 ( .A(n1079), .B(n1080), .Z(n1078) );
  NANDN U1075 ( .A(n1080), .B(n1079), .Z(n1075) );
  ANDN U1076 ( .B(B[79]), .A(n33), .Z(n993) );
  XNOR U1077 ( .A(n1001), .B(n1081), .Z(n994) );
  XNOR U1078 ( .A(n1000), .B(n998), .Z(n1081) );
  AND U1079 ( .A(n1082), .B(n1083), .Z(n998) );
  NANDN U1080 ( .A(n1084), .B(n1085), .Z(n1083) );
  OR U1081 ( .A(n1086), .B(n1087), .Z(n1085) );
  NAND U1082 ( .A(n1087), .B(n1086), .Z(n1082) );
  ANDN U1083 ( .B(B[80]), .A(n34), .Z(n1000) );
  XNOR U1084 ( .A(n1008), .B(n1088), .Z(n1001) );
  XNOR U1085 ( .A(n1007), .B(n1005), .Z(n1088) );
  AND U1086 ( .A(n1089), .B(n1090), .Z(n1005) );
  NANDN U1087 ( .A(n1091), .B(n1092), .Z(n1090) );
  NANDN U1088 ( .A(n1093), .B(n1094), .Z(n1092) );
  NANDN U1089 ( .A(n1094), .B(n1093), .Z(n1089) );
  ANDN U1090 ( .B(B[81]), .A(n35), .Z(n1007) );
  XNOR U1091 ( .A(n1015), .B(n1095), .Z(n1008) );
  XNOR U1092 ( .A(n1014), .B(n1012), .Z(n1095) );
  AND U1093 ( .A(n1096), .B(n1097), .Z(n1012) );
  NANDN U1094 ( .A(n1098), .B(n1099), .Z(n1097) );
  OR U1095 ( .A(n1100), .B(n1101), .Z(n1099) );
  NAND U1096 ( .A(n1101), .B(n1100), .Z(n1096) );
  ANDN U1097 ( .B(B[82]), .A(n36), .Z(n1014) );
  XNOR U1098 ( .A(n1022), .B(n1102), .Z(n1015) );
  XNOR U1099 ( .A(n1021), .B(n1019), .Z(n1102) );
  AND U1100 ( .A(n1103), .B(n1104), .Z(n1019) );
  NANDN U1101 ( .A(n1105), .B(n1106), .Z(n1104) );
  NANDN U1102 ( .A(n1107), .B(n1108), .Z(n1106) );
  NANDN U1103 ( .A(n1108), .B(n1107), .Z(n1103) );
  ANDN U1104 ( .B(B[83]), .A(n37), .Z(n1021) );
  XNOR U1105 ( .A(n1029), .B(n1109), .Z(n1022) );
  XNOR U1106 ( .A(n1028), .B(n1026), .Z(n1109) );
  AND U1107 ( .A(n1110), .B(n1111), .Z(n1026) );
  NANDN U1108 ( .A(n1112), .B(n1113), .Z(n1111) );
  OR U1109 ( .A(n1114), .B(n1115), .Z(n1113) );
  NAND U1110 ( .A(n1115), .B(n1114), .Z(n1110) );
  ANDN U1111 ( .B(B[84]), .A(n38), .Z(n1028) );
  XOR U1112 ( .A(n1033), .B(n1116), .Z(n1029) );
  XNOR U1113 ( .A(n1035), .B(n1036), .Z(n1116) );
  AND U1114 ( .A(n1117), .B(n1118), .Z(n1036) );
  NAND U1115 ( .A(n1119), .B(n1120), .Z(n1118) );
  NANDN U1116 ( .A(n1121), .B(n1122), .Z(n1119) );
  ANDN U1117 ( .B(B[85]), .A(n39), .Z(n1035) );
  XNOR U1118 ( .A(n1123), .B(n1124), .Z(n1033) );
  XNOR U1119 ( .A(n1125), .B(n20), .Z(n1124) );
  NAND U1120 ( .A(n1126), .B(n1127), .Z(n66) );
  NANDN U1121 ( .A(n1128), .B(n1129), .Z(n1127) );
  OR U1122 ( .A(n1130), .B(n1131), .Z(n1129) );
  NAND U1123 ( .A(n1131), .B(n1130), .Z(n1126) );
  XOR U1124 ( .A(n68), .B(n67), .Z(\A1[87] ) );
  XOR U1125 ( .A(n1131), .B(n1132), .Z(n67) );
  XNOR U1126 ( .A(n1130), .B(n1128), .Z(n1132) );
  AND U1127 ( .A(n1133), .B(n1134), .Z(n1128) );
  NANDN U1128 ( .A(n1135), .B(n1136), .Z(n1134) );
  NANDN U1129 ( .A(n1137), .B(n1138), .Z(n1136) );
  NANDN U1130 ( .A(n1138), .B(n1137), .Z(n1133) );
  ANDN U1131 ( .B(B[74]), .A(n29), .Z(n1130) );
  XNOR U1132 ( .A(n1052), .B(n1139), .Z(n1131) );
  XNOR U1133 ( .A(n1051), .B(n1049), .Z(n1139) );
  AND U1134 ( .A(n1140), .B(n1141), .Z(n1049) );
  NANDN U1135 ( .A(n1142), .B(n1143), .Z(n1141) );
  OR U1136 ( .A(n1144), .B(n1145), .Z(n1143) );
  NAND U1137 ( .A(n1145), .B(n1144), .Z(n1140) );
  ANDN U1138 ( .B(B[75]), .A(n30), .Z(n1051) );
  XNOR U1139 ( .A(n1059), .B(n1146), .Z(n1052) );
  XNOR U1140 ( .A(n1058), .B(n1056), .Z(n1146) );
  AND U1141 ( .A(n1147), .B(n1148), .Z(n1056) );
  NANDN U1142 ( .A(n1149), .B(n1150), .Z(n1148) );
  NANDN U1143 ( .A(n1151), .B(n1152), .Z(n1150) );
  NANDN U1144 ( .A(n1152), .B(n1151), .Z(n1147) );
  ANDN U1145 ( .B(B[76]), .A(n31), .Z(n1058) );
  XNOR U1146 ( .A(n1066), .B(n1153), .Z(n1059) );
  XNOR U1147 ( .A(n1065), .B(n1063), .Z(n1153) );
  AND U1148 ( .A(n1154), .B(n1155), .Z(n1063) );
  NANDN U1149 ( .A(n1156), .B(n1157), .Z(n1155) );
  OR U1150 ( .A(n1158), .B(n1159), .Z(n1157) );
  NAND U1151 ( .A(n1159), .B(n1158), .Z(n1154) );
  ANDN U1152 ( .B(B[77]), .A(n32), .Z(n1065) );
  XNOR U1153 ( .A(n1073), .B(n1160), .Z(n1066) );
  XNOR U1154 ( .A(n1072), .B(n1070), .Z(n1160) );
  AND U1155 ( .A(n1161), .B(n1162), .Z(n1070) );
  NANDN U1156 ( .A(n1163), .B(n1164), .Z(n1162) );
  NANDN U1157 ( .A(n1165), .B(n1166), .Z(n1164) );
  NANDN U1158 ( .A(n1166), .B(n1165), .Z(n1161) );
  ANDN U1159 ( .B(B[78]), .A(n33), .Z(n1072) );
  XNOR U1160 ( .A(n1080), .B(n1167), .Z(n1073) );
  XNOR U1161 ( .A(n1079), .B(n1077), .Z(n1167) );
  AND U1162 ( .A(n1168), .B(n1169), .Z(n1077) );
  NANDN U1163 ( .A(n1170), .B(n1171), .Z(n1169) );
  OR U1164 ( .A(n1172), .B(n1173), .Z(n1171) );
  NAND U1165 ( .A(n1173), .B(n1172), .Z(n1168) );
  ANDN U1166 ( .B(B[79]), .A(n34), .Z(n1079) );
  XNOR U1167 ( .A(n1087), .B(n1174), .Z(n1080) );
  XNOR U1168 ( .A(n1086), .B(n1084), .Z(n1174) );
  AND U1169 ( .A(n1175), .B(n1176), .Z(n1084) );
  NANDN U1170 ( .A(n1177), .B(n1178), .Z(n1176) );
  NANDN U1171 ( .A(n1179), .B(n1180), .Z(n1178) );
  NANDN U1172 ( .A(n1180), .B(n1179), .Z(n1175) );
  ANDN U1173 ( .B(B[80]), .A(n35), .Z(n1086) );
  XNOR U1174 ( .A(n1094), .B(n1181), .Z(n1087) );
  XNOR U1175 ( .A(n1093), .B(n1091), .Z(n1181) );
  AND U1176 ( .A(n1182), .B(n1183), .Z(n1091) );
  NANDN U1177 ( .A(n1184), .B(n1185), .Z(n1183) );
  OR U1178 ( .A(n1186), .B(n1187), .Z(n1185) );
  NAND U1179 ( .A(n1187), .B(n1186), .Z(n1182) );
  ANDN U1180 ( .B(B[81]), .A(n36), .Z(n1093) );
  XNOR U1181 ( .A(n1101), .B(n1188), .Z(n1094) );
  XNOR U1182 ( .A(n1100), .B(n1098), .Z(n1188) );
  AND U1183 ( .A(n1189), .B(n1190), .Z(n1098) );
  NANDN U1184 ( .A(n1191), .B(n1192), .Z(n1190) );
  NANDN U1185 ( .A(n1193), .B(n1194), .Z(n1192) );
  NANDN U1186 ( .A(n1194), .B(n1193), .Z(n1189) );
  ANDN U1187 ( .B(B[82]), .A(n37), .Z(n1100) );
  XNOR U1188 ( .A(n1108), .B(n1195), .Z(n1101) );
  XNOR U1189 ( .A(n1107), .B(n1105), .Z(n1195) );
  AND U1190 ( .A(n1196), .B(n1197), .Z(n1105) );
  NANDN U1191 ( .A(n1198), .B(n1199), .Z(n1197) );
  OR U1192 ( .A(n1200), .B(n1201), .Z(n1199) );
  NAND U1193 ( .A(n1201), .B(n1200), .Z(n1196) );
  ANDN U1194 ( .B(B[83]), .A(n38), .Z(n1107) );
  XNOR U1195 ( .A(n1115), .B(n1202), .Z(n1108) );
  XNOR U1196 ( .A(n1114), .B(n1112), .Z(n1202) );
  AND U1197 ( .A(n1203), .B(n1204), .Z(n1112) );
  NANDN U1198 ( .A(n1205), .B(n1206), .Z(n1204) );
  NANDN U1199 ( .A(n1207), .B(n1208), .Z(n1206) );
  NANDN U1200 ( .A(n1208), .B(n1207), .Z(n1203) );
  ANDN U1201 ( .B(B[84]), .A(n39), .Z(n1114) );
  XOR U1202 ( .A(n1120), .B(n1209), .Z(n1115) );
  XNOR U1203 ( .A(n1121), .B(n1122), .Z(n1209) );
  AND U1204 ( .A(n1210), .B(n1211), .Z(n1122) );
  NANDN U1205 ( .A(n1212), .B(n1213), .Z(n1211) );
  NANDN U1206 ( .A(n1214), .B(n1215), .Z(n1213) );
  ANDN U1207 ( .B(B[85]), .A(n40), .Z(n1121) );
  XNOR U1208 ( .A(n1216), .B(n1217), .Z(n1120) );
  XNOR U1209 ( .A(n1218), .B(n22), .Z(n1217) );
  NAND U1210 ( .A(n1219), .B(n1220), .Z(n68) );
  NANDN U1211 ( .A(n1221), .B(n1222), .Z(n1220) );
  OR U1212 ( .A(n1223), .B(n1224), .Z(n1222) );
  NAND U1213 ( .A(n1224), .B(n1223), .Z(n1219) );
  XOR U1214 ( .A(n70), .B(n69), .Z(\A1[86] ) );
  XOR U1215 ( .A(n1224), .B(n1225), .Z(n69) );
  XNOR U1216 ( .A(n1223), .B(n1221), .Z(n1225) );
  AND U1217 ( .A(n1226), .B(n1227), .Z(n1221) );
  NANDN U1218 ( .A(n1228), .B(n1229), .Z(n1227) );
  NANDN U1219 ( .A(n1230), .B(n1231), .Z(n1229) );
  NANDN U1220 ( .A(n1231), .B(n1230), .Z(n1226) );
  ANDN U1221 ( .B(B[73]), .A(n29), .Z(n1223) );
  XNOR U1222 ( .A(n1138), .B(n1232), .Z(n1224) );
  XNOR U1223 ( .A(n1137), .B(n1135), .Z(n1232) );
  AND U1224 ( .A(n1233), .B(n1234), .Z(n1135) );
  NANDN U1225 ( .A(n1235), .B(n1236), .Z(n1234) );
  OR U1226 ( .A(n1237), .B(n1238), .Z(n1236) );
  NAND U1227 ( .A(n1238), .B(n1237), .Z(n1233) );
  ANDN U1228 ( .B(B[74]), .A(n30), .Z(n1137) );
  XNOR U1229 ( .A(n1145), .B(n1239), .Z(n1138) );
  XNOR U1230 ( .A(n1144), .B(n1142), .Z(n1239) );
  AND U1231 ( .A(n1240), .B(n1241), .Z(n1142) );
  NANDN U1232 ( .A(n1242), .B(n1243), .Z(n1241) );
  NANDN U1233 ( .A(n1244), .B(n1245), .Z(n1243) );
  NANDN U1234 ( .A(n1245), .B(n1244), .Z(n1240) );
  ANDN U1235 ( .B(B[75]), .A(n31), .Z(n1144) );
  XNOR U1236 ( .A(n1152), .B(n1246), .Z(n1145) );
  XNOR U1237 ( .A(n1151), .B(n1149), .Z(n1246) );
  AND U1238 ( .A(n1247), .B(n1248), .Z(n1149) );
  NANDN U1239 ( .A(n1249), .B(n1250), .Z(n1248) );
  OR U1240 ( .A(n1251), .B(n1252), .Z(n1250) );
  NAND U1241 ( .A(n1252), .B(n1251), .Z(n1247) );
  ANDN U1242 ( .B(B[76]), .A(n32), .Z(n1151) );
  XNOR U1243 ( .A(n1159), .B(n1253), .Z(n1152) );
  XNOR U1244 ( .A(n1158), .B(n1156), .Z(n1253) );
  AND U1245 ( .A(n1254), .B(n1255), .Z(n1156) );
  NANDN U1246 ( .A(n1256), .B(n1257), .Z(n1255) );
  NANDN U1247 ( .A(n1258), .B(n1259), .Z(n1257) );
  NANDN U1248 ( .A(n1259), .B(n1258), .Z(n1254) );
  ANDN U1249 ( .B(B[77]), .A(n33), .Z(n1158) );
  XNOR U1250 ( .A(n1166), .B(n1260), .Z(n1159) );
  XNOR U1251 ( .A(n1165), .B(n1163), .Z(n1260) );
  AND U1252 ( .A(n1261), .B(n1262), .Z(n1163) );
  NANDN U1253 ( .A(n1263), .B(n1264), .Z(n1262) );
  OR U1254 ( .A(n1265), .B(n1266), .Z(n1264) );
  NAND U1255 ( .A(n1266), .B(n1265), .Z(n1261) );
  ANDN U1256 ( .B(B[78]), .A(n34), .Z(n1165) );
  XNOR U1257 ( .A(n1173), .B(n1267), .Z(n1166) );
  XNOR U1258 ( .A(n1172), .B(n1170), .Z(n1267) );
  AND U1259 ( .A(n1268), .B(n1269), .Z(n1170) );
  NANDN U1260 ( .A(n1270), .B(n1271), .Z(n1269) );
  NANDN U1261 ( .A(n1272), .B(n1273), .Z(n1271) );
  NANDN U1262 ( .A(n1273), .B(n1272), .Z(n1268) );
  ANDN U1263 ( .B(B[79]), .A(n35), .Z(n1172) );
  XNOR U1264 ( .A(n1180), .B(n1274), .Z(n1173) );
  XNOR U1265 ( .A(n1179), .B(n1177), .Z(n1274) );
  AND U1266 ( .A(n1275), .B(n1276), .Z(n1177) );
  NANDN U1267 ( .A(n1277), .B(n1278), .Z(n1276) );
  OR U1268 ( .A(n1279), .B(n1280), .Z(n1278) );
  NAND U1269 ( .A(n1280), .B(n1279), .Z(n1275) );
  ANDN U1270 ( .B(B[80]), .A(n36), .Z(n1179) );
  XNOR U1271 ( .A(n1187), .B(n1281), .Z(n1180) );
  XNOR U1272 ( .A(n1186), .B(n1184), .Z(n1281) );
  AND U1273 ( .A(n1282), .B(n1283), .Z(n1184) );
  NANDN U1274 ( .A(n1284), .B(n1285), .Z(n1283) );
  NANDN U1275 ( .A(n1286), .B(n1287), .Z(n1285) );
  NANDN U1276 ( .A(n1287), .B(n1286), .Z(n1282) );
  ANDN U1277 ( .B(B[81]), .A(n37), .Z(n1186) );
  XNOR U1278 ( .A(n1194), .B(n1288), .Z(n1187) );
  XNOR U1279 ( .A(n1193), .B(n1191), .Z(n1288) );
  AND U1280 ( .A(n1289), .B(n1290), .Z(n1191) );
  NANDN U1281 ( .A(n1291), .B(n1292), .Z(n1290) );
  OR U1282 ( .A(n1293), .B(n1294), .Z(n1292) );
  NAND U1283 ( .A(n1294), .B(n1293), .Z(n1289) );
  ANDN U1284 ( .B(B[82]), .A(n38), .Z(n1193) );
  XNOR U1285 ( .A(n1201), .B(n1295), .Z(n1194) );
  XNOR U1286 ( .A(n1200), .B(n1198), .Z(n1295) );
  AND U1287 ( .A(n1296), .B(n1297), .Z(n1198) );
  NANDN U1288 ( .A(n1298), .B(n1299), .Z(n1297) );
  NANDN U1289 ( .A(n1300), .B(n1301), .Z(n1299) );
  NANDN U1290 ( .A(n1301), .B(n1300), .Z(n1296) );
  ANDN U1291 ( .B(B[83]), .A(n39), .Z(n1200) );
  XNOR U1292 ( .A(n1208), .B(n1302), .Z(n1201) );
  XNOR U1293 ( .A(n1207), .B(n1205), .Z(n1302) );
  AND U1294 ( .A(n1303), .B(n1304), .Z(n1205) );
  NANDN U1295 ( .A(n1305), .B(n1306), .Z(n1304) );
  NANDN U1296 ( .A(n1307), .B(n1308), .Z(n1306) );
  NAND U1297 ( .A(n23), .B(n1307), .Z(n1303) );
  ANDN U1298 ( .B(B[84]), .A(n40), .Z(n1207) );
  XOR U1299 ( .A(n1212), .B(n1309), .Z(n1208) );
  XNOR U1300 ( .A(n1214), .B(n1215), .Z(n1309) );
  AND U1301 ( .A(n1310), .B(n1311), .Z(n1215) );
  NANDN U1302 ( .A(n1312), .B(n1313), .Z(n1311) );
  NANDN U1303 ( .A(n1314), .B(n1315), .Z(n1313) );
  NANDN U1304 ( .A(n1315), .B(n1314), .Z(n1310) );
  ANDN U1305 ( .B(B[85]), .A(n41), .Z(n1214) );
  XNOR U1306 ( .A(n1316), .B(n1317), .Z(n1212) );
  XOR U1307 ( .A(n1318), .B(n1319), .Z(n1317) );
  NAND U1308 ( .A(n1320), .B(n1321), .Z(n70) );
  NANDN U1309 ( .A(n1322), .B(n1323), .Z(n1321) );
  OR U1310 ( .A(n1324), .B(n1325), .Z(n1323) );
  NAND U1311 ( .A(n1325), .B(n1324), .Z(n1320) );
  XOR U1312 ( .A(n72), .B(n71), .Z(\A1[85] ) );
  XOR U1313 ( .A(n1325), .B(n1326), .Z(n71) );
  XNOR U1314 ( .A(n1324), .B(n1322), .Z(n1326) );
  AND U1315 ( .A(n1327), .B(n1328), .Z(n1322) );
  NANDN U1316 ( .A(n1329), .B(n1330), .Z(n1328) );
  NANDN U1317 ( .A(n1331), .B(n1332), .Z(n1330) );
  NANDN U1318 ( .A(n1332), .B(n1331), .Z(n1327) );
  ANDN U1319 ( .B(B[72]), .A(n29), .Z(n1324) );
  XNOR U1320 ( .A(n1231), .B(n1333), .Z(n1325) );
  XNOR U1321 ( .A(n1230), .B(n1228), .Z(n1333) );
  AND U1322 ( .A(n1334), .B(n1335), .Z(n1228) );
  NANDN U1323 ( .A(n1336), .B(n1337), .Z(n1335) );
  OR U1324 ( .A(n1338), .B(n1339), .Z(n1337) );
  NAND U1325 ( .A(n1339), .B(n1338), .Z(n1334) );
  ANDN U1326 ( .B(B[73]), .A(n30), .Z(n1230) );
  XNOR U1327 ( .A(n1238), .B(n1340), .Z(n1231) );
  XNOR U1328 ( .A(n1237), .B(n1235), .Z(n1340) );
  AND U1329 ( .A(n1341), .B(n1342), .Z(n1235) );
  NANDN U1330 ( .A(n1343), .B(n1344), .Z(n1342) );
  NANDN U1331 ( .A(n1345), .B(n1346), .Z(n1344) );
  NANDN U1332 ( .A(n1346), .B(n1345), .Z(n1341) );
  ANDN U1333 ( .B(B[74]), .A(n31), .Z(n1237) );
  XNOR U1334 ( .A(n1245), .B(n1347), .Z(n1238) );
  XNOR U1335 ( .A(n1244), .B(n1242), .Z(n1347) );
  AND U1336 ( .A(n1348), .B(n1349), .Z(n1242) );
  NANDN U1337 ( .A(n1350), .B(n1351), .Z(n1349) );
  OR U1338 ( .A(n1352), .B(n1353), .Z(n1351) );
  NAND U1339 ( .A(n1353), .B(n1352), .Z(n1348) );
  ANDN U1340 ( .B(B[75]), .A(n32), .Z(n1244) );
  XNOR U1341 ( .A(n1252), .B(n1354), .Z(n1245) );
  XNOR U1342 ( .A(n1251), .B(n1249), .Z(n1354) );
  AND U1343 ( .A(n1355), .B(n1356), .Z(n1249) );
  NANDN U1344 ( .A(n1357), .B(n1358), .Z(n1356) );
  NANDN U1345 ( .A(n1359), .B(n1360), .Z(n1358) );
  NANDN U1346 ( .A(n1360), .B(n1359), .Z(n1355) );
  ANDN U1347 ( .B(B[76]), .A(n33), .Z(n1251) );
  XNOR U1348 ( .A(n1259), .B(n1361), .Z(n1252) );
  XNOR U1349 ( .A(n1258), .B(n1256), .Z(n1361) );
  AND U1350 ( .A(n1362), .B(n1363), .Z(n1256) );
  NANDN U1351 ( .A(n1364), .B(n1365), .Z(n1363) );
  OR U1352 ( .A(n1366), .B(n1367), .Z(n1365) );
  NAND U1353 ( .A(n1367), .B(n1366), .Z(n1362) );
  ANDN U1354 ( .B(B[77]), .A(n34), .Z(n1258) );
  XNOR U1355 ( .A(n1266), .B(n1368), .Z(n1259) );
  XNOR U1356 ( .A(n1265), .B(n1263), .Z(n1368) );
  AND U1357 ( .A(n1369), .B(n1370), .Z(n1263) );
  NANDN U1358 ( .A(n1371), .B(n1372), .Z(n1370) );
  NANDN U1359 ( .A(n1373), .B(n1374), .Z(n1372) );
  NANDN U1360 ( .A(n1374), .B(n1373), .Z(n1369) );
  ANDN U1361 ( .B(B[78]), .A(n35), .Z(n1265) );
  XNOR U1362 ( .A(n1273), .B(n1375), .Z(n1266) );
  XNOR U1363 ( .A(n1272), .B(n1270), .Z(n1375) );
  AND U1364 ( .A(n1376), .B(n1377), .Z(n1270) );
  NANDN U1365 ( .A(n1378), .B(n1379), .Z(n1377) );
  OR U1366 ( .A(n1380), .B(n1381), .Z(n1379) );
  NAND U1367 ( .A(n1381), .B(n1380), .Z(n1376) );
  ANDN U1368 ( .B(B[79]), .A(n36), .Z(n1272) );
  XNOR U1369 ( .A(n1280), .B(n1382), .Z(n1273) );
  XNOR U1370 ( .A(n1279), .B(n1277), .Z(n1382) );
  AND U1371 ( .A(n1383), .B(n1384), .Z(n1277) );
  NANDN U1372 ( .A(n1385), .B(n1386), .Z(n1384) );
  NANDN U1373 ( .A(n1387), .B(n1388), .Z(n1386) );
  NANDN U1374 ( .A(n1388), .B(n1387), .Z(n1383) );
  ANDN U1375 ( .B(B[80]), .A(n37), .Z(n1279) );
  XNOR U1376 ( .A(n1287), .B(n1389), .Z(n1280) );
  XNOR U1377 ( .A(n1286), .B(n1284), .Z(n1389) );
  AND U1378 ( .A(n1390), .B(n1391), .Z(n1284) );
  NANDN U1379 ( .A(n1392), .B(n1393), .Z(n1391) );
  OR U1380 ( .A(n1394), .B(n1395), .Z(n1393) );
  NAND U1381 ( .A(n1395), .B(n1394), .Z(n1390) );
  ANDN U1382 ( .B(B[81]), .A(n38), .Z(n1286) );
  XNOR U1383 ( .A(n1294), .B(n1396), .Z(n1287) );
  XNOR U1384 ( .A(n1293), .B(n1291), .Z(n1396) );
  AND U1385 ( .A(n1397), .B(n1398), .Z(n1291) );
  NANDN U1386 ( .A(n1399), .B(n1400), .Z(n1398) );
  NANDN U1387 ( .A(n1401), .B(n1402), .Z(n1400) );
  NANDN U1388 ( .A(n1402), .B(n1401), .Z(n1397) );
  ANDN U1389 ( .B(B[82]), .A(n39), .Z(n1293) );
  XNOR U1390 ( .A(n1301), .B(n1403), .Z(n1294) );
  XNOR U1391 ( .A(n1300), .B(n1298), .Z(n1403) );
  AND U1392 ( .A(n1404), .B(n1405), .Z(n1298) );
  NANDN U1393 ( .A(n1406), .B(n1407), .Z(n1405) );
  OR U1394 ( .A(n1408), .B(n1409), .Z(n1407) );
  NAND U1395 ( .A(n1409), .B(n1408), .Z(n1404) );
  ANDN U1396 ( .B(B[83]), .A(n40), .Z(n1300) );
  XNOR U1397 ( .A(n23), .B(n1410), .Z(n1301) );
  XNOR U1398 ( .A(n1307), .B(n1305), .Z(n1410) );
  AND U1399 ( .A(n1411), .B(n1412), .Z(n1305) );
  NANDN U1400 ( .A(n1413), .B(n1414), .Z(n1412) );
  NAND U1401 ( .A(n1415), .B(n1416), .Z(n1414) );
  ANDN U1402 ( .B(B[84]), .A(n41), .Z(n1307) );
  XNOR U1403 ( .A(n1312), .B(n1417), .Z(n1308) );
  XOR U1404 ( .A(n1314), .B(n1315), .Z(n1417) );
  NAND U1405 ( .A(B[85]), .B(A[2]), .Z(n1315) );
  ANDN U1406 ( .B(n1418), .A(n1419), .Z(n1314) );
  AND U1407 ( .A(A[0]), .B(B[86]), .Z(n1418) );
  XNOR U1408 ( .A(n1420), .B(n1421), .Z(n1312) );
  NAND U1409 ( .A(B[87]), .B(A[0]), .Z(n1421) );
  NAND U1410 ( .A(n1422), .B(n1423), .Z(n72) );
  NANDN U1411 ( .A(n1424), .B(n1425), .Z(n1423) );
  OR U1412 ( .A(n1426), .B(n1427), .Z(n1425) );
  NAND U1413 ( .A(n1427), .B(n1426), .Z(n1422) );
  XOR U1414 ( .A(n74), .B(n73), .Z(\A1[84] ) );
  XOR U1415 ( .A(n1427), .B(n1428), .Z(n73) );
  XNOR U1416 ( .A(n1426), .B(n1424), .Z(n1428) );
  AND U1417 ( .A(n1429), .B(n1430), .Z(n1424) );
  NANDN U1418 ( .A(n1431), .B(n1432), .Z(n1430) );
  NANDN U1419 ( .A(n1433), .B(n1434), .Z(n1432) );
  NANDN U1420 ( .A(n1434), .B(n1433), .Z(n1429) );
  ANDN U1421 ( .B(B[71]), .A(n29), .Z(n1426) );
  XNOR U1422 ( .A(n1332), .B(n1435), .Z(n1427) );
  XNOR U1423 ( .A(n1331), .B(n1329), .Z(n1435) );
  AND U1424 ( .A(n1436), .B(n1437), .Z(n1329) );
  NANDN U1425 ( .A(n1438), .B(n1439), .Z(n1437) );
  OR U1426 ( .A(n1440), .B(n1441), .Z(n1439) );
  NAND U1427 ( .A(n1441), .B(n1440), .Z(n1436) );
  ANDN U1428 ( .B(B[72]), .A(n30), .Z(n1331) );
  XNOR U1429 ( .A(n1339), .B(n1442), .Z(n1332) );
  XNOR U1430 ( .A(n1338), .B(n1336), .Z(n1442) );
  AND U1431 ( .A(n1443), .B(n1444), .Z(n1336) );
  NANDN U1432 ( .A(n1445), .B(n1446), .Z(n1444) );
  NANDN U1433 ( .A(n1447), .B(n1448), .Z(n1446) );
  NANDN U1434 ( .A(n1448), .B(n1447), .Z(n1443) );
  ANDN U1435 ( .B(B[73]), .A(n31), .Z(n1338) );
  XNOR U1436 ( .A(n1346), .B(n1449), .Z(n1339) );
  XNOR U1437 ( .A(n1345), .B(n1343), .Z(n1449) );
  AND U1438 ( .A(n1450), .B(n1451), .Z(n1343) );
  NANDN U1439 ( .A(n1452), .B(n1453), .Z(n1451) );
  OR U1440 ( .A(n1454), .B(n1455), .Z(n1453) );
  NAND U1441 ( .A(n1455), .B(n1454), .Z(n1450) );
  ANDN U1442 ( .B(B[74]), .A(n32), .Z(n1345) );
  XNOR U1443 ( .A(n1353), .B(n1456), .Z(n1346) );
  XNOR U1444 ( .A(n1352), .B(n1350), .Z(n1456) );
  AND U1445 ( .A(n1457), .B(n1458), .Z(n1350) );
  NANDN U1446 ( .A(n1459), .B(n1460), .Z(n1458) );
  NANDN U1447 ( .A(n1461), .B(n1462), .Z(n1460) );
  NANDN U1448 ( .A(n1462), .B(n1461), .Z(n1457) );
  ANDN U1449 ( .B(B[75]), .A(n33), .Z(n1352) );
  XNOR U1450 ( .A(n1360), .B(n1463), .Z(n1353) );
  XNOR U1451 ( .A(n1359), .B(n1357), .Z(n1463) );
  AND U1452 ( .A(n1464), .B(n1465), .Z(n1357) );
  NANDN U1453 ( .A(n1466), .B(n1467), .Z(n1465) );
  OR U1454 ( .A(n1468), .B(n1469), .Z(n1467) );
  NAND U1455 ( .A(n1469), .B(n1468), .Z(n1464) );
  ANDN U1456 ( .B(B[76]), .A(n34), .Z(n1359) );
  XNOR U1457 ( .A(n1367), .B(n1470), .Z(n1360) );
  XNOR U1458 ( .A(n1366), .B(n1364), .Z(n1470) );
  AND U1459 ( .A(n1471), .B(n1472), .Z(n1364) );
  NANDN U1460 ( .A(n1473), .B(n1474), .Z(n1472) );
  NANDN U1461 ( .A(n1475), .B(n1476), .Z(n1474) );
  NANDN U1462 ( .A(n1476), .B(n1475), .Z(n1471) );
  ANDN U1463 ( .B(B[77]), .A(n35), .Z(n1366) );
  XNOR U1464 ( .A(n1374), .B(n1477), .Z(n1367) );
  XNOR U1465 ( .A(n1373), .B(n1371), .Z(n1477) );
  AND U1466 ( .A(n1478), .B(n1479), .Z(n1371) );
  NANDN U1467 ( .A(n1480), .B(n1481), .Z(n1479) );
  OR U1468 ( .A(n1482), .B(n1483), .Z(n1481) );
  NAND U1469 ( .A(n1483), .B(n1482), .Z(n1478) );
  ANDN U1470 ( .B(B[78]), .A(n36), .Z(n1373) );
  XNOR U1471 ( .A(n1381), .B(n1484), .Z(n1374) );
  XNOR U1472 ( .A(n1380), .B(n1378), .Z(n1484) );
  AND U1473 ( .A(n1485), .B(n1486), .Z(n1378) );
  NANDN U1474 ( .A(n1487), .B(n1488), .Z(n1486) );
  NANDN U1475 ( .A(n1489), .B(n1490), .Z(n1488) );
  NANDN U1476 ( .A(n1490), .B(n1489), .Z(n1485) );
  ANDN U1477 ( .B(B[79]), .A(n37), .Z(n1380) );
  XNOR U1478 ( .A(n1388), .B(n1491), .Z(n1381) );
  XNOR U1479 ( .A(n1387), .B(n1385), .Z(n1491) );
  AND U1480 ( .A(n1492), .B(n1493), .Z(n1385) );
  NANDN U1481 ( .A(n1494), .B(n1495), .Z(n1493) );
  OR U1482 ( .A(n1496), .B(n1497), .Z(n1495) );
  NAND U1483 ( .A(n1497), .B(n1496), .Z(n1492) );
  ANDN U1484 ( .B(B[80]), .A(n38), .Z(n1387) );
  XNOR U1485 ( .A(n1395), .B(n1498), .Z(n1388) );
  XNOR U1486 ( .A(n1394), .B(n1392), .Z(n1498) );
  AND U1487 ( .A(n1499), .B(n1500), .Z(n1392) );
  NANDN U1488 ( .A(n1501), .B(n1502), .Z(n1500) );
  NANDN U1489 ( .A(n1503), .B(n1504), .Z(n1502) );
  NANDN U1490 ( .A(n1504), .B(n1503), .Z(n1499) );
  ANDN U1491 ( .B(B[81]), .A(n39), .Z(n1394) );
  XNOR U1492 ( .A(n1402), .B(n1505), .Z(n1395) );
  XNOR U1493 ( .A(n1401), .B(n1399), .Z(n1505) );
  AND U1494 ( .A(n1506), .B(n1507), .Z(n1399) );
  NANDN U1495 ( .A(n1508), .B(n1509), .Z(n1507) );
  OR U1496 ( .A(n1510), .B(n1511), .Z(n1509) );
  NAND U1497 ( .A(n1511), .B(n1510), .Z(n1506) );
  ANDN U1498 ( .B(B[82]), .A(n40), .Z(n1401) );
  XNOR U1499 ( .A(n1409), .B(n1512), .Z(n1402) );
  XNOR U1500 ( .A(n1408), .B(n1406), .Z(n1512) );
  AND U1501 ( .A(n1513), .B(n1514), .Z(n1406) );
  NANDN U1502 ( .A(n1515), .B(n1516), .Z(n1514) );
  NAND U1503 ( .A(n1517), .B(n1518), .Z(n1516) );
  ANDN U1504 ( .B(B[83]), .A(n41), .Z(n1408) );
  XOR U1505 ( .A(n1415), .B(n1519), .Z(n1409) );
  XNOR U1506 ( .A(n1413), .B(n1416), .Z(n1519) );
  NAND U1507 ( .A(B[84]), .B(A[2]), .Z(n1416) );
  NAND U1508 ( .A(B[85]), .B(n1520), .Z(n1413) );
  ANDN U1509 ( .B(A[0]), .A(n1521), .Z(n1520) );
  XNOR U1510 ( .A(n1419), .B(n1522), .Z(n1415) );
  NAND U1511 ( .A(A[0]), .B(B[86]), .Z(n1522) );
  NAND U1512 ( .A(B[85]), .B(A[1]), .Z(n1419) );
  NAND U1513 ( .A(n1523), .B(n1524), .Z(n74) );
  NANDN U1514 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1515 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1516 ( .A(n1528), .B(n1527), .Z(n1523) );
  XOR U1517 ( .A(n76), .B(n75), .Z(\A1[83] ) );
  XOR U1518 ( .A(n1528), .B(n1529), .Z(n75) );
  XNOR U1519 ( .A(n1527), .B(n1525), .Z(n1529) );
  AND U1520 ( .A(n1530), .B(n1531), .Z(n1525) );
  NANDN U1521 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1522 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1523 ( .A(n1535), .B(n1534), .Z(n1530) );
  ANDN U1524 ( .B(B[70]), .A(n29), .Z(n1527) );
  XNOR U1525 ( .A(n1434), .B(n1536), .Z(n1528) );
  XNOR U1526 ( .A(n1433), .B(n1431), .Z(n1536) );
  AND U1527 ( .A(n1537), .B(n1538), .Z(n1431) );
  NANDN U1528 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1529 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1530 ( .A(n1542), .B(n1541), .Z(n1537) );
  ANDN U1531 ( .B(B[71]), .A(n30), .Z(n1433) );
  XNOR U1532 ( .A(n1441), .B(n1543), .Z(n1434) );
  XNOR U1533 ( .A(n1440), .B(n1438), .Z(n1543) );
  AND U1534 ( .A(n1544), .B(n1545), .Z(n1438) );
  NANDN U1535 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1536 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1537 ( .A(n1549), .B(n1548), .Z(n1544) );
  ANDN U1538 ( .B(B[72]), .A(n31), .Z(n1440) );
  XNOR U1539 ( .A(n1448), .B(n1550), .Z(n1441) );
  XNOR U1540 ( .A(n1447), .B(n1445), .Z(n1550) );
  AND U1541 ( .A(n1551), .B(n1552), .Z(n1445) );
  NANDN U1542 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1543 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1544 ( .A(n1556), .B(n1555), .Z(n1551) );
  ANDN U1545 ( .B(B[73]), .A(n32), .Z(n1447) );
  XNOR U1546 ( .A(n1455), .B(n1557), .Z(n1448) );
  XNOR U1547 ( .A(n1454), .B(n1452), .Z(n1557) );
  AND U1548 ( .A(n1558), .B(n1559), .Z(n1452) );
  NANDN U1549 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1550 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1551 ( .A(n1563), .B(n1562), .Z(n1558) );
  ANDN U1552 ( .B(B[74]), .A(n33), .Z(n1454) );
  XNOR U1553 ( .A(n1462), .B(n1564), .Z(n1455) );
  XNOR U1554 ( .A(n1461), .B(n1459), .Z(n1564) );
  AND U1555 ( .A(n1565), .B(n1566), .Z(n1459) );
  NANDN U1556 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1557 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1558 ( .A(n1570), .B(n1569), .Z(n1565) );
  ANDN U1559 ( .B(B[75]), .A(n34), .Z(n1461) );
  XNOR U1560 ( .A(n1469), .B(n1571), .Z(n1462) );
  XNOR U1561 ( .A(n1468), .B(n1466), .Z(n1571) );
  AND U1562 ( .A(n1572), .B(n1573), .Z(n1466) );
  NANDN U1563 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1564 ( .A(n1576), .B(n1577), .Z(n1575) );
  NANDN U1565 ( .A(n1577), .B(n1576), .Z(n1572) );
  ANDN U1566 ( .B(B[76]), .A(n35), .Z(n1468) );
  XNOR U1567 ( .A(n1476), .B(n1578), .Z(n1469) );
  XNOR U1568 ( .A(n1475), .B(n1473), .Z(n1578) );
  AND U1569 ( .A(n1579), .B(n1580), .Z(n1473) );
  NANDN U1570 ( .A(n1581), .B(n1582), .Z(n1580) );
  OR U1571 ( .A(n1583), .B(n1584), .Z(n1582) );
  NAND U1572 ( .A(n1584), .B(n1583), .Z(n1579) );
  ANDN U1573 ( .B(B[77]), .A(n36), .Z(n1475) );
  XNOR U1574 ( .A(n1483), .B(n1585), .Z(n1476) );
  XNOR U1575 ( .A(n1482), .B(n1480), .Z(n1585) );
  AND U1576 ( .A(n1586), .B(n1587), .Z(n1480) );
  NANDN U1577 ( .A(n1588), .B(n1589), .Z(n1587) );
  NANDN U1578 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1579 ( .A(n1591), .B(n1590), .Z(n1586) );
  ANDN U1580 ( .B(B[78]), .A(n37), .Z(n1482) );
  XNOR U1581 ( .A(n1490), .B(n1592), .Z(n1483) );
  XNOR U1582 ( .A(n1489), .B(n1487), .Z(n1592) );
  AND U1583 ( .A(n1593), .B(n1594), .Z(n1487) );
  NANDN U1584 ( .A(n1595), .B(n1596), .Z(n1594) );
  OR U1585 ( .A(n1597), .B(n1598), .Z(n1596) );
  NAND U1586 ( .A(n1598), .B(n1597), .Z(n1593) );
  ANDN U1587 ( .B(B[79]), .A(n38), .Z(n1489) );
  XNOR U1588 ( .A(n1497), .B(n1599), .Z(n1490) );
  XNOR U1589 ( .A(n1496), .B(n1494), .Z(n1599) );
  AND U1590 ( .A(n1600), .B(n1601), .Z(n1494) );
  NANDN U1591 ( .A(n1602), .B(n1603), .Z(n1601) );
  NANDN U1592 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1593 ( .A(n1605), .B(n1604), .Z(n1600) );
  ANDN U1594 ( .B(B[80]), .A(n39), .Z(n1496) );
  XNOR U1595 ( .A(n1504), .B(n1606), .Z(n1497) );
  XNOR U1596 ( .A(n1503), .B(n1501), .Z(n1606) );
  AND U1597 ( .A(n1607), .B(n1608), .Z(n1501) );
  NANDN U1598 ( .A(n1609), .B(n1610), .Z(n1608) );
  OR U1599 ( .A(n1611), .B(n1612), .Z(n1610) );
  NAND U1600 ( .A(n1612), .B(n1611), .Z(n1607) );
  ANDN U1601 ( .B(B[81]), .A(n40), .Z(n1503) );
  XNOR U1602 ( .A(n1511), .B(n1613), .Z(n1504) );
  XNOR U1603 ( .A(n1510), .B(n1508), .Z(n1613) );
  AND U1604 ( .A(n1614), .B(n1615), .Z(n1508) );
  NANDN U1605 ( .A(n1616), .B(n1617), .Z(n1615) );
  NAND U1606 ( .A(n1618), .B(n1619), .Z(n1617) );
  ANDN U1607 ( .B(B[82]), .A(n41), .Z(n1510) );
  XOR U1608 ( .A(n1517), .B(n1620), .Z(n1511) );
  XNOR U1609 ( .A(n1515), .B(n1518), .Z(n1620) );
  NAND U1610 ( .A(A[2]), .B(B[83]), .Z(n1518) );
  NANDN U1611 ( .A(n1621), .B(n1622), .Z(n1515) );
  AND U1612 ( .A(A[0]), .B(B[84]), .Z(n1622) );
  XNOR U1613 ( .A(n1521), .B(n1623), .Z(n1517) );
  NAND U1614 ( .A(B[85]), .B(A[0]), .Z(n1623) );
  NAND U1615 ( .A(B[84]), .B(A[1]), .Z(n1521) );
  NAND U1616 ( .A(n1624), .B(n1625), .Z(n76) );
  NANDN U1617 ( .A(n1626), .B(n1627), .Z(n1625) );
  OR U1618 ( .A(n1628), .B(n1629), .Z(n1627) );
  NAND U1619 ( .A(n1629), .B(n1628), .Z(n1624) );
  XOR U1620 ( .A(n78), .B(n77), .Z(\A1[82] ) );
  XOR U1621 ( .A(n1629), .B(n1630), .Z(n77) );
  XNOR U1622 ( .A(n1628), .B(n1626), .Z(n1630) );
  AND U1623 ( .A(n1631), .B(n1632), .Z(n1626) );
  NANDN U1624 ( .A(n1633), .B(n1634), .Z(n1632) );
  NANDN U1625 ( .A(n1635), .B(n1636), .Z(n1634) );
  NANDN U1626 ( .A(n1636), .B(n1635), .Z(n1631) );
  ANDN U1627 ( .B(B[69]), .A(n29), .Z(n1628) );
  XNOR U1628 ( .A(n1535), .B(n1637), .Z(n1629) );
  XNOR U1629 ( .A(n1534), .B(n1532), .Z(n1637) );
  AND U1630 ( .A(n1638), .B(n1639), .Z(n1532) );
  NANDN U1631 ( .A(n1640), .B(n1641), .Z(n1639) );
  OR U1632 ( .A(n1642), .B(n1643), .Z(n1641) );
  NAND U1633 ( .A(n1643), .B(n1642), .Z(n1638) );
  ANDN U1634 ( .B(B[70]), .A(n30), .Z(n1534) );
  XNOR U1635 ( .A(n1542), .B(n1644), .Z(n1535) );
  XNOR U1636 ( .A(n1541), .B(n1539), .Z(n1644) );
  AND U1637 ( .A(n1645), .B(n1646), .Z(n1539) );
  NANDN U1638 ( .A(n1647), .B(n1648), .Z(n1646) );
  NANDN U1639 ( .A(n1649), .B(n1650), .Z(n1648) );
  NANDN U1640 ( .A(n1650), .B(n1649), .Z(n1645) );
  ANDN U1641 ( .B(B[71]), .A(n31), .Z(n1541) );
  XNOR U1642 ( .A(n1549), .B(n1651), .Z(n1542) );
  XNOR U1643 ( .A(n1548), .B(n1546), .Z(n1651) );
  AND U1644 ( .A(n1652), .B(n1653), .Z(n1546) );
  NANDN U1645 ( .A(n1654), .B(n1655), .Z(n1653) );
  OR U1646 ( .A(n1656), .B(n1657), .Z(n1655) );
  NAND U1647 ( .A(n1657), .B(n1656), .Z(n1652) );
  ANDN U1648 ( .B(B[72]), .A(n32), .Z(n1548) );
  XNOR U1649 ( .A(n1556), .B(n1658), .Z(n1549) );
  XNOR U1650 ( .A(n1555), .B(n1553), .Z(n1658) );
  AND U1651 ( .A(n1659), .B(n1660), .Z(n1553) );
  NANDN U1652 ( .A(n1661), .B(n1662), .Z(n1660) );
  NANDN U1653 ( .A(n1663), .B(n1664), .Z(n1662) );
  NANDN U1654 ( .A(n1664), .B(n1663), .Z(n1659) );
  ANDN U1655 ( .B(B[73]), .A(n33), .Z(n1555) );
  XNOR U1656 ( .A(n1563), .B(n1665), .Z(n1556) );
  XNOR U1657 ( .A(n1562), .B(n1560), .Z(n1665) );
  AND U1658 ( .A(n1666), .B(n1667), .Z(n1560) );
  NANDN U1659 ( .A(n1668), .B(n1669), .Z(n1667) );
  OR U1660 ( .A(n1670), .B(n1671), .Z(n1669) );
  NAND U1661 ( .A(n1671), .B(n1670), .Z(n1666) );
  ANDN U1662 ( .B(B[74]), .A(n34), .Z(n1562) );
  XNOR U1663 ( .A(n1570), .B(n1672), .Z(n1563) );
  XNOR U1664 ( .A(n1569), .B(n1567), .Z(n1672) );
  AND U1665 ( .A(n1673), .B(n1674), .Z(n1567) );
  NANDN U1666 ( .A(n1675), .B(n1676), .Z(n1674) );
  NANDN U1667 ( .A(n1677), .B(n1678), .Z(n1676) );
  NANDN U1668 ( .A(n1678), .B(n1677), .Z(n1673) );
  ANDN U1669 ( .B(B[75]), .A(n35), .Z(n1569) );
  XNOR U1670 ( .A(n1577), .B(n1679), .Z(n1570) );
  XNOR U1671 ( .A(n1576), .B(n1574), .Z(n1679) );
  AND U1672 ( .A(n1680), .B(n1681), .Z(n1574) );
  NANDN U1673 ( .A(n1682), .B(n1683), .Z(n1681) );
  OR U1674 ( .A(n1684), .B(n1685), .Z(n1683) );
  NAND U1675 ( .A(n1685), .B(n1684), .Z(n1680) );
  ANDN U1676 ( .B(B[76]), .A(n36), .Z(n1576) );
  XNOR U1677 ( .A(n1584), .B(n1686), .Z(n1577) );
  XNOR U1678 ( .A(n1583), .B(n1581), .Z(n1686) );
  AND U1679 ( .A(n1687), .B(n1688), .Z(n1581) );
  NANDN U1680 ( .A(n1689), .B(n1690), .Z(n1688) );
  NANDN U1681 ( .A(n1691), .B(n1692), .Z(n1690) );
  NANDN U1682 ( .A(n1692), .B(n1691), .Z(n1687) );
  ANDN U1683 ( .B(B[77]), .A(n37), .Z(n1583) );
  XNOR U1684 ( .A(n1591), .B(n1693), .Z(n1584) );
  XNOR U1685 ( .A(n1590), .B(n1588), .Z(n1693) );
  AND U1686 ( .A(n1694), .B(n1695), .Z(n1588) );
  NANDN U1687 ( .A(n1696), .B(n1697), .Z(n1695) );
  OR U1688 ( .A(n1698), .B(n1699), .Z(n1697) );
  NAND U1689 ( .A(n1699), .B(n1698), .Z(n1694) );
  ANDN U1690 ( .B(B[78]), .A(n38), .Z(n1590) );
  XNOR U1691 ( .A(n1598), .B(n1700), .Z(n1591) );
  XNOR U1692 ( .A(n1597), .B(n1595), .Z(n1700) );
  AND U1693 ( .A(n1701), .B(n1702), .Z(n1595) );
  NANDN U1694 ( .A(n1703), .B(n1704), .Z(n1702) );
  NANDN U1695 ( .A(n1705), .B(n1706), .Z(n1704) );
  NANDN U1696 ( .A(n1706), .B(n1705), .Z(n1701) );
  ANDN U1697 ( .B(B[79]), .A(n39), .Z(n1597) );
  XNOR U1698 ( .A(n1605), .B(n1707), .Z(n1598) );
  XNOR U1699 ( .A(n1604), .B(n1602), .Z(n1707) );
  AND U1700 ( .A(n1708), .B(n1709), .Z(n1602) );
  NANDN U1701 ( .A(n1710), .B(n1711), .Z(n1709) );
  OR U1702 ( .A(n1712), .B(n1713), .Z(n1711) );
  NAND U1703 ( .A(n1713), .B(n1712), .Z(n1708) );
  ANDN U1704 ( .B(B[80]), .A(n40), .Z(n1604) );
  XNOR U1705 ( .A(n1612), .B(n1714), .Z(n1605) );
  XNOR U1706 ( .A(n1611), .B(n1609), .Z(n1714) );
  AND U1707 ( .A(n1715), .B(n1716), .Z(n1609) );
  NANDN U1708 ( .A(n1717), .B(n1718), .Z(n1716) );
  NAND U1709 ( .A(n1719), .B(n1720), .Z(n1718) );
  ANDN U1710 ( .B(B[81]), .A(n41), .Z(n1611) );
  XOR U1711 ( .A(n1618), .B(n1721), .Z(n1612) );
  XNOR U1712 ( .A(n1616), .B(n1619), .Z(n1721) );
  NAND U1713 ( .A(A[2]), .B(B[82]), .Z(n1619) );
  NANDN U1714 ( .A(n1722), .B(n1723), .Z(n1616) );
  AND U1715 ( .A(A[0]), .B(B[83]), .Z(n1723) );
  XNOR U1716 ( .A(n1621), .B(n1724), .Z(n1618) );
  NAND U1717 ( .A(A[0]), .B(B[84]), .Z(n1724) );
  NAND U1718 ( .A(B[83]), .B(A[1]), .Z(n1621) );
  NAND U1719 ( .A(n1725), .B(n1726), .Z(n78) );
  NANDN U1720 ( .A(n1727), .B(n1728), .Z(n1726) );
  OR U1721 ( .A(n1729), .B(n1730), .Z(n1728) );
  NAND U1722 ( .A(n1730), .B(n1729), .Z(n1725) );
  XOR U1723 ( .A(n80), .B(n79), .Z(\A1[81] ) );
  XOR U1724 ( .A(n1730), .B(n1731), .Z(n79) );
  XNOR U1725 ( .A(n1729), .B(n1727), .Z(n1731) );
  AND U1726 ( .A(n1732), .B(n1733), .Z(n1727) );
  NANDN U1727 ( .A(n1734), .B(n1735), .Z(n1733) );
  NANDN U1728 ( .A(n1736), .B(n1737), .Z(n1735) );
  NANDN U1729 ( .A(n1737), .B(n1736), .Z(n1732) );
  ANDN U1730 ( .B(B[68]), .A(n29), .Z(n1729) );
  XNOR U1731 ( .A(n1636), .B(n1738), .Z(n1730) );
  XNOR U1732 ( .A(n1635), .B(n1633), .Z(n1738) );
  AND U1733 ( .A(n1739), .B(n1740), .Z(n1633) );
  NANDN U1734 ( .A(n1741), .B(n1742), .Z(n1740) );
  OR U1735 ( .A(n1743), .B(n1744), .Z(n1742) );
  NAND U1736 ( .A(n1744), .B(n1743), .Z(n1739) );
  ANDN U1737 ( .B(B[69]), .A(n30), .Z(n1635) );
  XNOR U1738 ( .A(n1643), .B(n1745), .Z(n1636) );
  XNOR U1739 ( .A(n1642), .B(n1640), .Z(n1745) );
  AND U1740 ( .A(n1746), .B(n1747), .Z(n1640) );
  NANDN U1741 ( .A(n1748), .B(n1749), .Z(n1747) );
  NANDN U1742 ( .A(n1750), .B(n1751), .Z(n1749) );
  NANDN U1743 ( .A(n1751), .B(n1750), .Z(n1746) );
  ANDN U1744 ( .B(B[70]), .A(n31), .Z(n1642) );
  XNOR U1745 ( .A(n1650), .B(n1752), .Z(n1643) );
  XNOR U1746 ( .A(n1649), .B(n1647), .Z(n1752) );
  AND U1747 ( .A(n1753), .B(n1754), .Z(n1647) );
  NANDN U1748 ( .A(n1755), .B(n1756), .Z(n1754) );
  OR U1749 ( .A(n1757), .B(n1758), .Z(n1756) );
  NAND U1750 ( .A(n1758), .B(n1757), .Z(n1753) );
  ANDN U1751 ( .B(B[71]), .A(n32), .Z(n1649) );
  XNOR U1752 ( .A(n1657), .B(n1759), .Z(n1650) );
  XNOR U1753 ( .A(n1656), .B(n1654), .Z(n1759) );
  AND U1754 ( .A(n1760), .B(n1761), .Z(n1654) );
  NANDN U1755 ( .A(n1762), .B(n1763), .Z(n1761) );
  NANDN U1756 ( .A(n1764), .B(n1765), .Z(n1763) );
  NANDN U1757 ( .A(n1765), .B(n1764), .Z(n1760) );
  ANDN U1758 ( .B(B[72]), .A(n33), .Z(n1656) );
  XNOR U1759 ( .A(n1664), .B(n1766), .Z(n1657) );
  XNOR U1760 ( .A(n1663), .B(n1661), .Z(n1766) );
  AND U1761 ( .A(n1767), .B(n1768), .Z(n1661) );
  NANDN U1762 ( .A(n1769), .B(n1770), .Z(n1768) );
  OR U1763 ( .A(n1771), .B(n1772), .Z(n1770) );
  NAND U1764 ( .A(n1772), .B(n1771), .Z(n1767) );
  ANDN U1765 ( .B(B[73]), .A(n34), .Z(n1663) );
  XNOR U1766 ( .A(n1671), .B(n1773), .Z(n1664) );
  XNOR U1767 ( .A(n1670), .B(n1668), .Z(n1773) );
  AND U1768 ( .A(n1774), .B(n1775), .Z(n1668) );
  NANDN U1769 ( .A(n1776), .B(n1777), .Z(n1775) );
  NANDN U1770 ( .A(n1778), .B(n1779), .Z(n1777) );
  NANDN U1771 ( .A(n1779), .B(n1778), .Z(n1774) );
  ANDN U1772 ( .B(B[74]), .A(n35), .Z(n1670) );
  XNOR U1773 ( .A(n1678), .B(n1780), .Z(n1671) );
  XNOR U1774 ( .A(n1677), .B(n1675), .Z(n1780) );
  AND U1775 ( .A(n1781), .B(n1782), .Z(n1675) );
  NANDN U1776 ( .A(n1783), .B(n1784), .Z(n1782) );
  OR U1777 ( .A(n1785), .B(n1786), .Z(n1784) );
  NAND U1778 ( .A(n1786), .B(n1785), .Z(n1781) );
  ANDN U1779 ( .B(B[75]), .A(n36), .Z(n1677) );
  XNOR U1780 ( .A(n1685), .B(n1787), .Z(n1678) );
  XNOR U1781 ( .A(n1684), .B(n1682), .Z(n1787) );
  AND U1782 ( .A(n1788), .B(n1789), .Z(n1682) );
  NANDN U1783 ( .A(n1790), .B(n1791), .Z(n1789) );
  NANDN U1784 ( .A(n1792), .B(n1793), .Z(n1791) );
  NANDN U1785 ( .A(n1793), .B(n1792), .Z(n1788) );
  ANDN U1786 ( .B(B[76]), .A(n37), .Z(n1684) );
  XNOR U1787 ( .A(n1692), .B(n1794), .Z(n1685) );
  XNOR U1788 ( .A(n1691), .B(n1689), .Z(n1794) );
  AND U1789 ( .A(n1795), .B(n1796), .Z(n1689) );
  NANDN U1790 ( .A(n1797), .B(n1798), .Z(n1796) );
  OR U1791 ( .A(n1799), .B(n1800), .Z(n1798) );
  NAND U1792 ( .A(n1800), .B(n1799), .Z(n1795) );
  ANDN U1793 ( .B(B[77]), .A(n38), .Z(n1691) );
  XNOR U1794 ( .A(n1699), .B(n1801), .Z(n1692) );
  XNOR U1795 ( .A(n1698), .B(n1696), .Z(n1801) );
  AND U1796 ( .A(n1802), .B(n1803), .Z(n1696) );
  NANDN U1797 ( .A(n1804), .B(n1805), .Z(n1803) );
  NANDN U1798 ( .A(n1806), .B(n1807), .Z(n1805) );
  NANDN U1799 ( .A(n1807), .B(n1806), .Z(n1802) );
  ANDN U1800 ( .B(B[78]), .A(n39), .Z(n1698) );
  XNOR U1801 ( .A(n1706), .B(n1808), .Z(n1699) );
  XNOR U1802 ( .A(n1705), .B(n1703), .Z(n1808) );
  AND U1803 ( .A(n1809), .B(n1810), .Z(n1703) );
  NANDN U1804 ( .A(n1811), .B(n1812), .Z(n1810) );
  OR U1805 ( .A(n1813), .B(n1814), .Z(n1812) );
  NAND U1806 ( .A(n1814), .B(n1813), .Z(n1809) );
  ANDN U1807 ( .B(B[79]), .A(n40), .Z(n1705) );
  XNOR U1808 ( .A(n1713), .B(n1815), .Z(n1706) );
  XNOR U1809 ( .A(n1712), .B(n1710), .Z(n1815) );
  AND U1810 ( .A(n1816), .B(n1817), .Z(n1710) );
  NANDN U1811 ( .A(n1818), .B(n1819), .Z(n1817) );
  NAND U1812 ( .A(n1820), .B(n1821), .Z(n1819) );
  ANDN U1813 ( .B(B[80]), .A(n41), .Z(n1712) );
  XOR U1814 ( .A(n1719), .B(n1822), .Z(n1713) );
  XNOR U1815 ( .A(n1717), .B(n1720), .Z(n1822) );
  NAND U1816 ( .A(A[2]), .B(B[81]), .Z(n1720) );
  NANDN U1817 ( .A(n1823), .B(n1824), .Z(n1717) );
  AND U1818 ( .A(A[0]), .B(B[82]), .Z(n1824) );
  XNOR U1819 ( .A(n1722), .B(n1825), .Z(n1719) );
  NAND U1820 ( .A(A[0]), .B(B[83]), .Z(n1825) );
  NAND U1821 ( .A(B[82]), .B(A[1]), .Z(n1722) );
  NAND U1822 ( .A(n1826), .B(n1827), .Z(n80) );
  NANDN U1823 ( .A(n1828), .B(n1829), .Z(n1827) );
  OR U1824 ( .A(n1830), .B(n1831), .Z(n1829) );
  NAND U1825 ( .A(n1831), .B(n1830), .Z(n1826) );
  XOR U1826 ( .A(n82), .B(n81), .Z(\A1[80] ) );
  XOR U1827 ( .A(n1831), .B(n1832), .Z(n81) );
  XNOR U1828 ( .A(n1830), .B(n1828), .Z(n1832) );
  AND U1829 ( .A(n1833), .B(n1834), .Z(n1828) );
  NANDN U1830 ( .A(n1835), .B(n1836), .Z(n1834) );
  NANDN U1831 ( .A(n1837), .B(n1838), .Z(n1836) );
  NANDN U1832 ( .A(n1838), .B(n1837), .Z(n1833) );
  ANDN U1833 ( .B(B[67]), .A(n29), .Z(n1830) );
  XNOR U1834 ( .A(n1737), .B(n1839), .Z(n1831) );
  XNOR U1835 ( .A(n1736), .B(n1734), .Z(n1839) );
  AND U1836 ( .A(n1840), .B(n1841), .Z(n1734) );
  NANDN U1837 ( .A(n1842), .B(n1843), .Z(n1841) );
  OR U1838 ( .A(n1844), .B(n1845), .Z(n1843) );
  NAND U1839 ( .A(n1845), .B(n1844), .Z(n1840) );
  ANDN U1840 ( .B(B[68]), .A(n30), .Z(n1736) );
  XNOR U1841 ( .A(n1744), .B(n1846), .Z(n1737) );
  XNOR U1842 ( .A(n1743), .B(n1741), .Z(n1846) );
  AND U1843 ( .A(n1847), .B(n1848), .Z(n1741) );
  NANDN U1844 ( .A(n1849), .B(n1850), .Z(n1848) );
  NANDN U1845 ( .A(n1851), .B(n1852), .Z(n1850) );
  NANDN U1846 ( .A(n1852), .B(n1851), .Z(n1847) );
  ANDN U1847 ( .B(B[69]), .A(n31), .Z(n1743) );
  XNOR U1848 ( .A(n1751), .B(n1853), .Z(n1744) );
  XNOR U1849 ( .A(n1750), .B(n1748), .Z(n1853) );
  AND U1850 ( .A(n1854), .B(n1855), .Z(n1748) );
  NANDN U1851 ( .A(n1856), .B(n1857), .Z(n1855) );
  OR U1852 ( .A(n1858), .B(n1859), .Z(n1857) );
  NAND U1853 ( .A(n1859), .B(n1858), .Z(n1854) );
  ANDN U1854 ( .B(B[70]), .A(n32), .Z(n1750) );
  XNOR U1855 ( .A(n1758), .B(n1860), .Z(n1751) );
  XNOR U1856 ( .A(n1757), .B(n1755), .Z(n1860) );
  AND U1857 ( .A(n1861), .B(n1862), .Z(n1755) );
  NANDN U1858 ( .A(n1863), .B(n1864), .Z(n1862) );
  NANDN U1859 ( .A(n1865), .B(n1866), .Z(n1864) );
  NANDN U1860 ( .A(n1866), .B(n1865), .Z(n1861) );
  ANDN U1861 ( .B(B[71]), .A(n33), .Z(n1757) );
  XNOR U1862 ( .A(n1765), .B(n1867), .Z(n1758) );
  XNOR U1863 ( .A(n1764), .B(n1762), .Z(n1867) );
  AND U1864 ( .A(n1868), .B(n1869), .Z(n1762) );
  NANDN U1865 ( .A(n1870), .B(n1871), .Z(n1869) );
  OR U1866 ( .A(n1872), .B(n1873), .Z(n1871) );
  NAND U1867 ( .A(n1873), .B(n1872), .Z(n1868) );
  ANDN U1868 ( .B(B[72]), .A(n34), .Z(n1764) );
  XNOR U1869 ( .A(n1772), .B(n1874), .Z(n1765) );
  XNOR U1870 ( .A(n1771), .B(n1769), .Z(n1874) );
  AND U1871 ( .A(n1875), .B(n1876), .Z(n1769) );
  NANDN U1872 ( .A(n1877), .B(n1878), .Z(n1876) );
  NANDN U1873 ( .A(n1879), .B(n1880), .Z(n1878) );
  NANDN U1874 ( .A(n1880), .B(n1879), .Z(n1875) );
  ANDN U1875 ( .B(B[73]), .A(n35), .Z(n1771) );
  XNOR U1876 ( .A(n1779), .B(n1881), .Z(n1772) );
  XNOR U1877 ( .A(n1778), .B(n1776), .Z(n1881) );
  AND U1878 ( .A(n1882), .B(n1883), .Z(n1776) );
  NANDN U1879 ( .A(n1884), .B(n1885), .Z(n1883) );
  OR U1880 ( .A(n1886), .B(n1887), .Z(n1885) );
  NAND U1881 ( .A(n1887), .B(n1886), .Z(n1882) );
  ANDN U1882 ( .B(B[74]), .A(n36), .Z(n1778) );
  XNOR U1883 ( .A(n1786), .B(n1888), .Z(n1779) );
  XNOR U1884 ( .A(n1785), .B(n1783), .Z(n1888) );
  AND U1885 ( .A(n1889), .B(n1890), .Z(n1783) );
  NANDN U1886 ( .A(n1891), .B(n1892), .Z(n1890) );
  NANDN U1887 ( .A(n1893), .B(n1894), .Z(n1892) );
  NANDN U1888 ( .A(n1894), .B(n1893), .Z(n1889) );
  ANDN U1889 ( .B(B[75]), .A(n37), .Z(n1785) );
  XNOR U1890 ( .A(n1793), .B(n1895), .Z(n1786) );
  XNOR U1891 ( .A(n1792), .B(n1790), .Z(n1895) );
  AND U1892 ( .A(n1896), .B(n1897), .Z(n1790) );
  NANDN U1893 ( .A(n1898), .B(n1899), .Z(n1897) );
  OR U1894 ( .A(n1900), .B(n1901), .Z(n1899) );
  NAND U1895 ( .A(n1901), .B(n1900), .Z(n1896) );
  ANDN U1896 ( .B(B[76]), .A(n38), .Z(n1792) );
  XNOR U1897 ( .A(n1800), .B(n1902), .Z(n1793) );
  XNOR U1898 ( .A(n1799), .B(n1797), .Z(n1902) );
  AND U1899 ( .A(n1903), .B(n1904), .Z(n1797) );
  NANDN U1900 ( .A(n1905), .B(n1906), .Z(n1904) );
  NANDN U1901 ( .A(n1907), .B(n1908), .Z(n1906) );
  NANDN U1902 ( .A(n1908), .B(n1907), .Z(n1903) );
  ANDN U1903 ( .B(B[77]), .A(n39), .Z(n1799) );
  XNOR U1904 ( .A(n1807), .B(n1909), .Z(n1800) );
  XNOR U1905 ( .A(n1806), .B(n1804), .Z(n1909) );
  AND U1906 ( .A(n1910), .B(n1911), .Z(n1804) );
  NANDN U1907 ( .A(n1912), .B(n1913), .Z(n1911) );
  OR U1908 ( .A(n1914), .B(n1915), .Z(n1913) );
  NAND U1909 ( .A(n1915), .B(n1914), .Z(n1910) );
  ANDN U1910 ( .B(B[78]), .A(n40), .Z(n1806) );
  XNOR U1911 ( .A(n1814), .B(n1916), .Z(n1807) );
  XNOR U1912 ( .A(n1813), .B(n1811), .Z(n1916) );
  AND U1913 ( .A(n1917), .B(n1918), .Z(n1811) );
  NANDN U1914 ( .A(n1919), .B(n1920), .Z(n1918) );
  NAND U1915 ( .A(n1921), .B(n1922), .Z(n1920) );
  ANDN U1916 ( .B(B[79]), .A(n41), .Z(n1813) );
  XOR U1917 ( .A(n1820), .B(n1923), .Z(n1814) );
  XNOR U1918 ( .A(n1818), .B(n1821), .Z(n1923) );
  NAND U1919 ( .A(A[2]), .B(B[80]), .Z(n1821) );
  NANDN U1920 ( .A(n1924), .B(n1925), .Z(n1818) );
  AND U1921 ( .A(A[0]), .B(B[81]), .Z(n1925) );
  XNOR U1922 ( .A(n1823), .B(n1926), .Z(n1820) );
  NAND U1923 ( .A(A[0]), .B(B[82]), .Z(n1926) );
  NAND U1924 ( .A(B[81]), .B(A[1]), .Z(n1823) );
  NAND U1925 ( .A(n1927), .B(n1928), .Z(n82) );
  NANDN U1926 ( .A(n1929), .B(n1930), .Z(n1928) );
  OR U1927 ( .A(n1931), .B(n1932), .Z(n1930) );
  NAND U1928 ( .A(n1932), .B(n1931), .Z(n1927) );
  XOR U1929 ( .A(n1933), .B(n1934), .Z(\A1[7] ) );
  XNOR U1930 ( .A(n1935), .B(n25), .Z(n1934) );
  XOR U1931 ( .A(n84), .B(n83), .Z(\A1[79] ) );
  XOR U1932 ( .A(n1932), .B(n1936), .Z(n83) );
  XNOR U1933 ( .A(n1931), .B(n1929), .Z(n1936) );
  AND U1934 ( .A(n1937), .B(n1938), .Z(n1929) );
  NANDN U1935 ( .A(n1939), .B(n1940), .Z(n1938) );
  NANDN U1936 ( .A(n1941), .B(n1942), .Z(n1940) );
  NANDN U1937 ( .A(n1942), .B(n1941), .Z(n1937) );
  ANDN U1938 ( .B(B[66]), .A(n29), .Z(n1931) );
  XNOR U1939 ( .A(n1838), .B(n1943), .Z(n1932) );
  XNOR U1940 ( .A(n1837), .B(n1835), .Z(n1943) );
  AND U1941 ( .A(n1944), .B(n1945), .Z(n1835) );
  NANDN U1942 ( .A(n1946), .B(n1947), .Z(n1945) );
  OR U1943 ( .A(n1948), .B(n1949), .Z(n1947) );
  NAND U1944 ( .A(n1949), .B(n1948), .Z(n1944) );
  ANDN U1945 ( .B(B[67]), .A(n30), .Z(n1837) );
  XNOR U1946 ( .A(n1845), .B(n1950), .Z(n1838) );
  XNOR U1947 ( .A(n1844), .B(n1842), .Z(n1950) );
  AND U1948 ( .A(n1951), .B(n1952), .Z(n1842) );
  NANDN U1949 ( .A(n1953), .B(n1954), .Z(n1952) );
  NANDN U1950 ( .A(n1955), .B(n1956), .Z(n1954) );
  NANDN U1951 ( .A(n1956), .B(n1955), .Z(n1951) );
  ANDN U1952 ( .B(B[68]), .A(n31), .Z(n1844) );
  XNOR U1953 ( .A(n1852), .B(n1957), .Z(n1845) );
  XNOR U1954 ( .A(n1851), .B(n1849), .Z(n1957) );
  AND U1955 ( .A(n1958), .B(n1959), .Z(n1849) );
  NANDN U1956 ( .A(n1960), .B(n1961), .Z(n1959) );
  OR U1957 ( .A(n1962), .B(n1963), .Z(n1961) );
  NAND U1958 ( .A(n1963), .B(n1962), .Z(n1958) );
  ANDN U1959 ( .B(B[69]), .A(n32), .Z(n1851) );
  XNOR U1960 ( .A(n1859), .B(n1964), .Z(n1852) );
  XNOR U1961 ( .A(n1858), .B(n1856), .Z(n1964) );
  AND U1962 ( .A(n1965), .B(n1966), .Z(n1856) );
  NANDN U1963 ( .A(n1967), .B(n1968), .Z(n1966) );
  NANDN U1964 ( .A(n1969), .B(n1970), .Z(n1968) );
  NANDN U1965 ( .A(n1970), .B(n1969), .Z(n1965) );
  ANDN U1966 ( .B(B[70]), .A(n33), .Z(n1858) );
  XNOR U1967 ( .A(n1866), .B(n1971), .Z(n1859) );
  XNOR U1968 ( .A(n1865), .B(n1863), .Z(n1971) );
  AND U1969 ( .A(n1972), .B(n1973), .Z(n1863) );
  NANDN U1970 ( .A(n1974), .B(n1975), .Z(n1973) );
  OR U1971 ( .A(n1976), .B(n1977), .Z(n1975) );
  NAND U1972 ( .A(n1977), .B(n1976), .Z(n1972) );
  ANDN U1973 ( .B(B[71]), .A(n34), .Z(n1865) );
  XNOR U1974 ( .A(n1873), .B(n1978), .Z(n1866) );
  XNOR U1975 ( .A(n1872), .B(n1870), .Z(n1978) );
  AND U1976 ( .A(n1979), .B(n1980), .Z(n1870) );
  NANDN U1977 ( .A(n1981), .B(n1982), .Z(n1980) );
  NANDN U1978 ( .A(n1983), .B(n1984), .Z(n1982) );
  NANDN U1979 ( .A(n1984), .B(n1983), .Z(n1979) );
  ANDN U1980 ( .B(B[72]), .A(n35), .Z(n1872) );
  XNOR U1981 ( .A(n1880), .B(n1985), .Z(n1873) );
  XNOR U1982 ( .A(n1879), .B(n1877), .Z(n1985) );
  AND U1983 ( .A(n1986), .B(n1987), .Z(n1877) );
  NANDN U1984 ( .A(n1988), .B(n1989), .Z(n1987) );
  OR U1985 ( .A(n1990), .B(n1991), .Z(n1989) );
  NAND U1986 ( .A(n1991), .B(n1990), .Z(n1986) );
  ANDN U1987 ( .B(B[73]), .A(n36), .Z(n1879) );
  XNOR U1988 ( .A(n1887), .B(n1992), .Z(n1880) );
  XNOR U1989 ( .A(n1886), .B(n1884), .Z(n1992) );
  AND U1990 ( .A(n1993), .B(n1994), .Z(n1884) );
  NANDN U1991 ( .A(n1995), .B(n1996), .Z(n1994) );
  NANDN U1992 ( .A(n1997), .B(n1998), .Z(n1996) );
  NANDN U1993 ( .A(n1998), .B(n1997), .Z(n1993) );
  ANDN U1994 ( .B(B[74]), .A(n37), .Z(n1886) );
  XNOR U1995 ( .A(n1894), .B(n1999), .Z(n1887) );
  XNOR U1996 ( .A(n1893), .B(n1891), .Z(n1999) );
  AND U1997 ( .A(n2000), .B(n2001), .Z(n1891) );
  NANDN U1998 ( .A(n2002), .B(n2003), .Z(n2001) );
  OR U1999 ( .A(n2004), .B(n2005), .Z(n2003) );
  NAND U2000 ( .A(n2005), .B(n2004), .Z(n2000) );
  ANDN U2001 ( .B(B[75]), .A(n38), .Z(n1893) );
  XNOR U2002 ( .A(n1901), .B(n2006), .Z(n1894) );
  XNOR U2003 ( .A(n1900), .B(n1898), .Z(n2006) );
  AND U2004 ( .A(n2007), .B(n2008), .Z(n1898) );
  NANDN U2005 ( .A(n2009), .B(n2010), .Z(n2008) );
  NANDN U2006 ( .A(n2011), .B(n2012), .Z(n2010) );
  NANDN U2007 ( .A(n2012), .B(n2011), .Z(n2007) );
  ANDN U2008 ( .B(B[76]), .A(n39), .Z(n1900) );
  XNOR U2009 ( .A(n1908), .B(n2013), .Z(n1901) );
  XNOR U2010 ( .A(n1907), .B(n1905), .Z(n2013) );
  AND U2011 ( .A(n2014), .B(n2015), .Z(n1905) );
  NANDN U2012 ( .A(n2016), .B(n2017), .Z(n2015) );
  OR U2013 ( .A(n2018), .B(n2019), .Z(n2017) );
  NAND U2014 ( .A(n2019), .B(n2018), .Z(n2014) );
  ANDN U2015 ( .B(B[77]), .A(n40), .Z(n1907) );
  XNOR U2016 ( .A(n1915), .B(n2020), .Z(n1908) );
  XNOR U2017 ( .A(n1914), .B(n1912), .Z(n2020) );
  AND U2018 ( .A(n2021), .B(n2022), .Z(n1912) );
  NANDN U2019 ( .A(n2023), .B(n2024), .Z(n2022) );
  NAND U2020 ( .A(n2025), .B(n2026), .Z(n2024) );
  ANDN U2021 ( .B(B[78]), .A(n41), .Z(n1914) );
  XOR U2022 ( .A(n1921), .B(n2027), .Z(n1915) );
  XNOR U2023 ( .A(n1919), .B(n1922), .Z(n2027) );
  NAND U2024 ( .A(A[2]), .B(B[79]), .Z(n1922) );
  NANDN U2025 ( .A(n2028), .B(n2029), .Z(n1919) );
  AND U2026 ( .A(A[0]), .B(B[80]), .Z(n2029) );
  XNOR U2027 ( .A(n1924), .B(n2030), .Z(n1921) );
  NAND U2028 ( .A(A[0]), .B(B[81]), .Z(n2030) );
  NAND U2029 ( .A(B[80]), .B(A[1]), .Z(n1924) );
  NAND U2030 ( .A(n2031), .B(n2032), .Z(n84) );
  NANDN U2031 ( .A(n2033), .B(n2034), .Z(n2032) );
  OR U2032 ( .A(n2035), .B(n2036), .Z(n2034) );
  NAND U2033 ( .A(n2036), .B(n2035), .Z(n2031) );
  XOR U2034 ( .A(n86), .B(n85), .Z(\A1[78] ) );
  XOR U2035 ( .A(n2036), .B(n2037), .Z(n85) );
  XNOR U2036 ( .A(n2035), .B(n2033), .Z(n2037) );
  AND U2037 ( .A(n2038), .B(n2039), .Z(n2033) );
  NANDN U2038 ( .A(n2040), .B(n2041), .Z(n2039) );
  NANDN U2039 ( .A(n2042), .B(n2043), .Z(n2041) );
  NANDN U2040 ( .A(n2043), .B(n2042), .Z(n2038) );
  ANDN U2041 ( .B(B[65]), .A(n29), .Z(n2035) );
  XNOR U2042 ( .A(n1942), .B(n2044), .Z(n2036) );
  XNOR U2043 ( .A(n1941), .B(n1939), .Z(n2044) );
  AND U2044 ( .A(n2045), .B(n2046), .Z(n1939) );
  NANDN U2045 ( .A(n2047), .B(n2048), .Z(n2046) );
  OR U2046 ( .A(n2049), .B(n2050), .Z(n2048) );
  NAND U2047 ( .A(n2050), .B(n2049), .Z(n2045) );
  ANDN U2048 ( .B(B[66]), .A(n30), .Z(n1941) );
  XNOR U2049 ( .A(n1949), .B(n2051), .Z(n1942) );
  XNOR U2050 ( .A(n1948), .B(n1946), .Z(n2051) );
  AND U2051 ( .A(n2052), .B(n2053), .Z(n1946) );
  NANDN U2052 ( .A(n2054), .B(n2055), .Z(n2053) );
  NANDN U2053 ( .A(n2056), .B(n2057), .Z(n2055) );
  NANDN U2054 ( .A(n2057), .B(n2056), .Z(n2052) );
  ANDN U2055 ( .B(B[67]), .A(n31), .Z(n1948) );
  XNOR U2056 ( .A(n1956), .B(n2058), .Z(n1949) );
  XNOR U2057 ( .A(n1955), .B(n1953), .Z(n2058) );
  AND U2058 ( .A(n2059), .B(n2060), .Z(n1953) );
  NANDN U2059 ( .A(n2061), .B(n2062), .Z(n2060) );
  OR U2060 ( .A(n2063), .B(n2064), .Z(n2062) );
  NAND U2061 ( .A(n2064), .B(n2063), .Z(n2059) );
  ANDN U2062 ( .B(B[68]), .A(n32), .Z(n1955) );
  XNOR U2063 ( .A(n1963), .B(n2065), .Z(n1956) );
  XNOR U2064 ( .A(n1962), .B(n1960), .Z(n2065) );
  AND U2065 ( .A(n2066), .B(n2067), .Z(n1960) );
  NANDN U2066 ( .A(n2068), .B(n2069), .Z(n2067) );
  NANDN U2067 ( .A(n2070), .B(n2071), .Z(n2069) );
  NANDN U2068 ( .A(n2071), .B(n2070), .Z(n2066) );
  ANDN U2069 ( .B(B[69]), .A(n33), .Z(n1962) );
  XNOR U2070 ( .A(n1970), .B(n2072), .Z(n1963) );
  XNOR U2071 ( .A(n1969), .B(n1967), .Z(n2072) );
  AND U2072 ( .A(n2073), .B(n2074), .Z(n1967) );
  NANDN U2073 ( .A(n2075), .B(n2076), .Z(n2074) );
  OR U2074 ( .A(n2077), .B(n2078), .Z(n2076) );
  NAND U2075 ( .A(n2078), .B(n2077), .Z(n2073) );
  ANDN U2076 ( .B(B[70]), .A(n34), .Z(n1969) );
  XNOR U2077 ( .A(n1977), .B(n2079), .Z(n1970) );
  XNOR U2078 ( .A(n1976), .B(n1974), .Z(n2079) );
  AND U2079 ( .A(n2080), .B(n2081), .Z(n1974) );
  NANDN U2080 ( .A(n2082), .B(n2083), .Z(n2081) );
  NANDN U2081 ( .A(n2084), .B(n2085), .Z(n2083) );
  NANDN U2082 ( .A(n2085), .B(n2084), .Z(n2080) );
  ANDN U2083 ( .B(B[71]), .A(n35), .Z(n1976) );
  XNOR U2084 ( .A(n1984), .B(n2086), .Z(n1977) );
  XNOR U2085 ( .A(n1983), .B(n1981), .Z(n2086) );
  AND U2086 ( .A(n2087), .B(n2088), .Z(n1981) );
  NANDN U2087 ( .A(n2089), .B(n2090), .Z(n2088) );
  OR U2088 ( .A(n2091), .B(n2092), .Z(n2090) );
  NAND U2089 ( .A(n2092), .B(n2091), .Z(n2087) );
  ANDN U2090 ( .B(B[72]), .A(n36), .Z(n1983) );
  XNOR U2091 ( .A(n1991), .B(n2093), .Z(n1984) );
  XNOR U2092 ( .A(n1990), .B(n1988), .Z(n2093) );
  AND U2093 ( .A(n2094), .B(n2095), .Z(n1988) );
  NANDN U2094 ( .A(n2096), .B(n2097), .Z(n2095) );
  NANDN U2095 ( .A(n2098), .B(n2099), .Z(n2097) );
  NANDN U2096 ( .A(n2099), .B(n2098), .Z(n2094) );
  ANDN U2097 ( .B(B[73]), .A(n37), .Z(n1990) );
  XNOR U2098 ( .A(n1998), .B(n2100), .Z(n1991) );
  XNOR U2099 ( .A(n1997), .B(n1995), .Z(n2100) );
  AND U2100 ( .A(n2101), .B(n2102), .Z(n1995) );
  NANDN U2101 ( .A(n2103), .B(n2104), .Z(n2102) );
  OR U2102 ( .A(n2105), .B(n2106), .Z(n2104) );
  NAND U2103 ( .A(n2106), .B(n2105), .Z(n2101) );
  ANDN U2104 ( .B(B[74]), .A(n38), .Z(n1997) );
  XNOR U2105 ( .A(n2005), .B(n2107), .Z(n1998) );
  XNOR U2106 ( .A(n2004), .B(n2002), .Z(n2107) );
  AND U2107 ( .A(n2108), .B(n2109), .Z(n2002) );
  NANDN U2108 ( .A(n2110), .B(n2111), .Z(n2109) );
  NANDN U2109 ( .A(n2112), .B(n2113), .Z(n2111) );
  NANDN U2110 ( .A(n2113), .B(n2112), .Z(n2108) );
  ANDN U2111 ( .B(B[75]), .A(n39), .Z(n2004) );
  XNOR U2112 ( .A(n2012), .B(n2114), .Z(n2005) );
  XNOR U2113 ( .A(n2011), .B(n2009), .Z(n2114) );
  AND U2114 ( .A(n2115), .B(n2116), .Z(n2009) );
  NANDN U2115 ( .A(n2117), .B(n2118), .Z(n2116) );
  OR U2116 ( .A(n2119), .B(n2120), .Z(n2118) );
  NAND U2117 ( .A(n2120), .B(n2119), .Z(n2115) );
  ANDN U2118 ( .B(B[76]), .A(n40), .Z(n2011) );
  XNOR U2119 ( .A(n2019), .B(n2121), .Z(n2012) );
  XNOR U2120 ( .A(n2018), .B(n2016), .Z(n2121) );
  AND U2121 ( .A(n2122), .B(n2123), .Z(n2016) );
  NANDN U2122 ( .A(n2124), .B(n2125), .Z(n2123) );
  NAND U2123 ( .A(n2126), .B(n2127), .Z(n2125) );
  ANDN U2124 ( .B(B[77]), .A(n41), .Z(n2018) );
  XOR U2125 ( .A(n2025), .B(n2128), .Z(n2019) );
  XNOR U2126 ( .A(n2023), .B(n2026), .Z(n2128) );
  NAND U2127 ( .A(A[2]), .B(B[78]), .Z(n2026) );
  NANDN U2128 ( .A(n2129), .B(n2130), .Z(n2023) );
  AND U2129 ( .A(A[0]), .B(B[79]), .Z(n2130) );
  XNOR U2130 ( .A(n2028), .B(n2131), .Z(n2025) );
  NAND U2131 ( .A(A[0]), .B(B[80]), .Z(n2131) );
  NAND U2132 ( .A(B[79]), .B(A[1]), .Z(n2028) );
  NAND U2133 ( .A(n2132), .B(n2133), .Z(n86) );
  NANDN U2134 ( .A(n2134), .B(n2135), .Z(n2133) );
  OR U2135 ( .A(n2136), .B(n2137), .Z(n2135) );
  NAND U2136 ( .A(n2137), .B(n2136), .Z(n2132) );
  XOR U2137 ( .A(n88), .B(n87), .Z(\A1[77] ) );
  XOR U2138 ( .A(n2137), .B(n2138), .Z(n87) );
  XNOR U2139 ( .A(n2136), .B(n2134), .Z(n2138) );
  AND U2140 ( .A(n2139), .B(n2140), .Z(n2134) );
  NANDN U2141 ( .A(n2141), .B(n2142), .Z(n2140) );
  NANDN U2142 ( .A(n2143), .B(n2144), .Z(n2142) );
  NANDN U2143 ( .A(n2144), .B(n2143), .Z(n2139) );
  ANDN U2144 ( .B(B[64]), .A(n29), .Z(n2136) );
  XNOR U2145 ( .A(n2043), .B(n2145), .Z(n2137) );
  XNOR U2146 ( .A(n2042), .B(n2040), .Z(n2145) );
  AND U2147 ( .A(n2146), .B(n2147), .Z(n2040) );
  NANDN U2148 ( .A(n2148), .B(n2149), .Z(n2147) );
  OR U2149 ( .A(n2150), .B(n2151), .Z(n2149) );
  NAND U2150 ( .A(n2151), .B(n2150), .Z(n2146) );
  ANDN U2151 ( .B(B[65]), .A(n30), .Z(n2042) );
  XNOR U2152 ( .A(n2050), .B(n2152), .Z(n2043) );
  XNOR U2153 ( .A(n2049), .B(n2047), .Z(n2152) );
  AND U2154 ( .A(n2153), .B(n2154), .Z(n2047) );
  NANDN U2155 ( .A(n2155), .B(n2156), .Z(n2154) );
  NANDN U2156 ( .A(n2157), .B(n2158), .Z(n2156) );
  NANDN U2157 ( .A(n2158), .B(n2157), .Z(n2153) );
  ANDN U2158 ( .B(B[66]), .A(n31), .Z(n2049) );
  XNOR U2159 ( .A(n2057), .B(n2159), .Z(n2050) );
  XNOR U2160 ( .A(n2056), .B(n2054), .Z(n2159) );
  AND U2161 ( .A(n2160), .B(n2161), .Z(n2054) );
  NANDN U2162 ( .A(n2162), .B(n2163), .Z(n2161) );
  OR U2163 ( .A(n2164), .B(n2165), .Z(n2163) );
  NAND U2164 ( .A(n2165), .B(n2164), .Z(n2160) );
  ANDN U2165 ( .B(B[67]), .A(n32), .Z(n2056) );
  XNOR U2166 ( .A(n2064), .B(n2166), .Z(n2057) );
  XNOR U2167 ( .A(n2063), .B(n2061), .Z(n2166) );
  AND U2168 ( .A(n2167), .B(n2168), .Z(n2061) );
  NANDN U2169 ( .A(n2169), .B(n2170), .Z(n2168) );
  NANDN U2170 ( .A(n2171), .B(n2172), .Z(n2170) );
  NANDN U2171 ( .A(n2172), .B(n2171), .Z(n2167) );
  ANDN U2172 ( .B(B[68]), .A(n33), .Z(n2063) );
  XNOR U2173 ( .A(n2071), .B(n2173), .Z(n2064) );
  XNOR U2174 ( .A(n2070), .B(n2068), .Z(n2173) );
  AND U2175 ( .A(n2174), .B(n2175), .Z(n2068) );
  NANDN U2176 ( .A(n2176), .B(n2177), .Z(n2175) );
  OR U2177 ( .A(n2178), .B(n2179), .Z(n2177) );
  NAND U2178 ( .A(n2179), .B(n2178), .Z(n2174) );
  ANDN U2179 ( .B(B[69]), .A(n34), .Z(n2070) );
  XNOR U2180 ( .A(n2078), .B(n2180), .Z(n2071) );
  XNOR U2181 ( .A(n2077), .B(n2075), .Z(n2180) );
  AND U2182 ( .A(n2181), .B(n2182), .Z(n2075) );
  NANDN U2183 ( .A(n2183), .B(n2184), .Z(n2182) );
  NANDN U2184 ( .A(n2185), .B(n2186), .Z(n2184) );
  NANDN U2185 ( .A(n2186), .B(n2185), .Z(n2181) );
  ANDN U2186 ( .B(B[70]), .A(n35), .Z(n2077) );
  XNOR U2187 ( .A(n2085), .B(n2187), .Z(n2078) );
  XNOR U2188 ( .A(n2084), .B(n2082), .Z(n2187) );
  AND U2189 ( .A(n2188), .B(n2189), .Z(n2082) );
  NANDN U2190 ( .A(n2190), .B(n2191), .Z(n2189) );
  OR U2191 ( .A(n2192), .B(n2193), .Z(n2191) );
  NAND U2192 ( .A(n2193), .B(n2192), .Z(n2188) );
  ANDN U2193 ( .B(B[71]), .A(n36), .Z(n2084) );
  XNOR U2194 ( .A(n2092), .B(n2194), .Z(n2085) );
  XNOR U2195 ( .A(n2091), .B(n2089), .Z(n2194) );
  AND U2196 ( .A(n2195), .B(n2196), .Z(n2089) );
  NANDN U2197 ( .A(n2197), .B(n2198), .Z(n2196) );
  NANDN U2198 ( .A(n2199), .B(n2200), .Z(n2198) );
  NANDN U2199 ( .A(n2200), .B(n2199), .Z(n2195) );
  ANDN U2200 ( .B(B[72]), .A(n37), .Z(n2091) );
  XNOR U2201 ( .A(n2099), .B(n2201), .Z(n2092) );
  XNOR U2202 ( .A(n2098), .B(n2096), .Z(n2201) );
  AND U2203 ( .A(n2202), .B(n2203), .Z(n2096) );
  NANDN U2204 ( .A(n2204), .B(n2205), .Z(n2203) );
  OR U2205 ( .A(n2206), .B(n2207), .Z(n2205) );
  NAND U2206 ( .A(n2207), .B(n2206), .Z(n2202) );
  ANDN U2207 ( .B(B[73]), .A(n38), .Z(n2098) );
  XNOR U2208 ( .A(n2106), .B(n2208), .Z(n2099) );
  XNOR U2209 ( .A(n2105), .B(n2103), .Z(n2208) );
  AND U2210 ( .A(n2209), .B(n2210), .Z(n2103) );
  NANDN U2211 ( .A(n2211), .B(n2212), .Z(n2210) );
  NANDN U2212 ( .A(n2213), .B(n2214), .Z(n2212) );
  NANDN U2213 ( .A(n2214), .B(n2213), .Z(n2209) );
  ANDN U2214 ( .B(B[74]), .A(n39), .Z(n2105) );
  XNOR U2215 ( .A(n2113), .B(n2215), .Z(n2106) );
  XNOR U2216 ( .A(n2112), .B(n2110), .Z(n2215) );
  AND U2217 ( .A(n2216), .B(n2217), .Z(n2110) );
  NANDN U2218 ( .A(n2218), .B(n2219), .Z(n2217) );
  OR U2219 ( .A(n2220), .B(n2221), .Z(n2219) );
  NAND U2220 ( .A(n2221), .B(n2220), .Z(n2216) );
  ANDN U2221 ( .B(B[75]), .A(n40), .Z(n2112) );
  XNOR U2222 ( .A(n2120), .B(n2222), .Z(n2113) );
  XNOR U2223 ( .A(n2119), .B(n2117), .Z(n2222) );
  AND U2224 ( .A(n2223), .B(n2224), .Z(n2117) );
  NANDN U2225 ( .A(n2225), .B(n2226), .Z(n2224) );
  NAND U2226 ( .A(n2227), .B(n2228), .Z(n2226) );
  ANDN U2227 ( .B(B[76]), .A(n41), .Z(n2119) );
  XOR U2228 ( .A(n2126), .B(n2229), .Z(n2120) );
  XNOR U2229 ( .A(n2124), .B(n2127), .Z(n2229) );
  NAND U2230 ( .A(A[2]), .B(B[77]), .Z(n2127) );
  NANDN U2231 ( .A(n2230), .B(n2231), .Z(n2124) );
  AND U2232 ( .A(A[0]), .B(B[78]), .Z(n2231) );
  XNOR U2233 ( .A(n2129), .B(n2232), .Z(n2126) );
  NAND U2234 ( .A(A[0]), .B(B[79]), .Z(n2232) );
  NAND U2235 ( .A(B[78]), .B(A[1]), .Z(n2129) );
  NAND U2236 ( .A(n2233), .B(n2234), .Z(n88) );
  NANDN U2237 ( .A(n2235), .B(n2236), .Z(n2234) );
  OR U2238 ( .A(n2237), .B(n2238), .Z(n2236) );
  NAND U2239 ( .A(n2238), .B(n2237), .Z(n2233) );
  XOR U2240 ( .A(n90), .B(n89), .Z(\A1[76] ) );
  XOR U2241 ( .A(n2238), .B(n2239), .Z(n89) );
  XNOR U2242 ( .A(n2237), .B(n2235), .Z(n2239) );
  AND U2243 ( .A(n2240), .B(n2241), .Z(n2235) );
  NANDN U2244 ( .A(n2242), .B(n2243), .Z(n2241) );
  NANDN U2245 ( .A(n2244), .B(n2245), .Z(n2243) );
  NANDN U2246 ( .A(n2245), .B(n2244), .Z(n2240) );
  ANDN U2247 ( .B(B[63]), .A(n29), .Z(n2237) );
  XNOR U2248 ( .A(n2144), .B(n2246), .Z(n2238) );
  XNOR U2249 ( .A(n2143), .B(n2141), .Z(n2246) );
  AND U2250 ( .A(n2247), .B(n2248), .Z(n2141) );
  NANDN U2251 ( .A(n2249), .B(n2250), .Z(n2248) );
  OR U2252 ( .A(n2251), .B(n2252), .Z(n2250) );
  NAND U2253 ( .A(n2252), .B(n2251), .Z(n2247) );
  ANDN U2254 ( .B(B[64]), .A(n30), .Z(n2143) );
  XNOR U2255 ( .A(n2151), .B(n2253), .Z(n2144) );
  XNOR U2256 ( .A(n2150), .B(n2148), .Z(n2253) );
  AND U2257 ( .A(n2254), .B(n2255), .Z(n2148) );
  NANDN U2258 ( .A(n2256), .B(n2257), .Z(n2255) );
  NANDN U2259 ( .A(n2258), .B(n2259), .Z(n2257) );
  NANDN U2260 ( .A(n2259), .B(n2258), .Z(n2254) );
  ANDN U2261 ( .B(B[65]), .A(n31), .Z(n2150) );
  XNOR U2262 ( .A(n2158), .B(n2260), .Z(n2151) );
  XNOR U2263 ( .A(n2157), .B(n2155), .Z(n2260) );
  AND U2264 ( .A(n2261), .B(n2262), .Z(n2155) );
  NANDN U2265 ( .A(n2263), .B(n2264), .Z(n2262) );
  OR U2266 ( .A(n2265), .B(n2266), .Z(n2264) );
  NAND U2267 ( .A(n2266), .B(n2265), .Z(n2261) );
  ANDN U2268 ( .B(B[66]), .A(n32), .Z(n2157) );
  XNOR U2269 ( .A(n2165), .B(n2267), .Z(n2158) );
  XNOR U2270 ( .A(n2164), .B(n2162), .Z(n2267) );
  AND U2271 ( .A(n2268), .B(n2269), .Z(n2162) );
  NANDN U2272 ( .A(n2270), .B(n2271), .Z(n2269) );
  NANDN U2273 ( .A(n2272), .B(n2273), .Z(n2271) );
  NANDN U2274 ( .A(n2273), .B(n2272), .Z(n2268) );
  ANDN U2275 ( .B(B[67]), .A(n33), .Z(n2164) );
  XNOR U2276 ( .A(n2172), .B(n2274), .Z(n2165) );
  XNOR U2277 ( .A(n2171), .B(n2169), .Z(n2274) );
  AND U2278 ( .A(n2275), .B(n2276), .Z(n2169) );
  NANDN U2279 ( .A(n2277), .B(n2278), .Z(n2276) );
  OR U2280 ( .A(n2279), .B(n2280), .Z(n2278) );
  NAND U2281 ( .A(n2280), .B(n2279), .Z(n2275) );
  ANDN U2282 ( .B(B[68]), .A(n34), .Z(n2171) );
  XNOR U2283 ( .A(n2179), .B(n2281), .Z(n2172) );
  XNOR U2284 ( .A(n2178), .B(n2176), .Z(n2281) );
  AND U2285 ( .A(n2282), .B(n2283), .Z(n2176) );
  NANDN U2286 ( .A(n2284), .B(n2285), .Z(n2283) );
  NANDN U2287 ( .A(n2286), .B(n2287), .Z(n2285) );
  NANDN U2288 ( .A(n2287), .B(n2286), .Z(n2282) );
  ANDN U2289 ( .B(B[69]), .A(n35), .Z(n2178) );
  XNOR U2290 ( .A(n2186), .B(n2288), .Z(n2179) );
  XNOR U2291 ( .A(n2185), .B(n2183), .Z(n2288) );
  AND U2292 ( .A(n2289), .B(n2290), .Z(n2183) );
  NANDN U2293 ( .A(n2291), .B(n2292), .Z(n2290) );
  OR U2294 ( .A(n2293), .B(n2294), .Z(n2292) );
  NAND U2295 ( .A(n2294), .B(n2293), .Z(n2289) );
  ANDN U2296 ( .B(B[70]), .A(n36), .Z(n2185) );
  XNOR U2297 ( .A(n2193), .B(n2295), .Z(n2186) );
  XNOR U2298 ( .A(n2192), .B(n2190), .Z(n2295) );
  AND U2299 ( .A(n2296), .B(n2297), .Z(n2190) );
  NANDN U2300 ( .A(n2298), .B(n2299), .Z(n2297) );
  NANDN U2301 ( .A(n2300), .B(n2301), .Z(n2299) );
  NANDN U2302 ( .A(n2301), .B(n2300), .Z(n2296) );
  ANDN U2303 ( .B(B[71]), .A(n37), .Z(n2192) );
  XNOR U2304 ( .A(n2200), .B(n2302), .Z(n2193) );
  XNOR U2305 ( .A(n2199), .B(n2197), .Z(n2302) );
  AND U2306 ( .A(n2303), .B(n2304), .Z(n2197) );
  NANDN U2307 ( .A(n2305), .B(n2306), .Z(n2304) );
  OR U2308 ( .A(n2307), .B(n2308), .Z(n2306) );
  NAND U2309 ( .A(n2308), .B(n2307), .Z(n2303) );
  ANDN U2310 ( .B(B[72]), .A(n38), .Z(n2199) );
  XNOR U2311 ( .A(n2207), .B(n2309), .Z(n2200) );
  XNOR U2312 ( .A(n2206), .B(n2204), .Z(n2309) );
  AND U2313 ( .A(n2310), .B(n2311), .Z(n2204) );
  NANDN U2314 ( .A(n2312), .B(n2313), .Z(n2311) );
  NANDN U2315 ( .A(n2314), .B(n2315), .Z(n2313) );
  NANDN U2316 ( .A(n2315), .B(n2314), .Z(n2310) );
  ANDN U2317 ( .B(B[73]), .A(n39), .Z(n2206) );
  XNOR U2318 ( .A(n2214), .B(n2316), .Z(n2207) );
  XNOR U2319 ( .A(n2213), .B(n2211), .Z(n2316) );
  AND U2320 ( .A(n2317), .B(n2318), .Z(n2211) );
  NANDN U2321 ( .A(n2319), .B(n2320), .Z(n2318) );
  OR U2322 ( .A(n2321), .B(n2322), .Z(n2320) );
  NAND U2323 ( .A(n2322), .B(n2321), .Z(n2317) );
  ANDN U2324 ( .B(B[74]), .A(n40), .Z(n2213) );
  XNOR U2325 ( .A(n2221), .B(n2323), .Z(n2214) );
  XNOR U2326 ( .A(n2220), .B(n2218), .Z(n2323) );
  AND U2327 ( .A(n2324), .B(n2325), .Z(n2218) );
  NANDN U2328 ( .A(n2326), .B(n2327), .Z(n2325) );
  NAND U2329 ( .A(n2328), .B(n2329), .Z(n2327) );
  ANDN U2330 ( .B(B[75]), .A(n41), .Z(n2220) );
  XOR U2331 ( .A(n2227), .B(n2330), .Z(n2221) );
  XNOR U2332 ( .A(n2225), .B(n2228), .Z(n2330) );
  NAND U2333 ( .A(A[2]), .B(B[76]), .Z(n2228) );
  NANDN U2334 ( .A(n2331), .B(n2332), .Z(n2225) );
  AND U2335 ( .A(A[0]), .B(B[77]), .Z(n2332) );
  XNOR U2336 ( .A(n2230), .B(n2333), .Z(n2227) );
  NAND U2337 ( .A(A[0]), .B(B[78]), .Z(n2333) );
  NAND U2338 ( .A(B[77]), .B(A[1]), .Z(n2230) );
  NAND U2339 ( .A(n2334), .B(n2335), .Z(n90) );
  NANDN U2340 ( .A(n2336), .B(n2337), .Z(n2335) );
  OR U2341 ( .A(n2338), .B(n2339), .Z(n2337) );
  NAND U2342 ( .A(n2339), .B(n2338), .Z(n2334) );
  XOR U2343 ( .A(n92), .B(n91), .Z(\A1[75] ) );
  XOR U2344 ( .A(n2339), .B(n2340), .Z(n91) );
  XNOR U2345 ( .A(n2338), .B(n2336), .Z(n2340) );
  AND U2346 ( .A(n2341), .B(n2342), .Z(n2336) );
  NANDN U2347 ( .A(n2343), .B(n2344), .Z(n2342) );
  NANDN U2348 ( .A(n2345), .B(n2346), .Z(n2344) );
  NANDN U2349 ( .A(n2346), .B(n2345), .Z(n2341) );
  ANDN U2350 ( .B(B[62]), .A(n29), .Z(n2338) );
  XNOR U2351 ( .A(n2245), .B(n2347), .Z(n2339) );
  XNOR U2352 ( .A(n2244), .B(n2242), .Z(n2347) );
  AND U2353 ( .A(n2348), .B(n2349), .Z(n2242) );
  NANDN U2354 ( .A(n2350), .B(n2351), .Z(n2349) );
  OR U2355 ( .A(n2352), .B(n2353), .Z(n2351) );
  NAND U2356 ( .A(n2353), .B(n2352), .Z(n2348) );
  ANDN U2357 ( .B(B[63]), .A(n30), .Z(n2244) );
  XNOR U2358 ( .A(n2252), .B(n2354), .Z(n2245) );
  XNOR U2359 ( .A(n2251), .B(n2249), .Z(n2354) );
  AND U2360 ( .A(n2355), .B(n2356), .Z(n2249) );
  NANDN U2361 ( .A(n2357), .B(n2358), .Z(n2356) );
  NANDN U2362 ( .A(n2359), .B(n2360), .Z(n2358) );
  NANDN U2363 ( .A(n2360), .B(n2359), .Z(n2355) );
  ANDN U2364 ( .B(B[64]), .A(n31), .Z(n2251) );
  XNOR U2365 ( .A(n2259), .B(n2361), .Z(n2252) );
  XNOR U2366 ( .A(n2258), .B(n2256), .Z(n2361) );
  AND U2367 ( .A(n2362), .B(n2363), .Z(n2256) );
  NANDN U2368 ( .A(n2364), .B(n2365), .Z(n2363) );
  OR U2369 ( .A(n2366), .B(n2367), .Z(n2365) );
  NAND U2370 ( .A(n2367), .B(n2366), .Z(n2362) );
  ANDN U2371 ( .B(B[65]), .A(n32), .Z(n2258) );
  XNOR U2372 ( .A(n2266), .B(n2368), .Z(n2259) );
  XNOR U2373 ( .A(n2265), .B(n2263), .Z(n2368) );
  AND U2374 ( .A(n2369), .B(n2370), .Z(n2263) );
  NANDN U2375 ( .A(n2371), .B(n2372), .Z(n2370) );
  NANDN U2376 ( .A(n2373), .B(n2374), .Z(n2372) );
  NANDN U2377 ( .A(n2374), .B(n2373), .Z(n2369) );
  ANDN U2378 ( .B(B[66]), .A(n33), .Z(n2265) );
  XNOR U2379 ( .A(n2273), .B(n2375), .Z(n2266) );
  XNOR U2380 ( .A(n2272), .B(n2270), .Z(n2375) );
  AND U2381 ( .A(n2376), .B(n2377), .Z(n2270) );
  NANDN U2382 ( .A(n2378), .B(n2379), .Z(n2377) );
  OR U2383 ( .A(n2380), .B(n2381), .Z(n2379) );
  NAND U2384 ( .A(n2381), .B(n2380), .Z(n2376) );
  ANDN U2385 ( .B(B[67]), .A(n34), .Z(n2272) );
  XNOR U2386 ( .A(n2280), .B(n2382), .Z(n2273) );
  XNOR U2387 ( .A(n2279), .B(n2277), .Z(n2382) );
  AND U2388 ( .A(n2383), .B(n2384), .Z(n2277) );
  NANDN U2389 ( .A(n2385), .B(n2386), .Z(n2384) );
  NANDN U2390 ( .A(n2387), .B(n2388), .Z(n2386) );
  NANDN U2391 ( .A(n2388), .B(n2387), .Z(n2383) );
  ANDN U2392 ( .B(B[68]), .A(n35), .Z(n2279) );
  XNOR U2393 ( .A(n2287), .B(n2389), .Z(n2280) );
  XNOR U2394 ( .A(n2286), .B(n2284), .Z(n2389) );
  AND U2395 ( .A(n2390), .B(n2391), .Z(n2284) );
  NANDN U2396 ( .A(n2392), .B(n2393), .Z(n2391) );
  OR U2397 ( .A(n2394), .B(n2395), .Z(n2393) );
  NAND U2398 ( .A(n2395), .B(n2394), .Z(n2390) );
  ANDN U2399 ( .B(B[69]), .A(n36), .Z(n2286) );
  XNOR U2400 ( .A(n2294), .B(n2396), .Z(n2287) );
  XNOR U2401 ( .A(n2293), .B(n2291), .Z(n2396) );
  AND U2402 ( .A(n2397), .B(n2398), .Z(n2291) );
  NANDN U2403 ( .A(n2399), .B(n2400), .Z(n2398) );
  NANDN U2404 ( .A(n2401), .B(n2402), .Z(n2400) );
  NANDN U2405 ( .A(n2402), .B(n2401), .Z(n2397) );
  ANDN U2406 ( .B(B[70]), .A(n37), .Z(n2293) );
  XNOR U2407 ( .A(n2301), .B(n2403), .Z(n2294) );
  XNOR U2408 ( .A(n2300), .B(n2298), .Z(n2403) );
  AND U2409 ( .A(n2404), .B(n2405), .Z(n2298) );
  NANDN U2410 ( .A(n2406), .B(n2407), .Z(n2405) );
  OR U2411 ( .A(n2408), .B(n2409), .Z(n2407) );
  NAND U2412 ( .A(n2409), .B(n2408), .Z(n2404) );
  ANDN U2413 ( .B(B[71]), .A(n38), .Z(n2300) );
  XNOR U2414 ( .A(n2308), .B(n2410), .Z(n2301) );
  XNOR U2415 ( .A(n2307), .B(n2305), .Z(n2410) );
  AND U2416 ( .A(n2411), .B(n2412), .Z(n2305) );
  NANDN U2417 ( .A(n2413), .B(n2414), .Z(n2412) );
  NANDN U2418 ( .A(n2415), .B(n2416), .Z(n2414) );
  NANDN U2419 ( .A(n2416), .B(n2415), .Z(n2411) );
  ANDN U2420 ( .B(B[72]), .A(n39), .Z(n2307) );
  XNOR U2421 ( .A(n2315), .B(n2417), .Z(n2308) );
  XNOR U2422 ( .A(n2314), .B(n2312), .Z(n2417) );
  AND U2423 ( .A(n2418), .B(n2419), .Z(n2312) );
  NANDN U2424 ( .A(n2420), .B(n2421), .Z(n2419) );
  OR U2425 ( .A(n2422), .B(n2423), .Z(n2421) );
  NAND U2426 ( .A(n2423), .B(n2422), .Z(n2418) );
  ANDN U2427 ( .B(B[73]), .A(n40), .Z(n2314) );
  XNOR U2428 ( .A(n2322), .B(n2424), .Z(n2315) );
  XNOR U2429 ( .A(n2321), .B(n2319), .Z(n2424) );
  AND U2430 ( .A(n2425), .B(n2426), .Z(n2319) );
  NANDN U2431 ( .A(n2427), .B(n2428), .Z(n2426) );
  NAND U2432 ( .A(n2429), .B(n2430), .Z(n2428) );
  ANDN U2433 ( .B(B[74]), .A(n41), .Z(n2321) );
  XOR U2434 ( .A(n2328), .B(n2431), .Z(n2322) );
  XNOR U2435 ( .A(n2326), .B(n2329), .Z(n2431) );
  NAND U2436 ( .A(A[2]), .B(B[75]), .Z(n2329) );
  NANDN U2437 ( .A(n2432), .B(n2433), .Z(n2326) );
  AND U2438 ( .A(A[0]), .B(B[76]), .Z(n2433) );
  XNOR U2439 ( .A(n2331), .B(n2434), .Z(n2328) );
  NAND U2440 ( .A(A[0]), .B(B[77]), .Z(n2434) );
  NAND U2441 ( .A(B[76]), .B(A[1]), .Z(n2331) );
  NAND U2442 ( .A(n2435), .B(n2436), .Z(n92) );
  NANDN U2443 ( .A(n2437), .B(n2438), .Z(n2436) );
  OR U2444 ( .A(n2439), .B(n2440), .Z(n2438) );
  NAND U2445 ( .A(n2440), .B(n2439), .Z(n2435) );
  XOR U2446 ( .A(n94), .B(n93), .Z(\A1[74] ) );
  XOR U2447 ( .A(n2440), .B(n2441), .Z(n93) );
  XNOR U2448 ( .A(n2439), .B(n2437), .Z(n2441) );
  AND U2449 ( .A(n2442), .B(n2443), .Z(n2437) );
  NANDN U2450 ( .A(n2444), .B(n2445), .Z(n2443) );
  NANDN U2451 ( .A(n2446), .B(n2447), .Z(n2445) );
  NANDN U2452 ( .A(n2447), .B(n2446), .Z(n2442) );
  ANDN U2453 ( .B(B[61]), .A(n29), .Z(n2439) );
  XNOR U2454 ( .A(n2346), .B(n2448), .Z(n2440) );
  XNOR U2455 ( .A(n2345), .B(n2343), .Z(n2448) );
  AND U2456 ( .A(n2449), .B(n2450), .Z(n2343) );
  NANDN U2457 ( .A(n2451), .B(n2452), .Z(n2450) );
  OR U2458 ( .A(n2453), .B(n2454), .Z(n2452) );
  NAND U2459 ( .A(n2454), .B(n2453), .Z(n2449) );
  ANDN U2460 ( .B(B[62]), .A(n30), .Z(n2345) );
  XNOR U2461 ( .A(n2353), .B(n2455), .Z(n2346) );
  XNOR U2462 ( .A(n2352), .B(n2350), .Z(n2455) );
  AND U2463 ( .A(n2456), .B(n2457), .Z(n2350) );
  NANDN U2464 ( .A(n2458), .B(n2459), .Z(n2457) );
  NANDN U2465 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U2466 ( .A(n2461), .B(n2460), .Z(n2456) );
  ANDN U2467 ( .B(B[63]), .A(n31), .Z(n2352) );
  XNOR U2468 ( .A(n2360), .B(n2462), .Z(n2353) );
  XNOR U2469 ( .A(n2359), .B(n2357), .Z(n2462) );
  AND U2470 ( .A(n2463), .B(n2464), .Z(n2357) );
  NANDN U2471 ( .A(n2465), .B(n2466), .Z(n2464) );
  OR U2472 ( .A(n2467), .B(n2468), .Z(n2466) );
  NAND U2473 ( .A(n2468), .B(n2467), .Z(n2463) );
  ANDN U2474 ( .B(B[64]), .A(n32), .Z(n2359) );
  XNOR U2475 ( .A(n2367), .B(n2469), .Z(n2360) );
  XNOR U2476 ( .A(n2366), .B(n2364), .Z(n2469) );
  AND U2477 ( .A(n2470), .B(n2471), .Z(n2364) );
  NANDN U2478 ( .A(n2472), .B(n2473), .Z(n2471) );
  NANDN U2479 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U2480 ( .A(n2475), .B(n2474), .Z(n2470) );
  ANDN U2481 ( .B(B[65]), .A(n33), .Z(n2366) );
  XNOR U2482 ( .A(n2374), .B(n2476), .Z(n2367) );
  XNOR U2483 ( .A(n2373), .B(n2371), .Z(n2476) );
  AND U2484 ( .A(n2477), .B(n2478), .Z(n2371) );
  NANDN U2485 ( .A(n2479), .B(n2480), .Z(n2478) );
  OR U2486 ( .A(n2481), .B(n2482), .Z(n2480) );
  NAND U2487 ( .A(n2482), .B(n2481), .Z(n2477) );
  ANDN U2488 ( .B(B[66]), .A(n34), .Z(n2373) );
  XNOR U2489 ( .A(n2381), .B(n2483), .Z(n2374) );
  XNOR U2490 ( .A(n2380), .B(n2378), .Z(n2483) );
  AND U2491 ( .A(n2484), .B(n2485), .Z(n2378) );
  NANDN U2492 ( .A(n2486), .B(n2487), .Z(n2485) );
  NANDN U2493 ( .A(n2488), .B(n2489), .Z(n2487) );
  NANDN U2494 ( .A(n2489), .B(n2488), .Z(n2484) );
  ANDN U2495 ( .B(B[67]), .A(n35), .Z(n2380) );
  XNOR U2496 ( .A(n2388), .B(n2490), .Z(n2381) );
  XNOR U2497 ( .A(n2387), .B(n2385), .Z(n2490) );
  AND U2498 ( .A(n2491), .B(n2492), .Z(n2385) );
  NANDN U2499 ( .A(n2493), .B(n2494), .Z(n2492) );
  OR U2500 ( .A(n2495), .B(n2496), .Z(n2494) );
  NAND U2501 ( .A(n2496), .B(n2495), .Z(n2491) );
  ANDN U2502 ( .B(B[68]), .A(n36), .Z(n2387) );
  XNOR U2503 ( .A(n2395), .B(n2497), .Z(n2388) );
  XNOR U2504 ( .A(n2394), .B(n2392), .Z(n2497) );
  AND U2505 ( .A(n2498), .B(n2499), .Z(n2392) );
  NANDN U2506 ( .A(n2500), .B(n2501), .Z(n2499) );
  NANDN U2507 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U2508 ( .A(n2503), .B(n2502), .Z(n2498) );
  ANDN U2509 ( .B(B[69]), .A(n37), .Z(n2394) );
  XNOR U2510 ( .A(n2402), .B(n2504), .Z(n2395) );
  XNOR U2511 ( .A(n2401), .B(n2399), .Z(n2504) );
  AND U2512 ( .A(n2505), .B(n2506), .Z(n2399) );
  NANDN U2513 ( .A(n2507), .B(n2508), .Z(n2506) );
  OR U2514 ( .A(n2509), .B(n2510), .Z(n2508) );
  NAND U2515 ( .A(n2510), .B(n2509), .Z(n2505) );
  ANDN U2516 ( .B(B[70]), .A(n38), .Z(n2401) );
  XNOR U2517 ( .A(n2409), .B(n2511), .Z(n2402) );
  XNOR U2518 ( .A(n2408), .B(n2406), .Z(n2511) );
  AND U2519 ( .A(n2512), .B(n2513), .Z(n2406) );
  NANDN U2520 ( .A(n2514), .B(n2515), .Z(n2513) );
  NANDN U2521 ( .A(n2516), .B(n2517), .Z(n2515) );
  NANDN U2522 ( .A(n2517), .B(n2516), .Z(n2512) );
  ANDN U2523 ( .B(B[71]), .A(n39), .Z(n2408) );
  XNOR U2524 ( .A(n2416), .B(n2518), .Z(n2409) );
  XNOR U2525 ( .A(n2415), .B(n2413), .Z(n2518) );
  AND U2526 ( .A(n2519), .B(n2520), .Z(n2413) );
  NANDN U2527 ( .A(n2521), .B(n2522), .Z(n2520) );
  OR U2528 ( .A(n2523), .B(n2524), .Z(n2522) );
  NAND U2529 ( .A(n2524), .B(n2523), .Z(n2519) );
  ANDN U2530 ( .B(B[72]), .A(n40), .Z(n2415) );
  XNOR U2531 ( .A(n2423), .B(n2525), .Z(n2416) );
  XNOR U2532 ( .A(n2422), .B(n2420), .Z(n2525) );
  AND U2533 ( .A(n2526), .B(n2527), .Z(n2420) );
  NANDN U2534 ( .A(n2528), .B(n2529), .Z(n2527) );
  NAND U2535 ( .A(n2530), .B(n2531), .Z(n2529) );
  ANDN U2536 ( .B(B[73]), .A(n41), .Z(n2422) );
  XOR U2537 ( .A(n2429), .B(n2532), .Z(n2423) );
  XNOR U2538 ( .A(n2427), .B(n2430), .Z(n2532) );
  NAND U2539 ( .A(A[2]), .B(B[74]), .Z(n2430) );
  NANDN U2540 ( .A(n2533), .B(n2534), .Z(n2427) );
  AND U2541 ( .A(A[0]), .B(B[75]), .Z(n2534) );
  XNOR U2542 ( .A(n2432), .B(n2535), .Z(n2429) );
  NAND U2543 ( .A(A[0]), .B(B[76]), .Z(n2535) );
  NAND U2544 ( .A(B[75]), .B(A[1]), .Z(n2432) );
  NAND U2545 ( .A(n2536), .B(n2537), .Z(n94) );
  NANDN U2546 ( .A(n2538), .B(n2539), .Z(n2537) );
  OR U2547 ( .A(n2540), .B(n2541), .Z(n2539) );
  NAND U2548 ( .A(n2541), .B(n2540), .Z(n2536) );
  XOR U2549 ( .A(n96), .B(n95), .Z(\A1[73] ) );
  XOR U2550 ( .A(n2541), .B(n2542), .Z(n95) );
  XNOR U2551 ( .A(n2540), .B(n2538), .Z(n2542) );
  AND U2552 ( .A(n2543), .B(n2544), .Z(n2538) );
  NANDN U2553 ( .A(n2545), .B(n2546), .Z(n2544) );
  NANDN U2554 ( .A(n2547), .B(n2548), .Z(n2546) );
  NANDN U2555 ( .A(n2548), .B(n2547), .Z(n2543) );
  ANDN U2556 ( .B(B[60]), .A(n29), .Z(n2540) );
  XNOR U2557 ( .A(n2447), .B(n2549), .Z(n2541) );
  XNOR U2558 ( .A(n2446), .B(n2444), .Z(n2549) );
  AND U2559 ( .A(n2550), .B(n2551), .Z(n2444) );
  NANDN U2560 ( .A(n2552), .B(n2553), .Z(n2551) );
  OR U2561 ( .A(n2554), .B(n2555), .Z(n2553) );
  NAND U2562 ( .A(n2555), .B(n2554), .Z(n2550) );
  ANDN U2563 ( .B(B[61]), .A(n30), .Z(n2446) );
  XNOR U2564 ( .A(n2454), .B(n2556), .Z(n2447) );
  XNOR U2565 ( .A(n2453), .B(n2451), .Z(n2556) );
  AND U2566 ( .A(n2557), .B(n2558), .Z(n2451) );
  NANDN U2567 ( .A(n2559), .B(n2560), .Z(n2558) );
  NANDN U2568 ( .A(n2561), .B(n2562), .Z(n2560) );
  NANDN U2569 ( .A(n2562), .B(n2561), .Z(n2557) );
  ANDN U2570 ( .B(B[62]), .A(n31), .Z(n2453) );
  XNOR U2571 ( .A(n2461), .B(n2563), .Z(n2454) );
  XNOR U2572 ( .A(n2460), .B(n2458), .Z(n2563) );
  AND U2573 ( .A(n2564), .B(n2565), .Z(n2458) );
  NANDN U2574 ( .A(n2566), .B(n2567), .Z(n2565) );
  OR U2575 ( .A(n2568), .B(n2569), .Z(n2567) );
  NAND U2576 ( .A(n2569), .B(n2568), .Z(n2564) );
  ANDN U2577 ( .B(B[63]), .A(n32), .Z(n2460) );
  XNOR U2578 ( .A(n2468), .B(n2570), .Z(n2461) );
  XNOR U2579 ( .A(n2467), .B(n2465), .Z(n2570) );
  AND U2580 ( .A(n2571), .B(n2572), .Z(n2465) );
  NANDN U2581 ( .A(n2573), .B(n2574), .Z(n2572) );
  NANDN U2582 ( .A(n2575), .B(n2576), .Z(n2574) );
  NANDN U2583 ( .A(n2576), .B(n2575), .Z(n2571) );
  ANDN U2584 ( .B(B[64]), .A(n33), .Z(n2467) );
  XNOR U2585 ( .A(n2475), .B(n2577), .Z(n2468) );
  XNOR U2586 ( .A(n2474), .B(n2472), .Z(n2577) );
  AND U2587 ( .A(n2578), .B(n2579), .Z(n2472) );
  NANDN U2588 ( .A(n2580), .B(n2581), .Z(n2579) );
  OR U2589 ( .A(n2582), .B(n2583), .Z(n2581) );
  NAND U2590 ( .A(n2583), .B(n2582), .Z(n2578) );
  ANDN U2591 ( .B(B[65]), .A(n34), .Z(n2474) );
  XNOR U2592 ( .A(n2482), .B(n2584), .Z(n2475) );
  XNOR U2593 ( .A(n2481), .B(n2479), .Z(n2584) );
  AND U2594 ( .A(n2585), .B(n2586), .Z(n2479) );
  NANDN U2595 ( .A(n2587), .B(n2588), .Z(n2586) );
  NANDN U2596 ( .A(n2589), .B(n2590), .Z(n2588) );
  NANDN U2597 ( .A(n2590), .B(n2589), .Z(n2585) );
  ANDN U2598 ( .B(B[66]), .A(n35), .Z(n2481) );
  XNOR U2599 ( .A(n2489), .B(n2591), .Z(n2482) );
  XNOR U2600 ( .A(n2488), .B(n2486), .Z(n2591) );
  AND U2601 ( .A(n2592), .B(n2593), .Z(n2486) );
  NANDN U2602 ( .A(n2594), .B(n2595), .Z(n2593) );
  OR U2603 ( .A(n2596), .B(n2597), .Z(n2595) );
  NAND U2604 ( .A(n2597), .B(n2596), .Z(n2592) );
  ANDN U2605 ( .B(B[67]), .A(n36), .Z(n2488) );
  XNOR U2606 ( .A(n2496), .B(n2598), .Z(n2489) );
  XNOR U2607 ( .A(n2495), .B(n2493), .Z(n2598) );
  AND U2608 ( .A(n2599), .B(n2600), .Z(n2493) );
  NANDN U2609 ( .A(n2601), .B(n2602), .Z(n2600) );
  NANDN U2610 ( .A(n2603), .B(n2604), .Z(n2602) );
  NANDN U2611 ( .A(n2604), .B(n2603), .Z(n2599) );
  ANDN U2612 ( .B(B[68]), .A(n37), .Z(n2495) );
  XNOR U2613 ( .A(n2503), .B(n2605), .Z(n2496) );
  XNOR U2614 ( .A(n2502), .B(n2500), .Z(n2605) );
  AND U2615 ( .A(n2606), .B(n2607), .Z(n2500) );
  NANDN U2616 ( .A(n2608), .B(n2609), .Z(n2607) );
  OR U2617 ( .A(n2610), .B(n2611), .Z(n2609) );
  NAND U2618 ( .A(n2611), .B(n2610), .Z(n2606) );
  ANDN U2619 ( .B(B[69]), .A(n38), .Z(n2502) );
  XNOR U2620 ( .A(n2510), .B(n2612), .Z(n2503) );
  XNOR U2621 ( .A(n2509), .B(n2507), .Z(n2612) );
  AND U2622 ( .A(n2613), .B(n2614), .Z(n2507) );
  NANDN U2623 ( .A(n2615), .B(n2616), .Z(n2614) );
  NANDN U2624 ( .A(n2617), .B(n2618), .Z(n2616) );
  NANDN U2625 ( .A(n2618), .B(n2617), .Z(n2613) );
  ANDN U2626 ( .B(B[70]), .A(n39), .Z(n2509) );
  XNOR U2627 ( .A(n2517), .B(n2619), .Z(n2510) );
  XNOR U2628 ( .A(n2516), .B(n2514), .Z(n2619) );
  AND U2629 ( .A(n2620), .B(n2621), .Z(n2514) );
  NANDN U2630 ( .A(n2622), .B(n2623), .Z(n2621) );
  OR U2631 ( .A(n2624), .B(n2625), .Z(n2623) );
  NAND U2632 ( .A(n2625), .B(n2624), .Z(n2620) );
  ANDN U2633 ( .B(B[71]), .A(n40), .Z(n2516) );
  XNOR U2634 ( .A(n2524), .B(n2626), .Z(n2517) );
  XNOR U2635 ( .A(n2523), .B(n2521), .Z(n2626) );
  AND U2636 ( .A(n2627), .B(n2628), .Z(n2521) );
  NANDN U2637 ( .A(n2629), .B(n2630), .Z(n2628) );
  NAND U2638 ( .A(n2631), .B(n2632), .Z(n2630) );
  ANDN U2639 ( .B(B[72]), .A(n41), .Z(n2523) );
  XOR U2640 ( .A(n2530), .B(n2633), .Z(n2524) );
  XNOR U2641 ( .A(n2528), .B(n2531), .Z(n2633) );
  NAND U2642 ( .A(A[2]), .B(B[73]), .Z(n2531) );
  NANDN U2643 ( .A(n2634), .B(n2635), .Z(n2528) );
  AND U2644 ( .A(A[0]), .B(B[74]), .Z(n2635) );
  XNOR U2645 ( .A(n2533), .B(n2636), .Z(n2530) );
  NAND U2646 ( .A(A[0]), .B(B[75]), .Z(n2636) );
  NAND U2647 ( .A(B[74]), .B(A[1]), .Z(n2533) );
  NAND U2648 ( .A(n2637), .B(n2638), .Z(n96) );
  NANDN U2649 ( .A(n2639), .B(n2640), .Z(n2638) );
  OR U2650 ( .A(n2641), .B(n2642), .Z(n2640) );
  NAND U2651 ( .A(n2642), .B(n2641), .Z(n2637) );
  XOR U2652 ( .A(n98), .B(n97), .Z(\A1[72] ) );
  XOR U2653 ( .A(n2642), .B(n2643), .Z(n97) );
  XNOR U2654 ( .A(n2641), .B(n2639), .Z(n2643) );
  AND U2655 ( .A(n2644), .B(n2645), .Z(n2639) );
  NANDN U2656 ( .A(n2646), .B(n2647), .Z(n2645) );
  NANDN U2657 ( .A(n2648), .B(n2649), .Z(n2647) );
  NANDN U2658 ( .A(n2649), .B(n2648), .Z(n2644) );
  ANDN U2659 ( .B(B[59]), .A(n29), .Z(n2641) );
  XNOR U2660 ( .A(n2548), .B(n2650), .Z(n2642) );
  XNOR U2661 ( .A(n2547), .B(n2545), .Z(n2650) );
  AND U2662 ( .A(n2651), .B(n2652), .Z(n2545) );
  NANDN U2663 ( .A(n2653), .B(n2654), .Z(n2652) );
  OR U2664 ( .A(n2655), .B(n2656), .Z(n2654) );
  NAND U2665 ( .A(n2656), .B(n2655), .Z(n2651) );
  ANDN U2666 ( .B(B[60]), .A(n30), .Z(n2547) );
  XNOR U2667 ( .A(n2555), .B(n2657), .Z(n2548) );
  XNOR U2668 ( .A(n2554), .B(n2552), .Z(n2657) );
  AND U2669 ( .A(n2658), .B(n2659), .Z(n2552) );
  NANDN U2670 ( .A(n2660), .B(n2661), .Z(n2659) );
  NANDN U2671 ( .A(n2662), .B(n2663), .Z(n2661) );
  NANDN U2672 ( .A(n2663), .B(n2662), .Z(n2658) );
  ANDN U2673 ( .B(B[61]), .A(n31), .Z(n2554) );
  XNOR U2674 ( .A(n2562), .B(n2664), .Z(n2555) );
  XNOR U2675 ( .A(n2561), .B(n2559), .Z(n2664) );
  AND U2676 ( .A(n2665), .B(n2666), .Z(n2559) );
  NANDN U2677 ( .A(n2667), .B(n2668), .Z(n2666) );
  OR U2678 ( .A(n2669), .B(n2670), .Z(n2668) );
  NAND U2679 ( .A(n2670), .B(n2669), .Z(n2665) );
  ANDN U2680 ( .B(B[62]), .A(n32), .Z(n2561) );
  XNOR U2681 ( .A(n2569), .B(n2671), .Z(n2562) );
  XNOR U2682 ( .A(n2568), .B(n2566), .Z(n2671) );
  AND U2683 ( .A(n2672), .B(n2673), .Z(n2566) );
  NANDN U2684 ( .A(n2674), .B(n2675), .Z(n2673) );
  NANDN U2685 ( .A(n2676), .B(n2677), .Z(n2675) );
  NANDN U2686 ( .A(n2677), .B(n2676), .Z(n2672) );
  ANDN U2687 ( .B(B[63]), .A(n33), .Z(n2568) );
  XNOR U2688 ( .A(n2576), .B(n2678), .Z(n2569) );
  XNOR U2689 ( .A(n2575), .B(n2573), .Z(n2678) );
  AND U2690 ( .A(n2679), .B(n2680), .Z(n2573) );
  NANDN U2691 ( .A(n2681), .B(n2682), .Z(n2680) );
  OR U2692 ( .A(n2683), .B(n2684), .Z(n2682) );
  NAND U2693 ( .A(n2684), .B(n2683), .Z(n2679) );
  ANDN U2694 ( .B(B[64]), .A(n34), .Z(n2575) );
  XNOR U2695 ( .A(n2583), .B(n2685), .Z(n2576) );
  XNOR U2696 ( .A(n2582), .B(n2580), .Z(n2685) );
  AND U2697 ( .A(n2686), .B(n2687), .Z(n2580) );
  NANDN U2698 ( .A(n2688), .B(n2689), .Z(n2687) );
  NANDN U2699 ( .A(n2690), .B(n2691), .Z(n2689) );
  NANDN U2700 ( .A(n2691), .B(n2690), .Z(n2686) );
  ANDN U2701 ( .B(B[65]), .A(n35), .Z(n2582) );
  XNOR U2702 ( .A(n2590), .B(n2692), .Z(n2583) );
  XNOR U2703 ( .A(n2589), .B(n2587), .Z(n2692) );
  AND U2704 ( .A(n2693), .B(n2694), .Z(n2587) );
  NANDN U2705 ( .A(n2695), .B(n2696), .Z(n2694) );
  OR U2706 ( .A(n2697), .B(n2698), .Z(n2696) );
  NAND U2707 ( .A(n2698), .B(n2697), .Z(n2693) );
  ANDN U2708 ( .B(B[66]), .A(n36), .Z(n2589) );
  XNOR U2709 ( .A(n2597), .B(n2699), .Z(n2590) );
  XNOR U2710 ( .A(n2596), .B(n2594), .Z(n2699) );
  AND U2711 ( .A(n2700), .B(n2701), .Z(n2594) );
  NANDN U2712 ( .A(n2702), .B(n2703), .Z(n2701) );
  NANDN U2713 ( .A(n2704), .B(n2705), .Z(n2703) );
  NANDN U2714 ( .A(n2705), .B(n2704), .Z(n2700) );
  ANDN U2715 ( .B(B[67]), .A(n37), .Z(n2596) );
  XNOR U2716 ( .A(n2604), .B(n2706), .Z(n2597) );
  XNOR U2717 ( .A(n2603), .B(n2601), .Z(n2706) );
  AND U2718 ( .A(n2707), .B(n2708), .Z(n2601) );
  NANDN U2719 ( .A(n2709), .B(n2710), .Z(n2708) );
  OR U2720 ( .A(n2711), .B(n2712), .Z(n2710) );
  NAND U2721 ( .A(n2712), .B(n2711), .Z(n2707) );
  ANDN U2722 ( .B(B[68]), .A(n38), .Z(n2603) );
  XNOR U2723 ( .A(n2611), .B(n2713), .Z(n2604) );
  XNOR U2724 ( .A(n2610), .B(n2608), .Z(n2713) );
  AND U2725 ( .A(n2714), .B(n2715), .Z(n2608) );
  NANDN U2726 ( .A(n2716), .B(n2717), .Z(n2715) );
  NANDN U2727 ( .A(n2718), .B(n2719), .Z(n2717) );
  NANDN U2728 ( .A(n2719), .B(n2718), .Z(n2714) );
  ANDN U2729 ( .B(B[69]), .A(n39), .Z(n2610) );
  XNOR U2730 ( .A(n2618), .B(n2720), .Z(n2611) );
  XNOR U2731 ( .A(n2617), .B(n2615), .Z(n2720) );
  AND U2732 ( .A(n2721), .B(n2722), .Z(n2615) );
  NANDN U2733 ( .A(n2723), .B(n2724), .Z(n2722) );
  OR U2734 ( .A(n2725), .B(n2726), .Z(n2724) );
  NAND U2735 ( .A(n2726), .B(n2725), .Z(n2721) );
  ANDN U2736 ( .B(B[70]), .A(n40), .Z(n2617) );
  XNOR U2737 ( .A(n2625), .B(n2727), .Z(n2618) );
  XNOR U2738 ( .A(n2624), .B(n2622), .Z(n2727) );
  AND U2739 ( .A(n2728), .B(n2729), .Z(n2622) );
  NANDN U2740 ( .A(n2730), .B(n2731), .Z(n2729) );
  NAND U2741 ( .A(n2732), .B(n2733), .Z(n2731) );
  ANDN U2742 ( .B(B[71]), .A(n41), .Z(n2624) );
  XOR U2743 ( .A(n2631), .B(n2734), .Z(n2625) );
  XNOR U2744 ( .A(n2629), .B(n2632), .Z(n2734) );
  NAND U2745 ( .A(A[2]), .B(B[72]), .Z(n2632) );
  NANDN U2746 ( .A(n2735), .B(n2736), .Z(n2629) );
  AND U2747 ( .A(A[0]), .B(B[73]), .Z(n2736) );
  XNOR U2748 ( .A(n2634), .B(n2737), .Z(n2631) );
  NAND U2749 ( .A(A[0]), .B(B[74]), .Z(n2737) );
  NAND U2750 ( .A(B[73]), .B(A[1]), .Z(n2634) );
  NAND U2751 ( .A(n2738), .B(n2739), .Z(n98) );
  NANDN U2752 ( .A(n2740), .B(n2741), .Z(n2739) );
  OR U2753 ( .A(n2742), .B(n2743), .Z(n2741) );
  NAND U2754 ( .A(n2743), .B(n2742), .Z(n2738) );
  XOR U2755 ( .A(n100), .B(n99), .Z(\A1[71] ) );
  XOR U2756 ( .A(n2743), .B(n2744), .Z(n99) );
  XNOR U2757 ( .A(n2742), .B(n2740), .Z(n2744) );
  AND U2758 ( .A(n2745), .B(n2746), .Z(n2740) );
  NANDN U2759 ( .A(n2747), .B(n2748), .Z(n2746) );
  NANDN U2760 ( .A(n2749), .B(n2750), .Z(n2748) );
  NANDN U2761 ( .A(n2750), .B(n2749), .Z(n2745) );
  ANDN U2762 ( .B(B[58]), .A(n29), .Z(n2742) );
  XNOR U2763 ( .A(n2649), .B(n2751), .Z(n2743) );
  XNOR U2764 ( .A(n2648), .B(n2646), .Z(n2751) );
  AND U2765 ( .A(n2752), .B(n2753), .Z(n2646) );
  NANDN U2766 ( .A(n2754), .B(n2755), .Z(n2753) );
  OR U2767 ( .A(n2756), .B(n2757), .Z(n2755) );
  NAND U2768 ( .A(n2757), .B(n2756), .Z(n2752) );
  ANDN U2769 ( .B(B[59]), .A(n30), .Z(n2648) );
  XNOR U2770 ( .A(n2656), .B(n2758), .Z(n2649) );
  XNOR U2771 ( .A(n2655), .B(n2653), .Z(n2758) );
  AND U2772 ( .A(n2759), .B(n2760), .Z(n2653) );
  NANDN U2773 ( .A(n2761), .B(n2762), .Z(n2760) );
  NANDN U2774 ( .A(n2763), .B(n2764), .Z(n2762) );
  NANDN U2775 ( .A(n2764), .B(n2763), .Z(n2759) );
  ANDN U2776 ( .B(B[60]), .A(n31), .Z(n2655) );
  XNOR U2777 ( .A(n2663), .B(n2765), .Z(n2656) );
  XNOR U2778 ( .A(n2662), .B(n2660), .Z(n2765) );
  AND U2779 ( .A(n2766), .B(n2767), .Z(n2660) );
  NANDN U2780 ( .A(n2768), .B(n2769), .Z(n2767) );
  OR U2781 ( .A(n2770), .B(n2771), .Z(n2769) );
  NAND U2782 ( .A(n2771), .B(n2770), .Z(n2766) );
  ANDN U2783 ( .B(B[61]), .A(n32), .Z(n2662) );
  XNOR U2784 ( .A(n2670), .B(n2772), .Z(n2663) );
  XNOR U2785 ( .A(n2669), .B(n2667), .Z(n2772) );
  AND U2786 ( .A(n2773), .B(n2774), .Z(n2667) );
  NANDN U2787 ( .A(n2775), .B(n2776), .Z(n2774) );
  NANDN U2788 ( .A(n2777), .B(n2778), .Z(n2776) );
  NANDN U2789 ( .A(n2778), .B(n2777), .Z(n2773) );
  ANDN U2790 ( .B(B[62]), .A(n33), .Z(n2669) );
  XNOR U2791 ( .A(n2677), .B(n2779), .Z(n2670) );
  XNOR U2792 ( .A(n2676), .B(n2674), .Z(n2779) );
  AND U2793 ( .A(n2780), .B(n2781), .Z(n2674) );
  NANDN U2794 ( .A(n2782), .B(n2783), .Z(n2781) );
  OR U2795 ( .A(n2784), .B(n2785), .Z(n2783) );
  NAND U2796 ( .A(n2785), .B(n2784), .Z(n2780) );
  ANDN U2797 ( .B(B[63]), .A(n34), .Z(n2676) );
  XNOR U2798 ( .A(n2684), .B(n2786), .Z(n2677) );
  XNOR U2799 ( .A(n2683), .B(n2681), .Z(n2786) );
  AND U2800 ( .A(n2787), .B(n2788), .Z(n2681) );
  NANDN U2801 ( .A(n2789), .B(n2790), .Z(n2788) );
  NANDN U2802 ( .A(n2791), .B(n2792), .Z(n2790) );
  NANDN U2803 ( .A(n2792), .B(n2791), .Z(n2787) );
  ANDN U2804 ( .B(B[64]), .A(n35), .Z(n2683) );
  XNOR U2805 ( .A(n2691), .B(n2793), .Z(n2684) );
  XNOR U2806 ( .A(n2690), .B(n2688), .Z(n2793) );
  AND U2807 ( .A(n2794), .B(n2795), .Z(n2688) );
  NANDN U2808 ( .A(n2796), .B(n2797), .Z(n2795) );
  OR U2809 ( .A(n2798), .B(n2799), .Z(n2797) );
  NAND U2810 ( .A(n2799), .B(n2798), .Z(n2794) );
  ANDN U2811 ( .B(B[65]), .A(n36), .Z(n2690) );
  XNOR U2812 ( .A(n2698), .B(n2800), .Z(n2691) );
  XNOR U2813 ( .A(n2697), .B(n2695), .Z(n2800) );
  AND U2814 ( .A(n2801), .B(n2802), .Z(n2695) );
  NANDN U2815 ( .A(n2803), .B(n2804), .Z(n2802) );
  NANDN U2816 ( .A(n2805), .B(n2806), .Z(n2804) );
  NANDN U2817 ( .A(n2806), .B(n2805), .Z(n2801) );
  ANDN U2818 ( .B(B[66]), .A(n37), .Z(n2697) );
  XNOR U2819 ( .A(n2705), .B(n2807), .Z(n2698) );
  XNOR U2820 ( .A(n2704), .B(n2702), .Z(n2807) );
  AND U2821 ( .A(n2808), .B(n2809), .Z(n2702) );
  NANDN U2822 ( .A(n2810), .B(n2811), .Z(n2809) );
  OR U2823 ( .A(n2812), .B(n2813), .Z(n2811) );
  NAND U2824 ( .A(n2813), .B(n2812), .Z(n2808) );
  ANDN U2825 ( .B(B[67]), .A(n38), .Z(n2704) );
  XNOR U2826 ( .A(n2712), .B(n2814), .Z(n2705) );
  XNOR U2827 ( .A(n2711), .B(n2709), .Z(n2814) );
  AND U2828 ( .A(n2815), .B(n2816), .Z(n2709) );
  NANDN U2829 ( .A(n2817), .B(n2818), .Z(n2816) );
  NANDN U2830 ( .A(n2819), .B(n2820), .Z(n2818) );
  NANDN U2831 ( .A(n2820), .B(n2819), .Z(n2815) );
  ANDN U2832 ( .B(B[68]), .A(n39), .Z(n2711) );
  XNOR U2833 ( .A(n2719), .B(n2821), .Z(n2712) );
  XNOR U2834 ( .A(n2718), .B(n2716), .Z(n2821) );
  AND U2835 ( .A(n2822), .B(n2823), .Z(n2716) );
  NANDN U2836 ( .A(n2824), .B(n2825), .Z(n2823) );
  OR U2837 ( .A(n2826), .B(n2827), .Z(n2825) );
  NAND U2838 ( .A(n2827), .B(n2826), .Z(n2822) );
  ANDN U2839 ( .B(B[69]), .A(n40), .Z(n2718) );
  XNOR U2840 ( .A(n2726), .B(n2828), .Z(n2719) );
  XNOR U2841 ( .A(n2725), .B(n2723), .Z(n2828) );
  AND U2842 ( .A(n2829), .B(n2830), .Z(n2723) );
  NANDN U2843 ( .A(n2831), .B(n2832), .Z(n2830) );
  NAND U2844 ( .A(n2833), .B(n2834), .Z(n2832) );
  ANDN U2845 ( .B(B[70]), .A(n41), .Z(n2725) );
  XOR U2846 ( .A(n2732), .B(n2835), .Z(n2726) );
  XNOR U2847 ( .A(n2730), .B(n2733), .Z(n2835) );
  NAND U2848 ( .A(A[2]), .B(B[71]), .Z(n2733) );
  NANDN U2849 ( .A(n2836), .B(n2837), .Z(n2730) );
  AND U2850 ( .A(A[0]), .B(B[72]), .Z(n2837) );
  XNOR U2851 ( .A(n2735), .B(n2838), .Z(n2732) );
  NAND U2852 ( .A(A[0]), .B(B[73]), .Z(n2838) );
  NAND U2853 ( .A(B[72]), .B(A[1]), .Z(n2735) );
  NAND U2854 ( .A(n2839), .B(n2840), .Z(n100) );
  NANDN U2855 ( .A(n2841), .B(n2842), .Z(n2840) );
  OR U2856 ( .A(n2843), .B(n2844), .Z(n2842) );
  NAND U2857 ( .A(n2844), .B(n2843), .Z(n2839) );
  XOR U2858 ( .A(n102), .B(n101), .Z(\A1[70] ) );
  XOR U2859 ( .A(n2844), .B(n2845), .Z(n101) );
  XNOR U2860 ( .A(n2843), .B(n2841), .Z(n2845) );
  AND U2861 ( .A(n2846), .B(n2847), .Z(n2841) );
  NANDN U2862 ( .A(n2848), .B(n2849), .Z(n2847) );
  NANDN U2863 ( .A(n2850), .B(n2851), .Z(n2849) );
  NANDN U2864 ( .A(n2851), .B(n2850), .Z(n2846) );
  ANDN U2865 ( .B(B[57]), .A(n29), .Z(n2843) );
  XNOR U2866 ( .A(n2750), .B(n2852), .Z(n2844) );
  XNOR U2867 ( .A(n2749), .B(n2747), .Z(n2852) );
  AND U2868 ( .A(n2853), .B(n2854), .Z(n2747) );
  NANDN U2869 ( .A(n2855), .B(n2856), .Z(n2854) );
  OR U2870 ( .A(n2857), .B(n2858), .Z(n2856) );
  NAND U2871 ( .A(n2858), .B(n2857), .Z(n2853) );
  ANDN U2872 ( .B(B[58]), .A(n30), .Z(n2749) );
  XNOR U2873 ( .A(n2757), .B(n2859), .Z(n2750) );
  XNOR U2874 ( .A(n2756), .B(n2754), .Z(n2859) );
  AND U2875 ( .A(n2860), .B(n2861), .Z(n2754) );
  NANDN U2876 ( .A(n2862), .B(n2863), .Z(n2861) );
  NANDN U2877 ( .A(n2864), .B(n2865), .Z(n2863) );
  NANDN U2878 ( .A(n2865), .B(n2864), .Z(n2860) );
  ANDN U2879 ( .B(B[59]), .A(n31), .Z(n2756) );
  XNOR U2880 ( .A(n2764), .B(n2866), .Z(n2757) );
  XNOR U2881 ( .A(n2763), .B(n2761), .Z(n2866) );
  AND U2882 ( .A(n2867), .B(n2868), .Z(n2761) );
  NANDN U2883 ( .A(n2869), .B(n2870), .Z(n2868) );
  OR U2884 ( .A(n2871), .B(n2872), .Z(n2870) );
  NAND U2885 ( .A(n2872), .B(n2871), .Z(n2867) );
  ANDN U2886 ( .B(B[60]), .A(n32), .Z(n2763) );
  XNOR U2887 ( .A(n2771), .B(n2873), .Z(n2764) );
  XNOR U2888 ( .A(n2770), .B(n2768), .Z(n2873) );
  AND U2889 ( .A(n2874), .B(n2875), .Z(n2768) );
  NANDN U2890 ( .A(n2876), .B(n2877), .Z(n2875) );
  NANDN U2891 ( .A(n2878), .B(n2879), .Z(n2877) );
  NANDN U2892 ( .A(n2879), .B(n2878), .Z(n2874) );
  ANDN U2893 ( .B(B[61]), .A(n33), .Z(n2770) );
  XNOR U2894 ( .A(n2778), .B(n2880), .Z(n2771) );
  XNOR U2895 ( .A(n2777), .B(n2775), .Z(n2880) );
  AND U2896 ( .A(n2881), .B(n2882), .Z(n2775) );
  NANDN U2897 ( .A(n2883), .B(n2884), .Z(n2882) );
  OR U2898 ( .A(n2885), .B(n2886), .Z(n2884) );
  NAND U2899 ( .A(n2886), .B(n2885), .Z(n2881) );
  ANDN U2900 ( .B(B[62]), .A(n34), .Z(n2777) );
  XNOR U2901 ( .A(n2785), .B(n2887), .Z(n2778) );
  XNOR U2902 ( .A(n2784), .B(n2782), .Z(n2887) );
  AND U2903 ( .A(n2888), .B(n2889), .Z(n2782) );
  NANDN U2904 ( .A(n2890), .B(n2891), .Z(n2889) );
  NANDN U2905 ( .A(n2892), .B(n2893), .Z(n2891) );
  NANDN U2906 ( .A(n2893), .B(n2892), .Z(n2888) );
  ANDN U2907 ( .B(B[63]), .A(n35), .Z(n2784) );
  XNOR U2908 ( .A(n2792), .B(n2894), .Z(n2785) );
  XNOR U2909 ( .A(n2791), .B(n2789), .Z(n2894) );
  AND U2910 ( .A(n2895), .B(n2896), .Z(n2789) );
  NANDN U2911 ( .A(n2897), .B(n2898), .Z(n2896) );
  OR U2912 ( .A(n2899), .B(n2900), .Z(n2898) );
  NAND U2913 ( .A(n2900), .B(n2899), .Z(n2895) );
  ANDN U2914 ( .B(B[64]), .A(n36), .Z(n2791) );
  XNOR U2915 ( .A(n2799), .B(n2901), .Z(n2792) );
  XNOR U2916 ( .A(n2798), .B(n2796), .Z(n2901) );
  AND U2917 ( .A(n2902), .B(n2903), .Z(n2796) );
  NANDN U2918 ( .A(n2904), .B(n2905), .Z(n2903) );
  NANDN U2919 ( .A(n2906), .B(n2907), .Z(n2905) );
  NANDN U2920 ( .A(n2907), .B(n2906), .Z(n2902) );
  ANDN U2921 ( .B(B[65]), .A(n37), .Z(n2798) );
  XNOR U2922 ( .A(n2806), .B(n2908), .Z(n2799) );
  XNOR U2923 ( .A(n2805), .B(n2803), .Z(n2908) );
  AND U2924 ( .A(n2909), .B(n2910), .Z(n2803) );
  NANDN U2925 ( .A(n2911), .B(n2912), .Z(n2910) );
  OR U2926 ( .A(n2913), .B(n2914), .Z(n2912) );
  NAND U2927 ( .A(n2914), .B(n2913), .Z(n2909) );
  ANDN U2928 ( .B(B[66]), .A(n38), .Z(n2805) );
  XNOR U2929 ( .A(n2813), .B(n2915), .Z(n2806) );
  XNOR U2930 ( .A(n2812), .B(n2810), .Z(n2915) );
  AND U2931 ( .A(n2916), .B(n2917), .Z(n2810) );
  NANDN U2932 ( .A(n2918), .B(n2919), .Z(n2917) );
  NANDN U2933 ( .A(n2920), .B(n2921), .Z(n2919) );
  NANDN U2934 ( .A(n2921), .B(n2920), .Z(n2916) );
  ANDN U2935 ( .B(B[67]), .A(n39), .Z(n2812) );
  XNOR U2936 ( .A(n2820), .B(n2922), .Z(n2813) );
  XNOR U2937 ( .A(n2819), .B(n2817), .Z(n2922) );
  AND U2938 ( .A(n2923), .B(n2924), .Z(n2817) );
  NANDN U2939 ( .A(n2925), .B(n2926), .Z(n2924) );
  OR U2940 ( .A(n2927), .B(n2928), .Z(n2926) );
  NAND U2941 ( .A(n2928), .B(n2927), .Z(n2923) );
  ANDN U2942 ( .B(B[68]), .A(n40), .Z(n2819) );
  XNOR U2943 ( .A(n2827), .B(n2929), .Z(n2820) );
  XNOR U2944 ( .A(n2826), .B(n2824), .Z(n2929) );
  AND U2945 ( .A(n2930), .B(n2931), .Z(n2824) );
  NANDN U2946 ( .A(n2932), .B(n2933), .Z(n2931) );
  NAND U2947 ( .A(n2934), .B(n2935), .Z(n2933) );
  ANDN U2948 ( .B(B[69]), .A(n41), .Z(n2826) );
  XOR U2949 ( .A(n2833), .B(n2936), .Z(n2827) );
  XNOR U2950 ( .A(n2831), .B(n2834), .Z(n2936) );
  NAND U2951 ( .A(A[2]), .B(B[70]), .Z(n2834) );
  NANDN U2952 ( .A(n2937), .B(n2938), .Z(n2831) );
  AND U2953 ( .A(A[0]), .B(B[71]), .Z(n2938) );
  XNOR U2954 ( .A(n2836), .B(n2939), .Z(n2833) );
  NAND U2955 ( .A(A[0]), .B(B[72]), .Z(n2939) );
  NAND U2956 ( .A(B[71]), .B(A[1]), .Z(n2836) );
  NAND U2957 ( .A(n2940), .B(n2941), .Z(n102) );
  NANDN U2958 ( .A(n2942), .B(n2943), .Z(n2941) );
  OR U2959 ( .A(n2944), .B(n2945), .Z(n2943) );
  NAND U2960 ( .A(n2945), .B(n2944), .Z(n2940) );
  XNOR U2961 ( .A(n2946), .B(n2947), .Z(\A1[6] ) );
  XNOR U2962 ( .A(n2948), .B(n2949), .Z(n2947) );
  XOR U2963 ( .A(n104), .B(n103), .Z(\A1[69] ) );
  XOR U2964 ( .A(n2945), .B(n2950), .Z(n103) );
  XNOR U2965 ( .A(n2944), .B(n2942), .Z(n2950) );
  AND U2966 ( .A(n2951), .B(n2952), .Z(n2942) );
  NANDN U2967 ( .A(n2953), .B(n2954), .Z(n2952) );
  NANDN U2968 ( .A(n2955), .B(n2956), .Z(n2954) );
  NANDN U2969 ( .A(n2956), .B(n2955), .Z(n2951) );
  ANDN U2970 ( .B(B[56]), .A(n29), .Z(n2944) );
  XNOR U2971 ( .A(n2851), .B(n2957), .Z(n2945) );
  XNOR U2972 ( .A(n2850), .B(n2848), .Z(n2957) );
  AND U2973 ( .A(n2958), .B(n2959), .Z(n2848) );
  NANDN U2974 ( .A(n2960), .B(n2961), .Z(n2959) );
  OR U2975 ( .A(n2962), .B(n2963), .Z(n2961) );
  NAND U2976 ( .A(n2963), .B(n2962), .Z(n2958) );
  ANDN U2977 ( .B(B[57]), .A(n30), .Z(n2850) );
  XNOR U2978 ( .A(n2858), .B(n2964), .Z(n2851) );
  XNOR U2979 ( .A(n2857), .B(n2855), .Z(n2964) );
  AND U2980 ( .A(n2965), .B(n2966), .Z(n2855) );
  NANDN U2981 ( .A(n2967), .B(n2968), .Z(n2966) );
  NANDN U2982 ( .A(n2969), .B(n2970), .Z(n2968) );
  NANDN U2983 ( .A(n2970), .B(n2969), .Z(n2965) );
  ANDN U2984 ( .B(B[58]), .A(n31), .Z(n2857) );
  XNOR U2985 ( .A(n2865), .B(n2971), .Z(n2858) );
  XNOR U2986 ( .A(n2864), .B(n2862), .Z(n2971) );
  AND U2987 ( .A(n2972), .B(n2973), .Z(n2862) );
  NANDN U2988 ( .A(n2974), .B(n2975), .Z(n2973) );
  OR U2989 ( .A(n2976), .B(n2977), .Z(n2975) );
  NAND U2990 ( .A(n2977), .B(n2976), .Z(n2972) );
  ANDN U2991 ( .B(B[59]), .A(n32), .Z(n2864) );
  XNOR U2992 ( .A(n2872), .B(n2978), .Z(n2865) );
  XNOR U2993 ( .A(n2871), .B(n2869), .Z(n2978) );
  AND U2994 ( .A(n2979), .B(n2980), .Z(n2869) );
  NANDN U2995 ( .A(n2981), .B(n2982), .Z(n2980) );
  NANDN U2996 ( .A(n2983), .B(n2984), .Z(n2982) );
  NANDN U2997 ( .A(n2984), .B(n2983), .Z(n2979) );
  ANDN U2998 ( .B(B[60]), .A(n33), .Z(n2871) );
  XNOR U2999 ( .A(n2879), .B(n2985), .Z(n2872) );
  XNOR U3000 ( .A(n2878), .B(n2876), .Z(n2985) );
  AND U3001 ( .A(n2986), .B(n2987), .Z(n2876) );
  NANDN U3002 ( .A(n2988), .B(n2989), .Z(n2987) );
  OR U3003 ( .A(n2990), .B(n2991), .Z(n2989) );
  NAND U3004 ( .A(n2991), .B(n2990), .Z(n2986) );
  ANDN U3005 ( .B(B[61]), .A(n34), .Z(n2878) );
  XNOR U3006 ( .A(n2886), .B(n2992), .Z(n2879) );
  XNOR U3007 ( .A(n2885), .B(n2883), .Z(n2992) );
  AND U3008 ( .A(n2993), .B(n2994), .Z(n2883) );
  NANDN U3009 ( .A(n2995), .B(n2996), .Z(n2994) );
  NANDN U3010 ( .A(n2997), .B(n2998), .Z(n2996) );
  NANDN U3011 ( .A(n2998), .B(n2997), .Z(n2993) );
  ANDN U3012 ( .B(B[62]), .A(n35), .Z(n2885) );
  XNOR U3013 ( .A(n2893), .B(n2999), .Z(n2886) );
  XNOR U3014 ( .A(n2892), .B(n2890), .Z(n2999) );
  AND U3015 ( .A(n3000), .B(n3001), .Z(n2890) );
  NANDN U3016 ( .A(n3002), .B(n3003), .Z(n3001) );
  OR U3017 ( .A(n3004), .B(n3005), .Z(n3003) );
  NAND U3018 ( .A(n3005), .B(n3004), .Z(n3000) );
  ANDN U3019 ( .B(B[63]), .A(n36), .Z(n2892) );
  XNOR U3020 ( .A(n2900), .B(n3006), .Z(n2893) );
  XNOR U3021 ( .A(n2899), .B(n2897), .Z(n3006) );
  AND U3022 ( .A(n3007), .B(n3008), .Z(n2897) );
  NANDN U3023 ( .A(n3009), .B(n3010), .Z(n3008) );
  NANDN U3024 ( .A(n3011), .B(n3012), .Z(n3010) );
  NANDN U3025 ( .A(n3012), .B(n3011), .Z(n3007) );
  ANDN U3026 ( .B(B[64]), .A(n37), .Z(n2899) );
  XNOR U3027 ( .A(n2907), .B(n3013), .Z(n2900) );
  XNOR U3028 ( .A(n2906), .B(n2904), .Z(n3013) );
  AND U3029 ( .A(n3014), .B(n3015), .Z(n2904) );
  NANDN U3030 ( .A(n3016), .B(n3017), .Z(n3015) );
  OR U3031 ( .A(n3018), .B(n3019), .Z(n3017) );
  NAND U3032 ( .A(n3019), .B(n3018), .Z(n3014) );
  ANDN U3033 ( .B(B[65]), .A(n38), .Z(n2906) );
  XNOR U3034 ( .A(n2914), .B(n3020), .Z(n2907) );
  XNOR U3035 ( .A(n2913), .B(n2911), .Z(n3020) );
  AND U3036 ( .A(n3021), .B(n3022), .Z(n2911) );
  NANDN U3037 ( .A(n3023), .B(n3024), .Z(n3022) );
  NANDN U3038 ( .A(n3025), .B(n3026), .Z(n3024) );
  NANDN U3039 ( .A(n3026), .B(n3025), .Z(n3021) );
  ANDN U3040 ( .B(B[66]), .A(n39), .Z(n2913) );
  XNOR U3041 ( .A(n2921), .B(n3027), .Z(n2914) );
  XNOR U3042 ( .A(n2920), .B(n2918), .Z(n3027) );
  AND U3043 ( .A(n3028), .B(n3029), .Z(n2918) );
  NANDN U3044 ( .A(n3030), .B(n3031), .Z(n3029) );
  OR U3045 ( .A(n3032), .B(n3033), .Z(n3031) );
  NAND U3046 ( .A(n3033), .B(n3032), .Z(n3028) );
  ANDN U3047 ( .B(B[67]), .A(n40), .Z(n2920) );
  XNOR U3048 ( .A(n2928), .B(n3034), .Z(n2921) );
  XNOR U3049 ( .A(n2927), .B(n2925), .Z(n3034) );
  AND U3050 ( .A(n3035), .B(n3036), .Z(n2925) );
  NANDN U3051 ( .A(n3037), .B(n3038), .Z(n3036) );
  NAND U3052 ( .A(n3039), .B(n3040), .Z(n3038) );
  ANDN U3053 ( .B(B[68]), .A(n41), .Z(n2927) );
  XOR U3054 ( .A(n2934), .B(n3041), .Z(n2928) );
  XNOR U3055 ( .A(n2932), .B(n2935), .Z(n3041) );
  NAND U3056 ( .A(A[2]), .B(B[69]), .Z(n2935) );
  NANDN U3057 ( .A(n3042), .B(n3043), .Z(n2932) );
  AND U3058 ( .A(A[0]), .B(B[70]), .Z(n3043) );
  XNOR U3059 ( .A(n2937), .B(n3044), .Z(n2934) );
  NAND U3060 ( .A(A[0]), .B(B[71]), .Z(n3044) );
  NAND U3061 ( .A(B[70]), .B(A[1]), .Z(n2937) );
  NAND U3062 ( .A(n3045), .B(n3046), .Z(n104) );
  NANDN U3063 ( .A(n3047), .B(n3048), .Z(n3046) );
  OR U3064 ( .A(n3049), .B(n3050), .Z(n3048) );
  NAND U3065 ( .A(n3050), .B(n3049), .Z(n3045) );
  XOR U3066 ( .A(n106), .B(n105), .Z(\A1[68] ) );
  XOR U3067 ( .A(n3050), .B(n3051), .Z(n105) );
  XNOR U3068 ( .A(n3049), .B(n3047), .Z(n3051) );
  AND U3069 ( .A(n3052), .B(n3053), .Z(n3047) );
  NANDN U3070 ( .A(n3054), .B(n3055), .Z(n3053) );
  NANDN U3071 ( .A(n3056), .B(n3057), .Z(n3055) );
  NANDN U3072 ( .A(n3057), .B(n3056), .Z(n3052) );
  ANDN U3073 ( .B(B[55]), .A(n29), .Z(n3049) );
  XNOR U3074 ( .A(n2956), .B(n3058), .Z(n3050) );
  XNOR U3075 ( .A(n2955), .B(n2953), .Z(n3058) );
  AND U3076 ( .A(n3059), .B(n3060), .Z(n2953) );
  NANDN U3077 ( .A(n3061), .B(n3062), .Z(n3060) );
  OR U3078 ( .A(n3063), .B(n3064), .Z(n3062) );
  NAND U3079 ( .A(n3064), .B(n3063), .Z(n3059) );
  ANDN U3080 ( .B(B[56]), .A(n30), .Z(n2955) );
  XNOR U3081 ( .A(n2963), .B(n3065), .Z(n2956) );
  XNOR U3082 ( .A(n2962), .B(n2960), .Z(n3065) );
  AND U3083 ( .A(n3066), .B(n3067), .Z(n2960) );
  NANDN U3084 ( .A(n3068), .B(n3069), .Z(n3067) );
  NANDN U3085 ( .A(n3070), .B(n3071), .Z(n3069) );
  NANDN U3086 ( .A(n3071), .B(n3070), .Z(n3066) );
  ANDN U3087 ( .B(B[57]), .A(n31), .Z(n2962) );
  XNOR U3088 ( .A(n2970), .B(n3072), .Z(n2963) );
  XNOR U3089 ( .A(n2969), .B(n2967), .Z(n3072) );
  AND U3090 ( .A(n3073), .B(n3074), .Z(n2967) );
  NANDN U3091 ( .A(n3075), .B(n3076), .Z(n3074) );
  OR U3092 ( .A(n3077), .B(n3078), .Z(n3076) );
  NAND U3093 ( .A(n3078), .B(n3077), .Z(n3073) );
  ANDN U3094 ( .B(B[58]), .A(n32), .Z(n2969) );
  XNOR U3095 ( .A(n2977), .B(n3079), .Z(n2970) );
  XNOR U3096 ( .A(n2976), .B(n2974), .Z(n3079) );
  AND U3097 ( .A(n3080), .B(n3081), .Z(n2974) );
  NANDN U3098 ( .A(n3082), .B(n3083), .Z(n3081) );
  NANDN U3099 ( .A(n3084), .B(n3085), .Z(n3083) );
  NANDN U3100 ( .A(n3085), .B(n3084), .Z(n3080) );
  ANDN U3101 ( .B(B[59]), .A(n33), .Z(n2976) );
  XNOR U3102 ( .A(n2984), .B(n3086), .Z(n2977) );
  XNOR U3103 ( .A(n2983), .B(n2981), .Z(n3086) );
  AND U3104 ( .A(n3087), .B(n3088), .Z(n2981) );
  NANDN U3105 ( .A(n3089), .B(n3090), .Z(n3088) );
  OR U3106 ( .A(n3091), .B(n3092), .Z(n3090) );
  NAND U3107 ( .A(n3092), .B(n3091), .Z(n3087) );
  ANDN U3108 ( .B(B[60]), .A(n34), .Z(n2983) );
  XNOR U3109 ( .A(n2991), .B(n3093), .Z(n2984) );
  XNOR U3110 ( .A(n2990), .B(n2988), .Z(n3093) );
  AND U3111 ( .A(n3094), .B(n3095), .Z(n2988) );
  NANDN U3112 ( .A(n3096), .B(n3097), .Z(n3095) );
  NANDN U3113 ( .A(n3098), .B(n3099), .Z(n3097) );
  NANDN U3114 ( .A(n3099), .B(n3098), .Z(n3094) );
  ANDN U3115 ( .B(B[61]), .A(n35), .Z(n2990) );
  XNOR U3116 ( .A(n2998), .B(n3100), .Z(n2991) );
  XNOR U3117 ( .A(n2997), .B(n2995), .Z(n3100) );
  AND U3118 ( .A(n3101), .B(n3102), .Z(n2995) );
  NANDN U3119 ( .A(n3103), .B(n3104), .Z(n3102) );
  OR U3120 ( .A(n3105), .B(n3106), .Z(n3104) );
  NAND U3121 ( .A(n3106), .B(n3105), .Z(n3101) );
  ANDN U3122 ( .B(B[62]), .A(n36), .Z(n2997) );
  XNOR U3123 ( .A(n3005), .B(n3107), .Z(n2998) );
  XNOR U3124 ( .A(n3004), .B(n3002), .Z(n3107) );
  AND U3125 ( .A(n3108), .B(n3109), .Z(n3002) );
  NANDN U3126 ( .A(n3110), .B(n3111), .Z(n3109) );
  NANDN U3127 ( .A(n3112), .B(n3113), .Z(n3111) );
  NANDN U3128 ( .A(n3113), .B(n3112), .Z(n3108) );
  ANDN U3129 ( .B(B[63]), .A(n37), .Z(n3004) );
  XNOR U3130 ( .A(n3012), .B(n3114), .Z(n3005) );
  XNOR U3131 ( .A(n3011), .B(n3009), .Z(n3114) );
  AND U3132 ( .A(n3115), .B(n3116), .Z(n3009) );
  NANDN U3133 ( .A(n3117), .B(n3118), .Z(n3116) );
  OR U3134 ( .A(n3119), .B(n3120), .Z(n3118) );
  NAND U3135 ( .A(n3120), .B(n3119), .Z(n3115) );
  ANDN U3136 ( .B(B[64]), .A(n38), .Z(n3011) );
  XNOR U3137 ( .A(n3019), .B(n3121), .Z(n3012) );
  XNOR U3138 ( .A(n3018), .B(n3016), .Z(n3121) );
  AND U3139 ( .A(n3122), .B(n3123), .Z(n3016) );
  NANDN U3140 ( .A(n3124), .B(n3125), .Z(n3123) );
  NANDN U3141 ( .A(n3126), .B(n3127), .Z(n3125) );
  NANDN U3142 ( .A(n3127), .B(n3126), .Z(n3122) );
  ANDN U3143 ( .B(B[65]), .A(n39), .Z(n3018) );
  XNOR U3144 ( .A(n3026), .B(n3128), .Z(n3019) );
  XNOR U3145 ( .A(n3025), .B(n3023), .Z(n3128) );
  AND U3146 ( .A(n3129), .B(n3130), .Z(n3023) );
  NANDN U3147 ( .A(n3131), .B(n3132), .Z(n3130) );
  OR U3148 ( .A(n3133), .B(n3134), .Z(n3132) );
  NAND U3149 ( .A(n3134), .B(n3133), .Z(n3129) );
  ANDN U3150 ( .B(B[66]), .A(n40), .Z(n3025) );
  XNOR U3151 ( .A(n3033), .B(n3135), .Z(n3026) );
  XNOR U3152 ( .A(n3032), .B(n3030), .Z(n3135) );
  AND U3153 ( .A(n3136), .B(n3137), .Z(n3030) );
  NANDN U3154 ( .A(n3138), .B(n3139), .Z(n3137) );
  NAND U3155 ( .A(n3140), .B(n3141), .Z(n3139) );
  ANDN U3156 ( .B(B[67]), .A(n41), .Z(n3032) );
  XOR U3157 ( .A(n3039), .B(n3142), .Z(n3033) );
  XNOR U3158 ( .A(n3037), .B(n3040), .Z(n3142) );
  NAND U3159 ( .A(A[2]), .B(B[68]), .Z(n3040) );
  NANDN U3160 ( .A(n3143), .B(n3144), .Z(n3037) );
  AND U3161 ( .A(A[0]), .B(B[69]), .Z(n3144) );
  XNOR U3162 ( .A(n3042), .B(n3145), .Z(n3039) );
  NAND U3163 ( .A(A[0]), .B(B[70]), .Z(n3145) );
  NAND U3164 ( .A(B[69]), .B(A[1]), .Z(n3042) );
  NAND U3165 ( .A(n3146), .B(n3147), .Z(n106) );
  NANDN U3166 ( .A(n3148), .B(n3149), .Z(n3147) );
  OR U3167 ( .A(n3150), .B(n3151), .Z(n3149) );
  NAND U3168 ( .A(n3151), .B(n3150), .Z(n3146) );
  XOR U3169 ( .A(n108), .B(n107), .Z(\A1[67] ) );
  XOR U3170 ( .A(n3151), .B(n3152), .Z(n107) );
  XNOR U3171 ( .A(n3150), .B(n3148), .Z(n3152) );
  AND U3172 ( .A(n3153), .B(n3154), .Z(n3148) );
  NANDN U3173 ( .A(n3155), .B(n3156), .Z(n3154) );
  NANDN U3174 ( .A(n3157), .B(n3158), .Z(n3156) );
  NANDN U3175 ( .A(n3158), .B(n3157), .Z(n3153) );
  ANDN U3176 ( .B(B[54]), .A(n29), .Z(n3150) );
  XNOR U3177 ( .A(n3057), .B(n3159), .Z(n3151) );
  XNOR U3178 ( .A(n3056), .B(n3054), .Z(n3159) );
  AND U3179 ( .A(n3160), .B(n3161), .Z(n3054) );
  NANDN U3180 ( .A(n3162), .B(n3163), .Z(n3161) );
  OR U3181 ( .A(n3164), .B(n3165), .Z(n3163) );
  NAND U3182 ( .A(n3165), .B(n3164), .Z(n3160) );
  ANDN U3183 ( .B(B[55]), .A(n30), .Z(n3056) );
  XNOR U3184 ( .A(n3064), .B(n3166), .Z(n3057) );
  XNOR U3185 ( .A(n3063), .B(n3061), .Z(n3166) );
  AND U3186 ( .A(n3167), .B(n3168), .Z(n3061) );
  NANDN U3187 ( .A(n3169), .B(n3170), .Z(n3168) );
  NANDN U3188 ( .A(n3171), .B(n3172), .Z(n3170) );
  NANDN U3189 ( .A(n3172), .B(n3171), .Z(n3167) );
  ANDN U3190 ( .B(B[56]), .A(n31), .Z(n3063) );
  XNOR U3191 ( .A(n3071), .B(n3173), .Z(n3064) );
  XNOR U3192 ( .A(n3070), .B(n3068), .Z(n3173) );
  AND U3193 ( .A(n3174), .B(n3175), .Z(n3068) );
  NANDN U3194 ( .A(n3176), .B(n3177), .Z(n3175) );
  OR U3195 ( .A(n3178), .B(n3179), .Z(n3177) );
  NAND U3196 ( .A(n3179), .B(n3178), .Z(n3174) );
  ANDN U3197 ( .B(B[57]), .A(n32), .Z(n3070) );
  XNOR U3198 ( .A(n3078), .B(n3180), .Z(n3071) );
  XNOR U3199 ( .A(n3077), .B(n3075), .Z(n3180) );
  AND U3200 ( .A(n3181), .B(n3182), .Z(n3075) );
  NANDN U3201 ( .A(n3183), .B(n3184), .Z(n3182) );
  NANDN U3202 ( .A(n3185), .B(n3186), .Z(n3184) );
  NANDN U3203 ( .A(n3186), .B(n3185), .Z(n3181) );
  ANDN U3204 ( .B(B[58]), .A(n33), .Z(n3077) );
  XNOR U3205 ( .A(n3085), .B(n3187), .Z(n3078) );
  XNOR U3206 ( .A(n3084), .B(n3082), .Z(n3187) );
  AND U3207 ( .A(n3188), .B(n3189), .Z(n3082) );
  NANDN U3208 ( .A(n3190), .B(n3191), .Z(n3189) );
  OR U3209 ( .A(n3192), .B(n3193), .Z(n3191) );
  NAND U3210 ( .A(n3193), .B(n3192), .Z(n3188) );
  ANDN U3211 ( .B(B[59]), .A(n34), .Z(n3084) );
  XNOR U3212 ( .A(n3092), .B(n3194), .Z(n3085) );
  XNOR U3213 ( .A(n3091), .B(n3089), .Z(n3194) );
  AND U3214 ( .A(n3195), .B(n3196), .Z(n3089) );
  NANDN U3215 ( .A(n3197), .B(n3198), .Z(n3196) );
  NANDN U3216 ( .A(n3199), .B(n3200), .Z(n3198) );
  NANDN U3217 ( .A(n3200), .B(n3199), .Z(n3195) );
  ANDN U3218 ( .B(B[60]), .A(n35), .Z(n3091) );
  XNOR U3219 ( .A(n3099), .B(n3201), .Z(n3092) );
  XNOR U3220 ( .A(n3098), .B(n3096), .Z(n3201) );
  AND U3221 ( .A(n3202), .B(n3203), .Z(n3096) );
  NANDN U3222 ( .A(n3204), .B(n3205), .Z(n3203) );
  OR U3223 ( .A(n3206), .B(n3207), .Z(n3205) );
  NAND U3224 ( .A(n3207), .B(n3206), .Z(n3202) );
  ANDN U3225 ( .B(B[61]), .A(n36), .Z(n3098) );
  XNOR U3226 ( .A(n3106), .B(n3208), .Z(n3099) );
  XNOR U3227 ( .A(n3105), .B(n3103), .Z(n3208) );
  AND U3228 ( .A(n3209), .B(n3210), .Z(n3103) );
  NANDN U3229 ( .A(n3211), .B(n3212), .Z(n3210) );
  NANDN U3230 ( .A(n3213), .B(n3214), .Z(n3212) );
  NANDN U3231 ( .A(n3214), .B(n3213), .Z(n3209) );
  ANDN U3232 ( .B(B[62]), .A(n37), .Z(n3105) );
  XNOR U3233 ( .A(n3113), .B(n3215), .Z(n3106) );
  XNOR U3234 ( .A(n3112), .B(n3110), .Z(n3215) );
  AND U3235 ( .A(n3216), .B(n3217), .Z(n3110) );
  NANDN U3236 ( .A(n3218), .B(n3219), .Z(n3217) );
  OR U3237 ( .A(n3220), .B(n3221), .Z(n3219) );
  NAND U3238 ( .A(n3221), .B(n3220), .Z(n3216) );
  ANDN U3239 ( .B(B[63]), .A(n38), .Z(n3112) );
  XNOR U3240 ( .A(n3120), .B(n3222), .Z(n3113) );
  XNOR U3241 ( .A(n3119), .B(n3117), .Z(n3222) );
  AND U3242 ( .A(n3223), .B(n3224), .Z(n3117) );
  NANDN U3243 ( .A(n3225), .B(n3226), .Z(n3224) );
  NANDN U3244 ( .A(n3227), .B(n3228), .Z(n3226) );
  NANDN U3245 ( .A(n3228), .B(n3227), .Z(n3223) );
  ANDN U3246 ( .B(B[64]), .A(n39), .Z(n3119) );
  XNOR U3247 ( .A(n3127), .B(n3229), .Z(n3120) );
  XNOR U3248 ( .A(n3126), .B(n3124), .Z(n3229) );
  AND U3249 ( .A(n3230), .B(n3231), .Z(n3124) );
  NANDN U3250 ( .A(n3232), .B(n3233), .Z(n3231) );
  OR U3251 ( .A(n3234), .B(n3235), .Z(n3233) );
  NAND U3252 ( .A(n3235), .B(n3234), .Z(n3230) );
  ANDN U3253 ( .B(B[65]), .A(n40), .Z(n3126) );
  XNOR U3254 ( .A(n3134), .B(n3236), .Z(n3127) );
  XNOR U3255 ( .A(n3133), .B(n3131), .Z(n3236) );
  AND U3256 ( .A(n3237), .B(n3238), .Z(n3131) );
  NANDN U3257 ( .A(n3239), .B(n3240), .Z(n3238) );
  NAND U3258 ( .A(n3241), .B(n3242), .Z(n3240) );
  ANDN U3259 ( .B(B[66]), .A(n41), .Z(n3133) );
  XOR U3260 ( .A(n3140), .B(n3243), .Z(n3134) );
  XNOR U3261 ( .A(n3138), .B(n3141), .Z(n3243) );
  NAND U3262 ( .A(A[2]), .B(B[67]), .Z(n3141) );
  NANDN U3263 ( .A(n3244), .B(n3245), .Z(n3138) );
  AND U3264 ( .A(A[0]), .B(B[68]), .Z(n3245) );
  XNOR U3265 ( .A(n3143), .B(n3246), .Z(n3140) );
  NAND U3266 ( .A(A[0]), .B(B[69]), .Z(n3246) );
  NAND U3267 ( .A(B[68]), .B(A[1]), .Z(n3143) );
  NAND U3268 ( .A(n3247), .B(n3248), .Z(n108) );
  NANDN U3269 ( .A(n3249), .B(n3250), .Z(n3248) );
  OR U3270 ( .A(n3251), .B(n3252), .Z(n3250) );
  NAND U3271 ( .A(n3252), .B(n3251), .Z(n3247) );
  XOR U3272 ( .A(n110), .B(n109), .Z(\A1[66] ) );
  XOR U3273 ( .A(n3252), .B(n3253), .Z(n109) );
  XNOR U3274 ( .A(n3251), .B(n3249), .Z(n3253) );
  AND U3275 ( .A(n3254), .B(n3255), .Z(n3249) );
  NANDN U3276 ( .A(n3256), .B(n3257), .Z(n3255) );
  NANDN U3277 ( .A(n3258), .B(n3259), .Z(n3257) );
  NANDN U3278 ( .A(n3259), .B(n3258), .Z(n3254) );
  ANDN U3279 ( .B(B[53]), .A(n29), .Z(n3251) );
  XNOR U3280 ( .A(n3158), .B(n3260), .Z(n3252) );
  XNOR U3281 ( .A(n3157), .B(n3155), .Z(n3260) );
  AND U3282 ( .A(n3261), .B(n3262), .Z(n3155) );
  NANDN U3283 ( .A(n3263), .B(n3264), .Z(n3262) );
  OR U3284 ( .A(n3265), .B(n3266), .Z(n3264) );
  NAND U3285 ( .A(n3266), .B(n3265), .Z(n3261) );
  ANDN U3286 ( .B(B[54]), .A(n30), .Z(n3157) );
  XNOR U3287 ( .A(n3165), .B(n3267), .Z(n3158) );
  XNOR U3288 ( .A(n3164), .B(n3162), .Z(n3267) );
  AND U3289 ( .A(n3268), .B(n3269), .Z(n3162) );
  NANDN U3290 ( .A(n3270), .B(n3271), .Z(n3269) );
  NANDN U3291 ( .A(n3272), .B(n3273), .Z(n3271) );
  NANDN U3292 ( .A(n3273), .B(n3272), .Z(n3268) );
  ANDN U3293 ( .B(B[55]), .A(n31), .Z(n3164) );
  XNOR U3294 ( .A(n3172), .B(n3274), .Z(n3165) );
  XNOR U3295 ( .A(n3171), .B(n3169), .Z(n3274) );
  AND U3296 ( .A(n3275), .B(n3276), .Z(n3169) );
  NANDN U3297 ( .A(n3277), .B(n3278), .Z(n3276) );
  OR U3298 ( .A(n3279), .B(n3280), .Z(n3278) );
  NAND U3299 ( .A(n3280), .B(n3279), .Z(n3275) );
  ANDN U3300 ( .B(B[56]), .A(n32), .Z(n3171) );
  XNOR U3301 ( .A(n3179), .B(n3281), .Z(n3172) );
  XNOR U3302 ( .A(n3178), .B(n3176), .Z(n3281) );
  AND U3303 ( .A(n3282), .B(n3283), .Z(n3176) );
  NANDN U3304 ( .A(n3284), .B(n3285), .Z(n3283) );
  NANDN U3305 ( .A(n3286), .B(n3287), .Z(n3285) );
  NANDN U3306 ( .A(n3287), .B(n3286), .Z(n3282) );
  ANDN U3307 ( .B(B[57]), .A(n33), .Z(n3178) );
  XNOR U3308 ( .A(n3186), .B(n3288), .Z(n3179) );
  XNOR U3309 ( .A(n3185), .B(n3183), .Z(n3288) );
  AND U3310 ( .A(n3289), .B(n3290), .Z(n3183) );
  NANDN U3311 ( .A(n3291), .B(n3292), .Z(n3290) );
  OR U3312 ( .A(n3293), .B(n3294), .Z(n3292) );
  NAND U3313 ( .A(n3294), .B(n3293), .Z(n3289) );
  ANDN U3314 ( .B(B[58]), .A(n34), .Z(n3185) );
  XNOR U3315 ( .A(n3193), .B(n3295), .Z(n3186) );
  XNOR U3316 ( .A(n3192), .B(n3190), .Z(n3295) );
  AND U3317 ( .A(n3296), .B(n3297), .Z(n3190) );
  NANDN U3318 ( .A(n3298), .B(n3299), .Z(n3297) );
  NANDN U3319 ( .A(n3300), .B(n3301), .Z(n3299) );
  NANDN U3320 ( .A(n3301), .B(n3300), .Z(n3296) );
  ANDN U3321 ( .B(B[59]), .A(n35), .Z(n3192) );
  XNOR U3322 ( .A(n3200), .B(n3302), .Z(n3193) );
  XNOR U3323 ( .A(n3199), .B(n3197), .Z(n3302) );
  AND U3324 ( .A(n3303), .B(n3304), .Z(n3197) );
  NANDN U3325 ( .A(n3305), .B(n3306), .Z(n3304) );
  OR U3326 ( .A(n3307), .B(n3308), .Z(n3306) );
  NAND U3327 ( .A(n3308), .B(n3307), .Z(n3303) );
  ANDN U3328 ( .B(B[60]), .A(n36), .Z(n3199) );
  XNOR U3329 ( .A(n3207), .B(n3309), .Z(n3200) );
  XNOR U3330 ( .A(n3206), .B(n3204), .Z(n3309) );
  AND U3331 ( .A(n3310), .B(n3311), .Z(n3204) );
  NANDN U3332 ( .A(n3312), .B(n3313), .Z(n3311) );
  NANDN U3333 ( .A(n3314), .B(n3315), .Z(n3313) );
  NANDN U3334 ( .A(n3315), .B(n3314), .Z(n3310) );
  ANDN U3335 ( .B(B[61]), .A(n37), .Z(n3206) );
  XNOR U3336 ( .A(n3214), .B(n3316), .Z(n3207) );
  XNOR U3337 ( .A(n3213), .B(n3211), .Z(n3316) );
  AND U3338 ( .A(n3317), .B(n3318), .Z(n3211) );
  NANDN U3339 ( .A(n3319), .B(n3320), .Z(n3318) );
  OR U3340 ( .A(n3321), .B(n3322), .Z(n3320) );
  NAND U3341 ( .A(n3322), .B(n3321), .Z(n3317) );
  ANDN U3342 ( .B(B[62]), .A(n38), .Z(n3213) );
  XNOR U3343 ( .A(n3221), .B(n3323), .Z(n3214) );
  XNOR U3344 ( .A(n3220), .B(n3218), .Z(n3323) );
  AND U3345 ( .A(n3324), .B(n3325), .Z(n3218) );
  NANDN U3346 ( .A(n3326), .B(n3327), .Z(n3325) );
  NANDN U3347 ( .A(n3328), .B(n3329), .Z(n3327) );
  NANDN U3348 ( .A(n3329), .B(n3328), .Z(n3324) );
  ANDN U3349 ( .B(B[63]), .A(n39), .Z(n3220) );
  XNOR U3350 ( .A(n3228), .B(n3330), .Z(n3221) );
  XNOR U3351 ( .A(n3227), .B(n3225), .Z(n3330) );
  AND U3352 ( .A(n3331), .B(n3332), .Z(n3225) );
  NANDN U3353 ( .A(n3333), .B(n3334), .Z(n3332) );
  OR U3354 ( .A(n3335), .B(n3336), .Z(n3334) );
  NAND U3355 ( .A(n3336), .B(n3335), .Z(n3331) );
  ANDN U3356 ( .B(B[64]), .A(n40), .Z(n3227) );
  XNOR U3357 ( .A(n3235), .B(n3337), .Z(n3228) );
  XNOR U3358 ( .A(n3234), .B(n3232), .Z(n3337) );
  AND U3359 ( .A(n3338), .B(n3339), .Z(n3232) );
  NANDN U3360 ( .A(n3340), .B(n3341), .Z(n3339) );
  NAND U3361 ( .A(n3342), .B(n3343), .Z(n3341) );
  ANDN U3362 ( .B(B[65]), .A(n41), .Z(n3234) );
  XOR U3363 ( .A(n3241), .B(n3344), .Z(n3235) );
  XNOR U3364 ( .A(n3239), .B(n3242), .Z(n3344) );
  NAND U3365 ( .A(A[2]), .B(B[66]), .Z(n3242) );
  NANDN U3366 ( .A(n3345), .B(n3346), .Z(n3239) );
  AND U3367 ( .A(A[0]), .B(B[67]), .Z(n3346) );
  XNOR U3368 ( .A(n3244), .B(n3347), .Z(n3241) );
  NAND U3369 ( .A(A[0]), .B(B[68]), .Z(n3347) );
  NAND U3370 ( .A(B[67]), .B(A[1]), .Z(n3244) );
  NAND U3371 ( .A(n3348), .B(n3349), .Z(n110) );
  NANDN U3372 ( .A(n3350), .B(n3351), .Z(n3349) );
  OR U3373 ( .A(n3352), .B(n3353), .Z(n3351) );
  NAND U3374 ( .A(n3353), .B(n3352), .Z(n3348) );
  XOR U3375 ( .A(n112), .B(n111), .Z(\A1[65] ) );
  XOR U3376 ( .A(n3353), .B(n3354), .Z(n111) );
  XNOR U3377 ( .A(n3352), .B(n3350), .Z(n3354) );
  AND U3378 ( .A(n3355), .B(n3356), .Z(n3350) );
  NANDN U3379 ( .A(n3357), .B(n3358), .Z(n3356) );
  NANDN U3380 ( .A(n3359), .B(n3360), .Z(n3358) );
  NANDN U3381 ( .A(n3360), .B(n3359), .Z(n3355) );
  ANDN U3382 ( .B(B[52]), .A(n29), .Z(n3352) );
  XNOR U3383 ( .A(n3259), .B(n3361), .Z(n3353) );
  XNOR U3384 ( .A(n3258), .B(n3256), .Z(n3361) );
  AND U3385 ( .A(n3362), .B(n3363), .Z(n3256) );
  NANDN U3386 ( .A(n3364), .B(n3365), .Z(n3363) );
  OR U3387 ( .A(n3366), .B(n3367), .Z(n3365) );
  NAND U3388 ( .A(n3367), .B(n3366), .Z(n3362) );
  ANDN U3389 ( .B(B[53]), .A(n30), .Z(n3258) );
  XNOR U3390 ( .A(n3266), .B(n3368), .Z(n3259) );
  XNOR U3391 ( .A(n3265), .B(n3263), .Z(n3368) );
  AND U3392 ( .A(n3369), .B(n3370), .Z(n3263) );
  NANDN U3393 ( .A(n3371), .B(n3372), .Z(n3370) );
  NANDN U3394 ( .A(n3373), .B(n3374), .Z(n3372) );
  NANDN U3395 ( .A(n3374), .B(n3373), .Z(n3369) );
  ANDN U3396 ( .B(B[54]), .A(n31), .Z(n3265) );
  XNOR U3397 ( .A(n3273), .B(n3375), .Z(n3266) );
  XNOR U3398 ( .A(n3272), .B(n3270), .Z(n3375) );
  AND U3399 ( .A(n3376), .B(n3377), .Z(n3270) );
  NANDN U3400 ( .A(n3378), .B(n3379), .Z(n3377) );
  OR U3401 ( .A(n3380), .B(n3381), .Z(n3379) );
  NAND U3402 ( .A(n3381), .B(n3380), .Z(n3376) );
  ANDN U3403 ( .B(B[55]), .A(n32), .Z(n3272) );
  XNOR U3404 ( .A(n3280), .B(n3382), .Z(n3273) );
  XNOR U3405 ( .A(n3279), .B(n3277), .Z(n3382) );
  AND U3406 ( .A(n3383), .B(n3384), .Z(n3277) );
  NANDN U3407 ( .A(n3385), .B(n3386), .Z(n3384) );
  NANDN U3408 ( .A(n3387), .B(n3388), .Z(n3386) );
  NANDN U3409 ( .A(n3388), .B(n3387), .Z(n3383) );
  ANDN U3410 ( .B(B[56]), .A(n33), .Z(n3279) );
  XNOR U3411 ( .A(n3287), .B(n3389), .Z(n3280) );
  XNOR U3412 ( .A(n3286), .B(n3284), .Z(n3389) );
  AND U3413 ( .A(n3390), .B(n3391), .Z(n3284) );
  NANDN U3414 ( .A(n3392), .B(n3393), .Z(n3391) );
  OR U3415 ( .A(n3394), .B(n3395), .Z(n3393) );
  NAND U3416 ( .A(n3395), .B(n3394), .Z(n3390) );
  ANDN U3417 ( .B(B[57]), .A(n34), .Z(n3286) );
  XNOR U3418 ( .A(n3294), .B(n3396), .Z(n3287) );
  XNOR U3419 ( .A(n3293), .B(n3291), .Z(n3396) );
  AND U3420 ( .A(n3397), .B(n3398), .Z(n3291) );
  NANDN U3421 ( .A(n3399), .B(n3400), .Z(n3398) );
  NANDN U3422 ( .A(n3401), .B(n3402), .Z(n3400) );
  NANDN U3423 ( .A(n3402), .B(n3401), .Z(n3397) );
  ANDN U3424 ( .B(B[58]), .A(n35), .Z(n3293) );
  XNOR U3425 ( .A(n3301), .B(n3403), .Z(n3294) );
  XNOR U3426 ( .A(n3300), .B(n3298), .Z(n3403) );
  AND U3427 ( .A(n3404), .B(n3405), .Z(n3298) );
  NANDN U3428 ( .A(n3406), .B(n3407), .Z(n3405) );
  OR U3429 ( .A(n3408), .B(n3409), .Z(n3407) );
  NAND U3430 ( .A(n3409), .B(n3408), .Z(n3404) );
  ANDN U3431 ( .B(B[59]), .A(n36), .Z(n3300) );
  XNOR U3432 ( .A(n3308), .B(n3410), .Z(n3301) );
  XNOR U3433 ( .A(n3307), .B(n3305), .Z(n3410) );
  AND U3434 ( .A(n3411), .B(n3412), .Z(n3305) );
  NANDN U3435 ( .A(n3413), .B(n3414), .Z(n3412) );
  NANDN U3436 ( .A(n3415), .B(n3416), .Z(n3414) );
  NANDN U3437 ( .A(n3416), .B(n3415), .Z(n3411) );
  ANDN U3438 ( .B(B[60]), .A(n37), .Z(n3307) );
  XNOR U3439 ( .A(n3315), .B(n3417), .Z(n3308) );
  XNOR U3440 ( .A(n3314), .B(n3312), .Z(n3417) );
  AND U3441 ( .A(n3418), .B(n3419), .Z(n3312) );
  NANDN U3442 ( .A(n3420), .B(n3421), .Z(n3419) );
  OR U3443 ( .A(n3422), .B(n3423), .Z(n3421) );
  NAND U3444 ( .A(n3423), .B(n3422), .Z(n3418) );
  ANDN U3445 ( .B(B[61]), .A(n38), .Z(n3314) );
  XNOR U3446 ( .A(n3322), .B(n3424), .Z(n3315) );
  XNOR U3447 ( .A(n3321), .B(n3319), .Z(n3424) );
  AND U3448 ( .A(n3425), .B(n3426), .Z(n3319) );
  NANDN U3449 ( .A(n3427), .B(n3428), .Z(n3426) );
  NANDN U3450 ( .A(n3429), .B(n3430), .Z(n3428) );
  NANDN U3451 ( .A(n3430), .B(n3429), .Z(n3425) );
  ANDN U3452 ( .B(B[62]), .A(n39), .Z(n3321) );
  XNOR U3453 ( .A(n3329), .B(n3431), .Z(n3322) );
  XNOR U3454 ( .A(n3328), .B(n3326), .Z(n3431) );
  AND U3455 ( .A(n3432), .B(n3433), .Z(n3326) );
  NANDN U3456 ( .A(n3434), .B(n3435), .Z(n3433) );
  OR U3457 ( .A(n3436), .B(n3437), .Z(n3435) );
  NAND U3458 ( .A(n3437), .B(n3436), .Z(n3432) );
  ANDN U3459 ( .B(B[63]), .A(n40), .Z(n3328) );
  XNOR U3460 ( .A(n3336), .B(n3438), .Z(n3329) );
  XNOR U3461 ( .A(n3335), .B(n3333), .Z(n3438) );
  AND U3462 ( .A(n3439), .B(n3440), .Z(n3333) );
  NANDN U3463 ( .A(n3441), .B(n3442), .Z(n3440) );
  NAND U3464 ( .A(n3443), .B(n3444), .Z(n3442) );
  ANDN U3465 ( .B(B[64]), .A(n41), .Z(n3335) );
  XOR U3466 ( .A(n3342), .B(n3445), .Z(n3336) );
  XNOR U3467 ( .A(n3340), .B(n3343), .Z(n3445) );
  NAND U3468 ( .A(A[2]), .B(B[65]), .Z(n3343) );
  NANDN U3469 ( .A(n3446), .B(n3447), .Z(n3340) );
  AND U3470 ( .A(A[0]), .B(B[66]), .Z(n3447) );
  XNOR U3471 ( .A(n3345), .B(n3448), .Z(n3342) );
  NAND U3472 ( .A(A[0]), .B(B[67]), .Z(n3448) );
  NAND U3473 ( .A(B[66]), .B(A[1]), .Z(n3345) );
  NAND U3474 ( .A(n3449), .B(n3450), .Z(n112) );
  NANDN U3475 ( .A(n3451), .B(n3452), .Z(n3450) );
  OR U3476 ( .A(n3453), .B(n3454), .Z(n3452) );
  NAND U3477 ( .A(n3454), .B(n3453), .Z(n3449) );
  XOR U3478 ( .A(n114), .B(n113), .Z(\A1[64] ) );
  XOR U3479 ( .A(n3454), .B(n3455), .Z(n113) );
  XNOR U3480 ( .A(n3453), .B(n3451), .Z(n3455) );
  AND U3481 ( .A(n3456), .B(n3457), .Z(n3451) );
  NANDN U3482 ( .A(n3458), .B(n3459), .Z(n3457) );
  NANDN U3483 ( .A(n3460), .B(n3461), .Z(n3459) );
  NANDN U3484 ( .A(n3461), .B(n3460), .Z(n3456) );
  ANDN U3485 ( .B(B[51]), .A(n29), .Z(n3453) );
  XNOR U3486 ( .A(n3360), .B(n3462), .Z(n3454) );
  XNOR U3487 ( .A(n3359), .B(n3357), .Z(n3462) );
  AND U3488 ( .A(n3463), .B(n3464), .Z(n3357) );
  NANDN U3489 ( .A(n3465), .B(n3466), .Z(n3464) );
  OR U3490 ( .A(n3467), .B(n3468), .Z(n3466) );
  NAND U3491 ( .A(n3468), .B(n3467), .Z(n3463) );
  ANDN U3492 ( .B(B[52]), .A(n30), .Z(n3359) );
  XNOR U3493 ( .A(n3367), .B(n3469), .Z(n3360) );
  XNOR U3494 ( .A(n3366), .B(n3364), .Z(n3469) );
  AND U3495 ( .A(n3470), .B(n3471), .Z(n3364) );
  NANDN U3496 ( .A(n3472), .B(n3473), .Z(n3471) );
  NANDN U3497 ( .A(n3474), .B(n3475), .Z(n3473) );
  NANDN U3498 ( .A(n3475), .B(n3474), .Z(n3470) );
  ANDN U3499 ( .B(B[53]), .A(n31), .Z(n3366) );
  XNOR U3500 ( .A(n3374), .B(n3476), .Z(n3367) );
  XNOR U3501 ( .A(n3373), .B(n3371), .Z(n3476) );
  AND U3502 ( .A(n3477), .B(n3478), .Z(n3371) );
  NANDN U3503 ( .A(n3479), .B(n3480), .Z(n3478) );
  OR U3504 ( .A(n3481), .B(n3482), .Z(n3480) );
  NAND U3505 ( .A(n3482), .B(n3481), .Z(n3477) );
  ANDN U3506 ( .B(B[54]), .A(n32), .Z(n3373) );
  XNOR U3507 ( .A(n3381), .B(n3483), .Z(n3374) );
  XNOR U3508 ( .A(n3380), .B(n3378), .Z(n3483) );
  AND U3509 ( .A(n3484), .B(n3485), .Z(n3378) );
  NANDN U3510 ( .A(n3486), .B(n3487), .Z(n3485) );
  NANDN U3511 ( .A(n3488), .B(n3489), .Z(n3487) );
  NANDN U3512 ( .A(n3489), .B(n3488), .Z(n3484) );
  ANDN U3513 ( .B(B[55]), .A(n33), .Z(n3380) );
  XNOR U3514 ( .A(n3388), .B(n3490), .Z(n3381) );
  XNOR U3515 ( .A(n3387), .B(n3385), .Z(n3490) );
  AND U3516 ( .A(n3491), .B(n3492), .Z(n3385) );
  NANDN U3517 ( .A(n3493), .B(n3494), .Z(n3492) );
  OR U3518 ( .A(n3495), .B(n3496), .Z(n3494) );
  NAND U3519 ( .A(n3496), .B(n3495), .Z(n3491) );
  ANDN U3520 ( .B(B[56]), .A(n34), .Z(n3387) );
  XNOR U3521 ( .A(n3395), .B(n3497), .Z(n3388) );
  XNOR U3522 ( .A(n3394), .B(n3392), .Z(n3497) );
  AND U3523 ( .A(n3498), .B(n3499), .Z(n3392) );
  NANDN U3524 ( .A(n3500), .B(n3501), .Z(n3499) );
  NANDN U3525 ( .A(n3502), .B(n3503), .Z(n3501) );
  NANDN U3526 ( .A(n3503), .B(n3502), .Z(n3498) );
  ANDN U3527 ( .B(B[57]), .A(n35), .Z(n3394) );
  XNOR U3528 ( .A(n3402), .B(n3504), .Z(n3395) );
  XNOR U3529 ( .A(n3401), .B(n3399), .Z(n3504) );
  AND U3530 ( .A(n3505), .B(n3506), .Z(n3399) );
  NANDN U3531 ( .A(n3507), .B(n3508), .Z(n3506) );
  OR U3532 ( .A(n3509), .B(n3510), .Z(n3508) );
  NAND U3533 ( .A(n3510), .B(n3509), .Z(n3505) );
  ANDN U3534 ( .B(B[58]), .A(n36), .Z(n3401) );
  XNOR U3535 ( .A(n3409), .B(n3511), .Z(n3402) );
  XNOR U3536 ( .A(n3408), .B(n3406), .Z(n3511) );
  AND U3537 ( .A(n3512), .B(n3513), .Z(n3406) );
  NANDN U3538 ( .A(n3514), .B(n3515), .Z(n3513) );
  NANDN U3539 ( .A(n3516), .B(n3517), .Z(n3515) );
  NANDN U3540 ( .A(n3517), .B(n3516), .Z(n3512) );
  ANDN U3541 ( .B(B[59]), .A(n37), .Z(n3408) );
  XNOR U3542 ( .A(n3416), .B(n3518), .Z(n3409) );
  XNOR U3543 ( .A(n3415), .B(n3413), .Z(n3518) );
  AND U3544 ( .A(n3519), .B(n3520), .Z(n3413) );
  NANDN U3545 ( .A(n3521), .B(n3522), .Z(n3520) );
  OR U3546 ( .A(n3523), .B(n3524), .Z(n3522) );
  NAND U3547 ( .A(n3524), .B(n3523), .Z(n3519) );
  ANDN U3548 ( .B(B[60]), .A(n38), .Z(n3415) );
  XNOR U3549 ( .A(n3423), .B(n3525), .Z(n3416) );
  XNOR U3550 ( .A(n3422), .B(n3420), .Z(n3525) );
  AND U3551 ( .A(n3526), .B(n3527), .Z(n3420) );
  NANDN U3552 ( .A(n3528), .B(n3529), .Z(n3527) );
  NANDN U3553 ( .A(n3530), .B(n3531), .Z(n3529) );
  NANDN U3554 ( .A(n3531), .B(n3530), .Z(n3526) );
  ANDN U3555 ( .B(B[61]), .A(n39), .Z(n3422) );
  XNOR U3556 ( .A(n3430), .B(n3532), .Z(n3423) );
  XNOR U3557 ( .A(n3429), .B(n3427), .Z(n3532) );
  AND U3558 ( .A(n3533), .B(n3534), .Z(n3427) );
  NANDN U3559 ( .A(n3535), .B(n3536), .Z(n3534) );
  OR U3560 ( .A(n3537), .B(n3538), .Z(n3536) );
  NAND U3561 ( .A(n3538), .B(n3537), .Z(n3533) );
  ANDN U3562 ( .B(B[62]), .A(n40), .Z(n3429) );
  XNOR U3563 ( .A(n3437), .B(n3539), .Z(n3430) );
  XNOR U3564 ( .A(n3436), .B(n3434), .Z(n3539) );
  AND U3565 ( .A(n3540), .B(n3541), .Z(n3434) );
  NANDN U3566 ( .A(n3542), .B(n3543), .Z(n3541) );
  NAND U3567 ( .A(n3544), .B(n3545), .Z(n3543) );
  ANDN U3568 ( .B(B[63]), .A(n41), .Z(n3436) );
  XOR U3569 ( .A(n3443), .B(n3546), .Z(n3437) );
  XNOR U3570 ( .A(n3441), .B(n3444), .Z(n3546) );
  NAND U3571 ( .A(A[2]), .B(B[64]), .Z(n3444) );
  NANDN U3572 ( .A(n3547), .B(n3548), .Z(n3441) );
  AND U3573 ( .A(A[0]), .B(B[65]), .Z(n3548) );
  XNOR U3574 ( .A(n3446), .B(n3549), .Z(n3443) );
  NAND U3575 ( .A(A[0]), .B(B[66]), .Z(n3549) );
  NAND U3576 ( .A(B[65]), .B(A[1]), .Z(n3446) );
  NAND U3577 ( .A(n3550), .B(n3551), .Z(n114) );
  NANDN U3578 ( .A(n3552), .B(n3553), .Z(n3551) );
  OR U3579 ( .A(n3554), .B(n3555), .Z(n3553) );
  NAND U3580 ( .A(n3555), .B(n3554), .Z(n3550) );
  XOR U3581 ( .A(n116), .B(n115), .Z(\A1[63] ) );
  XOR U3582 ( .A(n3555), .B(n3556), .Z(n115) );
  XNOR U3583 ( .A(n3554), .B(n3552), .Z(n3556) );
  AND U3584 ( .A(n3557), .B(n3558), .Z(n3552) );
  NANDN U3585 ( .A(n3559), .B(n3560), .Z(n3558) );
  NANDN U3586 ( .A(n3561), .B(n3562), .Z(n3560) );
  NANDN U3587 ( .A(n3562), .B(n3561), .Z(n3557) );
  ANDN U3588 ( .B(B[50]), .A(n29), .Z(n3554) );
  XNOR U3589 ( .A(n3461), .B(n3563), .Z(n3555) );
  XNOR U3590 ( .A(n3460), .B(n3458), .Z(n3563) );
  AND U3591 ( .A(n3564), .B(n3565), .Z(n3458) );
  NANDN U3592 ( .A(n3566), .B(n3567), .Z(n3565) );
  OR U3593 ( .A(n3568), .B(n3569), .Z(n3567) );
  NAND U3594 ( .A(n3569), .B(n3568), .Z(n3564) );
  ANDN U3595 ( .B(B[51]), .A(n30), .Z(n3460) );
  XNOR U3596 ( .A(n3468), .B(n3570), .Z(n3461) );
  XNOR U3597 ( .A(n3467), .B(n3465), .Z(n3570) );
  AND U3598 ( .A(n3571), .B(n3572), .Z(n3465) );
  NANDN U3599 ( .A(n3573), .B(n3574), .Z(n3572) );
  NANDN U3600 ( .A(n3575), .B(n3576), .Z(n3574) );
  NANDN U3601 ( .A(n3576), .B(n3575), .Z(n3571) );
  ANDN U3602 ( .B(B[52]), .A(n31), .Z(n3467) );
  XNOR U3603 ( .A(n3475), .B(n3577), .Z(n3468) );
  XNOR U3604 ( .A(n3474), .B(n3472), .Z(n3577) );
  AND U3605 ( .A(n3578), .B(n3579), .Z(n3472) );
  NANDN U3606 ( .A(n3580), .B(n3581), .Z(n3579) );
  OR U3607 ( .A(n3582), .B(n3583), .Z(n3581) );
  NAND U3608 ( .A(n3583), .B(n3582), .Z(n3578) );
  ANDN U3609 ( .B(B[53]), .A(n32), .Z(n3474) );
  XNOR U3610 ( .A(n3482), .B(n3584), .Z(n3475) );
  XNOR U3611 ( .A(n3481), .B(n3479), .Z(n3584) );
  AND U3612 ( .A(n3585), .B(n3586), .Z(n3479) );
  NANDN U3613 ( .A(n3587), .B(n3588), .Z(n3586) );
  NANDN U3614 ( .A(n3589), .B(n3590), .Z(n3588) );
  NANDN U3615 ( .A(n3590), .B(n3589), .Z(n3585) );
  ANDN U3616 ( .B(B[54]), .A(n33), .Z(n3481) );
  XNOR U3617 ( .A(n3489), .B(n3591), .Z(n3482) );
  XNOR U3618 ( .A(n3488), .B(n3486), .Z(n3591) );
  AND U3619 ( .A(n3592), .B(n3593), .Z(n3486) );
  NANDN U3620 ( .A(n3594), .B(n3595), .Z(n3593) );
  OR U3621 ( .A(n3596), .B(n3597), .Z(n3595) );
  NAND U3622 ( .A(n3597), .B(n3596), .Z(n3592) );
  ANDN U3623 ( .B(B[55]), .A(n34), .Z(n3488) );
  XNOR U3624 ( .A(n3496), .B(n3598), .Z(n3489) );
  XNOR U3625 ( .A(n3495), .B(n3493), .Z(n3598) );
  AND U3626 ( .A(n3599), .B(n3600), .Z(n3493) );
  NANDN U3627 ( .A(n3601), .B(n3602), .Z(n3600) );
  NANDN U3628 ( .A(n3603), .B(n3604), .Z(n3602) );
  NANDN U3629 ( .A(n3604), .B(n3603), .Z(n3599) );
  ANDN U3630 ( .B(B[56]), .A(n35), .Z(n3495) );
  XNOR U3631 ( .A(n3503), .B(n3605), .Z(n3496) );
  XNOR U3632 ( .A(n3502), .B(n3500), .Z(n3605) );
  AND U3633 ( .A(n3606), .B(n3607), .Z(n3500) );
  NANDN U3634 ( .A(n3608), .B(n3609), .Z(n3607) );
  OR U3635 ( .A(n3610), .B(n3611), .Z(n3609) );
  NAND U3636 ( .A(n3611), .B(n3610), .Z(n3606) );
  ANDN U3637 ( .B(B[57]), .A(n36), .Z(n3502) );
  XNOR U3638 ( .A(n3510), .B(n3612), .Z(n3503) );
  XNOR U3639 ( .A(n3509), .B(n3507), .Z(n3612) );
  AND U3640 ( .A(n3613), .B(n3614), .Z(n3507) );
  NANDN U3641 ( .A(n3615), .B(n3616), .Z(n3614) );
  NANDN U3642 ( .A(n3617), .B(n3618), .Z(n3616) );
  NANDN U3643 ( .A(n3618), .B(n3617), .Z(n3613) );
  ANDN U3644 ( .B(B[58]), .A(n37), .Z(n3509) );
  XNOR U3645 ( .A(n3517), .B(n3619), .Z(n3510) );
  XNOR U3646 ( .A(n3516), .B(n3514), .Z(n3619) );
  AND U3647 ( .A(n3620), .B(n3621), .Z(n3514) );
  NANDN U3648 ( .A(n3622), .B(n3623), .Z(n3621) );
  OR U3649 ( .A(n3624), .B(n3625), .Z(n3623) );
  NAND U3650 ( .A(n3625), .B(n3624), .Z(n3620) );
  ANDN U3651 ( .B(B[59]), .A(n38), .Z(n3516) );
  XNOR U3652 ( .A(n3524), .B(n3626), .Z(n3517) );
  XNOR U3653 ( .A(n3523), .B(n3521), .Z(n3626) );
  AND U3654 ( .A(n3627), .B(n3628), .Z(n3521) );
  NANDN U3655 ( .A(n3629), .B(n3630), .Z(n3628) );
  NANDN U3656 ( .A(n3631), .B(n3632), .Z(n3630) );
  NANDN U3657 ( .A(n3632), .B(n3631), .Z(n3627) );
  ANDN U3658 ( .B(B[60]), .A(n39), .Z(n3523) );
  XNOR U3659 ( .A(n3531), .B(n3633), .Z(n3524) );
  XNOR U3660 ( .A(n3530), .B(n3528), .Z(n3633) );
  AND U3661 ( .A(n3634), .B(n3635), .Z(n3528) );
  NANDN U3662 ( .A(n3636), .B(n3637), .Z(n3635) );
  OR U3663 ( .A(n3638), .B(n3639), .Z(n3637) );
  NAND U3664 ( .A(n3639), .B(n3638), .Z(n3634) );
  ANDN U3665 ( .B(B[61]), .A(n40), .Z(n3530) );
  XNOR U3666 ( .A(n3538), .B(n3640), .Z(n3531) );
  XNOR U3667 ( .A(n3537), .B(n3535), .Z(n3640) );
  AND U3668 ( .A(n3641), .B(n3642), .Z(n3535) );
  NANDN U3669 ( .A(n3643), .B(n3644), .Z(n3642) );
  NAND U3670 ( .A(n3645), .B(n3646), .Z(n3644) );
  ANDN U3671 ( .B(B[62]), .A(n41), .Z(n3537) );
  XOR U3672 ( .A(n3544), .B(n3647), .Z(n3538) );
  XNOR U3673 ( .A(n3542), .B(n3545), .Z(n3647) );
  NAND U3674 ( .A(A[2]), .B(B[63]), .Z(n3545) );
  NANDN U3675 ( .A(n3648), .B(n3649), .Z(n3542) );
  AND U3676 ( .A(A[0]), .B(B[64]), .Z(n3649) );
  XNOR U3677 ( .A(n3547), .B(n3650), .Z(n3544) );
  NAND U3678 ( .A(A[0]), .B(B[65]), .Z(n3650) );
  NAND U3679 ( .A(B[64]), .B(A[1]), .Z(n3547) );
  NAND U3680 ( .A(n3651), .B(n3652), .Z(n116) );
  NANDN U3681 ( .A(n3653), .B(n3654), .Z(n3652) );
  OR U3682 ( .A(n3655), .B(n3656), .Z(n3654) );
  NAND U3683 ( .A(n3656), .B(n3655), .Z(n3651) );
  XOR U3684 ( .A(n118), .B(n117), .Z(\A1[62] ) );
  XOR U3685 ( .A(n3656), .B(n3657), .Z(n117) );
  XNOR U3686 ( .A(n3655), .B(n3653), .Z(n3657) );
  AND U3687 ( .A(n3658), .B(n3659), .Z(n3653) );
  NANDN U3688 ( .A(n3660), .B(n3661), .Z(n3659) );
  NANDN U3689 ( .A(n3662), .B(n3663), .Z(n3661) );
  NANDN U3690 ( .A(n3663), .B(n3662), .Z(n3658) );
  ANDN U3691 ( .B(B[49]), .A(n29), .Z(n3655) );
  XNOR U3692 ( .A(n3562), .B(n3664), .Z(n3656) );
  XNOR U3693 ( .A(n3561), .B(n3559), .Z(n3664) );
  AND U3694 ( .A(n3665), .B(n3666), .Z(n3559) );
  NANDN U3695 ( .A(n3667), .B(n3668), .Z(n3666) );
  OR U3696 ( .A(n3669), .B(n3670), .Z(n3668) );
  NAND U3697 ( .A(n3670), .B(n3669), .Z(n3665) );
  ANDN U3698 ( .B(B[50]), .A(n30), .Z(n3561) );
  XNOR U3699 ( .A(n3569), .B(n3671), .Z(n3562) );
  XNOR U3700 ( .A(n3568), .B(n3566), .Z(n3671) );
  AND U3701 ( .A(n3672), .B(n3673), .Z(n3566) );
  NANDN U3702 ( .A(n3674), .B(n3675), .Z(n3673) );
  NANDN U3703 ( .A(n3676), .B(n3677), .Z(n3675) );
  NANDN U3704 ( .A(n3677), .B(n3676), .Z(n3672) );
  ANDN U3705 ( .B(B[51]), .A(n31), .Z(n3568) );
  XNOR U3706 ( .A(n3576), .B(n3678), .Z(n3569) );
  XNOR U3707 ( .A(n3575), .B(n3573), .Z(n3678) );
  AND U3708 ( .A(n3679), .B(n3680), .Z(n3573) );
  NANDN U3709 ( .A(n3681), .B(n3682), .Z(n3680) );
  OR U3710 ( .A(n3683), .B(n3684), .Z(n3682) );
  NAND U3711 ( .A(n3684), .B(n3683), .Z(n3679) );
  ANDN U3712 ( .B(B[52]), .A(n32), .Z(n3575) );
  XNOR U3713 ( .A(n3583), .B(n3685), .Z(n3576) );
  XNOR U3714 ( .A(n3582), .B(n3580), .Z(n3685) );
  AND U3715 ( .A(n3686), .B(n3687), .Z(n3580) );
  NANDN U3716 ( .A(n3688), .B(n3689), .Z(n3687) );
  NANDN U3717 ( .A(n3690), .B(n3691), .Z(n3689) );
  NANDN U3718 ( .A(n3691), .B(n3690), .Z(n3686) );
  ANDN U3719 ( .B(B[53]), .A(n33), .Z(n3582) );
  XNOR U3720 ( .A(n3590), .B(n3692), .Z(n3583) );
  XNOR U3721 ( .A(n3589), .B(n3587), .Z(n3692) );
  AND U3722 ( .A(n3693), .B(n3694), .Z(n3587) );
  NANDN U3723 ( .A(n3695), .B(n3696), .Z(n3694) );
  OR U3724 ( .A(n3697), .B(n3698), .Z(n3696) );
  NAND U3725 ( .A(n3698), .B(n3697), .Z(n3693) );
  ANDN U3726 ( .B(B[54]), .A(n34), .Z(n3589) );
  XNOR U3727 ( .A(n3597), .B(n3699), .Z(n3590) );
  XNOR U3728 ( .A(n3596), .B(n3594), .Z(n3699) );
  AND U3729 ( .A(n3700), .B(n3701), .Z(n3594) );
  NANDN U3730 ( .A(n3702), .B(n3703), .Z(n3701) );
  NANDN U3731 ( .A(n3704), .B(n3705), .Z(n3703) );
  NANDN U3732 ( .A(n3705), .B(n3704), .Z(n3700) );
  ANDN U3733 ( .B(B[55]), .A(n35), .Z(n3596) );
  XNOR U3734 ( .A(n3604), .B(n3706), .Z(n3597) );
  XNOR U3735 ( .A(n3603), .B(n3601), .Z(n3706) );
  AND U3736 ( .A(n3707), .B(n3708), .Z(n3601) );
  NANDN U3737 ( .A(n3709), .B(n3710), .Z(n3708) );
  OR U3738 ( .A(n3711), .B(n3712), .Z(n3710) );
  NAND U3739 ( .A(n3712), .B(n3711), .Z(n3707) );
  ANDN U3740 ( .B(B[56]), .A(n36), .Z(n3603) );
  XNOR U3741 ( .A(n3611), .B(n3713), .Z(n3604) );
  XNOR U3742 ( .A(n3610), .B(n3608), .Z(n3713) );
  AND U3743 ( .A(n3714), .B(n3715), .Z(n3608) );
  NANDN U3744 ( .A(n3716), .B(n3717), .Z(n3715) );
  NANDN U3745 ( .A(n3718), .B(n3719), .Z(n3717) );
  NANDN U3746 ( .A(n3719), .B(n3718), .Z(n3714) );
  ANDN U3747 ( .B(B[57]), .A(n37), .Z(n3610) );
  XNOR U3748 ( .A(n3618), .B(n3720), .Z(n3611) );
  XNOR U3749 ( .A(n3617), .B(n3615), .Z(n3720) );
  AND U3750 ( .A(n3721), .B(n3722), .Z(n3615) );
  NANDN U3751 ( .A(n3723), .B(n3724), .Z(n3722) );
  OR U3752 ( .A(n3725), .B(n3726), .Z(n3724) );
  NAND U3753 ( .A(n3726), .B(n3725), .Z(n3721) );
  ANDN U3754 ( .B(B[58]), .A(n38), .Z(n3617) );
  XNOR U3755 ( .A(n3625), .B(n3727), .Z(n3618) );
  XNOR U3756 ( .A(n3624), .B(n3622), .Z(n3727) );
  AND U3757 ( .A(n3728), .B(n3729), .Z(n3622) );
  NANDN U3758 ( .A(n3730), .B(n3731), .Z(n3729) );
  NANDN U3759 ( .A(n3732), .B(n3733), .Z(n3731) );
  NANDN U3760 ( .A(n3733), .B(n3732), .Z(n3728) );
  ANDN U3761 ( .B(B[59]), .A(n39), .Z(n3624) );
  XNOR U3762 ( .A(n3632), .B(n3734), .Z(n3625) );
  XNOR U3763 ( .A(n3631), .B(n3629), .Z(n3734) );
  AND U3764 ( .A(n3735), .B(n3736), .Z(n3629) );
  NANDN U3765 ( .A(n3737), .B(n3738), .Z(n3736) );
  OR U3766 ( .A(n3739), .B(n3740), .Z(n3738) );
  NAND U3767 ( .A(n3740), .B(n3739), .Z(n3735) );
  ANDN U3768 ( .B(B[60]), .A(n40), .Z(n3631) );
  XNOR U3769 ( .A(n3639), .B(n3741), .Z(n3632) );
  XNOR U3770 ( .A(n3638), .B(n3636), .Z(n3741) );
  AND U3771 ( .A(n3742), .B(n3743), .Z(n3636) );
  NANDN U3772 ( .A(n3744), .B(n3745), .Z(n3743) );
  NAND U3773 ( .A(n3746), .B(n3747), .Z(n3745) );
  ANDN U3774 ( .B(B[61]), .A(n41), .Z(n3638) );
  XOR U3775 ( .A(n3645), .B(n3748), .Z(n3639) );
  XNOR U3776 ( .A(n3643), .B(n3646), .Z(n3748) );
  NAND U3777 ( .A(A[2]), .B(B[62]), .Z(n3646) );
  NANDN U3778 ( .A(n3749), .B(n3750), .Z(n3643) );
  AND U3779 ( .A(A[0]), .B(B[63]), .Z(n3750) );
  XNOR U3780 ( .A(n3648), .B(n3751), .Z(n3645) );
  NAND U3781 ( .A(A[0]), .B(B[64]), .Z(n3751) );
  NAND U3782 ( .A(B[63]), .B(A[1]), .Z(n3648) );
  NAND U3783 ( .A(n3752), .B(n3753), .Z(n118) );
  NANDN U3784 ( .A(n3754), .B(n3755), .Z(n3753) );
  OR U3785 ( .A(n3756), .B(n3757), .Z(n3755) );
  NAND U3786 ( .A(n3757), .B(n3756), .Z(n3752) );
  XOR U3787 ( .A(n120), .B(n119), .Z(\A1[61] ) );
  XOR U3788 ( .A(n3757), .B(n3758), .Z(n119) );
  XNOR U3789 ( .A(n3756), .B(n3754), .Z(n3758) );
  AND U3790 ( .A(n3759), .B(n3760), .Z(n3754) );
  NANDN U3791 ( .A(n3761), .B(n3762), .Z(n3760) );
  NANDN U3792 ( .A(n3763), .B(n3764), .Z(n3762) );
  NANDN U3793 ( .A(n3764), .B(n3763), .Z(n3759) );
  ANDN U3794 ( .B(B[48]), .A(n29), .Z(n3756) );
  XNOR U3795 ( .A(n3663), .B(n3765), .Z(n3757) );
  XNOR U3796 ( .A(n3662), .B(n3660), .Z(n3765) );
  AND U3797 ( .A(n3766), .B(n3767), .Z(n3660) );
  NANDN U3798 ( .A(n3768), .B(n3769), .Z(n3767) );
  OR U3799 ( .A(n3770), .B(n3771), .Z(n3769) );
  NAND U3800 ( .A(n3771), .B(n3770), .Z(n3766) );
  ANDN U3801 ( .B(B[49]), .A(n30), .Z(n3662) );
  XNOR U3802 ( .A(n3670), .B(n3772), .Z(n3663) );
  XNOR U3803 ( .A(n3669), .B(n3667), .Z(n3772) );
  AND U3804 ( .A(n3773), .B(n3774), .Z(n3667) );
  NANDN U3805 ( .A(n3775), .B(n3776), .Z(n3774) );
  NANDN U3806 ( .A(n3777), .B(n3778), .Z(n3776) );
  NANDN U3807 ( .A(n3778), .B(n3777), .Z(n3773) );
  ANDN U3808 ( .B(B[50]), .A(n31), .Z(n3669) );
  XNOR U3809 ( .A(n3677), .B(n3779), .Z(n3670) );
  XNOR U3810 ( .A(n3676), .B(n3674), .Z(n3779) );
  AND U3811 ( .A(n3780), .B(n3781), .Z(n3674) );
  NANDN U3812 ( .A(n3782), .B(n3783), .Z(n3781) );
  OR U3813 ( .A(n3784), .B(n3785), .Z(n3783) );
  NAND U3814 ( .A(n3785), .B(n3784), .Z(n3780) );
  ANDN U3815 ( .B(B[51]), .A(n32), .Z(n3676) );
  XNOR U3816 ( .A(n3684), .B(n3786), .Z(n3677) );
  XNOR U3817 ( .A(n3683), .B(n3681), .Z(n3786) );
  AND U3818 ( .A(n3787), .B(n3788), .Z(n3681) );
  NANDN U3819 ( .A(n3789), .B(n3790), .Z(n3788) );
  NANDN U3820 ( .A(n3791), .B(n3792), .Z(n3790) );
  NANDN U3821 ( .A(n3792), .B(n3791), .Z(n3787) );
  ANDN U3822 ( .B(B[52]), .A(n33), .Z(n3683) );
  XNOR U3823 ( .A(n3691), .B(n3793), .Z(n3684) );
  XNOR U3824 ( .A(n3690), .B(n3688), .Z(n3793) );
  AND U3825 ( .A(n3794), .B(n3795), .Z(n3688) );
  NANDN U3826 ( .A(n3796), .B(n3797), .Z(n3795) );
  OR U3827 ( .A(n3798), .B(n3799), .Z(n3797) );
  NAND U3828 ( .A(n3799), .B(n3798), .Z(n3794) );
  ANDN U3829 ( .B(B[53]), .A(n34), .Z(n3690) );
  XNOR U3830 ( .A(n3698), .B(n3800), .Z(n3691) );
  XNOR U3831 ( .A(n3697), .B(n3695), .Z(n3800) );
  AND U3832 ( .A(n3801), .B(n3802), .Z(n3695) );
  NANDN U3833 ( .A(n3803), .B(n3804), .Z(n3802) );
  NANDN U3834 ( .A(n3805), .B(n3806), .Z(n3804) );
  NANDN U3835 ( .A(n3806), .B(n3805), .Z(n3801) );
  ANDN U3836 ( .B(B[54]), .A(n35), .Z(n3697) );
  XNOR U3837 ( .A(n3705), .B(n3807), .Z(n3698) );
  XNOR U3838 ( .A(n3704), .B(n3702), .Z(n3807) );
  AND U3839 ( .A(n3808), .B(n3809), .Z(n3702) );
  NANDN U3840 ( .A(n3810), .B(n3811), .Z(n3809) );
  OR U3841 ( .A(n3812), .B(n3813), .Z(n3811) );
  NAND U3842 ( .A(n3813), .B(n3812), .Z(n3808) );
  ANDN U3843 ( .B(B[55]), .A(n36), .Z(n3704) );
  XNOR U3844 ( .A(n3712), .B(n3814), .Z(n3705) );
  XNOR U3845 ( .A(n3711), .B(n3709), .Z(n3814) );
  AND U3846 ( .A(n3815), .B(n3816), .Z(n3709) );
  NANDN U3847 ( .A(n3817), .B(n3818), .Z(n3816) );
  NANDN U3848 ( .A(n3819), .B(n3820), .Z(n3818) );
  NANDN U3849 ( .A(n3820), .B(n3819), .Z(n3815) );
  ANDN U3850 ( .B(B[56]), .A(n37), .Z(n3711) );
  XNOR U3851 ( .A(n3719), .B(n3821), .Z(n3712) );
  XNOR U3852 ( .A(n3718), .B(n3716), .Z(n3821) );
  AND U3853 ( .A(n3822), .B(n3823), .Z(n3716) );
  NANDN U3854 ( .A(n3824), .B(n3825), .Z(n3823) );
  OR U3855 ( .A(n3826), .B(n3827), .Z(n3825) );
  NAND U3856 ( .A(n3827), .B(n3826), .Z(n3822) );
  ANDN U3857 ( .B(B[57]), .A(n38), .Z(n3718) );
  XNOR U3858 ( .A(n3726), .B(n3828), .Z(n3719) );
  XNOR U3859 ( .A(n3725), .B(n3723), .Z(n3828) );
  AND U3860 ( .A(n3829), .B(n3830), .Z(n3723) );
  NANDN U3861 ( .A(n3831), .B(n3832), .Z(n3830) );
  NANDN U3862 ( .A(n3833), .B(n3834), .Z(n3832) );
  NANDN U3863 ( .A(n3834), .B(n3833), .Z(n3829) );
  ANDN U3864 ( .B(B[58]), .A(n39), .Z(n3725) );
  XNOR U3865 ( .A(n3733), .B(n3835), .Z(n3726) );
  XNOR U3866 ( .A(n3732), .B(n3730), .Z(n3835) );
  AND U3867 ( .A(n3836), .B(n3837), .Z(n3730) );
  NANDN U3868 ( .A(n3838), .B(n3839), .Z(n3837) );
  OR U3869 ( .A(n3840), .B(n3841), .Z(n3839) );
  NAND U3870 ( .A(n3841), .B(n3840), .Z(n3836) );
  ANDN U3871 ( .B(B[59]), .A(n40), .Z(n3732) );
  XNOR U3872 ( .A(n3740), .B(n3842), .Z(n3733) );
  XNOR U3873 ( .A(n3739), .B(n3737), .Z(n3842) );
  AND U3874 ( .A(n3843), .B(n3844), .Z(n3737) );
  NANDN U3875 ( .A(n3845), .B(n3846), .Z(n3844) );
  NAND U3876 ( .A(n3847), .B(n3848), .Z(n3846) );
  ANDN U3877 ( .B(B[60]), .A(n41), .Z(n3739) );
  XOR U3878 ( .A(n3746), .B(n3849), .Z(n3740) );
  XNOR U3879 ( .A(n3744), .B(n3747), .Z(n3849) );
  NAND U3880 ( .A(A[2]), .B(B[61]), .Z(n3747) );
  NANDN U3881 ( .A(n3850), .B(n3851), .Z(n3744) );
  AND U3882 ( .A(A[0]), .B(B[62]), .Z(n3851) );
  XNOR U3883 ( .A(n3749), .B(n3852), .Z(n3746) );
  NAND U3884 ( .A(A[0]), .B(B[63]), .Z(n3852) );
  NAND U3885 ( .A(B[62]), .B(A[1]), .Z(n3749) );
  NAND U3886 ( .A(n3853), .B(n3854), .Z(n120) );
  NANDN U3887 ( .A(n3855), .B(n3856), .Z(n3854) );
  OR U3888 ( .A(n3857), .B(n3858), .Z(n3856) );
  NAND U3889 ( .A(n3858), .B(n3857), .Z(n3853) );
  XOR U3890 ( .A(n122), .B(n121), .Z(\A1[60] ) );
  XOR U3891 ( .A(n3858), .B(n3859), .Z(n121) );
  XNOR U3892 ( .A(n3857), .B(n3855), .Z(n3859) );
  AND U3893 ( .A(n3860), .B(n3861), .Z(n3855) );
  NANDN U3894 ( .A(n3862), .B(n3863), .Z(n3861) );
  NANDN U3895 ( .A(n3864), .B(n3865), .Z(n3863) );
  NANDN U3896 ( .A(n3865), .B(n3864), .Z(n3860) );
  ANDN U3897 ( .B(B[47]), .A(n29), .Z(n3857) );
  XNOR U3898 ( .A(n3764), .B(n3866), .Z(n3858) );
  XNOR U3899 ( .A(n3763), .B(n3761), .Z(n3866) );
  AND U3900 ( .A(n3867), .B(n3868), .Z(n3761) );
  NANDN U3901 ( .A(n3869), .B(n3870), .Z(n3868) );
  OR U3902 ( .A(n3871), .B(n3872), .Z(n3870) );
  NAND U3903 ( .A(n3872), .B(n3871), .Z(n3867) );
  ANDN U3904 ( .B(B[48]), .A(n30), .Z(n3763) );
  XNOR U3905 ( .A(n3771), .B(n3873), .Z(n3764) );
  XNOR U3906 ( .A(n3770), .B(n3768), .Z(n3873) );
  AND U3907 ( .A(n3874), .B(n3875), .Z(n3768) );
  NANDN U3908 ( .A(n3876), .B(n3877), .Z(n3875) );
  NANDN U3909 ( .A(n3878), .B(n3879), .Z(n3877) );
  NANDN U3910 ( .A(n3879), .B(n3878), .Z(n3874) );
  ANDN U3911 ( .B(B[49]), .A(n31), .Z(n3770) );
  XNOR U3912 ( .A(n3778), .B(n3880), .Z(n3771) );
  XNOR U3913 ( .A(n3777), .B(n3775), .Z(n3880) );
  AND U3914 ( .A(n3881), .B(n3882), .Z(n3775) );
  NANDN U3915 ( .A(n3883), .B(n3884), .Z(n3882) );
  OR U3916 ( .A(n3885), .B(n3886), .Z(n3884) );
  NAND U3917 ( .A(n3886), .B(n3885), .Z(n3881) );
  ANDN U3918 ( .B(B[50]), .A(n32), .Z(n3777) );
  XNOR U3919 ( .A(n3785), .B(n3887), .Z(n3778) );
  XNOR U3920 ( .A(n3784), .B(n3782), .Z(n3887) );
  AND U3921 ( .A(n3888), .B(n3889), .Z(n3782) );
  NANDN U3922 ( .A(n3890), .B(n3891), .Z(n3889) );
  NANDN U3923 ( .A(n3892), .B(n3893), .Z(n3891) );
  NANDN U3924 ( .A(n3893), .B(n3892), .Z(n3888) );
  ANDN U3925 ( .B(B[51]), .A(n33), .Z(n3784) );
  XNOR U3926 ( .A(n3792), .B(n3894), .Z(n3785) );
  XNOR U3927 ( .A(n3791), .B(n3789), .Z(n3894) );
  AND U3928 ( .A(n3895), .B(n3896), .Z(n3789) );
  NANDN U3929 ( .A(n3897), .B(n3898), .Z(n3896) );
  OR U3930 ( .A(n3899), .B(n3900), .Z(n3898) );
  NAND U3931 ( .A(n3900), .B(n3899), .Z(n3895) );
  ANDN U3932 ( .B(B[52]), .A(n34), .Z(n3791) );
  XNOR U3933 ( .A(n3799), .B(n3901), .Z(n3792) );
  XNOR U3934 ( .A(n3798), .B(n3796), .Z(n3901) );
  AND U3935 ( .A(n3902), .B(n3903), .Z(n3796) );
  NANDN U3936 ( .A(n3904), .B(n3905), .Z(n3903) );
  NANDN U3937 ( .A(n3906), .B(n3907), .Z(n3905) );
  NANDN U3938 ( .A(n3907), .B(n3906), .Z(n3902) );
  ANDN U3939 ( .B(B[53]), .A(n35), .Z(n3798) );
  XNOR U3940 ( .A(n3806), .B(n3908), .Z(n3799) );
  XNOR U3941 ( .A(n3805), .B(n3803), .Z(n3908) );
  AND U3942 ( .A(n3909), .B(n3910), .Z(n3803) );
  NANDN U3943 ( .A(n3911), .B(n3912), .Z(n3910) );
  OR U3944 ( .A(n3913), .B(n3914), .Z(n3912) );
  NAND U3945 ( .A(n3914), .B(n3913), .Z(n3909) );
  ANDN U3946 ( .B(B[54]), .A(n36), .Z(n3805) );
  XNOR U3947 ( .A(n3813), .B(n3915), .Z(n3806) );
  XNOR U3948 ( .A(n3812), .B(n3810), .Z(n3915) );
  AND U3949 ( .A(n3916), .B(n3917), .Z(n3810) );
  NANDN U3950 ( .A(n3918), .B(n3919), .Z(n3917) );
  NANDN U3951 ( .A(n3920), .B(n3921), .Z(n3919) );
  NANDN U3952 ( .A(n3921), .B(n3920), .Z(n3916) );
  ANDN U3953 ( .B(B[55]), .A(n37), .Z(n3812) );
  XNOR U3954 ( .A(n3820), .B(n3922), .Z(n3813) );
  XNOR U3955 ( .A(n3819), .B(n3817), .Z(n3922) );
  AND U3956 ( .A(n3923), .B(n3924), .Z(n3817) );
  NANDN U3957 ( .A(n3925), .B(n3926), .Z(n3924) );
  OR U3958 ( .A(n3927), .B(n3928), .Z(n3926) );
  NAND U3959 ( .A(n3928), .B(n3927), .Z(n3923) );
  ANDN U3960 ( .B(B[56]), .A(n38), .Z(n3819) );
  XNOR U3961 ( .A(n3827), .B(n3929), .Z(n3820) );
  XNOR U3962 ( .A(n3826), .B(n3824), .Z(n3929) );
  AND U3963 ( .A(n3930), .B(n3931), .Z(n3824) );
  NANDN U3964 ( .A(n3932), .B(n3933), .Z(n3931) );
  NANDN U3965 ( .A(n3934), .B(n3935), .Z(n3933) );
  NANDN U3966 ( .A(n3935), .B(n3934), .Z(n3930) );
  ANDN U3967 ( .B(B[57]), .A(n39), .Z(n3826) );
  XNOR U3968 ( .A(n3834), .B(n3936), .Z(n3827) );
  XNOR U3969 ( .A(n3833), .B(n3831), .Z(n3936) );
  AND U3970 ( .A(n3937), .B(n3938), .Z(n3831) );
  NANDN U3971 ( .A(n3939), .B(n3940), .Z(n3938) );
  OR U3972 ( .A(n3941), .B(n3942), .Z(n3940) );
  NAND U3973 ( .A(n3942), .B(n3941), .Z(n3937) );
  ANDN U3974 ( .B(B[58]), .A(n40), .Z(n3833) );
  XNOR U3975 ( .A(n3841), .B(n3943), .Z(n3834) );
  XNOR U3976 ( .A(n3840), .B(n3838), .Z(n3943) );
  AND U3977 ( .A(n3944), .B(n3945), .Z(n3838) );
  NANDN U3978 ( .A(n3946), .B(n3947), .Z(n3945) );
  NAND U3979 ( .A(n3948), .B(n3949), .Z(n3947) );
  ANDN U3980 ( .B(B[59]), .A(n41), .Z(n3840) );
  XOR U3981 ( .A(n3847), .B(n3950), .Z(n3841) );
  XNOR U3982 ( .A(n3845), .B(n3848), .Z(n3950) );
  NAND U3983 ( .A(A[2]), .B(B[60]), .Z(n3848) );
  NANDN U3984 ( .A(n3951), .B(n3952), .Z(n3845) );
  AND U3985 ( .A(A[0]), .B(B[61]), .Z(n3952) );
  XNOR U3986 ( .A(n3850), .B(n3953), .Z(n3847) );
  NAND U3987 ( .A(A[0]), .B(B[62]), .Z(n3953) );
  NAND U3988 ( .A(B[61]), .B(A[1]), .Z(n3850) );
  NAND U3989 ( .A(n3954), .B(n3955), .Z(n122) );
  NANDN U3990 ( .A(n3956), .B(n3957), .Z(n3955) );
  OR U3991 ( .A(n3958), .B(n3959), .Z(n3957) );
  NAND U3992 ( .A(n3959), .B(n3958), .Z(n3954) );
  XOR U3993 ( .A(n3960), .B(n3961), .Z(\A1[5] ) );
  XNOR U3994 ( .A(n3962), .B(n26), .Z(n3961) );
  XOR U3995 ( .A(n124), .B(n123), .Z(\A1[59] ) );
  XOR U3996 ( .A(n3959), .B(n3963), .Z(n123) );
  XNOR U3997 ( .A(n3958), .B(n3956), .Z(n3963) );
  AND U3998 ( .A(n3964), .B(n3965), .Z(n3956) );
  NANDN U3999 ( .A(n3966), .B(n3967), .Z(n3965) );
  NANDN U4000 ( .A(n3968), .B(n3969), .Z(n3967) );
  NANDN U4001 ( .A(n3969), .B(n3968), .Z(n3964) );
  ANDN U4002 ( .B(B[46]), .A(n29), .Z(n3958) );
  XNOR U4003 ( .A(n3865), .B(n3970), .Z(n3959) );
  XNOR U4004 ( .A(n3864), .B(n3862), .Z(n3970) );
  AND U4005 ( .A(n3971), .B(n3972), .Z(n3862) );
  NANDN U4006 ( .A(n3973), .B(n3974), .Z(n3972) );
  OR U4007 ( .A(n3975), .B(n3976), .Z(n3974) );
  NAND U4008 ( .A(n3976), .B(n3975), .Z(n3971) );
  ANDN U4009 ( .B(B[47]), .A(n30), .Z(n3864) );
  XNOR U4010 ( .A(n3872), .B(n3977), .Z(n3865) );
  XNOR U4011 ( .A(n3871), .B(n3869), .Z(n3977) );
  AND U4012 ( .A(n3978), .B(n3979), .Z(n3869) );
  NANDN U4013 ( .A(n3980), .B(n3981), .Z(n3979) );
  NANDN U4014 ( .A(n3982), .B(n3983), .Z(n3981) );
  NANDN U4015 ( .A(n3983), .B(n3982), .Z(n3978) );
  ANDN U4016 ( .B(B[48]), .A(n31), .Z(n3871) );
  XNOR U4017 ( .A(n3879), .B(n3984), .Z(n3872) );
  XNOR U4018 ( .A(n3878), .B(n3876), .Z(n3984) );
  AND U4019 ( .A(n3985), .B(n3986), .Z(n3876) );
  NANDN U4020 ( .A(n3987), .B(n3988), .Z(n3986) );
  OR U4021 ( .A(n3989), .B(n3990), .Z(n3988) );
  NAND U4022 ( .A(n3990), .B(n3989), .Z(n3985) );
  ANDN U4023 ( .B(B[49]), .A(n32), .Z(n3878) );
  XNOR U4024 ( .A(n3886), .B(n3991), .Z(n3879) );
  XNOR U4025 ( .A(n3885), .B(n3883), .Z(n3991) );
  AND U4026 ( .A(n3992), .B(n3993), .Z(n3883) );
  NANDN U4027 ( .A(n3994), .B(n3995), .Z(n3993) );
  NANDN U4028 ( .A(n3996), .B(n3997), .Z(n3995) );
  NANDN U4029 ( .A(n3997), .B(n3996), .Z(n3992) );
  ANDN U4030 ( .B(B[50]), .A(n33), .Z(n3885) );
  XNOR U4031 ( .A(n3893), .B(n3998), .Z(n3886) );
  XNOR U4032 ( .A(n3892), .B(n3890), .Z(n3998) );
  AND U4033 ( .A(n3999), .B(n4000), .Z(n3890) );
  NANDN U4034 ( .A(n4001), .B(n4002), .Z(n4000) );
  OR U4035 ( .A(n4003), .B(n4004), .Z(n4002) );
  NAND U4036 ( .A(n4004), .B(n4003), .Z(n3999) );
  ANDN U4037 ( .B(B[51]), .A(n34), .Z(n3892) );
  XNOR U4038 ( .A(n3900), .B(n4005), .Z(n3893) );
  XNOR U4039 ( .A(n3899), .B(n3897), .Z(n4005) );
  AND U4040 ( .A(n4006), .B(n4007), .Z(n3897) );
  NANDN U4041 ( .A(n4008), .B(n4009), .Z(n4007) );
  NANDN U4042 ( .A(n4010), .B(n4011), .Z(n4009) );
  NANDN U4043 ( .A(n4011), .B(n4010), .Z(n4006) );
  ANDN U4044 ( .B(B[52]), .A(n35), .Z(n3899) );
  XNOR U4045 ( .A(n3907), .B(n4012), .Z(n3900) );
  XNOR U4046 ( .A(n3906), .B(n3904), .Z(n4012) );
  AND U4047 ( .A(n4013), .B(n4014), .Z(n3904) );
  NANDN U4048 ( .A(n4015), .B(n4016), .Z(n4014) );
  OR U4049 ( .A(n4017), .B(n4018), .Z(n4016) );
  NAND U4050 ( .A(n4018), .B(n4017), .Z(n4013) );
  ANDN U4051 ( .B(B[53]), .A(n36), .Z(n3906) );
  XNOR U4052 ( .A(n3914), .B(n4019), .Z(n3907) );
  XNOR U4053 ( .A(n3913), .B(n3911), .Z(n4019) );
  AND U4054 ( .A(n4020), .B(n4021), .Z(n3911) );
  NANDN U4055 ( .A(n4022), .B(n4023), .Z(n4021) );
  NANDN U4056 ( .A(n4024), .B(n4025), .Z(n4023) );
  NANDN U4057 ( .A(n4025), .B(n4024), .Z(n4020) );
  ANDN U4058 ( .B(B[54]), .A(n37), .Z(n3913) );
  XNOR U4059 ( .A(n3921), .B(n4026), .Z(n3914) );
  XNOR U4060 ( .A(n3920), .B(n3918), .Z(n4026) );
  AND U4061 ( .A(n4027), .B(n4028), .Z(n3918) );
  NANDN U4062 ( .A(n4029), .B(n4030), .Z(n4028) );
  OR U4063 ( .A(n4031), .B(n4032), .Z(n4030) );
  NAND U4064 ( .A(n4032), .B(n4031), .Z(n4027) );
  ANDN U4065 ( .B(B[55]), .A(n38), .Z(n3920) );
  XNOR U4066 ( .A(n3928), .B(n4033), .Z(n3921) );
  XNOR U4067 ( .A(n3927), .B(n3925), .Z(n4033) );
  AND U4068 ( .A(n4034), .B(n4035), .Z(n3925) );
  NANDN U4069 ( .A(n4036), .B(n4037), .Z(n4035) );
  NANDN U4070 ( .A(n4038), .B(n4039), .Z(n4037) );
  NANDN U4071 ( .A(n4039), .B(n4038), .Z(n4034) );
  ANDN U4072 ( .B(B[56]), .A(n39), .Z(n3927) );
  XNOR U4073 ( .A(n3935), .B(n4040), .Z(n3928) );
  XNOR U4074 ( .A(n3934), .B(n3932), .Z(n4040) );
  AND U4075 ( .A(n4041), .B(n4042), .Z(n3932) );
  NANDN U4076 ( .A(n4043), .B(n4044), .Z(n4042) );
  OR U4077 ( .A(n4045), .B(n4046), .Z(n4044) );
  NAND U4078 ( .A(n4046), .B(n4045), .Z(n4041) );
  ANDN U4079 ( .B(B[57]), .A(n40), .Z(n3934) );
  XNOR U4080 ( .A(n3942), .B(n4047), .Z(n3935) );
  XNOR U4081 ( .A(n3941), .B(n3939), .Z(n4047) );
  AND U4082 ( .A(n4048), .B(n4049), .Z(n3939) );
  NANDN U4083 ( .A(n4050), .B(n4051), .Z(n4049) );
  NAND U4084 ( .A(n4052), .B(n4053), .Z(n4051) );
  ANDN U4085 ( .B(B[58]), .A(n41), .Z(n3941) );
  XOR U4086 ( .A(n3948), .B(n4054), .Z(n3942) );
  XNOR U4087 ( .A(n3946), .B(n3949), .Z(n4054) );
  NAND U4088 ( .A(A[2]), .B(B[59]), .Z(n3949) );
  NANDN U4089 ( .A(n4055), .B(n4056), .Z(n3946) );
  AND U4090 ( .A(A[0]), .B(B[60]), .Z(n4056) );
  XNOR U4091 ( .A(n3951), .B(n4057), .Z(n3948) );
  NAND U4092 ( .A(A[0]), .B(B[61]), .Z(n4057) );
  NAND U4093 ( .A(B[60]), .B(A[1]), .Z(n3951) );
  NAND U4094 ( .A(n4058), .B(n4059), .Z(n124) );
  NANDN U4095 ( .A(n4060), .B(n4061), .Z(n4059) );
  OR U4096 ( .A(n4062), .B(n4063), .Z(n4061) );
  NAND U4097 ( .A(n4063), .B(n4062), .Z(n4058) );
  XOR U4098 ( .A(n126), .B(n125), .Z(\A1[58] ) );
  XOR U4099 ( .A(n4063), .B(n4064), .Z(n125) );
  XNOR U4100 ( .A(n4062), .B(n4060), .Z(n4064) );
  AND U4101 ( .A(n4065), .B(n4066), .Z(n4060) );
  NANDN U4102 ( .A(n4067), .B(n4068), .Z(n4066) );
  NANDN U4103 ( .A(n4069), .B(n4070), .Z(n4068) );
  NANDN U4104 ( .A(n4070), .B(n4069), .Z(n4065) );
  ANDN U4105 ( .B(B[45]), .A(n29), .Z(n4062) );
  XNOR U4106 ( .A(n3969), .B(n4071), .Z(n4063) );
  XNOR U4107 ( .A(n3968), .B(n3966), .Z(n4071) );
  AND U4108 ( .A(n4072), .B(n4073), .Z(n3966) );
  NANDN U4109 ( .A(n4074), .B(n4075), .Z(n4073) );
  OR U4110 ( .A(n4076), .B(n4077), .Z(n4075) );
  NAND U4111 ( .A(n4077), .B(n4076), .Z(n4072) );
  ANDN U4112 ( .B(B[46]), .A(n30), .Z(n3968) );
  XNOR U4113 ( .A(n3976), .B(n4078), .Z(n3969) );
  XNOR U4114 ( .A(n3975), .B(n3973), .Z(n4078) );
  AND U4115 ( .A(n4079), .B(n4080), .Z(n3973) );
  NANDN U4116 ( .A(n4081), .B(n4082), .Z(n4080) );
  NANDN U4117 ( .A(n4083), .B(n4084), .Z(n4082) );
  NANDN U4118 ( .A(n4084), .B(n4083), .Z(n4079) );
  ANDN U4119 ( .B(B[47]), .A(n31), .Z(n3975) );
  XNOR U4120 ( .A(n3983), .B(n4085), .Z(n3976) );
  XNOR U4121 ( .A(n3982), .B(n3980), .Z(n4085) );
  AND U4122 ( .A(n4086), .B(n4087), .Z(n3980) );
  NANDN U4123 ( .A(n4088), .B(n4089), .Z(n4087) );
  OR U4124 ( .A(n4090), .B(n4091), .Z(n4089) );
  NAND U4125 ( .A(n4091), .B(n4090), .Z(n4086) );
  ANDN U4126 ( .B(B[48]), .A(n32), .Z(n3982) );
  XNOR U4127 ( .A(n3990), .B(n4092), .Z(n3983) );
  XNOR U4128 ( .A(n3989), .B(n3987), .Z(n4092) );
  AND U4129 ( .A(n4093), .B(n4094), .Z(n3987) );
  NANDN U4130 ( .A(n4095), .B(n4096), .Z(n4094) );
  NANDN U4131 ( .A(n4097), .B(n4098), .Z(n4096) );
  NANDN U4132 ( .A(n4098), .B(n4097), .Z(n4093) );
  ANDN U4133 ( .B(B[49]), .A(n33), .Z(n3989) );
  XNOR U4134 ( .A(n3997), .B(n4099), .Z(n3990) );
  XNOR U4135 ( .A(n3996), .B(n3994), .Z(n4099) );
  AND U4136 ( .A(n4100), .B(n4101), .Z(n3994) );
  NANDN U4137 ( .A(n4102), .B(n4103), .Z(n4101) );
  OR U4138 ( .A(n4104), .B(n4105), .Z(n4103) );
  NAND U4139 ( .A(n4105), .B(n4104), .Z(n4100) );
  ANDN U4140 ( .B(B[50]), .A(n34), .Z(n3996) );
  XNOR U4141 ( .A(n4004), .B(n4106), .Z(n3997) );
  XNOR U4142 ( .A(n4003), .B(n4001), .Z(n4106) );
  AND U4143 ( .A(n4107), .B(n4108), .Z(n4001) );
  NANDN U4144 ( .A(n4109), .B(n4110), .Z(n4108) );
  NANDN U4145 ( .A(n4111), .B(n4112), .Z(n4110) );
  NANDN U4146 ( .A(n4112), .B(n4111), .Z(n4107) );
  ANDN U4147 ( .B(B[51]), .A(n35), .Z(n4003) );
  XNOR U4148 ( .A(n4011), .B(n4113), .Z(n4004) );
  XNOR U4149 ( .A(n4010), .B(n4008), .Z(n4113) );
  AND U4150 ( .A(n4114), .B(n4115), .Z(n4008) );
  NANDN U4151 ( .A(n4116), .B(n4117), .Z(n4115) );
  OR U4152 ( .A(n4118), .B(n4119), .Z(n4117) );
  NAND U4153 ( .A(n4119), .B(n4118), .Z(n4114) );
  ANDN U4154 ( .B(B[52]), .A(n36), .Z(n4010) );
  XNOR U4155 ( .A(n4018), .B(n4120), .Z(n4011) );
  XNOR U4156 ( .A(n4017), .B(n4015), .Z(n4120) );
  AND U4157 ( .A(n4121), .B(n4122), .Z(n4015) );
  NANDN U4158 ( .A(n4123), .B(n4124), .Z(n4122) );
  NANDN U4159 ( .A(n4125), .B(n4126), .Z(n4124) );
  NANDN U4160 ( .A(n4126), .B(n4125), .Z(n4121) );
  ANDN U4161 ( .B(B[53]), .A(n37), .Z(n4017) );
  XNOR U4162 ( .A(n4025), .B(n4127), .Z(n4018) );
  XNOR U4163 ( .A(n4024), .B(n4022), .Z(n4127) );
  AND U4164 ( .A(n4128), .B(n4129), .Z(n4022) );
  NANDN U4165 ( .A(n4130), .B(n4131), .Z(n4129) );
  OR U4166 ( .A(n4132), .B(n4133), .Z(n4131) );
  NAND U4167 ( .A(n4133), .B(n4132), .Z(n4128) );
  ANDN U4168 ( .B(B[54]), .A(n38), .Z(n4024) );
  XNOR U4169 ( .A(n4032), .B(n4134), .Z(n4025) );
  XNOR U4170 ( .A(n4031), .B(n4029), .Z(n4134) );
  AND U4171 ( .A(n4135), .B(n4136), .Z(n4029) );
  NANDN U4172 ( .A(n4137), .B(n4138), .Z(n4136) );
  NANDN U4173 ( .A(n4139), .B(n4140), .Z(n4138) );
  NANDN U4174 ( .A(n4140), .B(n4139), .Z(n4135) );
  ANDN U4175 ( .B(B[55]), .A(n39), .Z(n4031) );
  XNOR U4176 ( .A(n4039), .B(n4141), .Z(n4032) );
  XNOR U4177 ( .A(n4038), .B(n4036), .Z(n4141) );
  AND U4178 ( .A(n4142), .B(n4143), .Z(n4036) );
  NANDN U4179 ( .A(n4144), .B(n4145), .Z(n4143) );
  OR U4180 ( .A(n4146), .B(n4147), .Z(n4145) );
  NAND U4181 ( .A(n4147), .B(n4146), .Z(n4142) );
  ANDN U4182 ( .B(B[56]), .A(n40), .Z(n4038) );
  XNOR U4183 ( .A(n4046), .B(n4148), .Z(n4039) );
  XNOR U4184 ( .A(n4045), .B(n4043), .Z(n4148) );
  AND U4185 ( .A(n4149), .B(n4150), .Z(n4043) );
  NANDN U4186 ( .A(n4151), .B(n4152), .Z(n4150) );
  NAND U4187 ( .A(n4153), .B(n4154), .Z(n4152) );
  ANDN U4188 ( .B(B[57]), .A(n41), .Z(n4045) );
  XOR U4189 ( .A(n4052), .B(n4155), .Z(n4046) );
  XNOR U4190 ( .A(n4050), .B(n4053), .Z(n4155) );
  NAND U4191 ( .A(A[2]), .B(B[58]), .Z(n4053) );
  NANDN U4192 ( .A(n4156), .B(n4157), .Z(n4050) );
  AND U4193 ( .A(A[0]), .B(B[59]), .Z(n4157) );
  XNOR U4194 ( .A(n4055), .B(n4158), .Z(n4052) );
  NAND U4195 ( .A(A[0]), .B(B[60]), .Z(n4158) );
  NAND U4196 ( .A(B[59]), .B(A[1]), .Z(n4055) );
  NAND U4197 ( .A(n4159), .B(n4160), .Z(n126) );
  NANDN U4198 ( .A(n4161), .B(n4162), .Z(n4160) );
  OR U4199 ( .A(n4163), .B(n4164), .Z(n4162) );
  NAND U4200 ( .A(n4164), .B(n4163), .Z(n4159) );
  XOR U4201 ( .A(n128), .B(n127), .Z(\A1[57] ) );
  XOR U4202 ( .A(n4164), .B(n4165), .Z(n127) );
  XNOR U4203 ( .A(n4163), .B(n4161), .Z(n4165) );
  AND U4204 ( .A(n4166), .B(n4167), .Z(n4161) );
  NANDN U4205 ( .A(n4168), .B(n4169), .Z(n4167) );
  NANDN U4206 ( .A(n4170), .B(n4171), .Z(n4169) );
  NANDN U4207 ( .A(n4171), .B(n4170), .Z(n4166) );
  ANDN U4208 ( .B(B[44]), .A(n29), .Z(n4163) );
  XNOR U4209 ( .A(n4070), .B(n4172), .Z(n4164) );
  XNOR U4210 ( .A(n4069), .B(n4067), .Z(n4172) );
  AND U4211 ( .A(n4173), .B(n4174), .Z(n4067) );
  NANDN U4212 ( .A(n4175), .B(n4176), .Z(n4174) );
  OR U4213 ( .A(n4177), .B(n4178), .Z(n4176) );
  NAND U4214 ( .A(n4178), .B(n4177), .Z(n4173) );
  ANDN U4215 ( .B(B[45]), .A(n30), .Z(n4069) );
  XNOR U4216 ( .A(n4077), .B(n4179), .Z(n4070) );
  XNOR U4217 ( .A(n4076), .B(n4074), .Z(n4179) );
  AND U4218 ( .A(n4180), .B(n4181), .Z(n4074) );
  NANDN U4219 ( .A(n4182), .B(n4183), .Z(n4181) );
  NANDN U4220 ( .A(n4184), .B(n4185), .Z(n4183) );
  NANDN U4221 ( .A(n4185), .B(n4184), .Z(n4180) );
  ANDN U4222 ( .B(B[46]), .A(n31), .Z(n4076) );
  XNOR U4223 ( .A(n4084), .B(n4186), .Z(n4077) );
  XNOR U4224 ( .A(n4083), .B(n4081), .Z(n4186) );
  AND U4225 ( .A(n4187), .B(n4188), .Z(n4081) );
  NANDN U4226 ( .A(n4189), .B(n4190), .Z(n4188) );
  OR U4227 ( .A(n4191), .B(n4192), .Z(n4190) );
  NAND U4228 ( .A(n4192), .B(n4191), .Z(n4187) );
  ANDN U4229 ( .B(B[47]), .A(n32), .Z(n4083) );
  XNOR U4230 ( .A(n4091), .B(n4193), .Z(n4084) );
  XNOR U4231 ( .A(n4090), .B(n4088), .Z(n4193) );
  AND U4232 ( .A(n4194), .B(n4195), .Z(n4088) );
  NANDN U4233 ( .A(n4196), .B(n4197), .Z(n4195) );
  NANDN U4234 ( .A(n4198), .B(n4199), .Z(n4197) );
  NANDN U4235 ( .A(n4199), .B(n4198), .Z(n4194) );
  ANDN U4236 ( .B(B[48]), .A(n33), .Z(n4090) );
  XNOR U4237 ( .A(n4098), .B(n4200), .Z(n4091) );
  XNOR U4238 ( .A(n4097), .B(n4095), .Z(n4200) );
  AND U4239 ( .A(n4201), .B(n4202), .Z(n4095) );
  NANDN U4240 ( .A(n4203), .B(n4204), .Z(n4202) );
  OR U4241 ( .A(n4205), .B(n4206), .Z(n4204) );
  NAND U4242 ( .A(n4206), .B(n4205), .Z(n4201) );
  ANDN U4243 ( .B(B[49]), .A(n34), .Z(n4097) );
  XNOR U4244 ( .A(n4105), .B(n4207), .Z(n4098) );
  XNOR U4245 ( .A(n4104), .B(n4102), .Z(n4207) );
  AND U4246 ( .A(n4208), .B(n4209), .Z(n4102) );
  NANDN U4247 ( .A(n4210), .B(n4211), .Z(n4209) );
  NANDN U4248 ( .A(n4212), .B(n4213), .Z(n4211) );
  NANDN U4249 ( .A(n4213), .B(n4212), .Z(n4208) );
  ANDN U4250 ( .B(B[50]), .A(n35), .Z(n4104) );
  XNOR U4251 ( .A(n4112), .B(n4214), .Z(n4105) );
  XNOR U4252 ( .A(n4111), .B(n4109), .Z(n4214) );
  AND U4253 ( .A(n4215), .B(n4216), .Z(n4109) );
  NANDN U4254 ( .A(n4217), .B(n4218), .Z(n4216) );
  OR U4255 ( .A(n4219), .B(n4220), .Z(n4218) );
  NAND U4256 ( .A(n4220), .B(n4219), .Z(n4215) );
  ANDN U4257 ( .B(B[51]), .A(n36), .Z(n4111) );
  XNOR U4258 ( .A(n4119), .B(n4221), .Z(n4112) );
  XNOR U4259 ( .A(n4118), .B(n4116), .Z(n4221) );
  AND U4260 ( .A(n4222), .B(n4223), .Z(n4116) );
  NANDN U4261 ( .A(n4224), .B(n4225), .Z(n4223) );
  NANDN U4262 ( .A(n4226), .B(n4227), .Z(n4225) );
  NANDN U4263 ( .A(n4227), .B(n4226), .Z(n4222) );
  ANDN U4264 ( .B(B[52]), .A(n37), .Z(n4118) );
  XNOR U4265 ( .A(n4126), .B(n4228), .Z(n4119) );
  XNOR U4266 ( .A(n4125), .B(n4123), .Z(n4228) );
  AND U4267 ( .A(n4229), .B(n4230), .Z(n4123) );
  NANDN U4268 ( .A(n4231), .B(n4232), .Z(n4230) );
  OR U4269 ( .A(n4233), .B(n4234), .Z(n4232) );
  NAND U4270 ( .A(n4234), .B(n4233), .Z(n4229) );
  ANDN U4271 ( .B(B[53]), .A(n38), .Z(n4125) );
  XNOR U4272 ( .A(n4133), .B(n4235), .Z(n4126) );
  XNOR U4273 ( .A(n4132), .B(n4130), .Z(n4235) );
  AND U4274 ( .A(n4236), .B(n4237), .Z(n4130) );
  NANDN U4275 ( .A(n4238), .B(n4239), .Z(n4237) );
  NANDN U4276 ( .A(n4240), .B(n4241), .Z(n4239) );
  NANDN U4277 ( .A(n4241), .B(n4240), .Z(n4236) );
  ANDN U4278 ( .B(B[54]), .A(n39), .Z(n4132) );
  XNOR U4279 ( .A(n4140), .B(n4242), .Z(n4133) );
  XNOR U4280 ( .A(n4139), .B(n4137), .Z(n4242) );
  AND U4281 ( .A(n4243), .B(n4244), .Z(n4137) );
  NANDN U4282 ( .A(n4245), .B(n4246), .Z(n4244) );
  OR U4283 ( .A(n4247), .B(n4248), .Z(n4246) );
  NAND U4284 ( .A(n4248), .B(n4247), .Z(n4243) );
  ANDN U4285 ( .B(B[55]), .A(n40), .Z(n4139) );
  XNOR U4286 ( .A(n4147), .B(n4249), .Z(n4140) );
  XNOR U4287 ( .A(n4146), .B(n4144), .Z(n4249) );
  AND U4288 ( .A(n4250), .B(n4251), .Z(n4144) );
  NANDN U4289 ( .A(n4252), .B(n4253), .Z(n4251) );
  NAND U4290 ( .A(n4254), .B(n4255), .Z(n4253) );
  ANDN U4291 ( .B(B[56]), .A(n41), .Z(n4146) );
  XOR U4292 ( .A(n4153), .B(n4256), .Z(n4147) );
  XNOR U4293 ( .A(n4151), .B(n4154), .Z(n4256) );
  NAND U4294 ( .A(A[2]), .B(B[57]), .Z(n4154) );
  NANDN U4295 ( .A(n4257), .B(n4258), .Z(n4151) );
  AND U4296 ( .A(A[0]), .B(B[58]), .Z(n4258) );
  XNOR U4297 ( .A(n4156), .B(n4259), .Z(n4153) );
  NAND U4298 ( .A(A[0]), .B(B[59]), .Z(n4259) );
  NAND U4299 ( .A(B[58]), .B(A[1]), .Z(n4156) );
  NAND U4300 ( .A(n4260), .B(n4261), .Z(n128) );
  NANDN U4301 ( .A(n4262), .B(n4263), .Z(n4261) );
  OR U4302 ( .A(n4264), .B(n4265), .Z(n4263) );
  NAND U4303 ( .A(n4265), .B(n4264), .Z(n4260) );
  XOR U4304 ( .A(n130), .B(n129), .Z(\A1[56] ) );
  XOR U4305 ( .A(n4265), .B(n4266), .Z(n129) );
  XNOR U4306 ( .A(n4264), .B(n4262), .Z(n4266) );
  AND U4307 ( .A(n4267), .B(n4268), .Z(n4262) );
  NANDN U4308 ( .A(n4269), .B(n4270), .Z(n4268) );
  NANDN U4309 ( .A(n4271), .B(n4272), .Z(n4270) );
  NANDN U4310 ( .A(n4272), .B(n4271), .Z(n4267) );
  ANDN U4311 ( .B(B[43]), .A(n29), .Z(n4264) );
  XNOR U4312 ( .A(n4171), .B(n4273), .Z(n4265) );
  XNOR U4313 ( .A(n4170), .B(n4168), .Z(n4273) );
  AND U4314 ( .A(n4274), .B(n4275), .Z(n4168) );
  NANDN U4315 ( .A(n4276), .B(n4277), .Z(n4275) );
  OR U4316 ( .A(n4278), .B(n4279), .Z(n4277) );
  NAND U4317 ( .A(n4279), .B(n4278), .Z(n4274) );
  ANDN U4318 ( .B(B[44]), .A(n30), .Z(n4170) );
  XNOR U4319 ( .A(n4178), .B(n4280), .Z(n4171) );
  XNOR U4320 ( .A(n4177), .B(n4175), .Z(n4280) );
  AND U4321 ( .A(n4281), .B(n4282), .Z(n4175) );
  NANDN U4322 ( .A(n4283), .B(n4284), .Z(n4282) );
  NANDN U4323 ( .A(n4285), .B(n4286), .Z(n4284) );
  NANDN U4324 ( .A(n4286), .B(n4285), .Z(n4281) );
  ANDN U4325 ( .B(B[45]), .A(n31), .Z(n4177) );
  XNOR U4326 ( .A(n4185), .B(n4287), .Z(n4178) );
  XNOR U4327 ( .A(n4184), .B(n4182), .Z(n4287) );
  AND U4328 ( .A(n4288), .B(n4289), .Z(n4182) );
  NANDN U4329 ( .A(n4290), .B(n4291), .Z(n4289) );
  OR U4330 ( .A(n4292), .B(n4293), .Z(n4291) );
  NAND U4331 ( .A(n4293), .B(n4292), .Z(n4288) );
  ANDN U4332 ( .B(B[46]), .A(n32), .Z(n4184) );
  XNOR U4333 ( .A(n4192), .B(n4294), .Z(n4185) );
  XNOR U4334 ( .A(n4191), .B(n4189), .Z(n4294) );
  AND U4335 ( .A(n4295), .B(n4296), .Z(n4189) );
  NANDN U4336 ( .A(n4297), .B(n4298), .Z(n4296) );
  NANDN U4337 ( .A(n4299), .B(n4300), .Z(n4298) );
  NANDN U4338 ( .A(n4300), .B(n4299), .Z(n4295) );
  ANDN U4339 ( .B(B[47]), .A(n33), .Z(n4191) );
  XNOR U4340 ( .A(n4199), .B(n4301), .Z(n4192) );
  XNOR U4341 ( .A(n4198), .B(n4196), .Z(n4301) );
  AND U4342 ( .A(n4302), .B(n4303), .Z(n4196) );
  NANDN U4343 ( .A(n4304), .B(n4305), .Z(n4303) );
  OR U4344 ( .A(n4306), .B(n4307), .Z(n4305) );
  NAND U4345 ( .A(n4307), .B(n4306), .Z(n4302) );
  ANDN U4346 ( .B(B[48]), .A(n34), .Z(n4198) );
  XNOR U4347 ( .A(n4206), .B(n4308), .Z(n4199) );
  XNOR U4348 ( .A(n4205), .B(n4203), .Z(n4308) );
  AND U4349 ( .A(n4309), .B(n4310), .Z(n4203) );
  NANDN U4350 ( .A(n4311), .B(n4312), .Z(n4310) );
  NANDN U4351 ( .A(n4313), .B(n4314), .Z(n4312) );
  NANDN U4352 ( .A(n4314), .B(n4313), .Z(n4309) );
  ANDN U4353 ( .B(B[49]), .A(n35), .Z(n4205) );
  XNOR U4354 ( .A(n4213), .B(n4315), .Z(n4206) );
  XNOR U4355 ( .A(n4212), .B(n4210), .Z(n4315) );
  AND U4356 ( .A(n4316), .B(n4317), .Z(n4210) );
  NANDN U4357 ( .A(n4318), .B(n4319), .Z(n4317) );
  OR U4358 ( .A(n4320), .B(n4321), .Z(n4319) );
  NAND U4359 ( .A(n4321), .B(n4320), .Z(n4316) );
  ANDN U4360 ( .B(B[50]), .A(n36), .Z(n4212) );
  XNOR U4361 ( .A(n4220), .B(n4322), .Z(n4213) );
  XNOR U4362 ( .A(n4219), .B(n4217), .Z(n4322) );
  AND U4363 ( .A(n4323), .B(n4324), .Z(n4217) );
  NANDN U4364 ( .A(n4325), .B(n4326), .Z(n4324) );
  NANDN U4365 ( .A(n4327), .B(n4328), .Z(n4326) );
  NANDN U4366 ( .A(n4328), .B(n4327), .Z(n4323) );
  ANDN U4367 ( .B(B[51]), .A(n37), .Z(n4219) );
  XNOR U4368 ( .A(n4227), .B(n4329), .Z(n4220) );
  XNOR U4369 ( .A(n4226), .B(n4224), .Z(n4329) );
  AND U4370 ( .A(n4330), .B(n4331), .Z(n4224) );
  NANDN U4371 ( .A(n4332), .B(n4333), .Z(n4331) );
  OR U4372 ( .A(n4334), .B(n4335), .Z(n4333) );
  NAND U4373 ( .A(n4335), .B(n4334), .Z(n4330) );
  ANDN U4374 ( .B(B[52]), .A(n38), .Z(n4226) );
  XNOR U4375 ( .A(n4234), .B(n4336), .Z(n4227) );
  XNOR U4376 ( .A(n4233), .B(n4231), .Z(n4336) );
  AND U4377 ( .A(n4337), .B(n4338), .Z(n4231) );
  NANDN U4378 ( .A(n4339), .B(n4340), .Z(n4338) );
  NANDN U4379 ( .A(n4341), .B(n4342), .Z(n4340) );
  NANDN U4380 ( .A(n4342), .B(n4341), .Z(n4337) );
  ANDN U4381 ( .B(B[53]), .A(n39), .Z(n4233) );
  XNOR U4382 ( .A(n4241), .B(n4343), .Z(n4234) );
  XNOR U4383 ( .A(n4240), .B(n4238), .Z(n4343) );
  AND U4384 ( .A(n4344), .B(n4345), .Z(n4238) );
  NANDN U4385 ( .A(n4346), .B(n4347), .Z(n4345) );
  OR U4386 ( .A(n4348), .B(n4349), .Z(n4347) );
  NAND U4387 ( .A(n4349), .B(n4348), .Z(n4344) );
  ANDN U4388 ( .B(B[54]), .A(n40), .Z(n4240) );
  XNOR U4389 ( .A(n4248), .B(n4350), .Z(n4241) );
  XNOR U4390 ( .A(n4247), .B(n4245), .Z(n4350) );
  AND U4391 ( .A(n4351), .B(n4352), .Z(n4245) );
  NANDN U4392 ( .A(n4353), .B(n4354), .Z(n4352) );
  NAND U4393 ( .A(n4355), .B(n4356), .Z(n4354) );
  ANDN U4394 ( .B(B[55]), .A(n41), .Z(n4247) );
  XOR U4395 ( .A(n4254), .B(n4357), .Z(n4248) );
  XNOR U4396 ( .A(n4252), .B(n4255), .Z(n4357) );
  NAND U4397 ( .A(A[2]), .B(B[56]), .Z(n4255) );
  NANDN U4398 ( .A(n4358), .B(n4359), .Z(n4252) );
  AND U4399 ( .A(A[0]), .B(B[57]), .Z(n4359) );
  XNOR U4400 ( .A(n4257), .B(n4360), .Z(n4254) );
  NAND U4401 ( .A(A[0]), .B(B[58]), .Z(n4360) );
  NAND U4402 ( .A(B[57]), .B(A[1]), .Z(n4257) );
  NAND U4403 ( .A(n4361), .B(n4362), .Z(n130) );
  NANDN U4404 ( .A(n4363), .B(n4364), .Z(n4362) );
  OR U4405 ( .A(n4365), .B(n4366), .Z(n4364) );
  NAND U4406 ( .A(n4366), .B(n4365), .Z(n4361) );
  XOR U4407 ( .A(n132), .B(n131), .Z(\A1[55] ) );
  XOR U4408 ( .A(n4366), .B(n4367), .Z(n131) );
  XNOR U4409 ( .A(n4365), .B(n4363), .Z(n4367) );
  AND U4410 ( .A(n4368), .B(n4369), .Z(n4363) );
  NANDN U4411 ( .A(n4370), .B(n4371), .Z(n4369) );
  NANDN U4412 ( .A(n4372), .B(n4373), .Z(n4371) );
  NANDN U4413 ( .A(n4373), .B(n4372), .Z(n4368) );
  ANDN U4414 ( .B(B[42]), .A(n29), .Z(n4365) );
  XNOR U4415 ( .A(n4272), .B(n4374), .Z(n4366) );
  XNOR U4416 ( .A(n4271), .B(n4269), .Z(n4374) );
  AND U4417 ( .A(n4375), .B(n4376), .Z(n4269) );
  NANDN U4418 ( .A(n4377), .B(n4378), .Z(n4376) );
  OR U4419 ( .A(n4379), .B(n4380), .Z(n4378) );
  NAND U4420 ( .A(n4380), .B(n4379), .Z(n4375) );
  ANDN U4421 ( .B(B[43]), .A(n30), .Z(n4271) );
  XNOR U4422 ( .A(n4279), .B(n4381), .Z(n4272) );
  XNOR U4423 ( .A(n4278), .B(n4276), .Z(n4381) );
  AND U4424 ( .A(n4382), .B(n4383), .Z(n4276) );
  NANDN U4425 ( .A(n4384), .B(n4385), .Z(n4383) );
  NANDN U4426 ( .A(n4386), .B(n4387), .Z(n4385) );
  NANDN U4427 ( .A(n4387), .B(n4386), .Z(n4382) );
  ANDN U4428 ( .B(B[44]), .A(n31), .Z(n4278) );
  XNOR U4429 ( .A(n4286), .B(n4388), .Z(n4279) );
  XNOR U4430 ( .A(n4285), .B(n4283), .Z(n4388) );
  AND U4431 ( .A(n4389), .B(n4390), .Z(n4283) );
  NANDN U4432 ( .A(n4391), .B(n4392), .Z(n4390) );
  OR U4433 ( .A(n4393), .B(n4394), .Z(n4392) );
  NAND U4434 ( .A(n4394), .B(n4393), .Z(n4389) );
  ANDN U4435 ( .B(B[45]), .A(n32), .Z(n4285) );
  XNOR U4436 ( .A(n4293), .B(n4395), .Z(n4286) );
  XNOR U4437 ( .A(n4292), .B(n4290), .Z(n4395) );
  AND U4438 ( .A(n4396), .B(n4397), .Z(n4290) );
  NANDN U4439 ( .A(n4398), .B(n4399), .Z(n4397) );
  NANDN U4440 ( .A(n4400), .B(n4401), .Z(n4399) );
  NANDN U4441 ( .A(n4401), .B(n4400), .Z(n4396) );
  ANDN U4442 ( .B(B[46]), .A(n33), .Z(n4292) );
  XNOR U4443 ( .A(n4300), .B(n4402), .Z(n4293) );
  XNOR U4444 ( .A(n4299), .B(n4297), .Z(n4402) );
  AND U4445 ( .A(n4403), .B(n4404), .Z(n4297) );
  NANDN U4446 ( .A(n4405), .B(n4406), .Z(n4404) );
  OR U4447 ( .A(n4407), .B(n4408), .Z(n4406) );
  NAND U4448 ( .A(n4408), .B(n4407), .Z(n4403) );
  ANDN U4449 ( .B(B[47]), .A(n34), .Z(n4299) );
  XNOR U4450 ( .A(n4307), .B(n4409), .Z(n4300) );
  XNOR U4451 ( .A(n4306), .B(n4304), .Z(n4409) );
  AND U4452 ( .A(n4410), .B(n4411), .Z(n4304) );
  NANDN U4453 ( .A(n4412), .B(n4413), .Z(n4411) );
  NANDN U4454 ( .A(n4414), .B(n4415), .Z(n4413) );
  NANDN U4455 ( .A(n4415), .B(n4414), .Z(n4410) );
  ANDN U4456 ( .B(B[48]), .A(n35), .Z(n4306) );
  XNOR U4457 ( .A(n4314), .B(n4416), .Z(n4307) );
  XNOR U4458 ( .A(n4313), .B(n4311), .Z(n4416) );
  AND U4459 ( .A(n4417), .B(n4418), .Z(n4311) );
  NANDN U4460 ( .A(n4419), .B(n4420), .Z(n4418) );
  OR U4461 ( .A(n4421), .B(n4422), .Z(n4420) );
  NAND U4462 ( .A(n4422), .B(n4421), .Z(n4417) );
  ANDN U4463 ( .B(B[49]), .A(n36), .Z(n4313) );
  XNOR U4464 ( .A(n4321), .B(n4423), .Z(n4314) );
  XNOR U4465 ( .A(n4320), .B(n4318), .Z(n4423) );
  AND U4466 ( .A(n4424), .B(n4425), .Z(n4318) );
  NANDN U4467 ( .A(n4426), .B(n4427), .Z(n4425) );
  NANDN U4468 ( .A(n4428), .B(n4429), .Z(n4427) );
  NANDN U4469 ( .A(n4429), .B(n4428), .Z(n4424) );
  ANDN U4470 ( .B(B[50]), .A(n37), .Z(n4320) );
  XNOR U4471 ( .A(n4328), .B(n4430), .Z(n4321) );
  XNOR U4472 ( .A(n4327), .B(n4325), .Z(n4430) );
  AND U4473 ( .A(n4431), .B(n4432), .Z(n4325) );
  NANDN U4474 ( .A(n4433), .B(n4434), .Z(n4432) );
  OR U4475 ( .A(n4435), .B(n4436), .Z(n4434) );
  NAND U4476 ( .A(n4436), .B(n4435), .Z(n4431) );
  ANDN U4477 ( .B(B[51]), .A(n38), .Z(n4327) );
  XNOR U4478 ( .A(n4335), .B(n4437), .Z(n4328) );
  XNOR U4479 ( .A(n4334), .B(n4332), .Z(n4437) );
  AND U4480 ( .A(n4438), .B(n4439), .Z(n4332) );
  NANDN U4481 ( .A(n4440), .B(n4441), .Z(n4439) );
  NANDN U4482 ( .A(n4442), .B(n4443), .Z(n4441) );
  NANDN U4483 ( .A(n4443), .B(n4442), .Z(n4438) );
  ANDN U4484 ( .B(B[52]), .A(n39), .Z(n4334) );
  XNOR U4485 ( .A(n4342), .B(n4444), .Z(n4335) );
  XNOR U4486 ( .A(n4341), .B(n4339), .Z(n4444) );
  AND U4487 ( .A(n4445), .B(n4446), .Z(n4339) );
  NANDN U4488 ( .A(n4447), .B(n4448), .Z(n4446) );
  OR U4489 ( .A(n4449), .B(n4450), .Z(n4448) );
  NAND U4490 ( .A(n4450), .B(n4449), .Z(n4445) );
  ANDN U4491 ( .B(B[53]), .A(n40), .Z(n4341) );
  XNOR U4492 ( .A(n4349), .B(n4451), .Z(n4342) );
  XNOR U4493 ( .A(n4348), .B(n4346), .Z(n4451) );
  AND U4494 ( .A(n4452), .B(n4453), .Z(n4346) );
  NANDN U4495 ( .A(n4454), .B(n4455), .Z(n4453) );
  NAND U4496 ( .A(n4456), .B(n4457), .Z(n4455) );
  ANDN U4497 ( .B(B[54]), .A(n41), .Z(n4348) );
  XOR U4498 ( .A(n4355), .B(n4458), .Z(n4349) );
  XNOR U4499 ( .A(n4353), .B(n4356), .Z(n4458) );
  NAND U4500 ( .A(A[2]), .B(B[55]), .Z(n4356) );
  NANDN U4501 ( .A(n4459), .B(n4460), .Z(n4353) );
  AND U4502 ( .A(A[0]), .B(B[56]), .Z(n4460) );
  XNOR U4503 ( .A(n4358), .B(n4461), .Z(n4355) );
  NAND U4504 ( .A(A[0]), .B(B[57]), .Z(n4461) );
  NAND U4505 ( .A(B[56]), .B(A[1]), .Z(n4358) );
  NAND U4506 ( .A(n4462), .B(n4463), .Z(n132) );
  NANDN U4507 ( .A(n4464), .B(n4465), .Z(n4463) );
  OR U4508 ( .A(n4466), .B(n4467), .Z(n4465) );
  NAND U4509 ( .A(n4467), .B(n4466), .Z(n4462) );
  XOR U4510 ( .A(n134), .B(n133), .Z(\A1[54] ) );
  XOR U4511 ( .A(n4467), .B(n4468), .Z(n133) );
  XNOR U4512 ( .A(n4466), .B(n4464), .Z(n4468) );
  AND U4513 ( .A(n4469), .B(n4470), .Z(n4464) );
  NANDN U4514 ( .A(n4471), .B(n4472), .Z(n4470) );
  NANDN U4515 ( .A(n4473), .B(n4474), .Z(n4472) );
  NANDN U4516 ( .A(n4474), .B(n4473), .Z(n4469) );
  ANDN U4517 ( .B(B[41]), .A(n29), .Z(n4466) );
  XNOR U4518 ( .A(n4373), .B(n4475), .Z(n4467) );
  XNOR U4519 ( .A(n4372), .B(n4370), .Z(n4475) );
  AND U4520 ( .A(n4476), .B(n4477), .Z(n4370) );
  NANDN U4521 ( .A(n4478), .B(n4479), .Z(n4477) );
  OR U4522 ( .A(n4480), .B(n4481), .Z(n4479) );
  NAND U4523 ( .A(n4481), .B(n4480), .Z(n4476) );
  ANDN U4524 ( .B(B[42]), .A(n30), .Z(n4372) );
  XNOR U4525 ( .A(n4380), .B(n4482), .Z(n4373) );
  XNOR U4526 ( .A(n4379), .B(n4377), .Z(n4482) );
  AND U4527 ( .A(n4483), .B(n4484), .Z(n4377) );
  NANDN U4528 ( .A(n4485), .B(n4486), .Z(n4484) );
  NANDN U4529 ( .A(n4487), .B(n4488), .Z(n4486) );
  NANDN U4530 ( .A(n4488), .B(n4487), .Z(n4483) );
  ANDN U4531 ( .B(B[43]), .A(n31), .Z(n4379) );
  XNOR U4532 ( .A(n4387), .B(n4489), .Z(n4380) );
  XNOR U4533 ( .A(n4386), .B(n4384), .Z(n4489) );
  AND U4534 ( .A(n4490), .B(n4491), .Z(n4384) );
  NANDN U4535 ( .A(n4492), .B(n4493), .Z(n4491) );
  OR U4536 ( .A(n4494), .B(n4495), .Z(n4493) );
  NAND U4537 ( .A(n4495), .B(n4494), .Z(n4490) );
  ANDN U4538 ( .B(B[44]), .A(n32), .Z(n4386) );
  XNOR U4539 ( .A(n4394), .B(n4496), .Z(n4387) );
  XNOR U4540 ( .A(n4393), .B(n4391), .Z(n4496) );
  AND U4541 ( .A(n4497), .B(n4498), .Z(n4391) );
  NANDN U4542 ( .A(n4499), .B(n4500), .Z(n4498) );
  NANDN U4543 ( .A(n4501), .B(n4502), .Z(n4500) );
  NANDN U4544 ( .A(n4502), .B(n4501), .Z(n4497) );
  ANDN U4545 ( .B(B[45]), .A(n33), .Z(n4393) );
  XNOR U4546 ( .A(n4401), .B(n4503), .Z(n4394) );
  XNOR U4547 ( .A(n4400), .B(n4398), .Z(n4503) );
  AND U4548 ( .A(n4504), .B(n4505), .Z(n4398) );
  NANDN U4549 ( .A(n4506), .B(n4507), .Z(n4505) );
  OR U4550 ( .A(n4508), .B(n4509), .Z(n4507) );
  NAND U4551 ( .A(n4509), .B(n4508), .Z(n4504) );
  ANDN U4552 ( .B(B[46]), .A(n34), .Z(n4400) );
  XNOR U4553 ( .A(n4408), .B(n4510), .Z(n4401) );
  XNOR U4554 ( .A(n4407), .B(n4405), .Z(n4510) );
  AND U4555 ( .A(n4511), .B(n4512), .Z(n4405) );
  NANDN U4556 ( .A(n4513), .B(n4514), .Z(n4512) );
  NANDN U4557 ( .A(n4515), .B(n4516), .Z(n4514) );
  NANDN U4558 ( .A(n4516), .B(n4515), .Z(n4511) );
  ANDN U4559 ( .B(B[47]), .A(n35), .Z(n4407) );
  XNOR U4560 ( .A(n4415), .B(n4517), .Z(n4408) );
  XNOR U4561 ( .A(n4414), .B(n4412), .Z(n4517) );
  AND U4562 ( .A(n4518), .B(n4519), .Z(n4412) );
  NANDN U4563 ( .A(n4520), .B(n4521), .Z(n4519) );
  OR U4564 ( .A(n4522), .B(n4523), .Z(n4521) );
  NAND U4565 ( .A(n4523), .B(n4522), .Z(n4518) );
  ANDN U4566 ( .B(B[48]), .A(n36), .Z(n4414) );
  XNOR U4567 ( .A(n4422), .B(n4524), .Z(n4415) );
  XNOR U4568 ( .A(n4421), .B(n4419), .Z(n4524) );
  AND U4569 ( .A(n4525), .B(n4526), .Z(n4419) );
  NANDN U4570 ( .A(n4527), .B(n4528), .Z(n4526) );
  NANDN U4571 ( .A(n4529), .B(n4530), .Z(n4528) );
  NANDN U4572 ( .A(n4530), .B(n4529), .Z(n4525) );
  ANDN U4573 ( .B(B[49]), .A(n37), .Z(n4421) );
  XNOR U4574 ( .A(n4429), .B(n4531), .Z(n4422) );
  XNOR U4575 ( .A(n4428), .B(n4426), .Z(n4531) );
  AND U4576 ( .A(n4532), .B(n4533), .Z(n4426) );
  NANDN U4577 ( .A(n4534), .B(n4535), .Z(n4533) );
  OR U4578 ( .A(n4536), .B(n4537), .Z(n4535) );
  NAND U4579 ( .A(n4537), .B(n4536), .Z(n4532) );
  ANDN U4580 ( .B(B[50]), .A(n38), .Z(n4428) );
  XNOR U4581 ( .A(n4436), .B(n4538), .Z(n4429) );
  XNOR U4582 ( .A(n4435), .B(n4433), .Z(n4538) );
  AND U4583 ( .A(n4539), .B(n4540), .Z(n4433) );
  NANDN U4584 ( .A(n4541), .B(n4542), .Z(n4540) );
  NANDN U4585 ( .A(n4543), .B(n4544), .Z(n4542) );
  NANDN U4586 ( .A(n4544), .B(n4543), .Z(n4539) );
  ANDN U4587 ( .B(B[51]), .A(n39), .Z(n4435) );
  XNOR U4588 ( .A(n4443), .B(n4545), .Z(n4436) );
  XNOR U4589 ( .A(n4442), .B(n4440), .Z(n4545) );
  AND U4590 ( .A(n4546), .B(n4547), .Z(n4440) );
  NANDN U4591 ( .A(n4548), .B(n4549), .Z(n4547) );
  OR U4592 ( .A(n4550), .B(n4551), .Z(n4549) );
  NAND U4593 ( .A(n4551), .B(n4550), .Z(n4546) );
  ANDN U4594 ( .B(B[52]), .A(n40), .Z(n4442) );
  XNOR U4595 ( .A(n4450), .B(n4552), .Z(n4443) );
  XNOR U4596 ( .A(n4449), .B(n4447), .Z(n4552) );
  AND U4597 ( .A(n4553), .B(n4554), .Z(n4447) );
  NANDN U4598 ( .A(n4555), .B(n4556), .Z(n4554) );
  NAND U4599 ( .A(n4557), .B(n4558), .Z(n4556) );
  ANDN U4600 ( .B(B[53]), .A(n41), .Z(n4449) );
  XOR U4601 ( .A(n4456), .B(n4559), .Z(n4450) );
  XNOR U4602 ( .A(n4454), .B(n4457), .Z(n4559) );
  NAND U4603 ( .A(A[2]), .B(B[54]), .Z(n4457) );
  NANDN U4604 ( .A(n4560), .B(n4561), .Z(n4454) );
  AND U4605 ( .A(A[0]), .B(B[55]), .Z(n4561) );
  XNOR U4606 ( .A(n4459), .B(n4562), .Z(n4456) );
  NAND U4607 ( .A(A[0]), .B(B[56]), .Z(n4562) );
  NAND U4608 ( .A(B[55]), .B(A[1]), .Z(n4459) );
  NAND U4609 ( .A(n4563), .B(n4564), .Z(n134) );
  NANDN U4610 ( .A(n4565), .B(n4566), .Z(n4564) );
  OR U4611 ( .A(n4567), .B(n4568), .Z(n4566) );
  NAND U4612 ( .A(n4568), .B(n4567), .Z(n4563) );
  XOR U4613 ( .A(n136), .B(n135), .Z(\A1[53] ) );
  XOR U4614 ( .A(n4568), .B(n4569), .Z(n135) );
  XNOR U4615 ( .A(n4567), .B(n4565), .Z(n4569) );
  AND U4616 ( .A(n4570), .B(n4571), .Z(n4565) );
  NANDN U4617 ( .A(n4572), .B(n4573), .Z(n4571) );
  NANDN U4618 ( .A(n4574), .B(n4575), .Z(n4573) );
  NANDN U4619 ( .A(n4575), .B(n4574), .Z(n4570) );
  ANDN U4620 ( .B(B[40]), .A(n29), .Z(n4567) );
  XNOR U4621 ( .A(n4474), .B(n4576), .Z(n4568) );
  XNOR U4622 ( .A(n4473), .B(n4471), .Z(n4576) );
  AND U4623 ( .A(n4577), .B(n4578), .Z(n4471) );
  NANDN U4624 ( .A(n4579), .B(n4580), .Z(n4578) );
  OR U4625 ( .A(n4581), .B(n4582), .Z(n4580) );
  NAND U4626 ( .A(n4582), .B(n4581), .Z(n4577) );
  ANDN U4627 ( .B(B[41]), .A(n30), .Z(n4473) );
  XNOR U4628 ( .A(n4481), .B(n4583), .Z(n4474) );
  XNOR U4629 ( .A(n4480), .B(n4478), .Z(n4583) );
  AND U4630 ( .A(n4584), .B(n4585), .Z(n4478) );
  NANDN U4631 ( .A(n4586), .B(n4587), .Z(n4585) );
  NANDN U4632 ( .A(n4588), .B(n4589), .Z(n4587) );
  NANDN U4633 ( .A(n4589), .B(n4588), .Z(n4584) );
  ANDN U4634 ( .B(B[42]), .A(n31), .Z(n4480) );
  XNOR U4635 ( .A(n4488), .B(n4590), .Z(n4481) );
  XNOR U4636 ( .A(n4487), .B(n4485), .Z(n4590) );
  AND U4637 ( .A(n4591), .B(n4592), .Z(n4485) );
  NANDN U4638 ( .A(n4593), .B(n4594), .Z(n4592) );
  OR U4639 ( .A(n4595), .B(n4596), .Z(n4594) );
  NAND U4640 ( .A(n4596), .B(n4595), .Z(n4591) );
  ANDN U4641 ( .B(B[43]), .A(n32), .Z(n4487) );
  XNOR U4642 ( .A(n4495), .B(n4597), .Z(n4488) );
  XNOR U4643 ( .A(n4494), .B(n4492), .Z(n4597) );
  AND U4644 ( .A(n4598), .B(n4599), .Z(n4492) );
  NANDN U4645 ( .A(n4600), .B(n4601), .Z(n4599) );
  NANDN U4646 ( .A(n4602), .B(n4603), .Z(n4601) );
  NANDN U4647 ( .A(n4603), .B(n4602), .Z(n4598) );
  ANDN U4648 ( .B(B[44]), .A(n33), .Z(n4494) );
  XNOR U4649 ( .A(n4502), .B(n4604), .Z(n4495) );
  XNOR U4650 ( .A(n4501), .B(n4499), .Z(n4604) );
  AND U4651 ( .A(n4605), .B(n4606), .Z(n4499) );
  NANDN U4652 ( .A(n4607), .B(n4608), .Z(n4606) );
  OR U4653 ( .A(n4609), .B(n4610), .Z(n4608) );
  NAND U4654 ( .A(n4610), .B(n4609), .Z(n4605) );
  ANDN U4655 ( .B(B[45]), .A(n34), .Z(n4501) );
  XNOR U4656 ( .A(n4509), .B(n4611), .Z(n4502) );
  XNOR U4657 ( .A(n4508), .B(n4506), .Z(n4611) );
  AND U4658 ( .A(n4612), .B(n4613), .Z(n4506) );
  NANDN U4659 ( .A(n4614), .B(n4615), .Z(n4613) );
  NANDN U4660 ( .A(n4616), .B(n4617), .Z(n4615) );
  NANDN U4661 ( .A(n4617), .B(n4616), .Z(n4612) );
  ANDN U4662 ( .B(B[46]), .A(n35), .Z(n4508) );
  XNOR U4663 ( .A(n4516), .B(n4618), .Z(n4509) );
  XNOR U4664 ( .A(n4515), .B(n4513), .Z(n4618) );
  AND U4665 ( .A(n4619), .B(n4620), .Z(n4513) );
  NANDN U4666 ( .A(n4621), .B(n4622), .Z(n4620) );
  OR U4667 ( .A(n4623), .B(n4624), .Z(n4622) );
  NAND U4668 ( .A(n4624), .B(n4623), .Z(n4619) );
  ANDN U4669 ( .B(B[47]), .A(n36), .Z(n4515) );
  XNOR U4670 ( .A(n4523), .B(n4625), .Z(n4516) );
  XNOR U4671 ( .A(n4522), .B(n4520), .Z(n4625) );
  AND U4672 ( .A(n4626), .B(n4627), .Z(n4520) );
  NANDN U4673 ( .A(n4628), .B(n4629), .Z(n4627) );
  NANDN U4674 ( .A(n4630), .B(n4631), .Z(n4629) );
  NANDN U4675 ( .A(n4631), .B(n4630), .Z(n4626) );
  ANDN U4676 ( .B(B[48]), .A(n37), .Z(n4522) );
  XNOR U4677 ( .A(n4530), .B(n4632), .Z(n4523) );
  XNOR U4678 ( .A(n4529), .B(n4527), .Z(n4632) );
  AND U4679 ( .A(n4633), .B(n4634), .Z(n4527) );
  NANDN U4680 ( .A(n4635), .B(n4636), .Z(n4634) );
  OR U4681 ( .A(n4637), .B(n4638), .Z(n4636) );
  NAND U4682 ( .A(n4638), .B(n4637), .Z(n4633) );
  ANDN U4683 ( .B(B[49]), .A(n38), .Z(n4529) );
  XNOR U4684 ( .A(n4537), .B(n4639), .Z(n4530) );
  XNOR U4685 ( .A(n4536), .B(n4534), .Z(n4639) );
  AND U4686 ( .A(n4640), .B(n4641), .Z(n4534) );
  NANDN U4687 ( .A(n4642), .B(n4643), .Z(n4641) );
  NANDN U4688 ( .A(n4644), .B(n4645), .Z(n4643) );
  NANDN U4689 ( .A(n4645), .B(n4644), .Z(n4640) );
  ANDN U4690 ( .B(B[50]), .A(n39), .Z(n4536) );
  XNOR U4691 ( .A(n4544), .B(n4646), .Z(n4537) );
  XNOR U4692 ( .A(n4543), .B(n4541), .Z(n4646) );
  AND U4693 ( .A(n4647), .B(n4648), .Z(n4541) );
  NANDN U4694 ( .A(n4649), .B(n4650), .Z(n4648) );
  OR U4695 ( .A(n4651), .B(n4652), .Z(n4650) );
  NAND U4696 ( .A(n4652), .B(n4651), .Z(n4647) );
  ANDN U4697 ( .B(B[51]), .A(n40), .Z(n4543) );
  XNOR U4698 ( .A(n4551), .B(n4653), .Z(n4544) );
  XNOR U4699 ( .A(n4550), .B(n4548), .Z(n4653) );
  AND U4700 ( .A(n4654), .B(n4655), .Z(n4548) );
  NANDN U4701 ( .A(n4656), .B(n4657), .Z(n4655) );
  NAND U4702 ( .A(n4658), .B(n4659), .Z(n4657) );
  ANDN U4703 ( .B(B[52]), .A(n41), .Z(n4550) );
  XOR U4704 ( .A(n4557), .B(n4660), .Z(n4551) );
  XNOR U4705 ( .A(n4555), .B(n4558), .Z(n4660) );
  NAND U4706 ( .A(A[2]), .B(B[53]), .Z(n4558) );
  NANDN U4707 ( .A(n4661), .B(n4662), .Z(n4555) );
  AND U4708 ( .A(A[0]), .B(B[54]), .Z(n4662) );
  XNOR U4709 ( .A(n4560), .B(n4663), .Z(n4557) );
  NAND U4710 ( .A(A[0]), .B(B[55]), .Z(n4663) );
  NAND U4711 ( .A(B[54]), .B(A[1]), .Z(n4560) );
  NAND U4712 ( .A(n4664), .B(n4665), .Z(n136) );
  NANDN U4713 ( .A(n4666), .B(n4667), .Z(n4665) );
  OR U4714 ( .A(n4668), .B(n4669), .Z(n4667) );
  NAND U4715 ( .A(n4669), .B(n4668), .Z(n4664) );
  XOR U4716 ( .A(n138), .B(n137), .Z(\A1[52] ) );
  XOR U4717 ( .A(n4669), .B(n4670), .Z(n137) );
  XNOR U4718 ( .A(n4668), .B(n4666), .Z(n4670) );
  AND U4719 ( .A(n4671), .B(n4672), .Z(n4666) );
  NANDN U4720 ( .A(n4673), .B(n4674), .Z(n4672) );
  NANDN U4721 ( .A(n4675), .B(n4676), .Z(n4674) );
  NANDN U4722 ( .A(n4676), .B(n4675), .Z(n4671) );
  ANDN U4723 ( .B(B[39]), .A(n29), .Z(n4668) );
  XNOR U4724 ( .A(n4575), .B(n4677), .Z(n4669) );
  XNOR U4725 ( .A(n4574), .B(n4572), .Z(n4677) );
  AND U4726 ( .A(n4678), .B(n4679), .Z(n4572) );
  NANDN U4727 ( .A(n4680), .B(n4681), .Z(n4679) );
  OR U4728 ( .A(n4682), .B(n4683), .Z(n4681) );
  NAND U4729 ( .A(n4683), .B(n4682), .Z(n4678) );
  ANDN U4730 ( .B(B[40]), .A(n30), .Z(n4574) );
  XNOR U4731 ( .A(n4582), .B(n4684), .Z(n4575) );
  XNOR U4732 ( .A(n4581), .B(n4579), .Z(n4684) );
  AND U4733 ( .A(n4685), .B(n4686), .Z(n4579) );
  NANDN U4734 ( .A(n4687), .B(n4688), .Z(n4686) );
  NANDN U4735 ( .A(n4689), .B(n4690), .Z(n4688) );
  NANDN U4736 ( .A(n4690), .B(n4689), .Z(n4685) );
  ANDN U4737 ( .B(B[41]), .A(n31), .Z(n4581) );
  XNOR U4738 ( .A(n4589), .B(n4691), .Z(n4582) );
  XNOR U4739 ( .A(n4588), .B(n4586), .Z(n4691) );
  AND U4740 ( .A(n4692), .B(n4693), .Z(n4586) );
  NANDN U4741 ( .A(n4694), .B(n4695), .Z(n4693) );
  OR U4742 ( .A(n4696), .B(n4697), .Z(n4695) );
  NAND U4743 ( .A(n4697), .B(n4696), .Z(n4692) );
  ANDN U4744 ( .B(B[42]), .A(n32), .Z(n4588) );
  XNOR U4745 ( .A(n4596), .B(n4698), .Z(n4589) );
  XNOR U4746 ( .A(n4595), .B(n4593), .Z(n4698) );
  AND U4747 ( .A(n4699), .B(n4700), .Z(n4593) );
  NANDN U4748 ( .A(n4701), .B(n4702), .Z(n4700) );
  NANDN U4749 ( .A(n4703), .B(n4704), .Z(n4702) );
  NANDN U4750 ( .A(n4704), .B(n4703), .Z(n4699) );
  ANDN U4751 ( .B(B[43]), .A(n33), .Z(n4595) );
  XNOR U4752 ( .A(n4603), .B(n4705), .Z(n4596) );
  XNOR U4753 ( .A(n4602), .B(n4600), .Z(n4705) );
  AND U4754 ( .A(n4706), .B(n4707), .Z(n4600) );
  NANDN U4755 ( .A(n4708), .B(n4709), .Z(n4707) );
  OR U4756 ( .A(n4710), .B(n4711), .Z(n4709) );
  NAND U4757 ( .A(n4711), .B(n4710), .Z(n4706) );
  ANDN U4758 ( .B(B[44]), .A(n34), .Z(n4602) );
  XNOR U4759 ( .A(n4610), .B(n4712), .Z(n4603) );
  XNOR U4760 ( .A(n4609), .B(n4607), .Z(n4712) );
  AND U4761 ( .A(n4713), .B(n4714), .Z(n4607) );
  NANDN U4762 ( .A(n4715), .B(n4716), .Z(n4714) );
  NANDN U4763 ( .A(n4717), .B(n4718), .Z(n4716) );
  NANDN U4764 ( .A(n4718), .B(n4717), .Z(n4713) );
  ANDN U4765 ( .B(B[45]), .A(n35), .Z(n4609) );
  XNOR U4766 ( .A(n4617), .B(n4719), .Z(n4610) );
  XNOR U4767 ( .A(n4616), .B(n4614), .Z(n4719) );
  AND U4768 ( .A(n4720), .B(n4721), .Z(n4614) );
  NANDN U4769 ( .A(n4722), .B(n4723), .Z(n4721) );
  OR U4770 ( .A(n4724), .B(n4725), .Z(n4723) );
  NAND U4771 ( .A(n4725), .B(n4724), .Z(n4720) );
  ANDN U4772 ( .B(B[46]), .A(n36), .Z(n4616) );
  XNOR U4773 ( .A(n4624), .B(n4726), .Z(n4617) );
  XNOR U4774 ( .A(n4623), .B(n4621), .Z(n4726) );
  AND U4775 ( .A(n4727), .B(n4728), .Z(n4621) );
  NANDN U4776 ( .A(n4729), .B(n4730), .Z(n4728) );
  NANDN U4777 ( .A(n4731), .B(n4732), .Z(n4730) );
  NANDN U4778 ( .A(n4732), .B(n4731), .Z(n4727) );
  ANDN U4779 ( .B(B[47]), .A(n37), .Z(n4623) );
  XNOR U4780 ( .A(n4631), .B(n4733), .Z(n4624) );
  XNOR U4781 ( .A(n4630), .B(n4628), .Z(n4733) );
  AND U4782 ( .A(n4734), .B(n4735), .Z(n4628) );
  NANDN U4783 ( .A(n4736), .B(n4737), .Z(n4735) );
  OR U4784 ( .A(n4738), .B(n4739), .Z(n4737) );
  NAND U4785 ( .A(n4739), .B(n4738), .Z(n4734) );
  ANDN U4786 ( .B(B[48]), .A(n38), .Z(n4630) );
  XNOR U4787 ( .A(n4638), .B(n4740), .Z(n4631) );
  XNOR U4788 ( .A(n4637), .B(n4635), .Z(n4740) );
  AND U4789 ( .A(n4741), .B(n4742), .Z(n4635) );
  NANDN U4790 ( .A(n4743), .B(n4744), .Z(n4742) );
  NANDN U4791 ( .A(n4745), .B(n4746), .Z(n4744) );
  NANDN U4792 ( .A(n4746), .B(n4745), .Z(n4741) );
  ANDN U4793 ( .B(B[49]), .A(n39), .Z(n4637) );
  XNOR U4794 ( .A(n4645), .B(n4747), .Z(n4638) );
  XNOR U4795 ( .A(n4644), .B(n4642), .Z(n4747) );
  AND U4796 ( .A(n4748), .B(n4749), .Z(n4642) );
  NANDN U4797 ( .A(n4750), .B(n4751), .Z(n4749) );
  OR U4798 ( .A(n4752), .B(n4753), .Z(n4751) );
  NAND U4799 ( .A(n4753), .B(n4752), .Z(n4748) );
  ANDN U4800 ( .B(B[50]), .A(n40), .Z(n4644) );
  XNOR U4801 ( .A(n4652), .B(n4754), .Z(n4645) );
  XNOR U4802 ( .A(n4651), .B(n4649), .Z(n4754) );
  AND U4803 ( .A(n4755), .B(n4756), .Z(n4649) );
  NANDN U4804 ( .A(n4757), .B(n4758), .Z(n4756) );
  NAND U4805 ( .A(n4759), .B(n4760), .Z(n4758) );
  ANDN U4806 ( .B(B[51]), .A(n41), .Z(n4651) );
  XOR U4807 ( .A(n4658), .B(n4761), .Z(n4652) );
  XNOR U4808 ( .A(n4656), .B(n4659), .Z(n4761) );
  NAND U4809 ( .A(A[2]), .B(B[52]), .Z(n4659) );
  NANDN U4810 ( .A(n4762), .B(n4763), .Z(n4656) );
  AND U4811 ( .A(A[0]), .B(B[53]), .Z(n4763) );
  XNOR U4812 ( .A(n4661), .B(n4764), .Z(n4658) );
  NAND U4813 ( .A(A[0]), .B(B[54]), .Z(n4764) );
  NAND U4814 ( .A(B[53]), .B(A[1]), .Z(n4661) );
  NAND U4815 ( .A(n4765), .B(n4766), .Z(n138) );
  NANDN U4816 ( .A(n4767), .B(n4768), .Z(n4766) );
  OR U4817 ( .A(n4769), .B(n4770), .Z(n4768) );
  NAND U4818 ( .A(n4770), .B(n4769), .Z(n4765) );
  XOR U4819 ( .A(n140), .B(n139), .Z(\A1[51] ) );
  XOR U4820 ( .A(n4770), .B(n4771), .Z(n139) );
  XNOR U4821 ( .A(n4769), .B(n4767), .Z(n4771) );
  AND U4822 ( .A(n4772), .B(n4773), .Z(n4767) );
  NANDN U4823 ( .A(n4774), .B(n4775), .Z(n4773) );
  NANDN U4824 ( .A(n4776), .B(n4777), .Z(n4775) );
  NANDN U4825 ( .A(n4777), .B(n4776), .Z(n4772) );
  ANDN U4826 ( .B(B[38]), .A(n29), .Z(n4769) );
  XNOR U4827 ( .A(n4676), .B(n4778), .Z(n4770) );
  XNOR U4828 ( .A(n4675), .B(n4673), .Z(n4778) );
  AND U4829 ( .A(n4779), .B(n4780), .Z(n4673) );
  NANDN U4830 ( .A(n4781), .B(n4782), .Z(n4780) );
  OR U4831 ( .A(n4783), .B(n4784), .Z(n4782) );
  NAND U4832 ( .A(n4784), .B(n4783), .Z(n4779) );
  ANDN U4833 ( .B(B[39]), .A(n30), .Z(n4675) );
  XNOR U4834 ( .A(n4683), .B(n4785), .Z(n4676) );
  XNOR U4835 ( .A(n4682), .B(n4680), .Z(n4785) );
  AND U4836 ( .A(n4786), .B(n4787), .Z(n4680) );
  NANDN U4837 ( .A(n4788), .B(n4789), .Z(n4787) );
  NANDN U4838 ( .A(n4790), .B(n4791), .Z(n4789) );
  NANDN U4839 ( .A(n4791), .B(n4790), .Z(n4786) );
  ANDN U4840 ( .B(B[40]), .A(n31), .Z(n4682) );
  XNOR U4841 ( .A(n4690), .B(n4792), .Z(n4683) );
  XNOR U4842 ( .A(n4689), .B(n4687), .Z(n4792) );
  AND U4843 ( .A(n4793), .B(n4794), .Z(n4687) );
  NANDN U4844 ( .A(n4795), .B(n4796), .Z(n4794) );
  OR U4845 ( .A(n4797), .B(n4798), .Z(n4796) );
  NAND U4846 ( .A(n4798), .B(n4797), .Z(n4793) );
  ANDN U4847 ( .B(B[41]), .A(n32), .Z(n4689) );
  XNOR U4848 ( .A(n4697), .B(n4799), .Z(n4690) );
  XNOR U4849 ( .A(n4696), .B(n4694), .Z(n4799) );
  AND U4850 ( .A(n4800), .B(n4801), .Z(n4694) );
  NANDN U4851 ( .A(n4802), .B(n4803), .Z(n4801) );
  NANDN U4852 ( .A(n4804), .B(n4805), .Z(n4803) );
  NANDN U4853 ( .A(n4805), .B(n4804), .Z(n4800) );
  ANDN U4854 ( .B(B[42]), .A(n33), .Z(n4696) );
  XNOR U4855 ( .A(n4704), .B(n4806), .Z(n4697) );
  XNOR U4856 ( .A(n4703), .B(n4701), .Z(n4806) );
  AND U4857 ( .A(n4807), .B(n4808), .Z(n4701) );
  NANDN U4858 ( .A(n4809), .B(n4810), .Z(n4808) );
  OR U4859 ( .A(n4811), .B(n4812), .Z(n4810) );
  NAND U4860 ( .A(n4812), .B(n4811), .Z(n4807) );
  ANDN U4861 ( .B(B[43]), .A(n34), .Z(n4703) );
  XNOR U4862 ( .A(n4711), .B(n4813), .Z(n4704) );
  XNOR U4863 ( .A(n4710), .B(n4708), .Z(n4813) );
  AND U4864 ( .A(n4814), .B(n4815), .Z(n4708) );
  NANDN U4865 ( .A(n4816), .B(n4817), .Z(n4815) );
  NANDN U4866 ( .A(n4818), .B(n4819), .Z(n4817) );
  NANDN U4867 ( .A(n4819), .B(n4818), .Z(n4814) );
  ANDN U4868 ( .B(B[44]), .A(n35), .Z(n4710) );
  XNOR U4869 ( .A(n4718), .B(n4820), .Z(n4711) );
  XNOR U4870 ( .A(n4717), .B(n4715), .Z(n4820) );
  AND U4871 ( .A(n4821), .B(n4822), .Z(n4715) );
  NANDN U4872 ( .A(n4823), .B(n4824), .Z(n4822) );
  OR U4873 ( .A(n4825), .B(n4826), .Z(n4824) );
  NAND U4874 ( .A(n4826), .B(n4825), .Z(n4821) );
  ANDN U4875 ( .B(B[45]), .A(n36), .Z(n4717) );
  XNOR U4876 ( .A(n4725), .B(n4827), .Z(n4718) );
  XNOR U4877 ( .A(n4724), .B(n4722), .Z(n4827) );
  AND U4878 ( .A(n4828), .B(n4829), .Z(n4722) );
  NANDN U4879 ( .A(n4830), .B(n4831), .Z(n4829) );
  NANDN U4880 ( .A(n4832), .B(n4833), .Z(n4831) );
  NANDN U4881 ( .A(n4833), .B(n4832), .Z(n4828) );
  ANDN U4882 ( .B(B[46]), .A(n37), .Z(n4724) );
  XNOR U4883 ( .A(n4732), .B(n4834), .Z(n4725) );
  XNOR U4884 ( .A(n4731), .B(n4729), .Z(n4834) );
  AND U4885 ( .A(n4835), .B(n4836), .Z(n4729) );
  NANDN U4886 ( .A(n4837), .B(n4838), .Z(n4836) );
  OR U4887 ( .A(n4839), .B(n4840), .Z(n4838) );
  NAND U4888 ( .A(n4840), .B(n4839), .Z(n4835) );
  ANDN U4889 ( .B(B[47]), .A(n38), .Z(n4731) );
  XNOR U4890 ( .A(n4739), .B(n4841), .Z(n4732) );
  XNOR U4891 ( .A(n4738), .B(n4736), .Z(n4841) );
  AND U4892 ( .A(n4842), .B(n4843), .Z(n4736) );
  NANDN U4893 ( .A(n4844), .B(n4845), .Z(n4843) );
  NANDN U4894 ( .A(n4846), .B(n4847), .Z(n4845) );
  NANDN U4895 ( .A(n4847), .B(n4846), .Z(n4842) );
  ANDN U4896 ( .B(B[48]), .A(n39), .Z(n4738) );
  XNOR U4897 ( .A(n4746), .B(n4848), .Z(n4739) );
  XNOR U4898 ( .A(n4745), .B(n4743), .Z(n4848) );
  AND U4899 ( .A(n4849), .B(n4850), .Z(n4743) );
  NANDN U4900 ( .A(n4851), .B(n4852), .Z(n4850) );
  OR U4901 ( .A(n4853), .B(n4854), .Z(n4852) );
  NAND U4902 ( .A(n4854), .B(n4853), .Z(n4849) );
  ANDN U4903 ( .B(B[49]), .A(n40), .Z(n4745) );
  XNOR U4904 ( .A(n4753), .B(n4855), .Z(n4746) );
  XNOR U4905 ( .A(n4752), .B(n4750), .Z(n4855) );
  AND U4906 ( .A(n4856), .B(n4857), .Z(n4750) );
  NANDN U4907 ( .A(n4858), .B(n4859), .Z(n4857) );
  NAND U4908 ( .A(n4860), .B(n4861), .Z(n4859) );
  ANDN U4909 ( .B(B[50]), .A(n41), .Z(n4752) );
  XOR U4910 ( .A(n4759), .B(n4862), .Z(n4753) );
  XNOR U4911 ( .A(n4757), .B(n4760), .Z(n4862) );
  NAND U4912 ( .A(A[2]), .B(B[51]), .Z(n4760) );
  NANDN U4913 ( .A(n4863), .B(n4864), .Z(n4757) );
  AND U4914 ( .A(A[0]), .B(B[52]), .Z(n4864) );
  XNOR U4915 ( .A(n4762), .B(n4865), .Z(n4759) );
  NAND U4916 ( .A(A[0]), .B(B[53]), .Z(n4865) );
  NAND U4917 ( .A(B[52]), .B(A[1]), .Z(n4762) );
  NAND U4918 ( .A(n4866), .B(n4867), .Z(n140) );
  NANDN U4919 ( .A(n4868), .B(n4869), .Z(n4867) );
  OR U4920 ( .A(n4870), .B(n4871), .Z(n4869) );
  NAND U4921 ( .A(n4871), .B(n4870), .Z(n4866) );
  XOR U4922 ( .A(n142), .B(n141), .Z(\A1[50] ) );
  XOR U4923 ( .A(n4871), .B(n4872), .Z(n141) );
  XNOR U4924 ( .A(n4870), .B(n4868), .Z(n4872) );
  AND U4925 ( .A(n4873), .B(n4874), .Z(n4868) );
  NANDN U4926 ( .A(n4875), .B(n4876), .Z(n4874) );
  NANDN U4927 ( .A(n4877), .B(n4878), .Z(n4876) );
  NANDN U4928 ( .A(n4878), .B(n4877), .Z(n4873) );
  ANDN U4929 ( .B(B[37]), .A(n29), .Z(n4870) );
  XNOR U4930 ( .A(n4777), .B(n4879), .Z(n4871) );
  XNOR U4931 ( .A(n4776), .B(n4774), .Z(n4879) );
  AND U4932 ( .A(n4880), .B(n4881), .Z(n4774) );
  NANDN U4933 ( .A(n4882), .B(n4883), .Z(n4881) );
  OR U4934 ( .A(n4884), .B(n4885), .Z(n4883) );
  NAND U4935 ( .A(n4885), .B(n4884), .Z(n4880) );
  ANDN U4936 ( .B(B[38]), .A(n30), .Z(n4776) );
  XNOR U4937 ( .A(n4784), .B(n4886), .Z(n4777) );
  XNOR U4938 ( .A(n4783), .B(n4781), .Z(n4886) );
  AND U4939 ( .A(n4887), .B(n4888), .Z(n4781) );
  NANDN U4940 ( .A(n4889), .B(n4890), .Z(n4888) );
  NANDN U4941 ( .A(n4891), .B(n4892), .Z(n4890) );
  NANDN U4942 ( .A(n4892), .B(n4891), .Z(n4887) );
  ANDN U4943 ( .B(B[39]), .A(n31), .Z(n4783) );
  XNOR U4944 ( .A(n4791), .B(n4893), .Z(n4784) );
  XNOR U4945 ( .A(n4790), .B(n4788), .Z(n4893) );
  AND U4946 ( .A(n4894), .B(n4895), .Z(n4788) );
  NANDN U4947 ( .A(n4896), .B(n4897), .Z(n4895) );
  OR U4948 ( .A(n4898), .B(n4899), .Z(n4897) );
  NAND U4949 ( .A(n4899), .B(n4898), .Z(n4894) );
  ANDN U4950 ( .B(B[40]), .A(n32), .Z(n4790) );
  XNOR U4951 ( .A(n4798), .B(n4900), .Z(n4791) );
  XNOR U4952 ( .A(n4797), .B(n4795), .Z(n4900) );
  AND U4953 ( .A(n4901), .B(n4902), .Z(n4795) );
  NANDN U4954 ( .A(n4903), .B(n4904), .Z(n4902) );
  NANDN U4955 ( .A(n4905), .B(n4906), .Z(n4904) );
  NANDN U4956 ( .A(n4906), .B(n4905), .Z(n4901) );
  ANDN U4957 ( .B(B[41]), .A(n33), .Z(n4797) );
  XNOR U4958 ( .A(n4805), .B(n4907), .Z(n4798) );
  XNOR U4959 ( .A(n4804), .B(n4802), .Z(n4907) );
  AND U4960 ( .A(n4908), .B(n4909), .Z(n4802) );
  NANDN U4961 ( .A(n4910), .B(n4911), .Z(n4909) );
  OR U4962 ( .A(n4912), .B(n4913), .Z(n4911) );
  NAND U4963 ( .A(n4913), .B(n4912), .Z(n4908) );
  ANDN U4964 ( .B(B[42]), .A(n34), .Z(n4804) );
  XNOR U4965 ( .A(n4812), .B(n4914), .Z(n4805) );
  XNOR U4966 ( .A(n4811), .B(n4809), .Z(n4914) );
  AND U4967 ( .A(n4915), .B(n4916), .Z(n4809) );
  NANDN U4968 ( .A(n4917), .B(n4918), .Z(n4916) );
  NANDN U4969 ( .A(n4919), .B(n4920), .Z(n4918) );
  NANDN U4970 ( .A(n4920), .B(n4919), .Z(n4915) );
  ANDN U4971 ( .B(B[43]), .A(n35), .Z(n4811) );
  XNOR U4972 ( .A(n4819), .B(n4921), .Z(n4812) );
  XNOR U4973 ( .A(n4818), .B(n4816), .Z(n4921) );
  AND U4974 ( .A(n4922), .B(n4923), .Z(n4816) );
  NANDN U4975 ( .A(n4924), .B(n4925), .Z(n4923) );
  OR U4976 ( .A(n4926), .B(n4927), .Z(n4925) );
  NAND U4977 ( .A(n4927), .B(n4926), .Z(n4922) );
  ANDN U4978 ( .B(B[44]), .A(n36), .Z(n4818) );
  XNOR U4979 ( .A(n4826), .B(n4928), .Z(n4819) );
  XNOR U4980 ( .A(n4825), .B(n4823), .Z(n4928) );
  AND U4981 ( .A(n4929), .B(n4930), .Z(n4823) );
  NANDN U4982 ( .A(n4931), .B(n4932), .Z(n4930) );
  NANDN U4983 ( .A(n4933), .B(n4934), .Z(n4932) );
  NANDN U4984 ( .A(n4934), .B(n4933), .Z(n4929) );
  ANDN U4985 ( .B(B[45]), .A(n37), .Z(n4825) );
  XNOR U4986 ( .A(n4833), .B(n4935), .Z(n4826) );
  XNOR U4987 ( .A(n4832), .B(n4830), .Z(n4935) );
  AND U4988 ( .A(n4936), .B(n4937), .Z(n4830) );
  NANDN U4989 ( .A(n4938), .B(n4939), .Z(n4937) );
  OR U4990 ( .A(n4940), .B(n4941), .Z(n4939) );
  NAND U4991 ( .A(n4941), .B(n4940), .Z(n4936) );
  ANDN U4992 ( .B(B[46]), .A(n38), .Z(n4832) );
  XNOR U4993 ( .A(n4840), .B(n4942), .Z(n4833) );
  XNOR U4994 ( .A(n4839), .B(n4837), .Z(n4942) );
  AND U4995 ( .A(n4943), .B(n4944), .Z(n4837) );
  NANDN U4996 ( .A(n4945), .B(n4946), .Z(n4944) );
  NANDN U4997 ( .A(n4947), .B(n4948), .Z(n4946) );
  NANDN U4998 ( .A(n4948), .B(n4947), .Z(n4943) );
  ANDN U4999 ( .B(B[47]), .A(n39), .Z(n4839) );
  XNOR U5000 ( .A(n4847), .B(n4949), .Z(n4840) );
  XNOR U5001 ( .A(n4846), .B(n4844), .Z(n4949) );
  AND U5002 ( .A(n4950), .B(n4951), .Z(n4844) );
  NANDN U5003 ( .A(n4952), .B(n4953), .Z(n4951) );
  OR U5004 ( .A(n4954), .B(n4955), .Z(n4953) );
  NAND U5005 ( .A(n4955), .B(n4954), .Z(n4950) );
  ANDN U5006 ( .B(B[48]), .A(n40), .Z(n4846) );
  XNOR U5007 ( .A(n4854), .B(n4956), .Z(n4847) );
  XNOR U5008 ( .A(n4853), .B(n4851), .Z(n4956) );
  AND U5009 ( .A(n4957), .B(n4958), .Z(n4851) );
  NANDN U5010 ( .A(n4959), .B(n4960), .Z(n4958) );
  NAND U5011 ( .A(n4961), .B(n4962), .Z(n4960) );
  ANDN U5012 ( .B(B[49]), .A(n41), .Z(n4853) );
  XOR U5013 ( .A(n4860), .B(n4963), .Z(n4854) );
  XNOR U5014 ( .A(n4858), .B(n4861), .Z(n4963) );
  NAND U5015 ( .A(A[2]), .B(B[50]), .Z(n4861) );
  NANDN U5016 ( .A(n4964), .B(n4965), .Z(n4858) );
  AND U5017 ( .A(A[0]), .B(B[51]), .Z(n4965) );
  XNOR U5018 ( .A(n4863), .B(n4966), .Z(n4860) );
  NAND U5019 ( .A(A[0]), .B(B[52]), .Z(n4966) );
  NAND U5020 ( .A(B[51]), .B(A[1]), .Z(n4863) );
  NAND U5021 ( .A(n4967), .B(n4968), .Z(n142) );
  NANDN U5022 ( .A(n4969), .B(n4970), .Z(n4968) );
  OR U5023 ( .A(n4971), .B(n4972), .Z(n4970) );
  NAND U5024 ( .A(n4972), .B(n4971), .Z(n4967) );
  XNOR U5025 ( .A(n4973), .B(n4974), .Z(\A1[4] ) );
  XNOR U5026 ( .A(n4975), .B(n4976), .Z(n4974) );
  XOR U5027 ( .A(n144), .B(n143), .Z(\A1[49] ) );
  XOR U5028 ( .A(n4972), .B(n4977), .Z(n143) );
  XNOR U5029 ( .A(n4971), .B(n4969), .Z(n4977) );
  AND U5030 ( .A(n4978), .B(n4979), .Z(n4969) );
  NANDN U5031 ( .A(n4980), .B(n4981), .Z(n4979) );
  NANDN U5032 ( .A(n4982), .B(n4983), .Z(n4981) );
  NANDN U5033 ( .A(n4983), .B(n4982), .Z(n4978) );
  ANDN U5034 ( .B(B[36]), .A(n29), .Z(n4971) );
  XNOR U5035 ( .A(n4878), .B(n4984), .Z(n4972) );
  XNOR U5036 ( .A(n4877), .B(n4875), .Z(n4984) );
  AND U5037 ( .A(n4985), .B(n4986), .Z(n4875) );
  NANDN U5038 ( .A(n4987), .B(n4988), .Z(n4986) );
  OR U5039 ( .A(n4989), .B(n4990), .Z(n4988) );
  NAND U5040 ( .A(n4990), .B(n4989), .Z(n4985) );
  ANDN U5041 ( .B(B[37]), .A(n30), .Z(n4877) );
  XNOR U5042 ( .A(n4885), .B(n4991), .Z(n4878) );
  XNOR U5043 ( .A(n4884), .B(n4882), .Z(n4991) );
  AND U5044 ( .A(n4992), .B(n4993), .Z(n4882) );
  NANDN U5045 ( .A(n4994), .B(n4995), .Z(n4993) );
  NANDN U5046 ( .A(n4996), .B(n4997), .Z(n4995) );
  NANDN U5047 ( .A(n4997), .B(n4996), .Z(n4992) );
  ANDN U5048 ( .B(B[38]), .A(n31), .Z(n4884) );
  XNOR U5049 ( .A(n4892), .B(n4998), .Z(n4885) );
  XNOR U5050 ( .A(n4891), .B(n4889), .Z(n4998) );
  AND U5051 ( .A(n4999), .B(n5000), .Z(n4889) );
  NANDN U5052 ( .A(n5001), .B(n5002), .Z(n5000) );
  OR U5053 ( .A(n5003), .B(n5004), .Z(n5002) );
  NAND U5054 ( .A(n5004), .B(n5003), .Z(n4999) );
  ANDN U5055 ( .B(B[39]), .A(n32), .Z(n4891) );
  XNOR U5056 ( .A(n4899), .B(n5005), .Z(n4892) );
  XNOR U5057 ( .A(n4898), .B(n4896), .Z(n5005) );
  AND U5058 ( .A(n5006), .B(n5007), .Z(n4896) );
  NANDN U5059 ( .A(n5008), .B(n5009), .Z(n5007) );
  NANDN U5060 ( .A(n5010), .B(n5011), .Z(n5009) );
  NANDN U5061 ( .A(n5011), .B(n5010), .Z(n5006) );
  ANDN U5062 ( .B(B[40]), .A(n33), .Z(n4898) );
  XNOR U5063 ( .A(n4906), .B(n5012), .Z(n4899) );
  XNOR U5064 ( .A(n4905), .B(n4903), .Z(n5012) );
  AND U5065 ( .A(n5013), .B(n5014), .Z(n4903) );
  NANDN U5066 ( .A(n5015), .B(n5016), .Z(n5014) );
  OR U5067 ( .A(n5017), .B(n5018), .Z(n5016) );
  NAND U5068 ( .A(n5018), .B(n5017), .Z(n5013) );
  ANDN U5069 ( .B(B[41]), .A(n34), .Z(n4905) );
  XNOR U5070 ( .A(n4913), .B(n5019), .Z(n4906) );
  XNOR U5071 ( .A(n4912), .B(n4910), .Z(n5019) );
  AND U5072 ( .A(n5020), .B(n5021), .Z(n4910) );
  NANDN U5073 ( .A(n5022), .B(n5023), .Z(n5021) );
  NANDN U5074 ( .A(n5024), .B(n5025), .Z(n5023) );
  NANDN U5075 ( .A(n5025), .B(n5024), .Z(n5020) );
  ANDN U5076 ( .B(B[42]), .A(n35), .Z(n4912) );
  XNOR U5077 ( .A(n4920), .B(n5026), .Z(n4913) );
  XNOR U5078 ( .A(n4919), .B(n4917), .Z(n5026) );
  AND U5079 ( .A(n5027), .B(n5028), .Z(n4917) );
  NANDN U5080 ( .A(n5029), .B(n5030), .Z(n5028) );
  OR U5081 ( .A(n5031), .B(n5032), .Z(n5030) );
  NAND U5082 ( .A(n5032), .B(n5031), .Z(n5027) );
  ANDN U5083 ( .B(B[43]), .A(n36), .Z(n4919) );
  XNOR U5084 ( .A(n4927), .B(n5033), .Z(n4920) );
  XNOR U5085 ( .A(n4926), .B(n4924), .Z(n5033) );
  AND U5086 ( .A(n5034), .B(n5035), .Z(n4924) );
  NANDN U5087 ( .A(n5036), .B(n5037), .Z(n5035) );
  NANDN U5088 ( .A(n5038), .B(n5039), .Z(n5037) );
  NANDN U5089 ( .A(n5039), .B(n5038), .Z(n5034) );
  ANDN U5090 ( .B(B[44]), .A(n37), .Z(n4926) );
  XNOR U5091 ( .A(n4934), .B(n5040), .Z(n4927) );
  XNOR U5092 ( .A(n4933), .B(n4931), .Z(n5040) );
  AND U5093 ( .A(n5041), .B(n5042), .Z(n4931) );
  NANDN U5094 ( .A(n5043), .B(n5044), .Z(n5042) );
  OR U5095 ( .A(n5045), .B(n5046), .Z(n5044) );
  NAND U5096 ( .A(n5046), .B(n5045), .Z(n5041) );
  ANDN U5097 ( .B(B[45]), .A(n38), .Z(n4933) );
  XNOR U5098 ( .A(n4941), .B(n5047), .Z(n4934) );
  XNOR U5099 ( .A(n4940), .B(n4938), .Z(n5047) );
  AND U5100 ( .A(n5048), .B(n5049), .Z(n4938) );
  NANDN U5101 ( .A(n5050), .B(n5051), .Z(n5049) );
  NANDN U5102 ( .A(n5052), .B(n5053), .Z(n5051) );
  NANDN U5103 ( .A(n5053), .B(n5052), .Z(n5048) );
  ANDN U5104 ( .B(B[46]), .A(n39), .Z(n4940) );
  XNOR U5105 ( .A(n4948), .B(n5054), .Z(n4941) );
  XNOR U5106 ( .A(n4947), .B(n4945), .Z(n5054) );
  AND U5107 ( .A(n5055), .B(n5056), .Z(n4945) );
  NANDN U5108 ( .A(n5057), .B(n5058), .Z(n5056) );
  OR U5109 ( .A(n5059), .B(n5060), .Z(n5058) );
  NAND U5110 ( .A(n5060), .B(n5059), .Z(n5055) );
  ANDN U5111 ( .B(B[47]), .A(n40), .Z(n4947) );
  XNOR U5112 ( .A(n4955), .B(n5061), .Z(n4948) );
  XNOR U5113 ( .A(n4954), .B(n4952), .Z(n5061) );
  AND U5114 ( .A(n5062), .B(n5063), .Z(n4952) );
  NANDN U5115 ( .A(n5064), .B(n5065), .Z(n5063) );
  NAND U5116 ( .A(n5066), .B(n5067), .Z(n5065) );
  ANDN U5117 ( .B(B[48]), .A(n41), .Z(n4954) );
  XOR U5118 ( .A(n4961), .B(n5068), .Z(n4955) );
  XNOR U5119 ( .A(n4959), .B(n4962), .Z(n5068) );
  NAND U5120 ( .A(A[2]), .B(B[49]), .Z(n4962) );
  NANDN U5121 ( .A(n5069), .B(n5070), .Z(n4959) );
  AND U5122 ( .A(A[0]), .B(B[50]), .Z(n5070) );
  XNOR U5123 ( .A(n4964), .B(n5071), .Z(n4961) );
  NAND U5124 ( .A(A[0]), .B(B[51]), .Z(n5071) );
  NAND U5125 ( .A(B[50]), .B(A[1]), .Z(n4964) );
  NAND U5126 ( .A(n5072), .B(n5073), .Z(n144) );
  NANDN U5127 ( .A(n5074), .B(n5075), .Z(n5073) );
  OR U5128 ( .A(n5076), .B(n5077), .Z(n5075) );
  NAND U5129 ( .A(n5077), .B(n5076), .Z(n5072) );
  XOR U5130 ( .A(n146), .B(n145), .Z(\A1[48] ) );
  XOR U5131 ( .A(n5077), .B(n5078), .Z(n145) );
  XNOR U5132 ( .A(n5076), .B(n5074), .Z(n5078) );
  AND U5133 ( .A(n5079), .B(n5080), .Z(n5074) );
  NANDN U5134 ( .A(n5081), .B(n5082), .Z(n5080) );
  NANDN U5135 ( .A(n5083), .B(n5084), .Z(n5082) );
  NANDN U5136 ( .A(n5084), .B(n5083), .Z(n5079) );
  ANDN U5137 ( .B(B[35]), .A(n29), .Z(n5076) );
  XNOR U5138 ( .A(n4983), .B(n5085), .Z(n5077) );
  XNOR U5139 ( .A(n4982), .B(n4980), .Z(n5085) );
  AND U5140 ( .A(n5086), .B(n5087), .Z(n4980) );
  NANDN U5141 ( .A(n5088), .B(n5089), .Z(n5087) );
  OR U5142 ( .A(n5090), .B(n5091), .Z(n5089) );
  NAND U5143 ( .A(n5091), .B(n5090), .Z(n5086) );
  ANDN U5144 ( .B(B[36]), .A(n30), .Z(n4982) );
  XNOR U5145 ( .A(n4990), .B(n5092), .Z(n4983) );
  XNOR U5146 ( .A(n4989), .B(n4987), .Z(n5092) );
  AND U5147 ( .A(n5093), .B(n5094), .Z(n4987) );
  NANDN U5148 ( .A(n5095), .B(n5096), .Z(n5094) );
  NANDN U5149 ( .A(n5097), .B(n5098), .Z(n5096) );
  NANDN U5150 ( .A(n5098), .B(n5097), .Z(n5093) );
  ANDN U5151 ( .B(B[37]), .A(n31), .Z(n4989) );
  XNOR U5152 ( .A(n4997), .B(n5099), .Z(n4990) );
  XNOR U5153 ( .A(n4996), .B(n4994), .Z(n5099) );
  AND U5154 ( .A(n5100), .B(n5101), .Z(n4994) );
  NANDN U5155 ( .A(n5102), .B(n5103), .Z(n5101) );
  OR U5156 ( .A(n5104), .B(n5105), .Z(n5103) );
  NAND U5157 ( .A(n5105), .B(n5104), .Z(n5100) );
  ANDN U5158 ( .B(B[38]), .A(n32), .Z(n4996) );
  XNOR U5159 ( .A(n5004), .B(n5106), .Z(n4997) );
  XNOR U5160 ( .A(n5003), .B(n5001), .Z(n5106) );
  AND U5161 ( .A(n5107), .B(n5108), .Z(n5001) );
  NANDN U5162 ( .A(n5109), .B(n5110), .Z(n5108) );
  NANDN U5163 ( .A(n5111), .B(n5112), .Z(n5110) );
  NANDN U5164 ( .A(n5112), .B(n5111), .Z(n5107) );
  ANDN U5165 ( .B(B[39]), .A(n33), .Z(n5003) );
  XNOR U5166 ( .A(n5011), .B(n5113), .Z(n5004) );
  XNOR U5167 ( .A(n5010), .B(n5008), .Z(n5113) );
  AND U5168 ( .A(n5114), .B(n5115), .Z(n5008) );
  NANDN U5169 ( .A(n5116), .B(n5117), .Z(n5115) );
  OR U5170 ( .A(n5118), .B(n5119), .Z(n5117) );
  NAND U5171 ( .A(n5119), .B(n5118), .Z(n5114) );
  ANDN U5172 ( .B(B[40]), .A(n34), .Z(n5010) );
  XNOR U5173 ( .A(n5018), .B(n5120), .Z(n5011) );
  XNOR U5174 ( .A(n5017), .B(n5015), .Z(n5120) );
  AND U5175 ( .A(n5121), .B(n5122), .Z(n5015) );
  NANDN U5176 ( .A(n5123), .B(n5124), .Z(n5122) );
  NANDN U5177 ( .A(n5125), .B(n5126), .Z(n5124) );
  NANDN U5178 ( .A(n5126), .B(n5125), .Z(n5121) );
  ANDN U5179 ( .B(B[41]), .A(n35), .Z(n5017) );
  XNOR U5180 ( .A(n5025), .B(n5127), .Z(n5018) );
  XNOR U5181 ( .A(n5024), .B(n5022), .Z(n5127) );
  AND U5182 ( .A(n5128), .B(n5129), .Z(n5022) );
  NANDN U5183 ( .A(n5130), .B(n5131), .Z(n5129) );
  OR U5184 ( .A(n5132), .B(n5133), .Z(n5131) );
  NAND U5185 ( .A(n5133), .B(n5132), .Z(n5128) );
  ANDN U5186 ( .B(B[42]), .A(n36), .Z(n5024) );
  XNOR U5187 ( .A(n5032), .B(n5134), .Z(n5025) );
  XNOR U5188 ( .A(n5031), .B(n5029), .Z(n5134) );
  AND U5189 ( .A(n5135), .B(n5136), .Z(n5029) );
  NANDN U5190 ( .A(n5137), .B(n5138), .Z(n5136) );
  NANDN U5191 ( .A(n5139), .B(n5140), .Z(n5138) );
  NANDN U5192 ( .A(n5140), .B(n5139), .Z(n5135) );
  ANDN U5193 ( .B(B[43]), .A(n37), .Z(n5031) );
  XNOR U5194 ( .A(n5039), .B(n5141), .Z(n5032) );
  XNOR U5195 ( .A(n5038), .B(n5036), .Z(n5141) );
  AND U5196 ( .A(n5142), .B(n5143), .Z(n5036) );
  NANDN U5197 ( .A(n5144), .B(n5145), .Z(n5143) );
  OR U5198 ( .A(n5146), .B(n5147), .Z(n5145) );
  NAND U5199 ( .A(n5147), .B(n5146), .Z(n5142) );
  ANDN U5200 ( .B(B[44]), .A(n38), .Z(n5038) );
  XNOR U5201 ( .A(n5046), .B(n5148), .Z(n5039) );
  XNOR U5202 ( .A(n5045), .B(n5043), .Z(n5148) );
  AND U5203 ( .A(n5149), .B(n5150), .Z(n5043) );
  NANDN U5204 ( .A(n5151), .B(n5152), .Z(n5150) );
  NANDN U5205 ( .A(n5153), .B(n5154), .Z(n5152) );
  NANDN U5206 ( .A(n5154), .B(n5153), .Z(n5149) );
  ANDN U5207 ( .B(B[45]), .A(n39), .Z(n5045) );
  XNOR U5208 ( .A(n5053), .B(n5155), .Z(n5046) );
  XNOR U5209 ( .A(n5052), .B(n5050), .Z(n5155) );
  AND U5210 ( .A(n5156), .B(n5157), .Z(n5050) );
  NANDN U5211 ( .A(n5158), .B(n5159), .Z(n5157) );
  OR U5212 ( .A(n5160), .B(n5161), .Z(n5159) );
  NAND U5213 ( .A(n5161), .B(n5160), .Z(n5156) );
  ANDN U5214 ( .B(B[46]), .A(n40), .Z(n5052) );
  XNOR U5215 ( .A(n5060), .B(n5162), .Z(n5053) );
  XNOR U5216 ( .A(n5059), .B(n5057), .Z(n5162) );
  AND U5217 ( .A(n5163), .B(n5164), .Z(n5057) );
  NANDN U5218 ( .A(n5165), .B(n5166), .Z(n5164) );
  NAND U5219 ( .A(n5167), .B(n5168), .Z(n5166) );
  ANDN U5220 ( .B(B[47]), .A(n41), .Z(n5059) );
  XOR U5221 ( .A(n5066), .B(n5169), .Z(n5060) );
  XNOR U5222 ( .A(n5064), .B(n5067), .Z(n5169) );
  NAND U5223 ( .A(A[2]), .B(B[48]), .Z(n5067) );
  NANDN U5224 ( .A(n5170), .B(n5171), .Z(n5064) );
  AND U5225 ( .A(A[0]), .B(B[49]), .Z(n5171) );
  XNOR U5226 ( .A(n5069), .B(n5172), .Z(n5066) );
  NAND U5227 ( .A(A[0]), .B(B[50]), .Z(n5172) );
  NAND U5228 ( .A(B[49]), .B(A[1]), .Z(n5069) );
  NAND U5229 ( .A(n5173), .B(n5174), .Z(n146) );
  NANDN U5230 ( .A(n5175), .B(n5176), .Z(n5174) );
  OR U5231 ( .A(n5177), .B(n5178), .Z(n5176) );
  NAND U5232 ( .A(n5178), .B(n5177), .Z(n5173) );
  XOR U5233 ( .A(n148), .B(n147), .Z(\A1[47] ) );
  XOR U5234 ( .A(n5178), .B(n5179), .Z(n147) );
  XNOR U5235 ( .A(n5177), .B(n5175), .Z(n5179) );
  AND U5236 ( .A(n5180), .B(n5181), .Z(n5175) );
  NANDN U5237 ( .A(n5182), .B(n5183), .Z(n5181) );
  NANDN U5238 ( .A(n5184), .B(n5185), .Z(n5183) );
  NANDN U5239 ( .A(n5185), .B(n5184), .Z(n5180) );
  ANDN U5240 ( .B(B[34]), .A(n29), .Z(n5177) );
  XNOR U5241 ( .A(n5084), .B(n5186), .Z(n5178) );
  XNOR U5242 ( .A(n5083), .B(n5081), .Z(n5186) );
  AND U5243 ( .A(n5187), .B(n5188), .Z(n5081) );
  NANDN U5244 ( .A(n5189), .B(n5190), .Z(n5188) );
  OR U5245 ( .A(n5191), .B(n5192), .Z(n5190) );
  NAND U5246 ( .A(n5192), .B(n5191), .Z(n5187) );
  ANDN U5247 ( .B(B[35]), .A(n30), .Z(n5083) );
  XNOR U5248 ( .A(n5091), .B(n5193), .Z(n5084) );
  XNOR U5249 ( .A(n5090), .B(n5088), .Z(n5193) );
  AND U5250 ( .A(n5194), .B(n5195), .Z(n5088) );
  NANDN U5251 ( .A(n5196), .B(n5197), .Z(n5195) );
  NANDN U5252 ( .A(n5198), .B(n5199), .Z(n5197) );
  NANDN U5253 ( .A(n5199), .B(n5198), .Z(n5194) );
  ANDN U5254 ( .B(B[36]), .A(n31), .Z(n5090) );
  XNOR U5255 ( .A(n5098), .B(n5200), .Z(n5091) );
  XNOR U5256 ( .A(n5097), .B(n5095), .Z(n5200) );
  AND U5257 ( .A(n5201), .B(n5202), .Z(n5095) );
  NANDN U5258 ( .A(n5203), .B(n5204), .Z(n5202) );
  OR U5259 ( .A(n5205), .B(n5206), .Z(n5204) );
  NAND U5260 ( .A(n5206), .B(n5205), .Z(n5201) );
  ANDN U5261 ( .B(B[37]), .A(n32), .Z(n5097) );
  XNOR U5262 ( .A(n5105), .B(n5207), .Z(n5098) );
  XNOR U5263 ( .A(n5104), .B(n5102), .Z(n5207) );
  AND U5264 ( .A(n5208), .B(n5209), .Z(n5102) );
  NANDN U5265 ( .A(n5210), .B(n5211), .Z(n5209) );
  NANDN U5266 ( .A(n5212), .B(n5213), .Z(n5211) );
  NANDN U5267 ( .A(n5213), .B(n5212), .Z(n5208) );
  ANDN U5268 ( .B(B[38]), .A(n33), .Z(n5104) );
  XNOR U5269 ( .A(n5112), .B(n5214), .Z(n5105) );
  XNOR U5270 ( .A(n5111), .B(n5109), .Z(n5214) );
  AND U5271 ( .A(n5215), .B(n5216), .Z(n5109) );
  NANDN U5272 ( .A(n5217), .B(n5218), .Z(n5216) );
  OR U5273 ( .A(n5219), .B(n5220), .Z(n5218) );
  NAND U5274 ( .A(n5220), .B(n5219), .Z(n5215) );
  ANDN U5275 ( .B(B[39]), .A(n34), .Z(n5111) );
  XNOR U5276 ( .A(n5119), .B(n5221), .Z(n5112) );
  XNOR U5277 ( .A(n5118), .B(n5116), .Z(n5221) );
  AND U5278 ( .A(n5222), .B(n5223), .Z(n5116) );
  NANDN U5279 ( .A(n5224), .B(n5225), .Z(n5223) );
  NANDN U5280 ( .A(n5226), .B(n5227), .Z(n5225) );
  NANDN U5281 ( .A(n5227), .B(n5226), .Z(n5222) );
  ANDN U5282 ( .B(B[40]), .A(n35), .Z(n5118) );
  XNOR U5283 ( .A(n5126), .B(n5228), .Z(n5119) );
  XNOR U5284 ( .A(n5125), .B(n5123), .Z(n5228) );
  AND U5285 ( .A(n5229), .B(n5230), .Z(n5123) );
  NANDN U5286 ( .A(n5231), .B(n5232), .Z(n5230) );
  OR U5287 ( .A(n5233), .B(n5234), .Z(n5232) );
  NAND U5288 ( .A(n5234), .B(n5233), .Z(n5229) );
  ANDN U5289 ( .B(B[41]), .A(n36), .Z(n5125) );
  XNOR U5290 ( .A(n5133), .B(n5235), .Z(n5126) );
  XNOR U5291 ( .A(n5132), .B(n5130), .Z(n5235) );
  AND U5292 ( .A(n5236), .B(n5237), .Z(n5130) );
  NANDN U5293 ( .A(n5238), .B(n5239), .Z(n5237) );
  NANDN U5294 ( .A(n5240), .B(n5241), .Z(n5239) );
  NANDN U5295 ( .A(n5241), .B(n5240), .Z(n5236) );
  ANDN U5296 ( .B(B[42]), .A(n37), .Z(n5132) );
  XNOR U5297 ( .A(n5140), .B(n5242), .Z(n5133) );
  XNOR U5298 ( .A(n5139), .B(n5137), .Z(n5242) );
  AND U5299 ( .A(n5243), .B(n5244), .Z(n5137) );
  NANDN U5300 ( .A(n5245), .B(n5246), .Z(n5244) );
  OR U5301 ( .A(n5247), .B(n5248), .Z(n5246) );
  NAND U5302 ( .A(n5248), .B(n5247), .Z(n5243) );
  ANDN U5303 ( .B(B[43]), .A(n38), .Z(n5139) );
  XNOR U5304 ( .A(n5147), .B(n5249), .Z(n5140) );
  XNOR U5305 ( .A(n5146), .B(n5144), .Z(n5249) );
  AND U5306 ( .A(n5250), .B(n5251), .Z(n5144) );
  NANDN U5307 ( .A(n5252), .B(n5253), .Z(n5251) );
  NANDN U5308 ( .A(n5254), .B(n5255), .Z(n5253) );
  NANDN U5309 ( .A(n5255), .B(n5254), .Z(n5250) );
  ANDN U5310 ( .B(B[44]), .A(n39), .Z(n5146) );
  XNOR U5311 ( .A(n5154), .B(n5256), .Z(n5147) );
  XNOR U5312 ( .A(n5153), .B(n5151), .Z(n5256) );
  AND U5313 ( .A(n5257), .B(n5258), .Z(n5151) );
  NANDN U5314 ( .A(n5259), .B(n5260), .Z(n5258) );
  OR U5315 ( .A(n5261), .B(n5262), .Z(n5260) );
  NAND U5316 ( .A(n5262), .B(n5261), .Z(n5257) );
  ANDN U5317 ( .B(B[45]), .A(n40), .Z(n5153) );
  XNOR U5318 ( .A(n5161), .B(n5263), .Z(n5154) );
  XNOR U5319 ( .A(n5160), .B(n5158), .Z(n5263) );
  AND U5320 ( .A(n5264), .B(n5265), .Z(n5158) );
  NANDN U5321 ( .A(n5266), .B(n5267), .Z(n5265) );
  NAND U5322 ( .A(n5268), .B(n5269), .Z(n5267) );
  ANDN U5323 ( .B(B[46]), .A(n41), .Z(n5160) );
  XOR U5324 ( .A(n5167), .B(n5270), .Z(n5161) );
  XNOR U5325 ( .A(n5165), .B(n5168), .Z(n5270) );
  NAND U5326 ( .A(A[2]), .B(B[47]), .Z(n5168) );
  NANDN U5327 ( .A(n5271), .B(n5272), .Z(n5165) );
  AND U5328 ( .A(A[0]), .B(B[48]), .Z(n5272) );
  XNOR U5329 ( .A(n5170), .B(n5273), .Z(n5167) );
  NAND U5330 ( .A(A[0]), .B(B[49]), .Z(n5273) );
  NAND U5331 ( .A(B[48]), .B(A[1]), .Z(n5170) );
  NAND U5332 ( .A(n5274), .B(n5275), .Z(n148) );
  NANDN U5333 ( .A(n5276), .B(n5277), .Z(n5275) );
  OR U5334 ( .A(n5278), .B(n5279), .Z(n5277) );
  NAND U5335 ( .A(n5279), .B(n5278), .Z(n5274) );
  XOR U5336 ( .A(n150), .B(n149), .Z(\A1[46] ) );
  XOR U5337 ( .A(n5279), .B(n5280), .Z(n149) );
  XNOR U5338 ( .A(n5278), .B(n5276), .Z(n5280) );
  AND U5339 ( .A(n5281), .B(n5282), .Z(n5276) );
  NANDN U5340 ( .A(n5283), .B(n5284), .Z(n5282) );
  NANDN U5341 ( .A(n5285), .B(n5286), .Z(n5284) );
  NANDN U5342 ( .A(n5286), .B(n5285), .Z(n5281) );
  ANDN U5343 ( .B(B[33]), .A(n29), .Z(n5278) );
  XNOR U5344 ( .A(n5185), .B(n5287), .Z(n5279) );
  XNOR U5345 ( .A(n5184), .B(n5182), .Z(n5287) );
  AND U5346 ( .A(n5288), .B(n5289), .Z(n5182) );
  NANDN U5347 ( .A(n5290), .B(n5291), .Z(n5289) );
  OR U5348 ( .A(n5292), .B(n5293), .Z(n5291) );
  NAND U5349 ( .A(n5293), .B(n5292), .Z(n5288) );
  ANDN U5350 ( .B(B[34]), .A(n30), .Z(n5184) );
  XNOR U5351 ( .A(n5192), .B(n5294), .Z(n5185) );
  XNOR U5352 ( .A(n5191), .B(n5189), .Z(n5294) );
  AND U5353 ( .A(n5295), .B(n5296), .Z(n5189) );
  NANDN U5354 ( .A(n5297), .B(n5298), .Z(n5296) );
  NANDN U5355 ( .A(n5299), .B(n5300), .Z(n5298) );
  NANDN U5356 ( .A(n5300), .B(n5299), .Z(n5295) );
  ANDN U5357 ( .B(B[35]), .A(n31), .Z(n5191) );
  XNOR U5358 ( .A(n5199), .B(n5301), .Z(n5192) );
  XNOR U5359 ( .A(n5198), .B(n5196), .Z(n5301) );
  AND U5360 ( .A(n5302), .B(n5303), .Z(n5196) );
  NANDN U5361 ( .A(n5304), .B(n5305), .Z(n5303) );
  OR U5362 ( .A(n5306), .B(n5307), .Z(n5305) );
  NAND U5363 ( .A(n5307), .B(n5306), .Z(n5302) );
  ANDN U5364 ( .B(B[36]), .A(n32), .Z(n5198) );
  XNOR U5365 ( .A(n5206), .B(n5308), .Z(n5199) );
  XNOR U5366 ( .A(n5205), .B(n5203), .Z(n5308) );
  AND U5367 ( .A(n5309), .B(n5310), .Z(n5203) );
  NANDN U5368 ( .A(n5311), .B(n5312), .Z(n5310) );
  NANDN U5369 ( .A(n5313), .B(n5314), .Z(n5312) );
  NANDN U5370 ( .A(n5314), .B(n5313), .Z(n5309) );
  ANDN U5371 ( .B(B[37]), .A(n33), .Z(n5205) );
  XNOR U5372 ( .A(n5213), .B(n5315), .Z(n5206) );
  XNOR U5373 ( .A(n5212), .B(n5210), .Z(n5315) );
  AND U5374 ( .A(n5316), .B(n5317), .Z(n5210) );
  NANDN U5375 ( .A(n5318), .B(n5319), .Z(n5317) );
  OR U5376 ( .A(n5320), .B(n5321), .Z(n5319) );
  NAND U5377 ( .A(n5321), .B(n5320), .Z(n5316) );
  ANDN U5378 ( .B(B[38]), .A(n34), .Z(n5212) );
  XNOR U5379 ( .A(n5220), .B(n5322), .Z(n5213) );
  XNOR U5380 ( .A(n5219), .B(n5217), .Z(n5322) );
  AND U5381 ( .A(n5323), .B(n5324), .Z(n5217) );
  NANDN U5382 ( .A(n5325), .B(n5326), .Z(n5324) );
  NANDN U5383 ( .A(n5327), .B(n5328), .Z(n5326) );
  NANDN U5384 ( .A(n5328), .B(n5327), .Z(n5323) );
  ANDN U5385 ( .B(B[39]), .A(n35), .Z(n5219) );
  XNOR U5386 ( .A(n5227), .B(n5329), .Z(n5220) );
  XNOR U5387 ( .A(n5226), .B(n5224), .Z(n5329) );
  AND U5388 ( .A(n5330), .B(n5331), .Z(n5224) );
  NANDN U5389 ( .A(n5332), .B(n5333), .Z(n5331) );
  OR U5390 ( .A(n5334), .B(n5335), .Z(n5333) );
  NAND U5391 ( .A(n5335), .B(n5334), .Z(n5330) );
  ANDN U5392 ( .B(B[40]), .A(n36), .Z(n5226) );
  XNOR U5393 ( .A(n5234), .B(n5336), .Z(n5227) );
  XNOR U5394 ( .A(n5233), .B(n5231), .Z(n5336) );
  AND U5395 ( .A(n5337), .B(n5338), .Z(n5231) );
  NANDN U5396 ( .A(n5339), .B(n5340), .Z(n5338) );
  NANDN U5397 ( .A(n5341), .B(n5342), .Z(n5340) );
  NANDN U5398 ( .A(n5342), .B(n5341), .Z(n5337) );
  ANDN U5399 ( .B(B[41]), .A(n37), .Z(n5233) );
  XNOR U5400 ( .A(n5241), .B(n5343), .Z(n5234) );
  XNOR U5401 ( .A(n5240), .B(n5238), .Z(n5343) );
  AND U5402 ( .A(n5344), .B(n5345), .Z(n5238) );
  NANDN U5403 ( .A(n5346), .B(n5347), .Z(n5345) );
  OR U5404 ( .A(n5348), .B(n5349), .Z(n5347) );
  NAND U5405 ( .A(n5349), .B(n5348), .Z(n5344) );
  ANDN U5406 ( .B(B[42]), .A(n38), .Z(n5240) );
  XNOR U5407 ( .A(n5248), .B(n5350), .Z(n5241) );
  XNOR U5408 ( .A(n5247), .B(n5245), .Z(n5350) );
  AND U5409 ( .A(n5351), .B(n5352), .Z(n5245) );
  NANDN U5410 ( .A(n5353), .B(n5354), .Z(n5352) );
  NANDN U5411 ( .A(n5355), .B(n5356), .Z(n5354) );
  NANDN U5412 ( .A(n5356), .B(n5355), .Z(n5351) );
  ANDN U5413 ( .B(B[43]), .A(n39), .Z(n5247) );
  XNOR U5414 ( .A(n5255), .B(n5357), .Z(n5248) );
  XNOR U5415 ( .A(n5254), .B(n5252), .Z(n5357) );
  AND U5416 ( .A(n5358), .B(n5359), .Z(n5252) );
  NANDN U5417 ( .A(n5360), .B(n5361), .Z(n5359) );
  OR U5418 ( .A(n5362), .B(n5363), .Z(n5361) );
  NAND U5419 ( .A(n5363), .B(n5362), .Z(n5358) );
  ANDN U5420 ( .B(B[44]), .A(n40), .Z(n5254) );
  XNOR U5421 ( .A(n5262), .B(n5364), .Z(n5255) );
  XNOR U5422 ( .A(n5261), .B(n5259), .Z(n5364) );
  AND U5423 ( .A(n5365), .B(n5366), .Z(n5259) );
  NANDN U5424 ( .A(n5367), .B(n5368), .Z(n5366) );
  NAND U5425 ( .A(n5369), .B(n5370), .Z(n5368) );
  ANDN U5426 ( .B(B[45]), .A(n41), .Z(n5261) );
  XOR U5427 ( .A(n5268), .B(n5371), .Z(n5262) );
  XNOR U5428 ( .A(n5266), .B(n5269), .Z(n5371) );
  NAND U5429 ( .A(A[2]), .B(B[46]), .Z(n5269) );
  NANDN U5430 ( .A(n5372), .B(n5373), .Z(n5266) );
  AND U5431 ( .A(A[0]), .B(B[47]), .Z(n5373) );
  XNOR U5432 ( .A(n5271), .B(n5374), .Z(n5268) );
  NAND U5433 ( .A(A[0]), .B(B[48]), .Z(n5374) );
  NAND U5434 ( .A(B[47]), .B(A[1]), .Z(n5271) );
  NAND U5435 ( .A(n5375), .B(n5376), .Z(n150) );
  NANDN U5436 ( .A(n5377), .B(n5378), .Z(n5376) );
  OR U5437 ( .A(n5379), .B(n5380), .Z(n5378) );
  NAND U5438 ( .A(n5380), .B(n5379), .Z(n5375) );
  XOR U5439 ( .A(n152), .B(n151), .Z(\A1[45] ) );
  XOR U5440 ( .A(n5380), .B(n5381), .Z(n151) );
  XNOR U5441 ( .A(n5379), .B(n5377), .Z(n5381) );
  AND U5442 ( .A(n5382), .B(n5383), .Z(n5377) );
  NANDN U5443 ( .A(n5384), .B(n5385), .Z(n5383) );
  NANDN U5444 ( .A(n5386), .B(n5387), .Z(n5385) );
  NANDN U5445 ( .A(n5387), .B(n5386), .Z(n5382) );
  ANDN U5446 ( .B(B[32]), .A(n29), .Z(n5379) );
  XNOR U5447 ( .A(n5286), .B(n5388), .Z(n5380) );
  XNOR U5448 ( .A(n5285), .B(n5283), .Z(n5388) );
  AND U5449 ( .A(n5389), .B(n5390), .Z(n5283) );
  NANDN U5450 ( .A(n5391), .B(n5392), .Z(n5390) );
  OR U5451 ( .A(n5393), .B(n5394), .Z(n5392) );
  NAND U5452 ( .A(n5394), .B(n5393), .Z(n5389) );
  ANDN U5453 ( .B(B[33]), .A(n30), .Z(n5285) );
  XNOR U5454 ( .A(n5293), .B(n5395), .Z(n5286) );
  XNOR U5455 ( .A(n5292), .B(n5290), .Z(n5395) );
  AND U5456 ( .A(n5396), .B(n5397), .Z(n5290) );
  NANDN U5457 ( .A(n5398), .B(n5399), .Z(n5397) );
  NANDN U5458 ( .A(n5400), .B(n5401), .Z(n5399) );
  NANDN U5459 ( .A(n5401), .B(n5400), .Z(n5396) );
  ANDN U5460 ( .B(B[34]), .A(n31), .Z(n5292) );
  XNOR U5461 ( .A(n5300), .B(n5402), .Z(n5293) );
  XNOR U5462 ( .A(n5299), .B(n5297), .Z(n5402) );
  AND U5463 ( .A(n5403), .B(n5404), .Z(n5297) );
  NANDN U5464 ( .A(n5405), .B(n5406), .Z(n5404) );
  OR U5465 ( .A(n5407), .B(n5408), .Z(n5406) );
  NAND U5466 ( .A(n5408), .B(n5407), .Z(n5403) );
  ANDN U5467 ( .B(B[35]), .A(n32), .Z(n5299) );
  XNOR U5468 ( .A(n5307), .B(n5409), .Z(n5300) );
  XNOR U5469 ( .A(n5306), .B(n5304), .Z(n5409) );
  AND U5470 ( .A(n5410), .B(n5411), .Z(n5304) );
  NANDN U5471 ( .A(n5412), .B(n5413), .Z(n5411) );
  NANDN U5472 ( .A(n5414), .B(n5415), .Z(n5413) );
  NANDN U5473 ( .A(n5415), .B(n5414), .Z(n5410) );
  ANDN U5474 ( .B(B[36]), .A(n33), .Z(n5306) );
  XNOR U5475 ( .A(n5314), .B(n5416), .Z(n5307) );
  XNOR U5476 ( .A(n5313), .B(n5311), .Z(n5416) );
  AND U5477 ( .A(n5417), .B(n5418), .Z(n5311) );
  NANDN U5478 ( .A(n5419), .B(n5420), .Z(n5418) );
  OR U5479 ( .A(n5421), .B(n5422), .Z(n5420) );
  NAND U5480 ( .A(n5422), .B(n5421), .Z(n5417) );
  ANDN U5481 ( .B(B[37]), .A(n34), .Z(n5313) );
  XNOR U5482 ( .A(n5321), .B(n5423), .Z(n5314) );
  XNOR U5483 ( .A(n5320), .B(n5318), .Z(n5423) );
  AND U5484 ( .A(n5424), .B(n5425), .Z(n5318) );
  NANDN U5485 ( .A(n5426), .B(n5427), .Z(n5425) );
  NANDN U5486 ( .A(n5428), .B(n5429), .Z(n5427) );
  NANDN U5487 ( .A(n5429), .B(n5428), .Z(n5424) );
  ANDN U5488 ( .B(B[38]), .A(n35), .Z(n5320) );
  XNOR U5489 ( .A(n5328), .B(n5430), .Z(n5321) );
  XNOR U5490 ( .A(n5327), .B(n5325), .Z(n5430) );
  AND U5491 ( .A(n5431), .B(n5432), .Z(n5325) );
  NANDN U5492 ( .A(n5433), .B(n5434), .Z(n5432) );
  OR U5493 ( .A(n5435), .B(n5436), .Z(n5434) );
  NAND U5494 ( .A(n5436), .B(n5435), .Z(n5431) );
  ANDN U5495 ( .B(B[39]), .A(n36), .Z(n5327) );
  XNOR U5496 ( .A(n5335), .B(n5437), .Z(n5328) );
  XNOR U5497 ( .A(n5334), .B(n5332), .Z(n5437) );
  AND U5498 ( .A(n5438), .B(n5439), .Z(n5332) );
  NANDN U5499 ( .A(n5440), .B(n5441), .Z(n5439) );
  NANDN U5500 ( .A(n5442), .B(n5443), .Z(n5441) );
  NANDN U5501 ( .A(n5443), .B(n5442), .Z(n5438) );
  ANDN U5502 ( .B(B[40]), .A(n37), .Z(n5334) );
  XNOR U5503 ( .A(n5342), .B(n5444), .Z(n5335) );
  XNOR U5504 ( .A(n5341), .B(n5339), .Z(n5444) );
  AND U5505 ( .A(n5445), .B(n5446), .Z(n5339) );
  NANDN U5506 ( .A(n5447), .B(n5448), .Z(n5446) );
  OR U5507 ( .A(n5449), .B(n5450), .Z(n5448) );
  NAND U5508 ( .A(n5450), .B(n5449), .Z(n5445) );
  ANDN U5509 ( .B(B[41]), .A(n38), .Z(n5341) );
  XNOR U5510 ( .A(n5349), .B(n5451), .Z(n5342) );
  XNOR U5511 ( .A(n5348), .B(n5346), .Z(n5451) );
  AND U5512 ( .A(n5452), .B(n5453), .Z(n5346) );
  NANDN U5513 ( .A(n5454), .B(n5455), .Z(n5453) );
  NANDN U5514 ( .A(n5456), .B(n5457), .Z(n5455) );
  NANDN U5515 ( .A(n5457), .B(n5456), .Z(n5452) );
  ANDN U5516 ( .B(B[42]), .A(n39), .Z(n5348) );
  XNOR U5517 ( .A(n5356), .B(n5458), .Z(n5349) );
  XNOR U5518 ( .A(n5355), .B(n5353), .Z(n5458) );
  AND U5519 ( .A(n5459), .B(n5460), .Z(n5353) );
  NANDN U5520 ( .A(n5461), .B(n5462), .Z(n5460) );
  OR U5521 ( .A(n5463), .B(n5464), .Z(n5462) );
  NAND U5522 ( .A(n5464), .B(n5463), .Z(n5459) );
  ANDN U5523 ( .B(B[43]), .A(n40), .Z(n5355) );
  XNOR U5524 ( .A(n5363), .B(n5465), .Z(n5356) );
  XNOR U5525 ( .A(n5362), .B(n5360), .Z(n5465) );
  AND U5526 ( .A(n5466), .B(n5467), .Z(n5360) );
  NANDN U5527 ( .A(n5468), .B(n5469), .Z(n5467) );
  NAND U5528 ( .A(n5470), .B(n5471), .Z(n5469) );
  ANDN U5529 ( .B(B[44]), .A(n41), .Z(n5362) );
  XOR U5530 ( .A(n5369), .B(n5472), .Z(n5363) );
  XNOR U5531 ( .A(n5367), .B(n5370), .Z(n5472) );
  NAND U5532 ( .A(A[2]), .B(B[45]), .Z(n5370) );
  NANDN U5533 ( .A(n5473), .B(n5474), .Z(n5367) );
  AND U5534 ( .A(A[0]), .B(B[46]), .Z(n5474) );
  XNOR U5535 ( .A(n5372), .B(n5475), .Z(n5369) );
  NAND U5536 ( .A(A[0]), .B(B[47]), .Z(n5475) );
  NAND U5537 ( .A(B[46]), .B(A[1]), .Z(n5372) );
  NAND U5538 ( .A(n5476), .B(n5477), .Z(n152) );
  NANDN U5539 ( .A(n5478), .B(n5479), .Z(n5477) );
  OR U5540 ( .A(n5480), .B(n5481), .Z(n5479) );
  NAND U5541 ( .A(n5481), .B(n5480), .Z(n5476) );
  XOR U5542 ( .A(n154), .B(n153), .Z(\A1[44] ) );
  XOR U5543 ( .A(n5481), .B(n5482), .Z(n153) );
  XNOR U5544 ( .A(n5480), .B(n5478), .Z(n5482) );
  AND U5545 ( .A(n5483), .B(n5484), .Z(n5478) );
  NANDN U5546 ( .A(n5485), .B(n5486), .Z(n5484) );
  NANDN U5547 ( .A(n5487), .B(n5488), .Z(n5486) );
  NANDN U5548 ( .A(n5488), .B(n5487), .Z(n5483) );
  ANDN U5549 ( .B(B[31]), .A(n29), .Z(n5480) );
  XNOR U5550 ( .A(n5387), .B(n5489), .Z(n5481) );
  XNOR U5551 ( .A(n5386), .B(n5384), .Z(n5489) );
  AND U5552 ( .A(n5490), .B(n5491), .Z(n5384) );
  NANDN U5553 ( .A(n5492), .B(n5493), .Z(n5491) );
  OR U5554 ( .A(n5494), .B(n5495), .Z(n5493) );
  NAND U5555 ( .A(n5495), .B(n5494), .Z(n5490) );
  ANDN U5556 ( .B(B[32]), .A(n30), .Z(n5386) );
  XNOR U5557 ( .A(n5394), .B(n5496), .Z(n5387) );
  XNOR U5558 ( .A(n5393), .B(n5391), .Z(n5496) );
  AND U5559 ( .A(n5497), .B(n5498), .Z(n5391) );
  NANDN U5560 ( .A(n5499), .B(n5500), .Z(n5498) );
  NANDN U5561 ( .A(n5501), .B(n5502), .Z(n5500) );
  NANDN U5562 ( .A(n5502), .B(n5501), .Z(n5497) );
  ANDN U5563 ( .B(B[33]), .A(n31), .Z(n5393) );
  XNOR U5564 ( .A(n5401), .B(n5503), .Z(n5394) );
  XNOR U5565 ( .A(n5400), .B(n5398), .Z(n5503) );
  AND U5566 ( .A(n5504), .B(n5505), .Z(n5398) );
  NANDN U5567 ( .A(n5506), .B(n5507), .Z(n5505) );
  OR U5568 ( .A(n5508), .B(n5509), .Z(n5507) );
  NAND U5569 ( .A(n5509), .B(n5508), .Z(n5504) );
  ANDN U5570 ( .B(B[34]), .A(n32), .Z(n5400) );
  XNOR U5571 ( .A(n5408), .B(n5510), .Z(n5401) );
  XNOR U5572 ( .A(n5407), .B(n5405), .Z(n5510) );
  AND U5573 ( .A(n5511), .B(n5512), .Z(n5405) );
  NANDN U5574 ( .A(n5513), .B(n5514), .Z(n5512) );
  NANDN U5575 ( .A(n5515), .B(n5516), .Z(n5514) );
  NANDN U5576 ( .A(n5516), .B(n5515), .Z(n5511) );
  ANDN U5577 ( .B(B[35]), .A(n33), .Z(n5407) );
  XNOR U5578 ( .A(n5415), .B(n5517), .Z(n5408) );
  XNOR U5579 ( .A(n5414), .B(n5412), .Z(n5517) );
  AND U5580 ( .A(n5518), .B(n5519), .Z(n5412) );
  NANDN U5581 ( .A(n5520), .B(n5521), .Z(n5519) );
  OR U5582 ( .A(n5522), .B(n5523), .Z(n5521) );
  NAND U5583 ( .A(n5523), .B(n5522), .Z(n5518) );
  ANDN U5584 ( .B(B[36]), .A(n34), .Z(n5414) );
  XNOR U5585 ( .A(n5422), .B(n5524), .Z(n5415) );
  XNOR U5586 ( .A(n5421), .B(n5419), .Z(n5524) );
  AND U5587 ( .A(n5525), .B(n5526), .Z(n5419) );
  NANDN U5588 ( .A(n5527), .B(n5528), .Z(n5526) );
  NANDN U5589 ( .A(n5529), .B(n5530), .Z(n5528) );
  NANDN U5590 ( .A(n5530), .B(n5529), .Z(n5525) );
  ANDN U5591 ( .B(B[37]), .A(n35), .Z(n5421) );
  XNOR U5592 ( .A(n5429), .B(n5531), .Z(n5422) );
  XNOR U5593 ( .A(n5428), .B(n5426), .Z(n5531) );
  AND U5594 ( .A(n5532), .B(n5533), .Z(n5426) );
  NANDN U5595 ( .A(n5534), .B(n5535), .Z(n5533) );
  OR U5596 ( .A(n5536), .B(n5537), .Z(n5535) );
  NAND U5597 ( .A(n5537), .B(n5536), .Z(n5532) );
  ANDN U5598 ( .B(B[38]), .A(n36), .Z(n5428) );
  XNOR U5599 ( .A(n5436), .B(n5538), .Z(n5429) );
  XNOR U5600 ( .A(n5435), .B(n5433), .Z(n5538) );
  AND U5601 ( .A(n5539), .B(n5540), .Z(n5433) );
  NANDN U5602 ( .A(n5541), .B(n5542), .Z(n5540) );
  NANDN U5603 ( .A(n5543), .B(n5544), .Z(n5542) );
  NANDN U5604 ( .A(n5544), .B(n5543), .Z(n5539) );
  ANDN U5605 ( .B(B[39]), .A(n37), .Z(n5435) );
  XNOR U5606 ( .A(n5443), .B(n5545), .Z(n5436) );
  XNOR U5607 ( .A(n5442), .B(n5440), .Z(n5545) );
  AND U5608 ( .A(n5546), .B(n5547), .Z(n5440) );
  NANDN U5609 ( .A(n5548), .B(n5549), .Z(n5547) );
  OR U5610 ( .A(n5550), .B(n5551), .Z(n5549) );
  NAND U5611 ( .A(n5551), .B(n5550), .Z(n5546) );
  ANDN U5612 ( .B(B[40]), .A(n38), .Z(n5442) );
  XNOR U5613 ( .A(n5450), .B(n5552), .Z(n5443) );
  XNOR U5614 ( .A(n5449), .B(n5447), .Z(n5552) );
  AND U5615 ( .A(n5553), .B(n5554), .Z(n5447) );
  NANDN U5616 ( .A(n5555), .B(n5556), .Z(n5554) );
  NANDN U5617 ( .A(n5557), .B(n5558), .Z(n5556) );
  NANDN U5618 ( .A(n5558), .B(n5557), .Z(n5553) );
  ANDN U5619 ( .B(B[41]), .A(n39), .Z(n5449) );
  XNOR U5620 ( .A(n5457), .B(n5559), .Z(n5450) );
  XNOR U5621 ( .A(n5456), .B(n5454), .Z(n5559) );
  AND U5622 ( .A(n5560), .B(n5561), .Z(n5454) );
  NANDN U5623 ( .A(n5562), .B(n5563), .Z(n5561) );
  OR U5624 ( .A(n5564), .B(n5565), .Z(n5563) );
  NAND U5625 ( .A(n5565), .B(n5564), .Z(n5560) );
  ANDN U5626 ( .B(B[42]), .A(n40), .Z(n5456) );
  XNOR U5627 ( .A(n5464), .B(n5566), .Z(n5457) );
  XNOR U5628 ( .A(n5463), .B(n5461), .Z(n5566) );
  AND U5629 ( .A(n5567), .B(n5568), .Z(n5461) );
  NANDN U5630 ( .A(n5569), .B(n5570), .Z(n5568) );
  NAND U5631 ( .A(n5571), .B(n5572), .Z(n5570) );
  ANDN U5632 ( .B(B[43]), .A(n41), .Z(n5463) );
  XOR U5633 ( .A(n5470), .B(n5573), .Z(n5464) );
  XNOR U5634 ( .A(n5468), .B(n5471), .Z(n5573) );
  NAND U5635 ( .A(A[2]), .B(B[44]), .Z(n5471) );
  NANDN U5636 ( .A(n5574), .B(n5575), .Z(n5468) );
  AND U5637 ( .A(A[0]), .B(B[45]), .Z(n5575) );
  XNOR U5638 ( .A(n5473), .B(n5576), .Z(n5470) );
  NAND U5639 ( .A(A[0]), .B(B[46]), .Z(n5576) );
  NAND U5640 ( .A(B[45]), .B(A[1]), .Z(n5473) );
  NAND U5641 ( .A(n5577), .B(n5578), .Z(n154) );
  NANDN U5642 ( .A(n5579), .B(n5580), .Z(n5578) );
  OR U5643 ( .A(n5581), .B(n5582), .Z(n5580) );
  NAND U5644 ( .A(n5582), .B(n5581), .Z(n5577) );
  XOR U5645 ( .A(n156), .B(n155), .Z(\A1[43] ) );
  XOR U5646 ( .A(n5582), .B(n5583), .Z(n155) );
  XNOR U5647 ( .A(n5581), .B(n5579), .Z(n5583) );
  AND U5648 ( .A(n5584), .B(n5585), .Z(n5579) );
  NANDN U5649 ( .A(n5586), .B(n5587), .Z(n5585) );
  NANDN U5650 ( .A(n5588), .B(n5589), .Z(n5587) );
  NANDN U5651 ( .A(n5589), .B(n5588), .Z(n5584) );
  ANDN U5652 ( .B(B[30]), .A(n29), .Z(n5581) );
  XNOR U5653 ( .A(n5488), .B(n5590), .Z(n5582) );
  XNOR U5654 ( .A(n5487), .B(n5485), .Z(n5590) );
  AND U5655 ( .A(n5591), .B(n5592), .Z(n5485) );
  NANDN U5656 ( .A(n5593), .B(n5594), .Z(n5592) );
  OR U5657 ( .A(n5595), .B(n5596), .Z(n5594) );
  NAND U5658 ( .A(n5596), .B(n5595), .Z(n5591) );
  ANDN U5659 ( .B(B[31]), .A(n30), .Z(n5487) );
  XNOR U5660 ( .A(n5495), .B(n5597), .Z(n5488) );
  XNOR U5661 ( .A(n5494), .B(n5492), .Z(n5597) );
  AND U5662 ( .A(n5598), .B(n5599), .Z(n5492) );
  NANDN U5663 ( .A(n5600), .B(n5601), .Z(n5599) );
  NANDN U5664 ( .A(n5602), .B(n5603), .Z(n5601) );
  NANDN U5665 ( .A(n5603), .B(n5602), .Z(n5598) );
  ANDN U5666 ( .B(B[32]), .A(n31), .Z(n5494) );
  XNOR U5667 ( .A(n5502), .B(n5604), .Z(n5495) );
  XNOR U5668 ( .A(n5501), .B(n5499), .Z(n5604) );
  AND U5669 ( .A(n5605), .B(n5606), .Z(n5499) );
  NANDN U5670 ( .A(n5607), .B(n5608), .Z(n5606) );
  OR U5671 ( .A(n5609), .B(n5610), .Z(n5608) );
  NAND U5672 ( .A(n5610), .B(n5609), .Z(n5605) );
  ANDN U5673 ( .B(B[33]), .A(n32), .Z(n5501) );
  XNOR U5674 ( .A(n5509), .B(n5611), .Z(n5502) );
  XNOR U5675 ( .A(n5508), .B(n5506), .Z(n5611) );
  AND U5676 ( .A(n5612), .B(n5613), .Z(n5506) );
  NANDN U5677 ( .A(n5614), .B(n5615), .Z(n5613) );
  NANDN U5678 ( .A(n5616), .B(n5617), .Z(n5615) );
  NANDN U5679 ( .A(n5617), .B(n5616), .Z(n5612) );
  ANDN U5680 ( .B(B[34]), .A(n33), .Z(n5508) );
  XNOR U5681 ( .A(n5516), .B(n5618), .Z(n5509) );
  XNOR U5682 ( .A(n5515), .B(n5513), .Z(n5618) );
  AND U5683 ( .A(n5619), .B(n5620), .Z(n5513) );
  NANDN U5684 ( .A(n5621), .B(n5622), .Z(n5620) );
  OR U5685 ( .A(n5623), .B(n5624), .Z(n5622) );
  NAND U5686 ( .A(n5624), .B(n5623), .Z(n5619) );
  ANDN U5687 ( .B(B[35]), .A(n34), .Z(n5515) );
  XNOR U5688 ( .A(n5523), .B(n5625), .Z(n5516) );
  XNOR U5689 ( .A(n5522), .B(n5520), .Z(n5625) );
  AND U5690 ( .A(n5626), .B(n5627), .Z(n5520) );
  NANDN U5691 ( .A(n5628), .B(n5629), .Z(n5627) );
  NANDN U5692 ( .A(n5630), .B(n5631), .Z(n5629) );
  NANDN U5693 ( .A(n5631), .B(n5630), .Z(n5626) );
  ANDN U5694 ( .B(B[36]), .A(n35), .Z(n5522) );
  XNOR U5695 ( .A(n5530), .B(n5632), .Z(n5523) );
  XNOR U5696 ( .A(n5529), .B(n5527), .Z(n5632) );
  AND U5697 ( .A(n5633), .B(n5634), .Z(n5527) );
  NANDN U5698 ( .A(n5635), .B(n5636), .Z(n5634) );
  OR U5699 ( .A(n5637), .B(n5638), .Z(n5636) );
  NAND U5700 ( .A(n5638), .B(n5637), .Z(n5633) );
  ANDN U5701 ( .B(B[37]), .A(n36), .Z(n5529) );
  XNOR U5702 ( .A(n5537), .B(n5639), .Z(n5530) );
  XNOR U5703 ( .A(n5536), .B(n5534), .Z(n5639) );
  AND U5704 ( .A(n5640), .B(n5641), .Z(n5534) );
  NANDN U5705 ( .A(n5642), .B(n5643), .Z(n5641) );
  NANDN U5706 ( .A(n5644), .B(n5645), .Z(n5643) );
  NANDN U5707 ( .A(n5645), .B(n5644), .Z(n5640) );
  ANDN U5708 ( .B(B[38]), .A(n37), .Z(n5536) );
  XNOR U5709 ( .A(n5544), .B(n5646), .Z(n5537) );
  XNOR U5710 ( .A(n5543), .B(n5541), .Z(n5646) );
  AND U5711 ( .A(n5647), .B(n5648), .Z(n5541) );
  NANDN U5712 ( .A(n5649), .B(n5650), .Z(n5648) );
  OR U5713 ( .A(n5651), .B(n5652), .Z(n5650) );
  NAND U5714 ( .A(n5652), .B(n5651), .Z(n5647) );
  ANDN U5715 ( .B(B[39]), .A(n38), .Z(n5543) );
  XNOR U5716 ( .A(n5551), .B(n5653), .Z(n5544) );
  XNOR U5717 ( .A(n5550), .B(n5548), .Z(n5653) );
  AND U5718 ( .A(n5654), .B(n5655), .Z(n5548) );
  NANDN U5719 ( .A(n5656), .B(n5657), .Z(n5655) );
  NANDN U5720 ( .A(n5658), .B(n5659), .Z(n5657) );
  NANDN U5721 ( .A(n5659), .B(n5658), .Z(n5654) );
  ANDN U5722 ( .B(B[40]), .A(n39), .Z(n5550) );
  XNOR U5723 ( .A(n5558), .B(n5660), .Z(n5551) );
  XNOR U5724 ( .A(n5557), .B(n5555), .Z(n5660) );
  AND U5725 ( .A(n5661), .B(n5662), .Z(n5555) );
  NANDN U5726 ( .A(n5663), .B(n5664), .Z(n5662) );
  OR U5727 ( .A(n5665), .B(n5666), .Z(n5664) );
  NAND U5728 ( .A(n5666), .B(n5665), .Z(n5661) );
  ANDN U5729 ( .B(B[41]), .A(n40), .Z(n5557) );
  XNOR U5730 ( .A(n5565), .B(n5667), .Z(n5558) );
  XNOR U5731 ( .A(n5564), .B(n5562), .Z(n5667) );
  AND U5732 ( .A(n5668), .B(n5669), .Z(n5562) );
  NANDN U5733 ( .A(n5670), .B(n5671), .Z(n5669) );
  NAND U5734 ( .A(n5672), .B(n5673), .Z(n5671) );
  ANDN U5735 ( .B(B[42]), .A(n41), .Z(n5564) );
  XOR U5736 ( .A(n5571), .B(n5674), .Z(n5565) );
  XNOR U5737 ( .A(n5569), .B(n5572), .Z(n5674) );
  NAND U5738 ( .A(A[2]), .B(B[43]), .Z(n5572) );
  NANDN U5739 ( .A(n5675), .B(n5676), .Z(n5569) );
  AND U5740 ( .A(A[0]), .B(B[44]), .Z(n5676) );
  XNOR U5741 ( .A(n5574), .B(n5677), .Z(n5571) );
  NAND U5742 ( .A(A[0]), .B(B[45]), .Z(n5677) );
  NAND U5743 ( .A(B[44]), .B(A[1]), .Z(n5574) );
  NAND U5744 ( .A(n5678), .B(n5679), .Z(n156) );
  NANDN U5745 ( .A(n5680), .B(n5681), .Z(n5679) );
  OR U5746 ( .A(n5682), .B(n5683), .Z(n5681) );
  NAND U5747 ( .A(n5683), .B(n5682), .Z(n5678) );
  XOR U5748 ( .A(n158), .B(n157), .Z(\A1[42] ) );
  XOR U5749 ( .A(n5683), .B(n5684), .Z(n157) );
  XNOR U5750 ( .A(n5682), .B(n5680), .Z(n5684) );
  AND U5751 ( .A(n5685), .B(n5686), .Z(n5680) );
  NANDN U5752 ( .A(n5687), .B(n5688), .Z(n5686) );
  NANDN U5753 ( .A(n5689), .B(n5690), .Z(n5688) );
  NANDN U5754 ( .A(n5690), .B(n5689), .Z(n5685) );
  ANDN U5755 ( .B(B[29]), .A(n29), .Z(n5682) );
  XNOR U5756 ( .A(n5589), .B(n5691), .Z(n5683) );
  XNOR U5757 ( .A(n5588), .B(n5586), .Z(n5691) );
  AND U5758 ( .A(n5692), .B(n5693), .Z(n5586) );
  NANDN U5759 ( .A(n5694), .B(n5695), .Z(n5693) );
  OR U5760 ( .A(n5696), .B(n5697), .Z(n5695) );
  NAND U5761 ( .A(n5697), .B(n5696), .Z(n5692) );
  ANDN U5762 ( .B(B[30]), .A(n30), .Z(n5588) );
  XNOR U5763 ( .A(n5596), .B(n5698), .Z(n5589) );
  XNOR U5764 ( .A(n5595), .B(n5593), .Z(n5698) );
  AND U5765 ( .A(n5699), .B(n5700), .Z(n5593) );
  NANDN U5766 ( .A(n5701), .B(n5702), .Z(n5700) );
  NANDN U5767 ( .A(n5703), .B(n5704), .Z(n5702) );
  NANDN U5768 ( .A(n5704), .B(n5703), .Z(n5699) );
  ANDN U5769 ( .B(B[31]), .A(n31), .Z(n5595) );
  XNOR U5770 ( .A(n5603), .B(n5705), .Z(n5596) );
  XNOR U5771 ( .A(n5602), .B(n5600), .Z(n5705) );
  AND U5772 ( .A(n5706), .B(n5707), .Z(n5600) );
  NANDN U5773 ( .A(n5708), .B(n5709), .Z(n5707) );
  OR U5774 ( .A(n5710), .B(n5711), .Z(n5709) );
  NAND U5775 ( .A(n5711), .B(n5710), .Z(n5706) );
  ANDN U5776 ( .B(B[32]), .A(n32), .Z(n5602) );
  XNOR U5777 ( .A(n5610), .B(n5712), .Z(n5603) );
  XNOR U5778 ( .A(n5609), .B(n5607), .Z(n5712) );
  AND U5779 ( .A(n5713), .B(n5714), .Z(n5607) );
  NANDN U5780 ( .A(n5715), .B(n5716), .Z(n5714) );
  NANDN U5781 ( .A(n5717), .B(n5718), .Z(n5716) );
  NANDN U5782 ( .A(n5718), .B(n5717), .Z(n5713) );
  ANDN U5783 ( .B(B[33]), .A(n33), .Z(n5609) );
  XNOR U5784 ( .A(n5617), .B(n5719), .Z(n5610) );
  XNOR U5785 ( .A(n5616), .B(n5614), .Z(n5719) );
  AND U5786 ( .A(n5720), .B(n5721), .Z(n5614) );
  NANDN U5787 ( .A(n5722), .B(n5723), .Z(n5721) );
  OR U5788 ( .A(n5724), .B(n5725), .Z(n5723) );
  NAND U5789 ( .A(n5725), .B(n5724), .Z(n5720) );
  ANDN U5790 ( .B(B[34]), .A(n34), .Z(n5616) );
  XNOR U5791 ( .A(n5624), .B(n5726), .Z(n5617) );
  XNOR U5792 ( .A(n5623), .B(n5621), .Z(n5726) );
  AND U5793 ( .A(n5727), .B(n5728), .Z(n5621) );
  NANDN U5794 ( .A(n5729), .B(n5730), .Z(n5728) );
  NANDN U5795 ( .A(n5731), .B(n5732), .Z(n5730) );
  NANDN U5796 ( .A(n5732), .B(n5731), .Z(n5727) );
  ANDN U5797 ( .B(B[35]), .A(n35), .Z(n5623) );
  XNOR U5798 ( .A(n5631), .B(n5733), .Z(n5624) );
  XNOR U5799 ( .A(n5630), .B(n5628), .Z(n5733) );
  AND U5800 ( .A(n5734), .B(n5735), .Z(n5628) );
  NANDN U5801 ( .A(n5736), .B(n5737), .Z(n5735) );
  OR U5802 ( .A(n5738), .B(n5739), .Z(n5737) );
  NAND U5803 ( .A(n5739), .B(n5738), .Z(n5734) );
  ANDN U5804 ( .B(B[36]), .A(n36), .Z(n5630) );
  XNOR U5805 ( .A(n5638), .B(n5740), .Z(n5631) );
  XNOR U5806 ( .A(n5637), .B(n5635), .Z(n5740) );
  AND U5807 ( .A(n5741), .B(n5742), .Z(n5635) );
  NANDN U5808 ( .A(n5743), .B(n5744), .Z(n5742) );
  NANDN U5809 ( .A(n5745), .B(n5746), .Z(n5744) );
  NANDN U5810 ( .A(n5746), .B(n5745), .Z(n5741) );
  ANDN U5811 ( .B(B[37]), .A(n37), .Z(n5637) );
  XNOR U5812 ( .A(n5645), .B(n5747), .Z(n5638) );
  XNOR U5813 ( .A(n5644), .B(n5642), .Z(n5747) );
  AND U5814 ( .A(n5748), .B(n5749), .Z(n5642) );
  NANDN U5815 ( .A(n5750), .B(n5751), .Z(n5749) );
  OR U5816 ( .A(n5752), .B(n5753), .Z(n5751) );
  NAND U5817 ( .A(n5753), .B(n5752), .Z(n5748) );
  ANDN U5818 ( .B(B[38]), .A(n38), .Z(n5644) );
  XNOR U5819 ( .A(n5652), .B(n5754), .Z(n5645) );
  XNOR U5820 ( .A(n5651), .B(n5649), .Z(n5754) );
  AND U5821 ( .A(n5755), .B(n5756), .Z(n5649) );
  NANDN U5822 ( .A(n5757), .B(n5758), .Z(n5756) );
  NANDN U5823 ( .A(n5759), .B(n5760), .Z(n5758) );
  NANDN U5824 ( .A(n5760), .B(n5759), .Z(n5755) );
  ANDN U5825 ( .B(B[39]), .A(n39), .Z(n5651) );
  XNOR U5826 ( .A(n5659), .B(n5761), .Z(n5652) );
  XNOR U5827 ( .A(n5658), .B(n5656), .Z(n5761) );
  AND U5828 ( .A(n5762), .B(n5763), .Z(n5656) );
  NANDN U5829 ( .A(n5764), .B(n5765), .Z(n5763) );
  OR U5830 ( .A(n5766), .B(n5767), .Z(n5765) );
  NAND U5831 ( .A(n5767), .B(n5766), .Z(n5762) );
  ANDN U5832 ( .B(B[40]), .A(n40), .Z(n5658) );
  XNOR U5833 ( .A(n5666), .B(n5768), .Z(n5659) );
  XNOR U5834 ( .A(n5665), .B(n5663), .Z(n5768) );
  AND U5835 ( .A(n5769), .B(n5770), .Z(n5663) );
  NANDN U5836 ( .A(n5771), .B(n5772), .Z(n5770) );
  NAND U5837 ( .A(n5773), .B(n5774), .Z(n5772) );
  ANDN U5838 ( .B(B[41]), .A(n41), .Z(n5665) );
  XOR U5839 ( .A(n5672), .B(n5775), .Z(n5666) );
  XNOR U5840 ( .A(n5670), .B(n5673), .Z(n5775) );
  NAND U5841 ( .A(A[2]), .B(B[42]), .Z(n5673) );
  NANDN U5842 ( .A(n5776), .B(n5777), .Z(n5670) );
  AND U5843 ( .A(A[0]), .B(B[43]), .Z(n5777) );
  XNOR U5844 ( .A(n5675), .B(n5778), .Z(n5672) );
  NAND U5845 ( .A(A[0]), .B(B[44]), .Z(n5778) );
  NAND U5846 ( .A(B[43]), .B(A[1]), .Z(n5675) );
  NAND U5847 ( .A(n5779), .B(n5780), .Z(n158) );
  NANDN U5848 ( .A(n5781), .B(n5782), .Z(n5780) );
  OR U5849 ( .A(n5783), .B(n5784), .Z(n5782) );
  NAND U5850 ( .A(n5784), .B(n5783), .Z(n5779) );
  XOR U5851 ( .A(n160), .B(n159), .Z(\A1[41] ) );
  XOR U5852 ( .A(n5784), .B(n5785), .Z(n159) );
  XNOR U5853 ( .A(n5783), .B(n5781), .Z(n5785) );
  AND U5854 ( .A(n5786), .B(n5787), .Z(n5781) );
  NANDN U5855 ( .A(n5788), .B(n5789), .Z(n5787) );
  NANDN U5856 ( .A(n5790), .B(n5791), .Z(n5789) );
  NANDN U5857 ( .A(n5791), .B(n5790), .Z(n5786) );
  ANDN U5858 ( .B(B[28]), .A(n29), .Z(n5783) );
  XNOR U5859 ( .A(n5690), .B(n5792), .Z(n5784) );
  XNOR U5860 ( .A(n5689), .B(n5687), .Z(n5792) );
  AND U5861 ( .A(n5793), .B(n5794), .Z(n5687) );
  NANDN U5862 ( .A(n5795), .B(n5796), .Z(n5794) );
  OR U5863 ( .A(n5797), .B(n5798), .Z(n5796) );
  NAND U5864 ( .A(n5798), .B(n5797), .Z(n5793) );
  ANDN U5865 ( .B(B[29]), .A(n30), .Z(n5689) );
  XNOR U5866 ( .A(n5697), .B(n5799), .Z(n5690) );
  XNOR U5867 ( .A(n5696), .B(n5694), .Z(n5799) );
  AND U5868 ( .A(n5800), .B(n5801), .Z(n5694) );
  NANDN U5869 ( .A(n5802), .B(n5803), .Z(n5801) );
  NANDN U5870 ( .A(n5804), .B(n5805), .Z(n5803) );
  NANDN U5871 ( .A(n5805), .B(n5804), .Z(n5800) );
  ANDN U5872 ( .B(B[30]), .A(n31), .Z(n5696) );
  XNOR U5873 ( .A(n5704), .B(n5806), .Z(n5697) );
  XNOR U5874 ( .A(n5703), .B(n5701), .Z(n5806) );
  AND U5875 ( .A(n5807), .B(n5808), .Z(n5701) );
  NANDN U5876 ( .A(n5809), .B(n5810), .Z(n5808) );
  OR U5877 ( .A(n5811), .B(n5812), .Z(n5810) );
  NAND U5878 ( .A(n5812), .B(n5811), .Z(n5807) );
  ANDN U5879 ( .B(B[31]), .A(n32), .Z(n5703) );
  XNOR U5880 ( .A(n5711), .B(n5813), .Z(n5704) );
  XNOR U5881 ( .A(n5710), .B(n5708), .Z(n5813) );
  AND U5882 ( .A(n5814), .B(n5815), .Z(n5708) );
  NANDN U5883 ( .A(n5816), .B(n5817), .Z(n5815) );
  NANDN U5884 ( .A(n5818), .B(n5819), .Z(n5817) );
  NANDN U5885 ( .A(n5819), .B(n5818), .Z(n5814) );
  ANDN U5886 ( .B(B[32]), .A(n33), .Z(n5710) );
  XNOR U5887 ( .A(n5718), .B(n5820), .Z(n5711) );
  XNOR U5888 ( .A(n5717), .B(n5715), .Z(n5820) );
  AND U5889 ( .A(n5821), .B(n5822), .Z(n5715) );
  NANDN U5890 ( .A(n5823), .B(n5824), .Z(n5822) );
  OR U5891 ( .A(n5825), .B(n5826), .Z(n5824) );
  NAND U5892 ( .A(n5826), .B(n5825), .Z(n5821) );
  ANDN U5893 ( .B(B[33]), .A(n34), .Z(n5717) );
  XNOR U5894 ( .A(n5725), .B(n5827), .Z(n5718) );
  XNOR U5895 ( .A(n5724), .B(n5722), .Z(n5827) );
  AND U5896 ( .A(n5828), .B(n5829), .Z(n5722) );
  NANDN U5897 ( .A(n5830), .B(n5831), .Z(n5829) );
  NANDN U5898 ( .A(n5832), .B(n5833), .Z(n5831) );
  NANDN U5899 ( .A(n5833), .B(n5832), .Z(n5828) );
  ANDN U5900 ( .B(B[34]), .A(n35), .Z(n5724) );
  XNOR U5901 ( .A(n5732), .B(n5834), .Z(n5725) );
  XNOR U5902 ( .A(n5731), .B(n5729), .Z(n5834) );
  AND U5903 ( .A(n5835), .B(n5836), .Z(n5729) );
  NANDN U5904 ( .A(n5837), .B(n5838), .Z(n5836) );
  OR U5905 ( .A(n5839), .B(n5840), .Z(n5838) );
  NAND U5906 ( .A(n5840), .B(n5839), .Z(n5835) );
  ANDN U5907 ( .B(B[35]), .A(n36), .Z(n5731) );
  XNOR U5908 ( .A(n5739), .B(n5841), .Z(n5732) );
  XNOR U5909 ( .A(n5738), .B(n5736), .Z(n5841) );
  AND U5910 ( .A(n5842), .B(n5843), .Z(n5736) );
  NANDN U5911 ( .A(n5844), .B(n5845), .Z(n5843) );
  NANDN U5912 ( .A(n5846), .B(n5847), .Z(n5845) );
  NANDN U5913 ( .A(n5847), .B(n5846), .Z(n5842) );
  ANDN U5914 ( .B(B[36]), .A(n37), .Z(n5738) );
  XNOR U5915 ( .A(n5746), .B(n5848), .Z(n5739) );
  XNOR U5916 ( .A(n5745), .B(n5743), .Z(n5848) );
  AND U5917 ( .A(n5849), .B(n5850), .Z(n5743) );
  NANDN U5918 ( .A(n5851), .B(n5852), .Z(n5850) );
  OR U5919 ( .A(n5853), .B(n5854), .Z(n5852) );
  NAND U5920 ( .A(n5854), .B(n5853), .Z(n5849) );
  ANDN U5921 ( .B(B[37]), .A(n38), .Z(n5745) );
  XNOR U5922 ( .A(n5753), .B(n5855), .Z(n5746) );
  XNOR U5923 ( .A(n5752), .B(n5750), .Z(n5855) );
  AND U5924 ( .A(n5856), .B(n5857), .Z(n5750) );
  NANDN U5925 ( .A(n5858), .B(n5859), .Z(n5857) );
  NANDN U5926 ( .A(n5860), .B(n5861), .Z(n5859) );
  NANDN U5927 ( .A(n5861), .B(n5860), .Z(n5856) );
  ANDN U5928 ( .B(B[38]), .A(n39), .Z(n5752) );
  XNOR U5929 ( .A(n5760), .B(n5862), .Z(n5753) );
  XNOR U5930 ( .A(n5759), .B(n5757), .Z(n5862) );
  AND U5931 ( .A(n5863), .B(n5864), .Z(n5757) );
  NANDN U5932 ( .A(n5865), .B(n5866), .Z(n5864) );
  OR U5933 ( .A(n5867), .B(n5868), .Z(n5866) );
  NAND U5934 ( .A(n5868), .B(n5867), .Z(n5863) );
  ANDN U5935 ( .B(B[39]), .A(n40), .Z(n5759) );
  XNOR U5936 ( .A(n5767), .B(n5869), .Z(n5760) );
  XNOR U5937 ( .A(n5766), .B(n5764), .Z(n5869) );
  AND U5938 ( .A(n5870), .B(n5871), .Z(n5764) );
  NANDN U5939 ( .A(n5872), .B(n5873), .Z(n5871) );
  NAND U5940 ( .A(n5874), .B(n5875), .Z(n5873) );
  ANDN U5941 ( .B(B[40]), .A(n41), .Z(n5766) );
  XOR U5942 ( .A(n5773), .B(n5876), .Z(n5767) );
  XNOR U5943 ( .A(n5771), .B(n5774), .Z(n5876) );
  NAND U5944 ( .A(A[2]), .B(B[41]), .Z(n5774) );
  NANDN U5945 ( .A(n5877), .B(n5878), .Z(n5771) );
  AND U5946 ( .A(A[0]), .B(B[42]), .Z(n5878) );
  XNOR U5947 ( .A(n5776), .B(n5879), .Z(n5773) );
  NAND U5948 ( .A(A[0]), .B(B[43]), .Z(n5879) );
  NAND U5949 ( .A(B[42]), .B(A[1]), .Z(n5776) );
  NAND U5950 ( .A(n5880), .B(n5881), .Z(n160) );
  NANDN U5951 ( .A(n5882), .B(n5883), .Z(n5881) );
  OR U5952 ( .A(n5884), .B(n5885), .Z(n5883) );
  NAND U5953 ( .A(n5885), .B(n5884), .Z(n5880) );
  XOR U5954 ( .A(n162), .B(n161), .Z(\A1[40] ) );
  XOR U5955 ( .A(n5885), .B(n5886), .Z(n161) );
  XNOR U5956 ( .A(n5884), .B(n5882), .Z(n5886) );
  AND U5957 ( .A(n5887), .B(n5888), .Z(n5882) );
  NANDN U5958 ( .A(n5889), .B(n5890), .Z(n5888) );
  NANDN U5959 ( .A(n5891), .B(n5892), .Z(n5890) );
  NANDN U5960 ( .A(n5892), .B(n5891), .Z(n5887) );
  ANDN U5961 ( .B(B[27]), .A(n29), .Z(n5884) );
  XNOR U5962 ( .A(n5791), .B(n5893), .Z(n5885) );
  XNOR U5963 ( .A(n5790), .B(n5788), .Z(n5893) );
  AND U5964 ( .A(n5894), .B(n5895), .Z(n5788) );
  NANDN U5965 ( .A(n5896), .B(n5897), .Z(n5895) );
  OR U5966 ( .A(n5898), .B(n5899), .Z(n5897) );
  NAND U5967 ( .A(n5899), .B(n5898), .Z(n5894) );
  ANDN U5968 ( .B(B[28]), .A(n30), .Z(n5790) );
  XNOR U5969 ( .A(n5798), .B(n5900), .Z(n5791) );
  XNOR U5970 ( .A(n5797), .B(n5795), .Z(n5900) );
  AND U5971 ( .A(n5901), .B(n5902), .Z(n5795) );
  NANDN U5972 ( .A(n5903), .B(n5904), .Z(n5902) );
  NANDN U5973 ( .A(n5905), .B(n5906), .Z(n5904) );
  NANDN U5974 ( .A(n5906), .B(n5905), .Z(n5901) );
  ANDN U5975 ( .B(B[29]), .A(n31), .Z(n5797) );
  XNOR U5976 ( .A(n5805), .B(n5907), .Z(n5798) );
  XNOR U5977 ( .A(n5804), .B(n5802), .Z(n5907) );
  AND U5978 ( .A(n5908), .B(n5909), .Z(n5802) );
  NANDN U5979 ( .A(n5910), .B(n5911), .Z(n5909) );
  OR U5980 ( .A(n5912), .B(n5913), .Z(n5911) );
  NAND U5981 ( .A(n5913), .B(n5912), .Z(n5908) );
  ANDN U5982 ( .B(B[30]), .A(n32), .Z(n5804) );
  XNOR U5983 ( .A(n5812), .B(n5914), .Z(n5805) );
  XNOR U5984 ( .A(n5811), .B(n5809), .Z(n5914) );
  AND U5985 ( .A(n5915), .B(n5916), .Z(n5809) );
  NANDN U5986 ( .A(n5917), .B(n5918), .Z(n5916) );
  NANDN U5987 ( .A(n5919), .B(n5920), .Z(n5918) );
  NANDN U5988 ( .A(n5920), .B(n5919), .Z(n5915) );
  ANDN U5989 ( .B(B[31]), .A(n33), .Z(n5811) );
  XNOR U5990 ( .A(n5819), .B(n5921), .Z(n5812) );
  XNOR U5991 ( .A(n5818), .B(n5816), .Z(n5921) );
  AND U5992 ( .A(n5922), .B(n5923), .Z(n5816) );
  NANDN U5993 ( .A(n5924), .B(n5925), .Z(n5923) );
  OR U5994 ( .A(n5926), .B(n5927), .Z(n5925) );
  NAND U5995 ( .A(n5927), .B(n5926), .Z(n5922) );
  ANDN U5996 ( .B(B[32]), .A(n34), .Z(n5818) );
  XNOR U5997 ( .A(n5826), .B(n5928), .Z(n5819) );
  XNOR U5998 ( .A(n5825), .B(n5823), .Z(n5928) );
  AND U5999 ( .A(n5929), .B(n5930), .Z(n5823) );
  NANDN U6000 ( .A(n5931), .B(n5932), .Z(n5930) );
  NANDN U6001 ( .A(n5933), .B(n5934), .Z(n5932) );
  NANDN U6002 ( .A(n5934), .B(n5933), .Z(n5929) );
  ANDN U6003 ( .B(B[33]), .A(n35), .Z(n5825) );
  XNOR U6004 ( .A(n5833), .B(n5935), .Z(n5826) );
  XNOR U6005 ( .A(n5832), .B(n5830), .Z(n5935) );
  AND U6006 ( .A(n5936), .B(n5937), .Z(n5830) );
  NANDN U6007 ( .A(n5938), .B(n5939), .Z(n5937) );
  OR U6008 ( .A(n5940), .B(n5941), .Z(n5939) );
  NAND U6009 ( .A(n5941), .B(n5940), .Z(n5936) );
  ANDN U6010 ( .B(B[34]), .A(n36), .Z(n5832) );
  XNOR U6011 ( .A(n5840), .B(n5942), .Z(n5833) );
  XNOR U6012 ( .A(n5839), .B(n5837), .Z(n5942) );
  AND U6013 ( .A(n5943), .B(n5944), .Z(n5837) );
  NANDN U6014 ( .A(n5945), .B(n5946), .Z(n5944) );
  NANDN U6015 ( .A(n5947), .B(n5948), .Z(n5946) );
  NANDN U6016 ( .A(n5948), .B(n5947), .Z(n5943) );
  ANDN U6017 ( .B(B[35]), .A(n37), .Z(n5839) );
  XNOR U6018 ( .A(n5847), .B(n5949), .Z(n5840) );
  XNOR U6019 ( .A(n5846), .B(n5844), .Z(n5949) );
  AND U6020 ( .A(n5950), .B(n5951), .Z(n5844) );
  NANDN U6021 ( .A(n5952), .B(n5953), .Z(n5951) );
  OR U6022 ( .A(n5954), .B(n5955), .Z(n5953) );
  NAND U6023 ( .A(n5955), .B(n5954), .Z(n5950) );
  ANDN U6024 ( .B(B[36]), .A(n38), .Z(n5846) );
  XNOR U6025 ( .A(n5854), .B(n5956), .Z(n5847) );
  XNOR U6026 ( .A(n5853), .B(n5851), .Z(n5956) );
  AND U6027 ( .A(n5957), .B(n5958), .Z(n5851) );
  NANDN U6028 ( .A(n5959), .B(n5960), .Z(n5958) );
  NANDN U6029 ( .A(n5961), .B(n5962), .Z(n5960) );
  NANDN U6030 ( .A(n5962), .B(n5961), .Z(n5957) );
  ANDN U6031 ( .B(B[37]), .A(n39), .Z(n5853) );
  XNOR U6032 ( .A(n5861), .B(n5963), .Z(n5854) );
  XNOR U6033 ( .A(n5860), .B(n5858), .Z(n5963) );
  AND U6034 ( .A(n5964), .B(n5965), .Z(n5858) );
  NANDN U6035 ( .A(n5966), .B(n5967), .Z(n5965) );
  OR U6036 ( .A(n5968), .B(n5969), .Z(n5967) );
  NAND U6037 ( .A(n5969), .B(n5968), .Z(n5964) );
  ANDN U6038 ( .B(B[38]), .A(n40), .Z(n5860) );
  XNOR U6039 ( .A(n5868), .B(n5970), .Z(n5861) );
  XNOR U6040 ( .A(n5867), .B(n5865), .Z(n5970) );
  AND U6041 ( .A(n5971), .B(n5972), .Z(n5865) );
  NANDN U6042 ( .A(n5973), .B(n5974), .Z(n5972) );
  NAND U6043 ( .A(n5975), .B(n5976), .Z(n5974) );
  ANDN U6044 ( .B(B[39]), .A(n41), .Z(n5867) );
  XOR U6045 ( .A(n5874), .B(n5977), .Z(n5868) );
  XNOR U6046 ( .A(n5872), .B(n5875), .Z(n5977) );
  NAND U6047 ( .A(A[2]), .B(B[40]), .Z(n5875) );
  NANDN U6048 ( .A(n5978), .B(n5979), .Z(n5872) );
  AND U6049 ( .A(A[0]), .B(B[41]), .Z(n5979) );
  XNOR U6050 ( .A(n5877), .B(n5980), .Z(n5874) );
  NAND U6051 ( .A(A[0]), .B(B[42]), .Z(n5980) );
  NAND U6052 ( .A(B[41]), .B(A[1]), .Z(n5877) );
  NAND U6053 ( .A(n5981), .B(n5982), .Z(n162) );
  NANDN U6054 ( .A(n5983), .B(n5984), .Z(n5982) );
  OR U6055 ( .A(n5985), .B(n5986), .Z(n5984) );
  NAND U6056 ( .A(n5986), .B(n5985), .Z(n5981) );
  XOR U6057 ( .A(n5987), .B(n5988), .Z(\A1[3] ) );
  XNOR U6058 ( .A(n5989), .B(n27), .Z(n5988) );
  XOR U6059 ( .A(n164), .B(n163), .Z(\A1[39] ) );
  XOR U6060 ( .A(n5986), .B(n5990), .Z(n163) );
  XNOR U6061 ( .A(n5985), .B(n5983), .Z(n5990) );
  AND U6062 ( .A(n5991), .B(n5992), .Z(n5983) );
  NANDN U6063 ( .A(n5993), .B(n5994), .Z(n5992) );
  NANDN U6064 ( .A(n5995), .B(n5996), .Z(n5994) );
  NANDN U6065 ( .A(n5996), .B(n5995), .Z(n5991) );
  ANDN U6066 ( .B(B[26]), .A(n29), .Z(n5985) );
  XNOR U6067 ( .A(n5892), .B(n5997), .Z(n5986) );
  XNOR U6068 ( .A(n5891), .B(n5889), .Z(n5997) );
  AND U6069 ( .A(n5998), .B(n5999), .Z(n5889) );
  NANDN U6070 ( .A(n6000), .B(n6001), .Z(n5999) );
  OR U6071 ( .A(n6002), .B(n6003), .Z(n6001) );
  NAND U6072 ( .A(n6003), .B(n6002), .Z(n5998) );
  ANDN U6073 ( .B(B[27]), .A(n30), .Z(n5891) );
  XNOR U6074 ( .A(n5899), .B(n6004), .Z(n5892) );
  XNOR U6075 ( .A(n5898), .B(n5896), .Z(n6004) );
  AND U6076 ( .A(n6005), .B(n6006), .Z(n5896) );
  NANDN U6077 ( .A(n6007), .B(n6008), .Z(n6006) );
  NANDN U6078 ( .A(n6009), .B(n6010), .Z(n6008) );
  NANDN U6079 ( .A(n6010), .B(n6009), .Z(n6005) );
  ANDN U6080 ( .B(B[28]), .A(n31), .Z(n5898) );
  XNOR U6081 ( .A(n5906), .B(n6011), .Z(n5899) );
  XNOR U6082 ( .A(n5905), .B(n5903), .Z(n6011) );
  AND U6083 ( .A(n6012), .B(n6013), .Z(n5903) );
  NANDN U6084 ( .A(n6014), .B(n6015), .Z(n6013) );
  OR U6085 ( .A(n6016), .B(n6017), .Z(n6015) );
  NAND U6086 ( .A(n6017), .B(n6016), .Z(n6012) );
  ANDN U6087 ( .B(B[29]), .A(n32), .Z(n5905) );
  XNOR U6088 ( .A(n5913), .B(n6018), .Z(n5906) );
  XNOR U6089 ( .A(n5912), .B(n5910), .Z(n6018) );
  AND U6090 ( .A(n6019), .B(n6020), .Z(n5910) );
  NANDN U6091 ( .A(n6021), .B(n6022), .Z(n6020) );
  NANDN U6092 ( .A(n6023), .B(n6024), .Z(n6022) );
  NANDN U6093 ( .A(n6024), .B(n6023), .Z(n6019) );
  ANDN U6094 ( .B(B[30]), .A(n33), .Z(n5912) );
  XNOR U6095 ( .A(n5920), .B(n6025), .Z(n5913) );
  XNOR U6096 ( .A(n5919), .B(n5917), .Z(n6025) );
  AND U6097 ( .A(n6026), .B(n6027), .Z(n5917) );
  NANDN U6098 ( .A(n6028), .B(n6029), .Z(n6027) );
  OR U6099 ( .A(n6030), .B(n6031), .Z(n6029) );
  NAND U6100 ( .A(n6031), .B(n6030), .Z(n6026) );
  ANDN U6101 ( .B(B[31]), .A(n34), .Z(n5919) );
  XNOR U6102 ( .A(n5927), .B(n6032), .Z(n5920) );
  XNOR U6103 ( .A(n5926), .B(n5924), .Z(n6032) );
  AND U6104 ( .A(n6033), .B(n6034), .Z(n5924) );
  NANDN U6105 ( .A(n6035), .B(n6036), .Z(n6034) );
  NANDN U6106 ( .A(n6037), .B(n6038), .Z(n6036) );
  NANDN U6107 ( .A(n6038), .B(n6037), .Z(n6033) );
  ANDN U6108 ( .B(B[32]), .A(n35), .Z(n5926) );
  XNOR U6109 ( .A(n5934), .B(n6039), .Z(n5927) );
  XNOR U6110 ( .A(n5933), .B(n5931), .Z(n6039) );
  AND U6111 ( .A(n6040), .B(n6041), .Z(n5931) );
  NANDN U6112 ( .A(n6042), .B(n6043), .Z(n6041) );
  OR U6113 ( .A(n6044), .B(n6045), .Z(n6043) );
  NAND U6114 ( .A(n6045), .B(n6044), .Z(n6040) );
  ANDN U6115 ( .B(B[33]), .A(n36), .Z(n5933) );
  XNOR U6116 ( .A(n5941), .B(n6046), .Z(n5934) );
  XNOR U6117 ( .A(n5940), .B(n5938), .Z(n6046) );
  AND U6118 ( .A(n6047), .B(n6048), .Z(n5938) );
  NANDN U6119 ( .A(n6049), .B(n6050), .Z(n6048) );
  NANDN U6120 ( .A(n6051), .B(n6052), .Z(n6050) );
  NANDN U6121 ( .A(n6052), .B(n6051), .Z(n6047) );
  ANDN U6122 ( .B(B[34]), .A(n37), .Z(n5940) );
  XNOR U6123 ( .A(n5948), .B(n6053), .Z(n5941) );
  XNOR U6124 ( .A(n5947), .B(n5945), .Z(n6053) );
  AND U6125 ( .A(n6054), .B(n6055), .Z(n5945) );
  NANDN U6126 ( .A(n6056), .B(n6057), .Z(n6055) );
  OR U6127 ( .A(n6058), .B(n6059), .Z(n6057) );
  NAND U6128 ( .A(n6059), .B(n6058), .Z(n6054) );
  ANDN U6129 ( .B(B[35]), .A(n38), .Z(n5947) );
  XNOR U6130 ( .A(n5955), .B(n6060), .Z(n5948) );
  XNOR U6131 ( .A(n5954), .B(n5952), .Z(n6060) );
  AND U6132 ( .A(n6061), .B(n6062), .Z(n5952) );
  NANDN U6133 ( .A(n6063), .B(n6064), .Z(n6062) );
  NANDN U6134 ( .A(n6065), .B(n6066), .Z(n6064) );
  NANDN U6135 ( .A(n6066), .B(n6065), .Z(n6061) );
  ANDN U6136 ( .B(B[36]), .A(n39), .Z(n5954) );
  XNOR U6137 ( .A(n5962), .B(n6067), .Z(n5955) );
  XNOR U6138 ( .A(n5961), .B(n5959), .Z(n6067) );
  AND U6139 ( .A(n6068), .B(n6069), .Z(n5959) );
  NANDN U6140 ( .A(n6070), .B(n6071), .Z(n6069) );
  OR U6141 ( .A(n6072), .B(n6073), .Z(n6071) );
  NAND U6142 ( .A(n6073), .B(n6072), .Z(n6068) );
  ANDN U6143 ( .B(B[37]), .A(n40), .Z(n5961) );
  XNOR U6144 ( .A(n5969), .B(n6074), .Z(n5962) );
  XNOR U6145 ( .A(n5968), .B(n5966), .Z(n6074) );
  AND U6146 ( .A(n6075), .B(n6076), .Z(n5966) );
  NANDN U6147 ( .A(n6077), .B(n6078), .Z(n6076) );
  NAND U6148 ( .A(n6079), .B(n6080), .Z(n6078) );
  ANDN U6149 ( .B(B[38]), .A(n41), .Z(n5968) );
  XOR U6150 ( .A(n5975), .B(n6081), .Z(n5969) );
  XNOR U6151 ( .A(n5973), .B(n5976), .Z(n6081) );
  NAND U6152 ( .A(A[2]), .B(B[39]), .Z(n5976) );
  NANDN U6153 ( .A(n6082), .B(n6083), .Z(n5973) );
  AND U6154 ( .A(A[0]), .B(B[40]), .Z(n6083) );
  XNOR U6155 ( .A(n5978), .B(n6084), .Z(n5975) );
  NAND U6156 ( .A(A[0]), .B(B[41]), .Z(n6084) );
  NAND U6157 ( .A(B[40]), .B(A[1]), .Z(n5978) );
  NAND U6158 ( .A(n6085), .B(n6086), .Z(n164) );
  NANDN U6159 ( .A(n6087), .B(n6088), .Z(n6086) );
  OR U6160 ( .A(n6089), .B(n6090), .Z(n6088) );
  NAND U6161 ( .A(n6090), .B(n6089), .Z(n6085) );
  XOR U6162 ( .A(n166), .B(n165), .Z(\A1[38] ) );
  XOR U6163 ( .A(n6090), .B(n6091), .Z(n165) );
  XNOR U6164 ( .A(n6089), .B(n6087), .Z(n6091) );
  AND U6165 ( .A(n6092), .B(n6093), .Z(n6087) );
  NANDN U6166 ( .A(n6094), .B(n6095), .Z(n6093) );
  NANDN U6167 ( .A(n6096), .B(n6097), .Z(n6095) );
  NANDN U6168 ( .A(n6097), .B(n6096), .Z(n6092) );
  ANDN U6169 ( .B(B[25]), .A(n29), .Z(n6089) );
  XNOR U6170 ( .A(n5996), .B(n6098), .Z(n6090) );
  XNOR U6171 ( .A(n5995), .B(n5993), .Z(n6098) );
  AND U6172 ( .A(n6099), .B(n6100), .Z(n5993) );
  NANDN U6173 ( .A(n6101), .B(n6102), .Z(n6100) );
  OR U6174 ( .A(n6103), .B(n6104), .Z(n6102) );
  NAND U6175 ( .A(n6104), .B(n6103), .Z(n6099) );
  ANDN U6176 ( .B(B[26]), .A(n30), .Z(n5995) );
  XNOR U6177 ( .A(n6003), .B(n6105), .Z(n5996) );
  XNOR U6178 ( .A(n6002), .B(n6000), .Z(n6105) );
  AND U6179 ( .A(n6106), .B(n6107), .Z(n6000) );
  NANDN U6180 ( .A(n6108), .B(n6109), .Z(n6107) );
  NANDN U6181 ( .A(n6110), .B(n6111), .Z(n6109) );
  NANDN U6182 ( .A(n6111), .B(n6110), .Z(n6106) );
  ANDN U6183 ( .B(B[27]), .A(n31), .Z(n6002) );
  XNOR U6184 ( .A(n6010), .B(n6112), .Z(n6003) );
  XNOR U6185 ( .A(n6009), .B(n6007), .Z(n6112) );
  AND U6186 ( .A(n6113), .B(n6114), .Z(n6007) );
  NANDN U6187 ( .A(n6115), .B(n6116), .Z(n6114) );
  OR U6188 ( .A(n6117), .B(n6118), .Z(n6116) );
  NAND U6189 ( .A(n6118), .B(n6117), .Z(n6113) );
  ANDN U6190 ( .B(B[28]), .A(n32), .Z(n6009) );
  XNOR U6191 ( .A(n6017), .B(n6119), .Z(n6010) );
  XNOR U6192 ( .A(n6016), .B(n6014), .Z(n6119) );
  AND U6193 ( .A(n6120), .B(n6121), .Z(n6014) );
  NANDN U6194 ( .A(n6122), .B(n6123), .Z(n6121) );
  NANDN U6195 ( .A(n6124), .B(n6125), .Z(n6123) );
  NANDN U6196 ( .A(n6125), .B(n6124), .Z(n6120) );
  ANDN U6197 ( .B(B[29]), .A(n33), .Z(n6016) );
  XNOR U6198 ( .A(n6024), .B(n6126), .Z(n6017) );
  XNOR U6199 ( .A(n6023), .B(n6021), .Z(n6126) );
  AND U6200 ( .A(n6127), .B(n6128), .Z(n6021) );
  NANDN U6201 ( .A(n6129), .B(n6130), .Z(n6128) );
  OR U6202 ( .A(n6131), .B(n6132), .Z(n6130) );
  NAND U6203 ( .A(n6132), .B(n6131), .Z(n6127) );
  ANDN U6204 ( .B(B[30]), .A(n34), .Z(n6023) );
  XNOR U6205 ( .A(n6031), .B(n6133), .Z(n6024) );
  XNOR U6206 ( .A(n6030), .B(n6028), .Z(n6133) );
  AND U6207 ( .A(n6134), .B(n6135), .Z(n6028) );
  NANDN U6208 ( .A(n6136), .B(n6137), .Z(n6135) );
  NANDN U6209 ( .A(n6138), .B(n6139), .Z(n6137) );
  NANDN U6210 ( .A(n6139), .B(n6138), .Z(n6134) );
  ANDN U6211 ( .B(B[31]), .A(n35), .Z(n6030) );
  XNOR U6212 ( .A(n6038), .B(n6140), .Z(n6031) );
  XNOR U6213 ( .A(n6037), .B(n6035), .Z(n6140) );
  AND U6214 ( .A(n6141), .B(n6142), .Z(n6035) );
  NANDN U6215 ( .A(n6143), .B(n6144), .Z(n6142) );
  OR U6216 ( .A(n6145), .B(n6146), .Z(n6144) );
  NAND U6217 ( .A(n6146), .B(n6145), .Z(n6141) );
  ANDN U6218 ( .B(B[32]), .A(n36), .Z(n6037) );
  XNOR U6219 ( .A(n6045), .B(n6147), .Z(n6038) );
  XNOR U6220 ( .A(n6044), .B(n6042), .Z(n6147) );
  AND U6221 ( .A(n6148), .B(n6149), .Z(n6042) );
  NANDN U6222 ( .A(n6150), .B(n6151), .Z(n6149) );
  NANDN U6223 ( .A(n6152), .B(n6153), .Z(n6151) );
  NANDN U6224 ( .A(n6153), .B(n6152), .Z(n6148) );
  ANDN U6225 ( .B(B[33]), .A(n37), .Z(n6044) );
  XNOR U6226 ( .A(n6052), .B(n6154), .Z(n6045) );
  XNOR U6227 ( .A(n6051), .B(n6049), .Z(n6154) );
  AND U6228 ( .A(n6155), .B(n6156), .Z(n6049) );
  NANDN U6229 ( .A(n6157), .B(n6158), .Z(n6156) );
  OR U6230 ( .A(n6159), .B(n6160), .Z(n6158) );
  NAND U6231 ( .A(n6160), .B(n6159), .Z(n6155) );
  ANDN U6232 ( .B(B[34]), .A(n38), .Z(n6051) );
  XNOR U6233 ( .A(n6059), .B(n6161), .Z(n6052) );
  XNOR U6234 ( .A(n6058), .B(n6056), .Z(n6161) );
  AND U6235 ( .A(n6162), .B(n6163), .Z(n6056) );
  NANDN U6236 ( .A(n6164), .B(n6165), .Z(n6163) );
  NANDN U6237 ( .A(n6166), .B(n6167), .Z(n6165) );
  NANDN U6238 ( .A(n6167), .B(n6166), .Z(n6162) );
  ANDN U6239 ( .B(B[35]), .A(n39), .Z(n6058) );
  XNOR U6240 ( .A(n6066), .B(n6168), .Z(n6059) );
  XNOR U6241 ( .A(n6065), .B(n6063), .Z(n6168) );
  AND U6242 ( .A(n6169), .B(n6170), .Z(n6063) );
  NANDN U6243 ( .A(n6171), .B(n6172), .Z(n6170) );
  OR U6244 ( .A(n6173), .B(n6174), .Z(n6172) );
  NAND U6245 ( .A(n6174), .B(n6173), .Z(n6169) );
  ANDN U6246 ( .B(B[36]), .A(n40), .Z(n6065) );
  XNOR U6247 ( .A(n6073), .B(n6175), .Z(n6066) );
  XNOR U6248 ( .A(n6072), .B(n6070), .Z(n6175) );
  AND U6249 ( .A(n6176), .B(n6177), .Z(n6070) );
  NANDN U6250 ( .A(n6178), .B(n6179), .Z(n6177) );
  NAND U6251 ( .A(n6180), .B(n6181), .Z(n6179) );
  ANDN U6252 ( .B(B[37]), .A(n41), .Z(n6072) );
  XOR U6253 ( .A(n6079), .B(n6182), .Z(n6073) );
  XNOR U6254 ( .A(n6077), .B(n6080), .Z(n6182) );
  NAND U6255 ( .A(A[2]), .B(B[38]), .Z(n6080) );
  NANDN U6256 ( .A(n6183), .B(n6184), .Z(n6077) );
  AND U6257 ( .A(A[0]), .B(B[39]), .Z(n6184) );
  XNOR U6258 ( .A(n6082), .B(n6185), .Z(n6079) );
  NAND U6259 ( .A(A[0]), .B(B[40]), .Z(n6185) );
  NAND U6260 ( .A(B[39]), .B(A[1]), .Z(n6082) );
  NAND U6261 ( .A(n6186), .B(n6187), .Z(n166) );
  NANDN U6262 ( .A(n6188), .B(n6189), .Z(n6187) );
  OR U6263 ( .A(n6190), .B(n6191), .Z(n6189) );
  NAND U6264 ( .A(n6191), .B(n6190), .Z(n6186) );
  XOR U6265 ( .A(n168), .B(n167), .Z(\A1[37] ) );
  XOR U6266 ( .A(n6191), .B(n6192), .Z(n167) );
  XNOR U6267 ( .A(n6190), .B(n6188), .Z(n6192) );
  AND U6268 ( .A(n6193), .B(n6194), .Z(n6188) );
  NANDN U6269 ( .A(n6195), .B(n6196), .Z(n6194) );
  NANDN U6270 ( .A(n6197), .B(n6198), .Z(n6196) );
  NANDN U6271 ( .A(n6198), .B(n6197), .Z(n6193) );
  ANDN U6272 ( .B(B[24]), .A(n29), .Z(n6190) );
  XNOR U6273 ( .A(n6097), .B(n6199), .Z(n6191) );
  XNOR U6274 ( .A(n6096), .B(n6094), .Z(n6199) );
  AND U6275 ( .A(n6200), .B(n6201), .Z(n6094) );
  NANDN U6276 ( .A(n6202), .B(n6203), .Z(n6201) );
  OR U6277 ( .A(n6204), .B(n6205), .Z(n6203) );
  NAND U6278 ( .A(n6205), .B(n6204), .Z(n6200) );
  ANDN U6279 ( .B(B[25]), .A(n30), .Z(n6096) );
  XNOR U6280 ( .A(n6104), .B(n6206), .Z(n6097) );
  XNOR U6281 ( .A(n6103), .B(n6101), .Z(n6206) );
  AND U6282 ( .A(n6207), .B(n6208), .Z(n6101) );
  NANDN U6283 ( .A(n6209), .B(n6210), .Z(n6208) );
  NANDN U6284 ( .A(n6211), .B(n6212), .Z(n6210) );
  NANDN U6285 ( .A(n6212), .B(n6211), .Z(n6207) );
  ANDN U6286 ( .B(B[26]), .A(n31), .Z(n6103) );
  XNOR U6287 ( .A(n6111), .B(n6213), .Z(n6104) );
  XNOR U6288 ( .A(n6110), .B(n6108), .Z(n6213) );
  AND U6289 ( .A(n6214), .B(n6215), .Z(n6108) );
  NANDN U6290 ( .A(n6216), .B(n6217), .Z(n6215) );
  OR U6291 ( .A(n6218), .B(n6219), .Z(n6217) );
  NAND U6292 ( .A(n6219), .B(n6218), .Z(n6214) );
  ANDN U6293 ( .B(B[27]), .A(n32), .Z(n6110) );
  XNOR U6294 ( .A(n6118), .B(n6220), .Z(n6111) );
  XNOR U6295 ( .A(n6117), .B(n6115), .Z(n6220) );
  AND U6296 ( .A(n6221), .B(n6222), .Z(n6115) );
  NANDN U6297 ( .A(n6223), .B(n6224), .Z(n6222) );
  NANDN U6298 ( .A(n6225), .B(n6226), .Z(n6224) );
  NANDN U6299 ( .A(n6226), .B(n6225), .Z(n6221) );
  ANDN U6300 ( .B(B[28]), .A(n33), .Z(n6117) );
  XNOR U6301 ( .A(n6125), .B(n6227), .Z(n6118) );
  XNOR U6302 ( .A(n6124), .B(n6122), .Z(n6227) );
  AND U6303 ( .A(n6228), .B(n6229), .Z(n6122) );
  NANDN U6304 ( .A(n6230), .B(n6231), .Z(n6229) );
  OR U6305 ( .A(n6232), .B(n6233), .Z(n6231) );
  NAND U6306 ( .A(n6233), .B(n6232), .Z(n6228) );
  ANDN U6307 ( .B(B[29]), .A(n34), .Z(n6124) );
  XNOR U6308 ( .A(n6132), .B(n6234), .Z(n6125) );
  XNOR U6309 ( .A(n6131), .B(n6129), .Z(n6234) );
  AND U6310 ( .A(n6235), .B(n6236), .Z(n6129) );
  NANDN U6311 ( .A(n6237), .B(n6238), .Z(n6236) );
  NANDN U6312 ( .A(n6239), .B(n6240), .Z(n6238) );
  NANDN U6313 ( .A(n6240), .B(n6239), .Z(n6235) );
  ANDN U6314 ( .B(B[30]), .A(n35), .Z(n6131) );
  XNOR U6315 ( .A(n6139), .B(n6241), .Z(n6132) );
  XNOR U6316 ( .A(n6138), .B(n6136), .Z(n6241) );
  AND U6317 ( .A(n6242), .B(n6243), .Z(n6136) );
  NANDN U6318 ( .A(n6244), .B(n6245), .Z(n6243) );
  OR U6319 ( .A(n6246), .B(n6247), .Z(n6245) );
  NAND U6320 ( .A(n6247), .B(n6246), .Z(n6242) );
  ANDN U6321 ( .B(B[31]), .A(n36), .Z(n6138) );
  XNOR U6322 ( .A(n6146), .B(n6248), .Z(n6139) );
  XNOR U6323 ( .A(n6145), .B(n6143), .Z(n6248) );
  AND U6324 ( .A(n6249), .B(n6250), .Z(n6143) );
  NANDN U6325 ( .A(n6251), .B(n6252), .Z(n6250) );
  NANDN U6326 ( .A(n6253), .B(n6254), .Z(n6252) );
  NANDN U6327 ( .A(n6254), .B(n6253), .Z(n6249) );
  ANDN U6328 ( .B(B[32]), .A(n37), .Z(n6145) );
  XNOR U6329 ( .A(n6153), .B(n6255), .Z(n6146) );
  XNOR U6330 ( .A(n6152), .B(n6150), .Z(n6255) );
  AND U6331 ( .A(n6256), .B(n6257), .Z(n6150) );
  NANDN U6332 ( .A(n6258), .B(n6259), .Z(n6257) );
  OR U6333 ( .A(n6260), .B(n6261), .Z(n6259) );
  NAND U6334 ( .A(n6261), .B(n6260), .Z(n6256) );
  ANDN U6335 ( .B(B[33]), .A(n38), .Z(n6152) );
  XNOR U6336 ( .A(n6160), .B(n6262), .Z(n6153) );
  XNOR U6337 ( .A(n6159), .B(n6157), .Z(n6262) );
  AND U6338 ( .A(n6263), .B(n6264), .Z(n6157) );
  NANDN U6339 ( .A(n6265), .B(n6266), .Z(n6264) );
  NANDN U6340 ( .A(n6267), .B(n6268), .Z(n6266) );
  NANDN U6341 ( .A(n6268), .B(n6267), .Z(n6263) );
  ANDN U6342 ( .B(B[34]), .A(n39), .Z(n6159) );
  XNOR U6343 ( .A(n6167), .B(n6269), .Z(n6160) );
  XNOR U6344 ( .A(n6166), .B(n6164), .Z(n6269) );
  AND U6345 ( .A(n6270), .B(n6271), .Z(n6164) );
  NANDN U6346 ( .A(n6272), .B(n6273), .Z(n6271) );
  OR U6347 ( .A(n6274), .B(n6275), .Z(n6273) );
  NAND U6348 ( .A(n6275), .B(n6274), .Z(n6270) );
  ANDN U6349 ( .B(B[35]), .A(n40), .Z(n6166) );
  XNOR U6350 ( .A(n6174), .B(n6276), .Z(n6167) );
  XNOR U6351 ( .A(n6173), .B(n6171), .Z(n6276) );
  AND U6352 ( .A(n6277), .B(n6278), .Z(n6171) );
  NANDN U6353 ( .A(n6279), .B(n6280), .Z(n6278) );
  NAND U6354 ( .A(n6281), .B(n6282), .Z(n6280) );
  ANDN U6355 ( .B(B[36]), .A(n41), .Z(n6173) );
  XOR U6356 ( .A(n6180), .B(n6283), .Z(n6174) );
  XNOR U6357 ( .A(n6178), .B(n6181), .Z(n6283) );
  NAND U6358 ( .A(A[2]), .B(B[37]), .Z(n6181) );
  NANDN U6359 ( .A(n6284), .B(n6285), .Z(n6178) );
  AND U6360 ( .A(A[0]), .B(B[38]), .Z(n6285) );
  XNOR U6361 ( .A(n6183), .B(n6286), .Z(n6180) );
  NAND U6362 ( .A(A[0]), .B(B[39]), .Z(n6286) );
  NAND U6363 ( .A(B[38]), .B(A[1]), .Z(n6183) );
  NAND U6364 ( .A(n6287), .B(n6288), .Z(n168) );
  NANDN U6365 ( .A(n6289), .B(n6290), .Z(n6288) );
  OR U6366 ( .A(n6291), .B(n6292), .Z(n6290) );
  NAND U6367 ( .A(n6292), .B(n6291), .Z(n6287) );
  XOR U6368 ( .A(n170), .B(n169), .Z(\A1[36] ) );
  XOR U6369 ( .A(n6292), .B(n6293), .Z(n169) );
  XNOR U6370 ( .A(n6291), .B(n6289), .Z(n6293) );
  AND U6371 ( .A(n6294), .B(n6295), .Z(n6289) );
  NANDN U6372 ( .A(n6296), .B(n6297), .Z(n6295) );
  NANDN U6373 ( .A(n6298), .B(n6299), .Z(n6297) );
  NANDN U6374 ( .A(n6299), .B(n6298), .Z(n6294) );
  ANDN U6375 ( .B(B[23]), .A(n29), .Z(n6291) );
  XNOR U6376 ( .A(n6198), .B(n6300), .Z(n6292) );
  XNOR U6377 ( .A(n6197), .B(n6195), .Z(n6300) );
  AND U6378 ( .A(n6301), .B(n6302), .Z(n6195) );
  NANDN U6379 ( .A(n6303), .B(n6304), .Z(n6302) );
  OR U6380 ( .A(n6305), .B(n6306), .Z(n6304) );
  NAND U6381 ( .A(n6306), .B(n6305), .Z(n6301) );
  ANDN U6382 ( .B(B[24]), .A(n30), .Z(n6197) );
  XNOR U6383 ( .A(n6205), .B(n6307), .Z(n6198) );
  XNOR U6384 ( .A(n6204), .B(n6202), .Z(n6307) );
  AND U6385 ( .A(n6308), .B(n6309), .Z(n6202) );
  NANDN U6386 ( .A(n6310), .B(n6311), .Z(n6309) );
  NANDN U6387 ( .A(n6312), .B(n6313), .Z(n6311) );
  NANDN U6388 ( .A(n6313), .B(n6312), .Z(n6308) );
  ANDN U6389 ( .B(B[25]), .A(n31), .Z(n6204) );
  XNOR U6390 ( .A(n6212), .B(n6314), .Z(n6205) );
  XNOR U6391 ( .A(n6211), .B(n6209), .Z(n6314) );
  AND U6392 ( .A(n6315), .B(n6316), .Z(n6209) );
  NANDN U6393 ( .A(n6317), .B(n6318), .Z(n6316) );
  OR U6394 ( .A(n6319), .B(n6320), .Z(n6318) );
  NAND U6395 ( .A(n6320), .B(n6319), .Z(n6315) );
  ANDN U6396 ( .B(B[26]), .A(n32), .Z(n6211) );
  XNOR U6397 ( .A(n6219), .B(n6321), .Z(n6212) );
  XNOR U6398 ( .A(n6218), .B(n6216), .Z(n6321) );
  AND U6399 ( .A(n6322), .B(n6323), .Z(n6216) );
  NANDN U6400 ( .A(n6324), .B(n6325), .Z(n6323) );
  NANDN U6401 ( .A(n6326), .B(n6327), .Z(n6325) );
  NANDN U6402 ( .A(n6327), .B(n6326), .Z(n6322) );
  ANDN U6403 ( .B(B[27]), .A(n33), .Z(n6218) );
  XNOR U6404 ( .A(n6226), .B(n6328), .Z(n6219) );
  XNOR U6405 ( .A(n6225), .B(n6223), .Z(n6328) );
  AND U6406 ( .A(n6329), .B(n6330), .Z(n6223) );
  NANDN U6407 ( .A(n6331), .B(n6332), .Z(n6330) );
  OR U6408 ( .A(n6333), .B(n6334), .Z(n6332) );
  NAND U6409 ( .A(n6334), .B(n6333), .Z(n6329) );
  ANDN U6410 ( .B(B[28]), .A(n34), .Z(n6225) );
  XNOR U6411 ( .A(n6233), .B(n6335), .Z(n6226) );
  XNOR U6412 ( .A(n6232), .B(n6230), .Z(n6335) );
  AND U6413 ( .A(n6336), .B(n6337), .Z(n6230) );
  NANDN U6414 ( .A(n6338), .B(n6339), .Z(n6337) );
  NANDN U6415 ( .A(n6340), .B(n6341), .Z(n6339) );
  NANDN U6416 ( .A(n6341), .B(n6340), .Z(n6336) );
  ANDN U6417 ( .B(B[29]), .A(n35), .Z(n6232) );
  XNOR U6418 ( .A(n6240), .B(n6342), .Z(n6233) );
  XNOR U6419 ( .A(n6239), .B(n6237), .Z(n6342) );
  AND U6420 ( .A(n6343), .B(n6344), .Z(n6237) );
  NANDN U6421 ( .A(n6345), .B(n6346), .Z(n6344) );
  OR U6422 ( .A(n6347), .B(n6348), .Z(n6346) );
  NAND U6423 ( .A(n6348), .B(n6347), .Z(n6343) );
  ANDN U6424 ( .B(B[30]), .A(n36), .Z(n6239) );
  XNOR U6425 ( .A(n6247), .B(n6349), .Z(n6240) );
  XNOR U6426 ( .A(n6246), .B(n6244), .Z(n6349) );
  AND U6427 ( .A(n6350), .B(n6351), .Z(n6244) );
  NANDN U6428 ( .A(n6352), .B(n6353), .Z(n6351) );
  NANDN U6429 ( .A(n6354), .B(n6355), .Z(n6353) );
  NANDN U6430 ( .A(n6355), .B(n6354), .Z(n6350) );
  ANDN U6431 ( .B(B[31]), .A(n37), .Z(n6246) );
  XNOR U6432 ( .A(n6254), .B(n6356), .Z(n6247) );
  XNOR U6433 ( .A(n6253), .B(n6251), .Z(n6356) );
  AND U6434 ( .A(n6357), .B(n6358), .Z(n6251) );
  NANDN U6435 ( .A(n6359), .B(n6360), .Z(n6358) );
  OR U6436 ( .A(n6361), .B(n6362), .Z(n6360) );
  NAND U6437 ( .A(n6362), .B(n6361), .Z(n6357) );
  ANDN U6438 ( .B(B[32]), .A(n38), .Z(n6253) );
  XNOR U6439 ( .A(n6261), .B(n6363), .Z(n6254) );
  XNOR U6440 ( .A(n6260), .B(n6258), .Z(n6363) );
  AND U6441 ( .A(n6364), .B(n6365), .Z(n6258) );
  NANDN U6442 ( .A(n6366), .B(n6367), .Z(n6365) );
  NANDN U6443 ( .A(n6368), .B(n6369), .Z(n6367) );
  NANDN U6444 ( .A(n6369), .B(n6368), .Z(n6364) );
  ANDN U6445 ( .B(B[33]), .A(n39), .Z(n6260) );
  XNOR U6446 ( .A(n6268), .B(n6370), .Z(n6261) );
  XNOR U6447 ( .A(n6267), .B(n6265), .Z(n6370) );
  AND U6448 ( .A(n6371), .B(n6372), .Z(n6265) );
  NANDN U6449 ( .A(n6373), .B(n6374), .Z(n6372) );
  OR U6450 ( .A(n6375), .B(n6376), .Z(n6374) );
  NAND U6451 ( .A(n6376), .B(n6375), .Z(n6371) );
  ANDN U6452 ( .B(B[34]), .A(n40), .Z(n6267) );
  XNOR U6453 ( .A(n6275), .B(n6377), .Z(n6268) );
  XNOR U6454 ( .A(n6274), .B(n6272), .Z(n6377) );
  AND U6455 ( .A(n6378), .B(n6379), .Z(n6272) );
  NANDN U6456 ( .A(n6380), .B(n6381), .Z(n6379) );
  NAND U6457 ( .A(n6382), .B(n6383), .Z(n6381) );
  ANDN U6458 ( .B(B[35]), .A(n41), .Z(n6274) );
  XOR U6459 ( .A(n6281), .B(n6384), .Z(n6275) );
  XNOR U6460 ( .A(n6279), .B(n6282), .Z(n6384) );
  NAND U6461 ( .A(A[2]), .B(B[36]), .Z(n6282) );
  NANDN U6462 ( .A(n6385), .B(n6386), .Z(n6279) );
  AND U6463 ( .A(A[0]), .B(B[37]), .Z(n6386) );
  XNOR U6464 ( .A(n6284), .B(n6387), .Z(n6281) );
  NAND U6465 ( .A(A[0]), .B(B[38]), .Z(n6387) );
  NAND U6466 ( .A(B[37]), .B(A[1]), .Z(n6284) );
  NAND U6467 ( .A(n6388), .B(n6389), .Z(n170) );
  NANDN U6468 ( .A(n6390), .B(n6391), .Z(n6389) );
  OR U6469 ( .A(n6392), .B(n6393), .Z(n6391) );
  NAND U6470 ( .A(n6393), .B(n6392), .Z(n6388) );
  XOR U6471 ( .A(n172), .B(n171), .Z(\A1[35] ) );
  XOR U6472 ( .A(n6393), .B(n6394), .Z(n171) );
  XNOR U6473 ( .A(n6392), .B(n6390), .Z(n6394) );
  AND U6474 ( .A(n6395), .B(n6396), .Z(n6390) );
  NANDN U6475 ( .A(n6397), .B(n6398), .Z(n6396) );
  NANDN U6476 ( .A(n6399), .B(n6400), .Z(n6398) );
  NANDN U6477 ( .A(n6400), .B(n6399), .Z(n6395) );
  ANDN U6478 ( .B(B[22]), .A(n29), .Z(n6392) );
  XNOR U6479 ( .A(n6299), .B(n6401), .Z(n6393) );
  XNOR U6480 ( .A(n6298), .B(n6296), .Z(n6401) );
  AND U6481 ( .A(n6402), .B(n6403), .Z(n6296) );
  NANDN U6482 ( .A(n6404), .B(n6405), .Z(n6403) );
  OR U6483 ( .A(n6406), .B(n6407), .Z(n6405) );
  NAND U6484 ( .A(n6407), .B(n6406), .Z(n6402) );
  ANDN U6485 ( .B(B[23]), .A(n30), .Z(n6298) );
  XNOR U6486 ( .A(n6306), .B(n6408), .Z(n6299) );
  XNOR U6487 ( .A(n6305), .B(n6303), .Z(n6408) );
  AND U6488 ( .A(n6409), .B(n6410), .Z(n6303) );
  NANDN U6489 ( .A(n6411), .B(n6412), .Z(n6410) );
  NANDN U6490 ( .A(n6413), .B(n6414), .Z(n6412) );
  NANDN U6491 ( .A(n6414), .B(n6413), .Z(n6409) );
  ANDN U6492 ( .B(B[24]), .A(n31), .Z(n6305) );
  XNOR U6493 ( .A(n6313), .B(n6415), .Z(n6306) );
  XNOR U6494 ( .A(n6312), .B(n6310), .Z(n6415) );
  AND U6495 ( .A(n6416), .B(n6417), .Z(n6310) );
  NANDN U6496 ( .A(n6418), .B(n6419), .Z(n6417) );
  OR U6497 ( .A(n6420), .B(n6421), .Z(n6419) );
  NAND U6498 ( .A(n6421), .B(n6420), .Z(n6416) );
  ANDN U6499 ( .B(B[25]), .A(n32), .Z(n6312) );
  XNOR U6500 ( .A(n6320), .B(n6422), .Z(n6313) );
  XNOR U6501 ( .A(n6319), .B(n6317), .Z(n6422) );
  AND U6502 ( .A(n6423), .B(n6424), .Z(n6317) );
  NANDN U6503 ( .A(n6425), .B(n6426), .Z(n6424) );
  NANDN U6504 ( .A(n6427), .B(n6428), .Z(n6426) );
  NANDN U6505 ( .A(n6428), .B(n6427), .Z(n6423) );
  ANDN U6506 ( .B(B[26]), .A(n33), .Z(n6319) );
  XNOR U6507 ( .A(n6327), .B(n6429), .Z(n6320) );
  XNOR U6508 ( .A(n6326), .B(n6324), .Z(n6429) );
  AND U6509 ( .A(n6430), .B(n6431), .Z(n6324) );
  NANDN U6510 ( .A(n6432), .B(n6433), .Z(n6431) );
  OR U6511 ( .A(n6434), .B(n6435), .Z(n6433) );
  NAND U6512 ( .A(n6435), .B(n6434), .Z(n6430) );
  ANDN U6513 ( .B(B[27]), .A(n34), .Z(n6326) );
  XNOR U6514 ( .A(n6334), .B(n6436), .Z(n6327) );
  XNOR U6515 ( .A(n6333), .B(n6331), .Z(n6436) );
  AND U6516 ( .A(n6437), .B(n6438), .Z(n6331) );
  NANDN U6517 ( .A(n6439), .B(n6440), .Z(n6438) );
  NANDN U6518 ( .A(n6441), .B(n6442), .Z(n6440) );
  NANDN U6519 ( .A(n6442), .B(n6441), .Z(n6437) );
  ANDN U6520 ( .B(B[28]), .A(n35), .Z(n6333) );
  XNOR U6521 ( .A(n6341), .B(n6443), .Z(n6334) );
  XNOR U6522 ( .A(n6340), .B(n6338), .Z(n6443) );
  AND U6523 ( .A(n6444), .B(n6445), .Z(n6338) );
  NANDN U6524 ( .A(n6446), .B(n6447), .Z(n6445) );
  OR U6525 ( .A(n6448), .B(n6449), .Z(n6447) );
  NAND U6526 ( .A(n6449), .B(n6448), .Z(n6444) );
  ANDN U6527 ( .B(B[29]), .A(n36), .Z(n6340) );
  XNOR U6528 ( .A(n6348), .B(n6450), .Z(n6341) );
  XNOR U6529 ( .A(n6347), .B(n6345), .Z(n6450) );
  AND U6530 ( .A(n6451), .B(n6452), .Z(n6345) );
  NANDN U6531 ( .A(n6453), .B(n6454), .Z(n6452) );
  NANDN U6532 ( .A(n6455), .B(n6456), .Z(n6454) );
  NANDN U6533 ( .A(n6456), .B(n6455), .Z(n6451) );
  ANDN U6534 ( .B(B[30]), .A(n37), .Z(n6347) );
  XNOR U6535 ( .A(n6355), .B(n6457), .Z(n6348) );
  XNOR U6536 ( .A(n6354), .B(n6352), .Z(n6457) );
  AND U6537 ( .A(n6458), .B(n6459), .Z(n6352) );
  NANDN U6538 ( .A(n6460), .B(n6461), .Z(n6459) );
  OR U6539 ( .A(n6462), .B(n6463), .Z(n6461) );
  NAND U6540 ( .A(n6463), .B(n6462), .Z(n6458) );
  ANDN U6541 ( .B(B[31]), .A(n38), .Z(n6354) );
  XNOR U6542 ( .A(n6362), .B(n6464), .Z(n6355) );
  XNOR U6543 ( .A(n6361), .B(n6359), .Z(n6464) );
  AND U6544 ( .A(n6465), .B(n6466), .Z(n6359) );
  NANDN U6545 ( .A(n6467), .B(n6468), .Z(n6466) );
  NANDN U6546 ( .A(n6469), .B(n6470), .Z(n6468) );
  NANDN U6547 ( .A(n6470), .B(n6469), .Z(n6465) );
  ANDN U6548 ( .B(B[32]), .A(n39), .Z(n6361) );
  XNOR U6549 ( .A(n6369), .B(n6471), .Z(n6362) );
  XNOR U6550 ( .A(n6368), .B(n6366), .Z(n6471) );
  AND U6551 ( .A(n6472), .B(n6473), .Z(n6366) );
  NANDN U6552 ( .A(n6474), .B(n6475), .Z(n6473) );
  OR U6553 ( .A(n6476), .B(n6477), .Z(n6475) );
  NAND U6554 ( .A(n6477), .B(n6476), .Z(n6472) );
  ANDN U6555 ( .B(B[33]), .A(n40), .Z(n6368) );
  XNOR U6556 ( .A(n6376), .B(n6478), .Z(n6369) );
  XNOR U6557 ( .A(n6375), .B(n6373), .Z(n6478) );
  AND U6558 ( .A(n6479), .B(n6480), .Z(n6373) );
  NANDN U6559 ( .A(n6481), .B(n6482), .Z(n6480) );
  NAND U6560 ( .A(n6483), .B(n6484), .Z(n6482) );
  ANDN U6561 ( .B(B[34]), .A(n41), .Z(n6375) );
  XOR U6562 ( .A(n6382), .B(n6485), .Z(n6376) );
  XNOR U6563 ( .A(n6380), .B(n6383), .Z(n6485) );
  NAND U6564 ( .A(A[2]), .B(B[35]), .Z(n6383) );
  NANDN U6565 ( .A(n6486), .B(n6487), .Z(n6380) );
  AND U6566 ( .A(A[0]), .B(B[36]), .Z(n6487) );
  XNOR U6567 ( .A(n6385), .B(n6488), .Z(n6382) );
  NAND U6568 ( .A(A[0]), .B(B[37]), .Z(n6488) );
  NAND U6569 ( .A(B[36]), .B(A[1]), .Z(n6385) );
  NAND U6570 ( .A(n6489), .B(n6490), .Z(n172) );
  NANDN U6571 ( .A(n6491), .B(n6492), .Z(n6490) );
  OR U6572 ( .A(n6493), .B(n6494), .Z(n6492) );
  NAND U6573 ( .A(n6494), .B(n6493), .Z(n6489) );
  XOR U6574 ( .A(n174), .B(n173), .Z(\A1[34] ) );
  XOR U6575 ( .A(n6494), .B(n6495), .Z(n173) );
  XNOR U6576 ( .A(n6493), .B(n6491), .Z(n6495) );
  AND U6577 ( .A(n6496), .B(n6497), .Z(n6491) );
  NANDN U6578 ( .A(n6498), .B(n6499), .Z(n6497) );
  NANDN U6579 ( .A(n6500), .B(n6501), .Z(n6499) );
  NANDN U6580 ( .A(n6501), .B(n6500), .Z(n6496) );
  ANDN U6581 ( .B(B[21]), .A(n29), .Z(n6493) );
  XNOR U6582 ( .A(n6400), .B(n6502), .Z(n6494) );
  XNOR U6583 ( .A(n6399), .B(n6397), .Z(n6502) );
  AND U6584 ( .A(n6503), .B(n6504), .Z(n6397) );
  NANDN U6585 ( .A(n6505), .B(n6506), .Z(n6504) );
  OR U6586 ( .A(n6507), .B(n6508), .Z(n6506) );
  NAND U6587 ( .A(n6508), .B(n6507), .Z(n6503) );
  ANDN U6588 ( .B(B[22]), .A(n30), .Z(n6399) );
  XNOR U6589 ( .A(n6407), .B(n6509), .Z(n6400) );
  XNOR U6590 ( .A(n6406), .B(n6404), .Z(n6509) );
  AND U6591 ( .A(n6510), .B(n6511), .Z(n6404) );
  NANDN U6592 ( .A(n6512), .B(n6513), .Z(n6511) );
  NANDN U6593 ( .A(n6514), .B(n6515), .Z(n6513) );
  NANDN U6594 ( .A(n6515), .B(n6514), .Z(n6510) );
  ANDN U6595 ( .B(B[23]), .A(n31), .Z(n6406) );
  XNOR U6596 ( .A(n6414), .B(n6516), .Z(n6407) );
  XNOR U6597 ( .A(n6413), .B(n6411), .Z(n6516) );
  AND U6598 ( .A(n6517), .B(n6518), .Z(n6411) );
  NANDN U6599 ( .A(n6519), .B(n6520), .Z(n6518) );
  OR U6600 ( .A(n6521), .B(n6522), .Z(n6520) );
  NAND U6601 ( .A(n6522), .B(n6521), .Z(n6517) );
  ANDN U6602 ( .B(B[24]), .A(n32), .Z(n6413) );
  XNOR U6603 ( .A(n6421), .B(n6523), .Z(n6414) );
  XNOR U6604 ( .A(n6420), .B(n6418), .Z(n6523) );
  AND U6605 ( .A(n6524), .B(n6525), .Z(n6418) );
  NANDN U6606 ( .A(n6526), .B(n6527), .Z(n6525) );
  NANDN U6607 ( .A(n6528), .B(n6529), .Z(n6527) );
  NANDN U6608 ( .A(n6529), .B(n6528), .Z(n6524) );
  ANDN U6609 ( .B(B[25]), .A(n33), .Z(n6420) );
  XNOR U6610 ( .A(n6428), .B(n6530), .Z(n6421) );
  XNOR U6611 ( .A(n6427), .B(n6425), .Z(n6530) );
  AND U6612 ( .A(n6531), .B(n6532), .Z(n6425) );
  NANDN U6613 ( .A(n6533), .B(n6534), .Z(n6532) );
  OR U6614 ( .A(n6535), .B(n6536), .Z(n6534) );
  NAND U6615 ( .A(n6536), .B(n6535), .Z(n6531) );
  ANDN U6616 ( .B(B[26]), .A(n34), .Z(n6427) );
  XNOR U6617 ( .A(n6435), .B(n6537), .Z(n6428) );
  XNOR U6618 ( .A(n6434), .B(n6432), .Z(n6537) );
  AND U6619 ( .A(n6538), .B(n6539), .Z(n6432) );
  NANDN U6620 ( .A(n6540), .B(n6541), .Z(n6539) );
  NANDN U6621 ( .A(n6542), .B(n6543), .Z(n6541) );
  NANDN U6622 ( .A(n6543), .B(n6542), .Z(n6538) );
  ANDN U6623 ( .B(B[27]), .A(n35), .Z(n6434) );
  XNOR U6624 ( .A(n6442), .B(n6544), .Z(n6435) );
  XNOR U6625 ( .A(n6441), .B(n6439), .Z(n6544) );
  AND U6626 ( .A(n6545), .B(n6546), .Z(n6439) );
  NANDN U6627 ( .A(n6547), .B(n6548), .Z(n6546) );
  OR U6628 ( .A(n6549), .B(n6550), .Z(n6548) );
  NAND U6629 ( .A(n6550), .B(n6549), .Z(n6545) );
  ANDN U6630 ( .B(B[28]), .A(n36), .Z(n6441) );
  XNOR U6631 ( .A(n6449), .B(n6551), .Z(n6442) );
  XNOR U6632 ( .A(n6448), .B(n6446), .Z(n6551) );
  AND U6633 ( .A(n6552), .B(n6553), .Z(n6446) );
  NANDN U6634 ( .A(n6554), .B(n6555), .Z(n6553) );
  NANDN U6635 ( .A(n6556), .B(n6557), .Z(n6555) );
  NANDN U6636 ( .A(n6557), .B(n6556), .Z(n6552) );
  ANDN U6637 ( .B(B[29]), .A(n37), .Z(n6448) );
  XNOR U6638 ( .A(n6456), .B(n6558), .Z(n6449) );
  XNOR U6639 ( .A(n6455), .B(n6453), .Z(n6558) );
  AND U6640 ( .A(n6559), .B(n6560), .Z(n6453) );
  NANDN U6641 ( .A(n6561), .B(n6562), .Z(n6560) );
  OR U6642 ( .A(n6563), .B(n6564), .Z(n6562) );
  NAND U6643 ( .A(n6564), .B(n6563), .Z(n6559) );
  ANDN U6644 ( .B(B[30]), .A(n38), .Z(n6455) );
  XNOR U6645 ( .A(n6463), .B(n6565), .Z(n6456) );
  XNOR U6646 ( .A(n6462), .B(n6460), .Z(n6565) );
  AND U6647 ( .A(n6566), .B(n6567), .Z(n6460) );
  NANDN U6648 ( .A(n6568), .B(n6569), .Z(n6567) );
  NANDN U6649 ( .A(n6570), .B(n6571), .Z(n6569) );
  NANDN U6650 ( .A(n6571), .B(n6570), .Z(n6566) );
  ANDN U6651 ( .B(B[31]), .A(n39), .Z(n6462) );
  XNOR U6652 ( .A(n6470), .B(n6572), .Z(n6463) );
  XNOR U6653 ( .A(n6469), .B(n6467), .Z(n6572) );
  AND U6654 ( .A(n6573), .B(n6574), .Z(n6467) );
  NANDN U6655 ( .A(n6575), .B(n6576), .Z(n6574) );
  OR U6656 ( .A(n6577), .B(n6578), .Z(n6576) );
  NAND U6657 ( .A(n6578), .B(n6577), .Z(n6573) );
  ANDN U6658 ( .B(B[32]), .A(n40), .Z(n6469) );
  XNOR U6659 ( .A(n6477), .B(n6579), .Z(n6470) );
  XNOR U6660 ( .A(n6476), .B(n6474), .Z(n6579) );
  AND U6661 ( .A(n6580), .B(n6581), .Z(n6474) );
  NANDN U6662 ( .A(n6582), .B(n6583), .Z(n6581) );
  NAND U6663 ( .A(n6584), .B(n6585), .Z(n6583) );
  ANDN U6664 ( .B(B[33]), .A(n41), .Z(n6476) );
  XOR U6665 ( .A(n6483), .B(n6586), .Z(n6477) );
  XNOR U6666 ( .A(n6481), .B(n6484), .Z(n6586) );
  NAND U6667 ( .A(A[2]), .B(B[34]), .Z(n6484) );
  NANDN U6668 ( .A(n6587), .B(n6588), .Z(n6481) );
  AND U6669 ( .A(A[0]), .B(B[35]), .Z(n6588) );
  XNOR U6670 ( .A(n6486), .B(n6589), .Z(n6483) );
  NAND U6671 ( .A(A[0]), .B(B[36]), .Z(n6589) );
  NAND U6672 ( .A(B[35]), .B(A[1]), .Z(n6486) );
  NAND U6673 ( .A(n6590), .B(n6591), .Z(n174) );
  NANDN U6674 ( .A(n6592), .B(n6593), .Z(n6591) );
  OR U6675 ( .A(n6594), .B(n6595), .Z(n6593) );
  NAND U6676 ( .A(n6595), .B(n6594), .Z(n6590) );
  XOR U6677 ( .A(n176), .B(n175), .Z(\A1[33] ) );
  XOR U6678 ( .A(n6595), .B(n6596), .Z(n175) );
  XNOR U6679 ( .A(n6594), .B(n6592), .Z(n6596) );
  AND U6680 ( .A(n6597), .B(n6598), .Z(n6592) );
  NANDN U6681 ( .A(n6599), .B(n6600), .Z(n6598) );
  NANDN U6682 ( .A(n6601), .B(n6602), .Z(n6600) );
  NANDN U6683 ( .A(n6602), .B(n6601), .Z(n6597) );
  ANDN U6684 ( .B(B[20]), .A(n29), .Z(n6594) );
  XNOR U6685 ( .A(n6501), .B(n6603), .Z(n6595) );
  XNOR U6686 ( .A(n6500), .B(n6498), .Z(n6603) );
  AND U6687 ( .A(n6604), .B(n6605), .Z(n6498) );
  NANDN U6688 ( .A(n6606), .B(n6607), .Z(n6605) );
  OR U6689 ( .A(n6608), .B(n6609), .Z(n6607) );
  NAND U6690 ( .A(n6609), .B(n6608), .Z(n6604) );
  ANDN U6691 ( .B(B[21]), .A(n30), .Z(n6500) );
  XNOR U6692 ( .A(n6508), .B(n6610), .Z(n6501) );
  XNOR U6693 ( .A(n6507), .B(n6505), .Z(n6610) );
  AND U6694 ( .A(n6611), .B(n6612), .Z(n6505) );
  NANDN U6695 ( .A(n6613), .B(n6614), .Z(n6612) );
  NANDN U6696 ( .A(n6615), .B(n6616), .Z(n6614) );
  NANDN U6697 ( .A(n6616), .B(n6615), .Z(n6611) );
  ANDN U6698 ( .B(B[22]), .A(n31), .Z(n6507) );
  XNOR U6699 ( .A(n6515), .B(n6617), .Z(n6508) );
  XNOR U6700 ( .A(n6514), .B(n6512), .Z(n6617) );
  AND U6701 ( .A(n6618), .B(n6619), .Z(n6512) );
  NANDN U6702 ( .A(n6620), .B(n6621), .Z(n6619) );
  OR U6703 ( .A(n6622), .B(n6623), .Z(n6621) );
  NAND U6704 ( .A(n6623), .B(n6622), .Z(n6618) );
  ANDN U6705 ( .B(B[23]), .A(n32), .Z(n6514) );
  XNOR U6706 ( .A(n6522), .B(n6624), .Z(n6515) );
  XNOR U6707 ( .A(n6521), .B(n6519), .Z(n6624) );
  AND U6708 ( .A(n6625), .B(n6626), .Z(n6519) );
  NANDN U6709 ( .A(n6627), .B(n6628), .Z(n6626) );
  NANDN U6710 ( .A(n6629), .B(n6630), .Z(n6628) );
  NANDN U6711 ( .A(n6630), .B(n6629), .Z(n6625) );
  ANDN U6712 ( .B(B[24]), .A(n33), .Z(n6521) );
  XNOR U6713 ( .A(n6529), .B(n6631), .Z(n6522) );
  XNOR U6714 ( .A(n6528), .B(n6526), .Z(n6631) );
  AND U6715 ( .A(n6632), .B(n6633), .Z(n6526) );
  NANDN U6716 ( .A(n6634), .B(n6635), .Z(n6633) );
  OR U6717 ( .A(n6636), .B(n6637), .Z(n6635) );
  NAND U6718 ( .A(n6637), .B(n6636), .Z(n6632) );
  ANDN U6719 ( .B(B[25]), .A(n34), .Z(n6528) );
  XNOR U6720 ( .A(n6536), .B(n6638), .Z(n6529) );
  XNOR U6721 ( .A(n6535), .B(n6533), .Z(n6638) );
  AND U6722 ( .A(n6639), .B(n6640), .Z(n6533) );
  NANDN U6723 ( .A(n6641), .B(n6642), .Z(n6640) );
  NANDN U6724 ( .A(n6643), .B(n6644), .Z(n6642) );
  NANDN U6725 ( .A(n6644), .B(n6643), .Z(n6639) );
  ANDN U6726 ( .B(B[26]), .A(n35), .Z(n6535) );
  XNOR U6727 ( .A(n6543), .B(n6645), .Z(n6536) );
  XNOR U6728 ( .A(n6542), .B(n6540), .Z(n6645) );
  AND U6729 ( .A(n6646), .B(n6647), .Z(n6540) );
  NANDN U6730 ( .A(n6648), .B(n6649), .Z(n6647) );
  OR U6731 ( .A(n6650), .B(n6651), .Z(n6649) );
  NAND U6732 ( .A(n6651), .B(n6650), .Z(n6646) );
  ANDN U6733 ( .B(B[27]), .A(n36), .Z(n6542) );
  XNOR U6734 ( .A(n6550), .B(n6652), .Z(n6543) );
  XNOR U6735 ( .A(n6549), .B(n6547), .Z(n6652) );
  AND U6736 ( .A(n6653), .B(n6654), .Z(n6547) );
  NANDN U6737 ( .A(n6655), .B(n6656), .Z(n6654) );
  NANDN U6738 ( .A(n6657), .B(n6658), .Z(n6656) );
  NANDN U6739 ( .A(n6658), .B(n6657), .Z(n6653) );
  ANDN U6740 ( .B(B[28]), .A(n37), .Z(n6549) );
  XNOR U6741 ( .A(n6557), .B(n6659), .Z(n6550) );
  XNOR U6742 ( .A(n6556), .B(n6554), .Z(n6659) );
  AND U6743 ( .A(n6660), .B(n6661), .Z(n6554) );
  NANDN U6744 ( .A(n6662), .B(n6663), .Z(n6661) );
  OR U6745 ( .A(n6664), .B(n6665), .Z(n6663) );
  NAND U6746 ( .A(n6665), .B(n6664), .Z(n6660) );
  ANDN U6747 ( .B(B[29]), .A(n38), .Z(n6556) );
  XNOR U6748 ( .A(n6564), .B(n6666), .Z(n6557) );
  XNOR U6749 ( .A(n6563), .B(n6561), .Z(n6666) );
  AND U6750 ( .A(n6667), .B(n6668), .Z(n6561) );
  NANDN U6751 ( .A(n6669), .B(n6670), .Z(n6668) );
  NANDN U6752 ( .A(n6671), .B(n6672), .Z(n6670) );
  NANDN U6753 ( .A(n6672), .B(n6671), .Z(n6667) );
  ANDN U6754 ( .B(B[30]), .A(n39), .Z(n6563) );
  XNOR U6755 ( .A(n6571), .B(n6673), .Z(n6564) );
  XNOR U6756 ( .A(n6570), .B(n6568), .Z(n6673) );
  AND U6757 ( .A(n6674), .B(n6675), .Z(n6568) );
  NANDN U6758 ( .A(n6676), .B(n6677), .Z(n6675) );
  OR U6759 ( .A(n6678), .B(n6679), .Z(n6677) );
  NAND U6760 ( .A(n6679), .B(n6678), .Z(n6674) );
  ANDN U6761 ( .B(B[31]), .A(n40), .Z(n6570) );
  XNOR U6762 ( .A(n6578), .B(n6680), .Z(n6571) );
  XNOR U6763 ( .A(n6577), .B(n6575), .Z(n6680) );
  AND U6764 ( .A(n6681), .B(n6682), .Z(n6575) );
  NANDN U6765 ( .A(n6683), .B(n6684), .Z(n6682) );
  NAND U6766 ( .A(n6685), .B(n6686), .Z(n6684) );
  ANDN U6767 ( .B(B[32]), .A(n41), .Z(n6577) );
  XOR U6768 ( .A(n6584), .B(n6687), .Z(n6578) );
  XNOR U6769 ( .A(n6582), .B(n6585), .Z(n6687) );
  NAND U6770 ( .A(A[2]), .B(B[33]), .Z(n6585) );
  NANDN U6771 ( .A(n6688), .B(n6689), .Z(n6582) );
  AND U6772 ( .A(A[0]), .B(B[34]), .Z(n6689) );
  XNOR U6773 ( .A(n6587), .B(n6690), .Z(n6584) );
  NAND U6774 ( .A(A[0]), .B(B[35]), .Z(n6690) );
  NAND U6775 ( .A(B[34]), .B(A[1]), .Z(n6587) );
  NAND U6776 ( .A(n6691), .B(n6692), .Z(n176) );
  NANDN U6777 ( .A(n6693), .B(n6694), .Z(n6692) );
  OR U6778 ( .A(n6695), .B(n6696), .Z(n6694) );
  NAND U6779 ( .A(n6696), .B(n6695), .Z(n6691) );
  XOR U6780 ( .A(n178), .B(n177), .Z(\A1[32] ) );
  XOR U6781 ( .A(n6696), .B(n6697), .Z(n177) );
  XNOR U6782 ( .A(n6695), .B(n6693), .Z(n6697) );
  AND U6783 ( .A(n6698), .B(n6699), .Z(n6693) );
  NANDN U6784 ( .A(n6700), .B(n6701), .Z(n6699) );
  NANDN U6785 ( .A(n6702), .B(n6703), .Z(n6701) );
  NANDN U6786 ( .A(n6703), .B(n6702), .Z(n6698) );
  ANDN U6787 ( .B(B[19]), .A(n29), .Z(n6695) );
  XNOR U6788 ( .A(n6602), .B(n6704), .Z(n6696) );
  XNOR U6789 ( .A(n6601), .B(n6599), .Z(n6704) );
  AND U6790 ( .A(n6705), .B(n6706), .Z(n6599) );
  NANDN U6791 ( .A(n6707), .B(n6708), .Z(n6706) );
  OR U6792 ( .A(n6709), .B(n6710), .Z(n6708) );
  NAND U6793 ( .A(n6710), .B(n6709), .Z(n6705) );
  ANDN U6794 ( .B(B[20]), .A(n30), .Z(n6601) );
  XNOR U6795 ( .A(n6609), .B(n6711), .Z(n6602) );
  XNOR U6796 ( .A(n6608), .B(n6606), .Z(n6711) );
  AND U6797 ( .A(n6712), .B(n6713), .Z(n6606) );
  NANDN U6798 ( .A(n6714), .B(n6715), .Z(n6713) );
  NANDN U6799 ( .A(n6716), .B(n6717), .Z(n6715) );
  NANDN U6800 ( .A(n6717), .B(n6716), .Z(n6712) );
  ANDN U6801 ( .B(B[21]), .A(n31), .Z(n6608) );
  XNOR U6802 ( .A(n6616), .B(n6718), .Z(n6609) );
  XNOR U6803 ( .A(n6615), .B(n6613), .Z(n6718) );
  AND U6804 ( .A(n6719), .B(n6720), .Z(n6613) );
  NANDN U6805 ( .A(n6721), .B(n6722), .Z(n6720) );
  OR U6806 ( .A(n6723), .B(n6724), .Z(n6722) );
  NAND U6807 ( .A(n6724), .B(n6723), .Z(n6719) );
  ANDN U6808 ( .B(B[22]), .A(n32), .Z(n6615) );
  XNOR U6809 ( .A(n6623), .B(n6725), .Z(n6616) );
  XNOR U6810 ( .A(n6622), .B(n6620), .Z(n6725) );
  AND U6811 ( .A(n6726), .B(n6727), .Z(n6620) );
  NANDN U6812 ( .A(n6728), .B(n6729), .Z(n6727) );
  NANDN U6813 ( .A(n6730), .B(n6731), .Z(n6729) );
  NANDN U6814 ( .A(n6731), .B(n6730), .Z(n6726) );
  ANDN U6815 ( .B(B[23]), .A(n33), .Z(n6622) );
  XNOR U6816 ( .A(n6630), .B(n6732), .Z(n6623) );
  XNOR U6817 ( .A(n6629), .B(n6627), .Z(n6732) );
  AND U6818 ( .A(n6733), .B(n6734), .Z(n6627) );
  NANDN U6819 ( .A(n6735), .B(n6736), .Z(n6734) );
  OR U6820 ( .A(n6737), .B(n6738), .Z(n6736) );
  NAND U6821 ( .A(n6738), .B(n6737), .Z(n6733) );
  ANDN U6822 ( .B(B[24]), .A(n34), .Z(n6629) );
  XNOR U6823 ( .A(n6637), .B(n6739), .Z(n6630) );
  XNOR U6824 ( .A(n6636), .B(n6634), .Z(n6739) );
  AND U6825 ( .A(n6740), .B(n6741), .Z(n6634) );
  NANDN U6826 ( .A(n6742), .B(n6743), .Z(n6741) );
  NANDN U6827 ( .A(n6744), .B(n6745), .Z(n6743) );
  NANDN U6828 ( .A(n6745), .B(n6744), .Z(n6740) );
  ANDN U6829 ( .B(B[25]), .A(n35), .Z(n6636) );
  XNOR U6830 ( .A(n6644), .B(n6746), .Z(n6637) );
  XNOR U6831 ( .A(n6643), .B(n6641), .Z(n6746) );
  AND U6832 ( .A(n6747), .B(n6748), .Z(n6641) );
  NANDN U6833 ( .A(n6749), .B(n6750), .Z(n6748) );
  OR U6834 ( .A(n6751), .B(n6752), .Z(n6750) );
  NAND U6835 ( .A(n6752), .B(n6751), .Z(n6747) );
  ANDN U6836 ( .B(B[26]), .A(n36), .Z(n6643) );
  XNOR U6837 ( .A(n6651), .B(n6753), .Z(n6644) );
  XNOR U6838 ( .A(n6650), .B(n6648), .Z(n6753) );
  AND U6839 ( .A(n6754), .B(n6755), .Z(n6648) );
  NANDN U6840 ( .A(n6756), .B(n6757), .Z(n6755) );
  NANDN U6841 ( .A(n6758), .B(n6759), .Z(n6757) );
  NANDN U6842 ( .A(n6759), .B(n6758), .Z(n6754) );
  ANDN U6843 ( .B(B[27]), .A(n37), .Z(n6650) );
  XNOR U6844 ( .A(n6658), .B(n6760), .Z(n6651) );
  XNOR U6845 ( .A(n6657), .B(n6655), .Z(n6760) );
  AND U6846 ( .A(n6761), .B(n6762), .Z(n6655) );
  NANDN U6847 ( .A(n6763), .B(n6764), .Z(n6762) );
  OR U6848 ( .A(n6765), .B(n6766), .Z(n6764) );
  NAND U6849 ( .A(n6766), .B(n6765), .Z(n6761) );
  ANDN U6850 ( .B(B[28]), .A(n38), .Z(n6657) );
  XNOR U6851 ( .A(n6665), .B(n6767), .Z(n6658) );
  XNOR U6852 ( .A(n6664), .B(n6662), .Z(n6767) );
  AND U6853 ( .A(n6768), .B(n6769), .Z(n6662) );
  NANDN U6854 ( .A(n6770), .B(n6771), .Z(n6769) );
  NANDN U6855 ( .A(n6772), .B(n6773), .Z(n6771) );
  NANDN U6856 ( .A(n6773), .B(n6772), .Z(n6768) );
  ANDN U6857 ( .B(B[29]), .A(n39), .Z(n6664) );
  XNOR U6858 ( .A(n6672), .B(n6774), .Z(n6665) );
  XNOR U6859 ( .A(n6671), .B(n6669), .Z(n6774) );
  AND U6860 ( .A(n6775), .B(n6776), .Z(n6669) );
  NANDN U6861 ( .A(n6777), .B(n6778), .Z(n6776) );
  OR U6862 ( .A(n6779), .B(n6780), .Z(n6778) );
  NAND U6863 ( .A(n6780), .B(n6779), .Z(n6775) );
  ANDN U6864 ( .B(B[30]), .A(n40), .Z(n6671) );
  XNOR U6865 ( .A(n6679), .B(n6781), .Z(n6672) );
  XNOR U6866 ( .A(n6678), .B(n6676), .Z(n6781) );
  AND U6867 ( .A(n6782), .B(n6783), .Z(n6676) );
  NANDN U6868 ( .A(n6784), .B(n6785), .Z(n6783) );
  NAND U6869 ( .A(n6786), .B(n6787), .Z(n6785) );
  ANDN U6870 ( .B(B[31]), .A(n41), .Z(n6678) );
  XOR U6871 ( .A(n6685), .B(n6788), .Z(n6679) );
  XNOR U6872 ( .A(n6683), .B(n6686), .Z(n6788) );
  NAND U6873 ( .A(A[2]), .B(B[32]), .Z(n6686) );
  NANDN U6874 ( .A(n6789), .B(n6790), .Z(n6683) );
  AND U6875 ( .A(A[0]), .B(B[33]), .Z(n6790) );
  XNOR U6876 ( .A(n6688), .B(n6791), .Z(n6685) );
  NAND U6877 ( .A(A[0]), .B(B[34]), .Z(n6791) );
  NAND U6878 ( .A(B[33]), .B(A[1]), .Z(n6688) );
  NAND U6879 ( .A(n6792), .B(n6793), .Z(n178) );
  NANDN U6880 ( .A(n6794), .B(n6795), .Z(n6793) );
  OR U6881 ( .A(n6796), .B(n6797), .Z(n6795) );
  NAND U6882 ( .A(n6797), .B(n6796), .Z(n6792) );
  XOR U6883 ( .A(n180), .B(n179), .Z(\A1[31] ) );
  XOR U6884 ( .A(n6797), .B(n6798), .Z(n179) );
  XNOR U6885 ( .A(n6796), .B(n6794), .Z(n6798) );
  AND U6886 ( .A(n6799), .B(n6800), .Z(n6794) );
  NANDN U6887 ( .A(n6801), .B(n6802), .Z(n6800) );
  NANDN U6888 ( .A(n6803), .B(n6804), .Z(n6802) );
  NANDN U6889 ( .A(n6804), .B(n6803), .Z(n6799) );
  ANDN U6890 ( .B(B[18]), .A(n29), .Z(n6796) );
  XNOR U6891 ( .A(n6703), .B(n6805), .Z(n6797) );
  XNOR U6892 ( .A(n6702), .B(n6700), .Z(n6805) );
  AND U6893 ( .A(n6806), .B(n6807), .Z(n6700) );
  NANDN U6894 ( .A(n6808), .B(n6809), .Z(n6807) );
  OR U6895 ( .A(n6810), .B(n6811), .Z(n6809) );
  NAND U6896 ( .A(n6811), .B(n6810), .Z(n6806) );
  ANDN U6897 ( .B(B[19]), .A(n30), .Z(n6702) );
  XNOR U6898 ( .A(n6710), .B(n6812), .Z(n6703) );
  XNOR U6899 ( .A(n6709), .B(n6707), .Z(n6812) );
  AND U6900 ( .A(n6813), .B(n6814), .Z(n6707) );
  NANDN U6901 ( .A(n6815), .B(n6816), .Z(n6814) );
  NANDN U6902 ( .A(n6817), .B(n6818), .Z(n6816) );
  NANDN U6903 ( .A(n6818), .B(n6817), .Z(n6813) );
  ANDN U6904 ( .B(B[20]), .A(n31), .Z(n6709) );
  XNOR U6905 ( .A(n6717), .B(n6819), .Z(n6710) );
  XNOR U6906 ( .A(n6716), .B(n6714), .Z(n6819) );
  AND U6907 ( .A(n6820), .B(n6821), .Z(n6714) );
  NANDN U6908 ( .A(n6822), .B(n6823), .Z(n6821) );
  OR U6909 ( .A(n6824), .B(n6825), .Z(n6823) );
  NAND U6910 ( .A(n6825), .B(n6824), .Z(n6820) );
  ANDN U6911 ( .B(B[21]), .A(n32), .Z(n6716) );
  XNOR U6912 ( .A(n6724), .B(n6826), .Z(n6717) );
  XNOR U6913 ( .A(n6723), .B(n6721), .Z(n6826) );
  AND U6914 ( .A(n6827), .B(n6828), .Z(n6721) );
  NANDN U6915 ( .A(n6829), .B(n6830), .Z(n6828) );
  NANDN U6916 ( .A(n6831), .B(n6832), .Z(n6830) );
  NANDN U6917 ( .A(n6832), .B(n6831), .Z(n6827) );
  ANDN U6918 ( .B(B[22]), .A(n33), .Z(n6723) );
  XNOR U6919 ( .A(n6731), .B(n6833), .Z(n6724) );
  XNOR U6920 ( .A(n6730), .B(n6728), .Z(n6833) );
  AND U6921 ( .A(n6834), .B(n6835), .Z(n6728) );
  NANDN U6922 ( .A(n6836), .B(n6837), .Z(n6835) );
  OR U6923 ( .A(n6838), .B(n6839), .Z(n6837) );
  NAND U6924 ( .A(n6839), .B(n6838), .Z(n6834) );
  ANDN U6925 ( .B(B[23]), .A(n34), .Z(n6730) );
  XNOR U6926 ( .A(n6738), .B(n6840), .Z(n6731) );
  XNOR U6927 ( .A(n6737), .B(n6735), .Z(n6840) );
  AND U6928 ( .A(n6841), .B(n6842), .Z(n6735) );
  NANDN U6929 ( .A(n6843), .B(n6844), .Z(n6842) );
  NANDN U6930 ( .A(n6845), .B(n6846), .Z(n6844) );
  NANDN U6931 ( .A(n6846), .B(n6845), .Z(n6841) );
  ANDN U6932 ( .B(B[24]), .A(n35), .Z(n6737) );
  XNOR U6933 ( .A(n6745), .B(n6847), .Z(n6738) );
  XNOR U6934 ( .A(n6744), .B(n6742), .Z(n6847) );
  AND U6935 ( .A(n6848), .B(n6849), .Z(n6742) );
  NANDN U6936 ( .A(n6850), .B(n6851), .Z(n6849) );
  OR U6937 ( .A(n6852), .B(n6853), .Z(n6851) );
  NAND U6938 ( .A(n6853), .B(n6852), .Z(n6848) );
  ANDN U6939 ( .B(B[25]), .A(n36), .Z(n6744) );
  XNOR U6940 ( .A(n6752), .B(n6854), .Z(n6745) );
  XNOR U6941 ( .A(n6751), .B(n6749), .Z(n6854) );
  AND U6942 ( .A(n6855), .B(n6856), .Z(n6749) );
  NANDN U6943 ( .A(n6857), .B(n6858), .Z(n6856) );
  NANDN U6944 ( .A(n6859), .B(n6860), .Z(n6858) );
  NANDN U6945 ( .A(n6860), .B(n6859), .Z(n6855) );
  ANDN U6946 ( .B(B[26]), .A(n37), .Z(n6751) );
  XNOR U6947 ( .A(n6759), .B(n6861), .Z(n6752) );
  XNOR U6948 ( .A(n6758), .B(n6756), .Z(n6861) );
  AND U6949 ( .A(n6862), .B(n6863), .Z(n6756) );
  NANDN U6950 ( .A(n6864), .B(n6865), .Z(n6863) );
  OR U6951 ( .A(n6866), .B(n6867), .Z(n6865) );
  NAND U6952 ( .A(n6867), .B(n6866), .Z(n6862) );
  ANDN U6953 ( .B(B[27]), .A(n38), .Z(n6758) );
  XNOR U6954 ( .A(n6766), .B(n6868), .Z(n6759) );
  XNOR U6955 ( .A(n6765), .B(n6763), .Z(n6868) );
  AND U6956 ( .A(n6869), .B(n6870), .Z(n6763) );
  NANDN U6957 ( .A(n6871), .B(n6872), .Z(n6870) );
  NANDN U6958 ( .A(n6873), .B(n6874), .Z(n6872) );
  NANDN U6959 ( .A(n6874), .B(n6873), .Z(n6869) );
  ANDN U6960 ( .B(B[28]), .A(n39), .Z(n6765) );
  XNOR U6961 ( .A(n6773), .B(n6875), .Z(n6766) );
  XNOR U6962 ( .A(n6772), .B(n6770), .Z(n6875) );
  AND U6963 ( .A(n6876), .B(n6877), .Z(n6770) );
  NANDN U6964 ( .A(n6878), .B(n6879), .Z(n6877) );
  OR U6965 ( .A(n6880), .B(n6881), .Z(n6879) );
  NAND U6966 ( .A(n6881), .B(n6880), .Z(n6876) );
  ANDN U6967 ( .B(B[29]), .A(n40), .Z(n6772) );
  XNOR U6968 ( .A(n6780), .B(n6882), .Z(n6773) );
  XNOR U6969 ( .A(n6779), .B(n6777), .Z(n6882) );
  AND U6970 ( .A(n6883), .B(n6884), .Z(n6777) );
  NANDN U6971 ( .A(n6885), .B(n6886), .Z(n6884) );
  NAND U6972 ( .A(n6887), .B(n6888), .Z(n6886) );
  ANDN U6973 ( .B(B[30]), .A(n41), .Z(n6779) );
  XOR U6974 ( .A(n6786), .B(n6889), .Z(n6780) );
  XNOR U6975 ( .A(n6784), .B(n6787), .Z(n6889) );
  NAND U6976 ( .A(A[2]), .B(B[31]), .Z(n6787) );
  NANDN U6977 ( .A(n6890), .B(n6891), .Z(n6784) );
  AND U6978 ( .A(A[0]), .B(B[32]), .Z(n6891) );
  XNOR U6979 ( .A(n6789), .B(n6892), .Z(n6786) );
  NAND U6980 ( .A(A[0]), .B(B[33]), .Z(n6892) );
  NAND U6981 ( .A(B[32]), .B(A[1]), .Z(n6789) );
  NAND U6982 ( .A(n6893), .B(n6894), .Z(n180) );
  NANDN U6983 ( .A(n6895), .B(n6896), .Z(n6894) );
  OR U6984 ( .A(n6897), .B(n6898), .Z(n6896) );
  NAND U6985 ( .A(n6898), .B(n6897), .Z(n6893) );
  XOR U6986 ( .A(n182), .B(n181), .Z(\A1[30] ) );
  XOR U6987 ( .A(n6898), .B(n6899), .Z(n181) );
  XNOR U6988 ( .A(n6897), .B(n6895), .Z(n6899) );
  AND U6989 ( .A(n6900), .B(n6901), .Z(n6895) );
  NANDN U6990 ( .A(n6902), .B(n6903), .Z(n6901) );
  NANDN U6991 ( .A(n6904), .B(n6905), .Z(n6903) );
  NANDN U6992 ( .A(n6905), .B(n6904), .Z(n6900) );
  ANDN U6993 ( .B(B[17]), .A(n29), .Z(n6897) );
  XNOR U6994 ( .A(n6804), .B(n6906), .Z(n6898) );
  XNOR U6995 ( .A(n6803), .B(n6801), .Z(n6906) );
  AND U6996 ( .A(n6907), .B(n6908), .Z(n6801) );
  NANDN U6997 ( .A(n6909), .B(n6910), .Z(n6908) );
  OR U6998 ( .A(n6911), .B(n6912), .Z(n6910) );
  NAND U6999 ( .A(n6912), .B(n6911), .Z(n6907) );
  ANDN U7000 ( .B(B[18]), .A(n30), .Z(n6803) );
  XNOR U7001 ( .A(n6811), .B(n6913), .Z(n6804) );
  XNOR U7002 ( .A(n6810), .B(n6808), .Z(n6913) );
  AND U7003 ( .A(n6914), .B(n6915), .Z(n6808) );
  NANDN U7004 ( .A(n6916), .B(n6917), .Z(n6915) );
  NANDN U7005 ( .A(n6918), .B(n6919), .Z(n6917) );
  NANDN U7006 ( .A(n6919), .B(n6918), .Z(n6914) );
  ANDN U7007 ( .B(B[19]), .A(n31), .Z(n6810) );
  XNOR U7008 ( .A(n6818), .B(n6920), .Z(n6811) );
  XNOR U7009 ( .A(n6817), .B(n6815), .Z(n6920) );
  AND U7010 ( .A(n6921), .B(n6922), .Z(n6815) );
  NANDN U7011 ( .A(n6923), .B(n6924), .Z(n6922) );
  OR U7012 ( .A(n6925), .B(n6926), .Z(n6924) );
  NAND U7013 ( .A(n6926), .B(n6925), .Z(n6921) );
  ANDN U7014 ( .B(B[20]), .A(n32), .Z(n6817) );
  XNOR U7015 ( .A(n6825), .B(n6927), .Z(n6818) );
  XNOR U7016 ( .A(n6824), .B(n6822), .Z(n6927) );
  AND U7017 ( .A(n6928), .B(n6929), .Z(n6822) );
  NANDN U7018 ( .A(n6930), .B(n6931), .Z(n6929) );
  NANDN U7019 ( .A(n6932), .B(n6933), .Z(n6931) );
  NANDN U7020 ( .A(n6933), .B(n6932), .Z(n6928) );
  ANDN U7021 ( .B(B[21]), .A(n33), .Z(n6824) );
  XNOR U7022 ( .A(n6832), .B(n6934), .Z(n6825) );
  XNOR U7023 ( .A(n6831), .B(n6829), .Z(n6934) );
  AND U7024 ( .A(n6935), .B(n6936), .Z(n6829) );
  NANDN U7025 ( .A(n6937), .B(n6938), .Z(n6936) );
  OR U7026 ( .A(n6939), .B(n6940), .Z(n6938) );
  NAND U7027 ( .A(n6940), .B(n6939), .Z(n6935) );
  ANDN U7028 ( .B(B[22]), .A(n34), .Z(n6831) );
  XNOR U7029 ( .A(n6839), .B(n6941), .Z(n6832) );
  XNOR U7030 ( .A(n6838), .B(n6836), .Z(n6941) );
  AND U7031 ( .A(n6942), .B(n6943), .Z(n6836) );
  NANDN U7032 ( .A(n6944), .B(n6945), .Z(n6943) );
  NANDN U7033 ( .A(n6946), .B(n6947), .Z(n6945) );
  NANDN U7034 ( .A(n6947), .B(n6946), .Z(n6942) );
  ANDN U7035 ( .B(B[23]), .A(n35), .Z(n6838) );
  XNOR U7036 ( .A(n6846), .B(n6948), .Z(n6839) );
  XNOR U7037 ( .A(n6845), .B(n6843), .Z(n6948) );
  AND U7038 ( .A(n6949), .B(n6950), .Z(n6843) );
  NANDN U7039 ( .A(n6951), .B(n6952), .Z(n6950) );
  OR U7040 ( .A(n6953), .B(n6954), .Z(n6952) );
  NAND U7041 ( .A(n6954), .B(n6953), .Z(n6949) );
  ANDN U7042 ( .B(B[24]), .A(n36), .Z(n6845) );
  XNOR U7043 ( .A(n6853), .B(n6955), .Z(n6846) );
  XNOR U7044 ( .A(n6852), .B(n6850), .Z(n6955) );
  AND U7045 ( .A(n6956), .B(n6957), .Z(n6850) );
  NANDN U7046 ( .A(n6958), .B(n6959), .Z(n6957) );
  NANDN U7047 ( .A(n6960), .B(n6961), .Z(n6959) );
  NANDN U7048 ( .A(n6961), .B(n6960), .Z(n6956) );
  ANDN U7049 ( .B(B[25]), .A(n37), .Z(n6852) );
  XNOR U7050 ( .A(n6860), .B(n6962), .Z(n6853) );
  XNOR U7051 ( .A(n6859), .B(n6857), .Z(n6962) );
  AND U7052 ( .A(n6963), .B(n6964), .Z(n6857) );
  NANDN U7053 ( .A(n6965), .B(n6966), .Z(n6964) );
  OR U7054 ( .A(n6967), .B(n6968), .Z(n6966) );
  NAND U7055 ( .A(n6968), .B(n6967), .Z(n6963) );
  ANDN U7056 ( .B(B[26]), .A(n38), .Z(n6859) );
  XNOR U7057 ( .A(n6867), .B(n6969), .Z(n6860) );
  XNOR U7058 ( .A(n6866), .B(n6864), .Z(n6969) );
  AND U7059 ( .A(n6970), .B(n6971), .Z(n6864) );
  NANDN U7060 ( .A(n6972), .B(n6973), .Z(n6971) );
  NANDN U7061 ( .A(n6974), .B(n6975), .Z(n6973) );
  NANDN U7062 ( .A(n6975), .B(n6974), .Z(n6970) );
  ANDN U7063 ( .B(B[27]), .A(n39), .Z(n6866) );
  XNOR U7064 ( .A(n6874), .B(n6976), .Z(n6867) );
  XNOR U7065 ( .A(n6873), .B(n6871), .Z(n6976) );
  AND U7066 ( .A(n6977), .B(n6978), .Z(n6871) );
  NANDN U7067 ( .A(n6979), .B(n6980), .Z(n6978) );
  OR U7068 ( .A(n6981), .B(n6982), .Z(n6980) );
  NAND U7069 ( .A(n6982), .B(n6981), .Z(n6977) );
  ANDN U7070 ( .B(B[28]), .A(n40), .Z(n6873) );
  XNOR U7071 ( .A(n6881), .B(n6983), .Z(n6874) );
  XNOR U7072 ( .A(n6880), .B(n6878), .Z(n6983) );
  AND U7073 ( .A(n6984), .B(n6985), .Z(n6878) );
  NANDN U7074 ( .A(n6986), .B(n6987), .Z(n6985) );
  NAND U7075 ( .A(n6988), .B(n6989), .Z(n6987) );
  ANDN U7076 ( .B(B[29]), .A(n41), .Z(n6880) );
  XOR U7077 ( .A(n6887), .B(n6990), .Z(n6881) );
  XNOR U7078 ( .A(n6885), .B(n6888), .Z(n6990) );
  NAND U7079 ( .A(A[2]), .B(B[30]), .Z(n6888) );
  NANDN U7080 ( .A(n6991), .B(n6992), .Z(n6885) );
  AND U7081 ( .A(A[0]), .B(B[31]), .Z(n6992) );
  XNOR U7082 ( .A(n6890), .B(n6993), .Z(n6887) );
  NAND U7083 ( .A(A[0]), .B(B[32]), .Z(n6993) );
  NAND U7084 ( .A(B[31]), .B(A[1]), .Z(n6890) );
  NAND U7085 ( .A(n6994), .B(n6995), .Z(n182) );
  NANDN U7086 ( .A(n6996), .B(n6997), .Z(n6995) );
  OR U7087 ( .A(n6998), .B(n6999), .Z(n6997) );
  NAND U7088 ( .A(n6999), .B(n6998), .Z(n6994) );
  XNOR U7089 ( .A(n7000), .B(n7001), .Z(\A1[2] ) );
  XNOR U7090 ( .A(n7002), .B(n7003), .Z(n7001) );
  XOR U7091 ( .A(n184), .B(n183), .Z(\A1[29] ) );
  XOR U7092 ( .A(n6999), .B(n7004), .Z(n183) );
  XNOR U7093 ( .A(n6998), .B(n6996), .Z(n7004) );
  AND U7094 ( .A(n7005), .B(n7006), .Z(n6996) );
  NANDN U7095 ( .A(n7007), .B(n7008), .Z(n7006) );
  NANDN U7096 ( .A(n7009), .B(n7010), .Z(n7008) );
  NANDN U7097 ( .A(n7010), .B(n7009), .Z(n7005) );
  ANDN U7098 ( .B(B[16]), .A(n29), .Z(n6998) );
  XNOR U7099 ( .A(n6905), .B(n7011), .Z(n6999) );
  XNOR U7100 ( .A(n6904), .B(n6902), .Z(n7011) );
  AND U7101 ( .A(n7012), .B(n7013), .Z(n6902) );
  NANDN U7102 ( .A(n7014), .B(n7015), .Z(n7013) );
  OR U7103 ( .A(n7016), .B(n7017), .Z(n7015) );
  NAND U7104 ( .A(n7017), .B(n7016), .Z(n7012) );
  ANDN U7105 ( .B(B[17]), .A(n30), .Z(n6904) );
  XNOR U7106 ( .A(n6912), .B(n7018), .Z(n6905) );
  XNOR U7107 ( .A(n6911), .B(n6909), .Z(n7018) );
  AND U7108 ( .A(n7019), .B(n7020), .Z(n6909) );
  NANDN U7109 ( .A(n7021), .B(n7022), .Z(n7020) );
  NANDN U7110 ( .A(n7023), .B(n7024), .Z(n7022) );
  NANDN U7111 ( .A(n7024), .B(n7023), .Z(n7019) );
  ANDN U7112 ( .B(B[18]), .A(n31), .Z(n6911) );
  XNOR U7113 ( .A(n6919), .B(n7025), .Z(n6912) );
  XNOR U7114 ( .A(n6918), .B(n6916), .Z(n7025) );
  AND U7115 ( .A(n7026), .B(n7027), .Z(n6916) );
  NANDN U7116 ( .A(n7028), .B(n7029), .Z(n7027) );
  OR U7117 ( .A(n7030), .B(n7031), .Z(n7029) );
  NAND U7118 ( .A(n7031), .B(n7030), .Z(n7026) );
  ANDN U7119 ( .B(B[19]), .A(n32), .Z(n6918) );
  XNOR U7120 ( .A(n6926), .B(n7032), .Z(n6919) );
  XNOR U7121 ( .A(n6925), .B(n6923), .Z(n7032) );
  AND U7122 ( .A(n7033), .B(n7034), .Z(n6923) );
  NANDN U7123 ( .A(n7035), .B(n7036), .Z(n7034) );
  NANDN U7124 ( .A(n7037), .B(n7038), .Z(n7036) );
  NANDN U7125 ( .A(n7038), .B(n7037), .Z(n7033) );
  ANDN U7126 ( .B(B[20]), .A(n33), .Z(n6925) );
  XNOR U7127 ( .A(n6933), .B(n7039), .Z(n6926) );
  XNOR U7128 ( .A(n6932), .B(n6930), .Z(n7039) );
  AND U7129 ( .A(n7040), .B(n7041), .Z(n6930) );
  NANDN U7130 ( .A(n7042), .B(n7043), .Z(n7041) );
  OR U7131 ( .A(n7044), .B(n7045), .Z(n7043) );
  NAND U7132 ( .A(n7045), .B(n7044), .Z(n7040) );
  ANDN U7133 ( .B(B[21]), .A(n34), .Z(n6932) );
  XNOR U7134 ( .A(n6940), .B(n7046), .Z(n6933) );
  XNOR U7135 ( .A(n6939), .B(n6937), .Z(n7046) );
  AND U7136 ( .A(n7047), .B(n7048), .Z(n6937) );
  NANDN U7137 ( .A(n7049), .B(n7050), .Z(n7048) );
  NANDN U7138 ( .A(n7051), .B(n7052), .Z(n7050) );
  NANDN U7139 ( .A(n7052), .B(n7051), .Z(n7047) );
  ANDN U7140 ( .B(B[22]), .A(n35), .Z(n6939) );
  XNOR U7141 ( .A(n6947), .B(n7053), .Z(n6940) );
  XNOR U7142 ( .A(n6946), .B(n6944), .Z(n7053) );
  AND U7143 ( .A(n7054), .B(n7055), .Z(n6944) );
  NANDN U7144 ( .A(n7056), .B(n7057), .Z(n7055) );
  OR U7145 ( .A(n7058), .B(n7059), .Z(n7057) );
  NAND U7146 ( .A(n7059), .B(n7058), .Z(n7054) );
  ANDN U7147 ( .B(B[23]), .A(n36), .Z(n6946) );
  XNOR U7148 ( .A(n6954), .B(n7060), .Z(n6947) );
  XNOR U7149 ( .A(n6953), .B(n6951), .Z(n7060) );
  AND U7150 ( .A(n7061), .B(n7062), .Z(n6951) );
  NANDN U7151 ( .A(n7063), .B(n7064), .Z(n7062) );
  NANDN U7152 ( .A(n7065), .B(n7066), .Z(n7064) );
  NANDN U7153 ( .A(n7066), .B(n7065), .Z(n7061) );
  ANDN U7154 ( .B(B[24]), .A(n37), .Z(n6953) );
  XNOR U7155 ( .A(n6961), .B(n7067), .Z(n6954) );
  XNOR U7156 ( .A(n6960), .B(n6958), .Z(n7067) );
  AND U7157 ( .A(n7068), .B(n7069), .Z(n6958) );
  NANDN U7158 ( .A(n7070), .B(n7071), .Z(n7069) );
  OR U7159 ( .A(n7072), .B(n7073), .Z(n7071) );
  NAND U7160 ( .A(n7073), .B(n7072), .Z(n7068) );
  ANDN U7161 ( .B(B[25]), .A(n38), .Z(n6960) );
  XNOR U7162 ( .A(n6968), .B(n7074), .Z(n6961) );
  XNOR U7163 ( .A(n6967), .B(n6965), .Z(n7074) );
  AND U7164 ( .A(n7075), .B(n7076), .Z(n6965) );
  NANDN U7165 ( .A(n7077), .B(n7078), .Z(n7076) );
  NANDN U7166 ( .A(n7079), .B(n7080), .Z(n7078) );
  NANDN U7167 ( .A(n7080), .B(n7079), .Z(n7075) );
  ANDN U7168 ( .B(B[26]), .A(n39), .Z(n6967) );
  XNOR U7169 ( .A(n6975), .B(n7081), .Z(n6968) );
  XNOR U7170 ( .A(n6974), .B(n6972), .Z(n7081) );
  AND U7171 ( .A(n7082), .B(n7083), .Z(n6972) );
  NANDN U7172 ( .A(n7084), .B(n7085), .Z(n7083) );
  OR U7173 ( .A(n7086), .B(n7087), .Z(n7085) );
  NAND U7174 ( .A(n7087), .B(n7086), .Z(n7082) );
  ANDN U7175 ( .B(B[27]), .A(n40), .Z(n6974) );
  XNOR U7176 ( .A(n6982), .B(n7088), .Z(n6975) );
  XNOR U7177 ( .A(n6981), .B(n6979), .Z(n7088) );
  AND U7178 ( .A(n7089), .B(n7090), .Z(n6979) );
  NANDN U7179 ( .A(n7091), .B(n7092), .Z(n7090) );
  NAND U7180 ( .A(n7093), .B(n7094), .Z(n7092) );
  ANDN U7181 ( .B(B[28]), .A(n41), .Z(n6981) );
  XOR U7182 ( .A(n6988), .B(n7095), .Z(n6982) );
  XNOR U7183 ( .A(n6986), .B(n6989), .Z(n7095) );
  NAND U7184 ( .A(A[2]), .B(B[29]), .Z(n6989) );
  NANDN U7185 ( .A(n7096), .B(n7097), .Z(n6986) );
  AND U7186 ( .A(A[0]), .B(B[30]), .Z(n7097) );
  XNOR U7187 ( .A(n6991), .B(n7098), .Z(n6988) );
  NAND U7188 ( .A(A[0]), .B(B[31]), .Z(n7098) );
  NAND U7189 ( .A(B[30]), .B(A[1]), .Z(n6991) );
  NAND U7190 ( .A(n7099), .B(n7100), .Z(n184) );
  NANDN U7191 ( .A(n7101), .B(n7102), .Z(n7100) );
  OR U7192 ( .A(n7103), .B(n7104), .Z(n7102) );
  NAND U7193 ( .A(n7104), .B(n7103), .Z(n7099) );
  XOR U7194 ( .A(n186), .B(n185), .Z(\A1[28] ) );
  XOR U7195 ( .A(n7104), .B(n7105), .Z(n185) );
  XNOR U7196 ( .A(n7103), .B(n7101), .Z(n7105) );
  AND U7197 ( .A(n7106), .B(n7107), .Z(n7101) );
  NANDN U7198 ( .A(n7108), .B(n7109), .Z(n7107) );
  NANDN U7199 ( .A(n7110), .B(n7111), .Z(n7109) );
  NANDN U7200 ( .A(n7111), .B(n7110), .Z(n7106) );
  ANDN U7201 ( .B(B[15]), .A(n29), .Z(n7103) );
  XNOR U7202 ( .A(n7010), .B(n7112), .Z(n7104) );
  XNOR U7203 ( .A(n7009), .B(n7007), .Z(n7112) );
  AND U7204 ( .A(n7113), .B(n7114), .Z(n7007) );
  NANDN U7205 ( .A(n7115), .B(n7116), .Z(n7114) );
  OR U7206 ( .A(n7117), .B(n7118), .Z(n7116) );
  NAND U7207 ( .A(n7118), .B(n7117), .Z(n7113) );
  ANDN U7208 ( .B(B[16]), .A(n30), .Z(n7009) );
  XNOR U7209 ( .A(n7017), .B(n7119), .Z(n7010) );
  XNOR U7210 ( .A(n7016), .B(n7014), .Z(n7119) );
  AND U7211 ( .A(n7120), .B(n7121), .Z(n7014) );
  NANDN U7212 ( .A(n7122), .B(n7123), .Z(n7121) );
  NANDN U7213 ( .A(n7124), .B(n7125), .Z(n7123) );
  NANDN U7214 ( .A(n7125), .B(n7124), .Z(n7120) );
  ANDN U7215 ( .B(B[17]), .A(n31), .Z(n7016) );
  XNOR U7216 ( .A(n7024), .B(n7126), .Z(n7017) );
  XNOR U7217 ( .A(n7023), .B(n7021), .Z(n7126) );
  AND U7218 ( .A(n7127), .B(n7128), .Z(n7021) );
  NANDN U7219 ( .A(n7129), .B(n7130), .Z(n7128) );
  OR U7220 ( .A(n7131), .B(n7132), .Z(n7130) );
  NAND U7221 ( .A(n7132), .B(n7131), .Z(n7127) );
  ANDN U7222 ( .B(B[18]), .A(n32), .Z(n7023) );
  XNOR U7223 ( .A(n7031), .B(n7133), .Z(n7024) );
  XNOR U7224 ( .A(n7030), .B(n7028), .Z(n7133) );
  AND U7225 ( .A(n7134), .B(n7135), .Z(n7028) );
  NANDN U7226 ( .A(n7136), .B(n7137), .Z(n7135) );
  NANDN U7227 ( .A(n7138), .B(n7139), .Z(n7137) );
  NANDN U7228 ( .A(n7139), .B(n7138), .Z(n7134) );
  ANDN U7229 ( .B(B[19]), .A(n33), .Z(n7030) );
  XNOR U7230 ( .A(n7038), .B(n7140), .Z(n7031) );
  XNOR U7231 ( .A(n7037), .B(n7035), .Z(n7140) );
  AND U7232 ( .A(n7141), .B(n7142), .Z(n7035) );
  NANDN U7233 ( .A(n7143), .B(n7144), .Z(n7142) );
  OR U7234 ( .A(n7145), .B(n7146), .Z(n7144) );
  NAND U7235 ( .A(n7146), .B(n7145), .Z(n7141) );
  ANDN U7236 ( .B(B[20]), .A(n34), .Z(n7037) );
  XNOR U7237 ( .A(n7045), .B(n7147), .Z(n7038) );
  XNOR U7238 ( .A(n7044), .B(n7042), .Z(n7147) );
  AND U7239 ( .A(n7148), .B(n7149), .Z(n7042) );
  NANDN U7240 ( .A(n7150), .B(n7151), .Z(n7149) );
  NANDN U7241 ( .A(n7152), .B(n7153), .Z(n7151) );
  NANDN U7242 ( .A(n7153), .B(n7152), .Z(n7148) );
  ANDN U7243 ( .B(B[21]), .A(n35), .Z(n7044) );
  XNOR U7244 ( .A(n7052), .B(n7154), .Z(n7045) );
  XNOR U7245 ( .A(n7051), .B(n7049), .Z(n7154) );
  AND U7246 ( .A(n7155), .B(n7156), .Z(n7049) );
  NANDN U7247 ( .A(n7157), .B(n7158), .Z(n7156) );
  OR U7248 ( .A(n7159), .B(n7160), .Z(n7158) );
  NAND U7249 ( .A(n7160), .B(n7159), .Z(n7155) );
  ANDN U7250 ( .B(B[22]), .A(n36), .Z(n7051) );
  XNOR U7251 ( .A(n7059), .B(n7161), .Z(n7052) );
  XNOR U7252 ( .A(n7058), .B(n7056), .Z(n7161) );
  AND U7253 ( .A(n7162), .B(n7163), .Z(n7056) );
  NANDN U7254 ( .A(n7164), .B(n7165), .Z(n7163) );
  NANDN U7255 ( .A(n7166), .B(n7167), .Z(n7165) );
  NANDN U7256 ( .A(n7167), .B(n7166), .Z(n7162) );
  ANDN U7257 ( .B(B[23]), .A(n37), .Z(n7058) );
  XNOR U7258 ( .A(n7066), .B(n7168), .Z(n7059) );
  XNOR U7259 ( .A(n7065), .B(n7063), .Z(n7168) );
  AND U7260 ( .A(n7169), .B(n7170), .Z(n7063) );
  NANDN U7261 ( .A(n7171), .B(n7172), .Z(n7170) );
  OR U7262 ( .A(n7173), .B(n7174), .Z(n7172) );
  NAND U7263 ( .A(n7174), .B(n7173), .Z(n7169) );
  ANDN U7264 ( .B(B[24]), .A(n38), .Z(n7065) );
  XNOR U7265 ( .A(n7073), .B(n7175), .Z(n7066) );
  XNOR U7266 ( .A(n7072), .B(n7070), .Z(n7175) );
  AND U7267 ( .A(n7176), .B(n7177), .Z(n7070) );
  NANDN U7268 ( .A(n7178), .B(n7179), .Z(n7177) );
  NANDN U7269 ( .A(n7180), .B(n7181), .Z(n7179) );
  NANDN U7270 ( .A(n7181), .B(n7180), .Z(n7176) );
  ANDN U7271 ( .B(B[25]), .A(n39), .Z(n7072) );
  XNOR U7272 ( .A(n7080), .B(n7182), .Z(n7073) );
  XNOR U7273 ( .A(n7079), .B(n7077), .Z(n7182) );
  AND U7274 ( .A(n7183), .B(n7184), .Z(n7077) );
  NANDN U7275 ( .A(n7185), .B(n7186), .Z(n7184) );
  OR U7276 ( .A(n7187), .B(n7188), .Z(n7186) );
  NAND U7277 ( .A(n7188), .B(n7187), .Z(n7183) );
  ANDN U7278 ( .B(B[26]), .A(n40), .Z(n7079) );
  XNOR U7279 ( .A(n7087), .B(n7189), .Z(n7080) );
  XNOR U7280 ( .A(n7086), .B(n7084), .Z(n7189) );
  AND U7281 ( .A(n7190), .B(n7191), .Z(n7084) );
  NANDN U7282 ( .A(n7192), .B(n7193), .Z(n7191) );
  NAND U7283 ( .A(n7194), .B(n7195), .Z(n7193) );
  ANDN U7284 ( .B(B[27]), .A(n41), .Z(n7086) );
  XOR U7285 ( .A(n7093), .B(n7196), .Z(n7087) );
  XNOR U7286 ( .A(n7091), .B(n7094), .Z(n7196) );
  NAND U7287 ( .A(A[2]), .B(B[28]), .Z(n7094) );
  NANDN U7288 ( .A(n7197), .B(n7198), .Z(n7091) );
  AND U7289 ( .A(A[0]), .B(B[29]), .Z(n7198) );
  XNOR U7290 ( .A(n7096), .B(n7199), .Z(n7093) );
  NAND U7291 ( .A(A[0]), .B(B[30]), .Z(n7199) );
  NAND U7292 ( .A(B[29]), .B(A[1]), .Z(n7096) );
  NAND U7293 ( .A(n7200), .B(n7201), .Z(n186) );
  NANDN U7294 ( .A(n7202), .B(n7203), .Z(n7201) );
  OR U7295 ( .A(n7204), .B(n7205), .Z(n7203) );
  NAND U7296 ( .A(n7205), .B(n7204), .Z(n7200) );
  XOR U7297 ( .A(n188), .B(n187), .Z(\A1[27] ) );
  XOR U7298 ( .A(n7205), .B(n7206), .Z(n187) );
  XNOR U7299 ( .A(n7204), .B(n7202), .Z(n7206) );
  AND U7300 ( .A(n7207), .B(n7208), .Z(n7202) );
  NANDN U7301 ( .A(n7209), .B(n7210), .Z(n7208) );
  NANDN U7302 ( .A(n7211), .B(n7212), .Z(n7210) );
  NANDN U7303 ( .A(n7212), .B(n7211), .Z(n7207) );
  ANDN U7304 ( .B(B[14]), .A(n29), .Z(n7204) );
  XNOR U7305 ( .A(n7111), .B(n7213), .Z(n7205) );
  XNOR U7306 ( .A(n7110), .B(n7108), .Z(n7213) );
  AND U7307 ( .A(n7214), .B(n7215), .Z(n7108) );
  NANDN U7308 ( .A(n7216), .B(n7217), .Z(n7215) );
  OR U7309 ( .A(n7218), .B(n7219), .Z(n7217) );
  NAND U7310 ( .A(n7219), .B(n7218), .Z(n7214) );
  ANDN U7311 ( .B(B[15]), .A(n30), .Z(n7110) );
  XNOR U7312 ( .A(n7118), .B(n7220), .Z(n7111) );
  XNOR U7313 ( .A(n7117), .B(n7115), .Z(n7220) );
  AND U7314 ( .A(n7221), .B(n7222), .Z(n7115) );
  NANDN U7315 ( .A(n7223), .B(n7224), .Z(n7222) );
  NANDN U7316 ( .A(n7225), .B(n7226), .Z(n7224) );
  NANDN U7317 ( .A(n7226), .B(n7225), .Z(n7221) );
  ANDN U7318 ( .B(B[16]), .A(n31), .Z(n7117) );
  XNOR U7319 ( .A(n7125), .B(n7227), .Z(n7118) );
  XNOR U7320 ( .A(n7124), .B(n7122), .Z(n7227) );
  AND U7321 ( .A(n7228), .B(n7229), .Z(n7122) );
  NANDN U7322 ( .A(n7230), .B(n7231), .Z(n7229) );
  OR U7323 ( .A(n7232), .B(n7233), .Z(n7231) );
  NAND U7324 ( .A(n7233), .B(n7232), .Z(n7228) );
  ANDN U7325 ( .B(B[17]), .A(n32), .Z(n7124) );
  XNOR U7326 ( .A(n7132), .B(n7234), .Z(n7125) );
  XNOR U7327 ( .A(n7131), .B(n7129), .Z(n7234) );
  AND U7328 ( .A(n7235), .B(n7236), .Z(n7129) );
  NANDN U7329 ( .A(n7237), .B(n7238), .Z(n7236) );
  NANDN U7330 ( .A(n7239), .B(n7240), .Z(n7238) );
  NANDN U7331 ( .A(n7240), .B(n7239), .Z(n7235) );
  ANDN U7332 ( .B(B[18]), .A(n33), .Z(n7131) );
  XNOR U7333 ( .A(n7139), .B(n7241), .Z(n7132) );
  XNOR U7334 ( .A(n7138), .B(n7136), .Z(n7241) );
  AND U7335 ( .A(n7242), .B(n7243), .Z(n7136) );
  NANDN U7336 ( .A(n7244), .B(n7245), .Z(n7243) );
  OR U7337 ( .A(n7246), .B(n7247), .Z(n7245) );
  NAND U7338 ( .A(n7247), .B(n7246), .Z(n7242) );
  ANDN U7339 ( .B(B[19]), .A(n34), .Z(n7138) );
  XNOR U7340 ( .A(n7146), .B(n7248), .Z(n7139) );
  XNOR U7341 ( .A(n7145), .B(n7143), .Z(n7248) );
  AND U7342 ( .A(n7249), .B(n7250), .Z(n7143) );
  NANDN U7343 ( .A(n7251), .B(n7252), .Z(n7250) );
  NANDN U7344 ( .A(n7253), .B(n7254), .Z(n7252) );
  NANDN U7345 ( .A(n7254), .B(n7253), .Z(n7249) );
  ANDN U7346 ( .B(B[20]), .A(n35), .Z(n7145) );
  XNOR U7347 ( .A(n7153), .B(n7255), .Z(n7146) );
  XNOR U7348 ( .A(n7152), .B(n7150), .Z(n7255) );
  AND U7349 ( .A(n7256), .B(n7257), .Z(n7150) );
  NANDN U7350 ( .A(n7258), .B(n7259), .Z(n7257) );
  OR U7351 ( .A(n7260), .B(n7261), .Z(n7259) );
  NAND U7352 ( .A(n7261), .B(n7260), .Z(n7256) );
  ANDN U7353 ( .B(B[21]), .A(n36), .Z(n7152) );
  XNOR U7354 ( .A(n7160), .B(n7262), .Z(n7153) );
  XNOR U7355 ( .A(n7159), .B(n7157), .Z(n7262) );
  AND U7356 ( .A(n7263), .B(n7264), .Z(n7157) );
  NANDN U7357 ( .A(n7265), .B(n7266), .Z(n7264) );
  NANDN U7358 ( .A(n7267), .B(n7268), .Z(n7266) );
  NANDN U7359 ( .A(n7268), .B(n7267), .Z(n7263) );
  ANDN U7360 ( .B(B[22]), .A(n37), .Z(n7159) );
  XNOR U7361 ( .A(n7167), .B(n7269), .Z(n7160) );
  XNOR U7362 ( .A(n7166), .B(n7164), .Z(n7269) );
  AND U7363 ( .A(n7270), .B(n7271), .Z(n7164) );
  NANDN U7364 ( .A(n7272), .B(n7273), .Z(n7271) );
  OR U7365 ( .A(n7274), .B(n7275), .Z(n7273) );
  NAND U7366 ( .A(n7275), .B(n7274), .Z(n7270) );
  ANDN U7367 ( .B(B[23]), .A(n38), .Z(n7166) );
  XNOR U7368 ( .A(n7174), .B(n7276), .Z(n7167) );
  XNOR U7369 ( .A(n7173), .B(n7171), .Z(n7276) );
  AND U7370 ( .A(n7277), .B(n7278), .Z(n7171) );
  NANDN U7371 ( .A(n7279), .B(n7280), .Z(n7278) );
  NANDN U7372 ( .A(n7281), .B(n7282), .Z(n7280) );
  NANDN U7373 ( .A(n7282), .B(n7281), .Z(n7277) );
  ANDN U7374 ( .B(B[24]), .A(n39), .Z(n7173) );
  XNOR U7375 ( .A(n7181), .B(n7283), .Z(n7174) );
  XNOR U7376 ( .A(n7180), .B(n7178), .Z(n7283) );
  AND U7377 ( .A(n7284), .B(n7285), .Z(n7178) );
  NANDN U7378 ( .A(n7286), .B(n7287), .Z(n7285) );
  OR U7379 ( .A(n7288), .B(n7289), .Z(n7287) );
  NAND U7380 ( .A(n7289), .B(n7288), .Z(n7284) );
  ANDN U7381 ( .B(B[25]), .A(n40), .Z(n7180) );
  XNOR U7382 ( .A(n7188), .B(n7290), .Z(n7181) );
  XNOR U7383 ( .A(n7187), .B(n7185), .Z(n7290) );
  AND U7384 ( .A(n7291), .B(n7292), .Z(n7185) );
  NANDN U7385 ( .A(n7293), .B(n7294), .Z(n7292) );
  NAND U7386 ( .A(n7295), .B(n7296), .Z(n7294) );
  ANDN U7387 ( .B(B[26]), .A(n41), .Z(n7187) );
  XOR U7388 ( .A(n7194), .B(n7297), .Z(n7188) );
  XNOR U7389 ( .A(n7192), .B(n7195), .Z(n7297) );
  NAND U7390 ( .A(A[2]), .B(B[27]), .Z(n7195) );
  NANDN U7391 ( .A(n7298), .B(n7299), .Z(n7192) );
  AND U7392 ( .A(A[0]), .B(B[28]), .Z(n7299) );
  XNOR U7393 ( .A(n7197), .B(n7300), .Z(n7194) );
  NAND U7394 ( .A(A[0]), .B(B[29]), .Z(n7300) );
  NAND U7395 ( .A(B[28]), .B(A[1]), .Z(n7197) );
  NAND U7396 ( .A(n7301), .B(n7302), .Z(n188) );
  NANDN U7397 ( .A(n7303), .B(n7304), .Z(n7302) );
  OR U7398 ( .A(n7305), .B(n7306), .Z(n7304) );
  NAND U7399 ( .A(n7306), .B(n7305), .Z(n7301) );
  XOR U7400 ( .A(n190), .B(n189), .Z(\A1[26] ) );
  XOR U7401 ( .A(n7306), .B(n7307), .Z(n189) );
  XNOR U7402 ( .A(n7305), .B(n7303), .Z(n7307) );
  AND U7403 ( .A(n7308), .B(n7309), .Z(n7303) );
  NANDN U7404 ( .A(n7310), .B(n7311), .Z(n7309) );
  NANDN U7405 ( .A(n7312), .B(n7313), .Z(n7311) );
  NANDN U7406 ( .A(n7313), .B(n7312), .Z(n7308) );
  ANDN U7407 ( .B(B[13]), .A(n29), .Z(n7305) );
  XNOR U7408 ( .A(n7212), .B(n7314), .Z(n7306) );
  XNOR U7409 ( .A(n7211), .B(n7209), .Z(n7314) );
  AND U7410 ( .A(n7315), .B(n7316), .Z(n7209) );
  NANDN U7411 ( .A(n7317), .B(n7318), .Z(n7316) );
  OR U7412 ( .A(n7319), .B(n7320), .Z(n7318) );
  NAND U7413 ( .A(n7320), .B(n7319), .Z(n7315) );
  ANDN U7414 ( .B(B[14]), .A(n30), .Z(n7211) );
  XNOR U7415 ( .A(n7219), .B(n7321), .Z(n7212) );
  XNOR U7416 ( .A(n7218), .B(n7216), .Z(n7321) );
  AND U7417 ( .A(n7322), .B(n7323), .Z(n7216) );
  NANDN U7418 ( .A(n7324), .B(n7325), .Z(n7323) );
  NANDN U7419 ( .A(n7326), .B(n7327), .Z(n7325) );
  NANDN U7420 ( .A(n7327), .B(n7326), .Z(n7322) );
  ANDN U7421 ( .B(B[15]), .A(n31), .Z(n7218) );
  XNOR U7422 ( .A(n7226), .B(n7328), .Z(n7219) );
  XNOR U7423 ( .A(n7225), .B(n7223), .Z(n7328) );
  AND U7424 ( .A(n7329), .B(n7330), .Z(n7223) );
  NANDN U7425 ( .A(n7331), .B(n7332), .Z(n7330) );
  OR U7426 ( .A(n7333), .B(n7334), .Z(n7332) );
  NAND U7427 ( .A(n7334), .B(n7333), .Z(n7329) );
  ANDN U7428 ( .B(B[16]), .A(n32), .Z(n7225) );
  XNOR U7429 ( .A(n7233), .B(n7335), .Z(n7226) );
  XNOR U7430 ( .A(n7232), .B(n7230), .Z(n7335) );
  AND U7431 ( .A(n7336), .B(n7337), .Z(n7230) );
  NANDN U7432 ( .A(n7338), .B(n7339), .Z(n7337) );
  NANDN U7433 ( .A(n7340), .B(n7341), .Z(n7339) );
  NANDN U7434 ( .A(n7341), .B(n7340), .Z(n7336) );
  ANDN U7435 ( .B(B[17]), .A(n33), .Z(n7232) );
  XNOR U7436 ( .A(n7240), .B(n7342), .Z(n7233) );
  XNOR U7437 ( .A(n7239), .B(n7237), .Z(n7342) );
  AND U7438 ( .A(n7343), .B(n7344), .Z(n7237) );
  NANDN U7439 ( .A(n7345), .B(n7346), .Z(n7344) );
  OR U7440 ( .A(n7347), .B(n7348), .Z(n7346) );
  NAND U7441 ( .A(n7348), .B(n7347), .Z(n7343) );
  ANDN U7442 ( .B(B[18]), .A(n34), .Z(n7239) );
  XNOR U7443 ( .A(n7247), .B(n7349), .Z(n7240) );
  XNOR U7444 ( .A(n7246), .B(n7244), .Z(n7349) );
  AND U7445 ( .A(n7350), .B(n7351), .Z(n7244) );
  NANDN U7446 ( .A(n7352), .B(n7353), .Z(n7351) );
  NANDN U7447 ( .A(n7354), .B(n7355), .Z(n7353) );
  NANDN U7448 ( .A(n7355), .B(n7354), .Z(n7350) );
  ANDN U7449 ( .B(B[19]), .A(n35), .Z(n7246) );
  XNOR U7450 ( .A(n7254), .B(n7356), .Z(n7247) );
  XNOR U7451 ( .A(n7253), .B(n7251), .Z(n7356) );
  AND U7452 ( .A(n7357), .B(n7358), .Z(n7251) );
  NANDN U7453 ( .A(n7359), .B(n7360), .Z(n7358) );
  OR U7454 ( .A(n7361), .B(n7362), .Z(n7360) );
  NAND U7455 ( .A(n7362), .B(n7361), .Z(n7357) );
  ANDN U7456 ( .B(B[20]), .A(n36), .Z(n7253) );
  XNOR U7457 ( .A(n7261), .B(n7363), .Z(n7254) );
  XNOR U7458 ( .A(n7260), .B(n7258), .Z(n7363) );
  AND U7459 ( .A(n7364), .B(n7365), .Z(n7258) );
  NANDN U7460 ( .A(n7366), .B(n7367), .Z(n7365) );
  NANDN U7461 ( .A(n7368), .B(n7369), .Z(n7367) );
  NANDN U7462 ( .A(n7369), .B(n7368), .Z(n7364) );
  ANDN U7463 ( .B(B[21]), .A(n37), .Z(n7260) );
  XNOR U7464 ( .A(n7268), .B(n7370), .Z(n7261) );
  XNOR U7465 ( .A(n7267), .B(n7265), .Z(n7370) );
  AND U7466 ( .A(n7371), .B(n7372), .Z(n7265) );
  NANDN U7467 ( .A(n7373), .B(n7374), .Z(n7372) );
  OR U7468 ( .A(n7375), .B(n7376), .Z(n7374) );
  NAND U7469 ( .A(n7376), .B(n7375), .Z(n7371) );
  ANDN U7470 ( .B(B[22]), .A(n38), .Z(n7267) );
  XNOR U7471 ( .A(n7275), .B(n7377), .Z(n7268) );
  XNOR U7472 ( .A(n7274), .B(n7272), .Z(n7377) );
  AND U7473 ( .A(n7378), .B(n7379), .Z(n7272) );
  NANDN U7474 ( .A(n7380), .B(n7381), .Z(n7379) );
  NANDN U7475 ( .A(n7382), .B(n7383), .Z(n7381) );
  NANDN U7476 ( .A(n7383), .B(n7382), .Z(n7378) );
  ANDN U7477 ( .B(B[23]), .A(n39), .Z(n7274) );
  XNOR U7478 ( .A(n7282), .B(n7384), .Z(n7275) );
  XNOR U7479 ( .A(n7281), .B(n7279), .Z(n7384) );
  AND U7480 ( .A(n7385), .B(n7386), .Z(n7279) );
  NANDN U7481 ( .A(n7387), .B(n7388), .Z(n7386) );
  OR U7482 ( .A(n7389), .B(n7390), .Z(n7388) );
  NAND U7483 ( .A(n7390), .B(n7389), .Z(n7385) );
  ANDN U7484 ( .B(B[24]), .A(n40), .Z(n7281) );
  XNOR U7485 ( .A(n7289), .B(n7391), .Z(n7282) );
  XNOR U7486 ( .A(n7288), .B(n7286), .Z(n7391) );
  AND U7487 ( .A(n7392), .B(n7393), .Z(n7286) );
  NANDN U7488 ( .A(n7394), .B(n7395), .Z(n7393) );
  NAND U7489 ( .A(n7396), .B(n7397), .Z(n7395) );
  ANDN U7490 ( .B(B[25]), .A(n41), .Z(n7288) );
  XOR U7491 ( .A(n7295), .B(n7398), .Z(n7289) );
  XNOR U7492 ( .A(n7293), .B(n7296), .Z(n7398) );
  NAND U7493 ( .A(A[2]), .B(B[26]), .Z(n7296) );
  NANDN U7494 ( .A(n7399), .B(n7400), .Z(n7293) );
  AND U7495 ( .A(A[0]), .B(B[27]), .Z(n7400) );
  XNOR U7496 ( .A(n7298), .B(n7401), .Z(n7295) );
  NAND U7497 ( .A(A[0]), .B(B[28]), .Z(n7401) );
  NAND U7498 ( .A(B[27]), .B(A[1]), .Z(n7298) );
  NAND U7499 ( .A(n7402), .B(n7403), .Z(n190) );
  NANDN U7500 ( .A(n7404), .B(n7405), .Z(n7403) );
  OR U7501 ( .A(n7406), .B(n7407), .Z(n7405) );
  NAND U7502 ( .A(n7407), .B(n7406), .Z(n7402) );
  XNOR U7504 ( .A(n193), .B(n7408), .Z(\A1[268] ) );
  NAND U7505 ( .A(A[15]), .B(B[255]), .Z(n7408) );
  NAND U7506 ( .A(n7409), .B(n7410), .Z(n193) );
  NAND U7507 ( .A(n7411), .B(n7412), .Z(n7410) );
  NANDN U7508 ( .A(n7413), .B(n7414), .Z(n7411) );
  NANDN U7509 ( .A(n7414), .B(n7413), .Z(n7409) );
  XOR U7510 ( .A(n195), .B(n194), .Z(\A1[267] ) );
  XNOR U7511 ( .A(n7412), .B(n7415), .Z(n194) );
  XOR U7512 ( .A(n7413), .B(n7414), .Z(n7415) );
  NAND U7513 ( .A(A[14]), .B(B[255]), .Z(n7414) );
  AND U7514 ( .A(B[254]), .B(A[15]), .Z(n7413) );
  NAND U7515 ( .A(n7416), .B(n7417), .Z(n7412) );
  NAND U7516 ( .A(n7418), .B(n7419), .Z(n7417) );
  NANDN U7517 ( .A(n7420), .B(n7421), .Z(n7418) );
  NANDN U7518 ( .A(n7421), .B(n7420), .Z(n7416) );
  NAND U7519 ( .A(n7422), .B(n7423), .Z(n195) );
  NANDN U7520 ( .A(n7424), .B(n7425), .Z(n7423) );
  NAND U7521 ( .A(n7427), .B(n7426), .Z(n7422) );
  XOR U7522 ( .A(n197), .B(n196), .Z(\A1[266] ) );
  XOR U7523 ( .A(n7427), .B(n7428), .Z(n196) );
  XNOR U7524 ( .A(n7426), .B(n7424), .Z(n7428) );
  AND U7525 ( .A(n7429), .B(n7430), .Z(n7424) );
  NANDN U7526 ( .A(n7431), .B(n7432), .Z(n7430) );
  NANDN U7527 ( .A(n7433), .B(n7434), .Z(n7432) );
  NANDN U7528 ( .A(n7434), .B(n7433), .Z(n7429) );
  ANDN U7529 ( .B(B[253]), .A(n29), .Z(n7426) );
  XNOR U7530 ( .A(n7419), .B(n7435), .Z(n7427) );
  XOR U7531 ( .A(n7420), .B(n7421), .Z(n7435) );
  NAND U7532 ( .A(A[13]), .B(B[255]), .Z(n7421) );
  AND U7533 ( .A(B[254]), .B(A[14]), .Z(n7420) );
  NAND U7534 ( .A(n7436), .B(n7437), .Z(n7419) );
  NAND U7535 ( .A(n7438), .B(n7439), .Z(n7437) );
  NANDN U7536 ( .A(n7440), .B(n7441), .Z(n7438) );
  NANDN U7537 ( .A(n7441), .B(n7440), .Z(n7436) );
  NAND U7538 ( .A(n7442), .B(n7443), .Z(n197) );
  NANDN U7539 ( .A(n7444), .B(n7445), .Z(n7443) );
  OR U7540 ( .A(n7446), .B(n7447), .Z(n7445) );
  NAND U7541 ( .A(n7447), .B(n7446), .Z(n7442) );
  XOR U7542 ( .A(n199), .B(n198), .Z(\A1[265] ) );
  XOR U7543 ( .A(n7447), .B(n7448), .Z(n198) );
  XNOR U7544 ( .A(n7446), .B(n7444), .Z(n7448) );
  AND U7545 ( .A(n7449), .B(n7450), .Z(n7444) );
  NANDN U7546 ( .A(n7451), .B(n7452), .Z(n7450) );
  OR U7547 ( .A(n7453), .B(n7454), .Z(n7452) );
  NAND U7548 ( .A(n7454), .B(n7453), .Z(n7449) );
  ANDN U7549 ( .B(B[252]), .A(n29), .Z(n7446) );
  XNOR U7550 ( .A(n7434), .B(n7455), .Z(n7447) );
  XNOR U7551 ( .A(n7433), .B(n7431), .Z(n7455) );
  AND U7552 ( .A(n7456), .B(n7457), .Z(n7431) );
  NANDN U7553 ( .A(n7458), .B(n7459), .Z(n7457) );
  NANDN U7554 ( .A(n7460), .B(n7461), .Z(n7459) );
  NANDN U7555 ( .A(n7461), .B(n7460), .Z(n7456) );
  ANDN U7556 ( .B(B[253]), .A(n30), .Z(n7433) );
  XOR U7557 ( .A(n7439), .B(n7462), .Z(n7434) );
  XOR U7558 ( .A(n7440), .B(n7441), .Z(n7462) );
  NAND U7559 ( .A(A[12]), .B(B[255]), .Z(n7441) );
  AND U7560 ( .A(B[254]), .B(A[13]), .Z(n7440) );
  NAND U7561 ( .A(n7463), .B(n7464), .Z(n7439) );
  NAND U7562 ( .A(n7465), .B(n7466), .Z(n7464) );
  NANDN U7563 ( .A(n7467), .B(n7468), .Z(n7465) );
  NANDN U7564 ( .A(n7468), .B(n7467), .Z(n7463) );
  NAND U7565 ( .A(n7469), .B(n7470), .Z(n199) );
  NANDN U7566 ( .A(n7471), .B(n7472), .Z(n7470) );
  NAND U7567 ( .A(n7474), .B(n7473), .Z(n7469) );
  XOR U7568 ( .A(n201), .B(n200), .Z(\A1[264] ) );
  XOR U7569 ( .A(n7474), .B(n7475), .Z(n200) );
  XNOR U7570 ( .A(n7473), .B(n7471), .Z(n7475) );
  AND U7571 ( .A(n7476), .B(n7477), .Z(n7471) );
  NANDN U7572 ( .A(n7478), .B(n7479), .Z(n7477) );
  NANDN U7573 ( .A(n7480), .B(n7481), .Z(n7479) );
  NANDN U7574 ( .A(n7481), .B(n7480), .Z(n7476) );
  ANDN U7575 ( .B(B[251]), .A(n29), .Z(n7473) );
  XOR U7576 ( .A(n7454), .B(n7482), .Z(n7474) );
  XNOR U7577 ( .A(n7453), .B(n7451), .Z(n7482) );
  AND U7578 ( .A(n7483), .B(n7484), .Z(n7451) );
  NANDN U7579 ( .A(n7485), .B(n7486), .Z(n7484) );
  OR U7580 ( .A(n7487), .B(n7488), .Z(n7486) );
  NAND U7581 ( .A(n7488), .B(n7487), .Z(n7483) );
  ANDN U7582 ( .B(B[252]), .A(n30), .Z(n7453) );
  XNOR U7583 ( .A(n7461), .B(n7489), .Z(n7454) );
  XNOR U7584 ( .A(n7460), .B(n7458), .Z(n7489) );
  AND U7585 ( .A(n7490), .B(n7491), .Z(n7458) );
  NANDN U7586 ( .A(n7492), .B(n7493), .Z(n7491) );
  NANDN U7587 ( .A(n7494), .B(n7495), .Z(n7493) );
  NANDN U7588 ( .A(n7495), .B(n7494), .Z(n7490) );
  ANDN U7589 ( .B(B[253]), .A(n31), .Z(n7460) );
  XOR U7590 ( .A(n7466), .B(n7496), .Z(n7461) );
  XOR U7591 ( .A(n7467), .B(n7468), .Z(n7496) );
  NAND U7592 ( .A(A[11]), .B(B[255]), .Z(n7468) );
  AND U7593 ( .A(B[254]), .B(A[12]), .Z(n7467) );
  NAND U7594 ( .A(n7497), .B(n7498), .Z(n7466) );
  NAND U7595 ( .A(n7499), .B(n7500), .Z(n7498) );
  NANDN U7596 ( .A(n7501), .B(n7502), .Z(n7499) );
  NANDN U7597 ( .A(n7502), .B(n7501), .Z(n7497) );
  NAND U7598 ( .A(n7503), .B(n7504), .Z(n201) );
  NANDN U7599 ( .A(n7505), .B(n7506), .Z(n7504) );
  OR U7600 ( .A(n7507), .B(n7508), .Z(n7506) );
  NAND U7601 ( .A(n7508), .B(n7507), .Z(n7503) );
  XOR U7602 ( .A(n203), .B(n202), .Z(\A1[263] ) );
  XOR U7603 ( .A(n7508), .B(n7509), .Z(n202) );
  XNOR U7604 ( .A(n7507), .B(n7505), .Z(n7509) );
  AND U7605 ( .A(n7510), .B(n7511), .Z(n7505) );
  NANDN U7606 ( .A(n7512), .B(n7513), .Z(n7511) );
  OR U7607 ( .A(n7514), .B(n7515), .Z(n7513) );
  NAND U7608 ( .A(n7515), .B(n7514), .Z(n7510) );
  ANDN U7609 ( .B(B[250]), .A(n29), .Z(n7507) );
  XNOR U7610 ( .A(n7481), .B(n7516), .Z(n7508) );
  XNOR U7611 ( .A(n7480), .B(n7478), .Z(n7516) );
  AND U7612 ( .A(n7517), .B(n7518), .Z(n7478) );
  NANDN U7613 ( .A(n7519), .B(n7520), .Z(n7518) );
  NANDN U7614 ( .A(n7521), .B(n7522), .Z(n7520) );
  NANDN U7615 ( .A(n7522), .B(n7521), .Z(n7517) );
  ANDN U7616 ( .B(B[251]), .A(n30), .Z(n7480) );
  XNOR U7617 ( .A(n7488), .B(n7523), .Z(n7481) );
  XNOR U7618 ( .A(n7487), .B(n7485), .Z(n7523) );
  AND U7619 ( .A(n7524), .B(n7525), .Z(n7485) );
  NANDN U7620 ( .A(n7526), .B(n7527), .Z(n7525) );
  OR U7621 ( .A(n7528), .B(n7529), .Z(n7527) );
  NAND U7622 ( .A(n7529), .B(n7528), .Z(n7524) );
  ANDN U7623 ( .B(B[252]), .A(n31), .Z(n7487) );
  XNOR U7624 ( .A(n7495), .B(n7530), .Z(n7488) );
  XNOR U7625 ( .A(n7494), .B(n7492), .Z(n7530) );
  AND U7626 ( .A(n7531), .B(n7532), .Z(n7492) );
  NANDN U7627 ( .A(n7533), .B(n7534), .Z(n7532) );
  NANDN U7628 ( .A(n7535), .B(n7536), .Z(n7534) );
  NANDN U7629 ( .A(n7536), .B(n7535), .Z(n7531) );
  ANDN U7630 ( .B(B[253]), .A(n32), .Z(n7494) );
  XOR U7631 ( .A(n7500), .B(n7537), .Z(n7495) );
  XOR U7632 ( .A(n7501), .B(n7502), .Z(n7537) );
  NAND U7633 ( .A(A[10]), .B(B[255]), .Z(n7502) );
  AND U7634 ( .A(B[254]), .B(A[11]), .Z(n7501) );
  NAND U7635 ( .A(n7538), .B(n7539), .Z(n7500) );
  NAND U7636 ( .A(n7540), .B(n7541), .Z(n7539) );
  NANDN U7637 ( .A(n7542), .B(n7543), .Z(n7540) );
  NANDN U7638 ( .A(n7543), .B(n7542), .Z(n7538) );
  NAND U7639 ( .A(n7544), .B(n7545), .Z(n203) );
  NANDN U7640 ( .A(n7546), .B(n7547), .Z(n7545) );
  NAND U7641 ( .A(n7549), .B(n7548), .Z(n7544) );
  XOR U7642 ( .A(n205), .B(n204), .Z(\A1[262] ) );
  XOR U7643 ( .A(n7549), .B(n7550), .Z(n204) );
  XNOR U7644 ( .A(n7548), .B(n7546), .Z(n7550) );
  AND U7645 ( .A(n7551), .B(n7552), .Z(n7546) );
  NANDN U7646 ( .A(n7553), .B(n7554), .Z(n7552) );
  NANDN U7647 ( .A(n7555), .B(n7556), .Z(n7554) );
  NANDN U7648 ( .A(n7556), .B(n7555), .Z(n7551) );
  ANDN U7649 ( .B(B[249]), .A(n29), .Z(n7548) );
  XOR U7650 ( .A(n7515), .B(n7557), .Z(n7549) );
  XNOR U7651 ( .A(n7514), .B(n7512), .Z(n7557) );
  AND U7652 ( .A(n7558), .B(n7559), .Z(n7512) );
  NANDN U7653 ( .A(n7560), .B(n7561), .Z(n7559) );
  OR U7654 ( .A(n7562), .B(n7563), .Z(n7561) );
  NAND U7655 ( .A(n7563), .B(n7562), .Z(n7558) );
  ANDN U7656 ( .B(B[250]), .A(n30), .Z(n7514) );
  XNOR U7657 ( .A(n7522), .B(n7564), .Z(n7515) );
  XNOR U7658 ( .A(n7521), .B(n7519), .Z(n7564) );
  AND U7659 ( .A(n7565), .B(n7566), .Z(n7519) );
  NANDN U7660 ( .A(n7567), .B(n7568), .Z(n7566) );
  NANDN U7661 ( .A(n7569), .B(n7570), .Z(n7568) );
  NANDN U7662 ( .A(n7570), .B(n7569), .Z(n7565) );
  ANDN U7663 ( .B(B[251]), .A(n31), .Z(n7521) );
  XNOR U7664 ( .A(n7529), .B(n7571), .Z(n7522) );
  XNOR U7665 ( .A(n7528), .B(n7526), .Z(n7571) );
  AND U7666 ( .A(n7572), .B(n7573), .Z(n7526) );
  NANDN U7667 ( .A(n7574), .B(n7575), .Z(n7573) );
  OR U7668 ( .A(n7576), .B(n7577), .Z(n7575) );
  NAND U7669 ( .A(n7577), .B(n7576), .Z(n7572) );
  ANDN U7670 ( .B(B[252]), .A(n32), .Z(n7528) );
  XNOR U7671 ( .A(n7536), .B(n7578), .Z(n7529) );
  XNOR U7672 ( .A(n7535), .B(n7533), .Z(n7578) );
  AND U7673 ( .A(n7579), .B(n7580), .Z(n7533) );
  NANDN U7674 ( .A(n7581), .B(n7582), .Z(n7580) );
  NANDN U7675 ( .A(n7583), .B(n7584), .Z(n7582) );
  NANDN U7676 ( .A(n7584), .B(n7583), .Z(n7579) );
  ANDN U7677 ( .B(B[253]), .A(n33), .Z(n7535) );
  XOR U7678 ( .A(n7541), .B(n7585), .Z(n7536) );
  XOR U7679 ( .A(n7542), .B(n7543), .Z(n7585) );
  NAND U7680 ( .A(A[9]), .B(B[255]), .Z(n7543) );
  AND U7681 ( .A(B[254]), .B(A[10]), .Z(n7542) );
  NAND U7682 ( .A(n7586), .B(n7587), .Z(n7541) );
  NAND U7683 ( .A(n7588), .B(n7589), .Z(n7587) );
  NANDN U7684 ( .A(n7590), .B(n7591), .Z(n7588) );
  NANDN U7685 ( .A(n7591), .B(n7590), .Z(n7586) );
  NAND U7686 ( .A(n7592), .B(n7593), .Z(n205) );
  NANDN U7687 ( .A(n7594), .B(n7595), .Z(n7593) );
  OR U7688 ( .A(n7596), .B(n7597), .Z(n7595) );
  NAND U7689 ( .A(n7597), .B(n7596), .Z(n7592) );
  XOR U7690 ( .A(n207), .B(n206), .Z(\A1[261] ) );
  XOR U7691 ( .A(n7597), .B(n7598), .Z(n206) );
  XNOR U7692 ( .A(n7596), .B(n7594), .Z(n7598) );
  AND U7693 ( .A(n7599), .B(n7600), .Z(n7594) );
  NANDN U7694 ( .A(n7601), .B(n7602), .Z(n7600) );
  OR U7695 ( .A(n7603), .B(n7604), .Z(n7602) );
  NAND U7696 ( .A(n7604), .B(n7603), .Z(n7599) );
  ANDN U7697 ( .B(B[248]), .A(n29), .Z(n7596) );
  XNOR U7698 ( .A(n7556), .B(n7605), .Z(n7597) );
  XNOR U7699 ( .A(n7555), .B(n7553), .Z(n7605) );
  AND U7700 ( .A(n7606), .B(n7607), .Z(n7553) );
  NANDN U7701 ( .A(n7608), .B(n7609), .Z(n7607) );
  NANDN U7702 ( .A(n7610), .B(n7611), .Z(n7609) );
  NANDN U7703 ( .A(n7611), .B(n7610), .Z(n7606) );
  ANDN U7704 ( .B(B[249]), .A(n30), .Z(n7555) );
  XNOR U7705 ( .A(n7563), .B(n7612), .Z(n7556) );
  XNOR U7706 ( .A(n7562), .B(n7560), .Z(n7612) );
  AND U7707 ( .A(n7613), .B(n7614), .Z(n7560) );
  NANDN U7708 ( .A(n7615), .B(n7616), .Z(n7614) );
  OR U7709 ( .A(n7617), .B(n7618), .Z(n7616) );
  NAND U7710 ( .A(n7618), .B(n7617), .Z(n7613) );
  ANDN U7711 ( .B(B[250]), .A(n31), .Z(n7562) );
  XNOR U7712 ( .A(n7570), .B(n7619), .Z(n7563) );
  XNOR U7713 ( .A(n7569), .B(n7567), .Z(n7619) );
  AND U7714 ( .A(n7620), .B(n7621), .Z(n7567) );
  NANDN U7715 ( .A(n7622), .B(n7623), .Z(n7621) );
  NANDN U7716 ( .A(n7624), .B(n7625), .Z(n7623) );
  NANDN U7717 ( .A(n7625), .B(n7624), .Z(n7620) );
  ANDN U7718 ( .B(B[251]), .A(n32), .Z(n7569) );
  XNOR U7719 ( .A(n7577), .B(n7626), .Z(n7570) );
  XNOR U7720 ( .A(n7576), .B(n7574), .Z(n7626) );
  AND U7721 ( .A(n7627), .B(n7628), .Z(n7574) );
  NANDN U7722 ( .A(n7629), .B(n7630), .Z(n7628) );
  OR U7723 ( .A(n7631), .B(n7632), .Z(n7630) );
  NAND U7724 ( .A(n7632), .B(n7631), .Z(n7627) );
  ANDN U7725 ( .B(B[252]), .A(n33), .Z(n7576) );
  XNOR U7726 ( .A(n7584), .B(n7633), .Z(n7577) );
  XNOR U7727 ( .A(n7583), .B(n7581), .Z(n7633) );
  AND U7728 ( .A(n7634), .B(n7635), .Z(n7581) );
  NANDN U7729 ( .A(n7636), .B(n7637), .Z(n7635) );
  NANDN U7730 ( .A(n7638), .B(n7639), .Z(n7637) );
  NANDN U7731 ( .A(n7639), .B(n7638), .Z(n7634) );
  ANDN U7732 ( .B(B[253]), .A(n34), .Z(n7583) );
  XOR U7733 ( .A(n7589), .B(n7640), .Z(n7584) );
  XOR U7734 ( .A(n7590), .B(n7591), .Z(n7640) );
  NAND U7735 ( .A(A[8]), .B(B[255]), .Z(n7591) );
  AND U7736 ( .A(B[254]), .B(A[9]), .Z(n7590) );
  NAND U7737 ( .A(n7641), .B(n7642), .Z(n7589) );
  NAND U7738 ( .A(n7643), .B(n7644), .Z(n7642) );
  NANDN U7739 ( .A(n7645), .B(n7646), .Z(n7643) );
  NANDN U7740 ( .A(n7646), .B(n7645), .Z(n7641) );
  NAND U7741 ( .A(n7647), .B(n7648), .Z(n207) );
  NANDN U7742 ( .A(n7649), .B(n7650), .Z(n7648) );
  NAND U7743 ( .A(n7652), .B(n7651), .Z(n7647) );
  XOR U7744 ( .A(n209), .B(n208), .Z(\A1[260] ) );
  XOR U7745 ( .A(n7652), .B(n7653), .Z(n208) );
  XNOR U7746 ( .A(n7651), .B(n7649), .Z(n7653) );
  AND U7747 ( .A(n7654), .B(n7655), .Z(n7649) );
  NANDN U7748 ( .A(n7656), .B(n7657), .Z(n7655) );
  NANDN U7749 ( .A(n7658), .B(n7659), .Z(n7657) );
  NANDN U7750 ( .A(n7659), .B(n7658), .Z(n7654) );
  ANDN U7751 ( .B(B[247]), .A(n29), .Z(n7651) );
  XOR U7752 ( .A(n7604), .B(n7660), .Z(n7652) );
  XNOR U7753 ( .A(n7603), .B(n7601), .Z(n7660) );
  AND U7754 ( .A(n7661), .B(n7662), .Z(n7601) );
  NANDN U7755 ( .A(n7663), .B(n7664), .Z(n7662) );
  OR U7756 ( .A(n7665), .B(n7666), .Z(n7664) );
  NAND U7757 ( .A(n7666), .B(n7665), .Z(n7661) );
  ANDN U7758 ( .B(B[248]), .A(n30), .Z(n7603) );
  XNOR U7759 ( .A(n7611), .B(n7667), .Z(n7604) );
  XNOR U7760 ( .A(n7610), .B(n7608), .Z(n7667) );
  AND U7761 ( .A(n7668), .B(n7669), .Z(n7608) );
  NANDN U7762 ( .A(n7670), .B(n7671), .Z(n7669) );
  NANDN U7763 ( .A(n7672), .B(n7673), .Z(n7671) );
  NANDN U7764 ( .A(n7673), .B(n7672), .Z(n7668) );
  ANDN U7765 ( .B(B[249]), .A(n31), .Z(n7610) );
  XNOR U7766 ( .A(n7618), .B(n7674), .Z(n7611) );
  XNOR U7767 ( .A(n7617), .B(n7615), .Z(n7674) );
  AND U7768 ( .A(n7675), .B(n7676), .Z(n7615) );
  NANDN U7769 ( .A(n7677), .B(n7678), .Z(n7676) );
  OR U7770 ( .A(n7679), .B(n7680), .Z(n7678) );
  NAND U7771 ( .A(n7680), .B(n7679), .Z(n7675) );
  ANDN U7772 ( .B(B[250]), .A(n32), .Z(n7617) );
  XNOR U7773 ( .A(n7625), .B(n7681), .Z(n7618) );
  XNOR U7774 ( .A(n7624), .B(n7622), .Z(n7681) );
  AND U7775 ( .A(n7682), .B(n7683), .Z(n7622) );
  NANDN U7776 ( .A(n7684), .B(n7685), .Z(n7683) );
  NANDN U7777 ( .A(n7686), .B(n7687), .Z(n7685) );
  NANDN U7778 ( .A(n7687), .B(n7686), .Z(n7682) );
  ANDN U7779 ( .B(B[251]), .A(n33), .Z(n7624) );
  XNOR U7780 ( .A(n7632), .B(n7688), .Z(n7625) );
  XNOR U7781 ( .A(n7631), .B(n7629), .Z(n7688) );
  AND U7782 ( .A(n7689), .B(n7690), .Z(n7629) );
  NANDN U7783 ( .A(n7691), .B(n7692), .Z(n7690) );
  OR U7784 ( .A(n7693), .B(n7694), .Z(n7692) );
  NAND U7785 ( .A(n7694), .B(n7693), .Z(n7689) );
  ANDN U7786 ( .B(B[252]), .A(n34), .Z(n7631) );
  XNOR U7787 ( .A(n7639), .B(n7695), .Z(n7632) );
  XNOR U7788 ( .A(n7638), .B(n7636), .Z(n7695) );
  AND U7789 ( .A(n7696), .B(n7697), .Z(n7636) );
  NANDN U7790 ( .A(n7698), .B(n7699), .Z(n7697) );
  NANDN U7791 ( .A(n7700), .B(n7701), .Z(n7699) );
  NANDN U7792 ( .A(n7701), .B(n7700), .Z(n7696) );
  ANDN U7793 ( .B(B[253]), .A(n35), .Z(n7638) );
  XOR U7794 ( .A(n7644), .B(n7702), .Z(n7639) );
  XOR U7795 ( .A(n7645), .B(n7646), .Z(n7702) );
  NAND U7796 ( .A(A[7]), .B(B[255]), .Z(n7646) );
  AND U7797 ( .A(B[254]), .B(A[8]), .Z(n7645) );
  NAND U7798 ( .A(n7703), .B(n7704), .Z(n7644) );
  NAND U7799 ( .A(n7705), .B(n7706), .Z(n7704) );
  NANDN U7800 ( .A(n7707), .B(n7708), .Z(n7705) );
  NANDN U7801 ( .A(n7708), .B(n7707), .Z(n7703) );
  NAND U7802 ( .A(n7709), .B(n7710), .Z(n209) );
  NANDN U7803 ( .A(n7711), .B(n7712), .Z(n7710) );
  OR U7804 ( .A(n7713), .B(n7714), .Z(n7712) );
  NAND U7805 ( .A(n7714), .B(n7713), .Z(n7709) );
  XOR U7806 ( .A(n192), .B(n191), .Z(\A1[25] ) );
  XOR U7807 ( .A(n7407), .B(n7715), .Z(n191) );
  XNOR U7808 ( .A(n7406), .B(n7404), .Z(n7715) );
  AND U7809 ( .A(n7716), .B(n7717), .Z(n7404) );
  NANDN U7810 ( .A(n7718), .B(n7719), .Z(n7717) );
  NANDN U7811 ( .A(n7720), .B(n7721), .Z(n7719) );
  NANDN U7812 ( .A(n7721), .B(n7720), .Z(n7716) );
  ANDN U7813 ( .B(B[12]), .A(n29), .Z(n7406) );
  XNOR U7814 ( .A(n7313), .B(n7722), .Z(n7407) );
  XNOR U7815 ( .A(n7312), .B(n7310), .Z(n7722) );
  AND U7816 ( .A(n7723), .B(n7724), .Z(n7310) );
  NANDN U7817 ( .A(n7725), .B(n7726), .Z(n7724) );
  OR U7818 ( .A(n7727), .B(n7728), .Z(n7726) );
  NAND U7819 ( .A(n7728), .B(n7727), .Z(n7723) );
  ANDN U7820 ( .B(B[13]), .A(n30), .Z(n7312) );
  XNOR U7821 ( .A(n7320), .B(n7729), .Z(n7313) );
  XNOR U7822 ( .A(n7319), .B(n7317), .Z(n7729) );
  AND U7823 ( .A(n7730), .B(n7731), .Z(n7317) );
  NANDN U7824 ( .A(n7732), .B(n7733), .Z(n7731) );
  NANDN U7825 ( .A(n7734), .B(n7735), .Z(n7733) );
  NANDN U7826 ( .A(n7735), .B(n7734), .Z(n7730) );
  ANDN U7827 ( .B(B[14]), .A(n31), .Z(n7319) );
  XNOR U7828 ( .A(n7327), .B(n7736), .Z(n7320) );
  XNOR U7829 ( .A(n7326), .B(n7324), .Z(n7736) );
  AND U7830 ( .A(n7737), .B(n7738), .Z(n7324) );
  NANDN U7831 ( .A(n7739), .B(n7740), .Z(n7738) );
  OR U7832 ( .A(n7741), .B(n7742), .Z(n7740) );
  NAND U7833 ( .A(n7742), .B(n7741), .Z(n7737) );
  ANDN U7834 ( .B(B[15]), .A(n32), .Z(n7326) );
  XNOR U7835 ( .A(n7334), .B(n7743), .Z(n7327) );
  XNOR U7836 ( .A(n7333), .B(n7331), .Z(n7743) );
  AND U7837 ( .A(n7744), .B(n7745), .Z(n7331) );
  NANDN U7838 ( .A(n7746), .B(n7747), .Z(n7745) );
  NANDN U7839 ( .A(n7748), .B(n7749), .Z(n7747) );
  NANDN U7840 ( .A(n7749), .B(n7748), .Z(n7744) );
  ANDN U7841 ( .B(B[16]), .A(n33), .Z(n7333) );
  XNOR U7842 ( .A(n7341), .B(n7750), .Z(n7334) );
  XNOR U7843 ( .A(n7340), .B(n7338), .Z(n7750) );
  AND U7844 ( .A(n7751), .B(n7752), .Z(n7338) );
  NANDN U7845 ( .A(n7753), .B(n7754), .Z(n7752) );
  OR U7846 ( .A(n7755), .B(n7756), .Z(n7754) );
  NAND U7847 ( .A(n7756), .B(n7755), .Z(n7751) );
  ANDN U7848 ( .B(B[17]), .A(n34), .Z(n7340) );
  XNOR U7849 ( .A(n7348), .B(n7757), .Z(n7341) );
  XNOR U7850 ( .A(n7347), .B(n7345), .Z(n7757) );
  AND U7851 ( .A(n7758), .B(n7759), .Z(n7345) );
  NANDN U7852 ( .A(n7760), .B(n7761), .Z(n7759) );
  NANDN U7853 ( .A(n7762), .B(n7763), .Z(n7761) );
  NANDN U7854 ( .A(n7763), .B(n7762), .Z(n7758) );
  ANDN U7855 ( .B(B[18]), .A(n35), .Z(n7347) );
  XNOR U7856 ( .A(n7355), .B(n7764), .Z(n7348) );
  XNOR U7857 ( .A(n7354), .B(n7352), .Z(n7764) );
  AND U7858 ( .A(n7765), .B(n7766), .Z(n7352) );
  NANDN U7859 ( .A(n7767), .B(n7768), .Z(n7766) );
  OR U7860 ( .A(n7769), .B(n7770), .Z(n7768) );
  NAND U7861 ( .A(n7770), .B(n7769), .Z(n7765) );
  ANDN U7862 ( .B(B[19]), .A(n36), .Z(n7354) );
  XNOR U7863 ( .A(n7362), .B(n7771), .Z(n7355) );
  XNOR U7864 ( .A(n7361), .B(n7359), .Z(n7771) );
  AND U7865 ( .A(n7772), .B(n7773), .Z(n7359) );
  NANDN U7866 ( .A(n7774), .B(n7775), .Z(n7773) );
  NANDN U7867 ( .A(n7776), .B(n7777), .Z(n7775) );
  NANDN U7868 ( .A(n7777), .B(n7776), .Z(n7772) );
  ANDN U7869 ( .B(B[20]), .A(n37), .Z(n7361) );
  XNOR U7870 ( .A(n7369), .B(n7778), .Z(n7362) );
  XNOR U7871 ( .A(n7368), .B(n7366), .Z(n7778) );
  AND U7872 ( .A(n7779), .B(n7780), .Z(n7366) );
  NANDN U7873 ( .A(n7781), .B(n7782), .Z(n7780) );
  OR U7874 ( .A(n7783), .B(n7784), .Z(n7782) );
  NAND U7875 ( .A(n7784), .B(n7783), .Z(n7779) );
  ANDN U7876 ( .B(B[21]), .A(n38), .Z(n7368) );
  XNOR U7877 ( .A(n7376), .B(n7785), .Z(n7369) );
  XNOR U7878 ( .A(n7375), .B(n7373), .Z(n7785) );
  AND U7879 ( .A(n7786), .B(n7787), .Z(n7373) );
  NANDN U7880 ( .A(n7788), .B(n7789), .Z(n7787) );
  NANDN U7881 ( .A(n7790), .B(n7791), .Z(n7789) );
  NANDN U7882 ( .A(n7791), .B(n7790), .Z(n7786) );
  ANDN U7883 ( .B(B[22]), .A(n39), .Z(n7375) );
  XNOR U7884 ( .A(n7383), .B(n7792), .Z(n7376) );
  XNOR U7885 ( .A(n7382), .B(n7380), .Z(n7792) );
  AND U7886 ( .A(n7793), .B(n7794), .Z(n7380) );
  NANDN U7887 ( .A(n7795), .B(n7796), .Z(n7794) );
  OR U7888 ( .A(n7797), .B(n7798), .Z(n7796) );
  NAND U7889 ( .A(n7798), .B(n7797), .Z(n7793) );
  ANDN U7890 ( .B(B[23]), .A(n40), .Z(n7382) );
  XNOR U7891 ( .A(n7390), .B(n7799), .Z(n7383) );
  XNOR U7892 ( .A(n7389), .B(n7387), .Z(n7799) );
  AND U7893 ( .A(n7800), .B(n7801), .Z(n7387) );
  NANDN U7894 ( .A(n7802), .B(n7803), .Z(n7801) );
  NAND U7895 ( .A(n7804), .B(n7805), .Z(n7803) );
  ANDN U7896 ( .B(B[24]), .A(n41), .Z(n7389) );
  XOR U7897 ( .A(n7396), .B(n7806), .Z(n7390) );
  XNOR U7898 ( .A(n7394), .B(n7397), .Z(n7806) );
  NAND U7899 ( .A(A[2]), .B(B[25]), .Z(n7397) );
  NANDN U7900 ( .A(n7807), .B(n7808), .Z(n7394) );
  AND U7901 ( .A(A[0]), .B(B[26]), .Z(n7808) );
  XNOR U7902 ( .A(n7399), .B(n7809), .Z(n7396) );
  NAND U7903 ( .A(A[0]), .B(B[27]), .Z(n7809) );
  NAND U7904 ( .A(B[26]), .B(A[1]), .Z(n7399) );
  NAND U7905 ( .A(n7810), .B(n7811), .Z(n192) );
  NANDN U7906 ( .A(n7812), .B(n7813), .Z(n7811) );
  OR U7907 ( .A(n7814), .B(n7815), .Z(n7813) );
  NAND U7908 ( .A(n7815), .B(n7814), .Z(n7810) );
  XOR U7909 ( .A(n211), .B(n210), .Z(\A1[259] ) );
  XOR U7910 ( .A(n7714), .B(n7816), .Z(n210) );
  XNOR U7911 ( .A(n7713), .B(n7711), .Z(n7816) );
  AND U7912 ( .A(n7817), .B(n7818), .Z(n7711) );
  NANDN U7913 ( .A(n7819), .B(n7820), .Z(n7818) );
  OR U7914 ( .A(n7821), .B(n7822), .Z(n7820) );
  NAND U7915 ( .A(n7822), .B(n7821), .Z(n7817) );
  ANDN U7916 ( .B(B[246]), .A(n29), .Z(n7713) );
  XNOR U7917 ( .A(n7659), .B(n7823), .Z(n7714) );
  XNOR U7918 ( .A(n7658), .B(n7656), .Z(n7823) );
  AND U7919 ( .A(n7824), .B(n7825), .Z(n7656) );
  NANDN U7920 ( .A(n7826), .B(n7827), .Z(n7825) );
  NANDN U7921 ( .A(n7828), .B(n7829), .Z(n7827) );
  NANDN U7922 ( .A(n7829), .B(n7828), .Z(n7824) );
  ANDN U7923 ( .B(B[247]), .A(n30), .Z(n7658) );
  XNOR U7924 ( .A(n7666), .B(n7830), .Z(n7659) );
  XNOR U7925 ( .A(n7665), .B(n7663), .Z(n7830) );
  AND U7926 ( .A(n7831), .B(n7832), .Z(n7663) );
  NANDN U7927 ( .A(n7833), .B(n7834), .Z(n7832) );
  OR U7928 ( .A(n7835), .B(n7836), .Z(n7834) );
  NAND U7929 ( .A(n7836), .B(n7835), .Z(n7831) );
  ANDN U7930 ( .B(B[248]), .A(n31), .Z(n7665) );
  XNOR U7931 ( .A(n7673), .B(n7837), .Z(n7666) );
  XNOR U7932 ( .A(n7672), .B(n7670), .Z(n7837) );
  AND U7933 ( .A(n7838), .B(n7839), .Z(n7670) );
  NANDN U7934 ( .A(n7840), .B(n7841), .Z(n7839) );
  NANDN U7935 ( .A(n7842), .B(n7843), .Z(n7841) );
  NANDN U7936 ( .A(n7843), .B(n7842), .Z(n7838) );
  ANDN U7937 ( .B(B[249]), .A(n32), .Z(n7672) );
  XNOR U7938 ( .A(n7680), .B(n7844), .Z(n7673) );
  XNOR U7939 ( .A(n7679), .B(n7677), .Z(n7844) );
  AND U7940 ( .A(n7845), .B(n7846), .Z(n7677) );
  NANDN U7941 ( .A(n7847), .B(n7848), .Z(n7846) );
  OR U7942 ( .A(n7849), .B(n7850), .Z(n7848) );
  NAND U7943 ( .A(n7850), .B(n7849), .Z(n7845) );
  ANDN U7944 ( .B(B[250]), .A(n33), .Z(n7679) );
  XNOR U7945 ( .A(n7687), .B(n7851), .Z(n7680) );
  XNOR U7946 ( .A(n7686), .B(n7684), .Z(n7851) );
  AND U7947 ( .A(n7852), .B(n7853), .Z(n7684) );
  NANDN U7948 ( .A(n7854), .B(n7855), .Z(n7853) );
  NANDN U7949 ( .A(n7856), .B(n7857), .Z(n7855) );
  NANDN U7950 ( .A(n7857), .B(n7856), .Z(n7852) );
  ANDN U7951 ( .B(B[251]), .A(n34), .Z(n7686) );
  XNOR U7952 ( .A(n7694), .B(n7858), .Z(n7687) );
  XNOR U7953 ( .A(n7693), .B(n7691), .Z(n7858) );
  AND U7954 ( .A(n7859), .B(n7860), .Z(n7691) );
  NANDN U7955 ( .A(n7861), .B(n7862), .Z(n7860) );
  OR U7956 ( .A(n7863), .B(n7864), .Z(n7862) );
  NAND U7957 ( .A(n7864), .B(n7863), .Z(n7859) );
  ANDN U7958 ( .B(B[252]), .A(n35), .Z(n7693) );
  XNOR U7959 ( .A(n7701), .B(n7865), .Z(n7694) );
  XNOR U7960 ( .A(n7700), .B(n7698), .Z(n7865) );
  AND U7961 ( .A(n7866), .B(n7867), .Z(n7698) );
  NANDN U7962 ( .A(n7868), .B(n7869), .Z(n7867) );
  NANDN U7963 ( .A(n7870), .B(n7871), .Z(n7869) );
  NANDN U7964 ( .A(n7871), .B(n7870), .Z(n7866) );
  ANDN U7965 ( .B(B[253]), .A(n36), .Z(n7700) );
  XOR U7966 ( .A(n7706), .B(n7872), .Z(n7701) );
  XOR U7967 ( .A(n7707), .B(n7708), .Z(n7872) );
  NAND U7968 ( .A(A[6]), .B(B[255]), .Z(n7708) );
  AND U7969 ( .A(B[254]), .B(A[7]), .Z(n7707) );
  NAND U7970 ( .A(n7873), .B(n7874), .Z(n7706) );
  NAND U7971 ( .A(n7875), .B(n7876), .Z(n7874) );
  NANDN U7972 ( .A(n7877), .B(n7878), .Z(n7875) );
  NANDN U7973 ( .A(n7878), .B(n7877), .Z(n7873) );
  NAND U7974 ( .A(n7879), .B(n7880), .Z(n211) );
  NANDN U7975 ( .A(n7881), .B(n7882), .Z(n7880) );
  NAND U7976 ( .A(n7884), .B(n7883), .Z(n7879) );
  XOR U7977 ( .A(n215), .B(n214), .Z(\A1[258] ) );
  XOR U7978 ( .A(n7884), .B(n7885), .Z(n214) );
  XNOR U7979 ( .A(n7883), .B(n7881), .Z(n7885) );
  AND U7980 ( .A(n7886), .B(n7887), .Z(n7881) );
  NANDN U7981 ( .A(n7888), .B(n7889), .Z(n7887) );
  NANDN U7982 ( .A(n7890), .B(n7891), .Z(n7889) );
  NANDN U7983 ( .A(n7891), .B(n7890), .Z(n7886) );
  ANDN U7984 ( .B(B[245]), .A(n29), .Z(n7883) );
  XOR U7985 ( .A(n7822), .B(n7892), .Z(n7884) );
  XNOR U7986 ( .A(n7821), .B(n7819), .Z(n7892) );
  AND U7987 ( .A(n7893), .B(n7894), .Z(n7819) );
  NANDN U7988 ( .A(n7895), .B(n7896), .Z(n7894) );
  OR U7989 ( .A(n7897), .B(n7898), .Z(n7896) );
  NAND U7990 ( .A(n7898), .B(n7897), .Z(n7893) );
  ANDN U7991 ( .B(B[246]), .A(n30), .Z(n7821) );
  XNOR U7992 ( .A(n7829), .B(n7899), .Z(n7822) );
  XNOR U7993 ( .A(n7828), .B(n7826), .Z(n7899) );
  AND U7994 ( .A(n7900), .B(n7901), .Z(n7826) );
  NANDN U7995 ( .A(n7902), .B(n7903), .Z(n7901) );
  NANDN U7996 ( .A(n7904), .B(n7905), .Z(n7903) );
  NANDN U7997 ( .A(n7905), .B(n7904), .Z(n7900) );
  ANDN U7998 ( .B(B[247]), .A(n31), .Z(n7828) );
  XNOR U7999 ( .A(n7836), .B(n7906), .Z(n7829) );
  XNOR U8000 ( .A(n7835), .B(n7833), .Z(n7906) );
  AND U8001 ( .A(n7907), .B(n7908), .Z(n7833) );
  NANDN U8002 ( .A(n7909), .B(n7910), .Z(n7908) );
  OR U8003 ( .A(n7911), .B(n7912), .Z(n7910) );
  NAND U8004 ( .A(n7912), .B(n7911), .Z(n7907) );
  ANDN U8005 ( .B(B[248]), .A(n32), .Z(n7835) );
  XNOR U8006 ( .A(n7843), .B(n7913), .Z(n7836) );
  XNOR U8007 ( .A(n7842), .B(n7840), .Z(n7913) );
  AND U8008 ( .A(n7914), .B(n7915), .Z(n7840) );
  NANDN U8009 ( .A(n7916), .B(n7917), .Z(n7915) );
  NANDN U8010 ( .A(n7918), .B(n7919), .Z(n7917) );
  NANDN U8011 ( .A(n7919), .B(n7918), .Z(n7914) );
  ANDN U8012 ( .B(B[249]), .A(n33), .Z(n7842) );
  XNOR U8013 ( .A(n7850), .B(n7920), .Z(n7843) );
  XNOR U8014 ( .A(n7849), .B(n7847), .Z(n7920) );
  AND U8015 ( .A(n7921), .B(n7922), .Z(n7847) );
  NANDN U8016 ( .A(n7923), .B(n7924), .Z(n7922) );
  OR U8017 ( .A(n7925), .B(n7926), .Z(n7924) );
  NAND U8018 ( .A(n7926), .B(n7925), .Z(n7921) );
  ANDN U8019 ( .B(B[250]), .A(n34), .Z(n7849) );
  XNOR U8020 ( .A(n7857), .B(n7927), .Z(n7850) );
  XNOR U8021 ( .A(n7856), .B(n7854), .Z(n7927) );
  AND U8022 ( .A(n7928), .B(n7929), .Z(n7854) );
  NANDN U8023 ( .A(n7930), .B(n7931), .Z(n7929) );
  NANDN U8024 ( .A(n7932), .B(n7933), .Z(n7931) );
  NANDN U8025 ( .A(n7933), .B(n7932), .Z(n7928) );
  ANDN U8026 ( .B(B[251]), .A(n35), .Z(n7856) );
  XNOR U8027 ( .A(n7864), .B(n7934), .Z(n7857) );
  XNOR U8028 ( .A(n7863), .B(n7861), .Z(n7934) );
  AND U8029 ( .A(n7935), .B(n7936), .Z(n7861) );
  NANDN U8030 ( .A(n7937), .B(n7938), .Z(n7936) );
  OR U8031 ( .A(n7939), .B(n7940), .Z(n7938) );
  NAND U8032 ( .A(n7940), .B(n7939), .Z(n7935) );
  ANDN U8033 ( .B(B[252]), .A(n36), .Z(n7863) );
  XNOR U8034 ( .A(n7871), .B(n7941), .Z(n7864) );
  XNOR U8035 ( .A(n7870), .B(n7868), .Z(n7941) );
  AND U8036 ( .A(n7942), .B(n7943), .Z(n7868) );
  NANDN U8037 ( .A(n7944), .B(n7945), .Z(n7943) );
  NANDN U8038 ( .A(n7946), .B(n7947), .Z(n7945) );
  NANDN U8039 ( .A(n7947), .B(n7946), .Z(n7942) );
  ANDN U8040 ( .B(B[253]), .A(n37), .Z(n7870) );
  XOR U8041 ( .A(n7876), .B(n7948), .Z(n7871) );
  XOR U8042 ( .A(n7877), .B(n7878), .Z(n7948) );
  NAND U8043 ( .A(A[5]), .B(B[255]), .Z(n7878) );
  AND U8044 ( .A(B[254]), .B(A[6]), .Z(n7877) );
  NAND U8045 ( .A(n7949), .B(n7950), .Z(n7876) );
  NAND U8046 ( .A(n7951), .B(n7952), .Z(n7950) );
  NANDN U8047 ( .A(n7953), .B(n7954), .Z(n7951) );
  NANDN U8048 ( .A(n7954), .B(n7953), .Z(n7949) );
  NAND U8049 ( .A(n7955), .B(n7956), .Z(n215) );
  NANDN U8050 ( .A(n7957), .B(n7958), .Z(n7956) );
  OR U8051 ( .A(n7959), .B(n7960), .Z(n7958) );
  NAND U8052 ( .A(n7960), .B(n7959), .Z(n7955) );
  XOR U8053 ( .A(n217), .B(n216), .Z(\A1[257] ) );
  XOR U8054 ( .A(n7960), .B(n7961), .Z(n216) );
  XNOR U8055 ( .A(n7959), .B(n7957), .Z(n7961) );
  AND U8056 ( .A(n7962), .B(n7963), .Z(n7957) );
  NANDN U8057 ( .A(n7964), .B(n7965), .Z(n7963) );
  OR U8058 ( .A(n7966), .B(n7967), .Z(n7965) );
  NAND U8059 ( .A(n7967), .B(n7966), .Z(n7962) );
  ANDN U8060 ( .B(B[244]), .A(n29), .Z(n7959) );
  XNOR U8061 ( .A(n7891), .B(n7968), .Z(n7960) );
  XNOR U8062 ( .A(n7890), .B(n7888), .Z(n7968) );
  AND U8063 ( .A(n7969), .B(n7970), .Z(n7888) );
  NANDN U8064 ( .A(n7971), .B(n7972), .Z(n7970) );
  NANDN U8065 ( .A(n7973), .B(n7974), .Z(n7972) );
  NANDN U8066 ( .A(n7974), .B(n7973), .Z(n7969) );
  ANDN U8067 ( .B(B[245]), .A(n30), .Z(n7890) );
  XNOR U8068 ( .A(n7898), .B(n7975), .Z(n7891) );
  XNOR U8069 ( .A(n7897), .B(n7895), .Z(n7975) );
  AND U8070 ( .A(n7976), .B(n7977), .Z(n7895) );
  NANDN U8071 ( .A(n7978), .B(n7979), .Z(n7977) );
  OR U8072 ( .A(n7980), .B(n7981), .Z(n7979) );
  NAND U8073 ( .A(n7981), .B(n7980), .Z(n7976) );
  ANDN U8074 ( .B(B[246]), .A(n31), .Z(n7897) );
  XNOR U8075 ( .A(n7905), .B(n7982), .Z(n7898) );
  XNOR U8076 ( .A(n7904), .B(n7902), .Z(n7982) );
  AND U8077 ( .A(n7983), .B(n7984), .Z(n7902) );
  NANDN U8078 ( .A(n7985), .B(n7986), .Z(n7984) );
  NANDN U8079 ( .A(n7987), .B(n7988), .Z(n7986) );
  NANDN U8080 ( .A(n7988), .B(n7987), .Z(n7983) );
  ANDN U8081 ( .B(B[247]), .A(n32), .Z(n7904) );
  XNOR U8082 ( .A(n7912), .B(n7989), .Z(n7905) );
  XNOR U8083 ( .A(n7911), .B(n7909), .Z(n7989) );
  AND U8084 ( .A(n7990), .B(n7991), .Z(n7909) );
  NANDN U8085 ( .A(n7992), .B(n7993), .Z(n7991) );
  OR U8086 ( .A(n7994), .B(n7995), .Z(n7993) );
  NAND U8087 ( .A(n7995), .B(n7994), .Z(n7990) );
  ANDN U8088 ( .B(B[248]), .A(n33), .Z(n7911) );
  XNOR U8089 ( .A(n7919), .B(n7996), .Z(n7912) );
  XNOR U8090 ( .A(n7918), .B(n7916), .Z(n7996) );
  AND U8091 ( .A(n7997), .B(n7998), .Z(n7916) );
  NANDN U8092 ( .A(n7999), .B(n8000), .Z(n7998) );
  NANDN U8093 ( .A(n8001), .B(n8002), .Z(n8000) );
  NANDN U8094 ( .A(n8002), .B(n8001), .Z(n7997) );
  ANDN U8095 ( .B(B[249]), .A(n34), .Z(n7918) );
  XNOR U8096 ( .A(n7926), .B(n8003), .Z(n7919) );
  XNOR U8097 ( .A(n7925), .B(n7923), .Z(n8003) );
  AND U8098 ( .A(n8004), .B(n8005), .Z(n7923) );
  NANDN U8099 ( .A(n8006), .B(n8007), .Z(n8005) );
  OR U8100 ( .A(n8008), .B(n8009), .Z(n8007) );
  NAND U8101 ( .A(n8009), .B(n8008), .Z(n8004) );
  ANDN U8102 ( .B(B[250]), .A(n35), .Z(n7925) );
  XNOR U8103 ( .A(n7933), .B(n8010), .Z(n7926) );
  XNOR U8104 ( .A(n7932), .B(n7930), .Z(n8010) );
  AND U8105 ( .A(n8011), .B(n8012), .Z(n7930) );
  NANDN U8106 ( .A(n8013), .B(n8014), .Z(n8012) );
  NANDN U8107 ( .A(n8015), .B(n8016), .Z(n8014) );
  NANDN U8108 ( .A(n8016), .B(n8015), .Z(n8011) );
  ANDN U8109 ( .B(B[251]), .A(n36), .Z(n7932) );
  XNOR U8110 ( .A(n7940), .B(n8017), .Z(n7933) );
  XNOR U8111 ( .A(n7939), .B(n7937), .Z(n8017) );
  AND U8112 ( .A(n8018), .B(n8019), .Z(n7937) );
  NANDN U8113 ( .A(n8020), .B(n8021), .Z(n8019) );
  OR U8114 ( .A(n8022), .B(n8023), .Z(n8021) );
  NAND U8115 ( .A(n8023), .B(n8022), .Z(n8018) );
  ANDN U8116 ( .B(B[252]), .A(n37), .Z(n7939) );
  XNOR U8117 ( .A(n7947), .B(n8024), .Z(n7940) );
  XNOR U8118 ( .A(n7946), .B(n7944), .Z(n8024) );
  AND U8119 ( .A(n8025), .B(n8026), .Z(n7944) );
  NANDN U8120 ( .A(n8027), .B(n8028), .Z(n8026) );
  NANDN U8121 ( .A(n8029), .B(n8030), .Z(n8028) );
  NANDN U8122 ( .A(n8030), .B(n8029), .Z(n8025) );
  ANDN U8123 ( .B(B[253]), .A(n38), .Z(n7946) );
  XOR U8124 ( .A(n7952), .B(n8031), .Z(n7947) );
  XOR U8125 ( .A(n7953), .B(n7954), .Z(n8031) );
  NAND U8126 ( .A(A[4]), .B(B[255]), .Z(n7954) );
  AND U8127 ( .A(B[254]), .B(A[5]), .Z(n7953) );
  NAND U8128 ( .A(n8032), .B(n8033), .Z(n7952) );
  NAND U8129 ( .A(n8034), .B(n8035), .Z(n8033) );
  NANDN U8130 ( .A(n8036), .B(n8037), .Z(n8034) );
  NANDN U8131 ( .A(n8037), .B(n8036), .Z(n8032) );
  NAND U8132 ( .A(n8038), .B(n8039), .Z(n217) );
  NANDN U8133 ( .A(n8040), .B(n8041), .Z(n8039) );
  NAND U8134 ( .A(n8043), .B(n8042), .Z(n8038) );
  XOR U8135 ( .A(n219), .B(n218), .Z(\A1[256] ) );
  XOR U8136 ( .A(n8043), .B(n8044), .Z(n218) );
  XNOR U8137 ( .A(n8042), .B(n8040), .Z(n8044) );
  AND U8138 ( .A(n8045), .B(n8046), .Z(n8040) );
  NANDN U8139 ( .A(n8047), .B(n8048), .Z(n8046) );
  NANDN U8140 ( .A(n8049), .B(n8050), .Z(n8048) );
  NANDN U8141 ( .A(n8050), .B(n8049), .Z(n8045) );
  ANDN U8142 ( .B(B[243]), .A(n29), .Z(n8042) );
  XOR U8143 ( .A(n7967), .B(n8051), .Z(n8043) );
  XNOR U8144 ( .A(n7966), .B(n7964), .Z(n8051) );
  AND U8145 ( .A(n8052), .B(n8053), .Z(n7964) );
  NANDN U8146 ( .A(n8054), .B(n8055), .Z(n8053) );
  OR U8147 ( .A(n8056), .B(n8057), .Z(n8055) );
  NAND U8148 ( .A(n8057), .B(n8056), .Z(n8052) );
  ANDN U8149 ( .B(B[244]), .A(n30), .Z(n7966) );
  XNOR U8150 ( .A(n7974), .B(n8058), .Z(n7967) );
  XNOR U8151 ( .A(n7973), .B(n7971), .Z(n8058) );
  AND U8152 ( .A(n8059), .B(n8060), .Z(n7971) );
  NANDN U8153 ( .A(n8061), .B(n8062), .Z(n8060) );
  NANDN U8154 ( .A(n8063), .B(n8064), .Z(n8062) );
  NANDN U8155 ( .A(n8064), .B(n8063), .Z(n8059) );
  ANDN U8156 ( .B(B[245]), .A(n31), .Z(n7973) );
  XNOR U8157 ( .A(n7981), .B(n8065), .Z(n7974) );
  XNOR U8158 ( .A(n7980), .B(n7978), .Z(n8065) );
  AND U8159 ( .A(n8066), .B(n8067), .Z(n7978) );
  NANDN U8160 ( .A(n8068), .B(n8069), .Z(n8067) );
  OR U8161 ( .A(n8070), .B(n8071), .Z(n8069) );
  NAND U8162 ( .A(n8071), .B(n8070), .Z(n8066) );
  ANDN U8163 ( .B(B[246]), .A(n32), .Z(n7980) );
  XNOR U8164 ( .A(n7988), .B(n8072), .Z(n7981) );
  XNOR U8165 ( .A(n7987), .B(n7985), .Z(n8072) );
  AND U8166 ( .A(n8073), .B(n8074), .Z(n7985) );
  NANDN U8167 ( .A(n8075), .B(n8076), .Z(n8074) );
  NANDN U8168 ( .A(n8077), .B(n8078), .Z(n8076) );
  NANDN U8169 ( .A(n8078), .B(n8077), .Z(n8073) );
  ANDN U8170 ( .B(B[247]), .A(n33), .Z(n7987) );
  XNOR U8171 ( .A(n7995), .B(n8079), .Z(n7988) );
  XNOR U8172 ( .A(n7994), .B(n7992), .Z(n8079) );
  AND U8173 ( .A(n8080), .B(n8081), .Z(n7992) );
  NANDN U8174 ( .A(n8082), .B(n8083), .Z(n8081) );
  OR U8175 ( .A(n8084), .B(n8085), .Z(n8083) );
  NAND U8176 ( .A(n8085), .B(n8084), .Z(n8080) );
  ANDN U8177 ( .B(B[248]), .A(n34), .Z(n7994) );
  XNOR U8178 ( .A(n8002), .B(n8086), .Z(n7995) );
  XNOR U8179 ( .A(n8001), .B(n7999), .Z(n8086) );
  AND U8180 ( .A(n8087), .B(n8088), .Z(n7999) );
  NANDN U8181 ( .A(n8089), .B(n8090), .Z(n8088) );
  NANDN U8182 ( .A(n8091), .B(n8092), .Z(n8090) );
  NANDN U8183 ( .A(n8092), .B(n8091), .Z(n8087) );
  ANDN U8184 ( .B(B[249]), .A(n35), .Z(n8001) );
  XNOR U8185 ( .A(n8009), .B(n8093), .Z(n8002) );
  XNOR U8186 ( .A(n8008), .B(n8006), .Z(n8093) );
  AND U8187 ( .A(n8094), .B(n8095), .Z(n8006) );
  NANDN U8188 ( .A(n8096), .B(n8097), .Z(n8095) );
  OR U8189 ( .A(n8098), .B(n8099), .Z(n8097) );
  NAND U8190 ( .A(n8099), .B(n8098), .Z(n8094) );
  ANDN U8191 ( .B(B[250]), .A(n36), .Z(n8008) );
  XNOR U8192 ( .A(n8016), .B(n8100), .Z(n8009) );
  XNOR U8193 ( .A(n8015), .B(n8013), .Z(n8100) );
  AND U8194 ( .A(n8101), .B(n8102), .Z(n8013) );
  NANDN U8195 ( .A(n8103), .B(n8104), .Z(n8102) );
  NANDN U8196 ( .A(n8105), .B(n8106), .Z(n8104) );
  NANDN U8197 ( .A(n8106), .B(n8105), .Z(n8101) );
  ANDN U8198 ( .B(B[251]), .A(n37), .Z(n8015) );
  XNOR U8199 ( .A(n8023), .B(n8107), .Z(n8016) );
  XNOR U8200 ( .A(n8022), .B(n8020), .Z(n8107) );
  AND U8201 ( .A(n8108), .B(n8109), .Z(n8020) );
  NANDN U8202 ( .A(n8110), .B(n8111), .Z(n8109) );
  OR U8203 ( .A(n8112), .B(n8113), .Z(n8111) );
  NAND U8204 ( .A(n8113), .B(n8112), .Z(n8108) );
  ANDN U8205 ( .B(B[252]), .A(n38), .Z(n8022) );
  XNOR U8206 ( .A(n8030), .B(n8114), .Z(n8023) );
  XNOR U8207 ( .A(n8029), .B(n8027), .Z(n8114) );
  AND U8208 ( .A(n8115), .B(n8116), .Z(n8027) );
  NANDN U8209 ( .A(n8117), .B(n8118), .Z(n8116) );
  NANDN U8210 ( .A(n8119), .B(n8120), .Z(n8118) );
  NANDN U8211 ( .A(n8120), .B(n8119), .Z(n8115) );
  ANDN U8212 ( .B(B[253]), .A(n39), .Z(n8029) );
  XOR U8213 ( .A(n8035), .B(n8121), .Z(n8030) );
  XOR U8214 ( .A(n8036), .B(n8037), .Z(n8121) );
  NAND U8215 ( .A(A[3]), .B(B[255]), .Z(n8037) );
  AND U8216 ( .A(B[254]), .B(A[4]), .Z(n8036) );
  NAND U8217 ( .A(n8122), .B(n8123), .Z(n8035) );
  NANDN U8218 ( .A(n8125), .B(n8126), .Z(n8124) );
  NANDN U8219 ( .A(n8126), .B(n8125), .Z(n8122) );
  NAND U8220 ( .A(n8128), .B(n8129), .Z(n219) );
  NANDN U8221 ( .A(n8130), .B(n8131), .Z(n8129) );
  OR U8222 ( .A(n8132), .B(n8133), .Z(n8131) );
  NAND U8223 ( .A(n8133), .B(n8132), .Z(n8128) );
  XOR U8224 ( .A(n221), .B(n220), .Z(\A1[255] ) );
  XOR U8225 ( .A(n8133), .B(n8134), .Z(n220) );
  XNOR U8226 ( .A(n8132), .B(n8130), .Z(n8134) );
  AND U8227 ( .A(n8135), .B(n8136), .Z(n8130) );
  NANDN U8228 ( .A(n8137), .B(n8138), .Z(n8136) );
  NANDN U8229 ( .A(n8139), .B(n8140), .Z(n8138) );
  NANDN U8230 ( .A(n8140), .B(n8139), .Z(n8135) );
  ANDN U8231 ( .B(B[242]), .A(n29), .Z(n8132) );
  XNOR U8232 ( .A(n8050), .B(n8141), .Z(n8133) );
  XNOR U8233 ( .A(n8049), .B(n8047), .Z(n8141) );
  AND U8234 ( .A(n8142), .B(n8143), .Z(n8047) );
  NANDN U8235 ( .A(n8144), .B(n8145), .Z(n8143) );
  OR U8236 ( .A(n8146), .B(n8147), .Z(n8145) );
  NAND U8237 ( .A(n8147), .B(n8146), .Z(n8142) );
  ANDN U8238 ( .B(B[243]), .A(n30), .Z(n8049) );
  XNOR U8239 ( .A(n8057), .B(n8148), .Z(n8050) );
  XNOR U8240 ( .A(n8056), .B(n8054), .Z(n8148) );
  AND U8241 ( .A(n8149), .B(n8150), .Z(n8054) );
  NANDN U8242 ( .A(n8151), .B(n8152), .Z(n8150) );
  NANDN U8243 ( .A(n8153), .B(n8154), .Z(n8152) );
  NANDN U8244 ( .A(n8154), .B(n8153), .Z(n8149) );
  ANDN U8245 ( .B(B[244]), .A(n31), .Z(n8056) );
  XNOR U8246 ( .A(n8064), .B(n8155), .Z(n8057) );
  XNOR U8247 ( .A(n8063), .B(n8061), .Z(n8155) );
  AND U8248 ( .A(n8156), .B(n8157), .Z(n8061) );
  NANDN U8249 ( .A(n8158), .B(n8159), .Z(n8157) );
  OR U8250 ( .A(n8160), .B(n8161), .Z(n8159) );
  NAND U8251 ( .A(n8161), .B(n8160), .Z(n8156) );
  ANDN U8252 ( .B(B[245]), .A(n32), .Z(n8063) );
  XNOR U8253 ( .A(n8071), .B(n8162), .Z(n8064) );
  XNOR U8254 ( .A(n8070), .B(n8068), .Z(n8162) );
  AND U8255 ( .A(n8163), .B(n8164), .Z(n8068) );
  NANDN U8256 ( .A(n8165), .B(n8166), .Z(n8164) );
  NANDN U8257 ( .A(n8167), .B(n8168), .Z(n8166) );
  NANDN U8258 ( .A(n8168), .B(n8167), .Z(n8163) );
  ANDN U8259 ( .B(B[246]), .A(n33), .Z(n8070) );
  XNOR U8260 ( .A(n8078), .B(n8169), .Z(n8071) );
  XNOR U8261 ( .A(n8077), .B(n8075), .Z(n8169) );
  AND U8262 ( .A(n8170), .B(n8171), .Z(n8075) );
  NANDN U8263 ( .A(n8172), .B(n8173), .Z(n8171) );
  OR U8264 ( .A(n8174), .B(n8175), .Z(n8173) );
  NAND U8265 ( .A(n8175), .B(n8174), .Z(n8170) );
  ANDN U8266 ( .B(B[247]), .A(n34), .Z(n8077) );
  XNOR U8267 ( .A(n8085), .B(n8176), .Z(n8078) );
  XNOR U8268 ( .A(n8084), .B(n8082), .Z(n8176) );
  AND U8269 ( .A(n8177), .B(n8178), .Z(n8082) );
  NANDN U8270 ( .A(n8179), .B(n8180), .Z(n8178) );
  NANDN U8271 ( .A(n8181), .B(n8182), .Z(n8180) );
  NANDN U8272 ( .A(n8182), .B(n8181), .Z(n8177) );
  ANDN U8273 ( .B(B[248]), .A(n35), .Z(n8084) );
  XNOR U8274 ( .A(n8092), .B(n8183), .Z(n8085) );
  XNOR U8275 ( .A(n8091), .B(n8089), .Z(n8183) );
  AND U8276 ( .A(n8184), .B(n8185), .Z(n8089) );
  NANDN U8277 ( .A(n8186), .B(n8187), .Z(n8185) );
  OR U8278 ( .A(n8188), .B(n8189), .Z(n8187) );
  NAND U8279 ( .A(n8189), .B(n8188), .Z(n8184) );
  ANDN U8280 ( .B(B[249]), .A(n36), .Z(n8091) );
  XNOR U8281 ( .A(n8099), .B(n8190), .Z(n8092) );
  XNOR U8282 ( .A(n8098), .B(n8096), .Z(n8190) );
  AND U8283 ( .A(n8191), .B(n8192), .Z(n8096) );
  NANDN U8284 ( .A(n8193), .B(n8194), .Z(n8192) );
  NANDN U8285 ( .A(n8195), .B(n8196), .Z(n8194) );
  NANDN U8286 ( .A(n8196), .B(n8195), .Z(n8191) );
  ANDN U8287 ( .B(B[250]), .A(n37), .Z(n8098) );
  XNOR U8288 ( .A(n8106), .B(n8197), .Z(n8099) );
  XNOR U8289 ( .A(n8105), .B(n8103), .Z(n8197) );
  AND U8290 ( .A(n8198), .B(n8199), .Z(n8103) );
  NANDN U8291 ( .A(n8200), .B(n8201), .Z(n8199) );
  OR U8292 ( .A(n8202), .B(n8203), .Z(n8201) );
  NAND U8293 ( .A(n8203), .B(n8202), .Z(n8198) );
  ANDN U8294 ( .B(B[251]), .A(n38), .Z(n8105) );
  XNOR U8295 ( .A(n8113), .B(n8204), .Z(n8106) );
  XNOR U8296 ( .A(n8112), .B(n8110), .Z(n8204) );
  AND U8297 ( .A(n8205), .B(n8206), .Z(n8110) );
  NANDN U8298 ( .A(n8207), .B(n8208), .Z(n8206) );
  NANDN U8299 ( .A(n8209), .B(n8210), .Z(n8208) );
  NANDN U8300 ( .A(n8210), .B(n8209), .Z(n8205) );
  ANDN U8301 ( .B(B[252]), .A(n39), .Z(n8112) );
  XNOR U8302 ( .A(n8120), .B(n8211), .Z(n8113) );
  XNOR U8303 ( .A(n8119), .B(n8117), .Z(n8211) );
  AND U8304 ( .A(n8212), .B(n8213), .Z(n8117) );
  NANDN U8305 ( .A(n8214), .B(n8215), .Z(n8213) );
  NANDN U8306 ( .A(n8216), .B(n8217), .Z(n8215) );
  NAND U8307 ( .A(n2), .B(n8216), .Z(n8212) );
  ANDN U8308 ( .B(B[253]), .A(n40), .Z(n8119) );
  XNOR U8309 ( .A(n8127), .B(n8218), .Z(n8120) );
  XOR U8310 ( .A(n8125), .B(n8126), .Z(n8218) );
  NAND U8311 ( .A(B[255]), .B(A[2]), .Z(n8126) );
  AND U8312 ( .A(B[254]), .B(A[3]), .Z(n8125) );
  AND U8313 ( .A(n8219), .B(n8220), .Z(n8127) );
  OR U8314 ( .A(n8221), .B(n8222), .Z(n8219) );
  NAND U8315 ( .A(n8223), .B(n8224), .Z(n221) );
  NANDN U8316 ( .A(n8225), .B(n8226), .Z(n8224) );
  OR U8317 ( .A(n8227), .B(n8228), .Z(n8226) );
  NAND U8318 ( .A(n8228), .B(n8227), .Z(n8223) );
  XOR U8319 ( .A(n223), .B(n222), .Z(\A1[254] ) );
  XOR U8320 ( .A(n8228), .B(n8229), .Z(n222) );
  XNOR U8321 ( .A(n8227), .B(n8225), .Z(n8229) );
  AND U8322 ( .A(n8230), .B(n8231), .Z(n8225) );
  NANDN U8323 ( .A(n8232), .B(n8233), .Z(n8231) );
  NANDN U8324 ( .A(n8234), .B(n8235), .Z(n8233) );
  NANDN U8325 ( .A(n8235), .B(n8234), .Z(n8230) );
  ANDN U8326 ( .B(B[241]), .A(n29), .Z(n8227) );
  XNOR U8327 ( .A(n8140), .B(n8236), .Z(n8228) );
  XNOR U8328 ( .A(n8139), .B(n8137), .Z(n8236) );
  AND U8329 ( .A(n8237), .B(n8238), .Z(n8137) );
  NANDN U8330 ( .A(n8239), .B(n8240), .Z(n8238) );
  OR U8331 ( .A(n8241), .B(n8242), .Z(n8240) );
  NAND U8332 ( .A(n8242), .B(n8241), .Z(n8237) );
  ANDN U8333 ( .B(B[242]), .A(n30), .Z(n8139) );
  XNOR U8334 ( .A(n8147), .B(n8243), .Z(n8140) );
  XNOR U8335 ( .A(n8146), .B(n8144), .Z(n8243) );
  AND U8336 ( .A(n8244), .B(n8245), .Z(n8144) );
  NANDN U8337 ( .A(n8246), .B(n8247), .Z(n8245) );
  NANDN U8338 ( .A(n8248), .B(n8249), .Z(n8247) );
  NANDN U8339 ( .A(n8249), .B(n8248), .Z(n8244) );
  ANDN U8340 ( .B(B[243]), .A(n31), .Z(n8146) );
  XNOR U8341 ( .A(n8154), .B(n8250), .Z(n8147) );
  XNOR U8342 ( .A(n8153), .B(n8151), .Z(n8250) );
  AND U8343 ( .A(n8251), .B(n8252), .Z(n8151) );
  NANDN U8344 ( .A(n8253), .B(n8254), .Z(n8252) );
  OR U8345 ( .A(n8255), .B(n8256), .Z(n8254) );
  NAND U8346 ( .A(n8256), .B(n8255), .Z(n8251) );
  ANDN U8347 ( .B(B[244]), .A(n32), .Z(n8153) );
  XNOR U8348 ( .A(n8161), .B(n8257), .Z(n8154) );
  XNOR U8349 ( .A(n8160), .B(n8158), .Z(n8257) );
  AND U8350 ( .A(n8258), .B(n8259), .Z(n8158) );
  NANDN U8351 ( .A(n8260), .B(n8261), .Z(n8259) );
  NANDN U8352 ( .A(n8262), .B(n8263), .Z(n8261) );
  NANDN U8353 ( .A(n8263), .B(n8262), .Z(n8258) );
  ANDN U8354 ( .B(B[245]), .A(n33), .Z(n8160) );
  XNOR U8355 ( .A(n8168), .B(n8264), .Z(n8161) );
  XNOR U8356 ( .A(n8167), .B(n8165), .Z(n8264) );
  AND U8357 ( .A(n8265), .B(n8266), .Z(n8165) );
  NANDN U8358 ( .A(n8267), .B(n8268), .Z(n8266) );
  OR U8359 ( .A(n8269), .B(n8270), .Z(n8268) );
  NAND U8360 ( .A(n8270), .B(n8269), .Z(n8265) );
  ANDN U8361 ( .B(B[246]), .A(n34), .Z(n8167) );
  XNOR U8362 ( .A(n8175), .B(n8271), .Z(n8168) );
  XNOR U8363 ( .A(n8174), .B(n8172), .Z(n8271) );
  AND U8364 ( .A(n8272), .B(n8273), .Z(n8172) );
  NANDN U8365 ( .A(n8274), .B(n8275), .Z(n8273) );
  NANDN U8366 ( .A(n8276), .B(n8277), .Z(n8275) );
  NANDN U8367 ( .A(n8277), .B(n8276), .Z(n8272) );
  ANDN U8368 ( .B(B[247]), .A(n35), .Z(n8174) );
  XNOR U8369 ( .A(n8182), .B(n8278), .Z(n8175) );
  XNOR U8370 ( .A(n8181), .B(n8179), .Z(n8278) );
  AND U8371 ( .A(n8279), .B(n8280), .Z(n8179) );
  NANDN U8372 ( .A(n8281), .B(n8282), .Z(n8280) );
  OR U8373 ( .A(n8283), .B(n8284), .Z(n8282) );
  NAND U8374 ( .A(n8284), .B(n8283), .Z(n8279) );
  ANDN U8375 ( .B(B[248]), .A(n36), .Z(n8181) );
  XNOR U8376 ( .A(n8189), .B(n8285), .Z(n8182) );
  XNOR U8377 ( .A(n8188), .B(n8186), .Z(n8285) );
  AND U8378 ( .A(n8286), .B(n8287), .Z(n8186) );
  NANDN U8379 ( .A(n8288), .B(n8289), .Z(n8287) );
  NANDN U8380 ( .A(n8290), .B(n8291), .Z(n8289) );
  NANDN U8381 ( .A(n8291), .B(n8290), .Z(n8286) );
  ANDN U8382 ( .B(B[249]), .A(n37), .Z(n8188) );
  XNOR U8383 ( .A(n8196), .B(n8292), .Z(n8189) );
  XNOR U8384 ( .A(n8195), .B(n8193), .Z(n8292) );
  AND U8385 ( .A(n8293), .B(n8294), .Z(n8193) );
  NANDN U8386 ( .A(n8295), .B(n8296), .Z(n8294) );
  OR U8387 ( .A(n8297), .B(n8298), .Z(n8296) );
  NAND U8388 ( .A(n8298), .B(n8297), .Z(n8293) );
  ANDN U8389 ( .B(B[250]), .A(n38), .Z(n8195) );
  XNOR U8390 ( .A(n8203), .B(n8299), .Z(n8196) );
  XNOR U8391 ( .A(n8202), .B(n8200), .Z(n8299) );
  AND U8392 ( .A(n8300), .B(n8301), .Z(n8200) );
  NANDN U8393 ( .A(n8302), .B(n8303), .Z(n8301) );
  NANDN U8394 ( .A(n8304), .B(n8305), .Z(n8303) );
  NANDN U8395 ( .A(n8305), .B(n8304), .Z(n8300) );
  ANDN U8396 ( .B(B[251]), .A(n39), .Z(n8202) );
  XNOR U8397 ( .A(n8210), .B(n8306), .Z(n8203) );
  XNOR U8398 ( .A(n8209), .B(n8207), .Z(n8306) );
  AND U8399 ( .A(n8307), .B(n8308), .Z(n8207) );
  NANDN U8400 ( .A(n8309), .B(n8310), .Z(n8308) );
  OR U8401 ( .A(n8311), .B(n8312), .Z(n8310) );
  NAND U8402 ( .A(n8312), .B(n8311), .Z(n8307) );
  ANDN U8403 ( .B(B[252]), .A(n40), .Z(n8209) );
  XNOR U8404 ( .A(n2), .B(n8313), .Z(n8210) );
  XNOR U8405 ( .A(n8216), .B(n8214), .Z(n8313) );
  AND U8406 ( .A(n8314), .B(n8315), .Z(n8214) );
  NANDN U8407 ( .A(n8316), .B(n8317), .Z(n8315) );
  NAND U8408 ( .A(n8318), .B(n8319), .Z(n8317) );
  ANDN U8409 ( .B(B[253]), .A(n41), .Z(n8216) );
  XNOR U8410 ( .A(n8222), .B(n8320), .Z(n8217) );
  XNOR U8411 ( .A(n8220), .B(n8221), .Z(n8320) );
  NAND U8412 ( .A(A[2]), .B(B[254]), .Z(n8221) );
  ANDN U8413 ( .B(A[0]), .A(n8322), .Z(n8321) );
  NAND U8414 ( .A(B[255]), .B(A[1]), .Z(n8222) );
  NAND U8415 ( .A(n8323), .B(n8324), .Z(n223) );
  NANDN U8416 ( .A(n8325), .B(n8326), .Z(n8324) );
  OR U8417 ( .A(n8327), .B(n8328), .Z(n8326) );
  NAND U8418 ( .A(n8328), .B(n8327), .Z(n8323) );
  XOR U8419 ( .A(n225), .B(n224), .Z(\A1[253] ) );
  XOR U8420 ( .A(n8328), .B(n8329), .Z(n224) );
  XNOR U8421 ( .A(n8327), .B(n8325), .Z(n8329) );
  AND U8422 ( .A(n8330), .B(n8331), .Z(n8325) );
  NANDN U8423 ( .A(n8332), .B(n8333), .Z(n8331) );
  NANDN U8424 ( .A(n8334), .B(n8335), .Z(n8333) );
  NANDN U8425 ( .A(n8335), .B(n8334), .Z(n8330) );
  ANDN U8426 ( .B(B[240]), .A(n29), .Z(n8327) );
  XNOR U8427 ( .A(n8235), .B(n8336), .Z(n8328) );
  XNOR U8428 ( .A(n8234), .B(n8232), .Z(n8336) );
  AND U8429 ( .A(n8337), .B(n8338), .Z(n8232) );
  NANDN U8430 ( .A(n8339), .B(n8340), .Z(n8338) );
  OR U8431 ( .A(n8341), .B(n8342), .Z(n8340) );
  NAND U8432 ( .A(n8342), .B(n8341), .Z(n8337) );
  ANDN U8433 ( .B(B[241]), .A(n30), .Z(n8234) );
  XNOR U8434 ( .A(n8242), .B(n8343), .Z(n8235) );
  XNOR U8435 ( .A(n8241), .B(n8239), .Z(n8343) );
  AND U8436 ( .A(n8344), .B(n8345), .Z(n8239) );
  NANDN U8437 ( .A(n8346), .B(n8347), .Z(n8345) );
  NANDN U8438 ( .A(n8348), .B(n8349), .Z(n8347) );
  NANDN U8439 ( .A(n8349), .B(n8348), .Z(n8344) );
  ANDN U8440 ( .B(B[242]), .A(n31), .Z(n8241) );
  XNOR U8441 ( .A(n8249), .B(n8350), .Z(n8242) );
  XNOR U8442 ( .A(n8248), .B(n8246), .Z(n8350) );
  AND U8443 ( .A(n8351), .B(n8352), .Z(n8246) );
  NANDN U8444 ( .A(n8353), .B(n8354), .Z(n8352) );
  OR U8445 ( .A(n8355), .B(n8356), .Z(n8354) );
  NAND U8446 ( .A(n8356), .B(n8355), .Z(n8351) );
  ANDN U8447 ( .B(B[243]), .A(n32), .Z(n8248) );
  XNOR U8448 ( .A(n8256), .B(n8357), .Z(n8249) );
  XNOR U8449 ( .A(n8255), .B(n8253), .Z(n8357) );
  AND U8450 ( .A(n8358), .B(n8359), .Z(n8253) );
  NANDN U8451 ( .A(n8360), .B(n8361), .Z(n8359) );
  NANDN U8452 ( .A(n8362), .B(n8363), .Z(n8361) );
  NANDN U8453 ( .A(n8363), .B(n8362), .Z(n8358) );
  ANDN U8454 ( .B(B[244]), .A(n33), .Z(n8255) );
  XNOR U8455 ( .A(n8263), .B(n8364), .Z(n8256) );
  XNOR U8456 ( .A(n8262), .B(n8260), .Z(n8364) );
  AND U8457 ( .A(n8365), .B(n8366), .Z(n8260) );
  NANDN U8458 ( .A(n8367), .B(n8368), .Z(n8366) );
  OR U8459 ( .A(n8369), .B(n8370), .Z(n8368) );
  NAND U8460 ( .A(n8370), .B(n8369), .Z(n8365) );
  ANDN U8461 ( .B(B[245]), .A(n34), .Z(n8262) );
  XNOR U8462 ( .A(n8270), .B(n8371), .Z(n8263) );
  XNOR U8463 ( .A(n8269), .B(n8267), .Z(n8371) );
  AND U8464 ( .A(n8372), .B(n8373), .Z(n8267) );
  NANDN U8465 ( .A(n8374), .B(n8375), .Z(n8373) );
  NANDN U8466 ( .A(n8376), .B(n8377), .Z(n8375) );
  NANDN U8467 ( .A(n8377), .B(n8376), .Z(n8372) );
  ANDN U8468 ( .B(B[246]), .A(n35), .Z(n8269) );
  XNOR U8469 ( .A(n8277), .B(n8378), .Z(n8270) );
  XNOR U8470 ( .A(n8276), .B(n8274), .Z(n8378) );
  AND U8471 ( .A(n8379), .B(n8380), .Z(n8274) );
  NANDN U8472 ( .A(n8381), .B(n8382), .Z(n8380) );
  OR U8473 ( .A(n8383), .B(n8384), .Z(n8382) );
  NAND U8474 ( .A(n8384), .B(n8383), .Z(n8379) );
  ANDN U8475 ( .B(B[247]), .A(n36), .Z(n8276) );
  XNOR U8476 ( .A(n8284), .B(n8385), .Z(n8277) );
  XNOR U8477 ( .A(n8283), .B(n8281), .Z(n8385) );
  AND U8478 ( .A(n8386), .B(n8387), .Z(n8281) );
  NANDN U8479 ( .A(n8388), .B(n8389), .Z(n8387) );
  NANDN U8480 ( .A(n8390), .B(n8391), .Z(n8389) );
  NANDN U8481 ( .A(n8391), .B(n8390), .Z(n8386) );
  ANDN U8482 ( .B(B[248]), .A(n37), .Z(n8283) );
  XNOR U8483 ( .A(n8291), .B(n8392), .Z(n8284) );
  XNOR U8484 ( .A(n8290), .B(n8288), .Z(n8392) );
  AND U8485 ( .A(n8393), .B(n8394), .Z(n8288) );
  NANDN U8486 ( .A(n8395), .B(n8396), .Z(n8394) );
  OR U8487 ( .A(n8397), .B(n8398), .Z(n8396) );
  NAND U8488 ( .A(n8398), .B(n8397), .Z(n8393) );
  ANDN U8489 ( .B(B[249]), .A(n38), .Z(n8290) );
  XNOR U8490 ( .A(n8298), .B(n8399), .Z(n8291) );
  XNOR U8491 ( .A(n8297), .B(n8295), .Z(n8399) );
  AND U8492 ( .A(n8400), .B(n8401), .Z(n8295) );
  NANDN U8493 ( .A(n8402), .B(n8403), .Z(n8401) );
  NANDN U8494 ( .A(n8404), .B(n8405), .Z(n8403) );
  NANDN U8495 ( .A(n8405), .B(n8404), .Z(n8400) );
  ANDN U8496 ( .B(B[250]), .A(n39), .Z(n8297) );
  XNOR U8497 ( .A(n8305), .B(n8406), .Z(n8298) );
  XNOR U8498 ( .A(n8304), .B(n8302), .Z(n8406) );
  AND U8499 ( .A(n8407), .B(n8408), .Z(n8302) );
  NANDN U8500 ( .A(n8409), .B(n8410), .Z(n8408) );
  OR U8501 ( .A(n8411), .B(n8412), .Z(n8410) );
  NAND U8502 ( .A(n8412), .B(n8411), .Z(n8407) );
  ANDN U8503 ( .B(B[251]), .A(n40), .Z(n8304) );
  XNOR U8504 ( .A(n8312), .B(n8413), .Z(n8305) );
  XNOR U8505 ( .A(n8311), .B(n8309), .Z(n8413) );
  AND U8506 ( .A(n8414), .B(n8415), .Z(n8309) );
  NANDN U8507 ( .A(n8416), .B(n8417), .Z(n8415) );
  NAND U8508 ( .A(n8418), .B(n8419), .Z(n8417) );
  ANDN U8509 ( .B(B[252]), .A(n41), .Z(n8311) );
  XOR U8510 ( .A(n8318), .B(n8420), .Z(n8312) );
  XNOR U8511 ( .A(n8316), .B(n8319), .Z(n8420) );
  NAND U8512 ( .A(A[2]), .B(B[253]), .Z(n8319) );
  NANDN U8513 ( .A(n8421), .B(n8422), .Z(n8316) );
  AND U8514 ( .A(A[0]), .B(B[254]), .Z(n8422) );
  XNOR U8515 ( .A(n8322), .B(n8423), .Z(n8318) );
  NAND U8516 ( .A(B[255]), .B(A[0]), .Z(n8423) );
  NAND U8517 ( .A(B[254]), .B(A[1]), .Z(n8322) );
  NAND U8518 ( .A(n8424), .B(n8425), .Z(n225) );
  NANDN U8519 ( .A(n8426), .B(n8427), .Z(n8425) );
  OR U8520 ( .A(n8428), .B(n8429), .Z(n8427) );
  NAND U8521 ( .A(n8429), .B(n8428), .Z(n8424) );
  XOR U8522 ( .A(n227), .B(n226), .Z(\A1[252] ) );
  XOR U8523 ( .A(n8429), .B(n8430), .Z(n226) );
  XNOR U8524 ( .A(n8428), .B(n8426), .Z(n8430) );
  AND U8525 ( .A(n8431), .B(n8432), .Z(n8426) );
  NANDN U8526 ( .A(n8433), .B(n8434), .Z(n8432) );
  NANDN U8527 ( .A(n8435), .B(n8436), .Z(n8434) );
  NANDN U8528 ( .A(n8436), .B(n8435), .Z(n8431) );
  ANDN U8529 ( .B(B[239]), .A(n29), .Z(n8428) );
  XNOR U8530 ( .A(n8335), .B(n8437), .Z(n8429) );
  XNOR U8531 ( .A(n8334), .B(n8332), .Z(n8437) );
  AND U8532 ( .A(n8438), .B(n8439), .Z(n8332) );
  NANDN U8533 ( .A(n8440), .B(n8441), .Z(n8439) );
  OR U8534 ( .A(n8442), .B(n8443), .Z(n8441) );
  NAND U8535 ( .A(n8443), .B(n8442), .Z(n8438) );
  ANDN U8536 ( .B(B[240]), .A(n30), .Z(n8334) );
  XNOR U8537 ( .A(n8342), .B(n8444), .Z(n8335) );
  XNOR U8538 ( .A(n8341), .B(n8339), .Z(n8444) );
  AND U8539 ( .A(n8445), .B(n8446), .Z(n8339) );
  NANDN U8540 ( .A(n8447), .B(n8448), .Z(n8446) );
  NANDN U8541 ( .A(n8449), .B(n8450), .Z(n8448) );
  NANDN U8542 ( .A(n8450), .B(n8449), .Z(n8445) );
  ANDN U8543 ( .B(B[241]), .A(n31), .Z(n8341) );
  XNOR U8544 ( .A(n8349), .B(n8451), .Z(n8342) );
  XNOR U8545 ( .A(n8348), .B(n8346), .Z(n8451) );
  AND U8546 ( .A(n8452), .B(n8453), .Z(n8346) );
  NANDN U8547 ( .A(n8454), .B(n8455), .Z(n8453) );
  OR U8548 ( .A(n8456), .B(n8457), .Z(n8455) );
  NAND U8549 ( .A(n8457), .B(n8456), .Z(n8452) );
  ANDN U8550 ( .B(B[242]), .A(n32), .Z(n8348) );
  XNOR U8551 ( .A(n8356), .B(n8458), .Z(n8349) );
  XNOR U8552 ( .A(n8355), .B(n8353), .Z(n8458) );
  AND U8553 ( .A(n8459), .B(n8460), .Z(n8353) );
  NANDN U8554 ( .A(n8461), .B(n8462), .Z(n8460) );
  NANDN U8555 ( .A(n8463), .B(n8464), .Z(n8462) );
  NANDN U8556 ( .A(n8464), .B(n8463), .Z(n8459) );
  ANDN U8557 ( .B(B[243]), .A(n33), .Z(n8355) );
  XNOR U8558 ( .A(n8363), .B(n8465), .Z(n8356) );
  XNOR U8559 ( .A(n8362), .B(n8360), .Z(n8465) );
  AND U8560 ( .A(n8466), .B(n8467), .Z(n8360) );
  NANDN U8561 ( .A(n8468), .B(n8469), .Z(n8467) );
  OR U8562 ( .A(n8470), .B(n8471), .Z(n8469) );
  NAND U8563 ( .A(n8471), .B(n8470), .Z(n8466) );
  ANDN U8564 ( .B(B[244]), .A(n34), .Z(n8362) );
  XNOR U8565 ( .A(n8370), .B(n8472), .Z(n8363) );
  XNOR U8566 ( .A(n8369), .B(n8367), .Z(n8472) );
  AND U8567 ( .A(n8473), .B(n8474), .Z(n8367) );
  NANDN U8568 ( .A(n8475), .B(n8476), .Z(n8474) );
  NANDN U8569 ( .A(n8477), .B(n8478), .Z(n8476) );
  NANDN U8570 ( .A(n8478), .B(n8477), .Z(n8473) );
  ANDN U8571 ( .B(B[245]), .A(n35), .Z(n8369) );
  XNOR U8572 ( .A(n8377), .B(n8479), .Z(n8370) );
  XNOR U8573 ( .A(n8376), .B(n8374), .Z(n8479) );
  AND U8574 ( .A(n8480), .B(n8481), .Z(n8374) );
  NANDN U8575 ( .A(n8482), .B(n8483), .Z(n8481) );
  OR U8576 ( .A(n8484), .B(n8485), .Z(n8483) );
  NAND U8577 ( .A(n8485), .B(n8484), .Z(n8480) );
  ANDN U8578 ( .B(B[246]), .A(n36), .Z(n8376) );
  XNOR U8579 ( .A(n8384), .B(n8486), .Z(n8377) );
  XNOR U8580 ( .A(n8383), .B(n8381), .Z(n8486) );
  AND U8581 ( .A(n8487), .B(n8488), .Z(n8381) );
  NANDN U8582 ( .A(n8489), .B(n8490), .Z(n8488) );
  NANDN U8583 ( .A(n8491), .B(n8492), .Z(n8490) );
  NANDN U8584 ( .A(n8492), .B(n8491), .Z(n8487) );
  ANDN U8585 ( .B(B[247]), .A(n37), .Z(n8383) );
  XNOR U8586 ( .A(n8391), .B(n8493), .Z(n8384) );
  XNOR U8587 ( .A(n8390), .B(n8388), .Z(n8493) );
  AND U8588 ( .A(n8494), .B(n8495), .Z(n8388) );
  NANDN U8589 ( .A(n8496), .B(n8497), .Z(n8495) );
  OR U8590 ( .A(n8498), .B(n8499), .Z(n8497) );
  NAND U8591 ( .A(n8499), .B(n8498), .Z(n8494) );
  ANDN U8592 ( .B(B[248]), .A(n38), .Z(n8390) );
  XNOR U8593 ( .A(n8398), .B(n8500), .Z(n8391) );
  XNOR U8594 ( .A(n8397), .B(n8395), .Z(n8500) );
  AND U8595 ( .A(n8501), .B(n8502), .Z(n8395) );
  NANDN U8596 ( .A(n8503), .B(n8504), .Z(n8502) );
  NANDN U8597 ( .A(n8505), .B(n8506), .Z(n8504) );
  NANDN U8598 ( .A(n8506), .B(n8505), .Z(n8501) );
  ANDN U8599 ( .B(B[249]), .A(n39), .Z(n8397) );
  XNOR U8600 ( .A(n8405), .B(n8507), .Z(n8398) );
  XNOR U8601 ( .A(n8404), .B(n8402), .Z(n8507) );
  AND U8602 ( .A(n8508), .B(n8509), .Z(n8402) );
  NANDN U8603 ( .A(n8510), .B(n8511), .Z(n8509) );
  OR U8604 ( .A(n8512), .B(n8513), .Z(n8511) );
  NAND U8605 ( .A(n8513), .B(n8512), .Z(n8508) );
  ANDN U8606 ( .B(B[250]), .A(n40), .Z(n8404) );
  XNOR U8607 ( .A(n8412), .B(n8514), .Z(n8405) );
  XNOR U8608 ( .A(n8411), .B(n8409), .Z(n8514) );
  AND U8609 ( .A(n8515), .B(n8516), .Z(n8409) );
  NANDN U8610 ( .A(n8517), .B(n8518), .Z(n8516) );
  NAND U8611 ( .A(n8519), .B(n8520), .Z(n8518) );
  ANDN U8612 ( .B(B[251]), .A(n41), .Z(n8411) );
  XOR U8613 ( .A(n8418), .B(n8521), .Z(n8412) );
  XNOR U8614 ( .A(n8416), .B(n8419), .Z(n8521) );
  NAND U8615 ( .A(A[2]), .B(B[252]), .Z(n8419) );
  NANDN U8616 ( .A(n8522), .B(n8523), .Z(n8416) );
  AND U8617 ( .A(A[0]), .B(B[253]), .Z(n8523) );
  XNOR U8618 ( .A(n8421), .B(n8524), .Z(n8418) );
  NAND U8619 ( .A(A[0]), .B(B[254]), .Z(n8524) );
  NAND U8620 ( .A(B[253]), .B(A[1]), .Z(n8421) );
  NAND U8621 ( .A(n8525), .B(n8526), .Z(n227) );
  NANDN U8622 ( .A(n8527), .B(n8528), .Z(n8526) );
  OR U8623 ( .A(n8529), .B(n8530), .Z(n8528) );
  NAND U8624 ( .A(n8530), .B(n8529), .Z(n8525) );
  XOR U8625 ( .A(n229), .B(n228), .Z(\A1[251] ) );
  XOR U8626 ( .A(n8530), .B(n8531), .Z(n228) );
  XNOR U8627 ( .A(n8529), .B(n8527), .Z(n8531) );
  AND U8628 ( .A(n8532), .B(n8533), .Z(n8527) );
  NANDN U8629 ( .A(n8534), .B(n8535), .Z(n8533) );
  NANDN U8630 ( .A(n8536), .B(n8537), .Z(n8535) );
  NANDN U8631 ( .A(n8537), .B(n8536), .Z(n8532) );
  ANDN U8632 ( .B(B[238]), .A(n29), .Z(n8529) );
  XNOR U8633 ( .A(n8436), .B(n8538), .Z(n8530) );
  XNOR U8634 ( .A(n8435), .B(n8433), .Z(n8538) );
  AND U8635 ( .A(n8539), .B(n8540), .Z(n8433) );
  NANDN U8636 ( .A(n8541), .B(n8542), .Z(n8540) );
  OR U8637 ( .A(n8543), .B(n8544), .Z(n8542) );
  NAND U8638 ( .A(n8544), .B(n8543), .Z(n8539) );
  ANDN U8639 ( .B(B[239]), .A(n30), .Z(n8435) );
  XNOR U8640 ( .A(n8443), .B(n8545), .Z(n8436) );
  XNOR U8641 ( .A(n8442), .B(n8440), .Z(n8545) );
  AND U8642 ( .A(n8546), .B(n8547), .Z(n8440) );
  NANDN U8643 ( .A(n8548), .B(n8549), .Z(n8547) );
  NANDN U8644 ( .A(n8550), .B(n8551), .Z(n8549) );
  NANDN U8645 ( .A(n8551), .B(n8550), .Z(n8546) );
  ANDN U8646 ( .B(B[240]), .A(n31), .Z(n8442) );
  XNOR U8647 ( .A(n8450), .B(n8552), .Z(n8443) );
  XNOR U8648 ( .A(n8449), .B(n8447), .Z(n8552) );
  AND U8649 ( .A(n8553), .B(n8554), .Z(n8447) );
  NANDN U8650 ( .A(n8555), .B(n8556), .Z(n8554) );
  OR U8651 ( .A(n8557), .B(n8558), .Z(n8556) );
  NAND U8652 ( .A(n8558), .B(n8557), .Z(n8553) );
  ANDN U8653 ( .B(B[241]), .A(n32), .Z(n8449) );
  XNOR U8654 ( .A(n8457), .B(n8559), .Z(n8450) );
  XNOR U8655 ( .A(n8456), .B(n8454), .Z(n8559) );
  AND U8656 ( .A(n8560), .B(n8561), .Z(n8454) );
  NANDN U8657 ( .A(n8562), .B(n8563), .Z(n8561) );
  NANDN U8658 ( .A(n8564), .B(n8565), .Z(n8563) );
  NANDN U8659 ( .A(n8565), .B(n8564), .Z(n8560) );
  ANDN U8660 ( .B(B[242]), .A(n33), .Z(n8456) );
  XNOR U8661 ( .A(n8464), .B(n8566), .Z(n8457) );
  XNOR U8662 ( .A(n8463), .B(n8461), .Z(n8566) );
  AND U8663 ( .A(n8567), .B(n8568), .Z(n8461) );
  NANDN U8664 ( .A(n8569), .B(n8570), .Z(n8568) );
  OR U8665 ( .A(n8571), .B(n8572), .Z(n8570) );
  NAND U8666 ( .A(n8572), .B(n8571), .Z(n8567) );
  ANDN U8667 ( .B(B[243]), .A(n34), .Z(n8463) );
  XNOR U8668 ( .A(n8471), .B(n8573), .Z(n8464) );
  XNOR U8669 ( .A(n8470), .B(n8468), .Z(n8573) );
  AND U8670 ( .A(n8574), .B(n8575), .Z(n8468) );
  NANDN U8671 ( .A(n8576), .B(n8577), .Z(n8575) );
  NANDN U8672 ( .A(n8578), .B(n8579), .Z(n8577) );
  NANDN U8673 ( .A(n8579), .B(n8578), .Z(n8574) );
  ANDN U8674 ( .B(B[244]), .A(n35), .Z(n8470) );
  XNOR U8675 ( .A(n8478), .B(n8580), .Z(n8471) );
  XNOR U8676 ( .A(n8477), .B(n8475), .Z(n8580) );
  AND U8677 ( .A(n8581), .B(n8582), .Z(n8475) );
  NANDN U8678 ( .A(n8583), .B(n8584), .Z(n8582) );
  OR U8679 ( .A(n8585), .B(n8586), .Z(n8584) );
  NAND U8680 ( .A(n8586), .B(n8585), .Z(n8581) );
  ANDN U8681 ( .B(B[245]), .A(n36), .Z(n8477) );
  XNOR U8682 ( .A(n8485), .B(n8587), .Z(n8478) );
  XNOR U8683 ( .A(n8484), .B(n8482), .Z(n8587) );
  AND U8684 ( .A(n8588), .B(n8589), .Z(n8482) );
  NANDN U8685 ( .A(n8590), .B(n8591), .Z(n8589) );
  NANDN U8686 ( .A(n8592), .B(n8593), .Z(n8591) );
  NANDN U8687 ( .A(n8593), .B(n8592), .Z(n8588) );
  ANDN U8688 ( .B(B[246]), .A(n37), .Z(n8484) );
  XNOR U8689 ( .A(n8492), .B(n8594), .Z(n8485) );
  XNOR U8690 ( .A(n8491), .B(n8489), .Z(n8594) );
  AND U8691 ( .A(n8595), .B(n8596), .Z(n8489) );
  NANDN U8692 ( .A(n8597), .B(n8598), .Z(n8596) );
  OR U8693 ( .A(n8599), .B(n8600), .Z(n8598) );
  NAND U8694 ( .A(n8600), .B(n8599), .Z(n8595) );
  ANDN U8695 ( .B(B[247]), .A(n38), .Z(n8491) );
  XNOR U8696 ( .A(n8499), .B(n8601), .Z(n8492) );
  XNOR U8697 ( .A(n8498), .B(n8496), .Z(n8601) );
  AND U8698 ( .A(n8602), .B(n8603), .Z(n8496) );
  NANDN U8699 ( .A(n8604), .B(n8605), .Z(n8603) );
  NANDN U8700 ( .A(n8606), .B(n8607), .Z(n8605) );
  NANDN U8701 ( .A(n8607), .B(n8606), .Z(n8602) );
  ANDN U8702 ( .B(B[248]), .A(n39), .Z(n8498) );
  XNOR U8703 ( .A(n8506), .B(n8608), .Z(n8499) );
  XNOR U8704 ( .A(n8505), .B(n8503), .Z(n8608) );
  AND U8705 ( .A(n8609), .B(n8610), .Z(n8503) );
  NANDN U8706 ( .A(n8611), .B(n8612), .Z(n8610) );
  OR U8707 ( .A(n8613), .B(n8614), .Z(n8612) );
  NAND U8708 ( .A(n8614), .B(n8613), .Z(n8609) );
  ANDN U8709 ( .B(B[249]), .A(n40), .Z(n8505) );
  XNOR U8710 ( .A(n8513), .B(n8615), .Z(n8506) );
  XNOR U8711 ( .A(n8512), .B(n8510), .Z(n8615) );
  AND U8712 ( .A(n8616), .B(n8617), .Z(n8510) );
  NANDN U8713 ( .A(n8618), .B(n8619), .Z(n8617) );
  NAND U8714 ( .A(n8620), .B(n8621), .Z(n8619) );
  ANDN U8715 ( .B(B[250]), .A(n41), .Z(n8512) );
  XOR U8716 ( .A(n8519), .B(n8622), .Z(n8513) );
  XNOR U8717 ( .A(n8517), .B(n8520), .Z(n8622) );
  NAND U8718 ( .A(A[2]), .B(B[251]), .Z(n8520) );
  NANDN U8719 ( .A(n8623), .B(n8624), .Z(n8517) );
  AND U8720 ( .A(A[0]), .B(B[252]), .Z(n8624) );
  XNOR U8721 ( .A(n8522), .B(n8625), .Z(n8519) );
  NAND U8722 ( .A(A[0]), .B(B[253]), .Z(n8625) );
  NAND U8723 ( .A(B[252]), .B(A[1]), .Z(n8522) );
  NAND U8724 ( .A(n8626), .B(n8627), .Z(n229) );
  NANDN U8725 ( .A(n8628), .B(n8629), .Z(n8627) );
  OR U8726 ( .A(n8630), .B(n8631), .Z(n8629) );
  NAND U8727 ( .A(n8631), .B(n8630), .Z(n8626) );
  XOR U8728 ( .A(n231), .B(n230), .Z(\A1[250] ) );
  XOR U8729 ( .A(n8631), .B(n8632), .Z(n230) );
  XNOR U8730 ( .A(n8630), .B(n8628), .Z(n8632) );
  AND U8731 ( .A(n8633), .B(n8634), .Z(n8628) );
  NANDN U8732 ( .A(n8635), .B(n8636), .Z(n8634) );
  NANDN U8733 ( .A(n8637), .B(n8638), .Z(n8636) );
  NANDN U8734 ( .A(n8638), .B(n8637), .Z(n8633) );
  ANDN U8735 ( .B(B[237]), .A(n29), .Z(n8630) );
  XNOR U8736 ( .A(n8537), .B(n8639), .Z(n8631) );
  XNOR U8737 ( .A(n8536), .B(n8534), .Z(n8639) );
  AND U8738 ( .A(n8640), .B(n8641), .Z(n8534) );
  NANDN U8739 ( .A(n8642), .B(n8643), .Z(n8641) );
  OR U8740 ( .A(n8644), .B(n8645), .Z(n8643) );
  NAND U8741 ( .A(n8645), .B(n8644), .Z(n8640) );
  ANDN U8742 ( .B(B[238]), .A(n30), .Z(n8536) );
  XNOR U8743 ( .A(n8544), .B(n8646), .Z(n8537) );
  XNOR U8744 ( .A(n8543), .B(n8541), .Z(n8646) );
  AND U8745 ( .A(n8647), .B(n8648), .Z(n8541) );
  NANDN U8746 ( .A(n8649), .B(n8650), .Z(n8648) );
  NANDN U8747 ( .A(n8651), .B(n8652), .Z(n8650) );
  NANDN U8748 ( .A(n8652), .B(n8651), .Z(n8647) );
  ANDN U8749 ( .B(B[239]), .A(n31), .Z(n8543) );
  XNOR U8750 ( .A(n8551), .B(n8653), .Z(n8544) );
  XNOR U8751 ( .A(n8550), .B(n8548), .Z(n8653) );
  AND U8752 ( .A(n8654), .B(n8655), .Z(n8548) );
  NANDN U8753 ( .A(n8656), .B(n8657), .Z(n8655) );
  OR U8754 ( .A(n8658), .B(n8659), .Z(n8657) );
  NAND U8755 ( .A(n8659), .B(n8658), .Z(n8654) );
  ANDN U8756 ( .B(B[240]), .A(n32), .Z(n8550) );
  XNOR U8757 ( .A(n8558), .B(n8660), .Z(n8551) );
  XNOR U8758 ( .A(n8557), .B(n8555), .Z(n8660) );
  AND U8759 ( .A(n8661), .B(n8662), .Z(n8555) );
  NANDN U8760 ( .A(n8663), .B(n8664), .Z(n8662) );
  NANDN U8761 ( .A(n8665), .B(n8666), .Z(n8664) );
  NANDN U8762 ( .A(n8666), .B(n8665), .Z(n8661) );
  ANDN U8763 ( .B(B[241]), .A(n33), .Z(n8557) );
  XNOR U8764 ( .A(n8565), .B(n8667), .Z(n8558) );
  XNOR U8765 ( .A(n8564), .B(n8562), .Z(n8667) );
  AND U8766 ( .A(n8668), .B(n8669), .Z(n8562) );
  NANDN U8767 ( .A(n8670), .B(n8671), .Z(n8669) );
  OR U8768 ( .A(n8672), .B(n8673), .Z(n8671) );
  NAND U8769 ( .A(n8673), .B(n8672), .Z(n8668) );
  ANDN U8770 ( .B(B[242]), .A(n34), .Z(n8564) );
  XNOR U8771 ( .A(n8572), .B(n8674), .Z(n8565) );
  XNOR U8772 ( .A(n8571), .B(n8569), .Z(n8674) );
  AND U8773 ( .A(n8675), .B(n8676), .Z(n8569) );
  NANDN U8774 ( .A(n8677), .B(n8678), .Z(n8676) );
  NANDN U8775 ( .A(n8679), .B(n8680), .Z(n8678) );
  NANDN U8776 ( .A(n8680), .B(n8679), .Z(n8675) );
  ANDN U8777 ( .B(B[243]), .A(n35), .Z(n8571) );
  XNOR U8778 ( .A(n8579), .B(n8681), .Z(n8572) );
  XNOR U8779 ( .A(n8578), .B(n8576), .Z(n8681) );
  AND U8780 ( .A(n8682), .B(n8683), .Z(n8576) );
  NANDN U8781 ( .A(n8684), .B(n8685), .Z(n8683) );
  OR U8782 ( .A(n8686), .B(n8687), .Z(n8685) );
  NAND U8783 ( .A(n8687), .B(n8686), .Z(n8682) );
  ANDN U8784 ( .B(B[244]), .A(n36), .Z(n8578) );
  XNOR U8785 ( .A(n8586), .B(n8688), .Z(n8579) );
  XNOR U8786 ( .A(n8585), .B(n8583), .Z(n8688) );
  AND U8787 ( .A(n8689), .B(n8690), .Z(n8583) );
  NANDN U8788 ( .A(n8691), .B(n8692), .Z(n8690) );
  NANDN U8789 ( .A(n8693), .B(n8694), .Z(n8692) );
  NANDN U8790 ( .A(n8694), .B(n8693), .Z(n8689) );
  ANDN U8791 ( .B(B[245]), .A(n37), .Z(n8585) );
  XNOR U8792 ( .A(n8593), .B(n8695), .Z(n8586) );
  XNOR U8793 ( .A(n8592), .B(n8590), .Z(n8695) );
  AND U8794 ( .A(n8696), .B(n8697), .Z(n8590) );
  NANDN U8795 ( .A(n8698), .B(n8699), .Z(n8697) );
  OR U8796 ( .A(n8700), .B(n8701), .Z(n8699) );
  NAND U8797 ( .A(n8701), .B(n8700), .Z(n8696) );
  ANDN U8798 ( .B(B[246]), .A(n38), .Z(n8592) );
  XNOR U8799 ( .A(n8600), .B(n8702), .Z(n8593) );
  XNOR U8800 ( .A(n8599), .B(n8597), .Z(n8702) );
  AND U8801 ( .A(n8703), .B(n8704), .Z(n8597) );
  NANDN U8802 ( .A(n8705), .B(n8706), .Z(n8704) );
  NANDN U8803 ( .A(n8707), .B(n8708), .Z(n8706) );
  NANDN U8804 ( .A(n8708), .B(n8707), .Z(n8703) );
  ANDN U8805 ( .B(B[247]), .A(n39), .Z(n8599) );
  XNOR U8806 ( .A(n8607), .B(n8709), .Z(n8600) );
  XNOR U8807 ( .A(n8606), .B(n8604), .Z(n8709) );
  AND U8808 ( .A(n8710), .B(n8711), .Z(n8604) );
  NANDN U8809 ( .A(n8712), .B(n8713), .Z(n8711) );
  OR U8810 ( .A(n8714), .B(n8715), .Z(n8713) );
  NAND U8811 ( .A(n8715), .B(n8714), .Z(n8710) );
  ANDN U8812 ( .B(B[248]), .A(n40), .Z(n8606) );
  XNOR U8813 ( .A(n8614), .B(n8716), .Z(n8607) );
  XNOR U8814 ( .A(n8613), .B(n8611), .Z(n8716) );
  AND U8815 ( .A(n8717), .B(n8718), .Z(n8611) );
  NANDN U8816 ( .A(n8719), .B(n8720), .Z(n8718) );
  NAND U8817 ( .A(n8721), .B(n8722), .Z(n8720) );
  ANDN U8818 ( .B(B[249]), .A(n41), .Z(n8613) );
  XOR U8819 ( .A(n8620), .B(n8723), .Z(n8614) );
  XNOR U8820 ( .A(n8618), .B(n8621), .Z(n8723) );
  NAND U8821 ( .A(A[2]), .B(B[250]), .Z(n8621) );
  NANDN U8822 ( .A(n8724), .B(n8725), .Z(n8618) );
  AND U8823 ( .A(A[0]), .B(B[251]), .Z(n8725) );
  XNOR U8824 ( .A(n8623), .B(n8726), .Z(n8620) );
  NAND U8825 ( .A(A[0]), .B(B[252]), .Z(n8726) );
  NAND U8826 ( .A(B[251]), .B(A[1]), .Z(n8623) );
  NAND U8827 ( .A(n8727), .B(n8728), .Z(n231) );
  NANDN U8828 ( .A(n8729), .B(n8730), .Z(n8728) );
  OR U8829 ( .A(n8731), .B(n8732), .Z(n8730) );
  NAND U8830 ( .A(n8732), .B(n8731), .Z(n8727) );
  XOR U8831 ( .A(n213), .B(n212), .Z(\A1[24] ) );
  XOR U8832 ( .A(n7815), .B(n8733), .Z(n212) );
  XNOR U8833 ( .A(n7814), .B(n7812), .Z(n8733) );
  AND U8834 ( .A(n8734), .B(n8735), .Z(n7812) );
  NANDN U8835 ( .A(n8736), .B(n8737), .Z(n8735) );
  NANDN U8836 ( .A(n8738), .B(n8739), .Z(n8737) );
  NANDN U8837 ( .A(n8739), .B(n8738), .Z(n8734) );
  ANDN U8838 ( .B(B[11]), .A(n29), .Z(n7814) );
  XNOR U8839 ( .A(n7721), .B(n8740), .Z(n7815) );
  XNOR U8840 ( .A(n7720), .B(n7718), .Z(n8740) );
  AND U8841 ( .A(n8741), .B(n8742), .Z(n7718) );
  NANDN U8842 ( .A(n8743), .B(n8744), .Z(n8742) );
  OR U8843 ( .A(n8745), .B(n8746), .Z(n8744) );
  NAND U8844 ( .A(n8746), .B(n8745), .Z(n8741) );
  ANDN U8845 ( .B(B[12]), .A(n30), .Z(n7720) );
  XNOR U8846 ( .A(n7728), .B(n8747), .Z(n7721) );
  XNOR U8847 ( .A(n7727), .B(n7725), .Z(n8747) );
  AND U8848 ( .A(n8748), .B(n8749), .Z(n7725) );
  NANDN U8849 ( .A(n8750), .B(n8751), .Z(n8749) );
  NANDN U8850 ( .A(n8752), .B(n8753), .Z(n8751) );
  NANDN U8851 ( .A(n8753), .B(n8752), .Z(n8748) );
  ANDN U8852 ( .B(B[13]), .A(n31), .Z(n7727) );
  XNOR U8853 ( .A(n7735), .B(n8754), .Z(n7728) );
  XNOR U8854 ( .A(n7734), .B(n7732), .Z(n8754) );
  AND U8855 ( .A(n8755), .B(n8756), .Z(n7732) );
  NANDN U8856 ( .A(n8757), .B(n8758), .Z(n8756) );
  OR U8857 ( .A(n8759), .B(n8760), .Z(n8758) );
  NAND U8858 ( .A(n8760), .B(n8759), .Z(n8755) );
  ANDN U8859 ( .B(B[14]), .A(n32), .Z(n7734) );
  XNOR U8860 ( .A(n7742), .B(n8761), .Z(n7735) );
  XNOR U8861 ( .A(n7741), .B(n7739), .Z(n8761) );
  AND U8862 ( .A(n8762), .B(n8763), .Z(n7739) );
  NANDN U8863 ( .A(n8764), .B(n8765), .Z(n8763) );
  NANDN U8864 ( .A(n8766), .B(n8767), .Z(n8765) );
  NANDN U8865 ( .A(n8767), .B(n8766), .Z(n8762) );
  ANDN U8866 ( .B(B[15]), .A(n33), .Z(n7741) );
  XNOR U8867 ( .A(n7749), .B(n8768), .Z(n7742) );
  XNOR U8868 ( .A(n7748), .B(n7746), .Z(n8768) );
  AND U8869 ( .A(n8769), .B(n8770), .Z(n7746) );
  NANDN U8870 ( .A(n8771), .B(n8772), .Z(n8770) );
  OR U8871 ( .A(n8773), .B(n8774), .Z(n8772) );
  NAND U8872 ( .A(n8774), .B(n8773), .Z(n8769) );
  ANDN U8873 ( .B(B[16]), .A(n34), .Z(n7748) );
  XNOR U8874 ( .A(n7756), .B(n8775), .Z(n7749) );
  XNOR U8875 ( .A(n7755), .B(n7753), .Z(n8775) );
  AND U8876 ( .A(n8776), .B(n8777), .Z(n7753) );
  NANDN U8877 ( .A(n8778), .B(n8779), .Z(n8777) );
  NANDN U8878 ( .A(n8780), .B(n8781), .Z(n8779) );
  NANDN U8879 ( .A(n8781), .B(n8780), .Z(n8776) );
  ANDN U8880 ( .B(B[17]), .A(n35), .Z(n7755) );
  XNOR U8881 ( .A(n7763), .B(n8782), .Z(n7756) );
  XNOR U8882 ( .A(n7762), .B(n7760), .Z(n8782) );
  AND U8883 ( .A(n8783), .B(n8784), .Z(n7760) );
  NANDN U8884 ( .A(n8785), .B(n8786), .Z(n8784) );
  OR U8885 ( .A(n8787), .B(n8788), .Z(n8786) );
  NAND U8886 ( .A(n8788), .B(n8787), .Z(n8783) );
  ANDN U8887 ( .B(B[18]), .A(n36), .Z(n7762) );
  XNOR U8888 ( .A(n7770), .B(n8789), .Z(n7763) );
  XNOR U8889 ( .A(n7769), .B(n7767), .Z(n8789) );
  AND U8890 ( .A(n8790), .B(n8791), .Z(n7767) );
  NANDN U8891 ( .A(n8792), .B(n8793), .Z(n8791) );
  NANDN U8892 ( .A(n8794), .B(n8795), .Z(n8793) );
  NANDN U8893 ( .A(n8795), .B(n8794), .Z(n8790) );
  ANDN U8894 ( .B(B[19]), .A(n37), .Z(n7769) );
  XNOR U8895 ( .A(n7777), .B(n8796), .Z(n7770) );
  XNOR U8896 ( .A(n7776), .B(n7774), .Z(n8796) );
  AND U8897 ( .A(n8797), .B(n8798), .Z(n7774) );
  NANDN U8898 ( .A(n8799), .B(n8800), .Z(n8798) );
  OR U8899 ( .A(n8801), .B(n8802), .Z(n8800) );
  NAND U8900 ( .A(n8802), .B(n8801), .Z(n8797) );
  ANDN U8901 ( .B(B[20]), .A(n38), .Z(n7776) );
  XNOR U8902 ( .A(n7784), .B(n8803), .Z(n7777) );
  XNOR U8903 ( .A(n7783), .B(n7781), .Z(n8803) );
  AND U8904 ( .A(n8804), .B(n8805), .Z(n7781) );
  NANDN U8905 ( .A(n8806), .B(n8807), .Z(n8805) );
  NANDN U8906 ( .A(n8808), .B(n8809), .Z(n8807) );
  NANDN U8907 ( .A(n8809), .B(n8808), .Z(n8804) );
  ANDN U8908 ( .B(B[21]), .A(n39), .Z(n7783) );
  XNOR U8909 ( .A(n7791), .B(n8810), .Z(n7784) );
  XNOR U8910 ( .A(n7790), .B(n7788), .Z(n8810) );
  AND U8911 ( .A(n8811), .B(n8812), .Z(n7788) );
  NANDN U8912 ( .A(n8813), .B(n8814), .Z(n8812) );
  OR U8913 ( .A(n8815), .B(n8816), .Z(n8814) );
  NAND U8914 ( .A(n8816), .B(n8815), .Z(n8811) );
  ANDN U8915 ( .B(B[22]), .A(n40), .Z(n7790) );
  XNOR U8916 ( .A(n7798), .B(n8817), .Z(n7791) );
  XNOR U8917 ( .A(n7797), .B(n7795), .Z(n8817) );
  AND U8918 ( .A(n8818), .B(n8819), .Z(n7795) );
  NANDN U8919 ( .A(n8820), .B(n8821), .Z(n8819) );
  NAND U8920 ( .A(n8822), .B(n8823), .Z(n8821) );
  ANDN U8921 ( .B(B[23]), .A(n41), .Z(n7797) );
  XOR U8922 ( .A(n7804), .B(n8824), .Z(n7798) );
  XNOR U8923 ( .A(n7802), .B(n7805), .Z(n8824) );
  NAND U8924 ( .A(A[2]), .B(B[24]), .Z(n7805) );
  NANDN U8925 ( .A(n8825), .B(n8826), .Z(n7802) );
  AND U8926 ( .A(A[0]), .B(B[25]), .Z(n8826) );
  XNOR U8927 ( .A(n7807), .B(n8827), .Z(n7804) );
  NAND U8928 ( .A(A[0]), .B(B[26]), .Z(n8827) );
  NAND U8929 ( .A(B[25]), .B(A[1]), .Z(n7807) );
  NAND U8930 ( .A(n8828), .B(n8829), .Z(n213) );
  NANDN U8931 ( .A(n8830), .B(n8831), .Z(n8829) );
  OR U8932 ( .A(n8832), .B(n8833), .Z(n8831) );
  NAND U8933 ( .A(n8833), .B(n8832), .Z(n8828) );
  XOR U8934 ( .A(n233), .B(n232), .Z(\A1[249] ) );
  XOR U8935 ( .A(n8732), .B(n8834), .Z(n232) );
  XNOR U8936 ( .A(n8731), .B(n8729), .Z(n8834) );
  AND U8937 ( .A(n8835), .B(n8836), .Z(n8729) );
  NANDN U8938 ( .A(n8837), .B(n8838), .Z(n8836) );
  NANDN U8939 ( .A(n8839), .B(n8840), .Z(n8838) );
  NANDN U8940 ( .A(n8840), .B(n8839), .Z(n8835) );
  ANDN U8941 ( .B(B[236]), .A(n29), .Z(n8731) );
  XNOR U8942 ( .A(n8638), .B(n8841), .Z(n8732) );
  XNOR U8943 ( .A(n8637), .B(n8635), .Z(n8841) );
  AND U8944 ( .A(n8842), .B(n8843), .Z(n8635) );
  NANDN U8945 ( .A(n8844), .B(n8845), .Z(n8843) );
  OR U8946 ( .A(n8846), .B(n8847), .Z(n8845) );
  NAND U8947 ( .A(n8847), .B(n8846), .Z(n8842) );
  ANDN U8948 ( .B(B[237]), .A(n30), .Z(n8637) );
  XNOR U8949 ( .A(n8645), .B(n8848), .Z(n8638) );
  XNOR U8950 ( .A(n8644), .B(n8642), .Z(n8848) );
  AND U8951 ( .A(n8849), .B(n8850), .Z(n8642) );
  NANDN U8952 ( .A(n8851), .B(n8852), .Z(n8850) );
  NANDN U8953 ( .A(n8853), .B(n8854), .Z(n8852) );
  NANDN U8954 ( .A(n8854), .B(n8853), .Z(n8849) );
  ANDN U8955 ( .B(B[238]), .A(n31), .Z(n8644) );
  XNOR U8956 ( .A(n8652), .B(n8855), .Z(n8645) );
  XNOR U8957 ( .A(n8651), .B(n8649), .Z(n8855) );
  AND U8958 ( .A(n8856), .B(n8857), .Z(n8649) );
  NANDN U8959 ( .A(n8858), .B(n8859), .Z(n8857) );
  OR U8960 ( .A(n8860), .B(n8861), .Z(n8859) );
  NAND U8961 ( .A(n8861), .B(n8860), .Z(n8856) );
  ANDN U8962 ( .B(B[239]), .A(n32), .Z(n8651) );
  XNOR U8963 ( .A(n8659), .B(n8862), .Z(n8652) );
  XNOR U8964 ( .A(n8658), .B(n8656), .Z(n8862) );
  AND U8965 ( .A(n8863), .B(n8864), .Z(n8656) );
  NANDN U8966 ( .A(n8865), .B(n8866), .Z(n8864) );
  NANDN U8967 ( .A(n8867), .B(n8868), .Z(n8866) );
  NANDN U8968 ( .A(n8868), .B(n8867), .Z(n8863) );
  ANDN U8969 ( .B(B[240]), .A(n33), .Z(n8658) );
  XNOR U8970 ( .A(n8666), .B(n8869), .Z(n8659) );
  XNOR U8971 ( .A(n8665), .B(n8663), .Z(n8869) );
  AND U8972 ( .A(n8870), .B(n8871), .Z(n8663) );
  NANDN U8973 ( .A(n8872), .B(n8873), .Z(n8871) );
  OR U8974 ( .A(n8874), .B(n8875), .Z(n8873) );
  NAND U8975 ( .A(n8875), .B(n8874), .Z(n8870) );
  ANDN U8976 ( .B(B[241]), .A(n34), .Z(n8665) );
  XNOR U8977 ( .A(n8673), .B(n8876), .Z(n8666) );
  XNOR U8978 ( .A(n8672), .B(n8670), .Z(n8876) );
  AND U8979 ( .A(n8877), .B(n8878), .Z(n8670) );
  NANDN U8980 ( .A(n8879), .B(n8880), .Z(n8878) );
  NANDN U8981 ( .A(n8881), .B(n8882), .Z(n8880) );
  NANDN U8982 ( .A(n8882), .B(n8881), .Z(n8877) );
  ANDN U8983 ( .B(B[242]), .A(n35), .Z(n8672) );
  XNOR U8984 ( .A(n8680), .B(n8883), .Z(n8673) );
  XNOR U8985 ( .A(n8679), .B(n8677), .Z(n8883) );
  AND U8986 ( .A(n8884), .B(n8885), .Z(n8677) );
  NANDN U8987 ( .A(n8886), .B(n8887), .Z(n8885) );
  OR U8988 ( .A(n8888), .B(n8889), .Z(n8887) );
  NAND U8989 ( .A(n8889), .B(n8888), .Z(n8884) );
  ANDN U8990 ( .B(B[243]), .A(n36), .Z(n8679) );
  XNOR U8991 ( .A(n8687), .B(n8890), .Z(n8680) );
  XNOR U8992 ( .A(n8686), .B(n8684), .Z(n8890) );
  AND U8993 ( .A(n8891), .B(n8892), .Z(n8684) );
  NANDN U8994 ( .A(n8893), .B(n8894), .Z(n8892) );
  NANDN U8995 ( .A(n8895), .B(n8896), .Z(n8894) );
  NANDN U8996 ( .A(n8896), .B(n8895), .Z(n8891) );
  ANDN U8997 ( .B(B[244]), .A(n37), .Z(n8686) );
  XNOR U8998 ( .A(n8694), .B(n8897), .Z(n8687) );
  XNOR U8999 ( .A(n8693), .B(n8691), .Z(n8897) );
  AND U9000 ( .A(n8898), .B(n8899), .Z(n8691) );
  NANDN U9001 ( .A(n8900), .B(n8901), .Z(n8899) );
  OR U9002 ( .A(n8902), .B(n8903), .Z(n8901) );
  NAND U9003 ( .A(n8903), .B(n8902), .Z(n8898) );
  ANDN U9004 ( .B(B[245]), .A(n38), .Z(n8693) );
  XNOR U9005 ( .A(n8701), .B(n8904), .Z(n8694) );
  XNOR U9006 ( .A(n8700), .B(n8698), .Z(n8904) );
  AND U9007 ( .A(n8905), .B(n8906), .Z(n8698) );
  NANDN U9008 ( .A(n8907), .B(n8908), .Z(n8906) );
  NANDN U9009 ( .A(n8909), .B(n8910), .Z(n8908) );
  NANDN U9010 ( .A(n8910), .B(n8909), .Z(n8905) );
  ANDN U9011 ( .B(B[246]), .A(n39), .Z(n8700) );
  XNOR U9012 ( .A(n8708), .B(n8911), .Z(n8701) );
  XNOR U9013 ( .A(n8707), .B(n8705), .Z(n8911) );
  AND U9014 ( .A(n8912), .B(n8913), .Z(n8705) );
  NANDN U9015 ( .A(n8914), .B(n8915), .Z(n8913) );
  OR U9016 ( .A(n8916), .B(n8917), .Z(n8915) );
  NAND U9017 ( .A(n8917), .B(n8916), .Z(n8912) );
  ANDN U9018 ( .B(B[247]), .A(n40), .Z(n8707) );
  XNOR U9019 ( .A(n8715), .B(n8918), .Z(n8708) );
  XNOR U9020 ( .A(n8714), .B(n8712), .Z(n8918) );
  AND U9021 ( .A(n8919), .B(n8920), .Z(n8712) );
  NANDN U9022 ( .A(n8921), .B(n8922), .Z(n8920) );
  NAND U9023 ( .A(n8923), .B(n8924), .Z(n8922) );
  ANDN U9024 ( .B(B[248]), .A(n41), .Z(n8714) );
  XOR U9025 ( .A(n8721), .B(n8925), .Z(n8715) );
  XNOR U9026 ( .A(n8719), .B(n8722), .Z(n8925) );
  NAND U9027 ( .A(A[2]), .B(B[249]), .Z(n8722) );
  NANDN U9028 ( .A(n8926), .B(n8927), .Z(n8719) );
  AND U9029 ( .A(A[0]), .B(B[250]), .Z(n8927) );
  XNOR U9030 ( .A(n8724), .B(n8928), .Z(n8721) );
  NAND U9031 ( .A(A[0]), .B(B[251]), .Z(n8928) );
  NAND U9032 ( .A(B[250]), .B(A[1]), .Z(n8724) );
  NAND U9033 ( .A(n8929), .B(n8930), .Z(n233) );
  NANDN U9034 ( .A(n8931), .B(n8932), .Z(n8930) );
  OR U9035 ( .A(n8933), .B(n8934), .Z(n8932) );
  NAND U9036 ( .A(n8934), .B(n8933), .Z(n8929) );
  XOR U9037 ( .A(n237), .B(n236), .Z(\A1[248] ) );
  XOR U9038 ( .A(n8934), .B(n8935), .Z(n236) );
  XNOR U9039 ( .A(n8933), .B(n8931), .Z(n8935) );
  AND U9040 ( .A(n8936), .B(n8937), .Z(n8931) );
  NANDN U9041 ( .A(n8938), .B(n8939), .Z(n8937) );
  NANDN U9042 ( .A(n8940), .B(n8941), .Z(n8939) );
  NANDN U9043 ( .A(n8941), .B(n8940), .Z(n8936) );
  ANDN U9044 ( .B(B[235]), .A(n29), .Z(n8933) );
  XNOR U9045 ( .A(n8840), .B(n8942), .Z(n8934) );
  XNOR U9046 ( .A(n8839), .B(n8837), .Z(n8942) );
  AND U9047 ( .A(n8943), .B(n8944), .Z(n8837) );
  NANDN U9048 ( .A(n8945), .B(n8946), .Z(n8944) );
  OR U9049 ( .A(n8947), .B(n8948), .Z(n8946) );
  NAND U9050 ( .A(n8948), .B(n8947), .Z(n8943) );
  ANDN U9051 ( .B(B[236]), .A(n30), .Z(n8839) );
  XNOR U9052 ( .A(n8847), .B(n8949), .Z(n8840) );
  XNOR U9053 ( .A(n8846), .B(n8844), .Z(n8949) );
  AND U9054 ( .A(n8950), .B(n8951), .Z(n8844) );
  NANDN U9055 ( .A(n8952), .B(n8953), .Z(n8951) );
  NANDN U9056 ( .A(n8954), .B(n8955), .Z(n8953) );
  NANDN U9057 ( .A(n8955), .B(n8954), .Z(n8950) );
  ANDN U9058 ( .B(B[237]), .A(n31), .Z(n8846) );
  XNOR U9059 ( .A(n8854), .B(n8956), .Z(n8847) );
  XNOR U9060 ( .A(n8853), .B(n8851), .Z(n8956) );
  AND U9061 ( .A(n8957), .B(n8958), .Z(n8851) );
  NANDN U9062 ( .A(n8959), .B(n8960), .Z(n8958) );
  OR U9063 ( .A(n8961), .B(n8962), .Z(n8960) );
  NAND U9064 ( .A(n8962), .B(n8961), .Z(n8957) );
  ANDN U9065 ( .B(B[238]), .A(n32), .Z(n8853) );
  XNOR U9066 ( .A(n8861), .B(n8963), .Z(n8854) );
  XNOR U9067 ( .A(n8860), .B(n8858), .Z(n8963) );
  AND U9068 ( .A(n8964), .B(n8965), .Z(n8858) );
  NANDN U9069 ( .A(n8966), .B(n8967), .Z(n8965) );
  NANDN U9070 ( .A(n8968), .B(n8969), .Z(n8967) );
  NANDN U9071 ( .A(n8969), .B(n8968), .Z(n8964) );
  ANDN U9072 ( .B(B[239]), .A(n33), .Z(n8860) );
  XNOR U9073 ( .A(n8868), .B(n8970), .Z(n8861) );
  XNOR U9074 ( .A(n8867), .B(n8865), .Z(n8970) );
  AND U9075 ( .A(n8971), .B(n8972), .Z(n8865) );
  NANDN U9076 ( .A(n8973), .B(n8974), .Z(n8972) );
  OR U9077 ( .A(n8975), .B(n8976), .Z(n8974) );
  NAND U9078 ( .A(n8976), .B(n8975), .Z(n8971) );
  ANDN U9079 ( .B(B[240]), .A(n34), .Z(n8867) );
  XNOR U9080 ( .A(n8875), .B(n8977), .Z(n8868) );
  XNOR U9081 ( .A(n8874), .B(n8872), .Z(n8977) );
  AND U9082 ( .A(n8978), .B(n8979), .Z(n8872) );
  NANDN U9083 ( .A(n8980), .B(n8981), .Z(n8979) );
  NANDN U9084 ( .A(n8982), .B(n8983), .Z(n8981) );
  NANDN U9085 ( .A(n8983), .B(n8982), .Z(n8978) );
  ANDN U9086 ( .B(B[241]), .A(n35), .Z(n8874) );
  XNOR U9087 ( .A(n8882), .B(n8984), .Z(n8875) );
  XNOR U9088 ( .A(n8881), .B(n8879), .Z(n8984) );
  AND U9089 ( .A(n8985), .B(n8986), .Z(n8879) );
  NANDN U9090 ( .A(n8987), .B(n8988), .Z(n8986) );
  OR U9091 ( .A(n8989), .B(n8990), .Z(n8988) );
  NAND U9092 ( .A(n8990), .B(n8989), .Z(n8985) );
  ANDN U9093 ( .B(B[242]), .A(n36), .Z(n8881) );
  XNOR U9094 ( .A(n8889), .B(n8991), .Z(n8882) );
  XNOR U9095 ( .A(n8888), .B(n8886), .Z(n8991) );
  AND U9096 ( .A(n8992), .B(n8993), .Z(n8886) );
  NANDN U9097 ( .A(n8994), .B(n8995), .Z(n8993) );
  NANDN U9098 ( .A(n8996), .B(n8997), .Z(n8995) );
  NANDN U9099 ( .A(n8997), .B(n8996), .Z(n8992) );
  ANDN U9100 ( .B(B[243]), .A(n37), .Z(n8888) );
  XNOR U9101 ( .A(n8896), .B(n8998), .Z(n8889) );
  XNOR U9102 ( .A(n8895), .B(n8893), .Z(n8998) );
  AND U9103 ( .A(n8999), .B(n9000), .Z(n8893) );
  NANDN U9104 ( .A(n9001), .B(n9002), .Z(n9000) );
  OR U9105 ( .A(n9003), .B(n9004), .Z(n9002) );
  NAND U9106 ( .A(n9004), .B(n9003), .Z(n8999) );
  ANDN U9107 ( .B(B[244]), .A(n38), .Z(n8895) );
  XNOR U9108 ( .A(n8903), .B(n9005), .Z(n8896) );
  XNOR U9109 ( .A(n8902), .B(n8900), .Z(n9005) );
  AND U9110 ( .A(n9006), .B(n9007), .Z(n8900) );
  NANDN U9111 ( .A(n9008), .B(n9009), .Z(n9007) );
  NANDN U9112 ( .A(n9010), .B(n9011), .Z(n9009) );
  NANDN U9113 ( .A(n9011), .B(n9010), .Z(n9006) );
  ANDN U9114 ( .B(B[245]), .A(n39), .Z(n8902) );
  XNOR U9115 ( .A(n8910), .B(n9012), .Z(n8903) );
  XNOR U9116 ( .A(n8909), .B(n8907), .Z(n9012) );
  AND U9117 ( .A(n9013), .B(n9014), .Z(n8907) );
  NANDN U9118 ( .A(n9015), .B(n9016), .Z(n9014) );
  OR U9119 ( .A(n9017), .B(n9018), .Z(n9016) );
  NAND U9120 ( .A(n9018), .B(n9017), .Z(n9013) );
  ANDN U9121 ( .B(B[246]), .A(n40), .Z(n8909) );
  XNOR U9122 ( .A(n8917), .B(n9019), .Z(n8910) );
  XNOR U9123 ( .A(n8916), .B(n8914), .Z(n9019) );
  AND U9124 ( .A(n9020), .B(n9021), .Z(n8914) );
  NANDN U9125 ( .A(n9022), .B(n9023), .Z(n9021) );
  NAND U9126 ( .A(n9024), .B(n9025), .Z(n9023) );
  ANDN U9127 ( .B(B[247]), .A(n41), .Z(n8916) );
  XOR U9128 ( .A(n8923), .B(n9026), .Z(n8917) );
  XNOR U9129 ( .A(n8921), .B(n8924), .Z(n9026) );
  NAND U9130 ( .A(A[2]), .B(B[248]), .Z(n8924) );
  NANDN U9131 ( .A(n9027), .B(n9028), .Z(n8921) );
  AND U9132 ( .A(A[0]), .B(B[249]), .Z(n9028) );
  XNOR U9133 ( .A(n8926), .B(n9029), .Z(n8923) );
  NAND U9134 ( .A(A[0]), .B(B[250]), .Z(n9029) );
  NAND U9135 ( .A(B[249]), .B(A[1]), .Z(n8926) );
  NAND U9136 ( .A(n9030), .B(n9031), .Z(n237) );
  NANDN U9137 ( .A(n9032), .B(n9033), .Z(n9031) );
  OR U9138 ( .A(n9034), .B(n9035), .Z(n9033) );
  NAND U9139 ( .A(n9035), .B(n9034), .Z(n9030) );
  XOR U9140 ( .A(n239), .B(n238), .Z(\A1[247] ) );
  XOR U9141 ( .A(n9035), .B(n9036), .Z(n238) );
  XNOR U9142 ( .A(n9034), .B(n9032), .Z(n9036) );
  AND U9143 ( .A(n9037), .B(n9038), .Z(n9032) );
  NANDN U9144 ( .A(n9039), .B(n9040), .Z(n9038) );
  NANDN U9145 ( .A(n9041), .B(n9042), .Z(n9040) );
  NANDN U9146 ( .A(n9042), .B(n9041), .Z(n9037) );
  ANDN U9147 ( .B(B[234]), .A(n29), .Z(n9034) );
  XNOR U9148 ( .A(n8941), .B(n9043), .Z(n9035) );
  XNOR U9149 ( .A(n8940), .B(n8938), .Z(n9043) );
  AND U9150 ( .A(n9044), .B(n9045), .Z(n8938) );
  NANDN U9151 ( .A(n9046), .B(n9047), .Z(n9045) );
  OR U9152 ( .A(n9048), .B(n9049), .Z(n9047) );
  NAND U9153 ( .A(n9049), .B(n9048), .Z(n9044) );
  ANDN U9154 ( .B(B[235]), .A(n30), .Z(n8940) );
  XNOR U9155 ( .A(n8948), .B(n9050), .Z(n8941) );
  XNOR U9156 ( .A(n8947), .B(n8945), .Z(n9050) );
  AND U9157 ( .A(n9051), .B(n9052), .Z(n8945) );
  NANDN U9158 ( .A(n9053), .B(n9054), .Z(n9052) );
  NANDN U9159 ( .A(n9055), .B(n9056), .Z(n9054) );
  NANDN U9160 ( .A(n9056), .B(n9055), .Z(n9051) );
  ANDN U9161 ( .B(B[236]), .A(n31), .Z(n8947) );
  XNOR U9162 ( .A(n8955), .B(n9057), .Z(n8948) );
  XNOR U9163 ( .A(n8954), .B(n8952), .Z(n9057) );
  AND U9164 ( .A(n9058), .B(n9059), .Z(n8952) );
  NANDN U9165 ( .A(n9060), .B(n9061), .Z(n9059) );
  OR U9166 ( .A(n9062), .B(n9063), .Z(n9061) );
  NAND U9167 ( .A(n9063), .B(n9062), .Z(n9058) );
  ANDN U9168 ( .B(B[237]), .A(n32), .Z(n8954) );
  XNOR U9169 ( .A(n8962), .B(n9064), .Z(n8955) );
  XNOR U9170 ( .A(n8961), .B(n8959), .Z(n9064) );
  AND U9171 ( .A(n9065), .B(n9066), .Z(n8959) );
  NANDN U9172 ( .A(n9067), .B(n9068), .Z(n9066) );
  NANDN U9173 ( .A(n9069), .B(n9070), .Z(n9068) );
  NANDN U9174 ( .A(n9070), .B(n9069), .Z(n9065) );
  ANDN U9175 ( .B(B[238]), .A(n33), .Z(n8961) );
  XNOR U9176 ( .A(n8969), .B(n9071), .Z(n8962) );
  XNOR U9177 ( .A(n8968), .B(n8966), .Z(n9071) );
  AND U9178 ( .A(n9072), .B(n9073), .Z(n8966) );
  NANDN U9179 ( .A(n9074), .B(n9075), .Z(n9073) );
  OR U9180 ( .A(n9076), .B(n9077), .Z(n9075) );
  NAND U9181 ( .A(n9077), .B(n9076), .Z(n9072) );
  ANDN U9182 ( .B(B[239]), .A(n34), .Z(n8968) );
  XNOR U9183 ( .A(n8976), .B(n9078), .Z(n8969) );
  XNOR U9184 ( .A(n8975), .B(n8973), .Z(n9078) );
  AND U9185 ( .A(n9079), .B(n9080), .Z(n8973) );
  NANDN U9186 ( .A(n9081), .B(n9082), .Z(n9080) );
  NANDN U9187 ( .A(n9083), .B(n9084), .Z(n9082) );
  NANDN U9188 ( .A(n9084), .B(n9083), .Z(n9079) );
  ANDN U9189 ( .B(B[240]), .A(n35), .Z(n8975) );
  XNOR U9190 ( .A(n8983), .B(n9085), .Z(n8976) );
  XNOR U9191 ( .A(n8982), .B(n8980), .Z(n9085) );
  AND U9192 ( .A(n9086), .B(n9087), .Z(n8980) );
  NANDN U9193 ( .A(n9088), .B(n9089), .Z(n9087) );
  OR U9194 ( .A(n9090), .B(n9091), .Z(n9089) );
  NAND U9195 ( .A(n9091), .B(n9090), .Z(n9086) );
  ANDN U9196 ( .B(B[241]), .A(n36), .Z(n8982) );
  XNOR U9197 ( .A(n8990), .B(n9092), .Z(n8983) );
  XNOR U9198 ( .A(n8989), .B(n8987), .Z(n9092) );
  AND U9199 ( .A(n9093), .B(n9094), .Z(n8987) );
  NANDN U9200 ( .A(n9095), .B(n9096), .Z(n9094) );
  NANDN U9201 ( .A(n9097), .B(n9098), .Z(n9096) );
  NANDN U9202 ( .A(n9098), .B(n9097), .Z(n9093) );
  ANDN U9203 ( .B(B[242]), .A(n37), .Z(n8989) );
  XNOR U9204 ( .A(n8997), .B(n9099), .Z(n8990) );
  XNOR U9205 ( .A(n8996), .B(n8994), .Z(n9099) );
  AND U9206 ( .A(n9100), .B(n9101), .Z(n8994) );
  NANDN U9207 ( .A(n9102), .B(n9103), .Z(n9101) );
  OR U9208 ( .A(n9104), .B(n9105), .Z(n9103) );
  NAND U9209 ( .A(n9105), .B(n9104), .Z(n9100) );
  ANDN U9210 ( .B(B[243]), .A(n38), .Z(n8996) );
  XNOR U9211 ( .A(n9004), .B(n9106), .Z(n8997) );
  XNOR U9212 ( .A(n9003), .B(n9001), .Z(n9106) );
  AND U9213 ( .A(n9107), .B(n9108), .Z(n9001) );
  NANDN U9214 ( .A(n9109), .B(n9110), .Z(n9108) );
  NANDN U9215 ( .A(n9111), .B(n9112), .Z(n9110) );
  NANDN U9216 ( .A(n9112), .B(n9111), .Z(n9107) );
  ANDN U9217 ( .B(B[244]), .A(n39), .Z(n9003) );
  XNOR U9218 ( .A(n9011), .B(n9113), .Z(n9004) );
  XNOR U9219 ( .A(n9010), .B(n9008), .Z(n9113) );
  AND U9220 ( .A(n9114), .B(n9115), .Z(n9008) );
  NANDN U9221 ( .A(n9116), .B(n9117), .Z(n9115) );
  OR U9222 ( .A(n9118), .B(n9119), .Z(n9117) );
  NAND U9223 ( .A(n9119), .B(n9118), .Z(n9114) );
  ANDN U9224 ( .B(B[245]), .A(n40), .Z(n9010) );
  XNOR U9225 ( .A(n9018), .B(n9120), .Z(n9011) );
  XNOR U9226 ( .A(n9017), .B(n9015), .Z(n9120) );
  AND U9227 ( .A(n9121), .B(n9122), .Z(n9015) );
  NANDN U9228 ( .A(n9123), .B(n9124), .Z(n9122) );
  NAND U9229 ( .A(n9125), .B(n9126), .Z(n9124) );
  ANDN U9230 ( .B(B[246]), .A(n41), .Z(n9017) );
  XOR U9231 ( .A(n9024), .B(n9127), .Z(n9018) );
  XNOR U9232 ( .A(n9022), .B(n9025), .Z(n9127) );
  NAND U9233 ( .A(A[2]), .B(B[247]), .Z(n9025) );
  NANDN U9234 ( .A(n9128), .B(n9129), .Z(n9022) );
  AND U9235 ( .A(A[0]), .B(B[248]), .Z(n9129) );
  XNOR U9236 ( .A(n9027), .B(n9130), .Z(n9024) );
  NAND U9237 ( .A(A[0]), .B(B[249]), .Z(n9130) );
  NAND U9238 ( .A(B[248]), .B(A[1]), .Z(n9027) );
  NAND U9239 ( .A(n9131), .B(n9132), .Z(n239) );
  NANDN U9240 ( .A(n9133), .B(n9134), .Z(n9132) );
  OR U9241 ( .A(n9135), .B(n9136), .Z(n9134) );
  NAND U9242 ( .A(n9136), .B(n9135), .Z(n9131) );
  XOR U9243 ( .A(n241), .B(n240), .Z(\A1[246] ) );
  XOR U9244 ( .A(n9136), .B(n9137), .Z(n240) );
  XNOR U9245 ( .A(n9135), .B(n9133), .Z(n9137) );
  AND U9246 ( .A(n9138), .B(n9139), .Z(n9133) );
  NANDN U9247 ( .A(n9140), .B(n9141), .Z(n9139) );
  NANDN U9248 ( .A(n9142), .B(n9143), .Z(n9141) );
  NANDN U9249 ( .A(n9143), .B(n9142), .Z(n9138) );
  ANDN U9250 ( .B(B[233]), .A(n29), .Z(n9135) );
  XNOR U9251 ( .A(n9042), .B(n9144), .Z(n9136) );
  XNOR U9252 ( .A(n9041), .B(n9039), .Z(n9144) );
  AND U9253 ( .A(n9145), .B(n9146), .Z(n9039) );
  NANDN U9254 ( .A(n9147), .B(n9148), .Z(n9146) );
  OR U9255 ( .A(n9149), .B(n9150), .Z(n9148) );
  NAND U9256 ( .A(n9150), .B(n9149), .Z(n9145) );
  ANDN U9257 ( .B(B[234]), .A(n30), .Z(n9041) );
  XNOR U9258 ( .A(n9049), .B(n9151), .Z(n9042) );
  XNOR U9259 ( .A(n9048), .B(n9046), .Z(n9151) );
  AND U9260 ( .A(n9152), .B(n9153), .Z(n9046) );
  NANDN U9261 ( .A(n9154), .B(n9155), .Z(n9153) );
  NANDN U9262 ( .A(n9156), .B(n9157), .Z(n9155) );
  NANDN U9263 ( .A(n9157), .B(n9156), .Z(n9152) );
  ANDN U9264 ( .B(B[235]), .A(n31), .Z(n9048) );
  XNOR U9265 ( .A(n9056), .B(n9158), .Z(n9049) );
  XNOR U9266 ( .A(n9055), .B(n9053), .Z(n9158) );
  AND U9267 ( .A(n9159), .B(n9160), .Z(n9053) );
  NANDN U9268 ( .A(n9161), .B(n9162), .Z(n9160) );
  OR U9269 ( .A(n9163), .B(n9164), .Z(n9162) );
  NAND U9270 ( .A(n9164), .B(n9163), .Z(n9159) );
  ANDN U9271 ( .B(B[236]), .A(n32), .Z(n9055) );
  XNOR U9272 ( .A(n9063), .B(n9165), .Z(n9056) );
  XNOR U9273 ( .A(n9062), .B(n9060), .Z(n9165) );
  AND U9274 ( .A(n9166), .B(n9167), .Z(n9060) );
  NANDN U9275 ( .A(n9168), .B(n9169), .Z(n9167) );
  NANDN U9276 ( .A(n9170), .B(n9171), .Z(n9169) );
  NANDN U9277 ( .A(n9171), .B(n9170), .Z(n9166) );
  ANDN U9278 ( .B(B[237]), .A(n33), .Z(n9062) );
  XNOR U9279 ( .A(n9070), .B(n9172), .Z(n9063) );
  XNOR U9280 ( .A(n9069), .B(n9067), .Z(n9172) );
  AND U9281 ( .A(n9173), .B(n9174), .Z(n9067) );
  NANDN U9282 ( .A(n9175), .B(n9176), .Z(n9174) );
  OR U9283 ( .A(n9177), .B(n9178), .Z(n9176) );
  NAND U9284 ( .A(n9178), .B(n9177), .Z(n9173) );
  ANDN U9285 ( .B(B[238]), .A(n34), .Z(n9069) );
  XNOR U9286 ( .A(n9077), .B(n9179), .Z(n9070) );
  XNOR U9287 ( .A(n9076), .B(n9074), .Z(n9179) );
  AND U9288 ( .A(n9180), .B(n9181), .Z(n9074) );
  NANDN U9289 ( .A(n9182), .B(n9183), .Z(n9181) );
  NANDN U9290 ( .A(n9184), .B(n9185), .Z(n9183) );
  NANDN U9291 ( .A(n9185), .B(n9184), .Z(n9180) );
  ANDN U9292 ( .B(B[239]), .A(n35), .Z(n9076) );
  XNOR U9293 ( .A(n9084), .B(n9186), .Z(n9077) );
  XNOR U9294 ( .A(n9083), .B(n9081), .Z(n9186) );
  AND U9295 ( .A(n9187), .B(n9188), .Z(n9081) );
  NANDN U9296 ( .A(n9189), .B(n9190), .Z(n9188) );
  OR U9297 ( .A(n9191), .B(n9192), .Z(n9190) );
  NAND U9298 ( .A(n9192), .B(n9191), .Z(n9187) );
  ANDN U9299 ( .B(B[240]), .A(n36), .Z(n9083) );
  XNOR U9300 ( .A(n9091), .B(n9193), .Z(n9084) );
  XNOR U9301 ( .A(n9090), .B(n9088), .Z(n9193) );
  AND U9302 ( .A(n9194), .B(n9195), .Z(n9088) );
  NANDN U9303 ( .A(n9196), .B(n9197), .Z(n9195) );
  NANDN U9304 ( .A(n9198), .B(n9199), .Z(n9197) );
  NANDN U9305 ( .A(n9199), .B(n9198), .Z(n9194) );
  ANDN U9306 ( .B(B[241]), .A(n37), .Z(n9090) );
  XNOR U9307 ( .A(n9098), .B(n9200), .Z(n9091) );
  XNOR U9308 ( .A(n9097), .B(n9095), .Z(n9200) );
  AND U9309 ( .A(n9201), .B(n9202), .Z(n9095) );
  NANDN U9310 ( .A(n9203), .B(n9204), .Z(n9202) );
  OR U9311 ( .A(n9205), .B(n9206), .Z(n9204) );
  NAND U9312 ( .A(n9206), .B(n9205), .Z(n9201) );
  ANDN U9313 ( .B(B[242]), .A(n38), .Z(n9097) );
  XNOR U9314 ( .A(n9105), .B(n9207), .Z(n9098) );
  XNOR U9315 ( .A(n9104), .B(n9102), .Z(n9207) );
  AND U9316 ( .A(n9208), .B(n9209), .Z(n9102) );
  NANDN U9317 ( .A(n9210), .B(n9211), .Z(n9209) );
  NANDN U9318 ( .A(n9212), .B(n9213), .Z(n9211) );
  NANDN U9319 ( .A(n9213), .B(n9212), .Z(n9208) );
  ANDN U9320 ( .B(B[243]), .A(n39), .Z(n9104) );
  XNOR U9321 ( .A(n9112), .B(n9214), .Z(n9105) );
  XNOR U9322 ( .A(n9111), .B(n9109), .Z(n9214) );
  AND U9323 ( .A(n9215), .B(n9216), .Z(n9109) );
  NANDN U9324 ( .A(n9217), .B(n9218), .Z(n9216) );
  OR U9325 ( .A(n9219), .B(n9220), .Z(n9218) );
  NAND U9326 ( .A(n9220), .B(n9219), .Z(n9215) );
  ANDN U9327 ( .B(B[244]), .A(n40), .Z(n9111) );
  XNOR U9328 ( .A(n9119), .B(n9221), .Z(n9112) );
  XNOR U9329 ( .A(n9118), .B(n9116), .Z(n9221) );
  AND U9330 ( .A(n9222), .B(n9223), .Z(n9116) );
  NANDN U9331 ( .A(n9224), .B(n9225), .Z(n9223) );
  NAND U9332 ( .A(n9226), .B(n9227), .Z(n9225) );
  ANDN U9333 ( .B(B[245]), .A(n41), .Z(n9118) );
  XOR U9334 ( .A(n9125), .B(n9228), .Z(n9119) );
  XNOR U9335 ( .A(n9123), .B(n9126), .Z(n9228) );
  NAND U9336 ( .A(A[2]), .B(B[246]), .Z(n9126) );
  NANDN U9337 ( .A(n9229), .B(n9230), .Z(n9123) );
  AND U9338 ( .A(A[0]), .B(B[247]), .Z(n9230) );
  XNOR U9339 ( .A(n9128), .B(n9231), .Z(n9125) );
  NAND U9340 ( .A(A[0]), .B(B[248]), .Z(n9231) );
  NAND U9341 ( .A(B[247]), .B(A[1]), .Z(n9128) );
  NAND U9342 ( .A(n9232), .B(n9233), .Z(n241) );
  NANDN U9343 ( .A(n9234), .B(n9235), .Z(n9233) );
  OR U9344 ( .A(n9236), .B(n9237), .Z(n9235) );
  NAND U9345 ( .A(n9237), .B(n9236), .Z(n9232) );
  XOR U9346 ( .A(n243), .B(n242), .Z(\A1[245] ) );
  XOR U9347 ( .A(n9237), .B(n9238), .Z(n242) );
  XNOR U9348 ( .A(n9236), .B(n9234), .Z(n9238) );
  AND U9349 ( .A(n9239), .B(n9240), .Z(n9234) );
  NANDN U9350 ( .A(n9241), .B(n9242), .Z(n9240) );
  NANDN U9351 ( .A(n9243), .B(n9244), .Z(n9242) );
  NANDN U9352 ( .A(n9244), .B(n9243), .Z(n9239) );
  ANDN U9353 ( .B(B[232]), .A(n29), .Z(n9236) );
  XNOR U9354 ( .A(n9143), .B(n9245), .Z(n9237) );
  XNOR U9355 ( .A(n9142), .B(n9140), .Z(n9245) );
  AND U9356 ( .A(n9246), .B(n9247), .Z(n9140) );
  NANDN U9357 ( .A(n9248), .B(n9249), .Z(n9247) );
  OR U9358 ( .A(n9250), .B(n9251), .Z(n9249) );
  NAND U9359 ( .A(n9251), .B(n9250), .Z(n9246) );
  ANDN U9360 ( .B(B[233]), .A(n30), .Z(n9142) );
  XNOR U9361 ( .A(n9150), .B(n9252), .Z(n9143) );
  XNOR U9362 ( .A(n9149), .B(n9147), .Z(n9252) );
  AND U9363 ( .A(n9253), .B(n9254), .Z(n9147) );
  NANDN U9364 ( .A(n9255), .B(n9256), .Z(n9254) );
  NANDN U9365 ( .A(n9257), .B(n9258), .Z(n9256) );
  NANDN U9366 ( .A(n9258), .B(n9257), .Z(n9253) );
  ANDN U9367 ( .B(B[234]), .A(n31), .Z(n9149) );
  XNOR U9368 ( .A(n9157), .B(n9259), .Z(n9150) );
  XNOR U9369 ( .A(n9156), .B(n9154), .Z(n9259) );
  AND U9370 ( .A(n9260), .B(n9261), .Z(n9154) );
  NANDN U9371 ( .A(n9262), .B(n9263), .Z(n9261) );
  OR U9372 ( .A(n9264), .B(n9265), .Z(n9263) );
  NAND U9373 ( .A(n9265), .B(n9264), .Z(n9260) );
  ANDN U9374 ( .B(B[235]), .A(n32), .Z(n9156) );
  XNOR U9375 ( .A(n9164), .B(n9266), .Z(n9157) );
  XNOR U9376 ( .A(n9163), .B(n9161), .Z(n9266) );
  AND U9377 ( .A(n9267), .B(n9268), .Z(n9161) );
  NANDN U9378 ( .A(n9269), .B(n9270), .Z(n9268) );
  NANDN U9379 ( .A(n9271), .B(n9272), .Z(n9270) );
  NANDN U9380 ( .A(n9272), .B(n9271), .Z(n9267) );
  ANDN U9381 ( .B(B[236]), .A(n33), .Z(n9163) );
  XNOR U9382 ( .A(n9171), .B(n9273), .Z(n9164) );
  XNOR U9383 ( .A(n9170), .B(n9168), .Z(n9273) );
  AND U9384 ( .A(n9274), .B(n9275), .Z(n9168) );
  NANDN U9385 ( .A(n9276), .B(n9277), .Z(n9275) );
  OR U9386 ( .A(n9278), .B(n9279), .Z(n9277) );
  NAND U9387 ( .A(n9279), .B(n9278), .Z(n9274) );
  ANDN U9388 ( .B(B[237]), .A(n34), .Z(n9170) );
  XNOR U9389 ( .A(n9178), .B(n9280), .Z(n9171) );
  XNOR U9390 ( .A(n9177), .B(n9175), .Z(n9280) );
  AND U9391 ( .A(n9281), .B(n9282), .Z(n9175) );
  NANDN U9392 ( .A(n9283), .B(n9284), .Z(n9282) );
  NANDN U9393 ( .A(n9285), .B(n9286), .Z(n9284) );
  NANDN U9394 ( .A(n9286), .B(n9285), .Z(n9281) );
  ANDN U9395 ( .B(B[238]), .A(n35), .Z(n9177) );
  XNOR U9396 ( .A(n9185), .B(n9287), .Z(n9178) );
  XNOR U9397 ( .A(n9184), .B(n9182), .Z(n9287) );
  AND U9398 ( .A(n9288), .B(n9289), .Z(n9182) );
  NANDN U9399 ( .A(n9290), .B(n9291), .Z(n9289) );
  OR U9400 ( .A(n9292), .B(n9293), .Z(n9291) );
  NAND U9401 ( .A(n9293), .B(n9292), .Z(n9288) );
  ANDN U9402 ( .B(B[239]), .A(n36), .Z(n9184) );
  XNOR U9403 ( .A(n9192), .B(n9294), .Z(n9185) );
  XNOR U9404 ( .A(n9191), .B(n9189), .Z(n9294) );
  AND U9405 ( .A(n9295), .B(n9296), .Z(n9189) );
  NANDN U9406 ( .A(n9297), .B(n9298), .Z(n9296) );
  NANDN U9407 ( .A(n9299), .B(n9300), .Z(n9298) );
  NANDN U9408 ( .A(n9300), .B(n9299), .Z(n9295) );
  ANDN U9409 ( .B(B[240]), .A(n37), .Z(n9191) );
  XNOR U9410 ( .A(n9199), .B(n9301), .Z(n9192) );
  XNOR U9411 ( .A(n9198), .B(n9196), .Z(n9301) );
  AND U9412 ( .A(n9302), .B(n9303), .Z(n9196) );
  NANDN U9413 ( .A(n9304), .B(n9305), .Z(n9303) );
  OR U9414 ( .A(n9306), .B(n9307), .Z(n9305) );
  NAND U9415 ( .A(n9307), .B(n9306), .Z(n9302) );
  ANDN U9416 ( .B(B[241]), .A(n38), .Z(n9198) );
  XNOR U9417 ( .A(n9206), .B(n9308), .Z(n9199) );
  XNOR U9418 ( .A(n9205), .B(n9203), .Z(n9308) );
  AND U9419 ( .A(n9309), .B(n9310), .Z(n9203) );
  NANDN U9420 ( .A(n9311), .B(n9312), .Z(n9310) );
  NANDN U9421 ( .A(n9313), .B(n9314), .Z(n9312) );
  NANDN U9422 ( .A(n9314), .B(n9313), .Z(n9309) );
  ANDN U9423 ( .B(B[242]), .A(n39), .Z(n9205) );
  XNOR U9424 ( .A(n9213), .B(n9315), .Z(n9206) );
  XNOR U9425 ( .A(n9212), .B(n9210), .Z(n9315) );
  AND U9426 ( .A(n9316), .B(n9317), .Z(n9210) );
  NANDN U9427 ( .A(n9318), .B(n9319), .Z(n9317) );
  OR U9428 ( .A(n9320), .B(n9321), .Z(n9319) );
  NAND U9429 ( .A(n9321), .B(n9320), .Z(n9316) );
  ANDN U9430 ( .B(B[243]), .A(n40), .Z(n9212) );
  XNOR U9431 ( .A(n9220), .B(n9322), .Z(n9213) );
  XNOR U9432 ( .A(n9219), .B(n9217), .Z(n9322) );
  AND U9433 ( .A(n9323), .B(n9324), .Z(n9217) );
  NANDN U9434 ( .A(n9325), .B(n9326), .Z(n9324) );
  NAND U9435 ( .A(n9327), .B(n9328), .Z(n9326) );
  ANDN U9436 ( .B(B[244]), .A(n41), .Z(n9219) );
  XOR U9437 ( .A(n9226), .B(n9329), .Z(n9220) );
  XNOR U9438 ( .A(n9224), .B(n9227), .Z(n9329) );
  NAND U9439 ( .A(A[2]), .B(B[245]), .Z(n9227) );
  NANDN U9440 ( .A(n9330), .B(n9331), .Z(n9224) );
  AND U9441 ( .A(A[0]), .B(B[246]), .Z(n9331) );
  XNOR U9442 ( .A(n9229), .B(n9332), .Z(n9226) );
  NAND U9443 ( .A(A[0]), .B(B[247]), .Z(n9332) );
  NAND U9444 ( .A(B[246]), .B(A[1]), .Z(n9229) );
  NAND U9445 ( .A(n9333), .B(n9334), .Z(n243) );
  NANDN U9446 ( .A(n9335), .B(n9336), .Z(n9334) );
  OR U9447 ( .A(n9337), .B(n9338), .Z(n9336) );
  NAND U9448 ( .A(n9338), .B(n9337), .Z(n9333) );
  XOR U9449 ( .A(n245), .B(n244), .Z(\A1[244] ) );
  XOR U9450 ( .A(n9338), .B(n9339), .Z(n244) );
  XNOR U9451 ( .A(n9337), .B(n9335), .Z(n9339) );
  AND U9452 ( .A(n9340), .B(n9341), .Z(n9335) );
  NANDN U9453 ( .A(n9342), .B(n9343), .Z(n9341) );
  NANDN U9454 ( .A(n9344), .B(n9345), .Z(n9343) );
  NANDN U9455 ( .A(n9345), .B(n9344), .Z(n9340) );
  ANDN U9456 ( .B(B[231]), .A(n29), .Z(n9337) );
  XNOR U9457 ( .A(n9244), .B(n9346), .Z(n9338) );
  XNOR U9458 ( .A(n9243), .B(n9241), .Z(n9346) );
  AND U9459 ( .A(n9347), .B(n9348), .Z(n9241) );
  NANDN U9460 ( .A(n9349), .B(n9350), .Z(n9348) );
  OR U9461 ( .A(n9351), .B(n9352), .Z(n9350) );
  NAND U9462 ( .A(n9352), .B(n9351), .Z(n9347) );
  ANDN U9463 ( .B(B[232]), .A(n30), .Z(n9243) );
  XNOR U9464 ( .A(n9251), .B(n9353), .Z(n9244) );
  XNOR U9465 ( .A(n9250), .B(n9248), .Z(n9353) );
  AND U9466 ( .A(n9354), .B(n9355), .Z(n9248) );
  NANDN U9467 ( .A(n9356), .B(n9357), .Z(n9355) );
  NANDN U9468 ( .A(n9358), .B(n9359), .Z(n9357) );
  NANDN U9469 ( .A(n9359), .B(n9358), .Z(n9354) );
  ANDN U9470 ( .B(B[233]), .A(n31), .Z(n9250) );
  XNOR U9471 ( .A(n9258), .B(n9360), .Z(n9251) );
  XNOR U9472 ( .A(n9257), .B(n9255), .Z(n9360) );
  AND U9473 ( .A(n9361), .B(n9362), .Z(n9255) );
  NANDN U9474 ( .A(n9363), .B(n9364), .Z(n9362) );
  OR U9475 ( .A(n9365), .B(n9366), .Z(n9364) );
  NAND U9476 ( .A(n9366), .B(n9365), .Z(n9361) );
  ANDN U9477 ( .B(B[234]), .A(n32), .Z(n9257) );
  XNOR U9478 ( .A(n9265), .B(n9367), .Z(n9258) );
  XNOR U9479 ( .A(n9264), .B(n9262), .Z(n9367) );
  AND U9480 ( .A(n9368), .B(n9369), .Z(n9262) );
  NANDN U9481 ( .A(n9370), .B(n9371), .Z(n9369) );
  NANDN U9482 ( .A(n9372), .B(n9373), .Z(n9371) );
  NANDN U9483 ( .A(n9373), .B(n9372), .Z(n9368) );
  ANDN U9484 ( .B(B[235]), .A(n33), .Z(n9264) );
  XNOR U9485 ( .A(n9272), .B(n9374), .Z(n9265) );
  XNOR U9486 ( .A(n9271), .B(n9269), .Z(n9374) );
  AND U9487 ( .A(n9375), .B(n9376), .Z(n9269) );
  NANDN U9488 ( .A(n9377), .B(n9378), .Z(n9376) );
  OR U9489 ( .A(n9379), .B(n9380), .Z(n9378) );
  NAND U9490 ( .A(n9380), .B(n9379), .Z(n9375) );
  ANDN U9491 ( .B(B[236]), .A(n34), .Z(n9271) );
  XNOR U9492 ( .A(n9279), .B(n9381), .Z(n9272) );
  XNOR U9493 ( .A(n9278), .B(n9276), .Z(n9381) );
  AND U9494 ( .A(n9382), .B(n9383), .Z(n9276) );
  NANDN U9495 ( .A(n9384), .B(n9385), .Z(n9383) );
  NANDN U9496 ( .A(n9386), .B(n9387), .Z(n9385) );
  NANDN U9497 ( .A(n9387), .B(n9386), .Z(n9382) );
  ANDN U9498 ( .B(B[237]), .A(n35), .Z(n9278) );
  XNOR U9499 ( .A(n9286), .B(n9388), .Z(n9279) );
  XNOR U9500 ( .A(n9285), .B(n9283), .Z(n9388) );
  AND U9501 ( .A(n9389), .B(n9390), .Z(n9283) );
  NANDN U9502 ( .A(n9391), .B(n9392), .Z(n9390) );
  OR U9503 ( .A(n9393), .B(n9394), .Z(n9392) );
  NAND U9504 ( .A(n9394), .B(n9393), .Z(n9389) );
  ANDN U9505 ( .B(B[238]), .A(n36), .Z(n9285) );
  XNOR U9506 ( .A(n9293), .B(n9395), .Z(n9286) );
  XNOR U9507 ( .A(n9292), .B(n9290), .Z(n9395) );
  AND U9508 ( .A(n9396), .B(n9397), .Z(n9290) );
  NANDN U9509 ( .A(n9398), .B(n9399), .Z(n9397) );
  NANDN U9510 ( .A(n9400), .B(n9401), .Z(n9399) );
  NANDN U9511 ( .A(n9401), .B(n9400), .Z(n9396) );
  ANDN U9512 ( .B(B[239]), .A(n37), .Z(n9292) );
  XNOR U9513 ( .A(n9300), .B(n9402), .Z(n9293) );
  XNOR U9514 ( .A(n9299), .B(n9297), .Z(n9402) );
  AND U9515 ( .A(n9403), .B(n9404), .Z(n9297) );
  NANDN U9516 ( .A(n9405), .B(n9406), .Z(n9404) );
  OR U9517 ( .A(n9407), .B(n9408), .Z(n9406) );
  NAND U9518 ( .A(n9408), .B(n9407), .Z(n9403) );
  ANDN U9519 ( .B(B[240]), .A(n38), .Z(n9299) );
  XNOR U9520 ( .A(n9307), .B(n9409), .Z(n9300) );
  XNOR U9521 ( .A(n9306), .B(n9304), .Z(n9409) );
  AND U9522 ( .A(n9410), .B(n9411), .Z(n9304) );
  NANDN U9523 ( .A(n9412), .B(n9413), .Z(n9411) );
  NANDN U9524 ( .A(n9414), .B(n9415), .Z(n9413) );
  NANDN U9525 ( .A(n9415), .B(n9414), .Z(n9410) );
  ANDN U9526 ( .B(B[241]), .A(n39), .Z(n9306) );
  XNOR U9527 ( .A(n9314), .B(n9416), .Z(n9307) );
  XNOR U9528 ( .A(n9313), .B(n9311), .Z(n9416) );
  AND U9529 ( .A(n9417), .B(n9418), .Z(n9311) );
  NANDN U9530 ( .A(n9419), .B(n9420), .Z(n9418) );
  OR U9531 ( .A(n9421), .B(n9422), .Z(n9420) );
  NAND U9532 ( .A(n9422), .B(n9421), .Z(n9417) );
  ANDN U9533 ( .B(B[242]), .A(n40), .Z(n9313) );
  XNOR U9534 ( .A(n9321), .B(n9423), .Z(n9314) );
  XNOR U9535 ( .A(n9320), .B(n9318), .Z(n9423) );
  AND U9536 ( .A(n9424), .B(n9425), .Z(n9318) );
  NANDN U9537 ( .A(n9426), .B(n9427), .Z(n9425) );
  NAND U9538 ( .A(n9428), .B(n9429), .Z(n9427) );
  ANDN U9539 ( .B(B[243]), .A(n41), .Z(n9320) );
  XOR U9540 ( .A(n9327), .B(n9430), .Z(n9321) );
  XNOR U9541 ( .A(n9325), .B(n9328), .Z(n9430) );
  NAND U9542 ( .A(A[2]), .B(B[244]), .Z(n9328) );
  NANDN U9543 ( .A(n9431), .B(n9432), .Z(n9325) );
  AND U9544 ( .A(A[0]), .B(B[245]), .Z(n9432) );
  XNOR U9545 ( .A(n9330), .B(n9433), .Z(n9327) );
  NAND U9546 ( .A(A[0]), .B(B[246]), .Z(n9433) );
  NAND U9547 ( .A(B[245]), .B(A[1]), .Z(n9330) );
  NAND U9548 ( .A(n9434), .B(n9435), .Z(n245) );
  NANDN U9549 ( .A(n9436), .B(n9437), .Z(n9435) );
  OR U9550 ( .A(n9438), .B(n9439), .Z(n9437) );
  NAND U9551 ( .A(n9439), .B(n9438), .Z(n9434) );
  XOR U9552 ( .A(n247), .B(n246), .Z(\A1[243] ) );
  XOR U9553 ( .A(n9439), .B(n9440), .Z(n246) );
  XNOR U9554 ( .A(n9438), .B(n9436), .Z(n9440) );
  AND U9555 ( .A(n9441), .B(n9442), .Z(n9436) );
  NANDN U9556 ( .A(n9443), .B(n9444), .Z(n9442) );
  NANDN U9557 ( .A(n9445), .B(n9446), .Z(n9444) );
  NANDN U9558 ( .A(n9446), .B(n9445), .Z(n9441) );
  ANDN U9559 ( .B(B[230]), .A(n29), .Z(n9438) );
  XNOR U9560 ( .A(n9345), .B(n9447), .Z(n9439) );
  XNOR U9561 ( .A(n9344), .B(n9342), .Z(n9447) );
  AND U9562 ( .A(n9448), .B(n9449), .Z(n9342) );
  NANDN U9563 ( .A(n9450), .B(n9451), .Z(n9449) );
  OR U9564 ( .A(n9452), .B(n9453), .Z(n9451) );
  NAND U9565 ( .A(n9453), .B(n9452), .Z(n9448) );
  ANDN U9566 ( .B(B[231]), .A(n30), .Z(n9344) );
  XNOR U9567 ( .A(n9352), .B(n9454), .Z(n9345) );
  XNOR U9568 ( .A(n9351), .B(n9349), .Z(n9454) );
  AND U9569 ( .A(n9455), .B(n9456), .Z(n9349) );
  NANDN U9570 ( .A(n9457), .B(n9458), .Z(n9456) );
  NANDN U9571 ( .A(n9459), .B(n9460), .Z(n9458) );
  NANDN U9572 ( .A(n9460), .B(n9459), .Z(n9455) );
  ANDN U9573 ( .B(B[232]), .A(n31), .Z(n9351) );
  XNOR U9574 ( .A(n9359), .B(n9461), .Z(n9352) );
  XNOR U9575 ( .A(n9358), .B(n9356), .Z(n9461) );
  AND U9576 ( .A(n9462), .B(n9463), .Z(n9356) );
  NANDN U9577 ( .A(n9464), .B(n9465), .Z(n9463) );
  OR U9578 ( .A(n9466), .B(n9467), .Z(n9465) );
  NAND U9579 ( .A(n9467), .B(n9466), .Z(n9462) );
  ANDN U9580 ( .B(B[233]), .A(n32), .Z(n9358) );
  XNOR U9581 ( .A(n9366), .B(n9468), .Z(n9359) );
  XNOR U9582 ( .A(n9365), .B(n9363), .Z(n9468) );
  AND U9583 ( .A(n9469), .B(n9470), .Z(n9363) );
  NANDN U9584 ( .A(n9471), .B(n9472), .Z(n9470) );
  NANDN U9585 ( .A(n9473), .B(n9474), .Z(n9472) );
  NANDN U9586 ( .A(n9474), .B(n9473), .Z(n9469) );
  ANDN U9587 ( .B(B[234]), .A(n33), .Z(n9365) );
  XNOR U9588 ( .A(n9373), .B(n9475), .Z(n9366) );
  XNOR U9589 ( .A(n9372), .B(n9370), .Z(n9475) );
  AND U9590 ( .A(n9476), .B(n9477), .Z(n9370) );
  NANDN U9591 ( .A(n9478), .B(n9479), .Z(n9477) );
  OR U9592 ( .A(n9480), .B(n9481), .Z(n9479) );
  NAND U9593 ( .A(n9481), .B(n9480), .Z(n9476) );
  ANDN U9594 ( .B(B[235]), .A(n34), .Z(n9372) );
  XNOR U9595 ( .A(n9380), .B(n9482), .Z(n9373) );
  XNOR U9596 ( .A(n9379), .B(n9377), .Z(n9482) );
  AND U9597 ( .A(n9483), .B(n9484), .Z(n9377) );
  NANDN U9598 ( .A(n9485), .B(n9486), .Z(n9484) );
  NANDN U9599 ( .A(n9487), .B(n9488), .Z(n9486) );
  NANDN U9600 ( .A(n9488), .B(n9487), .Z(n9483) );
  ANDN U9601 ( .B(B[236]), .A(n35), .Z(n9379) );
  XNOR U9602 ( .A(n9387), .B(n9489), .Z(n9380) );
  XNOR U9603 ( .A(n9386), .B(n9384), .Z(n9489) );
  AND U9604 ( .A(n9490), .B(n9491), .Z(n9384) );
  NANDN U9605 ( .A(n9492), .B(n9493), .Z(n9491) );
  OR U9606 ( .A(n9494), .B(n9495), .Z(n9493) );
  NAND U9607 ( .A(n9495), .B(n9494), .Z(n9490) );
  ANDN U9608 ( .B(B[237]), .A(n36), .Z(n9386) );
  XNOR U9609 ( .A(n9394), .B(n9496), .Z(n9387) );
  XNOR U9610 ( .A(n9393), .B(n9391), .Z(n9496) );
  AND U9611 ( .A(n9497), .B(n9498), .Z(n9391) );
  NANDN U9612 ( .A(n9499), .B(n9500), .Z(n9498) );
  NANDN U9613 ( .A(n9501), .B(n9502), .Z(n9500) );
  NANDN U9614 ( .A(n9502), .B(n9501), .Z(n9497) );
  ANDN U9615 ( .B(B[238]), .A(n37), .Z(n9393) );
  XNOR U9616 ( .A(n9401), .B(n9503), .Z(n9394) );
  XNOR U9617 ( .A(n9400), .B(n9398), .Z(n9503) );
  AND U9618 ( .A(n9504), .B(n9505), .Z(n9398) );
  NANDN U9619 ( .A(n9506), .B(n9507), .Z(n9505) );
  OR U9620 ( .A(n9508), .B(n9509), .Z(n9507) );
  NAND U9621 ( .A(n9509), .B(n9508), .Z(n9504) );
  ANDN U9622 ( .B(B[239]), .A(n38), .Z(n9400) );
  XNOR U9623 ( .A(n9408), .B(n9510), .Z(n9401) );
  XNOR U9624 ( .A(n9407), .B(n9405), .Z(n9510) );
  AND U9625 ( .A(n9511), .B(n9512), .Z(n9405) );
  NANDN U9626 ( .A(n9513), .B(n9514), .Z(n9512) );
  NANDN U9627 ( .A(n9515), .B(n9516), .Z(n9514) );
  NANDN U9628 ( .A(n9516), .B(n9515), .Z(n9511) );
  ANDN U9629 ( .B(B[240]), .A(n39), .Z(n9407) );
  XNOR U9630 ( .A(n9415), .B(n9517), .Z(n9408) );
  XNOR U9631 ( .A(n9414), .B(n9412), .Z(n9517) );
  AND U9632 ( .A(n9518), .B(n9519), .Z(n9412) );
  NANDN U9633 ( .A(n9520), .B(n9521), .Z(n9519) );
  OR U9634 ( .A(n9522), .B(n9523), .Z(n9521) );
  NAND U9635 ( .A(n9523), .B(n9522), .Z(n9518) );
  ANDN U9636 ( .B(B[241]), .A(n40), .Z(n9414) );
  XNOR U9637 ( .A(n9422), .B(n9524), .Z(n9415) );
  XNOR U9638 ( .A(n9421), .B(n9419), .Z(n9524) );
  AND U9639 ( .A(n9525), .B(n9526), .Z(n9419) );
  NANDN U9640 ( .A(n9527), .B(n9528), .Z(n9526) );
  NAND U9641 ( .A(n9529), .B(n9530), .Z(n9528) );
  ANDN U9642 ( .B(B[242]), .A(n41), .Z(n9421) );
  XOR U9643 ( .A(n9428), .B(n9531), .Z(n9422) );
  XNOR U9644 ( .A(n9426), .B(n9429), .Z(n9531) );
  NAND U9645 ( .A(A[2]), .B(B[243]), .Z(n9429) );
  NANDN U9646 ( .A(n9532), .B(n9533), .Z(n9426) );
  AND U9647 ( .A(A[0]), .B(B[244]), .Z(n9533) );
  XNOR U9648 ( .A(n9431), .B(n9534), .Z(n9428) );
  NAND U9649 ( .A(A[0]), .B(B[245]), .Z(n9534) );
  NAND U9650 ( .A(B[244]), .B(A[1]), .Z(n9431) );
  NAND U9651 ( .A(n9535), .B(n9536), .Z(n247) );
  NANDN U9652 ( .A(n9537), .B(n9538), .Z(n9536) );
  OR U9653 ( .A(n9539), .B(n9540), .Z(n9538) );
  NAND U9654 ( .A(n9540), .B(n9539), .Z(n9535) );
  XOR U9655 ( .A(n249), .B(n248), .Z(\A1[242] ) );
  XOR U9656 ( .A(n9540), .B(n9541), .Z(n248) );
  XNOR U9657 ( .A(n9539), .B(n9537), .Z(n9541) );
  AND U9658 ( .A(n9542), .B(n9543), .Z(n9537) );
  NANDN U9659 ( .A(n9544), .B(n9545), .Z(n9543) );
  NANDN U9660 ( .A(n9546), .B(n9547), .Z(n9545) );
  NANDN U9661 ( .A(n9547), .B(n9546), .Z(n9542) );
  ANDN U9662 ( .B(B[229]), .A(n29), .Z(n9539) );
  XNOR U9663 ( .A(n9446), .B(n9548), .Z(n9540) );
  XNOR U9664 ( .A(n9445), .B(n9443), .Z(n9548) );
  AND U9665 ( .A(n9549), .B(n9550), .Z(n9443) );
  NANDN U9666 ( .A(n9551), .B(n9552), .Z(n9550) );
  OR U9667 ( .A(n9553), .B(n9554), .Z(n9552) );
  NAND U9668 ( .A(n9554), .B(n9553), .Z(n9549) );
  ANDN U9669 ( .B(B[230]), .A(n30), .Z(n9445) );
  XNOR U9670 ( .A(n9453), .B(n9555), .Z(n9446) );
  XNOR U9671 ( .A(n9452), .B(n9450), .Z(n9555) );
  AND U9672 ( .A(n9556), .B(n9557), .Z(n9450) );
  NANDN U9673 ( .A(n9558), .B(n9559), .Z(n9557) );
  NANDN U9674 ( .A(n9560), .B(n9561), .Z(n9559) );
  NANDN U9675 ( .A(n9561), .B(n9560), .Z(n9556) );
  ANDN U9676 ( .B(B[231]), .A(n31), .Z(n9452) );
  XNOR U9677 ( .A(n9460), .B(n9562), .Z(n9453) );
  XNOR U9678 ( .A(n9459), .B(n9457), .Z(n9562) );
  AND U9679 ( .A(n9563), .B(n9564), .Z(n9457) );
  NANDN U9680 ( .A(n9565), .B(n9566), .Z(n9564) );
  OR U9681 ( .A(n9567), .B(n9568), .Z(n9566) );
  NAND U9682 ( .A(n9568), .B(n9567), .Z(n9563) );
  ANDN U9683 ( .B(B[232]), .A(n32), .Z(n9459) );
  XNOR U9684 ( .A(n9467), .B(n9569), .Z(n9460) );
  XNOR U9685 ( .A(n9466), .B(n9464), .Z(n9569) );
  AND U9686 ( .A(n9570), .B(n9571), .Z(n9464) );
  NANDN U9687 ( .A(n9572), .B(n9573), .Z(n9571) );
  NANDN U9688 ( .A(n9574), .B(n9575), .Z(n9573) );
  NANDN U9689 ( .A(n9575), .B(n9574), .Z(n9570) );
  ANDN U9690 ( .B(B[233]), .A(n33), .Z(n9466) );
  XNOR U9691 ( .A(n9474), .B(n9576), .Z(n9467) );
  XNOR U9692 ( .A(n9473), .B(n9471), .Z(n9576) );
  AND U9693 ( .A(n9577), .B(n9578), .Z(n9471) );
  NANDN U9694 ( .A(n9579), .B(n9580), .Z(n9578) );
  OR U9695 ( .A(n9581), .B(n9582), .Z(n9580) );
  NAND U9696 ( .A(n9582), .B(n9581), .Z(n9577) );
  ANDN U9697 ( .B(B[234]), .A(n34), .Z(n9473) );
  XNOR U9698 ( .A(n9481), .B(n9583), .Z(n9474) );
  XNOR U9699 ( .A(n9480), .B(n9478), .Z(n9583) );
  AND U9700 ( .A(n9584), .B(n9585), .Z(n9478) );
  NANDN U9701 ( .A(n9586), .B(n9587), .Z(n9585) );
  NANDN U9702 ( .A(n9588), .B(n9589), .Z(n9587) );
  NANDN U9703 ( .A(n9589), .B(n9588), .Z(n9584) );
  ANDN U9704 ( .B(B[235]), .A(n35), .Z(n9480) );
  XNOR U9705 ( .A(n9488), .B(n9590), .Z(n9481) );
  XNOR U9706 ( .A(n9487), .B(n9485), .Z(n9590) );
  AND U9707 ( .A(n9591), .B(n9592), .Z(n9485) );
  NANDN U9708 ( .A(n9593), .B(n9594), .Z(n9592) );
  OR U9709 ( .A(n9595), .B(n9596), .Z(n9594) );
  NAND U9710 ( .A(n9596), .B(n9595), .Z(n9591) );
  ANDN U9711 ( .B(B[236]), .A(n36), .Z(n9487) );
  XNOR U9712 ( .A(n9495), .B(n9597), .Z(n9488) );
  XNOR U9713 ( .A(n9494), .B(n9492), .Z(n9597) );
  AND U9714 ( .A(n9598), .B(n9599), .Z(n9492) );
  NANDN U9715 ( .A(n9600), .B(n9601), .Z(n9599) );
  NANDN U9716 ( .A(n9602), .B(n9603), .Z(n9601) );
  NANDN U9717 ( .A(n9603), .B(n9602), .Z(n9598) );
  ANDN U9718 ( .B(B[237]), .A(n37), .Z(n9494) );
  XNOR U9719 ( .A(n9502), .B(n9604), .Z(n9495) );
  XNOR U9720 ( .A(n9501), .B(n9499), .Z(n9604) );
  AND U9721 ( .A(n9605), .B(n9606), .Z(n9499) );
  NANDN U9722 ( .A(n9607), .B(n9608), .Z(n9606) );
  OR U9723 ( .A(n9609), .B(n9610), .Z(n9608) );
  NAND U9724 ( .A(n9610), .B(n9609), .Z(n9605) );
  ANDN U9725 ( .B(B[238]), .A(n38), .Z(n9501) );
  XNOR U9726 ( .A(n9509), .B(n9611), .Z(n9502) );
  XNOR U9727 ( .A(n9508), .B(n9506), .Z(n9611) );
  AND U9728 ( .A(n9612), .B(n9613), .Z(n9506) );
  NANDN U9729 ( .A(n9614), .B(n9615), .Z(n9613) );
  NANDN U9730 ( .A(n9616), .B(n9617), .Z(n9615) );
  NANDN U9731 ( .A(n9617), .B(n9616), .Z(n9612) );
  ANDN U9732 ( .B(B[239]), .A(n39), .Z(n9508) );
  XNOR U9733 ( .A(n9516), .B(n9618), .Z(n9509) );
  XNOR U9734 ( .A(n9515), .B(n9513), .Z(n9618) );
  AND U9735 ( .A(n9619), .B(n9620), .Z(n9513) );
  NANDN U9736 ( .A(n9621), .B(n9622), .Z(n9620) );
  OR U9737 ( .A(n9623), .B(n9624), .Z(n9622) );
  NAND U9738 ( .A(n9624), .B(n9623), .Z(n9619) );
  ANDN U9739 ( .B(B[240]), .A(n40), .Z(n9515) );
  XNOR U9740 ( .A(n9523), .B(n9625), .Z(n9516) );
  XNOR U9741 ( .A(n9522), .B(n9520), .Z(n9625) );
  AND U9742 ( .A(n9626), .B(n9627), .Z(n9520) );
  NANDN U9743 ( .A(n9628), .B(n9629), .Z(n9627) );
  NAND U9744 ( .A(n9630), .B(n9631), .Z(n9629) );
  ANDN U9745 ( .B(B[241]), .A(n41), .Z(n9522) );
  XOR U9746 ( .A(n9529), .B(n9632), .Z(n9523) );
  XNOR U9747 ( .A(n9527), .B(n9530), .Z(n9632) );
  NAND U9748 ( .A(A[2]), .B(B[242]), .Z(n9530) );
  NANDN U9749 ( .A(n9633), .B(n9634), .Z(n9527) );
  AND U9750 ( .A(A[0]), .B(B[243]), .Z(n9634) );
  XNOR U9751 ( .A(n9532), .B(n9635), .Z(n9529) );
  NAND U9752 ( .A(A[0]), .B(B[244]), .Z(n9635) );
  NAND U9753 ( .A(B[243]), .B(A[1]), .Z(n9532) );
  NAND U9754 ( .A(n9636), .B(n9637), .Z(n249) );
  NANDN U9755 ( .A(n9638), .B(n9639), .Z(n9637) );
  OR U9756 ( .A(n9640), .B(n9641), .Z(n9639) );
  NAND U9757 ( .A(n9641), .B(n9640), .Z(n9636) );
  XOR U9758 ( .A(n251), .B(n250), .Z(\A1[241] ) );
  XOR U9759 ( .A(n9641), .B(n9642), .Z(n250) );
  XNOR U9760 ( .A(n9640), .B(n9638), .Z(n9642) );
  AND U9761 ( .A(n9643), .B(n9644), .Z(n9638) );
  NANDN U9762 ( .A(n9645), .B(n9646), .Z(n9644) );
  NANDN U9763 ( .A(n9647), .B(n9648), .Z(n9646) );
  NANDN U9764 ( .A(n9648), .B(n9647), .Z(n9643) );
  ANDN U9765 ( .B(B[228]), .A(n29), .Z(n9640) );
  XNOR U9766 ( .A(n9547), .B(n9649), .Z(n9641) );
  XNOR U9767 ( .A(n9546), .B(n9544), .Z(n9649) );
  AND U9768 ( .A(n9650), .B(n9651), .Z(n9544) );
  NANDN U9769 ( .A(n9652), .B(n9653), .Z(n9651) );
  OR U9770 ( .A(n9654), .B(n9655), .Z(n9653) );
  NAND U9771 ( .A(n9655), .B(n9654), .Z(n9650) );
  ANDN U9772 ( .B(B[229]), .A(n30), .Z(n9546) );
  XNOR U9773 ( .A(n9554), .B(n9656), .Z(n9547) );
  XNOR U9774 ( .A(n9553), .B(n9551), .Z(n9656) );
  AND U9775 ( .A(n9657), .B(n9658), .Z(n9551) );
  NANDN U9776 ( .A(n9659), .B(n9660), .Z(n9658) );
  NANDN U9777 ( .A(n9661), .B(n9662), .Z(n9660) );
  NANDN U9778 ( .A(n9662), .B(n9661), .Z(n9657) );
  ANDN U9779 ( .B(B[230]), .A(n31), .Z(n9553) );
  XNOR U9780 ( .A(n9561), .B(n9663), .Z(n9554) );
  XNOR U9781 ( .A(n9560), .B(n9558), .Z(n9663) );
  AND U9782 ( .A(n9664), .B(n9665), .Z(n9558) );
  NANDN U9783 ( .A(n9666), .B(n9667), .Z(n9665) );
  OR U9784 ( .A(n9668), .B(n9669), .Z(n9667) );
  NAND U9785 ( .A(n9669), .B(n9668), .Z(n9664) );
  ANDN U9786 ( .B(B[231]), .A(n32), .Z(n9560) );
  XNOR U9787 ( .A(n9568), .B(n9670), .Z(n9561) );
  XNOR U9788 ( .A(n9567), .B(n9565), .Z(n9670) );
  AND U9789 ( .A(n9671), .B(n9672), .Z(n9565) );
  NANDN U9790 ( .A(n9673), .B(n9674), .Z(n9672) );
  NANDN U9791 ( .A(n9675), .B(n9676), .Z(n9674) );
  NANDN U9792 ( .A(n9676), .B(n9675), .Z(n9671) );
  ANDN U9793 ( .B(B[232]), .A(n33), .Z(n9567) );
  XNOR U9794 ( .A(n9575), .B(n9677), .Z(n9568) );
  XNOR U9795 ( .A(n9574), .B(n9572), .Z(n9677) );
  AND U9796 ( .A(n9678), .B(n9679), .Z(n9572) );
  NANDN U9797 ( .A(n9680), .B(n9681), .Z(n9679) );
  OR U9798 ( .A(n9682), .B(n9683), .Z(n9681) );
  NAND U9799 ( .A(n9683), .B(n9682), .Z(n9678) );
  ANDN U9800 ( .B(B[233]), .A(n34), .Z(n9574) );
  XNOR U9801 ( .A(n9582), .B(n9684), .Z(n9575) );
  XNOR U9802 ( .A(n9581), .B(n9579), .Z(n9684) );
  AND U9803 ( .A(n9685), .B(n9686), .Z(n9579) );
  NANDN U9804 ( .A(n9687), .B(n9688), .Z(n9686) );
  NANDN U9805 ( .A(n9689), .B(n9690), .Z(n9688) );
  NANDN U9806 ( .A(n9690), .B(n9689), .Z(n9685) );
  ANDN U9807 ( .B(B[234]), .A(n35), .Z(n9581) );
  XNOR U9808 ( .A(n9589), .B(n9691), .Z(n9582) );
  XNOR U9809 ( .A(n9588), .B(n9586), .Z(n9691) );
  AND U9810 ( .A(n9692), .B(n9693), .Z(n9586) );
  NANDN U9811 ( .A(n9694), .B(n9695), .Z(n9693) );
  OR U9812 ( .A(n9696), .B(n9697), .Z(n9695) );
  NAND U9813 ( .A(n9697), .B(n9696), .Z(n9692) );
  ANDN U9814 ( .B(B[235]), .A(n36), .Z(n9588) );
  XNOR U9815 ( .A(n9596), .B(n9698), .Z(n9589) );
  XNOR U9816 ( .A(n9595), .B(n9593), .Z(n9698) );
  AND U9817 ( .A(n9699), .B(n9700), .Z(n9593) );
  NANDN U9818 ( .A(n9701), .B(n9702), .Z(n9700) );
  NANDN U9819 ( .A(n9703), .B(n9704), .Z(n9702) );
  NANDN U9820 ( .A(n9704), .B(n9703), .Z(n9699) );
  ANDN U9821 ( .B(B[236]), .A(n37), .Z(n9595) );
  XNOR U9822 ( .A(n9603), .B(n9705), .Z(n9596) );
  XNOR U9823 ( .A(n9602), .B(n9600), .Z(n9705) );
  AND U9824 ( .A(n9706), .B(n9707), .Z(n9600) );
  NANDN U9825 ( .A(n9708), .B(n9709), .Z(n9707) );
  OR U9826 ( .A(n9710), .B(n9711), .Z(n9709) );
  NAND U9827 ( .A(n9711), .B(n9710), .Z(n9706) );
  ANDN U9828 ( .B(B[237]), .A(n38), .Z(n9602) );
  XNOR U9829 ( .A(n9610), .B(n9712), .Z(n9603) );
  XNOR U9830 ( .A(n9609), .B(n9607), .Z(n9712) );
  AND U9831 ( .A(n9713), .B(n9714), .Z(n9607) );
  NANDN U9832 ( .A(n9715), .B(n9716), .Z(n9714) );
  NANDN U9833 ( .A(n9717), .B(n9718), .Z(n9716) );
  NANDN U9834 ( .A(n9718), .B(n9717), .Z(n9713) );
  ANDN U9835 ( .B(B[238]), .A(n39), .Z(n9609) );
  XNOR U9836 ( .A(n9617), .B(n9719), .Z(n9610) );
  XNOR U9837 ( .A(n9616), .B(n9614), .Z(n9719) );
  AND U9838 ( .A(n9720), .B(n9721), .Z(n9614) );
  NANDN U9839 ( .A(n9722), .B(n9723), .Z(n9721) );
  OR U9840 ( .A(n9724), .B(n9725), .Z(n9723) );
  NAND U9841 ( .A(n9725), .B(n9724), .Z(n9720) );
  ANDN U9842 ( .B(B[239]), .A(n40), .Z(n9616) );
  XNOR U9843 ( .A(n9624), .B(n9726), .Z(n9617) );
  XNOR U9844 ( .A(n9623), .B(n9621), .Z(n9726) );
  AND U9845 ( .A(n9727), .B(n9728), .Z(n9621) );
  NANDN U9846 ( .A(n9729), .B(n9730), .Z(n9728) );
  NAND U9847 ( .A(n9731), .B(n9732), .Z(n9730) );
  ANDN U9848 ( .B(B[240]), .A(n41), .Z(n9623) );
  XOR U9849 ( .A(n9630), .B(n9733), .Z(n9624) );
  XNOR U9850 ( .A(n9628), .B(n9631), .Z(n9733) );
  NAND U9851 ( .A(A[2]), .B(B[241]), .Z(n9631) );
  NANDN U9852 ( .A(n9734), .B(n9735), .Z(n9628) );
  AND U9853 ( .A(A[0]), .B(B[242]), .Z(n9735) );
  XNOR U9854 ( .A(n9633), .B(n9736), .Z(n9630) );
  NAND U9855 ( .A(A[0]), .B(B[243]), .Z(n9736) );
  NAND U9856 ( .A(B[242]), .B(A[1]), .Z(n9633) );
  NAND U9857 ( .A(n9737), .B(n9738), .Z(n251) );
  NANDN U9858 ( .A(n9739), .B(n9740), .Z(n9738) );
  OR U9859 ( .A(n9741), .B(n9742), .Z(n9740) );
  NAND U9860 ( .A(n9742), .B(n9741), .Z(n9737) );
  XOR U9861 ( .A(n253), .B(n252), .Z(\A1[240] ) );
  XOR U9862 ( .A(n9742), .B(n9743), .Z(n252) );
  XNOR U9863 ( .A(n9741), .B(n9739), .Z(n9743) );
  AND U9864 ( .A(n9744), .B(n9745), .Z(n9739) );
  NANDN U9865 ( .A(n9746), .B(n9747), .Z(n9745) );
  NANDN U9866 ( .A(n9748), .B(n9749), .Z(n9747) );
  NANDN U9867 ( .A(n9749), .B(n9748), .Z(n9744) );
  ANDN U9868 ( .B(B[227]), .A(n29), .Z(n9741) );
  XNOR U9869 ( .A(n9648), .B(n9750), .Z(n9742) );
  XNOR U9870 ( .A(n9647), .B(n9645), .Z(n9750) );
  AND U9871 ( .A(n9751), .B(n9752), .Z(n9645) );
  NANDN U9872 ( .A(n9753), .B(n9754), .Z(n9752) );
  OR U9873 ( .A(n9755), .B(n9756), .Z(n9754) );
  NAND U9874 ( .A(n9756), .B(n9755), .Z(n9751) );
  ANDN U9875 ( .B(B[228]), .A(n30), .Z(n9647) );
  XNOR U9876 ( .A(n9655), .B(n9757), .Z(n9648) );
  XNOR U9877 ( .A(n9654), .B(n9652), .Z(n9757) );
  AND U9878 ( .A(n9758), .B(n9759), .Z(n9652) );
  NANDN U9879 ( .A(n9760), .B(n9761), .Z(n9759) );
  NANDN U9880 ( .A(n9762), .B(n9763), .Z(n9761) );
  NANDN U9881 ( .A(n9763), .B(n9762), .Z(n9758) );
  ANDN U9882 ( .B(B[229]), .A(n31), .Z(n9654) );
  XNOR U9883 ( .A(n9662), .B(n9764), .Z(n9655) );
  XNOR U9884 ( .A(n9661), .B(n9659), .Z(n9764) );
  AND U9885 ( .A(n9765), .B(n9766), .Z(n9659) );
  NANDN U9886 ( .A(n9767), .B(n9768), .Z(n9766) );
  OR U9887 ( .A(n9769), .B(n9770), .Z(n9768) );
  NAND U9888 ( .A(n9770), .B(n9769), .Z(n9765) );
  ANDN U9889 ( .B(B[230]), .A(n32), .Z(n9661) );
  XNOR U9890 ( .A(n9669), .B(n9771), .Z(n9662) );
  XNOR U9891 ( .A(n9668), .B(n9666), .Z(n9771) );
  AND U9892 ( .A(n9772), .B(n9773), .Z(n9666) );
  NANDN U9893 ( .A(n9774), .B(n9775), .Z(n9773) );
  NANDN U9894 ( .A(n9776), .B(n9777), .Z(n9775) );
  NANDN U9895 ( .A(n9777), .B(n9776), .Z(n9772) );
  ANDN U9896 ( .B(B[231]), .A(n33), .Z(n9668) );
  XNOR U9897 ( .A(n9676), .B(n9778), .Z(n9669) );
  XNOR U9898 ( .A(n9675), .B(n9673), .Z(n9778) );
  AND U9899 ( .A(n9779), .B(n9780), .Z(n9673) );
  NANDN U9900 ( .A(n9781), .B(n9782), .Z(n9780) );
  OR U9901 ( .A(n9783), .B(n9784), .Z(n9782) );
  NAND U9902 ( .A(n9784), .B(n9783), .Z(n9779) );
  ANDN U9903 ( .B(B[232]), .A(n34), .Z(n9675) );
  XNOR U9904 ( .A(n9683), .B(n9785), .Z(n9676) );
  XNOR U9905 ( .A(n9682), .B(n9680), .Z(n9785) );
  AND U9906 ( .A(n9786), .B(n9787), .Z(n9680) );
  NANDN U9907 ( .A(n9788), .B(n9789), .Z(n9787) );
  NANDN U9908 ( .A(n9790), .B(n9791), .Z(n9789) );
  NANDN U9909 ( .A(n9791), .B(n9790), .Z(n9786) );
  ANDN U9910 ( .B(B[233]), .A(n35), .Z(n9682) );
  XNOR U9911 ( .A(n9690), .B(n9792), .Z(n9683) );
  XNOR U9912 ( .A(n9689), .B(n9687), .Z(n9792) );
  AND U9913 ( .A(n9793), .B(n9794), .Z(n9687) );
  NANDN U9914 ( .A(n9795), .B(n9796), .Z(n9794) );
  OR U9915 ( .A(n9797), .B(n9798), .Z(n9796) );
  NAND U9916 ( .A(n9798), .B(n9797), .Z(n9793) );
  ANDN U9917 ( .B(B[234]), .A(n36), .Z(n9689) );
  XNOR U9918 ( .A(n9697), .B(n9799), .Z(n9690) );
  XNOR U9919 ( .A(n9696), .B(n9694), .Z(n9799) );
  AND U9920 ( .A(n9800), .B(n9801), .Z(n9694) );
  NANDN U9921 ( .A(n9802), .B(n9803), .Z(n9801) );
  NANDN U9922 ( .A(n9804), .B(n9805), .Z(n9803) );
  NANDN U9923 ( .A(n9805), .B(n9804), .Z(n9800) );
  ANDN U9924 ( .B(B[235]), .A(n37), .Z(n9696) );
  XNOR U9925 ( .A(n9704), .B(n9806), .Z(n9697) );
  XNOR U9926 ( .A(n9703), .B(n9701), .Z(n9806) );
  AND U9927 ( .A(n9807), .B(n9808), .Z(n9701) );
  NANDN U9928 ( .A(n9809), .B(n9810), .Z(n9808) );
  OR U9929 ( .A(n9811), .B(n9812), .Z(n9810) );
  NAND U9930 ( .A(n9812), .B(n9811), .Z(n9807) );
  ANDN U9931 ( .B(B[236]), .A(n38), .Z(n9703) );
  XNOR U9932 ( .A(n9711), .B(n9813), .Z(n9704) );
  XNOR U9933 ( .A(n9710), .B(n9708), .Z(n9813) );
  AND U9934 ( .A(n9814), .B(n9815), .Z(n9708) );
  NANDN U9935 ( .A(n9816), .B(n9817), .Z(n9815) );
  NANDN U9936 ( .A(n9818), .B(n9819), .Z(n9817) );
  NANDN U9937 ( .A(n9819), .B(n9818), .Z(n9814) );
  ANDN U9938 ( .B(B[237]), .A(n39), .Z(n9710) );
  XNOR U9939 ( .A(n9718), .B(n9820), .Z(n9711) );
  XNOR U9940 ( .A(n9717), .B(n9715), .Z(n9820) );
  AND U9941 ( .A(n9821), .B(n9822), .Z(n9715) );
  NANDN U9942 ( .A(n9823), .B(n9824), .Z(n9822) );
  OR U9943 ( .A(n9825), .B(n9826), .Z(n9824) );
  NAND U9944 ( .A(n9826), .B(n9825), .Z(n9821) );
  ANDN U9945 ( .B(B[238]), .A(n40), .Z(n9717) );
  XNOR U9946 ( .A(n9725), .B(n9827), .Z(n9718) );
  XNOR U9947 ( .A(n9724), .B(n9722), .Z(n9827) );
  AND U9948 ( .A(n9828), .B(n9829), .Z(n9722) );
  NANDN U9949 ( .A(n9830), .B(n9831), .Z(n9829) );
  NAND U9950 ( .A(n9832), .B(n9833), .Z(n9831) );
  ANDN U9951 ( .B(B[239]), .A(n41), .Z(n9724) );
  XOR U9952 ( .A(n9731), .B(n9834), .Z(n9725) );
  XNOR U9953 ( .A(n9729), .B(n9732), .Z(n9834) );
  NAND U9954 ( .A(A[2]), .B(B[240]), .Z(n9732) );
  NANDN U9955 ( .A(n9835), .B(n9836), .Z(n9729) );
  AND U9956 ( .A(A[0]), .B(B[241]), .Z(n9836) );
  XNOR U9957 ( .A(n9734), .B(n9837), .Z(n9731) );
  NAND U9958 ( .A(A[0]), .B(B[242]), .Z(n9837) );
  NAND U9959 ( .A(B[241]), .B(A[1]), .Z(n9734) );
  NAND U9960 ( .A(n9838), .B(n9839), .Z(n253) );
  NANDN U9961 ( .A(n9840), .B(n9841), .Z(n9839) );
  OR U9962 ( .A(n9842), .B(n9843), .Z(n9841) );
  NAND U9963 ( .A(n9843), .B(n9842), .Z(n9838) );
  XOR U9964 ( .A(n235), .B(n234), .Z(\A1[23] ) );
  XOR U9965 ( .A(n8833), .B(n9844), .Z(n234) );
  XNOR U9966 ( .A(n8832), .B(n8830), .Z(n9844) );
  AND U9967 ( .A(n9845), .B(n9846), .Z(n8830) );
  NANDN U9968 ( .A(n9847), .B(n9848), .Z(n9846) );
  NANDN U9969 ( .A(n9849), .B(n9850), .Z(n9848) );
  NANDN U9970 ( .A(n9850), .B(n9849), .Z(n9845) );
  ANDN U9971 ( .B(B[10]), .A(n29), .Z(n8832) );
  XNOR U9972 ( .A(n8739), .B(n9851), .Z(n8833) );
  XNOR U9973 ( .A(n8738), .B(n8736), .Z(n9851) );
  AND U9974 ( .A(n9852), .B(n9853), .Z(n8736) );
  NANDN U9975 ( .A(n9854), .B(n9855), .Z(n9853) );
  OR U9976 ( .A(n9856), .B(n9857), .Z(n9855) );
  NAND U9977 ( .A(n9857), .B(n9856), .Z(n9852) );
  ANDN U9978 ( .B(B[11]), .A(n30), .Z(n8738) );
  XNOR U9979 ( .A(n8746), .B(n9858), .Z(n8739) );
  XNOR U9980 ( .A(n8745), .B(n8743), .Z(n9858) );
  AND U9981 ( .A(n9859), .B(n9860), .Z(n8743) );
  NANDN U9982 ( .A(n9861), .B(n9862), .Z(n9860) );
  NANDN U9983 ( .A(n9863), .B(n9864), .Z(n9862) );
  NANDN U9984 ( .A(n9864), .B(n9863), .Z(n9859) );
  ANDN U9985 ( .B(B[12]), .A(n31), .Z(n8745) );
  XNOR U9986 ( .A(n8753), .B(n9865), .Z(n8746) );
  XNOR U9987 ( .A(n8752), .B(n8750), .Z(n9865) );
  AND U9988 ( .A(n9866), .B(n9867), .Z(n8750) );
  NANDN U9989 ( .A(n9868), .B(n9869), .Z(n9867) );
  OR U9990 ( .A(n9870), .B(n9871), .Z(n9869) );
  NAND U9991 ( .A(n9871), .B(n9870), .Z(n9866) );
  ANDN U9992 ( .B(B[13]), .A(n32), .Z(n8752) );
  XNOR U9993 ( .A(n8760), .B(n9872), .Z(n8753) );
  XNOR U9994 ( .A(n8759), .B(n8757), .Z(n9872) );
  AND U9995 ( .A(n9873), .B(n9874), .Z(n8757) );
  NANDN U9996 ( .A(n9875), .B(n9876), .Z(n9874) );
  NANDN U9997 ( .A(n9877), .B(n9878), .Z(n9876) );
  NANDN U9998 ( .A(n9878), .B(n9877), .Z(n9873) );
  ANDN U9999 ( .B(B[14]), .A(n33), .Z(n8759) );
  XNOR U10000 ( .A(n8767), .B(n9879), .Z(n8760) );
  XNOR U10001 ( .A(n8766), .B(n8764), .Z(n9879) );
  AND U10002 ( .A(n9880), .B(n9881), .Z(n8764) );
  NANDN U10003 ( .A(n9882), .B(n9883), .Z(n9881) );
  OR U10004 ( .A(n9884), .B(n9885), .Z(n9883) );
  NAND U10005 ( .A(n9885), .B(n9884), .Z(n9880) );
  ANDN U10006 ( .B(B[15]), .A(n34), .Z(n8766) );
  XNOR U10007 ( .A(n8774), .B(n9886), .Z(n8767) );
  XNOR U10008 ( .A(n8773), .B(n8771), .Z(n9886) );
  AND U10009 ( .A(n9887), .B(n9888), .Z(n8771) );
  NANDN U10010 ( .A(n9889), .B(n9890), .Z(n9888) );
  NANDN U10011 ( .A(n9891), .B(n9892), .Z(n9890) );
  NANDN U10012 ( .A(n9892), .B(n9891), .Z(n9887) );
  ANDN U10013 ( .B(B[16]), .A(n35), .Z(n8773) );
  XNOR U10014 ( .A(n8781), .B(n9893), .Z(n8774) );
  XNOR U10015 ( .A(n8780), .B(n8778), .Z(n9893) );
  AND U10016 ( .A(n9894), .B(n9895), .Z(n8778) );
  NANDN U10017 ( .A(n9896), .B(n9897), .Z(n9895) );
  OR U10018 ( .A(n9898), .B(n9899), .Z(n9897) );
  NAND U10019 ( .A(n9899), .B(n9898), .Z(n9894) );
  ANDN U10020 ( .B(B[17]), .A(n36), .Z(n8780) );
  XNOR U10021 ( .A(n8788), .B(n9900), .Z(n8781) );
  XNOR U10022 ( .A(n8787), .B(n8785), .Z(n9900) );
  AND U10023 ( .A(n9901), .B(n9902), .Z(n8785) );
  NANDN U10024 ( .A(n9903), .B(n9904), .Z(n9902) );
  NANDN U10025 ( .A(n9905), .B(n9906), .Z(n9904) );
  NANDN U10026 ( .A(n9906), .B(n9905), .Z(n9901) );
  ANDN U10027 ( .B(B[18]), .A(n37), .Z(n8787) );
  XNOR U10028 ( .A(n8795), .B(n9907), .Z(n8788) );
  XNOR U10029 ( .A(n8794), .B(n8792), .Z(n9907) );
  AND U10030 ( .A(n9908), .B(n9909), .Z(n8792) );
  NANDN U10031 ( .A(n9910), .B(n9911), .Z(n9909) );
  OR U10032 ( .A(n9912), .B(n9913), .Z(n9911) );
  NAND U10033 ( .A(n9913), .B(n9912), .Z(n9908) );
  ANDN U10034 ( .B(B[19]), .A(n38), .Z(n8794) );
  XNOR U10035 ( .A(n8802), .B(n9914), .Z(n8795) );
  XNOR U10036 ( .A(n8801), .B(n8799), .Z(n9914) );
  AND U10037 ( .A(n9915), .B(n9916), .Z(n8799) );
  NANDN U10038 ( .A(n9917), .B(n9918), .Z(n9916) );
  NANDN U10039 ( .A(n9919), .B(n9920), .Z(n9918) );
  NANDN U10040 ( .A(n9920), .B(n9919), .Z(n9915) );
  ANDN U10041 ( .B(B[20]), .A(n39), .Z(n8801) );
  XNOR U10042 ( .A(n8809), .B(n9921), .Z(n8802) );
  XNOR U10043 ( .A(n8808), .B(n8806), .Z(n9921) );
  AND U10044 ( .A(n9922), .B(n9923), .Z(n8806) );
  NANDN U10045 ( .A(n9924), .B(n9925), .Z(n9923) );
  OR U10046 ( .A(n9926), .B(n9927), .Z(n9925) );
  NAND U10047 ( .A(n9927), .B(n9926), .Z(n9922) );
  ANDN U10048 ( .B(B[21]), .A(n40), .Z(n8808) );
  XNOR U10049 ( .A(n8816), .B(n9928), .Z(n8809) );
  XNOR U10050 ( .A(n8815), .B(n8813), .Z(n9928) );
  AND U10051 ( .A(n9929), .B(n9930), .Z(n8813) );
  NANDN U10052 ( .A(n9931), .B(n9932), .Z(n9930) );
  NAND U10053 ( .A(n9933), .B(n9934), .Z(n9932) );
  ANDN U10054 ( .B(B[22]), .A(n41), .Z(n8815) );
  XOR U10055 ( .A(n8822), .B(n9935), .Z(n8816) );
  XNOR U10056 ( .A(n8820), .B(n8823), .Z(n9935) );
  NAND U10057 ( .A(A[2]), .B(B[23]), .Z(n8823) );
  NANDN U10058 ( .A(n9936), .B(n9937), .Z(n8820) );
  AND U10059 ( .A(A[0]), .B(B[24]), .Z(n9937) );
  XNOR U10060 ( .A(n8825), .B(n9938), .Z(n8822) );
  NAND U10061 ( .A(A[0]), .B(B[25]), .Z(n9938) );
  NAND U10062 ( .A(B[24]), .B(A[1]), .Z(n8825) );
  NAND U10063 ( .A(n9939), .B(n9940), .Z(n235) );
  NANDN U10064 ( .A(n9941), .B(n9942), .Z(n9940) );
  OR U10065 ( .A(n9943), .B(n9944), .Z(n9942) );
  NAND U10066 ( .A(n9944), .B(n9943), .Z(n9939) );
  XOR U10067 ( .A(n255), .B(n254), .Z(\A1[239] ) );
  XOR U10068 ( .A(n9843), .B(n9945), .Z(n254) );
  XNOR U10069 ( .A(n9842), .B(n9840), .Z(n9945) );
  AND U10070 ( .A(n9946), .B(n9947), .Z(n9840) );
  NANDN U10071 ( .A(n9948), .B(n9949), .Z(n9947) );
  NANDN U10072 ( .A(n9950), .B(n9951), .Z(n9949) );
  NANDN U10073 ( .A(n9951), .B(n9950), .Z(n9946) );
  ANDN U10074 ( .B(B[226]), .A(n29), .Z(n9842) );
  XNOR U10075 ( .A(n9749), .B(n9952), .Z(n9843) );
  XNOR U10076 ( .A(n9748), .B(n9746), .Z(n9952) );
  AND U10077 ( .A(n9953), .B(n9954), .Z(n9746) );
  NANDN U10078 ( .A(n9955), .B(n9956), .Z(n9954) );
  OR U10079 ( .A(n9957), .B(n9958), .Z(n9956) );
  NAND U10080 ( .A(n9958), .B(n9957), .Z(n9953) );
  ANDN U10081 ( .B(B[227]), .A(n30), .Z(n9748) );
  XNOR U10082 ( .A(n9756), .B(n9959), .Z(n9749) );
  XNOR U10083 ( .A(n9755), .B(n9753), .Z(n9959) );
  AND U10084 ( .A(n9960), .B(n9961), .Z(n9753) );
  NANDN U10085 ( .A(n9962), .B(n9963), .Z(n9961) );
  NANDN U10086 ( .A(n9964), .B(n9965), .Z(n9963) );
  NANDN U10087 ( .A(n9965), .B(n9964), .Z(n9960) );
  ANDN U10088 ( .B(B[228]), .A(n31), .Z(n9755) );
  XNOR U10089 ( .A(n9763), .B(n9966), .Z(n9756) );
  XNOR U10090 ( .A(n9762), .B(n9760), .Z(n9966) );
  AND U10091 ( .A(n9967), .B(n9968), .Z(n9760) );
  NANDN U10092 ( .A(n9969), .B(n9970), .Z(n9968) );
  OR U10093 ( .A(n9971), .B(n9972), .Z(n9970) );
  NAND U10094 ( .A(n9972), .B(n9971), .Z(n9967) );
  ANDN U10095 ( .B(B[229]), .A(n32), .Z(n9762) );
  XNOR U10096 ( .A(n9770), .B(n9973), .Z(n9763) );
  XNOR U10097 ( .A(n9769), .B(n9767), .Z(n9973) );
  AND U10098 ( .A(n9974), .B(n9975), .Z(n9767) );
  NANDN U10099 ( .A(n9976), .B(n9977), .Z(n9975) );
  NANDN U10100 ( .A(n9978), .B(n9979), .Z(n9977) );
  NANDN U10101 ( .A(n9979), .B(n9978), .Z(n9974) );
  ANDN U10102 ( .B(B[230]), .A(n33), .Z(n9769) );
  XNOR U10103 ( .A(n9777), .B(n9980), .Z(n9770) );
  XNOR U10104 ( .A(n9776), .B(n9774), .Z(n9980) );
  AND U10105 ( .A(n9981), .B(n9982), .Z(n9774) );
  NANDN U10106 ( .A(n9983), .B(n9984), .Z(n9982) );
  OR U10107 ( .A(n9985), .B(n9986), .Z(n9984) );
  NAND U10108 ( .A(n9986), .B(n9985), .Z(n9981) );
  ANDN U10109 ( .B(B[231]), .A(n34), .Z(n9776) );
  XNOR U10110 ( .A(n9784), .B(n9987), .Z(n9777) );
  XNOR U10111 ( .A(n9783), .B(n9781), .Z(n9987) );
  AND U10112 ( .A(n9988), .B(n9989), .Z(n9781) );
  NANDN U10113 ( .A(n9990), .B(n9991), .Z(n9989) );
  NANDN U10114 ( .A(n9992), .B(n9993), .Z(n9991) );
  NANDN U10115 ( .A(n9993), .B(n9992), .Z(n9988) );
  ANDN U10116 ( .B(B[232]), .A(n35), .Z(n9783) );
  XNOR U10117 ( .A(n9791), .B(n9994), .Z(n9784) );
  XNOR U10118 ( .A(n9790), .B(n9788), .Z(n9994) );
  AND U10119 ( .A(n9995), .B(n9996), .Z(n9788) );
  NANDN U10120 ( .A(n9997), .B(n9998), .Z(n9996) );
  OR U10121 ( .A(n9999), .B(n10000), .Z(n9998) );
  NAND U10122 ( .A(n10000), .B(n9999), .Z(n9995) );
  ANDN U10123 ( .B(B[233]), .A(n36), .Z(n9790) );
  XNOR U10124 ( .A(n9798), .B(n10001), .Z(n9791) );
  XNOR U10125 ( .A(n9797), .B(n9795), .Z(n10001) );
  AND U10126 ( .A(n10002), .B(n10003), .Z(n9795) );
  NANDN U10127 ( .A(n10004), .B(n10005), .Z(n10003) );
  NANDN U10128 ( .A(n10006), .B(n10007), .Z(n10005) );
  NANDN U10129 ( .A(n10007), .B(n10006), .Z(n10002) );
  ANDN U10130 ( .B(B[234]), .A(n37), .Z(n9797) );
  XNOR U10131 ( .A(n9805), .B(n10008), .Z(n9798) );
  XNOR U10132 ( .A(n9804), .B(n9802), .Z(n10008) );
  AND U10133 ( .A(n10009), .B(n10010), .Z(n9802) );
  NANDN U10134 ( .A(n10011), .B(n10012), .Z(n10010) );
  OR U10135 ( .A(n10013), .B(n10014), .Z(n10012) );
  NAND U10136 ( .A(n10014), .B(n10013), .Z(n10009) );
  ANDN U10137 ( .B(B[235]), .A(n38), .Z(n9804) );
  XNOR U10138 ( .A(n9812), .B(n10015), .Z(n9805) );
  XNOR U10139 ( .A(n9811), .B(n9809), .Z(n10015) );
  AND U10140 ( .A(n10016), .B(n10017), .Z(n9809) );
  NANDN U10141 ( .A(n10018), .B(n10019), .Z(n10017) );
  NANDN U10142 ( .A(n10020), .B(n10021), .Z(n10019) );
  NANDN U10143 ( .A(n10021), .B(n10020), .Z(n10016) );
  ANDN U10144 ( .B(B[236]), .A(n39), .Z(n9811) );
  XNOR U10145 ( .A(n9819), .B(n10022), .Z(n9812) );
  XNOR U10146 ( .A(n9818), .B(n9816), .Z(n10022) );
  AND U10147 ( .A(n10023), .B(n10024), .Z(n9816) );
  NANDN U10148 ( .A(n10025), .B(n10026), .Z(n10024) );
  OR U10149 ( .A(n10027), .B(n10028), .Z(n10026) );
  NAND U10150 ( .A(n10028), .B(n10027), .Z(n10023) );
  ANDN U10151 ( .B(B[237]), .A(n40), .Z(n9818) );
  XNOR U10152 ( .A(n9826), .B(n10029), .Z(n9819) );
  XNOR U10153 ( .A(n9825), .B(n9823), .Z(n10029) );
  AND U10154 ( .A(n10030), .B(n10031), .Z(n9823) );
  NANDN U10155 ( .A(n10032), .B(n10033), .Z(n10031) );
  NAND U10156 ( .A(n10034), .B(n10035), .Z(n10033) );
  ANDN U10157 ( .B(B[238]), .A(n41), .Z(n9825) );
  XOR U10158 ( .A(n9832), .B(n10036), .Z(n9826) );
  XNOR U10159 ( .A(n9830), .B(n9833), .Z(n10036) );
  NAND U10160 ( .A(A[2]), .B(B[239]), .Z(n9833) );
  NANDN U10161 ( .A(n10037), .B(n10038), .Z(n9830) );
  AND U10162 ( .A(A[0]), .B(B[240]), .Z(n10038) );
  XNOR U10163 ( .A(n9835), .B(n10039), .Z(n9832) );
  NAND U10164 ( .A(A[0]), .B(B[241]), .Z(n10039) );
  NAND U10165 ( .A(B[240]), .B(A[1]), .Z(n9835) );
  NAND U10166 ( .A(n10040), .B(n10041), .Z(n255) );
  NANDN U10167 ( .A(n10042), .B(n10043), .Z(n10041) );
  OR U10168 ( .A(n10044), .B(n10045), .Z(n10043) );
  NAND U10169 ( .A(n10045), .B(n10044), .Z(n10040) );
  XOR U10170 ( .A(n259), .B(n258), .Z(\A1[238] ) );
  XOR U10171 ( .A(n10045), .B(n10046), .Z(n258) );
  XNOR U10172 ( .A(n10044), .B(n10042), .Z(n10046) );
  AND U10173 ( .A(n10047), .B(n10048), .Z(n10042) );
  NANDN U10174 ( .A(n10049), .B(n10050), .Z(n10048) );
  NANDN U10175 ( .A(n10051), .B(n10052), .Z(n10050) );
  NANDN U10176 ( .A(n10052), .B(n10051), .Z(n10047) );
  ANDN U10177 ( .B(B[225]), .A(n29), .Z(n10044) );
  XNOR U10178 ( .A(n9951), .B(n10053), .Z(n10045) );
  XNOR U10179 ( .A(n9950), .B(n9948), .Z(n10053) );
  AND U10180 ( .A(n10054), .B(n10055), .Z(n9948) );
  NANDN U10181 ( .A(n10056), .B(n10057), .Z(n10055) );
  OR U10182 ( .A(n10058), .B(n10059), .Z(n10057) );
  NAND U10183 ( .A(n10059), .B(n10058), .Z(n10054) );
  ANDN U10184 ( .B(B[226]), .A(n30), .Z(n9950) );
  XNOR U10185 ( .A(n9958), .B(n10060), .Z(n9951) );
  XNOR U10186 ( .A(n9957), .B(n9955), .Z(n10060) );
  AND U10187 ( .A(n10061), .B(n10062), .Z(n9955) );
  NANDN U10188 ( .A(n10063), .B(n10064), .Z(n10062) );
  NANDN U10189 ( .A(n10065), .B(n10066), .Z(n10064) );
  NANDN U10190 ( .A(n10066), .B(n10065), .Z(n10061) );
  ANDN U10191 ( .B(B[227]), .A(n31), .Z(n9957) );
  XNOR U10192 ( .A(n9965), .B(n10067), .Z(n9958) );
  XNOR U10193 ( .A(n9964), .B(n9962), .Z(n10067) );
  AND U10194 ( .A(n10068), .B(n10069), .Z(n9962) );
  NANDN U10195 ( .A(n10070), .B(n10071), .Z(n10069) );
  OR U10196 ( .A(n10072), .B(n10073), .Z(n10071) );
  NAND U10197 ( .A(n10073), .B(n10072), .Z(n10068) );
  ANDN U10198 ( .B(B[228]), .A(n32), .Z(n9964) );
  XNOR U10199 ( .A(n9972), .B(n10074), .Z(n9965) );
  XNOR U10200 ( .A(n9971), .B(n9969), .Z(n10074) );
  AND U10201 ( .A(n10075), .B(n10076), .Z(n9969) );
  NANDN U10202 ( .A(n10077), .B(n10078), .Z(n10076) );
  NANDN U10203 ( .A(n10079), .B(n10080), .Z(n10078) );
  NANDN U10204 ( .A(n10080), .B(n10079), .Z(n10075) );
  ANDN U10205 ( .B(B[229]), .A(n33), .Z(n9971) );
  XNOR U10206 ( .A(n9979), .B(n10081), .Z(n9972) );
  XNOR U10207 ( .A(n9978), .B(n9976), .Z(n10081) );
  AND U10208 ( .A(n10082), .B(n10083), .Z(n9976) );
  NANDN U10209 ( .A(n10084), .B(n10085), .Z(n10083) );
  OR U10210 ( .A(n10086), .B(n10087), .Z(n10085) );
  NAND U10211 ( .A(n10087), .B(n10086), .Z(n10082) );
  ANDN U10212 ( .B(B[230]), .A(n34), .Z(n9978) );
  XNOR U10213 ( .A(n9986), .B(n10088), .Z(n9979) );
  XNOR U10214 ( .A(n9985), .B(n9983), .Z(n10088) );
  AND U10215 ( .A(n10089), .B(n10090), .Z(n9983) );
  NANDN U10216 ( .A(n10091), .B(n10092), .Z(n10090) );
  NANDN U10217 ( .A(n10093), .B(n10094), .Z(n10092) );
  NANDN U10218 ( .A(n10094), .B(n10093), .Z(n10089) );
  ANDN U10219 ( .B(B[231]), .A(n35), .Z(n9985) );
  XNOR U10220 ( .A(n9993), .B(n10095), .Z(n9986) );
  XNOR U10221 ( .A(n9992), .B(n9990), .Z(n10095) );
  AND U10222 ( .A(n10096), .B(n10097), .Z(n9990) );
  NANDN U10223 ( .A(n10098), .B(n10099), .Z(n10097) );
  OR U10224 ( .A(n10100), .B(n10101), .Z(n10099) );
  NAND U10225 ( .A(n10101), .B(n10100), .Z(n10096) );
  ANDN U10226 ( .B(B[232]), .A(n36), .Z(n9992) );
  XNOR U10227 ( .A(n10000), .B(n10102), .Z(n9993) );
  XNOR U10228 ( .A(n9999), .B(n9997), .Z(n10102) );
  AND U10229 ( .A(n10103), .B(n10104), .Z(n9997) );
  NANDN U10230 ( .A(n10105), .B(n10106), .Z(n10104) );
  NANDN U10231 ( .A(n10107), .B(n10108), .Z(n10106) );
  NANDN U10232 ( .A(n10108), .B(n10107), .Z(n10103) );
  ANDN U10233 ( .B(B[233]), .A(n37), .Z(n9999) );
  XNOR U10234 ( .A(n10007), .B(n10109), .Z(n10000) );
  XNOR U10235 ( .A(n10006), .B(n10004), .Z(n10109) );
  AND U10236 ( .A(n10110), .B(n10111), .Z(n10004) );
  NANDN U10237 ( .A(n10112), .B(n10113), .Z(n10111) );
  OR U10238 ( .A(n10114), .B(n10115), .Z(n10113) );
  NAND U10239 ( .A(n10115), .B(n10114), .Z(n10110) );
  ANDN U10240 ( .B(B[234]), .A(n38), .Z(n10006) );
  XNOR U10241 ( .A(n10014), .B(n10116), .Z(n10007) );
  XNOR U10242 ( .A(n10013), .B(n10011), .Z(n10116) );
  AND U10243 ( .A(n10117), .B(n10118), .Z(n10011) );
  NANDN U10244 ( .A(n10119), .B(n10120), .Z(n10118) );
  NANDN U10245 ( .A(n10121), .B(n10122), .Z(n10120) );
  NANDN U10246 ( .A(n10122), .B(n10121), .Z(n10117) );
  ANDN U10247 ( .B(B[235]), .A(n39), .Z(n10013) );
  XNOR U10248 ( .A(n10021), .B(n10123), .Z(n10014) );
  XNOR U10249 ( .A(n10020), .B(n10018), .Z(n10123) );
  AND U10250 ( .A(n10124), .B(n10125), .Z(n10018) );
  NANDN U10251 ( .A(n10126), .B(n10127), .Z(n10125) );
  OR U10252 ( .A(n10128), .B(n10129), .Z(n10127) );
  NAND U10253 ( .A(n10129), .B(n10128), .Z(n10124) );
  ANDN U10254 ( .B(B[236]), .A(n40), .Z(n10020) );
  XNOR U10255 ( .A(n10028), .B(n10130), .Z(n10021) );
  XNOR U10256 ( .A(n10027), .B(n10025), .Z(n10130) );
  AND U10257 ( .A(n10131), .B(n10132), .Z(n10025) );
  NANDN U10258 ( .A(n10133), .B(n10134), .Z(n10132) );
  NAND U10259 ( .A(n10135), .B(n10136), .Z(n10134) );
  ANDN U10260 ( .B(B[237]), .A(n41), .Z(n10027) );
  XOR U10261 ( .A(n10034), .B(n10137), .Z(n10028) );
  XNOR U10262 ( .A(n10032), .B(n10035), .Z(n10137) );
  NAND U10263 ( .A(A[2]), .B(B[238]), .Z(n10035) );
  NANDN U10264 ( .A(n10138), .B(n10139), .Z(n10032) );
  AND U10265 ( .A(A[0]), .B(B[239]), .Z(n10139) );
  XNOR U10266 ( .A(n10037), .B(n10140), .Z(n10034) );
  NAND U10267 ( .A(A[0]), .B(B[240]), .Z(n10140) );
  NAND U10268 ( .A(B[239]), .B(A[1]), .Z(n10037) );
  NAND U10269 ( .A(n10141), .B(n10142), .Z(n259) );
  NANDN U10270 ( .A(n10143), .B(n10144), .Z(n10142) );
  OR U10271 ( .A(n10145), .B(n10146), .Z(n10144) );
  NAND U10272 ( .A(n10146), .B(n10145), .Z(n10141) );
  XOR U10273 ( .A(n261), .B(n260), .Z(\A1[237] ) );
  XOR U10274 ( .A(n10146), .B(n10147), .Z(n260) );
  XNOR U10275 ( .A(n10145), .B(n10143), .Z(n10147) );
  AND U10276 ( .A(n10148), .B(n10149), .Z(n10143) );
  NANDN U10277 ( .A(n10150), .B(n10151), .Z(n10149) );
  NANDN U10278 ( .A(n10152), .B(n10153), .Z(n10151) );
  NANDN U10279 ( .A(n10153), .B(n10152), .Z(n10148) );
  ANDN U10280 ( .B(B[224]), .A(n29), .Z(n10145) );
  XNOR U10281 ( .A(n10052), .B(n10154), .Z(n10146) );
  XNOR U10282 ( .A(n10051), .B(n10049), .Z(n10154) );
  AND U10283 ( .A(n10155), .B(n10156), .Z(n10049) );
  NANDN U10284 ( .A(n10157), .B(n10158), .Z(n10156) );
  OR U10285 ( .A(n10159), .B(n10160), .Z(n10158) );
  NAND U10286 ( .A(n10160), .B(n10159), .Z(n10155) );
  ANDN U10287 ( .B(B[225]), .A(n30), .Z(n10051) );
  XNOR U10288 ( .A(n10059), .B(n10161), .Z(n10052) );
  XNOR U10289 ( .A(n10058), .B(n10056), .Z(n10161) );
  AND U10290 ( .A(n10162), .B(n10163), .Z(n10056) );
  NANDN U10291 ( .A(n10164), .B(n10165), .Z(n10163) );
  NANDN U10292 ( .A(n10166), .B(n10167), .Z(n10165) );
  NANDN U10293 ( .A(n10167), .B(n10166), .Z(n10162) );
  ANDN U10294 ( .B(B[226]), .A(n31), .Z(n10058) );
  XNOR U10295 ( .A(n10066), .B(n10168), .Z(n10059) );
  XNOR U10296 ( .A(n10065), .B(n10063), .Z(n10168) );
  AND U10297 ( .A(n10169), .B(n10170), .Z(n10063) );
  NANDN U10298 ( .A(n10171), .B(n10172), .Z(n10170) );
  OR U10299 ( .A(n10173), .B(n10174), .Z(n10172) );
  NAND U10300 ( .A(n10174), .B(n10173), .Z(n10169) );
  ANDN U10301 ( .B(B[227]), .A(n32), .Z(n10065) );
  XNOR U10302 ( .A(n10073), .B(n10175), .Z(n10066) );
  XNOR U10303 ( .A(n10072), .B(n10070), .Z(n10175) );
  AND U10304 ( .A(n10176), .B(n10177), .Z(n10070) );
  NANDN U10305 ( .A(n10178), .B(n10179), .Z(n10177) );
  NANDN U10306 ( .A(n10180), .B(n10181), .Z(n10179) );
  NANDN U10307 ( .A(n10181), .B(n10180), .Z(n10176) );
  ANDN U10308 ( .B(B[228]), .A(n33), .Z(n10072) );
  XNOR U10309 ( .A(n10080), .B(n10182), .Z(n10073) );
  XNOR U10310 ( .A(n10079), .B(n10077), .Z(n10182) );
  AND U10311 ( .A(n10183), .B(n10184), .Z(n10077) );
  NANDN U10312 ( .A(n10185), .B(n10186), .Z(n10184) );
  OR U10313 ( .A(n10187), .B(n10188), .Z(n10186) );
  NAND U10314 ( .A(n10188), .B(n10187), .Z(n10183) );
  ANDN U10315 ( .B(B[229]), .A(n34), .Z(n10079) );
  XNOR U10316 ( .A(n10087), .B(n10189), .Z(n10080) );
  XNOR U10317 ( .A(n10086), .B(n10084), .Z(n10189) );
  AND U10318 ( .A(n10190), .B(n10191), .Z(n10084) );
  NANDN U10319 ( .A(n10192), .B(n10193), .Z(n10191) );
  NANDN U10320 ( .A(n10194), .B(n10195), .Z(n10193) );
  NANDN U10321 ( .A(n10195), .B(n10194), .Z(n10190) );
  ANDN U10322 ( .B(B[230]), .A(n35), .Z(n10086) );
  XNOR U10323 ( .A(n10094), .B(n10196), .Z(n10087) );
  XNOR U10324 ( .A(n10093), .B(n10091), .Z(n10196) );
  AND U10325 ( .A(n10197), .B(n10198), .Z(n10091) );
  NANDN U10326 ( .A(n10199), .B(n10200), .Z(n10198) );
  OR U10327 ( .A(n10201), .B(n10202), .Z(n10200) );
  NAND U10328 ( .A(n10202), .B(n10201), .Z(n10197) );
  ANDN U10329 ( .B(B[231]), .A(n36), .Z(n10093) );
  XNOR U10330 ( .A(n10101), .B(n10203), .Z(n10094) );
  XNOR U10331 ( .A(n10100), .B(n10098), .Z(n10203) );
  AND U10332 ( .A(n10204), .B(n10205), .Z(n10098) );
  NANDN U10333 ( .A(n10206), .B(n10207), .Z(n10205) );
  NANDN U10334 ( .A(n10208), .B(n10209), .Z(n10207) );
  NANDN U10335 ( .A(n10209), .B(n10208), .Z(n10204) );
  ANDN U10336 ( .B(B[232]), .A(n37), .Z(n10100) );
  XNOR U10337 ( .A(n10108), .B(n10210), .Z(n10101) );
  XNOR U10338 ( .A(n10107), .B(n10105), .Z(n10210) );
  AND U10339 ( .A(n10211), .B(n10212), .Z(n10105) );
  NANDN U10340 ( .A(n10213), .B(n10214), .Z(n10212) );
  OR U10341 ( .A(n10215), .B(n10216), .Z(n10214) );
  NAND U10342 ( .A(n10216), .B(n10215), .Z(n10211) );
  ANDN U10343 ( .B(B[233]), .A(n38), .Z(n10107) );
  XNOR U10344 ( .A(n10115), .B(n10217), .Z(n10108) );
  XNOR U10345 ( .A(n10114), .B(n10112), .Z(n10217) );
  AND U10346 ( .A(n10218), .B(n10219), .Z(n10112) );
  NANDN U10347 ( .A(n10220), .B(n10221), .Z(n10219) );
  NANDN U10348 ( .A(n10222), .B(n10223), .Z(n10221) );
  NANDN U10349 ( .A(n10223), .B(n10222), .Z(n10218) );
  ANDN U10350 ( .B(B[234]), .A(n39), .Z(n10114) );
  XNOR U10351 ( .A(n10122), .B(n10224), .Z(n10115) );
  XNOR U10352 ( .A(n10121), .B(n10119), .Z(n10224) );
  AND U10353 ( .A(n10225), .B(n10226), .Z(n10119) );
  NANDN U10354 ( .A(n10227), .B(n10228), .Z(n10226) );
  OR U10355 ( .A(n10229), .B(n10230), .Z(n10228) );
  NAND U10356 ( .A(n10230), .B(n10229), .Z(n10225) );
  ANDN U10357 ( .B(B[235]), .A(n40), .Z(n10121) );
  XNOR U10358 ( .A(n10129), .B(n10231), .Z(n10122) );
  XNOR U10359 ( .A(n10128), .B(n10126), .Z(n10231) );
  AND U10360 ( .A(n10232), .B(n10233), .Z(n10126) );
  NANDN U10361 ( .A(n10234), .B(n10235), .Z(n10233) );
  NAND U10362 ( .A(n10236), .B(n10237), .Z(n10235) );
  ANDN U10363 ( .B(B[236]), .A(n41), .Z(n10128) );
  XOR U10364 ( .A(n10135), .B(n10238), .Z(n10129) );
  XNOR U10365 ( .A(n10133), .B(n10136), .Z(n10238) );
  NAND U10366 ( .A(A[2]), .B(B[237]), .Z(n10136) );
  NANDN U10367 ( .A(n10239), .B(n10240), .Z(n10133) );
  AND U10368 ( .A(A[0]), .B(B[238]), .Z(n10240) );
  XNOR U10369 ( .A(n10138), .B(n10241), .Z(n10135) );
  NAND U10370 ( .A(A[0]), .B(B[239]), .Z(n10241) );
  NAND U10371 ( .A(B[238]), .B(A[1]), .Z(n10138) );
  NAND U10372 ( .A(n10242), .B(n10243), .Z(n261) );
  NANDN U10373 ( .A(n10244), .B(n10245), .Z(n10243) );
  OR U10374 ( .A(n10246), .B(n10247), .Z(n10245) );
  NAND U10375 ( .A(n10247), .B(n10246), .Z(n10242) );
  XOR U10376 ( .A(n263), .B(n262), .Z(\A1[236] ) );
  XOR U10377 ( .A(n10247), .B(n10248), .Z(n262) );
  XNOR U10378 ( .A(n10246), .B(n10244), .Z(n10248) );
  AND U10379 ( .A(n10249), .B(n10250), .Z(n10244) );
  NANDN U10380 ( .A(n10251), .B(n10252), .Z(n10250) );
  NANDN U10381 ( .A(n10253), .B(n10254), .Z(n10252) );
  NANDN U10382 ( .A(n10254), .B(n10253), .Z(n10249) );
  ANDN U10383 ( .B(B[223]), .A(n29), .Z(n10246) );
  XNOR U10384 ( .A(n10153), .B(n10255), .Z(n10247) );
  XNOR U10385 ( .A(n10152), .B(n10150), .Z(n10255) );
  AND U10386 ( .A(n10256), .B(n10257), .Z(n10150) );
  NANDN U10387 ( .A(n10258), .B(n10259), .Z(n10257) );
  OR U10388 ( .A(n10260), .B(n10261), .Z(n10259) );
  NAND U10389 ( .A(n10261), .B(n10260), .Z(n10256) );
  ANDN U10390 ( .B(B[224]), .A(n30), .Z(n10152) );
  XNOR U10391 ( .A(n10160), .B(n10262), .Z(n10153) );
  XNOR U10392 ( .A(n10159), .B(n10157), .Z(n10262) );
  AND U10393 ( .A(n10263), .B(n10264), .Z(n10157) );
  NANDN U10394 ( .A(n10265), .B(n10266), .Z(n10264) );
  NANDN U10395 ( .A(n10267), .B(n10268), .Z(n10266) );
  NANDN U10396 ( .A(n10268), .B(n10267), .Z(n10263) );
  ANDN U10397 ( .B(B[225]), .A(n31), .Z(n10159) );
  XNOR U10398 ( .A(n10167), .B(n10269), .Z(n10160) );
  XNOR U10399 ( .A(n10166), .B(n10164), .Z(n10269) );
  AND U10400 ( .A(n10270), .B(n10271), .Z(n10164) );
  NANDN U10401 ( .A(n10272), .B(n10273), .Z(n10271) );
  OR U10402 ( .A(n10274), .B(n10275), .Z(n10273) );
  NAND U10403 ( .A(n10275), .B(n10274), .Z(n10270) );
  ANDN U10404 ( .B(B[226]), .A(n32), .Z(n10166) );
  XNOR U10405 ( .A(n10174), .B(n10276), .Z(n10167) );
  XNOR U10406 ( .A(n10173), .B(n10171), .Z(n10276) );
  AND U10407 ( .A(n10277), .B(n10278), .Z(n10171) );
  NANDN U10408 ( .A(n10279), .B(n10280), .Z(n10278) );
  NANDN U10409 ( .A(n10281), .B(n10282), .Z(n10280) );
  NANDN U10410 ( .A(n10282), .B(n10281), .Z(n10277) );
  ANDN U10411 ( .B(B[227]), .A(n33), .Z(n10173) );
  XNOR U10412 ( .A(n10181), .B(n10283), .Z(n10174) );
  XNOR U10413 ( .A(n10180), .B(n10178), .Z(n10283) );
  AND U10414 ( .A(n10284), .B(n10285), .Z(n10178) );
  NANDN U10415 ( .A(n10286), .B(n10287), .Z(n10285) );
  OR U10416 ( .A(n10288), .B(n10289), .Z(n10287) );
  NAND U10417 ( .A(n10289), .B(n10288), .Z(n10284) );
  ANDN U10418 ( .B(B[228]), .A(n34), .Z(n10180) );
  XNOR U10419 ( .A(n10188), .B(n10290), .Z(n10181) );
  XNOR U10420 ( .A(n10187), .B(n10185), .Z(n10290) );
  AND U10421 ( .A(n10291), .B(n10292), .Z(n10185) );
  NANDN U10422 ( .A(n10293), .B(n10294), .Z(n10292) );
  NANDN U10423 ( .A(n10295), .B(n10296), .Z(n10294) );
  NANDN U10424 ( .A(n10296), .B(n10295), .Z(n10291) );
  ANDN U10425 ( .B(B[229]), .A(n35), .Z(n10187) );
  XNOR U10426 ( .A(n10195), .B(n10297), .Z(n10188) );
  XNOR U10427 ( .A(n10194), .B(n10192), .Z(n10297) );
  AND U10428 ( .A(n10298), .B(n10299), .Z(n10192) );
  NANDN U10429 ( .A(n10300), .B(n10301), .Z(n10299) );
  OR U10430 ( .A(n10302), .B(n10303), .Z(n10301) );
  NAND U10431 ( .A(n10303), .B(n10302), .Z(n10298) );
  ANDN U10432 ( .B(B[230]), .A(n36), .Z(n10194) );
  XNOR U10433 ( .A(n10202), .B(n10304), .Z(n10195) );
  XNOR U10434 ( .A(n10201), .B(n10199), .Z(n10304) );
  AND U10435 ( .A(n10305), .B(n10306), .Z(n10199) );
  NANDN U10436 ( .A(n10307), .B(n10308), .Z(n10306) );
  NANDN U10437 ( .A(n10309), .B(n10310), .Z(n10308) );
  NANDN U10438 ( .A(n10310), .B(n10309), .Z(n10305) );
  ANDN U10439 ( .B(B[231]), .A(n37), .Z(n10201) );
  XNOR U10440 ( .A(n10209), .B(n10311), .Z(n10202) );
  XNOR U10441 ( .A(n10208), .B(n10206), .Z(n10311) );
  AND U10442 ( .A(n10312), .B(n10313), .Z(n10206) );
  NANDN U10443 ( .A(n10314), .B(n10315), .Z(n10313) );
  OR U10444 ( .A(n10316), .B(n10317), .Z(n10315) );
  NAND U10445 ( .A(n10317), .B(n10316), .Z(n10312) );
  ANDN U10446 ( .B(B[232]), .A(n38), .Z(n10208) );
  XNOR U10447 ( .A(n10216), .B(n10318), .Z(n10209) );
  XNOR U10448 ( .A(n10215), .B(n10213), .Z(n10318) );
  AND U10449 ( .A(n10319), .B(n10320), .Z(n10213) );
  NANDN U10450 ( .A(n10321), .B(n10322), .Z(n10320) );
  NANDN U10451 ( .A(n10323), .B(n10324), .Z(n10322) );
  NANDN U10452 ( .A(n10324), .B(n10323), .Z(n10319) );
  ANDN U10453 ( .B(B[233]), .A(n39), .Z(n10215) );
  XNOR U10454 ( .A(n10223), .B(n10325), .Z(n10216) );
  XNOR U10455 ( .A(n10222), .B(n10220), .Z(n10325) );
  AND U10456 ( .A(n10326), .B(n10327), .Z(n10220) );
  NANDN U10457 ( .A(n10328), .B(n10329), .Z(n10327) );
  OR U10458 ( .A(n10330), .B(n10331), .Z(n10329) );
  NAND U10459 ( .A(n10331), .B(n10330), .Z(n10326) );
  ANDN U10460 ( .B(B[234]), .A(n40), .Z(n10222) );
  XNOR U10461 ( .A(n10230), .B(n10332), .Z(n10223) );
  XNOR U10462 ( .A(n10229), .B(n10227), .Z(n10332) );
  AND U10463 ( .A(n10333), .B(n10334), .Z(n10227) );
  NANDN U10464 ( .A(n10335), .B(n10336), .Z(n10334) );
  NAND U10465 ( .A(n10337), .B(n10338), .Z(n10336) );
  ANDN U10466 ( .B(B[235]), .A(n41), .Z(n10229) );
  XOR U10467 ( .A(n10236), .B(n10339), .Z(n10230) );
  XNOR U10468 ( .A(n10234), .B(n10237), .Z(n10339) );
  NAND U10469 ( .A(A[2]), .B(B[236]), .Z(n10237) );
  NANDN U10470 ( .A(n10340), .B(n10341), .Z(n10234) );
  AND U10471 ( .A(A[0]), .B(B[237]), .Z(n10341) );
  XNOR U10472 ( .A(n10239), .B(n10342), .Z(n10236) );
  NAND U10473 ( .A(A[0]), .B(B[238]), .Z(n10342) );
  NAND U10474 ( .A(B[237]), .B(A[1]), .Z(n10239) );
  NAND U10475 ( .A(n10343), .B(n10344), .Z(n263) );
  NANDN U10476 ( .A(n10345), .B(n10346), .Z(n10344) );
  OR U10477 ( .A(n10347), .B(n10348), .Z(n10346) );
  NAND U10478 ( .A(n10348), .B(n10347), .Z(n10343) );
  XOR U10479 ( .A(n265), .B(n264), .Z(\A1[235] ) );
  XOR U10480 ( .A(n10348), .B(n10349), .Z(n264) );
  XNOR U10481 ( .A(n10347), .B(n10345), .Z(n10349) );
  AND U10482 ( .A(n10350), .B(n10351), .Z(n10345) );
  NANDN U10483 ( .A(n10352), .B(n10353), .Z(n10351) );
  NANDN U10484 ( .A(n10354), .B(n10355), .Z(n10353) );
  NANDN U10485 ( .A(n10355), .B(n10354), .Z(n10350) );
  ANDN U10486 ( .B(B[222]), .A(n29), .Z(n10347) );
  XNOR U10487 ( .A(n10254), .B(n10356), .Z(n10348) );
  XNOR U10488 ( .A(n10253), .B(n10251), .Z(n10356) );
  AND U10489 ( .A(n10357), .B(n10358), .Z(n10251) );
  NANDN U10490 ( .A(n10359), .B(n10360), .Z(n10358) );
  OR U10491 ( .A(n10361), .B(n10362), .Z(n10360) );
  NAND U10492 ( .A(n10362), .B(n10361), .Z(n10357) );
  ANDN U10493 ( .B(B[223]), .A(n30), .Z(n10253) );
  XNOR U10494 ( .A(n10261), .B(n10363), .Z(n10254) );
  XNOR U10495 ( .A(n10260), .B(n10258), .Z(n10363) );
  AND U10496 ( .A(n10364), .B(n10365), .Z(n10258) );
  NANDN U10497 ( .A(n10366), .B(n10367), .Z(n10365) );
  NANDN U10498 ( .A(n10368), .B(n10369), .Z(n10367) );
  NANDN U10499 ( .A(n10369), .B(n10368), .Z(n10364) );
  ANDN U10500 ( .B(B[224]), .A(n31), .Z(n10260) );
  XNOR U10501 ( .A(n10268), .B(n10370), .Z(n10261) );
  XNOR U10502 ( .A(n10267), .B(n10265), .Z(n10370) );
  AND U10503 ( .A(n10371), .B(n10372), .Z(n10265) );
  NANDN U10504 ( .A(n10373), .B(n10374), .Z(n10372) );
  OR U10505 ( .A(n10375), .B(n10376), .Z(n10374) );
  NAND U10506 ( .A(n10376), .B(n10375), .Z(n10371) );
  ANDN U10507 ( .B(B[225]), .A(n32), .Z(n10267) );
  XNOR U10508 ( .A(n10275), .B(n10377), .Z(n10268) );
  XNOR U10509 ( .A(n10274), .B(n10272), .Z(n10377) );
  AND U10510 ( .A(n10378), .B(n10379), .Z(n10272) );
  NANDN U10511 ( .A(n10380), .B(n10381), .Z(n10379) );
  NANDN U10512 ( .A(n10382), .B(n10383), .Z(n10381) );
  NANDN U10513 ( .A(n10383), .B(n10382), .Z(n10378) );
  ANDN U10514 ( .B(B[226]), .A(n33), .Z(n10274) );
  XNOR U10515 ( .A(n10282), .B(n10384), .Z(n10275) );
  XNOR U10516 ( .A(n10281), .B(n10279), .Z(n10384) );
  AND U10517 ( .A(n10385), .B(n10386), .Z(n10279) );
  NANDN U10518 ( .A(n10387), .B(n10388), .Z(n10386) );
  OR U10519 ( .A(n10389), .B(n10390), .Z(n10388) );
  NAND U10520 ( .A(n10390), .B(n10389), .Z(n10385) );
  ANDN U10521 ( .B(B[227]), .A(n34), .Z(n10281) );
  XNOR U10522 ( .A(n10289), .B(n10391), .Z(n10282) );
  XNOR U10523 ( .A(n10288), .B(n10286), .Z(n10391) );
  AND U10524 ( .A(n10392), .B(n10393), .Z(n10286) );
  NANDN U10525 ( .A(n10394), .B(n10395), .Z(n10393) );
  NANDN U10526 ( .A(n10396), .B(n10397), .Z(n10395) );
  NANDN U10527 ( .A(n10397), .B(n10396), .Z(n10392) );
  ANDN U10528 ( .B(B[228]), .A(n35), .Z(n10288) );
  XNOR U10529 ( .A(n10296), .B(n10398), .Z(n10289) );
  XNOR U10530 ( .A(n10295), .B(n10293), .Z(n10398) );
  AND U10531 ( .A(n10399), .B(n10400), .Z(n10293) );
  NANDN U10532 ( .A(n10401), .B(n10402), .Z(n10400) );
  OR U10533 ( .A(n10403), .B(n10404), .Z(n10402) );
  NAND U10534 ( .A(n10404), .B(n10403), .Z(n10399) );
  ANDN U10535 ( .B(B[229]), .A(n36), .Z(n10295) );
  XNOR U10536 ( .A(n10303), .B(n10405), .Z(n10296) );
  XNOR U10537 ( .A(n10302), .B(n10300), .Z(n10405) );
  AND U10538 ( .A(n10406), .B(n10407), .Z(n10300) );
  NANDN U10539 ( .A(n10408), .B(n10409), .Z(n10407) );
  NANDN U10540 ( .A(n10410), .B(n10411), .Z(n10409) );
  NANDN U10541 ( .A(n10411), .B(n10410), .Z(n10406) );
  ANDN U10542 ( .B(B[230]), .A(n37), .Z(n10302) );
  XNOR U10543 ( .A(n10310), .B(n10412), .Z(n10303) );
  XNOR U10544 ( .A(n10309), .B(n10307), .Z(n10412) );
  AND U10545 ( .A(n10413), .B(n10414), .Z(n10307) );
  NANDN U10546 ( .A(n10415), .B(n10416), .Z(n10414) );
  OR U10547 ( .A(n10417), .B(n10418), .Z(n10416) );
  NAND U10548 ( .A(n10418), .B(n10417), .Z(n10413) );
  ANDN U10549 ( .B(B[231]), .A(n38), .Z(n10309) );
  XNOR U10550 ( .A(n10317), .B(n10419), .Z(n10310) );
  XNOR U10551 ( .A(n10316), .B(n10314), .Z(n10419) );
  AND U10552 ( .A(n10420), .B(n10421), .Z(n10314) );
  NANDN U10553 ( .A(n10422), .B(n10423), .Z(n10421) );
  NANDN U10554 ( .A(n10424), .B(n10425), .Z(n10423) );
  NANDN U10555 ( .A(n10425), .B(n10424), .Z(n10420) );
  ANDN U10556 ( .B(B[232]), .A(n39), .Z(n10316) );
  XNOR U10557 ( .A(n10324), .B(n10426), .Z(n10317) );
  XNOR U10558 ( .A(n10323), .B(n10321), .Z(n10426) );
  AND U10559 ( .A(n10427), .B(n10428), .Z(n10321) );
  NANDN U10560 ( .A(n10429), .B(n10430), .Z(n10428) );
  OR U10561 ( .A(n10431), .B(n10432), .Z(n10430) );
  NAND U10562 ( .A(n10432), .B(n10431), .Z(n10427) );
  ANDN U10563 ( .B(B[233]), .A(n40), .Z(n10323) );
  XNOR U10564 ( .A(n10331), .B(n10433), .Z(n10324) );
  XNOR U10565 ( .A(n10330), .B(n10328), .Z(n10433) );
  AND U10566 ( .A(n10434), .B(n10435), .Z(n10328) );
  NANDN U10567 ( .A(n10436), .B(n10437), .Z(n10435) );
  NAND U10568 ( .A(n10438), .B(n10439), .Z(n10437) );
  ANDN U10569 ( .B(B[234]), .A(n41), .Z(n10330) );
  XOR U10570 ( .A(n10337), .B(n10440), .Z(n10331) );
  XNOR U10571 ( .A(n10335), .B(n10338), .Z(n10440) );
  NAND U10572 ( .A(A[2]), .B(B[235]), .Z(n10338) );
  NANDN U10573 ( .A(n10441), .B(n10442), .Z(n10335) );
  AND U10574 ( .A(A[0]), .B(B[236]), .Z(n10442) );
  XNOR U10575 ( .A(n10340), .B(n10443), .Z(n10337) );
  NAND U10576 ( .A(A[0]), .B(B[237]), .Z(n10443) );
  NAND U10577 ( .A(B[236]), .B(A[1]), .Z(n10340) );
  NAND U10578 ( .A(n10444), .B(n10445), .Z(n265) );
  NANDN U10579 ( .A(n10446), .B(n10447), .Z(n10445) );
  OR U10580 ( .A(n10448), .B(n10449), .Z(n10447) );
  NAND U10581 ( .A(n10449), .B(n10448), .Z(n10444) );
  XOR U10582 ( .A(n267), .B(n266), .Z(\A1[234] ) );
  XOR U10583 ( .A(n10449), .B(n10450), .Z(n266) );
  XNOR U10584 ( .A(n10448), .B(n10446), .Z(n10450) );
  AND U10585 ( .A(n10451), .B(n10452), .Z(n10446) );
  NANDN U10586 ( .A(n10453), .B(n10454), .Z(n10452) );
  NANDN U10587 ( .A(n10455), .B(n10456), .Z(n10454) );
  NANDN U10588 ( .A(n10456), .B(n10455), .Z(n10451) );
  ANDN U10589 ( .B(B[221]), .A(n29), .Z(n10448) );
  XNOR U10590 ( .A(n10355), .B(n10457), .Z(n10449) );
  XNOR U10591 ( .A(n10354), .B(n10352), .Z(n10457) );
  AND U10592 ( .A(n10458), .B(n10459), .Z(n10352) );
  NANDN U10593 ( .A(n10460), .B(n10461), .Z(n10459) );
  OR U10594 ( .A(n10462), .B(n10463), .Z(n10461) );
  NAND U10595 ( .A(n10463), .B(n10462), .Z(n10458) );
  ANDN U10596 ( .B(B[222]), .A(n30), .Z(n10354) );
  XNOR U10597 ( .A(n10362), .B(n10464), .Z(n10355) );
  XNOR U10598 ( .A(n10361), .B(n10359), .Z(n10464) );
  AND U10599 ( .A(n10465), .B(n10466), .Z(n10359) );
  NANDN U10600 ( .A(n10467), .B(n10468), .Z(n10466) );
  NANDN U10601 ( .A(n10469), .B(n10470), .Z(n10468) );
  NANDN U10602 ( .A(n10470), .B(n10469), .Z(n10465) );
  ANDN U10603 ( .B(B[223]), .A(n31), .Z(n10361) );
  XNOR U10604 ( .A(n10369), .B(n10471), .Z(n10362) );
  XNOR U10605 ( .A(n10368), .B(n10366), .Z(n10471) );
  AND U10606 ( .A(n10472), .B(n10473), .Z(n10366) );
  NANDN U10607 ( .A(n10474), .B(n10475), .Z(n10473) );
  OR U10608 ( .A(n10476), .B(n10477), .Z(n10475) );
  NAND U10609 ( .A(n10477), .B(n10476), .Z(n10472) );
  ANDN U10610 ( .B(B[224]), .A(n32), .Z(n10368) );
  XNOR U10611 ( .A(n10376), .B(n10478), .Z(n10369) );
  XNOR U10612 ( .A(n10375), .B(n10373), .Z(n10478) );
  AND U10613 ( .A(n10479), .B(n10480), .Z(n10373) );
  NANDN U10614 ( .A(n10481), .B(n10482), .Z(n10480) );
  NANDN U10615 ( .A(n10483), .B(n10484), .Z(n10482) );
  NANDN U10616 ( .A(n10484), .B(n10483), .Z(n10479) );
  ANDN U10617 ( .B(B[225]), .A(n33), .Z(n10375) );
  XNOR U10618 ( .A(n10383), .B(n10485), .Z(n10376) );
  XNOR U10619 ( .A(n10382), .B(n10380), .Z(n10485) );
  AND U10620 ( .A(n10486), .B(n10487), .Z(n10380) );
  NANDN U10621 ( .A(n10488), .B(n10489), .Z(n10487) );
  OR U10622 ( .A(n10490), .B(n10491), .Z(n10489) );
  NAND U10623 ( .A(n10491), .B(n10490), .Z(n10486) );
  ANDN U10624 ( .B(B[226]), .A(n34), .Z(n10382) );
  XNOR U10625 ( .A(n10390), .B(n10492), .Z(n10383) );
  XNOR U10626 ( .A(n10389), .B(n10387), .Z(n10492) );
  AND U10627 ( .A(n10493), .B(n10494), .Z(n10387) );
  NANDN U10628 ( .A(n10495), .B(n10496), .Z(n10494) );
  NANDN U10629 ( .A(n10497), .B(n10498), .Z(n10496) );
  NANDN U10630 ( .A(n10498), .B(n10497), .Z(n10493) );
  ANDN U10631 ( .B(B[227]), .A(n35), .Z(n10389) );
  XNOR U10632 ( .A(n10397), .B(n10499), .Z(n10390) );
  XNOR U10633 ( .A(n10396), .B(n10394), .Z(n10499) );
  AND U10634 ( .A(n10500), .B(n10501), .Z(n10394) );
  NANDN U10635 ( .A(n10502), .B(n10503), .Z(n10501) );
  OR U10636 ( .A(n10504), .B(n10505), .Z(n10503) );
  NAND U10637 ( .A(n10505), .B(n10504), .Z(n10500) );
  ANDN U10638 ( .B(B[228]), .A(n36), .Z(n10396) );
  XNOR U10639 ( .A(n10404), .B(n10506), .Z(n10397) );
  XNOR U10640 ( .A(n10403), .B(n10401), .Z(n10506) );
  AND U10641 ( .A(n10507), .B(n10508), .Z(n10401) );
  NANDN U10642 ( .A(n10509), .B(n10510), .Z(n10508) );
  NANDN U10643 ( .A(n10511), .B(n10512), .Z(n10510) );
  NANDN U10644 ( .A(n10512), .B(n10511), .Z(n10507) );
  ANDN U10645 ( .B(B[229]), .A(n37), .Z(n10403) );
  XNOR U10646 ( .A(n10411), .B(n10513), .Z(n10404) );
  XNOR U10647 ( .A(n10410), .B(n10408), .Z(n10513) );
  AND U10648 ( .A(n10514), .B(n10515), .Z(n10408) );
  NANDN U10649 ( .A(n10516), .B(n10517), .Z(n10515) );
  OR U10650 ( .A(n10518), .B(n10519), .Z(n10517) );
  NAND U10651 ( .A(n10519), .B(n10518), .Z(n10514) );
  ANDN U10652 ( .B(B[230]), .A(n38), .Z(n10410) );
  XNOR U10653 ( .A(n10418), .B(n10520), .Z(n10411) );
  XNOR U10654 ( .A(n10417), .B(n10415), .Z(n10520) );
  AND U10655 ( .A(n10521), .B(n10522), .Z(n10415) );
  NANDN U10656 ( .A(n10523), .B(n10524), .Z(n10522) );
  NANDN U10657 ( .A(n10525), .B(n10526), .Z(n10524) );
  NANDN U10658 ( .A(n10526), .B(n10525), .Z(n10521) );
  ANDN U10659 ( .B(B[231]), .A(n39), .Z(n10417) );
  XNOR U10660 ( .A(n10425), .B(n10527), .Z(n10418) );
  XNOR U10661 ( .A(n10424), .B(n10422), .Z(n10527) );
  AND U10662 ( .A(n10528), .B(n10529), .Z(n10422) );
  NANDN U10663 ( .A(n10530), .B(n10531), .Z(n10529) );
  OR U10664 ( .A(n10532), .B(n10533), .Z(n10531) );
  NAND U10665 ( .A(n10533), .B(n10532), .Z(n10528) );
  ANDN U10666 ( .B(B[232]), .A(n40), .Z(n10424) );
  XNOR U10667 ( .A(n10432), .B(n10534), .Z(n10425) );
  XNOR U10668 ( .A(n10431), .B(n10429), .Z(n10534) );
  AND U10669 ( .A(n10535), .B(n10536), .Z(n10429) );
  NANDN U10670 ( .A(n10537), .B(n10538), .Z(n10536) );
  NAND U10671 ( .A(n10539), .B(n10540), .Z(n10538) );
  ANDN U10672 ( .B(B[233]), .A(n41), .Z(n10431) );
  XOR U10673 ( .A(n10438), .B(n10541), .Z(n10432) );
  XNOR U10674 ( .A(n10436), .B(n10439), .Z(n10541) );
  NAND U10675 ( .A(A[2]), .B(B[234]), .Z(n10439) );
  NANDN U10676 ( .A(n10542), .B(n10543), .Z(n10436) );
  AND U10677 ( .A(A[0]), .B(B[235]), .Z(n10543) );
  XNOR U10678 ( .A(n10441), .B(n10544), .Z(n10438) );
  NAND U10679 ( .A(A[0]), .B(B[236]), .Z(n10544) );
  NAND U10680 ( .A(B[235]), .B(A[1]), .Z(n10441) );
  NAND U10681 ( .A(n10545), .B(n10546), .Z(n267) );
  NANDN U10682 ( .A(n10547), .B(n10548), .Z(n10546) );
  OR U10683 ( .A(n10549), .B(n10550), .Z(n10548) );
  NAND U10684 ( .A(n10550), .B(n10549), .Z(n10545) );
  XOR U10685 ( .A(n269), .B(n268), .Z(\A1[233] ) );
  XOR U10686 ( .A(n10550), .B(n10551), .Z(n268) );
  XNOR U10687 ( .A(n10549), .B(n10547), .Z(n10551) );
  AND U10688 ( .A(n10552), .B(n10553), .Z(n10547) );
  NANDN U10689 ( .A(n10554), .B(n10555), .Z(n10553) );
  NANDN U10690 ( .A(n10556), .B(n10557), .Z(n10555) );
  NANDN U10691 ( .A(n10557), .B(n10556), .Z(n10552) );
  ANDN U10692 ( .B(B[220]), .A(n29), .Z(n10549) );
  XNOR U10693 ( .A(n10456), .B(n10558), .Z(n10550) );
  XNOR U10694 ( .A(n10455), .B(n10453), .Z(n10558) );
  AND U10695 ( .A(n10559), .B(n10560), .Z(n10453) );
  NANDN U10696 ( .A(n10561), .B(n10562), .Z(n10560) );
  OR U10697 ( .A(n10563), .B(n10564), .Z(n10562) );
  NAND U10698 ( .A(n10564), .B(n10563), .Z(n10559) );
  ANDN U10699 ( .B(B[221]), .A(n30), .Z(n10455) );
  XNOR U10700 ( .A(n10463), .B(n10565), .Z(n10456) );
  XNOR U10701 ( .A(n10462), .B(n10460), .Z(n10565) );
  AND U10702 ( .A(n10566), .B(n10567), .Z(n10460) );
  NANDN U10703 ( .A(n10568), .B(n10569), .Z(n10567) );
  NANDN U10704 ( .A(n10570), .B(n10571), .Z(n10569) );
  NANDN U10705 ( .A(n10571), .B(n10570), .Z(n10566) );
  ANDN U10706 ( .B(B[222]), .A(n31), .Z(n10462) );
  XNOR U10707 ( .A(n10470), .B(n10572), .Z(n10463) );
  XNOR U10708 ( .A(n10469), .B(n10467), .Z(n10572) );
  AND U10709 ( .A(n10573), .B(n10574), .Z(n10467) );
  NANDN U10710 ( .A(n10575), .B(n10576), .Z(n10574) );
  OR U10711 ( .A(n10577), .B(n10578), .Z(n10576) );
  NAND U10712 ( .A(n10578), .B(n10577), .Z(n10573) );
  ANDN U10713 ( .B(B[223]), .A(n32), .Z(n10469) );
  XNOR U10714 ( .A(n10477), .B(n10579), .Z(n10470) );
  XNOR U10715 ( .A(n10476), .B(n10474), .Z(n10579) );
  AND U10716 ( .A(n10580), .B(n10581), .Z(n10474) );
  NANDN U10717 ( .A(n10582), .B(n10583), .Z(n10581) );
  NANDN U10718 ( .A(n10584), .B(n10585), .Z(n10583) );
  NANDN U10719 ( .A(n10585), .B(n10584), .Z(n10580) );
  ANDN U10720 ( .B(B[224]), .A(n33), .Z(n10476) );
  XNOR U10721 ( .A(n10484), .B(n10586), .Z(n10477) );
  XNOR U10722 ( .A(n10483), .B(n10481), .Z(n10586) );
  AND U10723 ( .A(n10587), .B(n10588), .Z(n10481) );
  NANDN U10724 ( .A(n10589), .B(n10590), .Z(n10588) );
  OR U10725 ( .A(n10591), .B(n10592), .Z(n10590) );
  NAND U10726 ( .A(n10592), .B(n10591), .Z(n10587) );
  ANDN U10727 ( .B(B[225]), .A(n34), .Z(n10483) );
  XNOR U10728 ( .A(n10491), .B(n10593), .Z(n10484) );
  XNOR U10729 ( .A(n10490), .B(n10488), .Z(n10593) );
  AND U10730 ( .A(n10594), .B(n10595), .Z(n10488) );
  NANDN U10731 ( .A(n10596), .B(n10597), .Z(n10595) );
  NANDN U10732 ( .A(n10598), .B(n10599), .Z(n10597) );
  NANDN U10733 ( .A(n10599), .B(n10598), .Z(n10594) );
  ANDN U10734 ( .B(B[226]), .A(n35), .Z(n10490) );
  XNOR U10735 ( .A(n10498), .B(n10600), .Z(n10491) );
  XNOR U10736 ( .A(n10497), .B(n10495), .Z(n10600) );
  AND U10737 ( .A(n10601), .B(n10602), .Z(n10495) );
  NANDN U10738 ( .A(n10603), .B(n10604), .Z(n10602) );
  OR U10739 ( .A(n10605), .B(n10606), .Z(n10604) );
  NAND U10740 ( .A(n10606), .B(n10605), .Z(n10601) );
  ANDN U10741 ( .B(B[227]), .A(n36), .Z(n10497) );
  XNOR U10742 ( .A(n10505), .B(n10607), .Z(n10498) );
  XNOR U10743 ( .A(n10504), .B(n10502), .Z(n10607) );
  AND U10744 ( .A(n10608), .B(n10609), .Z(n10502) );
  NANDN U10745 ( .A(n10610), .B(n10611), .Z(n10609) );
  NANDN U10746 ( .A(n10612), .B(n10613), .Z(n10611) );
  NANDN U10747 ( .A(n10613), .B(n10612), .Z(n10608) );
  ANDN U10748 ( .B(B[228]), .A(n37), .Z(n10504) );
  XNOR U10749 ( .A(n10512), .B(n10614), .Z(n10505) );
  XNOR U10750 ( .A(n10511), .B(n10509), .Z(n10614) );
  AND U10751 ( .A(n10615), .B(n10616), .Z(n10509) );
  NANDN U10752 ( .A(n10617), .B(n10618), .Z(n10616) );
  OR U10753 ( .A(n10619), .B(n10620), .Z(n10618) );
  NAND U10754 ( .A(n10620), .B(n10619), .Z(n10615) );
  ANDN U10755 ( .B(B[229]), .A(n38), .Z(n10511) );
  XNOR U10756 ( .A(n10519), .B(n10621), .Z(n10512) );
  XNOR U10757 ( .A(n10518), .B(n10516), .Z(n10621) );
  AND U10758 ( .A(n10622), .B(n10623), .Z(n10516) );
  NANDN U10759 ( .A(n10624), .B(n10625), .Z(n10623) );
  NANDN U10760 ( .A(n10626), .B(n10627), .Z(n10625) );
  NANDN U10761 ( .A(n10627), .B(n10626), .Z(n10622) );
  ANDN U10762 ( .B(B[230]), .A(n39), .Z(n10518) );
  XNOR U10763 ( .A(n10526), .B(n10628), .Z(n10519) );
  XNOR U10764 ( .A(n10525), .B(n10523), .Z(n10628) );
  AND U10765 ( .A(n10629), .B(n10630), .Z(n10523) );
  NANDN U10766 ( .A(n10631), .B(n10632), .Z(n10630) );
  OR U10767 ( .A(n10633), .B(n10634), .Z(n10632) );
  NAND U10768 ( .A(n10634), .B(n10633), .Z(n10629) );
  ANDN U10769 ( .B(B[231]), .A(n40), .Z(n10525) );
  XNOR U10770 ( .A(n10533), .B(n10635), .Z(n10526) );
  XNOR U10771 ( .A(n10532), .B(n10530), .Z(n10635) );
  AND U10772 ( .A(n10636), .B(n10637), .Z(n10530) );
  NANDN U10773 ( .A(n10638), .B(n10639), .Z(n10637) );
  NAND U10774 ( .A(n10640), .B(n10641), .Z(n10639) );
  ANDN U10775 ( .B(B[232]), .A(n41), .Z(n10532) );
  XOR U10776 ( .A(n10539), .B(n10642), .Z(n10533) );
  XNOR U10777 ( .A(n10537), .B(n10540), .Z(n10642) );
  NAND U10778 ( .A(A[2]), .B(B[233]), .Z(n10540) );
  NANDN U10779 ( .A(n10643), .B(n10644), .Z(n10537) );
  AND U10780 ( .A(A[0]), .B(B[234]), .Z(n10644) );
  XNOR U10781 ( .A(n10542), .B(n10645), .Z(n10539) );
  NAND U10782 ( .A(A[0]), .B(B[235]), .Z(n10645) );
  NAND U10783 ( .A(B[234]), .B(A[1]), .Z(n10542) );
  NAND U10784 ( .A(n10646), .B(n10647), .Z(n269) );
  NANDN U10785 ( .A(n10648), .B(n10649), .Z(n10647) );
  OR U10786 ( .A(n10650), .B(n10651), .Z(n10649) );
  NAND U10787 ( .A(n10651), .B(n10650), .Z(n10646) );
  XOR U10788 ( .A(n271), .B(n270), .Z(\A1[232] ) );
  XOR U10789 ( .A(n10651), .B(n10652), .Z(n270) );
  XNOR U10790 ( .A(n10650), .B(n10648), .Z(n10652) );
  AND U10791 ( .A(n10653), .B(n10654), .Z(n10648) );
  NANDN U10792 ( .A(n10655), .B(n10656), .Z(n10654) );
  NANDN U10793 ( .A(n10657), .B(n10658), .Z(n10656) );
  NANDN U10794 ( .A(n10658), .B(n10657), .Z(n10653) );
  ANDN U10795 ( .B(B[219]), .A(n29), .Z(n10650) );
  XNOR U10796 ( .A(n10557), .B(n10659), .Z(n10651) );
  XNOR U10797 ( .A(n10556), .B(n10554), .Z(n10659) );
  AND U10798 ( .A(n10660), .B(n10661), .Z(n10554) );
  NANDN U10799 ( .A(n10662), .B(n10663), .Z(n10661) );
  OR U10800 ( .A(n10664), .B(n10665), .Z(n10663) );
  NAND U10801 ( .A(n10665), .B(n10664), .Z(n10660) );
  ANDN U10802 ( .B(B[220]), .A(n30), .Z(n10556) );
  XNOR U10803 ( .A(n10564), .B(n10666), .Z(n10557) );
  XNOR U10804 ( .A(n10563), .B(n10561), .Z(n10666) );
  AND U10805 ( .A(n10667), .B(n10668), .Z(n10561) );
  NANDN U10806 ( .A(n10669), .B(n10670), .Z(n10668) );
  NANDN U10807 ( .A(n10671), .B(n10672), .Z(n10670) );
  NANDN U10808 ( .A(n10672), .B(n10671), .Z(n10667) );
  ANDN U10809 ( .B(B[221]), .A(n31), .Z(n10563) );
  XNOR U10810 ( .A(n10571), .B(n10673), .Z(n10564) );
  XNOR U10811 ( .A(n10570), .B(n10568), .Z(n10673) );
  AND U10812 ( .A(n10674), .B(n10675), .Z(n10568) );
  NANDN U10813 ( .A(n10676), .B(n10677), .Z(n10675) );
  OR U10814 ( .A(n10678), .B(n10679), .Z(n10677) );
  NAND U10815 ( .A(n10679), .B(n10678), .Z(n10674) );
  ANDN U10816 ( .B(B[222]), .A(n32), .Z(n10570) );
  XNOR U10817 ( .A(n10578), .B(n10680), .Z(n10571) );
  XNOR U10818 ( .A(n10577), .B(n10575), .Z(n10680) );
  AND U10819 ( .A(n10681), .B(n10682), .Z(n10575) );
  NANDN U10820 ( .A(n10683), .B(n10684), .Z(n10682) );
  NANDN U10821 ( .A(n10685), .B(n10686), .Z(n10684) );
  NANDN U10822 ( .A(n10686), .B(n10685), .Z(n10681) );
  ANDN U10823 ( .B(B[223]), .A(n33), .Z(n10577) );
  XNOR U10824 ( .A(n10585), .B(n10687), .Z(n10578) );
  XNOR U10825 ( .A(n10584), .B(n10582), .Z(n10687) );
  AND U10826 ( .A(n10688), .B(n10689), .Z(n10582) );
  NANDN U10827 ( .A(n10690), .B(n10691), .Z(n10689) );
  OR U10828 ( .A(n10692), .B(n10693), .Z(n10691) );
  NAND U10829 ( .A(n10693), .B(n10692), .Z(n10688) );
  ANDN U10830 ( .B(B[224]), .A(n34), .Z(n10584) );
  XNOR U10831 ( .A(n10592), .B(n10694), .Z(n10585) );
  XNOR U10832 ( .A(n10591), .B(n10589), .Z(n10694) );
  AND U10833 ( .A(n10695), .B(n10696), .Z(n10589) );
  NANDN U10834 ( .A(n10697), .B(n10698), .Z(n10696) );
  NANDN U10835 ( .A(n10699), .B(n10700), .Z(n10698) );
  NANDN U10836 ( .A(n10700), .B(n10699), .Z(n10695) );
  ANDN U10837 ( .B(B[225]), .A(n35), .Z(n10591) );
  XNOR U10838 ( .A(n10599), .B(n10701), .Z(n10592) );
  XNOR U10839 ( .A(n10598), .B(n10596), .Z(n10701) );
  AND U10840 ( .A(n10702), .B(n10703), .Z(n10596) );
  NANDN U10841 ( .A(n10704), .B(n10705), .Z(n10703) );
  OR U10842 ( .A(n10706), .B(n10707), .Z(n10705) );
  NAND U10843 ( .A(n10707), .B(n10706), .Z(n10702) );
  ANDN U10844 ( .B(B[226]), .A(n36), .Z(n10598) );
  XNOR U10845 ( .A(n10606), .B(n10708), .Z(n10599) );
  XNOR U10846 ( .A(n10605), .B(n10603), .Z(n10708) );
  AND U10847 ( .A(n10709), .B(n10710), .Z(n10603) );
  NANDN U10848 ( .A(n10711), .B(n10712), .Z(n10710) );
  NANDN U10849 ( .A(n10713), .B(n10714), .Z(n10712) );
  NANDN U10850 ( .A(n10714), .B(n10713), .Z(n10709) );
  ANDN U10851 ( .B(B[227]), .A(n37), .Z(n10605) );
  XNOR U10852 ( .A(n10613), .B(n10715), .Z(n10606) );
  XNOR U10853 ( .A(n10612), .B(n10610), .Z(n10715) );
  AND U10854 ( .A(n10716), .B(n10717), .Z(n10610) );
  NANDN U10855 ( .A(n10718), .B(n10719), .Z(n10717) );
  OR U10856 ( .A(n10720), .B(n10721), .Z(n10719) );
  NAND U10857 ( .A(n10721), .B(n10720), .Z(n10716) );
  ANDN U10858 ( .B(B[228]), .A(n38), .Z(n10612) );
  XNOR U10859 ( .A(n10620), .B(n10722), .Z(n10613) );
  XNOR U10860 ( .A(n10619), .B(n10617), .Z(n10722) );
  AND U10861 ( .A(n10723), .B(n10724), .Z(n10617) );
  NANDN U10862 ( .A(n10725), .B(n10726), .Z(n10724) );
  NANDN U10863 ( .A(n10727), .B(n10728), .Z(n10726) );
  NANDN U10864 ( .A(n10728), .B(n10727), .Z(n10723) );
  ANDN U10865 ( .B(B[229]), .A(n39), .Z(n10619) );
  XNOR U10866 ( .A(n10627), .B(n10729), .Z(n10620) );
  XNOR U10867 ( .A(n10626), .B(n10624), .Z(n10729) );
  AND U10868 ( .A(n10730), .B(n10731), .Z(n10624) );
  NANDN U10869 ( .A(n10732), .B(n10733), .Z(n10731) );
  OR U10870 ( .A(n10734), .B(n10735), .Z(n10733) );
  NAND U10871 ( .A(n10735), .B(n10734), .Z(n10730) );
  ANDN U10872 ( .B(B[230]), .A(n40), .Z(n10626) );
  XNOR U10873 ( .A(n10634), .B(n10736), .Z(n10627) );
  XNOR U10874 ( .A(n10633), .B(n10631), .Z(n10736) );
  AND U10875 ( .A(n10737), .B(n10738), .Z(n10631) );
  NANDN U10876 ( .A(n10739), .B(n10740), .Z(n10738) );
  NAND U10877 ( .A(n10741), .B(n10742), .Z(n10740) );
  ANDN U10878 ( .B(B[231]), .A(n41), .Z(n10633) );
  XOR U10879 ( .A(n10640), .B(n10743), .Z(n10634) );
  XNOR U10880 ( .A(n10638), .B(n10641), .Z(n10743) );
  NAND U10881 ( .A(A[2]), .B(B[232]), .Z(n10641) );
  NANDN U10882 ( .A(n10744), .B(n10745), .Z(n10638) );
  AND U10883 ( .A(A[0]), .B(B[233]), .Z(n10745) );
  XNOR U10884 ( .A(n10643), .B(n10746), .Z(n10640) );
  NAND U10885 ( .A(A[0]), .B(B[234]), .Z(n10746) );
  NAND U10886 ( .A(B[233]), .B(A[1]), .Z(n10643) );
  NAND U10887 ( .A(n10747), .B(n10748), .Z(n271) );
  NANDN U10888 ( .A(n10749), .B(n10750), .Z(n10748) );
  OR U10889 ( .A(n10751), .B(n10752), .Z(n10750) );
  NAND U10890 ( .A(n10752), .B(n10751), .Z(n10747) );
  XOR U10891 ( .A(n273), .B(n272), .Z(\A1[231] ) );
  XOR U10892 ( .A(n10752), .B(n10753), .Z(n272) );
  XNOR U10893 ( .A(n10751), .B(n10749), .Z(n10753) );
  AND U10894 ( .A(n10754), .B(n10755), .Z(n10749) );
  NANDN U10895 ( .A(n10756), .B(n10757), .Z(n10755) );
  NANDN U10896 ( .A(n10758), .B(n10759), .Z(n10757) );
  NANDN U10897 ( .A(n10759), .B(n10758), .Z(n10754) );
  ANDN U10898 ( .B(B[218]), .A(n29), .Z(n10751) );
  XNOR U10899 ( .A(n10658), .B(n10760), .Z(n10752) );
  XNOR U10900 ( .A(n10657), .B(n10655), .Z(n10760) );
  AND U10901 ( .A(n10761), .B(n10762), .Z(n10655) );
  NANDN U10902 ( .A(n10763), .B(n10764), .Z(n10762) );
  OR U10903 ( .A(n10765), .B(n10766), .Z(n10764) );
  NAND U10904 ( .A(n10766), .B(n10765), .Z(n10761) );
  ANDN U10905 ( .B(B[219]), .A(n30), .Z(n10657) );
  XNOR U10906 ( .A(n10665), .B(n10767), .Z(n10658) );
  XNOR U10907 ( .A(n10664), .B(n10662), .Z(n10767) );
  AND U10908 ( .A(n10768), .B(n10769), .Z(n10662) );
  NANDN U10909 ( .A(n10770), .B(n10771), .Z(n10769) );
  NANDN U10910 ( .A(n10772), .B(n10773), .Z(n10771) );
  NANDN U10911 ( .A(n10773), .B(n10772), .Z(n10768) );
  ANDN U10912 ( .B(B[220]), .A(n31), .Z(n10664) );
  XNOR U10913 ( .A(n10672), .B(n10774), .Z(n10665) );
  XNOR U10914 ( .A(n10671), .B(n10669), .Z(n10774) );
  AND U10915 ( .A(n10775), .B(n10776), .Z(n10669) );
  NANDN U10916 ( .A(n10777), .B(n10778), .Z(n10776) );
  OR U10917 ( .A(n10779), .B(n10780), .Z(n10778) );
  NAND U10918 ( .A(n10780), .B(n10779), .Z(n10775) );
  ANDN U10919 ( .B(B[221]), .A(n32), .Z(n10671) );
  XNOR U10920 ( .A(n10679), .B(n10781), .Z(n10672) );
  XNOR U10921 ( .A(n10678), .B(n10676), .Z(n10781) );
  AND U10922 ( .A(n10782), .B(n10783), .Z(n10676) );
  NANDN U10923 ( .A(n10784), .B(n10785), .Z(n10783) );
  NANDN U10924 ( .A(n10786), .B(n10787), .Z(n10785) );
  NANDN U10925 ( .A(n10787), .B(n10786), .Z(n10782) );
  ANDN U10926 ( .B(B[222]), .A(n33), .Z(n10678) );
  XNOR U10927 ( .A(n10686), .B(n10788), .Z(n10679) );
  XNOR U10928 ( .A(n10685), .B(n10683), .Z(n10788) );
  AND U10929 ( .A(n10789), .B(n10790), .Z(n10683) );
  NANDN U10930 ( .A(n10791), .B(n10792), .Z(n10790) );
  OR U10931 ( .A(n10793), .B(n10794), .Z(n10792) );
  NAND U10932 ( .A(n10794), .B(n10793), .Z(n10789) );
  ANDN U10933 ( .B(B[223]), .A(n34), .Z(n10685) );
  XNOR U10934 ( .A(n10693), .B(n10795), .Z(n10686) );
  XNOR U10935 ( .A(n10692), .B(n10690), .Z(n10795) );
  AND U10936 ( .A(n10796), .B(n10797), .Z(n10690) );
  NANDN U10937 ( .A(n10798), .B(n10799), .Z(n10797) );
  NANDN U10938 ( .A(n10800), .B(n10801), .Z(n10799) );
  NANDN U10939 ( .A(n10801), .B(n10800), .Z(n10796) );
  ANDN U10940 ( .B(B[224]), .A(n35), .Z(n10692) );
  XNOR U10941 ( .A(n10700), .B(n10802), .Z(n10693) );
  XNOR U10942 ( .A(n10699), .B(n10697), .Z(n10802) );
  AND U10943 ( .A(n10803), .B(n10804), .Z(n10697) );
  NANDN U10944 ( .A(n10805), .B(n10806), .Z(n10804) );
  OR U10945 ( .A(n10807), .B(n10808), .Z(n10806) );
  NAND U10946 ( .A(n10808), .B(n10807), .Z(n10803) );
  ANDN U10947 ( .B(B[225]), .A(n36), .Z(n10699) );
  XNOR U10948 ( .A(n10707), .B(n10809), .Z(n10700) );
  XNOR U10949 ( .A(n10706), .B(n10704), .Z(n10809) );
  AND U10950 ( .A(n10810), .B(n10811), .Z(n10704) );
  NANDN U10951 ( .A(n10812), .B(n10813), .Z(n10811) );
  NANDN U10952 ( .A(n10814), .B(n10815), .Z(n10813) );
  NANDN U10953 ( .A(n10815), .B(n10814), .Z(n10810) );
  ANDN U10954 ( .B(B[226]), .A(n37), .Z(n10706) );
  XNOR U10955 ( .A(n10714), .B(n10816), .Z(n10707) );
  XNOR U10956 ( .A(n10713), .B(n10711), .Z(n10816) );
  AND U10957 ( .A(n10817), .B(n10818), .Z(n10711) );
  NANDN U10958 ( .A(n10819), .B(n10820), .Z(n10818) );
  OR U10959 ( .A(n10821), .B(n10822), .Z(n10820) );
  NAND U10960 ( .A(n10822), .B(n10821), .Z(n10817) );
  ANDN U10961 ( .B(B[227]), .A(n38), .Z(n10713) );
  XNOR U10962 ( .A(n10721), .B(n10823), .Z(n10714) );
  XNOR U10963 ( .A(n10720), .B(n10718), .Z(n10823) );
  AND U10964 ( .A(n10824), .B(n10825), .Z(n10718) );
  NANDN U10965 ( .A(n10826), .B(n10827), .Z(n10825) );
  NANDN U10966 ( .A(n10828), .B(n10829), .Z(n10827) );
  NANDN U10967 ( .A(n10829), .B(n10828), .Z(n10824) );
  ANDN U10968 ( .B(B[228]), .A(n39), .Z(n10720) );
  XNOR U10969 ( .A(n10728), .B(n10830), .Z(n10721) );
  XNOR U10970 ( .A(n10727), .B(n10725), .Z(n10830) );
  AND U10971 ( .A(n10831), .B(n10832), .Z(n10725) );
  NANDN U10972 ( .A(n10833), .B(n10834), .Z(n10832) );
  OR U10973 ( .A(n10835), .B(n10836), .Z(n10834) );
  NAND U10974 ( .A(n10836), .B(n10835), .Z(n10831) );
  ANDN U10975 ( .B(B[229]), .A(n40), .Z(n10727) );
  XNOR U10976 ( .A(n10735), .B(n10837), .Z(n10728) );
  XNOR U10977 ( .A(n10734), .B(n10732), .Z(n10837) );
  AND U10978 ( .A(n10838), .B(n10839), .Z(n10732) );
  NANDN U10979 ( .A(n10840), .B(n10841), .Z(n10839) );
  NAND U10980 ( .A(n10842), .B(n10843), .Z(n10841) );
  ANDN U10981 ( .B(B[230]), .A(n41), .Z(n10734) );
  XOR U10982 ( .A(n10741), .B(n10844), .Z(n10735) );
  XNOR U10983 ( .A(n10739), .B(n10742), .Z(n10844) );
  NAND U10984 ( .A(A[2]), .B(B[231]), .Z(n10742) );
  NANDN U10985 ( .A(n10845), .B(n10846), .Z(n10739) );
  AND U10986 ( .A(A[0]), .B(B[232]), .Z(n10846) );
  XNOR U10987 ( .A(n10744), .B(n10847), .Z(n10741) );
  NAND U10988 ( .A(A[0]), .B(B[233]), .Z(n10847) );
  NAND U10989 ( .A(B[232]), .B(A[1]), .Z(n10744) );
  NAND U10990 ( .A(n10848), .B(n10849), .Z(n273) );
  NANDN U10991 ( .A(n10850), .B(n10851), .Z(n10849) );
  OR U10992 ( .A(n10852), .B(n10853), .Z(n10851) );
  NAND U10993 ( .A(n10853), .B(n10852), .Z(n10848) );
  XOR U10994 ( .A(n275), .B(n274), .Z(\A1[230] ) );
  XOR U10995 ( .A(n10853), .B(n10854), .Z(n274) );
  XNOR U10996 ( .A(n10852), .B(n10850), .Z(n10854) );
  AND U10997 ( .A(n10855), .B(n10856), .Z(n10850) );
  NANDN U10998 ( .A(n10857), .B(n10858), .Z(n10856) );
  NANDN U10999 ( .A(n10859), .B(n10860), .Z(n10858) );
  NANDN U11000 ( .A(n10860), .B(n10859), .Z(n10855) );
  ANDN U11001 ( .B(B[217]), .A(n29), .Z(n10852) );
  XNOR U11002 ( .A(n10759), .B(n10861), .Z(n10853) );
  XNOR U11003 ( .A(n10758), .B(n10756), .Z(n10861) );
  AND U11004 ( .A(n10862), .B(n10863), .Z(n10756) );
  NANDN U11005 ( .A(n10864), .B(n10865), .Z(n10863) );
  OR U11006 ( .A(n10866), .B(n10867), .Z(n10865) );
  NAND U11007 ( .A(n10867), .B(n10866), .Z(n10862) );
  ANDN U11008 ( .B(B[218]), .A(n30), .Z(n10758) );
  XNOR U11009 ( .A(n10766), .B(n10868), .Z(n10759) );
  XNOR U11010 ( .A(n10765), .B(n10763), .Z(n10868) );
  AND U11011 ( .A(n10869), .B(n10870), .Z(n10763) );
  NANDN U11012 ( .A(n10871), .B(n10872), .Z(n10870) );
  NANDN U11013 ( .A(n10873), .B(n10874), .Z(n10872) );
  NANDN U11014 ( .A(n10874), .B(n10873), .Z(n10869) );
  ANDN U11015 ( .B(B[219]), .A(n31), .Z(n10765) );
  XNOR U11016 ( .A(n10773), .B(n10875), .Z(n10766) );
  XNOR U11017 ( .A(n10772), .B(n10770), .Z(n10875) );
  AND U11018 ( .A(n10876), .B(n10877), .Z(n10770) );
  NANDN U11019 ( .A(n10878), .B(n10879), .Z(n10877) );
  OR U11020 ( .A(n10880), .B(n10881), .Z(n10879) );
  NAND U11021 ( .A(n10881), .B(n10880), .Z(n10876) );
  ANDN U11022 ( .B(B[220]), .A(n32), .Z(n10772) );
  XNOR U11023 ( .A(n10780), .B(n10882), .Z(n10773) );
  XNOR U11024 ( .A(n10779), .B(n10777), .Z(n10882) );
  AND U11025 ( .A(n10883), .B(n10884), .Z(n10777) );
  NANDN U11026 ( .A(n10885), .B(n10886), .Z(n10884) );
  NANDN U11027 ( .A(n10887), .B(n10888), .Z(n10886) );
  NANDN U11028 ( .A(n10888), .B(n10887), .Z(n10883) );
  ANDN U11029 ( .B(B[221]), .A(n33), .Z(n10779) );
  XNOR U11030 ( .A(n10787), .B(n10889), .Z(n10780) );
  XNOR U11031 ( .A(n10786), .B(n10784), .Z(n10889) );
  AND U11032 ( .A(n10890), .B(n10891), .Z(n10784) );
  NANDN U11033 ( .A(n10892), .B(n10893), .Z(n10891) );
  OR U11034 ( .A(n10894), .B(n10895), .Z(n10893) );
  NAND U11035 ( .A(n10895), .B(n10894), .Z(n10890) );
  ANDN U11036 ( .B(B[222]), .A(n34), .Z(n10786) );
  XNOR U11037 ( .A(n10794), .B(n10896), .Z(n10787) );
  XNOR U11038 ( .A(n10793), .B(n10791), .Z(n10896) );
  AND U11039 ( .A(n10897), .B(n10898), .Z(n10791) );
  NANDN U11040 ( .A(n10899), .B(n10900), .Z(n10898) );
  NANDN U11041 ( .A(n10901), .B(n10902), .Z(n10900) );
  NANDN U11042 ( .A(n10902), .B(n10901), .Z(n10897) );
  ANDN U11043 ( .B(B[223]), .A(n35), .Z(n10793) );
  XNOR U11044 ( .A(n10801), .B(n10903), .Z(n10794) );
  XNOR U11045 ( .A(n10800), .B(n10798), .Z(n10903) );
  AND U11046 ( .A(n10904), .B(n10905), .Z(n10798) );
  NANDN U11047 ( .A(n10906), .B(n10907), .Z(n10905) );
  OR U11048 ( .A(n10908), .B(n10909), .Z(n10907) );
  NAND U11049 ( .A(n10909), .B(n10908), .Z(n10904) );
  ANDN U11050 ( .B(B[224]), .A(n36), .Z(n10800) );
  XNOR U11051 ( .A(n10808), .B(n10910), .Z(n10801) );
  XNOR U11052 ( .A(n10807), .B(n10805), .Z(n10910) );
  AND U11053 ( .A(n10911), .B(n10912), .Z(n10805) );
  NANDN U11054 ( .A(n10913), .B(n10914), .Z(n10912) );
  NANDN U11055 ( .A(n10915), .B(n10916), .Z(n10914) );
  NANDN U11056 ( .A(n10916), .B(n10915), .Z(n10911) );
  ANDN U11057 ( .B(B[225]), .A(n37), .Z(n10807) );
  XNOR U11058 ( .A(n10815), .B(n10917), .Z(n10808) );
  XNOR U11059 ( .A(n10814), .B(n10812), .Z(n10917) );
  AND U11060 ( .A(n10918), .B(n10919), .Z(n10812) );
  NANDN U11061 ( .A(n10920), .B(n10921), .Z(n10919) );
  OR U11062 ( .A(n10922), .B(n10923), .Z(n10921) );
  NAND U11063 ( .A(n10923), .B(n10922), .Z(n10918) );
  ANDN U11064 ( .B(B[226]), .A(n38), .Z(n10814) );
  XNOR U11065 ( .A(n10822), .B(n10924), .Z(n10815) );
  XNOR U11066 ( .A(n10821), .B(n10819), .Z(n10924) );
  AND U11067 ( .A(n10925), .B(n10926), .Z(n10819) );
  NANDN U11068 ( .A(n10927), .B(n10928), .Z(n10926) );
  NANDN U11069 ( .A(n10929), .B(n10930), .Z(n10928) );
  NANDN U11070 ( .A(n10930), .B(n10929), .Z(n10925) );
  ANDN U11071 ( .B(B[227]), .A(n39), .Z(n10821) );
  XNOR U11072 ( .A(n10829), .B(n10931), .Z(n10822) );
  XNOR U11073 ( .A(n10828), .B(n10826), .Z(n10931) );
  AND U11074 ( .A(n10932), .B(n10933), .Z(n10826) );
  NANDN U11075 ( .A(n10934), .B(n10935), .Z(n10933) );
  OR U11076 ( .A(n10936), .B(n10937), .Z(n10935) );
  NAND U11077 ( .A(n10937), .B(n10936), .Z(n10932) );
  ANDN U11078 ( .B(B[228]), .A(n40), .Z(n10828) );
  XNOR U11079 ( .A(n10836), .B(n10938), .Z(n10829) );
  XNOR U11080 ( .A(n10835), .B(n10833), .Z(n10938) );
  AND U11081 ( .A(n10939), .B(n10940), .Z(n10833) );
  NANDN U11082 ( .A(n10941), .B(n10942), .Z(n10940) );
  NAND U11083 ( .A(n10943), .B(n10944), .Z(n10942) );
  ANDN U11084 ( .B(B[229]), .A(n41), .Z(n10835) );
  XOR U11085 ( .A(n10842), .B(n10945), .Z(n10836) );
  XNOR U11086 ( .A(n10840), .B(n10843), .Z(n10945) );
  NAND U11087 ( .A(A[2]), .B(B[230]), .Z(n10843) );
  NANDN U11088 ( .A(n10946), .B(n10947), .Z(n10840) );
  AND U11089 ( .A(A[0]), .B(B[231]), .Z(n10947) );
  XNOR U11090 ( .A(n10845), .B(n10948), .Z(n10842) );
  NAND U11091 ( .A(A[0]), .B(B[232]), .Z(n10948) );
  NAND U11092 ( .A(B[231]), .B(A[1]), .Z(n10845) );
  NAND U11093 ( .A(n10949), .B(n10950), .Z(n275) );
  NANDN U11094 ( .A(n10951), .B(n10952), .Z(n10950) );
  OR U11095 ( .A(n10953), .B(n10954), .Z(n10952) );
  NAND U11096 ( .A(n10954), .B(n10953), .Z(n10949) );
  XOR U11097 ( .A(n257), .B(n256), .Z(\A1[22] ) );
  XOR U11098 ( .A(n9944), .B(n10955), .Z(n256) );
  XNOR U11099 ( .A(n9943), .B(n9941), .Z(n10955) );
  AND U11100 ( .A(n10956), .B(n10957), .Z(n9941) );
  NANDN U11101 ( .A(n10958), .B(n10959), .Z(n10957) );
  NANDN U11102 ( .A(n10960), .B(n10961), .Z(n10959) );
  NANDN U11103 ( .A(n10961), .B(n10960), .Z(n10956) );
  ANDN U11104 ( .B(B[9]), .A(n29), .Z(n9943) );
  XNOR U11105 ( .A(n9850), .B(n10962), .Z(n9944) );
  XNOR U11106 ( .A(n9849), .B(n9847), .Z(n10962) );
  AND U11107 ( .A(n10963), .B(n10964), .Z(n9847) );
  NANDN U11108 ( .A(n10965), .B(n10966), .Z(n10964) );
  OR U11109 ( .A(n10967), .B(n10968), .Z(n10966) );
  NAND U11110 ( .A(n10968), .B(n10967), .Z(n10963) );
  ANDN U11111 ( .B(B[10]), .A(n30), .Z(n9849) );
  XNOR U11112 ( .A(n9857), .B(n10969), .Z(n9850) );
  XNOR U11113 ( .A(n9856), .B(n9854), .Z(n10969) );
  AND U11114 ( .A(n10970), .B(n10971), .Z(n9854) );
  NANDN U11115 ( .A(n10972), .B(n10973), .Z(n10971) );
  NANDN U11116 ( .A(n10974), .B(n10975), .Z(n10973) );
  NANDN U11117 ( .A(n10975), .B(n10974), .Z(n10970) );
  ANDN U11118 ( .B(B[11]), .A(n31), .Z(n9856) );
  XNOR U11119 ( .A(n9864), .B(n10976), .Z(n9857) );
  XNOR U11120 ( .A(n9863), .B(n9861), .Z(n10976) );
  AND U11121 ( .A(n10977), .B(n10978), .Z(n9861) );
  NANDN U11122 ( .A(n10979), .B(n10980), .Z(n10978) );
  OR U11123 ( .A(n10981), .B(n10982), .Z(n10980) );
  NAND U11124 ( .A(n10982), .B(n10981), .Z(n10977) );
  ANDN U11125 ( .B(B[12]), .A(n32), .Z(n9863) );
  XNOR U11126 ( .A(n9871), .B(n10983), .Z(n9864) );
  XNOR U11127 ( .A(n9870), .B(n9868), .Z(n10983) );
  AND U11128 ( .A(n10984), .B(n10985), .Z(n9868) );
  NANDN U11129 ( .A(n10986), .B(n10987), .Z(n10985) );
  NANDN U11130 ( .A(n10988), .B(n10989), .Z(n10987) );
  NANDN U11131 ( .A(n10989), .B(n10988), .Z(n10984) );
  ANDN U11132 ( .B(B[13]), .A(n33), .Z(n9870) );
  XNOR U11133 ( .A(n9878), .B(n10990), .Z(n9871) );
  XNOR U11134 ( .A(n9877), .B(n9875), .Z(n10990) );
  AND U11135 ( .A(n10991), .B(n10992), .Z(n9875) );
  NANDN U11136 ( .A(n10993), .B(n10994), .Z(n10992) );
  OR U11137 ( .A(n10995), .B(n10996), .Z(n10994) );
  NAND U11138 ( .A(n10996), .B(n10995), .Z(n10991) );
  ANDN U11139 ( .B(B[14]), .A(n34), .Z(n9877) );
  XNOR U11140 ( .A(n9885), .B(n10997), .Z(n9878) );
  XNOR U11141 ( .A(n9884), .B(n9882), .Z(n10997) );
  AND U11142 ( .A(n10998), .B(n10999), .Z(n9882) );
  NANDN U11143 ( .A(n11000), .B(n11001), .Z(n10999) );
  NANDN U11144 ( .A(n11002), .B(n11003), .Z(n11001) );
  NANDN U11145 ( .A(n11003), .B(n11002), .Z(n10998) );
  ANDN U11146 ( .B(B[15]), .A(n35), .Z(n9884) );
  XNOR U11147 ( .A(n9892), .B(n11004), .Z(n9885) );
  XNOR U11148 ( .A(n9891), .B(n9889), .Z(n11004) );
  AND U11149 ( .A(n11005), .B(n11006), .Z(n9889) );
  NANDN U11150 ( .A(n11007), .B(n11008), .Z(n11006) );
  OR U11151 ( .A(n11009), .B(n11010), .Z(n11008) );
  NAND U11152 ( .A(n11010), .B(n11009), .Z(n11005) );
  ANDN U11153 ( .B(B[16]), .A(n36), .Z(n9891) );
  XNOR U11154 ( .A(n9899), .B(n11011), .Z(n9892) );
  XNOR U11155 ( .A(n9898), .B(n9896), .Z(n11011) );
  AND U11156 ( .A(n11012), .B(n11013), .Z(n9896) );
  NANDN U11157 ( .A(n11014), .B(n11015), .Z(n11013) );
  NANDN U11158 ( .A(n11016), .B(n11017), .Z(n11015) );
  NANDN U11159 ( .A(n11017), .B(n11016), .Z(n11012) );
  ANDN U11160 ( .B(B[17]), .A(n37), .Z(n9898) );
  XNOR U11161 ( .A(n9906), .B(n11018), .Z(n9899) );
  XNOR U11162 ( .A(n9905), .B(n9903), .Z(n11018) );
  AND U11163 ( .A(n11019), .B(n11020), .Z(n9903) );
  NANDN U11164 ( .A(n11021), .B(n11022), .Z(n11020) );
  OR U11165 ( .A(n11023), .B(n11024), .Z(n11022) );
  NAND U11166 ( .A(n11024), .B(n11023), .Z(n11019) );
  ANDN U11167 ( .B(B[18]), .A(n38), .Z(n9905) );
  XNOR U11168 ( .A(n9913), .B(n11025), .Z(n9906) );
  XNOR U11169 ( .A(n9912), .B(n9910), .Z(n11025) );
  AND U11170 ( .A(n11026), .B(n11027), .Z(n9910) );
  NANDN U11171 ( .A(n11028), .B(n11029), .Z(n11027) );
  NANDN U11172 ( .A(n11030), .B(n11031), .Z(n11029) );
  NANDN U11173 ( .A(n11031), .B(n11030), .Z(n11026) );
  ANDN U11174 ( .B(B[19]), .A(n39), .Z(n9912) );
  XNOR U11175 ( .A(n9920), .B(n11032), .Z(n9913) );
  XNOR U11176 ( .A(n9919), .B(n9917), .Z(n11032) );
  AND U11177 ( .A(n11033), .B(n11034), .Z(n9917) );
  NANDN U11178 ( .A(n11035), .B(n11036), .Z(n11034) );
  OR U11179 ( .A(n11037), .B(n11038), .Z(n11036) );
  NAND U11180 ( .A(n11038), .B(n11037), .Z(n11033) );
  ANDN U11181 ( .B(B[20]), .A(n40), .Z(n9919) );
  XNOR U11182 ( .A(n9927), .B(n11039), .Z(n9920) );
  XNOR U11183 ( .A(n9926), .B(n9924), .Z(n11039) );
  AND U11184 ( .A(n11040), .B(n11041), .Z(n9924) );
  NANDN U11185 ( .A(n11042), .B(n11043), .Z(n11041) );
  NAND U11186 ( .A(n11044), .B(n11045), .Z(n11043) );
  ANDN U11187 ( .B(B[21]), .A(n41), .Z(n9926) );
  XOR U11188 ( .A(n9933), .B(n11046), .Z(n9927) );
  XNOR U11189 ( .A(n9931), .B(n9934), .Z(n11046) );
  NAND U11190 ( .A(A[2]), .B(B[22]), .Z(n9934) );
  NANDN U11191 ( .A(n11047), .B(n11048), .Z(n9931) );
  AND U11192 ( .A(A[0]), .B(B[23]), .Z(n11048) );
  XNOR U11193 ( .A(n9936), .B(n11049), .Z(n9933) );
  NAND U11194 ( .A(A[0]), .B(B[24]), .Z(n11049) );
  NAND U11195 ( .A(B[23]), .B(A[1]), .Z(n9936) );
  NAND U11196 ( .A(n11050), .B(n11051), .Z(n257) );
  NANDN U11197 ( .A(n11052), .B(n11053), .Z(n11051) );
  OR U11198 ( .A(n11054), .B(n11055), .Z(n11053) );
  NAND U11199 ( .A(n11055), .B(n11054), .Z(n11050) );
  XOR U11200 ( .A(n277), .B(n276), .Z(\A1[229] ) );
  XOR U11201 ( .A(n10954), .B(n11056), .Z(n276) );
  XNOR U11202 ( .A(n10953), .B(n10951), .Z(n11056) );
  AND U11203 ( .A(n11057), .B(n11058), .Z(n10951) );
  NANDN U11204 ( .A(n11059), .B(n11060), .Z(n11058) );
  NANDN U11205 ( .A(n11061), .B(n11062), .Z(n11060) );
  NANDN U11206 ( .A(n11062), .B(n11061), .Z(n11057) );
  ANDN U11207 ( .B(B[216]), .A(n29), .Z(n10953) );
  XNOR U11208 ( .A(n10860), .B(n11063), .Z(n10954) );
  XNOR U11209 ( .A(n10859), .B(n10857), .Z(n11063) );
  AND U11210 ( .A(n11064), .B(n11065), .Z(n10857) );
  NANDN U11211 ( .A(n11066), .B(n11067), .Z(n11065) );
  OR U11212 ( .A(n11068), .B(n11069), .Z(n11067) );
  NAND U11213 ( .A(n11069), .B(n11068), .Z(n11064) );
  ANDN U11214 ( .B(B[217]), .A(n30), .Z(n10859) );
  XNOR U11215 ( .A(n10867), .B(n11070), .Z(n10860) );
  XNOR U11216 ( .A(n10866), .B(n10864), .Z(n11070) );
  AND U11217 ( .A(n11071), .B(n11072), .Z(n10864) );
  NANDN U11218 ( .A(n11073), .B(n11074), .Z(n11072) );
  NANDN U11219 ( .A(n11075), .B(n11076), .Z(n11074) );
  NANDN U11220 ( .A(n11076), .B(n11075), .Z(n11071) );
  ANDN U11221 ( .B(B[218]), .A(n31), .Z(n10866) );
  XNOR U11222 ( .A(n10874), .B(n11077), .Z(n10867) );
  XNOR U11223 ( .A(n10873), .B(n10871), .Z(n11077) );
  AND U11224 ( .A(n11078), .B(n11079), .Z(n10871) );
  NANDN U11225 ( .A(n11080), .B(n11081), .Z(n11079) );
  OR U11226 ( .A(n11082), .B(n11083), .Z(n11081) );
  NAND U11227 ( .A(n11083), .B(n11082), .Z(n11078) );
  ANDN U11228 ( .B(B[219]), .A(n32), .Z(n10873) );
  XNOR U11229 ( .A(n10881), .B(n11084), .Z(n10874) );
  XNOR U11230 ( .A(n10880), .B(n10878), .Z(n11084) );
  AND U11231 ( .A(n11085), .B(n11086), .Z(n10878) );
  NANDN U11232 ( .A(n11087), .B(n11088), .Z(n11086) );
  NANDN U11233 ( .A(n11089), .B(n11090), .Z(n11088) );
  NANDN U11234 ( .A(n11090), .B(n11089), .Z(n11085) );
  ANDN U11235 ( .B(B[220]), .A(n33), .Z(n10880) );
  XNOR U11236 ( .A(n10888), .B(n11091), .Z(n10881) );
  XNOR U11237 ( .A(n10887), .B(n10885), .Z(n11091) );
  AND U11238 ( .A(n11092), .B(n11093), .Z(n10885) );
  NANDN U11239 ( .A(n11094), .B(n11095), .Z(n11093) );
  OR U11240 ( .A(n11096), .B(n11097), .Z(n11095) );
  NAND U11241 ( .A(n11097), .B(n11096), .Z(n11092) );
  ANDN U11242 ( .B(B[221]), .A(n34), .Z(n10887) );
  XNOR U11243 ( .A(n10895), .B(n11098), .Z(n10888) );
  XNOR U11244 ( .A(n10894), .B(n10892), .Z(n11098) );
  AND U11245 ( .A(n11099), .B(n11100), .Z(n10892) );
  NANDN U11246 ( .A(n11101), .B(n11102), .Z(n11100) );
  NANDN U11247 ( .A(n11103), .B(n11104), .Z(n11102) );
  NANDN U11248 ( .A(n11104), .B(n11103), .Z(n11099) );
  ANDN U11249 ( .B(B[222]), .A(n35), .Z(n10894) );
  XNOR U11250 ( .A(n10902), .B(n11105), .Z(n10895) );
  XNOR U11251 ( .A(n10901), .B(n10899), .Z(n11105) );
  AND U11252 ( .A(n11106), .B(n11107), .Z(n10899) );
  NANDN U11253 ( .A(n11108), .B(n11109), .Z(n11107) );
  OR U11254 ( .A(n11110), .B(n11111), .Z(n11109) );
  NAND U11255 ( .A(n11111), .B(n11110), .Z(n11106) );
  ANDN U11256 ( .B(B[223]), .A(n36), .Z(n10901) );
  XNOR U11257 ( .A(n10909), .B(n11112), .Z(n10902) );
  XNOR U11258 ( .A(n10908), .B(n10906), .Z(n11112) );
  AND U11259 ( .A(n11113), .B(n11114), .Z(n10906) );
  NANDN U11260 ( .A(n11115), .B(n11116), .Z(n11114) );
  NANDN U11261 ( .A(n11117), .B(n11118), .Z(n11116) );
  NANDN U11262 ( .A(n11118), .B(n11117), .Z(n11113) );
  ANDN U11263 ( .B(B[224]), .A(n37), .Z(n10908) );
  XNOR U11264 ( .A(n10916), .B(n11119), .Z(n10909) );
  XNOR U11265 ( .A(n10915), .B(n10913), .Z(n11119) );
  AND U11266 ( .A(n11120), .B(n11121), .Z(n10913) );
  NANDN U11267 ( .A(n11122), .B(n11123), .Z(n11121) );
  OR U11268 ( .A(n11124), .B(n11125), .Z(n11123) );
  NAND U11269 ( .A(n11125), .B(n11124), .Z(n11120) );
  ANDN U11270 ( .B(B[225]), .A(n38), .Z(n10915) );
  XNOR U11271 ( .A(n10923), .B(n11126), .Z(n10916) );
  XNOR U11272 ( .A(n10922), .B(n10920), .Z(n11126) );
  AND U11273 ( .A(n11127), .B(n11128), .Z(n10920) );
  NANDN U11274 ( .A(n11129), .B(n11130), .Z(n11128) );
  NANDN U11275 ( .A(n11131), .B(n11132), .Z(n11130) );
  NANDN U11276 ( .A(n11132), .B(n11131), .Z(n11127) );
  ANDN U11277 ( .B(B[226]), .A(n39), .Z(n10922) );
  XNOR U11278 ( .A(n10930), .B(n11133), .Z(n10923) );
  XNOR U11279 ( .A(n10929), .B(n10927), .Z(n11133) );
  AND U11280 ( .A(n11134), .B(n11135), .Z(n10927) );
  NANDN U11281 ( .A(n11136), .B(n11137), .Z(n11135) );
  OR U11282 ( .A(n11138), .B(n11139), .Z(n11137) );
  NAND U11283 ( .A(n11139), .B(n11138), .Z(n11134) );
  ANDN U11284 ( .B(B[227]), .A(n40), .Z(n10929) );
  XNOR U11285 ( .A(n10937), .B(n11140), .Z(n10930) );
  XNOR U11286 ( .A(n10936), .B(n10934), .Z(n11140) );
  AND U11287 ( .A(n11141), .B(n11142), .Z(n10934) );
  NANDN U11288 ( .A(n11143), .B(n11144), .Z(n11142) );
  NAND U11289 ( .A(n11145), .B(n11146), .Z(n11144) );
  ANDN U11290 ( .B(B[228]), .A(n41), .Z(n10936) );
  XOR U11291 ( .A(n10943), .B(n11147), .Z(n10937) );
  XNOR U11292 ( .A(n10941), .B(n10944), .Z(n11147) );
  NAND U11293 ( .A(A[2]), .B(B[229]), .Z(n10944) );
  NANDN U11294 ( .A(n11148), .B(n11149), .Z(n10941) );
  AND U11295 ( .A(A[0]), .B(B[230]), .Z(n11149) );
  XNOR U11296 ( .A(n10946), .B(n11150), .Z(n10943) );
  NAND U11297 ( .A(A[0]), .B(B[231]), .Z(n11150) );
  NAND U11298 ( .A(B[230]), .B(A[1]), .Z(n10946) );
  NAND U11299 ( .A(n11151), .B(n11152), .Z(n277) );
  NANDN U11300 ( .A(n11153), .B(n11154), .Z(n11152) );
  OR U11301 ( .A(n11155), .B(n11156), .Z(n11154) );
  NAND U11302 ( .A(n11156), .B(n11155), .Z(n11151) );
  XOR U11303 ( .A(n281), .B(n280), .Z(\A1[228] ) );
  XOR U11304 ( .A(n11156), .B(n11157), .Z(n280) );
  XNOR U11305 ( .A(n11155), .B(n11153), .Z(n11157) );
  AND U11306 ( .A(n11158), .B(n11159), .Z(n11153) );
  NANDN U11307 ( .A(n11160), .B(n11161), .Z(n11159) );
  NANDN U11308 ( .A(n11162), .B(n11163), .Z(n11161) );
  NANDN U11309 ( .A(n11163), .B(n11162), .Z(n11158) );
  ANDN U11310 ( .B(B[215]), .A(n29), .Z(n11155) );
  XNOR U11311 ( .A(n11062), .B(n11164), .Z(n11156) );
  XNOR U11312 ( .A(n11061), .B(n11059), .Z(n11164) );
  AND U11313 ( .A(n11165), .B(n11166), .Z(n11059) );
  NANDN U11314 ( .A(n11167), .B(n11168), .Z(n11166) );
  OR U11315 ( .A(n11169), .B(n11170), .Z(n11168) );
  NAND U11316 ( .A(n11170), .B(n11169), .Z(n11165) );
  ANDN U11317 ( .B(B[216]), .A(n30), .Z(n11061) );
  XNOR U11318 ( .A(n11069), .B(n11171), .Z(n11062) );
  XNOR U11319 ( .A(n11068), .B(n11066), .Z(n11171) );
  AND U11320 ( .A(n11172), .B(n11173), .Z(n11066) );
  NANDN U11321 ( .A(n11174), .B(n11175), .Z(n11173) );
  NANDN U11322 ( .A(n11176), .B(n11177), .Z(n11175) );
  NANDN U11323 ( .A(n11177), .B(n11176), .Z(n11172) );
  ANDN U11324 ( .B(B[217]), .A(n31), .Z(n11068) );
  XNOR U11325 ( .A(n11076), .B(n11178), .Z(n11069) );
  XNOR U11326 ( .A(n11075), .B(n11073), .Z(n11178) );
  AND U11327 ( .A(n11179), .B(n11180), .Z(n11073) );
  NANDN U11328 ( .A(n11181), .B(n11182), .Z(n11180) );
  OR U11329 ( .A(n11183), .B(n11184), .Z(n11182) );
  NAND U11330 ( .A(n11184), .B(n11183), .Z(n11179) );
  ANDN U11331 ( .B(B[218]), .A(n32), .Z(n11075) );
  XNOR U11332 ( .A(n11083), .B(n11185), .Z(n11076) );
  XNOR U11333 ( .A(n11082), .B(n11080), .Z(n11185) );
  AND U11334 ( .A(n11186), .B(n11187), .Z(n11080) );
  NANDN U11335 ( .A(n11188), .B(n11189), .Z(n11187) );
  NANDN U11336 ( .A(n11190), .B(n11191), .Z(n11189) );
  NANDN U11337 ( .A(n11191), .B(n11190), .Z(n11186) );
  ANDN U11338 ( .B(B[219]), .A(n33), .Z(n11082) );
  XNOR U11339 ( .A(n11090), .B(n11192), .Z(n11083) );
  XNOR U11340 ( .A(n11089), .B(n11087), .Z(n11192) );
  AND U11341 ( .A(n11193), .B(n11194), .Z(n11087) );
  NANDN U11342 ( .A(n11195), .B(n11196), .Z(n11194) );
  OR U11343 ( .A(n11197), .B(n11198), .Z(n11196) );
  NAND U11344 ( .A(n11198), .B(n11197), .Z(n11193) );
  ANDN U11345 ( .B(B[220]), .A(n34), .Z(n11089) );
  XNOR U11346 ( .A(n11097), .B(n11199), .Z(n11090) );
  XNOR U11347 ( .A(n11096), .B(n11094), .Z(n11199) );
  AND U11348 ( .A(n11200), .B(n11201), .Z(n11094) );
  NANDN U11349 ( .A(n11202), .B(n11203), .Z(n11201) );
  NANDN U11350 ( .A(n11204), .B(n11205), .Z(n11203) );
  NANDN U11351 ( .A(n11205), .B(n11204), .Z(n11200) );
  ANDN U11352 ( .B(B[221]), .A(n35), .Z(n11096) );
  XNOR U11353 ( .A(n11104), .B(n11206), .Z(n11097) );
  XNOR U11354 ( .A(n11103), .B(n11101), .Z(n11206) );
  AND U11355 ( .A(n11207), .B(n11208), .Z(n11101) );
  NANDN U11356 ( .A(n11209), .B(n11210), .Z(n11208) );
  OR U11357 ( .A(n11211), .B(n11212), .Z(n11210) );
  NAND U11358 ( .A(n11212), .B(n11211), .Z(n11207) );
  ANDN U11359 ( .B(B[222]), .A(n36), .Z(n11103) );
  XNOR U11360 ( .A(n11111), .B(n11213), .Z(n11104) );
  XNOR U11361 ( .A(n11110), .B(n11108), .Z(n11213) );
  AND U11362 ( .A(n11214), .B(n11215), .Z(n11108) );
  NANDN U11363 ( .A(n11216), .B(n11217), .Z(n11215) );
  NANDN U11364 ( .A(n11218), .B(n11219), .Z(n11217) );
  NANDN U11365 ( .A(n11219), .B(n11218), .Z(n11214) );
  ANDN U11366 ( .B(B[223]), .A(n37), .Z(n11110) );
  XNOR U11367 ( .A(n11118), .B(n11220), .Z(n11111) );
  XNOR U11368 ( .A(n11117), .B(n11115), .Z(n11220) );
  AND U11369 ( .A(n11221), .B(n11222), .Z(n11115) );
  NANDN U11370 ( .A(n11223), .B(n11224), .Z(n11222) );
  OR U11371 ( .A(n11225), .B(n11226), .Z(n11224) );
  NAND U11372 ( .A(n11226), .B(n11225), .Z(n11221) );
  ANDN U11373 ( .B(B[224]), .A(n38), .Z(n11117) );
  XNOR U11374 ( .A(n11125), .B(n11227), .Z(n11118) );
  XNOR U11375 ( .A(n11124), .B(n11122), .Z(n11227) );
  AND U11376 ( .A(n11228), .B(n11229), .Z(n11122) );
  NANDN U11377 ( .A(n11230), .B(n11231), .Z(n11229) );
  NANDN U11378 ( .A(n11232), .B(n11233), .Z(n11231) );
  NANDN U11379 ( .A(n11233), .B(n11232), .Z(n11228) );
  ANDN U11380 ( .B(B[225]), .A(n39), .Z(n11124) );
  XNOR U11381 ( .A(n11132), .B(n11234), .Z(n11125) );
  XNOR U11382 ( .A(n11131), .B(n11129), .Z(n11234) );
  AND U11383 ( .A(n11235), .B(n11236), .Z(n11129) );
  NANDN U11384 ( .A(n11237), .B(n11238), .Z(n11236) );
  OR U11385 ( .A(n11239), .B(n11240), .Z(n11238) );
  NAND U11386 ( .A(n11240), .B(n11239), .Z(n11235) );
  ANDN U11387 ( .B(B[226]), .A(n40), .Z(n11131) );
  XNOR U11388 ( .A(n11139), .B(n11241), .Z(n11132) );
  XNOR U11389 ( .A(n11138), .B(n11136), .Z(n11241) );
  AND U11390 ( .A(n11242), .B(n11243), .Z(n11136) );
  NANDN U11391 ( .A(n11244), .B(n11245), .Z(n11243) );
  NAND U11392 ( .A(n11246), .B(n11247), .Z(n11245) );
  ANDN U11393 ( .B(B[227]), .A(n41), .Z(n11138) );
  XOR U11394 ( .A(n11145), .B(n11248), .Z(n11139) );
  XNOR U11395 ( .A(n11143), .B(n11146), .Z(n11248) );
  NAND U11396 ( .A(A[2]), .B(B[228]), .Z(n11146) );
  NANDN U11397 ( .A(n11249), .B(n11250), .Z(n11143) );
  AND U11398 ( .A(A[0]), .B(B[229]), .Z(n11250) );
  XNOR U11399 ( .A(n11148), .B(n11251), .Z(n11145) );
  NAND U11400 ( .A(A[0]), .B(B[230]), .Z(n11251) );
  NAND U11401 ( .A(B[229]), .B(A[1]), .Z(n11148) );
  NAND U11402 ( .A(n11252), .B(n11253), .Z(n281) );
  NANDN U11403 ( .A(n11254), .B(n11255), .Z(n11253) );
  OR U11404 ( .A(n11256), .B(n11257), .Z(n11255) );
  NAND U11405 ( .A(n11257), .B(n11256), .Z(n11252) );
  XOR U11406 ( .A(n283), .B(n282), .Z(\A1[227] ) );
  XOR U11407 ( .A(n11257), .B(n11258), .Z(n282) );
  XNOR U11408 ( .A(n11256), .B(n11254), .Z(n11258) );
  AND U11409 ( .A(n11259), .B(n11260), .Z(n11254) );
  NANDN U11410 ( .A(n11261), .B(n11262), .Z(n11260) );
  NANDN U11411 ( .A(n11263), .B(n11264), .Z(n11262) );
  NANDN U11412 ( .A(n11264), .B(n11263), .Z(n11259) );
  ANDN U11413 ( .B(B[214]), .A(n29), .Z(n11256) );
  XNOR U11414 ( .A(n11163), .B(n11265), .Z(n11257) );
  XNOR U11415 ( .A(n11162), .B(n11160), .Z(n11265) );
  AND U11416 ( .A(n11266), .B(n11267), .Z(n11160) );
  NANDN U11417 ( .A(n11268), .B(n11269), .Z(n11267) );
  OR U11418 ( .A(n11270), .B(n11271), .Z(n11269) );
  NAND U11419 ( .A(n11271), .B(n11270), .Z(n11266) );
  ANDN U11420 ( .B(B[215]), .A(n30), .Z(n11162) );
  XNOR U11421 ( .A(n11170), .B(n11272), .Z(n11163) );
  XNOR U11422 ( .A(n11169), .B(n11167), .Z(n11272) );
  AND U11423 ( .A(n11273), .B(n11274), .Z(n11167) );
  NANDN U11424 ( .A(n11275), .B(n11276), .Z(n11274) );
  NANDN U11425 ( .A(n11277), .B(n11278), .Z(n11276) );
  NANDN U11426 ( .A(n11278), .B(n11277), .Z(n11273) );
  ANDN U11427 ( .B(B[216]), .A(n31), .Z(n11169) );
  XNOR U11428 ( .A(n11177), .B(n11279), .Z(n11170) );
  XNOR U11429 ( .A(n11176), .B(n11174), .Z(n11279) );
  AND U11430 ( .A(n11280), .B(n11281), .Z(n11174) );
  NANDN U11431 ( .A(n11282), .B(n11283), .Z(n11281) );
  OR U11432 ( .A(n11284), .B(n11285), .Z(n11283) );
  NAND U11433 ( .A(n11285), .B(n11284), .Z(n11280) );
  ANDN U11434 ( .B(B[217]), .A(n32), .Z(n11176) );
  XNOR U11435 ( .A(n11184), .B(n11286), .Z(n11177) );
  XNOR U11436 ( .A(n11183), .B(n11181), .Z(n11286) );
  AND U11437 ( .A(n11287), .B(n11288), .Z(n11181) );
  NANDN U11438 ( .A(n11289), .B(n11290), .Z(n11288) );
  NANDN U11439 ( .A(n11291), .B(n11292), .Z(n11290) );
  NANDN U11440 ( .A(n11292), .B(n11291), .Z(n11287) );
  ANDN U11441 ( .B(B[218]), .A(n33), .Z(n11183) );
  XNOR U11442 ( .A(n11191), .B(n11293), .Z(n11184) );
  XNOR U11443 ( .A(n11190), .B(n11188), .Z(n11293) );
  AND U11444 ( .A(n11294), .B(n11295), .Z(n11188) );
  NANDN U11445 ( .A(n11296), .B(n11297), .Z(n11295) );
  OR U11446 ( .A(n11298), .B(n11299), .Z(n11297) );
  NAND U11447 ( .A(n11299), .B(n11298), .Z(n11294) );
  ANDN U11448 ( .B(B[219]), .A(n34), .Z(n11190) );
  XNOR U11449 ( .A(n11198), .B(n11300), .Z(n11191) );
  XNOR U11450 ( .A(n11197), .B(n11195), .Z(n11300) );
  AND U11451 ( .A(n11301), .B(n11302), .Z(n11195) );
  NANDN U11452 ( .A(n11303), .B(n11304), .Z(n11302) );
  NANDN U11453 ( .A(n11305), .B(n11306), .Z(n11304) );
  NANDN U11454 ( .A(n11306), .B(n11305), .Z(n11301) );
  ANDN U11455 ( .B(B[220]), .A(n35), .Z(n11197) );
  XNOR U11456 ( .A(n11205), .B(n11307), .Z(n11198) );
  XNOR U11457 ( .A(n11204), .B(n11202), .Z(n11307) );
  AND U11458 ( .A(n11308), .B(n11309), .Z(n11202) );
  NANDN U11459 ( .A(n11310), .B(n11311), .Z(n11309) );
  OR U11460 ( .A(n11312), .B(n11313), .Z(n11311) );
  NAND U11461 ( .A(n11313), .B(n11312), .Z(n11308) );
  ANDN U11462 ( .B(B[221]), .A(n36), .Z(n11204) );
  XNOR U11463 ( .A(n11212), .B(n11314), .Z(n11205) );
  XNOR U11464 ( .A(n11211), .B(n11209), .Z(n11314) );
  AND U11465 ( .A(n11315), .B(n11316), .Z(n11209) );
  NANDN U11466 ( .A(n11317), .B(n11318), .Z(n11316) );
  NANDN U11467 ( .A(n11319), .B(n11320), .Z(n11318) );
  NANDN U11468 ( .A(n11320), .B(n11319), .Z(n11315) );
  ANDN U11469 ( .B(B[222]), .A(n37), .Z(n11211) );
  XNOR U11470 ( .A(n11219), .B(n11321), .Z(n11212) );
  XNOR U11471 ( .A(n11218), .B(n11216), .Z(n11321) );
  AND U11472 ( .A(n11322), .B(n11323), .Z(n11216) );
  NANDN U11473 ( .A(n11324), .B(n11325), .Z(n11323) );
  OR U11474 ( .A(n11326), .B(n11327), .Z(n11325) );
  NAND U11475 ( .A(n11327), .B(n11326), .Z(n11322) );
  ANDN U11476 ( .B(B[223]), .A(n38), .Z(n11218) );
  XNOR U11477 ( .A(n11226), .B(n11328), .Z(n11219) );
  XNOR U11478 ( .A(n11225), .B(n11223), .Z(n11328) );
  AND U11479 ( .A(n11329), .B(n11330), .Z(n11223) );
  NANDN U11480 ( .A(n11331), .B(n11332), .Z(n11330) );
  NANDN U11481 ( .A(n11333), .B(n11334), .Z(n11332) );
  NANDN U11482 ( .A(n11334), .B(n11333), .Z(n11329) );
  ANDN U11483 ( .B(B[224]), .A(n39), .Z(n11225) );
  XNOR U11484 ( .A(n11233), .B(n11335), .Z(n11226) );
  XNOR U11485 ( .A(n11232), .B(n11230), .Z(n11335) );
  AND U11486 ( .A(n11336), .B(n11337), .Z(n11230) );
  NANDN U11487 ( .A(n11338), .B(n11339), .Z(n11337) );
  OR U11488 ( .A(n11340), .B(n11341), .Z(n11339) );
  NAND U11489 ( .A(n11341), .B(n11340), .Z(n11336) );
  ANDN U11490 ( .B(B[225]), .A(n40), .Z(n11232) );
  XNOR U11491 ( .A(n11240), .B(n11342), .Z(n11233) );
  XNOR U11492 ( .A(n11239), .B(n11237), .Z(n11342) );
  AND U11493 ( .A(n11343), .B(n11344), .Z(n11237) );
  NANDN U11494 ( .A(n11345), .B(n11346), .Z(n11344) );
  NAND U11495 ( .A(n11347), .B(n11348), .Z(n11346) );
  ANDN U11496 ( .B(B[226]), .A(n41), .Z(n11239) );
  XOR U11497 ( .A(n11246), .B(n11349), .Z(n11240) );
  XNOR U11498 ( .A(n11244), .B(n11247), .Z(n11349) );
  NAND U11499 ( .A(A[2]), .B(B[227]), .Z(n11247) );
  NANDN U11500 ( .A(n11350), .B(n11351), .Z(n11244) );
  AND U11501 ( .A(A[0]), .B(B[228]), .Z(n11351) );
  XNOR U11502 ( .A(n11249), .B(n11352), .Z(n11246) );
  NAND U11503 ( .A(A[0]), .B(B[229]), .Z(n11352) );
  NAND U11504 ( .A(B[228]), .B(A[1]), .Z(n11249) );
  NAND U11505 ( .A(n11353), .B(n11354), .Z(n283) );
  NANDN U11506 ( .A(n11355), .B(n11356), .Z(n11354) );
  OR U11507 ( .A(n11357), .B(n11358), .Z(n11356) );
  NAND U11508 ( .A(n11358), .B(n11357), .Z(n11353) );
  XOR U11509 ( .A(n285), .B(n284), .Z(\A1[226] ) );
  XOR U11510 ( .A(n11358), .B(n11359), .Z(n284) );
  XNOR U11511 ( .A(n11357), .B(n11355), .Z(n11359) );
  AND U11512 ( .A(n11360), .B(n11361), .Z(n11355) );
  NANDN U11513 ( .A(n11362), .B(n11363), .Z(n11361) );
  NANDN U11514 ( .A(n11364), .B(n11365), .Z(n11363) );
  NANDN U11515 ( .A(n11365), .B(n11364), .Z(n11360) );
  ANDN U11516 ( .B(B[213]), .A(n29), .Z(n11357) );
  XNOR U11517 ( .A(n11264), .B(n11366), .Z(n11358) );
  XNOR U11518 ( .A(n11263), .B(n11261), .Z(n11366) );
  AND U11519 ( .A(n11367), .B(n11368), .Z(n11261) );
  NANDN U11520 ( .A(n11369), .B(n11370), .Z(n11368) );
  OR U11521 ( .A(n11371), .B(n11372), .Z(n11370) );
  NAND U11522 ( .A(n11372), .B(n11371), .Z(n11367) );
  ANDN U11523 ( .B(B[214]), .A(n30), .Z(n11263) );
  XNOR U11524 ( .A(n11271), .B(n11373), .Z(n11264) );
  XNOR U11525 ( .A(n11270), .B(n11268), .Z(n11373) );
  AND U11526 ( .A(n11374), .B(n11375), .Z(n11268) );
  NANDN U11527 ( .A(n11376), .B(n11377), .Z(n11375) );
  NANDN U11528 ( .A(n11378), .B(n11379), .Z(n11377) );
  NANDN U11529 ( .A(n11379), .B(n11378), .Z(n11374) );
  ANDN U11530 ( .B(B[215]), .A(n31), .Z(n11270) );
  XNOR U11531 ( .A(n11278), .B(n11380), .Z(n11271) );
  XNOR U11532 ( .A(n11277), .B(n11275), .Z(n11380) );
  AND U11533 ( .A(n11381), .B(n11382), .Z(n11275) );
  NANDN U11534 ( .A(n11383), .B(n11384), .Z(n11382) );
  OR U11535 ( .A(n11385), .B(n11386), .Z(n11384) );
  NAND U11536 ( .A(n11386), .B(n11385), .Z(n11381) );
  ANDN U11537 ( .B(B[216]), .A(n32), .Z(n11277) );
  XNOR U11538 ( .A(n11285), .B(n11387), .Z(n11278) );
  XNOR U11539 ( .A(n11284), .B(n11282), .Z(n11387) );
  AND U11540 ( .A(n11388), .B(n11389), .Z(n11282) );
  NANDN U11541 ( .A(n11390), .B(n11391), .Z(n11389) );
  NANDN U11542 ( .A(n11392), .B(n11393), .Z(n11391) );
  NANDN U11543 ( .A(n11393), .B(n11392), .Z(n11388) );
  ANDN U11544 ( .B(B[217]), .A(n33), .Z(n11284) );
  XNOR U11545 ( .A(n11292), .B(n11394), .Z(n11285) );
  XNOR U11546 ( .A(n11291), .B(n11289), .Z(n11394) );
  AND U11547 ( .A(n11395), .B(n11396), .Z(n11289) );
  NANDN U11548 ( .A(n11397), .B(n11398), .Z(n11396) );
  OR U11549 ( .A(n11399), .B(n11400), .Z(n11398) );
  NAND U11550 ( .A(n11400), .B(n11399), .Z(n11395) );
  ANDN U11551 ( .B(B[218]), .A(n34), .Z(n11291) );
  XNOR U11552 ( .A(n11299), .B(n11401), .Z(n11292) );
  XNOR U11553 ( .A(n11298), .B(n11296), .Z(n11401) );
  AND U11554 ( .A(n11402), .B(n11403), .Z(n11296) );
  NANDN U11555 ( .A(n11404), .B(n11405), .Z(n11403) );
  NANDN U11556 ( .A(n11406), .B(n11407), .Z(n11405) );
  NANDN U11557 ( .A(n11407), .B(n11406), .Z(n11402) );
  ANDN U11558 ( .B(B[219]), .A(n35), .Z(n11298) );
  XNOR U11559 ( .A(n11306), .B(n11408), .Z(n11299) );
  XNOR U11560 ( .A(n11305), .B(n11303), .Z(n11408) );
  AND U11561 ( .A(n11409), .B(n11410), .Z(n11303) );
  NANDN U11562 ( .A(n11411), .B(n11412), .Z(n11410) );
  OR U11563 ( .A(n11413), .B(n11414), .Z(n11412) );
  NAND U11564 ( .A(n11414), .B(n11413), .Z(n11409) );
  ANDN U11565 ( .B(B[220]), .A(n36), .Z(n11305) );
  XNOR U11566 ( .A(n11313), .B(n11415), .Z(n11306) );
  XNOR U11567 ( .A(n11312), .B(n11310), .Z(n11415) );
  AND U11568 ( .A(n11416), .B(n11417), .Z(n11310) );
  NANDN U11569 ( .A(n11418), .B(n11419), .Z(n11417) );
  NANDN U11570 ( .A(n11420), .B(n11421), .Z(n11419) );
  NANDN U11571 ( .A(n11421), .B(n11420), .Z(n11416) );
  ANDN U11572 ( .B(B[221]), .A(n37), .Z(n11312) );
  XNOR U11573 ( .A(n11320), .B(n11422), .Z(n11313) );
  XNOR U11574 ( .A(n11319), .B(n11317), .Z(n11422) );
  AND U11575 ( .A(n11423), .B(n11424), .Z(n11317) );
  NANDN U11576 ( .A(n11425), .B(n11426), .Z(n11424) );
  OR U11577 ( .A(n11427), .B(n11428), .Z(n11426) );
  NAND U11578 ( .A(n11428), .B(n11427), .Z(n11423) );
  ANDN U11579 ( .B(B[222]), .A(n38), .Z(n11319) );
  XNOR U11580 ( .A(n11327), .B(n11429), .Z(n11320) );
  XNOR U11581 ( .A(n11326), .B(n11324), .Z(n11429) );
  AND U11582 ( .A(n11430), .B(n11431), .Z(n11324) );
  NANDN U11583 ( .A(n11432), .B(n11433), .Z(n11431) );
  NANDN U11584 ( .A(n11434), .B(n11435), .Z(n11433) );
  NANDN U11585 ( .A(n11435), .B(n11434), .Z(n11430) );
  ANDN U11586 ( .B(B[223]), .A(n39), .Z(n11326) );
  XNOR U11587 ( .A(n11334), .B(n11436), .Z(n11327) );
  XNOR U11588 ( .A(n11333), .B(n11331), .Z(n11436) );
  AND U11589 ( .A(n11437), .B(n11438), .Z(n11331) );
  NANDN U11590 ( .A(n11439), .B(n11440), .Z(n11438) );
  OR U11591 ( .A(n11441), .B(n11442), .Z(n11440) );
  NAND U11592 ( .A(n11442), .B(n11441), .Z(n11437) );
  ANDN U11593 ( .B(B[224]), .A(n40), .Z(n11333) );
  XNOR U11594 ( .A(n11341), .B(n11443), .Z(n11334) );
  XNOR U11595 ( .A(n11340), .B(n11338), .Z(n11443) );
  AND U11596 ( .A(n11444), .B(n11445), .Z(n11338) );
  NANDN U11597 ( .A(n11446), .B(n11447), .Z(n11445) );
  NAND U11598 ( .A(n11448), .B(n11449), .Z(n11447) );
  ANDN U11599 ( .B(B[225]), .A(n41), .Z(n11340) );
  XOR U11600 ( .A(n11347), .B(n11450), .Z(n11341) );
  XNOR U11601 ( .A(n11345), .B(n11348), .Z(n11450) );
  NAND U11602 ( .A(A[2]), .B(B[226]), .Z(n11348) );
  NANDN U11603 ( .A(n11451), .B(n11452), .Z(n11345) );
  AND U11604 ( .A(A[0]), .B(B[227]), .Z(n11452) );
  XNOR U11605 ( .A(n11350), .B(n11453), .Z(n11347) );
  NAND U11606 ( .A(A[0]), .B(B[228]), .Z(n11453) );
  NAND U11607 ( .A(B[227]), .B(A[1]), .Z(n11350) );
  NAND U11608 ( .A(n11454), .B(n11455), .Z(n285) );
  NANDN U11609 ( .A(n11456), .B(n11457), .Z(n11455) );
  OR U11610 ( .A(n11458), .B(n11459), .Z(n11457) );
  NAND U11611 ( .A(n11459), .B(n11458), .Z(n11454) );
  XOR U11612 ( .A(n287), .B(n286), .Z(\A1[225] ) );
  XOR U11613 ( .A(n11459), .B(n11460), .Z(n286) );
  XNOR U11614 ( .A(n11458), .B(n11456), .Z(n11460) );
  AND U11615 ( .A(n11461), .B(n11462), .Z(n11456) );
  NANDN U11616 ( .A(n11463), .B(n11464), .Z(n11462) );
  NANDN U11617 ( .A(n11465), .B(n11466), .Z(n11464) );
  NANDN U11618 ( .A(n11466), .B(n11465), .Z(n11461) );
  ANDN U11619 ( .B(B[212]), .A(n29), .Z(n11458) );
  XNOR U11620 ( .A(n11365), .B(n11467), .Z(n11459) );
  XNOR U11621 ( .A(n11364), .B(n11362), .Z(n11467) );
  AND U11622 ( .A(n11468), .B(n11469), .Z(n11362) );
  NANDN U11623 ( .A(n11470), .B(n11471), .Z(n11469) );
  OR U11624 ( .A(n11472), .B(n11473), .Z(n11471) );
  NAND U11625 ( .A(n11473), .B(n11472), .Z(n11468) );
  ANDN U11626 ( .B(B[213]), .A(n30), .Z(n11364) );
  XNOR U11627 ( .A(n11372), .B(n11474), .Z(n11365) );
  XNOR U11628 ( .A(n11371), .B(n11369), .Z(n11474) );
  AND U11629 ( .A(n11475), .B(n11476), .Z(n11369) );
  NANDN U11630 ( .A(n11477), .B(n11478), .Z(n11476) );
  NANDN U11631 ( .A(n11479), .B(n11480), .Z(n11478) );
  NANDN U11632 ( .A(n11480), .B(n11479), .Z(n11475) );
  ANDN U11633 ( .B(B[214]), .A(n31), .Z(n11371) );
  XNOR U11634 ( .A(n11379), .B(n11481), .Z(n11372) );
  XNOR U11635 ( .A(n11378), .B(n11376), .Z(n11481) );
  AND U11636 ( .A(n11482), .B(n11483), .Z(n11376) );
  NANDN U11637 ( .A(n11484), .B(n11485), .Z(n11483) );
  OR U11638 ( .A(n11486), .B(n11487), .Z(n11485) );
  NAND U11639 ( .A(n11487), .B(n11486), .Z(n11482) );
  ANDN U11640 ( .B(B[215]), .A(n32), .Z(n11378) );
  XNOR U11641 ( .A(n11386), .B(n11488), .Z(n11379) );
  XNOR U11642 ( .A(n11385), .B(n11383), .Z(n11488) );
  AND U11643 ( .A(n11489), .B(n11490), .Z(n11383) );
  NANDN U11644 ( .A(n11491), .B(n11492), .Z(n11490) );
  NANDN U11645 ( .A(n11493), .B(n11494), .Z(n11492) );
  NANDN U11646 ( .A(n11494), .B(n11493), .Z(n11489) );
  ANDN U11647 ( .B(B[216]), .A(n33), .Z(n11385) );
  XNOR U11648 ( .A(n11393), .B(n11495), .Z(n11386) );
  XNOR U11649 ( .A(n11392), .B(n11390), .Z(n11495) );
  AND U11650 ( .A(n11496), .B(n11497), .Z(n11390) );
  NANDN U11651 ( .A(n11498), .B(n11499), .Z(n11497) );
  OR U11652 ( .A(n11500), .B(n11501), .Z(n11499) );
  NAND U11653 ( .A(n11501), .B(n11500), .Z(n11496) );
  ANDN U11654 ( .B(B[217]), .A(n34), .Z(n11392) );
  XNOR U11655 ( .A(n11400), .B(n11502), .Z(n11393) );
  XNOR U11656 ( .A(n11399), .B(n11397), .Z(n11502) );
  AND U11657 ( .A(n11503), .B(n11504), .Z(n11397) );
  NANDN U11658 ( .A(n11505), .B(n11506), .Z(n11504) );
  NANDN U11659 ( .A(n11507), .B(n11508), .Z(n11506) );
  NANDN U11660 ( .A(n11508), .B(n11507), .Z(n11503) );
  ANDN U11661 ( .B(B[218]), .A(n35), .Z(n11399) );
  XNOR U11662 ( .A(n11407), .B(n11509), .Z(n11400) );
  XNOR U11663 ( .A(n11406), .B(n11404), .Z(n11509) );
  AND U11664 ( .A(n11510), .B(n11511), .Z(n11404) );
  NANDN U11665 ( .A(n11512), .B(n11513), .Z(n11511) );
  OR U11666 ( .A(n11514), .B(n11515), .Z(n11513) );
  NAND U11667 ( .A(n11515), .B(n11514), .Z(n11510) );
  ANDN U11668 ( .B(B[219]), .A(n36), .Z(n11406) );
  XNOR U11669 ( .A(n11414), .B(n11516), .Z(n11407) );
  XNOR U11670 ( .A(n11413), .B(n11411), .Z(n11516) );
  AND U11671 ( .A(n11517), .B(n11518), .Z(n11411) );
  NANDN U11672 ( .A(n11519), .B(n11520), .Z(n11518) );
  NANDN U11673 ( .A(n11521), .B(n11522), .Z(n11520) );
  NANDN U11674 ( .A(n11522), .B(n11521), .Z(n11517) );
  ANDN U11675 ( .B(B[220]), .A(n37), .Z(n11413) );
  XNOR U11676 ( .A(n11421), .B(n11523), .Z(n11414) );
  XNOR U11677 ( .A(n11420), .B(n11418), .Z(n11523) );
  AND U11678 ( .A(n11524), .B(n11525), .Z(n11418) );
  NANDN U11679 ( .A(n11526), .B(n11527), .Z(n11525) );
  OR U11680 ( .A(n11528), .B(n11529), .Z(n11527) );
  NAND U11681 ( .A(n11529), .B(n11528), .Z(n11524) );
  ANDN U11682 ( .B(B[221]), .A(n38), .Z(n11420) );
  XNOR U11683 ( .A(n11428), .B(n11530), .Z(n11421) );
  XNOR U11684 ( .A(n11427), .B(n11425), .Z(n11530) );
  AND U11685 ( .A(n11531), .B(n11532), .Z(n11425) );
  NANDN U11686 ( .A(n11533), .B(n11534), .Z(n11532) );
  NANDN U11687 ( .A(n11535), .B(n11536), .Z(n11534) );
  NANDN U11688 ( .A(n11536), .B(n11535), .Z(n11531) );
  ANDN U11689 ( .B(B[222]), .A(n39), .Z(n11427) );
  XNOR U11690 ( .A(n11435), .B(n11537), .Z(n11428) );
  XNOR U11691 ( .A(n11434), .B(n11432), .Z(n11537) );
  AND U11692 ( .A(n11538), .B(n11539), .Z(n11432) );
  NANDN U11693 ( .A(n11540), .B(n11541), .Z(n11539) );
  OR U11694 ( .A(n11542), .B(n11543), .Z(n11541) );
  NAND U11695 ( .A(n11543), .B(n11542), .Z(n11538) );
  ANDN U11696 ( .B(B[223]), .A(n40), .Z(n11434) );
  XNOR U11697 ( .A(n11442), .B(n11544), .Z(n11435) );
  XNOR U11698 ( .A(n11441), .B(n11439), .Z(n11544) );
  AND U11699 ( .A(n11545), .B(n11546), .Z(n11439) );
  NANDN U11700 ( .A(n11547), .B(n11548), .Z(n11546) );
  NAND U11701 ( .A(n11549), .B(n11550), .Z(n11548) );
  ANDN U11702 ( .B(B[224]), .A(n41), .Z(n11441) );
  XOR U11703 ( .A(n11448), .B(n11551), .Z(n11442) );
  XNOR U11704 ( .A(n11446), .B(n11449), .Z(n11551) );
  NAND U11705 ( .A(A[2]), .B(B[225]), .Z(n11449) );
  NANDN U11706 ( .A(n11552), .B(n11553), .Z(n11446) );
  AND U11707 ( .A(A[0]), .B(B[226]), .Z(n11553) );
  XNOR U11708 ( .A(n11451), .B(n11554), .Z(n11448) );
  NAND U11709 ( .A(A[0]), .B(B[227]), .Z(n11554) );
  NAND U11710 ( .A(B[226]), .B(A[1]), .Z(n11451) );
  NAND U11711 ( .A(n11555), .B(n11556), .Z(n287) );
  NANDN U11712 ( .A(n11557), .B(n11558), .Z(n11556) );
  OR U11713 ( .A(n11559), .B(n11560), .Z(n11558) );
  NAND U11714 ( .A(n11560), .B(n11559), .Z(n11555) );
  XOR U11715 ( .A(n289), .B(n288), .Z(\A1[224] ) );
  XOR U11716 ( .A(n11560), .B(n11561), .Z(n288) );
  XNOR U11717 ( .A(n11559), .B(n11557), .Z(n11561) );
  AND U11718 ( .A(n11562), .B(n11563), .Z(n11557) );
  NANDN U11719 ( .A(n11564), .B(n11565), .Z(n11563) );
  NANDN U11720 ( .A(n11566), .B(n11567), .Z(n11565) );
  NANDN U11721 ( .A(n11567), .B(n11566), .Z(n11562) );
  ANDN U11722 ( .B(B[211]), .A(n29), .Z(n11559) );
  XNOR U11723 ( .A(n11466), .B(n11568), .Z(n11560) );
  XNOR U11724 ( .A(n11465), .B(n11463), .Z(n11568) );
  AND U11725 ( .A(n11569), .B(n11570), .Z(n11463) );
  NANDN U11726 ( .A(n11571), .B(n11572), .Z(n11570) );
  OR U11727 ( .A(n11573), .B(n11574), .Z(n11572) );
  NAND U11728 ( .A(n11574), .B(n11573), .Z(n11569) );
  ANDN U11729 ( .B(B[212]), .A(n30), .Z(n11465) );
  XNOR U11730 ( .A(n11473), .B(n11575), .Z(n11466) );
  XNOR U11731 ( .A(n11472), .B(n11470), .Z(n11575) );
  AND U11732 ( .A(n11576), .B(n11577), .Z(n11470) );
  NANDN U11733 ( .A(n11578), .B(n11579), .Z(n11577) );
  NANDN U11734 ( .A(n11580), .B(n11581), .Z(n11579) );
  NANDN U11735 ( .A(n11581), .B(n11580), .Z(n11576) );
  ANDN U11736 ( .B(B[213]), .A(n31), .Z(n11472) );
  XNOR U11737 ( .A(n11480), .B(n11582), .Z(n11473) );
  XNOR U11738 ( .A(n11479), .B(n11477), .Z(n11582) );
  AND U11739 ( .A(n11583), .B(n11584), .Z(n11477) );
  NANDN U11740 ( .A(n11585), .B(n11586), .Z(n11584) );
  OR U11741 ( .A(n11587), .B(n11588), .Z(n11586) );
  NAND U11742 ( .A(n11588), .B(n11587), .Z(n11583) );
  ANDN U11743 ( .B(B[214]), .A(n32), .Z(n11479) );
  XNOR U11744 ( .A(n11487), .B(n11589), .Z(n11480) );
  XNOR U11745 ( .A(n11486), .B(n11484), .Z(n11589) );
  AND U11746 ( .A(n11590), .B(n11591), .Z(n11484) );
  NANDN U11747 ( .A(n11592), .B(n11593), .Z(n11591) );
  NANDN U11748 ( .A(n11594), .B(n11595), .Z(n11593) );
  NANDN U11749 ( .A(n11595), .B(n11594), .Z(n11590) );
  ANDN U11750 ( .B(B[215]), .A(n33), .Z(n11486) );
  XNOR U11751 ( .A(n11494), .B(n11596), .Z(n11487) );
  XNOR U11752 ( .A(n11493), .B(n11491), .Z(n11596) );
  AND U11753 ( .A(n11597), .B(n11598), .Z(n11491) );
  NANDN U11754 ( .A(n11599), .B(n11600), .Z(n11598) );
  OR U11755 ( .A(n11601), .B(n11602), .Z(n11600) );
  NAND U11756 ( .A(n11602), .B(n11601), .Z(n11597) );
  ANDN U11757 ( .B(B[216]), .A(n34), .Z(n11493) );
  XNOR U11758 ( .A(n11501), .B(n11603), .Z(n11494) );
  XNOR U11759 ( .A(n11500), .B(n11498), .Z(n11603) );
  AND U11760 ( .A(n11604), .B(n11605), .Z(n11498) );
  NANDN U11761 ( .A(n11606), .B(n11607), .Z(n11605) );
  NANDN U11762 ( .A(n11608), .B(n11609), .Z(n11607) );
  NANDN U11763 ( .A(n11609), .B(n11608), .Z(n11604) );
  ANDN U11764 ( .B(B[217]), .A(n35), .Z(n11500) );
  XNOR U11765 ( .A(n11508), .B(n11610), .Z(n11501) );
  XNOR U11766 ( .A(n11507), .B(n11505), .Z(n11610) );
  AND U11767 ( .A(n11611), .B(n11612), .Z(n11505) );
  NANDN U11768 ( .A(n11613), .B(n11614), .Z(n11612) );
  OR U11769 ( .A(n11615), .B(n11616), .Z(n11614) );
  NAND U11770 ( .A(n11616), .B(n11615), .Z(n11611) );
  ANDN U11771 ( .B(B[218]), .A(n36), .Z(n11507) );
  XNOR U11772 ( .A(n11515), .B(n11617), .Z(n11508) );
  XNOR U11773 ( .A(n11514), .B(n11512), .Z(n11617) );
  AND U11774 ( .A(n11618), .B(n11619), .Z(n11512) );
  NANDN U11775 ( .A(n11620), .B(n11621), .Z(n11619) );
  NANDN U11776 ( .A(n11622), .B(n11623), .Z(n11621) );
  NANDN U11777 ( .A(n11623), .B(n11622), .Z(n11618) );
  ANDN U11778 ( .B(B[219]), .A(n37), .Z(n11514) );
  XNOR U11779 ( .A(n11522), .B(n11624), .Z(n11515) );
  XNOR U11780 ( .A(n11521), .B(n11519), .Z(n11624) );
  AND U11781 ( .A(n11625), .B(n11626), .Z(n11519) );
  NANDN U11782 ( .A(n11627), .B(n11628), .Z(n11626) );
  OR U11783 ( .A(n11629), .B(n11630), .Z(n11628) );
  NAND U11784 ( .A(n11630), .B(n11629), .Z(n11625) );
  ANDN U11785 ( .B(B[220]), .A(n38), .Z(n11521) );
  XNOR U11786 ( .A(n11529), .B(n11631), .Z(n11522) );
  XNOR U11787 ( .A(n11528), .B(n11526), .Z(n11631) );
  AND U11788 ( .A(n11632), .B(n11633), .Z(n11526) );
  NANDN U11789 ( .A(n11634), .B(n11635), .Z(n11633) );
  NANDN U11790 ( .A(n11636), .B(n11637), .Z(n11635) );
  NANDN U11791 ( .A(n11637), .B(n11636), .Z(n11632) );
  ANDN U11792 ( .B(B[221]), .A(n39), .Z(n11528) );
  XNOR U11793 ( .A(n11536), .B(n11638), .Z(n11529) );
  XNOR U11794 ( .A(n11535), .B(n11533), .Z(n11638) );
  AND U11795 ( .A(n11639), .B(n11640), .Z(n11533) );
  NANDN U11796 ( .A(n11641), .B(n11642), .Z(n11640) );
  OR U11797 ( .A(n11643), .B(n11644), .Z(n11642) );
  NAND U11798 ( .A(n11644), .B(n11643), .Z(n11639) );
  ANDN U11799 ( .B(B[222]), .A(n40), .Z(n11535) );
  XNOR U11800 ( .A(n11543), .B(n11645), .Z(n11536) );
  XNOR U11801 ( .A(n11542), .B(n11540), .Z(n11645) );
  AND U11802 ( .A(n11646), .B(n11647), .Z(n11540) );
  NANDN U11803 ( .A(n11648), .B(n11649), .Z(n11647) );
  NAND U11804 ( .A(n11650), .B(n11651), .Z(n11649) );
  ANDN U11805 ( .B(B[223]), .A(n41), .Z(n11542) );
  XOR U11806 ( .A(n11549), .B(n11652), .Z(n11543) );
  XNOR U11807 ( .A(n11547), .B(n11550), .Z(n11652) );
  NAND U11808 ( .A(A[2]), .B(B[224]), .Z(n11550) );
  NANDN U11809 ( .A(n11653), .B(n11654), .Z(n11547) );
  AND U11810 ( .A(A[0]), .B(B[225]), .Z(n11654) );
  XNOR U11811 ( .A(n11552), .B(n11655), .Z(n11549) );
  NAND U11812 ( .A(A[0]), .B(B[226]), .Z(n11655) );
  NAND U11813 ( .A(B[225]), .B(A[1]), .Z(n11552) );
  NAND U11814 ( .A(n11656), .B(n11657), .Z(n289) );
  NANDN U11815 ( .A(n11658), .B(n11659), .Z(n11657) );
  OR U11816 ( .A(n11660), .B(n11661), .Z(n11659) );
  NAND U11817 ( .A(n11661), .B(n11660), .Z(n11656) );
  XOR U11818 ( .A(n291), .B(n290), .Z(\A1[223] ) );
  XOR U11819 ( .A(n11661), .B(n11662), .Z(n290) );
  XNOR U11820 ( .A(n11660), .B(n11658), .Z(n11662) );
  AND U11821 ( .A(n11663), .B(n11664), .Z(n11658) );
  NANDN U11822 ( .A(n11665), .B(n11666), .Z(n11664) );
  NANDN U11823 ( .A(n11667), .B(n11668), .Z(n11666) );
  NANDN U11824 ( .A(n11668), .B(n11667), .Z(n11663) );
  ANDN U11825 ( .B(B[210]), .A(n29), .Z(n11660) );
  XNOR U11826 ( .A(n11567), .B(n11669), .Z(n11661) );
  XNOR U11827 ( .A(n11566), .B(n11564), .Z(n11669) );
  AND U11828 ( .A(n11670), .B(n11671), .Z(n11564) );
  NANDN U11829 ( .A(n11672), .B(n11673), .Z(n11671) );
  OR U11830 ( .A(n11674), .B(n11675), .Z(n11673) );
  NAND U11831 ( .A(n11675), .B(n11674), .Z(n11670) );
  ANDN U11832 ( .B(B[211]), .A(n30), .Z(n11566) );
  XNOR U11833 ( .A(n11574), .B(n11676), .Z(n11567) );
  XNOR U11834 ( .A(n11573), .B(n11571), .Z(n11676) );
  AND U11835 ( .A(n11677), .B(n11678), .Z(n11571) );
  NANDN U11836 ( .A(n11679), .B(n11680), .Z(n11678) );
  NANDN U11837 ( .A(n11681), .B(n11682), .Z(n11680) );
  NANDN U11838 ( .A(n11682), .B(n11681), .Z(n11677) );
  ANDN U11839 ( .B(B[212]), .A(n31), .Z(n11573) );
  XNOR U11840 ( .A(n11581), .B(n11683), .Z(n11574) );
  XNOR U11841 ( .A(n11580), .B(n11578), .Z(n11683) );
  AND U11842 ( .A(n11684), .B(n11685), .Z(n11578) );
  NANDN U11843 ( .A(n11686), .B(n11687), .Z(n11685) );
  OR U11844 ( .A(n11688), .B(n11689), .Z(n11687) );
  NAND U11845 ( .A(n11689), .B(n11688), .Z(n11684) );
  ANDN U11846 ( .B(B[213]), .A(n32), .Z(n11580) );
  XNOR U11847 ( .A(n11588), .B(n11690), .Z(n11581) );
  XNOR U11848 ( .A(n11587), .B(n11585), .Z(n11690) );
  AND U11849 ( .A(n11691), .B(n11692), .Z(n11585) );
  NANDN U11850 ( .A(n11693), .B(n11694), .Z(n11692) );
  NANDN U11851 ( .A(n11695), .B(n11696), .Z(n11694) );
  NANDN U11852 ( .A(n11696), .B(n11695), .Z(n11691) );
  ANDN U11853 ( .B(B[214]), .A(n33), .Z(n11587) );
  XNOR U11854 ( .A(n11595), .B(n11697), .Z(n11588) );
  XNOR U11855 ( .A(n11594), .B(n11592), .Z(n11697) );
  AND U11856 ( .A(n11698), .B(n11699), .Z(n11592) );
  NANDN U11857 ( .A(n11700), .B(n11701), .Z(n11699) );
  OR U11858 ( .A(n11702), .B(n11703), .Z(n11701) );
  NAND U11859 ( .A(n11703), .B(n11702), .Z(n11698) );
  ANDN U11860 ( .B(B[215]), .A(n34), .Z(n11594) );
  XNOR U11861 ( .A(n11602), .B(n11704), .Z(n11595) );
  XNOR U11862 ( .A(n11601), .B(n11599), .Z(n11704) );
  AND U11863 ( .A(n11705), .B(n11706), .Z(n11599) );
  NANDN U11864 ( .A(n11707), .B(n11708), .Z(n11706) );
  NANDN U11865 ( .A(n11709), .B(n11710), .Z(n11708) );
  NANDN U11866 ( .A(n11710), .B(n11709), .Z(n11705) );
  ANDN U11867 ( .B(B[216]), .A(n35), .Z(n11601) );
  XNOR U11868 ( .A(n11609), .B(n11711), .Z(n11602) );
  XNOR U11869 ( .A(n11608), .B(n11606), .Z(n11711) );
  AND U11870 ( .A(n11712), .B(n11713), .Z(n11606) );
  NANDN U11871 ( .A(n11714), .B(n11715), .Z(n11713) );
  OR U11872 ( .A(n11716), .B(n11717), .Z(n11715) );
  NAND U11873 ( .A(n11717), .B(n11716), .Z(n11712) );
  ANDN U11874 ( .B(B[217]), .A(n36), .Z(n11608) );
  XNOR U11875 ( .A(n11616), .B(n11718), .Z(n11609) );
  XNOR U11876 ( .A(n11615), .B(n11613), .Z(n11718) );
  AND U11877 ( .A(n11719), .B(n11720), .Z(n11613) );
  NANDN U11878 ( .A(n11721), .B(n11722), .Z(n11720) );
  NANDN U11879 ( .A(n11723), .B(n11724), .Z(n11722) );
  NANDN U11880 ( .A(n11724), .B(n11723), .Z(n11719) );
  ANDN U11881 ( .B(B[218]), .A(n37), .Z(n11615) );
  XNOR U11882 ( .A(n11623), .B(n11725), .Z(n11616) );
  XNOR U11883 ( .A(n11622), .B(n11620), .Z(n11725) );
  AND U11884 ( .A(n11726), .B(n11727), .Z(n11620) );
  NANDN U11885 ( .A(n11728), .B(n11729), .Z(n11727) );
  OR U11886 ( .A(n11730), .B(n11731), .Z(n11729) );
  NAND U11887 ( .A(n11731), .B(n11730), .Z(n11726) );
  ANDN U11888 ( .B(B[219]), .A(n38), .Z(n11622) );
  XNOR U11889 ( .A(n11630), .B(n11732), .Z(n11623) );
  XNOR U11890 ( .A(n11629), .B(n11627), .Z(n11732) );
  AND U11891 ( .A(n11733), .B(n11734), .Z(n11627) );
  NANDN U11892 ( .A(n11735), .B(n11736), .Z(n11734) );
  NANDN U11893 ( .A(n11737), .B(n11738), .Z(n11736) );
  NANDN U11894 ( .A(n11738), .B(n11737), .Z(n11733) );
  ANDN U11895 ( .B(B[220]), .A(n39), .Z(n11629) );
  XNOR U11896 ( .A(n11637), .B(n11739), .Z(n11630) );
  XNOR U11897 ( .A(n11636), .B(n11634), .Z(n11739) );
  AND U11898 ( .A(n11740), .B(n11741), .Z(n11634) );
  NANDN U11899 ( .A(n11742), .B(n11743), .Z(n11741) );
  OR U11900 ( .A(n11744), .B(n11745), .Z(n11743) );
  NAND U11901 ( .A(n11745), .B(n11744), .Z(n11740) );
  ANDN U11902 ( .B(B[221]), .A(n40), .Z(n11636) );
  XNOR U11903 ( .A(n11644), .B(n11746), .Z(n11637) );
  XNOR U11904 ( .A(n11643), .B(n11641), .Z(n11746) );
  AND U11905 ( .A(n11747), .B(n11748), .Z(n11641) );
  NANDN U11906 ( .A(n11749), .B(n11750), .Z(n11748) );
  NAND U11907 ( .A(n11751), .B(n11752), .Z(n11750) );
  ANDN U11908 ( .B(B[222]), .A(n41), .Z(n11643) );
  XOR U11909 ( .A(n11650), .B(n11753), .Z(n11644) );
  XNOR U11910 ( .A(n11648), .B(n11651), .Z(n11753) );
  NAND U11911 ( .A(A[2]), .B(B[223]), .Z(n11651) );
  NANDN U11912 ( .A(n11754), .B(n11755), .Z(n11648) );
  AND U11913 ( .A(A[0]), .B(B[224]), .Z(n11755) );
  XNOR U11914 ( .A(n11653), .B(n11756), .Z(n11650) );
  NAND U11915 ( .A(A[0]), .B(B[225]), .Z(n11756) );
  NAND U11916 ( .A(B[224]), .B(A[1]), .Z(n11653) );
  NAND U11917 ( .A(n11757), .B(n11758), .Z(n291) );
  NANDN U11918 ( .A(n11759), .B(n11760), .Z(n11758) );
  OR U11919 ( .A(n11761), .B(n11762), .Z(n11760) );
  NAND U11920 ( .A(n11762), .B(n11761), .Z(n11757) );
  XOR U11921 ( .A(n293), .B(n292), .Z(\A1[222] ) );
  XOR U11922 ( .A(n11762), .B(n11763), .Z(n292) );
  XNOR U11923 ( .A(n11761), .B(n11759), .Z(n11763) );
  AND U11924 ( .A(n11764), .B(n11765), .Z(n11759) );
  NANDN U11925 ( .A(n11766), .B(n11767), .Z(n11765) );
  NANDN U11926 ( .A(n11768), .B(n11769), .Z(n11767) );
  NANDN U11927 ( .A(n11769), .B(n11768), .Z(n11764) );
  ANDN U11928 ( .B(B[209]), .A(n29), .Z(n11761) );
  XNOR U11929 ( .A(n11668), .B(n11770), .Z(n11762) );
  XNOR U11930 ( .A(n11667), .B(n11665), .Z(n11770) );
  AND U11931 ( .A(n11771), .B(n11772), .Z(n11665) );
  NANDN U11932 ( .A(n11773), .B(n11774), .Z(n11772) );
  OR U11933 ( .A(n11775), .B(n11776), .Z(n11774) );
  NAND U11934 ( .A(n11776), .B(n11775), .Z(n11771) );
  ANDN U11935 ( .B(B[210]), .A(n30), .Z(n11667) );
  XNOR U11936 ( .A(n11675), .B(n11777), .Z(n11668) );
  XNOR U11937 ( .A(n11674), .B(n11672), .Z(n11777) );
  AND U11938 ( .A(n11778), .B(n11779), .Z(n11672) );
  NANDN U11939 ( .A(n11780), .B(n11781), .Z(n11779) );
  NANDN U11940 ( .A(n11782), .B(n11783), .Z(n11781) );
  NANDN U11941 ( .A(n11783), .B(n11782), .Z(n11778) );
  ANDN U11942 ( .B(B[211]), .A(n31), .Z(n11674) );
  XNOR U11943 ( .A(n11682), .B(n11784), .Z(n11675) );
  XNOR U11944 ( .A(n11681), .B(n11679), .Z(n11784) );
  AND U11945 ( .A(n11785), .B(n11786), .Z(n11679) );
  NANDN U11946 ( .A(n11787), .B(n11788), .Z(n11786) );
  OR U11947 ( .A(n11789), .B(n11790), .Z(n11788) );
  NAND U11948 ( .A(n11790), .B(n11789), .Z(n11785) );
  ANDN U11949 ( .B(B[212]), .A(n32), .Z(n11681) );
  XNOR U11950 ( .A(n11689), .B(n11791), .Z(n11682) );
  XNOR U11951 ( .A(n11688), .B(n11686), .Z(n11791) );
  AND U11952 ( .A(n11792), .B(n11793), .Z(n11686) );
  NANDN U11953 ( .A(n11794), .B(n11795), .Z(n11793) );
  NANDN U11954 ( .A(n11796), .B(n11797), .Z(n11795) );
  NANDN U11955 ( .A(n11797), .B(n11796), .Z(n11792) );
  ANDN U11956 ( .B(B[213]), .A(n33), .Z(n11688) );
  XNOR U11957 ( .A(n11696), .B(n11798), .Z(n11689) );
  XNOR U11958 ( .A(n11695), .B(n11693), .Z(n11798) );
  AND U11959 ( .A(n11799), .B(n11800), .Z(n11693) );
  NANDN U11960 ( .A(n11801), .B(n11802), .Z(n11800) );
  OR U11961 ( .A(n11803), .B(n11804), .Z(n11802) );
  NAND U11962 ( .A(n11804), .B(n11803), .Z(n11799) );
  ANDN U11963 ( .B(B[214]), .A(n34), .Z(n11695) );
  XNOR U11964 ( .A(n11703), .B(n11805), .Z(n11696) );
  XNOR U11965 ( .A(n11702), .B(n11700), .Z(n11805) );
  AND U11966 ( .A(n11806), .B(n11807), .Z(n11700) );
  NANDN U11967 ( .A(n11808), .B(n11809), .Z(n11807) );
  NANDN U11968 ( .A(n11810), .B(n11811), .Z(n11809) );
  NANDN U11969 ( .A(n11811), .B(n11810), .Z(n11806) );
  ANDN U11970 ( .B(B[215]), .A(n35), .Z(n11702) );
  XNOR U11971 ( .A(n11710), .B(n11812), .Z(n11703) );
  XNOR U11972 ( .A(n11709), .B(n11707), .Z(n11812) );
  AND U11973 ( .A(n11813), .B(n11814), .Z(n11707) );
  NANDN U11974 ( .A(n11815), .B(n11816), .Z(n11814) );
  OR U11975 ( .A(n11817), .B(n11818), .Z(n11816) );
  NAND U11976 ( .A(n11818), .B(n11817), .Z(n11813) );
  ANDN U11977 ( .B(B[216]), .A(n36), .Z(n11709) );
  XNOR U11978 ( .A(n11717), .B(n11819), .Z(n11710) );
  XNOR U11979 ( .A(n11716), .B(n11714), .Z(n11819) );
  AND U11980 ( .A(n11820), .B(n11821), .Z(n11714) );
  NANDN U11981 ( .A(n11822), .B(n11823), .Z(n11821) );
  NANDN U11982 ( .A(n11824), .B(n11825), .Z(n11823) );
  NANDN U11983 ( .A(n11825), .B(n11824), .Z(n11820) );
  ANDN U11984 ( .B(B[217]), .A(n37), .Z(n11716) );
  XNOR U11985 ( .A(n11724), .B(n11826), .Z(n11717) );
  XNOR U11986 ( .A(n11723), .B(n11721), .Z(n11826) );
  AND U11987 ( .A(n11827), .B(n11828), .Z(n11721) );
  NANDN U11988 ( .A(n11829), .B(n11830), .Z(n11828) );
  OR U11989 ( .A(n11831), .B(n11832), .Z(n11830) );
  NAND U11990 ( .A(n11832), .B(n11831), .Z(n11827) );
  ANDN U11991 ( .B(B[218]), .A(n38), .Z(n11723) );
  XNOR U11992 ( .A(n11731), .B(n11833), .Z(n11724) );
  XNOR U11993 ( .A(n11730), .B(n11728), .Z(n11833) );
  AND U11994 ( .A(n11834), .B(n11835), .Z(n11728) );
  NANDN U11995 ( .A(n11836), .B(n11837), .Z(n11835) );
  NANDN U11996 ( .A(n11838), .B(n11839), .Z(n11837) );
  NANDN U11997 ( .A(n11839), .B(n11838), .Z(n11834) );
  ANDN U11998 ( .B(B[219]), .A(n39), .Z(n11730) );
  XNOR U11999 ( .A(n11738), .B(n11840), .Z(n11731) );
  XNOR U12000 ( .A(n11737), .B(n11735), .Z(n11840) );
  AND U12001 ( .A(n11841), .B(n11842), .Z(n11735) );
  NANDN U12002 ( .A(n11843), .B(n11844), .Z(n11842) );
  OR U12003 ( .A(n11845), .B(n11846), .Z(n11844) );
  NAND U12004 ( .A(n11846), .B(n11845), .Z(n11841) );
  ANDN U12005 ( .B(B[220]), .A(n40), .Z(n11737) );
  XNOR U12006 ( .A(n11745), .B(n11847), .Z(n11738) );
  XNOR U12007 ( .A(n11744), .B(n11742), .Z(n11847) );
  AND U12008 ( .A(n11848), .B(n11849), .Z(n11742) );
  NANDN U12009 ( .A(n11850), .B(n11851), .Z(n11849) );
  NAND U12010 ( .A(n11852), .B(n11853), .Z(n11851) );
  ANDN U12011 ( .B(B[221]), .A(n41), .Z(n11744) );
  XOR U12012 ( .A(n11751), .B(n11854), .Z(n11745) );
  XNOR U12013 ( .A(n11749), .B(n11752), .Z(n11854) );
  NAND U12014 ( .A(A[2]), .B(B[222]), .Z(n11752) );
  NANDN U12015 ( .A(n11855), .B(n11856), .Z(n11749) );
  AND U12016 ( .A(A[0]), .B(B[223]), .Z(n11856) );
  XNOR U12017 ( .A(n11754), .B(n11857), .Z(n11751) );
  NAND U12018 ( .A(A[0]), .B(B[224]), .Z(n11857) );
  NAND U12019 ( .A(B[223]), .B(A[1]), .Z(n11754) );
  NAND U12020 ( .A(n11858), .B(n11859), .Z(n293) );
  NANDN U12021 ( .A(n11860), .B(n11861), .Z(n11859) );
  OR U12022 ( .A(n11862), .B(n11863), .Z(n11861) );
  NAND U12023 ( .A(n11863), .B(n11862), .Z(n11858) );
  XOR U12024 ( .A(n295), .B(n294), .Z(\A1[221] ) );
  XOR U12025 ( .A(n11863), .B(n11864), .Z(n294) );
  XNOR U12026 ( .A(n11862), .B(n11860), .Z(n11864) );
  AND U12027 ( .A(n11865), .B(n11866), .Z(n11860) );
  NANDN U12028 ( .A(n11867), .B(n11868), .Z(n11866) );
  NANDN U12029 ( .A(n11869), .B(n11870), .Z(n11868) );
  NANDN U12030 ( .A(n11870), .B(n11869), .Z(n11865) );
  ANDN U12031 ( .B(B[208]), .A(n29), .Z(n11862) );
  XNOR U12032 ( .A(n11769), .B(n11871), .Z(n11863) );
  XNOR U12033 ( .A(n11768), .B(n11766), .Z(n11871) );
  AND U12034 ( .A(n11872), .B(n11873), .Z(n11766) );
  NANDN U12035 ( .A(n11874), .B(n11875), .Z(n11873) );
  OR U12036 ( .A(n11876), .B(n11877), .Z(n11875) );
  NAND U12037 ( .A(n11877), .B(n11876), .Z(n11872) );
  ANDN U12038 ( .B(B[209]), .A(n30), .Z(n11768) );
  XNOR U12039 ( .A(n11776), .B(n11878), .Z(n11769) );
  XNOR U12040 ( .A(n11775), .B(n11773), .Z(n11878) );
  AND U12041 ( .A(n11879), .B(n11880), .Z(n11773) );
  NANDN U12042 ( .A(n11881), .B(n11882), .Z(n11880) );
  NANDN U12043 ( .A(n11883), .B(n11884), .Z(n11882) );
  NANDN U12044 ( .A(n11884), .B(n11883), .Z(n11879) );
  ANDN U12045 ( .B(B[210]), .A(n31), .Z(n11775) );
  XNOR U12046 ( .A(n11783), .B(n11885), .Z(n11776) );
  XNOR U12047 ( .A(n11782), .B(n11780), .Z(n11885) );
  AND U12048 ( .A(n11886), .B(n11887), .Z(n11780) );
  NANDN U12049 ( .A(n11888), .B(n11889), .Z(n11887) );
  OR U12050 ( .A(n11890), .B(n11891), .Z(n11889) );
  NAND U12051 ( .A(n11891), .B(n11890), .Z(n11886) );
  ANDN U12052 ( .B(B[211]), .A(n32), .Z(n11782) );
  XNOR U12053 ( .A(n11790), .B(n11892), .Z(n11783) );
  XNOR U12054 ( .A(n11789), .B(n11787), .Z(n11892) );
  AND U12055 ( .A(n11893), .B(n11894), .Z(n11787) );
  NANDN U12056 ( .A(n11895), .B(n11896), .Z(n11894) );
  NANDN U12057 ( .A(n11897), .B(n11898), .Z(n11896) );
  NANDN U12058 ( .A(n11898), .B(n11897), .Z(n11893) );
  ANDN U12059 ( .B(B[212]), .A(n33), .Z(n11789) );
  XNOR U12060 ( .A(n11797), .B(n11899), .Z(n11790) );
  XNOR U12061 ( .A(n11796), .B(n11794), .Z(n11899) );
  AND U12062 ( .A(n11900), .B(n11901), .Z(n11794) );
  NANDN U12063 ( .A(n11902), .B(n11903), .Z(n11901) );
  OR U12064 ( .A(n11904), .B(n11905), .Z(n11903) );
  NAND U12065 ( .A(n11905), .B(n11904), .Z(n11900) );
  ANDN U12066 ( .B(B[213]), .A(n34), .Z(n11796) );
  XNOR U12067 ( .A(n11804), .B(n11906), .Z(n11797) );
  XNOR U12068 ( .A(n11803), .B(n11801), .Z(n11906) );
  AND U12069 ( .A(n11907), .B(n11908), .Z(n11801) );
  NANDN U12070 ( .A(n11909), .B(n11910), .Z(n11908) );
  NANDN U12071 ( .A(n11911), .B(n11912), .Z(n11910) );
  NANDN U12072 ( .A(n11912), .B(n11911), .Z(n11907) );
  ANDN U12073 ( .B(B[214]), .A(n35), .Z(n11803) );
  XNOR U12074 ( .A(n11811), .B(n11913), .Z(n11804) );
  XNOR U12075 ( .A(n11810), .B(n11808), .Z(n11913) );
  AND U12076 ( .A(n11914), .B(n11915), .Z(n11808) );
  NANDN U12077 ( .A(n11916), .B(n11917), .Z(n11915) );
  OR U12078 ( .A(n11918), .B(n11919), .Z(n11917) );
  NAND U12079 ( .A(n11919), .B(n11918), .Z(n11914) );
  ANDN U12080 ( .B(B[215]), .A(n36), .Z(n11810) );
  XNOR U12081 ( .A(n11818), .B(n11920), .Z(n11811) );
  XNOR U12082 ( .A(n11817), .B(n11815), .Z(n11920) );
  AND U12083 ( .A(n11921), .B(n11922), .Z(n11815) );
  NANDN U12084 ( .A(n11923), .B(n11924), .Z(n11922) );
  NANDN U12085 ( .A(n11925), .B(n11926), .Z(n11924) );
  NANDN U12086 ( .A(n11926), .B(n11925), .Z(n11921) );
  ANDN U12087 ( .B(B[216]), .A(n37), .Z(n11817) );
  XNOR U12088 ( .A(n11825), .B(n11927), .Z(n11818) );
  XNOR U12089 ( .A(n11824), .B(n11822), .Z(n11927) );
  AND U12090 ( .A(n11928), .B(n11929), .Z(n11822) );
  NANDN U12091 ( .A(n11930), .B(n11931), .Z(n11929) );
  OR U12092 ( .A(n11932), .B(n11933), .Z(n11931) );
  NAND U12093 ( .A(n11933), .B(n11932), .Z(n11928) );
  ANDN U12094 ( .B(B[217]), .A(n38), .Z(n11824) );
  XNOR U12095 ( .A(n11832), .B(n11934), .Z(n11825) );
  XNOR U12096 ( .A(n11831), .B(n11829), .Z(n11934) );
  AND U12097 ( .A(n11935), .B(n11936), .Z(n11829) );
  NANDN U12098 ( .A(n11937), .B(n11938), .Z(n11936) );
  NANDN U12099 ( .A(n11939), .B(n11940), .Z(n11938) );
  NANDN U12100 ( .A(n11940), .B(n11939), .Z(n11935) );
  ANDN U12101 ( .B(B[218]), .A(n39), .Z(n11831) );
  XNOR U12102 ( .A(n11839), .B(n11941), .Z(n11832) );
  XNOR U12103 ( .A(n11838), .B(n11836), .Z(n11941) );
  AND U12104 ( .A(n11942), .B(n11943), .Z(n11836) );
  NANDN U12105 ( .A(n11944), .B(n11945), .Z(n11943) );
  OR U12106 ( .A(n11946), .B(n11947), .Z(n11945) );
  NAND U12107 ( .A(n11947), .B(n11946), .Z(n11942) );
  ANDN U12108 ( .B(B[219]), .A(n40), .Z(n11838) );
  XNOR U12109 ( .A(n11846), .B(n11948), .Z(n11839) );
  XNOR U12110 ( .A(n11845), .B(n11843), .Z(n11948) );
  AND U12111 ( .A(n11949), .B(n11950), .Z(n11843) );
  NANDN U12112 ( .A(n11951), .B(n11952), .Z(n11950) );
  NAND U12113 ( .A(n11953), .B(n11954), .Z(n11952) );
  ANDN U12114 ( .B(B[220]), .A(n41), .Z(n11845) );
  XOR U12115 ( .A(n11852), .B(n11955), .Z(n11846) );
  XNOR U12116 ( .A(n11850), .B(n11853), .Z(n11955) );
  NAND U12117 ( .A(A[2]), .B(B[221]), .Z(n11853) );
  NANDN U12118 ( .A(n11956), .B(n11957), .Z(n11850) );
  AND U12119 ( .A(A[0]), .B(B[222]), .Z(n11957) );
  XNOR U12120 ( .A(n11855), .B(n11958), .Z(n11852) );
  NAND U12121 ( .A(A[0]), .B(B[223]), .Z(n11958) );
  NAND U12122 ( .A(B[222]), .B(A[1]), .Z(n11855) );
  NAND U12123 ( .A(n11959), .B(n11960), .Z(n295) );
  NANDN U12124 ( .A(n11961), .B(n11962), .Z(n11960) );
  OR U12125 ( .A(n11963), .B(n11964), .Z(n11962) );
  NAND U12126 ( .A(n11964), .B(n11963), .Z(n11959) );
  XOR U12127 ( .A(n297), .B(n296), .Z(\A1[220] ) );
  XOR U12128 ( .A(n11964), .B(n11965), .Z(n296) );
  XNOR U12129 ( .A(n11963), .B(n11961), .Z(n11965) );
  AND U12130 ( .A(n11966), .B(n11967), .Z(n11961) );
  NANDN U12131 ( .A(n11968), .B(n11969), .Z(n11967) );
  NANDN U12132 ( .A(n11970), .B(n11971), .Z(n11969) );
  NANDN U12133 ( .A(n11971), .B(n11970), .Z(n11966) );
  ANDN U12134 ( .B(B[207]), .A(n29), .Z(n11963) );
  XNOR U12135 ( .A(n11870), .B(n11972), .Z(n11964) );
  XNOR U12136 ( .A(n11869), .B(n11867), .Z(n11972) );
  AND U12137 ( .A(n11973), .B(n11974), .Z(n11867) );
  NANDN U12138 ( .A(n11975), .B(n11976), .Z(n11974) );
  OR U12139 ( .A(n11977), .B(n11978), .Z(n11976) );
  NAND U12140 ( .A(n11978), .B(n11977), .Z(n11973) );
  ANDN U12141 ( .B(B[208]), .A(n30), .Z(n11869) );
  XNOR U12142 ( .A(n11877), .B(n11979), .Z(n11870) );
  XNOR U12143 ( .A(n11876), .B(n11874), .Z(n11979) );
  AND U12144 ( .A(n11980), .B(n11981), .Z(n11874) );
  NANDN U12145 ( .A(n11982), .B(n11983), .Z(n11981) );
  NANDN U12146 ( .A(n11984), .B(n11985), .Z(n11983) );
  NANDN U12147 ( .A(n11985), .B(n11984), .Z(n11980) );
  ANDN U12148 ( .B(B[209]), .A(n31), .Z(n11876) );
  XNOR U12149 ( .A(n11884), .B(n11986), .Z(n11877) );
  XNOR U12150 ( .A(n11883), .B(n11881), .Z(n11986) );
  AND U12151 ( .A(n11987), .B(n11988), .Z(n11881) );
  NANDN U12152 ( .A(n11989), .B(n11990), .Z(n11988) );
  OR U12153 ( .A(n11991), .B(n11992), .Z(n11990) );
  NAND U12154 ( .A(n11992), .B(n11991), .Z(n11987) );
  ANDN U12155 ( .B(B[210]), .A(n32), .Z(n11883) );
  XNOR U12156 ( .A(n11891), .B(n11993), .Z(n11884) );
  XNOR U12157 ( .A(n11890), .B(n11888), .Z(n11993) );
  AND U12158 ( .A(n11994), .B(n11995), .Z(n11888) );
  NANDN U12159 ( .A(n11996), .B(n11997), .Z(n11995) );
  NANDN U12160 ( .A(n11998), .B(n11999), .Z(n11997) );
  NANDN U12161 ( .A(n11999), .B(n11998), .Z(n11994) );
  ANDN U12162 ( .B(B[211]), .A(n33), .Z(n11890) );
  XNOR U12163 ( .A(n11898), .B(n12000), .Z(n11891) );
  XNOR U12164 ( .A(n11897), .B(n11895), .Z(n12000) );
  AND U12165 ( .A(n12001), .B(n12002), .Z(n11895) );
  NANDN U12166 ( .A(n12003), .B(n12004), .Z(n12002) );
  OR U12167 ( .A(n12005), .B(n12006), .Z(n12004) );
  NAND U12168 ( .A(n12006), .B(n12005), .Z(n12001) );
  ANDN U12169 ( .B(B[212]), .A(n34), .Z(n11897) );
  XNOR U12170 ( .A(n11905), .B(n12007), .Z(n11898) );
  XNOR U12171 ( .A(n11904), .B(n11902), .Z(n12007) );
  AND U12172 ( .A(n12008), .B(n12009), .Z(n11902) );
  NANDN U12173 ( .A(n12010), .B(n12011), .Z(n12009) );
  NANDN U12174 ( .A(n12012), .B(n12013), .Z(n12011) );
  NANDN U12175 ( .A(n12013), .B(n12012), .Z(n12008) );
  ANDN U12176 ( .B(B[213]), .A(n35), .Z(n11904) );
  XNOR U12177 ( .A(n11912), .B(n12014), .Z(n11905) );
  XNOR U12178 ( .A(n11911), .B(n11909), .Z(n12014) );
  AND U12179 ( .A(n12015), .B(n12016), .Z(n11909) );
  NANDN U12180 ( .A(n12017), .B(n12018), .Z(n12016) );
  OR U12181 ( .A(n12019), .B(n12020), .Z(n12018) );
  NAND U12182 ( .A(n12020), .B(n12019), .Z(n12015) );
  ANDN U12183 ( .B(B[214]), .A(n36), .Z(n11911) );
  XNOR U12184 ( .A(n11919), .B(n12021), .Z(n11912) );
  XNOR U12185 ( .A(n11918), .B(n11916), .Z(n12021) );
  AND U12186 ( .A(n12022), .B(n12023), .Z(n11916) );
  NANDN U12187 ( .A(n12024), .B(n12025), .Z(n12023) );
  NANDN U12188 ( .A(n12026), .B(n12027), .Z(n12025) );
  NANDN U12189 ( .A(n12027), .B(n12026), .Z(n12022) );
  ANDN U12190 ( .B(B[215]), .A(n37), .Z(n11918) );
  XNOR U12191 ( .A(n11926), .B(n12028), .Z(n11919) );
  XNOR U12192 ( .A(n11925), .B(n11923), .Z(n12028) );
  AND U12193 ( .A(n12029), .B(n12030), .Z(n11923) );
  NANDN U12194 ( .A(n12031), .B(n12032), .Z(n12030) );
  OR U12195 ( .A(n12033), .B(n12034), .Z(n12032) );
  NAND U12196 ( .A(n12034), .B(n12033), .Z(n12029) );
  ANDN U12197 ( .B(B[216]), .A(n38), .Z(n11925) );
  XNOR U12198 ( .A(n11933), .B(n12035), .Z(n11926) );
  XNOR U12199 ( .A(n11932), .B(n11930), .Z(n12035) );
  AND U12200 ( .A(n12036), .B(n12037), .Z(n11930) );
  NANDN U12201 ( .A(n12038), .B(n12039), .Z(n12037) );
  NANDN U12202 ( .A(n12040), .B(n12041), .Z(n12039) );
  NANDN U12203 ( .A(n12041), .B(n12040), .Z(n12036) );
  ANDN U12204 ( .B(B[217]), .A(n39), .Z(n11932) );
  XNOR U12205 ( .A(n11940), .B(n12042), .Z(n11933) );
  XNOR U12206 ( .A(n11939), .B(n11937), .Z(n12042) );
  AND U12207 ( .A(n12043), .B(n12044), .Z(n11937) );
  NANDN U12208 ( .A(n12045), .B(n12046), .Z(n12044) );
  OR U12209 ( .A(n12047), .B(n12048), .Z(n12046) );
  NAND U12210 ( .A(n12048), .B(n12047), .Z(n12043) );
  ANDN U12211 ( .B(B[218]), .A(n40), .Z(n11939) );
  XNOR U12212 ( .A(n11947), .B(n12049), .Z(n11940) );
  XNOR U12213 ( .A(n11946), .B(n11944), .Z(n12049) );
  AND U12214 ( .A(n12050), .B(n12051), .Z(n11944) );
  NANDN U12215 ( .A(n12052), .B(n12053), .Z(n12051) );
  NAND U12216 ( .A(n12054), .B(n12055), .Z(n12053) );
  ANDN U12217 ( .B(B[219]), .A(n41), .Z(n11946) );
  XOR U12218 ( .A(n11953), .B(n12056), .Z(n11947) );
  XNOR U12219 ( .A(n11951), .B(n11954), .Z(n12056) );
  NAND U12220 ( .A(A[2]), .B(B[220]), .Z(n11954) );
  NANDN U12221 ( .A(n12057), .B(n12058), .Z(n11951) );
  AND U12222 ( .A(A[0]), .B(B[221]), .Z(n12058) );
  XNOR U12223 ( .A(n11956), .B(n12059), .Z(n11953) );
  NAND U12224 ( .A(A[0]), .B(B[222]), .Z(n12059) );
  NAND U12225 ( .A(B[221]), .B(A[1]), .Z(n11956) );
  NAND U12226 ( .A(n12060), .B(n12061), .Z(n297) );
  NANDN U12227 ( .A(n12062), .B(n12063), .Z(n12061) );
  OR U12228 ( .A(n12064), .B(n12065), .Z(n12063) );
  NAND U12229 ( .A(n12065), .B(n12064), .Z(n12060) );
  XOR U12230 ( .A(n279), .B(n278), .Z(\A1[21] ) );
  XOR U12231 ( .A(n11055), .B(n12066), .Z(n278) );
  XNOR U12232 ( .A(n11054), .B(n11052), .Z(n12066) );
  AND U12233 ( .A(n12067), .B(n12068), .Z(n11052) );
  NANDN U12234 ( .A(n12069), .B(n12070), .Z(n12068) );
  NANDN U12235 ( .A(n12071), .B(n12072), .Z(n12070) );
  NANDN U12236 ( .A(n12072), .B(n12071), .Z(n12067) );
  ANDN U12237 ( .B(B[8]), .A(n29), .Z(n11054) );
  XNOR U12238 ( .A(n10961), .B(n12073), .Z(n11055) );
  XNOR U12239 ( .A(n10960), .B(n10958), .Z(n12073) );
  AND U12240 ( .A(n12074), .B(n12075), .Z(n10958) );
  NANDN U12241 ( .A(n12076), .B(n12077), .Z(n12075) );
  OR U12242 ( .A(n12078), .B(n12079), .Z(n12077) );
  NAND U12243 ( .A(n12079), .B(n12078), .Z(n12074) );
  ANDN U12244 ( .B(B[9]), .A(n30), .Z(n10960) );
  XNOR U12245 ( .A(n10968), .B(n12080), .Z(n10961) );
  XNOR U12246 ( .A(n10967), .B(n10965), .Z(n12080) );
  AND U12247 ( .A(n12081), .B(n12082), .Z(n10965) );
  NANDN U12248 ( .A(n12083), .B(n12084), .Z(n12082) );
  NANDN U12249 ( .A(n12085), .B(n12086), .Z(n12084) );
  NANDN U12250 ( .A(n12086), .B(n12085), .Z(n12081) );
  ANDN U12251 ( .B(B[10]), .A(n31), .Z(n10967) );
  XNOR U12252 ( .A(n10975), .B(n12087), .Z(n10968) );
  XNOR U12253 ( .A(n10974), .B(n10972), .Z(n12087) );
  AND U12254 ( .A(n12088), .B(n12089), .Z(n10972) );
  NANDN U12255 ( .A(n12090), .B(n12091), .Z(n12089) );
  OR U12256 ( .A(n12092), .B(n12093), .Z(n12091) );
  NAND U12257 ( .A(n12093), .B(n12092), .Z(n12088) );
  ANDN U12258 ( .B(B[11]), .A(n32), .Z(n10974) );
  XNOR U12259 ( .A(n10982), .B(n12094), .Z(n10975) );
  XNOR U12260 ( .A(n10981), .B(n10979), .Z(n12094) );
  AND U12261 ( .A(n12095), .B(n12096), .Z(n10979) );
  NANDN U12262 ( .A(n12097), .B(n12098), .Z(n12096) );
  NANDN U12263 ( .A(n12099), .B(n12100), .Z(n12098) );
  NANDN U12264 ( .A(n12100), .B(n12099), .Z(n12095) );
  ANDN U12265 ( .B(B[12]), .A(n33), .Z(n10981) );
  XNOR U12266 ( .A(n10989), .B(n12101), .Z(n10982) );
  XNOR U12267 ( .A(n10988), .B(n10986), .Z(n12101) );
  AND U12268 ( .A(n12102), .B(n12103), .Z(n10986) );
  NANDN U12269 ( .A(n12104), .B(n12105), .Z(n12103) );
  OR U12270 ( .A(n12106), .B(n12107), .Z(n12105) );
  NAND U12271 ( .A(n12107), .B(n12106), .Z(n12102) );
  ANDN U12272 ( .B(B[13]), .A(n34), .Z(n10988) );
  XNOR U12273 ( .A(n10996), .B(n12108), .Z(n10989) );
  XNOR U12274 ( .A(n10995), .B(n10993), .Z(n12108) );
  AND U12275 ( .A(n12109), .B(n12110), .Z(n10993) );
  NANDN U12276 ( .A(n12111), .B(n12112), .Z(n12110) );
  NANDN U12277 ( .A(n12113), .B(n12114), .Z(n12112) );
  NANDN U12278 ( .A(n12114), .B(n12113), .Z(n12109) );
  ANDN U12279 ( .B(B[14]), .A(n35), .Z(n10995) );
  XNOR U12280 ( .A(n11003), .B(n12115), .Z(n10996) );
  XNOR U12281 ( .A(n11002), .B(n11000), .Z(n12115) );
  AND U12282 ( .A(n12116), .B(n12117), .Z(n11000) );
  NANDN U12283 ( .A(n12118), .B(n12119), .Z(n12117) );
  OR U12284 ( .A(n12120), .B(n12121), .Z(n12119) );
  NAND U12285 ( .A(n12121), .B(n12120), .Z(n12116) );
  ANDN U12286 ( .B(B[15]), .A(n36), .Z(n11002) );
  XNOR U12287 ( .A(n11010), .B(n12122), .Z(n11003) );
  XNOR U12288 ( .A(n11009), .B(n11007), .Z(n12122) );
  AND U12289 ( .A(n12123), .B(n12124), .Z(n11007) );
  NANDN U12290 ( .A(n12125), .B(n12126), .Z(n12124) );
  NANDN U12291 ( .A(n12127), .B(n12128), .Z(n12126) );
  NANDN U12292 ( .A(n12128), .B(n12127), .Z(n12123) );
  ANDN U12293 ( .B(B[16]), .A(n37), .Z(n11009) );
  XNOR U12294 ( .A(n11017), .B(n12129), .Z(n11010) );
  XNOR U12295 ( .A(n11016), .B(n11014), .Z(n12129) );
  AND U12296 ( .A(n12130), .B(n12131), .Z(n11014) );
  NANDN U12297 ( .A(n12132), .B(n12133), .Z(n12131) );
  OR U12298 ( .A(n12134), .B(n12135), .Z(n12133) );
  NAND U12299 ( .A(n12135), .B(n12134), .Z(n12130) );
  ANDN U12300 ( .B(B[17]), .A(n38), .Z(n11016) );
  XNOR U12301 ( .A(n11024), .B(n12136), .Z(n11017) );
  XNOR U12302 ( .A(n11023), .B(n11021), .Z(n12136) );
  AND U12303 ( .A(n12137), .B(n12138), .Z(n11021) );
  NANDN U12304 ( .A(n12139), .B(n12140), .Z(n12138) );
  NANDN U12305 ( .A(n12141), .B(n12142), .Z(n12140) );
  NANDN U12306 ( .A(n12142), .B(n12141), .Z(n12137) );
  ANDN U12307 ( .B(B[18]), .A(n39), .Z(n11023) );
  XNOR U12308 ( .A(n11031), .B(n12143), .Z(n11024) );
  XNOR U12309 ( .A(n11030), .B(n11028), .Z(n12143) );
  AND U12310 ( .A(n12144), .B(n12145), .Z(n11028) );
  NANDN U12311 ( .A(n12146), .B(n12147), .Z(n12145) );
  OR U12312 ( .A(n12148), .B(n12149), .Z(n12147) );
  NAND U12313 ( .A(n12149), .B(n12148), .Z(n12144) );
  ANDN U12314 ( .B(B[19]), .A(n40), .Z(n11030) );
  XNOR U12315 ( .A(n11038), .B(n12150), .Z(n11031) );
  XNOR U12316 ( .A(n11037), .B(n11035), .Z(n12150) );
  AND U12317 ( .A(n12151), .B(n12152), .Z(n11035) );
  NANDN U12318 ( .A(n12153), .B(n12154), .Z(n12152) );
  NAND U12319 ( .A(n12155), .B(n12156), .Z(n12154) );
  ANDN U12320 ( .B(B[20]), .A(n41), .Z(n11037) );
  XOR U12321 ( .A(n11044), .B(n12157), .Z(n11038) );
  XNOR U12322 ( .A(n11042), .B(n11045), .Z(n12157) );
  NAND U12323 ( .A(A[2]), .B(B[21]), .Z(n11045) );
  NANDN U12324 ( .A(n12158), .B(n12159), .Z(n11042) );
  AND U12325 ( .A(A[0]), .B(B[22]), .Z(n12159) );
  XNOR U12326 ( .A(n11047), .B(n12160), .Z(n11044) );
  NAND U12327 ( .A(A[0]), .B(B[23]), .Z(n12160) );
  NAND U12328 ( .A(B[22]), .B(A[1]), .Z(n11047) );
  NAND U12329 ( .A(n12161), .B(n12162), .Z(n279) );
  NANDN U12330 ( .A(n12163), .B(n12164), .Z(n12162) );
  OR U12331 ( .A(n12165), .B(n12166), .Z(n12164) );
  NAND U12332 ( .A(n12166), .B(n12165), .Z(n12161) );
  XOR U12333 ( .A(n299), .B(n298), .Z(\A1[219] ) );
  XOR U12334 ( .A(n12065), .B(n12167), .Z(n298) );
  XNOR U12335 ( .A(n12064), .B(n12062), .Z(n12167) );
  AND U12336 ( .A(n12168), .B(n12169), .Z(n12062) );
  NANDN U12337 ( .A(n12170), .B(n12171), .Z(n12169) );
  NANDN U12338 ( .A(n12172), .B(n12173), .Z(n12171) );
  NANDN U12339 ( .A(n12173), .B(n12172), .Z(n12168) );
  ANDN U12340 ( .B(B[206]), .A(n29), .Z(n12064) );
  XNOR U12341 ( .A(n11971), .B(n12174), .Z(n12065) );
  XNOR U12342 ( .A(n11970), .B(n11968), .Z(n12174) );
  AND U12343 ( .A(n12175), .B(n12176), .Z(n11968) );
  NANDN U12344 ( .A(n12177), .B(n12178), .Z(n12176) );
  OR U12345 ( .A(n12179), .B(n12180), .Z(n12178) );
  NAND U12346 ( .A(n12180), .B(n12179), .Z(n12175) );
  ANDN U12347 ( .B(B[207]), .A(n30), .Z(n11970) );
  XNOR U12348 ( .A(n11978), .B(n12181), .Z(n11971) );
  XNOR U12349 ( .A(n11977), .B(n11975), .Z(n12181) );
  AND U12350 ( .A(n12182), .B(n12183), .Z(n11975) );
  NANDN U12351 ( .A(n12184), .B(n12185), .Z(n12183) );
  NANDN U12352 ( .A(n12186), .B(n12187), .Z(n12185) );
  NANDN U12353 ( .A(n12187), .B(n12186), .Z(n12182) );
  ANDN U12354 ( .B(B[208]), .A(n31), .Z(n11977) );
  XNOR U12355 ( .A(n11985), .B(n12188), .Z(n11978) );
  XNOR U12356 ( .A(n11984), .B(n11982), .Z(n12188) );
  AND U12357 ( .A(n12189), .B(n12190), .Z(n11982) );
  NANDN U12358 ( .A(n12191), .B(n12192), .Z(n12190) );
  OR U12359 ( .A(n12193), .B(n12194), .Z(n12192) );
  NAND U12360 ( .A(n12194), .B(n12193), .Z(n12189) );
  ANDN U12361 ( .B(B[209]), .A(n32), .Z(n11984) );
  XNOR U12362 ( .A(n11992), .B(n12195), .Z(n11985) );
  XNOR U12363 ( .A(n11991), .B(n11989), .Z(n12195) );
  AND U12364 ( .A(n12196), .B(n12197), .Z(n11989) );
  NANDN U12365 ( .A(n12198), .B(n12199), .Z(n12197) );
  NANDN U12366 ( .A(n12200), .B(n12201), .Z(n12199) );
  NANDN U12367 ( .A(n12201), .B(n12200), .Z(n12196) );
  ANDN U12368 ( .B(B[210]), .A(n33), .Z(n11991) );
  XNOR U12369 ( .A(n11999), .B(n12202), .Z(n11992) );
  XNOR U12370 ( .A(n11998), .B(n11996), .Z(n12202) );
  AND U12371 ( .A(n12203), .B(n12204), .Z(n11996) );
  NANDN U12372 ( .A(n12205), .B(n12206), .Z(n12204) );
  OR U12373 ( .A(n12207), .B(n12208), .Z(n12206) );
  NAND U12374 ( .A(n12208), .B(n12207), .Z(n12203) );
  ANDN U12375 ( .B(B[211]), .A(n34), .Z(n11998) );
  XNOR U12376 ( .A(n12006), .B(n12209), .Z(n11999) );
  XNOR U12377 ( .A(n12005), .B(n12003), .Z(n12209) );
  AND U12378 ( .A(n12210), .B(n12211), .Z(n12003) );
  NANDN U12379 ( .A(n12212), .B(n12213), .Z(n12211) );
  NANDN U12380 ( .A(n12214), .B(n12215), .Z(n12213) );
  NANDN U12381 ( .A(n12215), .B(n12214), .Z(n12210) );
  ANDN U12382 ( .B(B[212]), .A(n35), .Z(n12005) );
  XNOR U12383 ( .A(n12013), .B(n12216), .Z(n12006) );
  XNOR U12384 ( .A(n12012), .B(n12010), .Z(n12216) );
  AND U12385 ( .A(n12217), .B(n12218), .Z(n12010) );
  NANDN U12386 ( .A(n12219), .B(n12220), .Z(n12218) );
  OR U12387 ( .A(n12221), .B(n12222), .Z(n12220) );
  NAND U12388 ( .A(n12222), .B(n12221), .Z(n12217) );
  ANDN U12389 ( .B(B[213]), .A(n36), .Z(n12012) );
  XNOR U12390 ( .A(n12020), .B(n12223), .Z(n12013) );
  XNOR U12391 ( .A(n12019), .B(n12017), .Z(n12223) );
  AND U12392 ( .A(n12224), .B(n12225), .Z(n12017) );
  NANDN U12393 ( .A(n12226), .B(n12227), .Z(n12225) );
  NANDN U12394 ( .A(n12228), .B(n12229), .Z(n12227) );
  NANDN U12395 ( .A(n12229), .B(n12228), .Z(n12224) );
  ANDN U12396 ( .B(B[214]), .A(n37), .Z(n12019) );
  XNOR U12397 ( .A(n12027), .B(n12230), .Z(n12020) );
  XNOR U12398 ( .A(n12026), .B(n12024), .Z(n12230) );
  AND U12399 ( .A(n12231), .B(n12232), .Z(n12024) );
  NANDN U12400 ( .A(n12233), .B(n12234), .Z(n12232) );
  OR U12401 ( .A(n12235), .B(n12236), .Z(n12234) );
  NAND U12402 ( .A(n12236), .B(n12235), .Z(n12231) );
  ANDN U12403 ( .B(B[215]), .A(n38), .Z(n12026) );
  XNOR U12404 ( .A(n12034), .B(n12237), .Z(n12027) );
  XNOR U12405 ( .A(n12033), .B(n12031), .Z(n12237) );
  AND U12406 ( .A(n12238), .B(n12239), .Z(n12031) );
  NANDN U12407 ( .A(n12240), .B(n12241), .Z(n12239) );
  NANDN U12408 ( .A(n12242), .B(n12243), .Z(n12241) );
  NANDN U12409 ( .A(n12243), .B(n12242), .Z(n12238) );
  ANDN U12410 ( .B(B[216]), .A(n39), .Z(n12033) );
  XNOR U12411 ( .A(n12041), .B(n12244), .Z(n12034) );
  XNOR U12412 ( .A(n12040), .B(n12038), .Z(n12244) );
  AND U12413 ( .A(n12245), .B(n12246), .Z(n12038) );
  NANDN U12414 ( .A(n12247), .B(n12248), .Z(n12246) );
  OR U12415 ( .A(n12249), .B(n12250), .Z(n12248) );
  NAND U12416 ( .A(n12250), .B(n12249), .Z(n12245) );
  ANDN U12417 ( .B(B[217]), .A(n40), .Z(n12040) );
  XNOR U12418 ( .A(n12048), .B(n12251), .Z(n12041) );
  XNOR U12419 ( .A(n12047), .B(n12045), .Z(n12251) );
  AND U12420 ( .A(n12252), .B(n12253), .Z(n12045) );
  NANDN U12421 ( .A(n12254), .B(n12255), .Z(n12253) );
  NAND U12422 ( .A(n12256), .B(n12257), .Z(n12255) );
  ANDN U12423 ( .B(B[218]), .A(n41), .Z(n12047) );
  XOR U12424 ( .A(n12054), .B(n12258), .Z(n12048) );
  XNOR U12425 ( .A(n12052), .B(n12055), .Z(n12258) );
  NAND U12426 ( .A(A[2]), .B(B[219]), .Z(n12055) );
  NANDN U12427 ( .A(n12259), .B(n12260), .Z(n12052) );
  AND U12428 ( .A(A[0]), .B(B[220]), .Z(n12260) );
  XNOR U12429 ( .A(n12057), .B(n12261), .Z(n12054) );
  NAND U12430 ( .A(A[0]), .B(B[221]), .Z(n12261) );
  NAND U12431 ( .A(B[220]), .B(A[1]), .Z(n12057) );
  NAND U12432 ( .A(n12262), .B(n12263), .Z(n299) );
  NANDN U12433 ( .A(n12264), .B(n12265), .Z(n12263) );
  OR U12434 ( .A(n12266), .B(n12267), .Z(n12265) );
  NAND U12435 ( .A(n12267), .B(n12266), .Z(n12262) );
  XOR U12436 ( .A(n303), .B(n302), .Z(\A1[218] ) );
  XOR U12437 ( .A(n12267), .B(n12268), .Z(n302) );
  XNOR U12438 ( .A(n12266), .B(n12264), .Z(n12268) );
  AND U12439 ( .A(n12269), .B(n12270), .Z(n12264) );
  NANDN U12440 ( .A(n12271), .B(n12272), .Z(n12270) );
  NANDN U12441 ( .A(n12273), .B(n12274), .Z(n12272) );
  NANDN U12442 ( .A(n12274), .B(n12273), .Z(n12269) );
  ANDN U12443 ( .B(B[205]), .A(n29), .Z(n12266) );
  XNOR U12444 ( .A(n12173), .B(n12275), .Z(n12267) );
  XNOR U12445 ( .A(n12172), .B(n12170), .Z(n12275) );
  AND U12446 ( .A(n12276), .B(n12277), .Z(n12170) );
  NANDN U12447 ( .A(n12278), .B(n12279), .Z(n12277) );
  OR U12448 ( .A(n12280), .B(n12281), .Z(n12279) );
  NAND U12449 ( .A(n12281), .B(n12280), .Z(n12276) );
  ANDN U12450 ( .B(B[206]), .A(n30), .Z(n12172) );
  XNOR U12451 ( .A(n12180), .B(n12282), .Z(n12173) );
  XNOR U12452 ( .A(n12179), .B(n12177), .Z(n12282) );
  AND U12453 ( .A(n12283), .B(n12284), .Z(n12177) );
  NANDN U12454 ( .A(n12285), .B(n12286), .Z(n12284) );
  NANDN U12455 ( .A(n12287), .B(n12288), .Z(n12286) );
  NANDN U12456 ( .A(n12288), .B(n12287), .Z(n12283) );
  ANDN U12457 ( .B(B[207]), .A(n31), .Z(n12179) );
  XNOR U12458 ( .A(n12187), .B(n12289), .Z(n12180) );
  XNOR U12459 ( .A(n12186), .B(n12184), .Z(n12289) );
  AND U12460 ( .A(n12290), .B(n12291), .Z(n12184) );
  NANDN U12461 ( .A(n12292), .B(n12293), .Z(n12291) );
  OR U12462 ( .A(n12294), .B(n12295), .Z(n12293) );
  NAND U12463 ( .A(n12295), .B(n12294), .Z(n12290) );
  ANDN U12464 ( .B(B[208]), .A(n32), .Z(n12186) );
  XNOR U12465 ( .A(n12194), .B(n12296), .Z(n12187) );
  XNOR U12466 ( .A(n12193), .B(n12191), .Z(n12296) );
  AND U12467 ( .A(n12297), .B(n12298), .Z(n12191) );
  NANDN U12468 ( .A(n12299), .B(n12300), .Z(n12298) );
  NANDN U12469 ( .A(n12301), .B(n12302), .Z(n12300) );
  NANDN U12470 ( .A(n12302), .B(n12301), .Z(n12297) );
  ANDN U12471 ( .B(B[209]), .A(n33), .Z(n12193) );
  XNOR U12472 ( .A(n12201), .B(n12303), .Z(n12194) );
  XNOR U12473 ( .A(n12200), .B(n12198), .Z(n12303) );
  AND U12474 ( .A(n12304), .B(n12305), .Z(n12198) );
  NANDN U12475 ( .A(n12306), .B(n12307), .Z(n12305) );
  OR U12476 ( .A(n12308), .B(n12309), .Z(n12307) );
  NAND U12477 ( .A(n12309), .B(n12308), .Z(n12304) );
  ANDN U12478 ( .B(B[210]), .A(n34), .Z(n12200) );
  XNOR U12479 ( .A(n12208), .B(n12310), .Z(n12201) );
  XNOR U12480 ( .A(n12207), .B(n12205), .Z(n12310) );
  AND U12481 ( .A(n12311), .B(n12312), .Z(n12205) );
  NANDN U12482 ( .A(n12313), .B(n12314), .Z(n12312) );
  NANDN U12483 ( .A(n12315), .B(n12316), .Z(n12314) );
  NANDN U12484 ( .A(n12316), .B(n12315), .Z(n12311) );
  ANDN U12485 ( .B(B[211]), .A(n35), .Z(n12207) );
  XNOR U12486 ( .A(n12215), .B(n12317), .Z(n12208) );
  XNOR U12487 ( .A(n12214), .B(n12212), .Z(n12317) );
  AND U12488 ( .A(n12318), .B(n12319), .Z(n12212) );
  NANDN U12489 ( .A(n12320), .B(n12321), .Z(n12319) );
  OR U12490 ( .A(n12322), .B(n12323), .Z(n12321) );
  NAND U12491 ( .A(n12323), .B(n12322), .Z(n12318) );
  ANDN U12492 ( .B(B[212]), .A(n36), .Z(n12214) );
  XNOR U12493 ( .A(n12222), .B(n12324), .Z(n12215) );
  XNOR U12494 ( .A(n12221), .B(n12219), .Z(n12324) );
  AND U12495 ( .A(n12325), .B(n12326), .Z(n12219) );
  NANDN U12496 ( .A(n12327), .B(n12328), .Z(n12326) );
  NANDN U12497 ( .A(n12329), .B(n12330), .Z(n12328) );
  NANDN U12498 ( .A(n12330), .B(n12329), .Z(n12325) );
  ANDN U12499 ( .B(B[213]), .A(n37), .Z(n12221) );
  XNOR U12500 ( .A(n12229), .B(n12331), .Z(n12222) );
  XNOR U12501 ( .A(n12228), .B(n12226), .Z(n12331) );
  AND U12502 ( .A(n12332), .B(n12333), .Z(n12226) );
  NANDN U12503 ( .A(n12334), .B(n12335), .Z(n12333) );
  OR U12504 ( .A(n12336), .B(n12337), .Z(n12335) );
  NAND U12505 ( .A(n12337), .B(n12336), .Z(n12332) );
  ANDN U12506 ( .B(B[214]), .A(n38), .Z(n12228) );
  XNOR U12507 ( .A(n12236), .B(n12338), .Z(n12229) );
  XNOR U12508 ( .A(n12235), .B(n12233), .Z(n12338) );
  AND U12509 ( .A(n12339), .B(n12340), .Z(n12233) );
  NANDN U12510 ( .A(n12341), .B(n12342), .Z(n12340) );
  NANDN U12511 ( .A(n12343), .B(n12344), .Z(n12342) );
  NANDN U12512 ( .A(n12344), .B(n12343), .Z(n12339) );
  ANDN U12513 ( .B(B[215]), .A(n39), .Z(n12235) );
  XNOR U12514 ( .A(n12243), .B(n12345), .Z(n12236) );
  XNOR U12515 ( .A(n12242), .B(n12240), .Z(n12345) );
  AND U12516 ( .A(n12346), .B(n12347), .Z(n12240) );
  NANDN U12517 ( .A(n12348), .B(n12349), .Z(n12347) );
  OR U12518 ( .A(n12350), .B(n12351), .Z(n12349) );
  NAND U12519 ( .A(n12351), .B(n12350), .Z(n12346) );
  ANDN U12520 ( .B(B[216]), .A(n40), .Z(n12242) );
  XNOR U12521 ( .A(n12250), .B(n12352), .Z(n12243) );
  XNOR U12522 ( .A(n12249), .B(n12247), .Z(n12352) );
  AND U12523 ( .A(n12353), .B(n12354), .Z(n12247) );
  NANDN U12524 ( .A(n12355), .B(n12356), .Z(n12354) );
  NAND U12525 ( .A(n12357), .B(n12358), .Z(n12356) );
  ANDN U12526 ( .B(B[217]), .A(n41), .Z(n12249) );
  XOR U12527 ( .A(n12256), .B(n12359), .Z(n12250) );
  XNOR U12528 ( .A(n12254), .B(n12257), .Z(n12359) );
  NAND U12529 ( .A(A[2]), .B(B[218]), .Z(n12257) );
  NANDN U12530 ( .A(n12360), .B(n12361), .Z(n12254) );
  AND U12531 ( .A(A[0]), .B(B[219]), .Z(n12361) );
  XNOR U12532 ( .A(n12259), .B(n12362), .Z(n12256) );
  NAND U12533 ( .A(A[0]), .B(B[220]), .Z(n12362) );
  NAND U12534 ( .A(B[219]), .B(A[1]), .Z(n12259) );
  NAND U12535 ( .A(n12363), .B(n12364), .Z(n303) );
  NANDN U12536 ( .A(n12365), .B(n12366), .Z(n12364) );
  OR U12537 ( .A(n12367), .B(n12368), .Z(n12366) );
  NAND U12538 ( .A(n12368), .B(n12367), .Z(n12363) );
  XOR U12539 ( .A(n305), .B(n304), .Z(\A1[217] ) );
  XOR U12540 ( .A(n12368), .B(n12369), .Z(n304) );
  XNOR U12541 ( .A(n12367), .B(n12365), .Z(n12369) );
  AND U12542 ( .A(n12370), .B(n12371), .Z(n12365) );
  NANDN U12543 ( .A(n12372), .B(n12373), .Z(n12371) );
  NANDN U12544 ( .A(n12374), .B(n12375), .Z(n12373) );
  NANDN U12545 ( .A(n12375), .B(n12374), .Z(n12370) );
  ANDN U12546 ( .B(B[204]), .A(n29), .Z(n12367) );
  XNOR U12547 ( .A(n12274), .B(n12376), .Z(n12368) );
  XNOR U12548 ( .A(n12273), .B(n12271), .Z(n12376) );
  AND U12549 ( .A(n12377), .B(n12378), .Z(n12271) );
  NANDN U12550 ( .A(n12379), .B(n12380), .Z(n12378) );
  OR U12551 ( .A(n12381), .B(n12382), .Z(n12380) );
  NAND U12552 ( .A(n12382), .B(n12381), .Z(n12377) );
  ANDN U12553 ( .B(B[205]), .A(n30), .Z(n12273) );
  XNOR U12554 ( .A(n12281), .B(n12383), .Z(n12274) );
  XNOR U12555 ( .A(n12280), .B(n12278), .Z(n12383) );
  AND U12556 ( .A(n12384), .B(n12385), .Z(n12278) );
  NANDN U12557 ( .A(n12386), .B(n12387), .Z(n12385) );
  NANDN U12558 ( .A(n12388), .B(n12389), .Z(n12387) );
  NANDN U12559 ( .A(n12389), .B(n12388), .Z(n12384) );
  ANDN U12560 ( .B(B[206]), .A(n31), .Z(n12280) );
  XNOR U12561 ( .A(n12288), .B(n12390), .Z(n12281) );
  XNOR U12562 ( .A(n12287), .B(n12285), .Z(n12390) );
  AND U12563 ( .A(n12391), .B(n12392), .Z(n12285) );
  NANDN U12564 ( .A(n12393), .B(n12394), .Z(n12392) );
  OR U12565 ( .A(n12395), .B(n12396), .Z(n12394) );
  NAND U12566 ( .A(n12396), .B(n12395), .Z(n12391) );
  ANDN U12567 ( .B(B[207]), .A(n32), .Z(n12287) );
  XNOR U12568 ( .A(n12295), .B(n12397), .Z(n12288) );
  XNOR U12569 ( .A(n12294), .B(n12292), .Z(n12397) );
  AND U12570 ( .A(n12398), .B(n12399), .Z(n12292) );
  NANDN U12571 ( .A(n12400), .B(n12401), .Z(n12399) );
  NANDN U12572 ( .A(n12402), .B(n12403), .Z(n12401) );
  NANDN U12573 ( .A(n12403), .B(n12402), .Z(n12398) );
  ANDN U12574 ( .B(B[208]), .A(n33), .Z(n12294) );
  XNOR U12575 ( .A(n12302), .B(n12404), .Z(n12295) );
  XNOR U12576 ( .A(n12301), .B(n12299), .Z(n12404) );
  AND U12577 ( .A(n12405), .B(n12406), .Z(n12299) );
  NANDN U12578 ( .A(n12407), .B(n12408), .Z(n12406) );
  OR U12579 ( .A(n12409), .B(n12410), .Z(n12408) );
  NAND U12580 ( .A(n12410), .B(n12409), .Z(n12405) );
  ANDN U12581 ( .B(B[209]), .A(n34), .Z(n12301) );
  XNOR U12582 ( .A(n12309), .B(n12411), .Z(n12302) );
  XNOR U12583 ( .A(n12308), .B(n12306), .Z(n12411) );
  AND U12584 ( .A(n12412), .B(n12413), .Z(n12306) );
  NANDN U12585 ( .A(n12414), .B(n12415), .Z(n12413) );
  NANDN U12586 ( .A(n12416), .B(n12417), .Z(n12415) );
  NANDN U12587 ( .A(n12417), .B(n12416), .Z(n12412) );
  ANDN U12588 ( .B(B[210]), .A(n35), .Z(n12308) );
  XNOR U12589 ( .A(n12316), .B(n12418), .Z(n12309) );
  XNOR U12590 ( .A(n12315), .B(n12313), .Z(n12418) );
  AND U12591 ( .A(n12419), .B(n12420), .Z(n12313) );
  NANDN U12592 ( .A(n12421), .B(n12422), .Z(n12420) );
  OR U12593 ( .A(n12423), .B(n12424), .Z(n12422) );
  NAND U12594 ( .A(n12424), .B(n12423), .Z(n12419) );
  ANDN U12595 ( .B(B[211]), .A(n36), .Z(n12315) );
  XNOR U12596 ( .A(n12323), .B(n12425), .Z(n12316) );
  XNOR U12597 ( .A(n12322), .B(n12320), .Z(n12425) );
  AND U12598 ( .A(n12426), .B(n12427), .Z(n12320) );
  NANDN U12599 ( .A(n12428), .B(n12429), .Z(n12427) );
  NANDN U12600 ( .A(n12430), .B(n12431), .Z(n12429) );
  NANDN U12601 ( .A(n12431), .B(n12430), .Z(n12426) );
  ANDN U12602 ( .B(B[212]), .A(n37), .Z(n12322) );
  XNOR U12603 ( .A(n12330), .B(n12432), .Z(n12323) );
  XNOR U12604 ( .A(n12329), .B(n12327), .Z(n12432) );
  AND U12605 ( .A(n12433), .B(n12434), .Z(n12327) );
  NANDN U12606 ( .A(n12435), .B(n12436), .Z(n12434) );
  OR U12607 ( .A(n12437), .B(n12438), .Z(n12436) );
  NAND U12608 ( .A(n12438), .B(n12437), .Z(n12433) );
  ANDN U12609 ( .B(B[213]), .A(n38), .Z(n12329) );
  XNOR U12610 ( .A(n12337), .B(n12439), .Z(n12330) );
  XNOR U12611 ( .A(n12336), .B(n12334), .Z(n12439) );
  AND U12612 ( .A(n12440), .B(n12441), .Z(n12334) );
  NANDN U12613 ( .A(n12442), .B(n12443), .Z(n12441) );
  NANDN U12614 ( .A(n12444), .B(n12445), .Z(n12443) );
  NANDN U12615 ( .A(n12445), .B(n12444), .Z(n12440) );
  ANDN U12616 ( .B(B[214]), .A(n39), .Z(n12336) );
  XNOR U12617 ( .A(n12344), .B(n12446), .Z(n12337) );
  XNOR U12618 ( .A(n12343), .B(n12341), .Z(n12446) );
  AND U12619 ( .A(n12447), .B(n12448), .Z(n12341) );
  NANDN U12620 ( .A(n12449), .B(n12450), .Z(n12448) );
  OR U12621 ( .A(n12451), .B(n12452), .Z(n12450) );
  NAND U12622 ( .A(n12452), .B(n12451), .Z(n12447) );
  ANDN U12623 ( .B(B[215]), .A(n40), .Z(n12343) );
  XNOR U12624 ( .A(n12351), .B(n12453), .Z(n12344) );
  XNOR U12625 ( .A(n12350), .B(n12348), .Z(n12453) );
  AND U12626 ( .A(n12454), .B(n12455), .Z(n12348) );
  NANDN U12627 ( .A(n12456), .B(n12457), .Z(n12455) );
  NAND U12628 ( .A(n12458), .B(n12459), .Z(n12457) );
  ANDN U12629 ( .B(B[216]), .A(n41), .Z(n12350) );
  XOR U12630 ( .A(n12357), .B(n12460), .Z(n12351) );
  XNOR U12631 ( .A(n12355), .B(n12358), .Z(n12460) );
  NAND U12632 ( .A(A[2]), .B(B[217]), .Z(n12358) );
  NANDN U12633 ( .A(n12461), .B(n12462), .Z(n12355) );
  AND U12634 ( .A(A[0]), .B(B[218]), .Z(n12462) );
  XNOR U12635 ( .A(n12360), .B(n12463), .Z(n12357) );
  NAND U12636 ( .A(A[0]), .B(B[219]), .Z(n12463) );
  NAND U12637 ( .A(B[218]), .B(A[1]), .Z(n12360) );
  NAND U12638 ( .A(n12464), .B(n12465), .Z(n305) );
  NANDN U12639 ( .A(n12466), .B(n12467), .Z(n12465) );
  OR U12640 ( .A(n12468), .B(n12469), .Z(n12467) );
  NAND U12641 ( .A(n12469), .B(n12468), .Z(n12464) );
  XOR U12642 ( .A(n307), .B(n306), .Z(\A1[216] ) );
  XOR U12643 ( .A(n12469), .B(n12470), .Z(n306) );
  XNOR U12644 ( .A(n12468), .B(n12466), .Z(n12470) );
  AND U12645 ( .A(n12471), .B(n12472), .Z(n12466) );
  NANDN U12646 ( .A(n12473), .B(n12474), .Z(n12472) );
  NANDN U12647 ( .A(n12475), .B(n12476), .Z(n12474) );
  NANDN U12648 ( .A(n12476), .B(n12475), .Z(n12471) );
  ANDN U12649 ( .B(B[203]), .A(n29), .Z(n12468) );
  XNOR U12650 ( .A(n12375), .B(n12477), .Z(n12469) );
  XNOR U12651 ( .A(n12374), .B(n12372), .Z(n12477) );
  AND U12652 ( .A(n12478), .B(n12479), .Z(n12372) );
  NANDN U12653 ( .A(n12480), .B(n12481), .Z(n12479) );
  OR U12654 ( .A(n12482), .B(n12483), .Z(n12481) );
  NAND U12655 ( .A(n12483), .B(n12482), .Z(n12478) );
  ANDN U12656 ( .B(B[204]), .A(n30), .Z(n12374) );
  XNOR U12657 ( .A(n12382), .B(n12484), .Z(n12375) );
  XNOR U12658 ( .A(n12381), .B(n12379), .Z(n12484) );
  AND U12659 ( .A(n12485), .B(n12486), .Z(n12379) );
  NANDN U12660 ( .A(n12487), .B(n12488), .Z(n12486) );
  NANDN U12661 ( .A(n12489), .B(n12490), .Z(n12488) );
  NANDN U12662 ( .A(n12490), .B(n12489), .Z(n12485) );
  ANDN U12663 ( .B(B[205]), .A(n31), .Z(n12381) );
  XNOR U12664 ( .A(n12389), .B(n12491), .Z(n12382) );
  XNOR U12665 ( .A(n12388), .B(n12386), .Z(n12491) );
  AND U12666 ( .A(n12492), .B(n12493), .Z(n12386) );
  NANDN U12667 ( .A(n12494), .B(n12495), .Z(n12493) );
  OR U12668 ( .A(n12496), .B(n12497), .Z(n12495) );
  NAND U12669 ( .A(n12497), .B(n12496), .Z(n12492) );
  ANDN U12670 ( .B(B[206]), .A(n32), .Z(n12388) );
  XNOR U12671 ( .A(n12396), .B(n12498), .Z(n12389) );
  XNOR U12672 ( .A(n12395), .B(n12393), .Z(n12498) );
  AND U12673 ( .A(n12499), .B(n12500), .Z(n12393) );
  NANDN U12674 ( .A(n12501), .B(n12502), .Z(n12500) );
  NANDN U12675 ( .A(n12503), .B(n12504), .Z(n12502) );
  NANDN U12676 ( .A(n12504), .B(n12503), .Z(n12499) );
  ANDN U12677 ( .B(B[207]), .A(n33), .Z(n12395) );
  XNOR U12678 ( .A(n12403), .B(n12505), .Z(n12396) );
  XNOR U12679 ( .A(n12402), .B(n12400), .Z(n12505) );
  AND U12680 ( .A(n12506), .B(n12507), .Z(n12400) );
  NANDN U12681 ( .A(n12508), .B(n12509), .Z(n12507) );
  OR U12682 ( .A(n12510), .B(n12511), .Z(n12509) );
  NAND U12683 ( .A(n12511), .B(n12510), .Z(n12506) );
  ANDN U12684 ( .B(B[208]), .A(n34), .Z(n12402) );
  XNOR U12685 ( .A(n12410), .B(n12512), .Z(n12403) );
  XNOR U12686 ( .A(n12409), .B(n12407), .Z(n12512) );
  AND U12687 ( .A(n12513), .B(n12514), .Z(n12407) );
  NANDN U12688 ( .A(n12515), .B(n12516), .Z(n12514) );
  NANDN U12689 ( .A(n12517), .B(n12518), .Z(n12516) );
  NANDN U12690 ( .A(n12518), .B(n12517), .Z(n12513) );
  ANDN U12691 ( .B(B[209]), .A(n35), .Z(n12409) );
  XNOR U12692 ( .A(n12417), .B(n12519), .Z(n12410) );
  XNOR U12693 ( .A(n12416), .B(n12414), .Z(n12519) );
  AND U12694 ( .A(n12520), .B(n12521), .Z(n12414) );
  NANDN U12695 ( .A(n12522), .B(n12523), .Z(n12521) );
  OR U12696 ( .A(n12524), .B(n12525), .Z(n12523) );
  NAND U12697 ( .A(n12525), .B(n12524), .Z(n12520) );
  ANDN U12698 ( .B(B[210]), .A(n36), .Z(n12416) );
  XNOR U12699 ( .A(n12424), .B(n12526), .Z(n12417) );
  XNOR U12700 ( .A(n12423), .B(n12421), .Z(n12526) );
  AND U12701 ( .A(n12527), .B(n12528), .Z(n12421) );
  NANDN U12702 ( .A(n12529), .B(n12530), .Z(n12528) );
  NANDN U12703 ( .A(n12531), .B(n12532), .Z(n12530) );
  NANDN U12704 ( .A(n12532), .B(n12531), .Z(n12527) );
  ANDN U12705 ( .B(B[211]), .A(n37), .Z(n12423) );
  XNOR U12706 ( .A(n12431), .B(n12533), .Z(n12424) );
  XNOR U12707 ( .A(n12430), .B(n12428), .Z(n12533) );
  AND U12708 ( .A(n12534), .B(n12535), .Z(n12428) );
  NANDN U12709 ( .A(n12536), .B(n12537), .Z(n12535) );
  OR U12710 ( .A(n12538), .B(n12539), .Z(n12537) );
  NAND U12711 ( .A(n12539), .B(n12538), .Z(n12534) );
  ANDN U12712 ( .B(B[212]), .A(n38), .Z(n12430) );
  XNOR U12713 ( .A(n12438), .B(n12540), .Z(n12431) );
  XNOR U12714 ( .A(n12437), .B(n12435), .Z(n12540) );
  AND U12715 ( .A(n12541), .B(n12542), .Z(n12435) );
  NANDN U12716 ( .A(n12543), .B(n12544), .Z(n12542) );
  NANDN U12717 ( .A(n12545), .B(n12546), .Z(n12544) );
  NANDN U12718 ( .A(n12546), .B(n12545), .Z(n12541) );
  ANDN U12719 ( .B(B[213]), .A(n39), .Z(n12437) );
  XNOR U12720 ( .A(n12445), .B(n12547), .Z(n12438) );
  XNOR U12721 ( .A(n12444), .B(n12442), .Z(n12547) );
  AND U12722 ( .A(n12548), .B(n12549), .Z(n12442) );
  NANDN U12723 ( .A(n12550), .B(n12551), .Z(n12549) );
  OR U12724 ( .A(n12552), .B(n12553), .Z(n12551) );
  NAND U12725 ( .A(n12553), .B(n12552), .Z(n12548) );
  ANDN U12726 ( .B(B[214]), .A(n40), .Z(n12444) );
  XNOR U12727 ( .A(n12452), .B(n12554), .Z(n12445) );
  XNOR U12728 ( .A(n12451), .B(n12449), .Z(n12554) );
  AND U12729 ( .A(n12555), .B(n12556), .Z(n12449) );
  NANDN U12730 ( .A(n12557), .B(n12558), .Z(n12556) );
  NAND U12731 ( .A(n12559), .B(n12560), .Z(n12558) );
  ANDN U12732 ( .B(B[215]), .A(n41), .Z(n12451) );
  XOR U12733 ( .A(n12458), .B(n12561), .Z(n12452) );
  XNOR U12734 ( .A(n12456), .B(n12459), .Z(n12561) );
  NAND U12735 ( .A(A[2]), .B(B[216]), .Z(n12459) );
  NANDN U12736 ( .A(n12562), .B(n12563), .Z(n12456) );
  AND U12737 ( .A(A[0]), .B(B[217]), .Z(n12563) );
  XNOR U12738 ( .A(n12461), .B(n12564), .Z(n12458) );
  NAND U12739 ( .A(A[0]), .B(B[218]), .Z(n12564) );
  NAND U12740 ( .A(B[217]), .B(A[1]), .Z(n12461) );
  NAND U12741 ( .A(n12565), .B(n12566), .Z(n307) );
  NANDN U12742 ( .A(n12567), .B(n12568), .Z(n12566) );
  OR U12743 ( .A(n12569), .B(n12570), .Z(n12568) );
  NAND U12744 ( .A(n12570), .B(n12569), .Z(n12565) );
  XOR U12745 ( .A(n309), .B(n308), .Z(\A1[215] ) );
  XOR U12746 ( .A(n12570), .B(n12571), .Z(n308) );
  XNOR U12747 ( .A(n12569), .B(n12567), .Z(n12571) );
  AND U12748 ( .A(n12572), .B(n12573), .Z(n12567) );
  NANDN U12749 ( .A(n12574), .B(n12575), .Z(n12573) );
  NANDN U12750 ( .A(n12576), .B(n12577), .Z(n12575) );
  NANDN U12751 ( .A(n12577), .B(n12576), .Z(n12572) );
  ANDN U12752 ( .B(B[202]), .A(n29), .Z(n12569) );
  XNOR U12753 ( .A(n12476), .B(n12578), .Z(n12570) );
  XNOR U12754 ( .A(n12475), .B(n12473), .Z(n12578) );
  AND U12755 ( .A(n12579), .B(n12580), .Z(n12473) );
  NANDN U12756 ( .A(n12581), .B(n12582), .Z(n12580) );
  OR U12757 ( .A(n12583), .B(n12584), .Z(n12582) );
  NAND U12758 ( .A(n12584), .B(n12583), .Z(n12579) );
  ANDN U12759 ( .B(B[203]), .A(n30), .Z(n12475) );
  XNOR U12760 ( .A(n12483), .B(n12585), .Z(n12476) );
  XNOR U12761 ( .A(n12482), .B(n12480), .Z(n12585) );
  AND U12762 ( .A(n12586), .B(n12587), .Z(n12480) );
  NANDN U12763 ( .A(n12588), .B(n12589), .Z(n12587) );
  NANDN U12764 ( .A(n12590), .B(n12591), .Z(n12589) );
  NANDN U12765 ( .A(n12591), .B(n12590), .Z(n12586) );
  ANDN U12766 ( .B(B[204]), .A(n31), .Z(n12482) );
  XNOR U12767 ( .A(n12490), .B(n12592), .Z(n12483) );
  XNOR U12768 ( .A(n12489), .B(n12487), .Z(n12592) );
  AND U12769 ( .A(n12593), .B(n12594), .Z(n12487) );
  NANDN U12770 ( .A(n12595), .B(n12596), .Z(n12594) );
  OR U12771 ( .A(n12597), .B(n12598), .Z(n12596) );
  NAND U12772 ( .A(n12598), .B(n12597), .Z(n12593) );
  ANDN U12773 ( .B(B[205]), .A(n32), .Z(n12489) );
  XNOR U12774 ( .A(n12497), .B(n12599), .Z(n12490) );
  XNOR U12775 ( .A(n12496), .B(n12494), .Z(n12599) );
  AND U12776 ( .A(n12600), .B(n12601), .Z(n12494) );
  NANDN U12777 ( .A(n12602), .B(n12603), .Z(n12601) );
  NANDN U12778 ( .A(n12604), .B(n12605), .Z(n12603) );
  NANDN U12779 ( .A(n12605), .B(n12604), .Z(n12600) );
  ANDN U12780 ( .B(B[206]), .A(n33), .Z(n12496) );
  XNOR U12781 ( .A(n12504), .B(n12606), .Z(n12497) );
  XNOR U12782 ( .A(n12503), .B(n12501), .Z(n12606) );
  AND U12783 ( .A(n12607), .B(n12608), .Z(n12501) );
  NANDN U12784 ( .A(n12609), .B(n12610), .Z(n12608) );
  OR U12785 ( .A(n12611), .B(n12612), .Z(n12610) );
  NAND U12786 ( .A(n12612), .B(n12611), .Z(n12607) );
  ANDN U12787 ( .B(B[207]), .A(n34), .Z(n12503) );
  XNOR U12788 ( .A(n12511), .B(n12613), .Z(n12504) );
  XNOR U12789 ( .A(n12510), .B(n12508), .Z(n12613) );
  AND U12790 ( .A(n12614), .B(n12615), .Z(n12508) );
  NANDN U12791 ( .A(n12616), .B(n12617), .Z(n12615) );
  NANDN U12792 ( .A(n12618), .B(n12619), .Z(n12617) );
  NANDN U12793 ( .A(n12619), .B(n12618), .Z(n12614) );
  ANDN U12794 ( .B(B[208]), .A(n35), .Z(n12510) );
  XNOR U12795 ( .A(n12518), .B(n12620), .Z(n12511) );
  XNOR U12796 ( .A(n12517), .B(n12515), .Z(n12620) );
  AND U12797 ( .A(n12621), .B(n12622), .Z(n12515) );
  NANDN U12798 ( .A(n12623), .B(n12624), .Z(n12622) );
  OR U12799 ( .A(n12625), .B(n12626), .Z(n12624) );
  NAND U12800 ( .A(n12626), .B(n12625), .Z(n12621) );
  ANDN U12801 ( .B(B[209]), .A(n36), .Z(n12517) );
  XNOR U12802 ( .A(n12525), .B(n12627), .Z(n12518) );
  XNOR U12803 ( .A(n12524), .B(n12522), .Z(n12627) );
  AND U12804 ( .A(n12628), .B(n12629), .Z(n12522) );
  NANDN U12805 ( .A(n12630), .B(n12631), .Z(n12629) );
  NANDN U12806 ( .A(n12632), .B(n12633), .Z(n12631) );
  NANDN U12807 ( .A(n12633), .B(n12632), .Z(n12628) );
  ANDN U12808 ( .B(B[210]), .A(n37), .Z(n12524) );
  XNOR U12809 ( .A(n12532), .B(n12634), .Z(n12525) );
  XNOR U12810 ( .A(n12531), .B(n12529), .Z(n12634) );
  AND U12811 ( .A(n12635), .B(n12636), .Z(n12529) );
  NANDN U12812 ( .A(n12637), .B(n12638), .Z(n12636) );
  OR U12813 ( .A(n12639), .B(n12640), .Z(n12638) );
  NAND U12814 ( .A(n12640), .B(n12639), .Z(n12635) );
  ANDN U12815 ( .B(B[211]), .A(n38), .Z(n12531) );
  XNOR U12816 ( .A(n12539), .B(n12641), .Z(n12532) );
  XNOR U12817 ( .A(n12538), .B(n12536), .Z(n12641) );
  AND U12818 ( .A(n12642), .B(n12643), .Z(n12536) );
  NANDN U12819 ( .A(n12644), .B(n12645), .Z(n12643) );
  NANDN U12820 ( .A(n12646), .B(n12647), .Z(n12645) );
  NANDN U12821 ( .A(n12647), .B(n12646), .Z(n12642) );
  ANDN U12822 ( .B(B[212]), .A(n39), .Z(n12538) );
  XNOR U12823 ( .A(n12546), .B(n12648), .Z(n12539) );
  XNOR U12824 ( .A(n12545), .B(n12543), .Z(n12648) );
  AND U12825 ( .A(n12649), .B(n12650), .Z(n12543) );
  NANDN U12826 ( .A(n12651), .B(n12652), .Z(n12650) );
  OR U12827 ( .A(n12653), .B(n12654), .Z(n12652) );
  NAND U12828 ( .A(n12654), .B(n12653), .Z(n12649) );
  ANDN U12829 ( .B(B[213]), .A(n40), .Z(n12545) );
  XNOR U12830 ( .A(n12553), .B(n12655), .Z(n12546) );
  XNOR U12831 ( .A(n12552), .B(n12550), .Z(n12655) );
  AND U12832 ( .A(n12656), .B(n12657), .Z(n12550) );
  NANDN U12833 ( .A(n12658), .B(n12659), .Z(n12657) );
  NAND U12834 ( .A(n12660), .B(n12661), .Z(n12659) );
  ANDN U12835 ( .B(B[214]), .A(n41), .Z(n12552) );
  XOR U12836 ( .A(n12559), .B(n12662), .Z(n12553) );
  XNOR U12837 ( .A(n12557), .B(n12560), .Z(n12662) );
  NAND U12838 ( .A(A[2]), .B(B[215]), .Z(n12560) );
  NANDN U12839 ( .A(n12663), .B(n12664), .Z(n12557) );
  AND U12840 ( .A(A[0]), .B(B[216]), .Z(n12664) );
  XNOR U12841 ( .A(n12562), .B(n12665), .Z(n12559) );
  NAND U12842 ( .A(A[0]), .B(B[217]), .Z(n12665) );
  NAND U12843 ( .A(B[216]), .B(A[1]), .Z(n12562) );
  NAND U12844 ( .A(n12666), .B(n12667), .Z(n309) );
  NANDN U12845 ( .A(n12668), .B(n12669), .Z(n12667) );
  OR U12846 ( .A(n12670), .B(n12671), .Z(n12669) );
  NAND U12847 ( .A(n12671), .B(n12670), .Z(n12666) );
  XOR U12848 ( .A(n311), .B(n310), .Z(\A1[214] ) );
  XOR U12849 ( .A(n12671), .B(n12672), .Z(n310) );
  XNOR U12850 ( .A(n12670), .B(n12668), .Z(n12672) );
  AND U12851 ( .A(n12673), .B(n12674), .Z(n12668) );
  NANDN U12852 ( .A(n12675), .B(n12676), .Z(n12674) );
  NANDN U12853 ( .A(n12677), .B(n12678), .Z(n12676) );
  NANDN U12854 ( .A(n12678), .B(n12677), .Z(n12673) );
  ANDN U12855 ( .B(B[201]), .A(n29), .Z(n12670) );
  XNOR U12856 ( .A(n12577), .B(n12679), .Z(n12671) );
  XNOR U12857 ( .A(n12576), .B(n12574), .Z(n12679) );
  AND U12858 ( .A(n12680), .B(n12681), .Z(n12574) );
  NANDN U12859 ( .A(n12682), .B(n12683), .Z(n12681) );
  OR U12860 ( .A(n12684), .B(n12685), .Z(n12683) );
  NAND U12861 ( .A(n12685), .B(n12684), .Z(n12680) );
  ANDN U12862 ( .B(B[202]), .A(n30), .Z(n12576) );
  XNOR U12863 ( .A(n12584), .B(n12686), .Z(n12577) );
  XNOR U12864 ( .A(n12583), .B(n12581), .Z(n12686) );
  AND U12865 ( .A(n12687), .B(n12688), .Z(n12581) );
  NANDN U12866 ( .A(n12689), .B(n12690), .Z(n12688) );
  NANDN U12867 ( .A(n12691), .B(n12692), .Z(n12690) );
  NANDN U12868 ( .A(n12692), .B(n12691), .Z(n12687) );
  ANDN U12869 ( .B(B[203]), .A(n31), .Z(n12583) );
  XNOR U12870 ( .A(n12591), .B(n12693), .Z(n12584) );
  XNOR U12871 ( .A(n12590), .B(n12588), .Z(n12693) );
  AND U12872 ( .A(n12694), .B(n12695), .Z(n12588) );
  NANDN U12873 ( .A(n12696), .B(n12697), .Z(n12695) );
  OR U12874 ( .A(n12698), .B(n12699), .Z(n12697) );
  NAND U12875 ( .A(n12699), .B(n12698), .Z(n12694) );
  ANDN U12876 ( .B(B[204]), .A(n32), .Z(n12590) );
  XNOR U12877 ( .A(n12598), .B(n12700), .Z(n12591) );
  XNOR U12878 ( .A(n12597), .B(n12595), .Z(n12700) );
  AND U12879 ( .A(n12701), .B(n12702), .Z(n12595) );
  NANDN U12880 ( .A(n12703), .B(n12704), .Z(n12702) );
  NANDN U12881 ( .A(n12705), .B(n12706), .Z(n12704) );
  NANDN U12882 ( .A(n12706), .B(n12705), .Z(n12701) );
  ANDN U12883 ( .B(B[205]), .A(n33), .Z(n12597) );
  XNOR U12884 ( .A(n12605), .B(n12707), .Z(n12598) );
  XNOR U12885 ( .A(n12604), .B(n12602), .Z(n12707) );
  AND U12886 ( .A(n12708), .B(n12709), .Z(n12602) );
  NANDN U12887 ( .A(n12710), .B(n12711), .Z(n12709) );
  OR U12888 ( .A(n12712), .B(n12713), .Z(n12711) );
  NAND U12889 ( .A(n12713), .B(n12712), .Z(n12708) );
  ANDN U12890 ( .B(B[206]), .A(n34), .Z(n12604) );
  XNOR U12891 ( .A(n12612), .B(n12714), .Z(n12605) );
  XNOR U12892 ( .A(n12611), .B(n12609), .Z(n12714) );
  AND U12893 ( .A(n12715), .B(n12716), .Z(n12609) );
  NANDN U12894 ( .A(n12717), .B(n12718), .Z(n12716) );
  NANDN U12895 ( .A(n12719), .B(n12720), .Z(n12718) );
  NANDN U12896 ( .A(n12720), .B(n12719), .Z(n12715) );
  ANDN U12897 ( .B(B[207]), .A(n35), .Z(n12611) );
  XNOR U12898 ( .A(n12619), .B(n12721), .Z(n12612) );
  XNOR U12899 ( .A(n12618), .B(n12616), .Z(n12721) );
  AND U12900 ( .A(n12722), .B(n12723), .Z(n12616) );
  NANDN U12901 ( .A(n12724), .B(n12725), .Z(n12723) );
  OR U12902 ( .A(n12726), .B(n12727), .Z(n12725) );
  NAND U12903 ( .A(n12727), .B(n12726), .Z(n12722) );
  ANDN U12904 ( .B(B[208]), .A(n36), .Z(n12618) );
  XNOR U12905 ( .A(n12626), .B(n12728), .Z(n12619) );
  XNOR U12906 ( .A(n12625), .B(n12623), .Z(n12728) );
  AND U12907 ( .A(n12729), .B(n12730), .Z(n12623) );
  NANDN U12908 ( .A(n12731), .B(n12732), .Z(n12730) );
  NANDN U12909 ( .A(n12733), .B(n12734), .Z(n12732) );
  NANDN U12910 ( .A(n12734), .B(n12733), .Z(n12729) );
  ANDN U12911 ( .B(B[209]), .A(n37), .Z(n12625) );
  XNOR U12912 ( .A(n12633), .B(n12735), .Z(n12626) );
  XNOR U12913 ( .A(n12632), .B(n12630), .Z(n12735) );
  AND U12914 ( .A(n12736), .B(n12737), .Z(n12630) );
  NANDN U12915 ( .A(n12738), .B(n12739), .Z(n12737) );
  OR U12916 ( .A(n12740), .B(n12741), .Z(n12739) );
  NAND U12917 ( .A(n12741), .B(n12740), .Z(n12736) );
  ANDN U12918 ( .B(B[210]), .A(n38), .Z(n12632) );
  XNOR U12919 ( .A(n12640), .B(n12742), .Z(n12633) );
  XNOR U12920 ( .A(n12639), .B(n12637), .Z(n12742) );
  AND U12921 ( .A(n12743), .B(n12744), .Z(n12637) );
  NANDN U12922 ( .A(n12745), .B(n12746), .Z(n12744) );
  NANDN U12923 ( .A(n12747), .B(n12748), .Z(n12746) );
  NANDN U12924 ( .A(n12748), .B(n12747), .Z(n12743) );
  ANDN U12925 ( .B(B[211]), .A(n39), .Z(n12639) );
  XNOR U12926 ( .A(n12647), .B(n12749), .Z(n12640) );
  XNOR U12927 ( .A(n12646), .B(n12644), .Z(n12749) );
  AND U12928 ( .A(n12750), .B(n12751), .Z(n12644) );
  NANDN U12929 ( .A(n12752), .B(n12753), .Z(n12751) );
  OR U12930 ( .A(n12754), .B(n12755), .Z(n12753) );
  NAND U12931 ( .A(n12755), .B(n12754), .Z(n12750) );
  ANDN U12932 ( .B(B[212]), .A(n40), .Z(n12646) );
  XNOR U12933 ( .A(n12654), .B(n12756), .Z(n12647) );
  XNOR U12934 ( .A(n12653), .B(n12651), .Z(n12756) );
  AND U12935 ( .A(n12757), .B(n12758), .Z(n12651) );
  NANDN U12936 ( .A(n12759), .B(n12760), .Z(n12758) );
  NAND U12937 ( .A(n12761), .B(n12762), .Z(n12760) );
  ANDN U12938 ( .B(B[213]), .A(n41), .Z(n12653) );
  XOR U12939 ( .A(n12660), .B(n12763), .Z(n12654) );
  XNOR U12940 ( .A(n12658), .B(n12661), .Z(n12763) );
  NAND U12941 ( .A(A[2]), .B(B[214]), .Z(n12661) );
  NANDN U12942 ( .A(n12764), .B(n12765), .Z(n12658) );
  AND U12943 ( .A(A[0]), .B(B[215]), .Z(n12765) );
  XNOR U12944 ( .A(n12663), .B(n12766), .Z(n12660) );
  NAND U12945 ( .A(A[0]), .B(B[216]), .Z(n12766) );
  NAND U12946 ( .A(B[215]), .B(A[1]), .Z(n12663) );
  NAND U12947 ( .A(n12767), .B(n12768), .Z(n311) );
  NANDN U12948 ( .A(n12769), .B(n12770), .Z(n12768) );
  OR U12949 ( .A(n12771), .B(n12772), .Z(n12770) );
  NAND U12950 ( .A(n12772), .B(n12771), .Z(n12767) );
  XOR U12951 ( .A(n313), .B(n312), .Z(\A1[213] ) );
  XOR U12952 ( .A(n12772), .B(n12773), .Z(n312) );
  XNOR U12953 ( .A(n12771), .B(n12769), .Z(n12773) );
  AND U12954 ( .A(n12774), .B(n12775), .Z(n12769) );
  NANDN U12955 ( .A(n12776), .B(n12777), .Z(n12775) );
  NANDN U12956 ( .A(n12778), .B(n12779), .Z(n12777) );
  NANDN U12957 ( .A(n12779), .B(n12778), .Z(n12774) );
  ANDN U12958 ( .B(B[200]), .A(n29), .Z(n12771) );
  XNOR U12959 ( .A(n12678), .B(n12780), .Z(n12772) );
  XNOR U12960 ( .A(n12677), .B(n12675), .Z(n12780) );
  AND U12961 ( .A(n12781), .B(n12782), .Z(n12675) );
  NANDN U12962 ( .A(n12783), .B(n12784), .Z(n12782) );
  OR U12963 ( .A(n12785), .B(n12786), .Z(n12784) );
  NAND U12964 ( .A(n12786), .B(n12785), .Z(n12781) );
  ANDN U12965 ( .B(B[201]), .A(n30), .Z(n12677) );
  XNOR U12966 ( .A(n12685), .B(n12787), .Z(n12678) );
  XNOR U12967 ( .A(n12684), .B(n12682), .Z(n12787) );
  AND U12968 ( .A(n12788), .B(n12789), .Z(n12682) );
  NANDN U12969 ( .A(n12790), .B(n12791), .Z(n12789) );
  NANDN U12970 ( .A(n12792), .B(n12793), .Z(n12791) );
  NANDN U12971 ( .A(n12793), .B(n12792), .Z(n12788) );
  ANDN U12972 ( .B(B[202]), .A(n31), .Z(n12684) );
  XNOR U12973 ( .A(n12692), .B(n12794), .Z(n12685) );
  XNOR U12974 ( .A(n12691), .B(n12689), .Z(n12794) );
  AND U12975 ( .A(n12795), .B(n12796), .Z(n12689) );
  NANDN U12976 ( .A(n12797), .B(n12798), .Z(n12796) );
  OR U12977 ( .A(n12799), .B(n12800), .Z(n12798) );
  NAND U12978 ( .A(n12800), .B(n12799), .Z(n12795) );
  ANDN U12979 ( .B(B[203]), .A(n32), .Z(n12691) );
  XNOR U12980 ( .A(n12699), .B(n12801), .Z(n12692) );
  XNOR U12981 ( .A(n12698), .B(n12696), .Z(n12801) );
  AND U12982 ( .A(n12802), .B(n12803), .Z(n12696) );
  NANDN U12983 ( .A(n12804), .B(n12805), .Z(n12803) );
  NANDN U12984 ( .A(n12806), .B(n12807), .Z(n12805) );
  NANDN U12985 ( .A(n12807), .B(n12806), .Z(n12802) );
  ANDN U12986 ( .B(B[204]), .A(n33), .Z(n12698) );
  XNOR U12987 ( .A(n12706), .B(n12808), .Z(n12699) );
  XNOR U12988 ( .A(n12705), .B(n12703), .Z(n12808) );
  AND U12989 ( .A(n12809), .B(n12810), .Z(n12703) );
  NANDN U12990 ( .A(n12811), .B(n12812), .Z(n12810) );
  OR U12991 ( .A(n12813), .B(n12814), .Z(n12812) );
  NAND U12992 ( .A(n12814), .B(n12813), .Z(n12809) );
  ANDN U12993 ( .B(B[205]), .A(n34), .Z(n12705) );
  XNOR U12994 ( .A(n12713), .B(n12815), .Z(n12706) );
  XNOR U12995 ( .A(n12712), .B(n12710), .Z(n12815) );
  AND U12996 ( .A(n12816), .B(n12817), .Z(n12710) );
  NANDN U12997 ( .A(n12818), .B(n12819), .Z(n12817) );
  NANDN U12998 ( .A(n12820), .B(n12821), .Z(n12819) );
  NANDN U12999 ( .A(n12821), .B(n12820), .Z(n12816) );
  ANDN U13000 ( .B(B[206]), .A(n35), .Z(n12712) );
  XNOR U13001 ( .A(n12720), .B(n12822), .Z(n12713) );
  XNOR U13002 ( .A(n12719), .B(n12717), .Z(n12822) );
  AND U13003 ( .A(n12823), .B(n12824), .Z(n12717) );
  NANDN U13004 ( .A(n12825), .B(n12826), .Z(n12824) );
  OR U13005 ( .A(n12827), .B(n12828), .Z(n12826) );
  NAND U13006 ( .A(n12828), .B(n12827), .Z(n12823) );
  ANDN U13007 ( .B(B[207]), .A(n36), .Z(n12719) );
  XNOR U13008 ( .A(n12727), .B(n12829), .Z(n12720) );
  XNOR U13009 ( .A(n12726), .B(n12724), .Z(n12829) );
  AND U13010 ( .A(n12830), .B(n12831), .Z(n12724) );
  NANDN U13011 ( .A(n12832), .B(n12833), .Z(n12831) );
  NANDN U13012 ( .A(n12834), .B(n12835), .Z(n12833) );
  NANDN U13013 ( .A(n12835), .B(n12834), .Z(n12830) );
  ANDN U13014 ( .B(B[208]), .A(n37), .Z(n12726) );
  XNOR U13015 ( .A(n12734), .B(n12836), .Z(n12727) );
  XNOR U13016 ( .A(n12733), .B(n12731), .Z(n12836) );
  AND U13017 ( .A(n12837), .B(n12838), .Z(n12731) );
  NANDN U13018 ( .A(n12839), .B(n12840), .Z(n12838) );
  OR U13019 ( .A(n12841), .B(n12842), .Z(n12840) );
  NAND U13020 ( .A(n12842), .B(n12841), .Z(n12837) );
  ANDN U13021 ( .B(B[209]), .A(n38), .Z(n12733) );
  XNOR U13022 ( .A(n12741), .B(n12843), .Z(n12734) );
  XNOR U13023 ( .A(n12740), .B(n12738), .Z(n12843) );
  AND U13024 ( .A(n12844), .B(n12845), .Z(n12738) );
  NANDN U13025 ( .A(n12846), .B(n12847), .Z(n12845) );
  NANDN U13026 ( .A(n12848), .B(n12849), .Z(n12847) );
  NANDN U13027 ( .A(n12849), .B(n12848), .Z(n12844) );
  ANDN U13028 ( .B(B[210]), .A(n39), .Z(n12740) );
  XNOR U13029 ( .A(n12748), .B(n12850), .Z(n12741) );
  XNOR U13030 ( .A(n12747), .B(n12745), .Z(n12850) );
  AND U13031 ( .A(n12851), .B(n12852), .Z(n12745) );
  NANDN U13032 ( .A(n12853), .B(n12854), .Z(n12852) );
  OR U13033 ( .A(n12855), .B(n12856), .Z(n12854) );
  NAND U13034 ( .A(n12856), .B(n12855), .Z(n12851) );
  ANDN U13035 ( .B(B[211]), .A(n40), .Z(n12747) );
  XNOR U13036 ( .A(n12755), .B(n12857), .Z(n12748) );
  XNOR U13037 ( .A(n12754), .B(n12752), .Z(n12857) );
  AND U13038 ( .A(n12858), .B(n12859), .Z(n12752) );
  NANDN U13039 ( .A(n12860), .B(n12861), .Z(n12859) );
  NAND U13040 ( .A(n12862), .B(n12863), .Z(n12861) );
  ANDN U13041 ( .B(B[212]), .A(n41), .Z(n12754) );
  XOR U13042 ( .A(n12761), .B(n12864), .Z(n12755) );
  XNOR U13043 ( .A(n12759), .B(n12762), .Z(n12864) );
  NAND U13044 ( .A(A[2]), .B(B[213]), .Z(n12762) );
  NANDN U13045 ( .A(n12865), .B(n12866), .Z(n12759) );
  AND U13046 ( .A(A[0]), .B(B[214]), .Z(n12866) );
  XNOR U13047 ( .A(n12764), .B(n12867), .Z(n12761) );
  NAND U13048 ( .A(A[0]), .B(B[215]), .Z(n12867) );
  NAND U13049 ( .A(B[214]), .B(A[1]), .Z(n12764) );
  NAND U13050 ( .A(n12868), .B(n12869), .Z(n313) );
  NANDN U13051 ( .A(n12870), .B(n12871), .Z(n12869) );
  OR U13052 ( .A(n12872), .B(n12873), .Z(n12871) );
  NAND U13053 ( .A(n12873), .B(n12872), .Z(n12868) );
  XOR U13054 ( .A(n315), .B(n314), .Z(\A1[212] ) );
  XOR U13055 ( .A(n12873), .B(n12874), .Z(n314) );
  XNOR U13056 ( .A(n12872), .B(n12870), .Z(n12874) );
  AND U13057 ( .A(n12875), .B(n12876), .Z(n12870) );
  NANDN U13058 ( .A(n12877), .B(n12878), .Z(n12876) );
  NANDN U13059 ( .A(n12879), .B(n12880), .Z(n12878) );
  NANDN U13060 ( .A(n12880), .B(n12879), .Z(n12875) );
  ANDN U13061 ( .B(B[199]), .A(n29), .Z(n12872) );
  XNOR U13062 ( .A(n12779), .B(n12881), .Z(n12873) );
  XNOR U13063 ( .A(n12778), .B(n12776), .Z(n12881) );
  AND U13064 ( .A(n12882), .B(n12883), .Z(n12776) );
  NANDN U13065 ( .A(n12884), .B(n12885), .Z(n12883) );
  OR U13066 ( .A(n12886), .B(n12887), .Z(n12885) );
  NAND U13067 ( .A(n12887), .B(n12886), .Z(n12882) );
  ANDN U13068 ( .B(B[200]), .A(n30), .Z(n12778) );
  XNOR U13069 ( .A(n12786), .B(n12888), .Z(n12779) );
  XNOR U13070 ( .A(n12785), .B(n12783), .Z(n12888) );
  AND U13071 ( .A(n12889), .B(n12890), .Z(n12783) );
  NANDN U13072 ( .A(n12891), .B(n12892), .Z(n12890) );
  NANDN U13073 ( .A(n12893), .B(n12894), .Z(n12892) );
  NANDN U13074 ( .A(n12894), .B(n12893), .Z(n12889) );
  ANDN U13075 ( .B(B[201]), .A(n31), .Z(n12785) );
  XNOR U13076 ( .A(n12793), .B(n12895), .Z(n12786) );
  XNOR U13077 ( .A(n12792), .B(n12790), .Z(n12895) );
  AND U13078 ( .A(n12896), .B(n12897), .Z(n12790) );
  NANDN U13079 ( .A(n12898), .B(n12899), .Z(n12897) );
  OR U13080 ( .A(n12900), .B(n12901), .Z(n12899) );
  NAND U13081 ( .A(n12901), .B(n12900), .Z(n12896) );
  ANDN U13082 ( .B(B[202]), .A(n32), .Z(n12792) );
  XNOR U13083 ( .A(n12800), .B(n12902), .Z(n12793) );
  XNOR U13084 ( .A(n12799), .B(n12797), .Z(n12902) );
  AND U13085 ( .A(n12903), .B(n12904), .Z(n12797) );
  NANDN U13086 ( .A(n12905), .B(n12906), .Z(n12904) );
  NANDN U13087 ( .A(n12907), .B(n12908), .Z(n12906) );
  NANDN U13088 ( .A(n12908), .B(n12907), .Z(n12903) );
  ANDN U13089 ( .B(B[203]), .A(n33), .Z(n12799) );
  XNOR U13090 ( .A(n12807), .B(n12909), .Z(n12800) );
  XNOR U13091 ( .A(n12806), .B(n12804), .Z(n12909) );
  AND U13092 ( .A(n12910), .B(n12911), .Z(n12804) );
  NANDN U13093 ( .A(n12912), .B(n12913), .Z(n12911) );
  OR U13094 ( .A(n12914), .B(n12915), .Z(n12913) );
  NAND U13095 ( .A(n12915), .B(n12914), .Z(n12910) );
  ANDN U13096 ( .B(B[204]), .A(n34), .Z(n12806) );
  XNOR U13097 ( .A(n12814), .B(n12916), .Z(n12807) );
  XNOR U13098 ( .A(n12813), .B(n12811), .Z(n12916) );
  AND U13099 ( .A(n12917), .B(n12918), .Z(n12811) );
  NANDN U13100 ( .A(n12919), .B(n12920), .Z(n12918) );
  NANDN U13101 ( .A(n12921), .B(n12922), .Z(n12920) );
  NANDN U13102 ( .A(n12922), .B(n12921), .Z(n12917) );
  ANDN U13103 ( .B(B[205]), .A(n35), .Z(n12813) );
  XNOR U13104 ( .A(n12821), .B(n12923), .Z(n12814) );
  XNOR U13105 ( .A(n12820), .B(n12818), .Z(n12923) );
  AND U13106 ( .A(n12924), .B(n12925), .Z(n12818) );
  NANDN U13107 ( .A(n12926), .B(n12927), .Z(n12925) );
  OR U13108 ( .A(n12928), .B(n12929), .Z(n12927) );
  NAND U13109 ( .A(n12929), .B(n12928), .Z(n12924) );
  ANDN U13110 ( .B(B[206]), .A(n36), .Z(n12820) );
  XNOR U13111 ( .A(n12828), .B(n12930), .Z(n12821) );
  XNOR U13112 ( .A(n12827), .B(n12825), .Z(n12930) );
  AND U13113 ( .A(n12931), .B(n12932), .Z(n12825) );
  NANDN U13114 ( .A(n12933), .B(n12934), .Z(n12932) );
  NANDN U13115 ( .A(n12935), .B(n12936), .Z(n12934) );
  NANDN U13116 ( .A(n12936), .B(n12935), .Z(n12931) );
  ANDN U13117 ( .B(B[207]), .A(n37), .Z(n12827) );
  XNOR U13118 ( .A(n12835), .B(n12937), .Z(n12828) );
  XNOR U13119 ( .A(n12834), .B(n12832), .Z(n12937) );
  AND U13120 ( .A(n12938), .B(n12939), .Z(n12832) );
  NANDN U13121 ( .A(n12940), .B(n12941), .Z(n12939) );
  OR U13122 ( .A(n12942), .B(n12943), .Z(n12941) );
  NAND U13123 ( .A(n12943), .B(n12942), .Z(n12938) );
  ANDN U13124 ( .B(B[208]), .A(n38), .Z(n12834) );
  XNOR U13125 ( .A(n12842), .B(n12944), .Z(n12835) );
  XNOR U13126 ( .A(n12841), .B(n12839), .Z(n12944) );
  AND U13127 ( .A(n12945), .B(n12946), .Z(n12839) );
  NANDN U13128 ( .A(n12947), .B(n12948), .Z(n12946) );
  NANDN U13129 ( .A(n12949), .B(n12950), .Z(n12948) );
  NANDN U13130 ( .A(n12950), .B(n12949), .Z(n12945) );
  ANDN U13131 ( .B(B[209]), .A(n39), .Z(n12841) );
  XNOR U13132 ( .A(n12849), .B(n12951), .Z(n12842) );
  XNOR U13133 ( .A(n12848), .B(n12846), .Z(n12951) );
  AND U13134 ( .A(n12952), .B(n12953), .Z(n12846) );
  NANDN U13135 ( .A(n12954), .B(n12955), .Z(n12953) );
  OR U13136 ( .A(n12956), .B(n12957), .Z(n12955) );
  NAND U13137 ( .A(n12957), .B(n12956), .Z(n12952) );
  ANDN U13138 ( .B(B[210]), .A(n40), .Z(n12848) );
  XNOR U13139 ( .A(n12856), .B(n12958), .Z(n12849) );
  XNOR U13140 ( .A(n12855), .B(n12853), .Z(n12958) );
  AND U13141 ( .A(n12959), .B(n12960), .Z(n12853) );
  NANDN U13142 ( .A(n12961), .B(n12962), .Z(n12960) );
  NAND U13143 ( .A(n12963), .B(n12964), .Z(n12962) );
  ANDN U13144 ( .B(B[211]), .A(n41), .Z(n12855) );
  XOR U13145 ( .A(n12862), .B(n12965), .Z(n12856) );
  XNOR U13146 ( .A(n12860), .B(n12863), .Z(n12965) );
  NAND U13147 ( .A(A[2]), .B(B[212]), .Z(n12863) );
  NANDN U13148 ( .A(n12966), .B(n12967), .Z(n12860) );
  AND U13149 ( .A(A[0]), .B(B[213]), .Z(n12967) );
  XNOR U13150 ( .A(n12865), .B(n12968), .Z(n12862) );
  NAND U13151 ( .A(A[0]), .B(B[214]), .Z(n12968) );
  NAND U13152 ( .A(B[213]), .B(A[1]), .Z(n12865) );
  NAND U13153 ( .A(n12969), .B(n12970), .Z(n315) );
  NANDN U13154 ( .A(n12971), .B(n12972), .Z(n12970) );
  OR U13155 ( .A(n12973), .B(n12974), .Z(n12972) );
  NAND U13156 ( .A(n12974), .B(n12973), .Z(n12969) );
  XOR U13157 ( .A(n317), .B(n316), .Z(\A1[211] ) );
  XOR U13158 ( .A(n12974), .B(n12975), .Z(n316) );
  XNOR U13159 ( .A(n12973), .B(n12971), .Z(n12975) );
  AND U13160 ( .A(n12976), .B(n12977), .Z(n12971) );
  NANDN U13161 ( .A(n12978), .B(n12979), .Z(n12977) );
  NANDN U13162 ( .A(n12980), .B(n12981), .Z(n12979) );
  NANDN U13163 ( .A(n12981), .B(n12980), .Z(n12976) );
  ANDN U13164 ( .B(B[198]), .A(n29), .Z(n12973) );
  XNOR U13165 ( .A(n12880), .B(n12982), .Z(n12974) );
  XNOR U13166 ( .A(n12879), .B(n12877), .Z(n12982) );
  AND U13167 ( .A(n12983), .B(n12984), .Z(n12877) );
  NANDN U13168 ( .A(n12985), .B(n12986), .Z(n12984) );
  OR U13169 ( .A(n12987), .B(n12988), .Z(n12986) );
  NAND U13170 ( .A(n12988), .B(n12987), .Z(n12983) );
  ANDN U13171 ( .B(B[199]), .A(n30), .Z(n12879) );
  XNOR U13172 ( .A(n12887), .B(n12989), .Z(n12880) );
  XNOR U13173 ( .A(n12886), .B(n12884), .Z(n12989) );
  AND U13174 ( .A(n12990), .B(n12991), .Z(n12884) );
  NANDN U13175 ( .A(n12992), .B(n12993), .Z(n12991) );
  NANDN U13176 ( .A(n12994), .B(n12995), .Z(n12993) );
  NANDN U13177 ( .A(n12995), .B(n12994), .Z(n12990) );
  ANDN U13178 ( .B(B[200]), .A(n31), .Z(n12886) );
  XNOR U13179 ( .A(n12894), .B(n12996), .Z(n12887) );
  XNOR U13180 ( .A(n12893), .B(n12891), .Z(n12996) );
  AND U13181 ( .A(n12997), .B(n12998), .Z(n12891) );
  NANDN U13182 ( .A(n12999), .B(n13000), .Z(n12998) );
  OR U13183 ( .A(n13001), .B(n13002), .Z(n13000) );
  NAND U13184 ( .A(n13002), .B(n13001), .Z(n12997) );
  ANDN U13185 ( .B(B[201]), .A(n32), .Z(n12893) );
  XNOR U13186 ( .A(n12901), .B(n13003), .Z(n12894) );
  XNOR U13187 ( .A(n12900), .B(n12898), .Z(n13003) );
  AND U13188 ( .A(n13004), .B(n13005), .Z(n12898) );
  NANDN U13189 ( .A(n13006), .B(n13007), .Z(n13005) );
  NANDN U13190 ( .A(n13008), .B(n13009), .Z(n13007) );
  NANDN U13191 ( .A(n13009), .B(n13008), .Z(n13004) );
  ANDN U13192 ( .B(B[202]), .A(n33), .Z(n12900) );
  XNOR U13193 ( .A(n12908), .B(n13010), .Z(n12901) );
  XNOR U13194 ( .A(n12907), .B(n12905), .Z(n13010) );
  AND U13195 ( .A(n13011), .B(n13012), .Z(n12905) );
  NANDN U13196 ( .A(n13013), .B(n13014), .Z(n13012) );
  OR U13197 ( .A(n13015), .B(n13016), .Z(n13014) );
  NAND U13198 ( .A(n13016), .B(n13015), .Z(n13011) );
  ANDN U13199 ( .B(B[203]), .A(n34), .Z(n12907) );
  XNOR U13200 ( .A(n12915), .B(n13017), .Z(n12908) );
  XNOR U13201 ( .A(n12914), .B(n12912), .Z(n13017) );
  AND U13202 ( .A(n13018), .B(n13019), .Z(n12912) );
  NANDN U13203 ( .A(n13020), .B(n13021), .Z(n13019) );
  NANDN U13204 ( .A(n13022), .B(n13023), .Z(n13021) );
  NANDN U13205 ( .A(n13023), .B(n13022), .Z(n13018) );
  ANDN U13206 ( .B(B[204]), .A(n35), .Z(n12914) );
  XNOR U13207 ( .A(n12922), .B(n13024), .Z(n12915) );
  XNOR U13208 ( .A(n12921), .B(n12919), .Z(n13024) );
  AND U13209 ( .A(n13025), .B(n13026), .Z(n12919) );
  NANDN U13210 ( .A(n13027), .B(n13028), .Z(n13026) );
  OR U13211 ( .A(n13029), .B(n13030), .Z(n13028) );
  NAND U13212 ( .A(n13030), .B(n13029), .Z(n13025) );
  ANDN U13213 ( .B(B[205]), .A(n36), .Z(n12921) );
  XNOR U13214 ( .A(n12929), .B(n13031), .Z(n12922) );
  XNOR U13215 ( .A(n12928), .B(n12926), .Z(n13031) );
  AND U13216 ( .A(n13032), .B(n13033), .Z(n12926) );
  NANDN U13217 ( .A(n13034), .B(n13035), .Z(n13033) );
  NANDN U13218 ( .A(n13036), .B(n13037), .Z(n13035) );
  NANDN U13219 ( .A(n13037), .B(n13036), .Z(n13032) );
  ANDN U13220 ( .B(B[206]), .A(n37), .Z(n12928) );
  XNOR U13221 ( .A(n12936), .B(n13038), .Z(n12929) );
  XNOR U13222 ( .A(n12935), .B(n12933), .Z(n13038) );
  AND U13223 ( .A(n13039), .B(n13040), .Z(n12933) );
  NANDN U13224 ( .A(n13041), .B(n13042), .Z(n13040) );
  OR U13225 ( .A(n13043), .B(n13044), .Z(n13042) );
  NAND U13226 ( .A(n13044), .B(n13043), .Z(n13039) );
  ANDN U13227 ( .B(B[207]), .A(n38), .Z(n12935) );
  XNOR U13228 ( .A(n12943), .B(n13045), .Z(n12936) );
  XNOR U13229 ( .A(n12942), .B(n12940), .Z(n13045) );
  AND U13230 ( .A(n13046), .B(n13047), .Z(n12940) );
  NANDN U13231 ( .A(n13048), .B(n13049), .Z(n13047) );
  NANDN U13232 ( .A(n13050), .B(n13051), .Z(n13049) );
  NANDN U13233 ( .A(n13051), .B(n13050), .Z(n13046) );
  ANDN U13234 ( .B(B[208]), .A(n39), .Z(n12942) );
  XNOR U13235 ( .A(n12950), .B(n13052), .Z(n12943) );
  XNOR U13236 ( .A(n12949), .B(n12947), .Z(n13052) );
  AND U13237 ( .A(n13053), .B(n13054), .Z(n12947) );
  NANDN U13238 ( .A(n13055), .B(n13056), .Z(n13054) );
  OR U13239 ( .A(n13057), .B(n13058), .Z(n13056) );
  NAND U13240 ( .A(n13058), .B(n13057), .Z(n13053) );
  ANDN U13241 ( .B(B[209]), .A(n40), .Z(n12949) );
  XNOR U13242 ( .A(n12957), .B(n13059), .Z(n12950) );
  XNOR U13243 ( .A(n12956), .B(n12954), .Z(n13059) );
  AND U13244 ( .A(n13060), .B(n13061), .Z(n12954) );
  NANDN U13245 ( .A(n13062), .B(n13063), .Z(n13061) );
  NAND U13246 ( .A(n13064), .B(n13065), .Z(n13063) );
  ANDN U13247 ( .B(B[210]), .A(n41), .Z(n12956) );
  XOR U13248 ( .A(n12963), .B(n13066), .Z(n12957) );
  XNOR U13249 ( .A(n12961), .B(n12964), .Z(n13066) );
  NAND U13250 ( .A(A[2]), .B(B[211]), .Z(n12964) );
  NANDN U13251 ( .A(n13067), .B(n13068), .Z(n12961) );
  AND U13252 ( .A(A[0]), .B(B[212]), .Z(n13068) );
  XNOR U13253 ( .A(n12966), .B(n13069), .Z(n12963) );
  NAND U13254 ( .A(A[0]), .B(B[213]), .Z(n13069) );
  NAND U13255 ( .A(B[212]), .B(A[1]), .Z(n12966) );
  NAND U13256 ( .A(n13070), .B(n13071), .Z(n317) );
  NANDN U13257 ( .A(n13072), .B(n13073), .Z(n13071) );
  OR U13258 ( .A(n13074), .B(n13075), .Z(n13073) );
  NAND U13259 ( .A(n13075), .B(n13074), .Z(n13070) );
  XOR U13260 ( .A(n319), .B(n318), .Z(\A1[210] ) );
  XOR U13261 ( .A(n13075), .B(n13076), .Z(n318) );
  XNOR U13262 ( .A(n13074), .B(n13072), .Z(n13076) );
  AND U13263 ( .A(n13077), .B(n13078), .Z(n13072) );
  NANDN U13264 ( .A(n13079), .B(n13080), .Z(n13078) );
  NANDN U13265 ( .A(n13081), .B(n13082), .Z(n13080) );
  NANDN U13266 ( .A(n13082), .B(n13081), .Z(n13077) );
  ANDN U13267 ( .B(B[197]), .A(n29), .Z(n13074) );
  XNOR U13268 ( .A(n12981), .B(n13083), .Z(n13075) );
  XNOR U13269 ( .A(n12980), .B(n12978), .Z(n13083) );
  AND U13270 ( .A(n13084), .B(n13085), .Z(n12978) );
  NANDN U13271 ( .A(n13086), .B(n13087), .Z(n13085) );
  OR U13272 ( .A(n13088), .B(n13089), .Z(n13087) );
  NAND U13273 ( .A(n13089), .B(n13088), .Z(n13084) );
  ANDN U13274 ( .B(B[198]), .A(n30), .Z(n12980) );
  XNOR U13275 ( .A(n12988), .B(n13090), .Z(n12981) );
  XNOR U13276 ( .A(n12987), .B(n12985), .Z(n13090) );
  AND U13277 ( .A(n13091), .B(n13092), .Z(n12985) );
  NANDN U13278 ( .A(n13093), .B(n13094), .Z(n13092) );
  NANDN U13279 ( .A(n13095), .B(n13096), .Z(n13094) );
  NANDN U13280 ( .A(n13096), .B(n13095), .Z(n13091) );
  ANDN U13281 ( .B(B[199]), .A(n31), .Z(n12987) );
  XNOR U13282 ( .A(n12995), .B(n13097), .Z(n12988) );
  XNOR U13283 ( .A(n12994), .B(n12992), .Z(n13097) );
  AND U13284 ( .A(n13098), .B(n13099), .Z(n12992) );
  NANDN U13285 ( .A(n13100), .B(n13101), .Z(n13099) );
  OR U13286 ( .A(n13102), .B(n13103), .Z(n13101) );
  NAND U13287 ( .A(n13103), .B(n13102), .Z(n13098) );
  ANDN U13288 ( .B(B[200]), .A(n32), .Z(n12994) );
  XNOR U13289 ( .A(n13002), .B(n13104), .Z(n12995) );
  XNOR U13290 ( .A(n13001), .B(n12999), .Z(n13104) );
  AND U13291 ( .A(n13105), .B(n13106), .Z(n12999) );
  NANDN U13292 ( .A(n13107), .B(n13108), .Z(n13106) );
  NANDN U13293 ( .A(n13109), .B(n13110), .Z(n13108) );
  NANDN U13294 ( .A(n13110), .B(n13109), .Z(n13105) );
  ANDN U13295 ( .B(B[201]), .A(n33), .Z(n13001) );
  XNOR U13296 ( .A(n13009), .B(n13111), .Z(n13002) );
  XNOR U13297 ( .A(n13008), .B(n13006), .Z(n13111) );
  AND U13298 ( .A(n13112), .B(n13113), .Z(n13006) );
  NANDN U13299 ( .A(n13114), .B(n13115), .Z(n13113) );
  OR U13300 ( .A(n13116), .B(n13117), .Z(n13115) );
  NAND U13301 ( .A(n13117), .B(n13116), .Z(n13112) );
  ANDN U13302 ( .B(B[202]), .A(n34), .Z(n13008) );
  XNOR U13303 ( .A(n13016), .B(n13118), .Z(n13009) );
  XNOR U13304 ( .A(n13015), .B(n13013), .Z(n13118) );
  AND U13305 ( .A(n13119), .B(n13120), .Z(n13013) );
  NANDN U13306 ( .A(n13121), .B(n13122), .Z(n13120) );
  NANDN U13307 ( .A(n13123), .B(n13124), .Z(n13122) );
  NANDN U13308 ( .A(n13124), .B(n13123), .Z(n13119) );
  ANDN U13309 ( .B(B[203]), .A(n35), .Z(n13015) );
  XNOR U13310 ( .A(n13023), .B(n13125), .Z(n13016) );
  XNOR U13311 ( .A(n13022), .B(n13020), .Z(n13125) );
  AND U13312 ( .A(n13126), .B(n13127), .Z(n13020) );
  NANDN U13313 ( .A(n13128), .B(n13129), .Z(n13127) );
  OR U13314 ( .A(n13130), .B(n13131), .Z(n13129) );
  NAND U13315 ( .A(n13131), .B(n13130), .Z(n13126) );
  ANDN U13316 ( .B(B[204]), .A(n36), .Z(n13022) );
  XNOR U13317 ( .A(n13030), .B(n13132), .Z(n13023) );
  XNOR U13318 ( .A(n13029), .B(n13027), .Z(n13132) );
  AND U13319 ( .A(n13133), .B(n13134), .Z(n13027) );
  NANDN U13320 ( .A(n13135), .B(n13136), .Z(n13134) );
  NANDN U13321 ( .A(n13137), .B(n13138), .Z(n13136) );
  NANDN U13322 ( .A(n13138), .B(n13137), .Z(n13133) );
  ANDN U13323 ( .B(B[205]), .A(n37), .Z(n13029) );
  XNOR U13324 ( .A(n13037), .B(n13139), .Z(n13030) );
  XNOR U13325 ( .A(n13036), .B(n13034), .Z(n13139) );
  AND U13326 ( .A(n13140), .B(n13141), .Z(n13034) );
  NANDN U13327 ( .A(n13142), .B(n13143), .Z(n13141) );
  OR U13328 ( .A(n13144), .B(n13145), .Z(n13143) );
  NAND U13329 ( .A(n13145), .B(n13144), .Z(n13140) );
  ANDN U13330 ( .B(B[206]), .A(n38), .Z(n13036) );
  XNOR U13331 ( .A(n13044), .B(n13146), .Z(n13037) );
  XNOR U13332 ( .A(n13043), .B(n13041), .Z(n13146) );
  AND U13333 ( .A(n13147), .B(n13148), .Z(n13041) );
  NANDN U13334 ( .A(n13149), .B(n13150), .Z(n13148) );
  NANDN U13335 ( .A(n13151), .B(n13152), .Z(n13150) );
  NANDN U13336 ( .A(n13152), .B(n13151), .Z(n13147) );
  ANDN U13337 ( .B(B[207]), .A(n39), .Z(n13043) );
  XNOR U13338 ( .A(n13051), .B(n13153), .Z(n13044) );
  XNOR U13339 ( .A(n13050), .B(n13048), .Z(n13153) );
  AND U13340 ( .A(n13154), .B(n13155), .Z(n13048) );
  NANDN U13341 ( .A(n13156), .B(n13157), .Z(n13155) );
  OR U13342 ( .A(n13158), .B(n13159), .Z(n13157) );
  NAND U13343 ( .A(n13159), .B(n13158), .Z(n13154) );
  ANDN U13344 ( .B(B[208]), .A(n40), .Z(n13050) );
  XNOR U13345 ( .A(n13058), .B(n13160), .Z(n13051) );
  XNOR U13346 ( .A(n13057), .B(n13055), .Z(n13160) );
  AND U13347 ( .A(n13161), .B(n13162), .Z(n13055) );
  NANDN U13348 ( .A(n13163), .B(n13164), .Z(n13162) );
  NAND U13349 ( .A(n13165), .B(n13166), .Z(n13164) );
  ANDN U13350 ( .B(B[209]), .A(n41), .Z(n13057) );
  XOR U13351 ( .A(n13064), .B(n13167), .Z(n13058) );
  XNOR U13352 ( .A(n13062), .B(n13065), .Z(n13167) );
  NAND U13353 ( .A(A[2]), .B(B[210]), .Z(n13065) );
  NANDN U13354 ( .A(n13168), .B(n13169), .Z(n13062) );
  AND U13355 ( .A(A[0]), .B(B[211]), .Z(n13169) );
  XNOR U13356 ( .A(n13067), .B(n13170), .Z(n13064) );
  NAND U13357 ( .A(A[0]), .B(B[212]), .Z(n13170) );
  NAND U13358 ( .A(B[211]), .B(A[1]), .Z(n13067) );
  NAND U13359 ( .A(n13171), .B(n13172), .Z(n319) );
  NANDN U13360 ( .A(n13173), .B(n13174), .Z(n13172) );
  OR U13361 ( .A(n13175), .B(n13176), .Z(n13174) );
  NAND U13362 ( .A(n13176), .B(n13175), .Z(n13171) );
  XOR U13363 ( .A(n301), .B(n300), .Z(\A1[20] ) );
  XOR U13364 ( .A(n12166), .B(n13177), .Z(n300) );
  XNOR U13365 ( .A(n12165), .B(n12163), .Z(n13177) );
  AND U13366 ( .A(n13178), .B(n13179), .Z(n12163) );
  NANDN U13367 ( .A(n13180), .B(n13181), .Z(n13179) );
  NANDN U13368 ( .A(n13182), .B(n13183), .Z(n13181) );
  NANDN U13369 ( .A(n13183), .B(n13182), .Z(n13178) );
  ANDN U13370 ( .B(B[7]), .A(n29), .Z(n12165) );
  XNOR U13371 ( .A(n12072), .B(n13184), .Z(n12166) );
  XNOR U13372 ( .A(n12071), .B(n12069), .Z(n13184) );
  AND U13373 ( .A(n13185), .B(n13186), .Z(n12069) );
  NANDN U13374 ( .A(n13187), .B(n13188), .Z(n13186) );
  OR U13375 ( .A(n13189), .B(n13190), .Z(n13188) );
  NAND U13376 ( .A(n13190), .B(n13189), .Z(n13185) );
  ANDN U13377 ( .B(B[8]), .A(n30), .Z(n12071) );
  XNOR U13378 ( .A(n12079), .B(n13191), .Z(n12072) );
  XNOR U13379 ( .A(n12078), .B(n12076), .Z(n13191) );
  AND U13380 ( .A(n13192), .B(n13193), .Z(n12076) );
  NANDN U13381 ( .A(n13194), .B(n13195), .Z(n13193) );
  NANDN U13382 ( .A(n13196), .B(n13197), .Z(n13195) );
  NANDN U13383 ( .A(n13197), .B(n13196), .Z(n13192) );
  ANDN U13384 ( .B(B[9]), .A(n31), .Z(n12078) );
  XNOR U13385 ( .A(n12086), .B(n13198), .Z(n12079) );
  XNOR U13386 ( .A(n12085), .B(n12083), .Z(n13198) );
  AND U13387 ( .A(n13199), .B(n13200), .Z(n12083) );
  NANDN U13388 ( .A(n13201), .B(n13202), .Z(n13200) );
  OR U13389 ( .A(n13203), .B(n13204), .Z(n13202) );
  NAND U13390 ( .A(n13204), .B(n13203), .Z(n13199) );
  ANDN U13391 ( .B(B[10]), .A(n32), .Z(n12085) );
  XNOR U13392 ( .A(n12093), .B(n13205), .Z(n12086) );
  XNOR U13393 ( .A(n12092), .B(n12090), .Z(n13205) );
  AND U13394 ( .A(n13206), .B(n13207), .Z(n12090) );
  NANDN U13395 ( .A(n13208), .B(n13209), .Z(n13207) );
  NANDN U13396 ( .A(n13210), .B(n13211), .Z(n13209) );
  NANDN U13397 ( .A(n13211), .B(n13210), .Z(n13206) );
  ANDN U13398 ( .B(B[11]), .A(n33), .Z(n12092) );
  XNOR U13399 ( .A(n12100), .B(n13212), .Z(n12093) );
  XNOR U13400 ( .A(n12099), .B(n12097), .Z(n13212) );
  AND U13401 ( .A(n13213), .B(n13214), .Z(n12097) );
  NANDN U13402 ( .A(n13215), .B(n13216), .Z(n13214) );
  OR U13403 ( .A(n13217), .B(n13218), .Z(n13216) );
  NAND U13404 ( .A(n13218), .B(n13217), .Z(n13213) );
  ANDN U13405 ( .B(B[12]), .A(n34), .Z(n12099) );
  XNOR U13406 ( .A(n12107), .B(n13219), .Z(n12100) );
  XNOR U13407 ( .A(n12106), .B(n12104), .Z(n13219) );
  AND U13408 ( .A(n13220), .B(n13221), .Z(n12104) );
  NANDN U13409 ( .A(n13222), .B(n13223), .Z(n13221) );
  NANDN U13410 ( .A(n13224), .B(n13225), .Z(n13223) );
  NANDN U13411 ( .A(n13225), .B(n13224), .Z(n13220) );
  ANDN U13412 ( .B(B[13]), .A(n35), .Z(n12106) );
  XNOR U13413 ( .A(n12114), .B(n13226), .Z(n12107) );
  XNOR U13414 ( .A(n12113), .B(n12111), .Z(n13226) );
  AND U13415 ( .A(n13227), .B(n13228), .Z(n12111) );
  NANDN U13416 ( .A(n13229), .B(n13230), .Z(n13228) );
  OR U13417 ( .A(n13231), .B(n13232), .Z(n13230) );
  NAND U13418 ( .A(n13232), .B(n13231), .Z(n13227) );
  ANDN U13419 ( .B(B[14]), .A(n36), .Z(n12113) );
  XNOR U13420 ( .A(n12121), .B(n13233), .Z(n12114) );
  XNOR U13421 ( .A(n12120), .B(n12118), .Z(n13233) );
  AND U13422 ( .A(n13234), .B(n13235), .Z(n12118) );
  NANDN U13423 ( .A(n13236), .B(n13237), .Z(n13235) );
  NANDN U13424 ( .A(n13238), .B(n13239), .Z(n13237) );
  NANDN U13425 ( .A(n13239), .B(n13238), .Z(n13234) );
  ANDN U13426 ( .B(B[15]), .A(n37), .Z(n12120) );
  XNOR U13427 ( .A(n12128), .B(n13240), .Z(n12121) );
  XNOR U13428 ( .A(n12127), .B(n12125), .Z(n13240) );
  AND U13429 ( .A(n13241), .B(n13242), .Z(n12125) );
  NANDN U13430 ( .A(n13243), .B(n13244), .Z(n13242) );
  OR U13431 ( .A(n13245), .B(n13246), .Z(n13244) );
  NAND U13432 ( .A(n13246), .B(n13245), .Z(n13241) );
  ANDN U13433 ( .B(B[16]), .A(n38), .Z(n12127) );
  XNOR U13434 ( .A(n12135), .B(n13247), .Z(n12128) );
  XNOR U13435 ( .A(n12134), .B(n12132), .Z(n13247) );
  AND U13436 ( .A(n13248), .B(n13249), .Z(n12132) );
  NANDN U13437 ( .A(n13250), .B(n13251), .Z(n13249) );
  NANDN U13438 ( .A(n13252), .B(n13253), .Z(n13251) );
  NANDN U13439 ( .A(n13253), .B(n13252), .Z(n13248) );
  ANDN U13440 ( .B(B[17]), .A(n39), .Z(n12134) );
  XNOR U13441 ( .A(n12142), .B(n13254), .Z(n12135) );
  XNOR U13442 ( .A(n12141), .B(n12139), .Z(n13254) );
  AND U13443 ( .A(n13255), .B(n13256), .Z(n12139) );
  NANDN U13444 ( .A(n13257), .B(n13258), .Z(n13256) );
  OR U13445 ( .A(n13259), .B(n13260), .Z(n13258) );
  NAND U13446 ( .A(n13260), .B(n13259), .Z(n13255) );
  ANDN U13447 ( .B(B[18]), .A(n40), .Z(n12141) );
  XNOR U13448 ( .A(n12149), .B(n13261), .Z(n12142) );
  XNOR U13449 ( .A(n12148), .B(n12146), .Z(n13261) );
  AND U13450 ( .A(n13262), .B(n13263), .Z(n12146) );
  NANDN U13451 ( .A(n13264), .B(n13265), .Z(n13263) );
  NAND U13452 ( .A(n13266), .B(n13267), .Z(n13265) );
  ANDN U13453 ( .B(B[19]), .A(n41), .Z(n12148) );
  XOR U13454 ( .A(n12155), .B(n13268), .Z(n12149) );
  XNOR U13455 ( .A(n12153), .B(n12156), .Z(n13268) );
  NAND U13456 ( .A(A[2]), .B(B[20]), .Z(n12156) );
  NANDN U13457 ( .A(n13269), .B(n13270), .Z(n12153) );
  AND U13458 ( .A(A[0]), .B(B[21]), .Z(n13270) );
  XNOR U13459 ( .A(n12158), .B(n13271), .Z(n12155) );
  NAND U13460 ( .A(A[0]), .B(B[22]), .Z(n13271) );
  NAND U13461 ( .A(B[21]), .B(A[1]), .Z(n12158) );
  NAND U13462 ( .A(n13272), .B(n13273), .Z(n301) );
  NANDN U13463 ( .A(n13274), .B(n13275), .Z(n13273) );
  OR U13464 ( .A(n13276), .B(n13277), .Z(n13275) );
  NAND U13465 ( .A(n13277), .B(n13276), .Z(n13272) );
  XOR U13466 ( .A(n321), .B(n320), .Z(\A1[209] ) );
  XOR U13467 ( .A(n13176), .B(n13278), .Z(n320) );
  XNOR U13468 ( .A(n13175), .B(n13173), .Z(n13278) );
  AND U13469 ( .A(n13279), .B(n13280), .Z(n13173) );
  NANDN U13470 ( .A(n13281), .B(n13282), .Z(n13280) );
  NANDN U13471 ( .A(n13283), .B(n13284), .Z(n13282) );
  NANDN U13472 ( .A(n13284), .B(n13283), .Z(n13279) );
  ANDN U13473 ( .B(B[196]), .A(n29), .Z(n13175) );
  XNOR U13474 ( .A(n13082), .B(n13285), .Z(n13176) );
  XNOR U13475 ( .A(n13081), .B(n13079), .Z(n13285) );
  AND U13476 ( .A(n13286), .B(n13287), .Z(n13079) );
  NANDN U13477 ( .A(n13288), .B(n13289), .Z(n13287) );
  OR U13478 ( .A(n13290), .B(n13291), .Z(n13289) );
  NAND U13479 ( .A(n13291), .B(n13290), .Z(n13286) );
  ANDN U13480 ( .B(B[197]), .A(n30), .Z(n13081) );
  XNOR U13481 ( .A(n13089), .B(n13292), .Z(n13082) );
  XNOR U13482 ( .A(n13088), .B(n13086), .Z(n13292) );
  AND U13483 ( .A(n13293), .B(n13294), .Z(n13086) );
  NANDN U13484 ( .A(n13295), .B(n13296), .Z(n13294) );
  NANDN U13485 ( .A(n13297), .B(n13298), .Z(n13296) );
  NANDN U13486 ( .A(n13298), .B(n13297), .Z(n13293) );
  ANDN U13487 ( .B(B[198]), .A(n31), .Z(n13088) );
  XNOR U13488 ( .A(n13096), .B(n13299), .Z(n13089) );
  XNOR U13489 ( .A(n13095), .B(n13093), .Z(n13299) );
  AND U13490 ( .A(n13300), .B(n13301), .Z(n13093) );
  NANDN U13491 ( .A(n13302), .B(n13303), .Z(n13301) );
  OR U13492 ( .A(n13304), .B(n13305), .Z(n13303) );
  NAND U13493 ( .A(n13305), .B(n13304), .Z(n13300) );
  ANDN U13494 ( .B(B[199]), .A(n32), .Z(n13095) );
  XNOR U13495 ( .A(n13103), .B(n13306), .Z(n13096) );
  XNOR U13496 ( .A(n13102), .B(n13100), .Z(n13306) );
  AND U13497 ( .A(n13307), .B(n13308), .Z(n13100) );
  NANDN U13498 ( .A(n13309), .B(n13310), .Z(n13308) );
  NANDN U13499 ( .A(n13311), .B(n13312), .Z(n13310) );
  NANDN U13500 ( .A(n13312), .B(n13311), .Z(n13307) );
  ANDN U13501 ( .B(B[200]), .A(n33), .Z(n13102) );
  XNOR U13502 ( .A(n13110), .B(n13313), .Z(n13103) );
  XNOR U13503 ( .A(n13109), .B(n13107), .Z(n13313) );
  AND U13504 ( .A(n13314), .B(n13315), .Z(n13107) );
  NANDN U13505 ( .A(n13316), .B(n13317), .Z(n13315) );
  OR U13506 ( .A(n13318), .B(n13319), .Z(n13317) );
  NAND U13507 ( .A(n13319), .B(n13318), .Z(n13314) );
  ANDN U13508 ( .B(B[201]), .A(n34), .Z(n13109) );
  XNOR U13509 ( .A(n13117), .B(n13320), .Z(n13110) );
  XNOR U13510 ( .A(n13116), .B(n13114), .Z(n13320) );
  AND U13511 ( .A(n13321), .B(n13322), .Z(n13114) );
  NANDN U13512 ( .A(n13323), .B(n13324), .Z(n13322) );
  NANDN U13513 ( .A(n13325), .B(n13326), .Z(n13324) );
  NANDN U13514 ( .A(n13326), .B(n13325), .Z(n13321) );
  ANDN U13515 ( .B(B[202]), .A(n35), .Z(n13116) );
  XNOR U13516 ( .A(n13124), .B(n13327), .Z(n13117) );
  XNOR U13517 ( .A(n13123), .B(n13121), .Z(n13327) );
  AND U13518 ( .A(n13328), .B(n13329), .Z(n13121) );
  NANDN U13519 ( .A(n13330), .B(n13331), .Z(n13329) );
  OR U13520 ( .A(n13332), .B(n13333), .Z(n13331) );
  NAND U13521 ( .A(n13333), .B(n13332), .Z(n13328) );
  ANDN U13522 ( .B(B[203]), .A(n36), .Z(n13123) );
  XNOR U13523 ( .A(n13131), .B(n13334), .Z(n13124) );
  XNOR U13524 ( .A(n13130), .B(n13128), .Z(n13334) );
  AND U13525 ( .A(n13335), .B(n13336), .Z(n13128) );
  NANDN U13526 ( .A(n13337), .B(n13338), .Z(n13336) );
  NANDN U13527 ( .A(n13339), .B(n13340), .Z(n13338) );
  NANDN U13528 ( .A(n13340), .B(n13339), .Z(n13335) );
  ANDN U13529 ( .B(B[204]), .A(n37), .Z(n13130) );
  XNOR U13530 ( .A(n13138), .B(n13341), .Z(n13131) );
  XNOR U13531 ( .A(n13137), .B(n13135), .Z(n13341) );
  AND U13532 ( .A(n13342), .B(n13343), .Z(n13135) );
  NANDN U13533 ( .A(n13344), .B(n13345), .Z(n13343) );
  OR U13534 ( .A(n13346), .B(n13347), .Z(n13345) );
  NAND U13535 ( .A(n13347), .B(n13346), .Z(n13342) );
  ANDN U13536 ( .B(B[205]), .A(n38), .Z(n13137) );
  XNOR U13537 ( .A(n13145), .B(n13348), .Z(n13138) );
  XNOR U13538 ( .A(n13144), .B(n13142), .Z(n13348) );
  AND U13539 ( .A(n13349), .B(n13350), .Z(n13142) );
  NANDN U13540 ( .A(n13351), .B(n13352), .Z(n13350) );
  NANDN U13541 ( .A(n13353), .B(n13354), .Z(n13352) );
  NANDN U13542 ( .A(n13354), .B(n13353), .Z(n13349) );
  ANDN U13543 ( .B(B[206]), .A(n39), .Z(n13144) );
  XNOR U13544 ( .A(n13152), .B(n13355), .Z(n13145) );
  XNOR U13545 ( .A(n13151), .B(n13149), .Z(n13355) );
  AND U13546 ( .A(n13356), .B(n13357), .Z(n13149) );
  NANDN U13547 ( .A(n13358), .B(n13359), .Z(n13357) );
  OR U13548 ( .A(n13360), .B(n13361), .Z(n13359) );
  NAND U13549 ( .A(n13361), .B(n13360), .Z(n13356) );
  ANDN U13550 ( .B(B[207]), .A(n40), .Z(n13151) );
  XNOR U13551 ( .A(n13159), .B(n13362), .Z(n13152) );
  XNOR U13552 ( .A(n13158), .B(n13156), .Z(n13362) );
  AND U13553 ( .A(n13363), .B(n13364), .Z(n13156) );
  NANDN U13554 ( .A(n13365), .B(n13366), .Z(n13364) );
  NAND U13555 ( .A(n13367), .B(n13368), .Z(n13366) );
  ANDN U13556 ( .B(B[208]), .A(n41), .Z(n13158) );
  XOR U13557 ( .A(n13165), .B(n13369), .Z(n13159) );
  XNOR U13558 ( .A(n13163), .B(n13166), .Z(n13369) );
  NAND U13559 ( .A(A[2]), .B(B[209]), .Z(n13166) );
  NANDN U13560 ( .A(n13370), .B(n13371), .Z(n13163) );
  AND U13561 ( .A(A[0]), .B(B[210]), .Z(n13371) );
  XNOR U13562 ( .A(n13168), .B(n13372), .Z(n13165) );
  NAND U13563 ( .A(A[0]), .B(B[211]), .Z(n13372) );
  NAND U13564 ( .A(B[210]), .B(A[1]), .Z(n13168) );
  NAND U13565 ( .A(n13373), .B(n13374), .Z(n321) );
  NANDN U13566 ( .A(n13375), .B(n13376), .Z(n13374) );
  OR U13567 ( .A(n13377), .B(n13378), .Z(n13376) );
  NAND U13568 ( .A(n13378), .B(n13377), .Z(n13373) );
  XOR U13569 ( .A(n325), .B(n324), .Z(\A1[208] ) );
  XOR U13570 ( .A(n13378), .B(n13379), .Z(n324) );
  XNOR U13571 ( .A(n13377), .B(n13375), .Z(n13379) );
  AND U13572 ( .A(n13380), .B(n13381), .Z(n13375) );
  NANDN U13573 ( .A(n13382), .B(n13383), .Z(n13381) );
  NANDN U13574 ( .A(n13384), .B(n13385), .Z(n13383) );
  NANDN U13575 ( .A(n13385), .B(n13384), .Z(n13380) );
  ANDN U13576 ( .B(B[195]), .A(n29), .Z(n13377) );
  XNOR U13577 ( .A(n13284), .B(n13386), .Z(n13378) );
  XNOR U13578 ( .A(n13283), .B(n13281), .Z(n13386) );
  AND U13579 ( .A(n13387), .B(n13388), .Z(n13281) );
  NANDN U13580 ( .A(n13389), .B(n13390), .Z(n13388) );
  OR U13581 ( .A(n13391), .B(n13392), .Z(n13390) );
  NAND U13582 ( .A(n13392), .B(n13391), .Z(n13387) );
  ANDN U13583 ( .B(B[196]), .A(n30), .Z(n13283) );
  XNOR U13584 ( .A(n13291), .B(n13393), .Z(n13284) );
  XNOR U13585 ( .A(n13290), .B(n13288), .Z(n13393) );
  AND U13586 ( .A(n13394), .B(n13395), .Z(n13288) );
  NANDN U13587 ( .A(n13396), .B(n13397), .Z(n13395) );
  NANDN U13588 ( .A(n13398), .B(n13399), .Z(n13397) );
  NANDN U13589 ( .A(n13399), .B(n13398), .Z(n13394) );
  ANDN U13590 ( .B(B[197]), .A(n31), .Z(n13290) );
  XNOR U13591 ( .A(n13298), .B(n13400), .Z(n13291) );
  XNOR U13592 ( .A(n13297), .B(n13295), .Z(n13400) );
  AND U13593 ( .A(n13401), .B(n13402), .Z(n13295) );
  NANDN U13594 ( .A(n13403), .B(n13404), .Z(n13402) );
  OR U13595 ( .A(n13405), .B(n13406), .Z(n13404) );
  NAND U13596 ( .A(n13406), .B(n13405), .Z(n13401) );
  ANDN U13597 ( .B(B[198]), .A(n32), .Z(n13297) );
  XNOR U13598 ( .A(n13305), .B(n13407), .Z(n13298) );
  XNOR U13599 ( .A(n13304), .B(n13302), .Z(n13407) );
  AND U13600 ( .A(n13408), .B(n13409), .Z(n13302) );
  NANDN U13601 ( .A(n13410), .B(n13411), .Z(n13409) );
  NANDN U13602 ( .A(n13412), .B(n13413), .Z(n13411) );
  NANDN U13603 ( .A(n13413), .B(n13412), .Z(n13408) );
  ANDN U13604 ( .B(B[199]), .A(n33), .Z(n13304) );
  XNOR U13605 ( .A(n13312), .B(n13414), .Z(n13305) );
  XNOR U13606 ( .A(n13311), .B(n13309), .Z(n13414) );
  AND U13607 ( .A(n13415), .B(n13416), .Z(n13309) );
  NANDN U13608 ( .A(n13417), .B(n13418), .Z(n13416) );
  OR U13609 ( .A(n13419), .B(n13420), .Z(n13418) );
  NAND U13610 ( .A(n13420), .B(n13419), .Z(n13415) );
  ANDN U13611 ( .B(B[200]), .A(n34), .Z(n13311) );
  XNOR U13612 ( .A(n13319), .B(n13421), .Z(n13312) );
  XNOR U13613 ( .A(n13318), .B(n13316), .Z(n13421) );
  AND U13614 ( .A(n13422), .B(n13423), .Z(n13316) );
  NANDN U13615 ( .A(n13424), .B(n13425), .Z(n13423) );
  NANDN U13616 ( .A(n13426), .B(n13427), .Z(n13425) );
  NANDN U13617 ( .A(n13427), .B(n13426), .Z(n13422) );
  ANDN U13618 ( .B(B[201]), .A(n35), .Z(n13318) );
  XNOR U13619 ( .A(n13326), .B(n13428), .Z(n13319) );
  XNOR U13620 ( .A(n13325), .B(n13323), .Z(n13428) );
  AND U13621 ( .A(n13429), .B(n13430), .Z(n13323) );
  NANDN U13622 ( .A(n13431), .B(n13432), .Z(n13430) );
  OR U13623 ( .A(n13433), .B(n13434), .Z(n13432) );
  NAND U13624 ( .A(n13434), .B(n13433), .Z(n13429) );
  ANDN U13625 ( .B(B[202]), .A(n36), .Z(n13325) );
  XNOR U13626 ( .A(n13333), .B(n13435), .Z(n13326) );
  XNOR U13627 ( .A(n13332), .B(n13330), .Z(n13435) );
  AND U13628 ( .A(n13436), .B(n13437), .Z(n13330) );
  NANDN U13629 ( .A(n13438), .B(n13439), .Z(n13437) );
  NANDN U13630 ( .A(n13440), .B(n13441), .Z(n13439) );
  NANDN U13631 ( .A(n13441), .B(n13440), .Z(n13436) );
  ANDN U13632 ( .B(B[203]), .A(n37), .Z(n13332) );
  XNOR U13633 ( .A(n13340), .B(n13442), .Z(n13333) );
  XNOR U13634 ( .A(n13339), .B(n13337), .Z(n13442) );
  AND U13635 ( .A(n13443), .B(n13444), .Z(n13337) );
  NANDN U13636 ( .A(n13445), .B(n13446), .Z(n13444) );
  OR U13637 ( .A(n13447), .B(n13448), .Z(n13446) );
  NAND U13638 ( .A(n13448), .B(n13447), .Z(n13443) );
  ANDN U13639 ( .B(B[204]), .A(n38), .Z(n13339) );
  XNOR U13640 ( .A(n13347), .B(n13449), .Z(n13340) );
  XNOR U13641 ( .A(n13346), .B(n13344), .Z(n13449) );
  AND U13642 ( .A(n13450), .B(n13451), .Z(n13344) );
  NANDN U13643 ( .A(n13452), .B(n13453), .Z(n13451) );
  NANDN U13644 ( .A(n13454), .B(n13455), .Z(n13453) );
  NANDN U13645 ( .A(n13455), .B(n13454), .Z(n13450) );
  ANDN U13646 ( .B(B[205]), .A(n39), .Z(n13346) );
  XNOR U13647 ( .A(n13354), .B(n13456), .Z(n13347) );
  XNOR U13648 ( .A(n13353), .B(n13351), .Z(n13456) );
  AND U13649 ( .A(n13457), .B(n13458), .Z(n13351) );
  NANDN U13650 ( .A(n13459), .B(n13460), .Z(n13458) );
  OR U13651 ( .A(n13461), .B(n13462), .Z(n13460) );
  NAND U13652 ( .A(n13462), .B(n13461), .Z(n13457) );
  ANDN U13653 ( .B(B[206]), .A(n40), .Z(n13353) );
  XNOR U13654 ( .A(n13361), .B(n13463), .Z(n13354) );
  XNOR U13655 ( .A(n13360), .B(n13358), .Z(n13463) );
  AND U13656 ( .A(n13464), .B(n13465), .Z(n13358) );
  NANDN U13657 ( .A(n13466), .B(n13467), .Z(n13465) );
  NAND U13658 ( .A(n13468), .B(n13469), .Z(n13467) );
  ANDN U13659 ( .B(B[207]), .A(n41), .Z(n13360) );
  XOR U13660 ( .A(n13367), .B(n13470), .Z(n13361) );
  XNOR U13661 ( .A(n13365), .B(n13368), .Z(n13470) );
  NAND U13662 ( .A(A[2]), .B(B[208]), .Z(n13368) );
  NANDN U13663 ( .A(n13471), .B(n13472), .Z(n13365) );
  AND U13664 ( .A(A[0]), .B(B[209]), .Z(n13472) );
  XNOR U13665 ( .A(n13370), .B(n13473), .Z(n13367) );
  NAND U13666 ( .A(A[0]), .B(B[210]), .Z(n13473) );
  NAND U13667 ( .A(B[209]), .B(A[1]), .Z(n13370) );
  NAND U13668 ( .A(n13474), .B(n13475), .Z(n325) );
  NANDN U13669 ( .A(n13476), .B(n13477), .Z(n13475) );
  OR U13670 ( .A(n13478), .B(n13479), .Z(n13477) );
  NAND U13671 ( .A(n13479), .B(n13478), .Z(n13474) );
  XOR U13672 ( .A(n327), .B(n326), .Z(\A1[207] ) );
  XOR U13673 ( .A(n13479), .B(n13480), .Z(n326) );
  XNOR U13674 ( .A(n13478), .B(n13476), .Z(n13480) );
  AND U13675 ( .A(n13481), .B(n13482), .Z(n13476) );
  NANDN U13676 ( .A(n13483), .B(n13484), .Z(n13482) );
  NANDN U13677 ( .A(n13485), .B(n13486), .Z(n13484) );
  NANDN U13678 ( .A(n13486), .B(n13485), .Z(n13481) );
  ANDN U13679 ( .B(B[194]), .A(n29), .Z(n13478) );
  XNOR U13680 ( .A(n13385), .B(n13487), .Z(n13479) );
  XNOR U13681 ( .A(n13384), .B(n13382), .Z(n13487) );
  AND U13682 ( .A(n13488), .B(n13489), .Z(n13382) );
  NANDN U13683 ( .A(n13490), .B(n13491), .Z(n13489) );
  OR U13684 ( .A(n13492), .B(n13493), .Z(n13491) );
  NAND U13685 ( .A(n13493), .B(n13492), .Z(n13488) );
  ANDN U13686 ( .B(B[195]), .A(n30), .Z(n13384) );
  XNOR U13687 ( .A(n13392), .B(n13494), .Z(n13385) );
  XNOR U13688 ( .A(n13391), .B(n13389), .Z(n13494) );
  AND U13689 ( .A(n13495), .B(n13496), .Z(n13389) );
  NANDN U13690 ( .A(n13497), .B(n13498), .Z(n13496) );
  NANDN U13691 ( .A(n13499), .B(n13500), .Z(n13498) );
  NANDN U13692 ( .A(n13500), .B(n13499), .Z(n13495) );
  ANDN U13693 ( .B(B[196]), .A(n31), .Z(n13391) );
  XNOR U13694 ( .A(n13399), .B(n13501), .Z(n13392) );
  XNOR U13695 ( .A(n13398), .B(n13396), .Z(n13501) );
  AND U13696 ( .A(n13502), .B(n13503), .Z(n13396) );
  NANDN U13697 ( .A(n13504), .B(n13505), .Z(n13503) );
  OR U13698 ( .A(n13506), .B(n13507), .Z(n13505) );
  NAND U13699 ( .A(n13507), .B(n13506), .Z(n13502) );
  ANDN U13700 ( .B(B[197]), .A(n32), .Z(n13398) );
  XNOR U13701 ( .A(n13406), .B(n13508), .Z(n13399) );
  XNOR U13702 ( .A(n13405), .B(n13403), .Z(n13508) );
  AND U13703 ( .A(n13509), .B(n13510), .Z(n13403) );
  NANDN U13704 ( .A(n13511), .B(n13512), .Z(n13510) );
  NANDN U13705 ( .A(n13513), .B(n13514), .Z(n13512) );
  NANDN U13706 ( .A(n13514), .B(n13513), .Z(n13509) );
  ANDN U13707 ( .B(B[198]), .A(n33), .Z(n13405) );
  XNOR U13708 ( .A(n13413), .B(n13515), .Z(n13406) );
  XNOR U13709 ( .A(n13412), .B(n13410), .Z(n13515) );
  AND U13710 ( .A(n13516), .B(n13517), .Z(n13410) );
  NANDN U13711 ( .A(n13518), .B(n13519), .Z(n13517) );
  OR U13712 ( .A(n13520), .B(n13521), .Z(n13519) );
  NAND U13713 ( .A(n13521), .B(n13520), .Z(n13516) );
  ANDN U13714 ( .B(B[199]), .A(n34), .Z(n13412) );
  XNOR U13715 ( .A(n13420), .B(n13522), .Z(n13413) );
  XNOR U13716 ( .A(n13419), .B(n13417), .Z(n13522) );
  AND U13717 ( .A(n13523), .B(n13524), .Z(n13417) );
  NANDN U13718 ( .A(n13525), .B(n13526), .Z(n13524) );
  NANDN U13719 ( .A(n13527), .B(n13528), .Z(n13526) );
  NANDN U13720 ( .A(n13528), .B(n13527), .Z(n13523) );
  ANDN U13721 ( .B(B[200]), .A(n35), .Z(n13419) );
  XNOR U13722 ( .A(n13427), .B(n13529), .Z(n13420) );
  XNOR U13723 ( .A(n13426), .B(n13424), .Z(n13529) );
  AND U13724 ( .A(n13530), .B(n13531), .Z(n13424) );
  NANDN U13725 ( .A(n13532), .B(n13533), .Z(n13531) );
  OR U13726 ( .A(n13534), .B(n13535), .Z(n13533) );
  NAND U13727 ( .A(n13535), .B(n13534), .Z(n13530) );
  ANDN U13728 ( .B(B[201]), .A(n36), .Z(n13426) );
  XNOR U13729 ( .A(n13434), .B(n13536), .Z(n13427) );
  XNOR U13730 ( .A(n13433), .B(n13431), .Z(n13536) );
  AND U13731 ( .A(n13537), .B(n13538), .Z(n13431) );
  NANDN U13732 ( .A(n13539), .B(n13540), .Z(n13538) );
  NANDN U13733 ( .A(n13541), .B(n13542), .Z(n13540) );
  NANDN U13734 ( .A(n13542), .B(n13541), .Z(n13537) );
  ANDN U13735 ( .B(B[202]), .A(n37), .Z(n13433) );
  XNOR U13736 ( .A(n13441), .B(n13543), .Z(n13434) );
  XNOR U13737 ( .A(n13440), .B(n13438), .Z(n13543) );
  AND U13738 ( .A(n13544), .B(n13545), .Z(n13438) );
  NANDN U13739 ( .A(n13546), .B(n13547), .Z(n13545) );
  OR U13740 ( .A(n13548), .B(n13549), .Z(n13547) );
  NAND U13741 ( .A(n13549), .B(n13548), .Z(n13544) );
  ANDN U13742 ( .B(B[203]), .A(n38), .Z(n13440) );
  XNOR U13743 ( .A(n13448), .B(n13550), .Z(n13441) );
  XNOR U13744 ( .A(n13447), .B(n13445), .Z(n13550) );
  AND U13745 ( .A(n13551), .B(n13552), .Z(n13445) );
  NANDN U13746 ( .A(n13553), .B(n13554), .Z(n13552) );
  NANDN U13747 ( .A(n13555), .B(n13556), .Z(n13554) );
  NANDN U13748 ( .A(n13556), .B(n13555), .Z(n13551) );
  ANDN U13749 ( .B(B[204]), .A(n39), .Z(n13447) );
  XNOR U13750 ( .A(n13455), .B(n13557), .Z(n13448) );
  XNOR U13751 ( .A(n13454), .B(n13452), .Z(n13557) );
  AND U13752 ( .A(n13558), .B(n13559), .Z(n13452) );
  NANDN U13753 ( .A(n13560), .B(n13561), .Z(n13559) );
  OR U13754 ( .A(n13562), .B(n13563), .Z(n13561) );
  NAND U13755 ( .A(n13563), .B(n13562), .Z(n13558) );
  ANDN U13756 ( .B(B[205]), .A(n40), .Z(n13454) );
  XNOR U13757 ( .A(n13462), .B(n13564), .Z(n13455) );
  XNOR U13758 ( .A(n13461), .B(n13459), .Z(n13564) );
  AND U13759 ( .A(n13565), .B(n13566), .Z(n13459) );
  NANDN U13760 ( .A(n13567), .B(n13568), .Z(n13566) );
  NAND U13761 ( .A(n13569), .B(n13570), .Z(n13568) );
  ANDN U13762 ( .B(B[206]), .A(n41), .Z(n13461) );
  XOR U13763 ( .A(n13468), .B(n13571), .Z(n13462) );
  XNOR U13764 ( .A(n13466), .B(n13469), .Z(n13571) );
  NAND U13765 ( .A(A[2]), .B(B[207]), .Z(n13469) );
  NANDN U13766 ( .A(n13572), .B(n13573), .Z(n13466) );
  AND U13767 ( .A(A[0]), .B(B[208]), .Z(n13573) );
  XNOR U13768 ( .A(n13471), .B(n13574), .Z(n13468) );
  NAND U13769 ( .A(A[0]), .B(B[209]), .Z(n13574) );
  NAND U13770 ( .A(B[208]), .B(A[1]), .Z(n13471) );
  NAND U13771 ( .A(n13575), .B(n13576), .Z(n327) );
  NANDN U13772 ( .A(n13577), .B(n13578), .Z(n13576) );
  OR U13773 ( .A(n13579), .B(n13580), .Z(n13578) );
  NAND U13774 ( .A(n13580), .B(n13579), .Z(n13575) );
  XOR U13775 ( .A(n329), .B(n328), .Z(\A1[206] ) );
  XOR U13776 ( .A(n13580), .B(n13581), .Z(n328) );
  XNOR U13777 ( .A(n13579), .B(n13577), .Z(n13581) );
  AND U13778 ( .A(n13582), .B(n13583), .Z(n13577) );
  NANDN U13779 ( .A(n13584), .B(n13585), .Z(n13583) );
  NANDN U13780 ( .A(n13586), .B(n13587), .Z(n13585) );
  NANDN U13781 ( .A(n13587), .B(n13586), .Z(n13582) );
  ANDN U13782 ( .B(B[193]), .A(n29), .Z(n13579) );
  XNOR U13783 ( .A(n13486), .B(n13588), .Z(n13580) );
  XNOR U13784 ( .A(n13485), .B(n13483), .Z(n13588) );
  AND U13785 ( .A(n13589), .B(n13590), .Z(n13483) );
  NANDN U13786 ( .A(n13591), .B(n13592), .Z(n13590) );
  OR U13787 ( .A(n13593), .B(n13594), .Z(n13592) );
  NAND U13788 ( .A(n13594), .B(n13593), .Z(n13589) );
  ANDN U13789 ( .B(B[194]), .A(n30), .Z(n13485) );
  XNOR U13790 ( .A(n13493), .B(n13595), .Z(n13486) );
  XNOR U13791 ( .A(n13492), .B(n13490), .Z(n13595) );
  AND U13792 ( .A(n13596), .B(n13597), .Z(n13490) );
  NANDN U13793 ( .A(n13598), .B(n13599), .Z(n13597) );
  NANDN U13794 ( .A(n13600), .B(n13601), .Z(n13599) );
  NANDN U13795 ( .A(n13601), .B(n13600), .Z(n13596) );
  ANDN U13796 ( .B(B[195]), .A(n31), .Z(n13492) );
  XNOR U13797 ( .A(n13500), .B(n13602), .Z(n13493) );
  XNOR U13798 ( .A(n13499), .B(n13497), .Z(n13602) );
  AND U13799 ( .A(n13603), .B(n13604), .Z(n13497) );
  NANDN U13800 ( .A(n13605), .B(n13606), .Z(n13604) );
  OR U13801 ( .A(n13607), .B(n13608), .Z(n13606) );
  NAND U13802 ( .A(n13608), .B(n13607), .Z(n13603) );
  ANDN U13803 ( .B(B[196]), .A(n32), .Z(n13499) );
  XNOR U13804 ( .A(n13507), .B(n13609), .Z(n13500) );
  XNOR U13805 ( .A(n13506), .B(n13504), .Z(n13609) );
  AND U13806 ( .A(n13610), .B(n13611), .Z(n13504) );
  NANDN U13807 ( .A(n13612), .B(n13613), .Z(n13611) );
  NANDN U13808 ( .A(n13614), .B(n13615), .Z(n13613) );
  NANDN U13809 ( .A(n13615), .B(n13614), .Z(n13610) );
  ANDN U13810 ( .B(B[197]), .A(n33), .Z(n13506) );
  XNOR U13811 ( .A(n13514), .B(n13616), .Z(n13507) );
  XNOR U13812 ( .A(n13513), .B(n13511), .Z(n13616) );
  AND U13813 ( .A(n13617), .B(n13618), .Z(n13511) );
  NANDN U13814 ( .A(n13619), .B(n13620), .Z(n13618) );
  OR U13815 ( .A(n13621), .B(n13622), .Z(n13620) );
  NAND U13816 ( .A(n13622), .B(n13621), .Z(n13617) );
  ANDN U13817 ( .B(B[198]), .A(n34), .Z(n13513) );
  XNOR U13818 ( .A(n13521), .B(n13623), .Z(n13514) );
  XNOR U13819 ( .A(n13520), .B(n13518), .Z(n13623) );
  AND U13820 ( .A(n13624), .B(n13625), .Z(n13518) );
  NANDN U13821 ( .A(n13626), .B(n13627), .Z(n13625) );
  NANDN U13822 ( .A(n13628), .B(n13629), .Z(n13627) );
  NANDN U13823 ( .A(n13629), .B(n13628), .Z(n13624) );
  ANDN U13824 ( .B(B[199]), .A(n35), .Z(n13520) );
  XNOR U13825 ( .A(n13528), .B(n13630), .Z(n13521) );
  XNOR U13826 ( .A(n13527), .B(n13525), .Z(n13630) );
  AND U13827 ( .A(n13631), .B(n13632), .Z(n13525) );
  NANDN U13828 ( .A(n13633), .B(n13634), .Z(n13632) );
  OR U13829 ( .A(n13635), .B(n13636), .Z(n13634) );
  NAND U13830 ( .A(n13636), .B(n13635), .Z(n13631) );
  ANDN U13831 ( .B(B[200]), .A(n36), .Z(n13527) );
  XNOR U13832 ( .A(n13535), .B(n13637), .Z(n13528) );
  XNOR U13833 ( .A(n13534), .B(n13532), .Z(n13637) );
  AND U13834 ( .A(n13638), .B(n13639), .Z(n13532) );
  NANDN U13835 ( .A(n13640), .B(n13641), .Z(n13639) );
  NANDN U13836 ( .A(n13642), .B(n13643), .Z(n13641) );
  NANDN U13837 ( .A(n13643), .B(n13642), .Z(n13638) );
  ANDN U13838 ( .B(B[201]), .A(n37), .Z(n13534) );
  XNOR U13839 ( .A(n13542), .B(n13644), .Z(n13535) );
  XNOR U13840 ( .A(n13541), .B(n13539), .Z(n13644) );
  AND U13841 ( .A(n13645), .B(n13646), .Z(n13539) );
  NANDN U13842 ( .A(n13647), .B(n13648), .Z(n13646) );
  OR U13843 ( .A(n13649), .B(n13650), .Z(n13648) );
  NAND U13844 ( .A(n13650), .B(n13649), .Z(n13645) );
  ANDN U13845 ( .B(B[202]), .A(n38), .Z(n13541) );
  XNOR U13846 ( .A(n13549), .B(n13651), .Z(n13542) );
  XNOR U13847 ( .A(n13548), .B(n13546), .Z(n13651) );
  AND U13848 ( .A(n13652), .B(n13653), .Z(n13546) );
  NANDN U13849 ( .A(n13654), .B(n13655), .Z(n13653) );
  NANDN U13850 ( .A(n13656), .B(n13657), .Z(n13655) );
  NANDN U13851 ( .A(n13657), .B(n13656), .Z(n13652) );
  ANDN U13852 ( .B(B[203]), .A(n39), .Z(n13548) );
  XNOR U13853 ( .A(n13556), .B(n13658), .Z(n13549) );
  XNOR U13854 ( .A(n13555), .B(n13553), .Z(n13658) );
  AND U13855 ( .A(n13659), .B(n13660), .Z(n13553) );
  NANDN U13856 ( .A(n13661), .B(n13662), .Z(n13660) );
  OR U13857 ( .A(n13663), .B(n13664), .Z(n13662) );
  NAND U13858 ( .A(n13664), .B(n13663), .Z(n13659) );
  ANDN U13859 ( .B(B[204]), .A(n40), .Z(n13555) );
  XNOR U13860 ( .A(n13563), .B(n13665), .Z(n13556) );
  XNOR U13861 ( .A(n13562), .B(n13560), .Z(n13665) );
  AND U13862 ( .A(n13666), .B(n13667), .Z(n13560) );
  NANDN U13863 ( .A(n13668), .B(n13669), .Z(n13667) );
  NAND U13864 ( .A(n13670), .B(n13671), .Z(n13669) );
  ANDN U13865 ( .B(B[205]), .A(n41), .Z(n13562) );
  XOR U13866 ( .A(n13569), .B(n13672), .Z(n13563) );
  XNOR U13867 ( .A(n13567), .B(n13570), .Z(n13672) );
  NAND U13868 ( .A(A[2]), .B(B[206]), .Z(n13570) );
  NANDN U13869 ( .A(n13673), .B(n13674), .Z(n13567) );
  AND U13870 ( .A(A[0]), .B(B[207]), .Z(n13674) );
  XNOR U13871 ( .A(n13572), .B(n13675), .Z(n13569) );
  NAND U13872 ( .A(A[0]), .B(B[208]), .Z(n13675) );
  NAND U13873 ( .A(B[207]), .B(A[1]), .Z(n13572) );
  NAND U13874 ( .A(n13676), .B(n13677), .Z(n329) );
  NANDN U13875 ( .A(n13678), .B(n13679), .Z(n13677) );
  OR U13876 ( .A(n13680), .B(n13681), .Z(n13679) );
  NAND U13877 ( .A(n13681), .B(n13680), .Z(n13676) );
  XOR U13878 ( .A(n331), .B(n330), .Z(\A1[205] ) );
  XOR U13879 ( .A(n13681), .B(n13682), .Z(n330) );
  XNOR U13880 ( .A(n13680), .B(n13678), .Z(n13682) );
  AND U13881 ( .A(n13683), .B(n13684), .Z(n13678) );
  NANDN U13882 ( .A(n13685), .B(n13686), .Z(n13684) );
  NANDN U13883 ( .A(n13687), .B(n13688), .Z(n13686) );
  NANDN U13884 ( .A(n13688), .B(n13687), .Z(n13683) );
  ANDN U13885 ( .B(B[192]), .A(n29), .Z(n13680) );
  XNOR U13886 ( .A(n13587), .B(n13689), .Z(n13681) );
  XNOR U13887 ( .A(n13586), .B(n13584), .Z(n13689) );
  AND U13888 ( .A(n13690), .B(n13691), .Z(n13584) );
  NANDN U13889 ( .A(n13692), .B(n13693), .Z(n13691) );
  OR U13890 ( .A(n13694), .B(n13695), .Z(n13693) );
  NAND U13891 ( .A(n13695), .B(n13694), .Z(n13690) );
  ANDN U13892 ( .B(B[193]), .A(n30), .Z(n13586) );
  XNOR U13893 ( .A(n13594), .B(n13696), .Z(n13587) );
  XNOR U13894 ( .A(n13593), .B(n13591), .Z(n13696) );
  AND U13895 ( .A(n13697), .B(n13698), .Z(n13591) );
  NANDN U13896 ( .A(n13699), .B(n13700), .Z(n13698) );
  NANDN U13897 ( .A(n13701), .B(n13702), .Z(n13700) );
  NANDN U13898 ( .A(n13702), .B(n13701), .Z(n13697) );
  ANDN U13899 ( .B(B[194]), .A(n31), .Z(n13593) );
  XNOR U13900 ( .A(n13601), .B(n13703), .Z(n13594) );
  XNOR U13901 ( .A(n13600), .B(n13598), .Z(n13703) );
  AND U13902 ( .A(n13704), .B(n13705), .Z(n13598) );
  NANDN U13903 ( .A(n13706), .B(n13707), .Z(n13705) );
  OR U13904 ( .A(n13708), .B(n13709), .Z(n13707) );
  NAND U13905 ( .A(n13709), .B(n13708), .Z(n13704) );
  ANDN U13906 ( .B(B[195]), .A(n32), .Z(n13600) );
  XNOR U13907 ( .A(n13608), .B(n13710), .Z(n13601) );
  XNOR U13908 ( .A(n13607), .B(n13605), .Z(n13710) );
  AND U13909 ( .A(n13711), .B(n13712), .Z(n13605) );
  NANDN U13910 ( .A(n13713), .B(n13714), .Z(n13712) );
  NANDN U13911 ( .A(n13715), .B(n13716), .Z(n13714) );
  NANDN U13912 ( .A(n13716), .B(n13715), .Z(n13711) );
  ANDN U13913 ( .B(B[196]), .A(n33), .Z(n13607) );
  XNOR U13914 ( .A(n13615), .B(n13717), .Z(n13608) );
  XNOR U13915 ( .A(n13614), .B(n13612), .Z(n13717) );
  AND U13916 ( .A(n13718), .B(n13719), .Z(n13612) );
  NANDN U13917 ( .A(n13720), .B(n13721), .Z(n13719) );
  OR U13918 ( .A(n13722), .B(n13723), .Z(n13721) );
  NAND U13919 ( .A(n13723), .B(n13722), .Z(n13718) );
  ANDN U13920 ( .B(B[197]), .A(n34), .Z(n13614) );
  XNOR U13921 ( .A(n13622), .B(n13724), .Z(n13615) );
  XNOR U13922 ( .A(n13621), .B(n13619), .Z(n13724) );
  AND U13923 ( .A(n13725), .B(n13726), .Z(n13619) );
  NANDN U13924 ( .A(n13727), .B(n13728), .Z(n13726) );
  NANDN U13925 ( .A(n13729), .B(n13730), .Z(n13728) );
  NANDN U13926 ( .A(n13730), .B(n13729), .Z(n13725) );
  ANDN U13927 ( .B(B[198]), .A(n35), .Z(n13621) );
  XNOR U13928 ( .A(n13629), .B(n13731), .Z(n13622) );
  XNOR U13929 ( .A(n13628), .B(n13626), .Z(n13731) );
  AND U13930 ( .A(n13732), .B(n13733), .Z(n13626) );
  NANDN U13931 ( .A(n13734), .B(n13735), .Z(n13733) );
  OR U13932 ( .A(n13736), .B(n13737), .Z(n13735) );
  NAND U13933 ( .A(n13737), .B(n13736), .Z(n13732) );
  ANDN U13934 ( .B(B[199]), .A(n36), .Z(n13628) );
  XNOR U13935 ( .A(n13636), .B(n13738), .Z(n13629) );
  XNOR U13936 ( .A(n13635), .B(n13633), .Z(n13738) );
  AND U13937 ( .A(n13739), .B(n13740), .Z(n13633) );
  NANDN U13938 ( .A(n13741), .B(n13742), .Z(n13740) );
  NANDN U13939 ( .A(n13743), .B(n13744), .Z(n13742) );
  NANDN U13940 ( .A(n13744), .B(n13743), .Z(n13739) );
  ANDN U13941 ( .B(B[200]), .A(n37), .Z(n13635) );
  XNOR U13942 ( .A(n13643), .B(n13745), .Z(n13636) );
  XNOR U13943 ( .A(n13642), .B(n13640), .Z(n13745) );
  AND U13944 ( .A(n13746), .B(n13747), .Z(n13640) );
  NANDN U13945 ( .A(n13748), .B(n13749), .Z(n13747) );
  OR U13946 ( .A(n13750), .B(n13751), .Z(n13749) );
  NAND U13947 ( .A(n13751), .B(n13750), .Z(n13746) );
  ANDN U13948 ( .B(B[201]), .A(n38), .Z(n13642) );
  XNOR U13949 ( .A(n13650), .B(n13752), .Z(n13643) );
  XNOR U13950 ( .A(n13649), .B(n13647), .Z(n13752) );
  AND U13951 ( .A(n13753), .B(n13754), .Z(n13647) );
  NANDN U13952 ( .A(n13755), .B(n13756), .Z(n13754) );
  NANDN U13953 ( .A(n13757), .B(n13758), .Z(n13756) );
  NANDN U13954 ( .A(n13758), .B(n13757), .Z(n13753) );
  ANDN U13955 ( .B(B[202]), .A(n39), .Z(n13649) );
  XNOR U13956 ( .A(n13657), .B(n13759), .Z(n13650) );
  XNOR U13957 ( .A(n13656), .B(n13654), .Z(n13759) );
  AND U13958 ( .A(n13760), .B(n13761), .Z(n13654) );
  NANDN U13959 ( .A(n13762), .B(n13763), .Z(n13761) );
  OR U13960 ( .A(n13764), .B(n13765), .Z(n13763) );
  NAND U13961 ( .A(n13765), .B(n13764), .Z(n13760) );
  ANDN U13962 ( .B(B[203]), .A(n40), .Z(n13656) );
  XNOR U13963 ( .A(n13664), .B(n13766), .Z(n13657) );
  XNOR U13964 ( .A(n13663), .B(n13661), .Z(n13766) );
  AND U13965 ( .A(n13767), .B(n13768), .Z(n13661) );
  NANDN U13966 ( .A(n13769), .B(n13770), .Z(n13768) );
  NAND U13967 ( .A(n13771), .B(n13772), .Z(n13770) );
  ANDN U13968 ( .B(B[204]), .A(n41), .Z(n13663) );
  XOR U13969 ( .A(n13670), .B(n13773), .Z(n13664) );
  XNOR U13970 ( .A(n13668), .B(n13671), .Z(n13773) );
  NAND U13971 ( .A(A[2]), .B(B[205]), .Z(n13671) );
  NANDN U13972 ( .A(n13774), .B(n13775), .Z(n13668) );
  AND U13973 ( .A(A[0]), .B(B[206]), .Z(n13775) );
  XNOR U13974 ( .A(n13673), .B(n13776), .Z(n13670) );
  NAND U13975 ( .A(A[0]), .B(B[207]), .Z(n13776) );
  NAND U13976 ( .A(B[206]), .B(A[1]), .Z(n13673) );
  NAND U13977 ( .A(n13777), .B(n13778), .Z(n331) );
  NANDN U13978 ( .A(n13779), .B(n13780), .Z(n13778) );
  OR U13979 ( .A(n13781), .B(n13782), .Z(n13780) );
  NAND U13980 ( .A(n13782), .B(n13781), .Z(n13777) );
  XOR U13981 ( .A(n333), .B(n332), .Z(\A1[204] ) );
  XOR U13982 ( .A(n13782), .B(n13783), .Z(n332) );
  XNOR U13983 ( .A(n13781), .B(n13779), .Z(n13783) );
  AND U13984 ( .A(n13784), .B(n13785), .Z(n13779) );
  NANDN U13985 ( .A(n13786), .B(n13787), .Z(n13785) );
  NANDN U13986 ( .A(n13788), .B(n13789), .Z(n13787) );
  NANDN U13987 ( .A(n13789), .B(n13788), .Z(n13784) );
  ANDN U13988 ( .B(B[191]), .A(n29), .Z(n13781) );
  XNOR U13989 ( .A(n13688), .B(n13790), .Z(n13782) );
  XNOR U13990 ( .A(n13687), .B(n13685), .Z(n13790) );
  AND U13991 ( .A(n13791), .B(n13792), .Z(n13685) );
  NANDN U13992 ( .A(n13793), .B(n13794), .Z(n13792) );
  OR U13993 ( .A(n13795), .B(n13796), .Z(n13794) );
  NAND U13994 ( .A(n13796), .B(n13795), .Z(n13791) );
  ANDN U13995 ( .B(B[192]), .A(n30), .Z(n13687) );
  XNOR U13996 ( .A(n13695), .B(n13797), .Z(n13688) );
  XNOR U13997 ( .A(n13694), .B(n13692), .Z(n13797) );
  AND U13998 ( .A(n13798), .B(n13799), .Z(n13692) );
  NANDN U13999 ( .A(n13800), .B(n13801), .Z(n13799) );
  NANDN U14000 ( .A(n13802), .B(n13803), .Z(n13801) );
  NANDN U14001 ( .A(n13803), .B(n13802), .Z(n13798) );
  ANDN U14002 ( .B(B[193]), .A(n31), .Z(n13694) );
  XNOR U14003 ( .A(n13702), .B(n13804), .Z(n13695) );
  XNOR U14004 ( .A(n13701), .B(n13699), .Z(n13804) );
  AND U14005 ( .A(n13805), .B(n13806), .Z(n13699) );
  NANDN U14006 ( .A(n13807), .B(n13808), .Z(n13806) );
  OR U14007 ( .A(n13809), .B(n13810), .Z(n13808) );
  NAND U14008 ( .A(n13810), .B(n13809), .Z(n13805) );
  ANDN U14009 ( .B(B[194]), .A(n32), .Z(n13701) );
  XNOR U14010 ( .A(n13709), .B(n13811), .Z(n13702) );
  XNOR U14011 ( .A(n13708), .B(n13706), .Z(n13811) );
  AND U14012 ( .A(n13812), .B(n13813), .Z(n13706) );
  NANDN U14013 ( .A(n13814), .B(n13815), .Z(n13813) );
  NANDN U14014 ( .A(n13816), .B(n13817), .Z(n13815) );
  NANDN U14015 ( .A(n13817), .B(n13816), .Z(n13812) );
  ANDN U14016 ( .B(B[195]), .A(n33), .Z(n13708) );
  XNOR U14017 ( .A(n13716), .B(n13818), .Z(n13709) );
  XNOR U14018 ( .A(n13715), .B(n13713), .Z(n13818) );
  AND U14019 ( .A(n13819), .B(n13820), .Z(n13713) );
  NANDN U14020 ( .A(n13821), .B(n13822), .Z(n13820) );
  OR U14021 ( .A(n13823), .B(n13824), .Z(n13822) );
  NAND U14022 ( .A(n13824), .B(n13823), .Z(n13819) );
  ANDN U14023 ( .B(B[196]), .A(n34), .Z(n13715) );
  XNOR U14024 ( .A(n13723), .B(n13825), .Z(n13716) );
  XNOR U14025 ( .A(n13722), .B(n13720), .Z(n13825) );
  AND U14026 ( .A(n13826), .B(n13827), .Z(n13720) );
  NANDN U14027 ( .A(n13828), .B(n13829), .Z(n13827) );
  NANDN U14028 ( .A(n13830), .B(n13831), .Z(n13829) );
  NANDN U14029 ( .A(n13831), .B(n13830), .Z(n13826) );
  ANDN U14030 ( .B(B[197]), .A(n35), .Z(n13722) );
  XNOR U14031 ( .A(n13730), .B(n13832), .Z(n13723) );
  XNOR U14032 ( .A(n13729), .B(n13727), .Z(n13832) );
  AND U14033 ( .A(n13833), .B(n13834), .Z(n13727) );
  NANDN U14034 ( .A(n13835), .B(n13836), .Z(n13834) );
  OR U14035 ( .A(n13837), .B(n13838), .Z(n13836) );
  NAND U14036 ( .A(n13838), .B(n13837), .Z(n13833) );
  ANDN U14037 ( .B(B[198]), .A(n36), .Z(n13729) );
  XNOR U14038 ( .A(n13737), .B(n13839), .Z(n13730) );
  XNOR U14039 ( .A(n13736), .B(n13734), .Z(n13839) );
  AND U14040 ( .A(n13840), .B(n13841), .Z(n13734) );
  NANDN U14041 ( .A(n13842), .B(n13843), .Z(n13841) );
  NANDN U14042 ( .A(n13844), .B(n13845), .Z(n13843) );
  NANDN U14043 ( .A(n13845), .B(n13844), .Z(n13840) );
  ANDN U14044 ( .B(B[199]), .A(n37), .Z(n13736) );
  XNOR U14045 ( .A(n13744), .B(n13846), .Z(n13737) );
  XNOR U14046 ( .A(n13743), .B(n13741), .Z(n13846) );
  AND U14047 ( .A(n13847), .B(n13848), .Z(n13741) );
  NANDN U14048 ( .A(n13849), .B(n13850), .Z(n13848) );
  OR U14049 ( .A(n13851), .B(n13852), .Z(n13850) );
  NAND U14050 ( .A(n13852), .B(n13851), .Z(n13847) );
  ANDN U14051 ( .B(B[200]), .A(n38), .Z(n13743) );
  XNOR U14052 ( .A(n13751), .B(n13853), .Z(n13744) );
  XNOR U14053 ( .A(n13750), .B(n13748), .Z(n13853) );
  AND U14054 ( .A(n13854), .B(n13855), .Z(n13748) );
  NANDN U14055 ( .A(n13856), .B(n13857), .Z(n13855) );
  NANDN U14056 ( .A(n13858), .B(n13859), .Z(n13857) );
  NANDN U14057 ( .A(n13859), .B(n13858), .Z(n13854) );
  ANDN U14058 ( .B(B[201]), .A(n39), .Z(n13750) );
  XNOR U14059 ( .A(n13758), .B(n13860), .Z(n13751) );
  XNOR U14060 ( .A(n13757), .B(n13755), .Z(n13860) );
  AND U14061 ( .A(n13861), .B(n13862), .Z(n13755) );
  NANDN U14062 ( .A(n13863), .B(n13864), .Z(n13862) );
  OR U14063 ( .A(n13865), .B(n13866), .Z(n13864) );
  NAND U14064 ( .A(n13866), .B(n13865), .Z(n13861) );
  ANDN U14065 ( .B(B[202]), .A(n40), .Z(n13757) );
  XNOR U14066 ( .A(n13765), .B(n13867), .Z(n13758) );
  XNOR U14067 ( .A(n13764), .B(n13762), .Z(n13867) );
  AND U14068 ( .A(n13868), .B(n13869), .Z(n13762) );
  NANDN U14069 ( .A(n13870), .B(n13871), .Z(n13869) );
  NAND U14070 ( .A(n13872), .B(n13873), .Z(n13871) );
  ANDN U14071 ( .B(B[203]), .A(n41), .Z(n13764) );
  XOR U14072 ( .A(n13771), .B(n13874), .Z(n13765) );
  XNOR U14073 ( .A(n13769), .B(n13772), .Z(n13874) );
  NAND U14074 ( .A(A[2]), .B(B[204]), .Z(n13772) );
  NANDN U14075 ( .A(n13875), .B(n13876), .Z(n13769) );
  AND U14076 ( .A(A[0]), .B(B[205]), .Z(n13876) );
  XNOR U14077 ( .A(n13774), .B(n13877), .Z(n13771) );
  NAND U14078 ( .A(A[0]), .B(B[206]), .Z(n13877) );
  NAND U14079 ( .A(B[205]), .B(A[1]), .Z(n13774) );
  NAND U14080 ( .A(n13878), .B(n13879), .Z(n333) );
  NANDN U14081 ( .A(n13880), .B(n13881), .Z(n13879) );
  OR U14082 ( .A(n13882), .B(n13883), .Z(n13881) );
  NAND U14083 ( .A(n13883), .B(n13882), .Z(n13878) );
  XOR U14084 ( .A(n335), .B(n334), .Z(\A1[203] ) );
  XOR U14085 ( .A(n13883), .B(n13884), .Z(n334) );
  XNOR U14086 ( .A(n13882), .B(n13880), .Z(n13884) );
  AND U14087 ( .A(n13885), .B(n13886), .Z(n13880) );
  NANDN U14088 ( .A(n13887), .B(n13888), .Z(n13886) );
  NANDN U14089 ( .A(n13889), .B(n13890), .Z(n13888) );
  NANDN U14090 ( .A(n13890), .B(n13889), .Z(n13885) );
  ANDN U14091 ( .B(B[190]), .A(n29), .Z(n13882) );
  XNOR U14092 ( .A(n13789), .B(n13891), .Z(n13883) );
  XNOR U14093 ( .A(n13788), .B(n13786), .Z(n13891) );
  AND U14094 ( .A(n13892), .B(n13893), .Z(n13786) );
  NANDN U14095 ( .A(n13894), .B(n13895), .Z(n13893) );
  OR U14096 ( .A(n13896), .B(n13897), .Z(n13895) );
  NAND U14097 ( .A(n13897), .B(n13896), .Z(n13892) );
  ANDN U14098 ( .B(B[191]), .A(n30), .Z(n13788) );
  XNOR U14099 ( .A(n13796), .B(n13898), .Z(n13789) );
  XNOR U14100 ( .A(n13795), .B(n13793), .Z(n13898) );
  AND U14101 ( .A(n13899), .B(n13900), .Z(n13793) );
  NANDN U14102 ( .A(n13901), .B(n13902), .Z(n13900) );
  NANDN U14103 ( .A(n13903), .B(n13904), .Z(n13902) );
  NANDN U14104 ( .A(n13904), .B(n13903), .Z(n13899) );
  ANDN U14105 ( .B(B[192]), .A(n31), .Z(n13795) );
  XNOR U14106 ( .A(n13803), .B(n13905), .Z(n13796) );
  XNOR U14107 ( .A(n13802), .B(n13800), .Z(n13905) );
  AND U14108 ( .A(n13906), .B(n13907), .Z(n13800) );
  NANDN U14109 ( .A(n13908), .B(n13909), .Z(n13907) );
  OR U14110 ( .A(n13910), .B(n13911), .Z(n13909) );
  NAND U14111 ( .A(n13911), .B(n13910), .Z(n13906) );
  ANDN U14112 ( .B(B[193]), .A(n32), .Z(n13802) );
  XNOR U14113 ( .A(n13810), .B(n13912), .Z(n13803) );
  XNOR U14114 ( .A(n13809), .B(n13807), .Z(n13912) );
  AND U14115 ( .A(n13913), .B(n13914), .Z(n13807) );
  NANDN U14116 ( .A(n13915), .B(n13916), .Z(n13914) );
  NANDN U14117 ( .A(n13917), .B(n13918), .Z(n13916) );
  NANDN U14118 ( .A(n13918), .B(n13917), .Z(n13913) );
  ANDN U14119 ( .B(B[194]), .A(n33), .Z(n13809) );
  XNOR U14120 ( .A(n13817), .B(n13919), .Z(n13810) );
  XNOR U14121 ( .A(n13816), .B(n13814), .Z(n13919) );
  AND U14122 ( .A(n13920), .B(n13921), .Z(n13814) );
  NANDN U14123 ( .A(n13922), .B(n13923), .Z(n13921) );
  OR U14124 ( .A(n13924), .B(n13925), .Z(n13923) );
  NAND U14125 ( .A(n13925), .B(n13924), .Z(n13920) );
  ANDN U14126 ( .B(B[195]), .A(n34), .Z(n13816) );
  XNOR U14127 ( .A(n13824), .B(n13926), .Z(n13817) );
  XNOR U14128 ( .A(n13823), .B(n13821), .Z(n13926) );
  AND U14129 ( .A(n13927), .B(n13928), .Z(n13821) );
  NANDN U14130 ( .A(n13929), .B(n13930), .Z(n13928) );
  NANDN U14131 ( .A(n13931), .B(n13932), .Z(n13930) );
  NANDN U14132 ( .A(n13932), .B(n13931), .Z(n13927) );
  ANDN U14133 ( .B(B[196]), .A(n35), .Z(n13823) );
  XNOR U14134 ( .A(n13831), .B(n13933), .Z(n13824) );
  XNOR U14135 ( .A(n13830), .B(n13828), .Z(n13933) );
  AND U14136 ( .A(n13934), .B(n13935), .Z(n13828) );
  NANDN U14137 ( .A(n13936), .B(n13937), .Z(n13935) );
  OR U14138 ( .A(n13938), .B(n13939), .Z(n13937) );
  NAND U14139 ( .A(n13939), .B(n13938), .Z(n13934) );
  ANDN U14140 ( .B(B[197]), .A(n36), .Z(n13830) );
  XNOR U14141 ( .A(n13838), .B(n13940), .Z(n13831) );
  XNOR U14142 ( .A(n13837), .B(n13835), .Z(n13940) );
  AND U14143 ( .A(n13941), .B(n13942), .Z(n13835) );
  NANDN U14144 ( .A(n13943), .B(n13944), .Z(n13942) );
  NANDN U14145 ( .A(n13945), .B(n13946), .Z(n13944) );
  NANDN U14146 ( .A(n13946), .B(n13945), .Z(n13941) );
  ANDN U14147 ( .B(B[198]), .A(n37), .Z(n13837) );
  XNOR U14148 ( .A(n13845), .B(n13947), .Z(n13838) );
  XNOR U14149 ( .A(n13844), .B(n13842), .Z(n13947) );
  AND U14150 ( .A(n13948), .B(n13949), .Z(n13842) );
  NANDN U14151 ( .A(n13950), .B(n13951), .Z(n13949) );
  OR U14152 ( .A(n13952), .B(n13953), .Z(n13951) );
  NAND U14153 ( .A(n13953), .B(n13952), .Z(n13948) );
  ANDN U14154 ( .B(B[199]), .A(n38), .Z(n13844) );
  XNOR U14155 ( .A(n13852), .B(n13954), .Z(n13845) );
  XNOR U14156 ( .A(n13851), .B(n13849), .Z(n13954) );
  AND U14157 ( .A(n13955), .B(n13956), .Z(n13849) );
  NANDN U14158 ( .A(n13957), .B(n13958), .Z(n13956) );
  NANDN U14159 ( .A(n13959), .B(n13960), .Z(n13958) );
  NANDN U14160 ( .A(n13960), .B(n13959), .Z(n13955) );
  ANDN U14161 ( .B(B[200]), .A(n39), .Z(n13851) );
  XNOR U14162 ( .A(n13859), .B(n13961), .Z(n13852) );
  XNOR U14163 ( .A(n13858), .B(n13856), .Z(n13961) );
  AND U14164 ( .A(n13962), .B(n13963), .Z(n13856) );
  NANDN U14165 ( .A(n13964), .B(n13965), .Z(n13963) );
  OR U14166 ( .A(n13966), .B(n13967), .Z(n13965) );
  NAND U14167 ( .A(n13967), .B(n13966), .Z(n13962) );
  ANDN U14168 ( .B(B[201]), .A(n40), .Z(n13858) );
  XNOR U14169 ( .A(n13866), .B(n13968), .Z(n13859) );
  XNOR U14170 ( .A(n13865), .B(n13863), .Z(n13968) );
  AND U14171 ( .A(n13969), .B(n13970), .Z(n13863) );
  NANDN U14172 ( .A(n13971), .B(n13972), .Z(n13970) );
  NAND U14173 ( .A(n13973), .B(n13974), .Z(n13972) );
  ANDN U14174 ( .B(B[202]), .A(n41), .Z(n13865) );
  XOR U14175 ( .A(n13872), .B(n13975), .Z(n13866) );
  XNOR U14176 ( .A(n13870), .B(n13873), .Z(n13975) );
  NAND U14177 ( .A(A[2]), .B(B[203]), .Z(n13873) );
  NANDN U14178 ( .A(n13976), .B(n13977), .Z(n13870) );
  AND U14179 ( .A(A[0]), .B(B[204]), .Z(n13977) );
  XNOR U14180 ( .A(n13875), .B(n13978), .Z(n13872) );
  NAND U14181 ( .A(A[0]), .B(B[205]), .Z(n13978) );
  NAND U14182 ( .A(B[204]), .B(A[1]), .Z(n13875) );
  NAND U14183 ( .A(n13979), .B(n13980), .Z(n335) );
  NANDN U14184 ( .A(n13981), .B(n13982), .Z(n13980) );
  OR U14185 ( .A(n13983), .B(n13984), .Z(n13982) );
  NAND U14186 ( .A(n13984), .B(n13983), .Z(n13979) );
  XOR U14187 ( .A(n337), .B(n336), .Z(\A1[202] ) );
  XOR U14188 ( .A(n13984), .B(n13985), .Z(n336) );
  XNOR U14189 ( .A(n13983), .B(n13981), .Z(n13985) );
  AND U14190 ( .A(n13986), .B(n13987), .Z(n13981) );
  NANDN U14191 ( .A(n13988), .B(n13989), .Z(n13987) );
  NANDN U14192 ( .A(n13990), .B(n13991), .Z(n13989) );
  NANDN U14193 ( .A(n13991), .B(n13990), .Z(n13986) );
  ANDN U14194 ( .B(B[189]), .A(n29), .Z(n13983) );
  XNOR U14195 ( .A(n13890), .B(n13992), .Z(n13984) );
  XNOR U14196 ( .A(n13889), .B(n13887), .Z(n13992) );
  AND U14197 ( .A(n13993), .B(n13994), .Z(n13887) );
  NANDN U14198 ( .A(n13995), .B(n13996), .Z(n13994) );
  OR U14199 ( .A(n13997), .B(n13998), .Z(n13996) );
  NAND U14200 ( .A(n13998), .B(n13997), .Z(n13993) );
  ANDN U14201 ( .B(B[190]), .A(n30), .Z(n13889) );
  XNOR U14202 ( .A(n13897), .B(n13999), .Z(n13890) );
  XNOR U14203 ( .A(n13896), .B(n13894), .Z(n13999) );
  AND U14204 ( .A(n14000), .B(n14001), .Z(n13894) );
  NANDN U14205 ( .A(n14002), .B(n14003), .Z(n14001) );
  NANDN U14206 ( .A(n14004), .B(n14005), .Z(n14003) );
  NANDN U14207 ( .A(n14005), .B(n14004), .Z(n14000) );
  ANDN U14208 ( .B(B[191]), .A(n31), .Z(n13896) );
  XNOR U14209 ( .A(n13904), .B(n14006), .Z(n13897) );
  XNOR U14210 ( .A(n13903), .B(n13901), .Z(n14006) );
  AND U14211 ( .A(n14007), .B(n14008), .Z(n13901) );
  NANDN U14212 ( .A(n14009), .B(n14010), .Z(n14008) );
  OR U14213 ( .A(n14011), .B(n14012), .Z(n14010) );
  NAND U14214 ( .A(n14012), .B(n14011), .Z(n14007) );
  ANDN U14215 ( .B(B[192]), .A(n32), .Z(n13903) );
  XNOR U14216 ( .A(n13911), .B(n14013), .Z(n13904) );
  XNOR U14217 ( .A(n13910), .B(n13908), .Z(n14013) );
  AND U14218 ( .A(n14014), .B(n14015), .Z(n13908) );
  NANDN U14219 ( .A(n14016), .B(n14017), .Z(n14015) );
  NANDN U14220 ( .A(n14018), .B(n14019), .Z(n14017) );
  NANDN U14221 ( .A(n14019), .B(n14018), .Z(n14014) );
  ANDN U14222 ( .B(B[193]), .A(n33), .Z(n13910) );
  XNOR U14223 ( .A(n13918), .B(n14020), .Z(n13911) );
  XNOR U14224 ( .A(n13917), .B(n13915), .Z(n14020) );
  AND U14225 ( .A(n14021), .B(n14022), .Z(n13915) );
  NANDN U14226 ( .A(n14023), .B(n14024), .Z(n14022) );
  OR U14227 ( .A(n14025), .B(n14026), .Z(n14024) );
  NAND U14228 ( .A(n14026), .B(n14025), .Z(n14021) );
  ANDN U14229 ( .B(B[194]), .A(n34), .Z(n13917) );
  XNOR U14230 ( .A(n13925), .B(n14027), .Z(n13918) );
  XNOR U14231 ( .A(n13924), .B(n13922), .Z(n14027) );
  AND U14232 ( .A(n14028), .B(n14029), .Z(n13922) );
  NANDN U14233 ( .A(n14030), .B(n14031), .Z(n14029) );
  NANDN U14234 ( .A(n14032), .B(n14033), .Z(n14031) );
  NANDN U14235 ( .A(n14033), .B(n14032), .Z(n14028) );
  ANDN U14236 ( .B(B[195]), .A(n35), .Z(n13924) );
  XNOR U14237 ( .A(n13932), .B(n14034), .Z(n13925) );
  XNOR U14238 ( .A(n13931), .B(n13929), .Z(n14034) );
  AND U14239 ( .A(n14035), .B(n14036), .Z(n13929) );
  NANDN U14240 ( .A(n14037), .B(n14038), .Z(n14036) );
  OR U14241 ( .A(n14039), .B(n14040), .Z(n14038) );
  NAND U14242 ( .A(n14040), .B(n14039), .Z(n14035) );
  ANDN U14243 ( .B(B[196]), .A(n36), .Z(n13931) );
  XNOR U14244 ( .A(n13939), .B(n14041), .Z(n13932) );
  XNOR U14245 ( .A(n13938), .B(n13936), .Z(n14041) );
  AND U14246 ( .A(n14042), .B(n14043), .Z(n13936) );
  NANDN U14247 ( .A(n14044), .B(n14045), .Z(n14043) );
  NANDN U14248 ( .A(n14046), .B(n14047), .Z(n14045) );
  NANDN U14249 ( .A(n14047), .B(n14046), .Z(n14042) );
  ANDN U14250 ( .B(B[197]), .A(n37), .Z(n13938) );
  XNOR U14251 ( .A(n13946), .B(n14048), .Z(n13939) );
  XNOR U14252 ( .A(n13945), .B(n13943), .Z(n14048) );
  AND U14253 ( .A(n14049), .B(n14050), .Z(n13943) );
  NANDN U14254 ( .A(n14051), .B(n14052), .Z(n14050) );
  OR U14255 ( .A(n14053), .B(n14054), .Z(n14052) );
  NAND U14256 ( .A(n14054), .B(n14053), .Z(n14049) );
  ANDN U14257 ( .B(B[198]), .A(n38), .Z(n13945) );
  XNOR U14258 ( .A(n13953), .B(n14055), .Z(n13946) );
  XNOR U14259 ( .A(n13952), .B(n13950), .Z(n14055) );
  AND U14260 ( .A(n14056), .B(n14057), .Z(n13950) );
  NANDN U14261 ( .A(n14058), .B(n14059), .Z(n14057) );
  NANDN U14262 ( .A(n14060), .B(n14061), .Z(n14059) );
  NANDN U14263 ( .A(n14061), .B(n14060), .Z(n14056) );
  ANDN U14264 ( .B(B[199]), .A(n39), .Z(n13952) );
  XNOR U14265 ( .A(n13960), .B(n14062), .Z(n13953) );
  XNOR U14266 ( .A(n13959), .B(n13957), .Z(n14062) );
  AND U14267 ( .A(n14063), .B(n14064), .Z(n13957) );
  NANDN U14268 ( .A(n14065), .B(n14066), .Z(n14064) );
  OR U14269 ( .A(n14067), .B(n14068), .Z(n14066) );
  NAND U14270 ( .A(n14068), .B(n14067), .Z(n14063) );
  ANDN U14271 ( .B(B[200]), .A(n40), .Z(n13959) );
  XNOR U14272 ( .A(n13967), .B(n14069), .Z(n13960) );
  XNOR U14273 ( .A(n13966), .B(n13964), .Z(n14069) );
  AND U14274 ( .A(n14070), .B(n14071), .Z(n13964) );
  NANDN U14275 ( .A(n14072), .B(n14073), .Z(n14071) );
  NAND U14276 ( .A(n14074), .B(n14075), .Z(n14073) );
  ANDN U14277 ( .B(B[201]), .A(n41), .Z(n13966) );
  XOR U14278 ( .A(n13973), .B(n14076), .Z(n13967) );
  XNOR U14279 ( .A(n13971), .B(n13974), .Z(n14076) );
  NAND U14280 ( .A(A[2]), .B(B[202]), .Z(n13974) );
  NANDN U14281 ( .A(n14077), .B(n14078), .Z(n13971) );
  AND U14282 ( .A(A[0]), .B(B[203]), .Z(n14078) );
  XNOR U14283 ( .A(n13976), .B(n14079), .Z(n13973) );
  NAND U14284 ( .A(A[0]), .B(B[204]), .Z(n14079) );
  NAND U14285 ( .A(B[203]), .B(A[1]), .Z(n13976) );
  NAND U14286 ( .A(n14080), .B(n14081), .Z(n337) );
  NANDN U14287 ( .A(n14082), .B(n14083), .Z(n14081) );
  OR U14288 ( .A(n14084), .B(n14085), .Z(n14083) );
  NAND U14289 ( .A(n14085), .B(n14084), .Z(n14080) );
  XOR U14290 ( .A(n339), .B(n338), .Z(\A1[201] ) );
  XOR U14291 ( .A(n14085), .B(n14086), .Z(n338) );
  XNOR U14292 ( .A(n14084), .B(n14082), .Z(n14086) );
  AND U14293 ( .A(n14087), .B(n14088), .Z(n14082) );
  NANDN U14294 ( .A(n14089), .B(n14090), .Z(n14088) );
  NANDN U14295 ( .A(n14091), .B(n14092), .Z(n14090) );
  NANDN U14296 ( .A(n14092), .B(n14091), .Z(n14087) );
  ANDN U14297 ( .B(B[188]), .A(n29), .Z(n14084) );
  XNOR U14298 ( .A(n13991), .B(n14093), .Z(n14085) );
  XNOR U14299 ( .A(n13990), .B(n13988), .Z(n14093) );
  AND U14300 ( .A(n14094), .B(n14095), .Z(n13988) );
  NANDN U14301 ( .A(n14096), .B(n14097), .Z(n14095) );
  OR U14302 ( .A(n14098), .B(n14099), .Z(n14097) );
  NAND U14303 ( .A(n14099), .B(n14098), .Z(n14094) );
  ANDN U14304 ( .B(B[189]), .A(n30), .Z(n13990) );
  XNOR U14305 ( .A(n13998), .B(n14100), .Z(n13991) );
  XNOR U14306 ( .A(n13997), .B(n13995), .Z(n14100) );
  AND U14307 ( .A(n14101), .B(n14102), .Z(n13995) );
  NANDN U14308 ( .A(n14103), .B(n14104), .Z(n14102) );
  NANDN U14309 ( .A(n14105), .B(n14106), .Z(n14104) );
  NANDN U14310 ( .A(n14106), .B(n14105), .Z(n14101) );
  ANDN U14311 ( .B(B[190]), .A(n31), .Z(n13997) );
  XNOR U14312 ( .A(n14005), .B(n14107), .Z(n13998) );
  XNOR U14313 ( .A(n14004), .B(n14002), .Z(n14107) );
  AND U14314 ( .A(n14108), .B(n14109), .Z(n14002) );
  NANDN U14315 ( .A(n14110), .B(n14111), .Z(n14109) );
  OR U14316 ( .A(n14112), .B(n14113), .Z(n14111) );
  NAND U14317 ( .A(n14113), .B(n14112), .Z(n14108) );
  ANDN U14318 ( .B(B[191]), .A(n32), .Z(n14004) );
  XNOR U14319 ( .A(n14012), .B(n14114), .Z(n14005) );
  XNOR U14320 ( .A(n14011), .B(n14009), .Z(n14114) );
  AND U14321 ( .A(n14115), .B(n14116), .Z(n14009) );
  NANDN U14322 ( .A(n14117), .B(n14118), .Z(n14116) );
  NANDN U14323 ( .A(n14119), .B(n14120), .Z(n14118) );
  NANDN U14324 ( .A(n14120), .B(n14119), .Z(n14115) );
  ANDN U14325 ( .B(B[192]), .A(n33), .Z(n14011) );
  XNOR U14326 ( .A(n14019), .B(n14121), .Z(n14012) );
  XNOR U14327 ( .A(n14018), .B(n14016), .Z(n14121) );
  AND U14328 ( .A(n14122), .B(n14123), .Z(n14016) );
  NANDN U14329 ( .A(n14124), .B(n14125), .Z(n14123) );
  OR U14330 ( .A(n14126), .B(n14127), .Z(n14125) );
  NAND U14331 ( .A(n14127), .B(n14126), .Z(n14122) );
  ANDN U14332 ( .B(B[193]), .A(n34), .Z(n14018) );
  XNOR U14333 ( .A(n14026), .B(n14128), .Z(n14019) );
  XNOR U14334 ( .A(n14025), .B(n14023), .Z(n14128) );
  AND U14335 ( .A(n14129), .B(n14130), .Z(n14023) );
  NANDN U14336 ( .A(n14131), .B(n14132), .Z(n14130) );
  NANDN U14337 ( .A(n14133), .B(n14134), .Z(n14132) );
  NANDN U14338 ( .A(n14134), .B(n14133), .Z(n14129) );
  ANDN U14339 ( .B(B[194]), .A(n35), .Z(n14025) );
  XNOR U14340 ( .A(n14033), .B(n14135), .Z(n14026) );
  XNOR U14341 ( .A(n14032), .B(n14030), .Z(n14135) );
  AND U14342 ( .A(n14136), .B(n14137), .Z(n14030) );
  NANDN U14343 ( .A(n14138), .B(n14139), .Z(n14137) );
  OR U14344 ( .A(n14140), .B(n14141), .Z(n14139) );
  NAND U14345 ( .A(n14141), .B(n14140), .Z(n14136) );
  ANDN U14346 ( .B(B[195]), .A(n36), .Z(n14032) );
  XNOR U14347 ( .A(n14040), .B(n14142), .Z(n14033) );
  XNOR U14348 ( .A(n14039), .B(n14037), .Z(n14142) );
  AND U14349 ( .A(n14143), .B(n14144), .Z(n14037) );
  NANDN U14350 ( .A(n14145), .B(n14146), .Z(n14144) );
  NANDN U14351 ( .A(n14147), .B(n14148), .Z(n14146) );
  NANDN U14352 ( .A(n14148), .B(n14147), .Z(n14143) );
  ANDN U14353 ( .B(B[196]), .A(n37), .Z(n14039) );
  XNOR U14354 ( .A(n14047), .B(n14149), .Z(n14040) );
  XNOR U14355 ( .A(n14046), .B(n14044), .Z(n14149) );
  AND U14356 ( .A(n14150), .B(n14151), .Z(n14044) );
  NANDN U14357 ( .A(n14152), .B(n14153), .Z(n14151) );
  OR U14358 ( .A(n14154), .B(n14155), .Z(n14153) );
  NAND U14359 ( .A(n14155), .B(n14154), .Z(n14150) );
  ANDN U14360 ( .B(B[197]), .A(n38), .Z(n14046) );
  XNOR U14361 ( .A(n14054), .B(n14156), .Z(n14047) );
  XNOR U14362 ( .A(n14053), .B(n14051), .Z(n14156) );
  AND U14363 ( .A(n14157), .B(n14158), .Z(n14051) );
  NANDN U14364 ( .A(n14159), .B(n14160), .Z(n14158) );
  NANDN U14365 ( .A(n14161), .B(n14162), .Z(n14160) );
  NANDN U14366 ( .A(n14162), .B(n14161), .Z(n14157) );
  ANDN U14367 ( .B(B[198]), .A(n39), .Z(n14053) );
  XNOR U14368 ( .A(n14061), .B(n14163), .Z(n14054) );
  XNOR U14369 ( .A(n14060), .B(n14058), .Z(n14163) );
  AND U14370 ( .A(n14164), .B(n14165), .Z(n14058) );
  NANDN U14371 ( .A(n14166), .B(n14167), .Z(n14165) );
  OR U14372 ( .A(n14168), .B(n14169), .Z(n14167) );
  NAND U14373 ( .A(n14169), .B(n14168), .Z(n14164) );
  ANDN U14374 ( .B(B[199]), .A(n40), .Z(n14060) );
  XNOR U14375 ( .A(n14068), .B(n14170), .Z(n14061) );
  XNOR U14376 ( .A(n14067), .B(n14065), .Z(n14170) );
  AND U14377 ( .A(n14171), .B(n14172), .Z(n14065) );
  NANDN U14378 ( .A(n14173), .B(n14174), .Z(n14172) );
  NAND U14379 ( .A(n14175), .B(n14176), .Z(n14174) );
  ANDN U14380 ( .B(B[200]), .A(n41), .Z(n14067) );
  XOR U14381 ( .A(n14074), .B(n14177), .Z(n14068) );
  XNOR U14382 ( .A(n14072), .B(n14075), .Z(n14177) );
  NAND U14383 ( .A(A[2]), .B(B[201]), .Z(n14075) );
  NANDN U14384 ( .A(n14178), .B(n14179), .Z(n14072) );
  AND U14385 ( .A(A[0]), .B(B[202]), .Z(n14179) );
  XNOR U14386 ( .A(n14077), .B(n14180), .Z(n14074) );
  NAND U14387 ( .A(A[0]), .B(B[203]), .Z(n14180) );
  NAND U14388 ( .A(B[202]), .B(A[1]), .Z(n14077) );
  NAND U14389 ( .A(n14181), .B(n14182), .Z(n339) );
  NANDN U14390 ( .A(n14183), .B(n14184), .Z(n14182) );
  OR U14391 ( .A(n14185), .B(n14186), .Z(n14184) );
  NAND U14392 ( .A(n14186), .B(n14185), .Z(n14181) );
  XOR U14393 ( .A(n341), .B(n340), .Z(\A1[200] ) );
  XOR U14394 ( .A(n14186), .B(n14187), .Z(n340) );
  XNOR U14395 ( .A(n14185), .B(n14183), .Z(n14187) );
  AND U14396 ( .A(n14188), .B(n14189), .Z(n14183) );
  NANDN U14397 ( .A(n14190), .B(n14191), .Z(n14189) );
  NANDN U14398 ( .A(n14192), .B(n14193), .Z(n14191) );
  NANDN U14399 ( .A(n14193), .B(n14192), .Z(n14188) );
  ANDN U14400 ( .B(B[187]), .A(n29), .Z(n14185) );
  XNOR U14401 ( .A(n14092), .B(n14194), .Z(n14186) );
  XNOR U14402 ( .A(n14091), .B(n14089), .Z(n14194) );
  AND U14403 ( .A(n14195), .B(n14196), .Z(n14089) );
  NANDN U14404 ( .A(n14197), .B(n14198), .Z(n14196) );
  OR U14405 ( .A(n14199), .B(n14200), .Z(n14198) );
  NAND U14406 ( .A(n14200), .B(n14199), .Z(n14195) );
  ANDN U14407 ( .B(B[188]), .A(n30), .Z(n14091) );
  XNOR U14408 ( .A(n14099), .B(n14201), .Z(n14092) );
  XNOR U14409 ( .A(n14098), .B(n14096), .Z(n14201) );
  AND U14410 ( .A(n14202), .B(n14203), .Z(n14096) );
  NANDN U14411 ( .A(n14204), .B(n14205), .Z(n14203) );
  NANDN U14412 ( .A(n14206), .B(n14207), .Z(n14205) );
  NANDN U14413 ( .A(n14207), .B(n14206), .Z(n14202) );
  ANDN U14414 ( .B(B[189]), .A(n31), .Z(n14098) );
  XNOR U14415 ( .A(n14106), .B(n14208), .Z(n14099) );
  XNOR U14416 ( .A(n14105), .B(n14103), .Z(n14208) );
  AND U14417 ( .A(n14209), .B(n14210), .Z(n14103) );
  NANDN U14418 ( .A(n14211), .B(n14212), .Z(n14210) );
  OR U14419 ( .A(n14213), .B(n14214), .Z(n14212) );
  NAND U14420 ( .A(n14214), .B(n14213), .Z(n14209) );
  ANDN U14421 ( .B(B[190]), .A(n32), .Z(n14105) );
  XNOR U14422 ( .A(n14113), .B(n14215), .Z(n14106) );
  XNOR U14423 ( .A(n14112), .B(n14110), .Z(n14215) );
  AND U14424 ( .A(n14216), .B(n14217), .Z(n14110) );
  NANDN U14425 ( .A(n14218), .B(n14219), .Z(n14217) );
  NANDN U14426 ( .A(n14220), .B(n14221), .Z(n14219) );
  NANDN U14427 ( .A(n14221), .B(n14220), .Z(n14216) );
  ANDN U14428 ( .B(B[191]), .A(n33), .Z(n14112) );
  XNOR U14429 ( .A(n14120), .B(n14222), .Z(n14113) );
  XNOR U14430 ( .A(n14119), .B(n14117), .Z(n14222) );
  AND U14431 ( .A(n14223), .B(n14224), .Z(n14117) );
  NANDN U14432 ( .A(n14225), .B(n14226), .Z(n14224) );
  OR U14433 ( .A(n14227), .B(n14228), .Z(n14226) );
  NAND U14434 ( .A(n14228), .B(n14227), .Z(n14223) );
  ANDN U14435 ( .B(B[192]), .A(n34), .Z(n14119) );
  XNOR U14436 ( .A(n14127), .B(n14229), .Z(n14120) );
  XNOR U14437 ( .A(n14126), .B(n14124), .Z(n14229) );
  AND U14438 ( .A(n14230), .B(n14231), .Z(n14124) );
  NANDN U14439 ( .A(n14232), .B(n14233), .Z(n14231) );
  NANDN U14440 ( .A(n14234), .B(n14235), .Z(n14233) );
  NANDN U14441 ( .A(n14235), .B(n14234), .Z(n14230) );
  ANDN U14442 ( .B(B[193]), .A(n35), .Z(n14126) );
  XNOR U14443 ( .A(n14134), .B(n14236), .Z(n14127) );
  XNOR U14444 ( .A(n14133), .B(n14131), .Z(n14236) );
  AND U14445 ( .A(n14237), .B(n14238), .Z(n14131) );
  NANDN U14446 ( .A(n14239), .B(n14240), .Z(n14238) );
  OR U14447 ( .A(n14241), .B(n14242), .Z(n14240) );
  NAND U14448 ( .A(n14242), .B(n14241), .Z(n14237) );
  ANDN U14449 ( .B(B[194]), .A(n36), .Z(n14133) );
  XNOR U14450 ( .A(n14141), .B(n14243), .Z(n14134) );
  XNOR U14451 ( .A(n14140), .B(n14138), .Z(n14243) );
  AND U14452 ( .A(n14244), .B(n14245), .Z(n14138) );
  NANDN U14453 ( .A(n14246), .B(n14247), .Z(n14245) );
  NANDN U14454 ( .A(n14248), .B(n14249), .Z(n14247) );
  NANDN U14455 ( .A(n14249), .B(n14248), .Z(n14244) );
  ANDN U14456 ( .B(B[195]), .A(n37), .Z(n14140) );
  XNOR U14457 ( .A(n14148), .B(n14250), .Z(n14141) );
  XNOR U14458 ( .A(n14147), .B(n14145), .Z(n14250) );
  AND U14459 ( .A(n14251), .B(n14252), .Z(n14145) );
  NANDN U14460 ( .A(n14253), .B(n14254), .Z(n14252) );
  OR U14461 ( .A(n14255), .B(n14256), .Z(n14254) );
  NAND U14462 ( .A(n14256), .B(n14255), .Z(n14251) );
  ANDN U14463 ( .B(B[196]), .A(n38), .Z(n14147) );
  XNOR U14464 ( .A(n14155), .B(n14257), .Z(n14148) );
  XNOR U14465 ( .A(n14154), .B(n14152), .Z(n14257) );
  AND U14466 ( .A(n14258), .B(n14259), .Z(n14152) );
  NANDN U14467 ( .A(n14260), .B(n14261), .Z(n14259) );
  NANDN U14468 ( .A(n14262), .B(n14263), .Z(n14261) );
  NANDN U14469 ( .A(n14263), .B(n14262), .Z(n14258) );
  ANDN U14470 ( .B(B[197]), .A(n39), .Z(n14154) );
  XNOR U14471 ( .A(n14162), .B(n14264), .Z(n14155) );
  XNOR U14472 ( .A(n14161), .B(n14159), .Z(n14264) );
  AND U14473 ( .A(n14265), .B(n14266), .Z(n14159) );
  NANDN U14474 ( .A(n14267), .B(n14268), .Z(n14266) );
  OR U14475 ( .A(n14269), .B(n14270), .Z(n14268) );
  NAND U14476 ( .A(n14270), .B(n14269), .Z(n14265) );
  ANDN U14477 ( .B(B[198]), .A(n40), .Z(n14161) );
  XNOR U14478 ( .A(n14169), .B(n14271), .Z(n14162) );
  XNOR U14479 ( .A(n14168), .B(n14166), .Z(n14271) );
  AND U14480 ( .A(n14272), .B(n14273), .Z(n14166) );
  NANDN U14481 ( .A(n14274), .B(n14275), .Z(n14273) );
  NAND U14482 ( .A(n14276), .B(n14277), .Z(n14275) );
  ANDN U14483 ( .B(B[199]), .A(n41), .Z(n14168) );
  XOR U14484 ( .A(n14175), .B(n14278), .Z(n14169) );
  XNOR U14485 ( .A(n14173), .B(n14176), .Z(n14278) );
  NAND U14486 ( .A(A[2]), .B(B[200]), .Z(n14176) );
  NANDN U14487 ( .A(n14279), .B(n14280), .Z(n14173) );
  AND U14488 ( .A(A[0]), .B(B[201]), .Z(n14280) );
  XNOR U14489 ( .A(n14178), .B(n14281), .Z(n14175) );
  NAND U14490 ( .A(A[0]), .B(B[202]), .Z(n14281) );
  NAND U14491 ( .A(B[201]), .B(A[1]), .Z(n14178) );
  NAND U14492 ( .A(n14282), .B(n14283), .Z(n341) );
  NANDN U14493 ( .A(n14284), .B(n14285), .Z(n14283) );
  OR U14494 ( .A(n14286), .B(n14287), .Z(n14285) );
  NAND U14495 ( .A(n14287), .B(n14286), .Z(n14282) );
  XOR U14496 ( .A(n14288), .B(n14289), .Z(\A1[1] ) );
  XNOR U14497 ( .A(n14290), .B(n14291), .Z(n14289) );
  XOR U14498 ( .A(n323), .B(n322), .Z(\A1[19] ) );
  XOR U14499 ( .A(n13277), .B(n14292), .Z(n322) );
  XNOR U14500 ( .A(n13276), .B(n13274), .Z(n14292) );
  AND U14501 ( .A(n14293), .B(n14294), .Z(n13274) );
  NANDN U14502 ( .A(n14295), .B(n14296), .Z(n14294) );
  NANDN U14503 ( .A(n14297), .B(n14298), .Z(n14296) );
  NANDN U14504 ( .A(n14298), .B(n14297), .Z(n14293) );
  ANDN U14505 ( .B(B[6]), .A(n29), .Z(n13276) );
  XNOR U14506 ( .A(n13183), .B(n14299), .Z(n13277) );
  XNOR U14507 ( .A(n13182), .B(n13180), .Z(n14299) );
  AND U14508 ( .A(n14300), .B(n14301), .Z(n13180) );
  NANDN U14509 ( .A(n14302), .B(n14303), .Z(n14301) );
  OR U14510 ( .A(n14304), .B(n14305), .Z(n14303) );
  NAND U14511 ( .A(n14305), .B(n14304), .Z(n14300) );
  ANDN U14512 ( .B(B[7]), .A(n30), .Z(n13182) );
  XNOR U14513 ( .A(n13190), .B(n14306), .Z(n13183) );
  XNOR U14514 ( .A(n13189), .B(n13187), .Z(n14306) );
  AND U14515 ( .A(n14307), .B(n14308), .Z(n13187) );
  NANDN U14516 ( .A(n14309), .B(n14310), .Z(n14308) );
  NANDN U14517 ( .A(n14311), .B(n14312), .Z(n14310) );
  NANDN U14518 ( .A(n14312), .B(n14311), .Z(n14307) );
  ANDN U14519 ( .B(B[8]), .A(n31), .Z(n13189) );
  XNOR U14520 ( .A(n13197), .B(n14313), .Z(n13190) );
  XNOR U14521 ( .A(n13196), .B(n13194), .Z(n14313) );
  AND U14522 ( .A(n14314), .B(n14315), .Z(n13194) );
  NANDN U14523 ( .A(n14316), .B(n14317), .Z(n14315) );
  OR U14524 ( .A(n14318), .B(n14319), .Z(n14317) );
  NAND U14525 ( .A(n14319), .B(n14318), .Z(n14314) );
  ANDN U14526 ( .B(B[9]), .A(n32), .Z(n13196) );
  XNOR U14527 ( .A(n13204), .B(n14320), .Z(n13197) );
  XNOR U14528 ( .A(n13203), .B(n13201), .Z(n14320) );
  AND U14529 ( .A(n14321), .B(n14322), .Z(n13201) );
  NANDN U14530 ( .A(n14323), .B(n14324), .Z(n14322) );
  NANDN U14531 ( .A(n14325), .B(n14326), .Z(n14324) );
  NANDN U14532 ( .A(n14326), .B(n14325), .Z(n14321) );
  ANDN U14533 ( .B(B[10]), .A(n33), .Z(n13203) );
  XNOR U14534 ( .A(n13211), .B(n14327), .Z(n13204) );
  XNOR U14535 ( .A(n13210), .B(n13208), .Z(n14327) );
  AND U14536 ( .A(n14328), .B(n14329), .Z(n13208) );
  NANDN U14537 ( .A(n14330), .B(n14331), .Z(n14329) );
  OR U14538 ( .A(n14332), .B(n14333), .Z(n14331) );
  NAND U14539 ( .A(n14333), .B(n14332), .Z(n14328) );
  ANDN U14540 ( .B(B[11]), .A(n34), .Z(n13210) );
  XNOR U14541 ( .A(n13218), .B(n14334), .Z(n13211) );
  XNOR U14542 ( .A(n13217), .B(n13215), .Z(n14334) );
  AND U14543 ( .A(n14335), .B(n14336), .Z(n13215) );
  NANDN U14544 ( .A(n14337), .B(n14338), .Z(n14336) );
  NANDN U14545 ( .A(n14339), .B(n14340), .Z(n14338) );
  NANDN U14546 ( .A(n14340), .B(n14339), .Z(n14335) );
  ANDN U14547 ( .B(B[12]), .A(n35), .Z(n13217) );
  XNOR U14548 ( .A(n13225), .B(n14341), .Z(n13218) );
  XNOR U14549 ( .A(n13224), .B(n13222), .Z(n14341) );
  AND U14550 ( .A(n14342), .B(n14343), .Z(n13222) );
  NANDN U14551 ( .A(n14344), .B(n14345), .Z(n14343) );
  OR U14552 ( .A(n14346), .B(n14347), .Z(n14345) );
  NAND U14553 ( .A(n14347), .B(n14346), .Z(n14342) );
  ANDN U14554 ( .B(B[13]), .A(n36), .Z(n13224) );
  XNOR U14555 ( .A(n13232), .B(n14348), .Z(n13225) );
  XNOR U14556 ( .A(n13231), .B(n13229), .Z(n14348) );
  AND U14557 ( .A(n14349), .B(n14350), .Z(n13229) );
  NANDN U14558 ( .A(n14351), .B(n14352), .Z(n14350) );
  NANDN U14559 ( .A(n14353), .B(n14354), .Z(n14352) );
  NANDN U14560 ( .A(n14354), .B(n14353), .Z(n14349) );
  ANDN U14561 ( .B(B[14]), .A(n37), .Z(n13231) );
  XNOR U14562 ( .A(n13239), .B(n14355), .Z(n13232) );
  XNOR U14563 ( .A(n13238), .B(n13236), .Z(n14355) );
  AND U14564 ( .A(n14356), .B(n14357), .Z(n13236) );
  NANDN U14565 ( .A(n14358), .B(n14359), .Z(n14357) );
  OR U14566 ( .A(n14360), .B(n14361), .Z(n14359) );
  NAND U14567 ( .A(n14361), .B(n14360), .Z(n14356) );
  ANDN U14568 ( .B(B[15]), .A(n38), .Z(n13238) );
  XNOR U14569 ( .A(n13246), .B(n14362), .Z(n13239) );
  XNOR U14570 ( .A(n13245), .B(n13243), .Z(n14362) );
  AND U14571 ( .A(n14363), .B(n14364), .Z(n13243) );
  NANDN U14572 ( .A(n14365), .B(n14366), .Z(n14364) );
  NANDN U14573 ( .A(n14367), .B(n14368), .Z(n14366) );
  NANDN U14574 ( .A(n14368), .B(n14367), .Z(n14363) );
  ANDN U14575 ( .B(B[16]), .A(n39), .Z(n13245) );
  XNOR U14576 ( .A(n13253), .B(n14369), .Z(n13246) );
  XNOR U14577 ( .A(n13252), .B(n13250), .Z(n14369) );
  AND U14578 ( .A(n14370), .B(n14371), .Z(n13250) );
  NANDN U14579 ( .A(n14372), .B(n14373), .Z(n14371) );
  OR U14580 ( .A(n14374), .B(n14375), .Z(n14373) );
  NAND U14581 ( .A(n14375), .B(n14374), .Z(n14370) );
  ANDN U14582 ( .B(B[17]), .A(n40), .Z(n13252) );
  XNOR U14583 ( .A(n13260), .B(n14376), .Z(n13253) );
  XNOR U14584 ( .A(n13259), .B(n13257), .Z(n14376) );
  AND U14585 ( .A(n14377), .B(n14378), .Z(n13257) );
  NANDN U14586 ( .A(n14379), .B(n14380), .Z(n14378) );
  NAND U14587 ( .A(n14381), .B(n14382), .Z(n14380) );
  ANDN U14588 ( .B(B[18]), .A(n41), .Z(n13259) );
  XOR U14589 ( .A(n13266), .B(n14383), .Z(n13260) );
  XNOR U14590 ( .A(n13264), .B(n13267), .Z(n14383) );
  NAND U14591 ( .A(A[2]), .B(B[19]), .Z(n13267) );
  NANDN U14592 ( .A(n14384), .B(n14385), .Z(n13264) );
  AND U14593 ( .A(A[0]), .B(B[20]), .Z(n14385) );
  XNOR U14594 ( .A(n13269), .B(n14386), .Z(n13266) );
  NAND U14595 ( .A(A[0]), .B(B[21]), .Z(n14386) );
  NAND U14596 ( .A(B[20]), .B(A[1]), .Z(n13269) );
  NAND U14597 ( .A(n14387), .B(n14388), .Z(n323) );
  NANDN U14598 ( .A(n14389), .B(n14390), .Z(n14388) );
  OR U14599 ( .A(n14391), .B(n14392), .Z(n14390) );
  NAND U14600 ( .A(n14392), .B(n14391), .Z(n14387) );
  XOR U14601 ( .A(n343), .B(n342), .Z(\A1[199] ) );
  XOR U14602 ( .A(n14287), .B(n14393), .Z(n342) );
  XNOR U14603 ( .A(n14286), .B(n14284), .Z(n14393) );
  AND U14604 ( .A(n14394), .B(n14395), .Z(n14284) );
  NANDN U14605 ( .A(n14396), .B(n14397), .Z(n14395) );
  NANDN U14606 ( .A(n14398), .B(n14399), .Z(n14397) );
  NANDN U14607 ( .A(n14399), .B(n14398), .Z(n14394) );
  ANDN U14608 ( .B(B[186]), .A(n29), .Z(n14286) );
  XNOR U14609 ( .A(n14193), .B(n14400), .Z(n14287) );
  XNOR U14610 ( .A(n14192), .B(n14190), .Z(n14400) );
  AND U14611 ( .A(n14401), .B(n14402), .Z(n14190) );
  NANDN U14612 ( .A(n14403), .B(n14404), .Z(n14402) );
  OR U14613 ( .A(n14405), .B(n14406), .Z(n14404) );
  NAND U14614 ( .A(n14406), .B(n14405), .Z(n14401) );
  ANDN U14615 ( .B(B[187]), .A(n30), .Z(n14192) );
  XNOR U14616 ( .A(n14200), .B(n14407), .Z(n14193) );
  XNOR U14617 ( .A(n14199), .B(n14197), .Z(n14407) );
  AND U14618 ( .A(n14408), .B(n14409), .Z(n14197) );
  NANDN U14619 ( .A(n14410), .B(n14411), .Z(n14409) );
  NANDN U14620 ( .A(n14412), .B(n14413), .Z(n14411) );
  NANDN U14621 ( .A(n14413), .B(n14412), .Z(n14408) );
  ANDN U14622 ( .B(B[188]), .A(n31), .Z(n14199) );
  XNOR U14623 ( .A(n14207), .B(n14414), .Z(n14200) );
  XNOR U14624 ( .A(n14206), .B(n14204), .Z(n14414) );
  AND U14625 ( .A(n14415), .B(n14416), .Z(n14204) );
  NANDN U14626 ( .A(n14417), .B(n14418), .Z(n14416) );
  OR U14627 ( .A(n14419), .B(n14420), .Z(n14418) );
  NAND U14628 ( .A(n14420), .B(n14419), .Z(n14415) );
  ANDN U14629 ( .B(B[189]), .A(n32), .Z(n14206) );
  XNOR U14630 ( .A(n14214), .B(n14421), .Z(n14207) );
  XNOR U14631 ( .A(n14213), .B(n14211), .Z(n14421) );
  AND U14632 ( .A(n14422), .B(n14423), .Z(n14211) );
  NANDN U14633 ( .A(n14424), .B(n14425), .Z(n14423) );
  NANDN U14634 ( .A(n14426), .B(n14427), .Z(n14425) );
  NANDN U14635 ( .A(n14427), .B(n14426), .Z(n14422) );
  ANDN U14636 ( .B(B[190]), .A(n33), .Z(n14213) );
  XNOR U14637 ( .A(n14221), .B(n14428), .Z(n14214) );
  XNOR U14638 ( .A(n14220), .B(n14218), .Z(n14428) );
  AND U14639 ( .A(n14429), .B(n14430), .Z(n14218) );
  NANDN U14640 ( .A(n14431), .B(n14432), .Z(n14430) );
  OR U14641 ( .A(n14433), .B(n14434), .Z(n14432) );
  NAND U14642 ( .A(n14434), .B(n14433), .Z(n14429) );
  ANDN U14643 ( .B(B[191]), .A(n34), .Z(n14220) );
  XNOR U14644 ( .A(n14228), .B(n14435), .Z(n14221) );
  XNOR U14645 ( .A(n14227), .B(n14225), .Z(n14435) );
  AND U14646 ( .A(n14436), .B(n14437), .Z(n14225) );
  NANDN U14647 ( .A(n14438), .B(n14439), .Z(n14437) );
  NANDN U14648 ( .A(n14440), .B(n14441), .Z(n14439) );
  NANDN U14649 ( .A(n14441), .B(n14440), .Z(n14436) );
  ANDN U14650 ( .B(B[192]), .A(n35), .Z(n14227) );
  XNOR U14651 ( .A(n14235), .B(n14442), .Z(n14228) );
  XNOR U14652 ( .A(n14234), .B(n14232), .Z(n14442) );
  AND U14653 ( .A(n14443), .B(n14444), .Z(n14232) );
  NANDN U14654 ( .A(n14445), .B(n14446), .Z(n14444) );
  OR U14655 ( .A(n14447), .B(n14448), .Z(n14446) );
  NAND U14656 ( .A(n14448), .B(n14447), .Z(n14443) );
  ANDN U14657 ( .B(B[193]), .A(n36), .Z(n14234) );
  XNOR U14658 ( .A(n14242), .B(n14449), .Z(n14235) );
  XNOR U14659 ( .A(n14241), .B(n14239), .Z(n14449) );
  AND U14660 ( .A(n14450), .B(n14451), .Z(n14239) );
  NANDN U14661 ( .A(n14452), .B(n14453), .Z(n14451) );
  NANDN U14662 ( .A(n14454), .B(n14455), .Z(n14453) );
  NANDN U14663 ( .A(n14455), .B(n14454), .Z(n14450) );
  ANDN U14664 ( .B(B[194]), .A(n37), .Z(n14241) );
  XNOR U14665 ( .A(n14249), .B(n14456), .Z(n14242) );
  XNOR U14666 ( .A(n14248), .B(n14246), .Z(n14456) );
  AND U14667 ( .A(n14457), .B(n14458), .Z(n14246) );
  NANDN U14668 ( .A(n14459), .B(n14460), .Z(n14458) );
  OR U14669 ( .A(n14461), .B(n14462), .Z(n14460) );
  NAND U14670 ( .A(n14462), .B(n14461), .Z(n14457) );
  ANDN U14671 ( .B(B[195]), .A(n38), .Z(n14248) );
  XNOR U14672 ( .A(n14256), .B(n14463), .Z(n14249) );
  XNOR U14673 ( .A(n14255), .B(n14253), .Z(n14463) );
  AND U14674 ( .A(n14464), .B(n14465), .Z(n14253) );
  NANDN U14675 ( .A(n14466), .B(n14467), .Z(n14465) );
  NANDN U14676 ( .A(n14468), .B(n14469), .Z(n14467) );
  NANDN U14677 ( .A(n14469), .B(n14468), .Z(n14464) );
  ANDN U14678 ( .B(B[196]), .A(n39), .Z(n14255) );
  XNOR U14679 ( .A(n14263), .B(n14470), .Z(n14256) );
  XNOR U14680 ( .A(n14262), .B(n14260), .Z(n14470) );
  AND U14681 ( .A(n14471), .B(n14472), .Z(n14260) );
  NANDN U14682 ( .A(n14473), .B(n14474), .Z(n14472) );
  OR U14683 ( .A(n14475), .B(n14476), .Z(n14474) );
  NAND U14684 ( .A(n14476), .B(n14475), .Z(n14471) );
  ANDN U14685 ( .B(B[197]), .A(n40), .Z(n14262) );
  XNOR U14686 ( .A(n14270), .B(n14477), .Z(n14263) );
  XNOR U14687 ( .A(n14269), .B(n14267), .Z(n14477) );
  AND U14688 ( .A(n14478), .B(n14479), .Z(n14267) );
  NANDN U14689 ( .A(n14480), .B(n14481), .Z(n14479) );
  NAND U14690 ( .A(n14482), .B(n14483), .Z(n14481) );
  ANDN U14691 ( .B(B[198]), .A(n41), .Z(n14269) );
  XOR U14692 ( .A(n14276), .B(n14484), .Z(n14270) );
  XNOR U14693 ( .A(n14274), .B(n14277), .Z(n14484) );
  NAND U14694 ( .A(A[2]), .B(B[199]), .Z(n14277) );
  NANDN U14695 ( .A(n14485), .B(n14486), .Z(n14274) );
  AND U14696 ( .A(A[0]), .B(B[200]), .Z(n14486) );
  XNOR U14697 ( .A(n14279), .B(n14487), .Z(n14276) );
  NAND U14698 ( .A(A[0]), .B(B[201]), .Z(n14487) );
  NAND U14699 ( .A(B[200]), .B(A[1]), .Z(n14279) );
  NAND U14700 ( .A(n14488), .B(n14489), .Z(n343) );
  NANDN U14701 ( .A(n14490), .B(n14491), .Z(n14489) );
  OR U14702 ( .A(n14492), .B(n14493), .Z(n14491) );
  NAND U14703 ( .A(n14493), .B(n14492), .Z(n14488) );
  XOR U14704 ( .A(n347), .B(n346), .Z(\A1[198] ) );
  XOR U14705 ( .A(n14493), .B(n14494), .Z(n346) );
  XNOR U14706 ( .A(n14492), .B(n14490), .Z(n14494) );
  AND U14707 ( .A(n14495), .B(n14496), .Z(n14490) );
  NANDN U14708 ( .A(n14497), .B(n14498), .Z(n14496) );
  NANDN U14709 ( .A(n14499), .B(n14500), .Z(n14498) );
  NANDN U14710 ( .A(n14500), .B(n14499), .Z(n14495) );
  ANDN U14711 ( .B(B[185]), .A(n29), .Z(n14492) );
  XNOR U14712 ( .A(n14399), .B(n14501), .Z(n14493) );
  XNOR U14713 ( .A(n14398), .B(n14396), .Z(n14501) );
  AND U14714 ( .A(n14502), .B(n14503), .Z(n14396) );
  NANDN U14715 ( .A(n14504), .B(n14505), .Z(n14503) );
  OR U14716 ( .A(n14506), .B(n14507), .Z(n14505) );
  NAND U14717 ( .A(n14507), .B(n14506), .Z(n14502) );
  ANDN U14718 ( .B(B[186]), .A(n30), .Z(n14398) );
  XNOR U14719 ( .A(n14406), .B(n14508), .Z(n14399) );
  XNOR U14720 ( .A(n14405), .B(n14403), .Z(n14508) );
  AND U14721 ( .A(n14509), .B(n14510), .Z(n14403) );
  NANDN U14722 ( .A(n14511), .B(n14512), .Z(n14510) );
  NANDN U14723 ( .A(n14513), .B(n14514), .Z(n14512) );
  NANDN U14724 ( .A(n14514), .B(n14513), .Z(n14509) );
  ANDN U14725 ( .B(B[187]), .A(n31), .Z(n14405) );
  XNOR U14726 ( .A(n14413), .B(n14515), .Z(n14406) );
  XNOR U14727 ( .A(n14412), .B(n14410), .Z(n14515) );
  AND U14728 ( .A(n14516), .B(n14517), .Z(n14410) );
  NANDN U14729 ( .A(n14518), .B(n14519), .Z(n14517) );
  OR U14730 ( .A(n14520), .B(n14521), .Z(n14519) );
  NAND U14731 ( .A(n14521), .B(n14520), .Z(n14516) );
  ANDN U14732 ( .B(B[188]), .A(n32), .Z(n14412) );
  XNOR U14733 ( .A(n14420), .B(n14522), .Z(n14413) );
  XNOR U14734 ( .A(n14419), .B(n14417), .Z(n14522) );
  AND U14735 ( .A(n14523), .B(n14524), .Z(n14417) );
  NANDN U14736 ( .A(n14525), .B(n14526), .Z(n14524) );
  NANDN U14737 ( .A(n14527), .B(n14528), .Z(n14526) );
  NANDN U14738 ( .A(n14528), .B(n14527), .Z(n14523) );
  ANDN U14739 ( .B(B[189]), .A(n33), .Z(n14419) );
  XNOR U14740 ( .A(n14427), .B(n14529), .Z(n14420) );
  XNOR U14741 ( .A(n14426), .B(n14424), .Z(n14529) );
  AND U14742 ( .A(n14530), .B(n14531), .Z(n14424) );
  NANDN U14743 ( .A(n14532), .B(n14533), .Z(n14531) );
  OR U14744 ( .A(n14534), .B(n14535), .Z(n14533) );
  NAND U14745 ( .A(n14535), .B(n14534), .Z(n14530) );
  ANDN U14746 ( .B(B[190]), .A(n34), .Z(n14426) );
  XNOR U14747 ( .A(n14434), .B(n14536), .Z(n14427) );
  XNOR U14748 ( .A(n14433), .B(n14431), .Z(n14536) );
  AND U14749 ( .A(n14537), .B(n14538), .Z(n14431) );
  NANDN U14750 ( .A(n14539), .B(n14540), .Z(n14538) );
  NANDN U14751 ( .A(n14541), .B(n14542), .Z(n14540) );
  NANDN U14752 ( .A(n14542), .B(n14541), .Z(n14537) );
  ANDN U14753 ( .B(B[191]), .A(n35), .Z(n14433) );
  XNOR U14754 ( .A(n14441), .B(n14543), .Z(n14434) );
  XNOR U14755 ( .A(n14440), .B(n14438), .Z(n14543) );
  AND U14756 ( .A(n14544), .B(n14545), .Z(n14438) );
  NANDN U14757 ( .A(n14546), .B(n14547), .Z(n14545) );
  OR U14758 ( .A(n14548), .B(n14549), .Z(n14547) );
  NAND U14759 ( .A(n14549), .B(n14548), .Z(n14544) );
  ANDN U14760 ( .B(B[192]), .A(n36), .Z(n14440) );
  XNOR U14761 ( .A(n14448), .B(n14550), .Z(n14441) );
  XNOR U14762 ( .A(n14447), .B(n14445), .Z(n14550) );
  AND U14763 ( .A(n14551), .B(n14552), .Z(n14445) );
  NANDN U14764 ( .A(n14553), .B(n14554), .Z(n14552) );
  NANDN U14765 ( .A(n14555), .B(n14556), .Z(n14554) );
  NANDN U14766 ( .A(n14556), .B(n14555), .Z(n14551) );
  ANDN U14767 ( .B(B[193]), .A(n37), .Z(n14447) );
  XNOR U14768 ( .A(n14455), .B(n14557), .Z(n14448) );
  XNOR U14769 ( .A(n14454), .B(n14452), .Z(n14557) );
  AND U14770 ( .A(n14558), .B(n14559), .Z(n14452) );
  NANDN U14771 ( .A(n14560), .B(n14561), .Z(n14559) );
  OR U14772 ( .A(n14562), .B(n14563), .Z(n14561) );
  NAND U14773 ( .A(n14563), .B(n14562), .Z(n14558) );
  ANDN U14774 ( .B(B[194]), .A(n38), .Z(n14454) );
  XNOR U14775 ( .A(n14462), .B(n14564), .Z(n14455) );
  XNOR U14776 ( .A(n14461), .B(n14459), .Z(n14564) );
  AND U14777 ( .A(n14565), .B(n14566), .Z(n14459) );
  NANDN U14778 ( .A(n14567), .B(n14568), .Z(n14566) );
  NANDN U14779 ( .A(n14569), .B(n14570), .Z(n14568) );
  NANDN U14780 ( .A(n14570), .B(n14569), .Z(n14565) );
  ANDN U14781 ( .B(B[195]), .A(n39), .Z(n14461) );
  XNOR U14782 ( .A(n14469), .B(n14571), .Z(n14462) );
  XNOR U14783 ( .A(n14468), .B(n14466), .Z(n14571) );
  AND U14784 ( .A(n14572), .B(n14573), .Z(n14466) );
  NANDN U14785 ( .A(n14574), .B(n14575), .Z(n14573) );
  OR U14786 ( .A(n14576), .B(n14577), .Z(n14575) );
  NAND U14787 ( .A(n14577), .B(n14576), .Z(n14572) );
  ANDN U14788 ( .B(B[196]), .A(n40), .Z(n14468) );
  XNOR U14789 ( .A(n14476), .B(n14578), .Z(n14469) );
  XNOR U14790 ( .A(n14475), .B(n14473), .Z(n14578) );
  AND U14791 ( .A(n14579), .B(n14580), .Z(n14473) );
  NANDN U14792 ( .A(n14581), .B(n14582), .Z(n14580) );
  NAND U14793 ( .A(n14583), .B(n14584), .Z(n14582) );
  ANDN U14794 ( .B(B[197]), .A(n41), .Z(n14475) );
  XOR U14795 ( .A(n14482), .B(n14585), .Z(n14476) );
  XNOR U14796 ( .A(n14480), .B(n14483), .Z(n14585) );
  NAND U14797 ( .A(A[2]), .B(B[198]), .Z(n14483) );
  NANDN U14798 ( .A(n14586), .B(n14587), .Z(n14480) );
  AND U14799 ( .A(A[0]), .B(B[199]), .Z(n14587) );
  XNOR U14800 ( .A(n14485), .B(n14588), .Z(n14482) );
  NAND U14801 ( .A(A[0]), .B(B[200]), .Z(n14588) );
  NAND U14802 ( .A(B[199]), .B(A[1]), .Z(n14485) );
  NAND U14803 ( .A(n14589), .B(n14590), .Z(n347) );
  NANDN U14804 ( .A(n14591), .B(n14592), .Z(n14590) );
  OR U14805 ( .A(n14593), .B(n14594), .Z(n14592) );
  NAND U14806 ( .A(n14594), .B(n14593), .Z(n14589) );
  XOR U14807 ( .A(n349), .B(n348), .Z(\A1[197] ) );
  XOR U14808 ( .A(n14594), .B(n14595), .Z(n348) );
  XNOR U14809 ( .A(n14593), .B(n14591), .Z(n14595) );
  AND U14810 ( .A(n14596), .B(n14597), .Z(n14591) );
  NANDN U14811 ( .A(n14598), .B(n14599), .Z(n14597) );
  NANDN U14812 ( .A(n14600), .B(n14601), .Z(n14599) );
  NANDN U14813 ( .A(n14601), .B(n14600), .Z(n14596) );
  ANDN U14814 ( .B(B[184]), .A(n29), .Z(n14593) );
  XNOR U14815 ( .A(n14500), .B(n14602), .Z(n14594) );
  XNOR U14816 ( .A(n14499), .B(n14497), .Z(n14602) );
  AND U14817 ( .A(n14603), .B(n14604), .Z(n14497) );
  NANDN U14818 ( .A(n14605), .B(n14606), .Z(n14604) );
  OR U14819 ( .A(n14607), .B(n14608), .Z(n14606) );
  NAND U14820 ( .A(n14608), .B(n14607), .Z(n14603) );
  ANDN U14821 ( .B(B[185]), .A(n30), .Z(n14499) );
  XNOR U14822 ( .A(n14507), .B(n14609), .Z(n14500) );
  XNOR U14823 ( .A(n14506), .B(n14504), .Z(n14609) );
  AND U14824 ( .A(n14610), .B(n14611), .Z(n14504) );
  NANDN U14825 ( .A(n14612), .B(n14613), .Z(n14611) );
  NANDN U14826 ( .A(n14614), .B(n14615), .Z(n14613) );
  NANDN U14827 ( .A(n14615), .B(n14614), .Z(n14610) );
  ANDN U14828 ( .B(B[186]), .A(n31), .Z(n14506) );
  XNOR U14829 ( .A(n14514), .B(n14616), .Z(n14507) );
  XNOR U14830 ( .A(n14513), .B(n14511), .Z(n14616) );
  AND U14831 ( .A(n14617), .B(n14618), .Z(n14511) );
  NANDN U14832 ( .A(n14619), .B(n14620), .Z(n14618) );
  OR U14833 ( .A(n14621), .B(n14622), .Z(n14620) );
  NAND U14834 ( .A(n14622), .B(n14621), .Z(n14617) );
  ANDN U14835 ( .B(B[187]), .A(n32), .Z(n14513) );
  XNOR U14836 ( .A(n14521), .B(n14623), .Z(n14514) );
  XNOR U14837 ( .A(n14520), .B(n14518), .Z(n14623) );
  AND U14838 ( .A(n14624), .B(n14625), .Z(n14518) );
  NANDN U14839 ( .A(n14626), .B(n14627), .Z(n14625) );
  NANDN U14840 ( .A(n14628), .B(n14629), .Z(n14627) );
  NANDN U14841 ( .A(n14629), .B(n14628), .Z(n14624) );
  ANDN U14842 ( .B(B[188]), .A(n33), .Z(n14520) );
  XNOR U14843 ( .A(n14528), .B(n14630), .Z(n14521) );
  XNOR U14844 ( .A(n14527), .B(n14525), .Z(n14630) );
  AND U14845 ( .A(n14631), .B(n14632), .Z(n14525) );
  NANDN U14846 ( .A(n14633), .B(n14634), .Z(n14632) );
  OR U14847 ( .A(n14635), .B(n14636), .Z(n14634) );
  NAND U14848 ( .A(n14636), .B(n14635), .Z(n14631) );
  ANDN U14849 ( .B(B[189]), .A(n34), .Z(n14527) );
  XNOR U14850 ( .A(n14535), .B(n14637), .Z(n14528) );
  XNOR U14851 ( .A(n14534), .B(n14532), .Z(n14637) );
  AND U14852 ( .A(n14638), .B(n14639), .Z(n14532) );
  NANDN U14853 ( .A(n14640), .B(n14641), .Z(n14639) );
  NANDN U14854 ( .A(n14642), .B(n14643), .Z(n14641) );
  NANDN U14855 ( .A(n14643), .B(n14642), .Z(n14638) );
  ANDN U14856 ( .B(B[190]), .A(n35), .Z(n14534) );
  XNOR U14857 ( .A(n14542), .B(n14644), .Z(n14535) );
  XNOR U14858 ( .A(n14541), .B(n14539), .Z(n14644) );
  AND U14859 ( .A(n14645), .B(n14646), .Z(n14539) );
  NANDN U14860 ( .A(n14647), .B(n14648), .Z(n14646) );
  OR U14861 ( .A(n14649), .B(n14650), .Z(n14648) );
  NAND U14862 ( .A(n14650), .B(n14649), .Z(n14645) );
  ANDN U14863 ( .B(B[191]), .A(n36), .Z(n14541) );
  XNOR U14864 ( .A(n14549), .B(n14651), .Z(n14542) );
  XNOR U14865 ( .A(n14548), .B(n14546), .Z(n14651) );
  AND U14866 ( .A(n14652), .B(n14653), .Z(n14546) );
  NANDN U14867 ( .A(n14654), .B(n14655), .Z(n14653) );
  NANDN U14868 ( .A(n14656), .B(n14657), .Z(n14655) );
  NANDN U14869 ( .A(n14657), .B(n14656), .Z(n14652) );
  ANDN U14870 ( .B(B[192]), .A(n37), .Z(n14548) );
  XNOR U14871 ( .A(n14556), .B(n14658), .Z(n14549) );
  XNOR U14872 ( .A(n14555), .B(n14553), .Z(n14658) );
  AND U14873 ( .A(n14659), .B(n14660), .Z(n14553) );
  NANDN U14874 ( .A(n14661), .B(n14662), .Z(n14660) );
  OR U14875 ( .A(n14663), .B(n14664), .Z(n14662) );
  NAND U14876 ( .A(n14664), .B(n14663), .Z(n14659) );
  ANDN U14877 ( .B(B[193]), .A(n38), .Z(n14555) );
  XNOR U14878 ( .A(n14563), .B(n14665), .Z(n14556) );
  XNOR U14879 ( .A(n14562), .B(n14560), .Z(n14665) );
  AND U14880 ( .A(n14666), .B(n14667), .Z(n14560) );
  NANDN U14881 ( .A(n14668), .B(n14669), .Z(n14667) );
  NANDN U14882 ( .A(n14670), .B(n14671), .Z(n14669) );
  NANDN U14883 ( .A(n14671), .B(n14670), .Z(n14666) );
  ANDN U14884 ( .B(B[194]), .A(n39), .Z(n14562) );
  XNOR U14885 ( .A(n14570), .B(n14672), .Z(n14563) );
  XNOR U14886 ( .A(n14569), .B(n14567), .Z(n14672) );
  AND U14887 ( .A(n14673), .B(n14674), .Z(n14567) );
  NANDN U14888 ( .A(n14675), .B(n14676), .Z(n14674) );
  OR U14889 ( .A(n14677), .B(n14678), .Z(n14676) );
  NAND U14890 ( .A(n14678), .B(n14677), .Z(n14673) );
  ANDN U14891 ( .B(B[195]), .A(n40), .Z(n14569) );
  XNOR U14892 ( .A(n14577), .B(n14679), .Z(n14570) );
  XNOR U14893 ( .A(n14576), .B(n14574), .Z(n14679) );
  AND U14894 ( .A(n14680), .B(n14681), .Z(n14574) );
  NANDN U14895 ( .A(n14682), .B(n14683), .Z(n14681) );
  NAND U14896 ( .A(n14684), .B(n14685), .Z(n14683) );
  ANDN U14897 ( .B(B[196]), .A(n41), .Z(n14576) );
  XOR U14898 ( .A(n14583), .B(n14686), .Z(n14577) );
  XNOR U14899 ( .A(n14581), .B(n14584), .Z(n14686) );
  NAND U14900 ( .A(A[2]), .B(B[197]), .Z(n14584) );
  NANDN U14901 ( .A(n14687), .B(n14688), .Z(n14581) );
  AND U14902 ( .A(A[0]), .B(B[198]), .Z(n14688) );
  XNOR U14903 ( .A(n14586), .B(n14689), .Z(n14583) );
  NAND U14904 ( .A(A[0]), .B(B[199]), .Z(n14689) );
  NAND U14905 ( .A(B[198]), .B(A[1]), .Z(n14586) );
  NAND U14906 ( .A(n14690), .B(n14691), .Z(n349) );
  NANDN U14907 ( .A(n14692), .B(n14693), .Z(n14691) );
  OR U14908 ( .A(n14694), .B(n14695), .Z(n14693) );
  NAND U14909 ( .A(n14695), .B(n14694), .Z(n14690) );
  XOR U14910 ( .A(n351), .B(n350), .Z(\A1[196] ) );
  XOR U14911 ( .A(n14695), .B(n14696), .Z(n350) );
  XNOR U14912 ( .A(n14694), .B(n14692), .Z(n14696) );
  AND U14913 ( .A(n14697), .B(n14698), .Z(n14692) );
  NANDN U14914 ( .A(n14699), .B(n14700), .Z(n14698) );
  NANDN U14915 ( .A(n14701), .B(n14702), .Z(n14700) );
  NANDN U14916 ( .A(n14702), .B(n14701), .Z(n14697) );
  ANDN U14917 ( .B(B[183]), .A(n29), .Z(n14694) );
  XNOR U14918 ( .A(n14601), .B(n14703), .Z(n14695) );
  XNOR U14919 ( .A(n14600), .B(n14598), .Z(n14703) );
  AND U14920 ( .A(n14704), .B(n14705), .Z(n14598) );
  NANDN U14921 ( .A(n14706), .B(n14707), .Z(n14705) );
  OR U14922 ( .A(n14708), .B(n14709), .Z(n14707) );
  NAND U14923 ( .A(n14709), .B(n14708), .Z(n14704) );
  ANDN U14924 ( .B(B[184]), .A(n30), .Z(n14600) );
  XNOR U14925 ( .A(n14608), .B(n14710), .Z(n14601) );
  XNOR U14926 ( .A(n14607), .B(n14605), .Z(n14710) );
  AND U14927 ( .A(n14711), .B(n14712), .Z(n14605) );
  NANDN U14928 ( .A(n14713), .B(n14714), .Z(n14712) );
  NANDN U14929 ( .A(n14715), .B(n14716), .Z(n14714) );
  NANDN U14930 ( .A(n14716), .B(n14715), .Z(n14711) );
  ANDN U14931 ( .B(B[185]), .A(n31), .Z(n14607) );
  XNOR U14932 ( .A(n14615), .B(n14717), .Z(n14608) );
  XNOR U14933 ( .A(n14614), .B(n14612), .Z(n14717) );
  AND U14934 ( .A(n14718), .B(n14719), .Z(n14612) );
  NANDN U14935 ( .A(n14720), .B(n14721), .Z(n14719) );
  OR U14936 ( .A(n14722), .B(n14723), .Z(n14721) );
  NAND U14937 ( .A(n14723), .B(n14722), .Z(n14718) );
  ANDN U14938 ( .B(B[186]), .A(n32), .Z(n14614) );
  XNOR U14939 ( .A(n14622), .B(n14724), .Z(n14615) );
  XNOR U14940 ( .A(n14621), .B(n14619), .Z(n14724) );
  AND U14941 ( .A(n14725), .B(n14726), .Z(n14619) );
  NANDN U14942 ( .A(n14727), .B(n14728), .Z(n14726) );
  NANDN U14943 ( .A(n14729), .B(n14730), .Z(n14728) );
  NANDN U14944 ( .A(n14730), .B(n14729), .Z(n14725) );
  ANDN U14945 ( .B(B[187]), .A(n33), .Z(n14621) );
  XNOR U14946 ( .A(n14629), .B(n14731), .Z(n14622) );
  XNOR U14947 ( .A(n14628), .B(n14626), .Z(n14731) );
  AND U14948 ( .A(n14732), .B(n14733), .Z(n14626) );
  NANDN U14949 ( .A(n14734), .B(n14735), .Z(n14733) );
  OR U14950 ( .A(n14736), .B(n14737), .Z(n14735) );
  NAND U14951 ( .A(n14737), .B(n14736), .Z(n14732) );
  ANDN U14952 ( .B(B[188]), .A(n34), .Z(n14628) );
  XNOR U14953 ( .A(n14636), .B(n14738), .Z(n14629) );
  XNOR U14954 ( .A(n14635), .B(n14633), .Z(n14738) );
  AND U14955 ( .A(n14739), .B(n14740), .Z(n14633) );
  NANDN U14956 ( .A(n14741), .B(n14742), .Z(n14740) );
  NANDN U14957 ( .A(n14743), .B(n14744), .Z(n14742) );
  NANDN U14958 ( .A(n14744), .B(n14743), .Z(n14739) );
  ANDN U14959 ( .B(B[189]), .A(n35), .Z(n14635) );
  XNOR U14960 ( .A(n14643), .B(n14745), .Z(n14636) );
  XNOR U14961 ( .A(n14642), .B(n14640), .Z(n14745) );
  AND U14962 ( .A(n14746), .B(n14747), .Z(n14640) );
  NANDN U14963 ( .A(n14748), .B(n14749), .Z(n14747) );
  OR U14964 ( .A(n14750), .B(n14751), .Z(n14749) );
  NAND U14965 ( .A(n14751), .B(n14750), .Z(n14746) );
  ANDN U14966 ( .B(B[190]), .A(n36), .Z(n14642) );
  XNOR U14967 ( .A(n14650), .B(n14752), .Z(n14643) );
  XNOR U14968 ( .A(n14649), .B(n14647), .Z(n14752) );
  AND U14969 ( .A(n14753), .B(n14754), .Z(n14647) );
  NANDN U14970 ( .A(n14755), .B(n14756), .Z(n14754) );
  NANDN U14971 ( .A(n14757), .B(n14758), .Z(n14756) );
  NANDN U14972 ( .A(n14758), .B(n14757), .Z(n14753) );
  ANDN U14973 ( .B(B[191]), .A(n37), .Z(n14649) );
  XNOR U14974 ( .A(n14657), .B(n14759), .Z(n14650) );
  XNOR U14975 ( .A(n14656), .B(n14654), .Z(n14759) );
  AND U14976 ( .A(n14760), .B(n14761), .Z(n14654) );
  NANDN U14977 ( .A(n14762), .B(n14763), .Z(n14761) );
  OR U14978 ( .A(n14764), .B(n14765), .Z(n14763) );
  NAND U14979 ( .A(n14765), .B(n14764), .Z(n14760) );
  ANDN U14980 ( .B(B[192]), .A(n38), .Z(n14656) );
  XNOR U14981 ( .A(n14664), .B(n14766), .Z(n14657) );
  XNOR U14982 ( .A(n14663), .B(n14661), .Z(n14766) );
  AND U14983 ( .A(n14767), .B(n14768), .Z(n14661) );
  NANDN U14984 ( .A(n14769), .B(n14770), .Z(n14768) );
  NANDN U14985 ( .A(n14771), .B(n14772), .Z(n14770) );
  NANDN U14986 ( .A(n14772), .B(n14771), .Z(n14767) );
  ANDN U14987 ( .B(B[193]), .A(n39), .Z(n14663) );
  XNOR U14988 ( .A(n14671), .B(n14773), .Z(n14664) );
  XNOR U14989 ( .A(n14670), .B(n14668), .Z(n14773) );
  AND U14990 ( .A(n14774), .B(n14775), .Z(n14668) );
  NANDN U14991 ( .A(n14776), .B(n14777), .Z(n14775) );
  OR U14992 ( .A(n14778), .B(n14779), .Z(n14777) );
  NAND U14993 ( .A(n14779), .B(n14778), .Z(n14774) );
  ANDN U14994 ( .B(B[194]), .A(n40), .Z(n14670) );
  XNOR U14995 ( .A(n14678), .B(n14780), .Z(n14671) );
  XNOR U14996 ( .A(n14677), .B(n14675), .Z(n14780) );
  AND U14997 ( .A(n14781), .B(n14782), .Z(n14675) );
  NANDN U14998 ( .A(n14783), .B(n14784), .Z(n14782) );
  NAND U14999 ( .A(n14785), .B(n14786), .Z(n14784) );
  ANDN U15000 ( .B(B[195]), .A(n41), .Z(n14677) );
  XOR U15001 ( .A(n14684), .B(n14787), .Z(n14678) );
  XNOR U15002 ( .A(n14682), .B(n14685), .Z(n14787) );
  NAND U15003 ( .A(A[2]), .B(B[196]), .Z(n14685) );
  NANDN U15004 ( .A(n14788), .B(n14789), .Z(n14682) );
  AND U15005 ( .A(A[0]), .B(B[197]), .Z(n14789) );
  XNOR U15006 ( .A(n14687), .B(n14790), .Z(n14684) );
  NAND U15007 ( .A(A[0]), .B(B[198]), .Z(n14790) );
  NAND U15008 ( .A(B[197]), .B(A[1]), .Z(n14687) );
  NAND U15009 ( .A(n14791), .B(n14792), .Z(n351) );
  NANDN U15010 ( .A(n14793), .B(n14794), .Z(n14792) );
  OR U15011 ( .A(n14795), .B(n14796), .Z(n14794) );
  NAND U15012 ( .A(n14796), .B(n14795), .Z(n14791) );
  XOR U15013 ( .A(n353), .B(n352), .Z(\A1[195] ) );
  XOR U15014 ( .A(n14796), .B(n14797), .Z(n352) );
  XNOR U15015 ( .A(n14795), .B(n14793), .Z(n14797) );
  AND U15016 ( .A(n14798), .B(n14799), .Z(n14793) );
  NANDN U15017 ( .A(n14800), .B(n14801), .Z(n14799) );
  NANDN U15018 ( .A(n14802), .B(n14803), .Z(n14801) );
  NANDN U15019 ( .A(n14803), .B(n14802), .Z(n14798) );
  ANDN U15020 ( .B(B[182]), .A(n29), .Z(n14795) );
  XNOR U15021 ( .A(n14702), .B(n14804), .Z(n14796) );
  XNOR U15022 ( .A(n14701), .B(n14699), .Z(n14804) );
  AND U15023 ( .A(n14805), .B(n14806), .Z(n14699) );
  NANDN U15024 ( .A(n14807), .B(n14808), .Z(n14806) );
  OR U15025 ( .A(n14809), .B(n14810), .Z(n14808) );
  NAND U15026 ( .A(n14810), .B(n14809), .Z(n14805) );
  ANDN U15027 ( .B(B[183]), .A(n30), .Z(n14701) );
  XNOR U15028 ( .A(n14709), .B(n14811), .Z(n14702) );
  XNOR U15029 ( .A(n14708), .B(n14706), .Z(n14811) );
  AND U15030 ( .A(n14812), .B(n14813), .Z(n14706) );
  NANDN U15031 ( .A(n14814), .B(n14815), .Z(n14813) );
  NANDN U15032 ( .A(n14816), .B(n14817), .Z(n14815) );
  NANDN U15033 ( .A(n14817), .B(n14816), .Z(n14812) );
  ANDN U15034 ( .B(B[184]), .A(n31), .Z(n14708) );
  XNOR U15035 ( .A(n14716), .B(n14818), .Z(n14709) );
  XNOR U15036 ( .A(n14715), .B(n14713), .Z(n14818) );
  AND U15037 ( .A(n14819), .B(n14820), .Z(n14713) );
  NANDN U15038 ( .A(n14821), .B(n14822), .Z(n14820) );
  OR U15039 ( .A(n14823), .B(n14824), .Z(n14822) );
  NAND U15040 ( .A(n14824), .B(n14823), .Z(n14819) );
  ANDN U15041 ( .B(B[185]), .A(n32), .Z(n14715) );
  XNOR U15042 ( .A(n14723), .B(n14825), .Z(n14716) );
  XNOR U15043 ( .A(n14722), .B(n14720), .Z(n14825) );
  AND U15044 ( .A(n14826), .B(n14827), .Z(n14720) );
  NANDN U15045 ( .A(n14828), .B(n14829), .Z(n14827) );
  NANDN U15046 ( .A(n14830), .B(n14831), .Z(n14829) );
  NANDN U15047 ( .A(n14831), .B(n14830), .Z(n14826) );
  ANDN U15048 ( .B(B[186]), .A(n33), .Z(n14722) );
  XNOR U15049 ( .A(n14730), .B(n14832), .Z(n14723) );
  XNOR U15050 ( .A(n14729), .B(n14727), .Z(n14832) );
  AND U15051 ( .A(n14833), .B(n14834), .Z(n14727) );
  NANDN U15052 ( .A(n14835), .B(n14836), .Z(n14834) );
  OR U15053 ( .A(n14837), .B(n14838), .Z(n14836) );
  NAND U15054 ( .A(n14838), .B(n14837), .Z(n14833) );
  ANDN U15055 ( .B(B[187]), .A(n34), .Z(n14729) );
  XNOR U15056 ( .A(n14737), .B(n14839), .Z(n14730) );
  XNOR U15057 ( .A(n14736), .B(n14734), .Z(n14839) );
  AND U15058 ( .A(n14840), .B(n14841), .Z(n14734) );
  NANDN U15059 ( .A(n14842), .B(n14843), .Z(n14841) );
  NANDN U15060 ( .A(n14844), .B(n14845), .Z(n14843) );
  NANDN U15061 ( .A(n14845), .B(n14844), .Z(n14840) );
  ANDN U15062 ( .B(B[188]), .A(n35), .Z(n14736) );
  XNOR U15063 ( .A(n14744), .B(n14846), .Z(n14737) );
  XNOR U15064 ( .A(n14743), .B(n14741), .Z(n14846) );
  AND U15065 ( .A(n14847), .B(n14848), .Z(n14741) );
  NANDN U15066 ( .A(n14849), .B(n14850), .Z(n14848) );
  OR U15067 ( .A(n14851), .B(n14852), .Z(n14850) );
  NAND U15068 ( .A(n14852), .B(n14851), .Z(n14847) );
  ANDN U15069 ( .B(B[189]), .A(n36), .Z(n14743) );
  XNOR U15070 ( .A(n14751), .B(n14853), .Z(n14744) );
  XNOR U15071 ( .A(n14750), .B(n14748), .Z(n14853) );
  AND U15072 ( .A(n14854), .B(n14855), .Z(n14748) );
  NANDN U15073 ( .A(n14856), .B(n14857), .Z(n14855) );
  NANDN U15074 ( .A(n14858), .B(n14859), .Z(n14857) );
  NANDN U15075 ( .A(n14859), .B(n14858), .Z(n14854) );
  ANDN U15076 ( .B(B[190]), .A(n37), .Z(n14750) );
  XNOR U15077 ( .A(n14758), .B(n14860), .Z(n14751) );
  XNOR U15078 ( .A(n14757), .B(n14755), .Z(n14860) );
  AND U15079 ( .A(n14861), .B(n14862), .Z(n14755) );
  NANDN U15080 ( .A(n14863), .B(n14864), .Z(n14862) );
  OR U15081 ( .A(n14865), .B(n14866), .Z(n14864) );
  NAND U15082 ( .A(n14866), .B(n14865), .Z(n14861) );
  ANDN U15083 ( .B(B[191]), .A(n38), .Z(n14757) );
  XNOR U15084 ( .A(n14765), .B(n14867), .Z(n14758) );
  XNOR U15085 ( .A(n14764), .B(n14762), .Z(n14867) );
  AND U15086 ( .A(n14868), .B(n14869), .Z(n14762) );
  NANDN U15087 ( .A(n14870), .B(n14871), .Z(n14869) );
  NANDN U15088 ( .A(n14872), .B(n14873), .Z(n14871) );
  NANDN U15089 ( .A(n14873), .B(n14872), .Z(n14868) );
  ANDN U15090 ( .B(B[192]), .A(n39), .Z(n14764) );
  XNOR U15091 ( .A(n14772), .B(n14874), .Z(n14765) );
  XNOR U15092 ( .A(n14771), .B(n14769), .Z(n14874) );
  AND U15093 ( .A(n14875), .B(n14876), .Z(n14769) );
  NANDN U15094 ( .A(n14877), .B(n14878), .Z(n14876) );
  OR U15095 ( .A(n14879), .B(n14880), .Z(n14878) );
  NAND U15096 ( .A(n14880), .B(n14879), .Z(n14875) );
  ANDN U15097 ( .B(B[193]), .A(n40), .Z(n14771) );
  XNOR U15098 ( .A(n14779), .B(n14881), .Z(n14772) );
  XNOR U15099 ( .A(n14778), .B(n14776), .Z(n14881) );
  AND U15100 ( .A(n14882), .B(n14883), .Z(n14776) );
  NANDN U15101 ( .A(n14884), .B(n14885), .Z(n14883) );
  NAND U15102 ( .A(n14886), .B(n14887), .Z(n14885) );
  ANDN U15103 ( .B(B[194]), .A(n41), .Z(n14778) );
  XOR U15104 ( .A(n14785), .B(n14888), .Z(n14779) );
  XNOR U15105 ( .A(n14783), .B(n14786), .Z(n14888) );
  NAND U15106 ( .A(A[2]), .B(B[195]), .Z(n14786) );
  NANDN U15107 ( .A(n14889), .B(n14890), .Z(n14783) );
  AND U15108 ( .A(A[0]), .B(B[196]), .Z(n14890) );
  XNOR U15109 ( .A(n14788), .B(n14891), .Z(n14785) );
  NAND U15110 ( .A(A[0]), .B(B[197]), .Z(n14891) );
  NAND U15111 ( .A(B[196]), .B(A[1]), .Z(n14788) );
  NAND U15112 ( .A(n14892), .B(n14893), .Z(n353) );
  NANDN U15113 ( .A(n14894), .B(n14895), .Z(n14893) );
  OR U15114 ( .A(n14896), .B(n14897), .Z(n14895) );
  NAND U15115 ( .A(n14897), .B(n14896), .Z(n14892) );
  XOR U15116 ( .A(n355), .B(n354), .Z(\A1[194] ) );
  XOR U15117 ( .A(n14897), .B(n14898), .Z(n354) );
  XNOR U15118 ( .A(n14896), .B(n14894), .Z(n14898) );
  AND U15119 ( .A(n14899), .B(n14900), .Z(n14894) );
  NANDN U15120 ( .A(n14901), .B(n14902), .Z(n14900) );
  NANDN U15121 ( .A(n14903), .B(n14904), .Z(n14902) );
  NANDN U15122 ( .A(n14904), .B(n14903), .Z(n14899) );
  ANDN U15123 ( .B(B[181]), .A(n29), .Z(n14896) );
  XNOR U15124 ( .A(n14803), .B(n14905), .Z(n14897) );
  XNOR U15125 ( .A(n14802), .B(n14800), .Z(n14905) );
  AND U15126 ( .A(n14906), .B(n14907), .Z(n14800) );
  NANDN U15127 ( .A(n14908), .B(n14909), .Z(n14907) );
  OR U15128 ( .A(n14910), .B(n14911), .Z(n14909) );
  NAND U15129 ( .A(n14911), .B(n14910), .Z(n14906) );
  ANDN U15130 ( .B(B[182]), .A(n30), .Z(n14802) );
  XNOR U15131 ( .A(n14810), .B(n14912), .Z(n14803) );
  XNOR U15132 ( .A(n14809), .B(n14807), .Z(n14912) );
  AND U15133 ( .A(n14913), .B(n14914), .Z(n14807) );
  NANDN U15134 ( .A(n14915), .B(n14916), .Z(n14914) );
  NANDN U15135 ( .A(n14917), .B(n14918), .Z(n14916) );
  NANDN U15136 ( .A(n14918), .B(n14917), .Z(n14913) );
  ANDN U15137 ( .B(B[183]), .A(n31), .Z(n14809) );
  XNOR U15138 ( .A(n14817), .B(n14919), .Z(n14810) );
  XNOR U15139 ( .A(n14816), .B(n14814), .Z(n14919) );
  AND U15140 ( .A(n14920), .B(n14921), .Z(n14814) );
  NANDN U15141 ( .A(n14922), .B(n14923), .Z(n14921) );
  OR U15142 ( .A(n14924), .B(n14925), .Z(n14923) );
  NAND U15143 ( .A(n14925), .B(n14924), .Z(n14920) );
  ANDN U15144 ( .B(B[184]), .A(n32), .Z(n14816) );
  XNOR U15145 ( .A(n14824), .B(n14926), .Z(n14817) );
  XNOR U15146 ( .A(n14823), .B(n14821), .Z(n14926) );
  AND U15147 ( .A(n14927), .B(n14928), .Z(n14821) );
  NANDN U15148 ( .A(n14929), .B(n14930), .Z(n14928) );
  NANDN U15149 ( .A(n14931), .B(n14932), .Z(n14930) );
  NANDN U15150 ( .A(n14932), .B(n14931), .Z(n14927) );
  ANDN U15151 ( .B(B[185]), .A(n33), .Z(n14823) );
  XNOR U15152 ( .A(n14831), .B(n14933), .Z(n14824) );
  XNOR U15153 ( .A(n14830), .B(n14828), .Z(n14933) );
  AND U15154 ( .A(n14934), .B(n14935), .Z(n14828) );
  NANDN U15155 ( .A(n14936), .B(n14937), .Z(n14935) );
  OR U15156 ( .A(n14938), .B(n14939), .Z(n14937) );
  NAND U15157 ( .A(n14939), .B(n14938), .Z(n14934) );
  ANDN U15158 ( .B(B[186]), .A(n34), .Z(n14830) );
  XNOR U15159 ( .A(n14838), .B(n14940), .Z(n14831) );
  XNOR U15160 ( .A(n14837), .B(n14835), .Z(n14940) );
  AND U15161 ( .A(n14941), .B(n14942), .Z(n14835) );
  NANDN U15162 ( .A(n14943), .B(n14944), .Z(n14942) );
  NANDN U15163 ( .A(n14945), .B(n14946), .Z(n14944) );
  NANDN U15164 ( .A(n14946), .B(n14945), .Z(n14941) );
  ANDN U15165 ( .B(B[187]), .A(n35), .Z(n14837) );
  XNOR U15166 ( .A(n14845), .B(n14947), .Z(n14838) );
  XNOR U15167 ( .A(n14844), .B(n14842), .Z(n14947) );
  AND U15168 ( .A(n14948), .B(n14949), .Z(n14842) );
  NANDN U15169 ( .A(n14950), .B(n14951), .Z(n14949) );
  OR U15170 ( .A(n14952), .B(n14953), .Z(n14951) );
  NAND U15171 ( .A(n14953), .B(n14952), .Z(n14948) );
  ANDN U15172 ( .B(B[188]), .A(n36), .Z(n14844) );
  XNOR U15173 ( .A(n14852), .B(n14954), .Z(n14845) );
  XNOR U15174 ( .A(n14851), .B(n14849), .Z(n14954) );
  AND U15175 ( .A(n14955), .B(n14956), .Z(n14849) );
  NANDN U15176 ( .A(n14957), .B(n14958), .Z(n14956) );
  NANDN U15177 ( .A(n14959), .B(n14960), .Z(n14958) );
  NANDN U15178 ( .A(n14960), .B(n14959), .Z(n14955) );
  ANDN U15179 ( .B(B[189]), .A(n37), .Z(n14851) );
  XNOR U15180 ( .A(n14859), .B(n14961), .Z(n14852) );
  XNOR U15181 ( .A(n14858), .B(n14856), .Z(n14961) );
  AND U15182 ( .A(n14962), .B(n14963), .Z(n14856) );
  NANDN U15183 ( .A(n14964), .B(n14965), .Z(n14963) );
  OR U15184 ( .A(n14966), .B(n14967), .Z(n14965) );
  NAND U15185 ( .A(n14967), .B(n14966), .Z(n14962) );
  ANDN U15186 ( .B(B[190]), .A(n38), .Z(n14858) );
  XNOR U15187 ( .A(n14866), .B(n14968), .Z(n14859) );
  XNOR U15188 ( .A(n14865), .B(n14863), .Z(n14968) );
  AND U15189 ( .A(n14969), .B(n14970), .Z(n14863) );
  NANDN U15190 ( .A(n14971), .B(n14972), .Z(n14970) );
  NANDN U15191 ( .A(n14973), .B(n14974), .Z(n14972) );
  NANDN U15192 ( .A(n14974), .B(n14973), .Z(n14969) );
  ANDN U15193 ( .B(B[191]), .A(n39), .Z(n14865) );
  XNOR U15194 ( .A(n14873), .B(n14975), .Z(n14866) );
  XNOR U15195 ( .A(n14872), .B(n14870), .Z(n14975) );
  AND U15196 ( .A(n14976), .B(n14977), .Z(n14870) );
  NANDN U15197 ( .A(n14978), .B(n14979), .Z(n14977) );
  OR U15198 ( .A(n14980), .B(n14981), .Z(n14979) );
  NAND U15199 ( .A(n14981), .B(n14980), .Z(n14976) );
  ANDN U15200 ( .B(B[192]), .A(n40), .Z(n14872) );
  XNOR U15201 ( .A(n14880), .B(n14982), .Z(n14873) );
  XNOR U15202 ( .A(n14879), .B(n14877), .Z(n14982) );
  AND U15203 ( .A(n14983), .B(n14984), .Z(n14877) );
  NANDN U15204 ( .A(n14985), .B(n14986), .Z(n14984) );
  NAND U15205 ( .A(n14987), .B(n14988), .Z(n14986) );
  ANDN U15206 ( .B(B[193]), .A(n41), .Z(n14879) );
  XOR U15207 ( .A(n14886), .B(n14989), .Z(n14880) );
  XNOR U15208 ( .A(n14884), .B(n14887), .Z(n14989) );
  NAND U15209 ( .A(A[2]), .B(B[194]), .Z(n14887) );
  NANDN U15210 ( .A(n14990), .B(n14991), .Z(n14884) );
  AND U15211 ( .A(A[0]), .B(B[195]), .Z(n14991) );
  XNOR U15212 ( .A(n14889), .B(n14992), .Z(n14886) );
  NAND U15213 ( .A(A[0]), .B(B[196]), .Z(n14992) );
  NAND U15214 ( .A(B[195]), .B(A[1]), .Z(n14889) );
  NAND U15215 ( .A(n14993), .B(n14994), .Z(n355) );
  NANDN U15216 ( .A(n14995), .B(n14996), .Z(n14994) );
  OR U15217 ( .A(n14997), .B(n14998), .Z(n14996) );
  NAND U15218 ( .A(n14998), .B(n14997), .Z(n14993) );
  XOR U15219 ( .A(n357), .B(n356), .Z(\A1[193] ) );
  XOR U15220 ( .A(n14998), .B(n14999), .Z(n356) );
  XNOR U15221 ( .A(n14997), .B(n14995), .Z(n14999) );
  AND U15222 ( .A(n15000), .B(n15001), .Z(n14995) );
  NANDN U15223 ( .A(n15002), .B(n15003), .Z(n15001) );
  NANDN U15224 ( .A(n15004), .B(n15005), .Z(n15003) );
  NANDN U15225 ( .A(n15005), .B(n15004), .Z(n15000) );
  ANDN U15226 ( .B(B[180]), .A(n29), .Z(n14997) );
  XNOR U15227 ( .A(n14904), .B(n15006), .Z(n14998) );
  XNOR U15228 ( .A(n14903), .B(n14901), .Z(n15006) );
  AND U15229 ( .A(n15007), .B(n15008), .Z(n14901) );
  NANDN U15230 ( .A(n15009), .B(n15010), .Z(n15008) );
  OR U15231 ( .A(n15011), .B(n15012), .Z(n15010) );
  NAND U15232 ( .A(n15012), .B(n15011), .Z(n15007) );
  ANDN U15233 ( .B(B[181]), .A(n30), .Z(n14903) );
  XNOR U15234 ( .A(n14911), .B(n15013), .Z(n14904) );
  XNOR U15235 ( .A(n14910), .B(n14908), .Z(n15013) );
  AND U15236 ( .A(n15014), .B(n15015), .Z(n14908) );
  NANDN U15237 ( .A(n15016), .B(n15017), .Z(n15015) );
  NANDN U15238 ( .A(n15018), .B(n15019), .Z(n15017) );
  NANDN U15239 ( .A(n15019), .B(n15018), .Z(n15014) );
  ANDN U15240 ( .B(B[182]), .A(n31), .Z(n14910) );
  XNOR U15241 ( .A(n14918), .B(n15020), .Z(n14911) );
  XNOR U15242 ( .A(n14917), .B(n14915), .Z(n15020) );
  AND U15243 ( .A(n15021), .B(n15022), .Z(n14915) );
  NANDN U15244 ( .A(n15023), .B(n15024), .Z(n15022) );
  OR U15245 ( .A(n15025), .B(n15026), .Z(n15024) );
  NAND U15246 ( .A(n15026), .B(n15025), .Z(n15021) );
  ANDN U15247 ( .B(B[183]), .A(n32), .Z(n14917) );
  XNOR U15248 ( .A(n14925), .B(n15027), .Z(n14918) );
  XNOR U15249 ( .A(n14924), .B(n14922), .Z(n15027) );
  AND U15250 ( .A(n15028), .B(n15029), .Z(n14922) );
  NANDN U15251 ( .A(n15030), .B(n15031), .Z(n15029) );
  NANDN U15252 ( .A(n15032), .B(n15033), .Z(n15031) );
  NANDN U15253 ( .A(n15033), .B(n15032), .Z(n15028) );
  ANDN U15254 ( .B(B[184]), .A(n33), .Z(n14924) );
  XNOR U15255 ( .A(n14932), .B(n15034), .Z(n14925) );
  XNOR U15256 ( .A(n14931), .B(n14929), .Z(n15034) );
  AND U15257 ( .A(n15035), .B(n15036), .Z(n14929) );
  NANDN U15258 ( .A(n15037), .B(n15038), .Z(n15036) );
  OR U15259 ( .A(n15039), .B(n15040), .Z(n15038) );
  NAND U15260 ( .A(n15040), .B(n15039), .Z(n15035) );
  ANDN U15261 ( .B(B[185]), .A(n34), .Z(n14931) );
  XNOR U15262 ( .A(n14939), .B(n15041), .Z(n14932) );
  XNOR U15263 ( .A(n14938), .B(n14936), .Z(n15041) );
  AND U15264 ( .A(n15042), .B(n15043), .Z(n14936) );
  NANDN U15265 ( .A(n15044), .B(n15045), .Z(n15043) );
  NANDN U15266 ( .A(n15046), .B(n15047), .Z(n15045) );
  NANDN U15267 ( .A(n15047), .B(n15046), .Z(n15042) );
  ANDN U15268 ( .B(B[186]), .A(n35), .Z(n14938) );
  XNOR U15269 ( .A(n14946), .B(n15048), .Z(n14939) );
  XNOR U15270 ( .A(n14945), .B(n14943), .Z(n15048) );
  AND U15271 ( .A(n15049), .B(n15050), .Z(n14943) );
  NANDN U15272 ( .A(n15051), .B(n15052), .Z(n15050) );
  OR U15273 ( .A(n15053), .B(n15054), .Z(n15052) );
  NAND U15274 ( .A(n15054), .B(n15053), .Z(n15049) );
  ANDN U15275 ( .B(B[187]), .A(n36), .Z(n14945) );
  XNOR U15276 ( .A(n14953), .B(n15055), .Z(n14946) );
  XNOR U15277 ( .A(n14952), .B(n14950), .Z(n15055) );
  AND U15278 ( .A(n15056), .B(n15057), .Z(n14950) );
  NANDN U15279 ( .A(n15058), .B(n15059), .Z(n15057) );
  NANDN U15280 ( .A(n15060), .B(n15061), .Z(n15059) );
  NANDN U15281 ( .A(n15061), .B(n15060), .Z(n15056) );
  ANDN U15282 ( .B(B[188]), .A(n37), .Z(n14952) );
  XNOR U15283 ( .A(n14960), .B(n15062), .Z(n14953) );
  XNOR U15284 ( .A(n14959), .B(n14957), .Z(n15062) );
  AND U15285 ( .A(n15063), .B(n15064), .Z(n14957) );
  NANDN U15286 ( .A(n15065), .B(n15066), .Z(n15064) );
  OR U15287 ( .A(n15067), .B(n15068), .Z(n15066) );
  NAND U15288 ( .A(n15068), .B(n15067), .Z(n15063) );
  ANDN U15289 ( .B(B[189]), .A(n38), .Z(n14959) );
  XNOR U15290 ( .A(n14967), .B(n15069), .Z(n14960) );
  XNOR U15291 ( .A(n14966), .B(n14964), .Z(n15069) );
  AND U15292 ( .A(n15070), .B(n15071), .Z(n14964) );
  NANDN U15293 ( .A(n15072), .B(n15073), .Z(n15071) );
  NANDN U15294 ( .A(n15074), .B(n15075), .Z(n15073) );
  NANDN U15295 ( .A(n15075), .B(n15074), .Z(n15070) );
  ANDN U15296 ( .B(B[190]), .A(n39), .Z(n14966) );
  XNOR U15297 ( .A(n14974), .B(n15076), .Z(n14967) );
  XNOR U15298 ( .A(n14973), .B(n14971), .Z(n15076) );
  AND U15299 ( .A(n15077), .B(n15078), .Z(n14971) );
  NANDN U15300 ( .A(n15079), .B(n15080), .Z(n15078) );
  OR U15301 ( .A(n15081), .B(n15082), .Z(n15080) );
  NAND U15302 ( .A(n15082), .B(n15081), .Z(n15077) );
  ANDN U15303 ( .B(B[191]), .A(n40), .Z(n14973) );
  XNOR U15304 ( .A(n14981), .B(n15083), .Z(n14974) );
  XNOR U15305 ( .A(n14980), .B(n14978), .Z(n15083) );
  AND U15306 ( .A(n15084), .B(n15085), .Z(n14978) );
  NANDN U15307 ( .A(n15086), .B(n15087), .Z(n15085) );
  NAND U15308 ( .A(n15088), .B(n15089), .Z(n15087) );
  ANDN U15309 ( .B(B[192]), .A(n41), .Z(n14980) );
  XOR U15310 ( .A(n14987), .B(n15090), .Z(n14981) );
  XNOR U15311 ( .A(n14985), .B(n14988), .Z(n15090) );
  NAND U15312 ( .A(A[2]), .B(B[193]), .Z(n14988) );
  NANDN U15313 ( .A(n15091), .B(n15092), .Z(n14985) );
  AND U15314 ( .A(A[0]), .B(B[194]), .Z(n15092) );
  XNOR U15315 ( .A(n14990), .B(n15093), .Z(n14987) );
  NAND U15316 ( .A(A[0]), .B(B[195]), .Z(n15093) );
  NAND U15317 ( .A(B[194]), .B(A[1]), .Z(n14990) );
  NAND U15318 ( .A(n15094), .B(n15095), .Z(n357) );
  NANDN U15319 ( .A(n15096), .B(n15097), .Z(n15095) );
  OR U15320 ( .A(n15098), .B(n15099), .Z(n15097) );
  NAND U15321 ( .A(n15099), .B(n15098), .Z(n15094) );
  XOR U15322 ( .A(n359), .B(n358), .Z(\A1[192] ) );
  XOR U15323 ( .A(n15099), .B(n15100), .Z(n358) );
  XNOR U15324 ( .A(n15098), .B(n15096), .Z(n15100) );
  AND U15325 ( .A(n15101), .B(n15102), .Z(n15096) );
  NANDN U15326 ( .A(n15103), .B(n15104), .Z(n15102) );
  NANDN U15327 ( .A(n15105), .B(n15106), .Z(n15104) );
  NANDN U15328 ( .A(n15106), .B(n15105), .Z(n15101) );
  ANDN U15329 ( .B(B[179]), .A(n29), .Z(n15098) );
  XNOR U15330 ( .A(n15005), .B(n15107), .Z(n15099) );
  XNOR U15331 ( .A(n15004), .B(n15002), .Z(n15107) );
  AND U15332 ( .A(n15108), .B(n15109), .Z(n15002) );
  NANDN U15333 ( .A(n15110), .B(n15111), .Z(n15109) );
  OR U15334 ( .A(n15112), .B(n15113), .Z(n15111) );
  NAND U15335 ( .A(n15113), .B(n15112), .Z(n15108) );
  ANDN U15336 ( .B(B[180]), .A(n30), .Z(n15004) );
  XNOR U15337 ( .A(n15012), .B(n15114), .Z(n15005) );
  XNOR U15338 ( .A(n15011), .B(n15009), .Z(n15114) );
  AND U15339 ( .A(n15115), .B(n15116), .Z(n15009) );
  NANDN U15340 ( .A(n15117), .B(n15118), .Z(n15116) );
  NANDN U15341 ( .A(n15119), .B(n15120), .Z(n15118) );
  NANDN U15342 ( .A(n15120), .B(n15119), .Z(n15115) );
  ANDN U15343 ( .B(B[181]), .A(n31), .Z(n15011) );
  XNOR U15344 ( .A(n15019), .B(n15121), .Z(n15012) );
  XNOR U15345 ( .A(n15018), .B(n15016), .Z(n15121) );
  AND U15346 ( .A(n15122), .B(n15123), .Z(n15016) );
  NANDN U15347 ( .A(n15124), .B(n15125), .Z(n15123) );
  OR U15348 ( .A(n15126), .B(n15127), .Z(n15125) );
  NAND U15349 ( .A(n15127), .B(n15126), .Z(n15122) );
  ANDN U15350 ( .B(B[182]), .A(n32), .Z(n15018) );
  XNOR U15351 ( .A(n15026), .B(n15128), .Z(n15019) );
  XNOR U15352 ( .A(n15025), .B(n15023), .Z(n15128) );
  AND U15353 ( .A(n15129), .B(n15130), .Z(n15023) );
  NANDN U15354 ( .A(n15131), .B(n15132), .Z(n15130) );
  NANDN U15355 ( .A(n15133), .B(n15134), .Z(n15132) );
  NANDN U15356 ( .A(n15134), .B(n15133), .Z(n15129) );
  ANDN U15357 ( .B(B[183]), .A(n33), .Z(n15025) );
  XNOR U15358 ( .A(n15033), .B(n15135), .Z(n15026) );
  XNOR U15359 ( .A(n15032), .B(n15030), .Z(n15135) );
  AND U15360 ( .A(n15136), .B(n15137), .Z(n15030) );
  NANDN U15361 ( .A(n15138), .B(n15139), .Z(n15137) );
  OR U15362 ( .A(n15140), .B(n15141), .Z(n15139) );
  NAND U15363 ( .A(n15141), .B(n15140), .Z(n15136) );
  ANDN U15364 ( .B(B[184]), .A(n34), .Z(n15032) );
  XNOR U15365 ( .A(n15040), .B(n15142), .Z(n15033) );
  XNOR U15366 ( .A(n15039), .B(n15037), .Z(n15142) );
  AND U15367 ( .A(n15143), .B(n15144), .Z(n15037) );
  NANDN U15368 ( .A(n15145), .B(n15146), .Z(n15144) );
  NANDN U15369 ( .A(n15147), .B(n15148), .Z(n15146) );
  NANDN U15370 ( .A(n15148), .B(n15147), .Z(n15143) );
  ANDN U15371 ( .B(B[185]), .A(n35), .Z(n15039) );
  XNOR U15372 ( .A(n15047), .B(n15149), .Z(n15040) );
  XNOR U15373 ( .A(n15046), .B(n15044), .Z(n15149) );
  AND U15374 ( .A(n15150), .B(n15151), .Z(n15044) );
  NANDN U15375 ( .A(n15152), .B(n15153), .Z(n15151) );
  OR U15376 ( .A(n15154), .B(n15155), .Z(n15153) );
  NAND U15377 ( .A(n15155), .B(n15154), .Z(n15150) );
  ANDN U15378 ( .B(B[186]), .A(n36), .Z(n15046) );
  XNOR U15379 ( .A(n15054), .B(n15156), .Z(n15047) );
  XNOR U15380 ( .A(n15053), .B(n15051), .Z(n15156) );
  AND U15381 ( .A(n15157), .B(n15158), .Z(n15051) );
  NANDN U15382 ( .A(n15159), .B(n15160), .Z(n15158) );
  NANDN U15383 ( .A(n15161), .B(n15162), .Z(n15160) );
  NANDN U15384 ( .A(n15162), .B(n15161), .Z(n15157) );
  ANDN U15385 ( .B(B[187]), .A(n37), .Z(n15053) );
  XNOR U15386 ( .A(n15061), .B(n15163), .Z(n15054) );
  XNOR U15387 ( .A(n15060), .B(n15058), .Z(n15163) );
  AND U15388 ( .A(n15164), .B(n15165), .Z(n15058) );
  NANDN U15389 ( .A(n15166), .B(n15167), .Z(n15165) );
  OR U15390 ( .A(n15168), .B(n15169), .Z(n15167) );
  NAND U15391 ( .A(n15169), .B(n15168), .Z(n15164) );
  ANDN U15392 ( .B(B[188]), .A(n38), .Z(n15060) );
  XNOR U15393 ( .A(n15068), .B(n15170), .Z(n15061) );
  XNOR U15394 ( .A(n15067), .B(n15065), .Z(n15170) );
  AND U15395 ( .A(n15171), .B(n15172), .Z(n15065) );
  NANDN U15396 ( .A(n15173), .B(n15174), .Z(n15172) );
  NANDN U15397 ( .A(n15175), .B(n15176), .Z(n15174) );
  NANDN U15398 ( .A(n15176), .B(n15175), .Z(n15171) );
  ANDN U15399 ( .B(B[189]), .A(n39), .Z(n15067) );
  XNOR U15400 ( .A(n15075), .B(n15177), .Z(n15068) );
  XNOR U15401 ( .A(n15074), .B(n15072), .Z(n15177) );
  AND U15402 ( .A(n15178), .B(n15179), .Z(n15072) );
  NANDN U15403 ( .A(n15180), .B(n15181), .Z(n15179) );
  OR U15404 ( .A(n15182), .B(n15183), .Z(n15181) );
  NAND U15405 ( .A(n15183), .B(n15182), .Z(n15178) );
  ANDN U15406 ( .B(B[190]), .A(n40), .Z(n15074) );
  XNOR U15407 ( .A(n15082), .B(n15184), .Z(n15075) );
  XNOR U15408 ( .A(n15081), .B(n15079), .Z(n15184) );
  AND U15409 ( .A(n15185), .B(n15186), .Z(n15079) );
  NANDN U15410 ( .A(n15187), .B(n15188), .Z(n15186) );
  NAND U15411 ( .A(n15189), .B(n15190), .Z(n15188) );
  ANDN U15412 ( .B(B[191]), .A(n41), .Z(n15081) );
  XOR U15413 ( .A(n15088), .B(n15191), .Z(n15082) );
  XNOR U15414 ( .A(n15086), .B(n15089), .Z(n15191) );
  NAND U15415 ( .A(A[2]), .B(B[192]), .Z(n15089) );
  NANDN U15416 ( .A(n15192), .B(n15193), .Z(n15086) );
  AND U15417 ( .A(A[0]), .B(B[193]), .Z(n15193) );
  XNOR U15418 ( .A(n15091), .B(n15194), .Z(n15088) );
  NAND U15419 ( .A(A[0]), .B(B[194]), .Z(n15194) );
  NAND U15420 ( .A(B[193]), .B(A[1]), .Z(n15091) );
  NAND U15421 ( .A(n15195), .B(n15196), .Z(n359) );
  NANDN U15422 ( .A(n15197), .B(n15198), .Z(n15196) );
  OR U15423 ( .A(n15199), .B(n15200), .Z(n15198) );
  NAND U15424 ( .A(n15200), .B(n15199), .Z(n15195) );
  XOR U15425 ( .A(n361), .B(n360), .Z(\A1[191] ) );
  XOR U15426 ( .A(n15200), .B(n15201), .Z(n360) );
  XNOR U15427 ( .A(n15199), .B(n15197), .Z(n15201) );
  AND U15428 ( .A(n15202), .B(n15203), .Z(n15197) );
  NANDN U15429 ( .A(n15204), .B(n15205), .Z(n15203) );
  NANDN U15430 ( .A(n15206), .B(n15207), .Z(n15205) );
  NANDN U15431 ( .A(n15207), .B(n15206), .Z(n15202) );
  ANDN U15432 ( .B(B[178]), .A(n29), .Z(n15199) );
  XNOR U15433 ( .A(n15106), .B(n15208), .Z(n15200) );
  XNOR U15434 ( .A(n15105), .B(n15103), .Z(n15208) );
  AND U15435 ( .A(n15209), .B(n15210), .Z(n15103) );
  NANDN U15436 ( .A(n15211), .B(n15212), .Z(n15210) );
  OR U15437 ( .A(n15213), .B(n15214), .Z(n15212) );
  NAND U15438 ( .A(n15214), .B(n15213), .Z(n15209) );
  ANDN U15439 ( .B(B[179]), .A(n30), .Z(n15105) );
  XNOR U15440 ( .A(n15113), .B(n15215), .Z(n15106) );
  XNOR U15441 ( .A(n15112), .B(n15110), .Z(n15215) );
  AND U15442 ( .A(n15216), .B(n15217), .Z(n15110) );
  NANDN U15443 ( .A(n15218), .B(n15219), .Z(n15217) );
  NANDN U15444 ( .A(n15220), .B(n15221), .Z(n15219) );
  NANDN U15445 ( .A(n15221), .B(n15220), .Z(n15216) );
  ANDN U15446 ( .B(B[180]), .A(n31), .Z(n15112) );
  XNOR U15447 ( .A(n15120), .B(n15222), .Z(n15113) );
  XNOR U15448 ( .A(n15119), .B(n15117), .Z(n15222) );
  AND U15449 ( .A(n15223), .B(n15224), .Z(n15117) );
  NANDN U15450 ( .A(n15225), .B(n15226), .Z(n15224) );
  OR U15451 ( .A(n15227), .B(n15228), .Z(n15226) );
  NAND U15452 ( .A(n15228), .B(n15227), .Z(n15223) );
  ANDN U15453 ( .B(B[181]), .A(n32), .Z(n15119) );
  XNOR U15454 ( .A(n15127), .B(n15229), .Z(n15120) );
  XNOR U15455 ( .A(n15126), .B(n15124), .Z(n15229) );
  AND U15456 ( .A(n15230), .B(n15231), .Z(n15124) );
  NANDN U15457 ( .A(n15232), .B(n15233), .Z(n15231) );
  NANDN U15458 ( .A(n15234), .B(n15235), .Z(n15233) );
  NANDN U15459 ( .A(n15235), .B(n15234), .Z(n15230) );
  ANDN U15460 ( .B(B[182]), .A(n33), .Z(n15126) );
  XNOR U15461 ( .A(n15134), .B(n15236), .Z(n15127) );
  XNOR U15462 ( .A(n15133), .B(n15131), .Z(n15236) );
  AND U15463 ( .A(n15237), .B(n15238), .Z(n15131) );
  NANDN U15464 ( .A(n15239), .B(n15240), .Z(n15238) );
  OR U15465 ( .A(n15241), .B(n15242), .Z(n15240) );
  NAND U15466 ( .A(n15242), .B(n15241), .Z(n15237) );
  ANDN U15467 ( .B(B[183]), .A(n34), .Z(n15133) );
  XNOR U15468 ( .A(n15141), .B(n15243), .Z(n15134) );
  XNOR U15469 ( .A(n15140), .B(n15138), .Z(n15243) );
  AND U15470 ( .A(n15244), .B(n15245), .Z(n15138) );
  NANDN U15471 ( .A(n15246), .B(n15247), .Z(n15245) );
  NANDN U15472 ( .A(n15248), .B(n15249), .Z(n15247) );
  NANDN U15473 ( .A(n15249), .B(n15248), .Z(n15244) );
  ANDN U15474 ( .B(B[184]), .A(n35), .Z(n15140) );
  XNOR U15475 ( .A(n15148), .B(n15250), .Z(n15141) );
  XNOR U15476 ( .A(n15147), .B(n15145), .Z(n15250) );
  AND U15477 ( .A(n15251), .B(n15252), .Z(n15145) );
  NANDN U15478 ( .A(n15253), .B(n15254), .Z(n15252) );
  OR U15479 ( .A(n15255), .B(n15256), .Z(n15254) );
  NAND U15480 ( .A(n15256), .B(n15255), .Z(n15251) );
  ANDN U15481 ( .B(B[185]), .A(n36), .Z(n15147) );
  XNOR U15482 ( .A(n15155), .B(n15257), .Z(n15148) );
  XNOR U15483 ( .A(n15154), .B(n15152), .Z(n15257) );
  AND U15484 ( .A(n15258), .B(n15259), .Z(n15152) );
  NANDN U15485 ( .A(n15260), .B(n15261), .Z(n15259) );
  NANDN U15486 ( .A(n15262), .B(n15263), .Z(n15261) );
  NANDN U15487 ( .A(n15263), .B(n15262), .Z(n15258) );
  ANDN U15488 ( .B(B[186]), .A(n37), .Z(n15154) );
  XNOR U15489 ( .A(n15162), .B(n15264), .Z(n15155) );
  XNOR U15490 ( .A(n15161), .B(n15159), .Z(n15264) );
  AND U15491 ( .A(n15265), .B(n15266), .Z(n15159) );
  NANDN U15492 ( .A(n15267), .B(n15268), .Z(n15266) );
  OR U15493 ( .A(n15269), .B(n15270), .Z(n15268) );
  NAND U15494 ( .A(n15270), .B(n15269), .Z(n15265) );
  ANDN U15495 ( .B(B[187]), .A(n38), .Z(n15161) );
  XNOR U15496 ( .A(n15169), .B(n15271), .Z(n15162) );
  XNOR U15497 ( .A(n15168), .B(n15166), .Z(n15271) );
  AND U15498 ( .A(n15272), .B(n15273), .Z(n15166) );
  NANDN U15499 ( .A(n15274), .B(n15275), .Z(n15273) );
  NANDN U15500 ( .A(n15276), .B(n15277), .Z(n15275) );
  NANDN U15501 ( .A(n15277), .B(n15276), .Z(n15272) );
  ANDN U15502 ( .B(B[188]), .A(n39), .Z(n15168) );
  XNOR U15503 ( .A(n15176), .B(n15278), .Z(n15169) );
  XNOR U15504 ( .A(n15175), .B(n15173), .Z(n15278) );
  AND U15505 ( .A(n15279), .B(n15280), .Z(n15173) );
  NANDN U15506 ( .A(n15281), .B(n15282), .Z(n15280) );
  OR U15507 ( .A(n15283), .B(n15284), .Z(n15282) );
  NAND U15508 ( .A(n15284), .B(n15283), .Z(n15279) );
  ANDN U15509 ( .B(B[189]), .A(n40), .Z(n15175) );
  XNOR U15510 ( .A(n15183), .B(n15285), .Z(n15176) );
  XNOR U15511 ( .A(n15182), .B(n15180), .Z(n15285) );
  AND U15512 ( .A(n15286), .B(n15287), .Z(n15180) );
  NANDN U15513 ( .A(n15288), .B(n15289), .Z(n15287) );
  NAND U15514 ( .A(n15290), .B(n15291), .Z(n15289) );
  ANDN U15515 ( .B(B[190]), .A(n41), .Z(n15182) );
  XOR U15516 ( .A(n15189), .B(n15292), .Z(n15183) );
  XNOR U15517 ( .A(n15187), .B(n15190), .Z(n15292) );
  NAND U15518 ( .A(A[2]), .B(B[191]), .Z(n15190) );
  NANDN U15519 ( .A(n15293), .B(n15294), .Z(n15187) );
  AND U15520 ( .A(A[0]), .B(B[192]), .Z(n15294) );
  XNOR U15521 ( .A(n15192), .B(n15295), .Z(n15189) );
  NAND U15522 ( .A(A[0]), .B(B[193]), .Z(n15295) );
  NAND U15523 ( .A(B[192]), .B(A[1]), .Z(n15192) );
  NAND U15524 ( .A(n15296), .B(n15297), .Z(n361) );
  NANDN U15525 ( .A(n15298), .B(n15299), .Z(n15297) );
  OR U15526 ( .A(n15300), .B(n15301), .Z(n15299) );
  NAND U15527 ( .A(n15301), .B(n15300), .Z(n15296) );
  XOR U15528 ( .A(n363), .B(n362), .Z(\A1[190] ) );
  XOR U15529 ( .A(n15301), .B(n15302), .Z(n362) );
  XNOR U15530 ( .A(n15300), .B(n15298), .Z(n15302) );
  AND U15531 ( .A(n15303), .B(n15304), .Z(n15298) );
  NANDN U15532 ( .A(n15305), .B(n15306), .Z(n15304) );
  NANDN U15533 ( .A(n15307), .B(n15308), .Z(n15306) );
  NANDN U15534 ( .A(n15308), .B(n15307), .Z(n15303) );
  ANDN U15535 ( .B(B[177]), .A(n29), .Z(n15300) );
  XNOR U15536 ( .A(n15207), .B(n15309), .Z(n15301) );
  XNOR U15537 ( .A(n15206), .B(n15204), .Z(n15309) );
  AND U15538 ( .A(n15310), .B(n15311), .Z(n15204) );
  NANDN U15539 ( .A(n15312), .B(n15313), .Z(n15311) );
  OR U15540 ( .A(n15314), .B(n15315), .Z(n15313) );
  NAND U15541 ( .A(n15315), .B(n15314), .Z(n15310) );
  ANDN U15542 ( .B(B[178]), .A(n30), .Z(n15206) );
  XNOR U15543 ( .A(n15214), .B(n15316), .Z(n15207) );
  XNOR U15544 ( .A(n15213), .B(n15211), .Z(n15316) );
  AND U15545 ( .A(n15317), .B(n15318), .Z(n15211) );
  NANDN U15546 ( .A(n15319), .B(n15320), .Z(n15318) );
  NANDN U15547 ( .A(n15321), .B(n15322), .Z(n15320) );
  NANDN U15548 ( .A(n15322), .B(n15321), .Z(n15317) );
  ANDN U15549 ( .B(B[179]), .A(n31), .Z(n15213) );
  XNOR U15550 ( .A(n15221), .B(n15323), .Z(n15214) );
  XNOR U15551 ( .A(n15220), .B(n15218), .Z(n15323) );
  AND U15552 ( .A(n15324), .B(n15325), .Z(n15218) );
  NANDN U15553 ( .A(n15326), .B(n15327), .Z(n15325) );
  OR U15554 ( .A(n15328), .B(n15329), .Z(n15327) );
  NAND U15555 ( .A(n15329), .B(n15328), .Z(n15324) );
  ANDN U15556 ( .B(B[180]), .A(n32), .Z(n15220) );
  XNOR U15557 ( .A(n15228), .B(n15330), .Z(n15221) );
  XNOR U15558 ( .A(n15227), .B(n15225), .Z(n15330) );
  AND U15559 ( .A(n15331), .B(n15332), .Z(n15225) );
  NANDN U15560 ( .A(n15333), .B(n15334), .Z(n15332) );
  NANDN U15561 ( .A(n15335), .B(n15336), .Z(n15334) );
  NANDN U15562 ( .A(n15336), .B(n15335), .Z(n15331) );
  ANDN U15563 ( .B(B[181]), .A(n33), .Z(n15227) );
  XNOR U15564 ( .A(n15235), .B(n15337), .Z(n15228) );
  XNOR U15565 ( .A(n15234), .B(n15232), .Z(n15337) );
  AND U15566 ( .A(n15338), .B(n15339), .Z(n15232) );
  NANDN U15567 ( .A(n15340), .B(n15341), .Z(n15339) );
  OR U15568 ( .A(n15342), .B(n15343), .Z(n15341) );
  NAND U15569 ( .A(n15343), .B(n15342), .Z(n15338) );
  ANDN U15570 ( .B(B[182]), .A(n34), .Z(n15234) );
  XNOR U15571 ( .A(n15242), .B(n15344), .Z(n15235) );
  XNOR U15572 ( .A(n15241), .B(n15239), .Z(n15344) );
  AND U15573 ( .A(n15345), .B(n15346), .Z(n15239) );
  NANDN U15574 ( .A(n15347), .B(n15348), .Z(n15346) );
  NANDN U15575 ( .A(n15349), .B(n15350), .Z(n15348) );
  NANDN U15576 ( .A(n15350), .B(n15349), .Z(n15345) );
  ANDN U15577 ( .B(B[183]), .A(n35), .Z(n15241) );
  XNOR U15578 ( .A(n15249), .B(n15351), .Z(n15242) );
  XNOR U15579 ( .A(n15248), .B(n15246), .Z(n15351) );
  AND U15580 ( .A(n15352), .B(n15353), .Z(n15246) );
  NANDN U15581 ( .A(n15354), .B(n15355), .Z(n15353) );
  OR U15582 ( .A(n15356), .B(n15357), .Z(n15355) );
  NAND U15583 ( .A(n15357), .B(n15356), .Z(n15352) );
  ANDN U15584 ( .B(B[184]), .A(n36), .Z(n15248) );
  XNOR U15585 ( .A(n15256), .B(n15358), .Z(n15249) );
  XNOR U15586 ( .A(n15255), .B(n15253), .Z(n15358) );
  AND U15587 ( .A(n15359), .B(n15360), .Z(n15253) );
  NANDN U15588 ( .A(n15361), .B(n15362), .Z(n15360) );
  NANDN U15589 ( .A(n15363), .B(n15364), .Z(n15362) );
  NANDN U15590 ( .A(n15364), .B(n15363), .Z(n15359) );
  ANDN U15591 ( .B(B[185]), .A(n37), .Z(n15255) );
  XNOR U15592 ( .A(n15263), .B(n15365), .Z(n15256) );
  XNOR U15593 ( .A(n15262), .B(n15260), .Z(n15365) );
  AND U15594 ( .A(n15366), .B(n15367), .Z(n15260) );
  NANDN U15595 ( .A(n15368), .B(n15369), .Z(n15367) );
  OR U15596 ( .A(n15370), .B(n15371), .Z(n15369) );
  NAND U15597 ( .A(n15371), .B(n15370), .Z(n15366) );
  ANDN U15598 ( .B(B[186]), .A(n38), .Z(n15262) );
  XNOR U15599 ( .A(n15270), .B(n15372), .Z(n15263) );
  XNOR U15600 ( .A(n15269), .B(n15267), .Z(n15372) );
  AND U15601 ( .A(n15373), .B(n15374), .Z(n15267) );
  NANDN U15602 ( .A(n15375), .B(n15376), .Z(n15374) );
  NANDN U15603 ( .A(n15377), .B(n15378), .Z(n15376) );
  NANDN U15604 ( .A(n15378), .B(n15377), .Z(n15373) );
  ANDN U15605 ( .B(B[187]), .A(n39), .Z(n15269) );
  XNOR U15606 ( .A(n15277), .B(n15379), .Z(n15270) );
  XNOR U15607 ( .A(n15276), .B(n15274), .Z(n15379) );
  AND U15608 ( .A(n15380), .B(n15381), .Z(n15274) );
  NANDN U15609 ( .A(n15382), .B(n15383), .Z(n15381) );
  OR U15610 ( .A(n15384), .B(n15385), .Z(n15383) );
  NAND U15611 ( .A(n15385), .B(n15384), .Z(n15380) );
  ANDN U15612 ( .B(B[188]), .A(n40), .Z(n15276) );
  XNOR U15613 ( .A(n15284), .B(n15386), .Z(n15277) );
  XNOR U15614 ( .A(n15283), .B(n15281), .Z(n15386) );
  AND U15615 ( .A(n15387), .B(n15388), .Z(n15281) );
  NANDN U15616 ( .A(n15389), .B(n15390), .Z(n15388) );
  NAND U15617 ( .A(n15391), .B(n15392), .Z(n15390) );
  ANDN U15618 ( .B(B[189]), .A(n41), .Z(n15283) );
  XOR U15619 ( .A(n15290), .B(n15393), .Z(n15284) );
  XNOR U15620 ( .A(n15288), .B(n15291), .Z(n15393) );
  NAND U15621 ( .A(A[2]), .B(B[190]), .Z(n15291) );
  NANDN U15622 ( .A(n15394), .B(n15395), .Z(n15288) );
  AND U15623 ( .A(A[0]), .B(B[191]), .Z(n15395) );
  XNOR U15624 ( .A(n15293), .B(n15396), .Z(n15290) );
  NAND U15625 ( .A(A[0]), .B(B[192]), .Z(n15396) );
  NAND U15626 ( .A(B[191]), .B(A[1]), .Z(n15293) );
  NAND U15627 ( .A(n15397), .B(n15398), .Z(n363) );
  NANDN U15628 ( .A(n15399), .B(n15400), .Z(n15398) );
  OR U15629 ( .A(n15401), .B(n15402), .Z(n15400) );
  NAND U15630 ( .A(n15402), .B(n15401), .Z(n15397) );
  XOR U15631 ( .A(n345), .B(n344), .Z(\A1[18] ) );
  XOR U15632 ( .A(n14392), .B(n15403), .Z(n344) );
  XNOR U15633 ( .A(n14391), .B(n14389), .Z(n15403) );
  AND U15634 ( .A(n15404), .B(n15405), .Z(n14389) );
  NANDN U15635 ( .A(n15406), .B(n15407), .Z(n15405) );
  NANDN U15636 ( .A(n15408), .B(n15409), .Z(n15407) );
  NANDN U15637 ( .A(n15409), .B(n15408), .Z(n15404) );
  ANDN U15638 ( .B(B[5]), .A(n29), .Z(n14391) );
  XNOR U15639 ( .A(n14298), .B(n15410), .Z(n14392) );
  XNOR U15640 ( .A(n14297), .B(n14295), .Z(n15410) );
  AND U15641 ( .A(n15411), .B(n15412), .Z(n14295) );
  NANDN U15642 ( .A(n15413), .B(n15414), .Z(n15412) );
  OR U15643 ( .A(n15415), .B(n15416), .Z(n15414) );
  NAND U15644 ( .A(n15416), .B(n15415), .Z(n15411) );
  ANDN U15645 ( .B(B[6]), .A(n30), .Z(n14297) );
  XNOR U15646 ( .A(n14305), .B(n15417), .Z(n14298) );
  XNOR U15647 ( .A(n14304), .B(n14302), .Z(n15417) );
  AND U15648 ( .A(n15418), .B(n15419), .Z(n14302) );
  NANDN U15649 ( .A(n15420), .B(n15421), .Z(n15419) );
  NANDN U15650 ( .A(n15422), .B(n15423), .Z(n15421) );
  NANDN U15651 ( .A(n15423), .B(n15422), .Z(n15418) );
  ANDN U15652 ( .B(B[7]), .A(n31), .Z(n14304) );
  XNOR U15653 ( .A(n14312), .B(n15424), .Z(n14305) );
  XNOR U15654 ( .A(n14311), .B(n14309), .Z(n15424) );
  AND U15655 ( .A(n15425), .B(n15426), .Z(n14309) );
  NANDN U15656 ( .A(n15427), .B(n15428), .Z(n15426) );
  OR U15657 ( .A(n15429), .B(n15430), .Z(n15428) );
  NAND U15658 ( .A(n15430), .B(n15429), .Z(n15425) );
  ANDN U15659 ( .B(B[8]), .A(n32), .Z(n14311) );
  XNOR U15660 ( .A(n14319), .B(n15431), .Z(n14312) );
  XNOR U15661 ( .A(n14318), .B(n14316), .Z(n15431) );
  AND U15662 ( .A(n15432), .B(n15433), .Z(n14316) );
  NANDN U15663 ( .A(n15434), .B(n15435), .Z(n15433) );
  NANDN U15664 ( .A(n15436), .B(n15437), .Z(n15435) );
  NANDN U15665 ( .A(n15437), .B(n15436), .Z(n15432) );
  ANDN U15666 ( .B(B[9]), .A(n33), .Z(n14318) );
  XNOR U15667 ( .A(n14326), .B(n15438), .Z(n14319) );
  XNOR U15668 ( .A(n14325), .B(n14323), .Z(n15438) );
  AND U15669 ( .A(n15439), .B(n15440), .Z(n14323) );
  NANDN U15670 ( .A(n15441), .B(n15442), .Z(n15440) );
  OR U15671 ( .A(n15443), .B(n15444), .Z(n15442) );
  NAND U15672 ( .A(n15444), .B(n15443), .Z(n15439) );
  ANDN U15673 ( .B(B[10]), .A(n34), .Z(n14325) );
  XNOR U15674 ( .A(n14333), .B(n15445), .Z(n14326) );
  XNOR U15675 ( .A(n14332), .B(n14330), .Z(n15445) );
  AND U15676 ( .A(n15446), .B(n15447), .Z(n14330) );
  NANDN U15677 ( .A(n15448), .B(n15449), .Z(n15447) );
  NANDN U15678 ( .A(n15450), .B(n15451), .Z(n15449) );
  NANDN U15679 ( .A(n15451), .B(n15450), .Z(n15446) );
  ANDN U15680 ( .B(B[11]), .A(n35), .Z(n14332) );
  XNOR U15681 ( .A(n14340), .B(n15452), .Z(n14333) );
  XNOR U15682 ( .A(n14339), .B(n14337), .Z(n15452) );
  AND U15683 ( .A(n15453), .B(n15454), .Z(n14337) );
  NANDN U15684 ( .A(n15455), .B(n15456), .Z(n15454) );
  OR U15685 ( .A(n15457), .B(n15458), .Z(n15456) );
  NAND U15686 ( .A(n15458), .B(n15457), .Z(n15453) );
  ANDN U15687 ( .B(B[12]), .A(n36), .Z(n14339) );
  XNOR U15688 ( .A(n14347), .B(n15459), .Z(n14340) );
  XNOR U15689 ( .A(n14346), .B(n14344), .Z(n15459) );
  AND U15690 ( .A(n15460), .B(n15461), .Z(n14344) );
  NANDN U15691 ( .A(n15462), .B(n15463), .Z(n15461) );
  NANDN U15692 ( .A(n15464), .B(n15465), .Z(n15463) );
  NANDN U15693 ( .A(n15465), .B(n15464), .Z(n15460) );
  ANDN U15694 ( .B(B[13]), .A(n37), .Z(n14346) );
  XNOR U15695 ( .A(n14354), .B(n15466), .Z(n14347) );
  XNOR U15696 ( .A(n14353), .B(n14351), .Z(n15466) );
  AND U15697 ( .A(n15467), .B(n15468), .Z(n14351) );
  NANDN U15698 ( .A(n15469), .B(n15470), .Z(n15468) );
  OR U15699 ( .A(n15471), .B(n15472), .Z(n15470) );
  NAND U15700 ( .A(n15472), .B(n15471), .Z(n15467) );
  ANDN U15701 ( .B(B[14]), .A(n38), .Z(n14353) );
  XNOR U15702 ( .A(n14361), .B(n15473), .Z(n14354) );
  XNOR U15703 ( .A(n14360), .B(n14358), .Z(n15473) );
  AND U15704 ( .A(n15474), .B(n15475), .Z(n14358) );
  NANDN U15705 ( .A(n15476), .B(n15477), .Z(n15475) );
  NANDN U15706 ( .A(n15478), .B(n15479), .Z(n15477) );
  NANDN U15707 ( .A(n15479), .B(n15478), .Z(n15474) );
  ANDN U15708 ( .B(B[15]), .A(n39), .Z(n14360) );
  XNOR U15709 ( .A(n14368), .B(n15480), .Z(n14361) );
  XNOR U15710 ( .A(n14367), .B(n14365), .Z(n15480) );
  AND U15711 ( .A(n15481), .B(n15482), .Z(n14365) );
  NANDN U15712 ( .A(n15483), .B(n15484), .Z(n15482) );
  OR U15713 ( .A(n15485), .B(n15486), .Z(n15484) );
  NAND U15714 ( .A(n15486), .B(n15485), .Z(n15481) );
  ANDN U15715 ( .B(B[16]), .A(n40), .Z(n14367) );
  XNOR U15716 ( .A(n14375), .B(n15487), .Z(n14368) );
  XNOR U15717 ( .A(n14374), .B(n14372), .Z(n15487) );
  AND U15718 ( .A(n15488), .B(n15489), .Z(n14372) );
  NANDN U15719 ( .A(n15490), .B(n15491), .Z(n15489) );
  NAND U15720 ( .A(n15492), .B(n15493), .Z(n15491) );
  ANDN U15721 ( .B(B[17]), .A(n41), .Z(n14374) );
  XOR U15722 ( .A(n14381), .B(n15494), .Z(n14375) );
  XNOR U15723 ( .A(n14379), .B(n14382), .Z(n15494) );
  NAND U15724 ( .A(A[2]), .B(B[18]), .Z(n14382) );
  NANDN U15725 ( .A(n15495), .B(n15496), .Z(n14379) );
  AND U15726 ( .A(A[0]), .B(B[19]), .Z(n15496) );
  XNOR U15727 ( .A(n14384), .B(n15497), .Z(n14381) );
  NAND U15728 ( .A(A[0]), .B(B[20]), .Z(n15497) );
  NAND U15729 ( .A(B[19]), .B(A[1]), .Z(n14384) );
  NAND U15730 ( .A(n15498), .B(n15499), .Z(n345) );
  NANDN U15731 ( .A(n15500), .B(n15501), .Z(n15499) );
  OR U15732 ( .A(n15502), .B(n15503), .Z(n15501) );
  NAND U15733 ( .A(n15503), .B(n15502), .Z(n15498) );
  XOR U15734 ( .A(n365), .B(n364), .Z(\A1[189] ) );
  XOR U15735 ( .A(n15402), .B(n15504), .Z(n364) );
  XNOR U15736 ( .A(n15401), .B(n15399), .Z(n15504) );
  AND U15737 ( .A(n15505), .B(n15506), .Z(n15399) );
  NANDN U15738 ( .A(n15507), .B(n15508), .Z(n15506) );
  NANDN U15739 ( .A(n15509), .B(n15510), .Z(n15508) );
  NANDN U15740 ( .A(n15510), .B(n15509), .Z(n15505) );
  ANDN U15741 ( .B(B[176]), .A(n29), .Z(n15401) );
  XNOR U15742 ( .A(n15308), .B(n15511), .Z(n15402) );
  XNOR U15743 ( .A(n15307), .B(n15305), .Z(n15511) );
  AND U15744 ( .A(n15512), .B(n15513), .Z(n15305) );
  NANDN U15745 ( .A(n15514), .B(n15515), .Z(n15513) );
  OR U15746 ( .A(n15516), .B(n15517), .Z(n15515) );
  NAND U15747 ( .A(n15517), .B(n15516), .Z(n15512) );
  ANDN U15748 ( .B(B[177]), .A(n30), .Z(n15307) );
  XNOR U15749 ( .A(n15315), .B(n15518), .Z(n15308) );
  XNOR U15750 ( .A(n15314), .B(n15312), .Z(n15518) );
  AND U15751 ( .A(n15519), .B(n15520), .Z(n15312) );
  NANDN U15752 ( .A(n15521), .B(n15522), .Z(n15520) );
  NANDN U15753 ( .A(n15523), .B(n15524), .Z(n15522) );
  NANDN U15754 ( .A(n15524), .B(n15523), .Z(n15519) );
  ANDN U15755 ( .B(B[178]), .A(n31), .Z(n15314) );
  XNOR U15756 ( .A(n15322), .B(n15525), .Z(n15315) );
  XNOR U15757 ( .A(n15321), .B(n15319), .Z(n15525) );
  AND U15758 ( .A(n15526), .B(n15527), .Z(n15319) );
  NANDN U15759 ( .A(n15528), .B(n15529), .Z(n15527) );
  OR U15760 ( .A(n15530), .B(n15531), .Z(n15529) );
  NAND U15761 ( .A(n15531), .B(n15530), .Z(n15526) );
  ANDN U15762 ( .B(B[179]), .A(n32), .Z(n15321) );
  XNOR U15763 ( .A(n15329), .B(n15532), .Z(n15322) );
  XNOR U15764 ( .A(n15328), .B(n15326), .Z(n15532) );
  AND U15765 ( .A(n15533), .B(n15534), .Z(n15326) );
  NANDN U15766 ( .A(n15535), .B(n15536), .Z(n15534) );
  NANDN U15767 ( .A(n15537), .B(n15538), .Z(n15536) );
  NANDN U15768 ( .A(n15538), .B(n15537), .Z(n15533) );
  ANDN U15769 ( .B(B[180]), .A(n33), .Z(n15328) );
  XNOR U15770 ( .A(n15336), .B(n15539), .Z(n15329) );
  XNOR U15771 ( .A(n15335), .B(n15333), .Z(n15539) );
  AND U15772 ( .A(n15540), .B(n15541), .Z(n15333) );
  NANDN U15773 ( .A(n15542), .B(n15543), .Z(n15541) );
  OR U15774 ( .A(n15544), .B(n15545), .Z(n15543) );
  NAND U15775 ( .A(n15545), .B(n15544), .Z(n15540) );
  ANDN U15776 ( .B(B[181]), .A(n34), .Z(n15335) );
  XNOR U15777 ( .A(n15343), .B(n15546), .Z(n15336) );
  XNOR U15778 ( .A(n15342), .B(n15340), .Z(n15546) );
  AND U15779 ( .A(n15547), .B(n15548), .Z(n15340) );
  NANDN U15780 ( .A(n15549), .B(n15550), .Z(n15548) );
  NANDN U15781 ( .A(n15551), .B(n15552), .Z(n15550) );
  NANDN U15782 ( .A(n15552), .B(n15551), .Z(n15547) );
  ANDN U15783 ( .B(B[182]), .A(n35), .Z(n15342) );
  XNOR U15784 ( .A(n15350), .B(n15553), .Z(n15343) );
  XNOR U15785 ( .A(n15349), .B(n15347), .Z(n15553) );
  AND U15786 ( .A(n15554), .B(n15555), .Z(n15347) );
  NANDN U15787 ( .A(n15556), .B(n15557), .Z(n15555) );
  OR U15788 ( .A(n15558), .B(n15559), .Z(n15557) );
  NAND U15789 ( .A(n15559), .B(n15558), .Z(n15554) );
  ANDN U15790 ( .B(B[183]), .A(n36), .Z(n15349) );
  XNOR U15791 ( .A(n15357), .B(n15560), .Z(n15350) );
  XNOR U15792 ( .A(n15356), .B(n15354), .Z(n15560) );
  AND U15793 ( .A(n15561), .B(n15562), .Z(n15354) );
  NANDN U15794 ( .A(n15563), .B(n15564), .Z(n15562) );
  NANDN U15795 ( .A(n15565), .B(n15566), .Z(n15564) );
  NANDN U15796 ( .A(n15566), .B(n15565), .Z(n15561) );
  ANDN U15797 ( .B(B[184]), .A(n37), .Z(n15356) );
  XNOR U15798 ( .A(n15364), .B(n15567), .Z(n15357) );
  XNOR U15799 ( .A(n15363), .B(n15361), .Z(n15567) );
  AND U15800 ( .A(n15568), .B(n15569), .Z(n15361) );
  NANDN U15801 ( .A(n15570), .B(n15571), .Z(n15569) );
  OR U15802 ( .A(n15572), .B(n15573), .Z(n15571) );
  NAND U15803 ( .A(n15573), .B(n15572), .Z(n15568) );
  ANDN U15804 ( .B(B[185]), .A(n38), .Z(n15363) );
  XNOR U15805 ( .A(n15371), .B(n15574), .Z(n15364) );
  XNOR U15806 ( .A(n15370), .B(n15368), .Z(n15574) );
  AND U15807 ( .A(n15575), .B(n15576), .Z(n15368) );
  NANDN U15808 ( .A(n15577), .B(n15578), .Z(n15576) );
  NANDN U15809 ( .A(n15579), .B(n15580), .Z(n15578) );
  NANDN U15810 ( .A(n15580), .B(n15579), .Z(n15575) );
  ANDN U15811 ( .B(B[186]), .A(n39), .Z(n15370) );
  XNOR U15812 ( .A(n15378), .B(n15581), .Z(n15371) );
  XNOR U15813 ( .A(n15377), .B(n15375), .Z(n15581) );
  AND U15814 ( .A(n15582), .B(n15583), .Z(n15375) );
  NANDN U15815 ( .A(n15584), .B(n15585), .Z(n15583) );
  OR U15816 ( .A(n15586), .B(n15587), .Z(n15585) );
  NAND U15817 ( .A(n15587), .B(n15586), .Z(n15582) );
  ANDN U15818 ( .B(B[187]), .A(n40), .Z(n15377) );
  XNOR U15819 ( .A(n15385), .B(n15588), .Z(n15378) );
  XNOR U15820 ( .A(n15384), .B(n15382), .Z(n15588) );
  AND U15821 ( .A(n15589), .B(n15590), .Z(n15382) );
  NANDN U15822 ( .A(n15591), .B(n15592), .Z(n15590) );
  NAND U15823 ( .A(n15593), .B(n15594), .Z(n15592) );
  ANDN U15824 ( .B(B[188]), .A(n41), .Z(n15384) );
  XOR U15825 ( .A(n15391), .B(n15595), .Z(n15385) );
  XNOR U15826 ( .A(n15389), .B(n15392), .Z(n15595) );
  NAND U15827 ( .A(A[2]), .B(B[189]), .Z(n15392) );
  NANDN U15828 ( .A(n15596), .B(n15597), .Z(n15389) );
  AND U15829 ( .A(A[0]), .B(B[190]), .Z(n15597) );
  XNOR U15830 ( .A(n15394), .B(n15598), .Z(n15391) );
  NAND U15831 ( .A(A[0]), .B(B[191]), .Z(n15598) );
  NAND U15832 ( .A(B[190]), .B(A[1]), .Z(n15394) );
  NAND U15833 ( .A(n15599), .B(n15600), .Z(n365) );
  NANDN U15834 ( .A(n15601), .B(n15602), .Z(n15600) );
  OR U15835 ( .A(n15603), .B(n15604), .Z(n15602) );
  NAND U15836 ( .A(n15604), .B(n15603), .Z(n15599) );
  XOR U15837 ( .A(n369), .B(n368), .Z(\A1[188] ) );
  XOR U15838 ( .A(n15604), .B(n15605), .Z(n368) );
  XNOR U15839 ( .A(n15603), .B(n15601), .Z(n15605) );
  AND U15840 ( .A(n15606), .B(n15607), .Z(n15601) );
  NANDN U15841 ( .A(n15608), .B(n15609), .Z(n15607) );
  NANDN U15842 ( .A(n15610), .B(n15611), .Z(n15609) );
  NANDN U15843 ( .A(n15611), .B(n15610), .Z(n15606) );
  ANDN U15844 ( .B(B[175]), .A(n29), .Z(n15603) );
  XNOR U15845 ( .A(n15510), .B(n15612), .Z(n15604) );
  XNOR U15846 ( .A(n15509), .B(n15507), .Z(n15612) );
  AND U15847 ( .A(n15613), .B(n15614), .Z(n15507) );
  NANDN U15848 ( .A(n15615), .B(n15616), .Z(n15614) );
  OR U15849 ( .A(n15617), .B(n15618), .Z(n15616) );
  NAND U15850 ( .A(n15618), .B(n15617), .Z(n15613) );
  ANDN U15851 ( .B(B[176]), .A(n30), .Z(n15509) );
  XNOR U15852 ( .A(n15517), .B(n15619), .Z(n15510) );
  XNOR U15853 ( .A(n15516), .B(n15514), .Z(n15619) );
  AND U15854 ( .A(n15620), .B(n15621), .Z(n15514) );
  NANDN U15855 ( .A(n15622), .B(n15623), .Z(n15621) );
  NANDN U15856 ( .A(n15624), .B(n15625), .Z(n15623) );
  NANDN U15857 ( .A(n15625), .B(n15624), .Z(n15620) );
  ANDN U15858 ( .B(B[177]), .A(n31), .Z(n15516) );
  XNOR U15859 ( .A(n15524), .B(n15626), .Z(n15517) );
  XNOR U15860 ( .A(n15523), .B(n15521), .Z(n15626) );
  AND U15861 ( .A(n15627), .B(n15628), .Z(n15521) );
  NANDN U15862 ( .A(n15629), .B(n15630), .Z(n15628) );
  OR U15863 ( .A(n15631), .B(n15632), .Z(n15630) );
  NAND U15864 ( .A(n15632), .B(n15631), .Z(n15627) );
  ANDN U15865 ( .B(B[178]), .A(n32), .Z(n15523) );
  XNOR U15866 ( .A(n15531), .B(n15633), .Z(n15524) );
  XNOR U15867 ( .A(n15530), .B(n15528), .Z(n15633) );
  AND U15868 ( .A(n15634), .B(n15635), .Z(n15528) );
  NANDN U15869 ( .A(n15636), .B(n15637), .Z(n15635) );
  NANDN U15870 ( .A(n15638), .B(n15639), .Z(n15637) );
  NANDN U15871 ( .A(n15639), .B(n15638), .Z(n15634) );
  ANDN U15872 ( .B(B[179]), .A(n33), .Z(n15530) );
  XNOR U15873 ( .A(n15538), .B(n15640), .Z(n15531) );
  XNOR U15874 ( .A(n15537), .B(n15535), .Z(n15640) );
  AND U15875 ( .A(n15641), .B(n15642), .Z(n15535) );
  NANDN U15876 ( .A(n15643), .B(n15644), .Z(n15642) );
  OR U15877 ( .A(n15645), .B(n15646), .Z(n15644) );
  NAND U15878 ( .A(n15646), .B(n15645), .Z(n15641) );
  ANDN U15879 ( .B(B[180]), .A(n34), .Z(n15537) );
  XNOR U15880 ( .A(n15545), .B(n15647), .Z(n15538) );
  XNOR U15881 ( .A(n15544), .B(n15542), .Z(n15647) );
  AND U15882 ( .A(n15648), .B(n15649), .Z(n15542) );
  NANDN U15883 ( .A(n15650), .B(n15651), .Z(n15649) );
  NANDN U15884 ( .A(n15652), .B(n15653), .Z(n15651) );
  NANDN U15885 ( .A(n15653), .B(n15652), .Z(n15648) );
  ANDN U15886 ( .B(B[181]), .A(n35), .Z(n15544) );
  XNOR U15887 ( .A(n15552), .B(n15654), .Z(n15545) );
  XNOR U15888 ( .A(n15551), .B(n15549), .Z(n15654) );
  AND U15889 ( .A(n15655), .B(n15656), .Z(n15549) );
  NANDN U15890 ( .A(n15657), .B(n15658), .Z(n15656) );
  OR U15891 ( .A(n15659), .B(n15660), .Z(n15658) );
  NAND U15892 ( .A(n15660), .B(n15659), .Z(n15655) );
  ANDN U15893 ( .B(B[182]), .A(n36), .Z(n15551) );
  XNOR U15894 ( .A(n15559), .B(n15661), .Z(n15552) );
  XNOR U15895 ( .A(n15558), .B(n15556), .Z(n15661) );
  AND U15896 ( .A(n15662), .B(n15663), .Z(n15556) );
  NANDN U15897 ( .A(n15664), .B(n15665), .Z(n15663) );
  NANDN U15898 ( .A(n15666), .B(n15667), .Z(n15665) );
  NANDN U15899 ( .A(n15667), .B(n15666), .Z(n15662) );
  ANDN U15900 ( .B(B[183]), .A(n37), .Z(n15558) );
  XNOR U15901 ( .A(n15566), .B(n15668), .Z(n15559) );
  XNOR U15902 ( .A(n15565), .B(n15563), .Z(n15668) );
  AND U15903 ( .A(n15669), .B(n15670), .Z(n15563) );
  NANDN U15904 ( .A(n15671), .B(n15672), .Z(n15670) );
  OR U15905 ( .A(n15673), .B(n15674), .Z(n15672) );
  NAND U15906 ( .A(n15674), .B(n15673), .Z(n15669) );
  ANDN U15907 ( .B(B[184]), .A(n38), .Z(n15565) );
  XNOR U15908 ( .A(n15573), .B(n15675), .Z(n15566) );
  XNOR U15909 ( .A(n15572), .B(n15570), .Z(n15675) );
  AND U15910 ( .A(n15676), .B(n15677), .Z(n15570) );
  NANDN U15911 ( .A(n15678), .B(n15679), .Z(n15677) );
  NANDN U15912 ( .A(n15680), .B(n15681), .Z(n15679) );
  NANDN U15913 ( .A(n15681), .B(n15680), .Z(n15676) );
  ANDN U15914 ( .B(B[185]), .A(n39), .Z(n15572) );
  XNOR U15915 ( .A(n15580), .B(n15682), .Z(n15573) );
  XNOR U15916 ( .A(n15579), .B(n15577), .Z(n15682) );
  AND U15917 ( .A(n15683), .B(n15684), .Z(n15577) );
  NANDN U15918 ( .A(n15685), .B(n15686), .Z(n15684) );
  OR U15919 ( .A(n15687), .B(n15688), .Z(n15686) );
  NAND U15920 ( .A(n15688), .B(n15687), .Z(n15683) );
  ANDN U15921 ( .B(B[186]), .A(n40), .Z(n15579) );
  XNOR U15922 ( .A(n15587), .B(n15689), .Z(n15580) );
  XNOR U15923 ( .A(n15586), .B(n15584), .Z(n15689) );
  AND U15924 ( .A(n15690), .B(n15691), .Z(n15584) );
  NANDN U15925 ( .A(n15692), .B(n15693), .Z(n15691) );
  NAND U15926 ( .A(n15694), .B(n15695), .Z(n15693) );
  ANDN U15927 ( .B(B[187]), .A(n41), .Z(n15586) );
  XOR U15928 ( .A(n15593), .B(n15696), .Z(n15587) );
  XNOR U15929 ( .A(n15591), .B(n15594), .Z(n15696) );
  NAND U15930 ( .A(A[2]), .B(B[188]), .Z(n15594) );
  NANDN U15931 ( .A(n15697), .B(n15698), .Z(n15591) );
  AND U15932 ( .A(A[0]), .B(B[189]), .Z(n15698) );
  XNOR U15933 ( .A(n15596), .B(n15699), .Z(n15593) );
  NAND U15934 ( .A(A[0]), .B(B[190]), .Z(n15699) );
  NAND U15935 ( .A(B[189]), .B(A[1]), .Z(n15596) );
  NAND U15936 ( .A(n15700), .B(n15701), .Z(n369) );
  NANDN U15937 ( .A(n15702), .B(n15703), .Z(n15701) );
  OR U15938 ( .A(n15704), .B(n15705), .Z(n15703) );
  NAND U15939 ( .A(n15705), .B(n15704), .Z(n15700) );
  XOR U15940 ( .A(n371), .B(n370), .Z(\A1[187] ) );
  XOR U15941 ( .A(n15705), .B(n15706), .Z(n370) );
  XNOR U15942 ( .A(n15704), .B(n15702), .Z(n15706) );
  AND U15943 ( .A(n15707), .B(n15708), .Z(n15702) );
  NANDN U15944 ( .A(n15709), .B(n15710), .Z(n15708) );
  NANDN U15945 ( .A(n15711), .B(n15712), .Z(n15710) );
  NANDN U15946 ( .A(n15712), .B(n15711), .Z(n15707) );
  ANDN U15947 ( .B(B[174]), .A(n29), .Z(n15704) );
  XNOR U15948 ( .A(n15611), .B(n15713), .Z(n15705) );
  XNOR U15949 ( .A(n15610), .B(n15608), .Z(n15713) );
  AND U15950 ( .A(n15714), .B(n15715), .Z(n15608) );
  NANDN U15951 ( .A(n15716), .B(n15717), .Z(n15715) );
  OR U15952 ( .A(n15718), .B(n15719), .Z(n15717) );
  NAND U15953 ( .A(n15719), .B(n15718), .Z(n15714) );
  ANDN U15954 ( .B(B[175]), .A(n30), .Z(n15610) );
  XNOR U15955 ( .A(n15618), .B(n15720), .Z(n15611) );
  XNOR U15956 ( .A(n15617), .B(n15615), .Z(n15720) );
  AND U15957 ( .A(n15721), .B(n15722), .Z(n15615) );
  NANDN U15958 ( .A(n15723), .B(n15724), .Z(n15722) );
  NANDN U15959 ( .A(n15725), .B(n15726), .Z(n15724) );
  NANDN U15960 ( .A(n15726), .B(n15725), .Z(n15721) );
  ANDN U15961 ( .B(B[176]), .A(n31), .Z(n15617) );
  XNOR U15962 ( .A(n15625), .B(n15727), .Z(n15618) );
  XNOR U15963 ( .A(n15624), .B(n15622), .Z(n15727) );
  AND U15964 ( .A(n15728), .B(n15729), .Z(n15622) );
  NANDN U15965 ( .A(n15730), .B(n15731), .Z(n15729) );
  OR U15966 ( .A(n15732), .B(n15733), .Z(n15731) );
  NAND U15967 ( .A(n15733), .B(n15732), .Z(n15728) );
  ANDN U15968 ( .B(B[177]), .A(n32), .Z(n15624) );
  XNOR U15969 ( .A(n15632), .B(n15734), .Z(n15625) );
  XNOR U15970 ( .A(n15631), .B(n15629), .Z(n15734) );
  AND U15971 ( .A(n15735), .B(n15736), .Z(n15629) );
  NANDN U15972 ( .A(n15737), .B(n15738), .Z(n15736) );
  NANDN U15973 ( .A(n15739), .B(n15740), .Z(n15738) );
  NANDN U15974 ( .A(n15740), .B(n15739), .Z(n15735) );
  ANDN U15975 ( .B(B[178]), .A(n33), .Z(n15631) );
  XNOR U15976 ( .A(n15639), .B(n15741), .Z(n15632) );
  XNOR U15977 ( .A(n15638), .B(n15636), .Z(n15741) );
  AND U15978 ( .A(n15742), .B(n15743), .Z(n15636) );
  NANDN U15979 ( .A(n15744), .B(n15745), .Z(n15743) );
  OR U15980 ( .A(n15746), .B(n15747), .Z(n15745) );
  NAND U15981 ( .A(n15747), .B(n15746), .Z(n15742) );
  ANDN U15982 ( .B(B[179]), .A(n34), .Z(n15638) );
  XNOR U15983 ( .A(n15646), .B(n15748), .Z(n15639) );
  XNOR U15984 ( .A(n15645), .B(n15643), .Z(n15748) );
  AND U15985 ( .A(n15749), .B(n15750), .Z(n15643) );
  NANDN U15986 ( .A(n15751), .B(n15752), .Z(n15750) );
  NANDN U15987 ( .A(n15753), .B(n15754), .Z(n15752) );
  NANDN U15988 ( .A(n15754), .B(n15753), .Z(n15749) );
  ANDN U15989 ( .B(B[180]), .A(n35), .Z(n15645) );
  XNOR U15990 ( .A(n15653), .B(n15755), .Z(n15646) );
  XNOR U15991 ( .A(n15652), .B(n15650), .Z(n15755) );
  AND U15992 ( .A(n15756), .B(n15757), .Z(n15650) );
  NANDN U15993 ( .A(n15758), .B(n15759), .Z(n15757) );
  OR U15994 ( .A(n15760), .B(n15761), .Z(n15759) );
  NAND U15995 ( .A(n15761), .B(n15760), .Z(n15756) );
  ANDN U15996 ( .B(B[181]), .A(n36), .Z(n15652) );
  XNOR U15997 ( .A(n15660), .B(n15762), .Z(n15653) );
  XNOR U15998 ( .A(n15659), .B(n15657), .Z(n15762) );
  AND U15999 ( .A(n15763), .B(n15764), .Z(n15657) );
  NANDN U16000 ( .A(n15765), .B(n15766), .Z(n15764) );
  NANDN U16001 ( .A(n15767), .B(n15768), .Z(n15766) );
  NANDN U16002 ( .A(n15768), .B(n15767), .Z(n15763) );
  ANDN U16003 ( .B(B[182]), .A(n37), .Z(n15659) );
  XNOR U16004 ( .A(n15667), .B(n15769), .Z(n15660) );
  XNOR U16005 ( .A(n15666), .B(n15664), .Z(n15769) );
  AND U16006 ( .A(n15770), .B(n15771), .Z(n15664) );
  NANDN U16007 ( .A(n15772), .B(n15773), .Z(n15771) );
  OR U16008 ( .A(n15774), .B(n15775), .Z(n15773) );
  NAND U16009 ( .A(n15775), .B(n15774), .Z(n15770) );
  ANDN U16010 ( .B(B[183]), .A(n38), .Z(n15666) );
  XNOR U16011 ( .A(n15674), .B(n15776), .Z(n15667) );
  XNOR U16012 ( .A(n15673), .B(n15671), .Z(n15776) );
  AND U16013 ( .A(n15777), .B(n15778), .Z(n15671) );
  NANDN U16014 ( .A(n15779), .B(n15780), .Z(n15778) );
  NANDN U16015 ( .A(n15781), .B(n15782), .Z(n15780) );
  NANDN U16016 ( .A(n15782), .B(n15781), .Z(n15777) );
  ANDN U16017 ( .B(B[184]), .A(n39), .Z(n15673) );
  XNOR U16018 ( .A(n15681), .B(n15783), .Z(n15674) );
  XNOR U16019 ( .A(n15680), .B(n15678), .Z(n15783) );
  AND U16020 ( .A(n15784), .B(n15785), .Z(n15678) );
  NANDN U16021 ( .A(n15786), .B(n15787), .Z(n15785) );
  OR U16022 ( .A(n15788), .B(n15789), .Z(n15787) );
  NAND U16023 ( .A(n15789), .B(n15788), .Z(n15784) );
  ANDN U16024 ( .B(B[185]), .A(n40), .Z(n15680) );
  XNOR U16025 ( .A(n15688), .B(n15790), .Z(n15681) );
  XNOR U16026 ( .A(n15687), .B(n15685), .Z(n15790) );
  AND U16027 ( .A(n15791), .B(n15792), .Z(n15685) );
  NANDN U16028 ( .A(n15793), .B(n15794), .Z(n15792) );
  NAND U16029 ( .A(n15795), .B(n15796), .Z(n15794) );
  ANDN U16030 ( .B(B[186]), .A(n41), .Z(n15687) );
  XOR U16031 ( .A(n15694), .B(n15797), .Z(n15688) );
  XNOR U16032 ( .A(n15692), .B(n15695), .Z(n15797) );
  NAND U16033 ( .A(A[2]), .B(B[187]), .Z(n15695) );
  NANDN U16034 ( .A(n15798), .B(n15799), .Z(n15692) );
  AND U16035 ( .A(A[0]), .B(B[188]), .Z(n15799) );
  XNOR U16036 ( .A(n15697), .B(n15800), .Z(n15694) );
  NAND U16037 ( .A(A[0]), .B(B[189]), .Z(n15800) );
  NAND U16038 ( .A(B[188]), .B(A[1]), .Z(n15697) );
  NAND U16039 ( .A(n15801), .B(n15802), .Z(n371) );
  NANDN U16040 ( .A(n15803), .B(n15804), .Z(n15802) );
  OR U16041 ( .A(n15805), .B(n15806), .Z(n15804) );
  NAND U16042 ( .A(n15806), .B(n15805), .Z(n15801) );
  XOR U16043 ( .A(n373), .B(n372), .Z(\A1[186] ) );
  XOR U16044 ( .A(n15806), .B(n15807), .Z(n372) );
  XNOR U16045 ( .A(n15805), .B(n15803), .Z(n15807) );
  AND U16046 ( .A(n15808), .B(n15809), .Z(n15803) );
  NANDN U16047 ( .A(n15810), .B(n15811), .Z(n15809) );
  NANDN U16048 ( .A(n15812), .B(n15813), .Z(n15811) );
  NANDN U16049 ( .A(n15813), .B(n15812), .Z(n15808) );
  ANDN U16050 ( .B(B[173]), .A(n29), .Z(n15805) );
  XNOR U16051 ( .A(n15712), .B(n15814), .Z(n15806) );
  XNOR U16052 ( .A(n15711), .B(n15709), .Z(n15814) );
  AND U16053 ( .A(n15815), .B(n15816), .Z(n15709) );
  NANDN U16054 ( .A(n15817), .B(n15818), .Z(n15816) );
  OR U16055 ( .A(n15819), .B(n15820), .Z(n15818) );
  NAND U16056 ( .A(n15820), .B(n15819), .Z(n15815) );
  ANDN U16057 ( .B(B[174]), .A(n30), .Z(n15711) );
  XNOR U16058 ( .A(n15719), .B(n15821), .Z(n15712) );
  XNOR U16059 ( .A(n15718), .B(n15716), .Z(n15821) );
  AND U16060 ( .A(n15822), .B(n15823), .Z(n15716) );
  NANDN U16061 ( .A(n15824), .B(n15825), .Z(n15823) );
  NANDN U16062 ( .A(n15826), .B(n15827), .Z(n15825) );
  NANDN U16063 ( .A(n15827), .B(n15826), .Z(n15822) );
  ANDN U16064 ( .B(B[175]), .A(n31), .Z(n15718) );
  XNOR U16065 ( .A(n15726), .B(n15828), .Z(n15719) );
  XNOR U16066 ( .A(n15725), .B(n15723), .Z(n15828) );
  AND U16067 ( .A(n15829), .B(n15830), .Z(n15723) );
  NANDN U16068 ( .A(n15831), .B(n15832), .Z(n15830) );
  OR U16069 ( .A(n15833), .B(n15834), .Z(n15832) );
  NAND U16070 ( .A(n15834), .B(n15833), .Z(n15829) );
  ANDN U16071 ( .B(B[176]), .A(n32), .Z(n15725) );
  XNOR U16072 ( .A(n15733), .B(n15835), .Z(n15726) );
  XNOR U16073 ( .A(n15732), .B(n15730), .Z(n15835) );
  AND U16074 ( .A(n15836), .B(n15837), .Z(n15730) );
  NANDN U16075 ( .A(n15838), .B(n15839), .Z(n15837) );
  NANDN U16076 ( .A(n15840), .B(n15841), .Z(n15839) );
  NANDN U16077 ( .A(n15841), .B(n15840), .Z(n15836) );
  ANDN U16078 ( .B(B[177]), .A(n33), .Z(n15732) );
  XNOR U16079 ( .A(n15740), .B(n15842), .Z(n15733) );
  XNOR U16080 ( .A(n15739), .B(n15737), .Z(n15842) );
  AND U16081 ( .A(n15843), .B(n15844), .Z(n15737) );
  NANDN U16082 ( .A(n15845), .B(n15846), .Z(n15844) );
  OR U16083 ( .A(n15847), .B(n15848), .Z(n15846) );
  NAND U16084 ( .A(n15848), .B(n15847), .Z(n15843) );
  ANDN U16085 ( .B(B[178]), .A(n34), .Z(n15739) );
  XNOR U16086 ( .A(n15747), .B(n15849), .Z(n15740) );
  XNOR U16087 ( .A(n15746), .B(n15744), .Z(n15849) );
  AND U16088 ( .A(n15850), .B(n15851), .Z(n15744) );
  NANDN U16089 ( .A(n15852), .B(n15853), .Z(n15851) );
  NANDN U16090 ( .A(n15854), .B(n15855), .Z(n15853) );
  NANDN U16091 ( .A(n15855), .B(n15854), .Z(n15850) );
  ANDN U16092 ( .B(B[179]), .A(n35), .Z(n15746) );
  XNOR U16093 ( .A(n15754), .B(n15856), .Z(n15747) );
  XNOR U16094 ( .A(n15753), .B(n15751), .Z(n15856) );
  AND U16095 ( .A(n15857), .B(n15858), .Z(n15751) );
  NANDN U16096 ( .A(n15859), .B(n15860), .Z(n15858) );
  OR U16097 ( .A(n15861), .B(n15862), .Z(n15860) );
  NAND U16098 ( .A(n15862), .B(n15861), .Z(n15857) );
  ANDN U16099 ( .B(B[180]), .A(n36), .Z(n15753) );
  XNOR U16100 ( .A(n15761), .B(n15863), .Z(n15754) );
  XNOR U16101 ( .A(n15760), .B(n15758), .Z(n15863) );
  AND U16102 ( .A(n15864), .B(n15865), .Z(n15758) );
  NANDN U16103 ( .A(n15866), .B(n15867), .Z(n15865) );
  NANDN U16104 ( .A(n15868), .B(n15869), .Z(n15867) );
  NANDN U16105 ( .A(n15869), .B(n15868), .Z(n15864) );
  ANDN U16106 ( .B(B[181]), .A(n37), .Z(n15760) );
  XNOR U16107 ( .A(n15768), .B(n15870), .Z(n15761) );
  XNOR U16108 ( .A(n15767), .B(n15765), .Z(n15870) );
  AND U16109 ( .A(n15871), .B(n15872), .Z(n15765) );
  NANDN U16110 ( .A(n15873), .B(n15874), .Z(n15872) );
  OR U16111 ( .A(n15875), .B(n15876), .Z(n15874) );
  NAND U16112 ( .A(n15876), .B(n15875), .Z(n15871) );
  ANDN U16113 ( .B(B[182]), .A(n38), .Z(n15767) );
  XNOR U16114 ( .A(n15775), .B(n15877), .Z(n15768) );
  XNOR U16115 ( .A(n15774), .B(n15772), .Z(n15877) );
  AND U16116 ( .A(n15878), .B(n15879), .Z(n15772) );
  NANDN U16117 ( .A(n15880), .B(n15881), .Z(n15879) );
  NANDN U16118 ( .A(n15882), .B(n15883), .Z(n15881) );
  NANDN U16119 ( .A(n15883), .B(n15882), .Z(n15878) );
  ANDN U16120 ( .B(B[183]), .A(n39), .Z(n15774) );
  XNOR U16121 ( .A(n15782), .B(n15884), .Z(n15775) );
  XNOR U16122 ( .A(n15781), .B(n15779), .Z(n15884) );
  AND U16123 ( .A(n15885), .B(n15886), .Z(n15779) );
  NANDN U16124 ( .A(n15887), .B(n15888), .Z(n15886) );
  OR U16125 ( .A(n15889), .B(n15890), .Z(n15888) );
  NAND U16126 ( .A(n15890), .B(n15889), .Z(n15885) );
  ANDN U16127 ( .B(B[184]), .A(n40), .Z(n15781) );
  XNOR U16128 ( .A(n15789), .B(n15891), .Z(n15782) );
  XNOR U16129 ( .A(n15788), .B(n15786), .Z(n15891) );
  AND U16130 ( .A(n15892), .B(n15893), .Z(n15786) );
  NANDN U16131 ( .A(n15894), .B(n15895), .Z(n15893) );
  NAND U16132 ( .A(n15896), .B(n15897), .Z(n15895) );
  ANDN U16133 ( .B(B[185]), .A(n41), .Z(n15788) );
  XOR U16134 ( .A(n15795), .B(n15898), .Z(n15789) );
  XNOR U16135 ( .A(n15793), .B(n15796), .Z(n15898) );
  NAND U16136 ( .A(A[2]), .B(B[186]), .Z(n15796) );
  NANDN U16137 ( .A(n15899), .B(n15900), .Z(n15793) );
  AND U16138 ( .A(A[0]), .B(B[187]), .Z(n15900) );
  XNOR U16139 ( .A(n15798), .B(n15901), .Z(n15795) );
  NAND U16140 ( .A(A[0]), .B(B[188]), .Z(n15901) );
  NAND U16141 ( .A(B[187]), .B(A[1]), .Z(n15798) );
  NAND U16142 ( .A(n15902), .B(n15903), .Z(n373) );
  NANDN U16143 ( .A(n15904), .B(n15905), .Z(n15903) );
  OR U16144 ( .A(n15906), .B(n15907), .Z(n15905) );
  NAND U16145 ( .A(n15907), .B(n15906), .Z(n15902) );
  XOR U16146 ( .A(n375), .B(n374), .Z(\A1[185] ) );
  XOR U16147 ( .A(n15907), .B(n15908), .Z(n374) );
  XNOR U16148 ( .A(n15906), .B(n15904), .Z(n15908) );
  AND U16149 ( .A(n15909), .B(n15910), .Z(n15904) );
  NANDN U16150 ( .A(n15911), .B(n15912), .Z(n15910) );
  NANDN U16151 ( .A(n15913), .B(n15914), .Z(n15912) );
  NANDN U16152 ( .A(n15914), .B(n15913), .Z(n15909) );
  ANDN U16153 ( .B(B[172]), .A(n29), .Z(n15906) );
  XNOR U16154 ( .A(n15813), .B(n15915), .Z(n15907) );
  XNOR U16155 ( .A(n15812), .B(n15810), .Z(n15915) );
  AND U16156 ( .A(n15916), .B(n15917), .Z(n15810) );
  NANDN U16157 ( .A(n15918), .B(n15919), .Z(n15917) );
  OR U16158 ( .A(n15920), .B(n15921), .Z(n15919) );
  NAND U16159 ( .A(n15921), .B(n15920), .Z(n15916) );
  ANDN U16160 ( .B(B[173]), .A(n30), .Z(n15812) );
  XNOR U16161 ( .A(n15820), .B(n15922), .Z(n15813) );
  XNOR U16162 ( .A(n15819), .B(n15817), .Z(n15922) );
  AND U16163 ( .A(n15923), .B(n15924), .Z(n15817) );
  NANDN U16164 ( .A(n15925), .B(n15926), .Z(n15924) );
  NANDN U16165 ( .A(n15927), .B(n15928), .Z(n15926) );
  NANDN U16166 ( .A(n15928), .B(n15927), .Z(n15923) );
  ANDN U16167 ( .B(B[174]), .A(n31), .Z(n15819) );
  XNOR U16168 ( .A(n15827), .B(n15929), .Z(n15820) );
  XNOR U16169 ( .A(n15826), .B(n15824), .Z(n15929) );
  AND U16170 ( .A(n15930), .B(n15931), .Z(n15824) );
  NANDN U16171 ( .A(n15932), .B(n15933), .Z(n15931) );
  OR U16172 ( .A(n15934), .B(n15935), .Z(n15933) );
  NAND U16173 ( .A(n15935), .B(n15934), .Z(n15930) );
  ANDN U16174 ( .B(B[175]), .A(n32), .Z(n15826) );
  XNOR U16175 ( .A(n15834), .B(n15936), .Z(n15827) );
  XNOR U16176 ( .A(n15833), .B(n15831), .Z(n15936) );
  AND U16177 ( .A(n15937), .B(n15938), .Z(n15831) );
  NANDN U16178 ( .A(n15939), .B(n15940), .Z(n15938) );
  NANDN U16179 ( .A(n15941), .B(n15942), .Z(n15940) );
  NANDN U16180 ( .A(n15942), .B(n15941), .Z(n15937) );
  ANDN U16181 ( .B(B[176]), .A(n33), .Z(n15833) );
  XNOR U16182 ( .A(n15841), .B(n15943), .Z(n15834) );
  XNOR U16183 ( .A(n15840), .B(n15838), .Z(n15943) );
  AND U16184 ( .A(n15944), .B(n15945), .Z(n15838) );
  NANDN U16185 ( .A(n15946), .B(n15947), .Z(n15945) );
  OR U16186 ( .A(n15948), .B(n15949), .Z(n15947) );
  NAND U16187 ( .A(n15949), .B(n15948), .Z(n15944) );
  ANDN U16188 ( .B(B[177]), .A(n34), .Z(n15840) );
  XNOR U16189 ( .A(n15848), .B(n15950), .Z(n15841) );
  XNOR U16190 ( .A(n15847), .B(n15845), .Z(n15950) );
  AND U16191 ( .A(n15951), .B(n15952), .Z(n15845) );
  NANDN U16192 ( .A(n15953), .B(n15954), .Z(n15952) );
  NANDN U16193 ( .A(n15955), .B(n15956), .Z(n15954) );
  NANDN U16194 ( .A(n15956), .B(n15955), .Z(n15951) );
  ANDN U16195 ( .B(B[178]), .A(n35), .Z(n15847) );
  XNOR U16196 ( .A(n15855), .B(n15957), .Z(n15848) );
  XNOR U16197 ( .A(n15854), .B(n15852), .Z(n15957) );
  AND U16198 ( .A(n15958), .B(n15959), .Z(n15852) );
  NANDN U16199 ( .A(n15960), .B(n15961), .Z(n15959) );
  OR U16200 ( .A(n15962), .B(n15963), .Z(n15961) );
  NAND U16201 ( .A(n15963), .B(n15962), .Z(n15958) );
  ANDN U16202 ( .B(B[179]), .A(n36), .Z(n15854) );
  XNOR U16203 ( .A(n15862), .B(n15964), .Z(n15855) );
  XNOR U16204 ( .A(n15861), .B(n15859), .Z(n15964) );
  AND U16205 ( .A(n15965), .B(n15966), .Z(n15859) );
  NANDN U16206 ( .A(n15967), .B(n15968), .Z(n15966) );
  NANDN U16207 ( .A(n15969), .B(n15970), .Z(n15968) );
  NANDN U16208 ( .A(n15970), .B(n15969), .Z(n15965) );
  ANDN U16209 ( .B(B[180]), .A(n37), .Z(n15861) );
  XNOR U16210 ( .A(n15869), .B(n15971), .Z(n15862) );
  XNOR U16211 ( .A(n15868), .B(n15866), .Z(n15971) );
  AND U16212 ( .A(n15972), .B(n15973), .Z(n15866) );
  NANDN U16213 ( .A(n15974), .B(n15975), .Z(n15973) );
  OR U16214 ( .A(n15976), .B(n15977), .Z(n15975) );
  NAND U16215 ( .A(n15977), .B(n15976), .Z(n15972) );
  ANDN U16216 ( .B(B[181]), .A(n38), .Z(n15868) );
  XNOR U16217 ( .A(n15876), .B(n15978), .Z(n15869) );
  XNOR U16218 ( .A(n15875), .B(n15873), .Z(n15978) );
  AND U16219 ( .A(n15979), .B(n15980), .Z(n15873) );
  NANDN U16220 ( .A(n15981), .B(n15982), .Z(n15980) );
  NANDN U16221 ( .A(n15983), .B(n15984), .Z(n15982) );
  NANDN U16222 ( .A(n15984), .B(n15983), .Z(n15979) );
  ANDN U16223 ( .B(B[182]), .A(n39), .Z(n15875) );
  XNOR U16224 ( .A(n15883), .B(n15985), .Z(n15876) );
  XNOR U16225 ( .A(n15882), .B(n15880), .Z(n15985) );
  AND U16226 ( .A(n15986), .B(n15987), .Z(n15880) );
  NANDN U16227 ( .A(n15988), .B(n15989), .Z(n15987) );
  OR U16228 ( .A(n15990), .B(n15991), .Z(n15989) );
  NAND U16229 ( .A(n15991), .B(n15990), .Z(n15986) );
  ANDN U16230 ( .B(B[183]), .A(n40), .Z(n15882) );
  XNOR U16231 ( .A(n15890), .B(n15992), .Z(n15883) );
  XNOR U16232 ( .A(n15889), .B(n15887), .Z(n15992) );
  AND U16233 ( .A(n15993), .B(n15994), .Z(n15887) );
  NANDN U16234 ( .A(n15995), .B(n15996), .Z(n15994) );
  NAND U16235 ( .A(n15997), .B(n15998), .Z(n15996) );
  ANDN U16236 ( .B(B[184]), .A(n41), .Z(n15889) );
  XOR U16237 ( .A(n15896), .B(n15999), .Z(n15890) );
  XNOR U16238 ( .A(n15894), .B(n15897), .Z(n15999) );
  NAND U16239 ( .A(A[2]), .B(B[185]), .Z(n15897) );
  NANDN U16240 ( .A(n16000), .B(n16001), .Z(n15894) );
  AND U16241 ( .A(A[0]), .B(B[186]), .Z(n16001) );
  XNOR U16242 ( .A(n15899), .B(n16002), .Z(n15896) );
  NAND U16243 ( .A(A[0]), .B(B[187]), .Z(n16002) );
  NAND U16244 ( .A(B[186]), .B(A[1]), .Z(n15899) );
  NAND U16245 ( .A(n16003), .B(n16004), .Z(n375) );
  NANDN U16246 ( .A(n16005), .B(n16006), .Z(n16004) );
  OR U16247 ( .A(n16007), .B(n16008), .Z(n16006) );
  NAND U16248 ( .A(n16008), .B(n16007), .Z(n16003) );
  XOR U16249 ( .A(n377), .B(n376), .Z(\A1[184] ) );
  XOR U16250 ( .A(n16008), .B(n16009), .Z(n376) );
  XNOR U16251 ( .A(n16007), .B(n16005), .Z(n16009) );
  AND U16252 ( .A(n16010), .B(n16011), .Z(n16005) );
  NANDN U16253 ( .A(n16012), .B(n16013), .Z(n16011) );
  NANDN U16254 ( .A(n16014), .B(n16015), .Z(n16013) );
  NANDN U16255 ( .A(n16015), .B(n16014), .Z(n16010) );
  ANDN U16256 ( .B(B[171]), .A(n29), .Z(n16007) );
  XNOR U16257 ( .A(n15914), .B(n16016), .Z(n16008) );
  XNOR U16258 ( .A(n15913), .B(n15911), .Z(n16016) );
  AND U16259 ( .A(n16017), .B(n16018), .Z(n15911) );
  NANDN U16260 ( .A(n16019), .B(n16020), .Z(n16018) );
  OR U16261 ( .A(n16021), .B(n16022), .Z(n16020) );
  NAND U16262 ( .A(n16022), .B(n16021), .Z(n16017) );
  ANDN U16263 ( .B(B[172]), .A(n30), .Z(n15913) );
  XNOR U16264 ( .A(n15921), .B(n16023), .Z(n15914) );
  XNOR U16265 ( .A(n15920), .B(n15918), .Z(n16023) );
  AND U16266 ( .A(n16024), .B(n16025), .Z(n15918) );
  NANDN U16267 ( .A(n16026), .B(n16027), .Z(n16025) );
  NANDN U16268 ( .A(n16028), .B(n16029), .Z(n16027) );
  NANDN U16269 ( .A(n16029), .B(n16028), .Z(n16024) );
  ANDN U16270 ( .B(B[173]), .A(n31), .Z(n15920) );
  XNOR U16271 ( .A(n15928), .B(n16030), .Z(n15921) );
  XNOR U16272 ( .A(n15927), .B(n15925), .Z(n16030) );
  AND U16273 ( .A(n16031), .B(n16032), .Z(n15925) );
  NANDN U16274 ( .A(n16033), .B(n16034), .Z(n16032) );
  OR U16275 ( .A(n16035), .B(n16036), .Z(n16034) );
  NAND U16276 ( .A(n16036), .B(n16035), .Z(n16031) );
  ANDN U16277 ( .B(B[174]), .A(n32), .Z(n15927) );
  XNOR U16278 ( .A(n15935), .B(n16037), .Z(n15928) );
  XNOR U16279 ( .A(n15934), .B(n15932), .Z(n16037) );
  AND U16280 ( .A(n16038), .B(n16039), .Z(n15932) );
  NANDN U16281 ( .A(n16040), .B(n16041), .Z(n16039) );
  NANDN U16282 ( .A(n16042), .B(n16043), .Z(n16041) );
  NANDN U16283 ( .A(n16043), .B(n16042), .Z(n16038) );
  ANDN U16284 ( .B(B[175]), .A(n33), .Z(n15934) );
  XNOR U16285 ( .A(n15942), .B(n16044), .Z(n15935) );
  XNOR U16286 ( .A(n15941), .B(n15939), .Z(n16044) );
  AND U16287 ( .A(n16045), .B(n16046), .Z(n15939) );
  NANDN U16288 ( .A(n16047), .B(n16048), .Z(n16046) );
  OR U16289 ( .A(n16049), .B(n16050), .Z(n16048) );
  NAND U16290 ( .A(n16050), .B(n16049), .Z(n16045) );
  ANDN U16291 ( .B(B[176]), .A(n34), .Z(n15941) );
  XNOR U16292 ( .A(n15949), .B(n16051), .Z(n15942) );
  XNOR U16293 ( .A(n15948), .B(n15946), .Z(n16051) );
  AND U16294 ( .A(n16052), .B(n16053), .Z(n15946) );
  NANDN U16295 ( .A(n16054), .B(n16055), .Z(n16053) );
  NANDN U16296 ( .A(n16056), .B(n16057), .Z(n16055) );
  NANDN U16297 ( .A(n16057), .B(n16056), .Z(n16052) );
  ANDN U16298 ( .B(B[177]), .A(n35), .Z(n15948) );
  XNOR U16299 ( .A(n15956), .B(n16058), .Z(n15949) );
  XNOR U16300 ( .A(n15955), .B(n15953), .Z(n16058) );
  AND U16301 ( .A(n16059), .B(n16060), .Z(n15953) );
  NANDN U16302 ( .A(n16061), .B(n16062), .Z(n16060) );
  OR U16303 ( .A(n16063), .B(n16064), .Z(n16062) );
  NAND U16304 ( .A(n16064), .B(n16063), .Z(n16059) );
  ANDN U16305 ( .B(B[178]), .A(n36), .Z(n15955) );
  XNOR U16306 ( .A(n15963), .B(n16065), .Z(n15956) );
  XNOR U16307 ( .A(n15962), .B(n15960), .Z(n16065) );
  AND U16308 ( .A(n16066), .B(n16067), .Z(n15960) );
  NANDN U16309 ( .A(n16068), .B(n16069), .Z(n16067) );
  NANDN U16310 ( .A(n16070), .B(n16071), .Z(n16069) );
  NANDN U16311 ( .A(n16071), .B(n16070), .Z(n16066) );
  ANDN U16312 ( .B(B[179]), .A(n37), .Z(n15962) );
  XNOR U16313 ( .A(n15970), .B(n16072), .Z(n15963) );
  XNOR U16314 ( .A(n15969), .B(n15967), .Z(n16072) );
  AND U16315 ( .A(n16073), .B(n16074), .Z(n15967) );
  NANDN U16316 ( .A(n16075), .B(n16076), .Z(n16074) );
  OR U16317 ( .A(n16077), .B(n16078), .Z(n16076) );
  NAND U16318 ( .A(n16078), .B(n16077), .Z(n16073) );
  ANDN U16319 ( .B(B[180]), .A(n38), .Z(n15969) );
  XNOR U16320 ( .A(n15977), .B(n16079), .Z(n15970) );
  XNOR U16321 ( .A(n15976), .B(n15974), .Z(n16079) );
  AND U16322 ( .A(n16080), .B(n16081), .Z(n15974) );
  NANDN U16323 ( .A(n16082), .B(n16083), .Z(n16081) );
  NANDN U16324 ( .A(n16084), .B(n16085), .Z(n16083) );
  NANDN U16325 ( .A(n16085), .B(n16084), .Z(n16080) );
  ANDN U16326 ( .B(B[181]), .A(n39), .Z(n15976) );
  XNOR U16327 ( .A(n15984), .B(n16086), .Z(n15977) );
  XNOR U16328 ( .A(n15983), .B(n15981), .Z(n16086) );
  AND U16329 ( .A(n16087), .B(n16088), .Z(n15981) );
  NANDN U16330 ( .A(n16089), .B(n16090), .Z(n16088) );
  OR U16331 ( .A(n16091), .B(n16092), .Z(n16090) );
  NAND U16332 ( .A(n16092), .B(n16091), .Z(n16087) );
  ANDN U16333 ( .B(B[182]), .A(n40), .Z(n15983) );
  XNOR U16334 ( .A(n15991), .B(n16093), .Z(n15984) );
  XNOR U16335 ( .A(n15990), .B(n15988), .Z(n16093) );
  AND U16336 ( .A(n16094), .B(n16095), .Z(n15988) );
  NANDN U16337 ( .A(n16096), .B(n16097), .Z(n16095) );
  NAND U16338 ( .A(n16098), .B(n16099), .Z(n16097) );
  ANDN U16339 ( .B(B[183]), .A(n41), .Z(n15990) );
  XOR U16340 ( .A(n15997), .B(n16100), .Z(n15991) );
  XNOR U16341 ( .A(n15995), .B(n15998), .Z(n16100) );
  NAND U16342 ( .A(A[2]), .B(B[184]), .Z(n15998) );
  NANDN U16343 ( .A(n16101), .B(n16102), .Z(n15995) );
  AND U16344 ( .A(A[0]), .B(B[185]), .Z(n16102) );
  XNOR U16345 ( .A(n16000), .B(n16103), .Z(n15997) );
  NAND U16346 ( .A(A[0]), .B(B[186]), .Z(n16103) );
  NAND U16347 ( .A(B[185]), .B(A[1]), .Z(n16000) );
  NAND U16348 ( .A(n16104), .B(n16105), .Z(n377) );
  NANDN U16349 ( .A(n16106), .B(n16107), .Z(n16105) );
  OR U16350 ( .A(n16108), .B(n16109), .Z(n16107) );
  NAND U16351 ( .A(n16109), .B(n16108), .Z(n16104) );
  XOR U16352 ( .A(n379), .B(n378), .Z(\A1[183] ) );
  XOR U16353 ( .A(n16109), .B(n16110), .Z(n378) );
  XNOR U16354 ( .A(n16108), .B(n16106), .Z(n16110) );
  AND U16355 ( .A(n16111), .B(n16112), .Z(n16106) );
  NANDN U16356 ( .A(n16113), .B(n16114), .Z(n16112) );
  NANDN U16357 ( .A(n16115), .B(n16116), .Z(n16114) );
  NANDN U16358 ( .A(n16116), .B(n16115), .Z(n16111) );
  ANDN U16359 ( .B(B[170]), .A(n29), .Z(n16108) );
  XNOR U16360 ( .A(n16015), .B(n16117), .Z(n16109) );
  XNOR U16361 ( .A(n16014), .B(n16012), .Z(n16117) );
  AND U16362 ( .A(n16118), .B(n16119), .Z(n16012) );
  NANDN U16363 ( .A(n16120), .B(n16121), .Z(n16119) );
  OR U16364 ( .A(n16122), .B(n16123), .Z(n16121) );
  NAND U16365 ( .A(n16123), .B(n16122), .Z(n16118) );
  ANDN U16366 ( .B(B[171]), .A(n30), .Z(n16014) );
  XNOR U16367 ( .A(n16022), .B(n16124), .Z(n16015) );
  XNOR U16368 ( .A(n16021), .B(n16019), .Z(n16124) );
  AND U16369 ( .A(n16125), .B(n16126), .Z(n16019) );
  NANDN U16370 ( .A(n16127), .B(n16128), .Z(n16126) );
  NANDN U16371 ( .A(n16129), .B(n16130), .Z(n16128) );
  NANDN U16372 ( .A(n16130), .B(n16129), .Z(n16125) );
  ANDN U16373 ( .B(B[172]), .A(n31), .Z(n16021) );
  XNOR U16374 ( .A(n16029), .B(n16131), .Z(n16022) );
  XNOR U16375 ( .A(n16028), .B(n16026), .Z(n16131) );
  AND U16376 ( .A(n16132), .B(n16133), .Z(n16026) );
  NANDN U16377 ( .A(n16134), .B(n16135), .Z(n16133) );
  OR U16378 ( .A(n16136), .B(n16137), .Z(n16135) );
  NAND U16379 ( .A(n16137), .B(n16136), .Z(n16132) );
  ANDN U16380 ( .B(B[173]), .A(n32), .Z(n16028) );
  XNOR U16381 ( .A(n16036), .B(n16138), .Z(n16029) );
  XNOR U16382 ( .A(n16035), .B(n16033), .Z(n16138) );
  AND U16383 ( .A(n16139), .B(n16140), .Z(n16033) );
  NANDN U16384 ( .A(n16141), .B(n16142), .Z(n16140) );
  NANDN U16385 ( .A(n16143), .B(n16144), .Z(n16142) );
  NANDN U16386 ( .A(n16144), .B(n16143), .Z(n16139) );
  ANDN U16387 ( .B(B[174]), .A(n33), .Z(n16035) );
  XNOR U16388 ( .A(n16043), .B(n16145), .Z(n16036) );
  XNOR U16389 ( .A(n16042), .B(n16040), .Z(n16145) );
  AND U16390 ( .A(n16146), .B(n16147), .Z(n16040) );
  NANDN U16391 ( .A(n16148), .B(n16149), .Z(n16147) );
  OR U16392 ( .A(n16150), .B(n16151), .Z(n16149) );
  NAND U16393 ( .A(n16151), .B(n16150), .Z(n16146) );
  ANDN U16394 ( .B(B[175]), .A(n34), .Z(n16042) );
  XNOR U16395 ( .A(n16050), .B(n16152), .Z(n16043) );
  XNOR U16396 ( .A(n16049), .B(n16047), .Z(n16152) );
  AND U16397 ( .A(n16153), .B(n16154), .Z(n16047) );
  NANDN U16398 ( .A(n16155), .B(n16156), .Z(n16154) );
  NANDN U16399 ( .A(n16157), .B(n16158), .Z(n16156) );
  NANDN U16400 ( .A(n16158), .B(n16157), .Z(n16153) );
  ANDN U16401 ( .B(B[176]), .A(n35), .Z(n16049) );
  XNOR U16402 ( .A(n16057), .B(n16159), .Z(n16050) );
  XNOR U16403 ( .A(n16056), .B(n16054), .Z(n16159) );
  AND U16404 ( .A(n16160), .B(n16161), .Z(n16054) );
  NANDN U16405 ( .A(n16162), .B(n16163), .Z(n16161) );
  OR U16406 ( .A(n16164), .B(n16165), .Z(n16163) );
  NAND U16407 ( .A(n16165), .B(n16164), .Z(n16160) );
  ANDN U16408 ( .B(B[177]), .A(n36), .Z(n16056) );
  XNOR U16409 ( .A(n16064), .B(n16166), .Z(n16057) );
  XNOR U16410 ( .A(n16063), .B(n16061), .Z(n16166) );
  AND U16411 ( .A(n16167), .B(n16168), .Z(n16061) );
  NANDN U16412 ( .A(n16169), .B(n16170), .Z(n16168) );
  NANDN U16413 ( .A(n16171), .B(n16172), .Z(n16170) );
  NANDN U16414 ( .A(n16172), .B(n16171), .Z(n16167) );
  ANDN U16415 ( .B(B[178]), .A(n37), .Z(n16063) );
  XNOR U16416 ( .A(n16071), .B(n16173), .Z(n16064) );
  XNOR U16417 ( .A(n16070), .B(n16068), .Z(n16173) );
  AND U16418 ( .A(n16174), .B(n16175), .Z(n16068) );
  NANDN U16419 ( .A(n16176), .B(n16177), .Z(n16175) );
  OR U16420 ( .A(n16178), .B(n16179), .Z(n16177) );
  NAND U16421 ( .A(n16179), .B(n16178), .Z(n16174) );
  ANDN U16422 ( .B(B[179]), .A(n38), .Z(n16070) );
  XNOR U16423 ( .A(n16078), .B(n16180), .Z(n16071) );
  XNOR U16424 ( .A(n16077), .B(n16075), .Z(n16180) );
  AND U16425 ( .A(n16181), .B(n16182), .Z(n16075) );
  NANDN U16426 ( .A(n16183), .B(n16184), .Z(n16182) );
  NANDN U16427 ( .A(n16185), .B(n16186), .Z(n16184) );
  NANDN U16428 ( .A(n16186), .B(n16185), .Z(n16181) );
  ANDN U16429 ( .B(B[180]), .A(n39), .Z(n16077) );
  XNOR U16430 ( .A(n16085), .B(n16187), .Z(n16078) );
  XNOR U16431 ( .A(n16084), .B(n16082), .Z(n16187) );
  AND U16432 ( .A(n16188), .B(n16189), .Z(n16082) );
  NANDN U16433 ( .A(n16190), .B(n16191), .Z(n16189) );
  OR U16434 ( .A(n16192), .B(n16193), .Z(n16191) );
  NAND U16435 ( .A(n16193), .B(n16192), .Z(n16188) );
  ANDN U16436 ( .B(B[181]), .A(n40), .Z(n16084) );
  XNOR U16437 ( .A(n16092), .B(n16194), .Z(n16085) );
  XNOR U16438 ( .A(n16091), .B(n16089), .Z(n16194) );
  AND U16439 ( .A(n16195), .B(n16196), .Z(n16089) );
  NANDN U16440 ( .A(n16197), .B(n16198), .Z(n16196) );
  NAND U16441 ( .A(n16199), .B(n16200), .Z(n16198) );
  ANDN U16442 ( .B(B[182]), .A(n41), .Z(n16091) );
  XOR U16443 ( .A(n16098), .B(n16201), .Z(n16092) );
  XNOR U16444 ( .A(n16096), .B(n16099), .Z(n16201) );
  NAND U16445 ( .A(A[2]), .B(B[183]), .Z(n16099) );
  NANDN U16446 ( .A(n16202), .B(n16203), .Z(n16096) );
  AND U16447 ( .A(A[0]), .B(B[184]), .Z(n16203) );
  XNOR U16448 ( .A(n16101), .B(n16204), .Z(n16098) );
  NAND U16449 ( .A(A[0]), .B(B[185]), .Z(n16204) );
  NAND U16450 ( .A(B[184]), .B(A[1]), .Z(n16101) );
  NAND U16451 ( .A(n16205), .B(n16206), .Z(n379) );
  NANDN U16452 ( .A(n16207), .B(n16208), .Z(n16206) );
  OR U16453 ( .A(n16209), .B(n16210), .Z(n16208) );
  NAND U16454 ( .A(n16210), .B(n16209), .Z(n16205) );
  XOR U16455 ( .A(n381), .B(n380), .Z(\A1[182] ) );
  XOR U16456 ( .A(n16210), .B(n16211), .Z(n380) );
  XNOR U16457 ( .A(n16209), .B(n16207), .Z(n16211) );
  AND U16458 ( .A(n16212), .B(n16213), .Z(n16207) );
  NANDN U16459 ( .A(n16214), .B(n16215), .Z(n16213) );
  NANDN U16460 ( .A(n16216), .B(n16217), .Z(n16215) );
  NANDN U16461 ( .A(n16217), .B(n16216), .Z(n16212) );
  ANDN U16462 ( .B(B[169]), .A(n29), .Z(n16209) );
  XNOR U16463 ( .A(n16116), .B(n16218), .Z(n16210) );
  XNOR U16464 ( .A(n16115), .B(n16113), .Z(n16218) );
  AND U16465 ( .A(n16219), .B(n16220), .Z(n16113) );
  NANDN U16466 ( .A(n16221), .B(n16222), .Z(n16220) );
  OR U16467 ( .A(n16223), .B(n16224), .Z(n16222) );
  NAND U16468 ( .A(n16224), .B(n16223), .Z(n16219) );
  ANDN U16469 ( .B(B[170]), .A(n30), .Z(n16115) );
  XNOR U16470 ( .A(n16123), .B(n16225), .Z(n16116) );
  XNOR U16471 ( .A(n16122), .B(n16120), .Z(n16225) );
  AND U16472 ( .A(n16226), .B(n16227), .Z(n16120) );
  NANDN U16473 ( .A(n16228), .B(n16229), .Z(n16227) );
  NANDN U16474 ( .A(n16230), .B(n16231), .Z(n16229) );
  NANDN U16475 ( .A(n16231), .B(n16230), .Z(n16226) );
  ANDN U16476 ( .B(B[171]), .A(n31), .Z(n16122) );
  XNOR U16477 ( .A(n16130), .B(n16232), .Z(n16123) );
  XNOR U16478 ( .A(n16129), .B(n16127), .Z(n16232) );
  AND U16479 ( .A(n16233), .B(n16234), .Z(n16127) );
  NANDN U16480 ( .A(n16235), .B(n16236), .Z(n16234) );
  OR U16481 ( .A(n16237), .B(n16238), .Z(n16236) );
  NAND U16482 ( .A(n16238), .B(n16237), .Z(n16233) );
  ANDN U16483 ( .B(B[172]), .A(n32), .Z(n16129) );
  XNOR U16484 ( .A(n16137), .B(n16239), .Z(n16130) );
  XNOR U16485 ( .A(n16136), .B(n16134), .Z(n16239) );
  AND U16486 ( .A(n16240), .B(n16241), .Z(n16134) );
  NANDN U16487 ( .A(n16242), .B(n16243), .Z(n16241) );
  NANDN U16488 ( .A(n16244), .B(n16245), .Z(n16243) );
  NANDN U16489 ( .A(n16245), .B(n16244), .Z(n16240) );
  ANDN U16490 ( .B(B[173]), .A(n33), .Z(n16136) );
  XNOR U16491 ( .A(n16144), .B(n16246), .Z(n16137) );
  XNOR U16492 ( .A(n16143), .B(n16141), .Z(n16246) );
  AND U16493 ( .A(n16247), .B(n16248), .Z(n16141) );
  NANDN U16494 ( .A(n16249), .B(n16250), .Z(n16248) );
  OR U16495 ( .A(n16251), .B(n16252), .Z(n16250) );
  NAND U16496 ( .A(n16252), .B(n16251), .Z(n16247) );
  ANDN U16497 ( .B(B[174]), .A(n34), .Z(n16143) );
  XNOR U16498 ( .A(n16151), .B(n16253), .Z(n16144) );
  XNOR U16499 ( .A(n16150), .B(n16148), .Z(n16253) );
  AND U16500 ( .A(n16254), .B(n16255), .Z(n16148) );
  NANDN U16501 ( .A(n16256), .B(n16257), .Z(n16255) );
  NANDN U16502 ( .A(n16258), .B(n16259), .Z(n16257) );
  NANDN U16503 ( .A(n16259), .B(n16258), .Z(n16254) );
  ANDN U16504 ( .B(B[175]), .A(n35), .Z(n16150) );
  XNOR U16505 ( .A(n16158), .B(n16260), .Z(n16151) );
  XNOR U16506 ( .A(n16157), .B(n16155), .Z(n16260) );
  AND U16507 ( .A(n16261), .B(n16262), .Z(n16155) );
  NANDN U16508 ( .A(n16263), .B(n16264), .Z(n16262) );
  OR U16509 ( .A(n16265), .B(n16266), .Z(n16264) );
  NAND U16510 ( .A(n16266), .B(n16265), .Z(n16261) );
  ANDN U16511 ( .B(B[176]), .A(n36), .Z(n16157) );
  XNOR U16512 ( .A(n16165), .B(n16267), .Z(n16158) );
  XNOR U16513 ( .A(n16164), .B(n16162), .Z(n16267) );
  AND U16514 ( .A(n16268), .B(n16269), .Z(n16162) );
  NANDN U16515 ( .A(n16270), .B(n16271), .Z(n16269) );
  NANDN U16516 ( .A(n16272), .B(n16273), .Z(n16271) );
  NANDN U16517 ( .A(n16273), .B(n16272), .Z(n16268) );
  ANDN U16518 ( .B(B[177]), .A(n37), .Z(n16164) );
  XNOR U16519 ( .A(n16172), .B(n16274), .Z(n16165) );
  XNOR U16520 ( .A(n16171), .B(n16169), .Z(n16274) );
  AND U16521 ( .A(n16275), .B(n16276), .Z(n16169) );
  NANDN U16522 ( .A(n16277), .B(n16278), .Z(n16276) );
  OR U16523 ( .A(n16279), .B(n16280), .Z(n16278) );
  NAND U16524 ( .A(n16280), .B(n16279), .Z(n16275) );
  ANDN U16525 ( .B(B[178]), .A(n38), .Z(n16171) );
  XNOR U16526 ( .A(n16179), .B(n16281), .Z(n16172) );
  XNOR U16527 ( .A(n16178), .B(n16176), .Z(n16281) );
  AND U16528 ( .A(n16282), .B(n16283), .Z(n16176) );
  NANDN U16529 ( .A(n16284), .B(n16285), .Z(n16283) );
  NANDN U16530 ( .A(n16286), .B(n16287), .Z(n16285) );
  NANDN U16531 ( .A(n16287), .B(n16286), .Z(n16282) );
  ANDN U16532 ( .B(B[179]), .A(n39), .Z(n16178) );
  XNOR U16533 ( .A(n16186), .B(n16288), .Z(n16179) );
  XNOR U16534 ( .A(n16185), .B(n16183), .Z(n16288) );
  AND U16535 ( .A(n16289), .B(n16290), .Z(n16183) );
  NANDN U16536 ( .A(n16291), .B(n16292), .Z(n16290) );
  OR U16537 ( .A(n16293), .B(n16294), .Z(n16292) );
  NAND U16538 ( .A(n16294), .B(n16293), .Z(n16289) );
  ANDN U16539 ( .B(B[180]), .A(n40), .Z(n16185) );
  XNOR U16540 ( .A(n16193), .B(n16295), .Z(n16186) );
  XNOR U16541 ( .A(n16192), .B(n16190), .Z(n16295) );
  AND U16542 ( .A(n16296), .B(n16297), .Z(n16190) );
  NANDN U16543 ( .A(n16298), .B(n16299), .Z(n16297) );
  NAND U16544 ( .A(n16300), .B(n16301), .Z(n16299) );
  ANDN U16545 ( .B(B[181]), .A(n41), .Z(n16192) );
  XOR U16546 ( .A(n16199), .B(n16302), .Z(n16193) );
  XNOR U16547 ( .A(n16197), .B(n16200), .Z(n16302) );
  NAND U16548 ( .A(A[2]), .B(B[182]), .Z(n16200) );
  NANDN U16549 ( .A(n16303), .B(n16304), .Z(n16197) );
  AND U16550 ( .A(A[0]), .B(B[183]), .Z(n16304) );
  XNOR U16551 ( .A(n16202), .B(n16305), .Z(n16199) );
  NAND U16552 ( .A(A[0]), .B(B[184]), .Z(n16305) );
  NAND U16553 ( .A(B[183]), .B(A[1]), .Z(n16202) );
  NAND U16554 ( .A(n16306), .B(n16307), .Z(n381) );
  NANDN U16555 ( .A(n16308), .B(n16309), .Z(n16307) );
  OR U16556 ( .A(n16310), .B(n16311), .Z(n16309) );
  NAND U16557 ( .A(n16311), .B(n16310), .Z(n16306) );
  XOR U16558 ( .A(n383), .B(n382), .Z(\A1[181] ) );
  XOR U16559 ( .A(n16311), .B(n16312), .Z(n382) );
  XNOR U16560 ( .A(n16310), .B(n16308), .Z(n16312) );
  AND U16561 ( .A(n16313), .B(n16314), .Z(n16308) );
  NANDN U16562 ( .A(n16315), .B(n16316), .Z(n16314) );
  NANDN U16563 ( .A(n16317), .B(n16318), .Z(n16316) );
  NANDN U16564 ( .A(n16318), .B(n16317), .Z(n16313) );
  ANDN U16565 ( .B(B[168]), .A(n29), .Z(n16310) );
  XNOR U16566 ( .A(n16217), .B(n16319), .Z(n16311) );
  XNOR U16567 ( .A(n16216), .B(n16214), .Z(n16319) );
  AND U16568 ( .A(n16320), .B(n16321), .Z(n16214) );
  NANDN U16569 ( .A(n16322), .B(n16323), .Z(n16321) );
  OR U16570 ( .A(n16324), .B(n16325), .Z(n16323) );
  NAND U16571 ( .A(n16325), .B(n16324), .Z(n16320) );
  ANDN U16572 ( .B(B[169]), .A(n30), .Z(n16216) );
  XNOR U16573 ( .A(n16224), .B(n16326), .Z(n16217) );
  XNOR U16574 ( .A(n16223), .B(n16221), .Z(n16326) );
  AND U16575 ( .A(n16327), .B(n16328), .Z(n16221) );
  NANDN U16576 ( .A(n16329), .B(n16330), .Z(n16328) );
  NANDN U16577 ( .A(n16331), .B(n16332), .Z(n16330) );
  NANDN U16578 ( .A(n16332), .B(n16331), .Z(n16327) );
  ANDN U16579 ( .B(B[170]), .A(n31), .Z(n16223) );
  XNOR U16580 ( .A(n16231), .B(n16333), .Z(n16224) );
  XNOR U16581 ( .A(n16230), .B(n16228), .Z(n16333) );
  AND U16582 ( .A(n16334), .B(n16335), .Z(n16228) );
  NANDN U16583 ( .A(n16336), .B(n16337), .Z(n16335) );
  OR U16584 ( .A(n16338), .B(n16339), .Z(n16337) );
  NAND U16585 ( .A(n16339), .B(n16338), .Z(n16334) );
  ANDN U16586 ( .B(B[171]), .A(n32), .Z(n16230) );
  XNOR U16587 ( .A(n16238), .B(n16340), .Z(n16231) );
  XNOR U16588 ( .A(n16237), .B(n16235), .Z(n16340) );
  AND U16589 ( .A(n16341), .B(n16342), .Z(n16235) );
  NANDN U16590 ( .A(n16343), .B(n16344), .Z(n16342) );
  NANDN U16591 ( .A(n16345), .B(n16346), .Z(n16344) );
  NANDN U16592 ( .A(n16346), .B(n16345), .Z(n16341) );
  ANDN U16593 ( .B(B[172]), .A(n33), .Z(n16237) );
  XNOR U16594 ( .A(n16245), .B(n16347), .Z(n16238) );
  XNOR U16595 ( .A(n16244), .B(n16242), .Z(n16347) );
  AND U16596 ( .A(n16348), .B(n16349), .Z(n16242) );
  NANDN U16597 ( .A(n16350), .B(n16351), .Z(n16349) );
  OR U16598 ( .A(n16352), .B(n16353), .Z(n16351) );
  NAND U16599 ( .A(n16353), .B(n16352), .Z(n16348) );
  ANDN U16600 ( .B(B[173]), .A(n34), .Z(n16244) );
  XNOR U16601 ( .A(n16252), .B(n16354), .Z(n16245) );
  XNOR U16602 ( .A(n16251), .B(n16249), .Z(n16354) );
  AND U16603 ( .A(n16355), .B(n16356), .Z(n16249) );
  NANDN U16604 ( .A(n16357), .B(n16358), .Z(n16356) );
  NANDN U16605 ( .A(n16359), .B(n16360), .Z(n16358) );
  NANDN U16606 ( .A(n16360), .B(n16359), .Z(n16355) );
  ANDN U16607 ( .B(B[174]), .A(n35), .Z(n16251) );
  XNOR U16608 ( .A(n16259), .B(n16361), .Z(n16252) );
  XNOR U16609 ( .A(n16258), .B(n16256), .Z(n16361) );
  AND U16610 ( .A(n16362), .B(n16363), .Z(n16256) );
  NANDN U16611 ( .A(n16364), .B(n16365), .Z(n16363) );
  OR U16612 ( .A(n16366), .B(n16367), .Z(n16365) );
  NAND U16613 ( .A(n16367), .B(n16366), .Z(n16362) );
  ANDN U16614 ( .B(B[175]), .A(n36), .Z(n16258) );
  XNOR U16615 ( .A(n16266), .B(n16368), .Z(n16259) );
  XNOR U16616 ( .A(n16265), .B(n16263), .Z(n16368) );
  AND U16617 ( .A(n16369), .B(n16370), .Z(n16263) );
  NANDN U16618 ( .A(n16371), .B(n16372), .Z(n16370) );
  NANDN U16619 ( .A(n16373), .B(n16374), .Z(n16372) );
  NANDN U16620 ( .A(n16374), .B(n16373), .Z(n16369) );
  ANDN U16621 ( .B(B[176]), .A(n37), .Z(n16265) );
  XNOR U16622 ( .A(n16273), .B(n16375), .Z(n16266) );
  XNOR U16623 ( .A(n16272), .B(n16270), .Z(n16375) );
  AND U16624 ( .A(n16376), .B(n16377), .Z(n16270) );
  NANDN U16625 ( .A(n16378), .B(n16379), .Z(n16377) );
  OR U16626 ( .A(n16380), .B(n16381), .Z(n16379) );
  NAND U16627 ( .A(n16381), .B(n16380), .Z(n16376) );
  ANDN U16628 ( .B(B[177]), .A(n38), .Z(n16272) );
  XNOR U16629 ( .A(n16280), .B(n16382), .Z(n16273) );
  XNOR U16630 ( .A(n16279), .B(n16277), .Z(n16382) );
  AND U16631 ( .A(n16383), .B(n16384), .Z(n16277) );
  NANDN U16632 ( .A(n16385), .B(n16386), .Z(n16384) );
  NANDN U16633 ( .A(n16387), .B(n16388), .Z(n16386) );
  NANDN U16634 ( .A(n16388), .B(n16387), .Z(n16383) );
  ANDN U16635 ( .B(B[178]), .A(n39), .Z(n16279) );
  XNOR U16636 ( .A(n16287), .B(n16389), .Z(n16280) );
  XNOR U16637 ( .A(n16286), .B(n16284), .Z(n16389) );
  AND U16638 ( .A(n16390), .B(n16391), .Z(n16284) );
  NANDN U16639 ( .A(n16392), .B(n16393), .Z(n16391) );
  OR U16640 ( .A(n16394), .B(n16395), .Z(n16393) );
  NAND U16641 ( .A(n16395), .B(n16394), .Z(n16390) );
  ANDN U16642 ( .B(B[179]), .A(n40), .Z(n16286) );
  XNOR U16643 ( .A(n16294), .B(n16396), .Z(n16287) );
  XNOR U16644 ( .A(n16293), .B(n16291), .Z(n16396) );
  AND U16645 ( .A(n16397), .B(n16398), .Z(n16291) );
  NANDN U16646 ( .A(n16399), .B(n16400), .Z(n16398) );
  NAND U16647 ( .A(n16401), .B(n16402), .Z(n16400) );
  ANDN U16648 ( .B(B[180]), .A(n41), .Z(n16293) );
  XOR U16649 ( .A(n16300), .B(n16403), .Z(n16294) );
  XNOR U16650 ( .A(n16298), .B(n16301), .Z(n16403) );
  NAND U16651 ( .A(A[2]), .B(B[181]), .Z(n16301) );
  NANDN U16652 ( .A(n16404), .B(n16405), .Z(n16298) );
  AND U16653 ( .A(A[0]), .B(B[182]), .Z(n16405) );
  XNOR U16654 ( .A(n16303), .B(n16406), .Z(n16300) );
  NAND U16655 ( .A(A[0]), .B(B[183]), .Z(n16406) );
  NAND U16656 ( .A(B[182]), .B(A[1]), .Z(n16303) );
  NAND U16657 ( .A(n16407), .B(n16408), .Z(n383) );
  NANDN U16658 ( .A(n16409), .B(n16410), .Z(n16408) );
  OR U16659 ( .A(n16411), .B(n16412), .Z(n16410) );
  NAND U16660 ( .A(n16412), .B(n16411), .Z(n16407) );
  XOR U16661 ( .A(n385), .B(n384), .Z(\A1[180] ) );
  XOR U16662 ( .A(n16412), .B(n16413), .Z(n384) );
  XNOR U16663 ( .A(n16411), .B(n16409), .Z(n16413) );
  AND U16664 ( .A(n16414), .B(n16415), .Z(n16409) );
  NANDN U16665 ( .A(n16416), .B(n16417), .Z(n16415) );
  NANDN U16666 ( .A(n16418), .B(n16419), .Z(n16417) );
  NANDN U16667 ( .A(n16419), .B(n16418), .Z(n16414) );
  ANDN U16668 ( .B(B[167]), .A(n29), .Z(n16411) );
  XNOR U16669 ( .A(n16318), .B(n16420), .Z(n16412) );
  XNOR U16670 ( .A(n16317), .B(n16315), .Z(n16420) );
  AND U16671 ( .A(n16421), .B(n16422), .Z(n16315) );
  NANDN U16672 ( .A(n16423), .B(n16424), .Z(n16422) );
  OR U16673 ( .A(n16425), .B(n16426), .Z(n16424) );
  NAND U16674 ( .A(n16426), .B(n16425), .Z(n16421) );
  ANDN U16675 ( .B(B[168]), .A(n30), .Z(n16317) );
  XNOR U16676 ( .A(n16325), .B(n16427), .Z(n16318) );
  XNOR U16677 ( .A(n16324), .B(n16322), .Z(n16427) );
  AND U16678 ( .A(n16428), .B(n16429), .Z(n16322) );
  NANDN U16679 ( .A(n16430), .B(n16431), .Z(n16429) );
  NANDN U16680 ( .A(n16432), .B(n16433), .Z(n16431) );
  NANDN U16681 ( .A(n16433), .B(n16432), .Z(n16428) );
  ANDN U16682 ( .B(B[169]), .A(n31), .Z(n16324) );
  XNOR U16683 ( .A(n16332), .B(n16434), .Z(n16325) );
  XNOR U16684 ( .A(n16331), .B(n16329), .Z(n16434) );
  AND U16685 ( .A(n16435), .B(n16436), .Z(n16329) );
  NANDN U16686 ( .A(n16437), .B(n16438), .Z(n16436) );
  OR U16687 ( .A(n16439), .B(n16440), .Z(n16438) );
  NAND U16688 ( .A(n16440), .B(n16439), .Z(n16435) );
  ANDN U16689 ( .B(B[170]), .A(n32), .Z(n16331) );
  XNOR U16690 ( .A(n16339), .B(n16441), .Z(n16332) );
  XNOR U16691 ( .A(n16338), .B(n16336), .Z(n16441) );
  AND U16692 ( .A(n16442), .B(n16443), .Z(n16336) );
  NANDN U16693 ( .A(n16444), .B(n16445), .Z(n16443) );
  NANDN U16694 ( .A(n16446), .B(n16447), .Z(n16445) );
  NANDN U16695 ( .A(n16447), .B(n16446), .Z(n16442) );
  ANDN U16696 ( .B(B[171]), .A(n33), .Z(n16338) );
  XNOR U16697 ( .A(n16346), .B(n16448), .Z(n16339) );
  XNOR U16698 ( .A(n16345), .B(n16343), .Z(n16448) );
  AND U16699 ( .A(n16449), .B(n16450), .Z(n16343) );
  NANDN U16700 ( .A(n16451), .B(n16452), .Z(n16450) );
  OR U16701 ( .A(n16453), .B(n16454), .Z(n16452) );
  NAND U16702 ( .A(n16454), .B(n16453), .Z(n16449) );
  ANDN U16703 ( .B(B[172]), .A(n34), .Z(n16345) );
  XNOR U16704 ( .A(n16353), .B(n16455), .Z(n16346) );
  XNOR U16705 ( .A(n16352), .B(n16350), .Z(n16455) );
  AND U16706 ( .A(n16456), .B(n16457), .Z(n16350) );
  NANDN U16707 ( .A(n16458), .B(n16459), .Z(n16457) );
  NANDN U16708 ( .A(n16460), .B(n16461), .Z(n16459) );
  NANDN U16709 ( .A(n16461), .B(n16460), .Z(n16456) );
  ANDN U16710 ( .B(B[173]), .A(n35), .Z(n16352) );
  XNOR U16711 ( .A(n16360), .B(n16462), .Z(n16353) );
  XNOR U16712 ( .A(n16359), .B(n16357), .Z(n16462) );
  AND U16713 ( .A(n16463), .B(n16464), .Z(n16357) );
  NANDN U16714 ( .A(n16465), .B(n16466), .Z(n16464) );
  OR U16715 ( .A(n16467), .B(n16468), .Z(n16466) );
  NAND U16716 ( .A(n16468), .B(n16467), .Z(n16463) );
  ANDN U16717 ( .B(B[174]), .A(n36), .Z(n16359) );
  XNOR U16718 ( .A(n16367), .B(n16469), .Z(n16360) );
  XNOR U16719 ( .A(n16366), .B(n16364), .Z(n16469) );
  AND U16720 ( .A(n16470), .B(n16471), .Z(n16364) );
  NANDN U16721 ( .A(n16472), .B(n16473), .Z(n16471) );
  NANDN U16722 ( .A(n16474), .B(n16475), .Z(n16473) );
  NANDN U16723 ( .A(n16475), .B(n16474), .Z(n16470) );
  ANDN U16724 ( .B(B[175]), .A(n37), .Z(n16366) );
  XNOR U16725 ( .A(n16374), .B(n16476), .Z(n16367) );
  XNOR U16726 ( .A(n16373), .B(n16371), .Z(n16476) );
  AND U16727 ( .A(n16477), .B(n16478), .Z(n16371) );
  NANDN U16728 ( .A(n16479), .B(n16480), .Z(n16478) );
  OR U16729 ( .A(n16481), .B(n16482), .Z(n16480) );
  NAND U16730 ( .A(n16482), .B(n16481), .Z(n16477) );
  ANDN U16731 ( .B(B[176]), .A(n38), .Z(n16373) );
  XNOR U16732 ( .A(n16381), .B(n16483), .Z(n16374) );
  XNOR U16733 ( .A(n16380), .B(n16378), .Z(n16483) );
  AND U16734 ( .A(n16484), .B(n16485), .Z(n16378) );
  NANDN U16735 ( .A(n16486), .B(n16487), .Z(n16485) );
  NANDN U16736 ( .A(n16488), .B(n16489), .Z(n16487) );
  NANDN U16737 ( .A(n16489), .B(n16488), .Z(n16484) );
  ANDN U16738 ( .B(B[177]), .A(n39), .Z(n16380) );
  XNOR U16739 ( .A(n16388), .B(n16490), .Z(n16381) );
  XNOR U16740 ( .A(n16387), .B(n16385), .Z(n16490) );
  AND U16741 ( .A(n16491), .B(n16492), .Z(n16385) );
  NANDN U16742 ( .A(n16493), .B(n16494), .Z(n16492) );
  OR U16743 ( .A(n16495), .B(n16496), .Z(n16494) );
  NAND U16744 ( .A(n16496), .B(n16495), .Z(n16491) );
  ANDN U16745 ( .B(B[178]), .A(n40), .Z(n16387) );
  XNOR U16746 ( .A(n16395), .B(n16497), .Z(n16388) );
  XNOR U16747 ( .A(n16394), .B(n16392), .Z(n16497) );
  AND U16748 ( .A(n16498), .B(n16499), .Z(n16392) );
  NANDN U16749 ( .A(n16500), .B(n16501), .Z(n16499) );
  NAND U16750 ( .A(n16502), .B(n16503), .Z(n16501) );
  ANDN U16751 ( .B(B[179]), .A(n41), .Z(n16394) );
  XOR U16752 ( .A(n16401), .B(n16504), .Z(n16395) );
  XNOR U16753 ( .A(n16399), .B(n16402), .Z(n16504) );
  NAND U16754 ( .A(A[2]), .B(B[180]), .Z(n16402) );
  NANDN U16755 ( .A(n16505), .B(n16506), .Z(n16399) );
  AND U16756 ( .A(A[0]), .B(B[181]), .Z(n16506) );
  XNOR U16757 ( .A(n16404), .B(n16507), .Z(n16401) );
  NAND U16758 ( .A(A[0]), .B(B[182]), .Z(n16507) );
  NAND U16759 ( .A(B[181]), .B(A[1]), .Z(n16404) );
  NAND U16760 ( .A(n16508), .B(n16509), .Z(n385) );
  NANDN U16761 ( .A(n16510), .B(n16511), .Z(n16509) );
  OR U16762 ( .A(n16512), .B(n16513), .Z(n16511) );
  NAND U16763 ( .A(n16513), .B(n16512), .Z(n16508) );
  XOR U16764 ( .A(n367), .B(n366), .Z(\A1[17] ) );
  XOR U16765 ( .A(n15503), .B(n16514), .Z(n366) );
  XNOR U16766 ( .A(n15502), .B(n15500), .Z(n16514) );
  AND U16767 ( .A(n16515), .B(n16516), .Z(n15500) );
  NANDN U16768 ( .A(n16517), .B(n16518), .Z(n16516) );
  NANDN U16769 ( .A(n16519), .B(n16520), .Z(n16518) );
  NANDN U16770 ( .A(n16520), .B(n16519), .Z(n16515) );
  ANDN U16771 ( .B(B[4]), .A(n29), .Z(n15502) );
  XNOR U16772 ( .A(n15409), .B(n16521), .Z(n15503) );
  XNOR U16773 ( .A(n15408), .B(n15406), .Z(n16521) );
  AND U16774 ( .A(n16522), .B(n16523), .Z(n15406) );
  NANDN U16775 ( .A(n16524), .B(n16525), .Z(n16523) );
  OR U16776 ( .A(n16526), .B(n16527), .Z(n16525) );
  NAND U16777 ( .A(n16527), .B(n16526), .Z(n16522) );
  ANDN U16778 ( .B(B[5]), .A(n30), .Z(n15408) );
  XNOR U16779 ( .A(n15416), .B(n16528), .Z(n15409) );
  XNOR U16780 ( .A(n15415), .B(n15413), .Z(n16528) );
  AND U16781 ( .A(n16529), .B(n16530), .Z(n15413) );
  NANDN U16782 ( .A(n16531), .B(n16532), .Z(n16530) );
  NANDN U16783 ( .A(n16533), .B(n16534), .Z(n16532) );
  NANDN U16784 ( .A(n16534), .B(n16533), .Z(n16529) );
  ANDN U16785 ( .B(B[6]), .A(n31), .Z(n15415) );
  XNOR U16786 ( .A(n15423), .B(n16535), .Z(n15416) );
  XNOR U16787 ( .A(n15422), .B(n15420), .Z(n16535) );
  AND U16788 ( .A(n16536), .B(n16537), .Z(n15420) );
  NANDN U16789 ( .A(n16538), .B(n16539), .Z(n16537) );
  OR U16790 ( .A(n16540), .B(n16541), .Z(n16539) );
  NAND U16791 ( .A(n16541), .B(n16540), .Z(n16536) );
  ANDN U16792 ( .B(B[7]), .A(n32), .Z(n15422) );
  XNOR U16793 ( .A(n15430), .B(n16542), .Z(n15423) );
  XNOR U16794 ( .A(n15429), .B(n15427), .Z(n16542) );
  AND U16795 ( .A(n16543), .B(n16544), .Z(n15427) );
  NANDN U16796 ( .A(n16545), .B(n16546), .Z(n16544) );
  NANDN U16797 ( .A(n16547), .B(n16548), .Z(n16546) );
  NANDN U16798 ( .A(n16548), .B(n16547), .Z(n16543) );
  ANDN U16799 ( .B(B[8]), .A(n33), .Z(n15429) );
  XNOR U16800 ( .A(n15437), .B(n16549), .Z(n15430) );
  XNOR U16801 ( .A(n15436), .B(n15434), .Z(n16549) );
  AND U16802 ( .A(n16550), .B(n16551), .Z(n15434) );
  NANDN U16803 ( .A(n16552), .B(n16553), .Z(n16551) );
  OR U16804 ( .A(n16554), .B(n16555), .Z(n16553) );
  NAND U16805 ( .A(n16555), .B(n16554), .Z(n16550) );
  ANDN U16806 ( .B(B[9]), .A(n34), .Z(n15436) );
  XNOR U16807 ( .A(n15444), .B(n16556), .Z(n15437) );
  XNOR U16808 ( .A(n15443), .B(n15441), .Z(n16556) );
  AND U16809 ( .A(n16557), .B(n16558), .Z(n15441) );
  NANDN U16810 ( .A(n16559), .B(n16560), .Z(n16558) );
  NANDN U16811 ( .A(n16561), .B(n16562), .Z(n16560) );
  NANDN U16812 ( .A(n16562), .B(n16561), .Z(n16557) );
  ANDN U16813 ( .B(B[10]), .A(n35), .Z(n15443) );
  XNOR U16814 ( .A(n15451), .B(n16563), .Z(n15444) );
  XNOR U16815 ( .A(n15450), .B(n15448), .Z(n16563) );
  AND U16816 ( .A(n16564), .B(n16565), .Z(n15448) );
  NANDN U16817 ( .A(n16566), .B(n16567), .Z(n16565) );
  OR U16818 ( .A(n16568), .B(n16569), .Z(n16567) );
  NAND U16819 ( .A(n16569), .B(n16568), .Z(n16564) );
  ANDN U16820 ( .B(B[11]), .A(n36), .Z(n15450) );
  XNOR U16821 ( .A(n15458), .B(n16570), .Z(n15451) );
  XNOR U16822 ( .A(n15457), .B(n15455), .Z(n16570) );
  AND U16823 ( .A(n16571), .B(n16572), .Z(n15455) );
  NANDN U16824 ( .A(n16573), .B(n16574), .Z(n16572) );
  NANDN U16825 ( .A(n16575), .B(n16576), .Z(n16574) );
  NANDN U16826 ( .A(n16576), .B(n16575), .Z(n16571) );
  ANDN U16827 ( .B(B[12]), .A(n37), .Z(n15457) );
  XNOR U16828 ( .A(n15465), .B(n16577), .Z(n15458) );
  XNOR U16829 ( .A(n15464), .B(n15462), .Z(n16577) );
  AND U16830 ( .A(n16578), .B(n16579), .Z(n15462) );
  NANDN U16831 ( .A(n16580), .B(n16581), .Z(n16579) );
  OR U16832 ( .A(n16582), .B(n16583), .Z(n16581) );
  NAND U16833 ( .A(n16583), .B(n16582), .Z(n16578) );
  ANDN U16834 ( .B(B[13]), .A(n38), .Z(n15464) );
  XNOR U16835 ( .A(n15472), .B(n16584), .Z(n15465) );
  XNOR U16836 ( .A(n15471), .B(n15469), .Z(n16584) );
  AND U16837 ( .A(n16585), .B(n16586), .Z(n15469) );
  NANDN U16838 ( .A(n16587), .B(n16588), .Z(n16586) );
  NANDN U16839 ( .A(n16589), .B(n16590), .Z(n16588) );
  NANDN U16840 ( .A(n16590), .B(n16589), .Z(n16585) );
  ANDN U16841 ( .B(B[14]), .A(n39), .Z(n15471) );
  XNOR U16842 ( .A(n15479), .B(n16591), .Z(n15472) );
  XNOR U16843 ( .A(n15478), .B(n15476), .Z(n16591) );
  AND U16844 ( .A(n16592), .B(n16593), .Z(n15476) );
  NANDN U16845 ( .A(n16594), .B(n16595), .Z(n16593) );
  OR U16846 ( .A(n16596), .B(n16597), .Z(n16595) );
  NAND U16847 ( .A(n16597), .B(n16596), .Z(n16592) );
  ANDN U16848 ( .B(B[15]), .A(n40), .Z(n15478) );
  XNOR U16849 ( .A(n15486), .B(n16598), .Z(n15479) );
  XNOR U16850 ( .A(n15485), .B(n15483), .Z(n16598) );
  AND U16851 ( .A(n16599), .B(n16600), .Z(n15483) );
  NANDN U16852 ( .A(n16601), .B(n16602), .Z(n16600) );
  NAND U16853 ( .A(n16603), .B(n16604), .Z(n16602) );
  ANDN U16854 ( .B(B[16]), .A(n41), .Z(n15485) );
  XOR U16855 ( .A(n15492), .B(n16605), .Z(n15486) );
  XNOR U16856 ( .A(n15490), .B(n15493), .Z(n16605) );
  NAND U16857 ( .A(A[2]), .B(B[17]), .Z(n15493) );
  NANDN U16858 ( .A(n16606), .B(n16607), .Z(n15490) );
  AND U16859 ( .A(A[0]), .B(B[18]), .Z(n16607) );
  XNOR U16860 ( .A(n15495), .B(n16608), .Z(n15492) );
  NAND U16861 ( .A(A[0]), .B(B[19]), .Z(n16608) );
  NAND U16862 ( .A(B[18]), .B(A[1]), .Z(n15495) );
  NAND U16863 ( .A(n16609), .B(n16610), .Z(n367) );
  NANDN U16864 ( .A(n16611), .B(n16612), .Z(n16610) );
  OR U16865 ( .A(n16613), .B(n16614), .Z(n16612) );
  NAND U16866 ( .A(n16614), .B(n16613), .Z(n16609) );
  XOR U16867 ( .A(n387), .B(n386), .Z(\A1[179] ) );
  XOR U16868 ( .A(n16513), .B(n16615), .Z(n386) );
  XNOR U16869 ( .A(n16512), .B(n16510), .Z(n16615) );
  AND U16870 ( .A(n16616), .B(n16617), .Z(n16510) );
  NANDN U16871 ( .A(n16618), .B(n16619), .Z(n16617) );
  NANDN U16872 ( .A(n16620), .B(n16621), .Z(n16619) );
  NANDN U16873 ( .A(n16621), .B(n16620), .Z(n16616) );
  ANDN U16874 ( .B(B[166]), .A(n29), .Z(n16512) );
  XNOR U16875 ( .A(n16419), .B(n16622), .Z(n16513) );
  XNOR U16876 ( .A(n16418), .B(n16416), .Z(n16622) );
  AND U16877 ( .A(n16623), .B(n16624), .Z(n16416) );
  NANDN U16878 ( .A(n16625), .B(n16626), .Z(n16624) );
  OR U16879 ( .A(n16627), .B(n16628), .Z(n16626) );
  NAND U16880 ( .A(n16628), .B(n16627), .Z(n16623) );
  ANDN U16881 ( .B(B[167]), .A(n30), .Z(n16418) );
  XNOR U16882 ( .A(n16426), .B(n16629), .Z(n16419) );
  XNOR U16883 ( .A(n16425), .B(n16423), .Z(n16629) );
  AND U16884 ( .A(n16630), .B(n16631), .Z(n16423) );
  NANDN U16885 ( .A(n16632), .B(n16633), .Z(n16631) );
  NANDN U16886 ( .A(n16634), .B(n16635), .Z(n16633) );
  NANDN U16887 ( .A(n16635), .B(n16634), .Z(n16630) );
  ANDN U16888 ( .B(B[168]), .A(n31), .Z(n16425) );
  XNOR U16889 ( .A(n16433), .B(n16636), .Z(n16426) );
  XNOR U16890 ( .A(n16432), .B(n16430), .Z(n16636) );
  AND U16891 ( .A(n16637), .B(n16638), .Z(n16430) );
  NANDN U16892 ( .A(n16639), .B(n16640), .Z(n16638) );
  OR U16893 ( .A(n16641), .B(n16642), .Z(n16640) );
  NAND U16894 ( .A(n16642), .B(n16641), .Z(n16637) );
  ANDN U16895 ( .B(B[169]), .A(n32), .Z(n16432) );
  XNOR U16896 ( .A(n16440), .B(n16643), .Z(n16433) );
  XNOR U16897 ( .A(n16439), .B(n16437), .Z(n16643) );
  AND U16898 ( .A(n16644), .B(n16645), .Z(n16437) );
  NANDN U16899 ( .A(n16646), .B(n16647), .Z(n16645) );
  NANDN U16900 ( .A(n16648), .B(n16649), .Z(n16647) );
  NANDN U16901 ( .A(n16649), .B(n16648), .Z(n16644) );
  ANDN U16902 ( .B(B[170]), .A(n33), .Z(n16439) );
  XNOR U16903 ( .A(n16447), .B(n16650), .Z(n16440) );
  XNOR U16904 ( .A(n16446), .B(n16444), .Z(n16650) );
  AND U16905 ( .A(n16651), .B(n16652), .Z(n16444) );
  NANDN U16906 ( .A(n16653), .B(n16654), .Z(n16652) );
  OR U16907 ( .A(n16655), .B(n16656), .Z(n16654) );
  NAND U16908 ( .A(n16656), .B(n16655), .Z(n16651) );
  ANDN U16909 ( .B(B[171]), .A(n34), .Z(n16446) );
  XNOR U16910 ( .A(n16454), .B(n16657), .Z(n16447) );
  XNOR U16911 ( .A(n16453), .B(n16451), .Z(n16657) );
  AND U16912 ( .A(n16658), .B(n16659), .Z(n16451) );
  NANDN U16913 ( .A(n16660), .B(n16661), .Z(n16659) );
  NANDN U16914 ( .A(n16662), .B(n16663), .Z(n16661) );
  NANDN U16915 ( .A(n16663), .B(n16662), .Z(n16658) );
  ANDN U16916 ( .B(B[172]), .A(n35), .Z(n16453) );
  XNOR U16917 ( .A(n16461), .B(n16664), .Z(n16454) );
  XNOR U16918 ( .A(n16460), .B(n16458), .Z(n16664) );
  AND U16919 ( .A(n16665), .B(n16666), .Z(n16458) );
  NANDN U16920 ( .A(n16667), .B(n16668), .Z(n16666) );
  OR U16921 ( .A(n16669), .B(n16670), .Z(n16668) );
  NAND U16922 ( .A(n16670), .B(n16669), .Z(n16665) );
  ANDN U16923 ( .B(B[173]), .A(n36), .Z(n16460) );
  XNOR U16924 ( .A(n16468), .B(n16671), .Z(n16461) );
  XNOR U16925 ( .A(n16467), .B(n16465), .Z(n16671) );
  AND U16926 ( .A(n16672), .B(n16673), .Z(n16465) );
  NANDN U16927 ( .A(n16674), .B(n16675), .Z(n16673) );
  NANDN U16928 ( .A(n16676), .B(n16677), .Z(n16675) );
  NANDN U16929 ( .A(n16677), .B(n16676), .Z(n16672) );
  ANDN U16930 ( .B(B[174]), .A(n37), .Z(n16467) );
  XNOR U16931 ( .A(n16475), .B(n16678), .Z(n16468) );
  XNOR U16932 ( .A(n16474), .B(n16472), .Z(n16678) );
  AND U16933 ( .A(n16679), .B(n16680), .Z(n16472) );
  NANDN U16934 ( .A(n16681), .B(n16682), .Z(n16680) );
  OR U16935 ( .A(n16683), .B(n16684), .Z(n16682) );
  NAND U16936 ( .A(n16684), .B(n16683), .Z(n16679) );
  ANDN U16937 ( .B(B[175]), .A(n38), .Z(n16474) );
  XNOR U16938 ( .A(n16482), .B(n16685), .Z(n16475) );
  XNOR U16939 ( .A(n16481), .B(n16479), .Z(n16685) );
  AND U16940 ( .A(n16686), .B(n16687), .Z(n16479) );
  NANDN U16941 ( .A(n16688), .B(n16689), .Z(n16687) );
  NANDN U16942 ( .A(n16690), .B(n16691), .Z(n16689) );
  NANDN U16943 ( .A(n16691), .B(n16690), .Z(n16686) );
  ANDN U16944 ( .B(B[176]), .A(n39), .Z(n16481) );
  XNOR U16945 ( .A(n16489), .B(n16692), .Z(n16482) );
  XNOR U16946 ( .A(n16488), .B(n16486), .Z(n16692) );
  AND U16947 ( .A(n16693), .B(n16694), .Z(n16486) );
  NANDN U16948 ( .A(n16695), .B(n16696), .Z(n16694) );
  OR U16949 ( .A(n16697), .B(n16698), .Z(n16696) );
  NAND U16950 ( .A(n16698), .B(n16697), .Z(n16693) );
  ANDN U16951 ( .B(B[177]), .A(n40), .Z(n16488) );
  XNOR U16952 ( .A(n16496), .B(n16699), .Z(n16489) );
  XNOR U16953 ( .A(n16495), .B(n16493), .Z(n16699) );
  AND U16954 ( .A(n16700), .B(n16701), .Z(n16493) );
  NANDN U16955 ( .A(n16702), .B(n16703), .Z(n16701) );
  NAND U16956 ( .A(n16704), .B(n16705), .Z(n16703) );
  ANDN U16957 ( .B(B[178]), .A(n41), .Z(n16495) );
  XOR U16958 ( .A(n16502), .B(n16706), .Z(n16496) );
  XNOR U16959 ( .A(n16500), .B(n16503), .Z(n16706) );
  NAND U16960 ( .A(A[2]), .B(B[179]), .Z(n16503) );
  NANDN U16961 ( .A(n16707), .B(n16708), .Z(n16500) );
  AND U16962 ( .A(A[0]), .B(B[180]), .Z(n16708) );
  XNOR U16963 ( .A(n16505), .B(n16709), .Z(n16502) );
  NAND U16964 ( .A(A[0]), .B(B[181]), .Z(n16709) );
  NAND U16965 ( .A(B[180]), .B(A[1]), .Z(n16505) );
  NAND U16966 ( .A(n16710), .B(n16711), .Z(n387) );
  NANDN U16967 ( .A(n16712), .B(n16713), .Z(n16711) );
  OR U16968 ( .A(n16714), .B(n16715), .Z(n16713) );
  NAND U16969 ( .A(n16715), .B(n16714), .Z(n16710) );
  XOR U16970 ( .A(n391), .B(n390), .Z(\A1[178] ) );
  XOR U16971 ( .A(n16715), .B(n16716), .Z(n390) );
  XNOR U16972 ( .A(n16714), .B(n16712), .Z(n16716) );
  AND U16973 ( .A(n16717), .B(n16718), .Z(n16712) );
  NANDN U16974 ( .A(n16719), .B(n16720), .Z(n16718) );
  NANDN U16975 ( .A(n16721), .B(n16722), .Z(n16720) );
  NANDN U16976 ( .A(n16722), .B(n16721), .Z(n16717) );
  ANDN U16977 ( .B(B[165]), .A(n29), .Z(n16714) );
  XNOR U16978 ( .A(n16621), .B(n16723), .Z(n16715) );
  XNOR U16979 ( .A(n16620), .B(n16618), .Z(n16723) );
  AND U16980 ( .A(n16724), .B(n16725), .Z(n16618) );
  NANDN U16981 ( .A(n16726), .B(n16727), .Z(n16725) );
  OR U16982 ( .A(n16728), .B(n16729), .Z(n16727) );
  NAND U16983 ( .A(n16729), .B(n16728), .Z(n16724) );
  ANDN U16984 ( .B(B[166]), .A(n30), .Z(n16620) );
  XNOR U16985 ( .A(n16628), .B(n16730), .Z(n16621) );
  XNOR U16986 ( .A(n16627), .B(n16625), .Z(n16730) );
  AND U16987 ( .A(n16731), .B(n16732), .Z(n16625) );
  NANDN U16988 ( .A(n16733), .B(n16734), .Z(n16732) );
  NANDN U16989 ( .A(n16735), .B(n16736), .Z(n16734) );
  NANDN U16990 ( .A(n16736), .B(n16735), .Z(n16731) );
  ANDN U16991 ( .B(B[167]), .A(n31), .Z(n16627) );
  XNOR U16992 ( .A(n16635), .B(n16737), .Z(n16628) );
  XNOR U16993 ( .A(n16634), .B(n16632), .Z(n16737) );
  AND U16994 ( .A(n16738), .B(n16739), .Z(n16632) );
  NANDN U16995 ( .A(n16740), .B(n16741), .Z(n16739) );
  OR U16996 ( .A(n16742), .B(n16743), .Z(n16741) );
  NAND U16997 ( .A(n16743), .B(n16742), .Z(n16738) );
  ANDN U16998 ( .B(B[168]), .A(n32), .Z(n16634) );
  XNOR U16999 ( .A(n16642), .B(n16744), .Z(n16635) );
  XNOR U17000 ( .A(n16641), .B(n16639), .Z(n16744) );
  AND U17001 ( .A(n16745), .B(n16746), .Z(n16639) );
  NANDN U17002 ( .A(n16747), .B(n16748), .Z(n16746) );
  NANDN U17003 ( .A(n16749), .B(n16750), .Z(n16748) );
  NANDN U17004 ( .A(n16750), .B(n16749), .Z(n16745) );
  ANDN U17005 ( .B(B[169]), .A(n33), .Z(n16641) );
  XNOR U17006 ( .A(n16649), .B(n16751), .Z(n16642) );
  XNOR U17007 ( .A(n16648), .B(n16646), .Z(n16751) );
  AND U17008 ( .A(n16752), .B(n16753), .Z(n16646) );
  NANDN U17009 ( .A(n16754), .B(n16755), .Z(n16753) );
  OR U17010 ( .A(n16756), .B(n16757), .Z(n16755) );
  NAND U17011 ( .A(n16757), .B(n16756), .Z(n16752) );
  ANDN U17012 ( .B(B[170]), .A(n34), .Z(n16648) );
  XNOR U17013 ( .A(n16656), .B(n16758), .Z(n16649) );
  XNOR U17014 ( .A(n16655), .B(n16653), .Z(n16758) );
  AND U17015 ( .A(n16759), .B(n16760), .Z(n16653) );
  NANDN U17016 ( .A(n16761), .B(n16762), .Z(n16760) );
  NANDN U17017 ( .A(n16763), .B(n16764), .Z(n16762) );
  NANDN U17018 ( .A(n16764), .B(n16763), .Z(n16759) );
  ANDN U17019 ( .B(B[171]), .A(n35), .Z(n16655) );
  XNOR U17020 ( .A(n16663), .B(n16765), .Z(n16656) );
  XNOR U17021 ( .A(n16662), .B(n16660), .Z(n16765) );
  AND U17022 ( .A(n16766), .B(n16767), .Z(n16660) );
  NANDN U17023 ( .A(n16768), .B(n16769), .Z(n16767) );
  OR U17024 ( .A(n16770), .B(n16771), .Z(n16769) );
  NAND U17025 ( .A(n16771), .B(n16770), .Z(n16766) );
  ANDN U17026 ( .B(B[172]), .A(n36), .Z(n16662) );
  XNOR U17027 ( .A(n16670), .B(n16772), .Z(n16663) );
  XNOR U17028 ( .A(n16669), .B(n16667), .Z(n16772) );
  AND U17029 ( .A(n16773), .B(n16774), .Z(n16667) );
  NANDN U17030 ( .A(n16775), .B(n16776), .Z(n16774) );
  NANDN U17031 ( .A(n16777), .B(n16778), .Z(n16776) );
  NANDN U17032 ( .A(n16778), .B(n16777), .Z(n16773) );
  ANDN U17033 ( .B(B[173]), .A(n37), .Z(n16669) );
  XNOR U17034 ( .A(n16677), .B(n16779), .Z(n16670) );
  XNOR U17035 ( .A(n16676), .B(n16674), .Z(n16779) );
  AND U17036 ( .A(n16780), .B(n16781), .Z(n16674) );
  NANDN U17037 ( .A(n16782), .B(n16783), .Z(n16781) );
  OR U17038 ( .A(n16784), .B(n16785), .Z(n16783) );
  NAND U17039 ( .A(n16785), .B(n16784), .Z(n16780) );
  ANDN U17040 ( .B(B[174]), .A(n38), .Z(n16676) );
  XNOR U17041 ( .A(n16684), .B(n16786), .Z(n16677) );
  XNOR U17042 ( .A(n16683), .B(n16681), .Z(n16786) );
  AND U17043 ( .A(n16787), .B(n16788), .Z(n16681) );
  NANDN U17044 ( .A(n16789), .B(n16790), .Z(n16788) );
  NANDN U17045 ( .A(n16791), .B(n16792), .Z(n16790) );
  NANDN U17046 ( .A(n16792), .B(n16791), .Z(n16787) );
  ANDN U17047 ( .B(B[175]), .A(n39), .Z(n16683) );
  XNOR U17048 ( .A(n16691), .B(n16793), .Z(n16684) );
  XNOR U17049 ( .A(n16690), .B(n16688), .Z(n16793) );
  AND U17050 ( .A(n16794), .B(n16795), .Z(n16688) );
  NANDN U17051 ( .A(n16796), .B(n16797), .Z(n16795) );
  OR U17052 ( .A(n16798), .B(n16799), .Z(n16797) );
  NAND U17053 ( .A(n16799), .B(n16798), .Z(n16794) );
  ANDN U17054 ( .B(B[176]), .A(n40), .Z(n16690) );
  XNOR U17055 ( .A(n16698), .B(n16800), .Z(n16691) );
  XNOR U17056 ( .A(n16697), .B(n16695), .Z(n16800) );
  AND U17057 ( .A(n16801), .B(n16802), .Z(n16695) );
  NANDN U17058 ( .A(n16803), .B(n16804), .Z(n16802) );
  NAND U17059 ( .A(n16805), .B(n16806), .Z(n16804) );
  ANDN U17060 ( .B(B[177]), .A(n41), .Z(n16697) );
  XOR U17061 ( .A(n16704), .B(n16807), .Z(n16698) );
  XNOR U17062 ( .A(n16702), .B(n16705), .Z(n16807) );
  NAND U17063 ( .A(A[2]), .B(B[178]), .Z(n16705) );
  NANDN U17064 ( .A(n16808), .B(n16809), .Z(n16702) );
  AND U17065 ( .A(A[0]), .B(B[179]), .Z(n16809) );
  XNOR U17066 ( .A(n16707), .B(n16810), .Z(n16704) );
  NAND U17067 ( .A(A[0]), .B(B[180]), .Z(n16810) );
  NAND U17068 ( .A(B[179]), .B(A[1]), .Z(n16707) );
  NAND U17069 ( .A(n16811), .B(n16812), .Z(n391) );
  NANDN U17070 ( .A(n16813), .B(n16814), .Z(n16812) );
  OR U17071 ( .A(n16815), .B(n16816), .Z(n16814) );
  NAND U17072 ( .A(n16816), .B(n16815), .Z(n16811) );
  XOR U17073 ( .A(n393), .B(n392), .Z(\A1[177] ) );
  XOR U17074 ( .A(n16816), .B(n16817), .Z(n392) );
  XNOR U17075 ( .A(n16815), .B(n16813), .Z(n16817) );
  AND U17076 ( .A(n16818), .B(n16819), .Z(n16813) );
  NANDN U17077 ( .A(n16820), .B(n16821), .Z(n16819) );
  NANDN U17078 ( .A(n16822), .B(n16823), .Z(n16821) );
  NANDN U17079 ( .A(n16823), .B(n16822), .Z(n16818) );
  ANDN U17080 ( .B(B[164]), .A(n29), .Z(n16815) );
  XNOR U17081 ( .A(n16722), .B(n16824), .Z(n16816) );
  XNOR U17082 ( .A(n16721), .B(n16719), .Z(n16824) );
  AND U17083 ( .A(n16825), .B(n16826), .Z(n16719) );
  NANDN U17084 ( .A(n16827), .B(n16828), .Z(n16826) );
  OR U17085 ( .A(n16829), .B(n16830), .Z(n16828) );
  NAND U17086 ( .A(n16830), .B(n16829), .Z(n16825) );
  ANDN U17087 ( .B(B[165]), .A(n30), .Z(n16721) );
  XNOR U17088 ( .A(n16729), .B(n16831), .Z(n16722) );
  XNOR U17089 ( .A(n16728), .B(n16726), .Z(n16831) );
  AND U17090 ( .A(n16832), .B(n16833), .Z(n16726) );
  NANDN U17091 ( .A(n16834), .B(n16835), .Z(n16833) );
  NANDN U17092 ( .A(n16836), .B(n16837), .Z(n16835) );
  NANDN U17093 ( .A(n16837), .B(n16836), .Z(n16832) );
  ANDN U17094 ( .B(B[166]), .A(n31), .Z(n16728) );
  XNOR U17095 ( .A(n16736), .B(n16838), .Z(n16729) );
  XNOR U17096 ( .A(n16735), .B(n16733), .Z(n16838) );
  AND U17097 ( .A(n16839), .B(n16840), .Z(n16733) );
  NANDN U17098 ( .A(n16841), .B(n16842), .Z(n16840) );
  OR U17099 ( .A(n16843), .B(n16844), .Z(n16842) );
  NAND U17100 ( .A(n16844), .B(n16843), .Z(n16839) );
  ANDN U17101 ( .B(B[167]), .A(n32), .Z(n16735) );
  XNOR U17102 ( .A(n16743), .B(n16845), .Z(n16736) );
  XNOR U17103 ( .A(n16742), .B(n16740), .Z(n16845) );
  AND U17104 ( .A(n16846), .B(n16847), .Z(n16740) );
  NANDN U17105 ( .A(n16848), .B(n16849), .Z(n16847) );
  NANDN U17106 ( .A(n16850), .B(n16851), .Z(n16849) );
  NANDN U17107 ( .A(n16851), .B(n16850), .Z(n16846) );
  ANDN U17108 ( .B(B[168]), .A(n33), .Z(n16742) );
  XNOR U17109 ( .A(n16750), .B(n16852), .Z(n16743) );
  XNOR U17110 ( .A(n16749), .B(n16747), .Z(n16852) );
  AND U17111 ( .A(n16853), .B(n16854), .Z(n16747) );
  NANDN U17112 ( .A(n16855), .B(n16856), .Z(n16854) );
  OR U17113 ( .A(n16857), .B(n16858), .Z(n16856) );
  NAND U17114 ( .A(n16858), .B(n16857), .Z(n16853) );
  ANDN U17115 ( .B(B[169]), .A(n34), .Z(n16749) );
  XNOR U17116 ( .A(n16757), .B(n16859), .Z(n16750) );
  XNOR U17117 ( .A(n16756), .B(n16754), .Z(n16859) );
  AND U17118 ( .A(n16860), .B(n16861), .Z(n16754) );
  NANDN U17119 ( .A(n16862), .B(n16863), .Z(n16861) );
  NANDN U17120 ( .A(n16864), .B(n16865), .Z(n16863) );
  NANDN U17121 ( .A(n16865), .B(n16864), .Z(n16860) );
  ANDN U17122 ( .B(B[170]), .A(n35), .Z(n16756) );
  XNOR U17123 ( .A(n16764), .B(n16866), .Z(n16757) );
  XNOR U17124 ( .A(n16763), .B(n16761), .Z(n16866) );
  AND U17125 ( .A(n16867), .B(n16868), .Z(n16761) );
  NANDN U17126 ( .A(n16869), .B(n16870), .Z(n16868) );
  OR U17127 ( .A(n16871), .B(n16872), .Z(n16870) );
  NAND U17128 ( .A(n16872), .B(n16871), .Z(n16867) );
  ANDN U17129 ( .B(B[171]), .A(n36), .Z(n16763) );
  XNOR U17130 ( .A(n16771), .B(n16873), .Z(n16764) );
  XNOR U17131 ( .A(n16770), .B(n16768), .Z(n16873) );
  AND U17132 ( .A(n16874), .B(n16875), .Z(n16768) );
  NANDN U17133 ( .A(n16876), .B(n16877), .Z(n16875) );
  NANDN U17134 ( .A(n16878), .B(n16879), .Z(n16877) );
  NANDN U17135 ( .A(n16879), .B(n16878), .Z(n16874) );
  ANDN U17136 ( .B(B[172]), .A(n37), .Z(n16770) );
  XNOR U17137 ( .A(n16778), .B(n16880), .Z(n16771) );
  XNOR U17138 ( .A(n16777), .B(n16775), .Z(n16880) );
  AND U17139 ( .A(n16881), .B(n16882), .Z(n16775) );
  NANDN U17140 ( .A(n16883), .B(n16884), .Z(n16882) );
  OR U17141 ( .A(n16885), .B(n16886), .Z(n16884) );
  NAND U17142 ( .A(n16886), .B(n16885), .Z(n16881) );
  ANDN U17143 ( .B(B[173]), .A(n38), .Z(n16777) );
  XNOR U17144 ( .A(n16785), .B(n16887), .Z(n16778) );
  XNOR U17145 ( .A(n16784), .B(n16782), .Z(n16887) );
  AND U17146 ( .A(n16888), .B(n16889), .Z(n16782) );
  NANDN U17147 ( .A(n16890), .B(n16891), .Z(n16889) );
  NANDN U17148 ( .A(n16892), .B(n16893), .Z(n16891) );
  NANDN U17149 ( .A(n16893), .B(n16892), .Z(n16888) );
  ANDN U17150 ( .B(B[174]), .A(n39), .Z(n16784) );
  XNOR U17151 ( .A(n16792), .B(n16894), .Z(n16785) );
  XNOR U17152 ( .A(n16791), .B(n16789), .Z(n16894) );
  AND U17153 ( .A(n16895), .B(n16896), .Z(n16789) );
  NANDN U17154 ( .A(n16897), .B(n16898), .Z(n16896) );
  OR U17155 ( .A(n16899), .B(n16900), .Z(n16898) );
  NAND U17156 ( .A(n16900), .B(n16899), .Z(n16895) );
  ANDN U17157 ( .B(B[175]), .A(n40), .Z(n16791) );
  XNOR U17158 ( .A(n16799), .B(n16901), .Z(n16792) );
  XNOR U17159 ( .A(n16798), .B(n16796), .Z(n16901) );
  AND U17160 ( .A(n16902), .B(n16903), .Z(n16796) );
  NANDN U17161 ( .A(n16904), .B(n16905), .Z(n16903) );
  NAND U17162 ( .A(n16906), .B(n16907), .Z(n16905) );
  ANDN U17163 ( .B(B[176]), .A(n41), .Z(n16798) );
  XOR U17164 ( .A(n16805), .B(n16908), .Z(n16799) );
  XNOR U17165 ( .A(n16803), .B(n16806), .Z(n16908) );
  NAND U17166 ( .A(A[2]), .B(B[177]), .Z(n16806) );
  NANDN U17167 ( .A(n16909), .B(n16910), .Z(n16803) );
  AND U17168 ( .A(A[0]), .B(B[178]), .Z(n16910) );
  XNOR U17169 ( .A(n16808), .B(n16911), .Z(n16805) );
  NAND U17170 ( .A(A[0]), .B(B[179]), .Z(n16911) );
  NAND U17171 ( .A(B[178]), .B(A[1]), .Z(n16808) );
  NAND U17172 ( .A(n16912), .B(n16913), .Z(n393) );
  NANDN U17173 ( .A(n16914), .B(n16915), .Z(n16913) );
  OR U17174 ( .A(n16916), .B(n16917), .Z(n16915) );
  NAND U17175 ( .A(n16917), .B(n16916), .Z(n16912) );
  XOR U17176 ( .A(n395), .B(n394), .Z(\A1[176] ) );
  XOR U17177 ( .A(n16917), .B(n16918), .Z(n394) );
  XNOR U17178 ( .A(n16916), .B(n16914), .Z(n16918) );
  AND U17179 ( .A(n16919), .B(n16920), .Z(n16914) );
  NANDN U17180 ( .A(n16921), .B(n16922), .Z(n16920) );
  NANDN U17181 ( .A(n16923), .B(n16924), .Z(n16922) );
  NANDN U17182 ( .A(n16924), .B(n16923), .Z(n16919) );
  ANDN U17183 ( .B(B[163]), .A(n29), .Z(n16916) );
  XNOR U17184 ( .A(n16823), .B(n16925), .Z(n16917) );
  XNOR U17185 ( .A(n16822), .B(n16820), .Z(n16925) );
  AND U17186 ( .A(n16926), .B(n16927), .Z(n16820) );
  NANDN U17187 ( .A(n16928), .B(n16929), .Z(n16927) );
  OR U17188 ( .A(n16930), .B(n16931), .Z(n16929) );
  NAND U17189 ( .A(n16931), .B(n16930), .Z(n16926) );
  ANDN U17190 ( .B(B[164]), .A(n30), .Z(n16822) );
  XNOR U17191 ( .A(n16830), .B(n16932), .Z(n16823) );
  XNOR U17192 ( .A(n16829), .B(n16827), .Z(n16932) );
  AND U17193 ( .A(n16933), .B(n16934), .Z(n16827) );
  NANDN U17194 ( .A(n16935), .B(n16936), .Z(n16934) );
  NANDN U17195 ( .A(n16937), .B(n16938), .Z(n16936) );
  NANDN U17196 ( .A(n16938), .B(n16937), .Z(n16933) );
  ANDN U17197 ( .B(B[165]), .A(n31), .Z(n16829) );
  XNOR U17198 ( .A(n16837), .B(n16939), .Z(n16830) );
  XNOR U17199 ( .A(n16836), .B(n16834), .Z(n16939) );
  AND U17200 ( .A(n16940), .B(n16941), .Z(n16834) );
  NANDN U17201 ( .A(n16942), .B(n16943), .Z(n16941) );
  OR U17202 ( .A(n16944), .B(n16945), .Z(n16943) );
  NAND U17203 ( .A(n16945), .B(n16944), .Z(n16940) );
  ANDN U17204 ( .B(B[166]), .A(n32), .Z(n16836) );
  XNOR U17205 ( .A(n16844), .B(n16946), .Z(n16837) );
  XNOR U17206 ( .A(n16843), .B(n16841), .Z(n16946) );
  AND U17207 ( .A(n16947), .B(n16948), .Z(n16841) );
  NANDN U17208 ( .A(n16949), .B(n16950), .Z(n16948) );
  NANDN U17209 ( .A(n16951), .B(n16952), .Z(n16950) );
  NANDN U17210 ( .A(n16952), .B(n16951), .Z(n16947) );
  ANDN U17211 ( .B(B[167]), .A(n33), .Z(n16843) );
  XNOR U17212 ( .A(n16851), .B(n16953), .Z(n16844) );
  XNOR U17213 ( .A(n16850), .B(n16848), .Z(n16953) );
  AND U17214 ( .A(n16954), .B(n16955), .Z(n16848) );
  NANDN U17215 ( .A(n16956), .B(n16957), .Z(n16955) );
  OR U17216 ( .A(n16958), .B(n16959), .Z(n16957) );
  NAND U17217 ( .A(n16959), .B(n16958), .Z(n16954) );
  ANDN U17218 ( .B(B[168]), .A(n34), .Z(n16850) );
  XNOR U17219 ( .A(n16858), .B(n16960), .Z(n16851) );
  XNOR U17220 ( .A(n16857), .B(n16855), .Z(n16960) );
  AND U17221 ( .A(n16961), .B(n16962), .Z(n16855) );
  NANDN U17222 ( .A(n16963), .B(n16964), .Z(n16962) );
  NANDN U17223 ( .A(n16965), .B(n16966), .Z(n16964) );
  NANDN U17224 ( .A(n16966), .B(n16965), .Z(n16961) );
  ANDN U17225 ( .B(B[169]), .A(n35), .Z(n16857) );
  XNOR U17226 ( .A(n16865), .B(n16967), .Z(n16858) );
  XNOR U17227 ( .A(n16864), .B(n16862), .Z(n16967) );
  AND U17228 ( .A(n16968), .B(n16969), .Z(n16862) );
  NANDN U17229 ( .A(n16970), .B(n16971), .Z(n16969) );
  OR U17230 ( .A(n16972), .B(n16973), .Z(n16971) );
  NAND U17231 ( .A(n16973), .B(n16972), .Z(n16968) );
  ANDN U17232 ( .B(B[170]), .A(n36), .Z(n16864) );
  XNOR U17233 ( .A(n16872), .B(n16974), .Z(n16865) );
  XNOR U17234 ( .A(n16871), .B(n16869), .Z(n16974) );
  AND U17235 ( .A(n16975), .B(n16976), .Z(n16869) );
  NANDN U17236 ( .A(n16977), .B(n16978), .Z(n16976) );
  NANDN U17237 ( .A(n16979), .B(n16980), .Z(n16978) );
  NANDN U17238 ( .A(n16980), .B(n16979), .Z(n16975) );
  ANDN U17239 ( .B(B[171]), .A(n37), .Z(n16871) );
  XNOR U17240 ( .A(n16879), .B(n16981), .Z(n16872) );
  XNOR U17241 ( .A(n16878), .B(n16876), .Z(n16981) );
  AND U17242 ( .A(n16982), .B(n16983), .Z(n16876) );
  NANDN U17243 ( .A(n16984), .B(n16985), .Z(n16983) );
  OR U17244 ( .A(n16986), .B(n16987), .Z(n16985) );
  NAND U17245 ( .A(n16987), .B(n16986), .Z(n16982) );
  ANDN U17246 ( .B(B[172]), .A(n38), .Z(n16878) );
  XNOR U17247 ( .A(n16886), .B(n16988), .Z(n16879) );
  XNOR U17248 ( .A(n16885), .B(n16883), .Z(n16988) );
  AND U17249 ( .A(n16989), .B(n16990), .Z(n16883) );
  NANDN U17250 ( .A(n16991), .B(n16992), .Z(n16990) );
  NANDN U17251 ( .A(n16993), .B(n16994), .Z(n16992) );
  NANDN U17252 ( .A(n16994), .B(n16993), .Z(n16989) );
  ANDN U17253 ( .B(B[173]), .A(n39), .Z(n16885) );
  XNOR U17254 ( .A(n16893), .B(n16995), .Z(n16886) );
  XNOR U17255 ( .A(n16892), .B(n16890), .Z(n16995) );
  AND U17256 ( .A(n16996), .B(n16997), .Z(n16890) );
  NANDN U17257 ( .A(n16998), .B(n16999), .Z(n16997) );
  OR U17258 ( .A(n17000), .B(n17001), .Z(n16999) );
  NAND U17259 ( .A(n17001), .B(n17000), .Z(n16996) );
  ANDN U17260 ( .B(B[174]), .A(n40), .Z(n16892) );
  XNOR U17261 ( .A(n16900), .B(n17002), .Z(n16893) );
  XNOR U17262 ( .A(n16899), .B(n16897), .Z(n17002) );
  AND U17263 ( .A(n17003), .B(n17004), .Z(n16897) );
  NANDN U17264 ( .A(n17005), .B(n17006), .Z(n17004) );
  NAND U17265 ( .A(n17007), .B(n17008), .Z(n17006) );
  ANDN U17266 ( .B(B[175]), .A(n41), .Z(n16899) );
  XOR U17267 ( .A(n16906), .B(n17009), .Z(n16900) );
  XNOR U17268 ( .A(n16904), .B(n16907), .Z(n17009) );
  NAND U17269 ( .A(A[2]), .B(B[176]), .Z(n16907) );
  NANDN U17270 ( .A(n17010), .B(n17011), .Z(n16904) );
  AND U17271 ( .A(A[0]), .B(B[177]), .Z(n17011) );
  XNOR U17272 ( .A(n16909), .B(n17012), .Z(n16906) );
  NAND U17273 ( .A(A[0]), .B(B[178]), .Z(n17012) );
  NAND U17274 ( .A(B[177]), .B(A[1]), .Z(n16909) );
  NAND U17275 ( .A(n17013), .B(n17014), .Z(n395) );
  NANDN U17276 ( .A(n17015), .B(n17016), .Z(n17014) );
  OR U17277 ( .A(n17017), .B(n17018), .Z(n17016) );
  NAND U17278 ( .A(n17018), .B(n17017), .Z(n17013) );
  XOR U17279 ( .A(n397), .B(n396), .Z(\A1[175] ) );
  XOR U17280 ( .A(n17018), .B(n17019), .Z(n396) );
  XNOR U17281 ( .A(n17017), .B(n17015), .Z(n17019) );
  AND U17282 ( .A(n17020), .B(n17021), .Z(n17015) );
  NANDN U17283 ( .A(n17022), .B(n17023), .Z(n17021) );
  NANDN U17284 ( .A(n17024), .B(n17025), .Z(n17023) );
  NANDN U17285 ( .A(n17025), .B(n17024), .Z(n17020) );
  ANDN U17286 ( .B(B[162]), .A(n29), .Z(n17017) );
  XNOR U17287 ( .A(n16924), .B(n17026), .Z(n17018) );
  XNOR U17288 ( .A(n16923), .B(n16921), .Z(n17026) );
  AND U17289 ( .A(n17027), .B(n17028), .Z(n16921) );
  NANDN U17290 ( .A(n17029), .B(n17030), .Z(n17028) );
  OR U17291 ( .A(n17031), .B(n17032), .Z(n17030) );
  NAND U17292 ( .A(n17032), .B(n17031), .Z(n17027) );
  ANDN U17293 ( .B(B[163]), .A(n30), .Z(n16923) );
  XNOR U17294 ( .A(n16931), .B(n17033), .Z(n16924) );
  XNOR U17295 ( .A(n16930), .B(n16928), .Z(n17033) );
  AND U17296 ( .A(n17034), .B(n17035), .Z(n16928) );
  NANDN U17297 ( .A(n17036), .B(n17037), .Z(n17035) );
  NANDN U17298 ( .A(n17038), .B(n17039), .Z(n17037) );
  NANDN U17299 ( .A(n17039), .B(n17038), .Z(n17034) );
  ANDN U17300 ( .B(B[164]), .A(n31), .Z(n16930) );
  XNOR U17301 ( .A(n16938), .B(n17040), .Z(n16931) );
  XNOR U17302 ( .A(n16937), .B(n16935), .Z(n17040) );
  AND U17303 ( .A(n17041), .B(n17042), .Z(n16935) );
  NANDN U17304 ( .A(n17043), .B(n17044), .Z(n17042) );
  OR U17305 ( .A(n17045), .B(n17046), .Z(n17044) );
  NAND U17306 ( .A(n17046), .B(n17045), .Z(n17041) );
  ANDN U17307 ( .B(B[165]), .A(n32), .Z(n16937) );
  XNOR U17308 ( .A(n16945), .B(n17047), .Z(n16938) );
  XNOR U17309 ( .A(n16944), .B(n16942), .Z(n17047) );
  AND U17310 ( .A(n17048), .B(n17049), .Z(n16942) );
  NANDN U17311 ( .A(n17050), .B(n17051), .Z(n17049) );
  NANDN U17312 ( .A(n17052), .B(n17053), .Z(n17051) );
  NANDN U17313 ( .A(n17053), .B(n17052), .Z(n17048) );
  ANDN U17314 ( .B(B[166]), .A(n33), .Z(n16944) );
  XNOR U17315 ( .A(n16952), .B(n17054), .Z(n16945) );
  XNOR U17316 ( .A(n16951), .B(n16949), .Z(n17054) );
  AND U17317 ( .A(n17055), .B(n17056), .Z(n16949) );
  NANDN U17318 ( .A(n17057), .B(n17058), .Z(n17056) );
  OR U17319 ( .A(n17059), .B(n17060), .Z(n17058) );
  NAND U17320 ( .A(n17060), .B(n17059), .Z(n17055) );
  ANDN U17321 ( .B(B[167]), .A(n34), .Z(n16951) );
  XNOR U17322 ( .A(n16959), .B(n17061), .Z(n16952) );
  XNOR U17323 ( .A(n16958), .B(n16956), .Z(n17061) );
  AND U17324 ( .A(n17062), .B(n17063), .Z(n16956) );
  NANDN U17325 ( .A(n17064), .B(n17065), .Z(n17063) );
  NANDN U17326 ( .A(n17066), .B(n17067), .Z(n17065) );
  NANDN U17327 ( .A(n17067), .B(n17066), .Z(n17062) );
  ANDN U17328 ( .B(B[168]), .A(n35), .Z(n16958) );
  XNOR U17329 ( .A(n16966), .B(n17068), .Z(n16959) );
  XNOR U17330 ( .A(n16965), .B(n16963), .Z(n17068) );
  AND U17331 ( .A(n17069), .B(n17070), .Z(n16963) );
  NANDN U17332 ( .A(n17071), .B(n17072), .Z(n17070) );
  OR U17333 ( .A(n17073), .B(n17074), .Z(n17072) );
  NAND U17334 ( .A(n17074), .B(n17073), .Z(n17069) );
  ANDN U17335 ( .B(B[169]), .A(n36), .Z(n16965) );
  XNOR U17336 ( .A(n16973), .B(n17075), .Z(n16966) );
  XNOR U17337 ( .A(n16972), .B(n16970), .Z(n17075) );
  AND U17338 ( .A(n17076), .B(n17077), .Z(n16970) );
  NANDN U17339 ( .A(n17078), .B(n17079), .Z(n17077) );
  NANDN U17340 ( .A(n17080), .B(n17081), .Z(n17079) );
  NANDN U17341 ( .A(n17081), .B(n17080), .Z(n17076) );
  ANDN U17342 ( .B(B[170]), .A(n37), .Z(n16972) );
  XNOR U17343 ( .A(n16980), .B(n17082), .Z(n16973) );
  XNOR U17344 ( .A(n16979), .B(n16977), .Z(n17082) );
  AND U17345 ( .A(n17083), .B(n17084), .Z(n16977) );
  NANDN U17346 ( .A(n17085), .B(n17086), .Z(n17084) );
  OR U17347 ( .A(n17087), .B(n17088), .Z(n17086) );
  NAND U17348 ( .A(n17088), .B(n17087), .Z(n17083) );
  ANDN U17349 ( .B(B[171]), .A(n38), .Z(n16979) );
  XNOR U17350 ( .A(n16987), .B(n17089), .Z(n16980) );
  XNOR U17351 ( .A(n16986), .B(n16984), .Z(n17089) );
  AND U17352 ( .A(n17090), .B(n17091), .Z(n16984) );
  NANDN U17353 ( .A(n17092), .B(n17093), .Z(n17091) );
  NANDN U17354 ( .A(n17094), .B(n17095), .Z(n17093) );
  NANDN U17355 ( .A(n17095), .B(n17094), .Z(n17090) );
  ANDN U17356 ( .B(B[172]), .A(n39), .Z(n16986) );
  XNOR U17357 ( .A(n16994), .B(n17096), .Z(n16987) );
  XNOR U17358 ( .A(n16993), .B(n16991), .Z(n17096) );
  AND U17359 ( .A(n17097), .B(n17098), .Z(n16991) );
  NANDN U17360 ( .A(n17099), .B(n17100), .Z(n17098) );
  OR U17361 ( .A(n17101), .B(n17102), .Z(n17100) );
  NAND U17362 ( .A(n17102), .B(n17101), .Z(n17097) );
  ANDN U17363 ( .B(B[173]), .A(n40), .Z(n16993) );
  XNOR U17364 ( .A(n17001), .B(n17103), .Z(n16994) );
  XNOR U17365 ( .A(n17000), .B(n16998), .Z(n17103) );
  AND U17366 ( .A(n17104), .B(n17105), .Z(n16998) );
  NANDN U17367 ( .A(n17106), .B(n17107), .Z(n17105) );
  NAND U17368 ( .A(n17108), .B(n17109), .Z(n17107) );
  ANDN U17369 ( .B(B[174]), .A(n41), .Z(n17000) );
  XOR U17370 ( .A(n17007), .B(n17110), .Z(n17001) );
  XNOR U17371 ( .A(n17005), .B(n17008), .Z(n17110) );
  NAND U17372 ( .A(A[2]), .B(B[175]), .Z(n17008) );
  NANDN U17373 ( .A(n17111), .B(n17112), .Z(n17005) );
  AND U17374 ( .A(A[0]), .B(B[176]), .Z(n17112) );
  XNOR U17375 ( .A(n17010), .B(n17113), .Z(n17007) );
  NAND U17376 ( .A(A[0]), .B(B[177]), .Z(n17113) );
  NAND U17377 ( .A(B[176]), .B(A[1]), .Z(n17010) );
  NAND U17378 ( .A(n17114), .B(n17115), .Z(n397) );
  NANDN U17379 ( .A(n17116), .B(n17117), .Z(n17115) );
  OR U17380 ( .A(n17118), .B(n17119), .Z(n17117) );
  NAND U17381 ( .A(n17119), .B(n17118), .Z(n17114) );
  XOR U17382 ( .A(n399), .B(n398), .Z(\A1[174] ) );
  XOR U17383 ( .A(n17119), .B(n17120), .Z(n398) );
  XNOR U17384 ( .A(n17118), .B(n17116), .Z(n17120) );
  AND U17385 ( .A(n17121), .B(n17122), .Z(n17116) );
  NANDN U17386 ( .A(n17123), .B(n17124), .Z(n17122) );
  NANDN U17387 ( .A(n17125), .B(n17126), .Z(n17124) );
  NANDN U17388 ( .A(n17126), .B(n17125), .Z(n17121) );
  ANDN U17389 ( .B(B[161]), .A(n29), .Z(n17118) );
  XNOR U17390 ( .A(n17025), .B(n17127), .Z(n17119) );
  XNOR U17391 ( .A(n17024), .B(n17022), .Z(n17127) );
  AND U17392 ( .A(n17128), .B(n17129), .Z(n17022) );
  NANDN U17393 ( .A(n17130), .B(n17131), .Z(n17129) );
  OR U17394 ( .A(n17132), .B(n17133), .Z(n17131) );
  NAND U17395 ( .A(n17133), .B(n17132), .Z(n17128) );
  ANDN U17396 ( .B(B[162]), .A(n30), .Z(n17024) );
  XNOR U17397 ( .A(n17032), .B(n17134), .Z(n17025) );
  XNOR U17398 ( .A(n17031), .B(n17029), .Z(n17134) );
  AND U17399 ( .A(n17135), .B(n17136), .Z(n17029) );
  NANDN U17400 ( .A(n17137), .B(n17138), .Z(n17136) );
  NANDN U17401 ( .A(n17139), .B(n17140), .Z(n17138) );
  NANDN U17402 ( .A(n17140), .B(n17139), .Z(n17135) );
  ANDN U17403 ( .B(B[163]), .A(n31), .Z(n17031) );
  XNOR U17404 ( .A(n17039), .B(n17141), .Z(n17032) );
  XNOR U17405 ( .A(n17038), .B(n17036), .Z(n17141) );
  AND U17406 ( .A(n17142), .B(n17143), .Z(n17036) );
  NANDN U17407 ( .A(n17144), .B(n17145), .Z(n17143) );
  OR U17408 ( .A(n17146), .B(n17147), .Z(n17145) );
  NAND U17409 ( .A(n17147), .B(n17146), .Z(n17142) );
  ANDN U17410 ( .B(B[164]), .A(n32), .Z(n17038) );
  XNOR U17411 ( .A(n17046), .B(n17148), .Z(n17039) );
  XNOR U17412 ( .A(n17045), .B(n17043), .Z(n17148) );
  AND U17413 ( .A(n17149), .B(n17150), .Z(n17043) );
  NANDN U17414 ( .A(n17151), .B(n17152), .Z(n17150) );
  NANDN U17415 ( .A(n17153), .B(n17154), .Z(n17152) );
  NANDN U17416 ( .A(n17154), .B(n17153), .Z(n17149) );
  ANDN U17417 ( .B(B[165]), .A(n33), .Z(n17045) );
  XNOR U17418 ( .A(n17053), .B(n17155), .Z(n17046) );
  XNOR U17419 ( .A(n17052), .B(n17050), .Z(n17155) );
  AND U17420 ( .A(n17156), .B(n17157), .Z(n17050) );
  NANDN U17421 ( .A(n17158), .B(n17159), .Z(n17157) );
  OR U17422 ( .A(n17160), .B(n17161), .Z(n17159) );
  NAND U17423 ( .A(n17161), .B(n17160), .Z(n17156) );
  ANDN U17424 ( .B(B[166]), .A(n34), .Z(n17052) );
  XNOR U17425 ( .A(n17060), .B(n17162), .Z(n17053) );
  XNOR U17426 ( .A(n17059), .B(n17057), .Z(n17162) );
  AND U17427 ( .A(n17163), .B(n17164), .Z(n17057) );
  NANDN U17428 ( .A(n17165), .B(n17166), .Z(n17164) );
  NANDN U17429 ( .A(n17167), .B(n17168), .Z(n17166) );
  NANDN U17430 ( .A(n17168), .B(n17167), .Z(n17163) );
  ANDN U17431 ( .B(B[167]), .A(n35), .Z(n17059) );
  XNOR U17432 ( .A(n17067), .B(n17169), .Z(n17060) );
  XNOR U17433 ( .A(n17066), .B(n17064), .Z(n17169) );
  AND U17434 ( .A(n17170), .B(n17171), .Z(n17064) );
  NANDN U17435 ( .A(n17172), .B(n17173), .Z(n17171) );
  OR U17436 ( .A(n17174), .B(n17175), .Z(n17173) );
  NAND U17437 ( .A(n17175), .B(n17174), .Z(n17170) );
  ANDN U17438 ( .B(B[168]), .A(n36), .Z(n17066) );
  XNOR U17439 ( .A(n17074), .B(n17176), .Z(n17067) );
  XNOR U17440 ( .A(n17073), .B(n17071), .Z(n17176) );
  AND U17441 ( .A(n17177), .B(n17178), .Z(n17071) );
  NANDN U17442 ( .A(n17179), .B(n17180), .Z(n17178) );
  NANDN U17443 ( .A(n17181), .B(n17182), .Z(n17180) );
  NANDN U17444 ( .A(n17182), .B(n17181), .Z(n17177) );
  ANDN U17445 ( .B(B[169]), .A(n37), .Z(n17073) );
  XNOR U17446 ( .A(n17081), .B(n17183), .Z(n17074) );
  XNOR U17447 ( .A(n17080), .B(n17078), .Z(n17183) );
  AND U17448 ( .A(n17184), .B(n17185), .Z(n17078) );
  NANDN U17449 ( .A(n17186), .B(n17187), .Z(n17185) );
  OR U17450 ( .A(n17188), .B(n17189), .Z(n17187) );
  NAND U17451 ( .A(n17189), .B(n17188), .Z(n17184) );
  ANDN U17452 ( .B(B[170]), .A(n38), .Z(n17080) );
  XNOR U17453 ( .A(n17088), .B(n17190), .Z(n17081) );
  XNOR U17454 ( .A(n17087), .B(n17085), .Z(n17190) );
  AND U17455 ( .A(n17191), .B(n17192), .Z(n17085) );
  NANDN U17456 ( .A(n17193), .B(n17194), .Z(n17192) );
  NANDN U17457 ( .A(n17195), .B(n17196), .Z(n17194) );
  NANDN U17458 ( .A(n17196), .B(n17195), .Z(n17191) );
  ANDN U17459 ( .B(B[171]), .A(n39), .Z(n17087) );
  XNOR U17460 ( .A(n17095), .B(n17197), .Z(n17088) );
  XNOR U17461 ( .A(n17094), .B(n17092), .Z(n17197) );
  AND U17462 ( .A(n17198), .B(n17199), .Z(n17092) );
  NANDN U17463 ( .A(n17200), .B(n17201), .Z(n17199) );
  OR U17464 ( .A(n17202), .B(n17203), .Z(n17201) );
  NAND U17465 ( .A(n17203), .B(n17202), .Z(n17198) );
  ANDN U17466 ( .B(B[172]), .A(n40), .Z(n17094) );
  XNOR U17467 ( .A(n17102), .B(n17204), .Z(n17095) );
  XNOR U17468 ( .A(n17101), .B(n17099), .Z(n17204) );
  AND U17469 ( .A(n17205), .B(n17206), .Z(n17099) );
  NANDN U17470 ( .A(n17207), .B(n17208), .Z(n17206) );
  NAND U17471 ( .A(n17209), .B(n17210), .Z(n17208) );
  ANDN U17472 ( .B(B[173]), .A(n41), .Z(n17101) );
  XOR U17473 ( .A(n17108), .B(n17211), .Z(n17102) );
  XNOR U17474 ( .A(n17106), .B(n17109), .Z(n17211) );
  NAND U17475 ( .A(A[2]), .B(B[174]), .Z(n17109) );
  NANDN U17476 ( .A(n17212), .B(n17213), .Z(n17106) );
  AND U17477 ( .A(A[0]), .B(B[175]), .Z(n17213) );
  XNOR U17478 ( .A(n17111), .B(n17214), .Z(n17108) );
  NAND U17479 ( .A(A[0]), .B(B[176]), .Z(n17214) );
  NAND U17480 ( .A(B[175]), .B(A[1]), .Z(n17111) );
  NAND U17481 ( .A(n17215), .B(n17216), .Z(n399) );
  NANDN U17482 ( .A(n17217), .B(n17218), .Z(n17216) );
  OR U17483 ( .A(n17219), .B(n17220), .Z(n17218) );
  NAND U17484 ( .A(n17220), .B(n17219), .Z(n17215) );
  XOR U17485 ( .A(n401), .B(n400), .Z(\A1[173] ) );
  XOR U17486 ( .A(n17220), .B(n17221), .Z(n400) );
  XNOR U17487 ( .A(n17219), .B(n17217), .Z(n17221) );
  AND U17488 ( .A(n17222), .B(n17223), .Z(n17217) );
  NANDN U17489 ( .A(n17224), .B(n17225), .Z(n17223) );
  NANDN U17490 ( .A(n17226), .B(n17227), .Z(n17225) );
  NANDN U17491 ( .A(n17227), .B(n17226), .Z(n17222) );
  ANDN U17492 ( .B(B[160]), .A(n29), .Z(n17219) );
  XNOR U17493 ( .A(n17126), .B(n17228), .Z(n17220) );
  XNOR U17494 ( .A(n17125), .B(n17123), .Z(n17228) );
  AND U17495 ( .A(n17229), .B(n17230), .Z(n17123) );
  NANDN U17496 ( .A(n17231), .B(n17232), .Z(n17230) );
  OR U17497 ( .A(n17233), .B(n17234), .Z(n17232) );
  NAND U17498 ( .A(n17234), .B(n17233), .Z(n17229) );
  ANDN U17499 ( .B(B[161]), .A(n30), .Z(n17125) );
  XNOR U17500 ( .A(n17133), .B(n17235), .Z(n17126) );
  XNOR U17501 ( .A(n17132), .B(n17130), .Z(n17235) );
  AND U17502 ( .A(n17236), .B(n17237), .Z(n17130) );
  NANDN U17503 ( .A(n17238), .B(n17239), .Z(n17237) );
  NANDN U17504 ( .A(n17240), .B(n17241), .Z(n17239) );
  NANDN U17505 ( .A(n17241), .B(n17240), .Z(n17236) );
  ANDN U17506 ( .B(B[162]), .A(n31), .Z(n17132) );
  XNOR U17507 ( .A(n17140), .B(n17242), .Z(n17133) );
  XNOR U17508 ( .A(n17139), .B(n17137), .Z(n17242) );
  AND U17509 ( .A(n17243), .B(n17244), .Z(n17137) );
  NANDN U17510 ( .A(n17245), .B(n17246), .Z(n17244) );
  OR U17511 ( .A(n17247), .B(n17248), .Z(n17246) );
  NAND U17512 ( .A(n17248), .B(n17247), .Z(n17243) );
  ANDN U17513 ( .B(B[163]), .A(n32), .Z(n17139) );
  XNOR U17514 ( .A(n17147), .B(n17249), .Z(n17140) );
  XNOR U17515 ( .A(n17146), .B(n17144), .Z(n17249) );
  AND U17516 ( .A(n17250), .B(n17251), .Z(n17144) );
  NANDN U17517 ( .A(n17252), .B(n17253), .Z(n17251) );
  NANDN U17518 ( .A(n17254), .B(n17255), .Z(n17253) );
  NANDN U17519 ( .A(n17255), .B(n17254), .Z(n17250) );
  ANDN U17520 ( .B(B[164]), .A(n33), .Z(n17146) );
  XNOR U17521 ( .A(n17154), .B(n17256), .Z(n17147) );
  XNOR U17522 ( .A(n17153), .B(n17151), .Z(n17256) );
  AND U17523 ( .A(n17257), .B(n17258), .Z(n17151) );
  NANDN U17524 ( .A(n17259), .B(n17260), .Z(n17258) );
  OR U17525 ( .A(n17261), .B(n17262), .Z(n17260) );
  NAND U17526 ( .A(n17262), .B(n17261), .Z(n17257) );
  ANDN U17527 ( .B(B[165]), .A(n34), .Z(n17153) );
  XNOR U17528 ( .A(n17161), .B(n17263), .Z(n17154) );
  XNOR U17529 ( .A(n17160), .B(n17158), .Z(n17263) );
  AND U17530 ( .A(n17264), .B(n17265), .Z(n17158) );
  NANDN U17531 ( .A(n17266), .B(n17267), .Z(n17265) );
  NANDN U17532 ( .A(n17268), .B(n17269), .Z(n17267) );
  NANDN U17533 ( .A(n17269), .B(n17268), .Z(n17264) );
  ANDN U17534 ( .B(B[166]), .A(n35), .Z(n17160) );
  XNOR U17535 ( .A(n17168), .B(n17270), .Z(n17161) );
  XNOR U17536 ( .A(n17167), .B(n17165), .Z(n17270) );
  AND U17537 ( .A(n17271), .B(n17272), .Z(n17165) );
  NANDN U17538 ( .A(n17273), .B(n17274), .Z(n17272) );
  OR U17539 ( .A(n17275), .B(n17276), .Z(n17274) );
  NAND U17540 ( .A(n17276), .B(n17275), .Z(n17271) );
  ANDN U17541 ( .B(B[167]), .A(n36), .Z(n17167) );
  XNOR U17542 ( .A(n17175), .B(n17277), .Z(n17168) );
  XNOR U17543 ( .A(n17174), .B(n17172), .Z(n17277) );
  AND U17544 ( .A(n17278), .B(n17279), .Z(n17172) );
  NANDN U17545 ( .A(n17280), .B(n17281), .Z(n17279) );
  NANDN U17546 ( .A(n17282), .B(n17283), .Z(n17281) );
  NANDN U17547 ( .A(n17283), .B(n17282), .Z(n17278) );
  ANDN U17548 ( .B(B[168]), .A(n37), .Z(n17174) );
  XNOR U17549 ( .A(n17182), .B(n17284), .Z(n17175) );
  XNOR U17550 ( .A(n17181), .B(n17179), .Z(n17284) );
  AND U17551 ( .A(n17285), .B(n17286), .Z(n17179) );
  NANDN U17552 ( .A(n17287), .B(n17288), .Z(n17286) );
  OR U17553 ( .A(n17289), .B(n17290), .Z(n17288) );
  NAND U17554 ( .A(n17290), .B(n17289), .Z(n17285) );
  ANDN U17555 ( .B(B[169]), .A(n38), .Z(n17181) );
  XNOR U17556 ( .A(n17189), .B(n17291), .Z(n17182) );
  XNOR U17557 ( .A(n17188), .B(n17186), .Z(n17291) );
  AND U17558 ( .A(n17292), .B(n17293), .Z(n17186) );
  NANDN U17559 ( .A(n17294), .B(n17295), .Z(n17293) );
  NANDN U17560 ( .A(n17296), .B(n17297), .Z(n17295) );
  NANDN U17561 ( .A(n17297), .B(n17296), .Z(n17292) );
  ANDN U17562 ( .B(B[170]), .A(n39), .Z(n17188) );
  XNOR U17563 ( .A(n17196), .B(n17298), .Z(n17189) );
  XNOR U17564 ( .A(n17195), .B(n17193), .Z(n17298) );
  AND U17565 ( .A(n17299), .B(n17300), .Z(n17193) );
  NANDN U17566 ( .A(n17301), .B(n17302), .Z(n17300) );
  OR U17567 ( .A(n17303), .B(n17304), .Z(n17302) );
  NAND U17568 ( .A(n17304), .B(n17303), .Z(n17299) );
  ANDN U17569 ( .B(B[171]), .A(n40), .Z(n17195) );
  XNOR U17570 ( .A(n17203), .B(n17305), .Z(n17196) );
  XNOR U17571 ( .A(n17202), .B(n17200), .Z(n17305) );
  AND U17572 ( .A(n17306), .B(n17307), .Z(n17200) );
  NANDN U17573 ( .A(n17308), .B(n17309), .Z(n17307) );
  NAND U17574 ( .A(n17310), .B(n17311), .Z(n17309) );
  ANDN U17575 ( .B(B[172]), .A(n41), .Z(n17202) );
  XOR U17576 ( .A(n17209), .B(n17312), .Z(n17203) );
  XNOR U17577 ( .A(n17207), .B(n17210), .Z(n17312) );
  NAND U17578 ( .A(A[2]), .B(B[173]), .Z(n17210) );
  NANDN U17579 ( .A(n17313), .B(n17314), .Z(n17207) );
  AND U17580 ( .A(A[0]), .B(B[174]), .Z(n17314) );
  XNOR U17581 ( .A(n17212), .B(n17315), .Z(n17209) );
  NAND U17582 ( .A(A[0]), .B(B[175]), .Z(n17315) );
  NAND U17583 ( .A(B[174]), .B(A[1]), .Z(n17212) );
  NAND U17584 ( .A(n17316), .B(n17317), .Z(n401) );
  NANDN U17585 ( .A(n17318), .B(n17319), .Z(n17317) );
  OR U17586 ( .A(n17320), .B(n17321), .Z(n17319) );
  NAND U17587 ( .A(n17321), .B(n17320), .Z(n17316) );
  XOR U17588 ( .A(n403), .B(n402), .Z(\A1[172] ) );
  XOR U17589 ( .A(n17321), .B(n17322), .Z(n402) );
  XNOR U17590 ( .A(n17320), .B(n17318), .Z(n17322) );
  AND U17591 ( .A(n17323), .B(n17324), .Z(n17318) );
  NANDN U17592 ( .A(n17325), .B(n17326), .Z(n17324) );
  NANDN U17593 ( .A(n17327), .B(n17328), .Z(n17326) );
  NANDN U17594 ( .A(n17328), .B(n17327), .Z(n17323) );
  ANDN U17595 ( .B(B[159]), .A(n29), .Z(n17320) );
  XNOR U17596 ( .A(n17227), .B(n17329), .Z(n17321) );
  XNOR U17597 ( .A(n17226), .B(n17224), .Z(n17329) );
  AND U17598 ( .A(n17330), .B(n17331), .Z(n17224) );
  NANDN U17599 ( .A(n17332), .B(n17333), .Z(n17331) );
  OR U17600 ( .A(n17334), .B(n17335), .Z(n17333) );
  NAND U17601 ( .A(n17335), .B(n17334), .Z(n17330) );
  ANDN U17602 ( .B(B[160]), .A(n30), .Z(n17226) );
  XNOR U17603 ( .A(n17234), .B(n17336), .Z(n17227) );
  XNOR U17604 ( .A(n17233), .B(n17231), .Z(n17336) );
  AND U17605 ( .A(n17337), .B(n17338), .Z(n17231) );
  NANDN U17606 ( .A(n17339), .B(n17340), .Z(n17338) );
  NANDN U17607 ( .A(n17341), .B(n17342), .Z(n17340) );
  NANDN U17608 ( .A(n17342), .B(n17341), .Z(n17337) );
  ANDN U17609 ( .B(B[161]), .A(n31), .Z(n17233) );
  XNOR U17610 ( .A(n17241), .B(n17343), .Z(n17234) );
  XNOR U17611 ( .A(n17240), .B(n17238), .Z(n17343) );
  AND U17612 ( .A(n17344), .B(n17345), .Z(n17238) );
  NANDN U17613 ( .A(n17346), .B(n17347), .Z(n17345) );
  OR U17614 ( .A(n17348), .B(n17349), .Z(n17347) );
  NAND U17615 ( .A(n17349), .B(n17348), .Z(n17344) );
  ANDN U17616 ( .B(B[162]), .A(n32), .Z(n17240) );
  XNOR U17617 ( .A(n17248), .B(n17350), .Z(n17241) );
  XNOR U17618 ( .A(n17247), .B(n17245), .Z(n17350) );
  AND U17619 ( .A(n17351), .B(n17352), .Z(n17245) );
  NANDN U17620 ( .A(n17353), .B(n17354), .Z(n17352) );
  NANDN U17621 ( .A(n17355), .B(n17356), .Z(n17354) );
  NANDN U17622 ( .A(n17356), .B(n17355), .Z(n17351) );
  ANDN U17623 ( .B(B[163]), .A(n33), .Z(n17247) );
  XNOR U17624 ( .A(n17255), .B(n17357), .Z(n17248) );
  XNOR U17625 ( .A(n17254), .B(n17252), .Z(n17357) );
  AND U17626 ( .A(n17358), .B(n17359), .Z(n17252) );
  NANDN U17627 ( .A(n17360), .B(n17361), .Z(n17359) );
  OR U17628 ( .A(n17362), .B(n17363), .Z(n17361) );
  NAND U17629 ( .A(n17363), .B(n17362), .Z(n17358) );
  ANDN U17630 ( .B(B[164]), .A(n34), .Z(n17254) );
  XNOR U17631 ( .A(n17262), .B(n17364), .Z(n17255) );
  XNOR U17632 ( .A(n17261), .B(n17259), .Z(n17364) );
  AND U17633 ( .A(n17365), .B(n17366), .Z(n17259) );
  NANDN U17634 ( .A(n17367), .B(n17368), .Z(n17366) );
  NANDN U17635 ( .A(n17369), .B(n17370), .Z(n17368) );
  NANDN U17636 ( .A(n17370), .B(n17369), .Z(n17365) );
  ANDN U17637 ( .B(B[165]), .A(n35), .Z(n17261) );
  XNOR U17638 ( .A(n17269), .B(n17371), .Z(n17262) );
  XNOR U17639 ( .A(n17268), .B(n17266), .Z(n17371) );
  AND U17640 ( .A(n17372), .B(n17373), .Z(n17266) );
  NANDN U17641 ( .A(n17374), .B(n17375), .Z(n17373) );
  OR U17642 ( .A(n17376), .B(n17377), .Z(n17375) );
  NAND U17643 ( .A(n17377), .B(n17376), .Z(n17372) );
  ANDN U17644 ( .B(B[166]), .A(n36), .Z(n17268) );
  XNOR U17645 ( .A(n17276), .B(n17378), .Z(n17269) );
  XNOR U17646 ( .A(n17275), .B(n17273), .Z(n17378) );
  AND U17647 ( .A(n17379), .B(n17380), .Z(n17273) );
  NANDN U17648 ( .A(n17381), .B(n17382), .Z(n17380) );
  NANDN U17649 ( .A(n17383), .B(n17384), .Z(n17382) );
  NANDN U17650 ( .A(n17384), .B(n17383), .Z(n17379) );
  ANDN U17651 ( .B(B[167]), .A(n37), .Z(n17275) );
  XNOR U17652 ( .A(n17283), .B(n17385), .Z(n17276) );
  XNOR U17653 ( .A(n17282), .B(n17280), .Z(n17385) );
  AND U17654 ( .A(n17386), .B(n17387), .Z(n17280) );
  NANDN U17655 ( .A(n17388), .B(n17389), .Z(n17387) );
  OR U17656 ( .A(n17390), .B(n17391), .Z(n17389) );
  NAND U17657 ( .A(n17391), .B(n17390), .Z(n17386) );
  ANDN U17658 ( .B(B[168]), .A(n38), .Z(n17282) );
  XNOR U17659 ( .A(n17290), .B(n17392), .Z(n17283) );
  XNOR U17660 ( .A(n17289), .B(n17287), .Z(n17392) );
  AND U17661 ( .A(n17393), .B(n17394), .Z(n17287) );
  NANDN U17662 ( .A(n17395), .B(n17396), .Z(n17394) );
  NANDN U17663 ( .A(n17397), .B(n17398), .Z(n17396) );
  NANDN U17664 ( .A(n17398), .B(n17397), .Z(n17393) );
  ANDN U17665 ( .B(B[169]), .A(n39), .Z(n17289) );
  XNOR U17666 ( .A(n17297), .B(n17399), .Z(n17290) );
  XNOR U17667 ( .A(n17296), .B(n17294), .Z(n17399) );
  AND U17668 ( .A(n17400), .B(n17401), .Z(n17294) );
  NANDN U17669 ( .A(n17402), .B(n17403), .Z(n17401) );
  OR U17670 ( .A(n17404), .B(n17405), .Z(n17403) );
  NAND U17671 ( .A(n17405), .B(n17404), .Z(n17400) );
  ANDN U17672 ( .B(B[170]), .A(n40), .Z(n17296) );
  XNOR U17673 ( .A(n17304), .B(n17406), .Z(n17297) );
  XNOR U17674 ( .A(n17303), .B(n17301), .Z(n17406) );
  AND U17675 ( .A(n17407), .B(n17408), .Z(n17301) );
  NANDN U17676 ( .A(n17409), .B(n17410), .Z(n17408) );
  NAND U17677 ( .A(n17411), .B(n17412), .Z(n17410) );
  ANDN U17678 ( .B(B[171]), .A(n41), .Z(n17303) );
  XOR U17679 ( .A(n17310), .B(n17413), .Z(n17304) );
  XNOR U17680 ( .A(n17308), .B(n17311), .Z(n17413) );
  NAND U17681 ( .A(A[2]), .B(B[172]), .Z(n17311) );
  NANDN U17682 ( .A(n17414), .B(n17415), .Z(n17308) );
  AND U17683 ( .A(A[0]), .B(B[173]), .Z(n17415) );
  XNOR U17684 ( .A(n17313), .B(n17416), .Z(n17310) );
  NAND U17685 ( .A(A[0]), .B(B[174]), .Z(n17416) );
  NAND U17686 ( .A(B[173]), .B(A[1]), .Z(n17313) );
  NAND U17687 ( .A(n17417), .B(n17418), .Z(n403) );
  NANDN U17688 ( .A(n17419), .B(n17420), .Z(n17418) );
  OR U17689 ( .A(n17421), .B(n17422), .Z(n17420) );
  NAND U17690 ( .A(n17422), .B(n17421), .Z(n17417) );
  XOR U17691 ( .A(n405), .B(n404), .Z(\A1[171] ) );
  XOR U17692 ( .A(n17422), .B(n17423), .Z(n404) );
  XNOR U17693 ( .A(n17421), .B(n17419), .Z(n17423) );
  AND U17694 ( .A(n17424), .B(n17425), .Z(n17419) );
  NANDN U17695 ( .A(n17426), .B(n17427), .Z(n17425) );
  NANDN U17696 ( .A(n17428), .B(n17429), .Z(n17427) );
  NANDN U17697 ( .A(n17429), .B(n17428), .Z(n17424) );
  ANDN U17698 ( .B(B[158]), .A(n29), .Z(n17421) );
  XNOR U17699 ( .A(n17328), .B(n17430), .Z(n17422) );
  XNOR U17700 ( .A(n17327), .B(n17325), .Z(n17430) );
  AND U17701 ( .A(n17431), .B(n17432), .Z(n17325) );
  NANDN U17702 ( .A(n17433), .B(n17434), .Z(n17432) );
  OR U17703 ( .A(n17435), .B(n17436), .Z(n17434) );
  NAND U17704 ( .A(n17436), .B(n17435), .Z(n17431) );
  ANDN U17705 ( .B(B[159]), .A(n30), .Z(n17327) );
  XNOR U17706 ( .A(n17335), .B(n17437), .Z(n17328) );
  XNOR U17707 ( .A(n17334), .B(n17332), .Z(n17437) );
  AND U17708 ( .A(n17438), .B(n17439), .Z(n17332) );
  NANDN U17709 ( .A(n17440), .B(n17441), .Z(n17439) );
  NANDN U17710 ( .A(n17442), .B(n17443), .Z(n17441) );
  NANDN U17711 ( .A(n17443), .B(n17442), .Z(n17438) );
  ANDN U17712 ( .B(B[160]), .A(n31), .Z(n17334) );
  XNOR U17713 ( .A(n17342), .B(n17444), .Z(n17335) );
  XNOR U17714 ( .A(n17341), .B(n17339), .Z(n17444) );
  AND U17715 ( .A(n17445), .B(n17446), .Z(n17339) );
  NANDN U17716 ( .A(n17447), .B(n17448), .Z(n17446) );
  OR U17717 ( .A(n17449), .B(n17450), .Z(n17448) );
  NAND U17718 ( .A(n17450), .B(n17449), .Z(n17445) );
  ANDN U17719 ( .B(B[161]), .A(n32), .Z(n17341) );
  XNOR U17720 ( .A(n17349), .B(n17451), .Z(n17342) );
  XNOR U17721 ( .A(n17348), .B(n17346), .Z(n17451) );
  AND U17722 ( .A(n17452), .B(n17453), .Z(n17346) );
  NANDN U17723 ( .A(n17454), .B(n17455), .Z(n17453) );
  NANDN U17724 ( .A(n17456), .B(n17457), .Z(n17455) );
  NANDN U17725 ( .A(n17457), .B(n17456), .Z(n17452) );
  ANDN U17726 ( .B(B[162]), .A(n33), .Z(n17348) );
  XNOR U17727 ( .A(n17356), .B(n17458), .Z(n17349) );
  XNOR U17728 ( .A(n17355), .B(n17353), .Z(n17458) );
  AND U17729 ( .A(n17459), .B(n17460), .Z(n17353) );
  NANDN U17730 ( .A(n17461), .B(n17462), .Z(n17460) );
  OR U17731 ( .A(n17463), .B(n17464), .Z(n17462) );
  NAND U17732 ( .A(n17464), .B(n17463), .Z(n17459) );
  ANDN U17733 ( .B(B[163]), .A(n34), .Z(n17355) );
  XNOR U17734 ( .A(n17363), .B(n17465), .Z(n17356) );
  XNOR U17735 ( .A(n17362), .B(n17360), .Z(n17465) );
  AND U17736 ( .A(n17466), .B(n17467), .Z(n17360) );
  NANDN U17737 ( .A(n17468), .B(n17469), .Z(n17467) );
  NANDN U17738 ( .A(n17470), .B(n17471), .Z(n17469) );
  NANDN U17739 ( .A(n17471), .B(n17470), .Z(n17466) );
  ANDN U17740 ( .B(B[164]), .A(n35), .Z(n17362) );
  XNOR U17741 ( .A(n17370), .B(n17472), .Z(n17363) );
  XNOR U17742 ( .A(n17369), .B(n17367), .Z(n17472) );
  AND U17743 ( .A(n17473), .B(n17474), .Z(n17367) );
  NANDN U17744 ( .A(n17475), .B(n17476), .Z(n17474) );
  OR U17745 ( .A(n17477), .B(n17478), .Z(n17476) );
  NAND U17746 ( .A(n17478), .B(n17477), .Z(n17473) );
  ANDN U17747 ( .B(B[165]), .A(n36), .Z(n17369) );
  XNOR U17748 ( .A(n17377), .B(n17479), .Z(n17370) );
  XNOR U17749 ( .A(n17376), .B(n17374), .Z(n17479) );
  AND U17750 ( .A(n17480), .B(n17481), .Z(n17374) );
  NANDN U17751 ( .A(n17482), .B(n17483), .Z(n17481) );
  NANDN U17752 ( .A(n17484), .B(n17485), .Z(n17483) );
  NANDN U17753 ( .A(n17485), .B(n17484), .Z(n17480) );
  ANDN U17754 ( .B(B[166]), .A(n37), .Z(n17376) );
  XNOR U17755 ( .A(n17384), .B(n17486), .Z(n17377) );
  XNOR U17756 ( .A(n17383), .B(n17381), .Z(n17486) );
  AND U17757 ( .A(n17487), .B(n17488), .Z(n17381) );
  NANDN U17758 ( .A(n17489), .B(n17490), .Z(n17488) );
  OR U17759 ( .A(n17491), .B(n17492), .Z(n17490) );
  NAND U17760 ( .A(n17492), .B(n17491), .Z(n17487) );
  ANDN U17761 ( .B(B[167]), .A(n38), .Z(n17383) );
  XNOR U17762 ( .A(n17391), .B(n17493), .Z(n17384) );
  XNOR U17763 ( .A(n17390), .B(n17388), .Z(n17493) );
  AND U17764 ( .A(n17494), .B(n17495), .Z(n17388) );
  NANDN U17765 ( .A(n17496), .B(n17497), .Z(n17495) );
  NANDN U17766 ( .A(n17498), .B(n17499), .Z(n17497) );
  NANDN U17767 ( .A(n17499), .B(n17498), .Z(n17494) );
  ANDN U17768 ( .B(B[168]), .A(n39), .Z(n17390) );
  XNOR U17769 ( .A(n17398), .B(n17500), .Z(n17391) );
  XNOR U17770 ( .A(n17397), .B(n17395), .Z(n17500) );
  AND U17771 ( .A(n17501), .B(n17502), .Z(n17395) );
  NANDN U17772 ( .A(n17503), .B(n17504), .Z(n17502) );
  OR U17773 ( .A(n17505), .B(n17506), .Z(n17504) );
  NAND U17774 ( .A(n17506), .B(n17505), .Z(n17501) );
  ANDN U17775 ( .B(B[169]), .A(n40), .Z(n17397) );
  XNOR U17776 ( .A(n17405), .B(n17507), .Z(n17398) );
  XNOR U17777 ( .A(n17404), .B(n17402), .Z(n17507) );
  AND U17778 ( .A(n17508), .B(n17509), .Z(n17402) );
  NANDN U17779 ( .A(n17510), .B(n17511), .Z(n17509) );
  NAND U17780 ( .A(n17512), .B(n17513), .Z(n17511) );
  ANDN U17781 ( .B(B[170]), .A(n41), .Z(n17404) );
  XOR U17782 ( .A(n17411), .B(n17514), .Z(n17405) );
  XNOR U17783 ( .A(n17409), .B(n17412), .Z(n17514) );
  NAND U17784 ( .A(A[2]), .B(B[171]), .Z(n17412) );
  NANDN U17785 ( .A(n17515), .B(n17516), .Z(n17409) );
  AND U17786 ( .A(A[0]), .B(B[172]), .Z(n17516) );
  XNOR U17787 ( .A(n17414), .B(n17517), .Z(n17411) );
  NAND U17788 ( .A(A[0]), .B(B[173]), .Z(n17517) );
  NAND U17789 ( .A(B[172]), .B(A[1]), .Z(n17414) );
  NAND U17790 ( .A(n17518), .B(n17519), .Z(n405) );
  NANDN U17791 ( .A(n17520), .B(n17521), .Z(n17519) );
  OR U17792 ( .A(n17522), .B(n17523), .Z(n17521) );
  NAND U17793 ( .A(n17523), .B(n17522), .Z(n17518) );
  XOR U17794 ( .A(n407), .B(n406), .Z(\A1[170] ) );
  XOR U17795 ( .A(n17523), .B(n17524), .Z(n406) );
  XNOR U17796 ( .A(n17522), .B(n17520), .Z(n17524) );
  AND U17797 ( .A(n17525), .B(n17526), .Z(n17520) );
  NANDN U17798 ( .A(n17527), .B(n17528), .Z(n17526) );
  NANDN U17799 ( .A(n17529), .B(n17530), .Z(n17528) );
  NANDN U17800 ( .A(n17530), .B(n17529), .Z(n17525) );
  ANDN U17801 ( .B(B[157]), .A(n29), .Z(n17522) );
  XNOR U17802 ( .A(n17429), .B(n17531), .Z(n17523) );
  XNOR U17803 ( .A(n17428), .B(n17426), .Z(n17531) );
  AND U17804 ( .A(n17532), .B(n17533), .Z(n17426) );
  NANDN U17805 ( .A(n17534), .B(n17535), .Z(n17533) );
  OR U17806 ( .A(n17536), .B(n17537), .Z(n17535) );
  NAND U17807 ( .A(n17537), .B(n17536), .Z(n17532) );
  ANDN U17808 ( .B(B[158]), .A(n30), .Z(n17428) );
  XNOR U17809 ( .A(n17436), .B(n17538), .Z(n17429) );
  XNOR U17810 ( .A(n17435), .B(n17433), .Z(n17538) );
  AND U17811 ( .A(n17539), .B(n17540), .Z(n17433) );
  NANDN U17812 ( .A(n17541), .B(n17542), .Z(n17540) );
  NANDN U17813 ( .A(n17543), .B(n17544), .Z(n17542) );
  NANDN U17814 ( .A(n17544), .B(n17543), .Z(n17539) );
  ANDN U17815 ( .B(B[159]), .A(n31), .Z(n17435) );
  XNOR U17816 ( .A(n17443), .B(n17545), .Z(n17436) );
  XNOR U17817 ( .A(n17442), .B(n17440), .Z(n17545) );
  AND U17818 ( .A(n17546), .B(n17547), .Z(n17440) );
  NANDN U17819 ( .A(n17548), .B(n17549), .Z(n17547) );
  OR U17820 ( .A(n17550), .B(n17551), .Z(n17549) );
  NAND U17821 ( .A(n17551), .B(n17550), .Z(n17546) );
  ANDN U17822 ( .B(B[160]), .A(n32), .Z(n17442) );
  XNOR U17823 ( .A(n17450), .B(n17552), .Z(n17443) );
  XNOR U17824 ( .A(n17449), .B(n17447), .Z(n17552) );
  AND U17825 ( .A(n17553), .B(n17554), .Z(n17447) );
  NANDN U17826 ( .A(n17555), .B(n17556), .Z(n17554) );
  NANDN U17827 ( .A(n17557), .B(n17558), .Z(n17556) );
  NANDN U17828 ( .A(n17558), .B(n17557), .Z(n17553) );
  ANDN U17829 ( .B(B[161]), .A(n33), .Z(n17449) );
  XNOR U17830 ( .A(n17457), .B(n17559), .Z(n17450) );
  XNOR U17831 ( .A(n17456), .B(n17454), .Z(n17559) );
  AND U17832 ( .A(n17560), .B(n17561), .Z(n17454) );
  NANDN U17833 ( .A(n17562), .B(n17563), .Z(n17561) );
  OR U17834 ( .A(n17564), .B(n17565), .Z(n17563) );
  NAND U17835 ( .A(n17565), .B(n17564), .Z(n17560) );
  ANDN U17836 ( .B(B[162]), .A(n34), .Z(n17456) );
  XNOR U17837 ( .A(n17464), .B(n17566), .Z(n17457) );
  XNOR U17838 ( .A(n17463), .B(n17461), .Z(n17566) );
  AND U17839 ( .A(n17567), .B(n17568), .Z(n17461) );
  NANDN U17840 ( .A(n17569), .B(n17570), .Z(n17568) );
  NANDN U17841 ( .A(n17571), .B(n17572), .Z(n17570) );
  NANDN U17842 ( .A(n17572), .B(n17571), .Z(n17567) );
  ANDN U17843 ( .B(B[163]), .A(n35), .Z(n17463) );
  XNOR U17844 ( .A(n17471), .B(n17573), .Z(n17464) );
  XNOR U17845 ( .A(n17470), .B(n17468), .Z(n17573) );
  AND U17846 ( .A(n17574), .B(n17575), .Z(n17468) );
  NANDN U17847 ( .A(n17576), .B(n17577), .Z(n17575) );
  OR U17848 ( .A(n17578), .B(n17579), .Z(n17577) );
  NAND U17849 ( .A(n17579), .B(n17578), .Z(n17574) );
  ANDN U17850 ( .B(B[164]), .A(n36), .Z(n17470) );
  XNOR U17851 ( .A(n17478), .B(n17580), .Z(n17471) );
  XNOR U17852 ( .A(n17477), .B(n17475), .Z(n17580) );
  AND U17853 ( .A(n17581), .B(n17582), .Z(n17475) );
  NANDN U17854 ( .A(n17583), .B(n17584), .Z(n17582) );
  NANDN U17855 ( .A(n17585), .B(n17586), .Z(n17584) );
  NANDN U17856 ( .A(n17586), .B(n17585), .Z(n17581) );
  ANDN U17857 ( .B(B[165]), .A(n37), .Z(n17477) );
  XNOR U17858 ( .A(n17485), .B(n17587), .Z(n17478) );
  XNOR U17859 ( .A(n17484), .B(n17482), .Z(n17587) );
  AND U17860 ( .A(n17588), .B(n17589), .Z(n17482) );
  NANDN U17861 ( .A(n17590), .B(n17591), .Z(n17589) );
  OR U17862 ( .A(n17592), .B(n17593), .Z(n17591) );
  NAND U17863 ( .A(n17593), .B(n17592), .Z(n17588) );
  ANDN U17864 ( .B(B[166]), .A(n38), .Z(n17484) );
  XNOR U17865 ( .A(n17492), .B(n17594), .Z(n17485) );
  XNOR U17866 ( .A(n17491), .B(n17489), .Z(n17594) );
  AND U17867 ( .A(n17595), .B(n17596), .Z(n17489) );
  NANDN U17868 ( .A(n17597), .B(n17598), .Z(n17596) );
  NANDN U17869 ( .A(n17599), .B(n17600), .Z(n17598) );
  NANDN U17870 ( .A(n17600), .B(n17599), .Z(n17595) );
  ANDN U17871 ( .B(B[167]), .A(n39), .Z(n17491) );
  XNOR U17872 ( .A(n17499), .B(n17601), .Z(n17492) );
  XNOR U17873 ( .A(n17498), .B(n17496), .Z(n17601) );
  AND U17874 ( .A(n17602), .B(n17603), .Z(n17496) );
  NANDN U17875 ( .A(n17604), .B(n17605), .Z(n17603) );
  OR U17876 ( .A(n17606), .B(n17607), .Z(n17605) );
  NAND U17877 ( .A(n17607), .B(n17606), .Z(n17602) );
  ANDN U17878 ( .B(B[168]), .A(n40), .Z(n17498) );
  XNOR U17879 ( .A(n17506), .B(n17608), .Z(n17499) );
  XNOR U17880 ( .A(n17505), .B(n17503), .Z(n17608) );
  AND U17881 ( .A(n17609), .B(n17610), .Z(n17503) );
  NANDN U17882 ( .A(n17611), .B(n17612), .Z(n17610) );
  NAND U17883 ( .A(n17613), .B(n17614), .Z(n17612) );
  ANDN U17884 ( .B(B[169]), .A(n41), .Z(n17505) );
  XOR U17885 ( .A(n17512), .B(n17615), .Z(n17506) );
  XNOR U17886 ( .A(n17510), .B(n17513), .Z(n17615) );
  NAND U17887 ( .A(A[2]), .B(B[170]), .Z(n17513) );
  NANDN U17888 ( .A(n17616), .B(n17617), .Z(n17510) );
  AND U17889 ( .A(A[0]), .B(B[171]), .Z(n17617) );
  XNOR U17890 ( .A(n17515), .B(n17618), .Z(n17512) );
  NAND U17891 ( .A(A[0]), .B(B[172]), .Z(n17618) );
  NAND U17892 ( .A(B[171]), .B(A[1]), .Z(n17515) );
  NAND U17893 ( .A(n17619), .B(n17620), .Z(n407) );
  NANDN U17894 ( .A(n17621), .B(n17622), .Z(n17620) );
  OR U17895 ( .A(n17623), .B(n17624), .Z(n17622) );
  NAND U17896 ( .A(n17624), .B(n17623), .Z(n17619) );
  XOR U17897 ( .A(n389), .B(n388), .Z(\A1[16] ) );
  XOR U17898 ( .A(n16614), .B(n17625), .Z(n388) );
  XNOR U17899 ( .A(n16613), .B(n16611), .Z(n17625) );
  AND U17900 ( .A(n17626), .B(n17627), .Z(n16611) );
  NANDN U17901 ( .A(n17628), .B(n17629), .Z(n17627) );
  NANDN U17902 ( .A(n17630), .B(n17631), .Z(n17629) );
  NANDN U17903 ( .A(n17631), .B(n17630), .Z(n17626) );
  ANDN U17904 ( .B(B[3]), .A(n29), .Z(n16613) );
  XNOR U17905 ( .A(n16520), .B(n17632), .Z(n16614) );
  XNOR U17906 ( .A(n16519), .B(n16517), .Z(n17632) );
  AND U17907 ( .A(n17633), .B(n17634), .Z(n16517) );
  NANDN U17908 ( .A(n17635), .B(n17636), .Z(n17634) );
  OR U17909 ( .A(n17637), .B(n17638), .Z(n17636) );
  NAND U17910 ( .A(n17638), .B(n17637), .Z(n17633) );
  ANDN U17911 ( .B(B[4]), .A(n30), .Z(n16519) );
  XNOR U17912 ( .A(n16527), .B(n17639), .Z(n16520) );
  XNOR U17913 ( .A(n16526), .B(n16524), .Z(n17639) );
  AND U17914 ( .A(n17640), .B(n17641), .Z(n16524) );
  NANDN U17915 ( .A(n17642), .B(n17643), .Z(n17641) );
  NANDN U17916 ( .A(n17644), .B(n17645), .Z(n17643) );
  NANDN U17917 ( .A(n17645), .B(n17644), .Z(n17640) );
  ANDN U17918 ( .B(B[5]), .A(n31), .Z(n16526) );
  XNOR U17919 ( .A(n16534), .B(n17646), .Z(n16527) );
  XNOR U17920 ( .A(n16533), .B(n16531), .Z(n17646) );
  AND U17921 ( .A(n17647), .B(n17648), .Z(n16531) );
  NANDN U17922 ( .A(n17649), .B(n17650), .Z(n17648) );
  OR U17923 ( .A(n17651), .B(n17652), .Z(n17650) );
  NAND U17924 ( .A(n17652), .B(n17651), .Z(n17647) );
  ANDN U17925 ( .B(B[6]), .A(n32), .Z(n16533) );
  XNOR U17926 ( .A(n16541), .B(n17653), .Z(n16534) );
  XNOR U17927 ( .A(n16540), .B(n16538), .Z(n17653) );
  AND U17928 ( .A(n17654), .B(n17655), .Z(n16538) );
  NANDN U17929 ( .A(n17656), .B(n17657), .Z(n17655) );
  NANDN U17930 ( .A(n17658), .B(n17659), .Z(n17657) );
  NANDN U17931 ( .A(n17659), .B(n17658), .Z(n17654) );
  ANDN U17932 ( .B(B[7]), .A(n33), .Z(n16540) );
  XNOR U17933 ( .A(n16548), .B(n17660), .Z(n16541) );
  XNOR U17934 ( .A(n16547), .B(n16545), .Z(n17660) );
  AND U17935 ( .A(n17661), .B(n17662), .Z(n16545) );
  NANDN U17936 ( .A(n17663), .B(n17664), .Z(n17662) );
  OR U17937 ( .A(n17665), .B(n17666), .Z(n17664) );
  NAND U17938 ( .A(n17666), .B(n17665), .Z(n17661) );
  ANDN U17939 ( .B(B[8]), .A(n34), .Z(n16547) );
  XNOR U17940 ( .A(n16555), .B(n17667), .Z(n16548) );
  XNOR U17941 ( .A(n16554), .B(n16552), .Z(n17667) );
  AND U17942 ( .A(n17668), .B(n17669), .Z(n16552) );
  NANDN U17943 ( .A(n17670), .B(n17671), .Z(n17669) );
  NANDN U17944 ( .A(n17672), .B(n17673), .Z(n17671) );
  NANDN U17945 ( .A(n17673), .B(n17672), .Z(n17668) );
  ANDN U17946 ( .B(B[9]), .A(n35), .Z(n16554) );
  XNOR U17947 ( .A(n16562), .B(n17674), .Z(n16555) );
  XNOR U17948 ( .A(n16561), .B(n16559), .Z(n17674) );
  AND U17949 ( .A(n17675), .B(n17676), .Z(n16559) );
  NANDN U17950 ( .A(n17677), .B(n17678), .Z(n17676) );
  OR U17951 ( .A(n17679), .B(n17680), .Z(n17678) );
  NAND U17952 ( .A(n17680), .B(n17679), .Z(n17675) );
  ANDN U17953 ( .B(B[10]), .A(n36), .Z(n16561) );
  XNOR U17954 ( .A(n16569), .B(n17681), .Z(n16562) );
  XNOR U17955 ( .A(n16568), .B(n16566), .Z(n17681) );
  AND U17956 ( .A(n17682), .B(n17683), .Z(n16566) );
  NANDN U17957 ( .A(n17684), .B(n17685), .Z(n17683) );
  NANDN U17958 ( .A(n17686), .B(n17687), .Z(n17685) );
  NANDN U17959 ( .A(n17687), .B(n17686), .Z(n17682) );
  ANDN U17960 ( .B(B[11]), .A(n37), .Z(n16568) );
  XNOR U17961 ( .A(n16576), .B(n17688), .Z(n16569) );
  XNOR U17962 ( .A(n16575), .B(n16573), .Z(n17688) );
  AND U17963 ( .A(n17689), .B(n17690), .Z(n16573) );
  NANDN U17964 ( .A(n17691), .B(n17692), .Z(n17690) );
  OR U17965 ( .A(n17693), .B(n17694), .Z(n17692) );
  NAND U17966 ( .A(n17694), .B(n17693), .Z(n17689) );
  ANDN U17967 ( .B(B[12]), .A(n38), .Z(n16575) );
  XNOR U17968 ( .A(n16583), .B(n17695), .Z(n16576) );
  XNOR U17969 ( .A(n16582), .B(n16580), .Z(n17695) );
  AND U17970 ( .A(n17696), .B(n17697), .Z(n16580) );
  NANDN U17971 ( .A(n17698), .B(n17699), .Z(n17697) );
  NANDN U17972 ( .A(n17700), .B(n17701), .Z(n17699) );
  NANDN U17973 ( .A(n17701), .B(n17700), .Z(n17696) );
  ANDN U17974 ( .B(B[13]), .A(n39), .Z(n16582) );
  XNOR U17975 ( .A(n16590), .B(n17702), .Z(n16583) );
  XNOR U17976 ( .A(n16589), .B(n16587), .Z(n17702) );
  AND U17977 ( .A(n17703), .B(n17704), .Z(n16587) );
  NANDN U17978 ( .A(n17705), .B(n17706), .Z(n17704) );
  OR U17979 ( .A(n17707), .B(n17708), .Z(n17706) );
  NAND U17980 ( .A(n17708), .B(n17707), .Z(n17703) );
  ANDN U17981 ( .B(B[14]), .A(n40), .Z(n16589) );
  XNOR U17982 ( .A(n16597), .B(n17709), .Z(n16590) );
  XNOR U17983 ( .A(n16596), .B(n16594), .Z(n17709) );
  AND U17984 ( .A(n17710), .B(n17711), .Z(n16594) );
  NANDN U17985 ( .A(n17712), .B(n17713), .Z(n17711) );
  NAND U17986 ( .A(n17714), .B(n17715), .Z(n17713) );
  ANDN U17987 ( .B(B[15]), .A(n41), .Z(n16596) );
  XOR U17988 ( .A(n16603), .B(n17716), .Z(n16597) );
  XNOR U17989 ( .A(n16601), .B(n16604), .Z(n17716) );
  NAND U17990 ( .A(A[2]), .B(B[16]), .Z(n16604) );
  NANDN U17991 ( .A(n17717), .B(n17718), .Z(n16601) );
  AND U17992 ( .A(A[0]), .B(B[17]), .Z(n17718) );
  XNOR U17993 ( .A(n16606), .B(n17719), .Z(n16603) );
  NAND U17994 ( .A(A[0]), .B(B[18]), .Z(n17719) );
  NAND U17995 ( .A(B[17]), .B(A[1]), .Z(n16606) );
  NAND U17996 ( .A(n17720), .B(n17721), .Z(n389) );
  NANDN U17997 ( .A(n17722), .B(n17723), .Z(n17721) );
  OR U17998 ( .A(n17724), .B(n17725), .Z(n17723) );
  NAND U17999 ( .A(n17725), .B(n17724), .Z(n17720) );
  XOR U18000 ( .A(n409), .B(n408), .Z(\A1[169] ) );
  XOR U18001 ( .A(n17624), .B(n17726), .Z(n408) );
  XNOR U18002 ( .A(n17623), .B(n17621), .Z(n17726) );
  AND U18003 ( .A(n17727), .B(n17728), .Z(n17621) );
  NANDN U18004 ( .A(n17729), .B(n17730), .Z(n17728) );
  NANDN U18005 ( .A(n17731), .B(n17732), .Z(n17730) );
  NANDN U18006 ( .A(n17732), .B(n17731), .Z(n17727) );
  ANDN U18007 ( .B(B[156]), .A(n29), .Z(n17623) );
  XNOR U18008 ( .A(n17530), .B(n17733), .Z(n17624) );
  XNOR U18009 ( .A(n17529), .B(n17527), .Z(n17733) );
  AND U18010 ( .A(n17734), .B(n17735), .Z(n17527) );
  NANDN U18011 ( .A(n17736), .B(n17737), .Z(n17735) );
  OR U18012 ( .A(n17738), .B(n17739), .Z(n17737) );
  NAND U18013 ( .A(n17739), .B(n17738), .Z(n17734) );
  ANDN U18014 ( .B(B[157]), .A(n30), .Z(n17529) );
  XNOR U18015 ( .A(n17537), .B(n17740), .Z(n17530) );
  XNOR U18016 ( .A(n17536), .B(n17534), .Z(n17740) );
  AND U18017 ( .A(n17741), .B(n17742), .Z(n17534) );
  NANDN U18018 ( .A(n17743), .B(n17744), .Z(n17742) );
  NANDN U18019 ( .A(n17745), .B(n17746), .Z(n17744) );
  NANDN U18020 ( .A(n17746), .B(n17745), .Z(n17741) );
  ANDN U18021 ( .B(B[158]), .A(n31), .Z(n17536) );
  XNOR U18022 ( .A(n17544), .B(n17747), .Z(n17537) );
  XNOR U18023 ( .A(n17543), .B(n17541), .Z(n17747) );
  AND U18024 ( .A(n17748), .B(n17749), .Z(n17541) );
  NANDN U18025 ( .A(n17750), .B(n17751), .Z(n17749) );
  OR U18026 ( .A(n17752), .B(n17753), .Z(n17751) );
  NAND U18027 ( .A(n17753), .B(n17752), .Z(n17748) );
  ANDN U18028 ( .B(B[159]), .A(n32), .Z(n17543) );
  XNOR U18029 ( .A(n17551), .B(n17754), .Z(n17544) );
  XNOR U18030 ( .A(n17550), .B(n17548), .Z(n17754) );
  AND U18031 ( .A(n17755), .B(n17756), .Z(n17548) );
  NANDN U18032 ( .A(n17757), .B(n17758), .Z(n17756) );
  NANDN U18033 ( .A(n17759), .B(n17760), .Z(n17758) );
  NANDN U18034 ( .A(n17760), .B(n17759), .Z(n17755) );
  ANDN U18035 ( .B(B[160]), .A(n33), .Z(n17550) );
  XNOR U18036 ( .A(n17558), .B(n17761), .Z(n17551) );
  XNOR U18037 ( .A(n17557), .B(n17555), .Z(n17761) );
  AND U18038 ( .A(n17762), .B(n17763), .Z(n17555) );
  NANDN U18039 ( .A(n17764), .B(n17765), .Z(n17763) );
  OR U18040 ( .A(n17766), .B(n17767), .Z(n17765) );
  NAND U18041 ( .A(n17767), .B(n17766), .Z(n17762) );
  ANDN U18042 ( .B(B[161]), .A(n34), .Z(n17557) );
  XNOR U18043 ( .A(n17565), .B(n17768), .Z(n17558) );
  XNOR U18044 ( .A(n17564), .B(n17562), .Z(n17768) );
  AND U18045 ( .A(n17769), .B(n17770), .Z(n17562) );
  NANDN U18046 ( .A(n17771), .B(n17772), .Z(n17770) );
  NANDN U18047 ( .A(n17773), .B(n17774), .Z(n17772) );
  NANDN U18048 ( .A(n17774), .B(n17773), .Z(n17769) );
  ANDN U18049 ( .B(B[162]), .A(n35), .Z(n17564) );
  XNOR U18050 ( .A(n17572), .B(n17775), .Z(n17565) );
  XNOR U18051 ( .A(n17571), .B(n17569), .Z(n17775) );
  AND U18052 ( .A(n17776), .B(n17777), .Z(n17569) );
  NANDN U18053 ( .A(n17778), .B(n17779), .Z(n17777) );
  OR U18054 ( .A(n17780), .B(n17781), .Z(n17779) );
  NAND U18055 ( .A(n17781), .B(n17780), .Z(n17776) );
  ANDN U18056 ( .B(B[163]), .A(n36), .Z(n17571) );
  XNOR U18057 ( .A(n17579), .B(n17782), .Z(n17572) );
  XNOR U18058 ( .A(n17578), .B(n17576), .Z(n17782) );
  AND U18059 ( .A(n17783), .B(n17784), .Z(n17576) );
  NANDN U18060 ( .A(n17785), .B(n17786), .Z(n17784) );
  NANDN U18061 ( .A(n17787), .B(n17788), .Z(n17786) );
  NANDN U18062 ( .A(n17788), .B(n17787), .Z(n17783) );
  ANDN U18063 ( .B(B[164]), .A(n37), .Z(n17578) );
  XNOR U18064 ( .A(n17586), .B(n17789), .Z(n17579) );
  XNOR U18065 ( .A(n17585), .B(n17583), .Z(n17789) );
  AND U18066 ( .A(n17790), .B(n17791), .Z(n17583) );
  NANDN U18067 ( .A(n17792), .B(n17793), .Z(n17791) );
  OR U18068 ( .A(n17794), .B(n17795), .Z(n17793) );
  NAND U18069 ( .A(n17795), .B(n17794), .Z(n17790) );
  ANDN U18070 ( .B(B[165]), .A(n38), .Z(n17585) );
  XNOR U18071 ( .A(n17593), .B(n17796), .Z(n17586) );
  XNOR U18072 ( .A(n17592), .B(n17590), .Z(n17796) );
  AND U18073 ( .A(n17797), .B(n17798), .Z(n17590) );
  NANDN U18074 ( .A(n17799), .B(n17800), .Z(n17798) );
  NANDN U18075 ( .A(n17801), .B(n17802), .Z(n17800) );
  NANDN U18076 ( .A(n17802), .B(n17801), .Z(n17797) );
  ANDN U18077 ( .B(B[166]), .A(n39), .Z(n17592) );
  XNOR U18078 ( .A(n17600), .B(n17803), .Z(n17593) );
  XNOR U18079 ( .A(n17599), .B(n17597), .Z(n17803) );
  AND U18080 ( .A(n17804), .B(n17805), .Z(n17597) );
  NANDN U18081 ( .A(n17806), .B(n17807), .Z(n17805) );
  OR U18082 ( .A(n17808), .B(n17809), .Z(n17807) );
  NAND U18083 ( .A(n17809), .B(n17808), .Z(n17804) );
  ANDN U18084 ( .B(B[167]), .A(n40), .Z(n17599) );
  XNOR U18085 ( .A(n17607), .B(n17810), .Z(n17600) );
  XNOR U18086 ( .A(n17606), .B(n17604), .Z(n17810) );
  AND U18087 ( .A(n17811), .B(n17812), .Z(n17604) );
  NANDN U18088 ( .A(n17813), .B(n17814), .Z(n17812) );
  NAND U18089 ( .A(n17815), .B(n17816), .Z(n17814) );
  ANDN U18090 ( .B(B[168]), .A(n41), .Z(n17606) );
  XOR U18091 ( .A(n17613), .B(n17817), .Z(n17607) );
  XNOR U18092 ( .A(n17611), .B(n17614), .Z(n17817) );
  NAND U18093 ( .A(A[2]), .B(B[169]), .Z(n17614) );
  NANDN U18094 ( .A(n17818), .B(n17819), .Z(n17611) );
  AND U18095 ( .A(A[0]), .B(B[170]), .Z(n17819) );
  XNOR U18096 ( .A(n17616), .B(n17820), .Z(n17613) );
  NAND U18097 ( .A(A[0]), .B(B[171]), .Z(n17820) );
  NAND U18098 ( .A(B[170]), .B(A[1]), .Z(n17616) );
  NAND U18099 ( .A(n17821), .B(n17822), .Z(n409) );
  NANDN U18100 ( .A(n17823), .B(n17824), .Z(n17822) );
  OR U18101 ( .A(n17825), .B(n17826), .Z(n17824) );
  NAND U18102 ( .A(n17826), .B(n17825), .Z(n17821) );
  XOR U18103 ( .A(n413), .B(n412), .Z(\A1[168] ) );
  XOR U18104 ( .A(n17826), .B(n17827), .Z(n412) );
  XNOR U18105 ( .A(n17825), .B(n17823), .Z(n17827) );
  AND U18106 ( .A(n17828), .B(n17829), .Z(n17823) );
  NANDN U18107 ( .A(n17830), .B(n17831), .Z(n17829) );
  NANDN U18108 ( .A(n17832), .B(n17833), .Z(n17831) );
  NANDN U18109 ( .A(n17833), .B(n17832), .Z(n17828) );
  ANDN U18110 ( .B(B[155]), .A(n29), .Z(n17825) );
  XNOR U18111 ( .A(n17732), .B(n17834), .Z(n17826) );
  XNOR U18112 ( .A(n17731), .B(n17729), .Z(n17834) );
  AND U18113 ( .A(n17835), .B(n17836), .Z(n17729) );
  NANDN U18114 ( .A(n17837), .B(n17838), .Z(n17836) );
  OR U18115 ( .A(n17839), .B(n17840), .Z(n17838) );
  NAND U18116 ( .A(n17840), .B(n17839), .Z(n17835) );
  ANDN U18117 ( .B(B[156]), .A(n30), .Z(n17731) );
  XNOR U18118 ( .A(n17739), .B(n17841), .Z(n17732) );
  XNOR U18119 ( .A(n17738), .B(n17736), .Z(n17841) );
  AND U18120 ( .A(n17842), .B(n17843), .Z(n17736) );
  NANDN U18121 ( .A(n17844), .B(n17845), .Z(n17843) );
  NANDN U18122 ( .A(n17846), .B(n17847), .Z(n17845) );
  NANDN U18123 ( .A(n17847), .B(n17846), .Z(n17842) );
  ANDN U18124 ( .B(B[157]), .A(n31), .Z(n17738) );
  XNOR U18125 ( .A(n17746), .B(n17848), .Z(n17739) );
  XNOR U18126 ( .A(n17745), .B(n17743), .Z(n17848) );
  AND U18127 ( .A(n17849), .B(n17850), .Z(n17743) );
  NANDN U18128 ( .A(n17851), .B(n17852), .Z(n17850) );
  OR U18129 ( .A(n17853), .B(n17854), .Z(n17852) );
  NAND U18130 ( .A(n17854), .B(n17853), .Z(n17849) );
  ANDN U18131 ( .B(B[158]), .A(n32), .Z(n17745) );
  XNOR U18132 ( .A(n17753), .B(n17855), .Z(n17746) );
  XNOR U18133 ( .A(n17752), .B(n17750), .Z(n17855) );
  AND U18134 ( .A(n17856), .B(n17857), .Z(n17750) );
  NANDN U18135 ( .A(n17858), .B(n17859), .Z(n17857) );
  NANDN U18136 ( .A(n17860), .B(n17861), .Z(n17859) );
  NANDN U18137 ( .A(n17861), .B(n17860), .Z(n17856) );
  ANDN U18138 ( .B(B[159]), .A(n33), .Z(n17752) );
  XNOR U18139 ( .A(n17760), .B(n17862), .Z(n17753) );
  XNOR U18140 ( .A(n17759), .B(n17757), .Z(n17862) );
  AND U18141 ( .A(n17863), .B(n17864), .Z(n17757) );
  NANDN U18142 ( .A(n17865), .B(n17866), .Z(n17864) );
  OR U18143 ( .A(n17867), .B(n17868), .Z(n17866) );
  NAND U18144 ( .A(n17868), .B(n17867), .Z(n17863) );
  ANDN U18145 ( .B(B[160]), .A(n34), .Z(n17759) );
  XNOR U18146 ( .A(n17767), .B(n17869), .Z(n17760) );
  XNOR U18147 ( .A(n17766), .B(n17764), .Z(n17869) );
  AND U18148 ( .A(n17870), .B(n17871), .Z(n17764) );
  NANDN U18149 ( .A(n17872), .B(n17873), .Z(n17871) );
  NANDN U18150 ( .A(n17874), .B(n17875), .Z(n17873) );
  NANDN U18151 ( .A(n17875), .B(n17874), .Z(n17870) );
  ANDN U18152 ( .B(B[161]), .A(n35), .Z(n17766) );
  XNOR U18153 ( .A(n17774), .B(n17876), .Z(n17767) );
  XNOR U18154 ( .A(n17773), .B(n17771), .Z(n17876) );
  AND U18155 ( .A(n17877), .B(n17878), .Z(n17771) );
  NANDN U18156 ( .A(n17879), .B(n17880), .Z(n17878) );
  OR U18157 ( .A(n17881), .B(n17882), .Z(n17880) );
  NAND U18158 ( .A(n17882), .B(n17881), .Z(n17877) );
  ANDN U18159 ( .B(B[162]), .A(n36), .Z(n17773) );
  XNOR U18160 ( .A(n17781), .B(n17883), .Z(n17774) );
  XNOR U18161 ( .A(n17780), .B(n17778), .Z(n17883) );
  AND U18162 ( .A(n17884), .B(n17885), .Z(n17778) );
  NANDN U18163 ( .A(n17886), .B(n17887), .Z(n17885) );
  NANDN U18164 ( .A(n17888), .B(n17889), .Z(n17887) );
  NANDN U18165 ( .A(n17889), .B(n17888), .Z(n17884) );
  ANDN U18166 ( .B(B[163]), .A(n37), .Z(n17780) );
  XNOR U18167 ( .A(n17788), .B(n17890), .Z(n17781) );
  XNOR U18168 ( .A(n17787), .B(n17785), .Z(n17890) );
  AND U18169 ( .A(n17891), .B(n17892), .Z(n17785) );
  NANDN U18170 ( .A(n17893), .B(n17894), .Z(n17892) );
  OR U18171 ( .A(n17895), .B(n17896), .Z(n17894) );
  NAND U18172 ( .A(n17896), .B(n17895), .Z(n17891) );
  ANDN U18173 ( .B(B[164]), .A(n38), .Z(n17787) );
  XNOR U18174 ( .A(n17795), .B(n17897), .Z(n17788) );
  XNOR U18175 ( .A(n17794), .B(n17792), .Z(n17897) );
  AND U18176 ( .A(n17898), .B(n17899), .Z(n17792) );
  NANDN U18177 ( .A(n17900), .B(n17901), .Z(n17899) );
  NANDN U18178 ( .A(n17902), .B(n17903), .Z(n17901) );
  NANDN U18179 ( .A(n17903), .B(n17902), .Z(n17898) );
  ANDN U18180 ( .B(B[165]), .A(n39), .Z(n17794) );
  XNOR U18181 ( .A(n17802), .B(n17904), .Z(n17795) );
  XNOR U18182 ( .A(n17801), .B(n17799), .Z(n17904) );
  AND U18183 ( .A(n17905), .B(n17906), .Z(n17799) );
  NANDN U18184 ( .A(n17907), .B(n17908), .Z(n17906) );
  OR U18185 ( .A(n17909), .B(n17910), .Z(n17908) );
  NAND U18186 ( .A(n17910), .B(n17909), .Z(n17905) );
  ANDN U18187 ( .B(B[166]), .A(n40), .Z(n17801) );
  XNOR U18188 ( .A(n17809), .B(n17911), .Z(n17802) );
  XNOR U18189 ( .A(n17808), .B(n17806), .Z(n17911) );
  AND U18190 ( .A(n17912), .B(n17913), .Z(n17806) );
  NANDN U18191 ( .A(n17914), .B(n17915), .Z(n17913) );
  NAND U18192 ( .A(n17916), .B(n17917), .Z(n17915) );
  ANDN U18193 ( .B(B[167]), .A(n41), .Z(n17808) );
  XOR U18194 ( .A(n17815), .B(n17918), .Z(n17809) );
  XNOR U18195 ( .A(n17813), .B(n17816), .Z(n17918) );
  NAND U18196 ( .A(A[2]), .B(B[168]), .Z(n17816) );
  NANDN U18197 ( .A(n17919), .B(n17920), .Z(n17813) );
  AND U18198 ( .A(A[0]), .B(B[169]), .Z(n17920) );
  XNOR U18199 ( .A(n17818), .B(n17921), .Z(n17815) );
  NAND U18200 ( .A(A[0]), .B(B[170]), .Z(n17921) );
  NAND U18201 ( .A(B[169]), .B(A[1]), .Z(n17818) );
  NAND U18202 ( .A(n17922), .B(n17923), .Z(n413) );
  NANDN U18203 ( .A(n17924), .B(n17925), .Z(n17923) );
  OR U18204 ( .A(n17926), .B(n17927), .Z(n17925) );
  NAND U18205 ( .A(n17927), .B(n17926), .Z(n17922) );
  XOR U18206 ( .A(n415), .B(n414), .Z(\A1[167] ) );
  XOR U18207 ( .A(n17927), .B(n17928), .Z(n414) );
  XNOR U18208 ( .A(n17926), .B(n17924), .Z(n17928) );
  AND U18209 ( .A(n17929), .B(n17930), .Z(n17924) );
  NANDN U18210 ( .A(n17931), .B(n17932), .Z(n17930) );
  NANDN U18211 ( .A(n17933), .B(n17934), .Z(n17932) );
  NANDN U18212 ( .A(n17934), .B(n17933), .Z(n17929) );
  ANDN U18213 ( .B(B[154]), .A(n29), .Z(n17926) );
  XNOR U18214 ( .A(n17833), .B(n17935), .Z(n17927) );
  XNOR U18215 ( .A(n17832), .B(n17830), .Z(n17935) );
  AND U18216 ( .A(n17936), .B(n17937), .Z(n17830) );
  NANDN U18217 ( .A(n17938), .B(n17939), .Z(n17937) );
  OR U18218 ( .A(n17940), .B(n17941), .Z(n17939) );
  NAND U18219 ( .A(n17941), .B(n17940), .Z(n17936) );
  ANDN U18220 ( .B(B[155]), .A(n30), .Z(n17832) );
  XNOR U18221 ( .A(n17840), .B(n17942), .Z(n17833) );
  XNOR U18222 ( .A(n17839), .B(n17837), .Z(n17942) );
  AND U18223 ( .A(n17943), .B(n17944), .Z(n17837) );
  NANDN U18224 ( .A(n17945), .B(n17946), .Z(n17944) );
  NANDN U18225 ( .A(n17947), .B(n17948), .Z(n17946) );
  NANDN U18226 ( .A(n17948), .B(n17947), .Z(n17943) );
  ANDN U18227 ( .B(B[156]), .A(n31), .Z(n17839) );
  XNOR U18228 ( .A(n17847), .B(n17949), .Z(n17840) );
  XNOR U18229 ( .A(n17846), .B(n17844), .Z(n17949) );
  AND U18230 ( .A(n17950), .B(n17951), .Z(n17844) );
  NANDN U18231 ( .A(n17952), .B(n17953), .Z(n17951) );
  OR U18232 ( .A(n17954), .B(n17955), .Z(n17953) );
  NAND U18233 ( .A(n17955), .B(n17954), .Z(n17950) );
  ANDN U18234 ( .B(B[157]), .A(n32), .Z(n17846) );
  XNOR U18235 ( .A(n17854), .B(n17956), .Z(n17847) );
  XNOR U18236 ( .A(n17853), .B(n17851), .Z(n17956) );
  AND U18237 ( .A(n17957), .B(n17958), .Z(n17851) );
  NANDN U18238 ( .A(n17959), .B(n17960), .Z(n17958) );
  NANDN U18239 ( .A(n17961), .B(n17962), .Z(n17960) );
  NANDN U18240 ( .A(n17962), .B(n17961), .Z(n17957) );
  ANDN U18241 ( .B(B[158]), .A(n33), .Z(n17853) );
  XNOR U18242 ( .A(n17861), .B(n17963), .Z(n17854) );
  XNOR U18243 ( .A(n17860), .B(n17858), .Z(n17963) );
  AND U18244 ( .A(n17964), .B(n17965), .Z(n17858) );
  NANDN U18245 ( .A(n17966), .B(n17967), .Z(n17965) );
  OR U18246 ( .A(n17968), .B(n17969), .Z(n17967) );
  NAND U18247 ( .A(n17969), .B(n17968), .Z(n17964) );
  ANDN U18248 ( .B(B[159]), .A(n34), .Z(n17860) );
  XNOR U18249 ( .A(n17868), .B(n17970), .Z(n17861) );
  XNOR U18250 ( .A(n17867), .B(n17865), .Z(n17970) );
  AND U18251 ( .A(n17971), .B(n17972), .Z(n17865) );
  NANDN U18252 ( .A(n17973), .B(n17974), .Z(n17972) );
  NANDN U18253 ( .A(n17975), .B(n17976), .Z(n17974) );
  NANDN U18254 ( .A(n17976), .B(n17975), .Z(n17971) );
  ANDN U18255 ( .B(B[160]), .A(n35), .Z(n17867) );
  XNOR U18256 ( .A(n17875), .B(n17977), .Z(n17868) );
  XNOR U18257 ( .A(n17874), .B(n17872), .Z(n17977) );
  AND U18258 ( .A(n17978), .B(n17979), .Z(n17872) );
  NANDN U18259 ( .A(n17980), .B(n17981), .Z(n17979) );
  OR U18260 ( .A(n17982), .B(n17983), .Z(n17981) );
  NAND U18261 ( .A(n17983), .B(n17982), .Z(n17978) );
  ANDN U18262 ( .B(B[161]), .A(n36), .Z(n17874) );
  XNOR U18263 ( .A(n17882), .B(n17984), .Z(n17875) );
  XNOR U18264 ( .A(n17881), .B(n17879), .Z(n17984) );
  AND U18265 ( .A(n17985), .B(n17986), .Z(n17879) );
  NANDN U18266 ( .A(n17987), .B(n17988), .Z(n17986) );
  NANDN U18267 ( .A(n17989), .B(n17990), .Z(n17988) );
  NANDN U18268 ( .A(n17990), .B(n17989), .Z(n17985) );
  ANDN U18269 ( .B(B[162]), .A(n37), .Z(n17881) );
  XNOR U18270 ( .A(n17889), .B(n17991), .Z(n17882) );
  XNOR U18271 ( .A(n17888), .B(n17886), .Z(n17991) );
  AND U18272 ( .A(n17992), .B(n17993), .Z(n17886) );
  NANDN U18273 ( .A(n17994), .B(n17995), .Z(n17993) );
  OR U18274 ( .A(n17996), .B(n17997), .Z(n17995) );
  NAND U18275 ( .A(n17997), .B(n17996), .Z(n17992) );
  ANDN U18276 ( .B(B[163]), .A(n38), .Z(n17888) );
  XNOR U18277 ( .A(n17896), .B(n17998), .Z(n17889) );
  XNOR U18278 ( .A(n17895), .B(n17893), .Z(n17998) );
  AND U18279 ( .A(n17999), .B(n18000), .Z(n17893) );
  NANDN U18280 ( .A(n18001), .B(n18002), .Z(n18000) );
  NANDN U18281 ( .A(n18003), .B(n18004), .Z(n18002) );
  NANDN U18282 ( .A(n18004), .B(n18003), .Z(n17999) );
  ANDN U18283 ( .B(B[164]), .A(n39), .Z(n17895) );
  XNOR U18284 ( .A(n17903), .B(n18005), .Z(n17896) );
  XNOR U18285 ( .A(n17902), .B(n17900), .Z(n18005) );
  AND U18286 ( .A(n18006), .B(n18007), .Z(n17900) );
  NANDN U18287 ( .A(n18008), .B(n18009), .Z(n18007) );
  OR U18288 ( .A(n18010), .B(n18011), .Z(n18009) );
  NAND U18289 ( .A(n18011), .B(n18010), .Z(n18006) );
  ANDN U18290 ( .B(B[165]), .A(n40), .Z(n17902) );
  XNOR U18291 ( .A(n17910), .B(n18012), .Z(n17903) );
  XNOR U18292 ( .A(n17909), .B(n17907), .Z(n18012) );
  AND U18293 ( .A(n18013), .B(n18014), .Z(n17907) );
  NANDN U18294 ( .A(n18015), .B(n18016), .Z(n18014) );
  NAND U18295 ( .A(n18017), .B(n18018), .Z(n18016) );
  ANDN U18296 ( .B(B[166]), .A(n41), .Z(n17909) );
  XOR U18297 ( .A(n17916), .B(n18019), .Z(n17910) );
  XNOR U18298 ( .A(n17914), .B(n17917), .Z(n18019) );
  NAND U18299 ( .A(A[2]), .B(B[167]), .Z(n17917) );
  NANDN U18300 ( .A(n18020), .B(n18021), .Z(n17914) );
  AND U18301 ( .A(A[0]), .B(B[168]), .Z(n18021) );
  XNOR U18302 ( .A(n17919), .B(n18022), .Z(n17916) );
  NAND U18303 ( .A(A[0]), .B(B[169]), .Z(n18022) );
  NAND U18304 ( .A(B[168]), .B(A[1]), .Z(n17919) );
  NAND U18305 ( .A(n18023), .B(n18024), .Z(n415) );
  NANDN U18306 ( .A(n18025), .B(n18026), .Z(n18024) );
  OR U18307 ( .A(n18027), .B(n18028), .Z(n18026) );
  NAND U18308 ( .A(n18028), .B(n18027), .Z(n18023) );
  XOR U18309 ( .A(n417), .B(n416), .Z(\A1[166] ) );
  XOR U18310 ( .A(n18028), .B(n18029), .Z(n416) );
  XNOR U18311 ( .A(n18027), .B(n18025), .Z(n18029) );
  AND U18312 ( .A(n18030), .B(n18031), .Z(n18025) );
  NANDN U18313 ( .A(n18032), .B(n18033), .Z(n18031) );
  NANDN U18314 ( .A(n18034), .B(n18035), .Z(n18033) );
  NANDN U18315 ( .A(n18035), .B(n18034), .Z(n18030) );
  ANDN U18316 ( .B(B[153]), .A(n29), .Z(n18027) );
  XNOR U18317 ( .A(n17934), .B(n18036), .Z(n18028) );
  XNOR U18318 ( .A(n17933), .B(n17931), .Z(n18036) );
  AND U18319 ( .A(n18037), .B(n18038), .Z(n17931) );
  NANDN U18320 ( .A(n18039), .B(n18040), .Z(n18038) );
  OR U18321 ( .A(n18041), .B(n18042), .Z(n18040) );
  NAND U18322 ( .A(n18042), .B(n18041), .Z(n18037) );
  ANDN U18323 ( .B(B[154]), .A(n30), .Z(n17933) );
  XNOR U18324 ( .A(n17941), .B(n18043), .Z(n17934) );
  XNOR U18325 ( .A(n17940), .B(n17938), .Z(n18043) );
  AND U18326 ( .A(n18044), .B(n18045), .Z(n17938) );
  NANDN U18327 ( .A(n18046), .B(n18047), .Z(n18045) );
  NANDN U18328 ( .A(n18048), .B(n18049), .Z(n18047) );
  NANDN U18329 ( .A(n18049), .B(n18048), .Z(n18044) );
  ANDN U18330 ( .B(B[155]), .A(n31), .Z(n17940) );
  XNOR U18331 ( .A(n17948), .B(n18050), .Z(n17941) );
  XNOR U18332 ( .A(n17947), .B(n17945), .Z(n18050) );
  AND U18333 ( .A(n18051), .B(n18052), .Z(n17945) );
  NANDN U18334 ( .A(n18053), .B(n18054), .Z(n18052) );
  OR U18335 ( .A(n18055), .B(n18056), .Z(n18054) );
  NAND U18336 ( .A(n18056), .B(n18055), .Z(n18051) );
  ANDN U18337 ( .B(B[156]), .A(n32), .Z(n17947) );
  XNOR U18338 ( .A(n17955), .B(n18057), .Z(n17948) );
  XNOR U18339 ( .A(n17954), .B(n17952), .Z(n18057) );
  AND U18340 ( .A(n18058), .B(n18059), .Z(n17952) );
  NANDN U18341 ( .A(n18060), .B(n18061), .Z(n18059) );
  NANDN U18342 ( .A(n18062), .B(n18063), .Z(n18061) );
  NANDN U18343 ( .A(n18063), .B(n18062), .Z(n18058) );
  ANDN U18344 ( .B(B[157]), .A(n33), .Z(n17954) );
  XNOR U18345 ( .A(n17962), .B(n18064), .Z(n17955) );
  XNOR U18346 ( .A(n17961), .B(n17959), .Z(n18064) );
  AND U18347 ( .A(n18065), .B(n18066), .Z(n17959) );
  NANDN U18348 ( .A(n18067), .B(n18068), .Z(n18066) );
  OR U18349 ( .A(n18069), .B(n18070), .Z(n18068) );
  NAND U18350 ( .A(n18070), .B(n18069), .Z(n18065) );
  ANDN U18351 ( .B(B[158]), .A(n34), .Z(n17961) );
  XNOR U18352 ( .A(n17969), .B(n18071), .Z(n17962) );
  XNOR U18353 ( .A(n17968), .B(n17966), .Z(n18071) );
  AND U18354 ( .A(n18072), .B(n18073), .Z(n17966) );
  NANDN U18355 ( .A(n18074), .B(n18075), .Z(n18073) );
  NANDN U18356 ( .A(n18076), .B(n18077), .Z(n18075) );
  NANDN U18357 ( .A(n18077), .B(n18076), .Z(n18072) );
  ANDN U18358 ( .B(B[159]), .A(n35), .Z(n17968) );
  XNOR U18359 ( .A(n17976), .B(n18078), .Z(n17969) );
  XNOR U18360 ( .A(n17975), .B(n17973), .Z(n18078) );
  AND U18361 ( .A(n18079), .B(n18080), .Z(n17973) );
  NANDN U18362 ( .A(n18081), .B(n18082), .Z(n18080) );
  OR U18363 ( .A(n18083), .B(n18084), .Z(n18082) );
  NAND U18364 ( .A(n18084), .B(n18083), .Z(n18079) );
  ANDN U18365 ( .B(B[160]), .A(n36), .Z(n17975) );
  XNOR U18366 ( .A(n17983), .B(n18085), .Z(n17976) );
  XNOR U18367 ( .A(n17982), .B(n17980), .Z(n18085) );
  AND U18368 ( .A(n18086), .B(n18087), .Z(n17980) );
  NANDN U18369 ( .A(n18088), .B(n18089), .Z(n18087) );
  NANDN U18370 ( .A(n18090), .B(n18091), .Z(n18089) );
  NANDN U18371 ( .A(n18091), .B(n18090), .Z(n18086) );
  ANDN U18372 ( .B(B[161]), .A(n37), .Z(n17982) );
  XNOR U18373 ( .A(n17990), .B(n18092), .Z(n17983) );
  XNOR U18374 ( .A(n17989), .B(n17987), .Z(n18092) );
  AND U18375 ( .A(n18093), .B(n18094), .Z(n17987) );
  NANDN U18376 ( .A(n18095), .B(n18096), .Z(n18094) );
  OR U18377 ( .A(n18097), .B(n18098), .Z(n18096) );
  NAND U18378 ( .A(n18098), .B(n18097), .Z(n18093) );
  ANDN U18379 ( .B(B[162]), .A(n38), .Z(n17989) );
  XNOR U18380 ( .A(n17997), .B(n18099), .Z(n17990) );
  XNOR U18381 ( .A(n17996), .B(n17994), .Z(n18099) );
  AND U18382 ( .A(n18100), .B(n18101), .Z(n17994) );
  NANDN U18383 ( .A(n18102), .B(n18103), .Z(n18101) );
  NANDN U18384 ( .A(n18104), .B(n18105), .Z(n18103) );
  NANDN U18385 ( .A(n18105), .B(n18104), .Z(n18100) );
  ANDN U18386 ( .B(B[163]), .A(n39), .Z(n17996) );
  XNOR U18387 ( .A(n18004), .B(n18106), .Z(n17997) );
  XNOR U18388 ( .A(n18003), .B(n18001), .Z(n18106) );
  AND U18389 ( .A(n18107), .B(n18108), .Z(n18001) );
  NANDN U18390 ( .A(n18109), .B(n18110), .Z(n18108) );
  OR U18391 ( .A(n18111), .B(n18112), .Z(n18110) );
  NAND U18392 ( .A(n18112), .B(n18111), .Z(n18107) );
  ANDN U18393 ( .B(B[164]), .A(n40), .Z(n18003) );
  XNOR U18394 ( .A(n18011), .B(n18113), .Z(n18004) );
  XNOR U18395 ( .A(n18010), .B(n18008), .Z(n18113) );
  AND U18396 ( .A(n18114), .B(n18115), .Z(n18008) );
  NANDN U18397 ( .A(n18116), .B(n18117), .Z(n18115) );
  NAND U18398 ( .A(n18118), .B(n18119), .Z(n18117) );
  ANDN U18399 ( .B(B[165]), .A(n41), .Z(n18010) );
  XOR U18400 ( .A(n18017), .B(n18120), .Z(n18011) );
  XNOR U18401 ( .A(n18015), .B(n18018), .Z(n18120) );
  NAND U18402 ( .A(A[2]), .B(B[166]), .Z(n18018) );
  NANDN U18403 ( .A(n18121), .B(n18122), .Z(n18015) );
  AND U18404 ( .A(A[0]), .B(B[167]), .Z(n18122) );
  XNOR U18405 ( .A(n18020), .B(n18123), .Z(n18017) );
  NAND U18406 ( .A(A[0]), .B(B[168]), .Z(n18123) );
  NAND U18407 ( .A(B[167]), .B(A[1]), .Z(n18020) );
  NAND U18408 ( .A(n18124), .B(n18125), .Z(n417) );
  NANDN U18409 ( .A(n18126), .B(n18127), .Z(n18125) );
  OR U18410 ( .A(n18128), .B(n18129), .Z(n18127) );
  NAND U18411 ( .A(n18129), .B(n18128), .Z(n18124) );
  XOR U18412 ( .A(n419), .B(n418), .Z(\A1[165] ) );
  XOR U18413 ( .A(n18129), .B(n18130), .Z(n418) );
  XNOR U18414 ( .A(n18128), .B(n18126), .Z(n18130) );
  AND U18415 ( .A(n18131), .B(n18132), .Z(n18126) );
  NANDN U18416 ( .A(n18133), .B(n18134), .Z(n18132) );
  NANDN U18417 ( .A(n18135), .B(n18136), .Z(n18134) );
  NANDN U18418 ( .A(n18136), .B(n18135), .Z(n18131) );
  ANDN U18419 ( .B(B[152]), .A(n29), .Z(n18128) );
  XNOR U18420 ( .A(n18035), .B(n18137), .Z(n18129) );
  XNOR U18421 ( .A(n18034), .B(n18032), .Z(n18137) );
  AND U18422 ( .A(n18138), .B(n18139), .Z(n18032) );
  NANDN U18423 ( .A(n18140), .B(n18141), .Z(n18139) );
  OR U18424 ( .A(n18142), .B(n18143), .Z(n18141) );
  NAND U18425 ( .A(n18143), .B(n18142), .Z(n18138) );
  ANDN U18426 ( .B(B[153]), .A(n30), .Z(n18034) );
  XNOR U18427 ( .A(n18042), .B(n18144), .Z(n18035) );
  XNOR U18428 ( .A(n18041), .B(n18039), .Z(n18144) );
  AND U18429 ( .A(n18145), .B(n18146), .Z(n18039) );
  NANDN U18430 ( .A(n18147), .B(n18148), .Z(n18146) );
  NANDN U18431 ( .A(n18149), .B(n18150), .Z(n18148) );
  NANDN U18432 ( .A(n18150), .B(n18149), .Z(n18145) );
  ANDN U18433 ( .B(B[154]), .A(n31), .Z(n18041) );
  XNOR U18434 ( .A(n18049), .B(n18151), .Z(n18042) );
  XNOR U18435 ( .A(n18048), .B(n18046), .Z(n18151) );
  AND U18436 ( .A(n18152), .B(n18153), .Z(n18046) );
  NANDN U18437 ( .A(n18154), .B(n18155), .Z(n18153) );
  OR U18438 ( .A(n18156), .B(n18157), .Z(n18155) );
  NAND U18439 ( .A(n18157), .B(n18156), .Z(n18152) );
  ANDN U18440 ( .B(B[155]), .A(n32), .Z(n18048) );
  XNOR U18441 ( .A(n18056), .B(n18158), .Z(n18049) );
  XNOR U18442 ( .A(n18055), .B(n18053), .Z(n18158) );
  AND U18443 ( .A(n18159), .B(n18160), .Z(n18053) );
  NANDN U18444 ( .A(n18161), .B(n18162), .Z(n18160) );
  NANDN U18445 ( .A(n18163), .B(n18164), .Z(n18162) );
  NANDN U18446 ( .A(n18164), .B(n18163), .Z(n18159) );
  ANDN U18447 ( .B(B[156]), .A(n33), .Z(n18055) );
  XNOR U18448 ( .A(n18063), .B(n18165), .Z(n18056) );
  XNOR U18449 ( .A(n18062), .B(n18060), .Z(n18165) );
  AND U18450 ( .A(n18166), .B(n18167), .Z(n18060) );
  NANDN U18451 ( .A(n18168), .B(n18169), .Z(n18167) );
  OR U18452 ( .A(n18170), .B(n18171), .Z(n18169) );
  NAND U18453 ( .A(n18171), .B(n18170), .Z(n18166) );
  ANDN U18454 ( .B(B[157]), .A(n34), .Z(n18062) );
  XNOR U18455 ( .A(n18070), .B(n18172), .Z(n18063) );
  XNOR U18456 ( .A(n18069), .B(n18067), .Z(n18172) );
  AND U18457 ( .A(n18173), .B(n18174), .Z(n18067) );
  NANDN U18458 ( .A(n18175), .B(n18176), .Z(n18174) );
  NANDN U18459 ( .A(n18177), .B(n18178), .Z(n18176) );
  NANDN U18460 ( .A(n18178), .B(n18177), .Z(n18173) );
  ANDN U18461 ( .B(B[158]), .A(n35), .Z(n18069) );
  XNOR U18462 ( .A(n18077), .B(n18179), .Z(n18070) );
  XNOR U18463 ( .A(n18076), .B(n18074), .Z(n18179) );
  AND U18464 ( .A(n18180), .B(n18181), .Z(n18074) );
  NANDN U18465 ( .A(n18182), .B(n18183), .Z(n18181) );
  OR U18466 ( .A(n18184), .B(n18185), .Z(n18183) );
  NAND U18467 ( .A(n18185), .B(n18184), .Z(n18180) );
  ANDN U18468 ( .B(B[159]), .A(n36), .Z(n18076) );
  XNOR U18469 ( .A(n18084), .B(n18186), .Z(n18077) );
  XNOR U18470 ( .A(n18083), .B(n18081), .Z(n18186) );
  AND U18471 ( .A(n18187), .B(n18188), .Z(n18081) );
  NANDN U18472 ( .A(n18189), .B(n18190), .Z(n18188) );
  NANDN U18473 ( .A(n18191), .B(n18192), .Z(n18190) );
  NANDN U18474 ( .A(n18192), .B(n18191), .Z(n18187) );
  ANDN U18475 ( .B(B[160]), .A(n37), .Z(n18083) );
  XNOR U18476 ( .A(n18091), .B(n18193), .Z(n18084) );
  XNOR U18477 ( .A(n18090), .B(n18088), .Z(n18193) );
  AND U18478 ( .A(n18194), .B(n18195), .Z(n18088) );
  NANDN U18479 ( .A(n18196), .B(n18197), .Z(n18195) );
  OR U18480 ( .A(n18198), .B(n18199), .Z(n18197) );
  NAND U18481 ( .A(n18199), .B(n18198), .Z(n18194) );
  ANDN U18482 ( .B(B[161]), .A(n38), .Z(n18090) );
  XNOR U18483 ( .A(n18098), .B(n18200), .Z(n18091) );
  XNOR U18484 ( .A(n18097), .B(n18095), .Z(n18200) );
  AND U18485 ( .A(n18201), .B(n18202), .Z(n18095) );
  NANDN U18486 ( .A(n18203), .B(n18204), .Z(n18202) );
  NANDN U18487 ( .A(n18205), .B(n18206), .Z(n18204) );
  NANDN U18488 ( .A(n18206), .B(n18205), .Z(n18201) );
  ANDN U18489 ( .B(B[162]), .A(n39), .Z(n18097) );
  XNOR U18490 ( .A(n18105), .B(n18207), .Z(n18098) );
  XNOR U18491 ( .A(n18104), .B(n18102), .Z(n18207) );
  AND U18492 ( .A(n18208), .B(n18209), .Z(n18102) );
  NANDN U18493 ( .A(n18210), .B(n18211), .Z(n18209) );
  OR U18494 ( .A(n18212), .B(n18213), .Z(n18211) );
  NAND U18495 ( .A(n18213), .B(n18212), .Z(n18208) );
  ANDN U18496 ( .B(B[163]), .A(n40), .Z(n18104) );
  XNOR U18497 ( .A(n18112), .B(n18214), .Z(n18105) );
  XNOR U18498 ( .A(n18111), .B(n18109), .Z(n18214) );
  AND U18499 ( .A(n18215), .B(n18216), .Z(n18109) );
  NANDN U18500 ( .A(n18217), .B(n18218), .Z(n18216) );
  NAND U18501 ( .A(n18219), .B(n18220), .Z(n18218) );
  ANDN U18502 ( .B(B[164]), .A(n41), .Z(n18111) );
  XOR U18503 ( .A(n18118), .B(n18221), .Z(n18112) );
  XNOR U18504 ( .A(n18116), .B(n18119), .Z(n18221) );
  NAND U18505 ( .A(A[2]), .B(B[165]), .Z(n18119) );
  NANDN U18506 ( .A(n18222), .B(n18223), .Z(n18116) );
  AND U18507 ( .A(A[0]), .B(B[166]), .Z(n18223) );
  XNOR U18508 ( .A(n18121), .B(n18224), .Z(n18118) );
  NAND U18509 ( .A(A[0]), .B(B[167]), .Z(n18224) );
  NAND U18510 ( .A(B[166]), .B(A[1]), .Z(n18121) );
  NAND U18511 ( .A(n18225), .B(n18226), .Z(n419) );
  NANDN U18512 ( .A(n18227), .B(n18228), .Z(n18226) );
  OR U18513 ( .A(n18229), .B(n18230), .Z(n18228) );
  NAND U18514 ( .A(n18230), .B(n18229), .Z(n18225) );
  XOR U18515 ( .A(n421), .B(n420), .Z(\A1[164] ) );
  XOR U18516 ( .A(n18230), .B(n18231), .Z(n420) );
  XNOR U18517 ( .A(n18229), .B(n18227), .Z(n18231) );
  AND U18518 ( .A(n18232), .B(n18233), .Z(n18227) );
  NANDN U18519 ( .A(n18234), .B(n18235), .Z(n18233) );
  NANDN U18520 ( .A(n18236), .B(n18237), .Z(n18235) );
  NANDN U18521 ( .A(n18237), .B(n18236), .Z(n18232) );
  ANDN U18522 ( .B(B[151]), .A(n29), .Z(n18229) );
  XNOR U18523 ( .A(n18136), .B(n18238), .Z(n18230) );
  XNOR U18524 ( .A(n18135), .B(n18133), .Z(n18238) );
  AND U18525 ( .A(n18239), .B(n18240), .Z(n18133) );
  NANDN U18526 ( .A(n18241), .B(n18242), .Z(n18240) );
  OR U18527 ( .A(n18243), .B(n18244), .Z(n18242) );
  NAND U18528 ( .A(n18244), .B(n18243), .Z(n18239) );
  ANDN U18529 ( .B(B[152]), .A(n30), .Z(n18135) );
  XNOR U18530 ( .A(n18143), .B(n18245), .Z(n18136) );
  XNOR U18531 ( .A(n18142), .B(n18140), .Z(n18245) );
  AND U18532 ( .A(n18246), .B(n18247), .Z(n18140) );
  NANDN U18533 ( .A(n18248), .B(n18249), .Z(n18247) );
  NANDN U18534 ( .A(n18250), .B(n18251), .Z(n18249) );
  NANDN U18535 ( .A(n18251), .B(n18250), .Z(n18246) );
  ANDN U18536 ( .B(B[153]), .A(n31), .Z(n18142) );
  XNOR U18537 ( .A(n18150), .B(n18252), .Z(n18143) );
  XNOR U18538 ( .A(n18149), .B(n18147), .Z(n18252) );
  AND U18539 ( .A(n18253), .B(n18254), .Z(n18147) );
  NANDN U18540 ( .A(n18255), .B(n18256), .Z(n18254) );
  OR U18541 ( .A(n18257), .B(n18258), .Z(n18256) );
  NAND U18542 ( .A(n18258), .B(n18257), .Z(n18253) );
  ANDN U18543 ( .B(B[154]), .A(n32), .Z(n18149) );
  XNOR U18544 ( .A(n18157), .B(n18259), .Z(n18150) );
  XNOR U18545 ( .A(n18156), .B(n18154), .Z(n18259) );
  AND U18546 ( .A(n18260), .B(n18261), .Z(n18154) );
  NANDN U18547 ( .A(n18262), .B(n18263), .Z(n18261) );
  NANDN U18548 ( .A(n18264), .B(n18265), .Z(n18263) );
  NANDN U18549 ( .A(n18265), .B(n18264), .Z(n18260) );
  ANDN U18550 ( .B(B[155]), .A(n33), .Z(n18156) );
  XNOR U18551 ( .A(n18164), .B(n18266), .Z(n18157) );
  XNOR U18552 ( .A(n18163), .B(n18161), .Z(n18266) );
  AND U18553 ( .A(n18267), .B(n18268), .Z(n18161) );
  NANDN U18554 ( .A(n18269), .B(n18270), .Z(n18268) );
  OR U18555 ( .A(n18271), .B(n18272), .Z(n18270) );
  NAND U18556 ( .A(n18272), .B(n18271), .Z(n18267) );
  ANDN U18557 ( .B(B[156]), .A(n34), .Z(n18163) );
  XNOR U18558 ( .A(n18171), .B(n18273), .Z(n18164) );
  XNOR U18559 ( .A(n18170), .B(n18168), .Z(n18273) );
  AND U18560 ( .A(n18274), .B(n18275), .Z(n18168) );
  NANDN U18561 ( .A(n18276), .B(n18277), .Z(n18275) );
  NANDN U18562 ( .A(n18278), .B(n18279), .Z(n18277) );
  NANDN U18563 ( .A(n18279), .B(n18278), .Z(n18274) );
  ANDN U18564 ( .B(B[157]), .A(n35), .Z(n18170) );
  XNOR U18565 ( .A(n18178), .B(n18280), .Z(n18171) );
  XNOR U18566 ( .A(n18177), .B(n18175), .Z(n18280) );
  AND U18567 ( .A(n18281), .B(n18282), .Z(n18175) );
  NANDN U18568 ( .A(n18283), .B(n18284), .Z(n18282) );
  OR U18569 ( .A(n18285), .B(n18286), .Z(n18284) );
  NAND U18570 ( .A(n18286), .B(n18285), .Z(n18281) );
  ANDN U18571 ( .B(B[158]), .A(n36), .Z(n18177) );
  XNOR U18572 ( .A(n18185), .B(n18287), .Z(n18178) );
  XNOR U18573 ( .A(n18184), .B(n18182), .Z(n18287) );
  AND U18574 ( .A(n18288), .B(n18289), .Z(n18182) );
  NANDN U18575 ( .A(n18290), .B(n18291), .Z(n18289) );
  NANDN U18576 ( .A(n18292), .B(n18293), .Z(n18291) );
  NANDN U18577 ( .A(n18293), .B(n18292), .Z(n18288) );
  ANDN U18578 ( .B(B[159]), .A(n37), .Z(n18184) );
  XNOR U18579 ( .A(n18192), .B(n18294), .Z(n18185) );
  XNOR U18580 ( .A(n18191), .B(n18189), .Z(n18294) );
  AND U18581 ( .A(n18295), .B(n18296), .Z(n18189) );
  NANDN U18582 ( .A(n18297), .B(n18298), .Z(n18296) );
  OR U18583 ( .A(n18299), .B(n18300), .Z(n18298) );
  NAND U18584 ( .A(n18300), .B(n18299), .Z(n18295) );
  ANDN U18585 ( .B(B[160]), .A(n38), .Z(n18191) );
  XNOR U18586 ( .A(n18199), .B(n18301), .Z(n18192) );
  XNOR U18587 ( .A(n18198), .B(n18196), .Z(n18301) );
  AND U18588 ( .A(n18302), .B(n18303), .Z(n18196) );
  NANDN U18589 ( .A(n18304), .B(n18305), .Z(n18303) );
  NANDN U18590 ( .A(n18306), .B(n18307), .Z(n18305) );
  NANDN U18591 ( .A(n18307), .B(n18306), .Z(n18302) );
  ANDN U18592 ( .B(B[161]), .A(n39), .Z(n18198) );
  XNOR U18593 ( .A(n18206), .B(n18308), .Z(n18199) );
  XNOR U18594 ( .A(n18205), .B(n18203), .Z(n18308) );
  AND U18595 ( .A(n18309), .B(n18310), .Z(n18203) );
  NANDN U18596 ( .A(n18311), .B(n18312), .Z(n18310) );
  OR U18597 ( .A(n18313), .B(n18314), .Z(n18312) );
  NAND U18598 ( .A(n18314), .B(n18313), .Z(n18309) );
  ANDN U18599 ( .B(B[162]), .A(n40), .Z(n18205) );
  XNOR U18600 ( .A(n18213), .B(n18315), .Z(n18206) );
  XNOR U18601 ( .A(n18212), .B(n18210), .Z(n18315) );
  AND U18602 ( .A(n18316), .B(n18317), .Z(n18210) );
  NANDN U18603 ( .A(n18318), .B(n18319), .Z(n18317) );
  NAND U18604 ( .A(n18320), .B(n18321), .Z(n18319) );
  ANDN U18605 ( .B(B[163]), .A(n41), .Z(n18212) );
  XOR U18606 ( .A(n18219), .B(n18322), .Z(n18213) );
  XNOR U18607 ( .A(n18217), .B(n18220), .Z(n18322) );
  NAND U18608 ( .A(A[2]), .B(B[164]), .Z(n18220) );
  NANDN U18609 ( .A(n18323), .B(n18324), .Z(n18217) );
  AND U18610 ( .A(A[0]), .B(B[165]), .Z(n18324) );
  XNOR U18611 ( .A(n18222), .B(n18325), .Z(n18219) );
  NAND U18612 ( .A(A[0]), .B(B[166]), .Z(n18325) );
  NAND U18613 ( .A(B[165]), .B(A[1]), .Z(n18222) );
  NAND U18614 ( .A(n18326), .B(n18327), .Z(n421) );
  NANDN U18615 ( .A(n18328), .B(n18329), .Z(n18327) );
  OR U18616 ( .A(n18330), .B(n18331), .Z(n18329) );
  NAND U18617 ( .A(n18331), .B(n18330), .Z(n18326) );
  XOR U18618 ( .A(n423), .B(n422), .Z(\A1[163] ) );
  XOR U18619 ( .A(n18331), .B(n18332), .Z(n422) );
  XNOR U18620 ( .A(n18330), .B(n18328), .Z(n18332) );
  AND U18621 ( .A(n18333), .B(n18334), .Z(n18328) );
  NANDN U18622 ( .A(n18335), .B(n18336), .Z(n18334) );
  NANDN U18623 ( .A(n18337), .B(n18338), .Z(n18336) );
  NANDN U18624 ( .A(n18338), .B(n18337), .Z(n18333) );
  ANDN U18625 ( .B(B[150]), .A(n29), .Z(n18330) );
  XNOR U18626 ( .A(n18237), .B(n18339), .Z(n18331) );
  XNOR U18627 ( .A(n18236), .B(n18234), .Z(n18339) );
  AND U18628 ( .A(n18340), .B(n18341), .Z(n18234) );
  NANDN U18629 ( .A(n18342), .B(n18343), .Z(n18341) );
  OR U18630 ( .A(n18344), .B(n18345), .Z(n18343) );
  NAND U18631 ( .A(n18345), .B(n18344), .Z(n18340) );
  ANDN U18632 ( .B(B[151]), .A(n30), .Z(n18236) );
  XNOR U18633 ( .A(n18244), .B(n18346), .Z(n18237) );
  XNOR U18634 ( .A(n18243), .B(n18241), .Z(n18346) );
  AND U18635 ( .A(n18347), .B(n18348), .Z(n18241) );
  NANDN U18636 ( .A(n18349), .B(n18350), .Z(n18348) );
  NANDN U18637 ( .A(n18351), .B(n18352), .Z(n18350) );
  NANDN U18638 ( .A(n18352), .B(n18351), .Z(n18347) );
  ANDN U18639 ( .B(B[152]), .A(n31), .Z(n18243) );
  XNOR U18640 ( .A(n18251), .B(n18353), .Z(n18244) );
  XNOR U18641 ( .A(n18250), .B(n18248), .Z(n18353) );
  AND U18642 ( .A(n18354), .B(n18355), .Z(n18248) );
  NANDN U18643 ( .A(n18356), .B(n18357), .Z(n18355) );
  OR U18644 ( .A(n18358), .B(n18359), .Z(n18357) );
  NAND U18645 ( .A(n18359), .B(n18358), .Z(n18354) );
  ANDN U18646 ( .B(B[153]), .A(n32), .Z(n18250) );
  XNOR U18647 ( .A(n18258), .B(n18360), .Z(n18251) );
  XNOR U18648 ( .A(n18257), .B(n18255), .Z(n18360) );
  AND U18649 ( .A(n18361), .B(n18362), .Z(n18255) );
  NANDN U18650 ( .A(n18363), .B(n18364), .Z(n18362) );
  NANDN U18651 ( .A(n18365), .B(n18366), .Z(n18364) );
  NANDN U18652 ( .A(n18366), .B(n18365), .Z(n18361) );
  ANDN U18653 ( .B(B[154]), .A(n33), .Z(n18257) );
  XNOR U18654 ( .A(n18265), .B(n18367), .Z(n18258) );
  XNOR U18655 ( .A(n18264), .B(n18262), .Z(n18367) );
  AND U18656 ( .A(n18368), .B(n18369), .Z(n18262) );
  NANDN U18657 ( .A(n18370), .B(n18371), .Z(n18369) );
  OR U18658 ( .A(n18372), .B(n18373), .Z(n18371) );
  NAND U18659 ( .A(n18373), .B(n18372), .Z(n18368) );
  ANDN U18660 ( .B(B[155]), .A(n34), .Z(n18264) );
  XNOR U18661 ( .A(n18272), .B(n18374), .Z(n18265) );
  XNOR U18662 ( .A(n18271), .B(n18269), .Z(n18374) );
  AND U18663 ( .A(n18375), .B(n18376), .Z(n18269) );
  NANDN U18664 ( .A(n18377), .B(n18378), .Z(n18376) );
  NANDN U18665 ( .A(n18379), .B(n18380), .Z(n18378) );
  NANDN U18666 ( .A(n18380), .B(n18379), .Z(n18375) );
  ANDN U18667 ( .B(B[156]), .A(n35), .Z(n18271) );
  XNOR U18668 ( .A(n18279), .B(n18381), .Z(n18272) );
  XNOR U18669 ( .A(n18278), .B(n18276), .Z(n18381) );
  AND U18670 ( .A(n18382), .B(n18383), .Z(n18276) );
  NANDN U18671 ( .A(n18384), .B(n18385), .Z(n18383) );
  OR U18672 ( .A(n18386), .B(n18387), .Z(n18385) );
  NAND U18673 ( .A(n18387), .B(n18386), .Z(n18382) );
  ANDN U18674 ( .B(B[157]), .A(n36), .Z(n18278) );
  XNOR U18675 ( .A(n18286), .B(n18388), .Z(n18279) );
  XNOR U18676 ( .A(n18285), .B(n18283), .Z(n18388) );
  AND U18677 ( .A(n18389), .B(n18390), .Z(n18283) );
  NANDN U18678 ( .A(n18391), .B(n18392), .Z(n18390) );
  NANDN U18679 ( .A(n18393), .B(n18394), .Z(n18392) );
  NANDN U18680 ( .A(n18394), .B(n18393), .Z(n18389) );
  ANDN U18681 ( .B(B[158]), .A(n37), .Z(n18285) );
  XNOR U18682 ( .A(n18293), .B(n18395), .Z(n18286) );
  XNOR U18683 ( .A(n18292), .B(n18290), .Z(n18395) );
  AND U18684 ( .A(n18396), .B(n18397), .Z(n18290) );
  NANDN U18685 ( .A(n18398), .B(n18399), .Z(n18397) );
  OR U18686 ( .A(n18400), .B(n18401), .Z(n18399) );
  NAND U18687 ( .A(n18401), .B(n18400), .Z(n18396) );
  ANDN U18688 ( .B(B[159]), .A(n38), .Z(n18292) );
  XNOR U18689 ( .A(n18300), .B(n18402), .Z(n18293) );
  XNOR U18690 ( .A(n18299), .B(n18297), .Z(n18402) );
  AND U18691 ( .A(n18403), .B(n18404), .Z(n18297) );
  NANDN U18692 ( .A(n18405), .B(n18406), .Z(n18404) );
  NANDN U18693 ( .A(n18407), .B(n18408), .Z(n18406) );
  NANDN U18694 ( .A(n18408), .B(n18407), .Z(n18403) );
  ANDN U18695 ( .B(B[160]), .A(n39), .Z(n18299) );
  XNOR U18696 ( .A(n18307), .B(n18409), .Z(n18300) );
  XNOR U18697 ( .A(n18306), .B(n18304), .Z(n18409) );
  AND U18698 ( .A(n18410), .B(n18411), .Z(n18304) );
  NANDN U18699 ( .A(n18412), .B(n18413), .Z(n18411) );
  OR U18700 ( .A(n18414), .B(n18415), .Z(n18413) );
  NAND U18701 ( .A(n18415), .B(n18414), .Z(n18410) );
  ANDN U18702 ( .B(B[161]), .A(n40), .Z(n18306) );
  XNOR U18703 ( .A(n18314), .B(n18416), .Z(n18307) );
  XNOR U18704 ( .A(n18313), .B(n18311), .Z(n18416) );
  AND U18705 ( .A(n18417), .B(n18418), .Z(n18311) );
  NANDN U18706 ( .A(n18419), .B(n18420), .Z(n18418) );
  NAND U18707 ( .A(n18421), .B(n18422), .Z(n18420) );
  ANDN U18708 ( .B(B[162]), .A(n41), .Z(n18313) );
  XOR U18709 ( .A(n18320), .B(n18423), .Z(n18314) );
  XNOR U18710 ( .A(n18318), .B(n18321), .Z(n18423) );
  NAND U18711 ( .A(A[2]), .B(B[163]), .Z(n18321) );
  NANDN U18712 ( .A(n18424), .B(n18425), .Z(n18318) );
  AND U18713 ( .A(A[0]), .B(B[164]), .Z(n18425) );
  XNOR U18714 ( .A(n18323), .B(n18426), .Z(n18320) );
  NAND U18715 ( .A(A[0]), .B(B[165]), .Z(n18426) );
  NAND U18716 ( .A(B[164]), .B(A[1]), .Z(n18323) );
  NAND U18717 ( .A(n18427), .B(n18428), .Z(n423) );
  NANDN U18718 ( .A(n18429), .B(n18430), .Z(n18428) );
  OR U18719 ( .A(n18431), .B(n18432), .Z(n18430) );
  NAND U18720 ( .A(n18432), .B(n18431), .Z(n18427) );
  XOR U18721 ( .A(n425), .B(n424), .Z(\A1[162] ) );
  XOR U18722 ( .A(n18432), .B(n18433), .Z(n424) );
  XNOR U18723 ( .A(n18431), .B(n18429), .Z(n18433) );
  AND U18724 ( .A(n18434), .B(n18435), .Z(n18429) );
  NANDN U18725 ( .A(n18436), .B(n18437), .Z(n18435) );
  NANDN U18726 ( .A(n18438), .B(n18439), .Z(n18437) );
  NANDN U18727 ( .A(n18439), .B(n18438), .Z(n18434) );
  ANDN U18728 ( .B(B[149]), .A(n29), .Z(n18431) );
  XNOR U18729 ( .A(n18338), .B(n18440), .Z(n18432) );
  XNOR U18730 ( .A(n18337), .B(n18335), .Z(n18440) );
  AND U18731 ( .A(n18441), .B(n18442), .Z(n18335) );
  NANDN U18732 ( .A(n18443), .B(n18444), .Z(n18442) );
  OR U18733 ( .A(n18445), .B(n18446), .Z(n18444) );
  NAND U18734 ( .A(n18446), .B(n18445), .Z(n18441) );
  ANDN U18735 ( .B(B[150]), .A(n30), .Z(n18337) );
  XNOR U18736 ( .A(n18345), .B(n18447), .Z(n18338) );
  XNOR U18737 ( .A(n18344), .B(n18342), .Z(n18447) );
  AND U18738 ( .A(n18448), .B(n18449), .Z(n18342) );
  NANDN U18739 ( .A(n18450), .B(n18451), .Z(n18449) );
  NANDN U18740 ( .A(n18452), .B(n18453), .Z(n18451) );
  NANDN U18741 ( .A(n18453), .B(n18452), .Z(n18448) );
  ANDN U18742 ( .B(B[151]), .A(n31), .Z(n18344) );
  XNOR U18743 ( .A(n18352), .B(n18454), .Z(n18345) );
  XNOR U18744 ( .A(n18351), .B(n18349), .Z(n18454) );
  AND U18745 ( .A(n18455), .B(n18456), .Z(n18349) );
  NANDN U18746 ( .A(n18457), .B(n18458), .Z(n18456) );
  OR U18747 ( .A(n18459), .B(n18460), .Z(n18458) );
  NAND U18748 ( .A(n18460), .B(n18459), .Z(n18455) );
  ANDN U18749 ( .B(B[152]), .A(n32), .Z(n18351) );
  XNOR U18750 ( .A(n18359), .B(n18461), .Z(n18352) );
  XNOR U18751 ( .A(n18358), .B(n18356), .Z(n18461) );
  AND U18752 ( .A(n18462), .B(n18463), .Z(n18356) );
  NANDN U18753 ( .A(n18464), .B(n18465), .Z(n18463) );
  NANDN U18754 ( .A(n18466), .B(n18467), .Z(n18465) );
  NANDN U18755 ( .A(n18467), .B(n18466), .Z(n18462) );
  ANDN U18756 ( .B(B[153]), .A(n33), .Z(n18358) );
  XNOR U18757 ( .A(n18366), .B(n18468), .Z(n18359) );
  XNOR U18758 ( .A(n18365), .B(n18363), .Z(n18468) );
  AND U18759 ( .A(n18469), .B(n18470), .Z(n18363) );
  NANDN U18760 ( .A(n18471), .B(n18472), .Z(n18470) );
  OR U18761 ( .A(n18473), .B(n18474), .Z(n18472) );
  NAND U18762 ( .A(n18474), .B(n18473), .Z(n18469) );
  ANDN U18763 ( .B(B[154]), .A(n34), .Z(n18365) );
  XNOR U18764 ( .A(n18373), .B(n18475), .Z(n18366) );
  XNOR U18765 ( .A(n18372), .B(n18370), .Z(n18475) );
  AND U18766 ( .A(n18476), .B(n18477), .Z(n18370) );
  NANDN U18767 ( .A(n18478), .B(n18479), .Z(n18477) );
  NANDN U18768 ( .A(n18480), .B(n18481), .Z(n18479) );
  NANDN U18769 ( .A(n18481), .B(n18480), .Z(n18476) );
  ANDN U18770 ( .B(B[155]), .A(n35), .Z(n18372) );
  XNOR U18771 ( .A(n18380), .B(n18482), .Z(n18373) );
  XNOR U18772 ( .A(n18379), .B(n18377), .Z(n18482) );
  AND U18773 ( .A(n18483), .B(n18484), .Z(n18377) );
  NANDN U18774 ( .A(n18485), .B(n18486), .Z(n18484) );
  OR U18775 ( .A(n18487), .B(n18488), .Z(n18486) );
  NAND U18776 ( .A(n18488), .B(n18487), .Z(n18483) );
  ANDN U18777 ( .B(B[156]), .A(n36), .Z(n18379) );
  XNOR U18778 ( .A(n18387), .B(n18489), .Z(n18380) );
  XNOR U18779 ( .A(n18386), .B(n18384), .Z(n18489) );
  AND U18780 ( .A(n18490), .B(n18491), .Z(n18384) );
  NANDN U18781 ( .A(n18492), .B(n18493), .Z(n18491) );
  NANDN U18782 ( .A(n18494), .B(n18495), .Z(n18493) );
  NANDN U18783 ( .A(n18495), .B(n18494), .Z(n18490) );
  ANDN U18784 ( .B(B[157]), .A(n37), .Z(n18386) );
  XNOR U18785 ( .A(n18394), .B(n18496), .Z(n18387) );
  XNOR U18786 ( .A(n18393), .B(n18391), .Z(n18496) );
  AND U18787 ( .A(n18497), .B(n18498), .Z(n18391) );
  NANDN U18788 ( .A(n18499), .B(n18500), .Z(n18498) );
  OR U18789 ( .A(n18501), .B(n18502), .Z(n18500) );
  NAND U18790 ( .A(n18502), .B(n18501), .Z(n18497) );
  ANDN U18791 ( .B(B[158]), .A(n38), .Z(n18393) );
  XNOR U18792 ( .A(n18401), .B(n18503), .Z(n18394) );
  XNOR U18793 ( .A(n18400), .B(n18398), .Z(n18503) );
  AND U18794 ( .A(n18504), .B(n18505), .Z(n18398) );
  NANDN U18795 ( .A(n18506), .B(n18507), .Z(n18505) );
  NANDN U18796 ( .A(n18508), .B(n18509), .Z(n18507) );
  NANDN U18797 ( .A(n18509), .B(n18508), .Z(n18504) );
  ANDN U18798 ( .B(B[159]), .A(n39), .Z(n18400) );
  XNOR U18799 ( .A(n18408), .B(n18510), .Z(n18401) );
  XNOR U18800 ( .A(n18407), .B(n18405), .Z(n18510) );
  AND U18801 ( .A(n18511), .B(n18512), .Z(n18405) );
  NANDN U18802 ( .A(n18513), .B(n18514), .Z(n18512) );
  OR U18803 ( .A(n18515), .B(n18516), .Z(n18514) );
  NAND U18804 ( .A(n18516), .B(n18515), .Z(n18511) );
  ANDN U18805 ( .B(B[160]), .A(n40), .Z(n18407) );
  XNOR U18806 ( .A(n18415), .B(n18517), .Z(n18408) );
  XNOR U18807 ( .A(n18414), .B(n18412), .Z(n18517) );
  AND U18808 ( .A(n18518), .B(n18519), .Z(n18412) );
  NANDN U18809 ( .A(n18520), .B(n18521), .Z(n18519) );
  NAND U18810 ( .A(n18522), .B(n18523), .Z(n18521) );
  ANDN U18811 ( .B(B[161]), .A(n41), .Z(n18414) );
  XOR U18812 ( .A(n18421), .B(n18524), .Z(n18415) );
  XNOR U18813 ( .A(n18419), .B(n18422), .Z(n18524) );
  NAND U18814 ( .A(A[2]), .B(B[162]), .Z(n18422) );
  NANDN U18815 ( .A(n18525), .B(n18526), .Z(n18419) );
  AND U18816 ( .A(A[0]), .B(B[163]), .Z(n18526) );
  XNOR U18817 ( .A(n18424), .B(n18527), .Z(n18421) );
  NAND U18818 ( .A(A[0]), .B(B[164]), .Z(n18527) );
  NAND U18819 ( .A(B[163]), .B(A[1]), .Z(n18424) );
  NAND U18820 ( .A(n18528), .B(n18529), .Z(n425) );
  NANDN U18821 ( .A(n18530), .B(n18531), .Z(n18529) );
  OR U18822 ( .A(n18532), .B(n18533), .Z(n18531) );
  NAND U18823 ( .A(n18533), .B(n18532), .Z(n18528) );
  XOR U18824 ( .A(n427), .B(n426), .Z(\A1[161] ) );
  XOR U18825 ( .A(n18533), .B(n18534), .Z(n426) );
  XNOR U18826 ( .A(n18532), .B(n18530), .Z(n18534) );
  AND U18827 ( .A(n18535), .B(n18536), .Z(n18530) );
  NANDN U18828 ( .A(n18537), .B(n18538), .Z(n18536) );
  NANDN U18829 ( .A(n18539), .B(n18540), .Z(n18538) );
  NANDN U18830 ( .A(n18540), .B(n18539), .Z(n18535) );
  ANDN U18831 ( .B(B[148]), .A(n29), .Z(n18532) );
  XNOR U18832 ( .A(n18439), .B(n18541), .Z(n18533) );
  XNOR U18833 ( .A(n18438), .B(n18436), .Z(n18541) );
  AND U18834 ( .A(n18542), .B(n18543), .Z(n18436) );
  NANDN U18835 ( .A(n18544), .B(n18545), .Z(n18543) );
  OR U18836 ( .A(n18546), .B(n18547), .Z(n18545) );
  NAND U18837 ( .A(n18547), .B(n18546), .Z(n18542) );
  ANDN U18838 ( .B(B[149]), .A(n30), .Z(n18438) );
  XNOR U18839 ( .A(n18446), .B(n18548), .Z(n18439) );
  XNOR U18840 ( .A(n18445), .B(n18443), .Z(n18548) );
  AND U18841 ( .A(n18549), .B(n18550), .Z(n18443) );
  NANDN U18842 ( .A(n18551), .B(n18552), .Z(n18550) );
  NANDN U18843 ( .A(n18553), .B(n18554), .Z(n18552) );
  NANDN U18844 ( .A(n18554), .B(n18553), .Z(n18549) );
  ANDN U18845 ( .B(B[150]), .A(n31), .Z(n18445) );
  XNOR U18846 ( .A(n18453), .B(n18555), .Z(n18446) );
  XNOR U18847 ( .A(n18452), .B(n18450), .Z(n18555) );
  AND U18848 ( .A(n18556), .B(n18557), .Z(n18450) );
  NANDN U18849 ( .A(n18558), .B(n18559), .Z(n18557) );
  OR U18850 ( .A(n18560), .B(n18561), .Z(n18559) );
  NAND U18851 ( .A(n18561), .B(n18560), .Z(n18556) );
  ANDN U18852 ( .B(B[151]), .A(n32), .Z(n18452) );
  XNOR U18853 ( .A(n18460), .B(n18562), .Z(n18453) );
  XNOR U18854 ( .A(n18459), .B(n18457), .Z(n18562) );
  AND U18855 ( .A(n18563), .B(n18564), .Z(n18457) );
  NANDN U18856 ( .A(n18565), .B(n18566), .Z(n18564) );
  NANDN U18857 ( .A(n18567), .B(n18568), .Z(n18566) );
  NANDN U18858 ( .A(n18568), .B(n18567), .Z(n18563) );
  ANDN U18859 ( .B(B[152]), .A(n33), .Z(n18459) );
  XNOR U18860 ( .A(n18467), .B(n18569), .Z(n18460) );
  XNOR U18861 ( .A(n18466), .B(n18464), .Z(n18569) );
  AND U18862 ( .A(n18570), .B(n18571), .Z(n18464) );
  NANDN U18863 ( .A(n18572), .B(n18573), .Z(n18571) );
  OR U18864 ( .A(n18574), .B(n18575), .Z(n18573) );
  NAND U18865 ( .A(n18575), .B(n18574), .Z(n18570) );
  ANDN U18866 ( .B(B[153]), .A(n34), .Z(n18466) );
  XNOR U18867 ( .A(n18474), .B(n18576), .Z(n18467) );
  XNOR U18868 ( .A(n18473), .B(n18471), .Z(n18576) );
  AND U18869 ( .A(n18577), .B(n18578), .Z(n18471) );
  NANDN U18870 ( .A(n18579), .B(n18580), .Z(n18578) );
  NANDN U18871 ( .A(n18581), .B(n18582), .Z(n18580) );
  NANDN U18872 ( .A(n18582), .B(n18581), .Z(n18577) );
  ANDN U18873 ( .B(B[154]), .A(n35), .Z(n18473) );
  XNOR U18874 ( .A(n18481), .B(n18583), .Z(n18474) );
  XNOR U18875 ( .A(n18480), .B(n18478), .Z(n18583) );
  AND U18876 ( .A(n18584), .B(n18585), .Z(n18478) );
  NANDN U18877 ( .A(n18586), .B(n18587), .Z(n18585) );
  OR U18878 ( .A(n18588), .B(n18589), .Z(n18587) );
  NAND U18879 ( .A(n18589), .B(n18588), .Z(n18584) );
  ANDN U18880 ( .B(B[155]), .A(n36), .Z(n18480) );
  XNOR U18881 ( .A(n18488), .B(n18590), .Z(n18481) );
  XNOR U18882 ( .A(n18487), .B(n18485), .Z(n18590) );
  AND U18883 ( .A(n18591), .B(n18592), .Z(n18485) );
  NANDN U18884 ( .A(n18593), .B(n18594), .Z(n18592) );
  NANDN U18885 ( .A(n18595), .B(n18596), .Z(n18594) );
  NANDN U18886 ( .A(n18596), .B(n18595), .Z(n18591) );
  ANDN U18887 ( .B(B[156]), .A(n37), .Z(n18487) );
  XNOR U18888 ( .A(n18495), .B(n18597), .Z(n18488) );
  XNOR U18889 ( .A(n18494), .B(n18492), .Z(n18597) );
  AND U18890 ( .A(n18598), .B(n18599), .Z(n18492) );
  NANDN U18891 ( .A(n18600), .B(n18601), .Z(n18599) );
  OR U18892 ( .A(n18602), .B(n18603), .Z(n18601) );
  NAND U18893 ( .A(n18603), .B(n18602), .Z(n18598) );
  ANDN U18894 ( .B(B[157]), .A(n38), .Z(n18494) );
  XNOR U18895 ( .A(n18502), .B(n18604), .Z(n18495) );
  XNOR U18896 ( .A(n18501), .B(n18499), .Z(n18604) );
  AND U18897 ( .A(n18605), .B(n18606), .Z(n18499) );
  NANDN U18898 ( .A(n18607), .B(n18608), .Z(n18606) );
  NANDN U18899 ( .A(n18609), .B(n18610), .Z(n18608) );
  NANDN U18900 ( .A(n18610), .B(n18609), .Z(n18605) );
  ANDN U18901 ( .B(B[158]), .A(n39), .Z(n18501) );
  XNOR U18902 ( .A(n18509), .B(n18611), .Z(n18502) );
  XNOR U18903 ( .A(n18508), .B(n18506), .Z(n18611) );
  AND U18904 ( .A(n18612), .B(n18613), .Z(n18506) );
  NANDN U18905 ( .A(n18614), .B(n18615), .Z(n18613) );
  OR U18906 ( .A(n18616), .B(n18617), .Z(n18615) );
  NAND U18907 ( .A(n18617), .B(n18616), .Z(n18612) );
  ANDN U18908 ( .B(B[159]), .A(n40), .Z(n18508) );
  XNOR U18909 ( .A(n18516), .B(n18618), .Z(n18509) );
  XNOR U18910 ( .A(n18515), .B(n18513), .Z(n18618) );
  AND U18911 ( .A(n18619), .B(n18620), .Z(n18513) );
  NANDN U18912 ( .A(n18621), .B(n18622), .Z(n18620) );
  NAND U18913 ( .A(n18623), .B(n18624), .Z(n18622) );
  ANDN U18914 ( .B(B[160]), .A(n41), .Z(n18515) );
  XOR U18915 ( .A(n18522), .B(n18625), .Z(n18516) );
  XNOR U18916 ( .A(n18520), .B(n18523), .Z(n18625) );
  NAND U18917 ( .A(A[2]), .B(B[161]), .Z(n18523) );
  NANDN U18918 ( .A(n18626), .B(n18627), .Z(n18520) );
  AND U18919 ( .A(A[0]), .B(B[162]), .Z(n18627) );
  XNOR U18920 ( .A(n18525), .B(n18628), .Z(n18522) );
  NAND U18921 ( .A(A[0]), .B(B[163]), .Z(n18628) );
  NAND U18922 ( .A(B[162]), .B(A[1]), .Z(n18525) );
  NAND U18923 ( .A(n18629), .B(n18630), .Z(n427) );
  NANDN U18924 ( .A(n18631), .B(n18632), .Z(n18630) );
  OR U18925 ( .A(n18633), .B(n18634), .Z(n18632) );
  NAND U18926 ( .A(n18634), .B(n18633), .Z(n18629) );
  XOR U18927 ( .A(n429), .B(n428), .Z(\A1[160] ) );
  XOR U18928 ( .A(n18634), .B(n18635), .Z(n428) );
  XNOR U18929 ( .A(n18633), .B(n18631), .Z(n18635) );
  AND U18930 ( .A(n18636), .B(n18637), .Z(n18631) );
  NANDN U18931 ( .A(n18638), .B(n18639), .Z(n18637) );
  NANDN U18932 ( .A(n18640), .B(n18641), .Z(n18639) );
  NANDN U18933 ( .A(n18641), .B(n18640), .Z(n18636) );
  ANDN U18934 ( .B(B[147]), .A(n29), .Z(n18633) );
  XNOR U18935 ( .A(n18540), .B(n18642), .Z(n18634) );
  XNOR U18936 ( .A(n18539), .B(n18537), .Z(n18642) );
  AND U18937 ( .A(n18643), .B(n18644), .Z(n18537) );
  NANDN U18938 ( .A(n18645), .B(n18646), .Z(n18644) );
  OR U18939 ( .A(n18647), .B(n18648), .Z(n18646) );
  NAND U18940 ( .A(n18648), .B(n18647), .Z(n18643) );
  ANDN U18941 ( .B(B[148]), .A(n30), .Z(n18539) );
  XNOR U18942 ( .A(n18547), .B(n18649), .Z(n18540) );
  XNOR U18943 ( .A(n18546), .B(n18544), .Z(n18649) );
  AND U18944 ( .A(n18650), .B(n18651), .Z(n18544) );
  NANDN U18945 ( .A(n18652), .B(n18653), .Z(n18651) );
  NANDN U18946 ( .A(n18654), .B(n18655), .Z(n18653) );
  NANDN U18947 ( .A(n18655), .B(n18654), .Z(n18650) );
  ANDN U18948 ( .B(B[149]), .A(n31), .Z(n18546) );
  XNOR U18949 ( .A(n18554), .B(n18656), .Z(n18547) );
  XNOR U18950 ( .A(n18553), .B(n18551), .Z(n18656) );
  AND U18951 ( .A(n18657), .B(n18658), .Z(n18551) );
  NANDN U18952 ( .A(n18659), .B(n18660), .Z(n18658) );
  OR U18953 ( .A(n18661), .B(n18662), .Z(n18660) );
  NAND U18954 ( .A(n18662), .B(n18661), .Z(n18657) );
  ANDN U18955 ( .B(B[150]), .A(n32), .Z(n18553) );
  XNOR U18956 ( .A(n18561), .B(n18663), .Z(n18554) );
  XNOR U18957 ( .A(n18560), .B(n18558), .Z(n18663) );
  AND U18958 ( .A(n18664), .B(n18665), .Z(n18558) );
  NANDN U18959 ( .A(n18666), .B(n18667), .Z(n18665) );
  NANDN U18960 ( .A(n18668), .B(n18669), .Z(n18667) );
  NANDN U18961 ( .A(n18669), .B(n18668), .Z(n18664) );
  ANDN U18962 ( .B(B[151]), .A(n33), .Z(n18560) );
  XNOR U18963 ( .A(n18568), .B(n18670), .Z(n18561) );
  XNOR U18964 ( .A(n18567), .B(n18565), .Z(n18670) );
  AND U18965 ( .A(n18671), .B(n18672), .Z(n18565) );
  NANDN U18966 ( .A(n18673), .B(n18674), .Z(n18672) );
  OR U18967 ( .A(n18675), .B(n18676), .Z(n18674) );
  NAND U18968 ( .A(n18676), .B(n18675), .Z(n18671) );
  ANDN U18969 ( .B(B[152]), .A(n34), .Z(n18567) );
  XNOR U18970 ( .A(n18575), .B(n18677), .Z(n18568) );
  XNOR U18971 ( .A(n18574), .B(n18572), .Z(n18677) );
  AND U18972 ( .A(n18678), .B(n18679), .Z(n18572) );
  NANDN U18973 ( .A(n18680), .B(n18681), .Z(n18679) );
  NANDN U18974 ( .A(n18682), .B(n18683), .Z(n18681) );
  NANDN U18975 ( .A(n18683), .B(n18682), .Z(n18678) );
  ANDN U18976 ( .B(B[153]), .A(n35), .Z(n18574) );
  XNOR U18977 ( .A(n18582), .B(n18684), .Z(n18575) );
  XNOR U18978 ( .A(n18581), .B(n18579), .Z(n18684) );
  AND U18979 ( .A(n18685), .B(n18686), .Z(n18579) );
  NANDN U18980 ( .A(n18687), .B(n18688), .Z(n18686) );
  OR U18981 ( .A(n18689), .B(n18690), .Z(n18688) );
  NAND U18982 ( .A(n18690), .B(n18689), .Z(n18685) );
  ANDN U18983 ( .B(B[154]), .A(n36), .Z(n18581) );
  XNOR U18984 ( .A(n18589), .B(n18691), .Z(n18582) );
  XNOR U18985 ( .A(n18588), .B(n18586), .Z(n18691) );
  AND U18986 ( .A(n18692), .B(n18693), .Z(n18586) );
  NANDN U18987 ( .A(n18694), .B(n18695), .Z(n18693) );
  NANDN U18988 ( .A(n18696), .B(n18697), .Z(n18695) );
  NANDN U18989 ( .A(n18697), .B(n18696), .Z(n18692) );
  ANDN U18990 ( .B(B[155]), .A(n37), .Z(n18588) );
  XNOR U18991 ( .A(n18596), .B(n18698), .Z(n18589) );
  XNOR U18992 ( .A(n18595), .B(n18593), .Z(n18698) );
  AND U18993 ( .A(n18699), .B(n18700), .Z(n18593) );
  NANDN U18994 ( .A(n18701), .B(n18702), .Z(n18700) );
  OR U18995 ( .A(n18703), .B(n18704), .Z(n18702) );
  NAND U18996 ( .A(n18704), .B(n18703), .Z(n18699) );
  ANDN U18997 ( .B(B[156]), .A(n38), .Z(n18595) );
  XNOR U18998 ( .A(n18603), .B(n18705), .Z(n18596) );
  XNOR U18999 ( .A(n18602), .B(n18600), .Z(n18705) );
  AND U19000 ( .A(n18706), .B(n18707), .Z(n18600) );
  NANDN U19001 ( .A(n18708), .B(n18709), .Z(n18707) );
  NANDN U19002 ( .A(n18710), .B(n18711), .Z(n18709) );
  NANDN U19003 ( .A(n18711), .B(n18710), .Z(n18706) );
  ANDN U19004 ( .B(B[157]), .A(n39), .Z(n18602) );
  XNOR U19005 ( .A(n18610), .B(n18712), .Z(n18603) );
  XNOR U19006 ( .A(n18609), .B(n18607), .Z(n18712) );
  AND U19007 ( .A(n18713), .B(n18714), .Z(n18607) );
  NANDN U19008 ( .A(n18715), .B(n18716), .Z(n18714) );
  OR U19009 ( .A(n18717), .B(n18718), .Z(n18716) );
  NAND U19010 ( .A(n18718), .B(n18717), .Z(n18713) );
  ANDN U19011 ( .B(B[158]), .A(n40), .Z(n18609) );
  XNOR U19012 ( .A(n18617), .B(n18719), .Z(n18610) );
  XNOR U19013 ( .A(n18616), .B(n18614), .Z(n18719) );
  AND U19014 ( .A(n18720), .B(n18721), .Z(n18614) );
  NANDN U19015 ( .A(n18722), .B(n18723), .Z(n18721) );
  NAND U19016 ( .A(n18724), .B(n18725), .Z(n18723) );
  ANDN U19017 ( .B(B[159]), .A(n41), .Z(n18616) );
  XOR U19018 ( .A(n18623), .B(n18726), .Z(n18617) );
  XNOR U19019 ( .A(n18621), .B(n18624), .Z(n18726) );
  NAND U19020 ( .A(A[2]), .B(B[160]), .Z(n18624) );
  NANDN U19021 ( .A(n18727), .B(n18728), .Z(n18621) );
  AND U19022 ( .A(A[0]), .B(B[161]), .Z(n18728) );
  XNOR U19023 ( .A(n18626), .B(n18729), .Z(n18623) );
  NAND U19024 ( .A(A[0]), .B(B[162]), .Z(n18729) );
  NAND U19025 ( .A(B[161]), .B(A[1]), .Z(n18626) );
  NAND U19026 ( .A(n18730), .B(n18731), .Z(n429) );
  NANDN U19027 ( .A(n18732), .B(n18733), .Z(n18731) );
  OR U19028 ( .A(n18734), .B(n18735), .Z(n18733) );
  NAND U19029 ( .A(n18735), .B(n18734), .Z(n18730) );
  XOR U19030 ( .A(n411), .B(n410), .Z(\A1[15] ) );
  XOR U19031 ( .A(n17725), .B(n18736), .Z(n410) );
  XNOR U19032 ( .A(n17724), .B(n17722), .Z(n18736) );
  AND U19033 ( .A(n18737), .B(n18738), .Z(n17722) );
  NANDN U19034 ( .A(n18739), .B(n18740), .Z(n18738) );
  NANDN U19035 ( .A(n18741), .B(n18742), .Z(n18740) );
  NANDN U19036 ( .A(n18742), .B(n18741), .Z(n18737) );
  ANDN U19037 ( .B(B[2]), .A(n29), .Z(n17724) );
  XNOR U19038 ( .A(n17631), .B(n18743), .Z(n17725) );
  XNOR U19039 ( .A(n17630), .B(n17628), .Z(n18743) );
  AND U19040 ( .A(n18744), .B(n18745), .Z(n17628) );
  NANDN U19041 ( .A(n18746), .B(n18747), .Z(n18745) );
  OR U19042 ( .A(n18748), .B(n18749), .Z(n18747) );
  NAND U19043 ( .A(n18749), .B(n18748), .Z(n18744) );
  ANDN U19044 ( .B(B[3]), .A(n30), .Z(n17630) );
  XNOR U19045 ( .A(n17638), .B(n18750), .Z(n17631) );
  XNOR U19046 ( .A(n17637), .B(n17635), .Z(n18750) );
  AND U19047 ( .A(n18751), .B(n18752), .Z(n17635) );
  NANDN U19048 ( .A(n18753), .B(n18754), .Z(n18752) );
  NANDN U19049 ( .A(n18755), .B(n18756), .Z(n18754) );
  NANDN U19050 ( .A(n18756), .B(n18755), .Z(n18751) );
  ANDN U19051 ( .B(B[4]), .A(n31), .Z(n17637) );
  XNOR U19052 ( .A(n17645), .B(n18757), .Z(n17638) );
  XNOR U19053 ( .A(n17644), .B(n17642), .Z(n18757) );
  AND U19054 ( .A(n18758), .B(n18759), .Z(n17642) );
  NANDN U19055 ( .A(n18760), .B(n18761), .Z(n18759) );
  OR U19056 ( .A(n18762), .B(n18763), .Z(n18761) );
  NAND U19057 ( .A(n18763), .B(n18762), .Z(n18758) );
  ANDN U19058 ( .B(B[5]), .A(n32), .Z(n17644) );
  XNOR U19059 ( .A(n17652), .B(n18764), .Z(n17645) );
  XNOR U19060 ( .A(n17651), .B(n17649), .Z(n18764) );
  AND U19061 ( .A(n18765), .B(n18766), .Z(n17649) );
  NANDN U19062 ( .A(n18767), .B(n18768), .Z(n18766) );
  NANDN U19063 ( .A(n18769), .B(n18770), .Z(n18768) );
  NANDN U19064 ( .A(n18770), .B(n18769), .Z(n18765) );
  ANDN U19065 ( .B(B[6]), .A(n33), .Z(n17651) );
  XNOR U19066 ( .A(n17659), .B(n18771), .Z(n17652) );
  XNOR U19067 ( .A(n17658), .B(n17656), .Z(n18771) );
  AND U19068 ( .A(n18772), .B(n18773), .Z(n17656) );
  NANDN U19069 ( .A(n18774), .B(n18775), .Z(n18773) );
  OR U19070 ( .A(n18776), .B(n18777), .Z(n18775) );
  NAND U19071 ( .A(n18777), .B(n18776), .Z(n18772) );
  ANDN U19072 ( .B(B[7]), .A(n34), .Z(n17658) );
  XNOR U19073 ( .A(n17666), .B(n18778), .Z(n17659) );
  XNOR U19074 ( .A(n17665), .B(n17663), .Z(n18778) );
  AND U19075 ( .A(n18779), .B(n18780), .Z(n17663) );
  NANDN U19076 ( .A(n18781), .B(n18782), .Z(n18780) );
  NANDN U19077 ( .A(n18783), .B(n18784), .Z(n18782) );
  NANDN U19078 ( .A(n18784), .B(n18783), .Z(n18779) );
  ANDN U19079 ( .B(B[8]), .A(n35), .Z(n17665) );
  XNOR U19080 ( .A(n17673), .B(n18785), .Z(n17666) );
  XNOR U19081 ( .A(n17672), .B(n17670), .Z(n18785) );
  AND U19082 ( .A(n18786), .B(n18787), .Z(n17670) );
  NANDN U19083 ( .A(n18788), .B(n18789), .Z(n18787) );
  OR U19084 ( .A(n18790), .B(n18791), .Z(n18789) );
  NAND U19085 ( .A(n18791), .B(n18790), .Z(n18786) );
  ANDN U19086 ( .B(B[9]), .A(n36), .Z(n17672) );
  XNOR U19087 ( .A(n17680), .B(n18792), .Z(n17673) );
  XNOR U19088 ( .A(n17679), .B(n17677), .Z(n18792) );
  AND U19089 ( .A(n18793), .B(n18794), .Z(n17677) );
  NANDN U19090 ( .A(n18795), .B(n18796), .Z(n18794) );
  NANDN U19091 ( .A(n18797), .B(n18798), .Z(n18796) );
  NANDN U19092 ( .A(n18798), .B(n18797), .Z(n18793) );
  ANDN U19093 ( .B(B[10]), .A(n37), .Z(n17679) );
  XNOR U19094 ( .A(n17687), .B(n18799), .Z(n17680) );
  XNOR U19095 ( .A(n17686), .B(n17684), .Z(n18799) );
  AND U19096 ( .A(n18800), .B(n18801), .Z(n17684) );
  NANDN U19097 ( .A(n18802), .B(n18803), .Z(n18801) );
  OR U19098 ( .A(n18804), .B(n18805), .Z(n18803) );
  NAND U19099 ( .A(n18805), .B(n18804), .Z(n18800) );
  ANDN U19100 ( .B(B[11]), .A(n38), .Z(n17686) );
  XNOR U19101 ( .A(n17694), .B(n18806), .Z(n17687) );
  XNOR U19102 ( .A(n17693), .B(n17691), .Z(n18806) );
  AND U19103 ( .A(n18807), .B(n18808), .Z(n17691) );
  NANDN U19104 ( .A(n18809), .B(n18810), .Z(n18808) );
  NANDN U19105 ( .A(n18811), .B(n18812), .Z(n18810) );
  NANDN U19106 ( .A(n18812), .B(n18811), .Z(n18807) );
  ANDN U19107 ( .B(B[12]), .A(n39), .Z(n17693) );
  XNOR U19108 ( .A(n17701), .B(n18813), .Z(n17694) );
  XNOR U19109 ( .A(n17700), .B(n17698), .Z(n18813) );
  AND U19110 ( .A(n18814), .B(n18815), .Z(n17698) );
  NANDN U19111 ( .A(n18816), .B(n18817), .Z(n18815) );
  OR U19112 ( .A(n18818), .B(n18819), .Z(n18817) );
  NAND U19113 ( .A(n18819), .B(n18818), .Z(n18814) );
  ANDN U19114 ( .B(B[13]), .A(n40), .Z(n17700) );
  XNOR U19115 ( .A(n17708), .B(n18820), .Z(n17701) );
  XNOR U19116 ( .A(n17707), .B(n17705), .Z(n18820) );
  AND U19117 ( .A(n18821), .B(n18822), .Z(n17705) );
  NANDN U19118 ( .A(n18823), .B(n18824), .Z(n18822) );
  NAND U19119 ( .A(n18825), .B(n18826), .Z(n18824) );
  ANDN U19120 ( .B(B[14]), .A(n41), .Z(n17707) );
  XOR U19121 ( .A(n17714), .B(n18827), .Z(n17708) );
  XNOR U19122 ( .A(n17712), .B(n17715), .Z(n18827) );
  NAND U19123 ( .A(A[2]), .B(B[15]), .Z(n17715) );
  NANDN U19124 ( .A(n18828), .B(n18829), .Z(n17712) );
  AND U19125 ( .A(A[0]), .B(B[16]), .Z(n18829) );
  XNOR U19126 ( .A(n17717), .B(n18830), .Z(n17714) );
  NAND U19127 ( .A(A[0]), .B(B[17]), .Z(n18830) );
  NAND U19128 ( .A(B[16]), .B(A[1]), .Z(n17717) );
  NAND U19129 ( .A(n18831), .B(n18832), .Z(n411) );
  NANDN U19130 ( .A(n18833), .B(n18834), .Z(n18832) );
  OR U19131 ( .A(n18835), .B(n18836), .Z(n18834) );
  NAND U19132 ( .A(n18836), .B(n18835), .Z(n18831) );
  XOR U19133 ( .A(n431), .B(n430), .Z(\A1[159] ) );
  XOR U19134 ( .A(n18735), .B(n18837), .Z(n430) );
  XNOR U19135 ( .A(n18734), .B(n18732), .Z(n18837) );
  AND U19136 ( .A(n18838), .B(n18839), .Z(n18732) );
  NANDN U19137 ( .A(n18840), .B(n18841), .Z(n18839) );
  NANDN U19138 ( .A(n18842), .B(n18843), .Z(n18841) );
  NANDN U19139 ( .A(n18843), .B(n18842), .Z(n18838) );
  ANDN U19140 ( .B(B[146]), .A(n29), .Z(n18734) );
  XNOR U19141 ( .A(n18641), .B(n18844), .Z(n18735) );
  XNOR U19142 ( .A(n18640), .B(n18638), .Z(n18844) );
  AND U19143 ( .A(n18845), .B(n18846), .Z(n18638) );
  NANDN U19144 ( .A(n18847), .B(n18848), .Z(n18846) );
  OR U19145 ( .A(n18849), .B(n18850), .Z(n18848) );
  NAND U19146 ( .A(n18850), .B(n18849), .Z(n18845) );
  ANDN U19147 ( .B(B[147]), .A(n30), .Z(n18640) );
  XNOR U19148 ( .A(n18648), .B(n18851), .Z(n18641) );
  XNOR U19149 ( .A(n18647), .B(n18645), .Z(n18851) );
  AND U19150 ( .A(n18852), .B(n18853), .Z(n18645) );
  NANDN U19151 ( .A(n18854), .B(n18855), .Z(n18853) );
  NANDN U19152 ( .A(n18856), .B(n18857), .Z(n18855) );
  NANDN U19153 ( .A(n18857), .B(n18856), .Z(n18852) );
  ANDN U19154 ( .B(B[148]), .A(n31), .Z(n18647) );
  XNOR U19155 ( .A(n18655), .B(n18858), .Z(n18648) );
  XNOR U19156 ( .A(n18654), .B(n18652), .Z(n18858) );
  AND U19157 ( .A(n18859), .B(n18860), .Z(n18652) );
  NANDN U19158 ( .A(n18861), .B(n18862), .Z(n18860) );
  OR U19159 ( .A(n18863), .B(n18864), .Z(n18862) );
  NAND U19160 ( .A(n18864), .B(n18863), .Z(n18859) );
  ANDN U19161 ( .B(B[149]), .A(n32), .Z(n18654) );
  XNOR U19162 ( .A(n18662), .B(n18865), .Z(n18655) );
  XNOR U19163 ( .A(n18661), .B(n18659), .Z(n18865) );
  AND U19164 ( .A(n18866), .B(n18867), .Z(n18659) );
  NANDN U19165 ( .A(n18868), .B(n18869), .Z(n18867) );
  NANDN U19166 ( .A(n18870), .B(n18871), .Z(n18869) );
  NANDN U19167 ( .A(n18871), .B(n18870), .Z(n18866) );
  ANDN U19168 ( .B(B[150]), .A(n33), .Z(n18661) );
  XNOR U19169 ( .A(n18669), .B(n18872), .Z(n18662) );
  XNOR U19170 ( .A(n18668), .B(n18666), .Z(n18872) );
  AND U19171 ( .A(n18873), .B(n18874), .Z(n18666) );
  NANDN U19172 ( .A(n18875), .B(n18876), .Z(n18874) );
  OR U19173 ( .A(n18877), .B(n18878), .Z(n18876) );
  NAND U19174 ( .A(n18878), .B(n18877), .Z(n18873) );
  ANDN U19175 ( .B(B[151]), .A(n34), .Z(n18668) );
  XNOR U19176 ( .A(n18676), .B(n18879), .Z(n18669) );
  XNOR U19177 ( .A(n18675), .B(n18673), .Z(n18879) );
  AND U19178 ( .A(n18880), .B(n18881), .Z(n18673) );
  NANDN U19179 ( .A(n18882), .B(n18883), .Z(n18881) );
  NANDN U19180 ( .A(n18884), .B(n18885), .Z(n18883) );
  NANDN U19181 ( .A(n18885), .B(n18884), .Z(n18880) );
  ANDN U19182 ( .B(B[152]), .A(n35), .Z(n18675) );
  XNOR U19183 ( .A(n18683), .B(n18886), .Z(n18676) );
  XNOR U19184 ( .A(n18682), .B(n18680), .Z(n18886) );
  AND U19185 ( .A(n18887), .B(n18888), .Z(n18680) );
  NANDN U19186 ( .A(n18889), .B(n18890), .Z(n18888) );
  OR U19187 ( .A(n18891), .B(n18892), .Z(n18890) );
  NAND U19188 ( .A(n18892), .B(n18891), .Z(n18887) );
  ANDN U19189 ( .B(B[153]), .A(n36), .Z(n18682) );
  XNOR U19190 ( .A(n18690), .B(n18893), .Z(n18683) );
  XNOR U19191 ( .A(n18689), .B(n18687), .Z(n18893) );
  AND U19192 ( .A(n18894), .B(n18895), .Z(n18687) );
  NANDN U19193 ( .A(n18896), .B(n18897), .Z(n18895) );
  NANDN U19194 ( .A(n18898), .B(n18899), .Z(n18897) );
  NANDN U19195 ( .A(n18899), .B(n18898), .Z(n18894) );
  ANDN U19196 ( .B(B[154]), .A(n37), .Z(n18689) );
  XNOR U19197 ( .A(n18697), .B(n18900), .Z(n18690) );
  XNOR U19198 ( .A(n18696), .B(n18694), .Z(n18900) );
  AND U19199 ( .A(n18901), .B(n18902), .Z(n18694) );
  NANDN U19200 ( .A(n18903), .B(n18904), .Z(n18902) );
  OR U19201 ( .A(n18905), .B(n18906), .Z(n18904) );
  NAND U19202 ( .A(n18906), .B(n18905), .Z(n18901) );
  ANDN U19203 ( .B(B[155]), .A(n38), .Z(n18696) );
  XNOR U19204 ( .A(n18704), .B(n18907), .Z(n18697) );
  XNOR U19205 ( .A(n18703), .B(n18701), .Z(n18907) );
  AND U19206 ( .A(n18908), .B(n18909), .Z(n18701) );
  NANDN U19207 ( .A(n18910), .B(n18911), .Z(n18909) );
  NANDN U19208 ( .A(n18912), .B(n18913), .Z(n18911) );
  NANDN U19209 ( .A(n18913), .B(n18912), .Z(n18908) );
  ANDN U19210 ( .B(B[156]), .A(n39), .Z(n18703) );
  XNOR U19211 ( .A(n18711), .B(n18914), .Z(n18704) );
  XNOR U19212 ( .A(n18710), .B(n18708), .Z(n18914) );
  AND U19213 ( .A(n18915), .B(n18916), .Z(n18708) );
  NANDN U19214 ( .A(n18917), .B(n18918), .Z(n18916) );
  OR U19215 ( .A(n18919), .B(n18920), .Z(n18918) );
  NAND U19216 ( .A(n18920), .B(n18919), .Z(n18915) );
  ANDN U19217 ( .B(B[157]), .A(n40), .Z(n18710) );
  XNOR U19218 ( .A(n18718), .B(n18921), .Z(n18711) );
  XNOR U19219 ( .A(n18717), .B(n18715), .Z(n18921) );
  AND U19220 ( .A(n18922), .B(n18923), .Z(n18715) );
  NANDN U19221 ( .A(n18924), .B(n18925), .Z(n18923) );
  NAND U19222 ( .A(n18926), .B(n18927), .Z(n18925) );
  ANDN U19223 ( .B(B[158]), .A(n41), .Z(n18717) );
  XOR U19224 ( .A(n18724), .B(n18928), .Z(n18718) );
  XNOR U19225 ( .A(n18722), .B(n18725), .Z(n18928) );
  NAND U19226 ( .A(A[2]), .B(B[159]), .Z(n18725) );
  NANDN U19227 ( .A(n18929), .B(n18930), .Z(n18722) );
  AND U19228 ( .A(A[0]), .B(B[160]), .Z(n18930) );
  XNOR U19229 ( .A(n18727), .B(n18931), .Z(n18724) );
  NAND U19230 ( .A(A[0]), .B(B[161]), .Z(n18931) );
  NAND U19231 ( .A(B[160]), .B(A[1]), .Z(n18727) );
  NAND U19232 ( .A(n18932), .B(n18933), .Z(n431) );
  NANDN U19233 ( .A(n18934), .B(n18935), .Z(n18933) );
  OR U19234 ( .A(n18936), .B(n18937), .Z(n18935) );
  NAND U19235 ( .A(n18937), .B(n18936), .Z(n18932) );
  XOR U19236 ( .A(n435), .B(n434), .Z(\A1[158] ) );
  XOR U19237 ( .A(n18937), .B(n18938), .Z(n434) );
  XNOR U19238 ( .A(n18936), .B(n18934), .Z(n18938) );
  AND U19239 ( .A(n18939), .B(n18940), .Z(n18934) );
  NANDN U19240 ( .A(n18941), .B(n18942), .Z(n18940) );
  NANDN U19241 ( .A(n18943), .B(n18944), .Z(n18942) );
  NANDN U19242 ( .A(n18944), .B(n18943), .Z(n18939) );
  ANDN U19243 ( .B(B[145]), .A(n29), .Z(n18936) );
  XNOR U19244 ( .A(n18843), .B(n18945), .Z(n18937) );
  XNOR U19245 ( .A(n18842), .B(n18840), .Z(n18945) );
  AND U19246 ( .A(n18946), .B(n18947), .Z(n18840) );
  NANDN U19247 ( .A(n18948), .B(n18949), .Z(n18947) );
  OR U19248 ( .A(n18950), .B(n18951), .Z(n18949) );
  NAND U19249 ( .A(n18951), .B(n18950), .Z(n18946) );
  ANDN U19250 ( .B(B[146]), .A(n30), .Z(n18842) );
  XNOR U19251 ( .A(n18850), .B(n18952), .Z(n18843) );
  XNOR U19252 ( .A(n18849), .B(n18847), .Z(n18952) );
  AND U19253 ( .A(n18953), .B(n18954), .Z(n18847) );
  NANDN U19254 ( .A(n18955), .B(n18956), .Z(n18954) );
  NANDN U19255 ( .A(n18957), .B(n18958), .Z(n18956) );
  NANDN U19256 ( .A(n18958), .B(n18957), .Z(n18953) );
  ANDN U19257 ( .B(B[147]), .A(n31), .Z(n18849) );
  XNOR U19258 ( .A(n18857), .B(n18959), .Z(n18850) );
  XNOR U19259 ( .A(n18856), .B(n18854), .Z(n18959) );
  AND U19260 ( .A(n18960), .B(n18961), .Z(n18854) );
  NANDN U19261 ( .A(n18962), .B(n18963), .Z(n18961) );
  OR U19262 ( .A(n18964), .B(n18965), .Z(n18963) );
  NAND U19263 ( .A(n18965), .B(n18964), .Z(n18960) );
  ANDN U19264 ( .B(B[148]), .A(n32), .Z(n18856) );
  XNOR U19265 ( .A(n18864), .B(n18966), .Z(n18857) );
  XNOR U19266 ( .A(n18863), .B(n18861), .Z(n18966) );
  AND U19267 ( .A(n18967), .B(n18968), .Z(n18861) );
  NANDN U19268 ( .A(n18969), .B(n18970), .Z(n18968) );
  NANDN U19269 ( .A(n18971), .B(n18972), .Z(n18970) );
  NANDN U19270 ( .A(n18972), .B(n18971), .Z(n18967) );
  ANDN U19271 ( .B(B[149]), .A(n33), .Z(n18863) );
  XNOR U19272 ( .A(n18871), .B(n18973), .Z(n18864) );
  XNOR U19273 ( .A(n18870), .B(n18868), .Z(n18973) );
  AND U19274 ( .A(n18974), .B(n18975), .Z(n18868) );
  NANDN U19275 ( .A(n18976), .B(n18977), .Z(n18975) );
  OR U19276 ( .A(n18978), .B(n18979), .Z(n18977) );
  NAND U19277 ( .A(n18979), .B(n18978), .Z(n18974) );
  ANDN U19278 ( .B(B[150]), .A(n34), .Z(n18870) );
  XNOR U19279 ( .A(n18878), .B(n18980), .Z(n18871) );
  XNOR U19280 ( .A(n18877), .B(n18875), .Z(n18980) );
  AND U19281 ( .A(n18981), .B(n18982), .Z(n18875) );
  NANDN U19282 ( .A(n18983), .B(n18984), .Z(n18982) );
  NANDN U19283 ( .A(n18985), .B(n18986), .Z(n18984) );
  NANDN U19284 ( .A(n18986), .B(n18985), .Z(n18981) );
  ANDN U19285 ( .B(B[151]), .A(n35), .Z(n18877) );
  XNOR U19286 ( .A(n18885), .B(n18987), .Z(n18878) );
  XNOR U19287 ( .A(n18884), .B(n18882), .Z(n18987) );
  AND U19288 ( .A(n18988), .B(n18989), .Z(n18882) );
  NANDN U19289 ( .A(n18990), .B(n18991), .Z(n18989) );
  OR U19290 ( .A(n18992), .B(n18993), .Z(n18991) );
  NAND U19291 ( .A(n18993), .B(n18992), .Z(n18988) );
  ANDN U19292 ( .B(B[152]), .A(n36), .Z(n18884) );
  XNOR U19293 ( .A(n18892), .B(n18994), .Z(n18885) );
  XNOR U19294 ( .A(n18891), .B(n18889), .Z(n18994) );
  AND U19295 ( .A(n18995), .B(n18996), .Z(n18889) );
  NANDN U19296 ( .A(n18997), .B(n18998), .Z(n18996) );
  NANDN U19297 ( .A(n18999), .B(n19000), .Z(n18998) );
  NANDN U19298 ( .A(n19000), .B(n18999), .Z(n18995) );
  ANDN U19299 ( .B(B[153]), .A(n37), .Z(n18891) );
  XNOR U19300 ( .A(n18899), .B(n19001), .Z(n18892) );
  XNOR U19301 ( .A(n18898), .B(n18896), .Z(n19001) );
  AND U19302 ( .A(n19002), .B(n19003), .Z(n18896) );
  NANDN U19303 ( .A(n19004), .B(n19005), .Z(n19003) );
  OR U19304 ( .A(n19006), .B(n19007), .Z(n19005) );
  NAND U19305 ( .A(n19007), .B(n19006), .Z(n19002) );
  ANDN U19306 ( .B(B[154]), .A(n38), .Z(n18898) );
  XNOR U19307 ( .A(n18906), .B(n19008), .Z(n18899) );
  XNOR U19308 ( .A(n18905), .B(n18903), .Z(n19008) );
  AND U19309 ( .A(n19009), .B(n19010), .Z(n18903) );
  NANDN U19310 ( .A(n19011), .B(n19012), .Z(n19010) );
  NANDN U19311 ( .A(n19013), .B(n19014), .Z(n19012) );
  NANDN U19312 ( .A(n19014), .B(n19013), .Z(n19009) );
  ANDN U19313 ( .B(B[155]), .A(n39), .Z(n18905) );
  XNOR U19314 ( .A(n18913), .B(n19015), .Z(n18906) );
  XNOR U19315 ( .A(n18912), .B(n18910), .Z(n19015) );
  AND U19316 ( .A(n19016), .B(n19017), .Z(n18910) );
  NANDN U19317 ( .A(n19018), .B(n19019), .Z(n19017) );
  OR U19318 ( .A(n19020), .B(n19021), .Z(n19019) );
  NAND U19319 ( .A(n19021), .B(n19020), .Z(n19016) );
  ANDN U19320 ( .B(B[156]), .A(n40), .Z(n18912) );
  XNOR U19321 ( .A(n18920), .B(n19022), .Z(n18913) );
  XNOR U19322 ( .A(n18919), .B(n18917), .Z(n19022) );
  AND U19323 ( .A(n19023), .B(n19024), .Z(n18917) );
  NANDN U19324 ( .A(n19025), .B(n19026), .Z(n19024) );
  NAND U19325 ( .A(n19027), .B(n19028), .Z(n19026) );
  ANDN U19326 ( .B(B[157]), .A(n41), .Z(n18919) );
  XOR U19327 ( .A(n18926), .B(n19029), .Z(n18920) );
  XNOR U19328 ( .A(n18924), .B(n18927), .Z(n19029) );
  NAND U19329 ( .A(A[2]), .B(B[158]), .Z(n18927) );
  NANDN U19330 ( .A(n19030), .B(n19031), .Z(n18924) );
  AND U19331 ( .A(A[0]), .B(B[159]), .Z(n19031) );
  XNOR U19332 ( .A(n18929), .B(n19032), .Z(n18926) );
  NAND U19333 ( .A(A[0]), .B(B[160]), .Z(n19032) );
  NAND U19334 ( .A(B[159]), .B(A[1]), .Z(n18929) );
  NAND U19335 ( .A(n19033), .B(n19034), .Z(n435) );
  NANDN U19336 ( .A(n19035), .B(n19036), .Z(n19034) );
  OR U19337 ( .A(n19037), .B(n19038), .Z(n19036) );
  NAND U19338 ( .A(n19038), .B(n19037), .Z(n19033) );
  XOR U19339 ( .A(n437), .B(n436), .Z(\A1[157] ) );
  XOR U19340 ( .A(n19038), .B(n19039), .Z(n436) );
  XNOR U19341 ( .A(n19037), .B(n19035), .Z(n19039) );
  AND U19342 ( .A(n19040), .B(n19041), .Z(n19035) );
  NANDN U19343 ( .A(n19042), .B(n19043), .Z(n19041) );
  NANDN U19344 ( .A(n19044), .B(n19045), .Z(n19043) );
  NANDN U19345 ( .A(n19045), .B(n19044), .Z(n19040) );
  ANDN U19346 ( .B(B[144]), .A(n29), .Z(n19037) );
  XNOR U19347 ( .A(n18944), .B(n19046), .Z(n19038) );
  XNOR U19348 ( .A(n18943), .B(n18941), .Z(n19046) );
  AND U19349 ( .A(n19047), .B(n19048), .Z(n18941) );
  NANDN U19350 ( .A(n19049), .B(n19050), .Z(n19048) );
  OR U19351 ( .A(n19051), .B(n19052), .Z(n19050) );
  NAND U19352 ( .A(n19052), .B(n19051), .Z(n19047) );
  ANDN U19353 ( .B(B[145]), .A(n30), .Z(n18943) );
  XNOR U19354 ( .A(n18951), .B(n19053), .Z(n18944) );
  XNOR U19355 ( .A(n18950), .B(n18948), .Z(n19053) );
  AND U19356 ( .A(n19054), .B(n19055), .Z(n18948) );
  NANDN U19357 ( .A(n19056), .B(n19057), .Z(n19055) );
  NANDN U19358 ( .A(n19058), .B(n19059), .Z(n19057) );
  NANDN U19359 ( .A(n19059), .B(n19058), .Z(n19054) );
  ANDN U19360 ( .B(B[146]), .A(n31), .Z(n18950) );
  XNOR U19361 ( .A(n18958), .B(n19060), .Z(n18951) );
  XNOR U19362 ( .A(n18957), .B(n18955), .Z(n19060) );
  AND U19363 ( .A(n19061), .B(n19062), .Z(n18955) );
  NANDN U19364 ( .A(n19063), .B(n19064), .Z(n19062) );
  OR U19365 ( .A(n19065), .B(n19066), .Z(n19064) );
  NAND U19366 ( .A(n19066), .B(n19065), .Z(n19061) );
  ANDN U19367 ( .B(B[147]), .A(n32), .Z(n18957) );
  XNOR U19368 ( .A(n18965), .B(n19067), .Z(n18958) );
  XNOR U19369 ( .A(n18964), .B(n18962), .Z(n19067) );
  AND U19370 ( .A(n19068), .B(n19069), .Z(n18962) );
  NANDN U19371 ( .A(n19070), .B(n19071), .Z(n19069) );
  NANDN U19372 ( .A(n19072), .B(n19073), .Z(n19071) );
  NANDN U19373 ( .A(n19073), .B(n19072), .Z(n19068) );
  ANDN U19374 ( .B(B[148]), .A(n33), .Z(n18964) );
  XNOR U19375 ( .A(n18972), .B(n19074), .Z(n18965) );
  XNOR U19376 ( .A(n18971), .B(n18969), .Z(n19074) );
  AND U19377 ( .A(n19075), .B(n19076), .Z(n18969) );
  NANDN U19378 ( .A(n19077), .B(n19078), .Z(n19076) );
  OR U19379 ( .A(n19079), .B(n19080), .Z(n19078) );
  NAND U19380 ( .A(n19080), .B(n19079), .Z(n19075) );
  ANDN U19381 ( .B(B[149]), .A(n34), .Z(n18971) );
  XNOR U19382 ( .A(n18979), .B(n19081), .Z(n18972) );
  XNOR U19383 ( .A(n18978), .B(n18976), .Z(n19081) );
  AND U19384 ( .A(n19082), .B(n19083), .Z(n18976) );
  NANDN U19385 ( .A(n19084), .B(n19085), .Z(n19083) );
  NANDN U19386 ( .A(n19086), .B(n19087), .Z(n19085) );
  NANDN U19387 ( .A(n19087), .B(n19086), .Z(n19082) );
  ANDN U19388 ( .B(B[150]), .A(n35), .Z(n18978) );
  XNOR U19389 ( .A(n18986), .B(n19088), .Z(n18979) );
  XNOR U19390 ( .A(n18985), .B(n18983), .Z(n19088) );
  AND U19391 ( .A(n19089), .B(n19090), .Z(n18983) );
  NANDN U19392 ( .A(n19091), .B(n19092), .Z(n19090) );
  OR U19393 ( .A(n19093), .B(n19094), .Z(n19092) );
  NAND U19394 ( .A(n19094), .B(n19093), .Z(n19089) );
  ANDN U19395 ( .B(B[151]), .A(n36), .Z(n18985) );
  XNOR U19396 ( .A(n18993), .B(n19095), .Z(n18986) );
  XNOR U19397 ( .A(n18992), .B(n18990), .Z(n19095) );
  AND U19398 ( .A(n19096), .B(n19097), .Z(n18990) );
  NANDN U19399 ( .A(n19098), .B(n19099), .Z(n19097) );
  NANDN U19400 ( .A(n19100), .B(n19101), .Z(n19099) );
  NANDN U19401 ( .A(n19101), .B(n19100), .Z(n19096) );
  ANDN U19402 ( .B(B[152]), .A(n37), .Z(n18992) );
  XNOR U19403 ( .A(n19000), .B(n19102), .Z(n18993) );
  XNOR U19404 ( .A(n18999), .B(n18997), .Z(n19102) );
  AND U19405 ( .A(n19103), .B(n19104), .Z(n18997) );
  NANDN U19406 ( .A(n19105), .B(n19106), .Z(n19104) );
  OR U19407 ( .A(n19107), .B(n19108), .Z(n19106) );
  NAND U19408 ( .A(n19108), .B(n19107), .Z(n19103) );
  ANDN U19409 ( .B(B[153]), .A(n38), .Z(n18999) );
  XNOR U19410 ( .A(n19007), .B(n19109), .Z(n19000) );
  XNOR U19411 ( .A(n19006), .B(n19004), .Z(n19109) );
  AND U19412 ( .A(n19110), .B(n19111), .Z(n19004) );
  NANDN U19413 ( .A(n19112), .B(n19113), .Z(n19111) );
  NANDN U19414 ( .A(n19114), .B(n19115), .Z(n19113) );
  NANDN U19415 ( .A(n19115), .B(n19114), .Z(n19110) );
  ANDN U19416 ( .B(B[154]), .A(n39), .Z(n19006) );
  XNOR U19417 ( .A(n19014), .B(n19116), .Z(n19007) );
  XNOR U19418 ( .A(n19013), .B(n19011), .Z(n19116) );
  AND U19419 ( .A(n19117), .B(n19118), .Z(n19011) );
  NANDN U19420 ( .A(n19119), .B(n19120), .Z(n19118) );
  OR U19421 ( .A(n19121), .B(n19122), .Z(n19120) );
  NAND U19422 ( .A(n19122), .B(n19121), .Z(n19117) );
  ANDN U19423 ( .B(B[155]), .A(n40), .Z(n19013) );
  XNOR U19424 ( .A(n19021), .B(n19123), .Z(n19014) );
  XNOR U19425 ( .A(n19020), .B(n19018), .Z(n19123) );
  AND U19426 ( .A(n19124), .B(n19125), .Z(n19018) );
  NANDN U19427 ( .A(n19126), .B(n19127), .Z(n19125) );
  NAND U19428 ( .A(n19128), .B(n19129), .Z(n19127) );
  ANDN U19429 ( .B(B[156]), .A(n41), .Z(n19020) );
  XOR U19430 ( .A(n19027), .B(n19130), .Z(n19021) );
  XNOR U19431 ( .A(n19025), .B(n19028), .Z(n19130) );
  NAND U19432 ( .A(A[2]), .B(B[157]), .Z(n19028) );
  NANDN U19433 ( .A(n19131), .B(n19132), .Z(n19025) );
  AND U19434 ( .A(A[0]), .B(B[158]), .Z(n19132) );
  XNOR U19435 ( .A(n19030), .B(n19133), .Z(n19027) );
  NAND U19436 ( .A(A[0]), .B(B[159]), .Z(n19133) );
  NAND U19437 ( .A(B[158]), .B(A[1]), .Z(n19030) );
  NAND U19438 ( .A(n19134), .B(n19135), .Z(n437) );
  NANDN U19439 ( .A(n19136), .B(n19137), .Z(n19135) );
  OR U19440 ( .A(n19138), .B(n19139), .Z(n19137) );
  NAND U19441 ( .A(n19139), .B(n19138), .Z(n19134) );
  XOR U19442 ( .A(n439), .B(n438), .Z(\A1[156] ) );
  XOR U19443 ( .A(n19139), .B(n19140), .Z(n438) );
  XNOR U19444 ( .A(n19138), .B(n19136), .Z(n19140) );
  AND U19445 ( .A(n19141), .B(n19142), .Z(n19136) );
  NANDN U19446 ( .A(n19143), .B(n19144), .Z(n19142) );
  NANDN U19447 ( .A(n19145), .B(n19146), .Z(n19144) );
  NANDN U19448 ( .A(n19146), .B(n19145), .Z(n19141) );
  ANDN U19449 ( .B(B[143]), .A(n29), .Z(n19138) );
  XNOR U19450 ( .A(n19045), .B(n19147), .Z(n19139) );
  XNOR U19451 ( .A(n19044), .B(n19042), .Z(n19147) );
  AND U19452 ( .A(n19148), .B(n19149), .Z(n19042) );
  NANDN U19453 ( .A(n19150), .B(n19151), .Z(n19149) );
  OR U19454 ( .A(n19152), .B(n19153), .Z(n19151) );
  NAND U19455 ( .A(n19153), .B(n19152), .Z(n19148) );
  ANDN U19456 ( .B(B[144]), .A(n30), .Z(n19044) );
  XNOR U19457 ( .A(n19052), .B(n19154), .Z(n19045) );
  XNOR U19458 ( .A(n19051), .B(n19049), .Z(n19154) );
  AND U19459 ( .A(n19155), .B(n19156), .Z(n19049) );
  NANDN U19460 ( .A(n19157), .B(n19158), .Z(n19156) );
  NANDN U19461 ( .A(n19159), .B(n19160), .Z(n19158) );
  NANDN U19462 ( .A(n19160), .B(n19159), .Z(n19155) );
  ANDN U19463 ( .B(B[145]), .A(n31), .Z(n19051) );
  XNOR U19464 ( .A(n19059), .B(n19161), .Z(n19052) );
  XNOR U19465 ( .A(n19058), .B(n19056), .Z(n19161) );
  AND U19466 ( .A(n19162), .B(n19163), .Z(n19056) );
  NANDN U19467 ( .A(n19164), .B(n19165), .Z(n19163) );
  OR U19468 ( .A(n19166), .B(n19167), .Z(n19165) );
  NAND U19469 ( .A(n19167), .B(n19166), .Z(n19162) );
  ANDN U19470 ( .B(B[146]), .A(n32), .Z(n19058) );
  XNOR U19471 ( .A(n19066), .B(n19168), .Z(n19059) );
  XNOR U19472 ( .A(n19065), .B(n19063), .Z(n19168) );
  AND U19473 ( .A(n19169), .B(n19170), .Z(n19063) );
  NANDN U19474 ( .A(n19171), .B(n19172), .Z(n19170) );
  NANDN U19475 ( .A(n19173), .B(n19174), .Z(n19172) );
  NANDN U19476 ( .A(n19174), .B(n19173), .Z(n19169) );
  ANDN U19477 ( .B(B[147]), .A(n33), .Z(n19065) );
  XNOR U19478 ( .A(n19073), .B(n19175), .Z(n19066) );
  XNOR U19479 ( .A(n19072), .B(n19070), .Z(n19175) );
  AND U19480 ( .A(n19176), .B(n19177), .Z(n19070) );
  NANDN U19481 ( .A(n19178), .B(n19179), .Z(n19177) );
  OR U19482 ( .A(n19180), .B(n19181), .Z(n19179) );
  NAND U19483 ( .A(n19181), .B(n19180), .Z(n19176) );
  ANDN U19484 ( .B(B[148]), .A(n34), .Z(n19072) );
  XNOR U19485 ( .A(n19080), .B(n19182), .Z(n19073) );
  XNOR U19486 ( .A(n19079), .B(n19077), .Z(n19182) );
  AND U19487 ( .A(n19183), .B(n19184), .Z(n19077) );
  NANDN U19488 ( .A(n19185), .B(n19186), .Z(n19184) );
  NANDN U19489 ( .A(n19187), .B(n19188), .Z(n19186) );
  NANDN U19490 ( .A(n19188), .B(n19187), .Z(n19183) );
  ANDN U19491 ( .B(B[149]), .A(n35), .Z(n19079) );
  XNOR U19492 ( .A(n19087), .B(n19189), .Z(n19080) );
  XNOR U19493 ( .A(n19086), .B(n19084), .Z(n19189) );
  AND U19494 ( .A(n19190), .B(n19191), .Z(n19084) );
  NANDN U19495 ( .A(n19192), .B(n19193), .Z(n19191) );
  OR U19496 ( .A(n19194), .B(n19195), .Z(n19193) );
  NAND U19497 ( .A(n19195), .B(n19194), .Z(n19190) );
  ANDN U19498 ( .B(B[150]), .A(n36), .Z(n19086) );
  XNOR U19499 ( .A(n19094), .B(n19196), .Z(n19087) );
  XNOR U19500 ( .A(n19093), .B(n19091), .Z(n19196) );
  AND U19501 ( .A(n19197), .B(n19198), .Z(n19091) );
  NANDN U19502 ( .A(n19199), .B(n19200), .Z(n19198) );
  NANDN U19503 ( .A(n19201), .B(n19202), .Z(n19200) );
  NANDN U19504 ( .A(n19202), .B(n19201), .Z(n19197) );
  ANDN U19505 ( .B(B[151]), .A(n37), .Z(n19093) );
  XNOR U19506 ( .A(n19101), .B(n19203), .Z(n19094) );
  XNOR U19507 ( .A(n19100), .B(n19098), .Z(n19203) );
  AND U19508 ( .A(n19204), .B(n19205), .Z(n19098) );
  NANDN U19509 ( .A(n19206), .B(n19207), .Z(n19205) );
  OR U19510 ( .A(n19208), .B(n19209), .Z(n19207) );
  NAND U19511 ( .A(n19209), .B(n19208), .Z(n19204) );
  ANDN U19512 ( .B(B[152]), .A(n38), .Z(n19100) );
  XNOR U19513 ( .A(n19108), .B(n19210), .Z(n19101) );
  XNOR U19514 ( .A(n19107), .B(n19105), .Z(n19210) );
  AND U19515 ( .A(n19211), .B(n19212), .Z(n19105) );
  NANDN U19516 ( .A(n19213), .B(n19214), .Z(n19212) );
  NANDN U19517 ( .A(n19215), .B(n19216), .Z(n19214) );
  NANDN U19518 ( .A(n19216), .B(n19215), .Z(n19211) );
  ANDN U19519 ( .B(B[153]), .A(n39), .Z(n19107) );
  XNOR U19520 ( .A(n19115), .B(n19217), .Z(n19108) );
  XNOR U19521 ( .A(n19114), .B(n19112), .Z(n19217) );
  AND U19522 ( .A(n19218), .B(n19219), .Z(n19112) );
  NANDN U19523 ( .A(n19220), .B(n19221), .Z(n19219) );
  OR U19524 ( .A(n19222), .B(n19223), .Z(n19221) );
  NAND U19525 ( .A(n19223), .B(n19222), .Z(n19218) );
  ANDN U19526 ( .B(B[154]), .A(n40), .Z(n19114) );
  XNOR U19527 ( .A(n19122), .B(n19224), .Z(n19115) );
  XNOR U19528 ( .A(n19121), .B(n19119), .Z(n19224) );
  AND U19529 ( .A(n19225), .B(n19226), .Z(n19119) );
  NANDN U19530 ( .A(n19227), .B(n19228), .Z(n19226) );
  NAND U19531 ( .A(n19229), .B(n19230), .Z(n19228) );
  ANDN U19532 ( .B(B[155]), .A(n41), .Z(n19121) );
  XOR U19533 ( .A(n19128), .B(n19231), .Z(n19122) );
  XNOR U19534 ( .A(n19126), .B(n19129), .Z(n19231) );
  NAND U19535 ( .A(A[2]), .B(B[156]), .Z(n19129) );
  NANDN U19536 ( .A(n19232), .B(n19233), .Z(n19126) );
  AND U19537 ( .A(A[0]), .B(B[157]), .Z(n19233) );
  XNOR U19538 ( .A(n19131), .B(n19234), .Z(n19128) );
  NAND U19539 ( .A(A[0]), .B(B[158]), .Z(n19234) );
  NAND U19540 ( .A(B[157]), .B(A[1]), .Z(n19131) );
  NAND U19541 ( .A(n19235), .B(n19236), .Z(n439) );
  NANDN U19542 ( .A(n19237), .B(n19238), .Z(n19236) );
  OR U19543 ( .A(n19239), .B(n19240), .Z(n19238) );
  NAND U19544 ( .A(n19240), .B(n19239), .Z(n19235) );
  XOR U19545 ( .A(n441), .B(n440), .Z(\A1[155] ) );
  XOR U19546 ( .A(n19240), .B(n19241), .Z(n440) );
  XNOR U19547 ( .A(n19239), .B(n19237), .Z(n19241) );
  AND U19548 ( .A(n19242), .B(n19243), .Z(n19237) );
  NANDN U19549 ( .A(n19244), .B(n19245), .Z(n19243) );
  NANDN U19550 ( .A(n19246), .B(n19247), .Z(n19245) );
  NANDN U19551 ( .A(n19247), .B(n19246), .Z(n19242) );
  ANDN U19552 ( .B(B[142]), .A(n29), .Z(n19239) );
  XNOR U19553 ( .A(n19146), .B(n19248), .Z(n19240) );
  XNOR U19554 ( .A(n19145), .B(n19143), .Z(n19248) );
  AND U19555 ( .A(n19249), .B(n19250), .Z(n19143) );
  NANDN U19556 ( .A(n19251), .B(n19252), .Z(n19250) );
  OR U19557 ( .A(n19253), .B(n19254), .Z(n19252) );
  NAND U19558 ( .A(n19254), .B(n19253), .Z(n19249) );
  ANDN U19559 ( .B(B[143]), .A(n30), .Z(n19145) );
  XNOR U19560 ( .A(n19153), .B(n19255), .Z(n19146) );
  XNOR U19561 ( .A(n19152), .B(n19150), .Z(n19255) );
  AND U19562 ( .A(n19256), .B(n19257), .Z(n19150) );
  NANDN U19563 ( .A(n19258), .B(n19259), .Z(n19257) );
  NANDN U19564 ( .A(n19260), .B(n19261), .Z(n19259) );
  NANDN U19565 ( .A(n19261), .B(n19260), .Z(n19256) );
  ANDN U19566 ( .B(B[144]), .A(n31), .Z(n19152) );
  XNOR U19567 ( .A(n19160), .B(n19262), .Z(n19153) );
  XNOR U19568 ( .A(n19159), .B(n19157), .Z(n19262) );
  AND U19569 ( .A(n19263), .B(n19264), .Z(n19157) );
  NANDN U19570 ( .A(n19265), .B(n19266), .Z(n19264) );
  OR U19571 ( .A(n19267), .B(n19268), .Z(n19266) );
  NAND U19572 ( .A(n19268), .B(n19267), .Z(n19263) );
  ANDN U19573 ( .B(B[145]), .A(n32), .Z(n19159) );
  XNOR U19574 ( .A(n19167), .B(n19269), .Z(n19160) );
  XNOR U19575 ( .A(n19166), .B(n19164), .Z(n19269) );
  AND U19576 ( .A(n19270), .B(n19271), .Z(n19164) );
  NANDN U19577 ( .A(n19272), .B(n19273), .Z(n19271) );
  NANDN U19578 ( .A(n19274), .B(n19275), .Z(n19273) );
  NANDN U19579 ( .A(n19275), .B(n19274), .Z(n19270) );
  ANDN U19580 ( .B(B[146]), .A(n33), .Z(n19166) );
  XNOR U19581 ( .A(n19174), .B(n19276), .Z(n19167) );
  XNOR U19582 ( .A(n19173), .B(n19171), .Z(n19276) );
  AND U19583 ( .A(n19277), .B(n19278), .Z(n19171) );
  NANDN U19584 ( .A(n19279), .B(n19280), .Z(n19278) );
  OR U19585 ( .A(n19281), .B(n19282), .Z(n19280) );
  NAND U19586 ( .A(n19282), .B(n19281), .Z(n19277) );
  ANDN U19587 ( .B(B[147]), .A(n34), .Z(n19173) );
  XNOR U19588 ( .A(n19181), .B(n19283), .Z(n19174) );
  XNOR U19589 ( .A(n19180), .B(n19178), .Z(n19283) );
  AND U19590 ( .A(n19284), .B(n19285), .Z(n19178) );
  NANDN U19591 ( .A(n19286), .B(n19287), .Z(n19285) );
  NANDN U19592 ( .A(n19288), .B(n19289), .Z(n19287) );
  NANDN U19593 ( .A(n19289), .B(n19288), .Z(n19284) );
  ANDN U19594 ( .B(B[148]), .A(n35), .Z(n19180) );
  XNOR U19595 ( .A(n19188), .B(n19290), .Z(n19181) );
  XNOR U19596 ( .A(n19187), .B(n19185), .Z(n19290) );
  AND U19597 ( .A(n19291), .B(n19292), .Z(n19185) );
  NANDN U19598 ( .A(n19293), .B(n19294), .Z(n19292) );
  OR U19599 ( .A(n19295), .B(n19296), .Z(n19294) );
  NAND U19600 ( .A(n19296), .B(n19295), .Z(n19291) );
  ANDN U19601 ( .B(B[149]), .A(n36), .Z(n19187) );
  XNOR U19602 ( .A(n19195), .B(n19297), .Z(n19188) );
  XNOR U19603 ( .A(n19194), .B(n19192), .Z(n19297) );
  AND U19604 ( .A(n19298), .B(n19299), .Z(n19192) );
  NANDN U19605 ( .A(n19300), .B(n19301), .Z(n19299) );
  NANDN U19606 ( .A(n19302), .B(n19303), .Z(n19301) );
  NANDN U19607 ( .A(n19303), .B(n19302), .Z(n19298) );
  ANDN U19608 ( .B(B[150]), .A(n37), .Z(n19194) );
  XNOR U19609 ( .A(n19202), .B(n19304), .Z(n19195) );
  XNOR U19610 ( .A(n19201), .B(n19199), .Z(n19304) );
  AND U19611 ( .A(n19305), .B(n19306), .Z(n19199) );
  NANDN U19612 ( .A(n19307), .B(n19308), .Z(n19306) );
  OR U19613 ( .A(n19309), .B(n19310), .Z(n19308) );
  NAND U19614 ( .A(n19310), .B(n19309), .Z(n19305) );
  ANDN U19615 ( .B(B[151]), .A(n38), .Z(n19201) );
  XNOR U19616 ( .A(n19209), .B(n19311), .Z(n19202) );
  XNOR U19617 ( .A(n19208), .B(n19206), .Z(n19311) );
  AND U19618 ( .A(n19312), .B(n19313), .Z(n19206) );
  NANDN U19619 ( .A(n19314), .B(n19315), .Z(n19313) );
  NANDN U19620 ( .A(n19316), .B(n19317), .Z(n19315) );
  NANDN U19621 ( .A(n19317), .B(n19316), .Z(n19312) );
  ANDN U19622 ( .B(B[152]), .A(n39), .Z(n19208) );
  XNOR U19623 ( .A(n19216), .B(n19318), .Z(n19209) );
  XNOR U19624 ( .A(n19215), .B(n19213), .Z(n19318) );
  AND U19625 ( .A(n19319), .B(n19320), .Z(n19213) );
  NANDN U19626 ( .A(n19321), .B(n19322), .Z(n19320) );
  OR U19627 ( .A(n19323), .B(n19324), .Z(n19322) );
  NAND U19628 ( .A(n19324), .B(n19323), .Z(n19319) );
  ANDN U19629 ( .B(B[153]), .A(n40), .Z(n19215) );
  XNOR U19630 ( .A(n19223), .B(n19325), .Z(n19216) );
  XNOR U19631 ( .A(n19222), .B(n19220), .Z(n19325) );
  AND U19632 ( .A(n19326), .B(n19327), .Z(n19220) );
  NANDN U19633 ( .A(n19328), .B(n19329), .Z(n19327) );
  NAND U19634 ( .A(n19330), .B(n19331), .Z(n19329) );
  ANDN U19635 ( .B(B[154]), .A(n41), .Z(n19222) );
  XOR U19636 ( .A(n19229), .B(n19332), .Z(n19223) );
  XNOR U19637 ( .A(n19227), .B(n19230), .Z(n19332) );
  NAND U19638 ( .A(A[2]), .B(B[155]), .Z(n19230) );
  NANDN U19639 ( .A(n19333), .B(n19334), .Z(n19227) );
  AND U19640 ( .A(A[0]), .B(B[156]), .Z(n19334) );
  XNOR U19641 ( .A(n19232), .B(n19335), .Z(n19229) );
  NAND U19642 ( .A(A[0]), .B(B[157]), .Z(n19335) );
  NAND U19643 ( .A(B[156]), .B(A[1]), .Z(n19232) );
  NAND U19644 ( .A(n19336), .B(n19337), .Z(n441) );
  NANDN U19645 ( .A(n19338), .B(n19339), .Z(n19337) );
  OR U19646 ( .A(n19340), .B(n19341), .Z(n19339) );
  NAND U19647 ( .A(n19341), .B(n19340), .Z(n19336) );
  XOR U19648 ( .A(n443), .B(n442), .Z(\A1[154] ) );
  XOR U19649 ( .A(n19341), .B(n19342), .Z(n442) );
  XNOR U19650 ( .A(n19340), .B(n19338), .Z(n19342) );
  AND U19651 ( .A(n19343), .B(n19344), .Z(n19338) );
  NANDN U19652 ( .A(n19345), .B(n19346), .Z(n19344) );
  NANDN U19653 ( .A(n19347), .B(n19348), .Z(n19346) );
  NANDN U19654 ( .A(n19348), .B(n19347), .Z(n19343) );
  ANDN U19655 ( .B(B[141]), .A(n29), .Z(n19340) );
  XNOR U19656 ( .A(n19247), .B(n19349), .Z(n19341) );
  XNOR U19657 ( .A(n19246), .B(n19244), .Z(n19349) );
  AND U19658 ( .A(n19350), .B(n19351), .Z(n19244) );
  NANDN U19659 ( .A(n19352), .B(n19353), .Z(n19351) );
  OR U19660 ( .A(n19354), .B(n19355), .Z(n19353) );
  NAND U19661 ( .A(n19355), .B(n19354), .Z(n19350) );
  ANDN U19662 ( .B(B[142]), .A(n30), .Z(n19246) );
  XNOR U19663 ( .A(n19254), .B(n19356), .Z(n19247) );
  XNOR U19664 ( .A(n19253), .B(n19251), .Z(n19356) );
  AND U19665 ( .A(n19357), .B(n19358), .Z(n19251) );
  NANDN U19666 ( .A(n19359), .B(n19360), .Z(n19358) );
  NANDN U19667 ( .A(n19361), .B(n19362), .Z(n19360) );
  NANDN U19668 ( .A(n19362), .B(n19361), .Z(n19357) );
  ANDN U19669 ( .B(B[143]), .A(n31), .Z(n19253) );
  XNOR U19670 ( .A(n19261), .B(n19363), .Z(n19254) );
  XNOR U19671 ( .A(n19260), .B(n19258), .Z(n19363) );
  AND U19672 ( .A(n19364), .B(n19365), .Z(n19258) );
  NANDN U19673 ( .A(n19366), .B(n19367), .Z(n19365) );
  OR U19674 ( .A(n19368), .B(n19369), .Z(n19367) );
  NAND U19675 ( .A(n19369), .B(n19368), .Z(n19364) );
  ANDN U19676 ( .B(B[144]), .A(n32), .Z(n19260) );
  XNOR U19677 ( .A(n19268), .B(n19370), .Z(n19261) );
  XNOR U19678 ( .A(n19267), .B(n19265), .Z(n19370) );
  AND U19679 ( .A(n19371), .B(n19372), .Z(n19265) );
  NANDN U19680 ( .A(n19373), .B(n19374), .Z(n19372) );
  NANDN U19681 ( .A(n19375), .B(n19376), .Z(n19374) );
  NANDN U19682 ( .A(n19376), .B(n19375), .Z(n19371) );
  ANDN U19683 ( .B(B[145]), .A(n33), .Z(n19267) );
  XNOR U19684 ( .A(n19275), .B(n19377), .Z(n19268) );
  XNOR U19685 ( .A(n19274), .B(n19272), .Z(n19377) );
  AND U19686 ( .A(n19378), .B(n19379), .Z(n19272) );
  NANDN U19687 ( .A(n19380), .B(n19381), .Z(n19379) );
  OR U19688 ( .A(n19382), .B(n19383), .Z(n19381) );
  NAND U19689 ( .A(n19383), .B(n19382), .Z(n19378) );
  ANDN U19690 ( .B(B[146]), .A(n34), .Z(n19274) );
  XNOR U19691 ( .A(n19282), .B(n19384), .Z(n19275) );
  XNOR U19692 ( .A(n19281), .B(n19279), .Z(n19384) );
  AND U19693 ( .A(n19385), .B(n19386), .Z(n19279) );
  NANDN U19694 ( .A(n19387), .B(n19388), .Z(n19386) );
  NANDN U19695 ( .A(n19389), .B(n19390), .Z(n19388) );
  NANDN U19696 ( .A(n19390), .B(n19389), .Z(n19385) );
  ANDN U19697 ( .B(B[147]), .A(n35), .Z(n19281) );
  XNOR U19698 ( .A(n19289), .B(n19391), .Z(n19282) );
  XNOR U19699 ( .A(n19288), .B(n19286), .Z(n19391) );
  AND U19700 ( .A(n19392), .B(n19393), .Z(n19286) );
  NANDN U19701 ( .A(n19394), .B(n19395), .Z(n19393) );
  OR U19702 ( .A(n19396), .B(n19397), .Z(n19395) );
  NAND U19703 ( .A(n19397), .B(n19396), .Z(n19392) );
  ANDN U19704 ( .B(B[148]), .A(n36), .Z(n19288) );
  XNOR U19705 ( .A(n19296), .B(n19398), .Z(n19289) );
  XNOR U19706 ( .A(n19295), .B(n19293), .Z(n19398) );
  AND U19707 ( .A(n19399), .B(n19400), .Z(n19293) );
  NANDN U19708 ( .A(n19401), .B(n19402), .Z(n19400) );
  NANDN U19709 ( .A(n19403), .B(n19404), .Z(n19402) );
  NANDN U19710 ( .A(n19404), .B(n19403), .Z(n19399) );
  ANDN U19711 ( .B(B[149]), .A(n37), .Z(n19295) );
  XNOR U19712 ( .A(n19303), .B(n19405), .Z(n19296) );
  XNOR U19713 ( .A(n19302), .B(n19300), .Z(n19405) );
  AND U19714 ( .A(n19406), .B(n19407), .Z(n19300) );
  NANDN U19715 ( .A(n19408), .B(n19409), .Z(n19407) );
  OR U19716 ( .A(n19410), .B(n19411), .Z(n19409) );
  NAND U19717 ( .A(n19411), .B(n19410), .Z(n19406) );
  ANDN U19718 ( .B(B[150]), .A(n38), .Z(n19302) );
  XNOR U19719 ( .A(n19310), .B(n19412), .Z(n19303) );
  XNOR U19720 ( .A(n19309), .B(n19307), .Z(n19412) );
  AND U19721 ( .A(n19413), .B(n19414), .Z(n19307) );
  NANDN U19722 ( .A(n19415), .B(n19416), .Z(n19414) );
  NANDN U19723 ( .A(n19417), .B(n19418), .Z(n19416) );
  NANDN U19724 ( .A(n19418), .B(n19417), .Z(n19413) );
  ANDN U19725 ( .B(B[151]), .A(n39), .Z(n19309) );
  XNOR U19726 ( .A(n19317), .B(n19419), .Z(n19310) );
  XNOR U19727 ( .A(n19316), .B(n19314), .Z(n19419) );
  AND U19728 ( .A(n19420), .B(n19421), .Z(n19314) );
  NANDN U19729 ( .A(n19422), .B(n19423), .Z(n19421) );
  OR U19730 ( .A(n19424), .B(n19425), .Z(n19423) );
  NAND U19731 ( .A(n19425), .B(n19424), .Z(n19420) );
  ANDN U19732 ( .B(B[152]), .A(n40), .Z(n19316) );
  XNOR U19733 ( .A(n19324), .B(n19426), .Z(n19317) );
  XNOR U19734 ( .A(n19323), .B(n19321), .Z(n19426) );
  AND U19735 ( .A(n19427), .B(n19428), .Z(n19321) );
  NANDN U19736 ( .A(n19429), .B(n19430), .Z(n19428) );
  NAND U19737 ( .A(n19431), .B(n19432), .Z(n19430) );
  ANDN U19738 ( .B(B[153]), .A(n41), .Z(n19323) );
  XOR U19739 ( .A(n19330), .B(n19433), .Z(n19324) );
  XNOR U19740 ( .A(n19328), .B(n19331), .Z(n19433) );
  NAND U19741 ( .A(A[2]), .B(B[154]), .Z(n19331) );
  NANDN U19742 ( .A(n19434), .B(n19435), .Z(n19328) );
  AND U19743 ( .A(A[0]), .B(B[155]), .Z(n19435) );
  XNOR U19744 ( .A(n19333), .B(n19436), .Z(n19330) );
  NAND U19745 ( .A(A[0]), .B(B[156]), .Z(n19436) );
  NAND U19746 ( .A(B[155]), .B(A[1]), .Z(n19333) );
  NAND U19747 ( .A(n19437), .B(n19438), .Z(n443) );
  NANDN U19748 ( .A(n19439), .B(n19440), .Z(n19438) );
  OR U19749 ( .A(n19441), .B(n19442), .Z(n19440) );
  NAND U19750 ( .A(n19442), .B(n19441), .Z(n19437) );
  XOR U19751 ( .A(n445), .B(n444), .Z(\A1[153] ) );
  XOR U19752 ( .A(n19442), .B(n19443), .Z(n444) );
  XNOR U19753 ( .A(n19441), .B(n19439), .Z(n19443) );
  AND U19754 ( .A(n19444), .B(n19445), .Z(n19439) );
  NANDN U19755 ( .A(n19446), .B(n19447), .Z(n19445) );
  NANDN U19756 ( .A(n19448), .B(n19449), .Z(n19447) );
  NANDN U19757 ( .A(n19449), .B(n19448), .Z(n19444) );
  ANDN U19758 ( .B(B[140]), .A(n29), .Z(n19441) );
  XNOR U19759 ( .A(n19348), .B(n19450), .Z(n19442) );
  XNOR U19760 ( .A(n19347), .B(n19345), .Z(n19450) );
  AND U19761 ( .A(n19451), .B(n19452), .Z(n19345) );
  NANDN U19762 ( .A(n19453), .B(n19454), .Z(n19452) );
  OR U19763 ( .A(n19455), .B(n19456), .Z(n19454) );
  NAND U19764 ( .A(n19456), .B(n19455), .Z(n19451) );
  ANDN U19765 ( .B(B[141]), .A(n30), .Z(n19347) );
  XNOR U19766 ( .A(n19355), .B(n19457), .Z(n19348) );
  XNOR U19767 ( .A(n19354), .B(n19352), .Z(n19457) );
  AND U19768 ( .A(n19458), .B(n19459), .Z(n19352) );
  NANDN U19769 ( .A(n19460), .B(n19461), .Z(n19459) );
  NANDN U19770 ( .A(n19462), .B(n19463), .Z(n19461) );
  NANDN U19771 ( .A(n19463), .B(n19462), .Z(n19458) );
  ANDN U19772 ( .B(B[142]), .A(n31), .Z(n19354) );
  XNOR U19773 ( .A(n19362), .B(n19464), .Z(n19355) );
  XNOR U19774 ( .A(n19361), .B(n19359), .Z(n19464) );
  AND U19775 ( .A(n19465), .B(n19466), .Z(n19359) );
  NANDN U19776 ( .A(n19467), .B(n19468), .Z(n19466) );
  OR U19777 ( .A(n19469), .B(n19470), .Z(n19468) );
  NAND U19778 ( .A(n19470), .B(n19469), .Z(n19465) );
  ANDN U19779 ( .B(B[143]), .A(n32), .Z(n19361) );
  XNOR U19780 ( .A(n19369), .B(n19471), .Z(n19362) );
  XNOR U19781 ( .A(n19368), .B(n19366), .Z(n19471) );
  AND U19782 ( .A(n19472), .B(n19473), .Z(n19366) );
  NANDN U19783 ( .A(n19474), .B(n19475), .Z(n19473) );
  NANDN U19784 ( .A(n19476), .B(n19477), .Z(n19475) );
  NANDN U19785 ( .A(n19477), .B(n19476), .Z(n19472) );
  ANDN U19786 ( .B(B[144]), .A(n33), .Z(n19368) );
  XNOR U19787 ( .A(n19376), .B(n19478), .Z(n19369) );
  XNOR U19788 ( .A(n19375), .B(n19373), .Z(n19478) );
  AND U19789 ( .A(n19479), .B(n19480), .Z(n19373) );
  NANDN U19790 ( .A(n19481), .B(n19482), .Z(n19480) );
  OR U19791 ( .A(n19483), .B(n19484), .Z(n19482) );
  NAND U19792 ( .A(n19484), .B(n19483), .Z(n19479) );
  ANDN U19793 ( .B(B[145]), .A(n34), .Z(n19375) );
  XNOR U19794 ( .A(n19383), .B(n19485), .Z(n19376) );
  XNOR U19795 ( .A(n19382), .B(n19380), .Z(n19485) );
  AND U19796 ( .A(n19486), .B(n19487), .Z(n19380) );
  NANDN U19797 ( .A(n19488), .B(n19489), .Z(n19487) );
  NANDN U19798 ( .A(n19490), .B(n19491), .Z(n19489) );
  NANDN U19799 ( .A(n19491), .B(n19490), .Z(n19486) );
  ANDN U19800 ( .B(B[146]), .A(n35), .Z(n19382) );
  XNOR U19801 ( .A(n19390), .B(n19492), .Z(n19383) );
  XNOR U19802 ( .A(n19389), .B(n19387), .Z(n19492) );
  AND U19803 ( .A(n19493), .B(n19494), .Z(n19387) );
  NANDN U19804 ( .A(n19495), .B(n19496), .Z(n19494) );
  OR U19805 ( .A(n19497), .B(n19498), .Z(n19496) );
  NAND U19806 ( .A(n19498), .B(n19497), .Z(n19493) );
  ANDN U19807 ( .B(B[147]), .A(n36), .Z(n19389) );
  XNOR U19808 ( .A(n19397), .B(n19499), .Z(n19390) );
  XNOR U19809 ( .A(n19396), .B(n19394), .Z(n19499) );
  AND U19810 ( .A(n19500), .B(n19501), .Z(n19394) );
  NANDN U19811 ( .A(n19502), .B(n19503), .Z(n19501) );
  NANDN U19812 ( .A(n19504), .B(n19505), .Z(n19503) );
  NANDN U19813 ( .A(n19505), .B(n19504), .Z(n19500) );
  ANDN U19814 ( .B(B[148]), .A(n37), .Z(n19396) );
  XNOR U19815 ( .A(n19404), .B(n19506), .Z(n19397) );
  XNOR U19816 ( .A(n19403), .B(n19401), .Z(n19506) );
  AND U19817 ( .A(n19507), .B(n19508), .Z(n19401) );
  NANDN U19818 ( .A(n19509), .B(n19510), .Z(n19508) );
  OR U19819 ( .A(n19511), .B(n19512), .Z(n19510) );
  NAND U19820 ( .A(n19512), .B(n19511), .Z(n19507) );
  ANDN U19821 ( .B(B[149]), .A(n38), .Z(n19403) );
  XNOR U19822 ( .A(n19411), .B(n19513), .Z(n19404) );
  XNOR U19823 ( .A(n19410), .B(n19408), .Z(n19513) );
  AND U19824 ( .A(n19514), .B(n19515), .Z(n19408) );
  NANDN U19825 ( .A(n19516), .B(n19517), .Z(n19515) );
  NANDN U19826 ( .A(n19518), .B(n19519), .Z(n19517) );
  NANDN U19827 ( .A(n19519), .B(n19518), .Z(n19514) );
  ANDN U19828 ( .B(B[150]), .A(n39), .Z(n19410) );
  XNOR U19829 ( .A(n19418), .B(n19520), .Z(n19411) );
  XNOR U19830 ( .A(n19417), .B(n19415), .Z(n19520) );
  AND U19831 ( .A(n19521), .B(n19522), .Z(n19415) );
  NANDN U19832 ( .A(n19523), .B(n19524), .Z(n19522) );
  OR U19833 ( .A(n19525), .B(n19526), .Z(n19524) );
  NAND U19834 ( .A(n19526), .B(n19525), .Z(n19521) );
  ANDN U19835 ( .B(B[151]), .A(n40), .Z(n19417) );
  XNOR U19836 ( .A(n19425), .B(n19527), .Z(n19418) );
  XNOR U19837 ( .A(n19424), .B(n19422), .Z(n19527) );
  AND U19838 ( .A(n19528), .B(n19529), .Z(n19422) );
  NANDN U19839 ( .A(n19530), .B(n19531), .Z(n19529) );
  NAND U19840 ( .A(n19532), .B(n19533), .Z(n19531) );
  ANDN U19841 ( .B(B[152]), .A(n41), .Z(n19424) );
  XOR U19842 ( .A(n19431), .B(n19534), .Z(n19425) );
  XNOR U19843 ( .A(n19429), .B(n19432), .Z(n19534) );
  NAND U19844 ( .A(A[2]), .B(B[153]), .Z(n19432) );
  NANDN U19845 ( .A(n19535), .B(n19536), .Z(n19429) );
  AND U19846 ( .A(A[0]), .B(B[154]), .Z(n19536) );
  XNOR U19847 ( .A(n19434), .B(n19537), .Z(n19431) );
  NAND U19848 ( .A(A[0]), .B(B[155]), .Z(n19537) );
  NAND U19849 ( .A(B[154]), .B(A[1]), .Z(n19434) );
  NAND U19850 ( .A(n19538), .B(n19539), .Z(n445) );
  NANDN U19851 ( .A(n19540), .B(n19541), .Z(n19539) );
  OR U19852 ( .A(n19542), .B(n19543), .Z(n19541) );
  NAND U19853 ( .A(n19543), .B(n19542), .Z(n19538) );
  XOR U19854 ( .A(n447), .B(n446), .Z(\A1[152] ) );
  XOR U19855 ( .A(n19543), .B(n19544), .Z(n446) );
  XNOR U19856 ( .A(n19542), .B(n19540), .Z(n19544) );
  AND U19857 ( .A(n19545), .B(n19546), .Z(n19540) );
  NANDN U19858 ( .A(n19547), .B(n19548), .Z(n19546) );
  NANDN U19859 ( .A(n19549), .B(n19550), .Z(n19548) );
  NANDN U19860 ( .A(n19550), .B(n19549), .Z(n19545) );
  ANDN U19861 ( .B(B[139]), .A(n29), .Z(n19542) );
  XNOR U19862 ( .A(n19449), .B(n19551), .Z(n19543) );
  XNOR U19863 ( .A(n19448), .B(n19446), .Z(n19551) );
  AND U19864 ( .A(n19552), .B(n19553), .Z(n19446) );
  NANDN U19865 ( .A(n19554), .B(n19555), .Z(n19553) );
  OR U19866 ( .A(n19556), .B(n19557), .Z(n19555) );
  NAND U19867 ( .A(n19557), .B(n19556), .Z(n19552) );
  ANDN U19868 ( .B(B[140]), .A(n30), .Z(n19448) );
  XNOR U19869 ( .A(n19456), .B(n19558), .Z(n19449) );
  XNOR U19870 ( .A(n19455), .B(n19453), .Z(n19558) );
  AND U19871 ( .A(n19559), .B(n19560), .Z(n19453) );
  NANDN U19872 ( .A(n19561), .B(n19562), .Z(n19560) );
  NANDN U19873 ( .A(n19563), .B(n19564), .Z(n19562) );
  NANDN U19874 ( .A(n19564), .B(n19563), .Z(n19559) );
  ANDN U19875 ( .B(B[141]), .A(n31), .Z(n19455) );
  XNOR U19876 ( .A(n19463), .B(n19565), .Z(n19456) );
  XNOR U19877 ( .A(n19462), .B(n19460), .Z(n19565) );
  AND U19878 ( .A(n19566), .B(n19567), .Z(n19460) );
  NANDN U19879 ( .A(n19568), .B(n19569), .Z(n19567) );
  OR U19880 ( .A(n19570), .B(n19571), .Z(n19569) );
  NAND U19881 ( .A(n19571), .B(n19570), .Z(n19566) );
  ANDN U19882 ( .B(B[142]), .A(n32), .Z(n19462) );
  XNOR U19883 ( .A(n19470), .B(n19572), .Z(n19463) );
  XNOR U19884 ( .A(n19469), .B(n19467), .Z(n19572) );
  AND U19885 ( .A(n19573), .B(n19574), .Z(n19467) );
  NANDN U19886 ( .A(n19575), .B(n19576), .Z(n19574) );
  NANDN U19887 ( .A(n19577), .B(n19578), .Z(n19576) );
  NANDN U19888 ( .A(n19578), .B(n19577), .Z(n19573) );
  ANDN U19889 ( .B(B[143]), .A(n33), .Z(n19469) );
  XNOR U19890 ( .A(n19477), .B(n19579), .Z(n19470) );
  XNOR U19891 ( .A(n19476), .B(n19474), .Z(n19579) );
  AND U19892 ( .A(n19580), .B(n19581), .Z(n19474) );
  NANDN U19893 ( .A(n19582), .B(n19583), .Z(n19581) );
  OR U19894 ( .A(n19584), .B(n19585), .Z(n19583) );
  NAND U19895 ( .A(n19585), .B(n19584), .Z(n19580) );
  ANDN U19896 ( .B(B[144]), .A(n34), .Z(n19476) );
  XNOR U19897 ( .A(n19484), .B(n19586), .Z(n19477) );
  XNOR U19898 ( .A(n19483), .B(n19481), .Z(n19586) );
  AND U19899 ( .A(n19587), .B(n19588), .Z(n19481) );
  NANDN U19900 ( .A(n19589), .B(n19590), .Z(n19588) );
  NANDN U19901 ( .A(n19591), .B(n19592), .Z(n19590) );
  NANDN U19902 ( .A(n19592), .B(n19591), .Z(n19587) );
  ANDN U19903 ( .B(B[145]), .A(n35), .Z(n19483) );
  XNOR U19904 ( .A(n19491), .B(n19593), .Z(n19484) );
  XNOR U19905 ( .A(n19490), .B(n19488), .Z(n19593) );
  AND U19906 ( .A(n19594), .B(n19595), .Z(n19488) );
  NANDN U19907 ( .A(n19596), .B(n19597), .Z(n19595) );
  OR U19908 ( .A(n19598), .B(n19599), .Z(n19597) );
  NAND U19909 ( .A(n19599), .B(n19598), .Z(n19594) );
  ANDN U19910 ( .B(B[146]), .A(n36), .Z(n19490) );
  XNOR U19911 ( .A(n19498), .B(n19600), .Z(n19491) );
  XNOR U19912 ( .A(n19497), .B(n19495), .Z(n19600) );
  AND U19913 ( .A(n19601), .B(n19602), .Z(n19495) );
  NANDN U19914 ( .A(n19603), .B(n19604), .Z(n19602) );
  NANDN U19915 ( .A(n19605), .B(n19606), .Z(n19604) );
  NANDN U19916 ( .A(n19606), .B(n19605), .Z(n19601) );
  ANDN U19917 ( .B(B[147]), .A(n37), .Z(n19497) );
  XNOR U19918 ( .A(n19505), .B(n19607), .Z(n19498) );
  XNOR U19919 ( .A(n19504), .B(n19502), .Z(n19607) );
  AND U19920 ( .A(n19608), .B(n19609), .Z(n19502) );
  NANDN U19921 ( .A(n19610), .B(n19611), .Z(n19609) );
  OR U19922 ( .A(n19612), .B(n19613), .Z(n19611) );
  NAND U19923 ( .A(n19613), .B(n19612), .Z(n19608) );
  ANDN U19924 ( .B(B[148]), .A(n38), .Z(n19504) );
  XNOR U19925 ( .A(n19512), .B(n19614), .Z(n19505) );
  XNOR U19926 ( .A(n19511), .B(n19509), .Z(n19614) );
  AND U19927 ( .A(n19615), .B(n19616), .Z(n19509) );
  NANDN U19928 ( .A(n19617), .B(n19618), .Z(n19616) );
  NANDN U19929 ( .A(n19619), .B(n19620), .Z(n19618) );
  NANDN U19930 ( .A(n19620), .B(n19619), .Z(n19615) );
  ANDN U19931 ( .B(B[149]), .A(n39), .Z(n19511) );
  XNOR U19932 ( .A(n19519), .B(n19621), .Z(n19512) );
  XNOR U19933 ( .A(n19518), .B(n19516), .Z(n19621) );
  AND U19934 ( .A(n19622), .B(n19623), .Z(n19516) );
  NANDN U19935 ( .A(n19624), .B(n19625), .Z(n19623) );
  OR U19936 ( .A(n19626), .B(n19627), .Z(n19625) );
  NAND U19937 ( .A(n19627), .B(n19626), .Z(n19622) );
  ANDN U19938 ( .B(B[150]), .A(n40), .Z(n19518) );
  XNOR U19939 ( .A(n19526), .B(n19628), .Z(n19519) );
  XNOR U19940 ( .A(n19525), .B(n19523), .Z(n19628) );
  AND U19941 ( .A(n19629), .B(n19630), .Z(n19523) );
  NANDN U19942 ( .A(n19631), .B(n19632), .Z(n19630) );
  NAND U19943 ( .A(n19633), .B(n19634), .Z(n19632) );
  ANDN U19944 ( .B(B[151]), .A(n41), .Z(n19525) );
  XOR U19945 ( .A(n19532), .B(n19635), .Z(n19526) );
  XNOR U19946 ( .A(n19530), .B(n19533), .Z(n19635) );
  NAND U19947 ( .A(A[2]), .B(B[152]), .Z(n19533) );
  NANDN U19948 ( .A(n19636), .B(n19637), .Z(n19530) );
  AND U19949 ( .A(A[0]), .B(B[153]), .Z(n19637) );
  XNOR U19950 ( .A(n19535), .B(n19638), .Z(n19532) );
  NAND U19951 ( .A(A[0]), .B(B[154]), .Z(n19638) );
  NAND U19952 ( .A(B[153]), .B(A[1]), .Z(n19535) );
  NAND U19953 ( .A(n19639), .B(n19640), .Z(n447) );
  NANDN U19954 ( .A(n19641), .B(n19642), .Z(n19640) );
  OR U19955 ( .A(n19643), .B(n19644), .Z(n19642) );
  NAND U19956 ( .A(n19644), .B(n19643), .Z(n19639) );
  XOR U19957 ( .A(n449), .B(n448), .Z(\A1[151] ) );
  XOR U19958 ( .A(n19644), .B(n19645), .Z(n448) );
  XNOR U19959 ( .A(n19643), .B(n19641), .Z(n19645) );
  AND U19960 ( .A(n19646), .B(n19647), .Z(n19641) );
  NANDN U19961 ( .A(n19648), .B(n19649), .Z(n19647) );
  NANDN U19962 ( .A(n19650), .B(n19651), .Z(n19649) );
  NANDN U19963 ( .A(n19651), .B(n19650), .Z(n19646) );
  ANDN U19964 ( .B(B[138]), .A(n29), .Z(n19643) );
  XNOR U19965 ( .A(n19550), .B(n19652), .Z(n19644) );
  XNOR U19966 ( .A(n19549), .B(n19547), .Z(n19652) );
  AND U19967 ( .A(n19653), .B(n19654), .Z(n19547) );
  NANDN U19968 ( .A(n19655), .B(n19656), .Z(n19654) );
  OR U19969 ( .A(n19657), .B(n19658), .Z(n19656) );
  NAND U19970 ( .A(n19658), .B(n19657), .Z(n19653) );
  ANDN U19971 ( .B(B[139]), .A(n30), .Z(n19549) );
  XNOR U19972 ( .A(n19557), .B(n19659), .Z(n19550) );
  XNOR U19973 ( .A(n19556), .B(n19554), .Z(n19659) );
  AND U19974 ( .A(n19660), .B(n19661), .Z(n19554) );
  NANDN U19975 ( .A(n19662), .B(n19663), .Z(n19661) );
  NANDN U19976 ( .A(n19664), .B(n19665), .Z(n19663) );
  NANDN U19977 ( .A(n19665), .B(n19664), .Z(n19660) );
  ANDN U19978 ( .B(B[140]), .A(n31), .Z(n19556) );
  XNOR U19979 ( .A(n19564), .B(n19666), .Z(n19557) );
  XNOR U19980 ( .A(n19563), .B(n19561), .Z(n19666) );
  AND U19981 ( .A(n19667), .B(n19668), .Z(n19561) );
  NANDN U19982 ( .A(n19669), .B(n19670), .Z(n19668) );
  OR U19983 ( .A(n19671), .B(n19672), .Z(n19670) );
  NAND U19984 ( .A(n19672), .B(n19671), .Z(n19667) );
  ANDN U19985 ( .B(B[141]), .A(n32), .Z(n19563) );
  XNOR U19986 ( .A(n19571), .B(n19673), .Z(n19564) );
  XNOR U19987 ( .A(n19570), .B(n19568), .Z(n19673) );
  AND U19988 ( .A(n19674), .B(n19675), .Z(n19568) );
  NANDN U19989 ( .A(n19676), .B(n19677), .Z(n19675) );
  NANDN U19990 ( .A(n19678), .B(n19679), .Z(n19677) );
  NANDN U19991 ( .A(n19679), .B(n19678), .Z(n19674) );
  ANDN U19992 ( .B(B[142]), .A(n33), .Z(n19570) );
  XNOR U19993 ( .A(n19578), .B(n19680), .Z(n19571) );
  XNOR U19994 ( .A(n19577), .B(n19575), .Z(n19680) );
  AND U19995 ( .A(n19681), .B(n19682), .Z(n19575) );
  NANDN U19996 ( .A(n19683), .B(n19684), .Z(n19682) );
  OR U19997 ( .A(n19685), .B(n19686), .Z(n19684) );
  NAND U19998 ( .A(n19686), .B(n19685), .Z(n19681) );
  ANDN U19999 ( .B(B[143]), .A(n34), .Z(n19577) );
  XNOR U20000 ( .A(n19585), .B(n19687), .Z(n19578) );
  XNOR U20001 ( .A(n19584), .B(n19582), .Z(n19687) );
  AND U20002 ( .A(n19688), .B(n19689), .Z(n19582) );
  NANDN U20003 ( .A(n19690), .B(n19691), .Z(n19689) );
  NANDN U20004 ( .A(n19692), .B(n19693), .Z(n19691) );
  NANDN U20005 ( .A(n19693), .B(n19692), .Z(n19688) );
  ANDN U20006 ( .B(B[144]), .A(n35), .Z(n19584) );
  XNOR U20007 ( .A(n19592), .B(n19694), .Z(n19585) );
  XNOR U20008 ( .A(n19591), .B(n19589), .Z(n19694) );
  AND U20009 ( .A(n19695), .B(n19696), .Z(n19589) );
  NANDN U20010 ( .A(n19697), .B(n19698), .Z(n19696) );
  OR U20011 ( .A(n19699), .B(n19700), .Z(n19698) );
  NAND U20012 ( .A(n19700), .B(n19699), .Z(n19695) );
  ANDN U20013 ( .B(B[145]), .A(n36), .Z(n19591) );
  XNOR U20014 ( .A(n19599), .B(n19701), .Z(n19592) );
  XNOR U20015 ( .A(n19598), .B(n19596), .Z(n19701) );
  AND U20016 ( .A(n19702), .B(n19703), .Z(n19596) );
  NANDN U20017 ( .A(n19704), .B(n19705), .Z(n19703) );
  NANDN U20018 ( .A(n19706), .B(n19707), .Z(n19705) );
  NANDN U20019 ( .A(n19707), .B(n19706), .Z(n19702) );
  ANDN U20020 ( .B(B[146]), .A(n37), .Z(n19598) );
  XNOR U20021 ( .A(n19606), .B(n19708), .Z(n19599) );
  XNOR U20022 ( .A(n19605), .B(n19603), .Z(n19708) );
  AND U20023 ( .A(n19709), .B(n19710), .Z(n19603) );
  NANDN U20024 ( .A(n19711), .B(n19712), .Z(n19710) );
  OR U20025 ( .A(n19713), .B(n19714), .Z(n19712) );
  NAND U20026 ( .A(n19714), .B(n19713), .Z(n19709) );
  ANDN U20027 ( .B(B[147]), .A(n38), .Z(n19605) );
  XNOR U20028 ( .A(n19613), .B(n19715), .Z(n19606) );
  XNOR U20029 ( .A(n19612), .B(n19610), .Z(n19715) );
  AND U20030 ( .A(n19716), .B(n19717), .Z(n19610) );
  NANDN U20031 ( .A(n19718), .B(n19719), .Z(n19717) );
  NANDN U20032 ( .A(n19720), .B(n19721), .Z(n19719) );
  NANDN U20033 ( .A(n19721), .B(n19720), .Z(n19716) );
  ANDN U20034 ( .B(B[148]), .A(n39), .Z(n19612) );
  XNOR U20035 ( .A(n19620), .B(n19722), .Z(n19613) );
  XNOR U20036 ( .A(n19619), .B(n19617), .Z(n19722) );
  AND U20037 ( .A(n19723), .B(n19724), .Z(n19617) );
  NANDN U20038 ( .A(n19725), .B(n19726), .Z(n19724) );
  OR U20039 ( .A(n19727), .B(n19728), .Z(n19726) );
  NAND U20040 ( .A(n19728), .B(n19727), .Z(n19723) );
  ANDN U20041 ( .B(B[149]), .A(n40), .Z(n19619) );
  XNOR U20042 ( .A(n19627), .B(n19729), .Z(n19620) );
  XNOR U20043 ( .A(n19626), .B(n19624), .Z(n19729) );
  AND U20044 ( .A(n19730), .B(n19731), .Z(n19624) );
  NANDN U20045 ( .A(n19732), .B(n19733), .Z(n19731) );
  NAND U20046 ( .A(n19734), .B(n19735), .Z(n19733) );
  ANDN U20047 ( .B(B[150]), .A(n41), .Z(n19626) );
  XOR U20048 ( .A(n19633), .B(n19736), .Z(n19627) );
  XNOR U20049 ( .A(n19631), .B(n19634), .Z(n19736) );
  NAND U20050 ( .A(A[2]), .B(B[151]), .Z(n19634) );
  NANDN U20051 ( .A(n19737), .B(n19738), .Z(n19631) );
  AND U20052 ( .A(A[0]), .B(B[152]), .Z(n19738) );
  XNOR U20053 ( .A(n19636), .B(n19739), .Z(n19633) );
  NAND U20054 ( .A(A[0]), .B(B[153]), .Z(n19739) );
  NAND U20055 ( .A(B[152]), .B(A[1]), .Z(n19636) );
  NAND U20056 ( .A(n19740), .B(n19741), .Z(n449) );
  NANDN U20057 ( .A(n19742), .B(n19743), .Z(n19741) );
  OR U20058 ( .A(n19744), .B(n19745), .Z(n19743) );
  NAND U20059 ( .A(n19745), .B(n19744), .Z(n19740) );
  XOR U20060 ( .A(n451), .B(n450), .Z(\A1[150] ) );
  XOR U20061 ( .A(n19745), .B(n19746), .Z(n450) );
  XNOR U20062 ( .A(n19744), .B(n19742), .Z(n19746) );
  AND U20063 ( .A(n19747), .B(n19748), .Z(n19742) );
  NANDN U20064 ( .A(n19749), .B(n19750), .Z(n19748) );
  NANDN U20065 ( .A(n19751), .B(n19752), .Z(n19750) );
  NANDN U20066 ( .A(n19752), .B(n19751), .Z(n19747) );
  ANDN U20067 ( .B(B[137]), .A(n29), .Z(n19744) );
  XNOR U20068 ( .A(n19651), .B(n19753), .Z(n19745) );
  XNOR U20069 ( .A(n19650), .B(n19648), .Z(n19753) );
  AND U20070 ( .A(n19754), .B(n19755), .Z(n19648) );
  NANDN U20071 ( .A(n19756), .B(n19757), .Z(n19755) );
  OR U20072 ( .A(n19758), .B(n19759), .Z(n19757) );
  NAND U20073 ( .A(n19759), .B(n19758), .Z(n19754) );
  ANDN U20074 ( .B(B[138]), .A(n30), .Z(n19650) );
  XNOR U20075 ( .A(n19658), .B(n19760), .Z(n19651) );
  XNOR U20076 ( .A(n19657), .B(n19655), .Z(n19760) );
  AND U20077 ( .A(n19761), .B(n19762), .Z(n19655) );
  NANDN U20078 ( .A(n19763), .B(n19764), .Z(n19762) );
  NANDN U20079 ( .A(n19765), .B(n19766), .Z(n19764) );
  NANDN U20080 ( .A(n19766), .B(n19765), .Z(n19761) );
  ANDN U20081 ( .B(B[139]), .A(n31), .Z(n19657) );
  XNOR U20082 ( .A(n19665), .B(n19767), .Z(n19658) );
  XNOR U20083 ( .A(n19664), .B(n19662), .Z(n19767) );
  AND U20084 ( .A(n19768), .B(n19769), .Z(n19662) );
  NANDN U20085 ( .A(n19770), .B(n19771), .Z(n19769) );
  OR U20086 ( .A(n19772), .B(n19773), .Z(n19771) );
  NAND U20087 ( .A(n19773), .B(n19772), .Z(n19768) );
  ANDN U20088 ( .B(B[140]), .A(n32), .Z(n19664) );
  XNOR U20089 ( .A(n19672), .B(n19774), .Z(n19665) );
  XNOR U20090 ( .A(n19671), .B(n19669), .Z(n19774) );
  AND U20091 ( .A(n19775), .B(n19776), .Z(n19669) );
  NANDN U20092 ( .A(n19777), .B(n19778), .Z(n19776) );
  NANDN U20093 ( .A(n19779), .B(n19780), .Z(n19778) );
  NANDN U20094 ( .A(n19780), .B(n19779), .Z(n19775) );
  ANDN U20095 ( .B(B[141]), .A(n33), .Z(n19671) );
  XNOR U20096 ( .A(n19679), .B(n19781), .Z(n19672) );
  XNOR U20097 ( .A(n19678), .B(n19676), .Z(n19781) );
  AND U20098 ( .A(n19782), .B(n19783), .Z(n19676) );
  NANDN U20099 ( .A(n19784), .B(n19785), .Z(n19783) );
  OR U20100 ( .A(n19786), .B(n19787), .Z(n19785) );
  NAND U20101 ( .A(n19787), .B(n19786), .Z(n19782) );
  ANDN U20102 ( .B(B[142]), .A(n34), .Z(n19678) );
  XNOR U20103 ( .A(n19686), .B(n19788), .Z(n19679) );
  XNOR U20104 ( .A(n19685), .B(n19683), .Z(n19788) );
  AND U20105 ( .A(n19789), .B(n19790), .Z(n19683) );
  NANDN U20106 ( .A(n19791), .B(n19792), .Z(n19790) );
  NANDN U20107 ( .A(n19793), .B(n19794), .Z(n19792) );
  NANDN U20108 ( .A(n19794), .B(n19793), .Z(n19789) );
  ANDN U20109 ( .B(B[143]), .A(n35), .Z(n19685) );
  XNOR U20110 ( .A(n19693), .B(n19795), .Z(n19686) );
  XNOR U20111 ( .A(n19692), .B(n19690), .Z(n19795) );
  AND U20112 ( .A(n19796), .B(n19797), .Z(n19690) );
  NANDN U20113 ( .A(n19798), .B(n19799), .Z(n19797) );
  OR U20114 ( .A(n19800), .B(n19801), .Z(n19799) );
  NAND U20115 ( .A(n19801), .B(n19800), .Z(n19796) );
  ANDN U20116 ( .B(B[144]), .A(n36), .Z(n19692) );
  XNOR U20117 ( .A(n19700), .B(n19802), .Z(n19693) );
  XNOR U20118 ( .A(n19699), .B(n19697), .Z(n19802) );
  AND U20119 ( .A(n19803), .B(n19804), .Z(n19697) );
  NANDN U20120 ( .A(n19805), .B(n19806), .Z(n19804) );
  NANDN U20121 ( .A(n19807), .B(n19808), .Z(n19806) );
  NANDN U20122 ( .A(n19808), .B(n19807), .Z(n19803) );
  ANDN U20123 ( .B(B[145]), .A(n37), .Z(n19699) );
  XNOR U20124 ( .A(n19707), .B(n19809), .Z(n19700) );
  XNOR U20125 ( .A(n19706), .B(n19704), .Z(n19809) );
  AND U20126 ( .A(n19810), .B(n19811), .Z(n19704) );
  NANDN U20127 ( .A(n19812), .B(n19813), .Z(n19811) );
  OR U20128 ( .A(n19814), .B(n19815), .Z(n19813) );
  NAND U20129 ( .A(n19815), .B(n19814), .Z(n19810) );
  ANDN U20130 ( .B(B[146]), .A(n38), .Z(n19706) );
  XNOR U20131 ( .A(n19714), .B(n19816), .Z(n19707) );
  XNOR U20132 ( .A(n19713), .B(n19711), .Z(n19816) );
  AND U20133 ( .A(n19817), .B(n19818), .Z(n19711) );
  NANDN U20134 ( .A(n19819), .B(n19820), .Z(n19818) );
  NANDN U20135 ( .A(n19821), .B(n19822), .Z(n19820) );
  NANDN U20136 ( .A(n19822), .B(n19821), .Z(n19817) );
  ANDN U20137 ( .B(B[147]), .A(n39), .Z(n19713) );
  XNOR U20138 ( .A(n19721), .B(n19823), .Z(n19714) );
  XNOR U20139 ( .A(n19720), .B(n19718), .Z(n19823) );
  AND U20140 ( .A(n19824), .B(n19825), .Z(n19718) );
  NANDN U20141 ( .A(n19826), .B(n19827), .Z(n19825) );
  OR U20142 ( .A(n19828), .B(n19829), .Z(n19827) );
  NAND U20143 ( .A(n19829), .B(n19828), .Z(n19824) );
  ANDN U20144 ( .B(B[148]), .A(n40), .Z(n19720) );
  XNOR U20145 ( .A(n19728), .B(n19830), .Z(n19721) );
  XNOR U20146 ( .A(n19727), .B(n19725), .Z(n19830) );
  AND U20147 ( .A(n19831), .B(n19832), .Z(n19725) );
  NANDN U20148 ( .A(n19833), .B(n19834), .Z(n19832) );
  NAND U20149 ( .A(n19835), .B(n19836), .Z(n19834) );
  ANDN U20150 ( .B(B[149]), .A(n41), .Z(n19727) );
  XOR U20151 ( .A(n19734), .B(n19837), .Z(n19728) );
  XNOR U20152 ( .A(n19732), .B(n19735), .Z(n19837) );
  NAND U20153 ( .A(A[2]), .B(B[150]), .Z(n19735) );
  NANDN U20154 ( .A(n19838), .B(n19839), .Z(n19732) );
  AND U20155 ( .A(A[0]), .B(B[151]), .Z(n19839) );
  XNOR U20156 ( .A(n19737), .B(n19840), .Z(n19734) );
  NAND U20157 ( .A(A[0]), .B(B[152]), .Z(n19840) );
  NAND U20158 ( .A(B[151]), .B(A[1]), .Z(n19737) );
  NAND U20159 ( .A(n19841), .B(n19842), .Z(n451) );
  NANDN U20160 ( .A(n19843), .B(n19844), .Z(n19842) );
  OR U20161 ( .A(n19845), .B(n19846), .Z(n19844) );
  NAND U20162 ( .A(n19846), .B(n19845), .Z(n19841) );
  XOR U20163 ( .A(n433), .B(n432), .Z(\A1[14] ) );
  XOR U20164 ( .A(n18836), .B(n19847), .Z(n432) );
  XNOR U20165 ( .A(n18835), .B(n18833), .Z(n19847) );
  AND U20166 ( .A(n19848), .B(n19849), .Z(n18833) );
  NANDN U20167 ( .A(n19850), .B(n19851), .Z(n19849) );
  NANDN U20168 ( .A(n19852), .B(n19853), .Z(n19851) );
  NANDN U20169 ( .A(n19853), .B(n19852), .Z(n19848) );
  ANDN U20170 ( .B(B[1]), .A(n29), .Z(n18835) );
  XNOR U20171 ( .A(n18742), .B(n19854), .Z(n18836) );
  XNOR U20172 ( .A(n18741), .B(n18739), .Z(n19854) );
  AND U20173 ( .A(n19855), .B(n19856), .Z(n18739) );
  NANDN U20174 ( .A(n19857), .B(n19858), .Z(n19856) );
  OR U20175 ( .A(n19859), .B(n19860), .Z(n19858) );
  NAND U20176 ( .A(n19860), .B(n19859), .Z(n19855) );
  ANDN U20177 ( .B(B[2]), .A(n30), .Z(n18741) );
  XNOR U20178 ( .A(n18749), .B(n19861), .Z(n18742) );
  XNOR U20179 ( .A(n18748), .B(n18746), .Z(n19861) );
  AND U20180 ( .A(n19862), .B(n19863), .Z(n18746) );
  NANDN U20181 ( .A(n19864), .B(n19865), .Z(n19863) );
  NANDN U20182 ( .A(n19866), .B(n19867), .Z(n19865) );
  NANDN U20183 ( .A(n19867), .B(n19866), .Z(n19862) );
  ANDN U20184 ( .B(B[3]), .A(n31), .Z(n18748) );
  XNOR U20185 ( .A(n18756), .B(n19868), .Z(n18749) );
  XNOR U20186 ( .A(n18755), .B(n18753), .Z(n19868) );
  AND U20187 ( .A(n19869), .B(n19870), .Z(n18753) );
  NANDN U20188 ( .A(n19871), .B(n19872), .Z(n19870) );
  OR U20189 ( .A(n19873), .B(n19874), .Z(n19872) );
  NAND U20190 ( .A(n19874), .B(n19873), .Z(n19869) );
  ANDN U20191 ( .B(B[4]), .A(n32), .Z(n18755) );
  XNOR U20192 ( .A(n18763), .B(n19875), .Z(n18756) );
  XNOR U20193 ( .A(n18762), .B(n18760), .Z(n19875) );
  AND U20194 ( .A(n19876), .B(n19877), .Z(n18760) );
  NANDN U20195 ( .A(n19878), .B(n19879), .Z(n19877) );
  NANDN U20196 ( .A(n19880), .B(n19881), .Z(n19879) );
  NANDN U20197 ( .A(n19881), .B(n19880), .Z(n19876) );
  ANDN U20198 ( .B(B[5]), .A(n33), .Z(n18762) );
  XNOR U20199 ( .A(n18770), .B(n19882), .Z(n18763) );
  XNOR U20200 ( .A(n18769), .B(n18767), .Z(n19882) );
  AND U20201 ( .A(n19883), .B(n19884), .Z(n18767) );
  NANDN U20202 ( .A(n19885), .B(n19886), .Z(n19884) );
  OR U20203 ( .A(n19887), .B(n19888), .Z(n19886) );
  NAND U20204 ( .A(n19888), .B(n19887), .Z(n19883) );
  ANDN U20205 ( .B(B[6]), .A(n34), .Z(n18769) );
  XNOR U20206 ( .A(n18777), .B(n19889), .Z(n18770) );
  XNOR U20207 ( .A(n18776), .B(n18774), .Z(n19889) );
  AND U20208 ( .A(n19890), .B(n19891), .Z(n18774) );
  NANDN U20209 ( .A(n19892), .B(n19893), .Z(n19891) );
  NANDN U20210 ( .A(n19894), .B(n19895), .Z(n19893) );
  NANDN U20211 ( .A(n19895), .B(n19894), .Z(n19890) );
  ANDN U20212 ( .B(B[7]), .A(n35), .Z(n18776) );
  XNOR U20213 ( .A(n18784), .B(n19896), .Z(n18777) );
  XNOR U20214 ( .A(n18783), .B(n18781), .Z(n19896) );
  AND U20215 ( .A(n19897), .B(n19898), .Z(n18781) );
  NANDN U20216 ( .A(n19899), .B(n19900), .Z(n19898) );
  OR U20217 ( .A(n19901), .B(n19902), .Z(n19900) );
  NAND U20218 ( .A(n19902), .B(n19901), .Z(n19897) );
  ANDN U20219 ( .B(B[8]), .A(n36), .Z(n18783) );
  XNOR U20220 ( .A(n18791), .B(n19903), .Z(n18784) );
  XNOR U20221 ( .A(n18790), .B(n18788), .Z(n19903) );
  AND U20222 ( .A(n19904), .B(n19905), .Z(n18788) );
  NANDN U20223 ( .A(n19906), .B(n19907), .Z(n19905) );
  NANDN U20224 ( .A(n19908), .B(n19909), .Z(n19907) );
  NANDN U20225 ( .A(n19909), .B(n19908), .Z(n19904) );
  ANDN U20226 ( .B(B[9]), .A(n37), .Z(n18790) );
  XNOR U20227 ( .A(n18798), .B(n19910), .Z(n18791) );
  XNOR U20228 ( .A(n18797), .B(n18795), .Z(n19910) );
  AND U20229 ( .A(n19911), .B(n19912), .Z(n18795) );
  NANDN U20230 ( .A(n19913), .B(n19914), .Z(n19912) );
  OR U20231 ( .A(n19915), .B(n19916), .Z(n19914) );
  NAND U20232 ( .A(n19916), .B(n19915), .Z(n19911) );
  ANDN U20233 ( .B(B[10]), .A(n38), .Z(n18797) );
  XNOR U20234 ( .A(n18805), .B(n19917), .Z(n18798) );
  XNOR U20235 ( .A(n18804), .B(n18802), .Z(n19917) );
  AND U20236 ( .A(n19918), .B(n19919), .Z(n18802) );
  NANDN U20237 ( .A(n19920), .B(n19921), .Z(n19919) );
  NANDN U20238 ( .A(n19922), .B(n19923), .Z(n19921) );
  NANDN U20239 ( .A(n19923), .B(n19922), .Z(n19918) );
  ANDN U20240 ( .B(B[11]), .A(n39), .Z(n18804) );
  XNOR U20241 ( .A(n18812), .B(n19924), .Z(n18805) );
  XNOR U20242 ( .A(n18811), .B(n18809), .Z(n19924) );
  AND U20243 ( .A(n19925), .B(n19926), .Z(n18809) );
  NANDN U20244 ( .A(n19927), .B(n19928), .Z(n19926) );
  OR U20245 ( .A(n19929), .B(n19930), .Z(n19928) );
  NAND U20246 ( .A(n19930), .B(n19929), .Z(n19925) );
  ANDN U20247 ( .B(B[12]), .A(n40), .Z(n18811) );
  XNOR U20248 ( .A(n18819), .B(n19931), .Z(n18812) );
  XNOR U20249 ( .A(n18818), .B(n18816), .Z(n19931) );
  AND U20250 ( .A(n19932), .B(n19933), .Z(n18816) );
  NANDN U20251 ( .A(n19934), .B(n19935), .Z(n19933) );
  NAND U20252 ( .A(n19936), .B(n19937), .Z(n19935) );
  ANDN U20253 ( .B(B[13]), .A(n41), .Z(n18818) );
  XOR U20254 ( .A(n18825), .B(n19938), .Z(n18819) );
  XNOR U20255 ( .A(n18823), .B(n18826), .Z(n19938) );
  NAND U20256 ( .A(A[2]), .B(B[14]), .Z(n18826) );
  NANDN U20257 ( .A(n19939), .B(n19940), .Z(n18823) );
  AND U20258 ( .A(A[0]), .B(B[15]), .Z(n19940) );
  XNOR U20259 ( .A(n18828), .B(n19941), .Z(n18825) );
  NAND U20260 ( .A(A[0]), .B(B[16]), .Z(n19941) );
  NAND U20261 ( .A(B[15]), .B(A[1]), .Z(n18828) );
  NAND U20262 ( .A(n19942), .B(n19943), .Z(n433) );
  NANDN U20263 ( .A(n19944), .B(n19945), .Z(n19943) );
  OR U20264 ( .A(n19946), .B(n19947), .Z(n19945) );
  NAND U20265 ( .A(n19947), .B(n19946), .Z(n19942) );
  XOR U20266 ( .A(n453), .B(n452), .Z(\A1[149] ) );
  XOR U20267 ( .A(n19846), .B(n19948), .Z(n452) );
  XNOR U20268 ( .A(n19845), .B(n19843), .Z(n19948) );
  AND U20269 ( .A(n19949), .B(n19950), .Z(n19843) );
  NANDN U20270 ( .A(n19951), .B(n19952), .Z(n19950) );
  NANDN U20271 ( .A(n19953), .B(n19954), .Z(n19952) );
  NANDN U20272 ( .A(n19954), .B(n19953), .Z(n19949) );
  ANDN U20273 ( .B(B[136]), .A(n29), .Z(n19845) );
  XNOR U20274 ( .A(n19752), .B(n19955), .Z(n19846) );
  XNOR U20275 ( .A(n19751), .B(n19749), .Z(n19955) );
  AND U20276 ( .A(n19956), .B(n19957), .Z(n19749) );
  NANDN U20277 ( .A(n19958), .B(n19959), .Z(n19957) );
  OR U20278 ( .A(n19960), .B(n19961), .Z(n19959) );
  NAND U20279 ( .A(n19961), .B(n19960), .Z(n19956) );
  ANDN U20280 ( .B(B[137]), .A(n30), .Z(n19751) );
  XNOR U20281 ( .A(n19759), .B(n19962), .Z(n19752) );
  XNOR U20282 ( .A(n19758), .B(n19756), .Z(n19962) );
  AND U20283 ( .A(n19963), .B(n19964), .Z(n19756) );
  NANDN U20284 ( .A(n19965), .B(n19966), .Z(n19964) );
  NANDN U20285 ( .A(n19967), .B(n19968), .Z(n19966) );
  NANDN U20286 ( .A(n19968), .B(n19967), .Z(n19963) );
  ANDN U20287 ( .B(B[138]), .A(n31), .Z(n19758) );
  XNOR U20288 ( .A(n19766), .B(n19969), .Z(n19759) );
  XNOR U20289 ( .A(n19765), .B(n19763), .Z(n19969) );
  AND U20290 ( .A(n19970), .B(n19971), .Z(n19763) );
  NANDN U20291 ( .A(n19972), .B(n19973), .Z(n19971) );
  OR U20292 ( .A(n19974), .B(n19975), .Z(n19973) );
  NAND U20293 ( .A(n19975), .B(n19974), .Z(n19970) );
  ANDN U20294 ( .B(B[139]), .A(n32), .Z(n19765) );
  XNOR U20295 ( .A(n19773), .B(n19976), .Z(n19766) );
  XNOR U20296 ( .A(n19772), .B(n19770), .Z(n19976) );
  AND U20297 ( .A(n19977), .B(n19978), .Z(n19770) );
  NANDN U20298 ( .A(n19979), .B(n19980), .Z(n19978) );
  NANDN U20299 ( .A(n19981), .B(n19982), .Z(n19980) );
  NANDN U20300 ( .A(n19982), .B(n19981), .Z(n19977) );
  ANDN U20301 ( .B(B[140]), .A(n33), .Z(n19772) );
  XNOR U20302 ( .A(n19780), .B(n19983), .Z(n19773) );
  XNOR U20303 ( .A(n19779), .B(n19777), .Z(n19983) );
  AND U20304 ( .A(n19984), .B(n19985), .Z(n19777) );
  NANDN U20305 ( .A(n19986), .B(n19987), .Z(n19985) );
  OR U20306 ( .A(n19988), .B(n19989), .Z(n19987) );
  NAND U20307 ( .A(n19989), .B(n19988), .Z(n19984) );
  ANDN U20308 ( .B(B[141]), .A(n34), .Z(n19779) );
  XNOR U20309 ( .A(n19787), .B(n19990), .Z(n19780) );
  XNOR U20310 ( .A(n19786), .B(n19784), .Z(n19990) );
  AND U20311 ( .A(n19991), .B(n19992), .Z(n19784) );
  NANDN U20312 ( .A(n19993), .B(n19994), .Z(n19992) );
  NANDN U20313 ( .A(n19995), .B(n19996), .Z(n19994) );
  NANDN U20314 ( .A(n19996), .B(n19995), .Z(n19991) );
  ANDN U20315 ( .B(B[142]), .A(n35), .Z(n19786) );
  XNOR U20316 ( .A(n19794), .B(n19997), .Z(n19787) );
  XNOR U20317 ( .A(n19793), .B(n19791), .Z(n19997) );
  AND U20318 ( .A(n19998), .B(n19999), .Z(n19791) );
  NANDN U20319 ( .A(n20000), .B(n20001), .Z(n19999) );
  OR U20320 ( .A(n20002), .B(n20003), .Z(n20001) );
  NAND U20321 ( .A(n20003), .B(n20002), .Z(n19998) );
  ANDN U20322 ( .B(B[143]), .A(n36), .Z(n19793) );
  XNOR U20323 ( .A(n19801), .B(n20004), .Z(n19794) );
  XNOR U20324 ( .A(n19800), .B(n19798), .Z(n20004) );
  AND U20325 ( .A(n20005), .B(n20006), .Z(n19798) );
  NANDN U20326 ( .A(n20007), .B(n20008), .Z(n20006) );
  NANDN U20327 ( .A(n20009), .B(n20010), .Z(n20008) );
  NANDN U20328 ( .A(n20010), .B(n20009), .Z(n20005) );
  ANDN U20329 ( .B(B[144]), .A(n37), .Z(n19800) );
  XNOR U20330 ( .A(n19808), .B(n20011), .Z(n19801) );
  XNOR U20331 ( .A(n19807), .B(n19805), .Z(n20011) );
  AND U20332 ( .A(n20012), .B(n20013), .Z(n19805) );
  NANDN U20333 ( .A(n20014), .B(n20015), .Z(n20013) );
  OR U20334 ( .A(n20016), .B(n20017), .Z(n20015) );
  NAND U20335 ( .A(n20017), .B(n20016), .Z(n20012) );
  ANDN U20336 ( .B(B[145]), .A(n38), .Z(n19807) );
  XNOR U20337 ( .A(n19815), .B(n20018), .Z(n19808) );
  XNOR U20338 ( .A(n19814), .B(n19812), .Z(n20018) );
  AND U20339 ( .A(n20019), .B(n20020), .Z(n19812) );
  NANDN U20340 ( .A(n20021), .B(n20022), .Z(n20020) );
  NANDN U20341 ( .A(n20023), .B(n20024), .Z(n20022) );
  NANDN U20342 ( .A(n20024), .B(n20023), .Z(n20019) );
  ANDN U20343 ( .B(B[146]), .A(n39), .Z(n19814) );
  XNOR U20344 ( .A(n19822), .B(n20025), .Z(n19815) );
  XNOR U20345 ( .A(n19821), .B(n19819), .Z(n20025) );
  AND U20346 ( .A(n20026), .B(n20027), .Z(n19819) );
  NANDN U20347 ( .A(n20028), .B(n20029), .Z(n20027) );
  OR U20348 ( .A(n20030), .B(n20031), .Z(n20029) );
  NAND U20349 ( .A(n20031), .B(n20030), .Z(n20026) );
  ANDN U20350 ( .B(B[147]), .A(n40), .Z(n19821) );
  XNOR U20351 ( .A(n19829), .B(n20032), .Z(n19822) );
  XNOR U20352 ( .A(n19828), .B(n19826), .Z(n20032) );
  AND U20353 ( .A(n20033), .B(n20034), .Z(n19826) );
  NANDN U20354 ( .A(n20035), .B(n20036), .Z(n20034) );
  NAND U20355 ( .A(n20037), .B(n20038), .Z(n20036) );
  ANDN U20356 ( .B(B[148]), .A(n41), .Z(n19828) );
  XOR U20357 ( .A(n19835), .B(n20039), .Z(n19829) );
  XNOR U20358 ( .A(n19833), .B(n19836), .Z(n20039) );
  NAND U20359 ( .A(A[2]), .B(B[149]), .Z(n19836) );
  NANDN U20360 ( .A(n20040), .B(n20041), .Z(n19833) );
  AND U20361 ( .A(A[0]), .B(B[150]), .Z(n20041) );
  XNOR U20362 ( .A(n19838), .B(n20042), .Z(n19835) );
  NAND U20363 ( .A(A[0]), .B(B[151]), .Z(n20042) );
  NAND U20364 ( .A(B[150]), .B(A[1]), .Z(n19838) );
  NAND U20365 ( .A(n20043), .B(n20044), .Z(n453) );
  NANDN U20366 ( .A(n20045), .B(n20046), .Z(n20044) );
  OR U20367 ( .A(n20047), .B(n20048), .Z(n20046) );
  NAND U20368 ( .A(n20048), .B(n20047), .Z(n20043) );
  XOR U20369 ( .A(n455), .B(n454), .Z(\A1[148] ) );
  XOR U20370 ( .A(n20048), .B(n20049), .Z(n454) );
  XNOR U20371 ( .A(n20047), .B(n20045), .Z(n20049) );
  AND U20372 ( .A(n20050), .B(n20051), .Z(n20045) );
  NANDN U20373 ( .A(n20052), .B(n20053), .Z(n20051) );
  NANDN U20374 ( .A(n20054), .B(n20055), .Z(n20053) );
  NANDN U20375 ( .A(n20055), .B(n20054), .Z(n20050) );
  ANDN U20376 ( .B(B[135]), .A(n29), .Z(n20047) );
  XNOR U20377 ( .A(n19954), .B(n20056), .Z(n20048) );
  XNOR U20378 ( .A(n19953), .B(n19951), .Z(n20056) );
  AND U20379 ( .A(n20057), .B(n20058), .Z(n19951) );
  NANDN U20380 ( .A(n20059), .B(n20060), .Z(n20058) );
  OR U20381 ( .A(n20061), .B(n20062), .Z(n20060) );
  NAND U20382 ( .A(n20062), .B(n20061), .Z(n20057) );
  ANDN U20383 ( .B(B[136]), .A(n30), .Z(n19953) );
  XNOR U20384 ( .A(n19961), .B(n20063), .Z(n19954) );
  XNOR U20385 ( .A(n19960), .B(n19958), .Z(n20063) );
  AND U20386 ( .A(n20064), .B(n20065), .Z(n19958) );
  NANDN U20387 ( .A(n20066), .B(n20067), .Z(n20065) );
  NANDN U20388 ( .A(n20068), .B(n20069), .Z(n20067) );
  NANDN U20389 ( .A(n20069), .B(n20068), .Z(n20064) );
  ANDN U20390 ( .B(B[137]), .A(n31), .Z(n19960) );
  XNOR U20391 ( .A(n19968), .B(n20070), .Z(n19961) );
  XNOR U20392 ( .A(n19967), .B(n19965), .Z(n20070) );
  AND U20393 ( .A(n20071), .B(n20072), .Z(n19965) );
  NANDN U20394 ( .A(n20073), .B(n20074), .Z(n20072) );
  OR U20395 ( .A(n20075), .B(n20076), .Z(n20074) );
  NAND U20396 ( .A(n20076), .B(n20075), .Z(n20071) );
  ANDN U20397 ( .B(B[138]), .A(n32), .Z(n19967) );
  XNOR U20398 ( .A(n19975), .B(n20077), .Z(n19968) );
  XNOR U20399 ( .A(n19974), .B(n19972), .Z(n20077) );
  AND U20400 ( .A(n20078), .B(n20079), .Z(n19972) );
  NANDN U20401 ( .A(n20080), .B(n20081), .Z(n20079) );
  NANDN U20402 ( .A(n20082), .B(n20083), .Z(n20081) );
  NANDN U20403 ( .A(n20083), .B(n20082), .Z(n20078) );
  ANDN U20404 ( .B(B[139]), .A(n33), .Z(n19974) );
  XNOR U20405 ( .A(n19982), .B(n20084), .Z(n19975) );
  XNOR U20406 ( .A(n19981), .B(n19979), .Z(n20084) );
  AND U20407 ( .A(n20085), .B(n20086), .Z(n19979) );
  NANDN U20408 ( .A(n20087), .B(n20088), .Z(n20086) );
  OR U20409 ( .A(n20089), .B(n20090), .Z(n20088) );
  NAND U20410 ( .A(n20090), .B(n20089), .Z(n20085) );
  ANDN U20411 ( .B(B[140]), .A(n34), .Z(n19981) );
  XNOR U20412 ( .A(n19989), .B(n20091), .Z(n19982) );
  XNOR U20413 ( .A(n19988), .B(n19986), .Z(n20091) );
  AND U20414 ( .A(n20092), .B(n20093), .Z(n19986) );
  NANDN U20415 ( .A(n20094), .B(n20095), .Z(n20093) );
  NANDN U20416 ( .A(n20096), .B(n20097), .Z(n20095) );
  NANDN U20417 ( .A(n20097), .B(n20096), .Z(n20092) );
  ANDN U20418 ( .B(B[141]), .A(n35), .Z(n19988) );
  XNOR U20419 ( .A(n19996), .B(n20098), .Z(n19989) );
  XNOR U20420 ( .A(n19995), .B(n19993), .Z(n20098) );
  AND U20421 ( .A(n20099), .B(n20100), .Z(n19993) );
  NANDN U20422 ( .A(n20101), .B(n20102), .Z(n20100) );
  OR U20423 ( .A(n20103), .B(n20104), .Z(n20102) );
  NAND U20424 ( .A(n20104), .B(n20103), .Z(n20099) );
  ANDN U20425 ( .B(B[142]), .A(n36), .Z(n19995) );
  XNOR U20426 ( .A(n20003), .B(n20105), .Z(n19996) );
  XNOR U20427 ( .A(n20002), .B(n20000), .Z(n20105) );
  AND U20428 ( .A(n20106), .B(n20107), .Z(n20000) );
  NANDN U20429 ( .A(n20108), .B(n20109), .Z(n20107) );
  NANDN U20430 ( .A(n20110), .B(n20111), .Z(n20109) );
  NANDN U20431 ( .A(n20111), .B(n20110), .Z(n20106) );
  ANDN U20432 ( .B(B[143]), .A(n37), .Z(n20002) );
  XNOR U20433 ( .A(n20010), .B(n20112), .Z(n20003) );
  XNOR U20434 ( .A(n20009), .B(n20007), .Z(n20112) );
  AND U20435 ( .A(n20113), .B(n20114), .Z(n20007) );
  NANDN U20436 ( .A(n20115), .B(n20116), .Z(n20114) );
  OR U20437 ( .A(n20117), .B(n20118), .Z(n20116) );
  NAND U20438 ( .A(n20118), .B(n20117), .Z(n20113) );
  ANDN U20439 ( .B(B[144]), .A(n38), .Z(n20009) );
  XNOR U20440 ( .A(n20017), .B(n20119), .Z(n20010) );
  XNOR U20441 ( .A(n20016), .B(n20014), .Z(n20119) );
  AND U20442 ( .A(n20120), .B(n20121), .Z(n20014) );
  NANDN U20443 ( .A(n20122), .B(n20123), .Z(n20121) );
  NANDN U20444 ( .A(n20124), .B(n20125), .Z(n20123) );
  NANDN U20445 ( .A(n20125), .B(n20124), .Z(n20120) );
  ANDN U20446 ( .B(B[145]), .A(n39), .Z(n20016) );
  XNOR U20447 ( .A(n20024), .B(n20126), .Z(n20017) );
  XNOR U20448 ( .A(n20023), .B(n20021), .Z(n20126) );
  AND U20449 ( .A(n20127), .B(n20128), .Z(n20021) );
  NANDN U20450 ( .A(n20129), .B(n20130), .Z(n20128) );
  OR U20451 ( .A(n20131), .B(n20132), .Z(n20130) );
  NAND U20452 ( .A(n20132), .B(n20131), .Z(n20127) );
  ANDN U20453 ( .B(B[146]), .A(n40), .Z(n20023) );
  XNOR U20454 ( .A(n20031), .B(n20133), .Z(n20024) );
  XNOR U20455 ( .A(n20030), .B(n20028), .Z(n20133) );
  AND U20456 ( .A(n20134), .B(n20135), .Z(n20028) );
  NANDN U20457 ( .A(n20136), .B(n20137), .Z(n20135) );
  NAND U20458 ( .A(n20138), .B(n20139), .Z(n20137) );
  ANDN U20459 ( .B(B[147]), .A(n41), .Z(n20030) );
  XOR U20460 ( .A(n20037), .B(n20140), .Z(n20031) );
  XNOR U20461 ( .A(n20035), .B(n20038), .Z(n20140) );
  NAND U20462 ( .A(A[2]), .B(B[148]), .Z(n20038) );
  NANDN U20463 ( .A(n20141), .B(n20142), .Z(n20035) );
  AND U20464 ( .A(A[0]), .B(B[149]), .Z(n20142) );
  XNOR U20465 ( .A(n20040), .B(n20143), .Z(n20037) );
  NAND U20466 ( .A(A[0]), .B(B[150]), .Z(n20143) );
  NAND U20467 ( .A(B[149]), .B(A[1]), .Z(n20040) );
  NAND U20468 ( .A(n20144), .B(n20145), .Z(n455) );
  NANDN U20469 ( .A(n20146), .B(n20147), .Z(n20145) );
  OR U20470 ( .A(n20148), .B(n20149), .Z(n20147) );
  NAND U20471 ( .A(n20149), .B(n20148), .Z(n20144) );
  XOR U20472 ( .A(n457), .B(n456), .Z(\A1[147] ) );
  XOR U20473 ( .A(n20149), .B(n20150), .Z(n456) );
  XNOR U20474 ( .A(n20148), .B(n20146), .Z(n20150) );
  AND U20475 ( .A(n20151), .B(n20152), .Z(n20146) );
  NANDN U20476 ( .A(n20153), .B(n20154), .Z(n20152) );
  NANDN U20477 ( .A(n20155), .B(n20156), .Z(n20154) );
  NANDN U20478 ( .A(n20156), .B(n20155), .Z(n20151) );
  ANDN U20479 ( .B(B[134]), .A(n29), .Z(n20148) );
  XNOR U20480 ( .A(n20055), .B(n20157), .Z(n20149) );
  XNOR U20481 ( .A(n20054), .B(n20052), .Z(n20157) );
  AND U20482 ( .A(n20158), .B(n20159), .Z(n20052) );
  NANDN U20483 ( .A(n20160), .B(n20161), .Z(n20159) );
  OR U20484 ( .A(n20162), .B(n20163), .Z(n20161) );
  NAND U20485 ( .A(n20163), .B(n20162), .Z(n20158) );
  ANDN U20486 ( .B(B[135]), .A(n30), .Z(n20054) );
  XNOR U20487 ( .A(n20062), .B(n20164), .Z(n20055) );
  XNOR U20488 ( .A(n20061), .B(n20059), .Z(n20164) );
  AND U20489 ( .A(n20165), .B(n20166), .Z(n20059) );
  NANDN U20490 ( .A(n20167), .B(n20168), .Z(n20166) );
  NANDN U20491 ( .A(n20169), .B(n20170), .Z(n20168) );
  NANDN U20492 ( .A(n20170), .B(n20169), .Z(n20165) );
  ANDN U20493 ( .B(B[136]), .A(n31), .Z(n20061) );
  XNOR U20494 ( .A(n20069), .B(n20171), .Z(n20062) );
  XNOR U20495 ( .A(n20068), .B(n20066), .Z(n20171) );
  AND U20496 ( .A(n20172), .B(n20173), .Z(n20066) );
  NANDN U20497 ( .A(n20174), .B(n20175), .Z(n20173) );
  OR U20498 ( .A(n20176), .B(n20177), .Z(n20175) );
  NAND U20499 ( .A(n20177), .B(n20176), .Z(n20172) );
  ANDN U20500 ( .B(B[137]), .A(n32), .Z(n20068) );
  XNOR U20501 ( .A(n20076), .B(n20178), .Z(n20069) );
  XNOR U20502 ( .A(n20075), .B(n20073), .Z(n20178) );
  AND U20503 ( .A(n20179), .B(n20180), .Z(n20073) );
  NANDN U20504 ( .A(n20181), .B(n20182), .Z(n20180) );
  NANDN U20505 ( .A(n20183), .B(n20184), .Z(n20182) );
  NANDN U20506 ( .A(n20184), .B(n20183), .Z(n20179) );
  ANDN U20507 ( .B(B[138]), .A(n33), .Z(n20075) );
  XNOR U20508 ( .A(n20083), .B(n20185), .Z(n20076) );
  XNOR U20509 ( .A(n20082), .B(n20080), .Z(n20185) );
  AND U20510 ( .A(n20186), .B(n20187), .Z(n20080) );
  NANDN U20511 ( .A(n20188), .B(n20189), .Z(n20187) );
  OR U20512 ( .A(n20190), .B(n20191), .Z(n20189) );
  NAND U20513 ( .A(n20191), .B(n20190), .Z(n20186) );
  ANDN U20514 ( .B(B[139]), .A(n34), .Z(n20082) );
  XNOR U20515 ( .A(n20090), .B(n20192), .Z(n20083) );
  XNOR U20516 ( .A(n20089), .B(n20087), .Z(n20192) );
  AND U20517 ( .A(n20193), .B(n20194), .Z(n20087) );
  NANDN U20518 ( .A(n20195), .B(n20196), .Z(n20194) );
  NANDN U20519 ( .A(n20197), .B(n20198), .Z(n20196) );
  NANDN U20520 ( .A(n20198), .B(n20197), .Z(n20193) );
  ANDN U20521 ( .B(B[140]), .A(n35), .Z(n20089) );
  XNOR U20522 ( .A(n20097), .B(n20199), .Z(n20090) );
  XNOR U20523 ( .A(n20096), .B(n20094), .Z(n20199) );
  AND U20524 ( .A(n20200), .B(n20201), .Z(n20094) );
  NANDN U20525 ( .A(n20202), .B(n20203), .Z(n20201) );
  OR U20526 ( .A(n20204), .B(n20205), .Z(n20203) );
  NAND U20527 ( .A(n20205), .B(n20204), .Z(n20200) );
  ANDN U20528 ( .B(B[141]), .A(n36), .Z(n20096) );
  XNOR U20529 ( .A(n20104), .B(n20206), .Z(n20097) );
  XNOR U20530 ( .A(n20103), .B(n20101), .Z(n20206) );
  AND U20531 ( .A(n20207), .B(n20208), .Z(n20101) );
  NANDN U20532 ( .A(n20209), .B(n20210), .Z(n20208) );
  NANDN U20533 ( .A(n20211), .B(n20212), .Z(n20210) );
  NANDN U20534 ( .A(n20212), .B(n20211), .Z(n20207) );
  ANDN U20535 ( .B(B[142]), .A(n37), .Z(n20103) );
  XNOR U20536 ( .A(n20111), .B(n20213), .Z(n20104) );
  XNOR U20537 ( .A(n20110), .B(n20108), .Z(n20213) );
  AND U20538 ( .A(n20214), .B(n20215), .Z(n20108) );
  NANDN U20539 ( .A(n20216), .B(n20217), .Z(n20215) );
  OR U20540 ( .A(n20218), .B(n20219), .Z(n20217) );
  NAND U20541 ( .A(n20219), .B(n20218), .Z(n20214) );
  ANDN U20542 ( .B(B[143]), .A(n38), .Z(n20110) );
  XNOR U20543 ( .A(n20118), .B(n20220), .Z(n20111) );
  XNOR U20544 ( .A(n20117), .B(n20115), .Z(n20220) );
  AND U20545 ( .A(n20221), .B(n20222), .Z(n20115) );
  NANDN U20546 ( .A(n20223), .B(n20224), .Z(n20222) );
  NANDN U20547 ( .A(n20225), .B(n20226), .Z(n20224) );
  NANDN U20548 ( .A(n20226), .B(n20225), .Z(n20221) );
  ANDN U20549 ( .B(B[144]), .A(n39), .Z(n20117) );
  XNOR U20550 ( .A(n20125), .B(n20227), .Z(n20118) );
  XNOR U20551 ( .A(n20124), .B(n20122), .Z(n20227) );
  AND U20552 ( .A(n20228), .B(n20229), .Z(n20122) );
  NANDN U20553 ( .A(n20230), .B(n20231), .Z(n20229) );
  OR U20554 ( .A(n20232), .B(n20233), .Z(n20231) );
  NAND U20555 ( .A(n20233), .B(n20232), .Z(n20228) );
  ANDN U20556 ( .B(B[145]), .A(n40), .Z(n20124) );
  XNOR U20557 ( .A(n20132), .B(n20234), .Z(n20125) );
  XNOR U20558 ( .A(n20131), .B(n20129), .Z(n20234) );
  AND U20559 ( .A(n20235), .B(n20236), .Z(n20129) );
  NANDN U20560 ( .A(n20237), .B(n20238), .Z(n20236) );
  NAND U20561 ( .A(n20239), .B(n20240), .Z(n20238) );
  ANDN U20562 ( .B(B[146]), .A(n41), .Z(n20131) );
  XOR U20563 ( .A(n20138), .B(n20241), .Z(n20132) );
  XNOR U20564 ( .A(n20136), .B(n20139), .Z(n20241) );
  NAND U20565 ( .A(A[2]), .B(B[147]), .Z(n20139) );
  NANDN U20566 ( .A(n20242), .B(n20243), .Z(n20136) );
  AND U20567 ( .A(A[0]), .B(B[148]), .Z(n20243) );
  XNOR U20568 ( .A(n20141), .B(n20244), .Z(n20138) );
  NAND U20569 ( .A(A[0]), .B(B[149]), .Z(n20244) );
  NAND U20570 ( .A(B[148]), .B(A[1]), .Z(n20141) );
  NAND U20571 ( .A(n20245), .B(n20246), .Z(n457) );
  NANDN U20572 ( .A(n20247), .B(n20248), .Z(n20246) );
  OR U20573 ( .A(n20249), .B(n20250), .Z(n20248) );
  NAND U20574 ( .A(n20250), .B(n20249), .Z(n20245) );
  XOR U20575 ( .A(n459), .B(n458), .Z(\A1[146] ) );
  XOR U20576 ( .A(n20250), .B(n20251), .Z(n458) );
  XNOR U20577 ( .A(n20249), .B(n20247), .Z(n20251) );
  AND U20578 ( .A(n20252), .B(n20253), .Z(n20247) );
  NANDN U20579 ( .A(n20254), .B(n20255), .Z(n20253) );
  NANDN U20580 ( .A(n20256), .B(n20257), .Z(n20255) );
  NANDN U20581 ( .A(n20257), .B(n20256), .Z(n20252) );
  ANDN U20582 ( .B(B[133]), .A(n29), .Z(n20249) );
  XNOR U20583 ( .A(n20156), .B(n20258), .Z(n20250) );
  XNOR U20584 ( .A(n20155), .B(n20153), .Z(n20258) );
  AND U20585 ( .A(n20259), .B(n20260), .Z(n20153) );
  NANDN U20586 ( .A(n20261), .B(n20262), .Z(n20260) );
  OR U20587 ( .A(n20263), .B(n20264), .Z(n20262) );
  NAND U20588 ( .A(n20264), .B(n20263), .Z(n20259) );
  ANDN U20589 ( .B(B[134]), .A(n30), .Z(n20155) );
  XNOR U20590 ( .A(n20163), .B(n20265), .Z(n20156) );
  XNOR U20591 ( .A(n20162), .B(n20160), .Z(n20265) );
  AND U20592 ( .A(n20266), .B(n20267), .Z(n20160) );
  NANDN U20593 ( .A(n20268), .B(n20269), .Z(n20267) );
  NANDN U20594 ( .A(n20270), .B(n20271), .Z(n20269) );
  NANDN U20595 ( .A(n20271), .B(n20270), .Z(n20266) );
  ANDN U20596 ( .B(B[135]), .A(n31), .Z(n20162) );
  XNOR U20597 ( .A(n20170), .B(n20272), .Z(n20163) );
  XNOR U20598 ( .A(n20169), .B(n20167), .Z(n20272) );
  AND U20599 ( .A(n20273), .B(n20274), .Z(n20167) );
  NANDN U20600 ( .A(n20275), .B(n20276), .Z(n20274) );
  OR U20601 ( .A(n20277), .B(n20278), .Z(n20276) );
  NAND U20602 ( .A(n20278), .B(n20277), .Z(n20273) );
  ANDN U20603 ( .B(B[136]), .A(n32), .Z(n20169) );
  XNOR U20604 ( .A(n20177), .B(n20279), .Z(n20170) );
  XNOR U20605 ( .A(n20176), .B(n20174), .Z(n20279) );
  AND U20606 ( .A(n20280), .B(n20281), .Z(n20174) );
  NANDN U20607 ( .A(n20282), .B(n20283), .Z(n20281) );
  NANDN U20608 ( .A(n20284), .B(n20285), .Z(n20283) );
  NANDN U20609 ( .A(n20285), .B(n20284), .Z(n20280) );
  ANDN U20610 ( .B(B[137]), .A(n33), .Z(n20176) );
  XNOR U20611 ( .A(n20184), .B(n20286), .Z(n20177) );
  XNOR U20612 ( .A(n20183), .B(n20181), .Z(n20286) );
  AND U20613 ( .A(n20287), .B(n20288), .Z(n20181) );
  NANDN U20614 ( .A(n20289), .B(n20290), .Z(n20288) );
  OR U20615 ( .A(n20291), .B(n20292), .Z(n20290) );
  NAND U20616 ( .A(n20292), .B(n20291), .Z(n20287) );
  ANDN U20617 ( .B(B[138]), .A(n34), .Z(n20183) );
  XNOR U20618 ( .A(n20191), .B(n20293), .Z(n20184) );
  XNOR U20619 ( .A(n20190), .B(n20188), .Z(n20293) );
  AND U20620 ( .A(n20294), .B(n20295), .Z(n20188) );
  NANDN U20621 ( .A(n20296), .B(n20297), .Z(n20295) );
  NANDN U20622 ( .A(n20298), .B(n20299), .Z(n20297) );
  NANDN U20623 ( .A(n20299), .B(n20298), .Z(n20294) );
  ANDN U20624 ( .B(B[139]), .A(n35), .Z(n20190) );
  XNOR U20625 ( .A(n20198), .B(n20300), .Z(n20191) );
  XNOR U20626 ( .A(n20197), .B(n20195), .Z(n20300) );
  AND U20627 ( .A(n20301), .B(n20302), .Z(n20195) );
  NANDN U20628 ( .A(n20303), .B(n20304), .Z(n20302) );
  OR U20629 ( .A(n20305), .B(n20306), .Z(n20304) );
  NAND U20630 ( .A(n20306), .B(n20305), .Z(n20301) );
  ANDN U20631 ( .B(B[140]), .A(n36), .Z(n20197) );
  XNOR U20632 ( .A(n20205), .B(n20307), .Z(n20198) );
  XNOR U20633 ( .A(n20204), .B(n20202), .Z(n20307) );
  AND U20634 ( .A(n20308), .B(n20309), .Z(n20202) );
  NANDN U20635 ( .A(n20310), .B(n20311), .Z(n20309) );
  NANDN U20636 ( .A(n20312), .B(n20313), .Z(n20311) );
  NANDN U20637 ( .A(n20313), .B(n20312), .Z(n20308) );
  ANDN U20638 ( .B(B[141]), .A(n37), .Z(n20204) );
  XNOR U20639 ( .A(n20212), .B(n20314), .Z(n20205) );
  XNOR U20640 ( .A(n20211), .B(n20209), .Z(n20314) );
  AND U20641 ( .A(n20315), .B(n20316), .Z(n20209) );
  NANDN U20642 ( .A(n20317), .B(n20318), .Z(n20316) );
  OR U20643 ( .A(n20319), .B(n20320), .Z(n20318) );
  NAND U20644 ( .A(n20320), .B(n20319), .Z(n20315) );
  ANDN U20645 ( .B(B[142]), .A(n38), .Z(n20211) );
  XNOR U20646 ( .A(n20219), .B(n20321), .Z(n20212) );
  XNOR U20647 ( .A(n20218), .B(n20216), .Z(n20321) );
  AND U20648 ( .A(n20322), .B(n20323), .Z(n20216) );
  NANDN U20649 ( .A(n20324), .B(n20325), .Z(n20323) );
  NANDN U20650 ( .A(n20326), .B(n20327), .Z(n20325) );
  NANDN U20651 ( .A(n20327), .B(n20326), .Z(n20322) );
  ANDN U20652 ( .B(B[143]), .A(n39), .Z(n20218) );
  XNOR U20653 ( .A(n20226), .B(n20328), .Z(n20219) );
  XNOR U20654 ( .A(n20225), .B(n20223), .Z(n20328) );
  AND U20655 ( .A(n20329), .B(n20330), .Z(n20223) );
  NANDN U20656 ( .A(n20331), .B(n20332), .Z(n20330) );
  OR U20657 ( .A(n20333), .B(n20334), .Z(n20332) );
  NAND U20658 ( .A(n20334), .B(n20333), .Z(n20329) );
  ANDN U20659 ( .B(B[144]), .A(n40), .Z(n20225) );
  XNOR U20660 ( .A(n20233), .B(n20335), .Z(n20226) );
  XNOR U20661 ( .A(n20232), .B(n20230), .Z(n20335) );
  AND U20662 ( .A(n20336), .B(n20337), .Z(n20230) );
  NANDN U20663 ( .A(n20338), .B(n20339), .Z(n20337) );
  NAND U20664 ( .A(n20340), .B(n20341), .Z(n20339) );
  ANDN U20665 ( .B(B[145]), .A(n41), .Z(n20232) );
  XOR U20666 ( .A(n20239), .B(n20342), .Z(n20233) );
  XNOR U20667 ( .A(n20237), .B(n20240), .Z(n20342) );
  NAND U20668 ( .A(A[2]), .B(B[146]), .Z(n20240) );
  NANDN U20669 ( .A(n20343), .B(n20344), .Z(n20237) );
  AND U20670 ( .A(A[0]), .B(B[147]), .Z(n20344) );
  XNOR U20671 ( .A(n20242), .B(n20345), .Z(n20239) );
  NAND U20672 ( .A(A[0]), .B(B[148]), .Z(n20345) );
  NAND U20673 ( .A(B[147]), .B(A[1]), .Z(n20242) );
  NAND U20674 ( .A(n20346), .B(n20347), .Z(n459) );
  NANDN U20675 ( .A(n20348), .B(n20349), .Z(n20347) );
  OR U20676 ( .A(n20350), .B(n20351), .Z(n20349) );
  NAND U20677 ( .A(n20351), .B(n20350), .Z(n20346) );
  XOR U20678 ( .A(n461), .B(n460), .Z(\A1[145] ) );
  XOR U20679 ( .A(n20351), .B(n20352), .Z(n460) );
  XNOR U20680 ( .A(n20350), .B(n20348), .Z(n20352) );
  AND U20681 ( .A(n20353), .B(n20354), .Z(n20348) );
  NANDN U20682 ( .A(n20355), .B(n20356), .Z(n20354) );
  NANDN U20683 ( .A(n20357), .B(n20358), .Z(n20356) );
  NANDN U20684 ( .A(n20358), .B(n20357), .Z(n20353) );
  ANDN U20685 ( .B(B[132]), .A(n29), .Z(n20350) );
  XNOR U20686 ( .A(n20257), .B(n20359), .Z(n20351) );
  XNOR U20687 ( .A(n20256), .B(n20254), .Z(n20359) );
  AND U20688 ( .A(n20360), .B(n20361), .Z(n20254) );
  NANDN U20689 ( .A(n20362), .B(n20363), .Z(n20361) );
  OR U20690 ( .A(n20364), .B(n20365), .Z(n20363) );
  NAND U20691 ( .A(n20365), .B(n20364), .Z(n20360) );
  ANDN U20692 ( .B(B[133]), .A(n30), .Z(n20256) );
  XNOR U20693 ( .A(n20264), .B(n20366), .Z(n20257) );
  XNOR U20694 ( .A(n20263), .B(n20261), .Z(n20366) );
  AND U20695 ( .A(n20367), .B(n20368), .Z(n20261) );
  NANDN U20696 ( .A(n20369), .B(n20370), .Z(n20368) );
  NANDN U20697 ( .A(n20371), .B(n20372), .Z(n20370) );
  NANDN U20698 ( .A(n20372), .B(n20371), .Z(n20367) );
  ANDN U20699 ( .B(B[134]), .A(n31), .Z(n20263) );
  XNOR U20700 ( .A(n20271), .B(n20373), .Z(n20264) );
  XNOR U20701 ( .A(n20270), .B(n20268), .Z(n20373) );
  AND U20702 ( .A(n20374), .B(n20375), .Z(n20268) );
  NANDN U20703 ( .A(n20376), .B(n20377), .Z(n20375) );
  OR U20704 ( .A(n20378), .B(n20379), .Z(n20377) );
  NAND U20705 ( .A(n20379), .B(n20378), .Z(n20374) );
  ANDN U20706 ( .B(B[135]), .A(n32), .Z(n20270) );
  XNOR U20707 ( .A(n20278), .B(n20380), .Z(n20271) );
  XNOR U20708 ( .A(n20277), .B(n20275), .Z(n20380) );
  AND U20709 ( .A(n20381), .B(n20382), .Z(n20275) );
  NANDN U20710 ( .A(n20383), .B(n20384), .Z(n20382) );
  NANDN U20711 ( .A(n20385), .B(n20386), .Z(n20384) );
  NANDN U20712 ( .A(n20386), .B(n20385), .Z(n20381) );
  ANDN U20713 ( .B(B[136]), .A(n33), .Z(n20277) );
  XNOR U20714 ( .A(n20285), .B(n20387), .Z(n20278) );
  XNOR U20715 ( .A(n20284), .B(n20282), .Z(n20387) );
  AND U20716 ( .A(n20388), .B(n20389), .Z(n20282) );
  NANDN U20717 ( .A(n20390), .B(n20391), .Z(n20389) );
  OR U20718 ( .A(n20392), .B(n20393), .Z(n20391) );
  NAND U20719 ( .A(n20393), .B(n20392), .Z(n20388) );
  ANDN U20720 ( .B(B[137]), .A(n34), .Z(n20284) );
  XNOR U20721 ( .A(n20292), .B(n20394), .Z(n20285) );
  XNOR U20722 ( .A(n20291), .B(n20289), .Z(n20394) );
  AND U20723 ( .A(n20395), .B(n20396), .Z(n20289) );
  NANDN U20724 ( .A(n20397), .B(n20398), .Z(n20396) );
  NANDN U20725 ( .A(n20399), .B(n20400), .Z(n20398) );
  NANDN U20726 ( .A(n20400), .B(n20399), .Z(n20395) );
  ANDN U20727 ( .B(B[138]), .A(n35), .Z(n20291) );
  XNOR U20728 ( .A(n20299), .B(n20401), .Z(n20292) );
  XNOR U20729 ( .A(n20298), .B(n20296), .Z(n20401) );
  AND U20730 ( .A(n20402), .B(n20403), .Z(n20296) );
  NANDN U20731 ( .A(n20404), .B(n20405), .Z(n20403) );
  OR U20732 ( .A(n20406), .B(n20407), .Z(n20405) );
  NAND U20733 ( .A(n20407), .B(n20406), .Z(n20402) );
  ANDN U20734 ( .B(B[139]), .A(n36), .Z(n20298) );
  XNOR U20735 ( .A(n20306), .B(n20408), .Z(n20299) );
  XNOR U20736 ( .A(n20305), .B(n20303), .Z(n20408) );
  AND U20737 ( .A(n20409), .B(n20410), .Z(n20303) );
  NANDN U20738 ( .A(n20411), .B(n20412), .Z(n20410) );
  NANDN U20739 ( .A(n20413), .B(n20414), .Z(n20412) );
  NANDN U20740 ( .A(n20414), .B(n20413), .Z(n20409) );
  ANDN U20741 ( .B(B[140]), .A(n37), .Z(n20305) );
  XNOR U20742 ( .A(n20313), .B(n20415), .Z(n20306) );
  XNOR U20743 ( .A(n20312), .B(n20310), .Z(n20415) );
  AND U20744 ( .A(n20416), .B(n20417), .Z(n20310) );
  NANDN U20745 ( .A(n20418), .B(n20419), .Z(n20417) );
  OR U20746 ( .A(n20420), .B(n20421), .Z(n20419) );
  NAND U20747 ( .A(n20421), .B(n20420), .Z(n20416) );
  ANDN U20748 ( .B(B[141]), .A(n38), .Z(n20312) );
  XNOR U20749 ( .A(n20320), .B(n20422), .Z(n20313) );
  XNOR U20750 ( .A(n20319), .B(n20317), .Z(n20422) );
  AND U20751 ( .A(n20423), .B(n20424), .Z(n20317) );
  NANDN U20752 ( .A(n20425), .B(n20426), .Z(n20424) );
  NANDN U20753 ( .A(n20427), .B(n20428), .Z(n20426) );
  NANDN U20754 ( .A(n20428), .B(n20427), .Z(n20423) );
  ANDN U20755 ( .B(B[142]), .A(n39), .Z(n20319) );
  XNOR U20756 ( .A(n20327), .B(n20429), .Z(n20320) );
  XNOR U20757 ( .A(n20326), .B(n20324), .Z(n20429) );
  AND U20758 ( .A(n20430), .B(n20431), .Z(n20324) );
  NANDN U20759 ( .A(n20432), .B(n20433), .Z(n20431) );
  OR U20760 ( .A(n20434), .B(n20435), .Z(n20433) );
  NAND U20761 ( .A(n20435), .B(n20434), .Z(n20430) );
  ANDN U20762 ( .B(B[143]), .A(n40), .Z(n20326) );
  XNOR U20763 ( .A(n20334), .B(n20436), .Z(n20327) );
  XNOR U20764 ( .A(n20333), .B(n20331), .Z(n20436) );
  AND U20765 ( .A(n20437), .B(n20438), .Z(n20331) );
  NANDN U20766 ( .A(n20439), .B(n20440), .Z(n20438) );
  NAND U20767 ( .A(n20441), .B(n20442), .Z(n20440) );
  ANDN U20768 ( .B(B[144]), .A(n41), .Z(n20333) );
  XOR U20769 ( .A(n20340), .B(n20443), .Z(n20334) );
  XNOR U20770 ( .A(n20338), .B(n20341), .Z(n20443) );
  NAND U20771 ( .A(A[2]), .B(B[145]), .Z(n20341) );
  NANDN U20772 ( .A(n20444), .B(n20445), .Z(n20338) );
  AND U20773 ( .A(A[0]), .B(B[146]), .Z(n20445) );
  XNOR U20774 ( .A(n20343), .B(n20446), .Z(n20340) );
  NAND U20775 ( .A(A[0]), .B(B[147]), .Z(n20446) );
  NAND U20776 ( .A(B[146]), .B(A[1]), .Z(n20343) );
  NAND U20777 ( .A(n20447), .B(n20448), .Z(n461) );
  NANDN U20778 ( .A(n20449), .B(n20450), .Z(n20448) );
  OR U20779 ( .A(n20451), .B(n20452), .Z(n20450) );
  NAND U20780 ( .A(n20452), .B(n20451), .Z(n20447) );
  XOR U20781 ( .A(n463), .B(n462), .Z(\A1[144] ) );
  XOR U20782 ( .A(n20452), .B(n20453), .Z(n462) );
  XNOR U20783 ( .A(n20451), .B(n20449), .Z(n20453) );
  AND U20784 ( .A(n20454), .B(n20455), .Z(n20449) );
  NANDN U20785 ( .A(n20456), .B(n20457), .Z(n20455) );
  NANDN U20786 ( .A(n20458), .B(n20459), .Z(n20457) );
  NANDN U20787 ( .A(n20459), .B(n20458), .Z(n20454) );
  ANDN U20788 ( .B(B[131]), .A(n29), .Z(n20451) );
  XNOR U20789 ( .A(n20358), .B(n20460), .Z(n20452) );
  XNOR U20790 ( .A(n20357), .B(n20355), .Z(n20460) );
  AND U20791 ( .A(n20461), .B(n20462), .Z(n20355) );
  NANDN U20792 ( .A(n20463), .B(n20464), .Z(n20462) );
  OR U20793 ( .A(n20465), .B(n20466), .Z(n20464) );
  NAND U20794 ( .A(n20466), .B(n20465), .Z(n20461) );
  ANDN U20795 ( .B(B[132]), .A(n30), .Z(n20357) );
  XNOR U20796 ( .A(n20365), .B(n20467), .Z(n20358) );
  XNOR U20797 ( .A(n20364), .B(n20362), .Z(n20467) );
  AND U20798 ( .A(n20468), .B(n20469), .Z(n20362) );
  NANDN U20799 ( .A(n20470), .B(n20471), .Z(n20469) );
  NANDN U20800 ( .A(n20472), .B(n20473), .Z(n20471) );
  NANDN U20801 ( .A(n20473), .B(n20472), .Z(n20468) );
  ANDN U20802 ( .B(B[133]), .A(n31), .Z(n20364) );
  XNOR U20803 ( .A(n20372), .B(n20474), .Z(n20365) );
  XNOR U20804 ( .A(n20371), .B(n20369), .Z(n20474) );
  AND U20805 ( .A(n20475), .B(n20476), .Z(n20369) );
  NANDN U20806 ( .A(n20477), .B(n20478), .Z(n20476) );
  OR U20807 ( .A(n20479), .B(n20480), .Z(n20478) );
  NAND U20808 ( .A(n20480), .B(n20479), .Z(n20475) );
  ANDN U20809 ( .B(B[134]), .A(n32), .Z(n20371) );
  XNOR U20810 ( .A(n20379), .B(n20481), .Z(n20372) );
  XNOR U20811 ( .A(n20378), .B(n20376), .Z(n20481) );
  AND U20812 ( .A(n20482), .B(n20483), .Z(n20376) );
  NANDN U20813 ( .A(n20484), .B(n20485), .Z(n20483) );
  NANDN U20814 ( .A(n20486), .B(n20487), .Z(n20485) );
  NANDN U20815 ( .A(n20487), .B(n20486), .Z(n20482) );
  ANDN U20816 ( .B(B[135]), .A(n33), .Z(n20378) );
  XNOR U20817 ( .A(n20386), .B(n20488), .Z(n20379) );
  XNOR U20818 ( .A(n20385), .B(n20383), .Z(n20488) );
  AND U20819 ( .A(n20489), .B(n20490), .Z(n20383) );
  NANDN U20820 ( .A(n20491), .B(n20492), .Z(n20490) );
  OR U20821 ( .A(n20493), .B(n20494), .Z(n20492) );
  NAND U20822 ( .A(n20494), .B(n20493), .Z(n20489) );
  ANDN U20823 ( .B(B[136]), .A(n34), .Z(n20385) );
  XNOR U20824 ( .A(n20393), .B(n20495), .Z(n20386) );
  XNOR U20825 ( .A(n20392), .B(n20390), .Z(n20495) );
  AND U20826 ( .A(n20496), .B(n20497), .Z(n20390) );
  NANDN U20827 ( .A(n20498), .B(n20499), .Z(n20497) );
  NANDN U20828 ( .A(n20500), .B(n20501), .Z(n20499) );
  NANDN U20829 ( .A(n20501), .B(n20500), .Z(n20496) );
  ANDN U20830 ( .B(B[137]), .A(n35), .Z(n20392) );
  XNOR U20831 ( .A(n20400), .B(n20502), .Z(n20393) );
  XNOR U20832 ( .A(n20399), .B(n20397), .Z(n20502) );
  AND U20833 ( .A(n20503), .B(n20504), .Z(n20397) );
  NANDN U20834 ( .A(n20505), .B(n20506), .Z(n20504) );
  OR U20835 ( .A(n20507), .B(n20508), .Z(n20506) );
  NAND U20836 ( .A(n20508), .B(n20507), .Z(n20503) );
  ANDN U20837 ( .B(B[138]), .A(n36), .Z(n20399) );
  XNOR U20838 ( .A(n20407), .B(n20509), .Z(n20400) );
  XNOR U20839 ( .A(n20406), .B(n20404), .Z(n20509) );
  AND U20840 ( .A(n20510), .B(n20511), .Z(n20404) );
  NANDN U20841 ( .A(n20512), .B(n20513), .Z(n20511) );
  NANDN U20842 ( .A(n20514), .B(n20515), .Z(n20513) );
  NANDN U20843 ( .A(n20515), .B(n20514), .Z(n20510) );
  ANDN U20844 ( .B(B[139]), .A(n37), .Z(n20406) );
  XNOR U20845 ( .A(n20414), .B(n20516), .Z(n20407) );
  XNOR U20846 ( .A(n20413), .B(n20411), .Z(n20516) );
  AND U20847 ( .A(n20517), .B(n20518), .Z(n20411) );
  NANDN U20848 ( .A(n20519), .B(n20520), .Z(n20518) );
  OR U20849 ( .A(n20521), .B(n20522), .Z(n20520) );
  NAND U20850 ( .A(n20522), .B(n20521), .Z(n20517) );
  ANDN U20851 ( .B(B[140]), .A(n38), .Z(n20413) );
  XNOR U20852 ( .A(n20421), .B(n20523), .Z(n20414) );
  XNOR U20853 ( .A(n20420), .B(n20418), .Z(n20523) );
  AND U20854 ( .A(n20524), .B(n20525), .Z(n20418) );
  NANDN U20855 ( .A(n20526), .B(n20527), .Z(n20525) );
  NANDN U20856 ( .A(n20528), .B(n20529), .Z(n20527) );
  NANDN U20857 ( .A(n20529), .B(n20528), .Z(n20524) );
  ANDN U20858 ( .B(B[141]), .A(n39), .Z(n20420) );
  XNOR U20859 ( .A(n20428), .B(n20530), .Z(n20421) );
  XNOR U20860 ( .A(n20427), .B(n20425), .Z(n20530) );
  AND U20861 ( .A(n20531), .B(n20532), .Z(n20425) );
  NANDN U20862 ( .A(n20533), .B(n20534), .Z(n20532) );
  OR U20863 ( .A(n20535), .B(n20536), .Z(n20534) );
  NAND U20864 ( .A(n20536), .B(n20535), .Z(n20531) );
  ANDN U20865 ( .B(B[142]), .A(n40), .Z(n20427) );
  XNOR U20866 ( .A(n20435), .B(n20537), .Z(n20428) );
  XNOR U20867 ( .A(n20434), .B(n20432), .Z(n20537) );
  AND U20868 ( .A(n20538), .B(n20539), .Z(n20432) );
  NANDN U20869 ( .A(n20540), .B(n20541), .Z(n20539) );
  NAND U20870 ( .A(n20542), .B(n20543), .Z(n20541) );
  ANDN U20871 ( .B(B[143]), .A(n41), .Z(n20434) );
  XOR U20872 ( .A(n20441), .B(n20544), .Z(n20435) );
  XNOR U20873 ( .A(n20439), .B(n20442), .Z(n20544) );
  NAND U20874 ( .A(A[2]), .B(B[144]), .Z(n20442) );
  NANDN U20875 ( .A(n20545), .B(n20546), .Z(n20439) );
  AND U20876 ( .A(A[0]), .B(B[145]), .Z(n20546) );
  XNOR U20877 ( .A(n20444), .B(n20547), .Z(n20441) );
  NAND U20878 ( .A(A[0]), .B(B[146]), .Z(n20547) );
  NAND U20879 ( .A(B[145]), .B(A[1]), .Z(n20444) );
  NAND U20880 ( .A(n20548), .B(n20549), .Z(n463) );
  NANDN U20881 ( .A(n20550), .B(n20551), .Z(n20549) );
  OR U20882 ( .A(n20552), .B(n20553), .Z(n20551) );
  NAND U20883 ( .A(n20553), .B(n20552), .Z(n20548) );
  XOR U20884 ( .A(n465), .B(n464), .Z(\A1[143] ) );
  XOR U20885 ( .A(n20553), .B(n20554), .Z(n464) );
  XNOR U20886 ( .A(n20552), .B(n20550), .Z(n20554) );
  AND U20887 ( .A(n20555), .B(n20556), .Z(n20550) );
  NANDN U20888 ( .A(n20557), .B(n20558), .Z(n20556) );
  NANDN U20889 ( .A(n20559), .B(n20560), .Z(n20558) );
  NANDN U20890 ( .A(n20560), .B(n20559), .Z(n20555) );
  ANDN U20891 ( .B(B[130]), .A(n29), .Z(n20552) );
  XNOR U20892 ( .A(n20459), .B(n20561), .Z(n20553) );
  XNOR U20893 ( .A(n20458), .B(n20456), .Z(n20561) );
  AND U20894 ( .A(n20562), .B(n20563), .Z(n20456) );
  NANDN U20895 ( .A(n20564), .B(n20565), .Z(n20563) );
  OR U20896 ( .A(n20566), .B(n20567), .Z(n20565) );
  NAND U20897 ( .A(n20567), .B(n20566), .Z(n20562) );
  ANDN U20898 ( .B(B[131]), .A(n30), .Z(n20458) );
  XNOR U20899 ( .A(n20466), .B(n20568), .Z(n20459) );
  XNOR U20900 ( .A(n20465), .B(n20463), .Z(n20568) );
  AND U20901 ( .A(n20569), .B(n20570), .Z(n20463) );
  NANDN U20902 ( .A(n20571), .B(n20572), .Z(n20570) );
  NANDN U20903 ( .A(n20573), .B(n20574), .Z(n20572) );
  NANDN U20904 ( .A(n20574), .B(n20573), .Z(n20569) );
  ANDN U20905 ( .B(B[132]), .A(n31), .Z(n20465) );
  XNOR U20906 ( .A(n20473), .B(n20575), .Z(n20466) );
  XNOR U20907 ( .A(n20472), .B(n20470), .Z(n20575) );
  AND U20908 ( .A(n20576), .B(n20577), .Z(n20470) );
  NANDN U20909 ( .A(n20578), .B(n20579), .Z(n20577) );
  OR U20910 ( .A(n20580), .B(n20581), .Z(n20579) );
  NAND U20911 ( .A(n20581), .B(n20580), .Z(n20576) );
  ANDN U20912 ( .B(B[133]), .A(n32), .Z(n20472) );
  XNOR U20913 ( .A(n20480), .B(n20582), .Z(n20473) );
  XNOR U20914 ( .A(n20479), .B(n20477), .Z(n20582) );
  AND U20915 ( .A(n20583), .B(n20584), .Z(n20477) );
  NANDN U20916 ( .A(n20585), .B(n20586), .Z(n20584) );
  NANDN U20917 ( .A(n20587), .B(n20588), .Z(n20586) );
  NANDN U20918 ( .A(n20588), .B(n20587), .Z(n20583) );
  ANDN U20919 ( .B(B[134]), .A(n33), .Z(n20479) );
  XNOR U20920 ( .A(n20487), .B(n20589), .Z(n20480) );
  XNOR U20921 ( .A(n20486), .B(n20484), .Z(n20589) );
  AND U20922 ( .A(n20590), .B(n20591), .Z(n20484) );
  NANDN U20923 ( .A(n20592), .B(n20593), .Z(n20591) );
  OR U20924 ( .A(n20594), .B(n20595), .Z(n20593) );
  NAND U20925 ( .A(n20595), .B(n20594), .Z(n20590) );
  ANDN U20926 ( .B(B[135]), .A(n34), .Z(n20486) );
  XNOR U20927 ( .A(n20494), .B(n20596), .Z(n20487) );
  XNOR U20928 ( .A(n20493), .B(n20491), .Z(n20596) );
  AND U20929 ( .A(n20597), .B(n20598), .Z(n20491) );
  NANDN U20930 ( .A(n20599), .B(n20600), .Z(n20598) );
  NANDN U20931 ( .A(n20601), .B(n20602), .Z(n20600) );
  NANDN U20932 ( .A(n20602), .B(n20601), .Z(n20597) );
  ANDN U20933 ( .B(B[136]), .A(n35), .Z(n20493) );
  XNOR U20934 ( .A(n20501), .B(n20603), .Z(n20494) );
  XNOR U20935 ( .A(n20500), .B(n20498), .Z(n20603) );
  AND U20936 ( .A(n20604), .B(n20605), .Z(n20498) );
  NANDN U20937 ( .A(n20606), .B(n20607), .Z(n20605) );
  OR U20938 ( .A(n20608), .B(n20609), .Z(n20607) );
  NAND U20939 ( .A(n20609), .B(n20608), .Z(n20604) );
  ANDN U20940 ( .B(B[137]), .A(n36), .Z(n20500) );
  XNOR U20941 ( .A(n20508), .B(n20610), .Z(n20501) );
  XNOR U20942 ( .A(n20507), .B(n20505), .Z(n20610) );
  AND U20943 ( .A(n20611), .B(n20612), .Z(n20505) );
  NANDN U20944 ( .A(n20613), .B(n20614), .Z(n20612) );
  NANDN U20945 ( .A(n20615), .B(n20616), .Z(n20614) );
  NANDN U20946 ( .A(n20616), .B(n20615), .Z(n20611) );
  ANDN U20947 ( .B(B[138]), .A(n37), .Z(n20507) );
  XNOR U20948 ( .A(n20515), .B(n20617), .Z(n20508) );
  XNOR U20949 ( .A(n20514), .B(n20512), .Z(n20617) );
  AND U20950 ( .A(n20618), .B(n20619), .Z(n20512) );
  NANDN U20951 ( .A(n20620), .B(n20621), .Z(n20619) );
  OR U20952 ( .A(n20622), .B(n20623), .Z(n20621) );
  NAND U20953 ( .A(n20623), .B(n20622), .Z(n20618) );
  ANDN U20954 ( .B(B[139]), .A(n38), .Z(n20514) );
  XNOR U20955 ( .A(n20522), .B(n20624), .Z(n20515) );
  XNOR U20956 ( .A(n20521), .B(n20519), .Z(n20624) );
  AND U20957 ( .A(n20625), .B(n20626), .Z(n20519) );
  NANDN U20958 ( .A(n20627), .B(n20628), .Z(n20626) );
  NANDN U20959 ( .A(n20629), .B(n20630), .Z(n20628) );
  NANDN U20960 ( .A(n20630), .B(n20629), .Z(n20625) );
  ANDN U20961 ( .B(B[140]), .A(n39), .Z(n20521) );
  XNOR U20962 ( .A(n20529), .B(n20631), .Z(n20522) );
  XNOR U20963 ( .A(n20528), .B(n20526), .Z(n20631) );
  AND U20964 ( .A(n20632), .B(n20633), .Z(n20526) );
  NANDN U20965 ( .A(n20634), .B(n20635), .Z(n20633) );
  OR U20966 ( .A(n20636), .B(n20637), .Z(n20635) );
  NAND U20967 ( .A(n20637), .B(n20636), .Z(n20632) );
  ANDN U20968 ( .B(B[141]), .A(n40), .Z(n20528) );
  XNOR U20969 ( .A(n20536), .B(n20638), .Z(n20529) );
  XNOR U20970 ( .A(n20535), .B(n20533), .Z(n20638) );
  AND U20971 ( .A(n20639), .B(n20640), .Z(n20533) );
  NANDN U20972 ( .A(n20641), .B(n20642), .Z(n20640) );
  NAND U20973 ( .A(n20643), .B(n20644), .Z(n20642) );
  ANDN U20974 ( .B(B[142]), .A(n41), .Z(n20535) );
  XOR U20975 ( .A(n20542), .B(n20645), .Z(n20536) );
  XNOR U20976 ( .A(n20540), .B(n20543), .Z(n20645) );
  NAND U20977 ( .A(A[2]), .B(B[143]), .Z(n20543) );
  NANDN U20978 ( .A(n20646), .B(n20647), .Z(n20540) );
  AND U20979 ( .A(A[0]), .B(B[144]), .Z(n20647) );
  XNOR U20980 ( .A(n20545), .B(n20648), .Z(n20542) );
  NAND U20981 ( .A(A[0]), .B(B[145]), .Z(n20648) );
  NAND U20982 ( .A(B[144]), .B(A[1]), .Z(n20545) );
  NAND U20983 ( .A(n20649), .B(n20650), .Z(n465) );
  NANDN U20984 ( .A(n20651), .B(n20652), .Z(n20650) );
  OR U20985 ( .A(n20653), .B(n20654), .Z(n20652) );
  NAND U20986 ( .A(n20654), .B(n20653), .Z(n20649) );
  XOR U20987 ( .A(n467), .B(n466), .Z(\A1[142] ) );
  XOR U20988 ( .A(n20654), .B(n20655), .Z(n466) );
  XNOR U20989 ( .A(n20653), .B(n20651), .Z(n20655) );
  AND U20990 ( .A(n20656), .B(n20657), .Z(n20651) );
  NANDN U20991 ( .A(n20658), .B(n20659), .Z(n20657) );
  NANDN U20992 ( .A(n20660), .B(n20661), .Z(n20659) );
  NANDN U20993 ( .A(n20661), .B(n20660), .Z(n20656) );
  ANDN U20994 ( .B(B[129]), .A(n29), .Z(n20653) );
  XNOR U20995 ( .A(n20560), .B(n20662), .Z(n20654) );
  XNOR U20996 ( .A(n20559), .B(n20557), .Z(n20662) );
  AND U20997 ( .A(n20663), .B(n20664), .Z(n20557) );
  NANDN U20998 ( .A(n20665), .B(n20666), .Z(n20664) );
  OR U20999 ( .A(n20667), .B(n20668), .Z(n20666) );
  NAND U21000 ( .A(n20668), .B(n20667), .Z(n20663) );
  ANDN U21001 ( .B(B[130]), .A(n30), .Z(n20559) );
  XNOR U21002 ( .A(n20567), .B(n20669), .Z(n20560) );
  XNOR U21003 ( .A(n20566), .B(n20564), .Z(n20669) );
  AND U21004 ( .A(n20670), .B(n20671), .Z(n20564) );
  NANDN U21005 ( .A(n20672), .B(n20673), .Z(n20671) );
  NANDN U21006 ( .A(n20674), .B(n20675), .Z(n20673) );
  NANDN U21007 ( .A(n20675), .B(n20674), .Z(n20670) );
  ANDN U21008 ( .B(B[131]), .A(n31), .Z(n20566) );
  XNOR U21009 ( .A(n20574), .B(n20676), .Z(n20567) );
  XNOR U21010 ( .A(n20573), .B(n20571), .Z(n20676) );
  AND U21011 ( .A(n20677), .B(n20678), .Z(n20571) );
  NANDN U21012 ( .A(n20679), .B(n20680), .Z(n20678) );
  OR U21013 ( .A(n20681), .B(n20682), .Z(n20680) );
  NAND U21014 ( .A(n20682), .B(n20681), .Z(n20677) );
  ANDN U21015 ( .B(B[132]), .A(n32), .Z(n20573) );
  XNOR U21016 ( .A(n20581), .B(n20683), .Z(n20574) );
  XNOR U21017 ( .A(n20580), .B(n20578), .Z(n20683) );
  AND U21018 ( .A(n20684), .B(n20685), .Z(n20578) );
  NANDN U21019 ( .A(n20686), .B(n20687), .Z(n20685) );
  NANDN U21020 ( .A(n20688), .B(n20689), .Z(n20687) );
  NANDN U21021 ( .A(n20689), .B(n20688), .Z(n20684) );
  ANDN U21022 ( .B(B[133]), .A(n33), .Z(n20580) );
  XNOR U21023 ( .A(n20588), .B(n20690), .Z(n20581) );
  XNOR U21024 ( .A(n20587), .B(n20585), .Z(n20690) );
  AND U21025 ( .A(n20691), .B(n20692), .Z(n20585) );
  NANDN U21026 ( .A(n20693), .B(n20694), .Z(n20692) );
  OR U21027 ( .A(n20695), .B(n20696), .Z(n20694) );
  NAND U21028 ( .A(n20696), .B(n20695), .Z(n20691) );
  ANDN U21029 ( .B(B[134]), .A(n34), .Z(n20587) );
  XNOR U21030 ( .A(n20595), .B(n20697), .Z(n20588) );
  XNOR U21031 ( .A(n20594), .B(n20592), .Z(n20697) );
  AND U21032 ( .A(n20698), .B(n20699), .Z(n20592) );
  NANDN U21033 ( .A(n20700), .B(n20701), .Z(n20699) );
  NANDN U21034 ( .A(n20702), .B(n20703), .Z(n20701) );
  NANDN U21035 ( .A(n20703), .B(n20702), .Z(n20698) );
  ANDN U21036 ( .B(B[135]), .A(n35), .Z(n20594) );
  XNOR U21037 ( .A(n20602), .B(n20704), .Z(n20595) );
  XNOR U21038 ( .A(n20601), .B(n20599), .Z(n20704) );
  AND U21039 ( .A(n20705), .B(n20706), .Z(n20599) );
  NANDN U21040 ( .A(n20707), .B(n20708), .Z(n20706) );
  OR U21041 ( .A(n20709), .B(n20710), .Z(n20708) );
  NAND U21042 ( .A(n20710), .B(n20709), .Z(n20705) );
  ANDN U21043 ( .B(B[136]), .A(n36), .Z(n20601) );
  XNOR U21044 ( .A(n20609), .B(n20711), .Z(n20602) );
  XNOR U21045 ( .A(n20608), .B(n20606), .Z(n20711) );
  AND U21046 ( .A(n20712), .B(n20713), .Z(n20606) );
  NANDN U21047 ( .A(n20714), .B(n20715), .Z(n20713) );
  NANDN U21048 ( .A(n20716), .B(n20717), .Z(n20715) );
  NANDN U21049 ( .A(n20717), .B(n20716), .Z(n20712) );
  ANDN U21050 ( .B(B[137]), .A(n37), .Z(n20608) );
  XNOR U21051 ( .A(n20616), .B(n20718), .Z(n20609) );
  XNOR U21052 ( .A(n20615), .B(n20613), .Z(n20718) );
  AND U21053 ( .A(n20719), .B(n20720), .Z(n20613) );
  NANDN U21054 ( .A(n20721), .B(n20722), .Z(n20720) );
  OR U21055 ( .A(n20723), .B(n20724), .Z(n20722) );
  NAND U21056 ( .A(n20724), .B(n20723), .Z(n20719) );
  ANDN U21057 ( .B(B[138]), .A(n38), .Z(n20615) );
  XNOR U21058 ( .A(n20623), .B(n20725), .Z(n20616) );
  XNOR U21059 ( .A(n20622), .B(n20620), .Z(n20725) );
  AND U21060 ( .A(n20726), .B(n20727), .Z(n20620) );
  NANDN U21061 ( .A(n20728), .B(n20729), .Z(n20727) );
  NANDN U21062 ( .A(n20730), .B(n20731), .Z(n20729) );
  NANDN U21063 ( .A(n20731), .B(n20730), .Z(n20726) );
  ANDN U21064 ( .B(B[139]), .A(n39), .Z(n20622) );
  XNOR U21065 ( .A(n20630), .B(n20732), .Z(n20623) );
  XNOR U21066 ( .A(n20629), .B(n20627), .Z(n20732) );
  AND U21067 ( .A(n20733), .B(n20734), .Z(n20627) );
  NANDN U21068 ( .A(n20735), .B(n20736), .Z(n20734) );
  OR U21069 ( .A(n20737), .B(n20738), .Z(n20736) );
  NAND U21070 ( .A(n20738), .B(n20737), .Z(n20733) );
  ANDN U21071 ( .B(B[140]), .A(n40), .Z(n20629) );
  XNOR U21072 ( .A(n20637), .B(n20739), .Z(n20630) );
  XNOR U21073 ( .A(n20636), .B(n20634), .Z(n20739) );
  AND U21074 ( .A(n20740), .B(n20741), .Z(n20634) );
  NANDN U21075 ( .A(n20742), .B(n20743), .Z(n20741) );
  NAND U21076 ( .A(n20744), .B(n20745), .Z(n20743) );
  ANDN U21077 ( .B(B[141]), .A(n41), .Z(n20636) );
  XOR U21078 ( .A(n20643), .B(n20746), .Z(n20637) );
  XNOR U21079 ( .A(n20641), .B(n20644), .Z(n20746) );
  NAND U21080 ( .A(A[2]), .B(B[142]), .Z(n20644) );
  NANDN U21081 ( .A(n20747), .B(n20748), .Z(n20641) );
  AND U21082 ( .A(A[0]), .B(B[143]), .Z(n20748) );
  XNOR U21083 ( .A(n20646), .B(n20749), .Z(n20643) );
  NAND U21084 ( .A(A[0]), .B(B[144]), .Z(n20749) );
  NAND U21085 ( .A(B[143]), .B(A[1]), .Z(n20646) );
  NAND U21086 ( .A(n20750), .B(n20751), .Z(n467) );
  NANDN U21087 ( .A(n20752), .B(n20753), .Z(n20751) );
  OR U21088 ( .A(n20754), .B(n20755), .Z(n20753) );
  NAND U21089 ( .A(n20755), .B(n20754), .Z(n20750) );
  XOR U21090 ( .A(n469), .B(n468), .Z(\A1[141] ) );
  XOR U21091 ( .A(n20755), .B(n20756), .Z(n468) );
  XNOR U21092 ( .A(n20754), .B(n20752), .Z(n20756) );
  AND U21093 ( .A(n20757), .B(n20758), .Z(n20752) );
  NANDN U21094 ( .A(n20759), .B(n20760), .Z(n20758) );
  NANDN U21095 ( .A(n20761), .B(n20762), .Z(n20760) );
  NANDN U21096 ( .A(n20762), .B(n20761), .Z(n20757) );
  ANDN U21097 ( .B(B[128]), .A(n29), .Z(n20754) );
  XNOR U21098 ( .A(n20661), .B(n20763), .Z(n20755) );
  XNOR U21099 ( .A(n20660), .B(n20658), .Z(n20763) );
  AND U21100 ( .A(n20764), .B(n20765), .Z(n20658) );
  NANDN U21101 ( .A(n20766), .B(n20767), .Z(n20765) );
  OR U21102 ( .A(n20768), .B(n20769), .Z(n20767) );
  NAND U21103 ( .A(n20769), .B(n20768), .Z(n20764) );
  ANDN U21104 ( .B(B[129]), .A(n30), .Z(n20660) );
  XNOR U21105 ( .A(n20668), .B(n20770), .Z(n20661) );
  XNOR U21106 ( .A(n20667), .B(n20665), .Z(n20770) );
  AND U21107 ( .A(n20771), .B(n20772), .Z(n20665) );
  NANDN U21108 ( .A(n20773), .B(n20774), .Z(n20772) );
  NANDN U21109 ( .A(n20775), .B(n20776), .Z(n20774) );
  NANDN U21110 ( .A(n20776), .B(n20775), .Z(n20771) );
  ANDN U21111 ( .B(B[130]), .A(n31), .Z(n20667) );
  XNOR U21112 ( .A(n20675), .B(n20777), .Z(n20668) );
  XNOR U21113 ( .A(n20674), .B(n20672), .Z(n20777) );
  AND U21114 ( .A(n20778), .B(n20779), .Z(n20672) );
  NANDN U21115 ( .A(n20780), .B(n20781), .Z(n20779) );
  OR U21116 ( .A(n20782), .B(n20783), .Z(n20781) );
  NAND U21117 ( .A(n20783), .B(n20782), .Z(n20778) );
  ANDN U21118 ( .B(B[131]), .A(n32), .Z(n20674) );
  XNOR U21119 ( .A(n20682), .B(n20784), .Z(n20675) );
  XNOR U21120 ( .A(n20681), .B(n20679), .Z(n20784) );
  AND U21121 ( .A(n20785), .B(n20786), .Z(n20679) );
  NANDN U21122 ( .A(n20787), .B(n20788), .Z(n20786) );
  NANDN U21123 ( .A(n20789), .B(n20790), .Z(n20788) );
  NANDN U21124 ( .A(n20790), .B(n20789), .Z(n20785) );
  ANDN U21125 ( .B(B[132]), .A(n33), .Z(n20681) );
  XNOR U21126 ( .A(n20689), .B(n20791), .Z(n20682) );
  XNOR U21127 ( .A(n20688), .B(n20686), .Z(n20791) );
  AND U21128 ( .A(n20792), .B(n20793), .Z(n20686) );
  NANDN U21129 ( .A(n20794), .B(n20795), .Z(n20793) );
  OR U21130 ( .A(n20796), .B(n20797), .Z(n20795) );
  NAND U21131 ( .A(n20797), .B(n20796), .Z(n20792) );
  ANDN U21132 ( .B(B[133]), .A(n34), .Z(n20688) );
  XNOR U21133 ( .A(n20696), .B(n20798), .Z(n20689) );
  XNOR U21134 ( .A(n20695), .B(n20693), .Z(n20798) );
  AND U21135 ( .A(n20799), .B(n20800), .Z(n20693) );
  NANDN U21136 ( .A(n20801), .B(n20802), .Z(n20800) );
  NANDN U21137 ( .A(n20803), .B(n20804), .Z(n20802) );
  NANDN U21138 ( .A(n20804), .B(n20803), .Z(n20799) );
  ANDN U21139 ( .B(B[134]), .A(n35), .Z(n20695) );
  XNOR U21140 ( .A(n20703), .B(n20805), .Z(n20696) );
  XNOR U21141 ( .A(n20702), .B(n20700), .Z(n20805) );
  AND U21142 ( .A(n20806), .B(n20807), .Z(n20700) );
  NANDN U21143 ( .A(n20808), .B(n20809), .Z(n20807) );
  OR U21144 ( .A(n20810), .B(n20811), .Z(n20809) );
  NAND U21145 ( .A(n20811), .B(n20810), .Z(n20806) );
  ANDN U21146 ( .B(B[135]), .A(n36), .Z(n20702) );
  XNOR U21147 ( .A(n20710), .B(n20812), .Z(n20703) );
  XNOR U21148 ( .A(n20709), .B(n20707), .Z(n20812) );
  AND U21149 ( .A(n20813), .B(n20814), .Z(n20707) );
  NANDN U21150 ( .A(n20815), .B(n20816), .Z(n20814) );
  NANDN U21151 ( .A(n20817), .B(n20818), .Z(n20816) );
  NANDN U21152 ( .A(n20818), .B(n20817), .Z(n20813) );
  ANDN U21153 ( .B(B[136]), .A(n37), .Z(n20709) );
  XNOR U21154 ( .A(n20717), .B(n20819), .Z(n20710) );
  XNOR U21155 ( .A(n20716), .B(n20714), .Z(n20819) );
  AND U21156 ( .A(n20820), .B(n20821), .Z(n20714) );
  NANDN U21157 ( .A(n20822), .B(n20823), .Z(n20821) );
  OR U21158 ( .A(n20824), .B(n20825), .Z(n20823) );
  NAND U21159 ( .A(n20825), .B(n20824), .Z(n20820) );
  ANDN U21160 ( .B(B[137]), .A(n38), .Z(n20716) );
  XNOR U21161 ( .A(n20724), .B(n20826), .Z(n20717) );
  XNOR U21162 ( .A(n20723), .B(n20721), .Z(n20826) );
  AND U21163 ( .A(n20827), .B(n20828), .Z(n20721) );
  NANDN U21164 ( .A(n20829), .B(n20830), .Z(n20828) );
  NANDN U21165 ( .A(n20831), .B(n20832), .Z(n20830) );
  NANDN U21166 ( .A(n20832), .B(n20831), .Z(n20827) );
  ANDN U21167 ( .B(B[138]), .A(n39), .Z(n20723) );
  XNOR U21168 ( .A(n20731), .B(n20833), .Z(n20724) );
  XNOR U21169 ( .A(n20730), .B(n20728), .Z(n20833) );
  AND U21170 ( .A(n20834), .B(n20835), .Z(n20728) );
  NANDN U21171 ( .A(n20836), .B(n20837), .Z(n20835) );
  OR U21172 ( .A(n20838), .B(n20839), .Z(n20837) );
  NAND U21173 ( .A(n20839), .B(n20838), .Z(n20834) );
  ANDN U21174 ( .B(B[139]), .A(n40), .Z(n20730) );
  XNOR U21175 ( .A(n20738), .B(n20840), .Z(n20731) );
  XNOR U21176 ( .A(n20737), .B(n20735), .Z(n20840) );
  AND U21177 ( .A(n20841), .B(n20842), .Z(n20735) );
  NANDN U21178 ( .A(n20843), .B(n20844), .Z(n20842) );
  NAND U21179 ( .A(n20845), .B(n20846), .Z(n20844) );
  ANDN U21180 ( .B(B[140]), .A(n41), .Z(n20737) );
  XOR U21181 ( .A(n20744), .B(n20847), .Z(n20738) );
  XNOR U21182 ( .A(n20742), .B(n20745), .Z(n20847) );
  NAND U21183 ( .A(A[2]), .B(B[141]), .Z(n20745) );
  NANDN U21184 ( .A(n20848), .B(n20849), .Z(n20742) );
  AND U21185 ( .A(A[0]), .B(B[142]), .Z(n20849) );
  XNOR U21186 ( .A(n20747), .B(n20850), .Z(n20744) );
  NAND U21187 ( .A(A[0]), .B(B[143]), .Z(n20850) );
  NAND U21188 ( .A(B[142]), .B(A[1]), .Z(n20747) );
  NAND U21189 ( .A(n20851), .B(n20852), .Z(n469) );
  NANDN U21190 ( .A(n20853), .B(n20854), .Z(n20852) );
  OR U21191 ( .A(n20855), .B(n20856), .Z(n20854) );
  NAND U21192 ( .A(n20856), .B(n20855), .Z(n20851) );
  XOR U21193 ( .A(n471), .B(n470), .Z(\A1[140] ) );
  XOR U21194 ( .A(n20856), .B(n20857), .Z(n470) );
  XNOR U21195 ( .A(n20855), .B(n20853), .Z(n20857) );
  AND U21196 ( .A(n20858), .B(n20859), .Z(n20853) );
  NANDN U21197 ( .A(n20860), .B(n20861), .Z(n20859) );
  NANDN U21198 ( .A(n20862), .B(n20863), .Z(n20861) );
  NANDN U21199 ( .A(n20863), .B(n20862), .Z(n20858) );
  ANDN U21200 ( .B(B[127]), .A(n29), .Z(n20855) );
  XNOR U21201 ( .A(n20762), .B(n20864), .Z(n20856) );
  XNOR U21202 ( .A(n20761), .B(n20759), .Z(n20864) );
  AND U21203 ( .A(n20865), .B(n20866), .Z(n20759) );
  NANDN U21204 ( .A(n20867), .B(n20868), .Z(n20866) );
  OR U21205 ( .A(n20869), .B(n20870), .Z(n20868) );
  NAND U21206 ( .A(n20870), .B(n20869), .Z(n20865) );
  ANDN U21207 ( .B(B[128]), .A(n30), .Z(n20761) );
  XNOR U21208 ( .A(n20769), .B(n20871), .Z(n20762) );
  XNOR U21209 ( .A(n20768), .B(n20766), .Z(n20871) );
  AND U21210 ( .A(n20872), .B(n20873), .Z(n20766) );
  NANDN U21211 ( .A(n20874), .B(n20875), .Z(n20873) );
  NANDN U21212 ( .A(n20876), .B(n20877), .Z(n20875) );
  NANDN U21213 ( .A(n20877), .B(n20876), .Z(n20872) );
  ANDN U21214 ( .B(B[129]), .A(n31), .Z(n20768) );
  XNOR U21215 ( .A(n20776), .B(n20878), .Z(n20769) );
  XNOR U21216 ( .A(n20775), .B(n20773), .Z(n20878) );
  AND U21217 ( .A(n20879), .B(n20880), .Z(n20773) );
  NANDN U21218 ( .A(n20881), .B(n20882), .Z(n20880) );
  OR U21219 ( .A(n20883), .B(n20884), .Z(n20882) );
  NAND U21220 ( .A(n20884), .B(n20883), .Z(n20879) );
  ANDN U21221 ( .B(B[130]), .A(n32), .Z(n20775) );
  XNOR U21222 ( .A(n20783), .B(n20885), .Z(n20776) );
  XNOR U21223 ( .A(n20782), .B(n20780), .Z(n20885) );
  AND U21224 ( .A(n20886), .B(n20887), .Z(n20780) );
  NANDN U21225 ( .A(n20888), .B(n20889), .Z(n20887) );
  NANDN U21226 ( .A(n20890), .B(n20891), .Z(n20889) );
  NANDN U21227 ( .A(n20891), .B(n20890), .Z(n20886) );
  ANDN U21228 ( .B(B[131]), .A(n33), .Z(n20782) );
  XNOR U21229 ( .A(n20790), .B(n20892), .Z(n20783) );
  XNOR U21230 ( .A(n20789), .B(n20787), .Z(n20892) );
  AND U21231 ( .A(n20893), .B(n20894), .Z(n20787) );
  NANDN U21232 ( .A(n20895), .B(n20896), .Z(n20894) );
  OR U21233 ( .A(n20897), .B(n20898), .Z(n20896) );
  NAND U21234 ( .A(n20898), .B(n20897), .Z(n20893) );
  ANDN U21235 ( .B(B[132]), .A(n34), .Z(n20789) );
  XNOR U21236 ( .A(n20797), .B(n20899), .Z(n20790) );
  XNOR U21237 ( .A(n20796), .B(n20794), .Z(n20899) );
  AND U21238 ( .A(n20900), .B(n20901), .Z(n20794) );
  NANDN U21239 ( .A(n20902), .B(n20903), .Z(n20901) );
  NANDN U21240 ( .A(n20904), .B(n20905), .Z(n20903) );
  NANDN U21241 ( .A(n20905), .B(n20904), .Z(n20900) );
  ANDN U21242 ( .B(B[133]), .A(n35), .Z(n20796) );
  XNOR U21243 ( .A(n20804), .B(n20906), .Z(n20797) );
  XNOR U21244 ( .A(n20803), .B(n20801), .Z(n20906) );
  AND U21245 ( .A(n20907), .B(n20908), .Z(n20801) );
  NANDN U21246 ( .A(n20909), .B(n20910), .Z(n20908) );
  OR U21247 ( .A(n20911), .B(n20912), .Z(n20910) );
  NAND U21248 ( .A(n20912), .B(n20911), .Z(n20907) );
  ANDN U21249 ( .B(B[134]), .A(n36), .Z(n20803) );
  XNOR U21250 ( .A(n20811), .B(n20913), .Z(n20804) );
  XNOR U21251 ( .A(n20810), .B(n20808), .Z(n20913) );
  AND U21252 ( .A(n20914), .B(n20915), .Z(n20808) );
  NANDN U21253 ( .A(n20916), .B(n20917), .Z(n20915) );
  NANDN U21254 ( .A(n20918), .B(n20919), .Z(n20917) );
  NANDN U21255 ( .A(n20919), .B(n20918), .Z(n20914) );
  ANDN U21256 ( .B(B[135]), .A(n37), .Z(n20810) );
  XNOR U21257 ( .A(n20818), .B(n20920), .Z(n20811) );
  XNOR U21258 ( .A(n20817), .B(n20815), .Z(n20920) );
  AND U21259 ( .A(n20921), .B(n20922), .Z(n20815) );
  NANDN U21260 ( .A(n20923), .B(n20924), .Z(n20922) );
  OR U21261 ( .A(n20925), .B(n20926), .Z(n20924) );
  NAND U21262 ( .A(n20926), .B(n20925), .Z(n20921) );
  ANDN U21263 ( .B(B[136]), .A(n38), .Z(n20817) );
  XNOR U21264 ( .A(n20825), .B(n20927), .Z(n20818) );
  XNOR U21265 ( .A(n20824), .B(n20822), .Z(n20927) );
  AND U21266 ( .A(n20928), .B(n20929), .Z(n20822) );
  NANDN U21267 ( .A(n20930), .B(n20931), .Z(n20929) );
  NANDN U21268 ( .A(n20932), .B(n20933), .Z(n20931) );
  NANDN U21269 ( .A(n20933), .B(n20932), .Z(n20928) );
  ANDN U21270 ( .B(B[137]), .A(n39), .Z(n20824) );
  XNOR U21271 ( .A(n20832), .B(n20934), .Z(n20825) );
  XNOR U21272 ( .A(n20831), .B(n20829), .Z(n20934) );
  AND U21273 ( .A(n20935), .B(n20936), .Z(n20829) );
  NANDN U21274 ( .A(n20937), .B(n20938), .Z(n20936) );
  OR U21275 ( .A(n20939), .B(n20940), .Z(n20938) );
  NAND U21276 ( .A(n20940), .B(n20939), .Z(n20935) );
  ANDN U21277 ( .B(B[138]), .A(n40), .Z(n20831) );
  XNOR U21278 ( .A(n20839), .B(n20941), .Z(n20832) );
  XNOR U21279 ( .A(n20838), .B(n20836), .Z(n20941) );
  AND U21280 ( .A(n20942), .B(n20943), .Z(n20836) );
  NANDN U21281 ( .A(n20944), .B(n20945), .Z(n20943) );
  NAND U21282 ( .A(n20946), .B(n20947), .Z(n20945) );
  ANDN U21283 ( .B(B[139]), .A(n41), .Z(n20838) );
  XOR U21284 ( .A(n20845), .B(n20948), .Z(n20839) );
  XNOR U21285 ( .A(n20843), .B(n20846), .Z(n20948) );
  NAND U21286 ( .A(A[2]), .B(B[140]), .Z(n20846) );
  NANDN U21287 ( .A(n20949), .B(n20950), .Z(n20843) );
  AND U21288 ( .A(A[0]), .B(B[141]), .Z(n20950) );
  XNOR U21289 ( .A(n20848), .B(n20951), .Z(n20845) );
  NAND U21290 ( .A(A[0]), .B(B[142]), .Z(n20951) );
  NAND U21291 ( .A(B[141]), .B(A[1]), .Z(n20848) );
  NAND U21292 ( .A(n20952), .B(n20953), .Z(n471) );
  NANDN U21293 ( .A(n20954), .B(n20955), .Z(n20953) );
  OR U21294 ( .A(n20956), .B(n20957), .Z(n20955) );
  NAND U21295 ( .A(n20957), .B(n20956), .Z(n20952) );
  XOR U21296 ( .A(n19947), .B(n20958), .Z(\A1[13] ) );
  XNOR U21297 ( .A(n19946), .B(n19944), .Z(n20958) );
  AND U21298 ( .A(n20959), .B(n20960), .Z(n19944) );
  NAND U21299 ( .A(n20961), .B(n20962), .Z(n20960) );
  NANDN U21300 ( .A(n20963), .B(n20964), .Z(n20961) );
  NANDN U21301 ( .A(n20964), .B(n20963), .Z(n20959) );
  ANDN U21302 ( .B(B[0]), .A(n29), .Z(n19946) );
  XNOR U21303 ( .A(n19853), .B(n20965), .Z(n19947) );
  XNOR U21304 ( .A(n19852), .B(n19850), .Z(n20965) );
  AND U21305 ( .A(n20966), .B(n20967), .Z(n19850) );
  NANDN U21306 ( .A(n20968), .B(n20969), .Z(n20967) );
  OR U21307 ( .A(n20970), .B(n20971), .Z(n20969) );
  NAND U21308 ( .A(n20971), .B(n20970), .Z(n20966) );
  ANDN U21309 ( .B(B[1]), .A(n30), .Z(n19852) );
  XNOR U21310 ( .A(n19860), .B(n20972), .Z(n19853) );
  XNOR U21311 ( .A(n19859), .B(n19857), .Z(n20972) );
  AND U21312 ( .A(n20973), .B(n20974), .Z(n19857) );
  NANDN U21313 ( .A(n20975), .B(n20976), .Z(n20974) );
  NANDN U21314 ( .A(n20977), .B(n20978), .Z(n20976) );
  NANDN U21315 ( .A(n20978), .B(n20977), .Z(n20973) );
  ANDN U21316 ( .B(B[2]), .A(n31), .Z(n19859) );
  XNOR U21317 ( .A(n19867), .B(n20979), .Z(n19860) );
  XNOR U21318 ( .A(n19866), .B(n19864), .Z(n20979) );
  AND U21319 ( .A(n20980), .B(n20981), .Z(n19864) );
  NANDN U21320 ( .A(n20982), .B(n20983), .Z(n20981) );
  OR U21321 ( .A(n20984), .B(n20985), .Z(n20983) );
  NAND U21322 ( .A(n20985), .B(n20984), .Z(n20980) );
  ANDN U21323 ( .B(B[3]), .A(n32), .Z(n19866) );
  XNOR U21324 ( .A(n19874), .B(n20986), .Z(n19867) );
  XNOR U21325 ( .A(n19873), .B(n19871), .Z(n20986) );
  AND U21326 ( .A(n20987), .B(n20988), .Z(n19871) );
  NANDN U21327 ( .A(n20989), .B(n20990), .Z(n20988) );
  NANDN U21328 ( .A(n20991), .B(n20992), .Z(n20990) );
  NANDN U21329 ( .A(n20992), .B(n20991), .Z(n20987) );
  ANDN U21330 ( .B(B[4]), .A(n33), .Z(n19873) );
  XNOR U21331 ( .A(n19881), .B(n20993), .Z(n19874) );
  XNOR U21332 ( .A(n19880), .B(n19878), .Z(n20993) );
  AND U21333 ( .A(n20994), .B(n20995), .Z(n19878) );
  NANDN U21334 ( .A(n20996), .B(n20997), .Z(n20995) );
  OR U21335 ( .A(n20998), .B(n20999), .Z(n20997) );
  NAND U21336 ( .A(n20999), .B(n20998), .Z(n20994) );
  ANDN U21337 ( .B(B[5]), .A(n34), .Z(n19880) );
  XNOR U21338 ( .A(n19888), .B(n21000), .Z(n19881) );
  XNOR U21339 ( .A(n19887), .B(n19885), .Z(n21000) );
  AND U21340 ( .A(n21001), .B(n21002), .Z(n19885) );
  NANDN U21341 ( .A(n21003), .B(n21004), .Z(n21002) );
  NANDN U21342 ( .A(n21005), .B(n21006), .Z(n21004) );
  NANDN U21343 ( .A(n21006), .B(n21005), .Z(n21001) );
  ANDN U21344 ( .B(B[6]), .A(n35), .Z(n19887) );
  XNOR U21345 ( .A(n19895), .B(n21007), .Z(n19888) );
  XNOR U21346 ( .A(n19894), .B(n19892), .Z(n21007) );
  AND U21347 ( .A(n21008), .B(n21009), .Z(n19892) );
  NANDN U21348 ( .A(n21010), .B(n21011), .Z(n21009) );
  OR U21349 ( .A(n21012), .B(n21013), .Z(n21011) );
  NAND U21350 ( .A(n21013), .B(n21012), .Z(n21008) );
  ANDN U21351 ( .B(B[7]), .A(n36), .Z(n19894) );
  XNOR U21352 ( .A(n19902), .B(n21014), .Z(n19895) );
  XNOR U21353 ( .A(n19901), .B(n19899), .Z(n21014) );
  AND U21354 ( .A(n21015), .B(n21016), .Z(n19899) );
  NANDN U21355 ( .A(n21017), .B(n21018), .Z(n21016) );
  NANDN U21356 ( .A(n21019), .B(n21020), .Z(n21018) );
  NANDN U21357 ( .A(n21020), .B(n21019), .Z(n21015) );
  ANDN U21358 ( .B(B[8]), .A(n37), .Z(n19901) );
  XNOR U21359 ( .A(n19909), .B(n21021), .Z(n19902) );
  XNOR U21360 ( .A(n19908), .B(n19906), .Z(n21021) );
  AND U21361 ( .A(n21022), .B(n21023), .Z(n19906) );
  NANDN U21362 ( .A(n21024), .B(n21025), .Z(n21023) );
  OR U21363 ( .A(n21026), .B(n21027), .Z(n21025) );
  NAND U21364 ( .A(n21027), .B(n21026), .Z(n21022) );
  ANDN U21365 ( .B(B[9]), .A(n38), .Z(n19908) );
  XNOR U21366 ( .A(n19916), .B(n21028), .Z(n19909) );
  XNOR U21367 ( .A(n19915), .B(n19913), .Z(n21028) );
  AND U21368 ( .A(n21029), .B(n21030), .Z(n19913) );
  NANDN U21369 ( .A(n21031), .B(n21032), .Z(n21030) );
  NANDN U21370 ( .A(n21033), .B(n21034), .Z(n21032) );
  NANDN U21371 ( .A(n21034), .B(n21033), .Z(n21029) );
  ANDN U21372 ( .B(B[10]), .A(n39), .Z(n19915) );
  XNOR U21373 ( .A(n19923), .B(n21035), .Z(n19916) );
  XNOR U21374 ( .A(n19922), .B(n19920), .Z(n21035) );
  AND U21375 ( .A(n21036), .B(n21037), .Z(n19920) );
  NANDN U21376 ( .A(n21038), .B(n21039), .Z(n21037) );
  OR U21377 ( .A(n21040), .B(n21041), .Z(n21039) );
  NAND U21378 ( .A(n21041), .B(n21040), .Z(n21036) );
  ANDN U21379 ( .B(B[11]), .A(n40), .Z(n19922) );
  XNOR U21380 ( .A(n19930), .B(n21042), .Z(n19923) );
  XNOR U21381 ( .A(n19929), .B(n19927), .Z(n21042) );
  AND U21382 ( .A(n21043), .B(n21044), .Z(n19927) );
  NANDN U21383 ( .A(n21045), .B(n21046), .Z(n21044) );
  NAND U21384 ( .A(n21047), .B(n21048), .Z(n21046) );
  ANDN U21385 ( .B(B[12]), .A(n41), .Z(n19929) );
  XOR U21386 ( .A(n19936), .B(n21049), .Z(n19930) );
  XNOR U21387 ( .A(n19934), .B(n19937), .Z(n21049) );
  NAND U21388 ( .A(A[2]), .B(B[13]), .Z(n19937) );
  NANDN U21389 ( .A(n21050), .B(n21051), .Z(n19934) );
  AND U21390 ( .A(A[0]), .B(B[14]), .Z(n21051) );
  XNOR U21391 ( .A(n19939), .B(n21052), .Z(n19936) );
  NAND U21392 ( .A(A[0]), .B(B[15]), .Z(n21052) );
  NAND U21393 ( .A(B[14]), .B(A[1]), .Z(n19939) );
  XOR U21394 ( .A(n473), .B(n472), .Z(\A1[139] ) );
  XOR U21395 ( .A(n20957), .B(n21053), .Z(n472) );
  XNOR U21396 ( .A(n20956), .B(n20954), .Z(n21053) );
  AND U21397 ( .A(n21054), .B(n21055), .Z(n20954) );
  NANDN U21398 ( .A(n21056), .B(n21057), .Z(n21055) );
  NANDN U21399 ( .A(n21058), .B(n21059), .Z(n21057) );
  NANDN U21400 ( .A(n21059), .B(n21058), .Z(n21054) );
  ANDN U21401 ( .B(B[126]), .A(n29), .Z(n20956) );
  XNOR U21402 ( .A(n20863), .B(n21060), .Z(n20957) );
  XNOR U21403 ( .A(n20862), .B(n20860), .Z(n21060) );
  AND U21404 ( .A(n21061), .B(n21062), .Z(n20860) );
  NANDN U21405 ( .A(n21063), .B(n21064), .Z(n21062) );
  OR U21406 ( .A(n21065), .B(n21066), .Z(n21064) );
  NAND U21407 ( .A(n21066), .B(n21065), .Z(n21061) );
  ANDN U21408 ( .B(B[127]), .A(n30), .Z(n20862) );
  XNOR U21409 ( .A(n20870), .B(n21067), .Z(n20863) );
  XNOR U21410 ( .A(n20869), .B(n20867), .Z(n21067) );
  AND U21411 ( .A(n21068), .B(n21069), .Z(n20867) );
  NANDN U21412 ( .A(n21070), .B(n21071), .Z(n21069) );
  NANDN U21413 ( .A(n21072), .B(n21073), .Z(n21071) );
  NANDN U21414 ( .A(n21073), .B(n21072), .Z(n21068) );
  ANDN U21415 ( .B(B[128]), .A(n31), .Z(n20869) );
  XNOR U21416 ( .A(n20877), .B(n21074), .Z(n20870) );
  XNOR U21417 ( .A(n20876), .B(n20874), .Z(n21074) );
  AND U21418 ( .A(n21075), .B(n21076), .Z(n20874) );
  NANDN U21419 ( .A(n21077), .B(n21078), .Z(n21076) );
  OR U21420 ( .A(n21079), .B(n21080), .Z(n21078) );
  NAND U21421 ( .A(n21080), .B(n21079), .Z(n21075) );
  ANDN U21422 ( .B(B[129]), .A(n32), .Z(n20876) );
  XNOR U21423 ( .A(n20884), .B(n21081), .Z(n20877) );
  XNOR U21424 ( .A(n20883), .B(n20881), .Z(n21081) );
  AND U21425 ( .A(n21082), .B(n21083), .Z(n20881) );
  NANDN U21426 ( .A(n21084), .B(n21085), .Z(n21083) );
  NANDN U21427 ( .A(n21086), .B(n21087), .Z(n21085) );
  NANDN U21428 ( .A(n21087), .B(n21086), .Z(n21082) );
  ANDN U21429 ( .B(B[130]), .A(n33), .Z(n20883) );
  XNOR U21430 ( .A(n20891), .B(n21088), .Z(n20884) );
  XNOR U21431 ( .A(n20890), .B(n20888), .Z(n21088) );
  AND U21432 ( .A(n21089), .B(n21090), .Z(n20888) );
  NANDN U21433 ( .A(n21091), .B(n21092), .Z(n21090) );
  OR U21434 ( .A(n21093), .B(n21094), .Z(n21092) );
  NAND U21435 ( .A(n21094), .B(n21093), .Z(n21089) );
  ANDN U21436 ( .B(B[131]), .A(n34), .Z(n20890) );
  XNOR U21437 ( .A(n20898), .B(n21095), .Z(n20891) );
  XNOR U21438 ( .A(n20897), .B(n20895), .Z(n21095) );
  AND U21439 ( .A(n21096), .B(n21097), .Z(n20895) );
  NANDN U21440 ( .A(n21098), .B(n21099), .Z(n21097) );
  NANDN U21441 ( .A(n21100), .B(n21101), .Z(n21099) );
  NANDN U21442 ( .A(n21101), .B(n21100), .Z(n21096) );
  ANDN U21443 ( .B(B[132]), .A(n35), .Z(n20897) );
  XNOR U21444 ( .A(n20905), .B(n21102), .Z(n20898) );
  XNOR U21445 ( .A(n20904), .B(n20902), .Z(n21102) );
  AND U21446 ( .A(n21103), .B(n21104), .Z(n20902) );
  NANDN U21447 ( .A(n21105), .B(n21106), .Z(n21104) );
  OR U21448 ( .A(n21107), .B(n21108), .Z(n21106) );
  NAND U21449 ( .A(n21108), .B(n21107), .Z(n21103) );
  ANDN U21450 ( .B(B[133]), .A(n36), .Z(n20904) );
  XNOR U21451 ( .A(n20912), .B(n21109), .Z(n20905) );
  XNOR U21452 ( .A(n20911), .B(n20909), .Z(n21109) );
  AND U21453 ( .A(n21110), .B(n21111), .Z(n20909) );
  NANDN U21454 ( .A(n21112), .B(n21113), .Z(n21111) );
  NANDN U21455 ( .A(n21114), .B(n21115), .Z(n21113) );
  NANDN U21456 ( .A(n21115), .B(n21114), .Z(n21110) );
  ANDN U21457 ( .B(B[134]), .A(n37), .Z(n20911) );
  XNOR U21458 ( .A(n20919), .B(n21116), .Z(n20912) );
  XNOR U21459 ( .A(n20918), .B(n20916), .Z(n21116) );
  AND U21460 ( .A(n21117), .B(n21118), .Z(n20916) );
  NANDN U21461 ( .A(n21119), .B(n21120), .Z(n21118) );
  OR U21462 ( .A(n21121), .B(n21122), .Z(n21120) );
  NAND U21463 ( .A(n21122), .B(n21121), .Z(n21117) );
  ANDN U21464 ( .B(B[135]), .A(n38), .Z(n20918) );
  XNOR U21465 ( .A(n20926), .B(n21123), .Z(n20919) );
  XNOR U21466 ( .A(n20925), .B(n20923), .Z(n21123) );
  AND U21467 ( .A(n21124), .B(n21125), .Z(n20923) );
  NANDN U21468 ( .A(n21126), .B(n21127), .Z(n21125) );
  NANDN U21469 ( .A(n21128), .B(n21129), .Z(n21127) );
  NANDN U21470 ( .A(n21129), .B(n21128), .Z(n21124) );
  ANDN U21471 ( .B(B[136]), .A(n39), .Z(n20925) );
  XNOR U21472 ( .A(n20933), .B(n21130), .Z(n20926) );
  XNOR U21473 ( .A(n20932), .B(n20930), .Z(n21130) );
  AND U21474 ( .A(n21131), .B(n21132), .Z(n20930) );
  NANDN U21475 ( .A(n21133), .B(n21134), .Z(n21132) );
  OR U21476 ( .A(n21135), .B(n21136), .Z(n21134) );
  NAND U21477 ( .A(n21136), .B(n21135), .Z(n21131) );
  ANDN U21478 ( .B(B[137]), .A(n40), .Z(n20932) );
  XNOR U21479 ( .A(n20940), .B(n21137), .Z(n20933) );
  XNOR U21480 ( .A(n20939), .B(n20937), .Z(n21137) );
  AND U21481 ( .A(n21138), .B(n21139), .Z(n20937) );
  NANDN U21482 ( .A(n21140), .B(n21141), .Z(n21139) );
  NAND U21483 ( .A(n21142), .B(n21143), .Z(n21141) );
  ANDN U21484 ( .B(B[138]), .A(n41), .Z(n20939) );
  XOR U21485 ( .A(n20946), .B(n21144), .Z(n20940) );
  XNOR U21486 ( .A(n20944), .B(n20947), .Z(n21144) );
  NAND U21487 ( .A(A[2]), .B(B[139]), .Z(n20947) );
  NANDN U21488 ( .A(n21145), .B(n21146), .Z(n20944) );
  AND U21489 ( .A(A[0]), .B(B[140]), .Z(n21146) );
  XNOR U21490 ( .A(n20949), .B(n21147), .Z(n20946) );
  NAND U21491 ( .A(A[0]), .B(B[141]), .Z(n21147) );
  NAND U21492 ( .A(B[140]), .B(A[1]), .Z(n20949) );
  NAND U21493 ( .A(n21148), .B(n21149), .Z(n473) );
  NANDN U21494 ( .A(n21150), .B(n21151), .Z(n21149) );
  OR U21495 ( .A(n21152), .B(n21153), .Z(n21151) );
  NAND U21496 ( .A(n21153), .B(n21152), .Z(n21148) );
  XOR U21497 ( .A(n475), .B(n474), .Z(\A1[138] ) );
  XOR U21498 ( .A(n21153), .B(n21154), .Z(n474) );
  XNOR U21499 ( .A(n21152), .B(n21150), .Z(n21154) );
  AND U21500 ( .A(n21155), .B(n21156), .Z(n21150) );
  NANDN U21501 ( .A(n21157), .B(n21158), .Z(n21156) );
  NANDN U21502 ( .A(n21159), .B(n21160), .Z(n21158) );
  NANDN U21503 ( .A(n21160), .B(n21159), .Z(n21155) );
  ANDN U21504 ( .B(B[125]), .A(n29), .Z(n21152) );
  XNOR U21505 ( .A(n21059), .B(n21161), .Z(n21153) );
  XNOR U21506 ( .A(n21058), .B(n21056), .Z(n21161) );
  AND U21507 ( .A(n21162), .B(n21163), .Z(n21056) );
  NANDN U21508 ( .A(n21164), .B(n21165), .Z(n21163) );
  OR U21509 ( .A(n21166), .B(n21167), .Z(n21165) );
  NAND U21510 ( .A(n21167), .B(n21166), .Z(n21162) );
  ANDN U21511 ( .B(B[126]), .A(n30), .Z(n21058) );
  XNOR U21512 ( .A(n21066), .B(n21168), .Z(n21059) );
  XNOR U21513 ( .A(n21065), .B(n21063), .Z(n21168) );
  AND U21514 ( .A(n21169), .B(n21170), .Z(n21063) );
  NANDN U21515 ( .A(n21171), .B(n21172), .Z(n21170) );
  NANDN U21516 ( .A(n21173), .B(n21174), .Z(n21172) );
  NANDN U21517 ( .A(n21174), .B(n21173), .Z(n21169) );
  ANDN U21518 ( .B(B[127]), .A(n31), .Z(n21065) );
  XNOR U21519 ( .A(n21073), .B(n21175), .Z(n21066) );
  XNOR U21520 ( .A(n21072), .B(n21070), .Z(n21175) );
  AND U21521 ( .A(n21176), .B(n21177), .Z(n21070) );
  NANDN U21522 ( .A(n21178), .B(n21179), .Z(n21177) );
  OR U21523 ( .A(n21180), .B(n21181), .Z(n21179) );
  NAND U21524 ( .A(n21181), .B(n21180), .Z(n21176) );
  ANDN U21525 ( .B(B[128]), .A(n32), .Z(n21072) );
  XNOR U21526 ( .A(n21080), .B(n21182), .Z(n21073) );
  XNOR U21527 ( .A(n21079), .B(n21077), .Z(n21182) );
  AND U21528 ( .A(n21183), .B(n21184), .Z(n21077) );
  NANDN U21529 ( .A(n21185), .B(n21186), .Z(n21184) );
  NANDN U21530 ( .A(n21187), .B(n21188), .Z(n21186) );
  NANDN U21531 ( .A(n21188), .B(n21187), .Z(n21183) );
  ANDN U21532 ( .B(B[129]), .A(n33), .Z(n21079) );
  XNOR U21533 ( .A(n21087), .B(n21189), .Z(n21080) );
  XNOR U21534 ( .A(n21086), .B(n21084), .Z(n21189) );
  AND U21535 ( .A(n21190), .B(n21191), .Z(n21084) );
  NANDN U21536 ( .A(n21192), .B(n21193), .Z(n21191) );
  OR U21537 ( .A(n21194), .B(n21195), .Z(n21193) );
  NAND U21538 ( .A(n21195), .B(n21194), .Z(n21190) );
  ANDN U21539 ( .B(B[130]), .A(n34), .Z(n21086) );
  XNOR U21540 ( .A(n21094), .B(n21196), .Z(n21087) );
  XNOR U21541 ( .A(n21093), .B(n21091), .Z(n21196) );
  AND U21542 ( .A(n21197), .B(n21198), .Z(n21091) );
  NANDN U21543 ( .A(n21199), .B(n21200), .Z(n21198) );
  NANDN U21544 ( .A(n21201), .B(n21202), .Z(n21200) );
  NANDN U21545 ( .A(n21202), .B(n21201), .Z(n21197) );
  ANDN U21546 ( .B(B[131]), .A(n35), .Z(n21093) );
  XNOR U21547 ( .A(n21101), .B(n21203), .Z(n21094) );
  XNOR U21548 ( .A(n21100), .B(n21098), .Z(n21203) );
  AND U21549 ( .A(n21204), .B(n21205), .Z(n21098) );
  NANDN U21550 ( .A(n21206), .B(n21207), .Z(n21205) );
  OR U21551 ( .A(n21208), .B(n21209), .Z(n21207) );
  NAND U21552 ( .A(n21209), .B(n21208), .Z(n21204) );
  ANDN U21553 ( .B(B[132]), .A(n36), .Z(n21100) );
  XNOR U21554 ( .A(n21108), .B(n21210), .Z(n21101) );
  XNOR U21555 ( .A(n21107), .B(n21105), .Z(n21210) );
  AND U21556 ( .A(n21211), .B(n21212), .Z(n21105) );
  NANDN U21557 ( .A(n21213), .B(n21214), .Z(n21212) );
  NANDN U21558 ( .A(n21215), .B(n21216), .Z(n21214) );
  NANDN U21559 ( .A(n21216), .B(n21215), .Z(n21211) );
  ANDN U21560 ( .B(B[133]), .A(n37), .Z(n21107) );
  XNOR U21561 ( .A(n21115), .B(n21217), .Z(n21108) );
  XNOR U21562 ( .A(n21114), .B(n21112), .Z(n21217) );
  AND U21563 ( .A(n21218), .B(n21219), .Z(n21112) );
  NANDN U21564 ( .A(n21220), .B(n21221), .Z(n21219) );
  OR U21565 ( .A(n21222), .B(n21223), .Z(n21221) );
  NAND U21566 ( .A(n21223), .B(n21222), .Z(n21218) );
  ANDN U21567 ( .B(B[134]), .A(n38), .Z(n21114) );
  XNOR U21568 ( .A(n21122), .B(n21224), .Z(n21115) );
  XNOR U21569 ( .A(n21121), .B(n21119), .Z(n21224) );
  AND U21570 ( .A(n21225), .B(n21226), .Z(n21119) );
  NANDN U21571 ( .A(n21227), .B(n21228), .Z(n21226) );
  NANDN U21572 ( .A(n21229), .B(n21230), .Z(n21228) );
  NANDN U21573 ( .A(n21230), .B(n21229), .Z(n21225) );
  ANDN U21574 ( .B(B[135]), .A(n39), .Z(n21121) );
  XNOR U21575 ( .A(n21129), .B(n21231), .Z(n21122) );
  XNOR U21576 ( .A(n21128), .B(n21126), .Z(n21231) );
  AND U21577 ( .A(n21232), .B(n21233), .Z(n21126) );
  NANDN U21578 ( .A(n21234), .B(n21235), .Z(n21233) );
  OR U21579 ( .A(n21236), .B(n21237), .Z(n21235) );
  NAND U21580 ( .A(n21237), .B(n21236), .Z(n21232) );
  ANDN U21581 ( .B(B[136]), .A(n40), .Z(n21128) );
  XNOR U21582 ( .A(n21136), .B(n21238), .Z(n21129) );
  XNOR U21583 ( .A(n21135), .B(n21133), .Z(n21238) );
  AND U21584 ( .A(n21239), .B(n21240), .Z(n21133) );
  NANDN U21585 ( .A(n21241), .B(n21242), .Z(n21240) );
  NAND U21586 ( .A(n21243), .B(n21244), .Z(n21242) );
  ANDN U21587 ( .B(B[137]), .A(n41), .Z(n21135) );
  XOR U21588 ( .A(n21142), .B(n21245), .Z(n21136) );
  XNOR U21589 ( .A(n21140), .B(n21143), .Z(n21245) );
  NAND U21590 ( .A(A[2]), .B(B[138]), .Z(n21143) );
  NANDN U21591 ( .A(n21246), .B(n21247), .Z(n21140) );
  AND U21592 ( .A(A[0]), .B(B[139]), .Z(n21247) );
  XNOR U21593 ( .A(n21145), .B(n21248), .Z(n21142) );
  NAND U21594 ( .A(A[0]), .B(B[140]), .Z(n21248) );
  NAND U21595 ( .A(B[139]), .B(A[1]), .Z(n21145) );
  NAND U21596 ( .A(n21249), .B(n21250), .Z(n475) );
  NANDN U21597 ( .A(n21251), .B(n21252), .Z(n21250) );
  OR U21598 ( .A(n21253), .B(n21254), .Z(n21252) );
  NAND U21599 ( .A(n21254), .B(n21253), .Z(n21249) );
  XOR U21600 ( .A(n477), .B(n476), .Z(\A1[137] ) );
  XOR U21601 ( .A(n21254), .B(n21255), .Z(n476) );
  XNOR U21602 ( .A(n21253), .B(n21251), .Z(n21255) );
  AND U21603 ( .A(n21256), .B(n21257), .Z(n21251) );
  NANDN U21604 ( .A(n21258), .B(n21259), .Z(n21257) );
  NANDN U21605 ( .A(n21260), .B(n21261), .Z(n21259) );
  NANDN U21606 ( .A(n21261), .B(n21260), .Z(n21256) );
  ANDN U21607 ( .B(B[124]), .A(n29), .Z(n21253) );
  XNOR U21608 ( .A(n21160), .B(n21262), .Z(n21254) );
  XNOR U21609 ( .A(n21159), .B(n21157), .Z(n21262) );
  AND U21610 ( .A(n21263), .B(n21264), .Z(n21157) );
  NANDN U21611 ( .A(n21265), .B(n21266), .Z(n21264) );
  OR U21612 ( .A(n21267), .B(n21268), .Z(n21266) );
  NAND U21613 ( .A(n21268), .B(n21267), .Z(n21263) );
  ANDN U21614 ( .B(B[125]), .A(n30), .Z(n21159) );
  XNOR U21615 ( .A(n21167), .B(n21269), .Z(n21160) );
  XNOR U21616 ( .A(n21166), .B(n21164), .Z(n21269) );
  AND U21617 ( .A(n21270), .B(n21271), .Z(n21164) );
  NANDN U21618 ( .A(n21272), .B(n21273), .Z(n21271) );
  NANDN U21619 ( .A(n21274), .B(n21275), .Z(n21273) );
  NANDN U21620 ( .A(n21275), .B(n21274), .Z(n21270) );
  ANDN U21621 ( .B(B[126]), .A(n31), .Z(n21166) );
  XNOR U21622 ( .A(n21174), .B(n21276), .Z(n21167) );
  XNOR U21623 ( .A(n21173), .B(n21171), .Z(n21276) );
  AND U21624 ( .A(n21277), .B(n21278), .Z(n21171) );
  NANDN U21625 ( .A(n21279), .B(n21280), .Z(n21278) );
  OR U21626 ( .A(n21281), .B(n21282), .Z(n21280) );
  NAND U21627 ( .A(n21282), .B(n21281), .Z(n21277) );
  ANDN U21628 ( .B(B[127]), .A(n32), .Z(n21173) );
  XNOR U21629 ( .A(n21181), .B(n21283), .Z(n21174) );
  XNOR U21630 ( .A(n21180), .B(n21178), .Z(n21283) );
  AND U21631 ( .A(n21284), .B(n21285), .Z(n21178) );
  NANDN U21632 ( .A(n21286), .B(n21287), .Z(n21285) );
  NANDN U21633 ( .A(n21288), .B(n21289), .Z(n21287) );
  NANDN U21634 ( .A(n21289), .B(n21288), .Z(n21284) );
  ANDN U21635 ( .B(B[128]), .A(n33), .Z(n21180) );
  XNOR U21636 ( .A(n21188), .B(n21290), .Z(n21181) );
  XNOR U21637 ( .A(n21187), .B(n21185), .Z(n21290) );
  AND U21638 ( .A(n21291), .B(n21292), .Z(n21185) );
  NANDN U21639 ( .A(n21293), .B(n21294), .Z(n21292) );
  OR U21640 ( .A(n21295), .B(n21296), .Z(n21294) );
  NAND U21641 ( .A(n21296), .B(n21295), .Z(n21291) );
  ANDN U21642 ( .B(B[129]), .A(n34), .Z(n21187) );
  XNOR U21643 ( .A(n21195), .B(n21297), .Z(n21188) );
  XNOR U21644 ( .A(n21194), .B(n21192), .Z(n21297) );
  AND U21645 ( .A(n21298), .B(n21299), .Z(n21192) );
  NANDN U21646 ( .A(n21300), .B(n21301), .Z(n21299) );
  NANDN U21647 ( .A(n21302), .B(n21303), .Z(n21301) );
  NANDN U21648 ( .A(n21303), .B(n21302), .Z(n21298) );
  ANDN U21649 ( .B(B[130]), .A(n35), .Z(n21194) );
  XNOR U21650 ( .A(n21202), .B(n21304), .Z(n21195) );
  XNOR U21651 ( .A(n21201), .B(n21199), .Z(n21304) );
  AND U21652 ( .A(n21305), .B(n21306), .Z(n21199) );
  NANDN U21653 ( .A(n21307), .B(n21308), .Z(n21306) );
  OR U21654 ( .A(n21309), .B(n21310), .Z(n21308) );
  NAND U21655 ( .A(n21310), .B(n21309), .Z(n21305) );
  ANDN U21656 ( .B(B[131]), .A(n36), .Z(n21201) );
  XNOR U21657 ( .A(n21209), .B(n21311), .Z(n21202) );
  XNOR U21658 ( .A(n21208), .B(n21206), .Z(n21311) );
  AND U21659 ( .A(n21312), .B(n21313), .Z(n21206) );
  NANDN U21660 ( .A(n21314), .B(n21315), .Z(n21313) );
  NANDN U21661 ( .A(n21316), .B(n21317), .Z(n21315) );
  NANDN U21662 ( .A(n21317), .B(n21316), .Z(n21312) );
  ANDN U21663 ( .B(B[132]), .A(n37), .Z(n21208) );
  XNOR U21664 ( .A(n21216), .B(n21318), .Z(n21209) );
  XNOR U21665 ( .A(n21215), .B(n21213), .Z(n21318) );
  AND U21666 ( .A(n21319), .B(n21320), .Z(n21213) );
  NANDN U21667 ( .A(n21321), .B(n21322), .Z(n21320) );
  OR U21668 ( .A(n21323), .B(n21324), .Z(n21322) );
  NAND U21669 ( .A(n21324), .B(n21323), .Z(n21319) );
  ANDN U21670 ( .B(B[133]), .A(n38), .Z(n21215) );
  XNOR U21671 ( .A(n21223), .B(n21325), .Z(n21216) );
  XNOR U21672 ( .A(n21222), .B(n21220), .Z(n21325) );
  AND U21673 ( .A(n21326), .B(n21327), .Z(n21220) );
  NANDN U21674 ( .A(n21328), .B(n21329), .Z(n21327) );
  NANDN U21675 ( .A(n21330), .B(n21331), .Z(n21329) );
  NANDN U21676 ( .A(n21331), .B(n21330), .Z(n21326) );
  ANDN U21677 ( .B(B[134]), .A(n39), .Z(n21222) );
  XNOR U21678 ( .A(n21230), .B(n21332), .Z(n21223) );
  XNOR U21679 ( .A(n21229), .B(n21227), .Z(n21332) );
  AND U21680 ( .A(n21333), .B(n21334), .Z(n21227) );
  NANDN U21681 ( .A(n21335), .B(n21336), .Z(n21334) );
  OR U21682 ( .A(n21337), .B(n21338), .Z(n21336) );
  NAND U21683 ( .A(n21338), .B(n21337), .Z(n21333) );
  ANDN U21684 ( .B(B[135]), .A(n40), .Z(n21229) );
  XNOR U21685 ( .A(n21237), .B(n21339), .Z(n21230) );
  XNOR U21686 ( .A(n21236), .B(n21234), .Z(n21339) );
  AND U21687 ( .A(n21340), .B(n21341), .Z(n21234) );
  NANDN U21688 ( .A(n21342), .B(n21343), .Z(n21341) );
  NAND U21689 ( .A(n21344), .B(n21345), .Z(n21343) );
  ANDN U21690 ( .B(B[136]), .A(n41), .Z(n21236) );
  XOR U21691 ( .A(n21243), .B(n21346), .Z(n21237) );
  XNOR U21692 ( .A(n21241), .B(n21244), .Z(n21346) );
  NAND U21693 ( .A(A[2]), .B(B[137]), .Z(n21244) );
  NANDN U21694 ( .A(n21347), .B(n21348), .Z(n21241) );
  AND U21695 ( .A(A[0]), .B(B[138]), .Z(n21348) );
  XNOR U21696 ( .A(n21246), .B(n21349), .Z(n21243) );
  NAND U21697 ( .A(A[0]), .B(B[139]), .Z(n21349) );
  NAND U21698 ( .A(B[138]), .B(A[1]), .Z(n21246) );
  NAND U21699 ( .A(n21350), .B(n21351), .Z(n477) );
  NANDN U21700 ( .A(n21352), .B(n21353), .Z(n21351) );
  OR U21701 ( .A(n21354), .B(n21355), .Z(n21353) );
  NAND U21702 ( .A(n21355), .B(n21354), .Z(n21350) );
  XOR U21703 ( .A(n479), .B(n478), .Z(\A1[136] ) );
  XOR U21704 ( .A(n21355), .B(n21356), .Z(n478) );
  XNOR U21705 ( .A(n21354), .B(n21352), .Z(n21356) );
  AND U21706 ( .A(n21357), .B(n21358), .Z(n21352) );
  NANDN U21707 ( .A(n21359), .B(n21360), .Z(n21358) );
  NANDN U21708 ( .A(n21361), .B(n21362), .Z(n21360) );
  NANDN U21709 ( .A(n21362), .B(n21361), .Z(n21357) );
  ANDN U21710 ( .B(B[123]), .A(n29), .Z(n21354) );
  XNOR U21711 ( .A(n21261), .B(n21363), .Z(n21355) );
  XNOR U21712 ( .A(n21260), .B(n21258), .Z(n21363) );
  AND U21713 ( .A(n21364), .B(n21365), .Z(n21258) );
  NANDN U21714 ( .A(n21366), .B(n21367), .Z(n21365) );
  OR U21715 ( .A(n21368), .B(n21369), .Z(n21367) );
  NAND U21716 ( .A(n21369), .B(n21368), .Z(n21364) );
  ANDN U21717 ( .B(B[124]), .A(n30), .Z(n21260) );
  XNOR U21718 ( .A(n21268), .B(n21370), .Z(n21261) );
  XNOR U21719 ( .A(n21267), .B(n21265), .Z(n21370) );
  AND U21720 ( .A(n21371), .B(n21372), .Z(n21265) );
  NANDN U21721 ( .A(n21373), .B(n21374), .Z(n21372) );
  NANDN U21722 ( .A(n21375), .B(n21376), .Z(n21374) );
  NANDN U21723 ( .A(n21376), .B(n21375), .Z(n21371) );
  ANDN U21724 ( .B(B[125]), .A(n31), .Z(n21267) );
  XNOR U21725 ( .A(n21275), .B(n21377), .Z(n21268) );
  XNOR U21726 ( .A(n21274), .B(n21272), .Z(n21377) );
  AND U21727 ( .A(n21378), .B(n21379), .Z(n21272) );
  NANDN U21728 ( .A(n21380), .B(n21381), .Z(n21379) );
  OR U21729 ( .A(n21382), .B(n21383), .Z(n21381) );
  NAND U21730 ( .A(n21383), .B(n21382), .Z(n21378) );
  ANDN U21731 ( .B(B[126]), .A(n32), .Z(n21274) );
  XNOR U21732 ( .A(n21282), .B(n21384), .Z(n21275) );
  XNOR U21733 ( .A(n21281), .B(n21279), .Z(n21384) );
  AND U21734 ( .A(n21385), .B(n21386), .Z(n21279) );
  NANDN U21735 ( .A(n21387), .B(n21388), .Z(n21386) );
  NANDN U21736 ( .A(n21389), .B(n21390), .Z(n21388) );
  NANDN U21737 ( .A(n21390), .B(n21389), .Z(n21385) );
  ANDN U21738 ( .B(B[127]), .A(n33), .Z(n21281) );
  XNOR U21739 ( .A(n21289), .B(n21391), .Z(n21282) );
  XNOR U21740 ( .A(n21288), .B(n21286), .Z(n21391) );
  AND U21741 ( .A(n21392), .B(n21393), .Z(n21286) );
  NANDN U21742 ( .A(n21394), .B(n21395), .Z(n21393) );
  OR U21743 ( .A(n21396), .B(n21397), .Z(n21395) );
  NAND U21744 ( .A(n21397), .B(n21396), .Z(n21392) );
  ANDN U21745 ( .B(B[128]), .A(n34), .Z(n21288) );
  XNOR U21746 ( .A(n21296), .B(n21398), .Z(n21289) );
  XNOR U21747 ( .A(n21295), .B(n21293), .Z(n21398) );
  AND U21748 ( .A(n21399), .B(n21400), .Z(n21293) );
  NANDN U21749 ( .A(n21401), .B(n21402), .Z(n21400) );
  NANDN U21750 ( .A(n21403), .B(n21404), .Z(n21402) );
  NANDN U21751 ( .A(n21404), .B(n21403), .Z(n21399) );
  ANDN U21752 ( .B(B[129]), .A(n35), .Z(n21295) );
  XNOR U21753 ( .A(n21303), .B(n21405), .Z(n21296) );
  XNOR U21754 ( .A(n21302), .B(n21300), .Z(n21405) );
  AND U21755 ( .A(n21406), .B(n21407), .Z(n21300) );
  NANDN U21756 ( .A(n21408), .B(n21409), .Z(n21407) );
  OR U21757 ( .A(n21410), .B(n21411), .Z(n21409) );
  NAND U21758 ( .A(n21411), .B(n21410), .Z(n21406) );
  ANDN U21759 ( .B(B[130]), .A(n36), .Z(n21302) );
  XNOR U21760 ( .A(n21310), .B(n21412), .Z(n21303) );
  XNOR U21761 ( .A(n21309), .B(n21307), .Z(n21412) );
  AND U21762 ( .A(n21413), .B(n21414), .Z(n21307) );
  NANDN U21763 ( .A(n21415), .B(n21416), .Z(n21414) );
  NANDN U21764 ( .A(n21417), .B(n21418), .Z(n21416) );
  NANDN U21765 ( .A(n21418), .B(n21417), .Z(n21413) );
  ANDN U21766 ( .B(B[131]), .A(n37), .Z(n21309) );
  XNOR U21767 ( .A(n21317), .B(n21419), .Z(n21310) );
  XNOR U21768 ( .A(n21316), .B(n21314), .Z(n21419) );
  AND U21769 ( .A(n21420), .B(n21421), .Z(n21314) );
  NANDN U21770 ( .A(n21422), .B(n21423), .Z(n21421) );
  OR U21771 ( .A(n21424), .B(n21425), .Z(n21423) );
  NAND U21772 ( .A(n21425), .B(n21424), .Z(n21420) );
  ANDN U21773 ( .B(B[132]), .A(n38), .Z(n21316) );
  XNOR U21774 ( .A(n21324), .B(n21426), .Z(n21317) );
  XNOR U21775 ( .A(n21323), .B(n21321), .Z(n21426) );
  AND U21776 ( .A(n21427), .B(n21428), .Z(n21321) );
  NANDN U21777 ( .A(n21429), .B(n21430), .Z(n21428) );
  NANDN U21778 ( .A(n21431), .B(n21432), .Z(n21430) );
  NANDN U21779 ( .A(n21432), .B(n21431), .Z(n21427) );
  ANDN U21780 ( .B(B[133]), .A(n39), .Z(n21323) );
  XNOR U21781 ( .A(n21331), .B(n21433), .Z(n21324) );
  XNOR U21782 ( .A(n21330), .B(n21328), .Z(n21433) );
  AND U21783 ( .A(n21434), .B(n21435), .Z(n21328) );
  NANDN U21784 ( .A(n21436), .B(n21437), .Z(n21435) );
  OR U21785 ( .A(n21438), .B(n21439), .Z(n21437) );
  NAND U21786 ( .A(n21439), .B(n21438), .Z(n21434) );
  ANDN U21787 ( .B(B[134]), .A(n40), .Z(n21330) );
  XNOR U21788 ( .A(n21338), .B(n21440), .Z(n21331) );
  XNOR U21789 ( .A(n21337), .B(n21335), .Z(n21440) );
  AND U21790 ( .A(n21441), .B(n21442), .Z(n21335) );
  NANDN U21791 ( .A(n21443), .B(n21444), .Z(n21442) );
  NAND U21792 ( .A(n21445), .B(n21446), .Z(n21444) );
  ANDN U21793 ( .B(B[135]), .A(n41), .Z(n21337) );
  XOR U21794 ( .A(n21344), .B(n21447), .Z(n21338) );
  XNOR U21795 ( .A(n21342), .B(n21345), .Z(n21447) );
  NAND U21796 ( .A(A[2]), .B(B[136]), .Z(n21345) );
  NANDN U21797 ( .A(n21448), .B(n21449), .Z(n21342) );
  AND U21798 ( .A(A[0]), .B(B[137]), .Z(n21449) );
  XNOR U21799 ( .A(n21347), .B(n21450), .Z(n21344) );
  NAND U21800 ( .A(A[0]), .B(B[138]), .Z(n21450) );
  NAND U21801 ( .A(B[137]), .B(A[1]), .Z(n21347) );
  NAND U21802 ( .A(n21451), .B(n21452), .Z(n479) );
  NANDN U21803 ( .A(n21453), .B(n21454), .Z(n21452) );
  OR U21804 ( .A(n21455), .B(n21456), .Z(n21454) );
  NAND U21805 ( .A(n21456), .B(n21455), .Z(n21451) );
  XOR U21806 ( .A(n481), .B(n480), .Z(\A1[135] ) );
  XOR U21807 ( .A(n21456), .B(n21457), .Z(n480) );
  XNOR U21808 ( .A(n21455), .B(n21453), .Z(n21457) );
  AND U21809 ( .A(n21458), .B(n21459), .Z(n21453) );
  NANDN U21810 ( .A(n21460), .B(n21461), .Z(n21459) );
  NANDN U21811 ( .A(n21462), .B(n21463), .Z(n21461) );
  NANDN U21812 ( .A(n21463), .B(n21462), .Z(n21458) );
  ANDN U21813 ( .B(B[122]), .A(n29), .Z(n21455) );
  XNOR U21814 ( .A(n21362), .B(n21464), .Z(n21456) );
  XNOR U21815 ( .A(n21361), .B(n21359), .Z(n21464) );
  AND U21816 ( .A(n21465), .B(n21466), .Z(n21359) );
  NANDN U21817 ( .A(n21467), .B(n21468), .Z(n21466) );
  OR U21818 ( .A(n21469), .B(n21470), .Z(n21468) );
  NAND U21819 ( .A(n21470), .B(n21469), .Z(n21465) );
  ANDN U21820 ( .B(B[123]), .A(n30), .Z(n21361) );
  XNOR U21821 ( .A(n21369), .B(n21471), .Z(n21362) );
  XNOR U21822 ( .A(n21368), .B(n21366), .Z(n21471) );
  AND U21823 ( .A(n21472), .B(n21473), .Z(n21366) );
  NANDN U21824 ( .A(n21474), .B(n21475), .Z(n21473) );
  NANDN U21825 ( .A(n21476), .B(n21477), .Z(n21475) );
  NANDN U21826 ( .A(n21477), .B(n21476), .Z(n21472) );
  ANDN U21827 ( .B(B[124]), .A(n31), .Z(n21368) );
  XNOR U21828 ( .A(n21376), .B(n21478), .Z(n21369) );
  XNOR U21829 ( .A(n21375), .B(n21373), .Z(n21478) );
  AND U21830 ( .A(n21479), .B(n21480), .Z(n21373) );
  NANDN U21831 ( .A(n21481), .B(n21482), .Z(n21480) );
  OR U21832 ( .A(n21483), .B(n21484), .Z(n21482) );
  NAND U21833 ( .A(n21484), .B(n21483), .Z(n21479) );
  ANDN U21834 ( .B(B[125]), .A(n32), .Z(n21375) );
  XNOR U21835 ( .A(n21383), .B(n21485), .Z(n21376) );
  XNOR U21836 ( .A(n21382), .B(n21380), .Z(n21485) );
  AND U21837 ( .A(n21486), .B(n21487), .Z(n21380) );
  NANDN U21838 ( .A(n21488), .B(n21489), .Z(n21487) );
  NANDN U21839 ( .A(n21490), .B(n21491), .Z(n21489) );
  NANDN U21840 ( .A(n21491), .B(n21490), .Z(n21486) );
  ANDN U21841 ( .B(B[126]), .A(n33), .Z(n21382) );
  XNOR U21842 ( .A(n21390), .B(n21492), .Z(n21383) );
  XNOR U21843 ( .A(n21389), .B(n21387), .Z(n21492) );
  AND U21844 ( .A(n21493), .B(n21494), .Z(n21387) );
  NANDN U21845 ( .A(n21495), .B(n21496), .Z(n21494) );
  OR U21846 ( .A(n21497), .B(n21498), .Z(n21496) );
  NAND U21847 ( .A(n21498), .B(n21497), .Z(n21493) );
  ANDN U21848 ( .B(B[127]), .A(n34), .Z(n21389) );
  XNOR U21849 ( .A(n21397), .B(n21499), .Z(n21390) );
  XNOR U21850 ( .A(n21396), .B(n21394), .Z(n21499) );
  AND U21851 ( .A(n21500), .B(n21501), .Z(n21394) );
  NANDN U21852 ( .A(n21502), .B(n21503), .Z(n21501) );
  NANDN U21853 ( .A(n21504), .B(n21505), .Z(n21503) );
  NANDN U21854 ( .A(n21505), .B(n21504), .Z(n21500) );
  ANDN U21855 ( .B(B[128]), .A(n35), .Z(n21396) );
  XNOR U21856 ( .A(n21404), .B(n21506), .Z(n21397) );
  XNOR U21857 ( .A(n21403), .B(n21401), .Z(n21506) );
  AND U21858 ( .A(n21507), .B(n21508), .Z(n21401) );
  NANDN U21859 ( .A(n21509), .B(n21510), .Z(n21508) );
  OR U21860 ( .A(n21511), .B(n21512), .Z(n21510) );
  NAND U21861 ( .A(n21512), .B(n21511), .Z(n21507) );
  ANDN U21862 ( .B(B[129]), .A(n36), .Z(n21403) );
  XNOR U21863 ( .A(n21411), .B(n21513), .Z(n21404) );
  XNOR U21864 ( .A(n21410), .B(n21408), .Z(n21513) );
  AND U21865 ( .A(n21514), .B(n21515), .Z(n21408) );
  NANDN U21866 ( .A(n21516), .B(n21517), .Z(n21515) );
  NANDN U21867 ( .A(n21518), .B(n21519), .Z(n21517) );
  NANDN U21868 ( .A(n21519), .B(n21518), .Z(n21514) );
  ANDN U21869 ( .B(B[130]), .A(n37), .Z(n21410) );
  XNOR U21870 ( .A(n21418), .B(n21520), .Z(n21411) );
  XNOR U21871 ( .A(n21417), .B(n21415), .Z(n21520) );
  AND U21872 ( .A(n21521), .B(n21522), .Z(n21415) );
  NANDN U21873 ( .A(n21523), .B(n21524), .Z(n21522) );
  OR U21874 ( .A(n21525), .B(n21526), .Z(n21524) );
  NAND U21875 ( .A(n21526), .B(n21525), .Z(n21521) );
  ANDN U21876 ( .B(B[131]), .A(n38), .Z(n21417) );
  XNOR U21877 ( .A(n21425), .B(n21527), .Z(n21418) );
  XNOR U21878 ( .A(n21424), .B(n21422), .Z(n21527) );
  AND U21879 ( .A(n21528), .B(n21529), .Z(n21422) );
  NANDN U21880 ( .A(n21530), .B(n21531), .Z(n21529) );
  NANDN U21881 ( .A(n21532), .B(n21533), .Z(n21531) );
  NANDN U21882 ( .A(n21533), .B(n21532), .Z(n21528) );
  ANDN U21883 ( .B(B[132]), .A(n39), .Z(n21424) );
  XNOR U21884 ( .A(n21432), .B(n21534), .Z(n21425) );
  XNOR U21885 ( .A(n21431), .B(n21429), .Z(n21534) );
  AND U21886 ( .A(n21535), .B(n21536), .Z(n21429) );
  NANDN U21887 ( .A(n21537), .B(n21538), .Z(n21536) );
  OR U21888 ( .A(n21539), .B(n21540), .Z(n21538) );
  NAND U21889 ( .A(n21540), .B(n21539), .Z(n21535) );
  ANDN U21890 ( .B(B[133]), .A(n40), .Z(n21431) );
  XNOR U21891 ( .A(n21439), .B(n21541), .Z(n21432) );
  XNOR U21892 ( .A(n21438), .B(n21436), .Z(n21541) );
  AND U21893 ( .A(n21542), .B(n21543), .Z(n21436) );
  NANDN U21894 ( .A(n21544), .B(n21545), .Z(n21543) );
  NAND U21895 ( .A(n21546), .B(n21547), .Z(n21545) );
  ANDN U21896 ( .B(B[134]), .A(n41), .Z(n21438) );
  XOR U21897 ( .A(n21445), .B(n21548), .Z(n21439) );
  XNOR U21898 ( .A(n21443), .B(n21446), .Z(n21548) );
  NAND U21899 ( .A(A[2]), .B(B[135]), .Z(n21446) );
  NANDN U21900 ( .A(n21549), .B(n21550), .Z(n21443) );
  AND U21901 ( .A(A[0]), .B(B[136]), .Z(n21550) );
  XNOR U21902 ( .A(n21448), .B(n21551), .Z(n21445) );
  NAND U21903 ( .A(A[0]), .B(B[137]), .Z(n21551) );
  NAND U21904 ( .A(B[136]), .B(A[1]), .Z(n21448) );
  NAND U21905 ( .A(n21552), .B(n21553), .Z(n481) );
  NANDN U21906 ( .A(n21554), .B(n21555), .Z(n21553) );
  OR U21907 ( .A(n21556), .B(n21557), .Z(n21555) );
  NAND U21908 ( .A(n21557), .B(n21556), .Z(n21552) );
  XOR U21909 ( .A(n483), .B(n482), .Z(\A1[134] ) );
  XOR U21910 ( .A(n21557), .B(n21558), .Z(n482) );
  XNOR U21911 ( .A(n21556), .B(n21554), .Z(n21558) );
  AND U21912 ( .A(n21559), .B(n21560), .Z(n21554) );
  NANDN U21913 ( .A(n21561), .B(n21562), .Z(n21560) );
  NANDN U21914 ( .A(n21563), .B(n21564), .Z(n21562) );
  NANDN U21915 ( .A(n21564), .B(n21563), .Z(n21559) );
  ANDN U21916 ( .B(B[121]), .A(n29), .Z(n21556) );
  XNOR U21917 ( .A(n21463), .B(n21565), .Z(n21557) );
  XNOR U21918 ( .A(n21462), .B(n21460), .Z(n21565) );
  AND U21919 ( .A(n21566), .B(n21567), .Z(n21460) );
  NANDN U21920 ( .A(n21568), .B(n21569), .Z(n21567) );
  OR U21921 ( .A(n21570), .B(n21571), .Z(n21569) );
  NAND U21922 ( .A(n21571), .B(n21570), .Z(n21566) );
  ANDN U21923 ( .B(B[122]), .A(n30), .Z(n21462) );
  XNOR U21924 ( .A(n21470), .B(n21572), .Z(n21463) );
  XNOR U21925 ( .A(n21469), .B(n21467), .Z(n21572) );
  AND U21926 ( .A(n21573), .B(n21574), .Z(n21467) );
  NANDN U21927 ( .A(n21575), .B(n21576), .Z(n21574) );
  NANDN U21928 ( .A(n21577), .B(n21578), .Z(n21576) );
  NANDN U21929 ( .A(n21578), .B(n21577), .Z(n21573) );
  ANDN U21930 ( .B(B[123]), .A(n31), .Z(n21469) );
  XNOR U21931 ( .A(n21477), .B(n21579), .Z(n21470) );
  XNOR U21932 ( .A(n21476), .B(n21474), .Z(n21579) );
  AND U21933 ( .A(n21580), .B(n21581), .Z(n21474) );
  NANDN U21934 ( .A(n21582), .B(n21583), .Z(n21581) );
  OR U21935 ( .A(n21584), .B(n21585), .Z(n21583) );
  NAND U21936 ( .A(n21585), .B(n21584), .Z(n21580) );
  ANDN U21937 ( .B(B[124]), .A(n32), .Z(n21476) );
  XNOR U21938 ( .A(n21484), .B(n21586), .Z(n21477) );
  XNOR U21939 ( .A(n21483), .B(n21481), .Z(n21586) );
  AND U21940 ( .A(n21587), .B(n21588), .Z(n21481) );
  NANDN U21941 ( .A(n21589), .B(n21590), .Z(n21588) );
  NANDN U21942 ( .A(n21591), .B(n21592), .Z(n21590) );
  NANDN U21943 ( .A(n21592), .B(n21591), .Z(n21587) );
  ANDN U21944 ( .B(B[125]), .A(n33), .Z(n21483) );
  XNOR U21945 ( .A(n21491), .B(n21593), .Z(n21484) );
  XNOR U21946 ( .A(n21490), .B(n21488), .Z(n21593) );
  AND U21947 ( .A(n21594), .B(n21595), .Z(n21488) );
  NANDN U21948 ( .A(n21596), .B(n21597), .Z(n21595) );
  OR U21949 ( .A(n21598), .B(n21599), .Z(n21597) );
  NAND U21950 ( .A(n21599), .B(n21598), .Z(n21594) );
  ANDN U21951 ( .B(B[126]), .A(n34), .Z(n21490) );
  XNOR U21952 ( .A(n21498), .B(n21600), .Z(n21491) );
  XNOR U21953 ( .A(n21497), .B(n21495), .Z(n21600) );
  AND U21954 ( .A(n21601), .B(n21602), .Z(n21495) );
  NANDN U21955 ( .A(n21603), .B(n21604), .Z(n21602) );
  NANDN U21956 ( .A(n21605), .B(n21606), .Z(n21604) );
  NANDN U21957 ( .A(n21606), .B(n21605), .Z(n21601) );
  ANDN U21958 ( .B(B[127]), .A(n35), .Z(n21497) );
  XNOR U21959 ( .A(n21505), .B(n21607), .Z(n21498) );
  XNOR U21960 ( .A(n21504), .B(n21502), .Z(n21607) );
  AND U21961 ( .A(n21608), .B(n21609), .Z(n21502) );
  NANDN U21962 ( .A(n21610), .B(n21611), .Z(n21609) );
  OR U21963 ( .A(n21612), .B(n21613), .Z(n21611) );
  NAND U21964 ( .A(n21613), .B(n21612), .Z(n21608) );
  ANDN U21965 ( .B(B[128]), .A(n36), .Z(n21504) );
  XNOR U21966 ( .A(n21512), .B(n21614), .Z(n21505) );
  XNOR U21967 ( .A(n21511), .B(n21509), .Z(n21614) );
  AND U21968 ( .A(n21615), .B(n21616), .Z(n21509) );
  NANDN U21969 ( .A(n21617), .B(n21618), .Z(n21616) );
  NANDN U21970 ( .A(n21619), .B(n21620), .Z(n21618) );
  NANDN U21971 ( .A(n21620), .B(n21619), .Z(n21615) );
  ANDN U21972 ( .B(B[129]), .A(n37), .Z(n21511) );
  XNOR U21973 ( .A(n21519), .B(n21621), .Z(n21512) );
  XNOR U21974 ( .A(n21518), .B(n21516), .Z(n21621) );
  AND U21975 ( .A(n21622), .B(n21623), .Z(n21516) );
  NANDN U21976 ( .A(n21624), .B(n21625), .Z(n21623) );
  OR U21977 ( .A(n21626), .B(n21627), .Z(n21625) );
  NAND U21978 ( .A(n21627), .B(n21626), .Z(n21622) );
  ANDN U21979 ( .B(B[130]), .A(n38), .Z(n21518) );
  XNOR U21980 ( .A(n21526), .B(n21628), .Z(n21519) );
  XNOR U21981 ( .A(n21525), .B(n21523), .Z(n21628) );
  AND U21982 ( .A(n21629), .B(n21630), .Z(n21523) );
  NANDN U21983 ( .A(n21631), .B(n21632), .Z(n21630) );
  NANDN U21984 ( .A(n21633), .B(n21634), .Z(n21632) );
  NANDN U21985 ( .A(n21634), .B(n21633), .Z(n21629) );
  ANDN U21986 ( .B(B[131]), .A(n39), .Z(n21525) );
  XNOR U21987 ( .A(n21533), .B(n21635), .Z(n21526) );
  XNOR U21988 ( .A(n21532), .B(n21530), .Z(n21635) );
  AND U21989 ( .A(n21636), .B(n21637), .Z(n21530) );
  NANDN U21990 ( .A(n21638), .B(n21639), .Z(n21637) );
  OR U21991 ( .A(n21640), .B(n21641), .Z(n21639) );
  NAND U21992 ( .A(n21641), .B(n21640), .Z(n21636) );
  ANDN U21993 ( .B(B[132]), .A(n40), .Z(n21532) );
  XNOR U21994 ( .A(n21540), .B(n21642), .Z(n21533) );
  XNOR U21995 ( .A(n21539), .B(n21537), .Z(n21642) );
  AND U21996 ( .A(n21643), .B(n21644), .Z(n21537) );
  NANDN U21997 ( .A(n21645), .B(n21646), .Z(n21644) );
  NAND U21998 ( .A(n21647), .B(n21648), .Z(n21646) );
  ANDN U21999 ( .B(B[133]), .A(n41), .Z(n21539) );
  XOR U22000 ( .A(n21546), .B(n21649), .Z(n21540) );
  XNOR U22001 ( .A(n21544), .B(n21547), .Z(n21649) );
  NAND U22002 ( .A(A[2]), .B(B[134]), .Z(n21547) );
  NANDN U22003 ( .A(n21650), .B(n21651), .Z(n21544) );
  AND U22004 ( .A(A[0]), .B(B[135]), .Z(n21651) );
  XNOR U22005 ( .A(n21549), .B(n21652), .Z(n21546) );
  NAND U22006 ( .A(A[0]), .B(B[136]), .Z(n21652) );
  NAND U22007 ( .A(B[135]), .B(A[1]), .Z(n21549) );
  NAND U22008 ( .A(n21653), .B(n21654), .Z(n483) );
  NANDN U22009 ( .A(n21655), .B(n21656), .Z(n21654) );
  OR U22010 ( .A(n21657), .B(n21658), .Z(n21656) );
  NAND U22011 ( .A(n21658), .B(n21657), .Z(n21653) );
  XOR U22012 ( .A(n485), .B(n484), .Z(\A1[133] ) );
  XOR U22013 ( .A(n21658), .B(n21659), .Z(n484) );
  XNOR U22014 ( .A(n21657), .B(n21655), .Z(n21659) );
  AND U22015 ( .A(n21660), .B(n21661), .Z(n21655) );
  NANDN U22016 ( .A(n21662), .B(n21663), .Z(n21661) );
  NANDN U22017 ( .A(n21664), .B(n21665), .Z(n21663) );
  NANDN U22018 ( .A(n21665), .B(n21664), .Z(n21660) );
  ANDN U22019 ( .B(B[120]), .A(n29), .Z(n21657) );
  XNOR U22020 ( .A(n21564), .B(n21666), .Z(n21658) );
  XNOR U22021 ( .A(n21563), .B(n21561), .Z(n21666) );
  AND U22022 ( .A(n21667), .B(n21668), .Z(n21561) );
  NANDN U22023 ( .A(n21669), .B(n21670), .Z(n21668) );
  OR U22024 ( .A(n21671), .B(n21672), .Z(n21670) );
  NAND U22025 ( .A(n21672), .B(n21671), .Z(n21667) );
  ANDN U22026 ( .B(B[121]), .A(n30), .Z(n21563) );
  XNOR U22027 ( .A(n21571), .B(n21673), .Z(n21564) );
  XNOR U22028 ( .A(n21570), .B(n21568), .Z(n21673) );
  AND U22029 ( .A(n21674), .B(n21675), .Z(n21568) );
  NANDN U22030 ( .A(n21676), .B(n21677), .Z(n21675) );
  NANDN U22031 ( .A(n21678), .B(n21679), .Z(n21677) );
  NANDN U22032 ( .A(n21679), .B(n21678), .Z(n21674) );
  ANDN U22033 ( .B(B[122]), .A(n31), .Z(n21570) );
  XNOR U22034 ( .A(n21578), .B(n21680), .Z(n21571) );
  XNOR U22035 ( .A(n21577), .B(n21575), .Z(n21680) );
  AND U22036 ( .A(n21681), .B(n21682), .Z(n21575) );
  NANDN U22037 ( .A(n21683), .B(n21684), .Z(n21682) );
  OR U22038 ( .A(n21685), .B(n21686), .Z(n21684) );
  NAND U22039 ( .A(n21686), .B(n21685), .Z(n21681) );
  ANDN U22040 ( .B(B[123]), .A(n32), .Z(n21577) );
  XNOR U22041 ( .A(n21585), .B(n21687), .Z(n21578) );
  XNOR U22042 ( .A(n21584), .B(n21582), .Z(n21687) );
  AND U22043 ( .A(n21688), .B(n21689), .Z(n21582) );
  NANDN U22044 ( .A(n21690), .B(n21691), .Z(n21689) );
  NANDN U22045 ( .A(n21692), .B(n21693), .Z(n21691) );
  NANDN U22046 ( .A(n21693), .B(n21692), .Z(n21688) );
  ANDN U22047 ( .B(B[124]), .A(n33), .Z(n21584) );
  XNOR U22048 ( .A(n21592), .B(n21694), .Z(n21585) );
  XNOR U22049 ( .A(n21591), .B(n21589), .Z(n21694) );
  AND U22050 ( .A(n21695), .B(n21696), .Z(n21589) );
  NANDN U22051 ( .A(n21697), .B(n21698), .Z(n21696) );
  OR U22052 ( .A(n21699), .B(n21700), .Z(n21698) );
  NAND U22053 ( .A(n21700), .B(n21699), .Z(n21695) );
  ANDN U22054 ( .B(B[125]), .A(n34), .Z(n21591) );
  XNOR U22055 ( .A(n21599), .B(n21701), .Z(n21592) );
  XNOR U22056 ( .A(n21598), .B(n21596), .Z(n21701) );
  AND U22057 ( .A(n21702), .B(n21703), .Z(n21596) );
  NANDN U22058 ( .A(n21704), .B(n21705), .Z(n21703) );
  NANDN U22059 ( .A(n21706), .B(n21707), .Z(n21705) );
  NANDN U22060 ( .A(n21707), .B(n21706), .Z(n21702) );
  ANDN U22061 ( .B(B[126]), .A(n35), .Z(n21598) );
  XNOR U22062 ( .A(n21606), .B(n21708), .Z(n21599) );
  XNOR U22063 ( .A(n21605), .B(n21603), .Z(n21708) );
  AND U22064 ( .A(n21709), .B(n21710), .Z(n21603) );
  NANDN U22065 ( .A(n21711), .B(n21712), .Z(n21710) );
  OR U22066 ( .A(n21713), .B(n21714), .Z(n21712) );
  NAND U22067 ( .A(n21714), .B(n21713), .Z(n21709) );
  ANDN U22068 ( .B(B[127]), .A(n36), .Z(n21605) );
  XNOR U22069 ( .A(n21613), .B(n21715), .Z(n21606) );
  XNOR U22070 ( .A(n21612), .B(n21610), .Z(n21715) );
  AND U22071 ( .A(n21716), .B(n21717), .Z(n21610) );
  NANDN U22072 ( .A(n21718), .B(n21719), .Z(n21717) );
  NANDN U22073 ( .A(n21720), .B(n21721), .Z(n21719) );
  NANDN U22074 ( .A(n21721), .B(n21720), .Z(n21716) );
  ANDN U22075 ( .B(B[128]), .A(n37), .Z(n21612) );
  XNOR U22076 ( .A(n21620), .B(n21722), .Z(n21613) );
  XNOR U22077 ( .A(n21619), .B(n21617), .Z(n21722) );
  AND U22078 ( .A(n21723), .B(n21724), .Z(n21617) );
  NANDN U22079 ( .A(n21725), .B(n21726), .Z(n21724) );
  OR U22080 ( .A(n21727), .B(n21728), .Z(n21726) );
  NAND U22081 ( .A(n21728), .B(n21727), .Z(n21723) );
  ANDN U22082 ( .B(B[129]), .A(n38), .Z(n21619) );
  XNOR U22083 ( .A(n21627), .B(n21729), .Z(n21620) );
  XNOR U22084 ( .A(n21626), .B(n21624), .Z(n21729) );
  AND U22085 ( .A(n21730), .B(n21731), .Z(n21624) );
  NANDN U22086 ( .A(n21732), .B(n21733), .Z(n21731) );
  NANDN U22087 ( .A(n21734), .B(n21735), .Z(n21733) );
  NANDN U22088 ( .A(n21735), .B(n21734), .Z(n21730) );
  ANDN U22089 ( .B(B[130]), .A(n39), .Z(n21626) );
  XNOR U22090 ( .A(n21634), .B(n21736), .Z(n21627) );
  XNOR U22091 ( .A(n21633), .B(n21631), .Z(n21736) );
  AND U22092 ( .A(n21737), .B(n21738), .Z(n21631) );
  NANDN U22093 ( .A(n21739), .B(n21740), .Z(n21738) );
  OR U22094 ( .A(n21741), .B(n21742), .Z(n21740) );
  NAND U22095 ( .A(n21742), .B(n21741), .Z(n21737) );
  ANDN U22096 ( .B(B[131]), .A(n40), .Z(n21633) );
  XNOR U22097 ( .A(n21641), .B(n21743), .Z(n21634) );
  XNOR U22098 ( .A(n21640), .B(n21638), .Z(n21743) );
  AND U22099 ( .A(n21744), .B(n21745), .Z(n21638) );
  NANDN U22100 ( .A(n21746), .B(n21747), .Z(n21745) );
  NAND U22101 ( .A(n21748), .B(n21749), .Z(n21747) );
  ANDN U22102 ( .B(B[132]), .A(n41), .Z(n21640) );
  XOR U22103 ( .A(n21647), .B(n21750), .Z(n21641) );
  XNOR U22104 ( .A(n21645), .B(n21648), .Z(n21750) );
  NAND U22105 ( .A(A[2]), .B(B[133]), .Z(n21648) );
  NANDN U22106 ( .A(n21751), .B(n21752), .Z(n21645) );
  AND U22107 ( .A(A[0]), .B(B[134]), .Z(n21752) );
  XNOR U22108 ( .A(n21650), .B(n21753), .Z(n21647) );
  NAND U22109 ( .A(A[0]), .B(B[135]), .Z(n21753) );
  NAND U22110 ( .A(B[134]), .B(A[1]), .Z(n21650) );
  NAND U22111 ( .A(n21754), .B(n21755), .Z(n485) );
  NANDN U22112 ( .A(n21756), .B(n21757), .Z(n21755) );
  OR U22113 ( .A(n21758), .B(n21759), .Z(n21757) );
  NAND U22114 ( .A(n21759), .B(n21758), .Z(n21754) );
  XOR U22115 ( .A(n487), .B(n486), .Z(\A1[132] ) );
  XOR U22116 ( .A(n21759), .B(n21760), .Z(n486) );
  XNOR U22117 ( .A(n21758), .B(n21756), .Z(n21760) );
  AND U22118 ( .A(n21761), .B(n21762), .Z(n21756) );
  NANDN U22119 ( .A(n21763), .B(n21764), .Z(n21762) );
  NANDN U22120 ( .A(n21765), .B(n21766), .Z(n21764) );
  NANDN U22121 ( .A(n21766), .B(n21765), .Z(n21761) );
  ANDN U22122 ( .B(B[119]), .A(n29), .Z(n21758) );
  XNOR U22123 ( .A(n21665), .B(n21767), .Z(n21759) );
  XNOR U22124 ( .A(n21664), .B(n21662), .Z(n21767) );
  AND U22125 ( .A(n21768), .B(n21769), .Z(n21662) );
  NANDN U22126 ( .A(n21770), .B(n21771), .Z(n21769) );
  OR U22127 ( .A(n21772), .B(n21773), .Z(n21771) );
  NAND U22128 ( .A(n21773), .B(n21772), .Z(n21768) );
  ANDN U22129 ( .B(B[120]), .A(n30), .Z(n21664) );
  XNOR U22130 ( .A(n21672), .B(n21774), .Z(n21665) );
  XNOR U22131 ( .A(n21671), .B(n21669), .Z(n21774) );
  AND U22132 ( .A(n21775), .B(n21776), .Z(n21669) );
  NANDN U22133 ( .A(n21777), .B(n21778), .Z(n21776) );
  NANDN U22134 ( .A(n21779), .B(n21780), .Z(n21778) );
  NANDN U22135 ( .A(n21780), .B(n21779), .Z(n21775) );
  ANDN U22136 ( .B(B[121]), .A(n31), .Z(n21671) );
  XNOR U22137 ( .A(n21679), .B(n21781), .Z(n21672) );
  XNOR U22138 ( .A(n21678), .B(n21676), .Z(n21781) );
  AND U22139 ( .A(n21782), .B(n21783), .Z(n21676) );
  NANDN U22140 ( .A(n21784), .B(n21785), .Z(n21783) );
  OR U22141 ( .A(n21786), .B(n21787), .Z(n21785) );
  NAND U22142 ( .A(n21787), .B(n21786), .Z(n21782) );
  ANDN U22143 ( .B(B[122]), .A(n32), .Z(n21678) );
  XNOR U22144 ( .A(n21686), .B(n21788), .Z(n21679) );
  XNOR U22145 ( .A(n21685), .B(n21683), .Z(n21788) );
  AND U22146 ( .A(n21789), .B(n21790), .Z(n21683) );
  NANDN U22147 ( .A(n21791), .B(n21792), .Z(n21790) );
  NANDN U22148 ( .A(n21793), .B(n21794), .Z(n21792) );
  NANDN U22149 ( .A(n21794), .B(n21793), .Z(n21789) );
  ANDN U22150 ( .B(B[123]), .A(n33), .Z(n21685) );
  XNOR U22151 ( .A(n21693), .B(n21795), .Z(n21686) );
  XNOR U22152 ( .A(n21692), .B(n21690), .Z(n21795) );
  AND U22153 ( .A(n21796), .B(n21797), .Z(n21690) );
  NANDN U22154 ( .A(n21798), .B(n21799), .Z(n21797) );
  OR U22155 ( .A(n21800), .B(n21801), .Z(n21799) );
  NAND U22156 ( .A(n21801), .B(n21800), .Z(n21796) );
  ANDN U22157 ( .B(B[124]), .A(n34), .Z(n21692) );
  XNOR U22158 ( .A(n21700), .B(n21802), .Z(n21693) );
  XNOR U22159 ( .A(n21699), .B(n21697), .Z(n21802) );
  AND U22160 ( .A(n21803), .B(n21804), .Z(n21697) );
  NANDN U22161 ( .A(n21805), .B(n21806), .Z(n21804) );
  NANDN U22162 ( .A(n21807), .B(n21808), .Z(n21806) );
  NANDN U22163 ( .A(n21808), .B(n21807), .Z(n21803) );
  ANDN U22164 ( .B(B[125]), .A(n35), .Z(n21699) );
  XNOR U22165 ( .A(n21707), .B(n21809), .Z(n21700) );
  XNOR U22166 ( .A(n21706), .B(n21704), .Z(n21809) );
  AND U22167 ( .A(n21810), .B(n21811), .Z(n21704) );
  NANDN U22168 ( .A(n21812), .B(n21813), .Z(n21811) );
  OR U22169 ( .A(n21814), .B(n21815), .Z(n21813) );
  NAND U22170 ( .A(n21815), .B(n21814), .Z(n21810) );
  ANDN U22171 ( .B(B[126]), .A(n36), .Z(n21706) );
  XNOR U22172 ( .A(n21714), .B(n21816), .Z(n21707) );
  XNOR U22173 ( .A(n21713), .B(n21711), .Z(n21816) );
  AND U22174 ( .A(n21817), .B(n21818), .Z(n21711) );
  NANDN U22175 ( .A(n21819), .B(n21820), .Z(n21818) );
  NANDN U22176 ( .A(n21821), .B(n21822), .Z(n21820) );
  NANDN U22177 ( .A(n21822), .B(n21821), .Z(n21817) );
  ANDN U22178 ( .B(B[127]), .A(n37), .Z(n21713) );
  XNOR U22179 ( .A(n21721), .B(n21823), .Z(n21714) );
  XNOR U22180 ( .A(n21720), .B(n21718), .Z(n21823) );
  AND U22181 ( .A(n21824), .B(n21825), .Z(n21718) );
  NANDN U22182 ( .A(n21826), .B(n21827), .Z(n21825) );
  OR U22183 ( .A(n21828), .B(n21829), .Z(n21827) );
  NAND U22184 ( .A(n21829), .B(n21828), .Z(n21824) );
  ANDN U22185 ( .B(B[128]), .A(n38), .Z(n21720) );
  XNOR U22186 ( .A(n21728), .B(n21830), .Z(n21721) );
  XNOR U22187 ( .A(n21727), .B(n21725), .Z(n21830) );
  AND U22188 ( .A(n21831), .B(n21832), .Z(n21725) );
  NANDN U22189 ( .A(n21833), .B(n21834), .Z(n21832) );
  NANDN U22190 ( .A(n21835), .B(n21836), .Z(n21834) );
  NANDN U22191 ( .A(n21836), .B(n21835), .Z(n21831) );
  ANDN U22192 ( .B(B[129]), .A(n39), .Z(n21727) );
  XNOR U22193 ( .A(n21735), .B(n21837), .Z(n21728) );
  XNOR U22194 ( .A(n21734), .B(n21732), .Z(n21837) );
  AND U22195 ( .A(n21838), .B(n21839), .Z(n21732) );
  NANDN U22196 ( .A(n21840), .B(n21841), .Z(n21839) );
  OR U22197 ( .A(n21842), .B(n21843), .Z(n21841) );
  NAND U22198 ( .A(n21843), .B(n21842), .Z(n21838) );
  ANDN U22199 ( .B(B[130]), .A(n40), .Z(n21734) );
  XNOR U22200 ( .A(n21742), .B(n21844), .Z(n21735) );
  XNOR U22201 ( .A(n21741), .B(n21739), .Z(n21844) );
  AND U22202 ( .A(n21845), .B(n21846), .Z(n21739) );
  NANDN U22203 ( .A(n21847), .B(n21848), .Z(n21846) );
  NAND U22204 ( .A(n21849), .B(n21850), .Z(n21848) );
  ANDN U22205 ( .B(B[131]), .A(n41), .Z(n21741) );
  XOR U22206 ( .A(n21748), .B(n21851), .Z(n21742) );
  XNOR U22207 ( .A(n21746), .B(n21749), .Z(n21851) );
  NAND U22208 ( .A(A[2]), .B(B[132]), .Z(n21749) );
  NANDN U22209 ( .A(n21852), .B(n21853), .Z(n21746) );
  AND U22210 ( .A(A[0]), .B(B[133]), .Z(n21853) );
  XNOR U22211 ( .A(n21751), .B(n21854), .Z(n21748) );
  NAND U22212 ( .A(A[0]), .B(B[134]), .Z(n21854) );
  NAND U22213 ( .A(B[133]), .B(A[1]), .Z(n21751) );
  NAND U22214 ( .A(n21855), .B(n21856), .Z(n487) );
  NANDN U22215 ( .A(n21857), .B(n21858), .Z(n21856) );
  OR U22216 ( .A(n21859), .B(n21860), .Z(n21858) );
  NAND U22217 ( .A(n21860), .B(n21859), .Z(n21855) );
  XOR U22218 ( .A(n489), .B(n488), .Z(\A1[131] ) );
  XOR U22219 ( .A(n21860), .B(n21861), .Z(n488) );
  XNOR U22220 ( .A(n21859), .B(n21857), .Z(n21861) );
  AND U22221 ( .A(n21862), .B(n21863), .Z(n21857) );
  NANDN U22222 ( .A(n21864), .B(n21865), .Z(n21863) );
  NANDN U22223 ( .A(n21866), .B(n21867), .Z(n21865) );
  NANDN U22224 ( .A(n21867), .B(n21866), .Z(n21862) );
  ANDN U22225 ( .B(B[118]), .A(n29), .Z(n21859) );
  XNOR U22226 ( .A(n21766), .B(n21868), .Z(n21860) );
  XNOR U22227 ( .A(n21765), .B(n21763), .Z(n21868) );
  AND U22228 ( .A(n21869), .B(n21870), .Z(n21763) );
  NANDN U22229 ( .A(n21871), .B(n21872), .Z(n21870) );
  OR U22230 ( .A(n21873), .B(n21874), .Z(n21872) );
  NAND U22231 ( .A(n21874), .B(n21873), .Z(n21869) );
  ANDN U22232 ( .B(B[119]), .A(n30), .Z(n21765) );
  XNOR U22233 ( .A(n21773), .B(n21875), .Z(n21766) );
  XNOR U22234 ( .A(n21772), .B(n21770), .Z(n21875) );
  AND U22235 ( .A(n21876), .B(n21877), .Z(n21770) );
  NANDN U22236 ( .A(n21878), .B(n21879), .Z(n21877) );
  NANDN U22237 ( .A(n21880), .B(n21881), .Z(n21879) );
  NANDN U22238 ( .A(n21881), .B(n21880), .Z(n21876) );
  ANDN U22239 ( .B(B[120]), .A(n31), .Z(n21772) );
  XNOR U22240 ( .A(n21780), .B(n21882), .Z(n21773) );
  XNOR U22241 ( .A(n21779), .B(n21777), .Z(n21882) );
  AND U22242 ( .A(n21883), .B(n21884), .Z(n21777) );
  NANDN U22243 ( .A(n21885), .B(n21886), .Z(n21884) );
  OR U22244 ( .A(n21887), .B(n21888), .Z(n21886) );
  NAND U22245 ( .A(n21888), .B(n21887), .Z(n21883) );
  ANDN U22246 ( .B(B[121]), .A(n32), .Z(n21779) );
  XNOR U22247 ( .A(n21787), .B(n21889), .Z(n21780) );
  XNOR U22248 ( .A(n21786), .B(n21784), .Z(n21889) );
  AND U22249 ( .A(n21890), .B(n21891), .Z(n21784) );
  NANDN U22250 ( .A(n21892), .B(n21893), .Z(n21891) );
  NANDN U22251 ( .A(n21894), .B(n21895), .Z(n21893) );
  NANDN U22252 ( .A(n21895), .B(n21894), .Z(n21890) );
  ANDN U22253 ( .B(B[122]), .A(n33), .Z(n21786) );
  XNOR U22254 ( .A(n21794), .B(n21896), .Z(n21787) );
  XNOR U22255 ( .A(n21793), .B(n21791), .Z(n21896) );
  AND U22256 ( .A(n21897), .B(n21898), .Z(n21791) );
  NANDN U22257 ( .A(n21899), .B(n21900), .Z(n21898) );
  OR U22258 ( .A(n21901), .B(n21902), .Z(n21900) );
  NAND U22259 ( .A(n21902), .B(n21901), .Z(n21897) );
  ANDN U22260 ( .B(B[123]), .A(n34), .Z(n21793) );
  XNOR U22261 ( .A(n21801), .B(n21903), .Z(n21794) );
  XNOR U22262 ( .A(n21800), .B(n21798), .Z(n21903) );
  AND U22263 ( .A(n21904), .B(n21905), .Z(n21798) );
  NANDN U22264 ( .A(n21906), .B(n21907), .Z(n21905) );
  NANDN U22265 ( .A(n21908), .B(n21909), .Z(n21907) );
  NANDN U22266 ( .A(n21909), .B(n21908), .Z(n21904) );
  ANDN U22267 ( .B(B[124]), .A(n35), .Z(n21800) );
  XNOR U22268 ( .A(n21808), .B(n21910), .Z(n21801) );
  XNOR U22269 ( .A(n21807), .B(n21805), .Z(n21910) );
  AND U22270 ( .A(n21911), .B(n21912), .Z(n21805) );
  NANDN U22271 ( .A(n21913), .B(n21914), .Z(n21912) );
  OR U22272 ( .A(n21915), .B(n21916), .Z(n21914) );
  NAND U22273 ( .A(n21916), .B(n21915), .Z(n21911) );
  ANDN U22274 ( .B(B[125]), .A(n36), .Z(n21807) );
  XNOR U22275 ( .A(n21815), .B(n21917), .Z(n21808) );
  XNOR U22276 ( .A(n21814), .B(n21812), .Z(n21917) );
  AND U22277 ( .A(n21918), .B(n21919), .Z(n21812) );
  NANDN U22278 ( .A(n21920), .B(n21921), .Z(n21919) );
  NANDN U22279 ( .A(n21922), .B(n21923), .Z(n21921) );
  NANDN U22280 ( .A(n21923), .B(n21922), .Z(n21918) );
  ANDN U22281 ( .B(B[126]), .A(n37), .Z(n21814) );
  XNOR U22282 ( .A(n21822), .B(n21924), .Z(n21815) );
  XNOR U22283 ( .A(n21821), .B(n21819), .Z(n21924) );
  AND U22284 ( .A(n21925), .B(n21926), .Z(n21819) );
  NANDN U22285 ( .A(n21927), .B(n21928), .Z(n21926) );
  OR U22286 ( .A(n21929), .B(n21930), .Z(n21928) );
  NAND U22287 ( .A(n21930), .B(n21929), .Z(n21925) );
  ANDN U22288 ( .B(B[127]), .A(n38), .Z(n21821) );
  XNOR U22289 ( .A(n21829), .B(n21931), .Z(n21822) );
  XNOR U22290 ( .A(n21828), .B(n21826), .Z(n21931) );
  AND U22291 ( .A(n21932), .B(n21933), .Z(n21826) );
  NANDN U22292 ( .A(n21934), .B(n21935), .Z(n21933) );
  NANDN U22293 ( .A(n21936), .B(n21937), .Z(n21935) );
  NANDN U22294 ( .A(n21937), .B(n21936), .Z(n21932) );
  ANDN U22295 ( .B(B[128]), .A(n39), .Z(n21828) );
  XNOR U22296 ( .A(n21836), .B(n21938), .Z(n21829) );
  XNOR U22297 ( .A(n21835), .B(n21833), .Z(n21938) );
  AND U22298 ( .A(n21939), .B(n21940), .Z(n21833) );
  NANDN U22299 ( .A(n21941), .B(n21942), .Z(n21940) );
  OR U22300 ( .A(n21943), .B(n21944), .Z(n21942) );
  NAND U22301 ( .A(n21944), .B(n21943), .Z(n21939) );
  ANDN U22302 ( .B(B[129]), .A(n40), .Z(n21835) );
  XNOR U22303 ( .A(n21843), .B(n21945), .Z(n21836) );
  XNOR U22304 ( .A(n21842), .B(n21840), .Z(n21945) );
  AND U22305 ( .A(n21946), .B(n21947), .Z(n21840) );
  NANDN U22306 ( .A(n21948), .B(n21949), .Z(n21947) );
  NAND U22307 ( .A(n21950), .B(n21951), .Z(n21949) );
  ANDN U22308 ( .B(B[130]), .A(n41), .Z(n21842) );
  XOR U22309 ( .A(n21849), .B(n21952), .Z(n21843) );
  XNOR U22310 ( .A(n21847), .B(n21850), .Z(n21952) );
  NAND U22311 ( .A(A[2]), .B(B[131]), .Z(n21850) );
  NANDN U22312 ( .A(n21953), .B(n21954), .Z(n21847) );
  AND U22313 ( .A(A[0]), .B(B[132]), .Z(n21954) );
  XNOR U22314 ( .A(n21852), .B(n21955), .Z(n21849) );
  NAND U22315 ( .A(A[0]), .B(B[133]), .Z(n21955) );
  NAND U22316 ( .A(B[132]), .B(A[1]), .Z(n21852) );
  NAND U22317 ( .A(n21956), .B(n21957), .Z(n489) );
  NANDN U22318 ( .A(n21958), .B(n21959), .Z(n21957) );
  OR U22319 ( .A(n21960), .B(n21961), .Z(n21959) );
  NAND U22320 ( .A(n21961), .B(n21960), .Z(n21956) );
  XOR U22321 ( .A(n491), .B(n490), .Z(\A1[130] ) );
  XOR U22322 ( .A(n21961), .B(n21962), .Z(n490) );
  XNOR U22323 ( .A(n21960), .B(n21958), .Z(n21962) );
  AND U22324 ( .A(n21963), .B(n21964), .Z(n21958) );
  NANDN U22325 ( .A(n21965), .B(n21966), .Z(n21964) );
  NANDN U22326 ( .A(n21967), .B(n21968), .Z(n21966) );
  NANDN U22327 ( .A(n21968), .B(n21967), .Z(n21963) );
  ANDN U22328 ( .B(B[117]), .A(n29), .Z(n21960) );
  XNOR U22329 ( .A(n21867), .B(n21969), .Z(n21961) );
  XNOR U22330 ( .A(n21866), .B(n21864), .Z(n21969) );
  AND U22331 ( .A(n21970), .B(n21971), .Z(n21864) );
  NANDN U22332 ( .A(n21972), .B(n21973), .Z(n21971) );
  OR U22333 ( .A(n21974), .B(n21975), .Z(n21973) );
  NAND U22334 ( .A(n21975), .B(n21974), .Z(n21970) );
  ANDN U22335 ( .B(B[118]), .A(n30), .Z(n21866) );
  XNOR U22336 ( .A(n21874), .B(n21976), .Z(n21867) );
  XNOR U22337 ( .A(n21873), .B(n21871), .Z(n21976) );
  AND U22338 ( .A(n21977), .B(n21978), .Z(n21871) );
  NANDN U22339 ( .A(n21979), .B(n21980), .Z(n21978) );
  NANDN U22340 ( .A(n21981), .B(n21982), .Z(n21980) );
  NANDN U22341 ( .A(n21982), .B(n21981), .Z(n21977) );
  ANDN U22342 ( .B(B[119]), .A(n31), .Z(n21873) );
  XNOR U22343 ( .A(n21881), .B(n21983), .Z(n21874) );
  XNOR U22344 ( .A(n21880), .B(n21878), .Z(n21983) );
  AND U22345 ( .A(n21984), .B(n21985), .Z(n21878) );
  NANDN U22346 ( .A(n21986), .B(n21987), .Z(n21985) );
  OR U22347 ( .A(n21988), .B(n21989), .Z(n21987) );
  NAND U22348 ( .A(n21989), .B(n21988), .Z(n21984) );
  ANDN U22349 ( .B(B[120]), .A(n32), .Z(n21880) );
  XNOR U22350 ( .A(n21888), .B(n21990), .Z(n21881) );
  XNOR U22351 ( .A(n21887), .B(n21885), .Z(n21990) );
  AND U22352 ( .A(n21991), .B(n21992), .Z(n21885) );
  NANDN U22353 ( .A(n21993), .B(n21994), .Z(n21992) );
  NANDN U22354 ( .A(n21995), .B(n21996), .Z(n21994) );
  NANDN U22355 ( .A(n21996), .B(n21995), .Z(n21991) );
  ANDN U22356 ( .B(B[121]), .A(n33), .Z(n21887) );
  XNOR U22357 ( .A(n21895), .B(n21997), .Z(n21888) );
  XNOR U22358 ( .A(n21894), .B(n21892), .Z(n21997) );
  AND U22359 ( .A(n21998), .B(n21999), .Z(n21892) );
  NANDN U22360 ( .A(n22000), .B(n22001), .Z(n21999) );
  OR U22361 ( .A(n22002), .B(n22003), .Z(n22001) );
  NAND U22362 ( .A(n22003), .B(n22002), .Z(n21998) );
  ANDN U22363 ( .B(B[122]), .A(n34), .Z(n21894) );
  XNOR U22364 ( .A(n21902), .B(n22004), .Z(n21895) );
  XNOR U22365 ( .A(n21901), .B(n21899), .Z(n22004) );
  AND U22366 ( .A(n22005), .B(n22006), .Z(n21899) );
  NANDN U22367 ( .A(n22007), .B(n22008), .Z(n22006) );
  NANDN U22368 ( .A(n22009), .B(n22010), .Z(n22008) );
  NANDN U22369 ( .A(n22010), .B(n22009), .Z(n22005) );
  ANDN U22370 ( .B(B[123]), .A(n35), .Z(n21901) );
  XNOR U22371 ( .A(n21909), .B(n22011), .Z(n21902) );
  XNOR U22372 ( .A(n21908), .B(n21906), .Z(n22011) );
  AND U22373 ( .A(n22012), .B(n22013), .Z(n21906) );
  NANDN U22374 ( .A(n22014), .B(n22015), .Z(n22013) );
  OR U22375 ( .A(n22016), .B(n22017), .Z(n22015) );
  NAND U22376 ( .A(n22017), .B(n22016), .Z(n22012) );
  ANDN U22377 ( .B(B[124]), .A(n36), .Z(n21908) );
  XNOR U22378 ( .A(n21916), .B(n22018), .Z(n21909) );
  XNOR U22379 ( .A(n21915), .B(n21913), .Z(n22018) );
  AND U22380 ( .A(n22019), .B(n22020), .Z(n21913) );
  NANDN U22381 ( .A(n22021), .B(n22022), .Z(n22020) );
  NANDN U22382 ( .A(n22023), .B(n22024), .Z(n22022) );
  NANDN U22383 ( .A(n22024), .B(n22023), .Z(n22019) );
  ANDN U22384 ( .B(B[125]), .A(n37), .Z(n21915) );
  XNOR U22385 ( .A(n21923), .B(n22025), .Z(n21916) );
  XNOR U22386 ( .A(n21922), .B(n21920), .Z(n22025) );
  AND U22387 ( .A(n22026), .B(n22027), .Z(n21920) );
  NANDN U22388 ( .A(n22028), .B(n22029), .Z(n22027) );
  OR U22389 ( .A(n22030), .B(n22031), .Z(n22029) );
  NAND U22390 ( .A(n22031), .B(n22030), .Z(n22026) );
  ANDN U22391 ( .B(B[126]), .A(n38), .Z(n21922) );
  XNOR U22392 ( .A(n21930), .B(n22032), .Z(n21923) );
  XNOR U22393 ( .A(n21929), .B(n21927), .Z(n22032) );
  AND U22394 ( .A(n22033), .B(n22034), .Z(n21927) );
  NANDN U22395 ( .A(n22035), .B(n22036), .Z(n22034) );
  NANDN U22396 ( .A(n22037), .B(n22038), .Z(n22036) );
  NANDN U22397 ( .A(n22038), .B(n22037), .Z(n22033) );
  ANDN U22398 ( .B(B[127]), .A(n39), .Z(n21929) );
  XNOR U22399 ( .A(n21937), .B(n22039), .Z(n21930) );
  XNOR U22400 ( .A(n21936), .B(n21934), .Z(n22039) );
  AND U22401 ( .A(n22040), .B(n22041), .Z(n21934) );
  NANDN U22402 ( .A(n22042), .B(n22043), .Z(n22041) );
  OR U22403 ( .A(n22044), .B(n22045), .Z(n22043) );
  NAND U22404 ( .A(n22045), .B(n22044), .Z(n22040) );
  ANDN U22405 ( .B(B[128]), .A(n40), .Z(n21936) );
  XNOR U22406 ( .A(n21944), .B(n22046), .Z(n21937) );
  XNOR U22407 ( .A(n21943), .B(n21941), .Z(n22046) );
  AND U22408 ( .A(n22047), .B(n22048), .Z(n21941) );
  NANDN U22409 ( .A(n22049), .B(n22050), .Z(n22048) );
  NAND U22410 ( .A(n22051), .B(n22052), .Z(n22050) );
  ANDN U22411 ( .B(B[129]), .A(n41), .Z(n21943) );
  XOR U22412 ( .A(n21950), .B(n22053), .Z(n21944) );
  XNOR U22413 ( .A(n21948), .B(n21951), .Z(n22053) );
  NAND U22414 ( .A(A[2]), .B(B[130]), .Z(n21951) );
  NANDN U22415 ( .A(n22054), .B(n22055), .Z(n21948) );
  AND U22416 ( .A(A[0]), .B(B[131]), .Z(n22055) );
  XNOR U22417 ( .A(n21953), .B(n22056), .Z(n21950) );
  NAND U22418 ( .A(A[0]), .B(B[132]), .Z(n22056) );
  NAND U22419 ( .A(B[131]), .B(A[1]), .Z(n21953) );
  NAND U22420 ( .A(n22057), .B(n22058), .Z(n491) );
  NANDN U22421 ( .A(n22059), .B(n22060), .Z(n22058) );
  OR U22422 ( .A(n22061), .B(n22062), .Z(n22060) );
  NAND U22423 ( .A(n22062), .B(n22061), .Z(n22057) );
  XOR U22424 ( .A(n20964), .B(n22063), .Z(\A1[12] ) );
  XNOR U22425 ( .A(n20963), .B(n20962), .Z(n22063) );
  NAND U22426 ( .A(n22064), .B(n22065), .Z(n20962) );
  NANDN U22427 ( .A(n22066), .B(n22067), .Z(n22065) );
  OR U22428 ( .A(n22068), .B(n22069), .Z(n22067) );
  NAND U22429 ( .A(n22069), .B(n22068), .Z(n22064) );
  ANDN U22430 ( .B(B[0]), .A(n30), .Z(n20963) );
  XNOR U22431 ( .A(n20971), .B(n22070), .Z(n20964) );
  XNOR U22432 ( .A(n20970), .B(n20968), .Z(n22070) );
  AND U22433 ( .A(n22071), .B(n22072), .Z(n20968) );
  NANDN U22434 ( .A(n22073), .B(n22074), .Z(n22072) );
  NANDN U22435 ( .A(n22075), .B(n22076), .Z(n22074) );
  NANDN U22436 ( .A(n22076), .B(n22075), .Z(n22071) );
  ANDN U22437 ( .B(B[1]), .A(n31), .Z(n20970) );
  XNOR U22438 ( .A(n20978), .B(n22077), .Z(n20971) );
  XNOR U22439 ( .A(n20977), .B(n20975), .Z(n22077) );
  AND U22440 ( .A(n22078), .B(n22079), .Z(n20975) );
  NANDN U22441 ( .A(n22080), .B(n22081), .Z(n22079) );
  OR U22442 ( .A(n22082), .B(n22083), .Z(n22081) );
  NAND U22443 ( .A(n22083), .B(n22082), .Z(n22078) );
  ANDN U22444 ( .B(B[2]), .A(n32), .Z(n20977) );
  XNOR U22445 ( .A(n20985), .B(n22084), .Z(n20978) );
  XNOR U22446 ( .A(n20984), .B(n20982), .Z(n22084) );
  AND U22447 ( .A(n22085), .B(n22086), .Z(n20982) );
  NANDN U22448 ( .A(n22087), .B(n22088), .Z(n22086) );
  NANDN U22449 ( .A(n22089), .B(n22090), .Z(n22088) );
  NANDN U22450 ( .A(n22090), .B(n22089), .Z(n22085) );
  ANDN U22451 ( .B(B[3]), .A(n33), .Z(n20984) );
  XNOR U22452 ( .A(n20992), .B(n22091), .Z(n20985) );
  XNOR U22453 ( .A(n20991), .B(n20989), .Z(n22091) );
  AND U22454 ( .A(n22092), .B(n22093), .Z(n20989) );
  NANDN U22455 ( .A(n22094), .B(n22095), .Z(n22093) );
  OR U22456 ( .A(n22096), .B(n22097), .Z(n22095) );
  NAND U22457 ( .A(n22097), .B(n22096), .Z(n22092) );
  ANDN U22458 ( .B(B[4]), .A(n34), .Z(n20991) );
  XNOR U22459 ( .A(n20999), .B(n22098), .Z(n20992) );
  XNOR U22460 ( .A(n20998), .B(n20996), .Z(n22098) );
  AND U22461 ( .A(n22099), .B(n22100), .Z(n20996) );
  NANDN U22462 ( .A(n22101), .B(n22102), .Z(n22100) );
  NANDN U22463 ( .A(n22103), .B(n22104), .Z(n22102) );
  NANDN U22464 ( .A(n22104), .B(n22103), .Z(n22099) );
  ANDN U22465 ( .B(B[5]), .A(n35), .Z(n20998) );
  XNOR U22466 ( .A(n21006), .B(n22105), .Z(n20999) );
  XNOR U22467 ( .A(n21005), .B(n21003), .Z(n22105) );
  AND U22468 ( .A(n22106), .B(n22107), .Z(n21003) );
  NANDN U22469 ( .A(n22108), .B(n22109), .Z(n22107) );
  OR U22470 ( .A(n22110), .B(n22111), .Z(n22109) );
  NAND U22471 ( .A(n22111), .B(n22110), .Z(n22106) );
  ANDN U22472 ( .B(B[6]), .A(n36), .Z(n21005) );
  XNOR U22473 ( .A(n21013), .B(n22112), .Z(n21006) );
  XNOR U22474 ( .A(n21012), .B(n21010), .Z(n22112) );
  AND U22475 ( .A(n22113), .B(n22114), .Z(n21010) );
  NANDN U22476 ( .A(n22115), .B(n22116), .Z(n22114) );
  NANDN U22477 ( .A(n22117), .B(n22118), .Z(n22116) );
  NANDN U22478 ( .A(n22118), .B(n22117), .Z(n22113) );
  ANDN U22479 ( .B(B[7]), .A(n37), .Z(n21012) );
  XNOR U22480 ( .A(n21020), .B(n22119), .Z(n21013) );
  XNOR U22481 ( .A(n21019), .B(n21017), .Z(n22119) );
  AND U22482 ( .A(n22120), .B(n22121), .Z(n21017) );
  NANDN U22483 ( .A(n22122), .B(n22123), .Z(n22121) );
  OR U22484 ( .A(n22124), .B(n22125), .Z(n22123) );
  NAND U22485 ( .A(n22125), .B(n22124), .Z(n22120) );
  ANDN U22486 ( .B(B[8]), .A(n38), .Z(n21019) );
  XNOR U22487 ( .A(n21027), .B(n22126), .Z(n21020) );
  XNOR U22488 ( .A(n21026), .B(n21024), .Z(n22126) );
  AND U22489 ( .A(n22127), .B(n22128), .Z(n21024) );
  NANDN U22490 ( .A(n22129), .B(n22130), .Z(n22128) );
  NANDN U22491 ( .A(n22131), .B(n22132), .Z(n22130) );
  NANDN U22492 ( .A(n22132), .B(n22131), .Z(n22127) );
  ANDN U22493 ( .B(B[9]), .A(n39), .Z(n21026) );
  XNOR U22494 ( .A(n21034), .B(n22133), .Z(n21027) );
  XNOR U22495 ( .A(n21033), .B(n21031), .Z(n22133) );
  AND U22496 ( .A(n22134), .B(n22135), .Z(n21031) );
  NANDN U22497 ( .A(n22136), .B(n22137), .Z(n22135) );
  OR U22498 ( .A(n22138), .B(n22139), .Z(n22137) );
  NAND U22499 ( .A(n22139), .B(n22138), .Z(n22134) );
  ANDN U22500 ( .B(B[10]), .A(n40), .Z(n21033) );
  XNOR U22501 ( .A(n21041), .B(n22140), .Z(n21034) );
  XNOR U22502 ( .A(n21040), .B(n21038), .Z(n22140) );
  AND U22503 ( .A(n22141), .B(n22142), .Z(n21038) );
  NANDN U22504 ( .A(n22143), .B(n22144), .Z(n22142) );
  NAND U22505 ( .A(n22145), .B(n22146), .Z(n22144) );
  ANDN U22506 ( .B(B[11]), .A(n41), .Z(n21040) );
  XOR U22507 ( .A(n21047), .B(n22147), .Z(n21041) );
  XNOR U22508 ( .A(n21045), .B(n21048), .Z(n22147) );
  NAND U22509 ( .A(A[2]), .B(B[12]), .Z(n21048) );
  NANDN U22510 ( .A(n22148), .B(n22149), .Z(n21045) );
  AND U22511 ( .A(A[0]), .B(B[13]), .Z(n22149) );
  XNOR U22512 ( .A(n21050), .B(n22150), .Z(n21047) );
  NAND U22513 ( .A(A[0]), .B(B[14]), .Z(n22150) );
  NAND U22514 ( .A(B[13]), .B(A[1]), .Z(n21050) );
  XOR U22515 ( .A(n493), .B(n492), .Z(\A1[129] ) );
  XOR U22516 ( .A(n22062), .B(n22151), .Z(n492) );
  XNOR U22517 ( .A(n22061), .B(n22059), .Z(n22151) );
  AND U22518 ( .A(n22152), .B(n22153), .Z(n22059) );
  NANDN U22519 ( .A(n22154), .B(n22155), .Z(n22153) );
  NANDN U22520 ( .A(n22156), .B(n22157), .Z(n22155) );
  NANDN U22521 ( .A(n22157), .B(n22156), .Z(n22152) );
  ANDN U22522 ( .B(B[116]), .A(n29), .Z(n22061) );
  XNOR U22523 ( .A(n21968), .B(n22158), .Z(n22062) );
  XNOR U22524 ( .A(n21967), .B(n21965), .Z(n22158) );
  AND U22525 ( .A(n22159), .B(n22160), .Z(n21965) );
  NANDN U22526 ( .A(n22161), .B(n22162), .Z(n22160) );
  OR U22527 ( .A(n22163), .B(n22164), .Z(n22162) );
  NAND U22528 ( .A(n22164), .B(n22163), .Z(n22159) );
  ANDN U22529 ( .B(B[117]), .A(n30), .Z(n21967) );
  XNOR U22530 ( .A(n21975), .B(n22165), .Z(n21968) );
  XNOR U22531 ( .A(n21974), .B(n21972), .Z(n22165) );
  AND U22532 ( .A(n22166), .B(n22167), .Z(n21972) );
  NANDN U22533 ( .A(n22168), .B(n22169), .Z(n22167) );
  NANDN U22534 ( .A(n22170), .B(n22171), .Z(n22169) );
  NANDN U22535 ( .A(n22171), .B(n22170), .Z(n22166) );
  ANDN U22536 ( .B(B[118]), .A(n31), .Z(n21974) );
  XNOR U22537 ( .A(n21982), .B(n22172), .Z(n21975) );
  XNOR U22538 ( .A(n21981), .B(n21979), .Z(n22172) );
  AND U22539 ( .A(n22173), .B(n22174), .Z(n21979) );
  NANDN U22540 ( .A(n22175), .B(n22176), .Z(n22174) );
  OR U22541 ( .A(n22177), .B(n22178), .Z(n22176) );
  NAND U22542 ( .A(n22178), .B(n22177), .Z(n22173) );
  ANDN U22543 ( .B(B[119]), .A(n32), .Z(n21981) );
  XNOR U22544 ( .A(n21989), .B(n22179), .Z(n21982) );
  XNOR U22545 ( .A(n21988), .B(n21986), .Z(n22179) );
  AND U22546 ( .A(n22180), .B(n22181), .Z(n21986) );
  NANDN U22547 ( .A(n22182), .B(n22183), .Z(n22181) );
  NANDN U22548 ( .A(n22184), .B(n22185), .Z(n22183) );
  NANDN U22549 ( .A(n22185), .B(n22184), .Z(n22180) );
  ANDN U22550 ( .B(B[120]), .A(n33), .Z(n21988) );
  XNOR U22551 ( .A(n21996), .B(n22186), .Z(n21989) );
  XNOR U22552 ( .A(n21995), .B(n21993), .Z(n22186) );
  AND U22553 ( .A(n22187), .B(n22188), .Z(n21993) );
  NANDN U22554 ( .A(n22189), .B(n22190), .Z(n22188) );
  OR U22555 ( .A(n22191), .B(n22192), .Z(n22190) );
  NAND U22556 ( .A(n22192), .B(n22191), .Z(n22187) );
  ANDN U22557 ( .B(B[121]), .A(n34), .Z(n21995) );
  XNOR U22558 ( .A(n22003), .B(n22193), .Z(n21996) );
  XNOR U22559 ( .A(n22002), .B(n22000), .Z(n22193) );
  AND U22560 ( .A(n22194), .B(n22195), .Z(n22000) );
  NANDN U22561 ( .A(n22196), .B(n22197), .Z(n22195) );
  NANDN U22562 ( .A(n22198), .B(n22199), .Z(n22197) );
  NANDN U22563 ( .A(n22199), .B(n22198), .Z(n22194) );
  ANDN U22564 ( .B(B[122]), .A(n35), .Z(n22002) );
  XNOR U22565 ( .A(n22010), .B(n22200), .Z(n22003) );
  XNOR U22566 ( .A(n22009), .B(n22007), .Z(n22200) );
  AND U22567 ( .A(n22201), .B(n22202), .Z(n22007) );
  NANDN U22568 ( .A(n22203), .B(n22204), .Z(n22202) );
  OR U22569 ( .A(n22205), .B(n22206), .Z(n22204) );
  NAND U22570 ( .A(n22206), .B(n22205), .Z(n22201) );
  ANDN U22571 ( .B(B[123]), .A(n36), .Z(n22009) );
  XNOR U22572 ( .A(n22017), .B(n22207), .Z(n22010) );
  XNOR U22573 ( .A(n22016), .B(n22014), .Z(n22207) );
  AND U22574 ( .A(n22208), .B(n22209), .Z(n22014) );
  NANDN U22575 ( .A(n22210), .B(n22211), .Z(n22209) );
  NANDN U22576 ( .A(n22212), .B(n22213), .Z(n22211) );
  NANDN U22577 ( .A(n22213), .B(n22212), .Z(n22208) );
  ANDN U22578 ( .B(B[124]), .A(n37), .Z(n22016) );
  XNOR U22579 ( .A(n22024), .B(n22214), .Z(n22017) );
  XNOR U22580 ( .A(n22023), .B(n22021), .Z(n22214) );
  AND U22581 ( .A(n22215), .B(n22216), .Z(n22021) );
  NANDN U22582 ( .A(n22217), .B(n22218), .Z(n22216) );
  OR U22583 ( .A(n22219), .B(n22220), .Z(n22218) );
  NAND U22584 ( .A(n22220), .B(n22219), .Z(n22215) );
  ANDN U22585 ( .B(B[125]), .A(n38), .Z(n22023) );
  XNOR U22586 ( .A(n22031), .B(n22221), .Z(n22024) );
  XNOR U22587 ( .A(n22030), .B(n22028), .Z(n22221) );
  AND U22588 ( .A(n22222), .B(n22223), .Z(n22028) );
  NANDN U22589 ( .A(n22224), .B(n22225), .Z(n22223) );
  NANDN U22590 ( .A(n22226), .B(n22227), .Z(n22225) );
  NANDN U22591 ( .A(n22227), .B(n22226), .Z(n22222) );
  ANDN U22592 ( .B(B[126]), .A(n39), .Z(n22030) );
  XNOR U22593 ( .A(n22038), .B(n22228), .Z(n22031) );
  XNOR U22594 ( .A(n22037), .B(n22035), .Z(n22228) );
  AND U22595 ( .A(n22229), .B(n22230), .Z(n22035) );
  NANDN U22596 ( .A(n22231), .B(n22232), .Z(n22230) );
  OR U22597 ( .A(n22233), .B(n22234), .Z(n22232) );
  NAND U22598 ( .A(n22234), .B(n22233), .Z(n22229) );
  ANDN U22599 ( .B(B[127]), .A(n40), .Z(n22037) );
  XNOR U22600 ( .A(n22045), .B(n22235), .Z(n22038) );
  XNOR U22601 ( .A(n22044), .B(n22042), .Z(n22235) );
  AND U22602 ( .A(n22236), .B(n22237), .Z(n22042) );
  NANDN U22603 ( .A(n22238), .B(n22239), .Z(n22237) );
  NAND U22604 ( .A(n22240), .B(n22241), .Z(n22239) );
  ANDN U22605 ( .B(B[128]), .A(n41), .Z(n22044) );
  XOR U22606 ( .A(n22051), .B(n22242), .Z(n22045) );
  XNOR U22607 ( .A(n22049), .B(n22052), .Z(n22242) );
  NAND U22608 ( .A(A[2]), .B(B[129]), .Z(n22052) );
  NANDN U22609 ( .A(n22243), .B(n22244), .Z(n22049) );
  AND U22610 ( .A(A[0]), .B(B[130]), .Z(n22244) );
  XNOR U22611 ( .A(n22054), .B(n22245), .Z(n22051) );
  NAND U22612 ( .A(A[0]), .B(B[131]), .Z(n22245) );
  NAND U22613 ( .A(B[130]), .B(A[1]), .Z(n22054) );
  NAND U22614 ( .A(n22246), .B(n22247), .Z(n493) );
  NANDN U22615 ( .A(n22248), .B(n22249), .Z(n22247) );
  OR U22616 ( .A(n22250), .B(n22251), .Z(n22249) );
  NAND U22617 ( .A(n22251), .B(n22250), .Z(n22246) );
  XOR U22618 ( .A(n495), .B(n494), .Z(\A1[128] ) );
  XOR U22619 ( .A(n22251), .B(n22252), .Z(n494) );
  XNOR U22620 ( .A(n22250), .B(n22248), .Z(n22252) );
  AND U22621 ( .A(n22253), .B(n22254), .Z(n22248) );
  NANDN U22622 ( .A(n22255), .B(n22256), .Z(n22254) );
  NANDN U22623 ( .A(n22257), .B(n22258), .Z(n22256) );
  NANDN U22624 ( .A(n22258), .B(n22257), .Z(n22253) );
  ANDN U22625 ( .B(B[115]), .A(n29), .Z(n22250) );
  XNOR U22626 ( .A(n22157), .B(n22259), .Z(n22251) );
  XNOR U22627 ( .A(n22156), .B(n22154), .Z(n22259) );
  AND U22628 ( .A(n22260), .B(n22261), .Z(n22154) );
  NANDN U22629 ( .A(n22262), .B(n22263), .Z(n22261) );
  OR U22630 ( .A(n22264), .B(n22265), .Z(n22263) );
  NAND U22631 ( .A(n22265), .B(n22264), .Z(n22260) );
  ANDN U22632 ( .B(B[116]), .A(n30), .Z(n22156) );
  XNOR U22633 ( .A(n22164), .B(n22266), .Z(n22157) );
  XNOR U22634 ( .A(n22163), .B(n22161), .Z(n22266) );
  AND U22635 ( .A(n22267), .B(n22268), .Z(n22161) );
  NANDN U22636 ( .A(n22269), .B(n22270), .Z(n22268) );
  NANDN U22637 ( .A(n22271), .B(n22272), .Z(n22270) );
  NANDN U22638 ( .A(n22272), .B(n22271), .Z(n22267) );
  ANDN U22639 ( .B(B[117]), .A(n31), .Z(n22163) );
  XNOR U22640 ( .A(n22171), .B(n22273), .Z(n22164) );
  XNOR U22641 ( .A(n22170), .B(n22168), .Z(n22273) );
  AND U22642 ( .A(n22274), .B(n22275), .Z(n22168) );
  NANDN U22643 ( .A(n22276), .B(n22277), .Z(n22275) );
  OR U22644 ( .A(n22278), .B(n22279), .Z(n22277) );
  NAND U22645 ( .A(n22279), .B(n22278), .Z(n22274) );
  ANDN U22646 ( .B(B[118]), .A(n32), .Z(n22170) );
  XNOR U22647 ( .A(n22178), .B(n22280), .Z(n22171) );
  XNOR U22648 ( .A(n22177), .B(n22175), .Z(n22280) );
  AND U22649 ( .A(n22281), .B(n22282), .Z(n22175) );
  NANDN U22650 ( .A(n22283), .B(n22284), .Z(n22282) );
  NANDN U22651 ( .A(n22285), .B(n22286), .Z(n22284) );
  NANDN U22652 ( .A(n22286), .B(n22285), .Z(n22281) );
  ANDN U22653 ( .B(B[119]), .A(n33), .Z(n22177) );
  XNOR U22654 ( .A(n22185), .B(n22287), .Z(n22178) );
  XNOR U22655 ( .A(n22184), .B(n22182), .Z(n22287) );
  AND U22656 ( .A(n22288), .B(n22289), .Z(n22182) );
  NANDN U22657 ( .A(n22290), .B(n22291), .Z(n22289) );
  OR U22658 ( .A(n22292), .B(n22293), .Z(n22291) );
  NAND U22659 ( .A(n22293), .B(n22292), .Z(n22288) );
  ANDN U22660 ( .B(B[120]), .A(n34), .Z(n22184) );
  XNOR U22661 ( .A(n22192), .B(n22294), .Z(n22185) );
  XNOR U22662 ( .A(n22191), .B(n22189), .Z(n22294) );
  AND U22663 ( .A(n22295), .B(n22296), .Z(n22189) );
  NANDN U22664 ( .A(n22297), .B(n22298), .Z(n22296) );
  NANDN U22665 ( .A(n22299), .B(n22300), .Z(n22298) );
  NANDN U22666 ( .A(n22300), .B(n22299), .Z(n22295) );
  ANDN U22667 ( .B(B[121]), .A(n35), .Z(n22191) );
  XNOR U22668 ( .A(n22199), .B(n22301), .Z(n22192) );
  XNOR U22669 ( .A(n22198), .B(n22196), .Z(n22301) );
  AND U22670 ( .A(n22302), .B(n22303), .Z(n22196) );
  NANDN U22671 ( .A(n22304), .B(n22305), .Z(n22303) );
  OR U22672 ( .A(n22306), .B(n22307), .Z(n22305) );
  NAND U22673 ( .A(n22307), .B(n22306), .Z(n22302) );
  ANDN U22674 ( .B(B[122]), .A(n36), .Z(n22198) );
  XNOR U22675 ( .A(n22206), .B(n22308), .Z(n22199) );
  XNOR U22676 ( .A(n22205), .B(n22203), .Z(n22308) );
  AND U22677 ( .A(n22309), .B(n22310), .Z(n22203) );
  NANDN U22678 ( .A(n22311), .B(n22312), .Z(n22310) );
  NANDN U22679 ( .A(n22313), .B(n22314), .Z(n22312) );
  NANDN U22680 ( .A(n22314), .B(n22313), .Z(n22309) );
  ANDN U22681 ( .B(B[123]), .A(n37), .Z(n22205) );
  XNOR U22682 ( .A(n22213), .B(n22315), .Z(n22206) );
  XNOR U22683 ( .A(n22212), .B(n22210), .Z(n22315) );
  AND U22684 ( .A(n22316), .B(n22317), .Z(n22210) );
  NANDN U22685 ( .A(n22318), .B(n22319), .Z(n22317) );
  OR U22686 ( .A(n22320), .B(n22321), .Z(n22319) );
  NAND U22687 ( .A(n22321), .B(n22320), .Z(n22316) );
  ANDN U22688 ( .B(B[124]), .A(n38), .Z(n22212) );
  XNOR U22689 ( .A(n22220), .B(n22322), .Z(n22213) );
  XNOR U22690 ( .A(n22219), .B(n22217), .Z(n22322) );
  AND U22691 ( .A(n22323), .B(n22324), .Z(n22217) );
  NANDN U22692 ( .A(n22325), .B(n22326), .Z(n22324) );
  NANDN U22693 ( .A(n22327), .B(n22328), .Z(n22326) );
  NANDN U22694 ( .A(n22328), .B(n22327), .Z(n22323) );
  ANDN U22695 ( .B(B[125]), .A(n39), .Z(n22219) );
  XNOR U22696 ( .A(n22227), .B(n22329), .Z(n22220) );
  XNOR U22697 ( .A(n22226), .B(n22224), .Z(n22329) );
  AND U22698 ( .A(n22330), .B(n22331), .Z(n22224) );
  NANDN U22699 ( .A(n22332), .B(n22333), .Z(n22331) );
  OR U22700 ( .A(n22334), .B(n22335), .Z(n22333) );
  NAND U22701 ( .A(n22335), .B(n22334), .Z(n22330) );
  ANDN U22702 ( .B(B[126]), .A(n40), .Z(n22226) );
  XNOR U22703 ( .A(n22234), .B(n22336), .Z(n22227) );
  XNOR U22704 ( .A(n22233), .B(n22231), .Z(n22336) );
  AND U22705 ( .A(n22337), .B(n22338), .Z(n22231) );
  NANDN U22706 ( .A(n22339), .B(n22340), .Z(n22338) );
  NAND U22707 ( .A(n22341), .B(n22342), .Z(n22340) );
  ANDN U22708 ( .B(B[127]), .A(n41), .Z(n22233) );
  XOR U22709 ( .A(n22240), .B(n22343), .Z(n22234) );
  XNOR U22710 ( .A(n22238), .B(n22241), .Z(n22343) );
  NAND U22711 ( .A(A[2]), .B(B[128]), .Z(n22241) );
  NANDN U22712 ( .A(n22344), .B(n22345), .Z(n22238) );
  AND U22713 ( .A(A[0]), .B(B[129]), .Z(n22345) );
  XNOR U22714 ( .A(n22243), .B(n22346), .Z(n22240) );
  NAND U22715 ( .A(A[0]), .B(B[130]), .Z(n22346) );
  NAND U22716 ( .A(B[129]), .B(A[1]), .Z(n22243) );
  NAND U22717 ( .A(n22347), .B(n22348), .Z(n495) );
  NANDN U22718 ( .A(n22349), .B(n22350), .Z(n22348) );
  OR U22719 ( .A(n22351), .B(n22352), .Z(n22350) );
  NAND U22720 ( .A(n22352), .B(n22351), .Z(n22347) );
  XOR U22721 ( .A(n497), .B(n496), .Z(\A1[127] ) );
  XOR U22722 ( .A(n22352), .B(n22353), .Z(n496) );
  XNOR U22723 ( .A(n22351), .B(n22349), .Z(n22353) );
  AND U22724 ( .A(n22354), .B(n22355), .Z(n22349) );
  NANDN U22725 ( .A(n22356), .B(n22357), .Z(n22355) );
  NANDN U22726 ( .A(n22358), .B(n22359), .Z(n22357) );
  NANDN U22727 ( .A(n22359), .B(n22358), .Z(n22354) );
  ANDN U22728 ( .B(B[114]), .A(n29), .Z(n22351) );
  XNOR U22729 ( .A(n22258), .B(n22360), .Z(n22352) );
  XNOR U22730 ( .A(n22257), .B(n22255), .Z(n22360) );
  AND U22731 ( .A(n22361), .B(n22362), .Z(n22255) );
  NANDN U22732 ( .A(n22363), .B(n22364), .Z(n22362) );
  OR U22733 ( .A(n22365), .B(n22366), .Z(n22364) );
  NAND U22734 ( .A(n22366), .B(n22365), .Z(n22361) );
  ANDN U22735 ( .B(B[115]), .A(n30), .Z(n22257) );
  XNOR U22736 ( .A(n22265), .B(n22367), .Z(n22258) );
  XNOR U22737 ( .A(n22264), .B(n22262), .Z(n22367) );
  AND U22738 ( .A(n22368), .B(n22369), .Z(n22262) );
  NANDN U22739 ( .A(n22370), .B(n22371), .Z(n22369) );
  NANDN U22740 ( .A(n22372), .B(n22373), .Z(n22371) );
  NANDN U22741 ( .A(n22373), .B(n22372), .Z(n22368) );
  ANDN U22742 ( .B(B[116]), .A(n31), .Z(n22264) );
  XNOR U22743 ( .A(n22272), .B(n22374), .Z(n22265) );
  XNOR U22744 ( .A(n22271), .B(n22269), .Z(n22374) );
  AND U22745 ( .A(n22375), .B(n22376), .Z(n22269) );
  NANDN U22746 ( .A(n22377), .B(n22378), .Z(n22376) );
  OR U22747 ( .A(n22379), .B(n22380), .Z(n22378) );
  NAND U22748 ( .A(n22380), .B(n22379), .Z(n22375) );
  ANDN U22749 ( .B(B[117]), .A(n32), .Z(n22271) );
  XNOR U22750 ( .A(n22279), .B(n22381), .Z(n22272) );
  XNOR U22751 ( .A(n22278), .B(n22276), .Z(n22381) );
  AND U22752 ( .A(n22382), .B(n22383), .Z(n22276) );
  NANDN U22753 ( .A(n22384), .B(n22385), .Z(n22383) );
  NANDN U22754 ( .A(n22386), .B(n22387), .Z(n22385) );
  NANDN U22755 ( .A(n22387), .B(n22386), .Z(n22382) );
  ANDN U22756 ( .B(B[118]), .A(n33), .Z(n22278) );
  XNOR U22757 ( .A(n22286), .B(n22388), .Z(n22279) );
  XNOR U22758 ( .A(n22285), .B(n22283), .Z(n22388) );
  AND U22759 ( .A(n22389), .B(n22390), .Z(n22283) );
  NANDN U22760 ( .A(n22391), .B(n22392), .Z(n22390) );
  OR U22761 ( .A(n22393), .B(n22394), .Z(n22392) );
  NAND U22762 ( .A(n22394), .B(n22393), .Z(n22389) );
  ANDN U22763 ( .B(B[119]), .A(n34), .Z(n22285) );
  XNOR U22764 ( .A(n22293), .B(n22395), .Z(n22286) );
  XNOR U22765 ( .A(n22292), .B(n22290), .Z(n22395) );
  AND U22766 ( .A(n22396), .B(n22397), .Z(n22290) );
  NANDN U22767 ( .A(n22398), .B(n22399), .Z(n22397) );
  NANDN U22768 ( .A(n22400), .B(n22401), .Z(n22399) );
  NANDN U22769 ( .A(n22401), .B(n22400), .Z(n22396) );
  ANDN U22770 ( .B(B[120]), .A(n35), .Z(n22292) );
  XNOR U22771 ( .A(n22300), .B(n22402), .Z(n22293) );
  XNOR U22772 ( .A(n22299), .B(n22297), .Z(n22402) );
  AND U22773 ( .A(n22403), .B(n22404), .Z(n22297) );
  NANDN U22774 ( .A(n22405), .B(n22406), .Z(n22404) );
  OR U22775 ( .A(n22407), .B(n22408), .Z(n22406) );
  NAND U22776 ( .A(n22408), .B(n22407), .Z(n22403) );
  ANDN U22777 ( .B(B[121]), .A(n36), .Z(n22299) );
  XNOR U22778 ( .A(n22307), .B(n22409), .Z(n22300) );
  XNOR U22779 ( .A(n22306), .B(n22304), .Z(n22409) );
  AND U22780 ( .A(n22410), .B(n22411), .Z(n22304) );
  NANDN U22781 ( .A(n22412), .B(n22413), .Z(n22411) );
  NANDN U22782 ( .A(n22414), .B(n22415), .Z(n22413) );
  NANDN U22783 ( .A(n22415), .B(n22414), .Z(n22410) );
  ANDN U22784 ( .B(B[122]), .A(n37), .Z(n22306) );
  XNOR U22785 ( .A(n22314), .B(n22416), .Z(n22307) );
  XNOR U22786 ( .A(n22313), .B(n22311), .Z(n22416) );
  AND U22787 ( .A(n22417), .B(n22418), .Z(n22311) );
  NANDN U22788 ( .A(n22419), .B(n22420), .Z(n22418) );
  OR U22789 ( .A(n22421), .B(n22422), .Z(n22420) );
  NAND U22790 ( .A(n22422), .B(n22421), .Z(n22417) );
  ANDN U22791 ( .B(B[123]), .A(n38), .Z(n22313) );
  XNOR U22792 ( .A(n22321), .B(n22423), .Z(n22314) );
  XNOR U22793 ( .A(n22320), .B(n22318), .Z(n22423) );
  AND U22794 ( .A(n22424), .B(n22425), .Z(n22318) );
  NANDN U22795 ( .A(n22426), .B(n22427), .Z(n22425) );
  NANDN U22796 ( .A(n22428), .B(n22429), .Z(n22427) );
  NANDN U22797 ( .A(n22429), .B(n22428), .Z(n22424) );
  ANDN U22798 ( .B(B[124]), .A(n39), .Z(n22320) );
  XNOR U22799 ( .A(n22328), .B(n22430), .Z(n22321) );
  XNOR U22800 ( .A(n22327), .B(n22325), .Z(n22430) );
  AND U22801 ( .A(n22431), .B(n22432), .Z(n22325) );
  NANDN U22802 ( .A(n22433), .B(n22434), .Z(n22432) );
  OR U22803 ( .A(n22435), .B(n22436), .Z(n22434) );
  NAND U22804 ( .A(n22436), .B(n22435), .Z(n22431) );
  ANDN U22805 ( .B(B[125]), .A(n40), .Z(n22327) );
  XNOR U22806 ( .A(n22335), .B(n22437), .Z(n22328) );
  XNOR U22807 ( .A(n22334), .B(n22332), .Z(n22437) );
  AND U22808 ( .A(n22438), .B(n22439), .Z(n22332) );
  NANDN U22809 ( .A(n22440), .B(n22441), .Z(n22439) );
  NAND U22810 ( .A(n22442), .B(n22443), .Z(n22441) );
  ANDN U22811 ( .B(B[126]), .A(n41), .Z(n22334) );
  XOR U22812 ( .A(n22341), .B(n22444), .Z(n22335) );
  XNOR U22813 ( .A(n22339), .B(n22342), .Z(n22444) );
  NAND U22814 ( .A(A[2]), .B(B[127]), .Z(n22342) );
  NANDN U22815 ( .A(n22445), .B(n22446), .Z(n22339) );
  AND U22816 ( .A(A[0]), .B(B[128]), .Z(n22446) );
  XNOR U22817 ( .A(n22344), .B(n22447), .Z(n22341) );
  NAND U22818 ( .A(A[0]), .B(B[129]), .Z(n22447) );
  NAND U22819 ( .A(B[128]), .B(A[1]), .Z(n22344) );
  NAND U22820 ( .A(n22448), .B(n22449), .Z(n497) );
  NANDN U22821 ( .A(n22450), .B(n22451), .Z(n22449) );
  OR U22822 ( .A(n22452), .B(n22453), .Z(n22451) );
  NAND U22823 ( .A(n22453), .B(n22452), .Z(n22448) );
  XOR U22824 ( .A(n499), .B(n498), .Z(\A1[126] ) );
  XOR U22825 ( .A(n22453), .B(n22454), .Z(n498) );
  XNOR U22826 ( .A(n22452), .B(n22450), .Z(n22454) );
  AND U22827 ( .A(n22455), .B(n22456), .Z(n22450) );
  NANDN U22828 ( .A(n22457), .B(n22458), .Z(n22456) );
  NANDN U22829 ( .A(n22459), .B(n22460), .Z(n22458) );
  NANDN U22830 ( .A(n22460), .B(n22459), .Z(n22455) );
  ANDN U22831 ( .B(B[113]), .A(n29), .Z(n22452) );
  XNOR U22832 ( .A(n22359), .B(n22461), .Z(n22453) );
  XNOR U22833 ( .A(n22358), .B(n22356), .Z(n22461) );
  AND U22834 ( .A(n22462), .B(n22463), .Z(n22356) );
  NANDN U22835 ( .A(n22464), .B(n22465), .Z(n22463) );
  OR U22836 ( .A(n22466), .B(n22467), .Z(n22465) );
  NAND U22837 ( .A(n22467), .B(n22466), .Z(n22462) );
  ANDN U22838 ( .B(B[114]), .A(n30), .Z(n22358) );
  XNOR U22839 ( .A(n22366), .B(n22468), .Z(n22359) );
  XNOR U22840 ( .A(n22365), .B(n22363), .Z(n22468) );
  AND U22841 ( .A(n22469), .B(n22470), .Z(n22363) );
  NANDN U22842 ( .A(n22471), .B(n22472), .Z(n22470) );
  NANDN U22843 ( .A(n22473), .B(n22474), .Z(n22472) );
  NANDN U22844 ( .A(n22474), .B(n22473), .Z(n22469) );
  ANDN U22845 ( .B(B[115]), .A(n31), .Z(n22365) );
  XNOR U22846 ( .A(n22373), .B(n22475), .Z(n22366) );
  XNOR U22847 ( .A(n22372), .B(n22370), .Z(n22475) );
  AND U22848 ( .A(n22476), .B(n22477), .Z(n22370) );
  NANDN U22849 ( .A(n22478), .B(n22479), .Z(n22477) );
  OR U22850 ( .A(n22480), .B(n22481), .Z(n22479) );
  NAND U22851 ( .A(n22481), .B(n22480), .Z(n22476) );
  ANDN U22852 ( .B(B[116]), .A(n32), .Z(n22372) );
  XNOR U22853 ( .A(n22380), .B(n22482), .Z(n22373) );
  XNOR U22854 ( .A(n22379), .B(n22377), .Z(n22482) );
  AND U22855 ( .A(n22483), .B(n22484), .Z(n22377) );
  NANDN U22856 ( .A(n22485), .B(n22486), .Z(n22484) );
  NANDN U22857 ( .A(n22487), .B(n22488), .Z(n22486) );
  NANDN U22858 ( .A(n22488), .B(n22487), .Z(n22483) );
  ANDN U22859 ( .B(B[117]), .A(n33), .Z(n22379) );
  XNOR U22860 ( .A(n22387), .B(n22489), .Z(n22380) );
  XNOR U22861 ( .A(n22386), .B(n22384), .Z(n22489) );
  AND U22862 ( .A(n22490), .B(n22491), .Z(n22384) );
  NANDN U22863 ( .A(n22492), .B(n22493), .Z(n22491) );
  OR U22864 ( .A(n22494), .B(n22495), .Z(n22493) );
  NAND U22865 ( .A(n22495), .B(n22494), .Z(n22490) );
  ANDN U22866 ( .B(B[118]), .A(n34), .Z(n22386) );
  XNOR U22867 ( .A(n22394), .B(n22496), .Z(n22387) );
  XNOR U22868 ( .A(n22393), .B(n22391), .Z(n22496) );
  AND U22869 ( .A(n22497), .B(n22498), .Z(n22391) );
  NANDN U22870 ( .A(n22499), .B(n22500), .Z(n22498) );
  NANDN U22871 ( .A(n22501), .B(n22502), .Z(n22500) );
  NANDN U22872 ( .A(n22502), .B(n22501), .Z(n22497) );
  ANDN U22873 ( .B(B[119]), .A(n35), .Z(n22393) );
  XNOR U22874 ( .A(n22401), .B(n22503), .Z(n22394) );
  XNOR U22875 ( .A(n22400), .B(n22398), .Z(n22503) );
  AND U22876 ( .A(n22504), .B(n22505), .Z(n22398) );
  NANDN U22877 ( .A(n22506), .B(n22507), .Z(n22505) );
  OR U22878 ( .A(n22508), .B(n22509), .Z(n22507) );
  NAND U22879 ( .A(n22509), .B(n22508), .Z(n22504) );
  ANDN U22880 ( .B(B[120]), .A(n36), .Z(n22400) );
  XNOR U22881 ( .A(n22408), .B(n22510), .Z(n22401) );
  XNOR U22882 ( .A(n22407), .B(n22405), .Z(n22510) );
  AND U22883 ( .A(n22511), .B(n22512), .Z(n22405) );
  NANDN U22884 ( .A(n22513), .B(n22514), .Z(n22512) );
  NANDN U22885 ( .A(n22515), .B(n22516), .Z(n22514) );
  NANDN U22886 ( .A(n22516), .B(n22515), .Z(n22511) );
  ANDN U22887 ( .B(B[121]), .A(n37), .Z(n22407) );
  XNOR U22888 ( .A(n22415), .B(n22517), .Z(n22408) );
  XNOR U22889 ( .A(n22414), .B(n22412), .Z(n22517) );
  AND U22890 ( .A(n22518), .B(n22519), .Z(n22412) );
  NANDN U22891 ( .A(n22520), .B(n22521), .Z(n22519) );
  OR U22892 ( .A(n22522), .B(n22523), .Z(n22521) );
  NAND U22893 ( .A(n22523), .B(n22522), .Z(n22518) );
  ANDN U22894 ( .B(B[122]), .A(n38), .Z(n22414) );
  XNOR U22895 ( .A(n22422), .B(n22524), .Z(n22415) );
  XNOR U22896 ( .A(n22421), .B(n22419), .Z(n22524) );
  AND U22897 ( .A(n22525), .B(n22526), .Z(n22419) );
  NANDN U22898 ( .A(n22527), .B(n22528), .Z(n22526) );
  NANDN U22899 ( .A(n22529), .B(n22530), .Z(n22528) );
  NANDN U22900 ( .A(n22530), .B(n22529), .Z(n22525) );
  ANDN U22901 ( .B(B[123]), .A(n39), .Z(n22421) );
  XNOR U22902 ( .A(n22429), .B(n22531), .Z(n22422) );
  XNOR U22903 ( .A(n22428), .B(n22426), .Z(n22531) );
  AND U22904 ( .A(n22532), .B(n22533), .Z(n22426) );
  NANDN U22905 ( .A(n22534), .B(n22535), .Z(n22533) );
  OR U22906 ( .A(n22536), .B(n22537), .Z(n22535) );
  NAND U22907 ( .A(n22537), .B(n22536), .Z(n22532) );
  ANDN U22908 ( .B(B[124]), .A(n40), .Z(n22428) );
  XNOR U22909 ( .A(n22436), .B(n22538), .Z(n22429) );
  XNOR U22910 ( .A(n22435), .B(n22433), .Z(n22538) );
  AND U22911 ( .A(n22539), .B(n22540), .Z(n22433) );
  NANDN U22912 ( .A(n22541), .B(n22542), .Z(n22540) );
  NAND U22913 ( .A(n22543), .B(n22544), .Z(n22542) );
  ANDN U22914 ( .B(B[125]), .A(n41), .Z(n22435) );
  XOR U22915 ( .A(n22442), .B(n22545), .Z(n22436) );
  XNOR U22916 ( .A(n22440), .B(n22443), .Z(n22545) );
  NAND U22917 ( .A(A[2]), .B(B[126]), .Z(n22443) );
  NANDN U22918 ( .A(n22546), .B(n22547), .Z(n22440) );
  AND U22919 ( .A(A[0]), .B(B[127]), .Z(n22547) );
  XNOR U22920 ( .A(n22445), .B(n22548), .Z(n22442) );
  NAND U22921 ( .A(A[0]), .B(B[128]), .Z(n22548) );
  NAND U22922 ( .A(B[127]), .B(A[1]), .Z(n22445) );
  NAND U22923 ( .A(n22549), .B(n22550), .Z(n499) );
  NANDN U22924 ( .A(n22551), .B(n22552), .Z(n22550) );
  OR U22925 ( .A(n22553), .B(n22554), .Z(n22552) );
  NAND U22926 ( .A(n22554), .B(n22553), .Z(n22549) );
  XOR U22927 ( .A(n501), .B(n500), .Z(\A1[125] ) );
  XOR U22928 ( .A(n22554), .B(n22555), .Z(n500) );
  XNOR U22929 ( .A(n22553), .B(n22551), .Z(n22555) );
  AND U22930 ( .A(n22556), .B(n22557), .Z(n22551) );
  NANDN U22931 ( .A(n22558), .B(n22559), .Z(n22557) );
  NANDN U22932 ( .A(n22560), .B(n22561), .Z(n22559) );
  NANDN U22933 ( .A(n22561), .B(n22560), .Z(n22556) );
  ANDN U22934 ( .B(B[112]), .A(n29), .Z(n22553) );
  XNOR U22935 ( .A(n22460), .B(n22562), .Z(n22554) );
  XNOR U22936 ( .A(n22459), .B(n22457), .Z(n22562) );
  AND U22937 ( .A(n22563), .B(n22564), .Z(n22457) );
  NANDN U22938 ( .A(n22565), .B(n22566), .Z(n22564) );
  OR U22939 ( .A(n22567), .B(n22568), .Z(n22566) );
  NAND U22940 ( .A(n22568), .B(n22567), .Z(n22563) );
  ANDN U22941 ( .B(B[113]), .A(n30), .Z(n22459) );
  XNOR U22942 ( .A(n22467), .B(n22569), .Z(n22460) );
  XNOR U22943 ( .A(n22466), .B(n22464), .Z(n22569) );
  AND U22944 ( .A(n22570), .B(n22571), .Z(n22464) );
  NANDN U22945 ( .A(n22572), .B(n22573), .Z(n22571) );
  NANDN U22946 ( .A(n22574), .B(n22575), .Z(n22573) );
  NANDN U22947 ( .A(n22575), .B(n22574), .Z(n22570) );
  ANDN U22948 ( .B(B[114]), .A(n31), .Z(n22466) );
  XNOR U22949 ( .A(n22474), .B(n22576), .Z(n22467) );
  XNOR U22950 ( .A(n22473), .B(n22471), .Z(n22576) );
  AND U22951 ( .A(n22577), .B(n22578), .Z(n22471) );
  NANDN U22952 ( .A(n22579), .B(n22580), .Z(n22578) );
  OR U22953 ( .A(n22581), .B(n22582), .Z(n22580) );
  NAND U22954 ( .A(n22582), .B(n22581), .Z(n22577) );
  ANDN U22955 ( .B(B[115]), .A(n32), .Z(n22473) );
  XNOR U22956 ( .A(n22481), .B(n22583), .Z(n22474) );
  XNOR U22957 ( .A(n22480), .B(n22478), .Z(n22583) );
  AND U22958 ( .A(n22584), .B(n22585), .Z(n22478) );
  NANDN U22959 ( .A(n22586), .B(n22587), .Z(n22585) );
  NANDN U22960 ( .A(n22588), .B(n22589), .Z(n22587) );
  NANDN U22961 ( .A(n22589), .B(n22588), .Z(n22584) );
  ANDN U22962 ( .B(B[116]), .A(n33), .Z(n22480) );
  XNOR U22963 ( .A(n22488), .B(n22590), .Z(n22481) );
  XNOR U22964 ( .A(n22487), .B(n22485), .Z(n22590) );
  AND U22965 ( .A(n22591), .B(n22592), .Z(n22485) );
  NANDN U22966 ( .A(n22593), .B(n22594), .Z(n22592) );
  OR U22967 ( .A(n22595), .B(n22596), .Z(n22594) );
  NAND U22968 ( .A(n22596), .B(n22595), .Z(n22591) );
  ANDN U22969 ( .B(B[117]), .A(n34), .Z(n22487) );
  XNOR U22970 ( .A(n22495), .B(n22597), .Z(n22488) );
  XNOR U22971 ( .A(n22494), .B(n22492), .Z(n22597) );
  AND U22972 ( .A(n22598), .B(n22599), .Z(n22492) );
  NANDN U22973 ( .A(n22600), .B(n22601), .Z(n22599) );
  NANDN U22974 ( .A(n22602), .B(n22603), .Z(n22601) );
  NANDN U22975 ( .A(n22603), .B(n22602), .Z(n22598) );
  ANDN U22976 ( .B(B[118]), .A(n35), .Z(n22494) );
  XNOR U22977 ( .A(n22502), .B(n22604), .Z(n22495) );
  XNOR U22978 ( .A(n22501), .B(n22499), .Z(n22604) );
  AND U22979 ( .A(n22605), .B(n22606), .Z(n22499) );
  NANDN U22980 ( .A(n22607), .B(n22608), .Z(n22606) );
  OR U22981 ( .A(n22609), .B(n22610), .Z(n22608) );
  NAND U22982 ( .A(n22610), .B(n22609), .Z(n22605) );
  ANDN U22983 ( .B(B[119]), .A(n36), .Z(n22501) );
  XNOR U22984 ( .A(n22509), .B(n22611), .Z(n22502) );
  XNOR U22985 ( .A(n22508), .B(n22506), .Z(n22611) );
  AND U22986 ( .A(n22612), .B(n22613), .Z(n22506) );
  NANDN U22987 ( .A(n22614), .B(n22615), .Z(n22613) );
  NANDN U22988 ( .A(n22616), .B(n22617), .Z(n22615) );
  NANDN U22989 ( .A(n22617), .B(n22616), .Z(n22612) );
  ANDN U22990 ( .B(B[120]), .A(n37), .Z(n22508) );
  XNOR U22991 ( .A(n22516), .B(n22618), .Z(n22509) );
  XNOR U22992 ( .A(n22515), .B(n22513), .Z(n22618) );
  AND U22993 ( .A(n22619), .B(n22620), .Z(n22513) );
  NANDN U22994 ( .A(n22621), .B(n22622), .Z(n22620) );
  OR U22995 ( .A(n22623), .B(n22624), .Z(n22622) );
  NAND U22996 ( .A(n22624), .B(n22623), .Z(n22619) );
  ANDN U22997 ( .B(B[121]), .A(n38), .Z(n22515) );
  XNOR U22998 ( .A(n22523), .B(n22625), .Z(n22516) );
  XNOR U22999 ( .A(n22522), .B(n22520), .Z(n22625) );
  AND U23000 ( .A(n22626), .B(n22627), .Z(n22520) );
  NANDN U23001 ( .A(n22628), .B(n22629), .Z(n22627) );
  NANDN U23002 ( .A(n22630), .B(n22631), .Z(n22629) );
  NANDN U23003 ( .A(n22631), .B(n22630), .Z(n22626) );
  ANDN U23004 ( .B(B[122]), .A(n39), .Z(n22522) );
  XNOR U23005 ( .A(n22530), .B(n22632), .Z(n22523) );
  XNOR U23006 ( .A(n22529), .B(n22527), .Z(n22632) );
  AND U23007 ( .A(n22633), .B(n22634), .Z(n22527) );
  NANDN U23008 ( .A(n22635), .B(n22636), .Z(n22634) );
  OR U23009 ( .A(n22637), .B(n22638), .Z(n22636) );
  NAND U23010 ( .A(n22638), .B(n22637), .Z(n22633) );
  ANDN U23011 ( .B(B[123]), .A(n40), .Z(n22529) );
  XNOR U23012 ( .A(n22537), .B(n22639), .Z(n22530) );
  XNOR U23013 ( .A(n22536), .B(n22534), .Z(n22639) );
  AND U23014 ( .A(n22640), .B(n22641), .Z(n22534) );
  NANDN U23015 ( .A(n22642), .B(n22643), .Z(n22641) );
  NAND U23016 ( .A(n22644), .B(n22645), .Z(n22643) );
  ANDN U23017 ( .B(B[124]), .A(n41), .Z(n22536) );
  XOR U23018 ( .A(n22543), .B(n22646), .Z(n22537) );
  XNOR U23019 ( .A(n22541), .B(n22544), .Z(n22646) );
  NAND U23020 ( .A(A[2]), .B(B[125]), .Z(n22544) );
  NANDN U23021 ( .A(n22647), .B(n22648), .Z(n22541) );
  AND U23022 ( .A(A[0]), .B(B[126]), .Z(n22648) );
  XNOR U23023 ( .A(n22546), .B(n22649), .Z(n22543) );
  NAND U23024 ( .A(A[0]), .B(B[127]), .Z(n22649) );
  NAND U23025 ( .A(B[126]), .B(A[1]), .Z(n22546) );
  NAND U23026 ( .A(n22650), .B(n22651), .Z(n501) );
  NANDN U23027 ( .A(n22652), .B(n22653), .Z(n22651) );
  OR U23028 ( .A(n22654), .B(n22655), .Z(n22653) );
  NAND U23029 ( .A(n22655), .B(n22654), .Z(n22650) );
  XOR U23030 ( .A(n503), .B(n502), .Z(\A1[124] ) );
  XOR U23031 ( .A(n22655), .B(n22656), .Z(n502) );
  XNOR U23032 ( .A(n22654), .B(n22652), .Z(n22656) );
  AND U23033 ( .A(n22657), .B(n22658), .Z(n22652) );
  NANDN U23034 ( .A(n22659), .B(n22660), .Z(n22658) );
  NANDN U23035 ( .A(n22661), .B(n22662), .Z(n22660) );
  NANDN U23036 ( .A(n22662), .B(n22661), .Z(n22657) );
  ANDN U23037 ( .B(B[111]), .A(n29), .Z(n22654) );
  XNOR U23038 ( .A(n22561), .B(n22663), .Z(n22655) );
  XNOR U23039 ( .A(n22560), .B(n22558), .Z(n22663) );
  AND U23040 ( .A(n22664), .B(n22665), .Z(n22558) );
  NANDN U23041 ( .A(n22666), .B(n22667), .Z(n22665) );
  OR U23042 ( .A(n22668), .B(n22669), .Z(n22667) );
  NAND U23043 ( .A(n22669), .B(n22668), .Z(n22664) );
  ANDN U23044 ( .B(B[112]), .A(n30), .Z(n22560) );
  XNOR U23045 ( .A(n22568), .B(n22670), .Z(n22561) );
  XNOR U23046 ( .A(n22567), .B(n22565), .Z(n22670) );
  AND U23047 ( .A(n22671), .B(n22672), .Z(n22565) );
  NANDN U23048 ( .A(n22673), .B(n22674), .Z(n22672) );
  NANDN U23049 ( .A(n22675), .B(n22676), .Z(n22674) );
  NANDN U23050 ( .A(n22676), .B(n22675), .Z(n22671) );
  ANDN U23051 ( .B(B[113]), .A(n31), .Z(n22567) );
  XNOR U23052 ( .A(n22575), .B(n22677), .Z(n22568) );
  XNOR U23053 ( .A(n22574), .B(n22572), .Z(n22677) );
  AND U23054 ( .A(n22678), .B(n22679), .Z(n22572) );
  NANDN U23055 ( .A(n22680), .B(n22681), .Z(n22679) );
  OR U23056 ( .A(n22682), .B(n22683), .Z(n22681) );
  NAND U23057 ( .A(n22683), .B(n22682), .Z(n22678) );
  ANDN U23058 ( .B(B[114]), .A(n32), .Z(n22574) );
  XNOR U23059 ( .A(n22582), .B(n22684), .Z(n22575) );
  XNOR U23060 ( .A(n22581), .B(n22579), .Z(n22684) );
  AND U23061 ( .A(n22685), .B(n22686), .Z(n22579) );
  NANDN U23062 ( .A(n22687), .B(n22688), .Z(n22686) );
  NANDN U23063 ( .A(n22689), .B(n22690), .Z(n22688) );
  NANDN U23064 ( .A(n22690), .B(n22689), .Z(n22685) );
  ANDN U23065 ( .B(B[115]), .A(n33), .Z(n22581) );
  XNOR U23066 ( .A(n22589), .B(n22691), .Z(n22582) );
  XNOR U23067 ( .A(n22588), .B(n22586), .Z(n22691) );
  AND U23068 ( .A(n22692), .B(n22693), .Z(n22586) );
  NANDN U23069 ( .A(n22694), .B(n22695), .Z(n22693) );
  OR U23070 ( .A(n22696), .B(n22697), .Z(n22695) );
  NAND U23071 ( .A(n22697), .B(n22696), .Z(n22692) );
  ANDN U23072 ( .B(B[116]), .A(n34), .Z(n22588) );
  XNOR U23073 ( .A(n22596), .B(n22698), .Z(n22589) );
  XNOR U23074 ( .A(n22595), .B(n22593), .Z(n22698) );
  AND U23075 ( .A(n22699), .B(n22700), .Z(n22593) );
  NANDN U23076 ( .A(n22701), .B(n22702), .Z(n22700) );
  NANDN U23077 ( .A(n22703), .B(n22704), .Z(n22702) );
  NANDN U23078 ( .A(n22704), .B(n22703), .Z(n22699) );
  ANDN U23079 ( .B(B[117]), .A(n35), .Z(n22595) );
  XNOR U23080 ( .A(n22603), .B(n22705), .Z(n22596) );
  XNOR U23081 ( .A(n22602), .B(n22600), .Z(n22705) );
  AND U23082 ( .A(n22706), .B(n22707), .Z(n22600) );
  NANDN U23083 ( .A(n22708), .B(n22709), .Z(n22707) );
  OR U23084 ( .A(n22710), .B(n22711), .Z(n22709) );
  NAND U23085 ( .A(n22711), .B(n22710), .Z(n22706) );
  ANDN U23086 ( .B(B[118]), .A(n36), .Z(n22602) );
  XNOR U23087 ( .A(n22610), .B(n22712), .Z(n22603) );
  XNOR U23088 ( .A(n22609), .B(n22607), .Z(n22712) );
  AND U23089 ( .A(n22713), .B(n22714), .Z(n22607) );
  NANDN U23090 ( .A(n22715), .B(n22716), .Z(n22714) );
  NANDN U23091 ( .A(n22717), .B(n22718), .Z(n22716) );
  NANDN U23092 ( .A(n22718), .B(n22717), .Z(n22713) );
  ANDN U23093 ( .B(B[119]), .A(n37), .Z(n22609) );
  XNOR U23094 ( .A(n22617), .B(n22719), .Z(n22610) );
  XNOR U23095 ( .A(n22616), .B(n22614), .Z(n22719) );
  AND U23096 ( .A(n22720), .B(n22721), .Z(n22614) );
  NANDN U23097 ( .A(n22722), .B(n22723), .Z(n22721) );
  OR U23098 ( .A(n22724), .B(n22725), .Z(n22723) );
  NAND U23099 ( .A(n22725), .B(n22724), .Z(n22720) );
  ANDN U23100 ( .B(B[120]), .A(n38), .Z(n22616) );
  XNOR U23101 ( .A(n22624), .B(n22726), .Z(n22617) );
  XNOR U23102 ( .A(n22623), .B(n22621), .Z(n22726) );
  AND U23103 ( .A(n22727), .B(n22728), .Z(n22621) );
  NANDN U23104 ( .A(n22729), .B(n22730), .Z(n22728) );
  NANDN U23105 ( .A(n22731), .B(n22732), .Z(n22730) );
  NANDN U23106 ( .A(n22732), .B(n22731), .Z(n22727) );
  ANDN U23107 ( .B(B[121]), .A(n39), .Z(n22623) );
  XNOR U23108 ( .A(n22631), .B(n22733), .Z(n22624) );
  XNOR U23109 ( .A(n22630), .B(n22628), .Z(n22733) );
  AND U23110 ( .A(n22734), .B(n22735), .Z(n22628) );
  NANDN U23111 ( .A(n22736), .B(n22737), .Z(n22735) );
  OR U23112 ( .A(n22738), .B(n22739), .Z(n22737) );
  NAND U23113 ( .A(n22739), .B(n22738), .Z(n22734) );
  ANDN U23114 ( .B(B[122]), .A(n40), .Z(n22630) );
  XNOR U23115 ( .A(n22638), .B(n22740), .Z(n22631) );
  XNOR U23116 ( .A(n22637), .B(n22635), .Z(n22740) );
  AND U23117 ( .A(n22741), .B(n22742), .Z(n22635) );
  NANDN U23118 ( .A(n22743), .B(n22744), .Z(n22742) );
  NAND U23119 ( .A(n22745), .B(n22746), .Z(n22744) );
  ANDN U23120 ( .B(B[123]), .A(n41), .Z(n22637) );
  XOR U23121 ( .A(n22644), .B(n22747), .Z(n22638) );
  XNOR U23122 ( .A(n22642), .B(n22645), .Z(n22747) );
  NAND U23123 ( .A(A[2]), .B(B[124]), .Z(n22645) );
  NANDN U23124 ( .A(n22748), .B(n22749), .Z(n22642) );
  AND U23125 ( .A(A[0]), .B(B[125]), .Z(n22749) );
  XNOR U23126 ( .A(n22647), .B(n22750), .Z(n22644) );
  NAND U23127 ( .A(A[0]), .B(B[126]), .Z(n22750) );
  NAND U23128 ( .A(B[125]), .B(A[1]), .Z(n22647) );
  NAND U23129 ( .A(n22751), .B(n22752), .Z(n503) );
  NANDN U23130 ( .A(n22753), .B(n22754), .Z(n22752) );
  OR U23131 ( .A(n22755), .B(n22756), .Z(n22754) );
  NAND U23132 ( .A(n22756), .B(n22755), .Z(n22751) );
  XOR U23133 ( .A(n505), .B(n504), .Z(\A1[123] ) );
  XOR U23134 ( .A(n22756), .B(n22757), .Z(n504) );
  XNOR U23135 ( .A(n22755), .B(n22753), .Z(n22757) );
  AND U23136 ( .A(n22758), .B(n22759), .Z(n22753) );
  NANDN U23137 ( .A(n22760), .B(n22761), .Z(n22759) );
  NANDN U23138 ( .A(n22762), .B(n22763), .Z(n22761) );
  NANDN U23139 ( .A(n22763), .B(n22762), .Z(n22758) );
  ANDN U23140 ( .B(B[110]), .A(n29), .Z(n22755) );
  XNOR U23141 ( .A(n22662), .B(n22764), .Z(n22756) );
  XNOR U23142 ( .A(n22661), .B(n22659), .Z(n22764) );
  AND U23143 ( .A(n22765), .B(n22766), .Z(n22659) );
  NANDN U23144 ( .A(n22767), .B(n22768), .Z(n22766) );
  OR U23145 ( .A(n22769), .B(n22770), .Z(n22768) );
  NAND U23146 ( .A(n22770), .B(n22769), .Z(n22765) );
  ANDN U23147 ( .B(B[111]), .A(n30), .Z(n22661) );
  XNOR U23148 ( .A(n22669), .B(n22771), .Z(n22662) );
  XNOR U23149 ( .A(n22668), .B(n22666), .Z(n22771) );
  AND U23150 ( .A(n22772), .B(n22773), .Z(n22666) );
  NANDN U23151 ( .A(n22774), .B(n22775), .Z(n22773) );
  NANDN U23152 ( .A(n22776), .B(n22777), .Z(n22775) );
  NANDN U23153 ( .A(n22777), .B(n22776), .Z(n22772) );
  ANDN U23154 ( .B(B[112]), .A(n31), .Z(n22668) );
  XNOR U23155 ( .A(n22676), .B(n22778), .Z(n22669) );
  XNOR U23156 ( .A(n22675), .B(n22673), .Z(n22778) );
  AND U23157 ( .A(n22779), .B(n22780), .Z(n22673) );
  NANDN U23158 ( .A(n22781), .B(n22782), .Z(n22780) );
  OR U23159 ( .A(n22783), .B(n22784), .Z(n22782) );
  NAND U23160 ( .A(n22784), .B(n22783), .Z(n22779) );
  ANDN U23161 ( .B(B[113]), .A(n32), .Z(n22675) );
  XNOR U23162 ( .A(n22683), .B(n22785), .Z(n22676) );
  XNOR U23163 ( .A(n22682), .B(n22680), .Z(n22785) );
  AND U23164 ( .A(n22786), .B(n22787), .Z(n22680) );
  NANDN U23165 ( .A(n22788), .B(n22789), .Z(n22787) );
  NANDN U23166 ( .A(n22790), .B(n22791), .Z(n22789) );
  NANDN U23167 ( .A(n22791), .B(n22790), .Z(n22786) );
  ANDN U23168 ( .B(B[114]), .A(n33), .Z(n22682) );
  XNOR U23169 ( .A(n22690), .B(n22792), .Z(n22683) );
  XNOR U23170 ( .A(n22689), .B(n22687), .Z(n22792) );
  AND U23171 ( .A(n22793), .B(n22794), .Z(n22687) );
  NANDN U23172 ( .A(n22795), .B(n22796), .Z(n22794) );
  OR U23173 ( .A(n22797), .B(n22798), .Z(n22796) );
  NAND U23174 ( .A(n22798), .B(n22797), .Z(n22793) );
  ANDN U23175 ( .B(B[115]), .A(n34), .Z(n22689) );
  XNOR U23176 ( .A(n22697), .B(n22799), .Z(n22690) );
  XNOR U23177 ( .A(n22696), .B(n22694), .Z(n22799) );
  AND U23178 ( .A(n22800), .B(n22801), .Z(n22694) );
  NANDN U23179 ( .A(n22802), .B(n22803), .Z(n22801) );
  NANDN U23180 ( .A(n22804), .B(n22805), .Z(n22803) );
  NANDN U23181 ( .A(n22805), .B(n22804), .Z(n22800) );
  ANDN U23182 ( .B(B[116]), .A(n35), .Z(n22696) );
  XNOR U23183 ( .A(n22704), .B(n22806), .Z(n22697) );
  XNOR U23184 ( .A(n22703), .B(n22701), .Z(n22806) );
  AND U23185 ( .A(n22807), .B(n22808), .Z(n22701) );
  NANDN U23186 ( .A(n22809), .B(n22810), .Z(n22808) );
  OR U23187 ( .A(n22811), .B(n22812), .Z(n22810) );
  NAND U23188 ( .A(n22812), .B(n22811), .Z(n22807) );
  ANDN U23189 ( .B(B[117]), .A(n36), .Z(n22703) );
  XNOR U23190 ( .A(n22711), .B(n22813), .Z(n22704) );
  XNOR U23191 ( .A(n22710), .B(n22708), .Z(n22813) );
  AND U23192 ( .A(n22814), .B(n22815), .Z(n22708) );
  NANDN U23193 ( .A(n22816), .B(n22817), .Z(n22815) );
  NANDN U23194 ( .A(n22818), .B(n22819), .Z(n22817) );
  NANDN U23195 ( .A(n22819), .B(n22818), .Z(n22814) );
  ANDN U23196 ( .B(B[118]), .A(n37), .Z(n22710) );
  XNOR U23197 ( .A(n22718), .B(n22820), .Z(n22711) );
  XNOR U23198 ( .A(n22717), .B(n22715), .Z(n22820) );
  AND U23199 ( .A(n22821), .B(n22822), .Z(n22715) );
  NANDN U23200 ( .A(n22823), .B(n22824), .Z(n22822) );
  OR U23201 ( .A(n22825), .B(n22826), .Z(n22824) );
  NAND U23202 ( .A(n22826), .B(n22825), .Z(n22821) );
  ANDN U23203 ( .B(B[119]), .A(n38), .Z(n22717) );
  XNOR U23204 ( .A(n22725), .B(n22827), .Z(n22718) );
  XNOR U23205 ( .A(n22724), .B(n22722), .Z(n22827) );
  AND U23206 ( .A(n22828), .B(n22829), .Z(n22722) );
  NANDN U23207 ( .A(n22830), .B(n22831), .Z(n22829) );
  NANDN U23208 ( .A(n22832), .B(n22833), .Z(n22831) );
  NANDN U23209 ( .A(n22833), .B(n22832), .Z(n22828) );
  ANDN U23210 ( .B(B[120]), .A(n39), .Z(n22724) );
  XNOR U23211 ( .A(n22732), .B(n22834), .Z(n22725) );
  XNOR U23212 ( .A(n22731), .B(n22729), .Z(n22834) );
  AND U23213 ( .A(n22835), .B(n22836), .Z(n22729) );
  NANDN U23214 ( .A(n22837), .B(n22838), .Z(n22836) );
  OR U23215 ( .A(n22839), .B(n22840), .Z(n22838) );
  NAND U23216 ( .A(n22840), .B(n22839), .Z(n22835) );
  ANDN U23217 ( .B(B[121]), .A(n40), .Z(n22731) );
  XNOR U23218 ( .A(n22739), .B(n22841), .Z(n22732) );
  XNOR U23219 ( .A(n22738), .B(n22736), .Z(n22841) );
  AND U23220 ( .A(n22842), .B(n22843), .Z(n22736) );
  NANDN U23221 ( .A(n22844), .B(n22845), .Z(n22843) );
  NAND U23222 ( .A(n22846), .B(n22847), .Z(n22845) );
  ANDN U23223 ( .B(B[122]), .A(n41), .Z(n22738) );
  XOR U23224 ( .A(n22745), .B(n22848), .Z(n22739) );
  XNOR U23225 ( .A(n22743), .B(n22746), .Z(n22848) );
  NAND U23226 ( .A(A[2]), .B(B[123]), .Z(n22746) );
  NANDN U23227 ( .A(n22849), .B(n22850), .Z(n22743) );
  AND U23228 ( .A(A[0]), .B(B[124]), .Z(n22850) );
  XNOR U23229 ( .A(n22748), .B(n22851), .Z(n22745) );
  NAND U23230 ( .A(A[0]), .B(B[125]), .Z(n22851) );
  NAND U23231 ( .A(B[124]), .B(A[1]), .Z(n22748) );
  NAND U23232 ( .A(n22852), .B(n22853), .Z(n505) );
  NANDN U23233 ( .A(n22854), .B(n22855), .Z(n22853) );
  OR U23234 ( .A(n22856), .B(n22857), .Z(n22855) );
  NAND U23235 ( .A(n22857), .B(n22856), .Z(n22852) );
  XOR U23236 ( .A(n507), .B(n506), .Z(\A1[122] ) );
  XOR U23237 ( .A(n22857), .B(n22858), .Z(n506) );
  XNOR U23238 ( .A(n22856), .B(n22854), .Z(n22858) );
  AND U23239 ( .A(n22859), .B(n22860), .Z(n22854) );
  NANDN U23240 ( .A(n22861), .B(n22862), .Z(n22860) );
  NANDN U23241 ( .A(n22863), .B(n22864), .Z(n22862) );
  NANDN U23242 ( .A(n22864), .B(n22863), .Z(n22859) );
  ANDN U23243 ( .B(B[109]), .A(n29), .Z(n22856) );
  XNOR U23244 ( .A(n22763), .B(n22865), .Z(n22857) );
  XNOR U23245 ( .A(n22762), .B(n22760), .Z(n22865) );
  AND U23246 ( .A(n22866), .B(n22867), .Z(n22760) );
  NANDN U23247 ( .A(n22868), .B(n22869), .Z(n22867) );
  OR U23248 ( .A(n22870), .B(n22871), .Z(n22869) );
  NAND U23249 ( .A(n22871), .B(n22870), .Z(n22866) );
  ANDN U23250 ( .B(B[110]), .A(n30), .Z(n22762) );
  XNOR U23251 ( .A(n22770), .B(n22872), .Z(n22763) );
  XNOR U23252 ( .A(n22769), .B(n22767), .Z(n22872) );
  AND U23253 ( .A(n22873), .B(n22874), .Z(n22767) );
  NANDN U23254 ( .A(n22875), .B(n22876), .Z(n22874) );
  NANDN U23255 ( .A(n22877), .B(n22878), .Z(n22876) );
  NANDN U23256 ( .A(n22878), .B(n22877), .Z(n22873) );
  ANDN U23257 ( .B(B[111]), .A(n31), .Z(n22769) );
  XNOR U23258 ( .A(n22777), .B(n22879), .Z(n22770) );
  XNOR U23259 ( .A(n22776), .B(n22774), .Z(n22879) );
  AND U23260 ( .A(n22880), .B(n22881), .Z(n22774) );
  NANDN U23261 ( .A(n22882), .B(n22883), .Z(n22881) );
  OR U23262 ( .A(n22884), .B(n22885), .Z(n22883) );
  NAND U23263 ( .A(n22885), .B(n22884), .Z(n22880) );
  ANDN U23264 ( .B(B[112]), .A(n32), .Z(n22776) );
  XNOR U23265 ( .A(n22784), .B(n22886), .Z(n22777) );
  XNOR U23266 ( .A(n22783), .B(n22781), .Z(n22886) );
  AND U23267 ( .A(n22887), .B(n22888), .Z(n22781) );
  NANDN U23268 ( .A(n22889), .B(n22890), .Z(n22888) );
  NANDN U23269 ( .A(n22891), .B(n22892), .Z(n22890) );
  NANDN U23270 ( .A(n22892), .B(n22891), .Z(n22887) );
  ANDN U23271 ( .B(B[113]), .A(n33), .Z(n22783) );
  XNOR U23272 ( .A(n22791), .B(n22893), .Z(n22784) );
  XNOR U23273 ( .A(n22790), .B(n22788), .Z(n22893) );
  AND U23274 ( .A(n22894), .B(n22895), .Z(n22788) );
  NANDN U23275 ( .A(n22896), .B(n22897), .Z(n22895) );
  OR U23276 ( .A(n22898), .B(n22899), .Z(n22897) );
  NAND U23277 ( .A(n22899), .B(n22898), .Z(n22894) );
  ANDN U23278 ( .B(B[114]), .A(n34), .Z(n22790) );
  XNOR U23279 ( .A(n22798), .B(n22900), .Z(n22791) );
  XNOR U23280 ( .A(n22797), .B(n22795), .Z(n22900) );
  AND U23281 ( .A(n22901), .B(n22902), .Z(n22795) );
  NANDN U23282 ( .A(n22903), .B(n22904), .Z(n22902) );
  NANDN U23283 ( .A(n22905), .B(n22906), .Z(n22904) );
  NANDN U23284 ( .A(n22906), .B(n22905), .Z(n22901) );
  ANDN U23285 ( .B(B[115]), .A(n35), .Z(n22797) );
  XNOR U23286 ( .A(n22805), .B(n22907), .Z(n22798) );
  XNOR U23287 ( .A(n22804), .B(n22802), .Z(n22907) );
  AND U23288 ( .A(n22908), .B(n22909), .Z(n22802) );
  NANDN U23289 ( .A(n22910), .B(n22911), .Z(n22909) );
  OR U23290 ( .A(n22912), .B(n22913), .Z(n22911) );
  NAND U23291 ( .A(n22913), .B(n22912), .Z(n22908) );
  ANDN U23292 ( .B(B[116]), .A(n36), .Z(n22804) );
  XNOR U23293 ( .A(n22812), .B(n22914), .Z(n22805) );
  XNOR U23294 ( .A(n22811), .B(n22809), .Z(n22914) );
  AND U23295 ( .A(n22915), .B(n22916), .Z(n22809) );
  NANDN U23296 ( .A(n22917), .B(n22918), .Z(n22916) );
  NANDN U23297 ( .A(n22919), .B(n22920), .Z(n22918) );
  NANDN U23298 ( .A(n22920), .B(n22919), .Z(n22915) );
  ANDN U23299 ( .B(B[117]), .A(n37), .Z(n22811) );
  XNOR U23300 ( .A(n22819), .B(n22921), .Z(n22812) );
  XNOR U23301 ( .A(n22818), .B(n22816), .Z(n22921) );
  AND U23302 ( .A(n22922), .B(n22923), .Z(n22816) );
  NANDN U23303 ( .A(n22924), .B(n22925), .Z(n22923) );
  OR U23304 ( .A(n22926), .B(n22927), .Z(n22925) );
  NAND U23305 ( .A(n22927), .B(n22926), .Z(n22922) );
  ANDN U23306 ( .B(B[118]), .A(n38), .Z(n22818) );
  XNOR U23307 ( .A(n22826), .B(n22928), .Z(n22819) );
  XNOR U23308 ( .A(n22825), .B(n22823), .Z(n22928) );
  AND U23309 ( .A(n22929), .B(n22930), .Z(n22823) );
  NANDN U23310 ( .A(n22931), .B(n22932), .Z(n22930) );
  NANDN U23311 ( .A(n22933), .B(n22934), .Z(n22932) );
  NANDN U23312 ( .A(n22934), .B(n22933), .Z(n22929) );
  ANDN U23313 ( .B(B[119]), .A(n39), .Z(n22825) );
  XNOR U23314 ( .A(n22833), .B(n22935), .Z(n22826) );
  XNOR U23315 ( .A(n22832), .B(n22830), .Z(n22935) );
  AND U23316 ( .A(n22936), .B(n22937), .Z(n22830) );
  NANDN U23317 ( .A(n22938), .B(n22939), .Z(n22937) );
  OR U23318 ( .A(n22940), .B(n22941), .Z(n22939) );
  NAND U23319 ( .A(n22941), .B(n22940), .Z(n22936) );
  ANDN U23320 ( .B(B[120]), .A(n40), .Z(n22832) );
  XNOR U23321 ( .A(n22840), .B(n22942), .Z(n22833) );
  XNOR U23322 ( .A(n22839), .B(n22837), .Z(n22942) );
  AND U23323 ( .A(n22943), .B(n22944), .Z(n22837) );
  NANDN U23324 ( .A(n22945), .B(n22946), .Z(n22944) );
  NAND U23325 ( .A(n22947), .B(n22948), .Z(n22946) );
  ANDN U23326 ( .B(B[121]), .A(n41), .Z(n22839) );
  XOR U23327 ( .A(n22846), .B(n22949), .Z(n22840) );
  XNOR U23328 ( .A(n22844), .B(n22847), .Z(n22949) );
  NAND U23329 ( .A(A[2]), .B(B[122]), .Z(n22847) );
  NANDN U23330 ( .A(n22950), .B(n22951), .Z(n22844) );
  AND U23331 ( .A(A[0]), .B(B[123]), .Z(n22951) );
  XNOR U23332 ( .A(n22849), .B(n22952), .Z(n22846) );
  NAND U23333 ( .A(A[0]), .B(B[124]), .Z(n22952) );
  NAND U23334 ( .A(B[123]), .B(A[1]), .Z(n22849) );
  NAND U23335 ( .A(n22953), .B(n22954), .Z(n507) );
  NANDN U23336 ( .A(n22955), .B(n22956), .Z(n22954) );
  OR U23337 ( .A(n22957), .B(n22958), .Z(n22956) );
  NAND U23338 ( .A(n22958), .B(n22957), .Z(n22953) );
  XOR U23339 ( .A(n509), .B(n508), .Z(\A1[121] ) );
  XOR U23340 ( .A(n22958), .B(n22959), .Z(n508) );
  XNOR U23341 ( .A(n22957), .B(n22955), .Z(n22959) );
  AND U23342 ( .A(n22960), .B(n22961), .Z(n22955) );
  NANDN U23343 ( .A(n22962), .B(n22963), .Z(n22961) );
  NANDN U23344 ( .A(n22964), .B(n22965), .Z(n22963) );
  NANDN U23345 ( .A(n22965), .B(n22964), .Z(n22960) );
  ANDN U23346 ( .B(B[108]), .A(n29), .Z(n22957) );
  XNOR U23347 ( .A(n22864), .B(n22966), .Z(n22958) );
  XNOR U23348 ( .A(n22863), .B(n22861), .Z(n22966) );
  AND U23349 ( .A(n22967), .B(n22968), .Z(n22861) );
  NANDN U23350 ( .A(n22969), .B(n22970), .Z(n22968) );
  OR U23351 ( .A(n22971), .B(n22972), .Z(n22970) );
  NAND U23352 ( .A(n22972), .B(n22971), .Z(n22967) );
  ANDN U23353 ( .B(B[109]), .A(n30), .Z(n22863) );
  XNOR U23354 ( .A(n22871), .B(n22973), .Z(n22864) );
  XNOR U23355 ( .A(n22870), .B(n22868), .Z(n22973) );
  AND U23356 ( .A(n22974), .B(n22975), .Z(n22868) );
  NANDN U23357 ( .A(n22976), .B(n22977), .Z(n22975) );
  NANDN U23358 ( .A(n22978), .B(n22979), .Z(n22977) );
  NANDN U23359 ( .A(n22979), .B(n22978), .Z(n22974) );
  ANDN U23360 ( .B(B[110]), .A(n31), .Z(n22870) );
  XNOR U23361 ( .A(n22878), .B(n22980), .Z(n22871) );
  XNOR U23362 ( .A(n22877), .B(n22875), .Z(n22980) );
  AND U23363 ( .A(n22981), .B(n22982), .Z(n22875) );
  NANDN U23364 ( .A(n22983), .B(n22984), .Z(n22982) );
  OR U23365 ( .A(n22985), .B(n22986), .Z(n22984) );
  NAND U23366 ( .A(n22986), .B(n22985), .Z(n22981) );
  ANDN U23367 ( .B(B[111]), .A(n32), .Z(n22877) );
  XNOR U23368 ( .A(n22885), .B(n22987), .Z(n22878) );
  XNOR U23369 ( .A(n22884), .B(n22882), .Z(n22987) );
  AND U23370 ( .A(n22988), .B(n22989), .Z(n22882) );
  NANDN U23371 ( .A(n22990), .B(n22991), .Z(n22989) );
  NANDN U23372 ( .A(n22992), .B(n22993), .Z(n22991) );
  NANDN U23373 ( .A(n22993), .B(n22992), .Z(n22988) );
  ANDN U23374 ( .B(B[112]), .A(n33), .Z(n22884) );
  XNOR U23375 ( .A(n22892), .B(n22994), .Z(n22885) );
  XNOR U23376 ( .A(n22891), .B(n22889), .Z(n22994) );
  AND U23377 ( .A(n22995), .B(n22996), .Z(n22889) );
  NANDN U23378 ( .A(n22997), .B(n22998), .Z(n22996) );
  OR U23379 ( .A(n22999), .B(n23000), .Z(n22998) );
  NAND U23380 ( .A(n23000), .B(n22999), .Z(n22995) );
  ANDN U23381 ( .B(B[113]), .A(n34), .Z(n22891) );
  XNOR U23382 ( .A(n22899), .B(n23001), .Z(n22892) );
  XNOR U23383 ( .A(n22898), .B(n22896), .Z(n23001) );
  AND U23384 ( .A(n23002), .B(n23003), .Z(n22896) );
  NANDN U23385 ( .A(n23004), .B(n23005), .Z(n23003) );
  NANDN U23386 ( .A(n23006), .B(n23007), .Z(n23005) );
  NANDN U23387 ( .A(n23007), .B(n23006), .Z(n23002) );
  ANDN U23388 ( .B(B[114]), .A(n35), .Z(n22898) );
  XNOR U23389 ( .A(n22906), .B(n23008), .Z(n22899) );
  XNOR U23390 ( .A(n22905), .B(n22903), .Z(n23008) );
  AND U23391 ( .A(n23009), .B(n23010), .Z(n22903) );
  NANDN U23392 ( .A(n23011), .B(n23012), .Z(n23010) );
  OR U23393 ( .A(n23013), .B(n23014), .Z(n23012) );
  NAND U23394 ( .A(n23014), .B(n23013), .Z(n23009) );
  ANDN U23395 ( .B(B[115]), .A(n36), .Z(n22905) );
  XNOR U23396 ( .A(n22913), .B(n23015), .Z(n22906) );
  XNOR U23397 ( .A(n22912), .B(n22910), .Z(n23015) );
  AND U23398 ( .A(n23016), .B(n23017), .Z(n22910) );
  NANDN U23399 ( .A(n23018), .B(n23019), .Z(n23017) );
  NANDN U23400 ( .A(n23020), .B(n23021), .Z(n23019) );
  NANDN U23401 ( .A(n23021), .B(n23020), .Z(n23016) );
  ANDN U23402 ( .B(B[116]), .A(n37), .Z(n22912) );
  XNOR U23403 ( .A(n22920), .B(n23022), .Z(n22913) );
  XNOR U23404 ( .A(n22919), .B(n22917), .Z(n23022) );
  AND U23405 ( .A(n23023), .B(n23024), .Z(n22917) );
  NANDN U23406 ( .A(n23025), .B(n23026), .Z(n23024) );
  OR U23407 ( .A(n23027), .B(n23028), .Z(n23026) );
  NAND U23408 ( .A(n23028), .B(n23027), .Z(n23023) );
  ANDN U23409 ( .B(B[117]), .A(n38), .Z(n22919) );
  XNOR U23410 ( .A(n22927), .B(n23029), .Z(n22920) );
  XNOR U23411 ( .A(n22926), .B(n22924), .Z(n23029) );
  AND U23412 ( .A(n23030), .B(n23031), .Z(n22924) );
  NANDN U23413 ( .A(n23032), .B(n23033), .Z(n23031) );
  NANDN U23414 ( .A(n23034), .B(n23035), .Z(n23033) );
  NANDN U23415 ( .A(n23035), .B(n23034), .Z(n23030) );
  ANDN U23416 ( .B(B[118]), .A(n39), .Z(n22926) );
  XNOR U23417 ( .A(n22934), .B(n23036), .Z(n22927) );
  XNOR U23418 ( .A(n22933), .B(n22931), .Z(n23036) );
  AND U23419 ( .A(n23037), .B(n23038), .Z(n22931) );
  NANDN U23420 ( .A(n23039), .B(n23040), .Z(n23038) );
  OR U23421 ( .A(n23041), .B(n23042), .Z(n23040) );
  NAND U23422 ( .A(n23042), .B(n23041), .Z(n23037) );
  ANDN U23423 ( .B(B[119]), .A(n40), .Z(n22933) );
  XNOR U23424 ( .A(n22941), .B(n23043), .Z(n22934) );
  XNOR U23425 ( .A(n22940), .B(n22938), .Z(n23043) );
  AND U23426 ( .A(n23044), .B(n23045), .Z(n22938) );
  NANDN U23427 ( .A(n23046), .B(n23047), .Z(n23045) );
  NAND U23428 ( .A(n23048), .B(n23049), .Z(n23047) );
  ANDN U23429 ( .B(B[120]), .A(n41), .Z(n22940) );
  XOR U23430 ( .A(n22947), .B(n23050), .Z(n22941) );
  XNOR U23431 ( .A(n22945), .B(n22948), .Z(n23050) );
  NAND U23432 ( .A(A[2]), .B(B[121]), .Z(n22948) );
  NANDN U23433 ( .A(n23051), .B(n23052), .Z(n22945) );
  AND U23434 ( .A(A[0]), .B(B[122]), .Z(n23052) );
  XNOR U23435 ( .A(n22950), .B(n23053), .Z(n22947) );
  NAND U23436 ( .A(A[0]), .B(B[123]), .Z(n23053) );
  NAND U23437 ( .A(B[122]), .B(A[1]), .Z(n22950) );
  NAND U23438 ( .A(n23054), .B(n23055), .Z(n509) );
  NANDN U23439 ( .A(n23056), .B(n23057), .Z(n23055) );
  OR U23440 ( .A(n23058), .B(n23059), .Z(n23057) );
  NAND U23441 ( .A(n23059), .B(n23058), .Z(n23054) );
  XOR U23442 ( .A(n511), .B(n510), .Z(\A1[120] ) );
  XOR U23443 ( .A(n23059), .B(n23060), .Z(n510) );
  XNOR U23444 ( .A(n23058), .B(n23056), .Z(n23060) );
  AND U23445 ( .A(n23061), .B(n23062), .Z(n23056) );
  NANDN U23446 ( .A(n23063), .B(n23064), .Z(n23062) );
  NANDN U23447 ( .A(n23065), .B(n23066), .Z(n23064) );
  NANDN U23448 ( .A(n23066), .B(n23065), .Z(n23061) );
  ANDN U23449 ( .B(B[107]), .A(n29), .Z(n23058) );
  XNOR U23450 ( .A(n22965), .B(n23067), .Z(n23059) );
  XNOR U23451 ( .A(n22964), .B(n22962), .Z(n23067) );
  AND U23452 ( .A(n23068), .B(n23069), .Z(n22962) );
  NANDN U23453 ( .A(n23070), .B(n23071), .Z(n23069) );
  OR U23454 ( .A(n23072), .B(n23073), .Z(n23071) );
  NAND U23455 ( .A(n23073), .B(n23072), .Z(n23068) );
  ANDN U23456 ( .B(B[108]), .A(n30), .Z(n22964) );
  XNOR U23457 ( .A(n22972), .B(n23074), .Z(n22965) );
  XNOR U23458 ( .A(n22971), .B(n22969), .Z(n23074) );
  AND U23459 ( .A(n23075), .B(n23076), .Z(n22969) );
  NANDN U23460 ( .A(n23077), .B(n23078), .Z(n23076) );
  NANDN U23461 ( .A(n23079), .B(n23080), .Z(n23078) );
  NANDN U23462 ( .A(n23080), .B(n23079), .Z(n23075) );
  ANDN U23463 ( .B(B[109]), .A(n31), .Z(n22971) );
  XNOR U23464 ( .A(n22979), .B(n23081), .Z(n22972) );
  XNOR U23465 ( .A(n22978), .B(n22976), .Z(n23081) );
  AND U23466 ( .A(n23082), .B(n23083), .Z(n22976) );
  NANDN U23467 ( .A(n23084), .B(n23085), .Z(n23083) );
  OR U23468 ( .A(n23086), .B(n23087), .Z(n23085) );
  NAND U23469 ( .A(n23087), .B(n23086), .Z(n23082) );
  ANDN U23470 ( .B(B[110]), .A(n32), .Z(n22978) );
  XNOR U23471 ( .A(n22986), .B(n23088), .Z(n22979) );
  XNOR U23472 ( .A(n22985), .B(n22983), .Z(n23088) );
  AND U23473 ( .A(n23089), .B(n23090), .Z(n22983) );
  NANDN U23474 ( .A(n23091), .B(n23092), .Z(n23090) );
  NANDN U23475 ( .A(n23093), .B(n23094), .Z(n23092) );
  NANDN U23476 ( .A(n23094), .B(n23093), .Z(n23089) );
  ANDN U23477 ( .B(B[111]), .A(n33), .Z(n22985) );
  XNOR U23478 ( .A(n22993), .B(n23095), .Z(n22986) );
  XNOR U23479 ( .A(n22992), .B(n22990), .Z(n23095) );
  AND U23480 ( .A(n23096), .B(n23097), .Z(n22990) );
  NANDN U23481 ( .A(n23098), .B(n23099), .Z(n23097) );
  OR U23482 ( .A(n23100), .B(n23101), .Z(n23099) );
  NAND U23483 ( .A(n23101), .B(n23100), .Z(n23096) );
  ANDN U23484 ( .B(B[112]), .A(n34), .Z(n22992) );
  XNOR U23485 ( .A(n23000), .B(n23102), .Z(n22993) );
  XNOR U23486 ( .A(n22999), .B(n22997), .Z(n23102) );
  AND U23487 ( .A(n23103), .B(n23104), .Z(n22997) );
  NANDN U23488 ( .A(n23105), .B(n23106), .Z(n23104) );
  NANDN U23489 ( .A(n23107), .B(n23108), .Z(n23106) );
  NANDN U23490 ( .A(n23108), .B(n23107), .Z(n23103) );
  ANDN U23491 ( .B(B[113]), .A(n35), .Z(n22999) );
  XNOR U23492 ( .A(n23007), .B(n23109), .Z(n23000) );
  XNOR U23493 ( .A(n23006), .B(n23004), .Z(n23109) );
  AND U23494 ( .A(n23110), .B(n23111), .Z(n23004) );
  NANDN U23495 ( .A(n23112), .B(n23113), .Z(n23111) );
  OR U23496 ( .A(n23114), .B(n23115), .Z(n23113) );
  NAND U23497 ( .A(n23115), .B(n23114), .Z(n23110) );
  ANDN U23498 ( .B(B[114]), .A(n36), .Z(n23006) );
  XNOR U23499 ( .A(n23014), .B(n23116), .Z(n23007) );
  XNOR U23500 ( .A(n23013), .B(n23011), .Z(n23116) );
  AND U23501 ( .A(n23117), .B(n23118), .Z(n23011) );
  NANDN U23502 ( .A(n23119), .B(n23120), .Z(n23118) );
  NANDN U23503 ( .A(n23121), .B(n23122), .Z(n23120) );
  NANDN U23504 ( .A(n23122), .B(n23121), .Z(n23117) );
  ANDN U23505 ( .B(B[115]), .A(n37), .Z(n23013) );
  XNOR U23506 ( .A(n23021), .B(n23123), .Z(n23014) );
  XNOR U23507 ( .A(n23020), .B(n23018), .Z(n23123) );
  AND U23508 ( .A(n23124), .B(n23125), .Z(n23018) );
  NANDN U23509 ( .A(n23126), .B(n23127), .Z(n23125) );
  OR U23510 ( .A(n23128), .B(n23129), .Z(n23127) );
  NAND U23511 ( .A(n23129), .B(n23128), .Z(n23124) );
  ANDN U23512 ( .B(B[116]), .A(n38), .Z(n23020) );
  XNOR U23513 ( .A(n23028), .B(n23130), .Z(n23021) );
  XNOR U23514 ( .A(n23027), .B(n23025), .Z(n23130) );
  AND U23515 ( .A(n23131), .B(n23132), .Z(n23025) );
  NANDN U23516 ( .A(n23133), .B(n23134), .Z(n23132) );
  NANDN U23517 ( .A(n23135), .B(n23136), .Z(n23134) );
  NANDN U23518 ( .A(n23136), .B(n23135), .Z(n23131) );
  ANDN U23519 ( .B(B[117]), .A(n39), .Z(n23027) );
  XNOR U23520 ( .A(n23035), .B(n23137), .Z(n23028) );
  XNOR U23521 ( .A(n23034), .B(n23032), .Z(n23137) );
  AND U23522 ( .A(n23138), .B(n23139), .Z(n23032) );
  NANDN U23523 ( .A(n23140), .B(n23141), .Z(n23139) );
  OR U23524 ( .A(n23142), .B(n23143), .Z(n23141) );
  NAND U23525 ( .A(n23143), .B(n23142), .Z(n23138) );
  ANDN U23526 ( .B(B[118]), .A(n40), .Z(n23034) );
  XNOR U23527 ( .A(n23042), .B(n23144), .Z(n23035) );
  XNOR U23528 ( .A(n23041), .B(n23039), .Z(n23144) );
  AND U23529 ( .A(n23145), .B(n23146), .Z(n23039) );
  NANDN U23530 ( .A(n23147), .B(n23148), .Z(n23146) );
  NAND U23531 ( .A(n23149), .B(n23150), .Z(n23148) );
  ANDN U23532 ( .B(B[119]), .A(n41), .Z(n23041) );
  XOR U23533 ( .A(n23048), .B(n23151), .Z(n23042) );
  XNOR U23534 ( .A(n23046), .B(n23049), .Z(n23151) );
  NAND U23535 ( .A(A[2]), .B(B[120]), .Z(n23049) );
  NANDN U23536 ( .A(n23152), .B(n23153), .Z(n23046) );
  AND U23537 ( .A(A[0]), .B(B[121]), .Z(n23153) );
  XNOR U23538 ( .A(n23051), .B(n23154), .Z(n23048) );
  NAND U23539 ( .A(A[0]), .B(B[122]), .Z(n23154) );
  NAND U23540 ( .A(B[121]), .B(A[1]), .Z(n23051) );
  NAND U23541 ( .A(n23155), .B(n23156), .Z(n511) );
  NANDN U23542 ( .A(n23157), .B(n23158), .Z(n23156) );
  OR U23543 ( .A(n23159), .B(n23160), .Z(n23158) );
  NAND U23544 ( .A(n23160), .B(n23159), .Z(n23155) );
  XOR U23545 ( .A(n22069), .B(n23161), .Z(\A1[11] ) );
  XNOR U23546 ( .A(n22068), .B(n22066), .Z(n23161) );
  AND U23547 ( .A(n23162), .B(n23163), .Z(n22066) );
  NANDN U23548 ( .A(n23164), .B(n23165), .Z(n23163) );
  NANDN U23549 ( .A(n23166), .B(n23167), .Z(n23165) );
  NANDN U23550 ( .A(n23167), .B(n23166), .Z(n23162) );
  ANDN U23551 ( .B(B[0]), .A(n31), .Z(n22068) );
  XNOR U23552 ( .A(n22076), .B(n23168), .Z(n22069) );
  XNOR U23553 ( .A(n22075), .B(n22073), .Z(n23168) );
  AND U23554 ( .A(n23169), .B(n23170), .Z(n22073) );
  NANDN U23555 ( .A(n23171), .B(n23172), .Z(n23170) );
  OR U23556 ( .A(n23173), .B(n23174), .Z(n23172) );
  NAND U23557 ( .A(n23174), .B(n23173), .Z(n23169) );
  ANDN U23558 ( .B(B[1]), .A(n32), .Z(n22075) );
  XNOR U23559 ( .A(n22083), .B(n23175), .Z(n22076) );
  XNOR U23560 ( .A(n22082), .B(n22080), .Z(n23175) );
  AND U23561 ( .A(n23176), .B(n23177), .Z(n22080) );
  NANDN U23562 ( .A(n23178), .B(n23179), .Z(n23177) );
  NANDN U23563 ( .A(n23180), .B(n23181), .Z(n23179) );
  NANDN U23564 ( .A(n23181), .B(n23180), .Z(n23176) );
  ANDN U23565 ( .B(B[2]), .A(n33), .Z(n22082) );
  XNOR U23566 ( .A(n22090), .B(n23182), .Z(n22083) );
  XNOR U23567 ( .A(n22089), .B(n22087), .Z(n23182) );
  AND U23568 ( .A(n23183), .B(n23184), .Z(n22087) );
  NANDN U23569 ( .A(n23185), .B(n23186), .Z(n23184) );
  OR U23570 ( .A(n23187), .B(n23188), .Z(n23186) );
  NAND U23571 ( .A(n23188), .B(n23187), .Z(n23183) );
  ANDN U23572 ( .B(B[3]), .A(n34), .Z(n22089) );
  XNOR U23573 ( .A(n22097), .B(n23189), .Z(n22090) );
  XNOR U23574 ( .A(n22096), .B(n22094), .Z(n23189) );
  AND U23575 ( .A(n23190), .B(n23191), .Z(n22094) );
  NANDN U23576 ( .A(n23192), .B(n23193), .Z(n23191) );
  NANDN U23577 ( .A(n23194), .B(n23195), .Z(n23193) );
  NANDN U23578 ( .A(n23195), .B(n23194), .Z(n23190) );
  ANDN U23579 ( .B(B[4]), .A(n35), .Z(n22096) );
  XNOR U23580 ( .A(n22104), .B(n23196), .Z(n22097) );
  XNOR U23581 ( .A(n22103), .B(n22101), .Z(n23196) );
  AND U23582 ( .A(n23197), .B(n23198), .Z(n22101) );
  NANDN U23583 ( .A(n23199), .B(n23200), .Z(n23198) );
  OR U23584 ( .A(n23201), .B(n23202), .Z(n23200) );
  NAND U23585 ( .A(n23202), .B(n23201), .Z(n23197) );
  ANDN U23586 ( .B(B[5]), .A(n36), .Z(n22103) );
  XNOR U23587 ( .A(n22111), .B(n23203), .Z(n22104) );
  XNOR U23588 ( .A(n22110), .B(n22108), .Z(n23203) );
  AND U23589 ( .A(n23204), .B(n23205), .Z(n22108) );
  NANDN U23590 ( .A(n23206), .B(n23207), .Z(n23205) );
  NANDN U23591 ( .A(n23208), .B(n23209), .Z(n23207) );
  NANDN U23592 ( .A(n23209), .B(n23208), .Z(n23204) );
  ANDN U23593 ( .B(B[6]), .A(n37), .Z(n22110) );
  XNOR U23594 ( .A(n22118), .B(n23210), .Z(n22111) );
  XNOR U23595 ( .A(n22117), .B(n22115), .Z(n23210) );
  AND U23596 ( .A(n23211), .B(n23212), .Z(n22115) );
  NANDN U23597 ( .A(n23213), .B(n23214), .Z(n23212) );
  OR U23598 ( .A(n23215), .B(n23216), .Z(n23214) );
  NAND U23599 ( .A(n23216), .B(n23215), .Z(n23211) );
  ANDN U23600 ( .B(B[7]), .A(n38), .Z(n22117) );
  XNOR U23601 ( .A(n22125), .B(n23217), .Z(n22118) );
  XNOR U23602 ( .A(n22124), .B(n22122), .Z(n23217) );
  AND U23603 ( .A(n23218), .B(n23219), .Z(n22122) );
  NANDN U23604 ( .A(n23220), .B(n23221), .Z(n23219) );
  NANDN U23605 ( .A(n23222), .B(n23223), .Z(n23221) );
  NANDN U23606 ( .A(n23223), .B(n23222), .Z(n23218) );
  ANDN U23607 ( .B(B[8]), .A(n39), .Z(n22124) );
  XNOR U23608 ( .A(n22132), .B(n23224), .Z(n22125) );
  XNOR U23609 ( .A(n22131), .B(n22129), .Z(n23224) );
  AND U23610 ( .A(n23225), .B(n23226), .Z(n22129) );
  NANDN U23611 ( .A(n23227), .B(n23228), .Z(n23226) );
  OR U23612 ( .A(n23229), .B(n23230), .Z(n23228) );
  NAND U23613 ( .A(n23230), .B(n23229), .Z(n23225) );
  ANDN U23614 ( .B(B[9]), .A(n40), .Z(n22131) );
  XNOR U23615 ( .A(n22139), .B(n23231), .Z(n22132) );
  XNOR U23616 ( .A(n22138), .B(n22136), .Z(n23231) );
  AND U23617 ( .A(n23232), .B(n23233), .Z(n22136) );
  NANDN U23618 ( .A(n23234), .B(n23235), .Z(n23233) );
  NAND U23619 ( .A(n23236), .B(n23237), .Z(n23235) );
  ANDN U23620 ( .B(B[10]), .A(n41), .Z(n22138) );
  XOR U23621 ( .A(n22145), .B(n23238), .Z(n22139) );
  XNOR U23622 ( .A(n22143), .B(n22146), .Z(n23238) );
  NAND U23623 ( .A(A[2]), .B(B[11]), .Z(n22146) );
  NANDN U23624 ( .A(n23239), .B(n23240), .Z(n22143) );
  AND U23625 ( .A(A[0]), .B(B[12]), .Z(n23240) );
  XNOR U23626 ( .A(n22148), .B(n23241), .Z(n22145) );
  NAND U23627 ( .A(A[0]), .B(B[13]), .Z(n23241) );
  NAND U23628 ( .A(B[12]), .B(A[1]), .Z(n22148) );
  XOR U23629 ( .A(n513), .B(n512), .Z(\A1[119] ) );
  XOR U23630 ( .A(n23160), .B(n23242), .Z(n512) );
  XNOR U23631 ( .A(n23159), .B(n23157), .Z(n23242) );
  AND U23632 ( .A(n23243), .B(n23244), .Z(n23157) );
  NANDN U23633 ( .A(n23245), .B(n23246), .Z(n23244) );
  NANDN U23634 ( .A(n23247), .B(n23248), .Z(n23246) );
  NANDN U23635 ( .A(n23248), .B(n23247), .Z(n23243) );
  ANDN U23636 ( .B(B[106]), .A(n29), .Z(n23159) );
  XNOR U23637 ( .A(n23066), .B(n23249), .Z(n23160) );
  XNOR U23638 ( .A(n23065), .B(n23063), .Z(n23249) );
  AND U23639 ( .A(n23250), .B(n23251), .Z(n23063) );
  NANDN U23640 ( .A(n23252), .B(n23253), .Z(n23251) );
  OR U23641 ( .A(n23254), .B(n23255), .Z(n23253) );
  NAND U23642 ( .A(n23255), .B(n23254), .Z(n23250) );
  ANDN U23643 ( .B(B[107]), .A(n30), .Z(n23065) );
  XNOR U23644 ( .A(n23073), .B(n23256), .Z(n23066) );
  XNOR U23645 ( .A(n23072), .B(n23070), .Z(n23256) );
  AND U23646 ( .A(n23257), .B(n23258), .Z(n23070) );
  NANDN U23647 ( .A(n23259), .B(n23260), .Z(n23258) );
  NANDN U23648 ( .A(n23261), .B(n23262), .Z(n23260) );
  NANDN U23649 ( .A(n23262), .B(n23261), .Z(n23257) );
  ANDN U23650 ( .B(B[108]), .A(n31), .Z(n23072) );
  XNOR U23651 ( .A(n23080), .B(n23263), .Z(n23073) );
  XNOR U23652 ( .A(n23079), .B(n23077), .Z(n23263) );
  AND U23653 ( .A(n23264), .B(n23265), .Z(n23077) );
  NANDN U23654 ( .A(n23266), .B(n23267), .Z(n23265) );
  OR U23655 ( .A(n23268), .B(n23269), .Z(n23267) );
  NAND U23656 ( .A(n23269), .B(n23268), .Z(n23264) );
  ANDN U23657 ( .B(B[109]), .A(n32), .Z(n23079) );
  XNOR U23658 ( .A(n23087), .B(n23270), .Z(n23080) );
  XNOR U23659 ( .A(n23086), .B(n23084), .Z(n23270) );
  AND U23660 ( .A(n23271), .B(n23272), .Z(n23084) );
  NANDN U23661 ( .A(n23273), .B(n23274), .Z(n23272) );
  NANDN U23662 ( .A(n23275), .B(n23276), .Z(n23274) );
  NANDN U23663 ( .A(n23276), .B(n23275), .Z(n23271) );
  ANDN U23664 ( .B(B[110]), .A(n33), .Z(n23086) );
  XNOR U23665 ( .A(n23094), .B(n23277), .Z(n23087) );
  XNOR U23666 ( .A(n23093), .B(n23091), .Z(n23277) );
  AND U23667 ( .A(n23278), .B(n23279), .Z(n23091) );
  NANDN U23668 ( .A(n23280), .B(n23281), .Z(n23279) );
  OR U23669 ( .A(n23282), .B(n23283), .Z(n23281) );
  NAND U23670 ( .A(n23283), .B(n23282), .Z(n23278) );
  ANDN U23671 ( .B(B[111]), .A(n34), .Z(n23093) );
  XNOR U23672 ( .A(n23101), .B(n23284), .Z(n23094) );
  XNOR U23673 ( .A(n23100), .B(n23098), .Z(n23284) );
  AND U23674 ( .A(n23285), .B(n23286), .Z(n23098) );
  NANDN U23675 ( .A(n23287), .B(n23288), .Z(n23286) );
  NANDN U23676 ( .A(n23289), .B(n23290), .Z(n23288) );
  NANDN U23677 ( .A(n23290), .B(n23289), .Z(n23285) );
  ANDN U23678 ( .B(B[112]), .A(n35), .Z(n23100) );
  XNOR U23679 ( .A(n23108), .B(n23291), .Z(n23101) );
  XNOR U23680 ( .A(n23107), .B(n23105), .Z(n23291) );
  AND U23681 ( .A(n23292), .B(n23293), .Z(n23105) );
  NANDN U23682 ( .A(n23294), .B(n23295), .Z(n23293) );
  OR U23683 ( .A(n23296), .B(n23297), .Z(n23295) );
  NAND U23684 ( .A(n23297), .B(n23296), .Z(n23292) );
  ANDN U23685 ( .B(B[113]), .A(n36), .Z(n23107) );
  XNOR U23686 ( .A(n23115), .B(n23298), .Z(n23108) );
  XNOR U23687 ( .A(n23114), .B(n23112), .Z(n23298) );
  AND U23688 ( .A(n23299), .B(n23300), .Z(n23112) );
  NANDN U23689 ( .A(n23301), .B(n23302), .Z(n23300) );
  NANDN U23690 ( .A(n23303), .B(n23304), .Z(n23302) );
  NANDN U23691 ( .A(n23304), .B(n23303), .Z(n23299) );
  ANDN U23692 ( .B(B[114]), .A(n37), .Z(n23114) );
  XNOR U23693 ( .A(n23122), .B(n23305), .Z(n23115) );
  XNOR U23694 ( .A(n23121), .B(n23119), .Z(n23305) );
  AND U23695 ( .A(n23306), .B(n23307), .Z(n23119) );
  NANDN U23696 ( .A(n23308), .B(n23309), .Z(n23307) );
  OR U23697 ( .A(n23310), .B(n23311), .Z(n23309) );
  NAND U23698 ( .A(n23311), .B(n23310), .Z(n23306) );
  ANDN U23699 ( .B(B[115]), .A(n38), .Z(n23121) );
  XNOR U23700 ( .A(n23129), .B(n23312), .Z(n23122) );
  XNOR U23701 ( .A(n23128), .B(n23126), .Z(n23312) );
  AND U23702 ( .A(n23313), .B(n23314), .Z(n23126) );
  NANDN U23703 ( .A(n23315), .B(n23316), .Z(n23314) );
  NANDN U23704 ( .A(n23317), .B(n23318), .Z(n23316) );
  NANDN U23705 ( .A(n23318), .B(n23317), .Z(n23313) );
  ANDN U23706 ( .B(B[116]), .A(n39), .Z(n23128) );
  XNOR U23707 ( .A(n23136), .B(n23319), .Z(n23129) );
  XNOR U23708 ( .A(n23135), .B(n23133), .Z(n23319) );
  AND U23709 ( .A(n23320), .B(n23321), .Z(n23133) );
  NANDN U23710 ( .A(n23322), .B(n23323), .Z(n23321) );
  OR U23711 ( .A(n23324), .B(n23325), .Z(n23323) );
  NAND U23712 ( .A(n23325), .B(n23324), .Z(n23320) );
  ANDN U23713 ( .B(B[117]), .A(n40), .Z(n23135) );
  XNOR U23714 ( .A(n23143), .B(n23326), .Z(n23136) );
  XNOR U23715 ( .A(n23142), .B(n23140), .Z(n23326) );
  AND U23716 ( .A(n23327), .B(n23328), .Z(n23140) );
  NANDN U23717 ( .A(n23329), .B(n23330), .Z(n23328) );
  NAND U23718 ( .A(n23331), .B(n23332), .Z(n23330) );
  ANDN U23719 ( .B(B[118]), .A(n41), .Z(n23142) );
  XOR U23720 ( .A(n23149), .B(n23333), .Z(n23143) );
  XNOR U23721 ( .A(n23147), .B(n23150), .Z(n23333) );
  NAND U23722 ( .A(A[2]), .B(B[119]), .Z(n23150) );
  NANDN U23723 ( .A(n23334), .B(n23335), .Z(n23147) );
  AND U23724 ( .A(A[0]), .B(B[120]), .Z(n23335) );
  XNOR U23725 ( .A(n23152), .B(n23336), .Z(n23149) );
  NAND U23726 ( .A(A[0]), .B(B[121]), .Z(n23336) );
  NAND U23727 ( .A(B[120]), .B(A[1]), .Z(n23152) );
  NAND U23728 ( .A(n23337), .B(n23338), .Z(n513) );
  NANDN U23729 ( .A(n23339), .B(n23340), .Z(n23338) );
  OR U23730 ( .A(n23341), .B(n23342), .Z(n23340) );
  NAND U23731 ( .A(n23342), .B(n23341), .Z(n23337) );
  XOR U23732 ( .A(n515), .B(n514), .Z(\A1[118] ) );
  XOR U23733 ( .A(n23342), .B(n23343), .Z(n514) );
  XNOR U23734 ( .A(n23341), .B(n23339), .Z(n23343) );
  AND U23735 ( .A(n23344), .B(n23345), .Z(n23339) );
  NANDN U23736 ( .A(n23346), .B(n23347), .Z(n23345) );
  NANDN U23737 ( .A(n23348), .B(n23349), .Z(n23347) );
  NANDN U23738 ( .A(n23349), .B(n23348), .Z(n23344) );
  ANDN U23739 ( .B(B[105]), .A(n29), .Z(n23341) );
  XNOR U23740 ( .A(n23248), .B(n23350), .Z(n23342) );
  XNOR U23741 ( .A(n23247), .B(n23245), .Z(n23350) );
  AND U23742 ( .A(n23351), .B(n23352), .Z(n23245) );
  NANDN U23743 ( .A(n23353), .B(n23354), .Z(n23352) );
  OR U23744 ( .A(n23355), .B(n23356), .Z(n23354) );
  NAND U23745 ( .A(n23356), .B(n23355), .Z(n23351) );
  ANDN U23746 ( .B(B[106]), .A(n30), .Z(n23247) );
  XNOR U23747 ( .A(n23255), .B(n23357), .Z(n23248) );
  XNOR U23748 ( .A(n23254), .B(n23252), .Z(n23357) );
  AND U23749 ( .A(n23358), .B(n23359), .Z(n23252) );
  NANDN U23750 ( .A(n23360), .B(n23361), .Z(n23359) );
  NANDN U23751 ( .A(n23362), .B(n23363), .Z(n23361) );
  NANDN U23752 ( .A(n23363), .B(n23362), .Z(n23358) );
  ANDN U23753 ( .B(B[107]), .A(n31), .Z(n23254) );
  XNOR U23754 ( .A(n23262), .B(n23364), .Z(n23255) );
  XNOR U23755 ( .A(n23261), .B(n23259), .Z(n23364) );
  AND U23756 ( .A(n23365), .B(n23366), .Z(n23259) );
  NANDN U23757 ( .A(n23367), .B(n23368), .Z(n23366) );
  OR U23758 ( .A(n23369), .B(n23370), .Z(n23368) );
  NAND U23759 ( .A(n23370), .B(n23369), .Z(n23365) );
  ANDN U23760 ( .B(B[108]), .A(n32), .Z(n23261) );
  XNOR U23761 ( .A(n23269), .B(n23371), .Z(n23262) );
  XNOR U23762 ( .A(n23268), .B(n23266), .Z(n23371) );
  AND U23763 ( .A(n23372), .B(n23373), .Z(n23266) );
  NANDN U23764 ( .A(n23374), .B(n23375), .Z(n23373) );
  NANDN U23765 ( .A(n23376), .B(n23377), .Z(n23375) );
  NANDN U23766 ( .A(n23377), .B(n23376), .Z(n23372) );
  ANDN U23767 ( .B(B[109]), .A(n33), .Z(n23268) );
  XNOR U23768 ( .A(n23276), .B(n23378), .Z(n23269) );
  XNOR U23769 ( .A(n23275), .B(n23273), .Z(n23378) );
  AND U23770 ( .A(n23379), .B(n23380), .Z(n23273) );
  NANDN U23771 ( .A(n23381), .B(n23382), .Z(n23380) );
  OR U23772 ( .A(n23383), .B(n23384), .Z(n23382) );
  NAND U23773 ( .A(n23384), .B(n23383), .Z(n23379) );
  ANDN U23774 ( .B(B[110]), .A(n34), .Z(n23275) );
  XNOR U23775 ( .A(n23283), .B(n23385), .Z(n23276) );
  XNOR U23776 ( .A(n23282), .B(n23280), .Z(n23385) );
  AND U23777 ( .A(n23386), .B(n23387), .Z(n23280) );
  NANDN U23778 ( .A(n23388), .B(n23389), .Z(n23387) );
  NANDN U23779 ( .A(n23390), .B(n23391), .Z(n23389) );
  NANDN U23780 ( .A(n23391), .B(n23390), .Z(n23386) );
  ANDN U23781 ( .B(B[111]), .A(n35), .Z(n23282) );
  XNOR U23782 ( .A(n23290), .B(n23392), .Z(n23283) );
  XNOR U23783 ( .A(n23289), .B(n23287), .Z(n23392) );
  AND U23784 ( .A(n23393), .B(n23394), .Z(n23287) );
  NANDN U23785 ( .A(n23395), .B(n23396), .Z(n23394) );
  OR U23786 ( .A(n23397), .B(n23398), .Z(n23396) );
  NAND U23787 ( .A(n23398), .B(n23397), .Z(n23393) );
  ANDN U23788 ( .B(B[112]), .A(n36), .Z(n23289) );
  XNOR U23789 ( .A(n23297), .B(n23399), .Z(n23290) );
  XNOR U23790 ( .A(n23296), .B(n23294), .Z(n23399) );
  AND U23791 ( .A(n23400), .B(n23401), .Z(n23294) );
  NANDN U23792 ( .A(n23402), .B(n23403), .Z(n23401) );
  NANDN U23793 ( .A(n23404), .B(n23405), .Z(n23403) );
  NANDN U23794 ( .A(n23405), .B(n23404), .Z(n23400) );
  ANDN U23795 ( .B(B[113]), .A(n37), .Z(n23296) );
  XNOR U23796 ( .A(n23304), .B(n23406), .Z(n23297) );
  XNOR U23797 ( .A(n23303), .B(n23301), .Z(n23406) );
  AND U23798 ( .A(n23407), .B(n23408), .Z(n23301) );
  NANDN U23799 ( .A(n23409), .B(n23410), .Z(n23408) );
  OR U23800 ( .A(n23411), .B(n23412), .Z(n23410) );
  NAND U23801 ( .A(n23412), .B(n23411), .Z(n23407) );
  ANDN U23802 ( .B(B[114]), .A(n38), .Z(n23303) );
  XNOR U23803 ( .A(n23311), .B(n23413), .Z(n23304) );
  XNOR U23804 ( .A(n23310), .B(n23308), .Z(n23413) );
  AND U23805 ( .A(n23414), .B(n23415), .Z(n23308) );
  NANDN U23806 ( .A(n23416), .B(n23417), .Z(n23415) );
  NANDN U23807 ( .A(n23418), .B(n23419), .Z(n23417) );
  NANDN U23808 ( .A(n23419), .B(n23418), .Z(n23414) );
  ANDN U23809 ( .B(B[115]), .A(n39), .Z(n23310) );
  XNOR U23810 ( .A(n23318), .B(n23420), .Z(n23311) );
  XNOR U23811 ( .A(n23317), .B(n23315), .Z(n23420) );
  AND U23812 ( .A(n23421), .B(n23422), .Z(n23315) );
  NANDN U23813 ( .A(n23423), .B(n23424), .Z(n23422) );
  OR U23814 ( .A(n23425), .B(n23426), .Z(n23424) );
  NAND U23815 ( .A(n23426), .B(n23425), .Z(n23421) );
  ANDN U23816 ( .B(B[116]), .A(n40), .Z(n23317) );
  XNOR U23817 ( .A(n23325), .B(n23427), .Z(n23318) );
  XNOR U23818 ( .A(n23324), .B(n23322), .Z(n23427) );
  AND U23819 ( .A(n23428), .B(n23429), .Z(n23322) );
  NANDN U23820 ( .A(n23430), .B(n23431), .Z(n23429) );
  NAND U23821 ( .A(n23432), .B(n23433), .Z(n23431) );
  ANDN U23822 ( .B(B[117]), .A(n41), .Z(n23324) );
  XOR U23823 ( .A(n23331), .B(n23434), .Z(n23325) );
  XNOR U23824 ( .A(n23329), .B(n23332), .Z(n23434) );
  NAND U23825 ( .A(A[2]), .B(B[118]), .Z(n23332) );
  NANDN U23826 ( .A(n23435), .B(n23436), .Z(n23329) );
  AND U23827 ( .A(A[0]), .B(B[119]), .Z(n23436) );
  XNOR U23828 ( .A(n23334), .B(n23437), .Z(n23331) );
  NAND U23829 ( .A(A[0]), .B(B[120]), .Z(n23437) );
  NAND U23830 ( .A(B[119]), .B(A[1]), .Z(n23334) );
  NAND U23831 ( .A(n23438), .B(n23439), .Z(n515) );
  NANDN U23832 ( .A(n23440), .B(n23441), .Z(n23439) );
  OR U23833 ( .A(n23442), .B(n23443), .Z(n23441) );
  NAND U23834 ( .A(n23443), .B(n23442), .Z(n23438) );
  XOR U23835 ( .A(n517), .B(n516), .Z(\A1[117] ) );
  XOR U23836 ( .A(n23443), .B(n23444), .Z(n516) );
  XNOR U23837 ( .A(n23442), .B(n23440), .Z(n23444) );
  AND U23838 ( .A(n23445), .B(n23446), .Z(n23440) );
  NANDN U23839 ( .A(n23447), .B(n23448), .Z(n23446) );
  NANDN U23840 ( .A(n23449), .B(n23450), .Z(n23448) );
  NANDN U23841 ( .A(n23450), .B(n23449), .Z(n23445) );
  ANDN U23842 ( .B(B[104]), .A(n29), .Z(n23442) );
  XNOR U23843 ( .A(n23349), .B(n23451), .Z(n23443) );
  XNOR U23844 ( .A(n23348), .B(n23346), .Z(n23451) );
  AND U23845 ( .A(n23452), .B(n23453), .Z(n23346) );
  NANDN U23846 ( .A(n23454), .B(n23455), .Z(n23453) );
  OR U23847 ( .A(n23456), .B(n23457), .Z(n23455) );
  NAND U23848 ( .A(n23457), .B(n23456), .Z(n23452) );
  ANDN U23849 ( .B(B[105]), .A(n30), .Z(n23348) );
  XNOR U23850 ( .A(n23356), .B(n23458), .Z(n23349) );
  XNOR U23851 ( .A(n23355), .B(n23353), .Z(n23458) );
  AND U23852 ( .A(n23459), .B(n23460), .Z(n23353) );
  NANDN U23853 ( .A(n23461), .B(n23462), .Z(n23460) );
  NANDN U23854 ( .A(n23463), .B(n23464), .Z(n23462) );
  NANDN U23855 ( .A(n23464), .B(n23463), .Z(n23459) );
  ANDN U23856 ( .B(B[106]), .A(n31), .Z(n23355) );
  XNOR U23857 ( .A(n23363), .B(n23465), .Z(n23356) );
  XNOR U23858 ( .A(n23362), .B(n23360), .Z(n23465) );
  AND U23859 ( .A(n23466), .B(n23467), .Z(n23360) );
  NANDN U23860 ( .A(n23468), .B(n23469), .Z(n23467) );
  OR U23861 ( .A(n23470), .B(n23471), .Z(n23469) );
  NAND U23862 ( .A(n23471), .B(n23470), .Z(n23466) );
  ANDN U23863 ( .B(B[107]), .A(n32), .Z(n23362) );
  XNOR U23864 ( .A(n23370), .B(n23472), .Z(n23363) );
  XNOR U23865 ( .A(n23369), .B(n23367), .Z(n23472) );
  AND U23866 ( .A(n23473), .B(n23474), .Z(n23367) );
  NANDN U23867 ( .A(n23475), .B(n23476), .Z(n23474) );
  NANDN U23868 ( .A(n23477), .B(n23478), .Z(n23476) );
  NANDN U23869 ( .A(n23478), .B(n23477), .Z(n23473) );
  ANDN U23870 ( .B(B[108]), .A(n33), .Z(n23369) );
  XNOR U23871 ( .A(n23377), .B(n23479), .Z(n23370) );
  XNOR U23872 ( .A(n23376), .B(n23374), .Z(n23479) );
  AND U23873 ( .A(n23480), .B(n23481), .Z(n23374) );
  NANDN U23874 ( .A(n23482), .B(n23483), .Z(n23481) );
  OR U23875 ( .A(n23484), .B(n23485), .Z(n23483) );
  NAND U23876 ( .A(n23485), .B(n23484), .Z(n23480) );
  ANDN U23877 ( .B(B[109]), .A(n34), .Z(n23376) );
  XNOR U23878 ( .A(n23384), .B(n23486), .Z(n23377) );
  XNOR U23879 ( .A(n23383), .B(n23381), .Z(n23486) );
  AND U23880 ( .A(n23487), .B(n23488), .Z(n23381) );
  NANDN U23881 ( .A(n23489), .B(n23490), .Z(n23488) );
  NANDN U23882 ( .A(n23491), .B(n23492), .Z(n23490) );
  NANDN U23883 ( .A(n23492), .B(n23491), .Z(n23487) );
  ANDN U23884 ( .B(B[110]), .A(n35), .Z(n23383) );
  XNOR U23885 ( .A(n23391), .B(n23493), .Z(n23384) );
  XNOR U23886 ( .A(n23390), .B(n23388), .Z(n23493) );
  AND U23887 ( .A(n23494), .B(n23495), .Z(n23388) );
  NANDN U23888 ( .A(n23496), .B(n23497), .Z(n23495) );
  OR U23889 ( .A(n23498), .B(n23499), .Z(n23497) );
  NAND U23890 ( .A(n23499), .B(n23498), .Z(n23494) );
  ANDN U23891 ( .B(B[111]), .A(n36), .Z(n23390) );
  XNOR U23892 ( .A(n23398), .B(n23500), .Z(n23391) );
  XNOR U23893 ( .A(n23397), .B(n23395), .Z(n23500) );
  AND U23894 ( .A(n23501), .B(n23502), .Z(n23395) );
  NANDN U23895 ( .A(n23503), .B(n23504), .Z(n23502) );
  NANDN U23896 ( .A(n23505), .B(n23506), .Z(n23504) );
  NANDN U23897 ( .A(n23506), .B(n23505), .Z(n23501) );
  ANDN U23898 ( .B(B[112]), .A(n37), .Z(n23397) );
  XNOR U23899 ( .A(n23405), .B(n23507), .Z(n23398) );
  XNOR U23900 ( .A(n23404), .B(n23402), .Z(n23507) );
  AND U23901 ( .A(n23508), .B(n23509), .Z(n23402) );
  NANDN U23902 ( .A(n23510), .B(n23511), .Z(n23509) );
  OR U23903 ( .A(n23512), .B(n23513), .Z(n23511) );
  NAND U23904 ( .A(n23513), .B(n23512), .Z(n23508) );
  ANDN U23905 ( .B(B[113]), .A(n38), .Z(n23404) );
  XNOR U23906 ( .A(n23412), .B(n23514), .Z(n23405) );
  XNOR U23907 ( .A(n23411), .B(n23409), .Z(n23514) );
  AND U23908 ( .A(n23515), .B(n23516), .Z(n23409) );
  NANDN U23909 ( .A(n23517), .B(n23518), .Z(n23516) );
  NANDN U23910 ( .A(n23519), .B(n23520), .Z(n23518) );
  NANDN U23911 ( .A(n23520), .B(n23519), .Z(n23515) );
  ANDN U23912 ( .B(B[114]), .A(n39), .Z(n23411) );
  XNOR U23913 ( .A(n23419), .B(n23521), .Z(n23412) );
  XNOR U23914 ( .A(n23418), .B(n23416), .Z(n23521) );
  AND U23915 ( .A(n23522), .B(n23523), .Z(n23416) );
  NANDN U23916 ( .A(n23524), .B(n23525), .Z(n23523) );
  OR U23917 ( .A(n23526), .B(n23527), .Z(n23525) );
  NAND U23918 ( .A(n23527), .B(n23526), .Z(n23522) );
  ANDN U23919 ( .B(B[115]), .A(n40), .Z(n23418) );
  XNOR U23920 ( .A(n23426), .B(n23528), .Z(n23419) );
  XNOR U23921 ( .A(n23425), .B(n23423), .Z(n23528) );
  AND U23922 ( .A(n23529), .B(n23530), .Z(n23423) );
  NANDN U23923 ( .A(n23531), .B(n23532), .Z(n23530) );
  NAND U23924 ( .A(n23533), .B(n23534), .Z(n23532) );
  ANDN U23925 ( .B(B[116]), .A(n41), .Z(n23425) );
  XOR U23926 ( .A(n23432), .B(n23535), .Z(n23426) );
  XNOR U23927 ( .A(n23430), .B(n23433), .Z(n23535) );
  NAND U23928 ( .A(A[2]), .B(B[117]), .Z(n23433) );
  NANDN U23929 ( .A(n23536), .B(n23537), .Z(n23430) );
  AND U23930 ( .A(A[0]), .B(B[118]), .Z(n23537) );
  XNOR U23931 ( .A(n23435), .B(n23538), .Z(n23432) );
  NAND U23932 ( .A(A[0]), .B(B[119]), .Z(n23538) );
  NAND U23933 ( .A(B[118]), .B(A[1]), .Z(n23435) );
  NAND U23934 ( .A(n23539), .B(n23540), .Z(n517) );
  NANDN U23935 ( .A(n23541), .B(n23542), .Z(n23540) );
  OR U23936 ( .A(n23543), .B(n23544), .Z(n23542) );
  NAND U23937 ( .A(n23544), .B(n23543), .Z(n23539) );
  XOR U23938 ( .A(n519), .B(n518), .Z(\A1[116] ) );
  XOR U23939 ( .A(n23544), .B(n23545), .Z(n518) );
  XNOR U23940 ( .A(n23543), .B(n23541), .Z(n23545) );
  AND U23941 ( .A(n23546), .B(n23547), .Z(n23541) );
  NANDN U23942 ( .A(n23548), .B(n23549), .Z(n23547) );
  NANDN U23943 ( .A(n23550), .B(n23551), .Z(n23549) );
  NANDN U23944 ( .A(n23551), .B(n23550), .Z(n23546) );
  ANDN U23945 ( .B(B[103]), .A(n29), .Z(n23543) );
  XNOR U23946 ( .A(n23450), .B(n23552), .Z(n23544) );
  XNOR U23947 ( .A(n23449), .B(n23447), .Z(n23552) );
  AND U23948 ( .A(n23553), .B(n23554), .Z(n23447) );
  NANDN U23949 ( .A(n23555), .B(n23556), .Z(n23554) );
  OR U23950 ( .A(n23557), .B(n23558), .Z(n23556) );
  NAND U23951 ( .A(n23558), .B(n23557), .Z(n23553) );
  ANDN U23952 ( .B(B[104]), .A(n30), .Z(n23449) );
  XNOR U23953 ( .A(n23457), .B(n23559), .Z(n23450) );
  XNOR U23954 ( .A(n23456), .B(n23454), .Z(n23559) );
  AND U23955 ( .A(n23560), .B(n23561), .Z(n23454) );
  NANDN U23956 ( .A(n23562), .B(n23563), .Z(n23561) );
  NANDN U23957 ( .A(n23564), .B(n23565), .Z(n23563) );
  NANDN U23958 ( .A(n23565), .B(n23564), .Z(n23560) );
  ANDN U23959 ( .B(B[105]), .A(n31), .Z(n23456) );
  XNOR U23960 ( .A(n23464), .B(n23566), .Z(n23457) );
  XNOR U23961 ( .A(n23463), .B(n23461), .Z(n23566) );
  AND U23962 ( .A(n23567), .B(n23568), .Z(n23461) );
  NANDN U23963 ( .A(n23569), .B(n23570), .Z(n23568) );
  OR U23964 ( .A(n23571), .B(n23572), .Z(n23570) );
  NAND U23965 ( .A(n23572), .B(n23571), .Z(n23567) );
  ANDN U23966 ( .B(B[106]), .A(n32), .Z(n23463) );
  XNOR U23967 ( .A(n23471), .B(n23573), .Z(n23464) );
  XNOR U23968 ( .A(n23470), .B(n23468), .Z(n23573) );
  AND U23969 ( .A(n23574), .B(n23575), .Z(n23468) );
  NANDN U23970 ( .A(n23576), .B(n23577), .Z(n23575) );
  NANDN U23971 ( .A(n23578), .B(n23579), .Z(n23577) );
  NANDN U23972 ( .A(n23579), .B(n23578), .Z(n23574) );
  ANDN U23973 ( .B(B[107]), .A(n33), .Z(n23470) );
  XNOR U23974 ( .A(n23478), .B(n23580), .Z(n23471) );
  XNOR U23975 ( .A(n23477), .B(n23475), .Z(n23580) );
  AND U23976 ( .A(n23581), .B(n23582), .Z(n23475) );
  NANDN U23977 ( .A(n23583), .B(n23584), .Z(n23582) );
  OR U23978 ( .A(n23585), .B(n23586), .Z(n23584) );
  NAND U23979 ( .A(n23586), .B(n23585), .Z(n23581) );
  ANDN U23980 ( .B(B[108]), .A(n34), .Z(n23477) );
  XNOR U23981 ( .A(n23485), .B(n23587), .Z(n23478) );
  XNOR U23982 ( .A(n23484), .B(n23482), .Z(n23587) );
  AND U23983 ( .A(n23588), .B(n23589), .Z(n23482) );
  NANDN U23984 ( .A(n23590), .B(n23591), .Z(n23589) );
  NANDN U23985 ( .A(n23592), .B(n23593), .Z(n23591) );
  NANDN U23986 ( .A(n23593), .B(n23592), .Z(n23588) );
  ANDN U23987 ( .B(B[109]), .A(n35), .Z(n23484) );
  XNOR U23988 ( .A(n23492), .B(n23594), .Z(n23485) );
  XNOR U23989 ( .A(n23491), .B(n23489), .Z(n23594) );
  AND U23990 ( .A(n23595), .B(n23596), .Z(n23489) );
  NANDN U23991 ( .A(n23597), .B(n23598), .Z(n23596) );
  OR U23992 ( .A(n23599), .B(n23600), .Z(n23598) );
  NAND U23993 ( .A(n23600), .B(n23599), .Z(n23595) );
  ANDN U23994 ( .B(B[110]), .A(n36), .Z(n23491) );
  XNOR U23995 ( .A(n23499), .B(n23601), .Z(n23492) );
  XNOR U23996 ( .A(n23498), .B(n23496), .Z(n23601) );
  AND U23997 ( .A(n23602), .B(n23603), .Z(n23496) );
  NANDN U23998 ( .A(n23604), .B(n23605), .Z(n23603) );
  NANDN U23999 ( .A(n23606), .B(n23607), .Z(n23605) );
  NANDN U24000 ( .A(n23607), .B(n23606), .Z(n23602) );
  ANDN U24001 ( .B(B[111]), .A(n37), .Z(n23498) );
  XNOR U24002 ( .A(n23506), .B(n23608), .Z(n23499) );
  XNOR U24003 ( .A(n23505), .B(n23503), .Z(n23608) );
  AND U24004 ( .A(n23609), .B(n23610), .Z(n23503) );
  NANDN U24005 ( .A(n23611), .B(n23612), .Z(n23610) );
  OR U24006 ( .A(n23613), .B(n23614), .Z(n23612) );
  NAND U24007 ( .A(n23614), .B(n23613), .Z(n23609) );
  ANDN U24008 ( .B(B[112]), .A(n38), .Z(n23505) );
  XNOR U24009 ( .A(n23513), .B(n23615), .Z(n23506) );
  XNOR U24010 ( .A(n23512), .B(n23510), .Z(n23615) );
  AND U24011 ( .A(n23616), .B(n23617), .Z(n23510) );
  NANDN U24012 ( .A(n23618), .B(n23619), .Z(n23617) );
  NANDN U24013 ( .A(n23620), .B(n23621), .Z(n23619) );
  NANDN U24014 ( .A(n23621), .B(n23620), .Z(n23616) );
  ANDN U24015 ( .B(B[113]), .A(n39), .Z(n23512) );
  XNOR U24016 ( .A(n23520), .B(n23622), .Z(n23513) );
  XNOR U24017 ( .A(n23519), .B(n23517), .Z(n23622) );
  AND U24018 ( .A(n23623), .B(n23624), .Z(n23517) );
  NANDN U24019 ( .A(n23625), .B(n23626), .Z(n23624) );
  OR U24020 ( .A(n23627), .B(n23628), .Z(n23626) );
  NAND U24021 ( .A(n23628), .B(n23627), .Z(n23623) );
  ANDN U24022 ( .B(B[114]), .A(n40), .Z(n23519) );
  XNOR U24023 ( .A(n23527), .B(n23629), .Z(n23520) );
  XNOR U24024 ( .A(n23526), .B(n23524), .Z(n23629) );
  AND U24025 ( .A(n23630), .B(n23631), .Z(n23524) );
  NANDN U24026 ( .A(n23632), .B(n23633), .Z(n23631) );
  NAND U24027 ( .A(n23634), .B(n23635), .Z(n23633) );
  ANDN U24028 ( .B(B[115]), .A(n41), .Z(n23526) );
  XOR U24029 ( .A(n23533), .B(n23636), .Z(n23527) );
  XNOR U24030 ( .A(n23531), .B(n23534), .Z(n23636) );
  NAND U24031 ( .A(A[2]), .B(B[116]), .Z(n23534) );
  NANDN U24032 ( .A(n23637), .B(n23638), .Z(n23531) );
  AND U24033 ( .A(A[0]), .B(B[117]), .Z(n23638) );
  XNOR U24034 ( .A(n23536), .B(n23639), .Z(n23533) );
  NAND U24035 ( .A(A[0]), .B(B[118]), .Z(n23639) );
  NAND U24036 ( .A(B[117]), .B(A[1]), .Z(n23536) );
  NAND U24037 ( .A(n23640), .B(n23641), .Z(n519) );
  NANDN U24038 ( .A(n23642), .B(n23643), .Z(n23641) );
  OR U24039 ( .A(n23644), .B(n23645), .Z(n23643) );
  NAND U24040 ( .A(n23645), .B(n23644), .Z(n23640) );
  XOR U24041 ( .A(n521), .B(n520), .Z(\A1[115] ) );
  XOR U24042 ( .A(n23645), .B(n23646), .Z(n520) );
  XNOR U24043 ( .A(n23644), .B(n23642), .Z(n23646) );
  AND U24044 ( .A(n23647), .B(n23648), .Z(n23642) );
  NANDN U24045 ( .A(n23649), .B(n23650), .Z(n23648) );
  NANDN U24046 ( .A(n23651), .B(n23652), .Z(n23650) );
  NANDN U24047 ( .A(n23652), .B(n23651), .Z(n23647) );
  ANDN U24048 ( .B(B[102]), .A(n29), .Z(n23644) );
  XNOR U24049 ( .A(n23551), .B(n23653), .Z(n23645) );
  XNOR U24050 ( .A(n23550), .B(n23548), .Z(n23653) );
  AND U24051 ( .A(n23654), .B(n23655), .Z(n23548) );
  NANDN U24052 ( .A(n23656), .B(n23657), .Z(n23655) );
  OR U24053 ( .A(n23658), .B(n23659), .Z(n23657) );
  NAND U24054 ( .A(n23659), .B(n23658), .Z(n23654) );
  ANDN U24055 ( .B(B[103]), .A(n30), .Z(n23550) );
  XNOR U24056 ( .A(n23558), .B(n23660), .Z(n23551) );
  XNOR U24057 ( .A(n23557), .B(n23555), .Z(n23660) );
  AND U24058 ( .A(n23661), .B(n23662), .Z(n23555) );
  NANDN U24059 ( .A(n23663), .B(n23664), .Z(n23662) );
  NANDN U24060 ( .A(n23665), .B(n23666), .Z(n23664) );
  NANDN U24061 ( .A(n23666), .B(n23665), .Z(n23661) );
  ANDN U24062 ( .B(B[104]), .A(n31), .Z(n23557) );
  XNOR U24063 ( .A(n23565), .B(n23667), .Z(n23558) );
  XNOR U24064 ( .A(n23564), .B(n23562), .Z(n23667) );
  AND U24065 ( .A(n23668), .B(n23669), .Z(n23562) );
  NANDN U24066 ( .A(n23670), .B(n23671), .Z(n23669) );
  OR U24067 ( .A(n23672), .B(n23673), .Z(n23671) );
  NAND U24068 ( .A(n23673), .B(n23672), .Z(n23668) );
  ANDN U24069 ( .B(B[105]), .A(n32), .Z(n23564) );
  XNOR U24070 ( .A(n23572), .B(n23674), .Z(n23565) );
  XNOR U24071 ( .A(n23571), .B(n23569), .Z(n23674) );
  AND U24072 ( .A(n23675), .B(n23676), .Z(n23569) );
  NANDN U24073 ( .A(n23677), .B(n23678), .Z(n23676) );
  NANDN U24074 ( .A(n23679), .B(n23680), .Z(n23678) );
  NANDN U24075 ( .A(n23680), .B(n23679), .Z(n23675) );
  ANDN U24076 ( .B(B[106]), .A(n33), .Z(n23571) );
  XNOR U24077 ( .A(n23579), .B(n23681), .Z(n23572) );
  XNOR U24078 ( .A(n23578), .B(n23576), .Z(n23681) );
  AND U24079 ( .A(n23682), .B(n23683), .Z(n23576) );
  NANDN U24080 ( .A(n23684), .B(n23685), .Z(n23683) );
  OR U24081 ( .A(n23686), .B(n23687), .Z(n23685) );
  NAND U24082 ( .A(n23687), .B(n23686), .Z(n23682) );
  ANDN U24083 ( .B(B[107]), .A(n34), .Z(n23578) );
  XNOR U24084 ( .A(n23586), .B(n23688), .Z(n23579) );
  XNOR U24085 ( .A(n23585), .B(n23583), .Z(n23688) );
  AND U24086 ( .A(n23689), .B(n23690), .Z(n23583) );
  NANDN U24087 ( .A(n23691), .B(n23692), .Z(n23690) );
  NANDN U24088 ( .A(n23693), .B(n23694), .Z(n23692) );
  NANDN U24089 ( .A(n23694), .B(n23693), .Z(n23689) );
  ANDN U24090 ( .B(B[108]), .A(n35), .Z(n23585) );
  XNOR U24091 ( .A(n23593), .B(n23695), .Z(n23586) );
  XNOR U24092 ( .A(n23592), .B(n23590), .Z(n23695) );
  AND U24093 ( .A(n23696), .B(n23697), .Z(n23590) );
  NANDN U24094 ( .A(n23698), .B(n23699), .Z(n23697) );
  OR U24095 ( .A(n23700), .B(n23701), .Z(n23699) );
  NAND U24096 ( .A(n23701), .B(n23700), .Z(n23696) );
  ANDN U24097 ( .B(B[109]), .A(n36), .Z(n23592) );
  XNOR U24098 ( .A(n23600), .B(n23702), .Z(n23593) );
  XNOR U24099 ( .A(n23599), .B(n23597), .Z(n23702) );
  AND U24100 ( .A(n23703), .B(n23704), .Z(n23597) );
  NANDN U24101 ( .A(n23705), .B(n23706), .Z(n23704) );
  NANDN U24102 ( .A(n23707), .B(n23708), .Z(n23706) );
  NANDN U24103 ( .A(n23708), .B(n23707), .Z(n23703) );
  ANDN U24104 ( .B(B[110]), .A(n37), .Z(n23599) );
  XNOR U24105 ( .A(n23607), .B(n23709), .Z(n23600) );
  XNOR U24106 ( .A(n23606), .B(n23604), .Z(n23709) );
  AND U24107 ( .A(n23710), .B(n23711), .Z(n23604) );
  NANDN U24108 ( .A(n23712), .B(n23713), .Z(n23711) );
  OR U24109 ( .A(n23714), .B(n23715), .Z(n23713) );
  NAND U24110 ( .A(n23715), .B(n23714), .Z(n23710) );
  ANDN U24111 ( .B(B[111]), .A(n38), .Z(n23606) );
  XNOR U24112 ( .A(n23614), .B(n23716), .Z(n23607) );
  XNOR U24113 ( .A(n23613), .B(n23611), .Z(n23716) );
  AND U24114 ( .A(n23717), .B(n23718), .Z(n23611) );
  NANDN U24115 ( .A(n23719), .B(n23720), .Z(n23718) );
  NANDN U24116 ( .A(n23721), .B(n23722), .Z(n23720) );
  NANDN U24117 ( .A(n23722), .B(n23721), .Z(n23717) );
  ANDN U24118 ( .B(B[112]), .A(n39), .Z(n23613) );
  XNOR U24119 ( .A(n23621), .B(n23723), .Z(n23614) );
  XNOR U24120 ( .A(n23620), .B(n23618), .Z(n23723) );
  AND U24121 ( .A(n23724), .B(n23725), .Z(n23618) );
  NANDN U24122 ( .A(n23726), .B(n23727), .Z(n23725) );
  OR U24123 ( .A(n23728), .B(n23729), .Z(n23727) );
  NAND U24124 ( .A(n23729), .B(n23728), .Z(n23724) );
  ANDN U24125 ( .B(B[113]), .A(n40), .Z(n23620) );
  XNOR U24126 ( .A(n23628), .B(n23730), .Z(n23621) );
  XNOR U24127 ( .A(n23627), .B(n23625), .Z(n23730) );
  AND U24128 ( .A(n23731), .B(n23732), .Z(n23625) );
  NANDN U24129 ( .A(n23733), .B(n23734), .Z(n23732) );
  NAND U24130 ( .A(n23735), .B(n23736), .Z(n23734) );
  ANDN U24131 ( .B(B[114]), .A(n41), .Z(n23627) );
  XOR U24132 ( .A(n23634), .B(n23737), .Z(n23628) );
  XNOR U24133 ( .A(n23632), .B(n23635), .Z(n23737) );
  NAND U24134 ( .A(A[2]), .B(B[115]), .Z(n23635) );
  NANDN U24135 ( .A(n23738), .B(n23739), .Z(n23632) );
  AND U24136 ( .A(A[0]), .B(B[116]), .Z(n23739) );
  XNOR U24137 ( .A(n23637), .B(n23740), .Z(n23634) );
  NAND U24138 ( .A(A[0]), .B(B[117]), .Z(n23740) );
  NAND U24139 ( .A(B[116]), .B(A[1]), .Z(n23637) );
  NAND U24140 ( .A(n23741), .B(n23742), .Z(n521) );
  NANDN U24141 ( .A(n23743), .B(n23744), .Z(n23742) );
  OR U24142 ( .A(n23745), .B(n23746), .Z(n23744) );
  NAND U24143 ( .A(n23746), .B(n23745), .Z(n23741) );
  XOR U24144 ( .A(n523), .B(n522), .Z(\A1[114] ) );
  XOR U24145 ( .A(n23746), .B(n23747), .Z(n522) );
  XNOR U24146 ( .A(n23745), .B(n23743), .Z(n23747) );
  AND U24147 ( .A(n23748), .B(n23749), .Z(n23743) );
  NANDN U24148 ( .A(n23750), .B(n23751), .Z(n23749) );
  NANDN U24149 ( .A(n23752), .B(n23753), .Z(n23751) );
  NANDN U24150 ( .A(n23753), .B(n23752), .Z(n23748) );
  ANDN U24151 ( .B(B[101]), .A(n29), .Z(n23745) );
  XNOR U24152 ( .A(n23652), .B(n23754), .Z(n23746) );
  XNOR U24153 ( .A(n23651), .B(n23649), .Z(n23754) );
  AND U24154 ( .A(n23755), .B(n23756), .Z(n23649) );
  NANDN U24155 ( .A(n23757), .B(n23758), .Z(n23756) );
  OR U24156 ( .A(n23759), .B(n23760), .Z(n23758) );
  NAND U24157 ( .A(n23760), .B(n23759), .Z(n23755) );
  ANDN U24158 ( .B(B[102]), .A(n30), .Z(n23651) );
  XNOR U24159 ( .A(n23659), .B(n23761), .Z(n23652) );
  XNOR U24160 ( .A(n23658), .B(n23656), .Z(n23761) );
  AND U24161 ( .A(n23762), .B(n23763), .Z(n23656) );
  NANDN U24162 ( .A(n23764), .B(n23765), .Z(n23763) );
  NANDN U24163 ( .A(n23766), .B(n23767), .Z(n23765) );
  NANDN U24164 ( .A(n23767), .B(n23766), .Z(n23762) );
  ANDN U24165 ( .B(B[103]), .A(n31), .Z(n23658) );
  XNOR U24166 ( .A(n23666), .B(n23768), .Z(n23659) );
  XNOR U24167 ( .A(n23665), .B(n23663), .Z(n23768) );
  AND U24168 ( .A(n23769), .B(n23770), .Z(n23663) );
  NANDN U24169 ( .A(n23771), .B(n23772), .Z(n23770) );
  OR U24170 ( .A(n23773), .B(n23774), .Z(n23772) );
  NAND U24171 ( .A(n23774), .B(n23773), .Z(n23769) );
  ANDN U24172 ( .B(B[104]), .A(n32), .Z(n23665) );
  XNOR U24173 ( .A(n23673), .B(n23775), .Z(n23666) );
  XNOR U24174 ( .A(n23672), .B(n23670), .Z(n23775) );
  AND U24175 ( .A(n23776), .B(n23777), .Z(n23670) );
  NANDN U24176 ( .A(n23778), .B(n23779), .Z(n23777) );
  NANDN U24177 ( .A(n23780), .B(n23781), .Z(n23779) );
  NANDN U24178 ( .A(n23781), .B(n23780), .Z(n23776) );
  ANDN U24179 ( .B(B[105]), .A(n33), .Z(n23672) );
  XNOR U24180 ( .A(n23680), .B(n23782), .Z(n23673) );
  XNOR U24181 ( .A(n23679), .B(n23677), .Z(n23782) );
  AND U24182 ( .A(n23783), .B(n23784), .Z(n23677) );
  NANDN U24183 ( .A(n23785), .B(n23786), .Z(n23784) );
  OR U24184 ( .A(n23787), .B(n23788), .Z(n23786) );
  NAND U24185 ( .A(n23788), .B(n23787), .Z(n23783) );
  ANDN U24186 ( .B(B[106]), .A(n34), .Z(n23679) );
  XNOR U24187 ( .A(n23687), .B(n23789), .Z(n23680) );
  XNOR U24188 ( .A(n23686), .B(n23684), .Z(n23789) );
  AND U24189 ( .A(n23790), .B(n23791), .Z(n23684) );
  NANDN U24190 ( .A(n23792), .B(n23793), .Z(n23791) );
  NANDN U24191 ( .A(n23794), .B(n23795), .Z(n23793) );
  NANDN U24192 ( .A(n23795), .B(n23794), .Z(n23790) );
  ANDN U24193 ( .B(B[107]), .A(n35), .Z(n23686) );
  XNOR U24194 ( .A(n23694), .B(n23796), .Z(n23687) );
  XNOR U24195 ( .A(n23693), .B(n23691), .Z(n23796) );
  AND U24196 ( .A(n23797), .B(n23798), .Z(n23691) );
  NANDN U24197 ( .A(n23799), .B(n23800), .Z(n23798) );
  OR U24198 ( .A(n23801), .B(n23802), .Z(n23800) );
  NAND U24199 ( .A(n23802), .B(n23801), .Z(n23797) );
  ANDN U24200 ( .B(B[108]), .A(n36), .Z(n23693) );
  XNOR U24201 ( .A(n23701), .B(n23803), .Z(n23694) );
  XNOR U24202 ( .A(n23700), .B(n23698), .Z(n23803) );
  AND U24203 ( .A(n23804), .B(n23805), .Z(n23698) );
  NANDN U24204 ( .A(n23806), .B(n23807), .Z(n23805) );
  NANDN U24205 ( .A(n23808), .B(n23809), .Z(n23807) );
  NANDN U24206 ( .A(n23809), .B(n23808), .Z(n23804) );
  ANDN U24207 ( .B(B[109]), .A(n37), .Z(n23700) );
  XNOR U24208 ( .A(n23708), .B(n23810), .Z(n23701) );
  XNOR U24209 ( .A(n23707), .B(n23705), .Z(n23810) );
  AND U24210 ( .A(n23811), .B(n23812), .Z(n23705) );
  NANDN U24211 ( .A(n23813), .B(n23814), .Z(n23812) );
  OR U24212 ( .A(n23815), .B(n23816), .Z(n23814) );
  NAND U24213 ( .A(n23816), .B(n23815), .Z(n23811) );
  ANDN U24214 ( .B(B[110]), .A(n38), .Z(n23707) );
  XNOR U24215 ( .A(n23715), .B(n23817), .Z(n23708) );
  XNOR U24216 ( .A(n23714), .B(n23712), .Z(n23817) );
  AND U24217 ( .A(n23818), .B(n23819), .Z(n23712) );
  NANDN U24218 ( .A(n23820), .B(n23821), .Z(n23819) );
  NANDN U24219 ( .A(n23822), .B(n23823), .Z(n23821) );
  NANDN U24220 ( .A(n23823), .B(n23822), .Z(n23818) );
  ANDN U24221 ( .B(B[111]), .A(n39), .Z(n23714) );
  XNOR U24222 ( .A(n23722), .B(n23824), .Z(n23715) );
  XNOR U24223 ( .A(n23721), .B(n23719), .Z(n23824) );
  AND U24224 ( .A(n23825), .B(n23826), .Z(n23719) );
  NANDN U24225 ( .A(n23827), .B(n23828), .Z(n23826) );
  OR U24226 ( .A(n23829), .B(n23830), .Z(n23828) );
  NAND U24227 ( .A(n23830), .B(n23829), .Z(n23825) );
  ANDN U24228 ( .B(B[112]), .A(n40), .Z(n23721) );
  XNOR U24229 ( .A(n23729), .B(n23831), .Z(n23722) );
  XNOR U24230 ( .A(n23728), .B(n23726), .Z(n23831) );
  AND U24231 ( .A(n23832), .B(n23833), .Z(n23726) );
  NANDN U24232 ( .A(n23834), .B(n23835), .Z(n23833) );
  NAND U24233 ( .A(n23836), .B(n23837), .Z(n23835) );
  ANDN U24234 ( .B(B[113]), .A(n41), .Z(n23728) );
  XOR U24235 ( .A(n23735), .B(n23838), .Z(n23729) );
  XNOR U24236 ( .A(n23733), .B(n23736), .Z(n23838) );
  NAND U24237 ( .A(A[2]), .B(B[114]), .Z(n23736) );
  NANDN U24238 ( .A(n23839), .B(n23840), .Z(n23733) );
  AND U24239 ( .A(A[0]), .B(B[115]), .Z(n23840) );
  XNOR U24240 ( .A(n23738), .B(n23841), .Z(n23735) );
  NAND U24241 ( .A(A[0]), .B(B[116]), .Z(n23841) );
  NAND U24242 ( .A(B[115]), .B(A[1]), .Z(n23738) );
  NAND U24243 ( .A(n23842), .B(n23843), .Z(n523) );
  NANDN U24244 ( .A(n23844), .B(n23845), .Z(n23843) );
  OR U24245 ( .A(n23846), .B(n23847), .Z(n23845) );
  NAND U24246 ( .A(n23847), .B(n23846), .Z(n23842) );
  XOR U24247 ( .A(n525), .B(n524), .Z(\A1[113] ) );
  XOR U24248 ( .A(n23847), .B(n23848), .Z(n524) );
  XNOR U24249 ( .A(n23846), .B(n23844), .Z(n23848) );
  AND U24250 ( .A(n23849), .B(n23850), .Z(n23844) );
  NANDN U24251 ( .A(n23851), .B(n23852), .Z(n23850) );
  NANDN U24252 ( .A(n23853), .B(n23854), .Z(n23852) );
  NANDN U24253 ( .A(n23854), .B(n23853), .Z(n23849) );
  ANDN U24254 ( .B(A[15]), .A(n3), .Z(n23846) );
  XNOR U24255 ( .A(n23753), .B(n23855), .Z(n23847) );
  XNOR U24256 ( .A(n23752), .B(n23750), .Z(n23855) );
  AND U24257 ( .A(n23856), .B(n23857), .Z(n23750) );
  NANDN U24258 ( .A(n23858), .B(n23859), .Z(n23857) );
  OR U24259 ( .A(n23860), .B(n23861), .Z(n23859) );
  NAND U24260 ( .A(n23861), .B(n23860), .Z(n23856) );
  ANDN U24261 ( .B(B[101]), .A(n30), .Z(n23752) );
  XNOR U24262 ( .A(n23760), .B(n23862), .Z(n23753) );
  XNOR U24263 ( .A(n23759), .B(n23757), .Z(n23862) );
  AND U24264 ( .A(n23863), .B(n23864), .Z(n23757) );
  NANDN U24265 ( .A(n23865), .B(n23866), .Z(n23864) );
  NANDN U24266 ( .A(n23867), .B(n23868), .Z(n23866) );
  NANDN U24267 ( .A(n23868), .B(n23867), .Z(n23863) );
  ANDN U24268 ( .B(B[102]), .A(n31), .Z(n23759) );
  XNOR U24269 ( .A(n23767), .B(n23869), .Z(n23760) );
  XNOR U24270 ( .A(n23766), .B(n23764), .Z(n23869) );
  AND U24271 ( .A(n23870), .B(n23871), .Z(n23764) );
  NANDN U24272 ( .A(n23872), .B(n23873), .Z(n23871) );
  OR U24273 ( .A(n23874), .B(n23875), .Z(n23873) );
  NAND U24274 ( .A(n23875), .B(n23874), .Z(n23870) );
  ANDN U24275 ( .B(B[103]), .A(n32), .Z(n23766) );
  XNOR U24276 ( .A(n23774), .B(n23876), .Z(n23767) );
  XNOR U24277 ( .A(n23773), .B(n23771), .Z(n23876) );
  AND U24278 ( .A(n23877), .B(n23878), .Z(n23771) );
  NANDN U24279 ( .A(n23879), .B(n23880), .Z(n23878) );
  NANDN U24280 ( .A(n23881), .B(n23882), .Z(n23880) );
  NANDN U24281 ( .A(n23882), .B(n23881), .Z(n23877) );
  ANDN U24282 ( .B(B[104]), .A(n33), .Z(n23773) );
  XNOR U24283 ( .A(n23781), .B(n23883), .Z(n23774) );
  XNOR U24284 ( .A(n23780), .B(n23778), .Z(n23883) );
  AND U24285 ( .A(n23884), .B(n23885), .Z(n23778) );
  NANDN U24286 ( .A(n23886), .B(n23887), .Z(n23885) );
  OR U24287 ( .A(n23888), .B(n23889), .Z(n23887) );
  NAND U24288 ( .A(n23889), .B(n23888), .Z(n23884) );
  ANDN U24289 ( .B(B[105]), .A(n34), .Z(n23780) );
  XNOR U24290 ( .A(n23788), .B(n23890), .Z(n23781) );
  XNOR U24291 ( .A(n23787), .B(n23785), .Z(n23890) );
  AND U24292 ( .A(n23891), .B(n23892), .Z(n23785) );
  NANDN U24293 ( .A(n23893), .B(n23894), .Z(n23892) );
  NANDN U24294 ( .A(n23895), .B(n23896), .Z(n23894) );
  NANDN U24295 ( .A(n23896), .B(n23895), .Z(n23891) );
  ANDN U24296 ( .B(B[106]), .A(n35), .Z(n23787) );
  XNOR U24297 ( .A(n23795), .B(n23897), .Z(n23788) );
  XNOR U24298 ( .A(n23794), .B(n23792), .Z(n23897) );
  AND U24299 ( .A(n23898), .B(n23899), .Z(n23792) );
  NANDN U24300 ( .A(n23900), .B(n23901), .Z(n23899) );
  OR U24301 ( .A(n23902), .B(n23903), .Z(n23901) );
  NAND U24302 ( .A(n23903), .B(n23902), .Z(n23898) );
  ANDN U24303 ( .B(B[107]), .A(n36), .Z(n23794) );
  XNOR U24304 ( .A(n23802), .B(n23904), .Z(n23795) );
  XNOR U24305 ( .A(n23801), .B(n23799), .Z(n23904) );
  AND U24306 ( .A(n23905), .B(n23906), .Z(n23799) );
  NANDN U24307 ( .A(n23907), .B(n23908), .Z(n23906) );
  NANDN U24308 ( .A(n23909), .B(n23910), .Z(n23908) );
  NANDN U24309 ( .A(n23910), .B(n23909), .Z(n23905) );
  ANDN U24310 ( .B(B[108]), .A(n37), .Z(n23801) );
  XNOR U24311 ( .A(n23809), .B(n23911), .Z(n23802) );
  XNOR U24312 ( .A(n23808), .B(n23806), .Z(n23911) );
  AND U24313 ( .A(n23912), .B(n23913), .Z(n23806) );
  NANDN U24314 ( .A(n23914), .B(n23915), .Z(n23913) );
  OR U24315 ( .A(n23916), .B(n23917), .Z(n23915) );
  NAND U24316 ( .A(n23917), .B(n23916), .Z(n23912) );
  ANDN U24317 ( .B(B[109]), .A(n38), .Z(n23808) );
  XNOR U24318 ( .A(n23816), .B(n23918), .Z(n23809) );
  XNOR U24319 ( .A(n23815), .B(n23813), .Z(n23918) );
  AND U24320 ( .A(n23919), .B(n23920), .Z(n23813) );
  NANDN U24321 ( .A(n23921), .B(n23922), .Z(n23920) );
  NANDN U24322 ( .A(n23923), .B(n23924), .Z(n23922) );
  NANDN U24323 ( .A(n23924), .B(n23923), .Z(n23919) );
  ANDN U24324 ( .B(B[110]), .A(n39), .Z(n23815) );
  XNOR U24325 ( .A(n23823), .B(n23925), .Z(n23816) );
  XNOR U24326 ( .A(n23822), .B(n23820), .Z(n23925) );
  AND U24327 ( .A(n23926), .B(n23927), .Z(n23820) );
  NANDN U24328 ( .A(n23928), .B(n23929), .Z(n23927) );
  OR U24329 ( .A(n23930), .B(n23931), .Z(n23929) );
  NAND U24330 ( .A(n23931), .B(n23930), .Z(n23926) );
  ANDN U24331 ( .B(B[111]), .A(n40), .Z(n23822) );
  XNOR U24332 ( .A(n23830), .B(n23932), .Z(n23823) );
  XNOR U24333 ( .A(n23829), .B(n23827), .Z(n23932) );
  AND U24334 ( .A(n23933), .B(n23934), .Z(n23827) );
  NANDN U24335 ( .A(n23935), .B(n23936), .Z(n23934) );
  NAND U24336 ( .A(n23937), .B(n23938), .Z(n23936) );
  ANDN U24337 ( .B(B[112]), .A(n41), .Z(n23829) );
  XOR U24338 ( .A(n23836), .B(n23939), .Z(n23830) );
  XNOR U24339 ( .A(n23834), .B(n23837), .Z(n23939) );
  NAND U24340 ( .A(A[2]), .B(B[113]), .Z(n23837) );
  NANDN U24341 ( .A(n23940), .B(n23941), .Z(n23834) );
  AND U24342 ( .A(A[0]), .B(B[114]), .Z(n23941) );
  XNOR U24343 ( .A(n23839), .B(n23942), .Z(n23836) );
  NAND U24344 ( .A(A[0]), .B(B[115]), .Z(n23942) );
  NAND U24345 ( .A(B[114]), .B(A[1]), .Z(n23839) );
  NAND U24346 ( .A(n23943), .B(n23944), .Z(n525) );
  NANDN U24347 ( .A(n23945), .B(n23946), .Z(n23944) );
  OR U24348 ( .A(n23947), .B(n23948), .Z(n23946) );
  NAND U24349 ( .A(n23948), .B(n23947), .Z(n23943) );
  XOR U24350 ( .A(n527), .B(n526), .Z(\A1[112] ) );
  XOR U24351 ( .A(n23948), .B(n23949), .Z(n526) );
  XNOR U24352 ( .A(n23947), .B(n23945), .Z(n23949) );
  AND U24353 ( .A(n23950), .B(n23951), .Z(n23945) );
  NANDN U24354 ( .A(n23952), .B(n23953), .Z(n23951) );
  NANDN U24355 ( .A(n23954), .B(n23955), .Z(n23953) );
  NANDN U24356 ( .A(n23955), .B(n23954), .Z(n23950) );
  ANDN U24357 ( .B(A[15]), .A(n5), .Z(n23947) );
  XNOR U24358 ( .A(n23854), .B(n23956), .Z(n23948) );
  XNOR U24359 ( .A(n23853), .B(n23851), .Z(n23956) );
  AND U24360 ( .A(n23957), .B(n23958), .Z(n23851) );
  NANDN U24361 ( .A(n23959), .B(n23960), .Z(n23958) );
  OR U24362 ( .A(n23961), .B(n23962), .Z(n23960) );
  NAND U24363 ( .A(n23962), .B(n23961), .Z(n23957) );
  ANDN U24364 ( .B(A[14]), .A(n3), .Z(n23853) );
  XNOR U24365 ( .A(n23861), .B(n23963), .Z(n23854) );
  XNOR U24366 ( .A(n23860), .B(n23858), .Z(n23963) );
  AND U24367 ( .A(n23964), .B(n23965), .Z(n23858) );
  NANDN U24368 ( .A(n23966), .B(n23967), .Z(n23965) );
  NANDN U24369 ( .A(n23968), .B(n23969), .Z(n23967) );
  NANDN U24370 ( .A(n23969), .B(n23968), .Z(n23964) );
  ANDN U24371 ( .B(B[101]), .A(n31), .Z(n23860) );
  XNOR U24372 ( .A(n23868), .B(n23970), .Z(n23861) );
  XNOR U24373 ( .A(n23867), .B(n23865), .Z(n23970) );
  AND U24374 ( .A(n23971), .B(n23972), .Z(n23865) );
  NANDN U24375 ( .A(n23973), .B(n23974), .Z(n23972) );
  OR U24376 ( .A(n23975), .B(n23976), .Z(n23974) );
  NAND U24377 ( .A(n23976), .B(n23975), .Z(n23971) );
  ANDN U24378 ( .B(B[102]), .A(n32), .Z(n23867) );
  XNOR U24379 ( .A(n23875), .B(n23977), .Z(n23868) );
  XNOR U24380 ( .A(n23874), .B(n23872), .Z(n23977) );
  AND U24381 ( .A(n23978), .B(n23979), .Z(n23872) );
  NANDN U24382 ( .A(n23980), .B(n23981), .Z(n23979) );
  NANDN U24383 ( .A(n23982), .B(n23983), .Z(n23981) );
  NANDN U24384 ( .A(n23983), .B(n23982), .Z(n23978) );
  ANDN U24385 ( .B(B[103]), .A(n33), .Z(n23874) );
  XNOR U24386 ( .A(n23882), .B(n23984), .Z(n23875) );
  XNOR U24387 ( .A(n23881), .B(n23879), .Z(n23984) );
  AND U24388 ( .A(n23985), .B(n23986), .Z(n23879) );
  NANDN U24389 ( .A(n23987), .B(n23988), .Z(n23986) );
  OR U24390 ( .A(n23989), .B(n23990), .Z(n23988) );
  NAND U24391 ( .A(n23990), .B(n23989), .Z(n23985) );
  ANDN U24392 ( .B(B[104]), .A(n34), .Z(n23881) );
  XNOR U24393 ( .A(n23889), .B(n23991), .Z(n23882) );
  XNOR U24394 ( .A(n23888), .B(n23886), .Z(n23991) );
  AND U24395 ( .A(n23992), .B(n23993), .Z(n23886) );
  NANDN U24396 ( .A(n23994), .B(n23995), .Z(n23993) );
  NANDN U24397 ( .A(n23996), .B(n23997), .Z(n23995) );
  NANDN U24398 ( .A(n23997), .B(n23996), .Z(n23992) );
  ANDN U24399 ( .B(B[105]), .A(n35), .Z(n23888) );
  XNOR U24400 ( .A(n23896), .B(n23998), .Z(n23889) );
  XNOR U24401 ( .A(n23895), .B(n23893), .Z(n23998) );
  AND U24402 ( .A(n23999), .B(n24000), .Z(n23893) );
  NANDN U24403 ( .A(n24001), .B(n24002), .Z(n24000) );
  OR U24404 ( .A(n24003), .B(n24004), .Z(n24002) );
  NAND U24405 ( .A(n24004), .B(n24003), .Z(n23999) );
  ANDN U24406 ( .B(B[106]), .A(n36), .Z(n23895) );
  XNOR U24407 ( .A(n23903), .B(n24005), .Z(n23896) );
  XNOR U24408 ( .A(n23902), .B(n23900), .Z(n24005) );
  AND U24409 ( .A(n24006), .B(n24007), .Z(n23900) );
  NANDN U24410 ( .A(n24008), .B(n24009), .Z(n24007) );
  NANDN U24411 ( .A(n24010), .B(n24011), .Z(n24009) );
  NANDN U24412 ( .A(n24011), .B(n24010), .Z(n24006) );
  ANDN U24413 ( .B(B[107]), .A(n37), .Z(n23902) );
  XNOR U24414 ( .A(n23910), .B(n24012), .Z(n23903) );
  XNOR U24415 ( .A(n23909), .B(n23907), .Z(n24012) );
  AND U24416 ( .A(n24013), .B(n24014), .Z(n23907) );
  NANDN U24417 ( .A(n24015), .B(n24016), .Z(n24014) );
  OR U24418 ( .A(n24017), .B(n24018), .Z(n24016) );
  NAND U24419 ( .A(n24018), .B(n24017), .Z(n24013) );
  ANDN U24420 ( .B(B[108]), .A(n38), .Z(n23909) );
  XNOR U24421 ( .A(n23917), .B(n24019), .Z(n23910) );
  XNOR U24422 ( .A(n23916), .B(n23914), .Z(n24019) );
  AND U24423 ( .A(n24020), .B(n24021), .Z(n23914) );
  NANDN U24424 ( .A(n24022), .B(n24023), .Z(n24021) );
  NANDN U24425 ( .A(n24024), .B(n24025), .Z(n24023) );
  NANDN U24426 ( .A(n24025), .B(n24024), .Z(n24020) );
  ANDN U24427 ( .B(B[109]), .A(n39), .Z(n23916) );
  XNOR U24428 ( .A(n23924), .B(n24026), .Z(n23917) );
  XNOR U24429 ( .A(n23923), .B(n23921), .Z(n24026) );
  AND U24430 ( .A(n24027), .B(n24028), .Z(n23921) );
  NANDN U24431 ( .A(n24029), .B(n24030), .Z(n24028) );
  OR U24432 ( .A(n24031), .B(n24032), .Z(n24030) );
  NAND U24433 ( .A(n24032), .B(n24031), .Z(n24027) );
  ANDN U24434 ( .B(B[110]), .A(n40), .Z(n23923) );
  XNOR U24435 ( .A(n23931), .B(n24033), .Z(n23924) );
  XNOR U24436 ( .A(n23930), .B(n23928), .Z(n24033) );
  AND U24437 ( .A(n24034), .B(n24035), .Z(n23928) );
  NANDN U24438 ( .A(n24036), .B(n24037), .Z(n24035) );
  NAND U24439 ( .A(n24038), .B(n24039), .Z(n24037) );
  ANDN U24440 ( .B(B[111]), .A(n41), .Z(n23930) );
  XOR U24441 ( .A(n23937), .B(n24040), .Z(n23931) );
  XNOR U24442 ( .A(n23935), .B(n23938), .Z(n24040) );
  NAND U24443 ( .A(A[2]), .B(B[112]), .Z(n23938) );
  NANDN U24444 ( .A(n24041), .B(n24042), .Z(n23935) );
  AND U24445 ( .A(A[0]), .B(B[113]), .Z(n24042) );
  XNOR U24446 ( .A(n23940), .B(n24043), .Z(n23937) );
  NAND U24447 ( .A(A[0]), .B(B[114]), .Z(n24043) );
  NAND U24448 ( .A(B[113]), .B(A[1]), .Z(n23940) );
  NAND U24449 ( .A(n24044), .B(n24045), .Z(n527) );
  NANDN U24450 ( .A(n24046), .B(n24047), .Z(n24045) );
  OR U24451 ( .A(n24048), .B(n24049), .Z(n24047) );
  NAND U24452 ( .A(n24049), .B(n24048), .Z(n24044) );
  XOR U24453 ( .A(n529), .B(n528), .Z(\A1[111] ) );
  XOR U24454 ( .A(n24049), .B(n24050), .Z(n528) );
  XNOR U24455 ( .A(n24048), .B(n24046), .Z(n24050) );
  AND U24456 ( .A(n24051), .B(n24052), .Z(n24046) );
  NANDN U24457 ( .A(n24053), .B(n24054), .Z(n24052) );
  NANDN U24458 ( .A(n24055), .B(n24056), .Z(n24054) );
  NANDN U24459 ( .A(n24056), .B(n24055), .Z(n24051) );
  ANDN U24460 ( .B(B[98]), .A(n29), .Z(n24048) );
  XNOR U24461 ( .A(n23955), .B(n24057), .Z(n24049) );
  XNOR U24462 ( .A(n23954), .B(n23952), .Z(n24057) );
  AND U24463 ( .A(n24058), .B(n24059), .Z(n23952) );
  NANDN U24464 ( .A(n24060), .B(n24061), .Z(n24059) );
  OR U24465 ( .A(n24062), .B(n24063), .Z(n24061) );
  NAND U24466 ( .A(n24063), .B(n24062), .Z(n24058) );
  ANDN U24467 ( .B(A[14]), .A(n5), .Z(n23954) );
  XNOR U24468 ( .A(n23962), .B(n24064), .Z(n23955) );
  XNOR U24469 ( .A(n23961), .B(n23959), .Z(n24064) );
  AND U24470 ( .A(n24065), .B(n24066), .Z(n23959) );
  NANDN U24471 ( .A(n24067), .B(n24068), .Z(n24066) );
  NANDN U24472 ( .A(n24069), .B(n24070), .Z(n24068) );
  NANDN U24473 ( .A(n24070), .B(n24069), .Z(n24065) );
  ANDN U24474 ( .B(A[13]), .A(n3), .Z(n23961) );
  XNOR U24475 ( .A(n23969), .B(n24071), .Z(n23962) );
  XNOR U24476 ( .A(n23968), .B(n23966), .Z(n24071) );
  AND U24477 ( .A(n24072), .B(n24073), .Z(n23966) );
  NANDN U24478 ( .A(n24074), .B(n24075), .Z(n24073) );
  OR U24479 ( .A(n24076), .B(n24077), .Z(n24075) );
  NAND U24480 ( .A(n24077), .B(n24076), .Z(n24072) );
  ANDN U24481 ( .B(B[101]), .A(n32), .Z(n23968) );
  XNOR U24482 ( .A(n23976), .B(n24078), .Z(n23969) );
  XNOR U24483 ( .A(n23975), .B(n23973), .Z(n24078) );
  AND U24484 ( .A(n24079), .B(n24080), .Z(n23973) );
  NANDN U24485 ( .A(n24081), .B(n24082), .Z(n24080) );
  NANDN U24486 ( .A(n24083), .B(n24084), .Z(n24082) );
  NANDN U24487 ( .A(n24084), .B(n24083), .Z(n24079) );
  ANDN U24488 ( .B(B[102]), .A(n33), .Z(n23975) );
  XNOR U24489 ( .A(n23983), .B(n24085), .Z(n23976) );
  XNOR U24490 ( .A(n23982), .B(n23980), .Z(n24085) );
  AND U24491 ( .A(n24086), .B(n24087), .Z(n23980) );
  NANDN U24492 ( .A(n24088), .B(n24089), .Z(n24087) );
  OR U24493 ( .A(n24090), .B(n24091), .Z(n24089) );
  NAND U24494 ( .A(n24091), .B(n24090), .Z(n24086) );
  ANDN U24495 ( .B(B[103]), .A(n34), .Z(n23982) );
  XNOR U24496 ( .A(n23990), .B(n24092), .Z(n23983) );
  XNOR U24497 ( .A(n23989), .B(n23987), .Z(n24092) );
  AND U24498 ( .A(n24093), .B(n24094), .Z(n23987) );
  NANDN U24499 ( .A(n24095), .B(n24096), .Z(n24094) );
  NANDN U24500 ( .A(n24097), .B(n24098), .Z(n24096) );
  NANDN U24501 ( .A(n24098), .B(n24097), .Z(n24093) );
  ANDN U24502 ( .B(B[104]), .A(n35), .Z(n23989) );
  XNOR U24503 ( .A(n23997), .B(n24099), .Z(n23990) );
  XNOR U24504 ( .A(n23996), .B(n23994), .Z(n24099) );
  AND U24505 ( .A(n24100), .B(n24101), .Z(n23994) );
  NANDN U24506 ( .A(n24102), .B(n24103), .Z(n24101) );
  OR U24507 ( .A(n24104), .B(n24105), .Z(n24103) );
  NAND U24508 ( .A(n24105), .B(n24104), .Z(n24100) );
  ANDN U24509 ( .B(B[105]), .A(n36), .Z(n23996) );
  XNOR U24510 ( .A(n24004), .B(n24106), .Z(n23997) );
  XNOR U24511 ( .A(n24003), .B(n24001), .Z(n24106) );
  AND U24512 ( .A(n24107), .B(n24108), .Z(n24001) );
  NANDN U24513 ( .A(n24109), .B(n24110), .Z(n24108) );
  NANDN U24514 ( .A(n24111), .B(n24112), .Z(n24110) );
  NANDN U24515 ( .A(n24112), .B(n24111), .Z(n24107) );
  ANDN U24516 ( .B(B[106]), .A(n37), .Z(n24003) );
  XNOR U24517 ( .A(n24011), .B(n24113), .Z(n24004) );
  XNOR U24518 ( .A(n24010), .B(n24008), .Z(n24113) );
  AND U24519 ( .A(n24114), .B(n24115), .Z(n24008) );
  NANDN U24520 ( .A(n24116), .B(n24117), .Z(n24115) );
  OR U24521 ( .A(n24118), .B(n24119), .Z(n24117) );
  NAND U24522 ( .A(n24119), .B(n24118), .Z(n24114) );
  ANDN U24523 ( .B(B[107]), .A(n38), .Z(n24010) );
  XNOR U24524 ( .A(n24018), .B(n24120), .Z(n24011) );
  XNOR U24525 ( .A(n24017), .B(n24015), .Z(n24120) );
  AND U24526 ( .A(n24121), .B(n24122), .Z(n24015) );
  NANDN U24527 ( .A(n24123), .B(n24124), .Z(n24122) );
  NANDN U24528 ( .A(n24125), .B(n24126), .Z(n24124) );
  NANDN U24529 ( .A(n24126), .B(n24125), .Z(n24121) );
  ANDN U24530 ( .B(B[108]), .A(n39), .Z(n24017) );
  XNOR U24531 ( .A(n24025), .B(n24127), .Z(n24018) );
  XNOR U24532 ( .A(n24024), .B(n24022), .Z(n24127) );
  AND U24533 ( .A(n24128), .B(n24129), .Z(n24022) );
  NANDN U24534 ( .A(n24130), .B(n24131), .Z(n24129) );
  OR U24535 ( .A(n24132), .B(n24133), .Z(n24131) );
  NAND U24536 ( .A(n24133), .B(n24132), .Z(n24128) );
  ANDN U24537 ( .B(B[109]), .A(n40), .Z(n24024) );
  XNOR U24538 ( .A(n24032), .B(n24134), .Z(n24025) );
  XNOR U24539 ( .A(n24031), .B(n24029), .Z(n24134) );
  AND U24540 ( .A(n24135), .B(n24136), .Z(n24029) );
  NANDN U24541 ( .A(n24137), .B(n24138), .Z(n24136) );
  NAND U24542 ( .A(n24139), .B(n24140), .Z(n24138) );
  ANDN U24543 ( .B(B[110]), .A(n41), .Z(n24031) );
  XOR U24544 ( .A(n24038), .B(n24141), .Z(n24032) );
  XNOR U24545 ( .A(n24036), .B(n24039), .Z(n24141) );
  NAND U24546 ( .A(A[2]), .B(B[111]), .Z(n24039) );
  NANDN U24547 ( .A(n24142), .B(n24143), .Z(n24036) );
  AND U24548 ( .A(A[0]), .B(B[112]), .Z(n24143) );
  XNOR U24549 ( .A(n24041), .B(n24144), .Z(n24038) );
  NAND U24550 ( .A(A[0]), .B(B[113]), .Z(n24144) );
  NAND U24551 ( .A(B[112]), .B(A[1]), .Z(n24041) );
  NAND U24552 ( .A(n24145), .B(n24146), .Z(n529) );
  NANDN U24553 ( .A(n24147), .B(n24148), .Z(n24146) );
  OR U24554 ( .A(n24149), .B(n24150), .Z(n24148) );
  NAND U24555 ( .A(n24150), .B(n24149), .Z(n24145) );
  XOR U24556 ( .A(n531), .B(n530), .Z(\A1[110] ) );
  XOR U24557 ( .A(n24150), .B(n24151), .Z(n530) );
  XNOR U24558 ( .A(n24149), .B(n24147), .Z(n24151) );
  AND U24559 ( .A(n24152), .B(n24153), .Z(n24147) );
  NANDN U24560 ( .A(n24154), .B(n24155), .Z(n24153) );
  NANDN U24561 ( .A(n24156), .B(n24157), .Z(n24155) );
  NANDN U24562 ( .A(n24157), .B(n24156), .Z(n24152) );
  ANDN U24563 ( .B(B[97]), .A(n29), .Z(n24149) );
  XNOR U24564 ( .A(n24056), .B(n24158), .Z(n24150) );
  XNOR U24565 ( .A(n24055), .B(n24053), .Z(n24158) );
  AND U24566 ( .A(n24159), .B(n24160), .Z(n24053) );
  NANDN U24567 ( .A(n24161), .B(n24162), .Z(n24160) );
  OR U24568 ( .A(n24163), .B(n24164), .Z(n24162) );
  NAND U24569 ( .A(n24164), .B(n24163), .Z(n24159) );
  ANDN U24570 ( .B(B[98]), .A(n30), .Z(n24055) );
  XNOR U24571 ( .A(n24063), .B(n24165), .Z(n24056) );
  XNOR U24572 ( .A(n24062), .B(n24060), .Z(n24165) );
  AND U24573 ( .A(n24166), .B(n24167), .Z(n24060) );
  NANDN U24574 ( .A(n24168), .B(n24169), .Z(n24167) );
  NANDN U24575 ( .A(n24170), .B(n24171), .Z(n24169) );
  NANDN U24576 ( .A(n24171), .B(n24170), .Z(n24166) );
  ANDN U24577 ( .B(A[13]), .A(n5), .Z(n24062) );
  XNOR U24578 ( .A(n24070), .B(n24172), .Z(n24063) );
  XNOR U24579 ( .A(n24069), .B(n24067), .Z(n24172) );
  AND U24580 ( .A(n24173), .B(n24174), .Z(n24067) );
  NANDN U24581 ( .A(n24175), .B(n24176), .Z(n24174) );
  OR U24582 ( .A(n24177), .B(n24178), .Z(n24176) );
  NAND U24583 ( .A(n24178), .B(n24177), .Z(n24173) );
  ANDN U24584 ( .B(A[12]), .A(n3), .Z(n24069) );
  XNOR U24585 ( .A(n24077), .B(n24179), .Z(n24070) );
  XNOR U24586 ( .A(n24076), .B(n24074), .Z(n24179) );
  AND U24587 ( .A(n24180), .B(n24181), .Z(n24074) );
  NANDN U24588 ( .A(n24182), .B(n24183), .Z(n24181) );
  NANDN U24589 ( .A(n24184), .B(n24185), .Z(n24183) );
  NANDN U24590 ( .A(n24185), .B(n24184), .Z(n24180) );
  ANDN U24591 ( .B(B[101]), .A(n33), .Z(n24076) );
  XNOR U24592 ( .A(n24084), .B(n24186), .Z(n24077) );
  XNOR U24593 ( .A(n24083), .B(n24081), .Z(n24186) );
  AND U24594 ( .A(n24187), .B(n24188), .Z(n24081) );
  NANDN U24595 ( .A(n24189), .B(n24190), .Z(n24188) );
  OR U24596 ( .A(n24191), .B(n24192), .Z(n24190) );
  NAND U24597 ( .A(n24192), .B(n24191), .Z(n24187) );
  ANDN U24598 ( .B(B[102]), .A(n34), .Z(n24083) );
  XNOR U24599 ( .A(n24091), .B(n24193), .Z(n24084) );
  XNOR U24600 ( .A(n24090), .B(n24088), .Z(n24193) );
  AND U24601 ( .A(n24194), .B(n24195), .Z(n24088) );
  NANDN U24602 ( .A(n24196), .B(n24197), .Z(n24195) );
  NANDN U24603 ( .A(n24198), .B(n24199), .Z(n24197) );
  NANDN U24604 ( .A(n24199), .B(n24198), .Z(n24194) );
  ANDN U24605 ( .B(B[103]), .A(n35), .Z(n24090) );
  XNOR U24606 ( .A(n24098), .B(n24200), .Z(n24091) );
  XNOR U24607 ( .A(n24097), .B(n24095), .Z(n24200) );
  AND U24608 ( .A(n24201), .B(n24202), .Z(n24095) );
  NANDN U24609 ( .A(n24203), .B(n24204), .Z(n24202) );
  OR U24610 ( .A(n24205), .B(n24206), .Z(n24204) );
  NAND U24611 ( .A(n24206), .B(n24205), .Z(n24201) );
  ANDN U24612 ( .B(B[104]), .A(n36), .Z(n24097) );
  XNOR U24613 ( .A(n24105), .B(n24207), .Z(n24098) );
  XNOR U24614 ( .A(n24104), .B(n24102), .Z(n24207) );
  AND U24615 ( .A(n24208), .B(n24209), .Z(n24102) );
  NANDN U24616 ( .A(n24210), .B(n24211), .Z(n24209) );
  NANDN U24617 ( .A(n24212), .B(n24213), .Z(n24211) );
  NANDN U24618 ( .A(n24213), .B(n24212), .Z(n24208) );
  ANDN U24619 ( .B(B[105]), .A(n37), .Z(n24104) );
  XNOR U24620 ( .A(n24112), .B(n24214), .Z(n24105) );
  XNOR U24621 ( .A(n24111), .B(n24109), .Z(n24214) );
  AND U24622 ( .A(n24215), .B(n24216), .Z(n24109) );
  NANDN U24623 ( .A(n24217), .B(n24218), .Z(n24216) );
  OR U24624 ( .A(n24219), .B(n24220), .Z(n24218) );
  NAND U24625 ( .A(n24220), .B(n24219), .Z(n24215) );
  ANDN U24626 ( .B(B[106]), .A(n38), .Z(n24111) );
  XNOR U24627 ( .A(n24119), .B(n24221), .Z(n24112) );
  XNOR U24628 ( .A(n24118), .B(n24116), .Z(n24221) );
  AND U24629 ( .A(n24222), .B(n24223), .Z(n24116) );
  NANDN U24630 ( .A(n24224), .B(n24225), .Z(n24223) );
  NANDN U24631 ( .A(n24226), .B(n24227), .Z(n24225) );
  NANDN U24632 ( .A(n24227), .B(n24226), .Z(n24222) );
  ANDN U24633 ( .B(B[107]), .A(n39), .Z(n24118) );
  XNOR U24634 ( .A(n24126), .B(n24228), .Z(n24119) );
  XNOR U24635 ( .A(n24125), .B(n24123), .Z(n24228) );
  AND U24636 ( .A(n24229), .B(n24230), .Z(n24123) );
  NANDN U24637 ( .A(n24231), .B(n24232), .Z(n24230) );
  OR U24638 ( .A(n24233), .B(n24234), .Z(n24232) );
  NAND U24639 ( .A(n24234), .B(n24233), .Z(n24229) );
  ANDN U24640 ( .B(B[108]), .A(n40), .Z(n24125) );
  XNOR U24641 ( .A(n24133), .B(n24235), .Z(n24126) );
  XNOR U24642 ( .A(n24132), .B(n24130), .Z(n24235) );
  AND U24643 ( .A(n24236), .B(n24237), .Z(n24130) );
  NANDN U24644 ( .A(n24238), .B(n24239), .Z(n24237) );
  NAND U24645 ( .A(n24240), .B(n24241), .Z(n24239) );
  ANDN U24646 ( .B(B[109]), .A(n41), .Z(n24132) );
  XOR U24647 ( .A(n24139), .B(n24242), .Z(n24133) );
  XNOR U24648 ( .A(n24137), .B(n24140), .Z(n24242) );
  NAND U24649 ( .A(A[2]), .B(B[110]), .Z(n24140) );
  NANDN U24650 ( .A(n24243), .B(n24244), .Z(n24137) );
  AND U24651 ( .A(A[0]), .B(B[111]), .Z(n24244) );
  XNOR U24652 ( .A(n24142), .B(n24245), .Z(n24139) );
  NAND U24653 ( .A(A[0]), .B(B[112]), .Z(n24245) );
  NAND U24654 ( .A(B[111]), .B(A[1]), .Z(n24142) );
  NAND U24655 ( .A(n24246), .B(n24247), .Z(n531) );
  NANDN U24656 ( .A(n24248), .B(n24249), .Z(n24247) );
  OR U24657 ( .A(n24250), .B(n24251), .Z(n24249) );
  NAND U24658 ( .A(n24251), .B(n24250), .Z(n24246) );
  XNOR U24659 ( .A(n23166), .B(n24252), .Z(\A1[10] ) );
  XNOR U24660 ( .A(n23164), .B(n23167), .Z(n24252) );
  AND U24661 ( .A(n24253), .B(n24254), .Z(n23167) );
  NANDN U24662 ( .A(n556), .B(n24255), .Z(n24254) );
  NANDN U24663 ( .A(n554), .B(n24256), .Z(n24255) );
  NAND U24664 ( .A(A[11]), .B(B[0]), .Z(n556) );
  NAND U24665 ( .A(n24), .B(n554), .Z(n24253) );
  XOR U24666 ( .A(n24257), .B(n24258), .Z(n554) );
  XNOR U24667 ( .A(n24259), .B(n24260), .Z(n24258) );
  AND U24668 ( .A(n24261), .B(n24262), .Z(n24256) );
  NANDN U24669 ( .A(n965), .B(n24263), .Z(n24262) );
  NANDN U24670 ( .A(n963), .B(n966), .Z(n24263) );
  NAND U24671 ( .A(A[10]), .B(B[0]), .Z(n965) );
  NANDN U24672 ( .A(n966), .B(n963), .Z(n24261) );
  XOR U24673 ( .A(n24264), .B(n24265), .Z(n963) );
  XNOR U24674 ( .A(n24266), .B(n24267), .Z(n24265) );
  AND U24675 ( .A(n24268), .B(n24269), .Z(n966) );
  NANDN U24676 ( .A(n1935), .B(n24270), .Z(n24269) );
  NANDN U24677 ( .A(n1933), .B(n24271), .Z(n24270) );
  NAND U24678 ( .A(A[9]), .B(B[0]), .Z(n1935) );
  NAND U24679 ( .A(n25), .B(n1933), .Z(n24268) );
  XOR U24680 ( .A(n24272), .B(n24273), .Z(n1933) );
  XNOR U24681 ( .A(n24274), .B(n24275), .Z(n24273) );
  AND U24682 ( .A(n24276), .B(n24277), .Z(n24271) );
  NANDN U24683 ( .A(n2948), .B(n24278), .Z(n24277) );
  NANDN U24684 ( .A(n2946), .B(n2949), .Z(n24278) );
  NAND U24685 ( .A(A[8]), .B(B[0]), .Z(n2948) );
  NANDN U24686 ( .A(n2949), .B(n2946), .Z(n24276) );
  XOR U24687 ( .A(n24279), .B(n24280), .Z(n2946) );
  XNOR U24688 ( .A(n24281), .B(n24282), .Z(n24280) );
  AND U24689 ( .A(n24283), .B(n24284), .Z(n2949) );
  NANDN U24690 ( .A(n3962), .B(n24285), .Z(n24284) );
  NANDN U24691 ( .A(n3960), .B(n24286), .Z(n24285) );
  NAND U24692 ( .A(A[7]), .B(B[0]), .Z(n3962) );
  NAND U24693 ( .A(n26), .B(n3960), .Z(n24283) );
  XOR U24694 ( .A(n24287), .B(n24288), .Z(n3960) );
  XNOR U24695 ( .A(n24289), .B(n24290), .Z(n24288) );
  AND U24696 ( .A(n24291), .B(n24292), .Z(n24286) );
  NANDN U24697 ( .A(n4975), .B(n24293), .Z(n24292) );
  NANDN U24698 ( .A(n4973), .B(n4976), .Z(n24293) );
  NAND U24699 ( .A(A[6]), .B(B[0]), .Z(n4975) );
  NANDN U24700 ( .A(n4976), .B(n4973), .Z(n24291) );
  XOR U24701 ( .A(n24294), .B(n24295), .Z(n4973) );
  XNOR U24702 ( .A(n24296), .B(n24297), .Z(n24295) );
  AND U24703 ( .A(n24298), .B(n24299), .Z(n4976) );
  NANDN U24704 ( .A(n5989), .B(n24300), .Z(n24299) );
  NANDN U24705 ( .A(n5987), .B(n24301), .Z(n24300) );
  NAND U24706 ( .A(A[5]), .B(B[0]), .Z(n5989) );
  NAND U24707 ( .A(n27), .B(n5987), .Z(n24298) );
  XOR U24708 ( .A(n24302), .B(n24303), .Z(n5987) );
  XNOR U24709 ( .A(n24304), .B(n24305), .Z(n24303) );
  AND U24710 ( .A(n24306), .B(n24307), .Z(n24301) );
  NANDN U24711 ( .A(n7002), .B(n24308), .Z(n24307) );
  NANDN U24712 ( .A(n7000), .B(n7003), .Z(n24308) );
  NAND U24713 ( .A(A[4]), .B(B[0]), .Z(n7002) );
  NANDN U24714 ( .A(n7003), .B(n7000), .Z(n24306) );
  XOR U24715 ( .A(n24309), .B(n24310), .Z(n7000) );
  XNOR U24716 ( .A(n24311), .B(n24312), .Z(n24310) );
  AND U24717 ( .A(n24313), .B(n24314), .Z(n7003) );
  NANDN U24718 ( .A(n14291), .B(n24315), .Z(n24314) );
  OR U24719 ( .A(n14290), .B(n14288), .Z(n24315) );
  AND U24720 ( .A(n24316), .B(n24317), .Z(n14291) );
  NANDN U24721 ( .A(n24318), .B(n24319), .Z(n24317) );
  OR U24722 ( .A(n24320), .B(n28), .Z(n24319) );
  NAND U24723 ( .A(n28), .B(n24320), .Z(n24316) );
  NAND U24724 ( .A(n14288), .B(n14290), .Z(n24313) );
  ANDN U24725 ( .B(B[0]), .A(n41), .Z(n14290) );
  XOR U24726 ( .A(n24322), .B(n24323), .Z(n14288) );
  XNOR U24727 ( .A(n24324), .B(n24325), .Z(n24323) );
  NAND U24728 ( .A(A[12]), .B(B[0]), .Z(n23164) );
  XOR U24729 ( .A(n23174), .B(n24326), .Z(n23166) );
  XNOR U24730 ( .A(n23173), .B(n23171), .Z(n24326) );
  AND U24731 ( .A(n24327), .B(n24328), .Z(n23171) );
  NANDN U24732 ( .A(n24260), .B(n24329), .Z(n24328) );
  AND U24733 ( .A(n24330), .B(n24331), .Z(n24260) );
  NANDN U24734 ( .A(n24267), .B(n24332), .Z(n24331) );
  OR U24735 ( .A(n24266), .B(n24264), .Z(n24332) );
  AND U24736 ( .A(n24333), .B(n24334), .Z(n24267) );
  NANDN U24737 ( .A(n24275), .B(n24335), .Z(n24334) );
  AND U24738 ( .A(n24336), .B(n24337), .Z(n24275) );
  NANDN U24739 ( .A(n24282), .B(n24338), .Z(n24337) );
  OR U24740 ( .A(n24281), .B(n24279), .Z(n24338) );
  AND U24741 ( .A(n24339), .B(n24340), .Z(n24282) );
  NANDN U24742 ( .A(n24290), .B(n24341), .Z(n24340) );
  AND U24743 ( .A(n24342), .B(n24343), .Z(n24290) );
  NANDN U24744 ( .A(n24297), .B(n24344), .Z(n24343) );
  OR U24745 ( .A(n24296), .B(n24294), .Z(n24344) );
  AND U24746 ( .A(n24345), .B(n24346), .Z(n24297) );
  NANDN U24747 ( .A(n24305), .B(n24347), .Z(n24346) );
  AND U24748 ( .A(n24348), .B(n24349), .Z(n24305) );
  NANDN U24749 ( .A(n24312), .B(n24350), .Z(n24349) );
  OR U24750 ( .A(n24311), .B(n24309), .Z(n24350) );
  AND U24751 ( .A(n24351), .B(n24352), .Z(n24312) );
  NANDN U24752 ( .A(n24324), .B(n24353), .Z(n24352) );
  NAND U24753 ( .A(n24322), .B(n24325), .Z(n24353) );
  NANDN U24754 ( .A(n24354), .B(n24355), .Z(n24324) );
  AND U24755 ( .A(A[0]), .B(B[2]), .Z(n24355) );
  XNOR U24756 ( .A(n24356), .B(n24357), .Z(n24322) );
  NAND U24757 ( .A(A[0]), .B(B[3]), .Z(n24357) );
  NAND U24758 ( .A(B[1]), .B(A[2]), .Z(n24325) );
  NAND U24759 ( .A(n24309), .B(n24311), .Z(n24348) );
  ANDN U24760 ( .B(B[1]), .A(n41), .Z(n24311) );
  XOR U24761 ( .A(n24358), .B(n24359), .Z(n24309) );
  XNOR U24762 ( .A(n24360), .B(n24361), .Z(n24359) );
  NAND U24763 ( .A(n24302), .B(n24304), .Z(n24345) );
  ANDN U24764 ( .B(B[1]), .A(n40), .Z(n24304) );
  XOR U24765 ( .A(n24362), .B(n24363), .Z(n24302) );
  XNOR U24766 ( .A(n24364), .B(n24365), .Z(n24363) );
  NAND U24767 ( .A(n24294), .B(n24296), .Z(n24342) );
  ANDN U24768 ( .B(B[1]), .A(n39), .Z(n24296) );
  XNOR U24769 ( .A(n24366), .B(n24367), .Z(n24294) );
  XNOR U24770 ( .A(n24368), .B(n24369), .Z(n24367) );
  NAND U24771 ( .A(n24287), .B(n24289), .Z(n24339) );
  ANDN U24772 ( .B(B[1]), .A(n38), .Z(n24289) );
  XOR U24773 ( .A(n24370), .B(n24371), .Z(n24287) );
  XNOR U24774 ( .A(n24372), .B(n24373), .Z(n24371) );
  NAND U24775 ( .A(n24279), .B(n24281), .Z(n24336) );
  ANDN U24776 ( .B(B[1]), .A(n37), .Z(n24281) );
  XNOR U24777 ( .A(n24374), .B(n24375), .Z(n24279) );
  XNOR U24778 ( .A(n24376), .B(n24377), .Z(n24375) );
  NAND U24779 ( .A(n24272), .B(n24274), .Z(n24333) );
  ANDN U24780 ( .B(B[1]), .A(n36), .Z(n24274) );
  XOR U24781 ( .A(n24378), .B(n24379), .Z(n24272) );
  XNOR U24782 ( .A(n24380), .B(n24381), .Z(n24379) );
  NAND U24783 ( .A(n24264), .B(n24266), .Z(n24330) );
  ANDN U24784 ( .B(B[1]), .A(n35), .Z(n24266) );
  XNOR U24785 ( .A(n24382), .B(n24383), .Z(n24264) );
  XNOR U24786 ( .A(n24384), .B(n24385), .Z(n24383) );
  NAND U24787 ( .A(n24257), .B(n24259), .Z(n24327) );
  ANDN U24788 ( .B(B[1]), .A(n34), .Z(n24259) );
  XOR U24789 ( .A(n24386), .B(n24387), .Z(n24257) );
  XNOR U24790 ( .A(n24388), .B(n24389), .Z(n24387) );
  ANDN U24791 ( .B(B[1]), .A(n33), .Z(n23173) );
  XNOR U24792 ( .A(n23181), .B(n24390), .Z(n23174) );
  XNOR U24793 ( .A(n23180), .B(n23178), .Z(n24390) );
  AND U24794 ( .A(n24391), .B(n24392), .Z(n23178) );
  NANDN U24795 ( .A(n24389), .B(n24393), .Z(n24392) );
  OR U24796 ( .A(n24388), .B(n24386), .Z(n24393) );
  AND U24797 ( .A(n24394), .B(n24395), .Z(n24389) );
  NANDN U24798 ( .A(n24385), .B(n24396), .Z(n24395) );
  NANDN U24799 ( .A(n24384), .B(n24382), .Z(n24396) );
  AND U24800 ( .A(n24397), .B(n24398), .Z(n24385) );
  NANDN U24801 ( .A(n24381), .B(n24399), .Z(n24398) );
  OR U24802 ( .A(n24380), .B(n24378), .Z(n24399) );
  AND U24803 ( .A(n24400), .B(n24401), .Z(n24381) );
  NANDN U24804 ( .A(n24377), .B(n24402), .Z(n24401) );
  NANDN U24805 ( .A(n24376), .B(n24374), .Z(n24402) );
  AND U24806 ( .A(n24403), .B(n24404), .Z(n24377) );
  NANDN U24807 ( .A(n24373), .B(n24405), .Z(n24404) );
  OR U24808 ( .A(n24372), .B(n24370), .Z(n24405) );
  AND U24809 ( .A(n24406), .B(n24407), .Z(n24373) );
  NANDN U24810 ( .A(n24369), .B(n24408), .Z(n24407) );
  NANDN U24811 ( .A(n24368), .B(n24366), .Z(n24408) );
  AND U24812 ( .A(n24409), .B(n24410), .Z(n24369) );
  NANDN U24813 ( .A(n24365), .B(n24411), .Z(n24410) );
  OR U24814 ( .A(n24364), .B(n24362), .Z(n24411) );
  AND U24815 ( .A(n24412), .B(n24413), .Z(n24365) );
  NANDN U24816 ( .A(n24360), .B(n24414), .Z(n24413) );
  NAND U24817 ( .A(n24358), .B(n24361), .Z(n24414) );
  NANDN U24818 ( .A(n24356), .B(n24415), .Z(n24360) );
  AND U24819 ( .A(A[0]), .B(B[3]), .Z(n24415) );
  NAND U24820 ( .A(B[2]), .B(A[1]), .Z(n24356) );
  XNOR U24821 ( .A(n24416), .B(n24417), .Z(n24358) );
  NAND U24822 ( .A(A[0]), .B(B[4]), .Z(n24417) );
  NAND U24823 ( .A(A[2]), .B(B[2]), .Z(n24361) );
  NAND U24824 ( .A(n24362), .B(n24364), .Z(n24409) );
  ANDN U24825 ( .B(B[2]), .A(n41), .Z(n24364) );
  XOR U24826 ( .A(n24418), .B(n24419), .Z(n24362) );
  XNOR U24827 ( .A(n24420), .B(n24421), .Z(n24419) );
  NANDN U24828 ( .A(n24366), .B(n24368), .Z(n24406) );
  ANDN U24829 ( .B(B[2]), .A(n40), .Z(n24368) );
  XNOR U24830 ( .A(n24422), .B(n24423), .Z(n24366) );
  XNOR U24831 ( .A(n24424), .B(n24425), .Z(n24423) );
  NAND U24832 ( .A(n24370), .B(n24372), .Z(n24403) );
  ANDN U24833 ( .B(B[2]), .A(n39), .Z(n24372) );
  XNOR U24834 ( .A(n24426), .B(n24427), .Z(n24370) );
  XNOR U24835 ( .A(n24428), .B(n24429), .Z(n24427) );
  NANDN U24836 ( .A(n24374), .B(n24376), .Z(n24400) );
  ANDN U24837 ( .B(B[2]), .A(n38), .Z(n24376) );
  XNOR U24838 ( .A(n24430), .B(n24431), .Z(n24374) );
  XNOR U24839 ( .A(n24432), .B(n24433), .Z(n24431) );
  NAND U24840 ( .A(n24378), .B(n24380), .Z(n24397) );
  ANDN U24841 ( .B(B[2]), .A(n37), .Z(n24380) );
  XNOR U24842 ( .A(n24434), .B(n24435), .Z(n24378) );
  XNOR U24843 ( .A(n24436), .B(n24437), .Z(n24435) );
  NANDN U24844 ( .A(n24382), .B(n24384), .Z(n24394) );
  ANDN U24845 ( .B(B[2]), .A(n36), .Z(n24384) );
  XNOR U24846 ( .A(n24438), .B(n24439), .Z(n24382) );
  XNOR U24847 ( .A(n24440), .B(n24441), .Z(n24439) );
  NAND U24848 ( .A(n24386), .B(n24388), .Z(n24391) );
  ANDN U24849 ( .B(B[2]), .A(n35), .Z(n24388) );
  XNOR U24850 ( .A(n24442), .B(n24443), .Z(n24386) );
  XNOR U24851 ( .A(n24444), .B(n24445), .Z(n24443) );
  ANDN U24852 ( .B(B[2]), .A(n34), .Z(n23180) );
  XNOR U24853 ( .A(n23188), .B(n24446), .Z(n23181) );
  XNOR U24854 ( .A(n23187), .B(n23185), .Z(n24446) );
  AND U24855 ( .A(n24447), .B(n24448), .Z(n23185) );
  NANDN U24856 ( .A(n24445), .B(n24449), .Z(n24448) );
  NANDN U24857 ( .A(n24444), .B(n24442), .Z(n24449) );
  AND U24858 ( .A(n24450), .B(n24451), .Z(n24445) );
  NANDN U24859 ( .A(n24441), .B(n24452), .Z(n24451) );
  OR U24860 ( .A(n24440), .B(n24438), .Z(n24452) );
  AND U24861 ( .A(n24453), .B(n24454), .Z(n24441) );
  NANDN U24862 ( .A(n24437), .B(n24455), .Z(n24454) );
  NANDN U24863 ( .A(n24436), .B(n24434), .Z(n24455) );
  AND U24864 ( .A(n24456), .B(n24457), .Z(n24437) );
  NANDN U24865 ( .A(n24433), .B(n24458), .Z(n24457) );
  OR U24866 ( .A(n24432), .B(n24430), .Z(n24458) );
  AND U24867 ( .A(n24459), .B(n24460), .Z(n24433) );
  NANDN U24868 ( .A(n24429), .B(n24461), .Z(n24460) );
  NANDN U24869 ( .A(n24428), .B(n24426), .Z(n24461) );
  AND U24870 ( .A(n24462), .B(n24463), .Z(n24429) );
  NANDN U24871 ( .A(n24425), .B(n24464), .Z(n24463) );
  OR U24872 ( .A(n24424), .B(n24422), .Z(n24464) );
  AND U24873 ( .A(n24465), .B(n24466), .Z(n24425) );
  NANDN U24874 ( .A(n24420), .B(n24467), .Z(n24466) );
  NAND U24875 ( .A(n24418), .B(n24421), .Z(n24467) );
  NANDN U24876 ( .A(n24416), .B(n24468), .Z(n24420) );
  AND U24877 ( .A(A[0]), .B(B[4]), .Z(n24468) );
  NAND U24878 ( .A(B[3]), .B(A[1]), .Z(n24416) );
  XNOR U24879 ( .A(n24469), .B(n24470), .Z(n24418) );
  NAND U24880 ( .A(A[0]), .B(B[5]), .Z(n24470) );
  NAND U24881 ( .A(A[2]), .B(B[3]), .Z(n24421) );
  NAND U24882 ( .A(n24422), .B(n24424), .Z(n24462) );
  ANDN U24883 ( .B(B[3]), .A(n41), .Z(n24424) );
  XOR U24884 ( .A(n24471), .B(n24472), .Z(n24422) );
  XNOR U24885 ( .A(n24473), .B(n24474), .Z(n24472) );
  NANDN U24886 ( .A(n24426), .B(n24428), .Z(n24459) );
  ANDN U24887 ( .B(B[3]), .A(n40), .Z(n24428) );
  XNOR U24888 ( .A(n24475), .B(n24476), .Z(n24426) );
  XNOR U24889 ( .A(n24477), .B(n24478), .Z(n24476) );
  NAND U24890 ( .A(n24430), .B(n24432), .Z(n24456) );
  ANDN U24891 ( .B(B[3]), .A(n39), .Z(n24432) );
  XNOR U24892 ( .A(n24479), .B(n24480), .Z(n24430) );
  XNOR U24893 ( .A(n24481), .B(n24482), .Z(n24480) );
  NANDN U24894 ( .A(n24434), .B(n24436), .Z(n24453) );
  ANDN U24895 ( .B(B[3]), .A(n38), .Z(n24436) );
  XNOR U24896 ( .A(n24483), .B(n24484), .Z(n24434) );
  XNOR U24897 ( .A(n24485), .B(n24486), .Z(n24484) );
  NAND U24898 ( .A(n24438), .B(n24440), .Z(n24450) );
  ANDN U24899 ( .B(B[3]), .A(n37), .Z(n24440) );
  XNOR U24900 ( .A(n24487), .B(n24488), .Z(n24438) );
  XNOR U24901 ( .A(n24489), .B(n24490), .Z(n24488) );
  NANDN U24902 ( .A(n24442), .B(n24444), .Z(n24447) );
  ANDN U24903 ( .B(B[3]), .A(n36), .Z(n24444) );
  XNOR U24904 ( .A(n24491), .B(n24492), .Z(n24442) );
  XNOR U24905 ( .A(n24493), .B(n24494), .Z(n24492) );
  ANDN U24906 ( .B(B[3]), .A(n35), .Z(n23187) );
  XNOR U24907 ( .A(n23195), .B(n24495), .Z(n23188) );
  XNOR U24908 ( .A(n23194), .B(n23192), .Z(n24495) );
  AND U24909 ( .A(n24496), .B(n24497), .Z(n23192) );
  NANDN U24910 ( .A(n24494), .B(n24498), .Z(n24497) );
  OR U24911 ( .A(n24493), .B(n24491), .Z(n24498) );
  AND U24912 ( .A(n24499), .B(n24500), .Z(n24494) );
  NANDN U24913 ( .A(n24490), .B(n24501), .Z(n24500) );
  NANDN U24914 ( .A(n24489), .B(n24487), .Z(n24501) );
  AND U24915 ( .A(n24502), .B(n24503), .Z(n24490) );
  NANDN U24916 ( .A(n24486), .B(n24504), .Z(n24503) );
  OR U24917 ( .A(n24485), .B(n24483), .Z(n24504) );
  AND U24918 ( .A(n24505), .B(n24506), .Z(n24486) );
  NANDN U24919 ( .A(n24482), .B(n24507), .Z(n24506) );
  NANDN U24920 ( .A(n24481), .B(n24479), .Z(n24507) );
  AND U24921 ( .A(n24508), .B(n24509), .Z(n24482) );
  NANDN U24922 ( .A(n24478), .B(n24510), .Z(n24509) );
  OR U24923 ( .A(n24477), .B(n24475), .Z(n24510) );
  AND U24924 ( .A(n24511), .B(n24512), .Z(n24478) );
  NANDN U24925 ( .A(n24473), .B(n24513), .Z(n24512) );
  NAND U24926 ( .A(n24471), .B(n24474), .Z(n24513) );
  NANDN U24927 ( .A(n24469), .B(n24514), .Z(n24473) );
  AND U24928 ( .A(A[0]), .B(B[5]), .Z(n24514) );
  NAND U24929 ( .A(B[4]), .B(A[1]), .Z(n24469) );
  XNOR U24930 ( .A(n24515), .B(n24516), .Z(n24471) );
  NAND U24931 ( .A(A[0]), .B(B[6]), .Z(n24516) );
  NAND U24932 ( .A(A[2]), .B(B[4]), .Z(n24474) );
  NAND U24933 ( .A(n24475), .B(n24477), .Z(n24508) );
  ANDN U24934 ( .B(B[4]), .A(n41), .Z(n24477) );
  XOR U24935 ( .A(n24517), .B(n24518), .Z(n24475) );
  XNOR U24936 ( .A(n24519), .B(n24520), .Z(n24518) );
  NANDN U24937 ( .A(n24479), .B(n24481), .Z(n24505) );
  ANDN U24938 ( .B(B[4]), .A(n40), .Z(n24481) );
  XNOR U24939 ( .A(n24521), .B(n24522), .Z(n24479) );
  XNOR U24940 ( .A(n24523), .B(n24524), .Z(n24522) );
  NAND U24941 ( .A(n24483), .B(n24485), .Z(n24502) );
  ANDN U24942 ( .B(B[4]), .A(n39), .Z(n24485) );
  XNOR U24943 ( .A(n24525), .B(n24526), .Z(n24483) );
  XNOR U24944 ( .A(n24527), .B(n24528), .Z(n24526) );
  NANDN U24945 ( .A(n24487), .B(n24489), .Z(n24499) );
  ANDN U24946 ( .B(B[4]), .A(n38), .Z(n24489) );
  XNOR U24947 ( .A(n24529), .B(n24530), .Z(n24487) );
  XNOR U24948 ( .A(n24531), .B(n24532), .Z(n24530) );
  NAND U24949 ( .A(n24491), .B(n24493), .Z(n24496) );
  ANDN U24950 ( .B(B[4]), .A(n37), .Z(n24493) );
  XNOR U24951 ( .A(n24533), .B(n24534), .Z(n24491) );
  XNOR U24952 ( .A(n24535), .B(n24536), .Z(n24534) );
  ANDN U24953 ( .B(B[4]), .A(n36), .Z(n23194) );
  XNOR U24954 ( .A(n23202), .B(n24537), .Z(n23195) );
  XNOR U24955 ( .A(n23201), .B(n23199), .Z(n24537) );
  AND U24956 ( .A(n24538), .B(n24539), .Z(n23199) );
  NANDN U24957 ( .A(n24536), .B(n24540), .Z(n24539) );
  NANDN U24958 ( .A(n24535), .B(n24533), .Z(n24540) );
  AND U24959 ( .A(n24541), .B(n24542), .Z(n24536) );
  NANDN U24960 ( .A(n24532), .B(n24543), .Z(n24542) );
  OR U24961 ( .A(n24531), .B(n24529), .Z(n24543) );
  AND U24962 ( .A(n24544), .B(n24545), .Z(n24532) );
  NANDN U24963 ( .A(n24528), .B(n24546), .Z(n24545) );
  NANDN U24964 ( .A(n24527), .B(n24525), .Z(n24546) );
  AND U24965 ( .A(n24547), .B(n24548), .Z(n24528) );
  NANDN U24966 ( .A(n24524), .B(n24549), .Z(n24548) );
  OR U24967 ( .A(n24523), .B(n24521), .Z(n24549) );
  AND U24968 ( .A(n24550), .B(n24551), .Z(n24524) );
  NANDN U24969 ( .A(n24519), .B(n24552), .Z(n24551) );
  NAND U24970 ( .A(n24517), .B(n24520), .Z(n24552) );
  NANDN U24971 ( .A(n24515), .B(n24553), .Z(n24519) );
  AND U24972 ( .A(A[0]), .B(B[6]), .Z(n24553) );
  NAND U24973 ( .A(B[5]), .B(A[1]), .Z(n24515) );
  XNOR U24974 ( .A(n24554), .B(n24555), .Z(n24517) );
  NAND U24975 ( .A(A[0]), .B(B[7]), .Z(n24555) );
  NAND U24976 ( .A(A[2]), .B(B[5]), .Z(n24520) );
  NAND U24977 ( .A(n24521), .B(n24523), .Z(n24547) );
  ANDN U24978 ( .B(B[5]), .A(n41), .Z(n24523) );
  XOR U24979 ( .A(n24556), .B(n24557), .Z(n24521) );
  XNOR U24980 ( .A(n24558), .B(n24559), .Z(n24557) );
  NANDN U24981 ( .A(n24525), .B(n24527), .Z(n24544) );
  ANDN U24982 ( .B(B[5]), .A(n40), .Z(n24527) );
  XNOR U24983 ( .A(n24560), .B(n24561), .Z(n24525) );
  XNOR U24984 ( .A(n24562), .B(n24563), .Z(n24561) );
  NAND U24985 ( .A(n24529), .B(n24531), .Z(n24541) );
  ANDN U24986 ( .B(B[5]), .A(n39), .Z(n24531) );
  XNOR U24987 ( .A(n24564), .B(n24565), .Z(n24529) );
  XNOR U24988 ( .A(n24566), .B(n24567), .Z(n24565) );
  NANDN U24989 ( .A(n24533), .B(n24535), .Z(n24538) );
  ANDN U24990 ( .B(B[5]), .A(n38), .Z(n24535) );
  XNOR U24991 ( .A(n24568), .B(n24569), .Z(n24533) );
  XNOR U24992 ( .A(n24570), .B(n24571), .Z(n24569) );
  ANDN U24993 ( .B(B[5]), .A(n37), .Z(n23201) );
  XNOR U24994 ( .A(n23209), .B(n24572), .Z(n23202) );
  XNOR U24995 ( .A(n23208), .B(n23206), .Z(n24572) );
  AND U24996 ( .A(n24573), .B(n24574), .Z(n23206) );
  NANDN U24997 ( .A(n24571), .B(n24575), .Z(n24574) );
  OR U24998 ( .A(n24570), .B(n24568), .Z(n24575) );
  AND U24999 ( .A(n24576), .B(n24577), .Z(n24571) );
  NANDN U25000 ( .A(n24567), .B(n24578), .Z(n24577) );
  NANDN U25001 ( .A(n24566), .B(n24564), .Z(n24578) );
  AND U25002 ( .A(n24579), .B(n24580), .Z(n24567) );
  NANDN U25003 ( .A(n24563), .B(n24581), .Z(n24580) );
  OR U25004 ( .A(n24562), .B(n24560), .Z(n24581) );
  AND U25005 ( .A(n24582), .B(n24583), .Z(n24563) );
  NANDN U25006 ( .A(n24558), .B(n24584), .Z(n24583) );
  NAND U25007 ( .A(n24556), .B(n24559), .Z(n24584) );
  NANDN U25008 ( .A(n24554), .B(n24585), .Z(n24558) );
  AND U25009 ( .A(A[0]), .B(B[7]), .Z(n24585) );
  NAND U25010 ( .A(B[6]), .B(A[1]), .Z(n24554) );
  XNOR U25011 ( .A(n24586), .B(n24587), .Z(n24556) );
  NAND U25012 ( .A(A[0]), .B(B[8]), .Z(n24587) );
  NAND U25013 ( .A(A[2]), .B(B[6]), .Z(n24559) );
  NAND U25014 ( .A(n24560), .B(n24562), .Z(n24579) );
  ANDN U25015 ( .B(B[6]), .A(n41), .Z(n24562) );
  XOR U25016 ( .A(n24588), .B(n24589), .Z(n24560) );
  XNOR U25017 ( .A(n24590), .B(n24591), .Z(n24589) );
  NANDN U25018 ( .A(n24564), .B(n24566), .Z(n24576) );
  ANDN U25019 ( .B(B[6]), .A(n40), .Z(n24566) );
  XNOR U25020 ( .A(n24592), .B(n24593), .Z(n24564) );
  XNOR U25021 ( .A(n24594), .B(n24595), .Z(n24593) );
  NAND U25022 ( .A(n24568), .B(n24570), .Z(n24573) );
  ANDN U25023 ( .B(B[6]), .A(n39), .Z(n24570) );
  XNOR U25024 ( .A(n24596), .B(n24597), .Z(n24568) );
  XNOR U25025 ( .A(n24598), .B(n24599), .Z(n24597) );
  ANDN U25026 ( .B(B[6]), .A(n38), .Z(n23208) );
  XNOR U25027 ( .A(n23216), .B(n24600), .Z(n23209) );
  XNOR U25028 ( .A(n23215), .B(n23213), .Z(n24600) );
  AND U25029 ( .A(n24601), .B(n24602), .Z(n23213) );
  NANDN U25030 ( .A(n24599), .B(n24603), .Z(n24602) );
  NANDN U25031 ( .A(n24598), .B(n24596), .Z(n24603) );
  AND U25032 ( .A(n24604), .B(n24605), .Z(n24599) );
  NANDN U25033 ( .A(n24595), .B(n24606), .Z(n24605) );
  OR U25034 ( .A(n24594), .B(n24592), .Z(n24606) );
  AND U25035 ( .A(n24607), .B(n24608), .Z(n24595) );
  NANDN U25036 ( .A(n24590), .B(n24609), .Z(n24608) );
  NAND U25037 ( .A(n24588), .B(n24591), .Z(n24609) );
  NANDN U25038 ( .A(n24586), .B(n24610), .Z(n24590) );
  AND U25039 ( .A(A[0]), .B(B[8]), .Z(n24610) );
  NAND U25040 ( .A(B[7]), .B(A[1]), .Z(n24586) );
  XNOR U25041 ( .A(n24611), .B(n24612), .Z(n24588) );
  NAND U25042 ( .A(A[0]), .B(B[9]), .Z(n24612) );
  NAND U25043 ( .A(A[2]), .B(B[7]), .Z(n24591) );
  NAND U25044 ( .A(n24592), .B(n24594), .Z(n24604) );
  ANDN U25045 ( .B(B[7]), .A(n41), .Z(n24594) );
  XOR U25046 ( .A(n24613), .B(n24614), .Z(n24592) );
  XNOR U25047 ( .A(n24615), .B(n24616), .Z(n24614) );
  NANDN U25048 ( .A(n24596), .B(n24598), .Z(n24601) );
  ANDN U25049 ( .B(B[7]), .A(n40), .Z(n24598) );
  XNOR U25050 ( .A(n24617), .B(n24618), .Z(n24596) );
  XNOR U25051 ( .A(n24619), .B(n24620), .Z(n24618) );
  ANDN U25052 ( .B(B[7]), .A(n39), .Z(n23215) );
  XNOR U25053 ( .A(n23223), .B(n24621), .Z(n23216) );
  XNOR U25054 ( .A(n23222), .B(n23220), .Z(n24621) );
  AND U25055 ( .A(n24622), .B(n24623), .Z(n23220) );
  NANDN U25056 ( .A(n24620), .B(n24624), .Z(n24623) );
  OR U25057 ( .A(n24619), .B(n24617), .Z(n24624) );
  AND U25058 ( .A(n24625), .B(n24626), .Z(n24620) );
  NANDN U25059 ( .A(n24615), .B(n24627), .Z(n24626) );
  NAND U25060 ( .A(n24613), .B(n24616), .Z(n24627) );
  NANDN U25061 ( .A(n24611), .B(n24628), .Z(n24615) );
  AND U25062 ( .A(A[0]), .B(B[9]), .Z(n24628) );
  NAND U25063 ( .A(B[8]), .B(A[1]), .Z(n24611) );
  XNOR U25064 ( .A(n24629), .B(n24630), .Z(n24613) );
  NAND U25065 ( .A(A[0]), .B(B[10]), .Z(n24630) );
  NAND U25066 ( .A(A[2]), .B(B[8]), .Z(n24616) );
  NAND U25067 ( .A(n24617), .B(n24619), .Z(n24622) );
  ANDN U25068 ( .B(B[8]), .A(n41), .Z(n24619) );
  XOR U25069 ( .A(n24631), .B(n24632), .Z(n24617) );
  XNOR U25070 ( .A(n24633), .B(n24634), .Z(n24632) );
  ANDN U25071 ( .B(B[8]), .A(n40), .Z(n23222) );
  XNOR U25072 ( .A(n23230), .B(n24635), .Z(n23223) );
  XNOR U25073 ( .A(n23229), .B(n23227), .Z(n24635) );
  AND U25074 ( .A(n24636), .B(n24637), .Z(n23227) );
  NANDN U25075 ( .A(n24633), .B(n24638), .Z(n24637) );
  NAND U25076 ( .A(n24631), .B(n24634), .Z(n24638) );
  NANDN U25077 ( .A(n24629), .B(n24639), .Z(n24633) );
  AND U25078 ( .A(A[0]), .B(B[10]), .Z(n24639) );
  NAND U25079 ( .A(B[9]), .B(A[1]), .Z(n24629) );
  XNOR U25080 ( .A(n24640), .B(n24641), .Z(n24631) );
  NAND U25081 ( .A(A[0]), .B(B[11]), .Z(n24641) );
  NAND U25082 ( .A(A[2]), .B(B[9]), .Z(n24634) );
  ANDN U25083 ( .B(B[9]), .A(n41), .Z(n23229) );
  XOR U25084 ( .A(n23236), .B(n24642), .Z(n23230) );
  XNOR U25085 ( .A(n23234), .B(n23237), .Z(n24642) );
  NAND U25086 ( .A(A[2]), .B(B[10]), .Z(n23237) );
  NANDN U25087 ( .A(n24640), .B(n24643), .Z(n23234) );
  AND U25088 ( .A(A[0]), .B(B[11]), .Z(n24643) );
  NAND U25089 ( .A(B[10]), .B(A[1]), .Z(n24640) );
  XNOR U25090 ( .A(n23239), .B(n24644), .Z(n23236) );
  NAND U25091 ( .A(A[0]), .B(B[12]), .Z(n24644) );
  NAND U25092 ( .A(B[11]), .B(A[1]), .Z(n23239) );
  XOR U25093 ( .A(n533), .B(n532), .Z(\A1[109] ) );
  XOR U25094 ( .A(n24251), .B(n24645), .Z(n532) );
  XNOR U25095 ( .A(n24250), .B(n24248), .Z(n24645) );
  AND U25096 ( .A(n24646), .B(n24647), .Z(n24248) );
  NANDN U25097 ( .A(n24648), .B(n24649), .Z(n24647) );
  NANDN U25098 ( .A(n24650), .B(n24651), .Z(n24649) );
  NANDN U25099 ( .A(n24651), .B(n24650), .Z(n24646) );
  ANDN U25100 ( .B(B[96]), .A(n29), .Z(n24250) );
  XNOR U25101 ( .A(n24157), .B(n24652), .Z(n24251) );
  XNOR U25102 ( .A(n24156), .B(n24154), .Z(n24652) );
  AND U25103 ( .A(n24653), .B(n24654), .Z(n24154) );
  NANDN U25104 ( .A(n24655), .B(n24656), .Z(n24654) );
  OR U25105 ( .A(n24657), .B(n24658), .Z(n24656) );
  NAND U25106 ( .A(n24658), .B(n24657), .Z(n24653) );
  ANDN U25107 ( .B(B[97]), .A(n30), .Z(n24156) );
  XNOR U25108 ( .A(n24164), .B(n24659), .Z(n24157) );
  XNOR U25109 ( .A(n24163), .B(n24161), .Z(n24659) );
  AND U25110 ( .A(n24660), .B(n24661), .Z(n24161) );
  NANDN U25111 ( .A(n24662), .B(n24663), .Z(n24661) );
  NANDN U25112 ( .A(n24664), .B(n24665), .Z(n24663) );
  NANDN U25113 ( .A(n24665), .B(n24664), .Z(n24660) );
  ANDN U25114 ( .B(B[98]), .A(n31), .Z(n24163) );
  XNOR U25115 ( .A(n24171), .B(n24666), .Z(n24164) );
  XNOR U25116 ( .A(n24170), .B(n24168), .Z(n24666) );
  AND U25117 ( .A(n24667), .B(n24668), .Z(n24168) );
  NANDN U25118 ( .A(n24669), .B(n24670), .Z(n24668) );
  OR U25119 ( .A(n24671), .B(n24672), .Z(n24670) );
  NAND U25120 ( .A(n24672), .B(n24671), .Z(n24667) );
  ANDN U25121 ( .B(A[12]), .A(n5), .Z(n24170) );
  XNOR U25122 ( .A(n24178), .B(n24673), .Z(n24171) );
  XNOR U25123 ( .A(n24177), .B(n24175), .Z(n24673) );
  AND U25124 ( .A(n24674), .B(n24675), .Z(n24175) );
  NANDN U25125 ( .A(n24676), .B(n24677), .Z(n24675) );
  NANDN U25126 ( .A(n24678), .B(n24679), .Z(n24677) );
  NANDN U25127 ( .A(n24679), .B(n24678), .Z(n24674) );
  ANDN U25128 ( .B(A[11]), .A(n3), .Z(n24177) );
  XNOR U25129 ( .A(n24185), .B(n24680), .Z(n24178) );
  XNOR U25130 ( .A(n24184), .B(n24182), .Z(n24680) );
  AND U25131 ( .A(n24681), .B(n24682), .Z(n24182) );
  NANDN U25132 ( .A(n24683), .B(n24684), .Z(n24682) );
  OR U25133 ( .A(n24685), .B(n24686), .Z(n24684) );
  NAND U25134 ( .A(n24686), .B(n24685), .Z(n24681) );
  ANDN U25135 ( .B(B[101]), .A(n34), .Z(n24184) );
  XNOR U25136 ( .A(n24192), .B(n24687), .Z(n24185) );
  XNOR U25137 ( .A(n24191), .B(n24189), .Z(n24687) );
  AND U25138 ( .A(n24688), .B(n24689), .Z(n24189) );
  NANDN U25139 ( .A(n24690), .B(n24691), .Z(n24689) );
  NANDN U25140 ( .A(n24692), .B(n24693), .Z(n24691) );
  NANDN U25141 ( .A(n24693), .B(n24692), .Z(n24688) );
  ANDN U25142 ( .B(B[102]), .A(n35), .Z(n24191) );
  XNOR U25143 ( .A(n24199), .B(n24694), .Z(n24192) );
  XNOR U25144 ( .A(n24198), .B(n24196), .Z(n24694) );
  AND U25145 ( .A(n24695), .B(n24696), .Z(n24196) );
  NANDN U25146 ( .A(n24697), .B(n24698), .Z(n24696) );
  OR U25147 ( .A(n24699), .B(n24700), .Z(n24698) );
  NAND U25148 ( .A(n24700), .B(n24699), .Z(n24695) );
  ANDN U25149 ( .B(B[103]), .A(n36), .Z(n24198) );
  XNOR U25150 ( .A(n24206), .B(n24701), .Z(n24199) );
  XNOR U25151 ( .A(n24205), .B(n24203), .Z(n24701) );
  AND U25152 ( .A(n24702), .B(n24703), .Z(n24203) );
  NANDN U25153 ( .A(n24704), .B(n24705), .Z(n24703) );
  NANDN U25154 ( .A(n24706), .B(n24707), .Z(n24705) );
  NANDN U25155 ( .A(n24707), .B(n24706), .Z(n24702) );
  ANDN U25156 ( .B(B[104]), .A(n37), .Z(n24205) );
  XNOR U25157 ( .A(n24213), .B(n24708), .Z(n24206) );
  XNOR U25158 ( .A(n24212), .B(n24210), .Z(n24708) );
  AND U25159 ( .A(n24709), .B(n24710), .Z(n24210) );
  NANDN U25160 ( .A(n24711), .B(n24712), .Z(n24710) );
  OR U25161 ( .A(n24713), .B(n24714), .Z(n24712) );
  NAND U25162 ( .A(n24714), .B(n24713), .Z(n24709) );
  ANDN U25163 ( .B(B[105]), .A(n38), .Z(n24212) );
  XNOR U25164 ( .A(n24220), .B(n24715), .Z(n24213) );
  XNOR U25165 ( .A(n24219), .B(n24217), .Z(n24715) );
  AND U25166 ( .A(n24716), .B(n24717), .Z(n24217) );
  NANDN U25167 ( .A(n24718), .B(n24719), .Z(n24717) );
  NANDN U25168 ( .A(n24720), .B(n24721), .Z(n24719) );
  NANDN U25169 ( .A(n24721), .B(n24720), .Z(n24716) );
  ANDN U25170 ( .B(B[106]), .A(n39), .Z(n24219) );
  XNOR U25171 ( .A(n24227), .B(n24722), .Z(n24220) );
  XNOR U25172 ( .A(n24226), .B(n24224), .Z(n24722) );
  AND U25173 ( .A(n24723), .B(n24724), .Z(n24224) );
  NANDN U25174 ( .A(n24725), .B(n24726), .Z(n24724) );
  OR U25175 ( .A(n24727), .B(n24728), .Z(n24726) );
  NAND U25176 ( .A(n24728), .B(n24727), .Z(n24723) );
  ANDN U25177 ( .B(B[107]), .A(n40), .Z(n24226) );
  XNOR U25178 ( .A(n24234), .B(n24729), .Z(n24227) );
  XNOR U25179 ( .A(n24233), .B(n24231), .Z(n24729) );
  AND U25180 ( .A(n24730), .B(n24731), .Z(n24231) );
  NANDN U25181 ( .A(n24732), .B(n24733), .Z(n24731) );
  NAND U25182 ( .A(n24734), .B(n24735), .Z(n24733) );
  ANDN U25183 ( .B(B[108]), .A(n41), .Z(n24233) );
  XOR U25184 ( .A(n24240), .B(n24736), .Z(n24234) );
  XNOR U25185 ( .A(n24238), .B(n24241), .Z(n24736) );
  NAND U25186 ( .A(A[2]), .B(B[109]), .Z(n24241) );
  NANDN U25187 ( .A(n24737), .B(n24738), .Z(n24238) );
  AND U25188 ( .A(A[0]), .B(B[110]), .Z(n24738) );
  XNOR U25189 ( .A(n24243), .B(n24739), .Z(n24240) );
  NAND U25190 ( .A(A[0]), .B(B[111]), .Z(n24739) );
  NAND U25191 ( .A(B[110]), .B(A[1]), .Z(n24243) );
  NAND U25192 ( .A(n24740), .B(n24741), .Z(n533) );
  NANDN U25193 ( .A(n24742), .B(n24743), .Z(n24741) );
  OR U25194 ( .A(n24744), .B(n24745), .Z(n24743) );
  NAND U25195 ( .A(n24745), .B(n24744), .Z(n24740) );
  XOR U25196 ( .A(n535), .B(n534), .Z(\A1[108] ) );
  XOR U25197 ( .A(n24745), .B(n24746), .Z(n534) );
  XNOR U25198 ( .A(n24744), .B(n24742), .Z(n24746) );
  AND U25199 ( .A(n24747), .B(n24748), .Z(n24742) );
  NANDN U25200 ( .A(n24749), .B(n24750), .Z(n24748) );
  NANDN U25201 ( .A(n24751), .B(n24752), .Z(n24750) );
  NANDN U25202 ( .A(n24752), .B(n24751), .Z(n24747) );
  ANDN U25203 ( .B(B[95]), .A(n29), .Z(n24744) );
  XNOR U25204 ( .A(n24651), .B(n24753), .Z(n24745) );
  XNOR U25205 ( .A(n24650), .B(n24648), .Z(n24753) );
  AND U25206 ( .A(n24754), .B(n24755), .Z(n24648) );
  NANDN U25207 ( .A(n24756), .B(n24757), .Z(n24755) );
  OR U25208 ( .A(n24758), .B(n24759), .Z(n24757) );
  NAND U25209 ( .A(n24759), .B(n24758), .Z(n24754) );
  ANDN U25210 ( .B(B[96]), .A(n30), .Z(n24650) );
  XNOR U25211 ( .A(n24658), .B(n24760), .Z(n24651) );
  XNOR U25212 ( .A(n24657), .B(n24655), .Z(n24760) );
  AND U25213 ( .A(n24761), .B(n24762), .Z(n24655) );
  NANDN U25214 ( .A(n24763), .B(n24764), .Z(n24762) );
  NANDN U25215 ( .A(n24765), .B(n24766), .Z(n24764) );
  NANDN U25216 ( .A(n24766), .B(n24765), .Z(n24761) );
  ANDN U25217 ( .B(A[13]), .A(n8), .Z(n24657) );
  XNOR U25218 ( .A(n24665), .B(n24767), .Z(n24658) );
  XNOR U25219 ( .A(n24664), .B(n24662), .Z(n24767) );
  AND U25220 ( .A(n24768), .B(n24769), .Z(n24662) );
  NANDN U25221 ( .A(n24770), .B(n24771), .Z(n24769) );
  OR U25222 ( .A(n24772), .B(n24773), .Z(n24771) );
  NAND U25223 ( .A(n24773), .B(n24772), .Z(n24768) );
  ANDN U25224 ( .B(B[98]), .A(n32), .Z(n24664) );
  XNOR U25225 ( .A(n24672), .B(n24774), .Z(n24665) );
  XNOR U25226 ( .A(n24671), .B(n24669), .Z(n24774) );
  AND U25227 ( .A(n24775), .B(n24776), .Z(n24669) );
  NANDN U25228 ( .A(n24777), .B(n24778), .Z(n24776) );
  NANDN U25229 ( .A(n24779), .B(n24780), .Z(n24778) );
  NANDN U25230 ( .A(n24780), .B(n24779), .Z(n24775) );
  ANDN U25231 ( .B(A[11]), .A(n5), .Z(n24671) );
  XNOR U25232 ( .A(n24679), .B(n24781), .Z(n24672) );
  XNOR U25233 ( .A(n24678), .B(n24676), .Z(n24781) );
  AND U25234 ( .A(n24782), .B(n24783), .Z(n24676) );
  NANDN U25235 ( .A(n24784), .B(n24785), .Z(n24783) );
  OR U25236 ( .A(n24786), .B(n24787), .Z(n24785) );
  NAND U25237 ( .A(n24787), .B(n24786), .Z(n24782) );
  ANDN U25238 ( .B(A[10]), .A(n3), .Z(n24678) );
  XNOR U25239 ( .A(n24686), .B(n24788), .Z(n24679) );
  XNOR U25240 ( .A(n24685), .B(n24683), .Z(n24788) );
  AND U25241 ( .A(n24789), .B(n24790), .Z(n24683) );
  NANDN U25242 ( .A(n24791), .B(n24792), .Z(n24790) );
  NANDN U25243 ( .A(n24793), .B(n24794), .Z(n24792) );
  NANDN U25244 ( .A(n24794), .B(n24793), .Z(n24789) );
  ANDN U25245 ( .B(B[101]), .A(n35), .Z(n24685) );
  XNOR U25246 ( .A(n24693), .B(n24795), .Z(n24686) );
  XNOR U25247 ( .A(n24692), .B(n24690), .Z(n24795) );
  AND U25248 ( .A(n24796), .B(n24797), .Z(n24690) );
  NANDN U25249 ( .A(n24798), .B(n24799), .Z(n24797) );
  OR U25250 ( .A(n24800), .B(n24801), .Z(n24799) );
  NAND U25251 ( .A(n24801), .B(n24800), .Z(n24796) );
  ANDN U25252 ( .B(B[102]), .A(n36), .Z(n24692) );
  XNOR U25253 ( .A(n24700), .B(n24802), .Z(n24693) );
  XNOR U25254 ( .A(n24699), .B(n24697), .Z(n24802) );
  AND U25255 ( .A(n24803), .B(n24804), .Z(n24697) );
  NANDN U25256 ( .A(n24805), .B(n24806), .Z(n24804) );
  NANDN U25257 ( .A(n24807), .B(n24808), .Z(n24806) );
  NANDN U25258 ( .A(n24808), .B(n24807), .Z(n24803) );
  ANDN U25259 ( .B(B[103]), .A(n37), .Z(n24699) );
  XNOR U25260 ( .A(n24707), .B(n24809), .Z(n24700) );
  XNOR U25261 ( .A(n24706), .B(n24704), .Z(n24809) );
  AND U25262 ( .A(n24810), .B(n24811), .Z(n24704) );
  NANDN U25263 ( .A(n24812), .B(n24813), .Z(n24811) );
  OR U25264 ( .A(n24814), .B(n24815), .Z(n24813) );
  NAND U25265 ( .A(n24815), .B(n24814), .Z(n24810) );
  ANDN U25266 ( .B(B[104]), .A(n38), .Z(n24706) );
  XNOR U25267 ( .A(n24714), .B(n24816), .Z(n24707) );
  XNOR U25268 ( .A(n24713), .B(n24711), .Z(n24816) );
  AND U25269 ( .A(n24817), .B(n24818), .Z(n24711) );
  NANDN U25270 ( .A(n24819), .B(n24820), .Z(n24818) );
  NANDN U25271 ( .A(n24821), .B(n24822), .Z(n24820) );
  NANDN U25272 ( .A(n24822), .B(n24821), .Z(n24817) );
  ANDN U25273 ( .B(B[105]), .A(n39), .Z(n24713) );
  XNOR U25274 ( .A(n24721), .B(n24823), .Z(n24714) );
  XNOR U25275 ( .A(n24720), .B(n24718), .Z(n24823) );
  AND U25276 ( .A(n24824), .B(n24825), .Z(n24718) );
  NANDN U25277 ( .A(n24826), .B(n24827), .Z(n24825) );
  OR U25278 ( .A(n24828), .B(n24829), .Z(n24827) );
  NAND U25279 ( .A(n24829), .B(n24828), .Z(n24824) );
  ANDN U25280 ( .B(B[106]), .A(n40), .Z(n24720) );
  XNOR U25281 ( .A(n24728), .B(n24830), .Z(n24721) );
  XNOR U25282 ( .A(n24727), .B(n24725), .Z(n24830) );
  AND U25283 ( .A(n24831), .B(n24832), .Z(n24725) );
  NANDN U25284 ( .A(n24833), .B(n24834), .Z(n24832) );
  NAND U25285 ( .A(n24835), .B(n24836), .Z(n24834) );
  ANDN U25286 ( .B(B[107]), .A(n41), .Z(n24727) );
  XOR U25287 ( .A(n24734), .B(n24837), .Z(n24728) );
  XNOR U25288 ( .A(n24732), .B(n24735), .Z(n24837) );
  NAND U25289 ( .A(A[2]), .B(B[108]), .Z(n24735) );
  NANDN U25290 ( .A(n24838), .B(n24839), .Z(n24732) );
  AND U25291 ( .A(A[0]), .B(B[109]), .Z(n24839) );
  XNOR U25292 ( .A(n24737), .B(n24840), .Z(n24734) );
  NAND U25293 ( .A(A[0]), .B(B[110]), .Z(n24840) );
  NAND U25294 ( .A(B[109]), .B(A[1]), .Z(n24737) );
  NAND U25295 ( .A(n24841), .B(n24842), .Z(n535) );
  NANDN U25296 ( .A(n24843), .B(n24844), .Z(n24842) );
  OR U25297 ( .A(n24845), .B(n24846), .Z(n24844) );
  NAND U25298 ( .A(n24846), .B(n24845), .Z(n24841) );
  XOR U25299 ( .A(n537), .B(n536), .Z(\A1[107] ) );
  XOR U25300 ( .A(n24846), .B(n24847), .Z(n536) );
  XNOR U25301 ( .A(n24845), .B(n24843), .Z(n24847) );
  AND U25302 ( .A(n24848), .B(n24849), .Z(n24843) );
  NANDN U25303 ( .A(n24850), .B(n24851), .Z(n24849) );
  NANDN U25304 ( .A(n24852), .B(n24853), .Z(n24851) );
  NANDN U25305 ( .A(n24853), .B(n24852), .Z(n24848) );
  ANDN U25306 ( .B(B[94]), .A(n29), .Z(n24845) );
  XNOR U25307 ( .A(n24752), .B(n24854), .Z(n24846) );
  XNOR U25308 ( .A(n24751), .B(n24749), .Z(n24854) );
  AND U25309 ( .A(n24855), .B(n24856), .Z(n24749) );
  NANDN U25310 ( .A(n24857), .B(n24858), .Z(n24856) );
  OR U25311 ( .A(n24859), .B(n24860), .Z(n24858) );
  NAND U25312 ( .A(n24860), .B(n24859), .Z(n24855) );
  ANDN U25313 ( .B(B[95]), .A(n30), .Z(n24751) );
  XNOR U25314 ( .A(n24759), .B(n24861), .Z(n24752) );
  XNOR U25315 ( .A(n24758), .B(n24756), .Z(n24861) );
  AND U25316 ( .A(n24862), .B(n24863), .Z(n24756) );
  NANDN U25317 ( .A(n24864), .B(n24865), .Z(n24863) );
  NANDN U25318 ( .A(n24866), .B(n24867), .Z(n24865) );
  NANDN U25319 ( .A(n24867), .B(n24866), .Z(n24862) );
  ANDN U25320 ( .B(B[96]), .A(n31), .Z(n24758) );
  XNOR U25321 ( .A(n24766), .B(n24868), .Z(n24759) );
  XNOR U25322 ( .A(n24765), .B(n24763), .Z(n24868) );
  AND U25323 ( .A(n24869), .B(n24870), .Z(n24763) );
  NANDN U25324 ( .A(n24871), .B(n24872), .Z(n24870) );
  OR U25325 ( .A(n24873), .B(n24874), .Z(n24872) );
  NAND U25326 ( .A(n24874), .B(n24873), .Z(n24869) );
  ANDN U25327 ( .B(A[12]), .A(n8), .Z(n24765) );
  XNOR U25328 ( .A(n24773), .B(n24875), .Z(n24766) );
  XNOR U25329 ( .A(n24772), .B(n24770), .Z(n24875) );
  AND U25330 ( .A(n24876), .B(n24877), .Z(n24770) );
  NANDN U25331 ( .A(n24878), .B(n24879), .Z(n24877) );
  NANDN U25332 ( .A(n24880), .B(n24881), .Z(n24879) );
  NANDN U25333 ( .A(n24881), .B(n24880), .Z(n24876) );
  ANDN U25334 ( .B(B[98]), .A(n33), .Z(n24772) );
  XNOR U25335 ( .A(n24780), .B(n24882), .Z(n24773) );
  XNOR U25336 ( .A(n24779), .B(n24777), .Z(n24882) );
  AND U25337 ( .A(n24883), .B(n24884), .Z(n24777) );
  NANDN U25338 ( .A(n24885), .B(n24886), .Z(n24884) );
  OR U25339 ( .A(n24887), .B(n24888), .Z(n24886) );
  NAND U25340 ( .A(n24888), .B(n24887), .Z(n24883) );
  ANDN U25341 ( .B(A[10]), .A(n5), .Z(n24779) );
  XNOR U25342 ( .A(n24787), .B(n24889), .Z(n24780) );
  XNOR U25343 ( .A(n24786), .B(n24784), .Z(n24889) );
  AND U25344 ( .A(n24890), .B(n24891), .Z(n24784) );
  NANDN U25345 ( .A(n24892), .B(n24893), .Z(n24891) );
  NANDN U25346 ( .A(n24894), .B(n24895), .Z(n24893) );
  NANDN U25347 ( .A(n24895), .B(n24894), .Z(n24890) );
  ANDN U25348 ( .B(A[9]), .A(n3), .Z(n24786) );
  XNOR U25349 ( .A(n24794), .B(n24896), .Z(n24787) );
  XNOR U25350 ( .A(n24793), .B(n24791), .Z(n24896) );
  AND U25351 ( .A(n24897), .B(n24898), .Z(n24791) );
  NANDN U25352 ( .A(n24899), .B(n24900), .Z(n24898) );
  OR U25353 ( .A(n24901), .B(n24902), .Z(n24900) );
  NAND U25354 ( .A(n24902), .B(n24901), .Z(n24897) );
  ANDN U25355 ( .B(B[101]), .A(n36), .Z(n24793) );
  XNOR U25356 ( .A(n24801), .B(n24903), .Z(n24794) );
  XNOR U25357 ( .A(n24800), .B(n24798), .Z(n24903) );
  AND U25358 ( .A(n24904), .B(n24905), .Z(n24798) );
  NANDN U25359 ( .A(n24906), .B(n24907), .Z(n24905) );
  NANDN U25360 ( .A(n24908), .B(n24909), .Z(n24907) );
  NANDN U25361 ( .A(n24909), .B(n24908), .Z(n24904) );
  ANDN U25362 ( .B(B[102]), .A(n37), .Z(n24800) );
  XNOR U25363 ( .A(n24808), .B(n24910), .Z(n24801) );
  XNOR U25364 ( .A(n24807), .B(n24805), .Z(n24910) );
  AND U25365 ( .A(n24911), .B(n24912), .Z(n24805) );
  NANDN U25366 ( .A(n24913), .B(n24914), .Z(n24912) );
  OR U25367 ( .A(n24915), .B(n24916), .Z(n24914) );
  NAND U25368 ( .A(n24916), .B(n24915), .Z(n24911) );
  ANDN U25369 ( .B(B[103]), .A(n38), .Z(n24807) );
  XNOR U25370 ( .A(n24815), .B(n24917), .Z(n24808) );
  XNOR U25371 ( .A(n24814), .B(n24812), .Z(n24917) );
  AND U25372 ( .A(n24918), .B(n24919), .Z(n24812) );
  NANDN U25373 ( .A(n24920), .B(n24921), .Z(n24919) );
  NANDN U25374 ( .A(n24922), .B(n24923), .Z(n24921) );
  NANDN U25375 ( .A(n24923), .B(n24922), .Z(n24918) );
  ANDN U25376 ( .B(B[104]), .A(n39), .Z(n24814) );
  XNOR U25377 ( .A(n24822), .B(n24924), .Z(n24815) );
  XNOR U25378 ( .A(n24821), .B(n24819), .Z(n24924) );
  AND U25379 ( .A(n24925), .B(n24926), .Z(n24819) );
  NANDN U25380 ( .A(n24927), .B(n24928), .Z(n24926) );
  OR U25381 ( .A(n24929), .B(n24930), .Z(n24928) );
  NAND U25382 ( .A(n24930), .B(n24929), .Z(n24925) );
  ANDN U25383 ( .B(B[105]), .A(n40), .Z(n24821) );
  XNOR U25384 ( .A(n24829), .B(n24931), .Z(n24822) );
  XNOR U25385 ( .A(n24828), .B(n24826), .Z(n24931) );
  AND U25386 ( .A(n24932), .B(n24933), .Z(n24826) );
  NANDN U25387 ( .A(n24934), .B(n24935), .Z(n24933) );
  NAND U25388 ( .A(n24936), .B(n24937), .Z(n24935) );
  ANDN U25389 ( .B(B[106]), .A(n41), .Z(n24828) );
  XOR U25390 ( .A(n24835), .B(n24938), .Z(n24829) );
  XNOR U25391 ( .A(n24833), .B(n24836), .Z(n24938) );
  NAND U25392 ( .A(A[2]), .B(B[107]), .Z(n24836) );
  NANDN U25393 ( .A(n24939), .B(n24940), .Z(n24833) );
  AND U25394 ( .A(A[0]), .B(B[108]), .Z(n24940) );
  XNOR U25395 ( .A(n24838), .B(n24941), .Z(n24835) );
  NAND U25396 ( .A(A[0]), .B(B[109]), .Z(n24941) );
  NAND U25397 ( .A(B[108]), .B(A[1]), .Z(n24838) );
  NAND U25398 ( .A(n24942), .B(n24943), .Z(n537) );
  NANDN U25399 ( .A(n24944), .B(n24945), .Z(n24943) );
  OR U25400 ( .A(n24946), .B(n24947), .Z(n24945) );
  NAND U25401 ( .A(n24947), .B(n24946), .Z(n24942) );
  XOR U25402 ( .A(n539), .B(n538), .Z(\A1[106] ) );
  XOR U25403 ( .A(n24947), .B(n24948), .Z(n538) );
  XNOR U25404 ( .A(n24946), .B(n24944), .Z(n24948) );
  AND U25405 ( .A(n24949), .B(n24950), .Z(n24944) );
  NANDN U25406 ( .A(n24951), .B(n24952), .Z(n24950) );
  NANDN U25407 ( .A(n24953), .B(n24954), .Z(n24952) );
  NANDN U25408 ( .A(n24954), .B(n24953), .Z(n24949) );
  ANDN U25409 ( .B(B[93]), .A(n29), .Z(n24946) );
  XNOR U25410 ( .A(n24853), .B(n24955), .Z(n24947) );
  XNOR U25411 ( .A(n24852), .B(n24850), .Z(n24955) );
  AND U25412 ( .A(n24956), .B(n24957), .Z(n24850) );
  NANDN U25413 ( .A(n24958), .B(n24959), .Z(n24957) );
  OR U25414 ( .A(n24960), .B(n24961), .Z(n24959) );
  NAND U25415 ( .A(n24961), .B(n24960), .Z(n24956) );
  ANDN U25416 ( .B(B[94]), .A(n30), .Z(n24852) );
  XNOR U25417 ( .A(n24860), .B(n24962), .Z(n24853) );
  XNOR U25418 ( .A(n24859), .B(n24857), .Z(n24962) );
  AND U25419 ( .A(n24963), .B(n24964), .Z(n24857) );
  NANDN U25420 ( .A(n24965), .B(n24966), .Z(n24964) );
  NANDN U25421 ( .A(n24967), .B(n24968), .Z(n24966) );
  NANDN U25422 ( .A(n24968), .B(n24967), .Z(n24963) );
  ANDN U25423 ( .B(B[95]), .A(n31), .Z(n24859) );
  XNOR U25424 ( .A(n24867), .B(n24969), .Z(n24860) );
  XNOR U25425 ( .A(n24866), .B(n24864), .Z(n24969) );
  AND U25426 ( .A(n24970), .B(n24971), .Z(n24864) );
  NANDN U25427 ( .A(n24972), .B(n24973), .Z(n24971) );
  OR U25428 ( .A(n24974), .B(n24975), .Z(n24973) );
  NAND U25429 ( .A(n24975), .B(n24974), .Z(n24970) );
  ANDN U25430 ( .B(A[12]), .A(n10), .Z(n24866) );
  XNOR U25431 ( .A(n24874), .B(n24976), .Z(n24867) );
  XNOR U25432 ( .A(n24873), .B(n24871), .Z(n24976) );
  AND U25433 ( .A(n24977), .B(n24978), .Z(n24871) );
  NANDN U25434 ( .A(n24979), .B(n24980), .Z(n24978) );
  NANDN U25435 ( .A(n24981), .B(n24982), .Z(n24980) );
  NANDN U25436 ( .A(n24982), .B(n24981), .Z(n24977) );
  ANDN U25437 ( .B(A[11]), .A(n8), .Z(n24873) );
  XNOR U25438 ( .A(n24881), .B(n24983), .Z(n24874) );
  XNOR U25439 ( .A(n24880), .B(n24878), .Z(n24983) );
  AND U25440 ( .A(n24984), .B(n24985), .Z(n24878) );
  NANDN U25441 ( .A(n24986), .B(n24987), .Z(n24985) );
  OR U25442 ( .A(n24988), .B(n24989), .Z(n24987) );
  NAND U25443 ( .A(n24989), .B(n24988), .Z(n24984) );
  ANDN U25444 ( .B(B[98]), .A(n34), .Z(n24880) );
  XNOR U25445 ( .A(n24888), .B(n24990), .Z(n24881) );
  XNOR U25446 ( .A(n24887), .B(n24885), .Z(n24990) );
  AND U25447 ( .A(n24991), .B(n24992), .Z(n24885) );
  NANDN U25448 ( .A(n24993), .B(n24994), .Z(n24992) );
  NANDN U25449 ( .A(n24995), .B(n24996), .Z(n24994) );
  NANDN U25450 ( .A(n24996), .B(n24995), .Z(n24991) );
  ANDN U25451 ( .B(A[9]), .A(n5), .Z(n24887) );
  XNOR U25452 ( .A(n24895), .B(n24997), .Z(n24888) );
  XNOR U25453 ( .A(n24894), .B(n24892), .Z(n24997) );
  AND U25454 ( .A(n24998), .B(n24999), .Z(n24892) );
  NANDN U25455 ( .A(n25000), .B(n25001), .Z(n24999) );
  OR U25456 ( .A(n25002), .B(n25003), .Z(n25001) );
  NAND U25457 ( .A(n25003), .B(n25002), .Z(n24998) );
  ANDN U25458 ( .B(A[8]), .A(n3), .Z(n24894) );
  XNOR U25459 ( .A(n24902), .B(n25004), .Z(n24895) );
  XNOR U25460 ( .A(n24901), .B(n24899), .Z(n25004) );
  AND U25461 ( .A(n25005), .B(n25006), .Z(n24899) );
  NANDN U25462 ( .A(n25007), .B(n25008), .Z(n25006) );
  NANDN U25463 ( .A(n25009), .B(n25010), .Z(n25008) );
  NANDN U25464 ( .A(n25010), .B(n25009), .Z(n25005) );
  ANDN U25465 ( .B(B[101]), .A(n37), .Z(n24901) );
  XNOR U25466 ( .A(n24909), .B(n25011), .Z(n24902) );
  XNOR U25467 ( .A(n24908), .B(n24906), .Z(n25011) );
  AND U25468 ( .A(n25012), .B(n25013), .Z(n24906) );
  NANDN U25469 ( .A(n25014), .B(n25015), .Z(n25013) );
  OR U25470 ( .A(n25016), .B(n25017), .Z(n25015) );
  NAND U25471 ( .A(n25017), .B(n25016), .Z(n25012) );
  ANDN U25472 ( .B(B[102]), .A(n38), .Z(n24908) );
  XNOR U25473 ( .A(n24916), .B(n25018), .Z(n24909) );
  XNOR U25474 ( .A(n24915), .B(n24913), .Z(n25018) );
  AND U25475 ( .A(n25019), .B(n25020), .Z(n24913) );
  NANDN U25476 ( .A(n25021), .B(n25022), .Z(n25020) );
  NANDN U25477 ( .A(n25023), .B(n25024), .Z(n25022) );
  NANDN U25478 ( .A(n25024), .B(n25023), .Z(n25019) );
  ANDN U25479 ( .B(B[103]), .A(n39), .Z(n24915) );
  XNOR U25480 ( .A(n24923), .B(n25025), .Z(n24916) );
  XNOR U25481 ( .A(n24922), .B(n24920), .Z(n25025) );
  AND U25482 ( .A(n25026), .B(n25027), .Z(n24920) );
  NANDN U25483 ( .A(n25028), .B(n25029), .Z(n25027) );
  OR U25484 ( .A(n25030), .B(n25031), .Z(n25029) );
  NAND U25485 ( .A(n25031), .B(n25030), .Z(n25026) );
  ANDN U25486 ( .B(B[104]), .A(n40), .Z(n24922) );
  XNOR U25487 ( .A(n24930), .B(n25032), .Z(n24923) );
  XNOR U25488 ( .A(n24929), .B(n24927), .Z(n25032) );
  AND U25489 ( .A(n25033), .B(n25034), .Z(n24927) );
  NANDN U25490 ( .A(n25035), .B(n25036), .Z(n25034) );
  NAND U25491 ( .A(n25037), .B(n25038), .Z(n25036) );
  ANDN U25492 ( .B(B[105]), .A(n41), .Z(n24929) );
  XOR U25493 ( .A(n24936), .B(n25039), .Z(n24930) );
  XNOR U25494 ( .A(n24934), .B(n24937), .Z(n25039) );
  NAND U25495 ( .A(A[2]), .B(B[106]), .Z(n24937) );
  NANDN U25496 ( .A(n25040), .B(n25041), .Z(n24934) );
  AND U25497 ( .A(A[0]), .B(B[107]), .Z(n25041) );
  XNOR U25498 ( .A(n24939), .B(n25042), .Z(n24936) );
  NAND U25499 ( .A(A[0]), .B(B[108]), .Z(n25042) );
  NAND U25500 ( .A(B[107]), .B(A[1]), .Z(n24939) );
  NAND U25501 ( .A(n25043), .B(n25044), .Z(n539) );
  NANDN U25502 ( .A(n25045), .B(n25046), .Z(n25044) );
  OR U25503 ( .A(n25047), .B(n25048), .Z(n25046) );
  NAND U25504 ( .A(n25048), .B(n25047), .Z(n25043) );
  XOR U25505 ( .A(n541), .B(n540), .Z(\A1[105] ) );
  XOR U25506 ( .A(n25048), .B(n25049), .Z(n540) );
  XNOR U25507 ( .A(n25047), .B(n25045), .Z(n25049) );
  AND U25508 ( .A(n25050), .B(n25051), .Z(n25045) );
  NANDN U25509 ( .A(n25052), .B(n25053), .Z(n25051) );
  NANDN U25510 ( .A(n25054), .B(n25055), .Z(n25053) );
  NANDN U25511 ( .A(n25055), .B(n25054), .Z(n25050) );
  ANDN U25512 ( .B(B[92]), .A(n29), .Z(n25047) );
  XNOR U25513 ( .A(n24954), .B(n25056), .Z(n25048) );
  XNOR U25514 ( .A(n24953), .B(n24951), .Z(n25056) );
  AND U25515 ( .A(n25057), .B(n25058), .Z(n24951) );
  NANDN U25516 ( .A(n25059), .B(n25060), .Z(n25058) );
  OR U25517 ( .A(n25061), .B(n25062), .Z(n25060) );
  NAND U25518 ( .A(n25062), .B(n25061), .Z(n25057) );
  ANDN U25519 ( .B(B[93]), .A(n30), .Z(n24953) );
  XNOR U25520 ( .A(n24961), .B(n25063), .Z(n24954) );
  XNOR U25521 ( .A(n24960), .B(n24958), .Z(n25063) );
  AND U25522 ( .A(n25064), .B(n25065), .Z(n24958) );
  NANDN U25523 ( .A(n25066), .B(n25067), .Z(n25065) );
  NANDN U25524 ( .A(n25068), .B(n25069), .Z(n25067) );
  NANDN U25525 ( .A(n25069), .B(n25068), .Z(n25064) );
  ANDN U25526 ( .B(B[94]), .A(n31), .Z(n24960) );
  XNOR U25527 ( .A(n24968), .B(n25070), .Z(n24961) );
  XNOR U25528 ( .A(n24967), .B(n24965), .Z(n25070) );
  AND U25529 ( .A(n25071), .B(n25072), .Z(n24965) );
  NANDN U25530 ( .A(n25073), .B(n25074), .Z(n25072) );
  OR U25531 ( .A(n25075), .B(n25076), .Z(n25074) );
  NAND U25532 ( .A(n25076), .B(n25075), .Z(n25071) );
  ANDN U25533 ( .B(B[95]), .A(n32), .Z(n24967) );
  XNOR U25534 ( .A(n24975), .B(n25077), .Z(n24968) );
  XNOR U25535 ( .A(n24974), .B(n24972), .Z(n25077) );
  AND U25536 ( .A(n25078), .B(n25079), .Z(n24972) );
  NANDN U25537 ( .A(n25080), .B(n25081), .Z(n25079) );
  NANDN U25538 ( .A(n25082), .B(n25083), .Z(n25081) );
  NANDN U25539 ( .A(n25083), .B(n25082), .Z(n25078) );
  ANDN U25540 ( .B(A[11]), .A(n10), .Z(n24974) );
  XNOR U25541 ( .A(n24982), .B(n25084), .Z(n24975) );
  XNOR U25542 ( .A(n24981), .B(n24979), .Z(n25084) );
  AND U25543 ( .A(n25085), .B(n25086), .Z(n24979) );
  NANDN U25544 ( .A(n25087), .B(n25088), .Z(n25086) );
  OR U25545 ( .A(n25089), .B(n25090), .Z(n25088) );
  NAND U25546 ( .A(n25090), .B(n25089), .Z(n25085) );
  ANDN U25547 ( .B(A[10]), .A(n8), .Z(n24981) );
  XNOR U25548 ( .A(n24989), .B(n25091), .Z(n24982) );
  XNOR U25549 ( .A(n24988), .B(n24986), .Z(n25091) );
  AND U25550 ( .A(n25092), .B(n25093), .Z(n24986) );
  NANDN U25551 ( .A(n25094), .B(n25095), .Z(n25093) );
  NANDN U25552 ( .A(n25096), .B(n25097), .Z(n25095) );
  NANDN U25553 ( .A(n25097), .B(n25096), .Z(n25092) );
  ANDN U25554 ( .B(B[98]), .A(n35), .Z(n24988) );
  XNOR U25555 ( .A(n24996), .B(n25098), .Z(n24989) );
  XNOR U25556 ( .A(n24995), .B(n24993), .Z(n25098) );
  AND U25557 ( .A(n25099), .B(n25100), .Z(n24993) );
  NANDN U25558 ( .A(n25101), .B(n25102), .Z(n25100) );
  OR U25559 ( .A(n25103), .B(n25104), .Z(n25102) );
  NAND U25560 ( .A(n25104), .B(n25103), .Z(n25099) );
  ANDN U25561 ( .B(A[8]), .A(n5), .Z(n24995) );
  XNOR U25562 ( .A(n25003), .B(n25105), .Z(n24996) );
  XNOR U25563 ( .A(n25002), .B(n25000), .Z(n25105) );
  AND U25564 ( .A(n25106), .B(n25107), .Z(n25000) );
  NANDN U25565 ( .A(n25108), .B(n25109), .Z(n25107) );
  NANDN U25566 ( .A(n25110), .B(n25111), .Z(n25109) );
  NANDN U25567 ( .A(n25111), .B(n25110), .Z(n25106) );
  ANDN U25568 ( .B(A[7]), .A(n3), .Z(n25002) );
  XNOR U25569 ( .A(n25010), .B(n25112), .Z(n25003) );
  XNOR U25570 ( .A(n25009), .B(n25007), .Z(n25112) );
  AND U25571 ( .A(n25113), .B(n25114), .Z(n25007) );
  NANDN U25572 ( .A(n25115), .B(n25116), .Z(n25114) );
  OR U25573 ( .A(n25117), .B(n25118), .Z(n25116) );
  NAND U25574 ( .A(n25118), .B(n25117), .Z(n25113) );
  ANDN U25575 ( .B(B[101]), .A(n38), .Z(n25009) );
  XNOR U25576 ( .A(n25017), .B(n25119), .Z(n25010) );
  XNOR U25577 ( .A(n25016), .B(n25014), .Z(n25119) );
  AND U25578 ( .A(n25120), .B(n25121), .Z(n25014) );
  NANDN U25579 ( .A(n25122), .B(n25123), .Z(n25121) );
  NANDN U25580 ( .A(n25124), .B(n25125), .Z(n25123) );
  NANDN U25581 ( .A(n25125), .B(n25124), .Z(n25120) );
  ANDN U25582 ( .B(B[102]), .A(n39), .Z(n25016) );
  XNOR U25583 ( .A(n25024), .B(n25126), .Z(n25017) );
  XNOR U25584 ( .A(n25023), .B(n25021), .Z(n25126) );
  AND U25585 ( .A(n25127), .B(n25128), .Z(n25021) );
  NANDN U25586 ( .A(n25129), .B(n25130), .Z(n25128) );
  OR U25587 ( .A(n25131), .B(n25132), .Z(n25130) );
  NAND U25588 ( .A(n25132), .B(n25131), .Z(n25127) );
  ANDN U25589 ( .B(B[103]), .A(n40), .Z(n25023) );
  XNOR U25590 ( .A(n25031), .B(n25133), .Z(n25024) );
  XNOR U25591 ( .A(n25030), .B(n25028), .Z(n25133) );
  AND U25592 ( .A(n25134), .B(n25135), .Z(n25028) );
  NANDN U25593 ( .A(n25136), .B(n25137), .Z(n25135) );
  NAND U25594 ( .A(n25138), .B(n25139), .Z(n25137) );
  ANDN U25595 ( .B(B[104]), .A(n41), .Z(n25030) );
  XOR U25596 ( .A(n25037), .B(n25140), .Z(n25031) );
  XNOR U25597 ( .A(n25035), .B(n25038), .Z(n25140) );
  NAND U25598 ( .A(A[2]), .B(B[105]), .Z(n25038) );
  NANDN U25599 ( .A(n25141), .B(n25142), .Z(n25035) );
  AND U25600 ( .A(A[0]), .B(B[106]), .Z(n25142) );
  XNOR U25601 ( .A(n25040), .B(n25143), .Z(n25037) );
  NAND U25602 ( .A(A[0]), .B(B[107]), .Z(n25143) );
  NAND U25603 ( .A(B[106]), .B(A[1]), .Z(n25040) );
  NAND U25604 ( .A(n25144), .B(n25145), .Z(n541) );
  NANDN U25605 ( .A(n25146), .B(n25147), .Z(n25145) );
  OR U25606 ( .A(n25148), .B(n25149), .Z(n25147) );
  NAND U25607 ( .A(n25149), .B(n25148), .Z(n25144) );
  XOR U25608 ( .A(n543), .B(n542), .Z(\A1[104] ) );
  XOR U25609 ( .A(n25149), .B(n25150), .Z(n542) );
  XNOR U25610 ( .A(n25148), .B(n25146), .Z(n25150) );
  AND U25611 ( .A(n25151), .B(n25152), .Z(n25146) );
  NANDN U25612 ( .A(n25153), .B(n25154), .Z(n25152) );
  NANDN U25613 ( .A(n25155), .B(n25156), .Z(n25154) );
  NANDN U25614 ( .A(n25156), .B(n25155), .Z(n25151) );
  ANDN U25615 ( .B(B[91]), .A(n29), .Z(n25148) );
  XNOR U25616 ( .A(n25055), .B(n25157), .Z(n25149) );
  XNOR U25617 ( .A(n25054), .B(n25052), .Z(n25157) );
  AND U25618 ( .A(n25158), .B(n25159), .Z(n25052) );
  NANDN U25619 ( .A(n25160), .B(n25161), .Z(n25159) );
  OR U25620 ( .A(n25162), .B(n25163), .Z(n25161) );
  NAND U25621 ( .A(n25163), .B(n25162), .Z(n25158) );
  ANDN U25622 ( .B(B[92]), .A(n30), .Z(n25054) );
  XNOR U25623 ( .A(n25062), .B(n25164), .Z(n25055) );
  XNOR U25624 ( .A(n25061), .B(n25059), .Z(n25164) );
  AND U25625 ( .A(n25165), .B(n25166), .Z(n25059) );
  NANDN U25626 ( .A(n25167), .B(n25168), .Z(n25166) );
  NANDN U25627 ( .A(n25169), .B(n25170), .Z(n25168) );
  NANDN U25628 ( .A(n25170), .B(n25169), .Z(n25165) );
  ANDN U25629 ( .B(B[93]), .A(n31), .Z(n25061) );
  XNOR U25630 ( .A(n25069), .B(n25171), .Z(n25062) );
  XNOR U25631 ( .A(n25068), .B(n25066), .Z(n25171) );
  AND U25632 ( .A(n25172), .B(n25173), .Z(n25066) );
  NANDN U25633 ( .A(n25174), .B(n25175), .Z(n25173) );
  OR U25634 ( .A(n25176), .B(n25177), .Z(n25175) );
  NAND U25635 ( .A(n25177), .B(n25176), .Z(n25172) );
  ANDN U25636 ( .B(B[94]), .A(n32), .Z(n25068) );
  XNOR U25637 ( .A(n25076), .B(n25178), .Z(n25069) );
  XNOR U25638 ( .A(n25075), .B(n25073), .Z(n25178) );
  AND U25639 ( .A(n25179), .B(n25180), .Z(n25073) );
  NANDN U25640 ( .A(n25181), .B(n25182), .Z(n25180) );
  NANDN U25641 ( .A(n25183), .B(n25184), .Z(n25182) );
  NANDN U25642 ( .A(n25184), .B(n25183), .Z(n25179) );
  ANDN U25643 ( .B(A[11]), .A(n12), .Z(n25075) );
  XNOR U25644 ( .A(n25083), .B(n25185), .Z(n25076) );
  XNOR U25645 ( .A(n25082), .B(n25080), .Z(n25185) );
  AND U25646 ( .A(n25186), .B(n25187), .Z(n25080) );
  NANDN U25647 ( .A(n25188), .B(n25189), .Z(n25187) );
  OR U25648 ( .A(n25190), .B(n25191), .Z(n25189) );
  NAND U25649 ( .A(n25191), .B(n25190), .Z(n25186) );
  ANDN U25650 ( .B(A[10]), .A(n10), .Z(n25082) );
  XNOR U25651 ( .A(n25090), .B(n25192), .Z(n25083) );
  XNOR U25652 ( .A(n25089), .B(n25087), .Z(n25192) );
  AND U25653 ( .A(n25193), .B(n25194), .Z(n25087) );
  NANDN U25654 ( .A(n25195), .B(n25196), .Z(n25194) );
  NANDN U25655 ( .A(n25197), .B(n25198), .Z(n25196) );
  NANDN U25656 ( .A(n25198), .B(n25197), .Z(n25193) );
  ANDN U25657 ( .B(A[9]), .A(n8), .Z(n25089) );
  XNOR U25658 ( .A(n25097), .B(n25199), .Z(n25090) );
  XNOR U25659 ( .A(n25096), .B(n25094), .Z(n25199) );
  AND U25660 ( .A(n25200), .B(n25201), .Z(n25094) );
  NANDN U25661 ( .A(n25202), .B(n25203), .Z(n25201) );
  OR U25662 ( .A(n25204), .B(n25205), .Z(n25203) );
  NAND U25663 ( .A(n25205), .B(n25204), .Z(n25200) );
  ANDN U25664 ( .B(B[98]), .A(n36), .Z(n25096) );
  XNOR U25665 ( .A(n25104), .B(n25206), .Z(n25097) );
  XNOR U25666 ( .A(n25103), .B(n25101), .Z(n25206) );
  AND U25667 ( .A(n25207), .B(n25208), .Z(n25101) );
  NANDN U25668 ( .A(n25209), .B(n25210), .Z(n25208) );
  NANDN U25669 ( .A(n25211), .B(n25212), .Z(n25210) );
  NANDN U25670 ( .A(n25212), .B(n25211), .Z(n25207) );
  ANDN U25671 ( .B(A[7]), .A(n5), .Z(n25103) );
  XNOR U25672 ( .A(n25111), .B(n25213), .Z(n25104) );
  XNOR U25673 ( .A(n25110), .B(n25108), .Z(n25213) );
  AND U25674 ( .A(n25214), .B(n25215), .Z(n25108) );
  NANDN U25675 ( .A(n25216), .B(n25217), .Z(n25215) );
  OR U25676 ( .A(n25218), .B(n25219), .Z(n25217) );
  NAND U25677 ( .A(n25219), .B(n25218), .Z(n25214) );
  ANDN U25678 ( .B(A[6]), .A(n3), .Z(n25110) );
  XNOR U25679 ( .A(n25118), .B(n25220), .Z(n25111) );
  XNOR U25680 ( .A(n25117), .B(n25115), .Z(n25220) );
  AND U25681 ( .A(n25221), .B(n25222), .Z(n25115) );
  NANDN U25682 ( .A(n25223), .B(n25224), .Z(n25222) );
  NANDN U25683 ( .A(n25225), .B(n25226), .Z(n25224) );
  NANDN U25684 ( .A(n25226), .B(n25225), .Z(n25221) );
  ANDN U25685 ( .B(B[101]), .A(n39), .Z(n25117) );
  XNOR U25686 ( .A(n25125), .B(n25227), .Z(n25118) );
  XNOR U25687 ( .A(n25124), .B(n25122), .Z(n25227) );
  AND U25688 ( .A(n25228), .B(n25229), .Z(n25122) );
  NANDN U25689 ( .A(n25230), .B(n25231), .Z(n25229) );
  OR U25690 ( .A(n25232), .B(n25233), .Z(n25231) );
  NAND U25691 ( .A(n25233), .B(n25232), .Z(n25228) );
  ANDN U25692 ( .B(B[102]), .A(n40), .Z(n25124) );
  XNOR U25693 ( .A(n25132), .B(n25234), .Z(n25125) );
  XNOR U25694 ( .A(n25131), .B(n25129), .Z(n25234) );
  AND U25695 ( .A(n25235), .B(n25236), .Z(n25129) );
  NANDN U25696 ( .A(n25237), .B(n25238), .Z(n25236) );
  NAND U25697 ( .A(n25239), .B(n25240), .Z(n25238) );
  ANDN U25698 ( .B(B[103]), .A(n41), .Z(n25131) );
  XOR U25699 ( .A(n25138), .B(n25241), .Z(n25132) );
  XNOR U25700 ( .A(n25136), .B(n25139), .Z(n25241) );
  NAND U25701 ( .A(A[2]), .B(B[104]), .Z(n25139) );
  NANDN U25702 ( .A(n25242), .B(n25243), .Z(n25136) );
  AND U25703 ( .A(A[0]), .B(B[105]), .Z(n25243) );
  XNOR U25704 ( .A(n25141), .B(n25244), .Z(n25138) );
  NAND U25705 ( .A(A[0]), .B(B[106]), .Z(n25244) );
  NAND U25706 ( .A(B[105]), .B(A[1]), .Z(n25141) );
  NAND U25707 ( .A(n25245), .B(n25246), .Z(n543) );
  NANDN U25708 ( .A(n25247), .B(n25248), .Z(n25246) );
  OR U25709 ( .A(n25249), .B(n25250), .Z(n25248) );
  NAND U25710 ( .A(n25250), .B(n25249), .Z(n25245) );
  XOR U25711 ( .A(n545), .B(n544), .Z(\A1[103] ) );
  XOR U25712 ( .A(n25250), .B(n25251), .Z(n544) );
  XNOR U25713 ( .A(n25249), .B(n25247), .Z(n25251) );
  AND U25714 ( .A(n25252), .B(n25253), .Z(n25247) );
  NANDN U25715 ( .A(n25254), .B(n25255), .Z(n25253) );
  NANDN U25716 ( .A(n25256), .B(n25257), .Z(n25255) );
  NANDN U25717 ( .A(n25257), .B(n25256), .Z(n25252) );
  ANDN U25718 ( .B(B[90]), .A(n29), .Z(n25249) );
  XNOR U25719 ( .A(n25156), .B(n25258), .Z(n25250) );
  XNOR U25720 ( .A(n25155), .B(n25153), .Z(n25258) );
  AND U25721 ( .A(n25259), .B(n25260), .Z(n25153) );
  NANDN U25722 ( .A(n25261), .B(n25262), .Z(n25260) );
  OR U25723 ( .A(n25263), .B(n25264), .Z(n25262) );
  NAND U25724 ( .A(n25264), .B(n25263), .Z(n25259) );
  ANDN U25725 ( .B(B[91]), .A(n30), .Z(n25155) );
  XNOR U25726 ( .A(n25163), .B(n25265), .Z(n25156) );
  XNOR U25727 ( .A(n25162), .B(n25160), .Z(n25265) );
  AND U25728 ( .A(n25266), .B(n25267), .Z(n25160) );
  NANDN U25729 ( .A(n25268), .B(n25269), .Z(n25267) );
  NANDN U25730 ( .A(n25270), .B(n25271), .Z(n25269) );
  NANDN U25731 ( .A(n25271), .B(n25270), .Z(n25266) );
  ANDN U25732 ( .B(B[92]), .A(n31), .Z(n25162) );
  XNOR U25733 ( .A(n25170), .B(n25272), .Z(n25163) );
  XNOR U25734 ( .A(n25169), .B(n25167), .Z(n25272) );
  AND U25735 ( .A(n25273), .B(n25274), .Z(n25167) );
  NANDN U25736 ( .A(n25275), .B(n25276), .Z(n25274) );
  OR U25737 ( .A(n25277), .B(n25278), .Z(n25276) );
  NAND U25738 ( .A(n25278), .B(n25277), .Z(n25273) );
  ANDN U25739 ( .B(B[93]), .A(n32), .Z(n25169) );
  XNOR U25740 ( .A(n25177), .B(n25279), .Z(n25170) );
  XNOR U25741 ( .A(n25176), .B(n25174), .Z(n25279) );
  AND U25742 ( .A(n25280), .B(n25281), .Z(n25174) );
  NANDN U25743 ( .A(n25282), .B(n25283), .Z(n25281) );
  NANDN U25744 ( .A(n25284), .B(n25285), .Z(n25283) );
  NANDN U25745 ( .A(n25285), .B(n25284), .Z(n25280) );
  ANDN U25746 ( .B(B[94]), .A(n33), .Z(n25176) );
  XNOR U25747 ( .A(n25184), .B(n25286), .Z(n25177) );
  XNOR U25748 ( .A(n25183), .B(n25181), .Z(n25286) );
  AND U25749 ( .A(n25287), .B(n25288), .Z(n25181) );
  NANDN U25750 ( .A(n25289), .B(n25290), .Z(n25288) );
  OR U25751 ( .A(n25291), .B(n25292), .Z(n25290) );
  NAND U25752 ( .A(n25292), .B(n25291), .Z(n25287) );
  ANDN U25753 ( .B(A[10]), .A(n12), .Z(n25183) );
  XNOR U25754 ( .A(n25191), .B(n25293), .Z(n25184) );
  XNOR U25755 ( .A(n25190), .B(n25188), .Z(n25293) );
  AND U25756 ( .A(n25294), .B(n25295), .Z(n25188) );
  NANDN U25757 ( .A(n25296), .B(n25297), .Z(n25295) );
  NANDN U25758 ( .A(n25298), .B(n25299), .Z(n25297) );
  NANDN U25759 ( .A(n25299), .B(n25298), .Z(n25294) );
  ANDN U25760 ( .B(A[9]), .A(n10), .Z(n25190) );
  XNOR U25761 ( .A(n25198), .B(n25300), .Z(n25191) );
  XNOR U25762 ( .A(n25197), .B(n25195), .Z(n25300) );
  AND U25763 ( .A(n25301), .B(n25302), .Z(n25195) );
  NANDN U25764 ( .A(n25303), .B(n25304), .Z(n25302) );
  OR U25765 ( .A(n25305), .B(n25306), .Z(n25304) );
  NAND U25766 ( .A(n25306), .B(n25305), .Z(n25301) );
  ANDN U25767 ( .B(A[8]), .A(n8), .Z(n25197) );
  XNOR U25768 ( .A(n25205), .B(n25307), .Z(n25198) );
  XNOR U25769 ( .A(n25204), .B(n25202), .Z(n25307) );
  AND U25770 ( .A(n25308), .B(n25309), .Z(n25202) );
  NANDN U25771 ( .A(n25310), .B(n25311), .Z(n25309) );
  NANDN U25772 ( .A(n25312), .B(n25313), .Z(n25311) );
  NANDN U25773 ( .A(n25313), .B(n25312), .Z(n25308) );
  ANDN U25774 ( .B(B[98]), .A(n37), .Z(n25204) );
  XNOR U25775 ( .A(n25212), .B(n25314), .Z(n25205) );
  XNOR U25776 ( .A(n25211), .B(n25209), .Z(n25314) );
  AND U25777 ( .A(n25315), .B(n25316), .Z(n25209) );
  NANDN U25778 ( .A(n25317), .B(n25318), .Z(n25316) );
  OR U25779 ( .A(n25319), .B(n25320), .Z(n25318) );
  NAND U25780 ( .A(n25320), .B(n25319), .Z(n25315) );
  ANDN U25781 ( .B(A[6]), .A(n5), .Z(n25211) );
  XNOR U25782 ( .A(n25219), .B(n25321), .Z(n25212) );
  XNOR U25783 ( .A(n25218), .B(n25216), .Z(n25321) );
  AND U25784 ( .A(n25322), .B(n25323), .Z(n25216) );
  NANDN U25785 ( .A(n25324), .B(n25325), .Z(n25323) );
  NANDN U25786 ( .A(n25326), .B(n25327), .Z(n25325) );
  NANDN U25787 ( .A(n25327), .B(n25326), .Z(n25322) );
  ANDN U25788 ( .B(A[5]), .A(n3), .Z(n25218) );
  XNOR U25789 ( .A(n25226), .B(n25328), .Z(n25219) );
  XNOR U25790 ( .A(n25225), .B(n25223), .Z(n25328) );
  AND U25791 ( .A(n25329), .B(n25330), .Z(n25223) );
  NANDN U25792 ( .A(n25331), .B(n25332), .Z(n25330) );
  OR U25793 ( .A(n25333), .B(n25334), .Z(n25332) );
  NAND U25794 ( .A(n25334), .B(n25333), .Z(n25329) );
  ANDN U25795 ( .B(B[101]), .A(n40), .Z(n25225) );
  XNOR U25796 ( .A(n25233), .B(n25335), .Z(n25226) );
  XNOR U25797 ( .A(n25232), .B(n25230), .Z(n25335) );
  AND U25798 ( .A(n25336), .B(n25337), .Z(n25230) );
  NANDN U25799 ( .A(n25338), .B(n25339), .Z(n25337) );
  NAND U25800 ( .A(n25340), .B(n25341), .Z(n25339) );
  ANDN U25801 ( .B(B[102]), .A(n41), .Z(n25232) );
  XOR U25802 ( .A(n25239), .B(n25342), .Z(n25233) );
  XNOR U25803 ( .A(n25237), .B(n25240), .Z(n25342) );
  NAND U25804 ( .A(A[2]), .B(B[103]), .Z(n25240) );
  NANDN U25805 ( .A(n25343), .B(n25344), .Z(n25237) );
  AND U25806 ( .A(A[0]), .B(B[104]), .Z(n25344) );
  XNOR U25807 ( .A(n25242), .B(n25345), .Z(n25239) );
  NAND U25808 ( .A(A[0]), .B(B[105]), .Z(n25345) );
  NAND U25809 ( .A(B[104]), .B(A[1]), .Z(n25242) );
  NAND U25810 ( .A(n25346), .B(n25347), .Z(n545) );
  NANDN U25811 ( .A(n25348), .B(n25349), .Z(n25347) );
  OR U25812 ( .A(n25350), .B(n25351), .Z(n25349) );
  NAND U25813 ( .A(n25351), .B(n25350), .Z(n25346) );
  XOR U25814 ( .A(n547), .B(n546), .Z(\A1[102] ) );
  XOR U25815 ( .A(n25351), .B(n25352), .Z(n546) );
  XNOR U25816 ( .A(n25350), .B(n25348), .Z(n25352) );
  AND U25817 ( .A(n25353), .B(n25354), .Z(n25348) );
  NANDN U25818 ( .A(n25355), .B(n25356), .Z(n25354) );
  NANDN U25819 ( .A(n25357), .B(n25358), .Z(n25356) );
  NANDN U25820 ( .A(n25358), .B(n25357), .Z(n25353) );
  ANDN U25821 ( .B(B[89]), .A(n29), .Z(n25350) );
  XNOR U25822 ( .A(n25257), .B(n25359), .Z(n25351) );
  XNOR U25823 ( .A(n25256), .B(n25254), .Z(n25359) );
  AND U25824 ( .A(n25360), .B(n25361), .Z(n25254) );
  NANDN U25825 ( .A(n25362), .B(n25363), .Z(n25361) );
  OR U25826 ( .A(n25364), .B(n25365), .Z(n25363) );
  NAND U25827 ( .A(n25365), .B(n25364), .Z(n25360) );
  ANDN U25828 ( .B(B[90]), .A(n30), .Z(n25256) );
  XNOR U25829 ( .A(n25264), .B(n25366), .Z(n25257) );
  XNOR U25830 ( .A(n25263), .B(n25261), .Z(n25366) );
  AND U25831 ( .A(n25367), .B(n25368), .Z(n25261) );
  NANDN U25832 ( .A(n25369), .B(n25370), .Z(n25368) );
  NANDN U25833 ( .A(n25371), .B(n25372), .Z(n25370) );
  NANDN U25834 ( .A(n25372), .B(n25371), .Z(n25367) );
  ANDN U25835 ( .B(B[91]), .A(n31), .Z(n25263) );
  XNOR U25836 ( .A(n25271), .B(n25373), .Z(n25264) );
  XNOR U25837 ( .A(n25270), .B(n25268), .Z(n25373) );
  AND U25838 ( .A(n25374), .B(n25375), .Z(n25268) );
  NANDN U25839 ( .A(n25376), .B(n25377), .Z(n25375) );
  OR U25840 ( .A(n25378), .B(n25379), .Z(n25377) );
  NAND U25841 ( .A(n25379), .B(n25378), .Z(n25374) );
  ANDN U25842 ( .B(B[92]), .A(n32), .Z(n25270) );
  XNOR U25843 ( .A(n25278), .B(n25380), .Z(n25271) );
  XNOR U25844 ( .A(n25277), .B(n25275), .Z(n25380) );
  AND U25845 ( .A(n25381), .B(n25382), .Z(n25275) );
  NANDN U25846 ( .A(n25383), .B(n25384), .Z(n25382) );
  NANDN U25847 ( .A(n25385), .B(n25386), .Z(n25384) );
  NANDN U25848 ( .A(n25386), .B(n25385), .Z(n25381) );
  ANDN U25849 ( .B(B[93]), .A(n33), .Z(n25277) );
  XNOR U25850 ( .A(n25285), .B(n25387), .Z(n25278) );
  XNOR U25851 ( .A(n25284), .B(n25282), .Z(n25387) );
  AND U25852 ( .A(n25388), .B(n25389), .Z(n25282) );
  NANDN U25853 ( .A(n25390), .B(n25391), .Z(n25389) );
  OR U25854 ( .A(n25392), .B(n25393), .Z(n25391) );
  NAND U25855 ( .A(n25393), .B(n25392), .Z(n25388) );
  ANDN U25856 ( .B(A[10]), .A(n14), .Z(n25284) );
  XNOR U25857 ( .A(n25292), .B(n25394), .Z(n25285) );
  XNOR U25858 ( .A(n25291), .B(n25289), .Z(n25394) );
  AND U25859 ( .A(n25395), .B(n25396), .Z(n25289) );
  NANDN U25860 ( .A(n25397), .B(n25398), .Z(n25396) );
  NANDN U25861 ( .A(n25399), .B(n25400), .Z(n25398) );
  NANDN U25862 ( .A(n25400), .B(n25399), .Z(n25395) );
  ANDN U25863 ( .B(A[9]), .A(n12), .Z(n25291) );
  XNOR U25864 ( .A(n25299), .B(n25401), .Z(n25292) );
  XNOR U25865 ( .A(n25298), .B(n25296), .Z(n25401) );
  AND U25866 ( .A(n25402), .B(n25403), .Z(n25296) );
  NANDN U25867 ( .A(n25404), .B(n25405), .Z(n25403) );
  OR U25868 ( .A(n25406), .B(n25407), .Z(n25405) );
  NAND U25869 ( .A(n25407), .B(n25406), .Z(n25402) );
  ANDN U25870 ( .B(A[8]), .A(n10), .Z(n25298) );
  XNOR U25871 ( .A(n25306), .B(n25408), .Z(n25299) );
  XNOR U25872 ( .A(n25305), .B(n25303), .Z(n25408) );
  AND U25873 ( .A(n25409), .B(n25410), .Z(n25303) );
  NANDN U25874 ( .A(n25411), .B(n25412), .Z(n25410) );
  NANDN U25875 ( .A(n25413), .B(n25414), .Z(n25412) );
  NANDN U25876 ( .A(n25414), .B(n25413), .Z(n25409) );
  ANDN U25877 ( .B(A[7]), .A(n8), .Z(n25305) );
  XNOR U25878 ( .A(n25313), .B(n25415), .Z(n25306) );
  XNOR U25879 ( .A(n25312), .B(n25310), .Z(n25415) );
  AND U25880 ( .A(n25416), .B(n25417), .Z(n25310) );
  NANDN U25881 ( .A(n25418), .B(n25419), .Z(n25417) );
  OR U25882 ( .A(n25420), .B(n25421), .Z(n25419) );
  NAND U25883 ( .A(n25421), .B(n25420), .Z(n25416) );
  ANDN U25884 ( .B(B[98]), .A(n38), .Z(n25312) );
  XNOR U25885 ( .A(n25320), .B(n25422), .Z(n25313) );
  XNOR U25886 ( .A(n25319), .B(n25317), .Z(n25422) );
  AND U25887 ( .A(n25423), .B(n25424), .Z(n25317) );
  NANDN U25888 ( .A(n25425), .B(n25426), .Z(n25424) );
  NANDN U25889 ( .A(n25427), .B(n25428), .Z(n25426) );
  NANDN U25890 ( .A(n25428), .B(n25427), .Z(n25423) );
  ANDN U25891 ( .B(A[5]), .A(n5), .Z(n25319) );
  XNOR U25892 ( .A(n25327), .B(n25429), .Z(n25320) );
  XNOR U25893 ( .A(n25326), .B(n25324), .Z(n25429) );
  AND U25894 ( .A(n25430), .B(n25431), .Z(n25324) );
  NANDN U25895 ( .A(n25432), .B(n25433), .Z(n25431) );
  OR U25896 ( .A(n25434), .B(n25435), .Z(n25433) );
  NAND U25897 ( .A(n25435), .B(n25434), .Z(n25430) );
  ANDN U25898 ( .B(A[4]), .A(n3), .Z(n25326) );
  XNOR U25899 ( .A(n25334), .B(n25436), .Z(n25327) );
  XNOR U25900 ( .A(n25333), .B(n25331), .Z(n25436) );
  AND U25901 ( .A(n25437), .B(n25438), .Z(n25331) );
  NANDN U25902 ( .A(n25439), .B(n25440), .Z(n25438) );
  NAND U25903 ( .A(n25441), .B(n25442), .Z(n25440) );
  ANDN U25904 ( .B(B[101]), .A(n41), .Z(n25333) );
  XOR U25905 ( .A(n25340), .B(n25443), .Z(n25334) );
  XNOR U25906 ( .A(n25338), .B(n25341), .Z(n25443) );
  NAND U25907 ( .A(A[2]), .B(B[102]), .Z(n25341) );
  NANDN U25908 ( .A(n25444), .B(n25445), .Z(n25338) );
  AND U25909 ( .A(A[0]), .B(B[103]), .Z(n25445) );
  XNOR U25910 ( .A(n25343), .B(n25446), .Z(n25340) );
  NAND U25911 ( .A(A[0]), .B(B[104]), .Z(n25446) );
  NAND U25912 ( .A(B[103]), .B(A[1]), .Z(n25343) );
  NAND U25913 ( .A(n25447), .B(n25448), .Z(n547) );
  NANDN U25914 ( .A(n25449), .B(n25450), .Z(n25448) );
  OR U25915 ( .A(n25451), .B(n25452), .Z(n25450) );
  NAND U25916 ( .A(n25452), .B(n25451), .Z(n25447) );
  XOR U25917 ( .A(n549), .B(n548), .Z(\A1[101] ) );
  XOR U25918 ( .A(n25452), .B(n25453), .Z(n548) );
  XNOR U25919 ( .A(n25451), .B(n25449), .Z(n25453) );
  AND U25920 ( .A(n25454), .B(n25455), .Z(n25449) );
  NANDN U25921 ( .A(n25456), .B(n25457), .Z(n25455) );
  NANDN U25922 ( .A(n25458), .B(n25459), .Z(n25457) );
  NANDN U25923 ( .A(n25459), .B(n25458), .Z(n25454) );
  ANDN U25924 ( .B(B[88]), .A(n29), .Z(n25451) );
  XNOR U25925 ( .A(n25358), .B(n25460), .Z(n25452) );
  XNOR U25926 ( .A(n25357), .B(n25355), .Z(n25460) );
  AND U25927 ( .A(n25461), .B(n25462), .Z(n25355) );
  NANDN U25928 ( .A(n25463), .B(n25464), .Z(n25462) );
  OR U25929 ( .A(n25465), .B(n25466), .Z(n25464) );
  NAND U25930 ( .A(n25466), .B(n25465), .Z(n25461) );
  ANDN U25931 ( .B(B[89]), .A(n30), .Z(n25357) );
  XNOR U25932 ( .A(n25365), .B(n25467), .Z(n25358) );
  XNOR U25933 ( .A(n25364), .B(n25362), .Z(n25467) );
  AND U25934 ( .A(n25468), .B(n25469), .Z(n25362) );
  NANDN U25935 ( .A(n25470), .B(n25471), .Z(n25469) );
  NANDN U25936 ( .A(n25472), .B(n25473), .Z(n25471) );
  NANDN U25937 ( .A(n25473), .B(n25472), .Z(n25468) );
  ANDN U25938 ( .B(B[90]), .A(n31), .Z(n25364) );
  XNOR U25939 ( .A(n25372), .B(n25474), .Z(n25365) );
  XNOR U25940 ( .A(n25371), .B(n25369), .Z(n25474) );
  AND U25941 ( .A(n25475), .B(n25476), .Z(n25369) );
  NANDN U25942 ( .A(n25477), .B(n25478), .Z(n25476) );
  OR U25943 ( .A(n25479), .B(n25480), .Z(n25478) );
  NAND U25944 ( .A(n25480), .B(n25479), .Z(n25475) );
  ANDN U25945 ( .B(B[91]), .A(n32), .Z(n25371) );
  XNOR U25946 ( .A(n25379), .B(n25481), .Z(n25372) );
  XNOR U25947 ( .A(n25378), .B(n25376), .Z(n25481) );
  AND U25948 ( .A(n25482), .B(n25483), .Z(n25376) );
  NANDN U25949 ( .A(n25484), .B(n25485), .Z(n25483) );
  NANDN U25950 ( .A(n25486), .B(n25487), .Z(n25485) );
  NANDN U25951 ( .A(n25487), .B(n25486), .Z(n25482) );
  ANDN U25952 ( .B(B[92]), .A(n33), .Z(n25378) );
  XNOR U25953 ( .A(n25386), .B(n25488), .Z(n25379) );
  XNOR U25954 ( .A(n25385), .B(n25383), .Z(n25488) );
  AND U25955 ( .A(n25489), .B(n25490), .Z(n25383) );
  NANDN U25956 ( .A(n25491), .B(n25492), .Z(n25490) );
  OR U25957 ( .A(n25493), .B(n25494), .Z(n25492) );
  NAND U25958 ( .A(n25494), .B(n25493), .Z(n25489) );
  ANDN U25959 ( .B(B[93]), .A(n34), .Z(n25385) );
  XNOR U25960 ( .A(n25393), .B(n25495), .Z(n25386) );
  XNOR U25961 ( .A(n25392), .B(n25390), .Z(n25495) );
  AND U25962 ( .A(n25496), .B(n25497), .Z(n25390) );
  NANDN U25963 ( .A(n25498), .B(n25499), .Z(n25497) );
  NANDN U25964 ( .A(n25500), .B(n25501), .Z(n25499) );
  NANDN U25965 ( .A(n25501), .B(n25500), .Z(n25496) );
  ANDN U25966 ( .B(A[9]), .A(n14), .Z(n25392) );
  XNOR U25967 ( .A(n25400), .B(n25502), .Z(n25393) );
  XNOR U25968 ( .A(n25399), .B(n25397), .Z(n25502) );
  AND U25969 ( .A(n25503), .B(n25504), .Z(n25397) );
  NANDN U25970 ( .A(n25505), .B(n25506), .Z(n25504) );
  OR U25971 ( .A(n25507), .B(n25508), .Z(n25506) );
  NAND U25972 ( .A(n25508), .B(n25507), .Z(n25503) );
  ANDN U25973 ( .B(A[8]), .A(n12), .Z(n25399) );
  XNOR U25974 ( .A(n25407), .B(n25509), .Z(n25400) );
  XNOR U25975 ( .A(n25406), .B(n25404), .Z(n25509) );
  AND U25976 ( .A(n25510), .B(n25511), .Z(n25404) );
  NANDN U25977 ( .A(n25512), .B(n25513), .Z(n25511) );
  NANDN U25978 ( .A(n25514), .B(n25515), .Z(n25513) );
  NANDN U25979 ( .A(n25515), .B(n25514), .Z(n25510) );
  ANDN U25980 ( .B(A[7]), .A(n10), .Z(n25406) );
  XNOR U25981 ( .A(n25414), .B(n25516), .Z(n25407) );
  XNOR U25982 ( .A(n25413), .B(n25411), .Z(n25516) );
  AND U25983 ( .A(n25517), .B(n25518), .Z(n25411) );
  NANDN U25984 ( .A(n25519), .B(n25520), .Z(n25518) );
  OR U25985 ( .A(n25521), .B(n25522), .Z(n25520) );
  NAND U25986 ( .A(n25522), .B(n25521), .Z(n25517) );
  ANDN U25987 ( .B(A[6]), .A(n8), .Z(n25413) );
  XNOR U25988 ( .A(n25421), .B(n25523), .Z(n25414) );
  XNOR U25989 ( .A(n25420), .B(n25418), .Z(n25523) );
  AND U25990 ( .A(n25524), .B(n25525), .Z(n25418) );
  NANDN U25991 ( .A(n25526), .B(n25527), .Z(n25525) );
  NANDN U25992 ( .A(n25528), .B(n25529), .Z(n25527) );
  NANDN U25993 ( .A(n25529), .B(n25528), .Z(n25524) );
  ANDN U25994 ( .B(B[98]), .A(n39), .Z(n25420) );
  XNOR U25995 ( .A(n25428), .B(n25530), .Z(n25421) );
  XNOR U25996 ( .A(n25427), .B(n25425), .Z(n25530) );
  AND U25997 ( .A(n25531), .B(n25532), .Z(n25425) );
  NANDN U25998 ( .A(n25533), .B(n25534), .Z(n25532) );
  OR U25999 ( .A(n25535), .B(n25536), .Z(n25534) );
  NAND U26000 ( .A(n25536), .B(n25535), .Z(n25531) );
  ANDN U26001 ( .B(A[4]), .A(n5), .Z(n25427) );
  XNOR U26002 ( .A(n25435), .B(n25537), .Z(n25428) );
  XNOR U26003 ( .A(n25434), .B(n25432), .Z(n25537) );
  AND U26004 ( .A(n25538), .B(n25539), .Z(n25432) );
  NANDN U26005 ( .A(n25540), .B(n25541), .Z(n25539) );
  NAND U26006 ( .A(n25542), .B(n25543), .Z(n25541) );
  ANDN U26007 ( .B(A[3]), .A(n3), .Z(n25434) );
  XOR U26008 ( .A(n25441), .B(n25544), .Z(n25435) );
  XNOR U26009 ( .A(n25439), .B(n25442), .Z(n25544) );
  NAND U26010 ( .A(A[2]), .B(B[101]), .Z(n25442) );
  NANDN U26011 ( .A(n25545), .B(n25546), .Z(n25439) );
  AND U26012 ( .A(A[0]), .B(B[102]), .Z(n25546) );
  XNOR U26013 ( .A(n25444), .B(n25547), .Z(n25441) );
  NAND U26014 ( .A(A[0]), .B(B[103]), .Z(n25547) );
  NAND U26015 ( .A(B[102]), .B(A[1]), .Z(n25444) );
  NAND U26016 ( .A(n25548), .B(n25549), .Z(n549) );
  NANDN U26017 ( .A(n25550), .B(n25551), .Z(n25549) );
  OR U26018 ( .A(n25552), .B(n25553), .Z(n25551) );
  NAND U26019 ( .A(n25553), .B(n25552), .Z(n25548) );
  XOR U26020 ( .A(n551), .B(n550), .Z(\A1[100] ) );
  XOR U26021 ( .A(n25553), .B(n25554), .Z(n550) );
  XNOR U26022 ( .A(n25552), .B(n25550), .Z(n25554) );
  AND U26023 ( .A(n25555), .B(n25556), .Z(n25550) );
  NANDN U26024 ( .A(n25557), .B(n25558), .Z(n25556) );
  NAND U26025 ( .A(n25560), .B(n25559), .Z(n25555) );
  ANDN U26026 ( .B(B[87]), .A(n29), .Z(n25552) );
  XNOR U26027 ( .A(n25459), .B(n25561), .Z(n25553) );
  XNOR U26028 ( .A(n25458), .B(n25456), .Z(n25561) );
  AND U26029 ( .A(n25562), .B(n25563), .Z(n25456) );
  NANDN U26030 ( .A(n25564), .B(n25565), .Z(n25563) );
  OR U26031 ( .A(n25566), .B(n25567), .Z(n25565) );
  NAND U26032 ( .A(n25567), .B(n25566), .Z(n25562) );
  ANDN U26033 ( .B(B[88]), .A(n30), .Z(n25458) );
  XNOR U26034 ( .A(n25466), .B(n25568), .Z(n25459) );
  XNOR U26035 ( .A(n25465), .B(n25463), .Z(n25568) );
  AND U26036 ( .A(n25569), .B(n25570), .Z(n25463) );
  NANDN U26037 ( .A(n25571), .B(n25572), .Z(n25570) );
  NANDN U26038 ( .A(n25573), .B(n25574), .Z(n25572) );
  NANDN U26039 ( .A(n25574), .B(n25573), .Z(n25569) );
  ANDN U26040 ( .B(B[89]), .A(n31), .Z(n25465) );
  XNOR U26041 ( .A(n25473), .B(n25575), .Z(n25466) );
  XNOR U26042 ( .A(n25472), .B(n25470), .Z(n25575) );
  AND U26043 ( .A(n25576), .B(n25577), .Z(n25470) );
  NANDN U26044 ( .A(n25578), .B(n25579), .Z(n25577) );
  OR U26045 ( .A(n25580), .B(n25581), .Z(n25579) );
  NAND U26046 ( .A(n25581), .B(n25580), .Z(n25576) );
  ANDN U26047 ( .B(B[90]), .A(n32), .Z(n25472) );
  XNOR U26048 ( .A(n25480), .B(n25582), .Z(n25473) );
  XNOR U26049 ( .A(n25479), .B(n25477), .Z(n25582) );
  AND U26050 ( .A(n25583), .B(n25584), .Z(n25477) );
  NANDN U26051 ( .A(n25585), .B(n25586), .Z(n25584) );
  NANDN U26052 ( .A(n25587), .B(n25588), .Z(n25586) );
  NANDN U26053 ( .A(n25588), .B(n25587), .Z(n25583) );
  ANDN U26054 ( .B(B[91]), .A(n33), .Z(n25479) );
  XNOR U26055 ( .A(n25487), .B(n25589), .Z(n25480) );
  XNOR U26056 ( .A(n25486), .B(n25484), .Z(n25589) );
  AND U26057 ( .A(n25590), .B(n25591), .Z(n25484) );
  NANDN U26058 ( .A(n25592), .B(n25593), .Z(n25591) );
  OR U26059 ( .A(n25594), .B(n25595), .Z(n25593) );
  NAND U26060 ( .A(n25595), .B(n25594), .Z(n25590) );
  ANDN U26061 ( .B(B[92]), .A(n34), .Z(n25486) );
  XNOR U26062 ( .A(n25494), .B(n25596), .Z(n25487) );
  XNOR U26063 ( .A(n25493), .B(n25491), .Z(n25596) );
  AND U26064 ( .A(n25597), .B(n25598), .Z(n25491) );
  NANDN U26065 ( .A(n25599), .B(n25600), .Z(n25598) );
  NANDN U26066 ( .A(n25601), .B(n25602), .Z(n25600) );
  NANDN U26067 ( .A(n25602), .B(n25601), .Z(n25597) );
  ANDN U26068 ( .B(A[9]), .A(n16), .Z(n25493) );
  XNOR U26069 ( .A(n25501), .B(n25603), .Z(n25494) );
  XNOR U26070 ( .A(n25500), .B(n25498), .Z(n25603) );
  AND U26071 ( .A(n25604), .B(n25605), .Z(n25498) );
  NANDN U26072 ( .A(n25606), .B(n25607), .Z(n25605) );
  OR U26073 ( .A(n25608), .B(n25609), .Z(n25607) );
  NAND U26074 ( .A(n25609), .B(n25608), .Z(n25604) );
  ANDN U26075 ( .B(A[8]), .A(n14), .Z(n25500) );
  XNOR U26076 ( .A(n25508), .B(n25610), .Z(n25501) );
  XNOR U26077 ( .A(n25507), .B(n25505), .Z(n25610) );
  AND U26078 ( .A(n25611), .B(n25612), .Z(n25505) );
  NANDN U26079 ( .A(n25613), .B(n25614), .Z(n25612) );
  NANDN U26080 ( .A(n25615), .B(n25616), .Z(n25614) );
  NANDN U26081 ( .A(n25616), .B(n25615), .Z(n25611) );
  ANDN U26082 ( .B(A[7]), .A(n12), .Z(n25507) );
  XNOR U26083 ( .A(n25515), .B(n25617), .Z(n25508) );
  XNOR U26084 ( .A(n25514), .B(n25512), .Z(n25617) );
  AND U26085 ( .A(n25618), .B(n25619), .Z(n25512) );
  NANDN U26086 ( .A(n25620), .B(n25621), .Z(n25619) );
  OR U26087 ( .A(n25622), .B(n25623), .Z(n25621) );
  NAND U26088 ( .A(n25623), .B(n25622), .Z(n25618) );
  ANDN U26089 ( .B(A[6]), .A(n10), .Z(n25514) );
  XNOR U26090 ( .A(n25522), .B(n25624), .Z(n25515) );
  XNOR U26091 ( .A(n25521), .B(n25519), .Z(n25624) );
  AND U26092 ( .A(n25625), .B(n25626), .Z(n25519) );
  NANDN U26093 ( .A(n25627), .B(n25628), .Z(n25626) );
  NANDN U26094 ( .A(n25629), .B(n25630), .Z(n25628) );
  NANDN U26095 ( .A(n25630), .B(n25629), .Z(n25625) );
  ANDN U26096 ( .B(A[5]), .A(n8), .Z(n25521) );
  XNOR U26097 ( .A(n25529), .B(n25631), .Z(n25522) );
  XNOR U26098 ( .A(n25528), .B(n25526), .Z(n25631) );
  AND U26099 ( .A(n25632), .B(n25633), .Z(n25526) );
  NANDN U26100 ( .A(n25634), .B(n25635), .Z(n25633) );
  OR U26101 ( .A(n25636), .B(n25637), .Z(n25635) );
  NAND U26102 ( .A(n25637), .B(n25636), .Z(n25632) );
  ANDN U26103 ( .B(B[98]), .A(n40), .Z(n25528) );
  XNOR U26104 ( .A(n25536), .B(n25638), .Z(n25529) );
  XNOR U26105 ( .A(n25535), .B(n25533), .Z(n25638) );
  AND U26106 ( .A(n25639), .B(n25640), .Z(n25533) );
  NANDN U26107 ( .A(n25641), .B(n25642), .Z(n25640) );
  NAND U26108 ( .A(n25643), .B(n25644), .Z(n25642) );
  ANDN U26109 ( .B(A[3]), .A(n5), .Z(n25535) );
  XOR U26110 ( .A(n25542), .B(n25645), .Z(n25536) );
  XNOR U26111 ( .A(n25540), .B(n25543), .Z(n25645) );
  NAND U26112 ( .A(B[100]), .B(A[2]), .Z(n25543) );
  NANDN U26113 ( .A(n25646), .B(n25647), .Z(n25540) );
  AND U26114 ( .A(A[0]), .B(B[101]), .Z(n25647) );
  XNOR U26115 ( .A(n25545), .B(n25648), .Z(n25542) );
  NAND U26116 ( .A(A[0]), .B(B[102]), .Z(n25648) );
  NAND U26117 ( .A(B[101]), .B(A[1]), .Z(n25545) );
  NAND U26118 ( .A(n25649), .B(n25650), .Z(n551) );
  NANDN U26119 ( .A(n559), .B(n25651), .Z(n25650) );
  NANDN U26120 ( .A(n557), .B(n25652), .Z(n25651) );
  NAND U26121 ( .A(A[15]), .B(B[86]), .Z(n559) );
  NAND U26122 ( .A(n4), .B(n557), .Z(n25649) );
  XOR U26123 ( .A(n25560), .B(n25653), .Z(n557) );
  XNOR U26124 ( .A(n25559), .B(n25557), .Z(n25653) );
  AND U26125 ( .A(n25654), .B(n25655), .Z(n25557) );
  NANDN U26126 ( .A(n25656), .B(n25657), .Z(n25655) );
  OR U26127 ( .A(n25658), .B(n25659), .Z(n25657) );
  NAND U26128 ( .A(n25659), .B(n25658), .Z(n25654) );
  ANDN U26129 ( .B(B[87]), .A(n30), .Z(n25559) );
  XOR U26130 ( .A(n25567), .B(n25660), .Z(n25560) );
  XNOR U26131 ( .A(n25566), .B(n25564), .Z(n25660) );
  AND U26132 ( .A(n25661), .B(n25662), .Z(n25564) );
  NANDN U26133 ( .A(n25663), .B(n25664), .Z(n25662) );
  NANDN U26134 ( .A(n25665), .B(n25666), .Z(n25664) );
  ANDN U26135 ( .B(B[88]), .A(n31), .Z(n25566) );
  XNOR U26136 ( .A(n25574), .B(n25667), .Z(n25567) );
  XNOR U26137 ( .A(n25573), .B(n25571), .Z(n25667) );
  AND U26138 ( .A(n25668), .B(n25669), .Z(n25571) );
  NANDN U26139 ( .A(n25670), .B(n25671), .Z(n25669) );
  OR U26140 ( .A(n25672), .B(n25673), .Z(n25671) );
  NAND U26141 ( .A(n25673), .B(n25672), .Z(n25668) );
  ANDN U26142 ( .B(B[89]), .A(n32), .Z(n25573) );
  XNOR U26143 ( .A(n25581), .B(n25674), .Z(n25574) );
  XNOR U26144 ( .A(n25580), .B(n25578), .Z(n25674) );
  AND U26145 ( .A(n25675), .B(n25676), .Z(n25578) );
  NANDN U26146 ( .A(n25677), .B(n25678), .Z(n25676) );
  NANDN U26147 ( .A(n25679), .B(n25680), .Z(n25678) );
  ANDN U26148 ( .B(B[90]), .A(n33), .Z(n25580) );
  XNOR U26149 ( .A(n25588), .B(n25681), .Z(n25581) );
  XNOR U26150 ( .A(n25587), .B(n25585), .Z(n25681) );
  AND U26151 ( .A(n25682), .B(n25683), .Z(n25585) );
  NANDN U26152 ( .A(n25684), .B(n25685), .Z(n25683) );
  OR U26153 ( .A(n25686), .B(n25687), .Z(n25685) );
  NAND U26154 ( .A(n25687), .B(n25686), .Z(n25682) );
  ANDN U26155 ( .B(B[91]), .A(n34), .Z(n25587) );
  XNOR U26156 ( .A(n25595), .B(n25688), .Z(n25588) );
  XNOR U26157 ( .A(n25594), .B(n25592), .Z(n25688) );
  AND U26158 ( .A(n25689), .B(n25690), .Z(n25592) );
  NANDN U26159 ( .A(n25691), .B(n25692), .Z(n25690) );
  NANDN U26160 ( .A(n25693), .B(n25694), .Z(n25692) );
  ANDN U26161 ( .B(B[92]), .A(n35), .Z(n25594) );
  XNOR U26162 ( .A(n25602), .B(n25695), .Z(n25595) );
  XNOR U26163 ( .A(n25601), .B(n25599), .Z(n25695) );
  AND U26164 ( .A(n25696), .B(n25697), .Z(n25599) );
  NANDN U26165 ( .A(n25698), .B(n25699), .Z(n25697) );
  OR U26166 ( .A(n25700), .B(n25701), .Z(n25699) );
  NAND U26167 ( .A(n25701), .B(n25700), .Z(n25696) );
  ANDN U26168 ( .B(A[8]), .A(n16), .Z(n25601) );
  XNOR U26169 ( .A(n25609), .B(n25702), .Z(n25602) );
  XNOR U26170 ( .A(n25608), .B(n25606), .Z(n25702) );
  AND U26171 ( .A(n25703), .B(n25704), .Z(n25606) );
  NANDN U26172 ( .A(n25705), .B(n25706), .Z(n25704) );
  NANDN U26173 ( .A(n25707), .B(n25708), .Z(n25706) );
  ANDN U26174 ( .B(A[7]), .A(n14), .Z(n25608) );
  XNOR U26175 ( .A(n25616), .B(n25709), .Z(n25609) );
  XNOR U26176 ( .A(n25615), .B(n25613), .Z(n25709) );
  AND U26177 ( .A(n25710), .B(n25711), .Z(n25613) );
  NANDN U26178 ( .A(n25712), .B(n25713), .Z(n25711) );
  OR U26179 ( .A(n25714), .B(n25715), .Z(n25713) );
  NAND U26180 ( .A(n25715), .B(n25714), .Z(n25710) );
  ANDN U26181 ( .B(A[6]), .A(n12), .Z(n25615) );
  XNOR U26182 ( .A(n25623), .B(n25716), .Z(n25616) );
  XNOR U26183 ( .A(n25622), .B(n25620), .Z(n25716) );
  AND U26184 ( .A(n25717), .B(n25718), .Z(n25620) );
  NANDN U26185 ( .A(n25719), .B(n25720), .Z(n25718) );
  NANDN U26186 ( .A(n25721), .B(n25722), .Z(n25720) );
  ANDN U26187 ( .B(A[5]), .A(n10), .Z(n25622) );
  XNOR U26188 ( .A(n25630), .B(n25723), .Z(n25623) );
  XNOR U26189 ( .A(n25629), .B(n25627), .Z(n25723) );
  AND U26190 ( .A(n25724), .B(n25725), .Z(n25627) );
  NANDN U26191 ( .A(n25726), .B(n25727), .Z(n25725) );
  OR U26192 ( .A(n25728), .B(n25729), .Z(n25727) );
  NAND U26193 ( .A(n25729), .B(n25728), .Z(n25724) );
  ANDN U26194 ( .B(A[4]), .A(n8), .Z(n25629) );
  XNOR U26195 ( .A(n25637), .B(n25730), .Z(n25630) );
  XNOR U26196 ( .A(n25636), .B(n25634), .Z(n25730) );
  AND U26197 ( .A(n25731), .B(n25732), .Z(n25634) );
  NANDN U26198 ( .A(n25733), .B(n25734), .Z(n25732) );
  NANDN U26199 ( .A(n25735), .B(n25736), .Z(n25734) );
  NANDN U26200 ( .A(n25736), .B(n25735), .Z(n25731) );
  ANDN U26201 ( .B(B[98]), .A(n41), .Z(n25636) );
  XOR U26202 ( .A(n25643), .B(n25737), .Z(n25637) );
  XNOR U26203 ( .A(n25641), .B(n25644), .Z(n25737) );
  NAND U26204 ( .A(B[99]), .B(A[2]), .Z(n25644) );
  NANDN U26205 ( .A(n25738), .B(n25739), .Z(n25641) );
  AND U26206 ( .A(A[0]), .B(B[100]), .Z(n25739) );
  XNOR U26207 ( .A(n25646), .B(n25740), .Z(n25643) );
  NAND U26208 ( .A(A[0]), .B(B[101]), .Z(n25740) );
  NAND U26209 ( .A(B[100]), .B(A[1]), .Z(n25646) );
  AND U26210 ( .A(n25741), .B(n25742), .Z(n25652) );
  NANDN U26211 ( .A(n575), .B(n25743), .Z(n25742) );
  NAND U26212 ( .A(n576), .B(n573), .Z(n25743) );
  NAND U26213 ( .A(A[14]), .B(B[86]), .Z(n575) );
  AND U26214 ( .A(n25744), .B(n25745), .Z(n576) );
  NANDN U26215 ( .A(n599), .B(n25746), .Z(n25745) );
  NANDN U26216 ( .A(n597), .B(n25747), .Z(n25746) );
  NAND U26217 ( .A(A[13]), .B(B[86]), .Z(n599) );
  NAND U26218 ( .A(n6), .B(n597), .Z(n25744) );
  XOR U26219 ( .A(n25748), .B(n25749), .Z(n597) );
  XNOR U26220 ( .A(n25750), .B(n25751), .Z(n25749) );
  AND U26221 ( .A(n25752), .B(n25753), .Z(n25747) );
  NANDN U26222 ( .A(n629), .B(n25754), .Z(n25753) );
  NANDN U26223 ( .A(n627), .B(n25755), .Z(n25754) );
  NAND U26224 ( .A(A[12]), .B(B[86]), .Z(n629) );
  NAND U26225 ( .A(n7), .B(n627), .Z(n25752) );
  XOR U26226 ( .A(n25756), .B(n25757), .Z(n627) );
  XNOR U26227 ( .A(n25758), .B(n25759), .Z(n25757) );
  AND U26228 ( .A(n25760), .B(n25761), .Z(n25755) );
  NANDN U26229 ( .A(n666), .B(n25762), .Z(n25761) );
  NANDN U26230 ( .A(n664), .B(n25763), .Z(n25762) );
  NAND U26231 ( .A(A[11]), .B(B[86]), .Z(n666) );
  NAND U26232 ( .A(n9), .B(n664), .Z(n25760) );
  XOR U26233 ( .A(n25764), .B(n25765), .Z(n664) );
  XNOR U26234 ( .A(n25766), .B(n25767), .Z(n25765) );
  AND U26235 ( .A(n25768), .B(n25769), .Z(n25763) );
  NANDN U26236 ( .A(n710), .B(n25770), .Z(n25769) );
  NANDN U26237 ( .A(n708), .B(n25771), .Z(n25770) );
  NAND U26238 ( .A(A[10]), .B(B[86]), .Z(n710) );
  NAND U26239 ( .A(n11), .B(n708), .Z(n25768) );
  XOR U26240 ( .A(n25772), .B(n25773), .Z(n708) );
  XNOR U26241 ( .A(n25774), .B(n25775), .Z(n25773) );
  AND U26242 ( .A(n25776), .B(n25777), .Z(n25771) );
  NANDN U26243 ( .A(n761), .B(n25778), .Z(n25777) );
  NANDN U26244 ( .A(n759), .B(n25779), .Z(n25778) );
  NAND U26245 ( .A(A[9]), .B(B[86]), .Z(n761) );
  NAND U26246 ( .A(n13), .B(n759), .Z(n25776) );
  XOR U26247 ( .A(n25780), .B(n25781), .Z(n759) );
  XNOR U26248 ( .A(n25782), .B(n25783), .Z(n25781) );
  AND U26249 ( .A(n25784), .B(n25785), .Z(n25779) );
  NANDN U26250 ( .A(n819), .B(n25786), .Z(n25785) );
  NANDN U26251 ( .A(n817), .B(n25787), .Z(n25786) );
  NAND U26252 ( .A(A[8]), .B(B[86]), .Z(n819) );
  NAND U26253 ( .A(n15), .B(n817), .Z(n25784) );
  XOR U26254 ( .A(n25788), .B(n25789), .Z(n817) );
  XNOR U26255 ( .A(n25790), .B(n25791), .Z(n25789) );
  AND U26256 ( .A(n25792), .B(n25793), .Z(n25787) );
  NANDN U26257 ( .A(n884), .B(n25794), .Z(n25793) );
  NANDN U26258 ( .A(n882), .B(n25795), .Z(n25794) );
  NAND U26259 ( .A(A[7]), .B(B[86]), .Z(n884) );
  NAND U26260 ( .A(n17), .B(n882), .Z(n25792) );
  XOR U26261 ( .A(n25796), .B(n25797), .Z(n882) );
  XNOR U26262 ( .A(n25798), .B(n25799), .Z(n25797) );
  AND U26263 ( .A(n25800), .B(n25801), .Z(n25795) );
  NANDN U26264 ( .A(n956), .B(n25802), .Z(n25801) );
  NANDN U26265 ( .A(n954), .B(n25803), .Z(n25802) );
  NAND U26266 ( .A(A[6]), .B(B[86]), .Z(n956) );
  NAND U26267 ( .A(n18), .B(n954), .Z(n25800) );
  XOR U26268 ( .A(n25804), .B(n25805), .Z(n954) );
  XNOR U26269 ( .A(n25806), .B(n25807), .Z(n25805) );
  AND U26270 ( .A(n25808), .B(n25809), .Z(n25803) );
  NANDN U26271 ( .A(n1039), .B(n25810), .Z(n25809) );
  NANDN U26272 ( .A(n1037), .B(n25811), .Z(n25810) );
  NAND U26273 ( .A(A[5]), .B(B[86]), .Z(n1039) );
  NAND U26274 ( .A(n19), .B(n1037), .Z(n25808) );
  XOR U26275 ( .A(n25812), .B(n25813), .Z(n1037) );
  XNOR U26276 ( .A(n25814), .B(n25815), .Z(n25813) );
  AND U26277 ( .A(n25816), .B(n25817), .Z(n25811) );
  NANDN U26278 ( .A(n1125), .B(n25818), .Z(n25817) );
  NANDN U26279 ( .A(n1123), .B(n25819), .Z(n25818) );
  NAND U26280 ( .A(A[4]), .B(B[86]), .Z(n1125) );
  NAND U26281 ( .A(n20), .B(n1123), .Z(n25816) );
  XOR U26282 ( .A(n25820), .B(n25821), .Z(n1123) );
  XNOR U26283 ( .A(n25822), .B(n25823), .Z(n25821) );
  AND U26284 ( .A(n25824), .B(n25825), .Z(n25819) );
  NANDN U26285 ( .A(n1218), .B(n25826), .Z(n25825) );
  NAND U26286 ( .A(n25827), .B(n1216), .Z(n25826) );
  NAND U26287 ( .A(A[3]), .B(B[86]), .Z(n1218) );
  NANDN U26288 ( .A(n1216), .B(n22), .Z(n25824) );
  AND U26289 ( .A(n25828), .B(n25829), .Z(n25827) );
  NANDN U26290 ( .A(n1318), .B(n25830), .Z(n25829) );
  NANDN U26291 ( .A(n1319), .B(n1316), .Z(n25830) );
  NAND U26292 ( .A(B[86]), .B(A[2]), .Z(n1318) );
  ANDN U26293 ( .B(n25831), .A(n1420), .Z(n1319) );
  NAND U26294 ( .A(B[86]), .B(A[1]), .Z(n1420) );
  AND U26295 ( .A(A[0]), .B(B[87]), .Z(n25831) );
  XNOR U26296 ( .A(n25832), .B(n25833), .Z(n1316) );
  NAND U26297 ( .A(B[88]), .B(A[0]), .Z(n25833) );
  XOR U26298 ( .A(n21), .B(n25834), .Z(n1216) );
  XNOR U26299 ( .A(n25835), .B(n25836), .Z(n25834) );
  XNOR U26300 ( .A(n25659), .B(n25837), .Z(n573) );
  XNOR U26301 ( .A(n25658), .B(n25656), .Z(n25837) );
  AND U26302 ( .A(n25838), .B(n25839), .Z(n25656) );
  NANDN U26303 ( .A(n25751), .B(n25840), .Z(n25839) );
  AND U26304 ( .A(n25841), .B(n25842), .Z(n25751) );
  NANDN U26305 ( .A(n25759), .B(n25843), .Z(n25842) );
  OR U26306 ( .A(n25758), .B(n25756), .Z(n25843) );
  AND U26307 ( .A(n25844), .B(n25845), .Z(n25759) );
  NANDN U26308 ( .A(n25767), .B(n25846), .Z(n25845) );
  AND U26309 ( .A(n25847), .B(n25848), .Z(n25767) );
  NANDN U26310 ( .A(n25775), .B(n25849), .Z(n25848) );
  OR U26311 ( .A(n25774), .B(n25772), .Z(n25849) );
  AND U26312 ( .A(n25850), .B(n25851), .Z(n25775) );
  NANDN U26313 ( .A(n25783), .B(n25852), .Z(n25851) );
  AND U26314 ( .A(n25853), .B(n25854), .Z(n25783) );
  NANDN U26315 ( .A(n25791), .B(n25855), .Z(n25854) );
  OR U26316 ( .A(n25790), .B(n25788), .Z(n25855) );
  AND U26317 ( .A(n25856), .B(n25857), .Z(n25791) );
  NANDN U26318 ( .A(n25799), .B(n25858), .Z(n25857) );
  AND U26319 ( .A(n25859), .B(n25860), .Z(n25799) );
  NANDN U26320 ( .A(n25807), .B(n25861), .Z(n25860) );
  OR U26321 ( .A(n25806), .B(n25804), .Z(n25861) );
  AND U26322 ( .A(n25862), .B(n25863), .Z(n25807) );
  NANDN U26323 ( .A(n25815), .B(n25864), .Z(n25863) );
  AND U26324 ( .A(n25865), .B(n25866), .Z(n25815) );
  NANDN U26325 ( .A(n25823), .B(n25867), .Z(n25866) );
  OR U26326 ( .A(n25822), .B(n25820), .Z(n25867) );
  AND U26327 ( .A(n25868), .B(n25869), .Z(n25823) );
  NANDN U26328 ( .A(n25835), .B(n25870), .Z(n25869) );
  NAND U26329 ( .A(n25871), .B(n25836), .Z(n25870) );
  NANDN U26330 ( .A(n25832), .B(n25872), .Z(n25835) );
  AND U26331 ( .A(A[0]), .B(B[88]), .Z(n25872) );
  NAND U26332 ( .A(B[87]), .B(A[1]), .Z(n25832) );
  NANDN U26333 ( .A(n25836), .B(n21), .Z(n25868) );
  XNOR U26334 ( .A(n25873), .B(n25874), .Z(n25871) );
  NAND U26335 ( .A(B[89]), .B(A[0]), .Z(n25874) );
  NAND U26336 ( .A(B[87]), .B(A[2]), .Z(n25836) );
  NAND U26337 ( .A(n25820), .B(n25822), .Z(n25865) );
  ANDN U26338 ( .B(B[87]), .A(n41), .Z(n25822) );
  XOR U26339 ( .A(n25875), .B(n25876), .Z(n25820) );
  XNOR U26340 ( .A(n25877), .B(n25878), .Z(n25876) );
  NAND U26341 ( .A(n25812), .B(n25814), .Z(n25862) );
  ANDN U26342 ( .B(B[87]), .A(n40), .Z(n25814) );
  XOR U26343 ( .A(n25879), .B(n25880), .Z(n25812) );
  XNOR U26344 ( .A(n25881), .B(n25882), .Z(n25880) );
  NAND U26345 ( .A(n25804), .B(n25806), .Z(n25859) );
  ANDN U26346 ( .B(B[87]), .A(n39), .Z(n25806) );
  XNOR U26347 ( .A(n25883), .B(n25884), .Z(n25804) );
  XNOR U26348 ( .A(n25885), .B(n25886), .Z(n25884) );
  NAND U26349 ( .A(n25796), .B(n25798), .Z(n25856) );
  ANDN U26350 ( .B(B[87]), .A(n38), .Z(n25798) );
  XOR U26351 ( .A(n25887), .B(n25888), .Z(n25796) );
  XNOR U26352 ( .A(n25889), .B(n25890), .Z(n25888) );
  NAND U26353 ( .A(n25788), .B(n25790), .Z(n25853) );
  ANDN U26354 ( .B(B[87]), .A(n37), .Z(n25790) );
  XNOR U26355 ( .A(n25891), .B(n25892), .Z(n25788) );
  XNOR U26356 ( .A(n25893), .B(n25894), .Z(n25892) );
  NAND U26357 ( .A(n25780), .B(n25782), .Z(n25850) );
  ANDN U26358 ( .B(B[87]), .A(n36), .Z(n25782) );
  XOR U26359 ( .A(n25895), .B(n25896), .Z(n25780) );
  XNOR U26360 ( .A(n25897), .B(n25898), .Z(n25896) );
  NAND U26361 ( .A(n25772), .B(n25774), .Z(n25847) );
  ANDN U26362 ( .B(B[87]), .A(n35), .Z(n25774) );
  XNOR U26363 ( .A(n25899), .B(n25900), .Z(n25772) );
  XNOR U26364 ( .A(n25901), .B(n25902), .Z(n25900) );
  NAND U26365 ( .A(n25764), .B(n25766), .Z(n25844) );
  ANDN U26366 ( .B(B[87]), .A(n34), .Z(n25766) );
  XOR U26367 ( .A(n25903), .B(n25904), .Z(n25764) );
  XNOR U26368 ( .A(n25905), .B(n25906), .Z(n25904) );
  NAND U26369 ( .A(n25756), .B(n25758), .Z(n25841) );
  ANDN U26370 ( .B(B[87]), .A(n33), .Z(n25758) );
  XNOR U26371 ( .A(n25907), .B(n25908), .Z(n25756) );
  XNOR U26372 ( .A(n25909), .B(n25910), .Z(n25908) );
  NAND U26373 ( .A(n25748), .B(n25750), .Z(n25838) );
  ANDN U26374 ( .B(B[87]), .A(n32), .Z(n25750) );
  XOR U26375 ( .A(n25911), .B(n25912), .Z(n25748) );
  XNOR U26376 ( .A(n25913), .B(n25914), .Z(n25912) );
  ANDN U26377 ( .B(B[87]), .A(n31), .Z(n25658) );
  XNOR U26378 ( .A(n25666), .B(n25915), .Z(n25659) );
  XNOR U26379 ( .A(n25665), .B(n25663), .Z(n25915) );
  AND U26380 ( .A(n25916), .B(n25917), .Z(n25663) );
  NANDN U26381 ( .A(n25914), .B(n25918), .Z(n25917) );
  OR U26382 ( .A(n25913), .B(n25911), .Z(n25918) );
  AND U26383 ( .A(n25919), .B(n25920), .Z(n25914) );
  NANDN U26384 ( .A(n25910), .B(n25921), .Z(n25920) );
  NANDN U26385 ( .A(n25909), .B(n25907), .Z(n25921) );
  AND U26386 ( .A(n25922), .B(n25923), .Z(n25910) );
  NANDN U26387 ( .A(n25906), .B(n25924), .Z(n25923) );
  OR U26388 ( .A(n25905), .B(n25903), .Z(n25924) );
  AND U26389 ( .A(n25925), .B(n25926), .Z(n25906) );
  NANDN U26390 ( .A(n25902), .B(n25927), .Z(n25926) );
  NANDN U26391 ( .A(n25901), .B(n25899), .Z(n25927) );
  AND U26392 ( .A(n25928), .B(n25929), .Z(n25902) );
  NANDN U26393 ( .A(n25898), .B(n25930), .Z(n25929) );
  OR U26394 ( .A(n25897), .B(n25895), .Z(n25930) );
  AND U26395 ( .A(n25931), .B(n25932), .Z(n25898) );
  NANDN U26396 ( .A(n25894), .B(n25933), .Z(n25932) );
  NANDN U26397 ( .A(n25893), .B(n25891), .Z(n25933) );
  AND U26398 ( .A(n25934), .B(n25935), .Z(n25894) );
  NANDN U26399 ( .A(n25890), .B(n25936), .Z(n25935) );
  OR U26400 ( .A(n25889), .B(n25887), .Z(n25936) );
  AND U26401 ( .A(n25937), .B(n25938), .Z(n25890) );
  NANDN U26402 ( .A(n25886), .B(n25939), .Z(n25938) );
  NANDN U26403 ( .A(n25885), .B(n25883), .Z(n25939) );
  AND U26404 ( .A(n25940), .B(n25941), .Z(n25886) );
  NANDN U26405 ( .A(n25882), .B(n25942), .Z(n25941) );
  OR U26406 ( .A(n25881), .B(n25879), .Z(n25942) );
  AND U26407 ( .A(n25943), .B(n25944), .Z(n25882) );
  NANDN U26408 ( .A(n25877), .B(n25945), .Z(n25944) );
  NAND U26409 ( .A(n25875), .B(n25878), .Z(n25945) );
  NANDN U26410 ( .A(n25873), .B(n25946), .Z(n25877) );
  AND U26411 ( .A(A[0]), .B(B[89]), .Z(n25946) );
  NAND U26412 ( .A(B[88]), .B(A[1]), .Z(n25873) );
  XNOR U26413 ( .A(n25947), .B(n25948), .Z(n25875) );
  NAND U26414 ( .A(B[90]), .B(A[0]), .Z(n25948) );
  NAND U26415 ( .A(B[88]), .B(A[2]), .Z(n25878) );
  NAND U26416 ( .A(n25879), .B(n25881), .Z(n25940) );
  ANDN U26417 ( .B(B[88]), .A(n41), .Z(n25881) );
  XOR U26418 ( .A(n25949), .B(n25950), .Z(n25879) );
  XNOR U26419 ( .A(n25951), .B(n25952), .Z(n25950) );
  NANDN U26420 ( .A(n25883), .B(n25885), .Z(n25937) );
  ANDN U26421 ( .B(B[88]), .A(n40), .Z(n25885) );
  XNOR U26422 ( .A(n25953), .B(n25954), .Z(n25883) );
  XNOR U26423 ( .A(n25955), .B(n25956), .Z(n25954) );
  NAND U26424 ( .A(n25887), .B(n25889), .Z(n25934) );
  ANDN U26425 ( .B(B[88]), .A(n39), .Z(n25889) );
  XNOR U26426 ( .A(n25957), .B(n25958), .Z(n25887) );
  XNOR U26427 ( .A(n25959), .B(n25960), .Z(n25958) );
  NANDN U26428 ( .A(n25891), .B(n25893), .Z(n25931) );
  ANDN U26429 ( .B(B[88]), .A(n38), .Z(n25893) );
  XNOR U26430 ( .A(n25961), .B(n25962), .Z(n25891) );
  XNOR U26431 ( .A(n25963), .B(n25964), .Z(n25962) );
  NAND U26432 ( .A(n25895), .B(n25897), .Z(n25928) );
  ANDN U26433 ( .B(B[88]), .A(n37), .Z(n25897) );
  XNOR U26434 ( .A(n25965), .B(n25966), .Z(n25895) );
  XNOR U26435 ( .A(n25967), .B(n25968), .Z(n25966) );
  NANDN U26436 ( .A(n25899), .B(n25901), .Z(n25925) );
  ANDN U26437 ( .B(B[88]), .A(n36), .Z(n25901) );
  XNOR U26438 ( .A(n25969), .B(n25970), .Z(n25899) );
  XNOR U26439 ( .A(n25971), .B(n25972), .Z(n25970) );
  NAND U26440 ( .A(n25903), .B(n25905), .Z(n25922) );
  ANDN U26441 ( .B(B[88]), .A(n35), .Z(n25905) );
  XNOR U26442 ( .A(n25973), .B(n25974), .Z(n25903) );
  XNOR U26443 ( .A(n25975), .B(n25976), .Z(n25974) );
  NANDN U26444 ( .A(n25907), .B(n25909), .Z(n25919) );
  ANDN U26445 ( .B(B[88]), .A(n34), .Z(n25909) );
  XNOR U26446 ( .A(n25977), .B(n25978), .Z(n25907) );
  XNOR U26447 ( .A(n25979), .B(n25980), .Z(n25978) );
  NAND U26448 ( .A(n25911), .B(n25913), .Z(n25916) );
  ANDN U26449 ( .B(B[88]), .A(n33), .Z(n25913) );
  XNOR U26450 ( .A(n25981), .B(n25982), .Z(n25911) );
  XNOR U26451 ( .A(n25983), .B(n25984), .Z(n25982) );
  ANDN U26452 ( .B(B[88]), .A(n32), .Z(n25665) );
  XNOR U26453 ( .A(n25673), .B(n25985), .Z(n25666) );
  XNOR U26454 ( .A(n25672), .B(n25670), .Z(n25985) );
  AND U26455 ( .A(n25986), .B(n25987), .Z(n25670) );
  NANDN U26456 ( .A(n25984), .B(n25988), .Z(n25987) );
  NANDN U26457 ( .A(n25983), .B(n25981), .Z(n25988) );
  AND U26458 ( .A(n25989), .B(n25990), .Z(n25984) );
  NANDN U26459 ( .A(n25980), .B(n25991), .Z(n25990) );
  OR U26460 ( .A(n25979), .B(n25977), .Z(n25991) );
  AND U26461 ( .A(n25992), .B(n25993), .Z(n25980) );
  NANDN U26462 ( .A(n25976), .B(n25994), .Z(n25993) );
  NANDN U26463 ( .A(n25975), .B(n25973), .Z(n25994) );
  AND U26464 ( .A(n25995), .B(n25996), .Z(n25976) );
  NANDN U26465 ( .A(n25972), .B(n25997), .Z(n25996) );
  OR U26466 ( .A(n25971), .B(n25969), .Z(n25997) );
  AND U26467 ( .A(n25998), .B(n25999), .Z(n25972) );
  NANDN U26468 ( .A(n25968), .B(n26000), .Z(n25999) );
  NANDN U26469 ( .A(n25967), .B(n25965), .Z(n26000) );
  AND U26470 ( .A(n26001), .B(n26002), .Z(n25968) );
  NANDN U26471 ( .A(n25964), .B(n26003), .Z(n26002) );
  OR U26472 ( .A(n25963), .B(n25961), .Z(n26003) );
  AND U26473 ( .A(n26004), .B(n26005), .Z(n25964) );
  NANDN U26474 ( .A(n25960), .B(n26006), .Z(n26005) );
  NANDN U26475 ( .A(n25959), .B(n25957), .Z(n26006) );
  AND U26476 ( .A(n26007), .B(n26008), .Z(n25960) );
  NANDN U26477 ( .A(n25956), .B(n26009), .Z(n26008) );
  OR U26478 ( .A(n25955), .B(n25953), .Z(n26009) );
  AND U26479 ( .A(n26010), .B(n26011), .Z(n25956) );
  NANDN U26480 ( .A(n25951), .B(n26012), .Z(n26011) );
  NAND U26481 ( .A(n25949), .B(n25952), .Z(n26012) );
  NANDN U26482 ( .A(n25947), .B(n26013), .Z(n25951) );
  AND U26483 ( .A(A[0]), .B(B[90]), .Z(n26013) );
  NAND U26484 ( .A(B[89]), .B(A[1]), .Z(n25947) );
  XNOR U26485 ( .A(n26014), .B(n26015), .Z(n25949) );
  NAND U26486 ( .A(B[91]), .B(A[0]), .Z(n26015) );
  NAND U26487 ( .A(B[89]), .B(A[2]), .Z(n25952) );
  NAND U26488 ( .A(n25953), .B(n25955), .Z(n26007) );
  ANDN U26489 ( .B(B[89]), .A(n41), .Z(n25955) );
  XOR U26490 ( .A(n26016), .B(n26017), .Z(n25953) );
  XNOR U26491 ( .A(n26018), .B(n26019), .Z(n26017) );
  NANDN U26492 ( .A(n25957), .B(n25959), .Z(n26004) );
  ANDN U26493 ( .B(B[89]), .A(n40), .Z(n25959) );
  XNOR U26494 ( .A(n26020), .B(n26021), .Z(n25957) );
  XNOR U26495 ( .A(n26022), .B(n26023), .Z(n26021) );
  NAND U26496 ( .A(n25961), .B(n25963), .Z(n26001) );
  ANDN U26497 ( .B(B[89]), .A(n39), .Z(n25963) );
  XNOR U26498 ( .A(n26024), .B(n26025), .Z(n25961) );
  XNOR U26499 ( .A(n26026), .B(n26027), .Z(n26025) );
  NANDN U26500 ( .A(n25965), .B(n25967), .Z(n25998) );
  ANDN U26501 ( .B(B[89]), .A(n38), .Z(n25967) );
  XNOR U26502 ( .A(n26028), .B(n26029), .Z(n25965) );
  XNOR U26503 ( .A(n26030), .B(n26031), .Z(n26029) );
  NAND U26504 ( .A(n25969), .B(n25971), .Z(n25995) );
  ANDN U26505 ( .B(B[89]), .A(n37), .Z(n25971) );
  XNOR U26506 ( .A(n26032), .B(n26033), .Z(n25969) );
  XNOR U26507 ( .A(n26034), .B(n26035), .Z(n26033) );
  NANDN U26508 ( .A(n25973), .B(n25975), .Z(n25992) );
  ANDN U26509 ( .B(B[89]), .A(n36), .Z(n25975) );
  XNOR U26510 ( .A(n26036), .B(n26037), .Z(n25973) );
  XNOR U26511 ( .A(n26038), .B(n26039), .Z(n26037) );
  NAND U26512 ( .A(n25977), .B(n25979), .Z(n25989) );
  ANDN U26513 ( .B(B[89]), .A(n35), .Z(n25979) );
  XNOR U26514 ( .A(n26040), .B(n26041), .Z(n25977) );
  XNOR U26515 ( .A(n26042), .B(n26043), .Z(n26041) );
  NANDN U26516 ( .A(n25981), .B(n25983), .Z(n25986) );
  ANDN U26517 ( .B(B[89]), .A(n34), .Z(n25983) );
  XNOR U26518 ( .A(n26044), .B(n26045), .Z(n25981) );
  XNOR U26519 ( .A(n26046), .B(n26047), .Z(n26045) );
  ANDN U26520 ( .B(B[89]), .A(n33), .Z(n25672) );
  XNOR U26521 ( .A(n25680), .B(n26048), .Z(n25673) );
  XNOR U26522 ( .A(n25679), .B(n25677), .Z(n26048) );
  AND U26523 ( .A(n26049), .B(n26050), .Z(n25677) );
  NANDN U26524 ( .A(n26047), .B(n26051), .Z(n26050) );
  OR U26525 ( .A(n26046), .B(n26044), .Z(n26051) );
  AND U26526 ( .A(n26052), .B(n26053), .Z(n26047) );
  NANDN U26527 ( .A(n26043), .B(n26054), .Z(n26053) );
  NANDN U26528 ( .A(n26042), .B(n26040), .Z(n26054) );
  AND U26529 ( .A(n26055), .B(n26056), .Z(n26043) );
  NANDN U26530 ( .A(n26039), .B(n26057), .Z(n26056) );
  OR U26531 ( .A(n26038), .B(n26036), .Z(n26057) );
  AND U26532 ( .A(n26058), .B(n26059), .Z(n26039) );
  NANDN U26533 ( .A(n26035), .B(n26060), .Z(n26059) );
  NANDN U26534 ( .A(n26034), .B(n26032), .Z(n26060) );
  AND U26535 ( .A(n26061), .B(n26062), .Z(n26035) );
  NANDN U26536 ( .A(n26031), .B(n26063), .Z(n26062) );
  OR U26537 ( .A(n26030), .B(n26028), .Z(n26063) );
  AND U26538 ( .A(n26064), .B(n26065), .Z(n26031) );
  NANDN U26539 ( .A(n26027), .B(n26066), .Z(n26065) );
  NANDN U26540 ( .A(n26026), .B(n26024), .Z(n26066) );
  AND U26541 ( .A(n26067), .B(n26068), .Z(n26027) );
  NANDN U26542 ( .A(n26023), .B(n26069), .Z(n26068) );
  OR U26543 ( .A(n26022), .B(n26020), .Z(n26069) );
  AND U26544 ( .A(n26070), .B(n26071), .Z(n26023) );
  NANDN U26545 ( .A(n26018), .B(n26072), .Z(n26071) );
  NAND U26546 ( .A(n26016), .B(n26019), .Z(n26072) );
  NANDN U26547 ( .A(n26014), .B(n26073), .Z(n26018) );
  AND U26548 ( .A(A[0]), .B(B[91]), .Z(n26073) );
  NAND U26549 ( .A(B[90]), .B(A[1]), .Z(n26014) );
  XNOR U26550 ( .A(n26074), .B(n26075), .Z(n26016) );
  NAND U26551 ( .A(B[92]), .B(A[0]), .Z(n26075) );
  NAND U26552 ( .A(B[90]), .B(A[2]), .Z(n26019) );
  NAND U26553 ( .A(n26020), .B(n26022), .Z(n26067) );
  ANDN U26554 ( .B(B[90]), .A(n41), .Z(n26022) );
  XOR U26555 ( .A(n26076), .B(n26077), .Z(n26020) );
  XNOR U26556 ( .A(n26078), .B(n26079), .Z(n26077) );
  NANDN U26557 ( .A(n26024), .B(n26026), .Z(n26064) );
  ANDN U26558 ( .B(B[90]), .A(n40), .Z(n26026) );
  XNOR U26559 ( .A(n26080), .B(n26081), .Z(n26024) );
  XNOR U26560 ( .A(n26082), .B(n26083), .Z(n26081) );
  NAND U26561 ( .A(n26028), .B(n26030), .Z(n26061) );
  ANDN U26562 ( .B(B[90]), .A(n39), .Z(n26030) );
  XNOR U26563 ( .A(n26084), .B(n26085), .Z(n26028) );
  XNOR U26564 ( .A(n26086), .B(n26087), .Z(n26085) );
  NANDN U26565 ( .A(n26032), .B(n26034), .Z(n26058) );
  ANDN U26566 ( .B(B[90]), .A(n38), .Z(n26034) );
  XNOR U26567 ( .A(n26088), .B(n26089), .Z(n26032) );
  XNOR U26568 ( .A(n26090), .B(n26091), .Z(n26089) );
  NAND U26569 ( .A(n26036), .B(n26038), .Z(n26055) );
  ANDN U26570 ( .B(B[90]), .A(n37), .Z(n26038) );
  XNOR U26571 ( .A(n26092), .B(n26093), .Z(n26036) );
  XNOR U26572 ( .A(n26094), .B(n26095), .Z(n26093) );
  NANDN U26573 ( .A(n26040), .B(n26042), .Z(n26052) );
  ANDN U26574 ( .B(B[90]), .A(n36), .Z(n26042) );
  XNOR U26575 ( .A(n26096), .B(n26097), .Z(n26040) );
  XNOR U26576 ( .A(n26098), .B(n26099), .Z(n26097) );
  NAND U26577 ( .A(n26044), .B(n26046), .Z(n26049) );
  ANDN U26578 ( .B(B[90]), .A(n35), .Z(n26046) );
  XNOR U26579 ( .A(n26100), .B(n26101), .Z(n26044) );
  XNOR U26580 ( .A(n26102), .B(n26103), .Z(n26101) );
  ANDN U26581 ( .B(B[90]), .A(n34), .Z(n25679) );
  XNOR U26582 ( .A(n25687), .B(n26104), .Z(n25680) );
  XNOR U26583 ( .A(n25686), .B(n25684), .Z(n26104) );
  AND U26584 ( .A(n26105), .B(n26106), .Z(n25684) );
  NANDN U26585 ( .A(n26103), .B(n26107), .Z(n26106) );
  NANDN U26586 ( .A(n26102), .B(n26100), .Z(n26107) );
  AND U26587 ( .A(n26108), .B(n26109), .Z(n26103) );
  NANDN U26588 ( .A(n26099), .B(n26110), .Z(n26109) );
  OR U26589 ( .A(n26098), .B(n26096), .Z(n26110) );
  AND U26590 ( .A(n26111), .B(n26112), .Z(n26099) );
  NANDN U26591 ( .A(n26095), .B(n26113), .Z(n26112) );
  NANDN U26592 ( .A(n26094), .B(n26092), .Z(n26113) );
  AND U26593 ( .A(n26114), .B(n26115), .Z(n26095) );
  NANDN U26594 ( .A(n26091), .B(n26116), .Z(n26115) );
  OR U26595 ( .A(n26090), .B(n26088), .Z(n26116) );
  AND U26596 ( .A(n26117), .B(n26118), .Z(n26091) );
  NANDN U26597 ( .A(n26087), .B(n26119), .Z(n26118) );
  NANDN U26598 ( .A(n26086), .B(n26084), .Z(n26119) );
  AND U26599 ( .A(n26120), .B(n26121), .Z(n26087) );
  NANDN U26600 ( .A(n26083), .B(n26122), .Z(n26121) );
  OR U26601 ( .A(n26082), .B(n26080), .Z(n26122) );
  AND U26602 ( .A(n26123), .B(n26124), .Z(n26083) );
  NANDN U26603 ( .A(n26078), .B(n26125), .Z(n26124) );
  NAND U26604 ( .A(n26076), .B(n26079), .Z(n26125) );
  NANDN U26605 ( .A(n26074), .B(n26126), .Z(n26078) );
  AND U26606 ( .A(A[0]), .B(B[92]), .Z(n26126) );
  NAND U26607 ( .A(B[91]), .B(A[1]), .Z(n26074) );
  XNOR U26608 ( .A(n26127), .B(n26128), .Z(n26076) );
  NAND U26609 ( .A(B[93]), .B(A[0]), .Z(n26128) );
  NAND U26610 ( .A(B[91]), .B(A[2]), .Z(n26079) );
  NAND U26611 ( .A(n26080), .B(n26082), .Z(n26120) );
  ANDN U26612 ( .B(B[91]), .A(n41), .Z(n26082) );
  XOR U26613 ( .A(n26129), .B(n26130), .Z(n26080) );
  XNOR U26614 ( .A(n26131), .B(n26132), .Z(n26130) );
  NANDN U26615 ( .A(n26084), .B(n26086), .Z(n26117) );
  ANDN U26616 ( .B(B[91]), .A(n40), .Z(n26086) );
  XNOR U26617 ( .A(n26133), .B(n26134), .Z(n26084) );
  XNOR U26618 ( .A(n26135), .B(n26136), .Z(n26134) );
  NAND U26619 ( .A(n26088), .B(n26090), .Z(n26114) );
  ANDN U26620 ( .B(B[91]), .A(n39), .Z(n26090) );
  XNOR U26621 ( .A(n26137), .B(n26138), .Z(n26088) );
  XNOR U26622 ( .A(n26139), .B(n26140), .Z(n26138) );
  NANDN U26623 ( .A(n26092), .B(n26094), .Z(n26111) );
  ANDN U26624 ( .B(B[91]), .A(n38), .Z(n26094) );
  XNOR U26625 ( .A(n26141), .B(n26142), .Z(n26092) );
  XNOR U26626 ( .A(n26143), .B(n26144), .Z(n26142) );
  NAND U26627 ( .A(n26096), .B(n26098), .Z(n26108) );
  ANDN U26628 ( .B(B[91]), .A(n37), .Z(n26098) );
  XNOR U26629 ( .A(n26145), .B(n26146), .Z(n26096) );
  XNOR U26630 ( .A(n26147), .B(n26148), .Z(n26146) );
  NANDN U26631 ( .A(n26100), .B(n26102), .Z(n26105) );
  ANDN U26632 ( .B(B[91]), .A(n36), .Z(n26102) );
  XNOR U26633 ( .A(n26149), .B(n26150), .Z(n26100) );
  XNOR U26634 ( .A(n26151), .B(n26152), .Z(n26150) );
  ANDN U26635 ( .B(B[91]), .A(n35), .Z(n25686) );
  XNOR U26636 ( .A(n25694), .B(n26153), .Z(n25687) );
  XNOR U26637 ( .A(n25693), .B(n25691), .Z(n26153) );
  AND U26638 ( .A(n26154), .B(n26155), .Z(n25691) );
  NANDN U26639 ( .A(n26152), .B(n26156), .Z(n26155) );
  OR U26640 ( .A(n26151), .B(n26149), .Z(n26156) );
  AND U26641 ( .A(n26157), .B(n26158), .Z(n26152) );
  NANDN U26642 ( .A(n26148), .B(n26159), .Z(n26158) );
  NANDN U26643 ( .A(n26147), .B(n26145), .Z(n26159) );
  AND U26644 ( .A(n26160), .B(n26161), .Z(n26148) );
  NANDN U26645 ( .A(n26144), .B(n26162), .Z(n26161) );
  OR U26646 ( .A(n26143), .B(n26141), .Z(n26162) );
  AND U26647 ( .A(n26163), .B(n26164), .Z(n26144) );
  NANDN U26648 ( .A(n26140), .B(n26165), .Z(n26164) );
  NANDN U26649 ( .A(n26139), .B(n26137), .Z(n26165) );
  AND U26650 ( .A(n26166), .B(n26167), .Z(n26140) );
  NANDN U26651 ( .A(n26136), .B(n26168), .Z(n26167) );
  OR U26652 ( .A(n26135), .B(n26133), .Z(n26168) );
  AND U26653 ( .A(n26169), .B(n26170), .Z(n26136) );
  NANDN U26654 ( .A(n26131), .B(n26171), .Z(n26170) );
  NAND U26655 ( .A(n26129), .B(n26132), .Z(n26171) );
  NANDN U26656 ( .A(n26127), .B(n26172), .Z(n26131) );
  AND U26657 ( .A(A[0]), .B(B[93]), .Z(n26172) );
  NAND U26658 ( .A(B[92]), .B(A[1]), .Z(n26127) );
  XNOR U26659 ( .A(n26173), .B(n26174), .Z(n26129) );
  NAND U26660 ( .A(B[94]), .B(A[0]), .Z(n26174) );
  NAND U26661 ( .A(B[92]), .B(A[2]), .Z(n26132) );
  NAND U26662 ( .A(n26133), .B(n26135), .Z(n26166) );
  ANDN U26663 ( .B(B[92]), .A(n41), .Z(n26135) );
  XOR U26664 ( .A(n26175), .B(n26176), .Z(n26133) );
  XNOR U26665 ( .A(n26177), .B(n26178), .Z(n26176) );
  NANDN U26666 ( .A(n26137), .B(n26139), .Z(n26163) );
  ANDN U26667 ( .B(B[92]), .A(n40), .Z(n26139) );
  XNOR U26668 ( .A(n26179), .B(n26180), .Z(n26137) );
  XNOR U26669 ( .A(n26181), .B(n26182), .Z(n26180) );
  NAND U26670 ( .A(n26141), .B(n26143), .Z(n26160) );
  ANDN U26671 ( .B(B[92]), .A(n39), .Z(n26143) );
  XNOR U26672 ( .A(n26183), .B(n26184), .Z(n26141) );
  XNOR U26673 ( .A(n26185), .B(n26186), .Z(n26184) );
  NANDN U26674 ( .A(n26145), .B(n26147), .Z(n26157) );
  ANDN U26675 ( .B(B[92]), .A(n38), .Z(n26147) );
  XNOR U26676 ( .A(n26187), .B(n26188), .Z(n26145) );
  XNOR U26677 ( .A(n26189), .B(n26190), .Z(n26188) );
  NAND U26678 ( .A(n26149), .B(n26151), .Z(n26154) );
  ANDN U26679 ( .B(B[92]), .A(n37), .Z(n26151) );
  XNOR U26680 ( .A(n26191), .B(n26192), .Z(n26149) );
  XNOR U26681 ( .A(n26193), .B(n26194), .Z(n26192) );
  ANDN U26682 ( .B(B[92]), .A(n36), .Z(n25693) );
  XNOR U26683 ( .A(n25701), .B(n26195), .Z(n25694) );
  XNOR U26684 ( .A(n25700), .B(n25698), .Z(n26195) );
  AND U26685 ( .A(n26196), .B(n26197), .Z(n25698) );
  NANDN U26686 ( .A(n26194), .B(n26198), .Z(n26197) );
  NANDN U26687 ( .A(n26193), .B(n26191), .Z(n26198) );
  AND U26688 ( .A(n26199), .B(n26200), .Z(n26194) );
  NANDN U26689 ( .A(n26190), .B(n26201), .Z(n26200) );
  OR U26690 ( .A(n26189), .B(n26187), .Z(n26201) );
  AND U26691 ( .A(n26202), .B(n26203), .Z(n26190) );
  NANDN U26692 ( .A(n26186), .B(n26204), .Z(n26203) );
  NANDN U26693 ( .A(n26185), .B(n26183), .Z(n26204) );
  AND U26694 ( .A(n26205), .B(n26206), .Z(n26186) );
  NANDN U26695 ( .A(n26182), .B(n26207), .Z(n26206) );
  OR U26696 ( .A(n26181), .B(n26179), .Z(n26207) );
  AND U26697 ( .A(n26208), .B(n26209), .Z(n26182) );
  NANDN U26698 ( .A(n26177), .B(n26210), .Z(n26209) );
  NAND U26699 ( .A(n26175), .B(n26178), .Z(n26210) );
  NANDN U26700 ( .A(n26173), .B(n26211), .Z(n26177) );
  AND U26701 ( .A(A[0]), .B(B[94]), .Z(n26211) );
  NAND U26702 ( .A(B[93]), .B(A[1]), .Z(n26173) );
  XNOR U26703 ( .A(n26212), .B(n26213), .Z(n26175) );
  NAND U26704 ( .A(B[95]), .B(A[0]), .Z(n26213) );
  NAND U26705 ( .A(B[93]), .B(A[2]), .Z(n26178) );
  NAND U26706 ( .A(n26179), .B(n26181), .Z(n26205) );
  ANDN U26707 ( .B(A[3]), .A(n16), .Z(n26181) );
  XOR U26708 ( .A(n26214), .B(n26215), .Z(n26179) );
  XNOR U26709 ( .A(n26216), .B(n26217), .Z(n26215) );
  NANDN U26710 ( .A(n26183), .B(n26185), .Z(n26202) );
  ANDN U26711 ( .B(A[4]), .A(n16), .Z(n26185) );
  XNOR U26712 ( .A(n26218), .B(n26219), .Z(n26183) );
  XNOR U26713 ( .A(n26220), .B(n26221), .Z(n26219) );
  NAND U26714 ( .A(n26187), .B(n26189), .Z(n26199) );
  ANDN U26715 ( .B(A[5]), .A(n16), .Z(n26189) );
  XNOR U26716 ( .A(n26222), .B(n26223), .Z(n26187) );
  XNOR U26717 ( .A(n26224), .B(n26225), .Z(n26223) );
  NANDN U26718 ( .A(n26191), .B(n26193), .Z(n26196) );
  ANDN U26719 ( .B(A[6]), .A(n16), .Z(n26193) );
  XNOR U26720 ( .A(n26226), .B(n26227), .Z(n26191) );
  XNOR U26721 ( .A(n26228), .B(n26229), .Z(n26227) );
  ANDN U26722 ( .B(A[7]), .A(n16), .Z(n25700) );
  XNOR U26723 ( .A(n25708), .B(n26230), .Z(n25701) );
  XNOR U26724 ( .A(n25707), .B(n25705), .Z(n26230) );
  AND U26725 ( .A(n26231), .B(n26232), .Z(n25705) );
  NANDN U26726 ( .A(n26229), .B(n26233), .Z(n26232) );
  OR U26727 ( .A(n26228), .B(n26226), .Z(n26233) );
  AND U26728 ( .A(n26234), .B(n26235), .Z(n26229) );
  NANDN U26729 ( .A(n26225), .B(n26236), .Z(n26235) );
  NANDN U26730 ( .A(n26224), .B(n26222), .Z(n26236) );
  AND U26731 ( .A(n26237), .B(n26238), .Z(n26225) );
  NANDN U26732 ( .A(n26221), .B(n26239), .Z(n26238) );
  OR U26733 ( .A(n26220), .B(n26218), .Z(n26239) );
  AND U26734 ( .A(n26240), .B(n26241), .Z(n26221) );
  NANDN U26735 ( .A(n26216), .B(n26242), .Z(n26241) );
  NAND U26736 ( .A(n26214), .B(n26217), .Z(n26242) );
  NANDN U26737 ( .A(n26212), .B(n26243), .Z(n26216) );
  AND U26738 ( .A(A[0]), .B(B[95]), .Z(n26243) );
  NAND U26739 ( .A(B[94]), .B(A[1]), .Z(n26212) );
  XNOR U26740 ( .A(n26244), .B(n26245), .Z(n26214) );
  NAND U26741 ( .A(B[96]), .B(A[0]), .Z(n26245) );
  NAND U26742 ( .A(B[94]), .B(A[2]), .Z(n26217) );
  NAND U26743 ( .A(n26218), .B(n26220), .Z(n26237) );
  ANDN U26744 ( .B(A[3]), .A(n14), .Z(n26220) );
  XOR U26745 ( .A(n26246), .B(n26247), .Z(n26218) );
  XNOR U26746 ( .A(n26248), .B(n26249), .Z(n26247) );
  NANDN U26747 ( .A(n26222), .B(n26224), .Z(n26234) );
  ANDN U26748 ( .B(A[4]), .A(n14), .Z(n26224) );
  XNOR U26749 ( .A(n26250), .B(n26251), .Z(n26222) );
  XNOR U26750 ( .A(n26252), .B(n26253), .Z(n26251) );
  NAND U26751 ( .A(n26226), .B(n26228), .Z(n26231) );
  ANDN U26752 ( .B(A[5]), .A(n14), .Z(n26228) );
  XNOR U26753 ( .A(n26254), .B(n26255), .Z(n26226) );
  XNOR U26754 ( .A(n26256), .B(n26257), .Z(n26255) );
  ANDN U26755 ( .B(A[6]), .A(n14), .Z(n25707) );
  XNOR U26756 ( .A(n25715), .B(n26258), .Z(n25708) );
  XNOR U26757 ( .A(n25714), .B(n25712), .Z(n26258) );
  AND U26758 ( .A(n26259), .B(n26260), .Z(n25712) );
  NANDN U26759 ( .A(n26257), .B(n26261), .Z(n26260) );
  NANDN U26760 ( .A(n26256), .B(n26254), .Z(n26261) );
  AND U26761 ( .A(n26262), .B(n26263), .Z(n26257) );
  NANDN U26762 ( .A(n26253), .B(n26264), .Z(n26263) );
  OR U26763 ( .A(n26252), .B(n26250), .Z(n26264) );
  AND U26764 ( .A(n26265), .B(n26266), .Z(n26253) );
  NANDN U26765 ( .A(n26248), .B(n26267), .Z(n26266) );
  NAND U26766 ( .A(n26246), .B(n26249), .Z(n26267) );
  NANDN U26767 ( .A(n26244), .B(n26268), .Z(n26248) );
  AND U26768 ( .A(A[0]), .B(B[96]), .Z(n26268) );
  NAND U26769 ( .A(B[95]), .B(A[1]), .Z(n26244) );
  XNOR U26770 ( .A(n26269), .B(n26270), .Z(n26246) );
  NAND U26771 ( .A(B[97]), .B(A[0]), .Z(n26270) );
  NAND U26772 ( .A(B[95]), .B(A[2]), .Z(n26249) );
  NAND U26773 ( .A(n26250), .B(n26252), .Z(n26262) );
  ANDN U26774 ( .B(A[3]), .A(n12), .Z(n26252) );
  XOR U26775 ( .A(n26271), .B(n26272), .Z(n26250) );
  XNOR U26776 ( .A(n26273), .B(n26274), .Z(n26272) );
  NANDN U26777 ( .A(n26254), .B(n26256), .Z(n26259) );
  ANDN U26778 ( .B(A[4]), .A(n12), .Z(n26256) );
  XNOR U26779 ( .A(n26275), .B(n26276), .Z(n26254) );
  XNOR U26780 ( .A(n26277), .B(n26278), .Z(n26276) );
  ANDN U26781 ( .B(A[5]), .A(n12), .Z(n25714) );
  XNOR U26782 ( .A(n25722), .B(n26279), .Z(n25715) );
  XNOR U26783 ( .A(n25721), .B(n25719), .Z(n26279) );
  AND U26784 ( .A(n26280), .B(n26281), .Z(n25719) );
  NANDN U26785 ( .A(n26278), .B(n26282), .Z(n26281) );
  OR U26786 ( .A(n26277), .B(n26275), .Z(n26282) );
  AND U26787 ( .A(n26283), .B(n26284), .Z(n26278) );
  NANDN U26788 ( .A(n26273), .B(n26285), .Z(n26284) );
  NAND U26789 ( .A(n26271), .B(n26274), .Z(n26285) );
  NANDN U26790 ( .A(n26269), .B(n26286), .Z(n26273) );
  AND U26791 ( .A(A[0]), .B(B[97]), .Z(n26286) );
  NAND U26792 ( .A(B[96]), .B(A[1]), .Z(n26269) );
  XNOR U26793 ( .A(n26287), .B(n26288), .Z(n26271) );
  NAND U26794 ( .A(B[98]), .B(A[0]), .Z(n26288) );
  NAND U26795 ( .A(B[96]), .B(A[2]), .Z(n26274) );
  NAND U26796 ( .A(n26275), .B(n26277), .Z(n26280) );
  ANDN U26797 ( .B(A[3]), .A(n10), .Z(n26277) );
  XOR U26798 ( .A(n26289), .B(n26290), .Z(n26275) );
  XNOR U26799 ( .A(n26291), .B(n26292), .Z(n26290) );
  ANDN U26800 ( .B(A[4]), .A(n10), .Z(n25721) );
  XNOR U26801 ( .A(n25729), .B(n26293), .Z(n25722) );
  XNOR U26802 ( .A(n25728), .B(n25726), .Z(n26293) );
  AND U26803 ( .A(n26294), .B(n26295), .Z(n25726) );
  NANDN U26804 ( .A(n26291), .B(n26296), .Z(n26295) );
  NAND U26805 ( .A(n26289), .B(n26292), .Z(n26296) );
  NANDN U26806 ( .A(n26287), .B(n26297), .Z(n26291) );
  AND U26807 ( .A(A[0]), .B(B[98]), .Z(n26297) );
  NAND U26808 ( .A(B[97]), .B(A[1]), .Z(n26287) );
  XNOR U26809 ( .A(n26298), .B(n26299), .Z(n26289) );
  NAND U26810 ( .A(B[99]), .B(A[0]), .Z(n26299) );
  NAND U26811 ( .A(B[97]), .B(A[2]), .Z(n26292) );
  ANDN U26812 ( .B(A[3]), .A(n8), .Z(n25728) );
  XNOR U26813 ( .A(n25735), .B(n26300), .Z(n25729) );
  XNOR U26814 ( .A(n25733), .B(n25736), .Z(n26300) );
  NAND U26815 ( .A(B[98]), .B(A[2]), .Z(n25736) );
  NANDN U26816 ( .A(n26298), .B(n26301), .Z(n25733) );
  AND U26817 ( .A(A[0]), .B(B[99]), .Z(n26301) );
  NAND U26818 ( .A(B[98]), .B(A[1]), .Z(n26298) );
  XOR U26819 ( .A(n25738), .B(n26302), .Z(n25735) );
  NAND U26820 ( .A(B[100]), .B(A[0]), .Z(n26302) );
  NAND U26821 ( .A(B[99]), .B(A[1]), .Z(n25738) );
  XNOR U26822 ( .A(n24321), .B(n26303), .Z(\A1[0] ) );
  XNOR U26823 ( .A(n24318), .B(n24320), .Z(n26303) );
  ANDN U26824 ( .B(n44), .A(n43), .Z(n24320) );
  NAND U26825 ( .A(B[0]), .B(A[1]), .Z(n43) );
  AND U26826 ( .A(A[0]), .B(B[1]), .Z(n44) );
  NAND U26827 ( .A(B[0]), .B(A[2]), .Z(n24318) );
  XNOR U26828 ( .A(n24354), .B(n26304), .Z(n24321) );
  NAND U26829 ( .A(A[0]), .B(B[2]), .Z(n26304) );
  NAND U26830 ( .A(B[1]), .B(A[1]), .Z(n24354) );
endmodule


module mult_N256_CC16 ( clk, rst, a, b, c );
  input [255:0] a;
  input [15:0] b;
  output [255:0] c;
  input clk, rst;

  wire   [255:16] swire;
  wire   [511:256] sreg;
  wire   [255:0] clocal;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;

  DFF \sreg_reg[256]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[257]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[258]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[259]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[260]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[261]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[262]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[263]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[264]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[265]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[266]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[267]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[268]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[269]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[270]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[271]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[272]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[273]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[274]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[275]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[276]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[277]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[278]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[279]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[280]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[281]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[282]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[283]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[284]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[285]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[286]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[287]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[288]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[289]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[290]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[291]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[292]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[293]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[294]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[295]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[296]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[297]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[298]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[299]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[300]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[301]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[302]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[303]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[304]  ( .D(swire[64]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[305]  ( .D(swire[65]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[306]  ( .D(swire[66]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[307]  ( .D(swire[67]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[308]  ( .D(swire[68]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[309]  ( .D(swire[69]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[310]  ( .D(swire[70]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[311]  ( .D(swire[71]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[312]  ( .D(swire[72]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[313]  ( .D(swire[73]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[314]  ( .D(swire[74]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[315]  ( .D(swire[75]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[316]  ( .D(swire[76]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[317]  ( .D(swire[77]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[318]  ( .D(swire[78]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[319]  ( .D(swire[79]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[320]  ( .D(swire[80]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[321]  ( .D(swire[81]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[322]  ( .D(swire[82]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[323]  ( .D(swire[83]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[324]  ( .D(swire[84]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[325]  ( .D(swire[85]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[326]  ( .D(swire[86]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[327]  ( .D(swire[87]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[328]  ( .D(swire[88]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[329]  ( .D(swire[89]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[330]  ( .D(swire[90]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[331]  ( .D(swire[91]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[332]  ( .D(swire[92]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[333]  ( .D(swire[93]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[334]  ( .D(swire[94]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[335]  ( .D(swire[95]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[336]  ( .D(swire[96]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[337]  ( .D(swire[97]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[338]  ( .D(swire[98]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[339]  ( .D(swire[99]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[340]  ( .D(swire[100]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[341]  ( .D(swire[101]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[342]  ( .D(swire[102]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[343]  ( .D(swire[103]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[344]  ( .D(swire[104]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[345]  ( .D(swire[105]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[346]  ( .D(swire[106]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[347]  ( .D(swire[107]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[348]  ( .D(swire[108]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[349]  ( .D(swire[109]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[350]  ( .D(swire[110]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[351]  ( .D(swire[111]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[352]  ( .D(swire[112]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[353]  ( .D(swire[113]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[354]  ( .D(swire[114]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[355]  ( .D(swire[115]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[356]  ( .D(swire[116]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[357]  ( .D(swire[117]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[358]  ( .D(swire[118]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[359]  ( .D(swire[119]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[360]  ( .D(swire[120]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[361]  ( .D(swire[121]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[362]  ( .D(swire[122]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[363]  ( .D(swire[123]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[364]  ( .D(swire[124]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[365]  ( .D(swire[125]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[366]  ( .D(swire[126]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[367]  ( .D(swire[127]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[368]  ( .D(swire[128]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[369]  ( .D(swire[129]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[370]  ( .D(swire[130]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[371]  ( .D(swire[131]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[372]  ( .D(swire[132]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[373]  ( .D(swire[133]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[374]  ( .D(swire[134]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[375]  ( .D(swire[135]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[376]  ( .D(swire[136]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[377]  ( .D(swire[137]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[378]  ( .D(swire[138]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[379]  ( .D(swire[139]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[380]  ( .D(swire[140]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[381]  ( .D(swire[141]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[382]  ( .D(swire[142]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[383]  ( .D(swire[143]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[384]  ( .D(swire[144]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[385]  ( .D(swire[145]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[386]  ( .D(swire[146]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[387]  ( .D(swire[147]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[388]  ( .D(swire[148]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[389]  ( .D(swire[149]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[390]  ( .D(swire[150]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[391]  ( .D(swire[151]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[392]  ( .D(swire[152]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[393]  ( .D(swire[153]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[394]  ( .D(swire[154]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[395]  ( .D(swire[155]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[396]  ( .D(swire[156]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[397]  ( .D(swire[157]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[398]  ( .D(swire[158]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[399]  ( .D(swire[159]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[400]  ( .D(swire[160]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[401]  ( .D(swire[161]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[402]  ( .D(swire[162]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[403]  ( .D(swire[163]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[404]  ( .D(swire[164]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[405]  ( .D(swire[165]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[406]  ( .D(swire[166]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[407]  ( .D(swire[167]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[408]  ( .D(swire[168]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[409]  ( .D(swire[169]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[410]  ( .D(swire[170]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[411]  ( .D(swire[171]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[412]  ( .D(swire[172]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[413]  ( .D(swire[173]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[414]  ( .D(swire[174]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[415]  ( .D(swire[175]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[416]  ( .D(swire[176]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[417]  ( .D(swire[177]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[418]  ( .D(swire[178]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[419]  ( .D(swire[179]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[420]  ( .D(swire[180]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[421]  ( .D(swire[181]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[422]  ( .D(swire[182]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[423]  ( .D(swire[183]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[424]  ( .D(swire[184]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[425]  ( .D(swire[185]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[426]  ( .D(swire[186]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[427]  ( .D(swire[187]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[428]  ( .D(swire[188]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[429]  ( .D(swire[189]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[430]  ( .D(swire[190]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[431]  ( .D(swire[191]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[432]  ( .D(swire[192]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[433]  ( .D(swire[193]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[434]  ( .D(swire[194]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[435]  ( .D(swire[195]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[436]  ( .D(swire[196]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[437]  ( .D(swire[197]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[438]  ( .D(swire[198]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[439]  ( .D(swire[199]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[440]  ( .D(swire[200]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[441]  ( .D(swire[201]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[442]  ( .D(swire[202]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[443]  ( .D(swire[203]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[444]  ( .D(swire[204]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[445]  ( .D(swire[205]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[446]  ( .D(swire[206]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[447]  ( .D(swire[207]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[448]  ( .D(swire[208]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[449]  ( .D(swire[209]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[450]  ( .D(swire[210]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[451]  ( .D(swire[211]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[452]  ( .D(swire[212]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[453]  ( .D(swire[213]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[454]  ( .D(swire[214]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[455]  ( .D(swire[215]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[456]  ( .D(swire[216]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[457]  ( .D(swire[217]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[458]  ( .D(swire[218]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[459]  ( .D(swire[219]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[460]  ( .D(swire[220]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[461]  ( .D(swire[221]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[462]  ( .D(swire[222]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[463]  ( .D(swire[223]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[464]  ( .D(swire[224]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[465]  ( .D(swire[225]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[466]  ( .D(swire[226]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[467]  ( .D(swire[227]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[468]  ( .D(swire[228]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[469]  ( .D(swire[229]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[470]  ( .D(swire[230]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[471]  ( .D(swire[231]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[472]  ( .D(swire[232]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[473]  ( .D(swire[233]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[474]  ( .D(swire[234]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[475]  ( .D(swire[235]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[476]  ( .D(swire[236]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[477]  ( .D(swire[237]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[478]  ( .D(swire[238]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[479]  ( .D(swire[239]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[480]  ( .D(swire[240]), .CLK(clk), .RST(rst), .Q(sreg[480]) );
  DFF \sreg_reg[481]  ( .D(swire[241]), .CLK(clk), .RST(rst), .Q(sreg[481]) );
  DFF \sreg_reg[482]  ( .D(swire[242]), .CLK(clk), .RST(rst), .Q(sreg[482]) );
  DFF \sreg_reg[483]  ( .D(swire[243]), .CLK(clk), .RST(rst), .Q(sreg[483]) );
  DFF \sreg_reg[484]  ( .D(swire[244]), .CLK(clk), .RST(rst), .Q(sreg[484]) );
  DFF \sreg_reg[485]  ( .D(swire[245]), .CLK(clk), .RST(rst), .Q(sreg[485]) );
  DFF \sreg_reg[486]  ( .D(swire[246]), .CLK(clk), .RST(rst), .Q(sreg[486]) );
  DFF \sreg_reg[487]  ( .D(swire[247]), .CLK(clk), .RST(rst), .Q(sreg[487]) );
  DFF \sreg_reg[488]  ( .D(swire[248]), .CLK(clk), .RST(rst), .Q(sreg[488]) );
  DFF \sreg_reg[489]  ( .D(swire[249]), .CLK(clk), .RST(rst), .Q(sreg[489]) );
  DFF \sreg_reg[490]  ( .D(swire[250]), .CLK(clk), .RST(rst), .Q(sreg[490]) );
  DFF \sreg_reg[491]  ( .D(swire[251]), .CLK(clk), .RST(rst), .Q(sreg[491]) );
  DFF \sreg_reg[492]  ( .D(swire[252]), .CLK(clk), .RST(rst), .Q(sreg[492]) );
  DFF \sreg_reg[493]  ( .D(swire[253]), .CLK(clk), .RST(rst), .Q(sreg[493]) );
  DFF \sreg_reg[494]  ( .D(swire[254]), .CLK(clk), .RST(rst), .Q(sreg[494]) );
  DFF \sreg_reg[495]  ( .D(swire[255]), .CLK(clk), .RST(rst), .Q(sreg[495]) );
  DFF \sreg_reg[255]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[239]) );
  DFF \sreg_reg[254]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[238]) );
  DFF \sreg_reg[253]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[237]) );
  DFF \sreg_reg[252]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[236]) );
  DFF \sreg_reg[251]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[235]) );
  DFF \sreg_reg[250]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[234]) );
  DFF \sreg_reg[249]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[233]) );
  DFF \sreg_reg[248]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[232]) );
  DFF \sreg_reg[247]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[231]) );
  DFF \sreg_reg[246]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[230]) );
  DFF \sreg_reg[245]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[229]) );
  DFF \sreg_reg[244]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[228]) );
  DFF \sreg_reg[243]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[227]) );
  DFF \sreg_reg[242]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[226]) );
  DFF \sreg_reg[241]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[225]) );
  DFF \sreg_reg[240]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[224]) );
  DFF \sreg_reg[239]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[238]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[237]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[236]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[235]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[234]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[233]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[232]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[231]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[230]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[229]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[228]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[227]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[226]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[225]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[224]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[223]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[222]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[221]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[220]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[219]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[218]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[217]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[216]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[215]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[214]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[213]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[212]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[211]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[210]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[209]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[208]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[207]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[206]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[205]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[204]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[203]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[202]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[201]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[200]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[199]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[198]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[197]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[196]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[195]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[194]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[193]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[192]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[191]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[190]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[189]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[188]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[187]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[186]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[185]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[184]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[183]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[182]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[181]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[180]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[179]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[178]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[177]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[176]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[175]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[174]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[173]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[172]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[171]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[170]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[169]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[168]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[167]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[166]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[165]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[164]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[163]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[162]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[161]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[160]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[159]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[158]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[157]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[156]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[155]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[154]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[153]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[152]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[151]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[150]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[149]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[148]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[147]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[146]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[145]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[144]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[143]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[142]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[141]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[140]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[139]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[138]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[137]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[136]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[135]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[134]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[133]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[132]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[131]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[130]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[129]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[128]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[0]) );
  ADD_N256 ADD_ ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, sreg[495:256]}), .B(clocal), 
        .CI(1'b0), .S({swire, c[255:240]}) );
  mult_N256_CC16_DW02_mult_0 mult_44 ( .A(b), .B(a), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, clocal}) );
endmodule

