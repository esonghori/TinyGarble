
module hamming_N16000_CC16_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49;

  XOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[8]) );
  XNOR U4 ( .A(B[8]), .B(A[8]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U14 ( .A(B[3]), .B(A[3]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U16 ( .A(B[2]), .B(A[2]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[1]) );
  XOR U18 ( .A(B[1]), .B(A[1]), .Z(n18) );
  XOR U19 ( .A(A[13]), .B(n19), .Z(SUM[13]) );
  ANDN U20 ( .B(A[12]), .A(n20), .Z(n19) );
  XNOR U21 ( .A(A[12]), .B(n20), .Z(SUM[12]) );
  NAND U22 ( .A(n21), .B(A[11]), .Z(n20) );
  XOR U23 ( .A(A[11]), .B(n21), .Z(SUM[11]) );
  ANDN U24 ( .B(A[10]), .A(n22), .Z(n21) );
  XNOR U25 ( .A(A[10]), .B(n22), .Z(SUM[10]) );
  AND U26 ( .A(n23), .B(n24), .Z(n22) );
  NAND U27 ( .A(n25), .B(B[9]), .Z(n24) );
  NANDN U28 ( .A(A[9]), .B(n1), .Z(n25) );
  NANDN U29 ( .A(n1), .B(A[9]), .Z(n23) );
  AND U30 ( .A(n26), .B(n27), .Z(n1) );
  NAND U31 ( .A(n28), .B(B[8]), .Z(n27) );
  NANDN U32 ( .A(A[8]), .B(n3), .Z(n28) );
  NANDN U33 ( .A(n3), .B(A[8]), .Z(n26) );
  AND U34 ( .A(n29), .B(n30), .Z(n3) );
  NAND U35 ( .A(n31), .B(B[7]), .Z(n30) );
  NANDN U36 ( .A(A[7]), .B(n5), .Z(n31) );
  NANDN U37 ( .A(n5), .B(A[7]), .Z(n29) );
  AND U38 ( .A(n32), .B(n33), .Z(n5) );
  NAND U39 ( .A(n34), .B(B[6]), .Z(n33) );
  NANDN U40 ( .A(A[6]), .B(n7), .Z(n34) );
  NANDN U41 ( .A(n7), .B(A[6]), .Z(n32) );
  AND U42 ( .A(n35), .B(n36), .Z(n7) );
  NAND U43 ( .A(n37), .B(B[5]), .Z(n36) );
  NANDN U44 ( .A(A[5]), .B(n9), .Z(n37) );
  NANDN U45 ( .A(n9), .B(A[5]), .Z(n35) );
  AND U46 ( .A(n38), .B(n39), .Z(n9) );
  NAND U47 ( .A(n40), .B(B[4]), .Z(n39) );
  NANDN U48 ( .A(A[4]), .B(n11), .Z(n40) );
  NANDN U49 ( .A(n11), .B(A[4]), .Z(n38) );
  AND U50 ( .A(n41), .B(n42), .Z(n11) );
  NAND U51 ( .A(n43), .B(B[3]), .Z(n42) );
  NANDN U52 ( .A(A[3]), .B(n13), .Z(n43) );
  NANDN U53 ( .A(n13), .B(A[3]), .Z(n41) );
  AND U54 ( .A(n44), .B(n45), .Z(n13) );
  NAND U55 ( .A(n46), .B(B[2]), .Z(n45) );
  NANDN U56 ( .A(A[2]), .B(n15), .Z(n46) );
  NANDN U57 ( .A(n15), .B(A[2]), .Z(n44) );
  AND U58 ( .A(n47), .B(n48), .Z(n15) );
  NAND U59 ( .A(n49), .B(B[1]), .Z(n48) );
  OR U60 ( .A(n17), .B(A[1]), .Z(n49) );
  NAND U61 ( .A(n17), .B(A[1]), .Z(n47) );
  AND U62 ( .A(B[0]), .B(A[0]), .Z(n17) );
  XOR U63 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_1 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42;

  IV U1 ( .A(B[9]), .Z(n1) );
  XOR U2 ( .A(n2), .B(n1), .Z(SUM[9]) );
  AND U3 ( .A(n3), .B(n4), .Z(n2) );
  NAND U4 ( .A(n5), .B(B[8]), .Z(n4) );
  NANDN U5 ( .A(A[8]), .B(n6), .Z(n5) );
  NANDN U6 ( .A(n6), .B(A[8]), .Z(n3) );
  XOR U7 ( .A(n6), .B(n7), .Z(SUM[8]) );
  XNOR U8 ( .A(B[8]), .B(A[8]), .Z(n7) );
  AND U9 ( .A(n8), .B(n9), .Z(n6) );
  NAND U10 ( .A(n10), .B(B[7]), .Z(n9) );
  NANDN U11 ( .A(A[7]), .B(n11), .Z(n10) );
  NANDN U12 ( .A(n11), .B(A[7]), .Z(n8) );
  XOR U13 ( .A(n11), .B(n12), .Z(SUM[7]) );
  XNOR U14 ( .A(B[7]), .B(A[7]), .Z(n12) );
  AND U15 ( .A(n13), .B(n14), .Z(n11) );
  NAND U16 ( .A(n15), .B(B[6]), .Z(n14) );
  NANDN U17 ( .A(A[6]), .B(n16), .Z(n15) );
  NANDN U18 ( .A(n16), .B(A[6]), .Z(n13) );
  XOR U19 ( .A(n16), .B(n17), .Z(SUM[6]) );
  XNOR U20 ( .A(B[6]), .B(A[6]), .Z(n17) );
  AND U21 ( .A(n18), .B(n19), .Z(n16) );
  NAND U22 ( .A(n20), .B(B[5]), .Z(n19) );
  NANDN U23 ( .A(A[5]), .B(n21), .Z(n20) );
  NANDN U24 ( .A(n21), .B(A[5]), .Z(n18) );
  XOR U25 ( .A(n21), .B(n22), .Z(SUM[5]) );
  XNOR U26 ( .A(B[5]), .B(A[5]), .Z(n22) );
  AND U27 ( .A(n23), .B(n24), .Z(n21) );
  NAND U28 ( .A(n25), .B(B[4]), .Z(n24) );
  NANDN U29 ( .A(A[4]), .B(n26), .Z(n25) );
  NANDN U30 ( .A(n26), .B(A[4]), .Z(n23) );
  XOR U31 ( .A(n26), .B(n27), .Z(SUM[4]) );
  XNOR U32 ( .A(B[4]), .B(A[4]), .Z(n27) );
  AND U33 ( .A(n28), .B(n29), .Z(n26) );
  NAND U34 ( .A(n30), .B(B[3]), .Z(n29) );
  NANDN U35 ( .A(A[3]), .B(n31), .Z(n30) );
  NANDN U36 ( .A(n31), .B(A[3]), .Z(n28) );
  XOR U37 ( .A(n31), .B(n32), .Z(SUM[3]) );
  XNOR U38 ( .A(B[3]), .B(A[3]), .Z(n32) );
  AND U39 ( .A(n33), .B(n34), .Z(n31) );
  NAND U40 ( .A(n35), .B(B[2]), .Z(n34) );
  NANDN U41 ( .A(A[2]), .B(n36), .Z(n35) );
  NANDN U42 ( .A(n36), .B(A[2]), .Z(n33) );
  XOR U43 ( .A(n36), .B(n37), .Z(SUM[2]) );
  XNOR U44 ( .A(B[2]), .B(A[2]), .Z(n37) );
  AND U45 ( .A(n38), .B(n39), .Z(n36) );
  NAND U46 ( .A(n40), .B(B[1]), .Z(n39) );
  OR U47 ( .A(n41), .B(A[1]), .Z(n40) );
  NAND U48 ( .A(n41), .B(A[1]), .Z(n38) );
  XOR U49 ( .A(n41), .B(n42), .Z(SUM[1]) );
  XOR U50 ( .A(B[1]), .B(A[1]), .Z(n42) );
  AND U51 ( .A(B[0]), .B(A[0]), .Z(n41) );
  XOR U52 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_2 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[9]) );
  NAND U2 ( .A(n4), .B(B[8]), .Z(n3) );
  NANDN U3 ( .A(A[8]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[8]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[8]) );
  XNOR U6 ( .A(B[8]), .B(A[8]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[7]), .Z(n8) );
  NANDN U9 ( .A(A[7]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[7]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[7]) );
  XNOR U12 ( .A(B[7]), .B(A[7]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[6]), .Z(n13) );
  NANDN U15 ( .A(A[6]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[6]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[6]) );
  XNOR U18 ( .A(B[6]), .B(A[6]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[5]), .Z(n18) );
  NANDN U21 ( .A(A[5]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[5]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[5]) );
  XNOR U24 ( .A(B[5]), .B(A[5]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[4]), .Z(n23) );
  NANDN U27 ( .A(A[4]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(n25), .B(A[4]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[4]) );
  XNOR U30 ( .A(B[4]), .B(A[4]), .Z(n26) );
  AND U31 ( .A(n27), .B(n28), .Z(n25) );
  NAND U32 ( .A(n29), .B(B[3]), .Z(n28) );
  NANDN U33 ( .A(A[3]), .B(n30), .Z(n29) );
  NANDN U34 ( .A(n30), .B(A[3]), .Z(n27) );
  XOR U35 ( .A(n30), .B(n31), .Z(SUM[3]) );
  XNOR U36 ( .A(B[3]), .B(A[3]), .Z(n31) );
  AND U37 ( .A(n32), .B(n33), .Z(n30) );
  NAND U38 ( .A(n34), .B(B[2]), .Z(n33) );
  NANDN U39 ( .A(A[2]), .B(n35), .Z(n34) );
  NANDN U40 ( .A(n35), .B(A[2]), .Z(n32) );
  XOR U41 ( .A(n35), .B(n36), .Z(SUM[2]) );
  XNOR U42 ( .A(B[2]), .B(A[2]), .Z(n36) );
  AND U43 ( .A(n37), .B(n38), .Z(n35) );
  NAND U44 ( .A(n39), .B(B[1]), .Z(n38) );
  OR U45 ( .A(n40), .B(A[1]), .Z(n39) );
  NAND U46 ( .A(n40), .B(A[1]), .Z(n37) );
  XOR U47 ( .A(n40), .B(n41), .Z(SUM[1]) );
  XOR U48 ( .A(B[1]), .B(A[1]), .Z(n41) );
  AND U49 ( .A(B[0]), .B(A[0]), .Z(n40) );
  XOR U50 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_3 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[8]) );
  NAND U2 ( .A(n4), .B(B[7]), .Z(n3) );
  NANDN U3 ( .A(A[7]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[7]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[6]), .Z(n8) );
  NANDN U9 ( .A(A[6]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[6]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[6]) );
  XNOR U12 ( .A(B[6]), .B(A[6]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U15 ( .A(A[5]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[5]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[5]) );
  XNOR U18 ( .A(B[5]), .B(A[5]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[4]), .Z(n18) );
  NANDN U21 ( .A(A[4]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[4]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[4]) );
  XNOR U24 ( .A(B[4]), .B(A[4]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[3]), .Z(n23) );
  NANDN U27 ( .A(A[3]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(n25), .B(A[3]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[3]) );
  XNOR U30 ( .A(B[3]), .B(A[3]), .Z(n26) );
  AND U31 ( .A(n27), .B(n28), .Z(n25) );
  NAND U32 ( .A(n29), .B(B[2]), .Z(n28) );
  NANDN U33 ( .A(A[2]), .B(n30), .Z(n29) );
  NANDN U34 ( .A(n30), .B(A[2]), .Z(n27) );
  XOR U35 ( .A(n30), .B(n31), .Z(SUM[2]) );
  XNOR U36 ( .A(B[2]), .B(A[2]), .Z(n31) );
  AND U37 ( .A(n32), .B(n33), .Z(n30) );
  NAND U38 ( .A(n34), .B(B[1]), .Z(n33) );
  OR U39 ( .A(n35), .B(A[1]), .Z(n34) );
  NAND U40 ( .A(n35), .B(A[1]), .Z(n32) );
  XOR U41 ( .A(n35), .B(n36), .Z(SUM[1]) );
  XOR U42 ( .A(B[1]), .B(A[1]), .Z(n36) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n35) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_4 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[8]) );
  NAND U2 ( .A(n4), .B(B[7]), .Z(n3) );
  NANDN U3 ( .A(A[7]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[7]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[7]) );
  XNOR U6 ( .A(B[7]), .B(A[7]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[6]), .Z(n8) );
  NANDN U9 ( .A(A[6]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[6]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[6]) );
  XNOR U12 ( .A(B[6]), .B(A[6]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[5]), .Z(n13) );
  NANDN U15 ( .A(A[5]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[5]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[5]) );
  XNOR U18 ( .A(B[5]), .B(A[5]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[4]), .Z(n18) );
  NANDN U21 ( .A(A[4]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[4]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[4]) );
  XNOR U24 ( .A(B[4]), .B(A[4]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[3]), .Z(n23) );
  NANDN U27 ( .A(A[3]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(n25), .B(A[3]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[3]) );
  XNOR U30 ( .A(B[3]), .B(A[3]), .Z(n26) );
  AND U31 ( .A(n27), .B(n28), .Z(n25) );
  NAND U32 ( .A(n29), .B(B[2]), .Z(n28) );
  NANDN U33 ( .A(A[2]), .B(n30), .Z(n29) );
  NANDN U34 ( .A(n30), .B(A[2]), .Z(n27) );
  XOR U35 ( .A(n30), .B(n31), .Z(SUM[2]) );
  XNOR U36 ( .A(B[2]), .B(A[2]), .Z(n31) );
  AND U37 ( .A(n32), .B(n33), .Z(n30) );
  NAND U38 ( .A(n34), .B(B[1]), .Z(n33) );
  OR U39 ( .A(n35), .B(A[1]), .Z(n34) );
  NAND U40 ( .A(n35), .B(A[1]), .Z(n32) );
  XOR U41 ( .A(n35), .B(n36), .Z(SUM[1]) );
  XOR U42 ( .A(B[1]), .B(A[1]), .Z(n36) );
  AND U43 ( .A(B[0]), .B(A[0]), .Z(n35) );
  XOR U44 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_5 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34;

  AND U1 ( .A(n3), .B(B[7]), .Z(SUM[8]) );
  IV U2 ( .A(B[7]), .Z(n2) );
  IV U3 ( .A(n4), .Z(n3) );
  XOR U4 ( .A(n4), .B(n2), .Z(SUM[7]) );
  AND U5 ( .A(n5), .B(n6), .Z(n4) );
  NAND U6 ( .A(n7), .B(B[6]), .Z(n6) );
  NANDN U7 ( .A(A[6]), .B(n8), .Z(n7) );
  NANDN U8 ( .A(n8), .B(A[6]), .Z(n5) );
  XOR U9 ( .A(n8), .B(n9), .Z(SUM[6]) );
  XNOR U10 ( .A(B[6]), .B(A[6]), .Z(n9) );
  AND U11 ( .A(n10), .B(n11), .Z(n8) );
  NAND U12 ( .A(n12), .B(B[5]), .Z(n11) );
  NANDN U13 ( .A(A[5]), .B(n13), .Z(n12) );
  NANDN U14 ( .A(n13), .B(A[5]), .Z(n10) );
  XOR U15 ( .A(n13), .B(n14), .Z(SUM[5]) );
  XNOR U16 ( .A(B[5]), .B(A[5]), .Z(n14) );
  AND U17 ( .A(n15), .B(n16), .Z(n13) );
  NAND U18 ( .A(n17), .B(B[4]), .Z(n16) );
  NANDN U19 ( .A(A[4]), .B(n18), .Z(n17) );
  NANDN U20 ( .A(n18), .B(A[4]), .Z(n15) );
  XOR U21 ( .A(n18), .B(n19), .Z(SUM[4]) );
  XNOR U22 ( .A(B[4]), .B(A[4]), .Z(n19) );
  AND U23 ( .A(n20), .B(n21), .Z(n18) );
  NAND U24 ( .A(n22), .B(B[3]), .Z(n21) );
  NANDN U25 ( .A(A[3]), .B(n23), .Z(n22) );
  NANDN U26 ( .A(n23), .B(A[3]), .Z(n20) );
  XOR U27 ( .A(n23), .B(n24), .Z(SUM[3]) );
  XNOR U28 ( .A(B[3]), .B(A[3]), .Z(n24) );
  AND U29 ( .A(n25), .B(n26), .Z(n23) );
  NAND U30 ( .A(n27), .B(B[2]), .Z(n26) );
  NANDN U31 ( .A(A[2]), .B(n28), .Z(n27) );
  NANDN U32 ( .A(n28), .B(A[2]), .Z(n25) );
  XOR U33 ( .A(n28), .B(n29), .Z(SUM[2]) );
  XNOR U34 ( .A(B[2]), .B(A[2]), .Z(n29) );
  AND U35 ( .A(n30), .B(n31), .Z(n28) );
  NAND U36 ( .A(n32), .B(B[1]), .Z(n31) );
  OR U37 ( .A(n33), .B(A[1]), .Z(n32) );
  NAND U38 ( .A(n33), .B(A[1]), .Z(n30) );
  XOR U39 ( .A(n33), .B(n34), .Z(SUM[1]) );
  XOR U40 ( .A(B[1]), .B(A[1]), .Z(n34) );
  AND U41 ( .A(B[0]), .B(A[0]), .Z(n33) );
  XOR U42 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_6 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[7]) );
  NAND U2 ( .A(n4), .B(B[6]), .Z(n3) );
  NANDN U3 ( .A(A[6]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[6]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[5]), .Z(n8) );
  NANDN U9 ( .A(A[5]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[5]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U12 ( .A(B[5]), .B(A[5]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[4]), .Z(n13) );
  NANDN U15 ( .A(A[4]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[4]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[4]) );
  XNOR U18 ( .A(B[4]), .B(A[4]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[3]), .Z(n18) );
  NANDN U21 ( .A(A[3]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[3]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[3]) );
  XNOR U24 ( .A(B[3]), .B(A[3]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[2]), .Z(n23) );
  NANDN U27 ( .A(A[2]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(n25), .B(A[2]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[2]) );
  XNOR U30 ( .A(B[2]), .B(A[2]), .Z(n26) );
  AND U31 ( .A(n27), .B(n28), .Z(n25) );
  NAND U32 ( .A(n29), .B(B[1]), .Z(n28) );
  OR U33 ( .A(n30), .B(A[1]), .Z(n29) );
  NAND U34 ( .A(n30), .B(A[1]), .Z(n27) );
  XOR U35 ( .A(n30), .B(n31), .Z(SUM[1]) );
  XOR U36 ( .A(B[1]), .B(A[1]), .Z(n31) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n30) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_7 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[7]) );
  NAND U2 ( .A(n4), .B(B[6]), .Z(n3) );
  NANDN U3 ( .A(A[6]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[6]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[5]), .Z(n8) );
  NANDN U9 ( .A(A[5]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[5]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U12 ( .A(B[5]), .B(A[5]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[4]), .Z(n13) );
  NANDN U15 ( .A(A[4]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[4]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[4]) );
  XNOR U18 ( .A(B[4]), .B(A[4]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[3]), .Z(n18) );
  NANDN U21 ( .A(A[3]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[3]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[3]) );
  XNOR U24 ( .A(B[3]), .B(A[3]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[2]), .Z(n23) );
  NANDN U27 ( .A(A[2]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(n25), .B(A[2]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[2]) );
  XNOR U30 ( .A(B[2]), .B(A[2]), .Z(n26) );
  AND U31 ( .A(n27), .B(n28), .Z(n25) );
  NAND U32 ( .A(n29), .B(B[1]), .Z(n28) );
  OR U33 ( .A(n30), .B(A[1]), .Z(n29) );
  NAND U34 ( .A(n30), .B(A[1]), .Z(n27) );
  XOR U35 ( .A(n30), .B(n31), .Z(SUM[1]) );
  XOR U36 ( .A(B[1]), .B(A[1]), .Z(n31) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n30) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_8 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[7]) );
  NAND U2 ( .A(n4), .B(B[6]), .Z(n3) );
  NANDN U3 ( .A(A[6]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[6]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[5]), .Z(n8) );
  NANDN U9 ( .A(A[5]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[5]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U12 ( .A(B[5]), .B(A[5]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[4]), .Z(n13) );
  NANDN U15 ( .A(A[4]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[4]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[4]) );
  XNOR U18 ( .A(B[4]), .B(A[4]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[3]), .Z(n18) );
  NANDN U21 ( .A(A[3]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[3]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[3]) );
  XNOR U24 ( .A(B[3]), .B(A[3]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[2]), .Z(n23) );
  NANDN U27 ( .A(A[2]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(n25), .B(A[2]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[2]) );
  XNOR U30 ( .A(B[2]), .B(A[2]), .Z(n26) );
  AND U31 ( .A(n27), .B(n28), .Z(n25) );
  NAND U32 ( .A(n29), .B(B[1]), .Z(n28) );
  OR U33 ( .A(n30), .B(A[1]), .Z(n29) );
  NAND U34 ( .A(n30), .B(A[1]), .Z(n27) );
  XOR U35 ( .A(n30), .B(n31), .Z(SUM[1]) );
  XOR U36 ( .A(B[1]), .B(A[1]), .Z(n31) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n30) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_9 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[7]) );
  NAND U2 ( .A(n4), .B(B[6]), .Z(n3) );
  NANDN U3 ( .A(A[6]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[6]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[5]), .Z(n8) );
  NANDN U9 ( .A(A[5]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[5]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U12 ( .A(B[5]), .B(A[5]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[4]), .Z(n13) );
  NANDN U15 ( .A(A[4]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[4]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[4]) );
  XNOR U18 ( .A(B[4]), .B(A[4]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[3]), .Z(n18) );
  NANDN U21 ( .A(A[3]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[3]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[3]) );
  XNOR U24 ( .A(B[3]), .B(A[3]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[2]), .Z(n23) );
  NANDN U27 ( .A(A[2]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(n25), .B(A[2]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[2]) );
  XNOR U30 ( .A(B[2]), .B(A[2]), .Z(n26) );
  AND U31 ( .A(n27), .B(n28), .Z(n25) );
  NAND U32 ( .A(n29), .B(B[1]), .Z(n28) );
  OR U33 ( .A(n30), .B(A[1]), .Z(n29) );
  NAND U34 ( .A(n30), .B(A[1]), .Z(n27) );
  XOR U35 ( .A(n30), .B(n31), .Z(SUM[1]) );
  XOR U36 ( .A(B[1]), .B(A[1]), .Z(n31) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n30) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_10 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29;

  AND U1 ( .A(n2), .B(B[6]), .Z(SUM[7]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[6]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[6]) );
  AND U5 ( .A(n5), .B(n6), .Z(n4) );
  NAND U6 ( .A(n7), .B(B[5]), .Z(n6) );
  NANDN U7 ( .A(A[5]), .B(n8), .Z(n7) );
  NANDN U8 ( .A(n8), .B(A[5]), .Z(n5) );
  XOR U9 ( .A(n8), .B(n9), .Z(SUM[5]) );
  XNOR U10 ( .A(B[5]), .B(A[5]), .Z(n9) );
  AND U11 ( .A(n10), .B(n11), .Z(n8) );
  NAND U12 ( .A(n12), .B(B[4]), .Z(n11) );
  NANDN U13 ( .A(A[4]), .B(n13), .Z(n12) );
  NANDN U14 ( .A(n13), .B(A[4]), .Z(n10) );
  XOR U15 ( .A(n13), .B(n14), .Z(SUM[4]) );
  XNOR U16 ( .A(B[4]), .B(A[4]), .Z(n14) );
  AND U17 ( .A(n15), .B(n16), .Z(n13) );
  NAND U18 ( .A(n17), .B(B[3]), .Z(n16) );
  NANDN U19 ( .A(A[3]), .B(n18), .Z(n17) );
  NANDN U20 ( .A(n18), .B(A[3]), .Z(n15) );
  XOR U21 ( .A(n18), .B(n19), .Z(SUM[3]) );
  XNOR U22 ( .A(B[3]), .B(A[3]), .Z(n19) );
  AND U23 ( .A(n20), .B(n21), .Z(n18) );
  NAND U24 ( .A(n22), .B(B[2]), .Z(n21) );
  NANDN U25 ( .A(A[2]), .B(n23), .Z(n22) );
  NANDN U26 ( .A(n23), .B(A[2]), .Z(n20) );
  XOR U27 ( .A(n23), .B(n24), .Z(SUM[2]) );
  XNOR U28 ( .A(B[2]), .B(A[2]), .Z(n24) );
  AND U29 ( .A(n25), .B(n26), .Z(n23) );
  NAND U30 ( .A(n27), .B(B[1]), .Z(n26) );
  OR U31 ( .A(n28), .B(A[1]), .Z(n27) );
  NAND U32 ( .A(n28), .B(A[1]), .Z(n25) );
  XOR U33 ( .A(n28), .B(n29), .Z(SUM[1]) );
  XOR U34 ( .A(B[1]), .B(A[1]), .Z(n29) );
  AND U35 ( .A(B[0]), .B(A[0]), .Z(n28) );
  XOR U36 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_11 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_12 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_13 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_14 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_15 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_16 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_17 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_18 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_19 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_20 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_21 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_22 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_23 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_24 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_25 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_26 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_27 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_28 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_29 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_30 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_31 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_32 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_33 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_34 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_35 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_36 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_37 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_38 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_39 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_40 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16_DW01_add_41 ( A, B, CI, SUM, CO );
  input [9:0] A;
  input [9:0] B;
  output [9:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC16 ( clk, rst, x, y, o );
  input [999:0] x;
  input [999:0] y;
  output [13:0] o;
  input clk, rst;
  wire   N5784, N5785, N5786, N5787, N5788, N5794, N5795, N5796, N5797, N5798,
         N5804, N5805, N5806, N5807, N5808, N5814, N5815, N5816, N5817, N5818,
         N5824, N5825, N5826, N5827, N5828, N5834, N5835, N5836, N5837, N5838,
         N5844, N5845, N5846, N5847, N5848, N5854, N5855, N5856, N5857, N5858,
         N5864, N5865, N5866, N5867, N5868, N5874, N5875, N5876, N5877, N5878,
         N5884, N5885, N5886, N5887, N5888, N5894, N5895, N5896, N5897, N5898,
         N5904, N5905, N5906, N5907, N5908, N5914, N5915, N5916, N5917, N5918,
         N5924, N5925, N5926, N5927, N5928, N5934, N5935, N5936, N5937, N5938,
         N5944, N5945, N5946, N5947, N5948, N5954, N5955, N5956, N5957, N5958,
         N5964, N5965, N5966, N5967, N5968, N5974, N5975, N5976, N5977, N5978,
         N5984, N5985, N5986, N5987, N5988, N5994, N5995, N5996, N5997, N5998,
         N6004, N6005, N6006, N6007, N6008, N6014, N6015, N6016, N6017, N6018,
         N6024, N6025, N6026, N6027, N6028, N6034, N6035, N6036, N6037, N6038,
         N6044, N6045, N6046, N6047, N6048, N6054, N6055, N6056, N6057, N6058,
         N6064, N6065, N6066, N6067, N6068, N6074, N6075, N6076, N6077, N6078,
         N6084, N6085, N6086, N6087, N6088, N6094, N6095, N6096, N6097, N6098,
         N6104, N6105, N6106, N6107, N6108, N6114, N6115, N6116, N6117, N6118,
         N6124, N6125, N6126, N6127, N6128, N6134, N6135, N6136, N6137, N6138,
         N6144, N6145, N6146, N6147, N6148, N6154, N6155, N6156, N6157, N6158,
         N6164, N6165, N6166, N6167, N6168, N6174, N6175, N6176, N6177, N6178,
         N6184, N6185, N6186, N6187, N6188, N6194, N6195, N6196, N6197, N6198,
         N6204, N6205, N6206, N6207, N6208, N6209, N6214, N6215, N6216, N6217,
         N6218, N6219, N6224, N6225, N6226, N6227, N6228, N6229, N6234, N6235,
         N6236, N6237, N6238, N6239, N6244, N6245, N6246, N6247, N6248, N6249,
         N6254, N6255, N6256, N6257, N6258, N6259, N6264, N6265, N6266, N6267,
         N6268, N6269, N6274, N6275, N6276, N6277, N6278, N6279, N6284, N6285,
         N6286, N6287, N6288, N6289, N6294, N6295, N6296, N6297, N6298, N6299,
         N6304, N6305, N6306, N6307, N6308, N6309, N6314, N6315, N6316, N6317,
         N6318, N6319, N6324, N6325, N6326, N6327, N6328, N6329, N6334, N6335,
         N6336, N6337, N6338, N6339, N6344, N6345, N6346, N6347, N6348, N6349,
         N6354, N6355, N6356, N6357, N6358, N6359, N6364, N6365, N6366, N6367,
         N6368, N6369, N6374, N6375, N6376, N6377, N6378, N6379, N6384, N6385,
         N6386, N6387, N6388, N6389, N6394, N6395, N6396, N6397, N6398, N6399,
         N6404, N6405, N6406, N6407, N6408, N6409, N6414, N6415, N6416, N6417,
         N6418, N6419, N6420, N6424, N6425, N6426, N6427, N6428, N6429, N6430,
         N6434, N6435, N6436, N6437, N6438, N6439, N6440, N6444, N6445, N6446,
         N6447, N6448, N6449, N6450, N6454, N6455, N6456, N6457, N6458, N6459,
         N6460, N6464, N6465, N6466, N6467, N6468, N6469, N6470, N6474, N6475,
         N6476, N6477, N6478, N6479, N6480, N6484, N6485, N6486, N6487, N6488,
         N6489, N6490, N6494, N6495, N6496, N6497, N6498, N6499, N6500, N6504,
         N6505, N6506, N6507, N6508, N6509, N6510, N6514, N6515, N6516, N6517,
         N6518, N6519, N6520, N6521, N6524, N6525, N6526, N6527, N6528, N6529,
         N6530, N6531, N6534, N6535, N6536, N6537, N6538, N6539, N6540, N6541,
         N6544, N6545, N6546, N6547, N6548, N6549, N6550, N6551, N6554, N6555,
         N6556, N6557, N6558, N6559, N6560, N6561, N6564, N6565, N6566, N6567,
         N6568, N6569, N6570, N6571, N6572, N6574, N6575, N6576, N6577, N6578,
         N6579, N6580, N6581, N6582, N6584, N6585, N6586, N6587, N6588, N6589,
         N6590, N6591, N6592, N6594, N6595, N6596, N6597, N6598, N6599, N6600,
         N6601, N6602, N6603, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798;
  wire   [9:0] olocal;
  wire   [13:0] oglobal;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  hamming_N16000_CC16_DW01_add_0 add_97 ( .A(oglobal), .B({1'b0, 1'b0, 1'b0, 
        1'b0, olocal}), .CI(1'b0), .SUM(o) );
  hamming_N16000_CC16_DW01_add_1 add_334_root_add_47_I1000 ( .A({1'b0, N6592, 
        N6591, N6590, N6589, N6588, N6587, N6586, N6585, N6584}), .B({N6603, 
        N6602, N6601, N6600, N6599, N6598, N6597, N6596, N6595, N6594}), .CI(
        1'b0), .SUM(olocal) );
  hamming_N16000_CC16_DW01_add_2 add_335_root_add_47_I1000 ( .A({1'b0, N6572, 
        N6571, N6570, N6569, N6568, N6567, N6566, N6565, N6564}), .B({1'b0, 
        N6582, N6581, N6580, N6579, N6578, N6577, N6576, N6575, N6574}), .CI(
        1'b0), .SUM({N6603, N6602, N6601, N6600, N6599, N6598, N6597, N6596, 
        N6595, N6594}) );
  hamming_N16000_CC16_DW01_add_3 add_336_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        N6551, N6550, N6549, N6548, N6547, N6546, N6545, N6544}), .B({1'b0, 
        1'b0, N6561, N6560, N6559, N6558, N6557, N6556, N6555, N6554}), .CI(
        1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, N6592, N6591, N6590, N6589, 
        N6588, N6587, N6586, N6585, N6584}) );
  hamming_N16000_CC16_DW01_add_4 add_337_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        N6531, N6530, N6529, N6528, N6527, N6526, N6525, N6524}), .B({1'b0, 
        1'b0, N6541, N6540, N6539, N6538, N6537, N6536, N6535, N6534}), .CI(
        1'b0), .SUM({SYNOPSYS_UNCONNECTED__1, N6582, N6581, N6580, N6579, 
        N6578, N6577, N6576, N6575, N6574}) );
  hamming_N16000_CC16_DW01_add_5 add_338_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, N6510, N6509, N6508, N6507, N6506, N6505, N6504}), .B({1'b0, 
        1'b0, N6521, N6520, N6519, N6518, N6517, N6516, N6515, N6514}), .CI(
        1'b0), .SUM({SYNOPSYS_UNCONNECTED__2, N6572, N6571, N6570, N6569, 
        N6568, N6567, N6566, N6565, N6564}) );
  hamming_N16000_CC16_DW01_add_6 add_339_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, N6490, N6489, N6488, N6487, N6486, N6485, N6484}), .B({1'b0, 
        1'b0, 1'b0, N6500, N6499, N6498, N6497, N6496, N6495, N6494}), .CI(
        1'b0), .SUM({SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, N6561, 
        N6560, N6559, N6558, N6557, N6556, N6555, N6554}) );
  hamming_N16000_CC16_DW01_add_7 add_340_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, N6470, N6469, N6468, N6467, N6466, N6465, N6464}), .B({1'b0, 
        1'b0, 1'b0, N6480, N6479, N6478, N6477, N6476, N6475, N6474}), .CI(
        1'b0), .SUM({SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, N6551, 
        N6550, N6549, N6548, N6547, N6546, N6545, N6544}) );
  hamming_N16000_CC16_DW01_add_8 add_341_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, N6450, N6449, N6448, N6447, N6446, N6445, N6444}), .B({1'b0, 
        1'b0, 1'b0, N6460, N6459, N6458, N6457, N6456, N6455, N6454}), .CI(
        1'b0), .SUM({SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, N6541, 
        N6540, N6539, N6538, N6537, N6536, N6535, N6534}) );
  hamming_N16000_CC16_DW01_add_9 add_342_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, N6430, N6429, N6428, N6427, N6426, N6425, N6424}), .B({1'b0, 
        1'b0, 1'b0, N6440, N6439, N6438, N6437, N6436, N6435, N6434}), .CI(
        1'b0), .SUM({SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, N6531, 
        N6530, N6529, N6528, N6527, N6526, N6525, N6524}) );
  hamming_N16000_CC16_DW01_add_10 add_343_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N6409, N6408, N6407, N6406, N6405, N6404}), .B({1'b0, 1'b0, 
        1'b0, N6420, N6419, N6418, N6417, N6416, N6415, N6414}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, N6521, N6520, 
        N6519, N6518, N6517, N6516, N6515, N6514}) );
  hamming_N16000_CC16_DW01_add_11 add_344_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N6389, N6388, N6387, N6386, N6385, N6384}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, N6399, N6398, N6397, N6396, N6395, N6394}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, N6510, N6509, N6508, N6507, N6506, N6505, 
        N6504}) );
  hamming_N16000_CC16_DW01_add_12 add_345_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N6369, N6368, N6367, N6366, N6365, N6364}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, N6379, N6378, N6377, N6376, N6375, N6374}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, N6500, N6499, N6498, N6497, N6496, N6495, 
        N6494}) );
  hamming_N16000_CC16_DW01_add_13 add_346_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N6349, N6348, N6347, N6346, N6345, N6344}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, N6359, N6358, N6357, N6356, N6355, N6354}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, N6490, N6489, N6488, N6487, N6486, N6485, 
        N6484}) );
  hamming_N16000_CC16_DW01_add_14 add_347_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N6329, N6328, N6327, N6326, N6325, N6324}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, N6339, N6338, N6337, N6336, N6335, N6334}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, N6480, N6479, N6478, N6477, N6476, N6475, 
        N6474}) );
  hamming_N16000_CC16_DW01_add_15 add_348_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N6309, N6308, N6307, N6306, N6305, N6304}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, N6319, N6318, N6317, N6316, N6315, N6314}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, N6470, N6469, N6468, N6467, N6466, N6465, 
        N6464}) );
  hamming_N16000_CC16_DW01_add_16 add_349_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N6289, N6288, N6287, N6286, N6285, N6284}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, N6299, N6298, N6297, N6296, N6295, N6294}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, N6460, N6459, N6458, N6457, N6456, N6455, 
        N6454}) );
  hamming_N16000_CC16_DW01_add_17 add_350_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N6269, N6268, N6267, N6266, N6265, N6264}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, N6279, N6278, N6277, N6276, N6275, N6274}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, N6450, N6449, N6448, N6447, N6446, N6445, 
        N6444}) );
  hamming_N16000_CC16_DW01_add_18 add_351_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N6249, N6248, N6247, N6246, N6245, N6244}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, N6259, N6258, N6257, N6256, N6255, N6254}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, N6440, N6439, N6438, N6437, N6436, N6435, 
        N6434}) );
  hamming_N16000_CC16_DW01_add_19 add_352_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N6229, N6228, N6227, N6226, N6225, N6224}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, N6239, N6238, N6237, N6236, N6235, N6234}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, N6430, N6429, N6428, N6427, N6426, N6425, 
        N6424}) );
  hamming_N16000_CC16_DW01_add_20 add_353_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N6209, N6208, N6207, N6206, N6205, N6204}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, N6219, N6218, N6217, N6216, N6215, N6214}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, N6420, N6419, N6418, N6417, N6416, N6415, 
        N6414}) );
  hamming_N16000_CC16_DW01_add_21 add_354_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6188, N6187, N6186, N6185, N6184}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6198, N6197, N6196, N6195, N6194}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, N6409, N6408, 
        N6407, N6406, N6405, N6404}) );
  hamming_N16000_CC16_DW01_add_22 add_355_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6168, N6167, N6166, N6165, N6164}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6178, N6177, N6176, N6175, N6174}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, N6399, N6398, 
        N6397, N6396, N6395, N6394}) );
  hamming_N16000_CC16_DW01_add_23 add_356_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6148, N6147, N6146, N6145, N6144}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6158, N6157, N6156, N6155, N6154}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, N6389, N6388, 
        N6387, N6386, N6385, N6384}) );
  hamming_N16000_CC16_DW01_add_24 add_357_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6128, N6127, N6126, N6125, N6124}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6138, N6137, N6136, N6135, N6134}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, N6379, N6378, 
        N6377, N6376, N6375, N6374}) );
  hamming_N16000_CC16_DW01_add_25 add_358_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6108, N6107, N6106, N6105, N6104}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6118, N6117, N6116, N6115, N6114}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, N6369, N6368, 
        N6367, N6366, N6365, N6364}) );
  hamming_N16000_CC16_DW01_add_26 add_359_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6088, N6087, N6086, N6085, N6084}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6098, N6097, N6096, N6095, N6094}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, N6359, N6358, 
        N6357, N6356, N6355, N6354}) );
  hamming_N16000_CC16_DW01_add_27 add_360_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6068, N6067, N6066, N6065, N6064}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6078, N6077, N6076, N6075, N6074}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, N6349, N6348, 
        N6347, N6346, N6345, N6344}) );
  hamming_N16000_CC16_DW01_add_28 add_361_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6048, N6047, N6046, N6045, N6044}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6058, N6057, N6056, N6055, N6054}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        SYNOPSYS_UNCONNECTED__73, SYNOPSYS_UNCONNECTED__74, N6339, N6338, 
        N6337, N6336, N6335, N6334}) );
  hamming_N16000_CC16_DW01_add_29 add_362_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6028, N6027, N6026, N6025, N6024}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6038, N6037, N6036, N6035, N6034}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__75, SYNOPSYS_UNCONNECTED__76, 
        SYNOPSYS_UNCONNECTED__77, SYNOPSYS_UNCONNECTED__78, N6329, N6328, 
        N6327, N6326, N6325, N6324}) );
  hamming_N16000_CC16_DW01_add_30 add_363_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6008, N6007, N6006, N6005, N6004}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N6018, N6017, N6016, N6015, N6014}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__79, SYNOPSYS_UNCONNECTED__80, 
        SYNOPSYS_UNCONNECTED__81, SYNOPSYS_UNCONNECTED__82, N6319, N6318, 
        N6317, N6316, N6315, N6314}) );
  hamming_N16000_CC16_DW01_add_31 add_364_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5988, N5987, N5986, N5985, N5984}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5998, N5997, N5996, N5995, N5994}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__83, SYNOPSYS_UNCONNECTED__84, 
        SYNOPSYS_UNCONNECTED__85, SYNOPSYS_UNCONNECTED__86, N6309, N6308, 
        N6307, N6306, N6305, N6304}) );
  hamming_N16000_CC16_DW01_add_32 add_365_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5968, N5967, N5966, N5965, N5964}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5978, N5977, N5976, N5975, N5974}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__87, SYNOPSYS_UNCONNECTED__88, 
        SYNOPSYS_UNCONNECTED__89, SYNOPSYS_UNCONNECTED__90, N6299, N6298, 
        N6297, N6296, N6295, N6294}) );
  hamming_N16000_CC16_DW01_add_33 add_366_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5948, N5947, N5946, N5945, N5944}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5958, N5957, N5956, N5955, N5954}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__91, SYNOPSYS_UNCONNECTED__92, 
        SYNOPSYS_UNCONNECTED__93, SYNOPSYS_UNCONNECTED__94, N6289, N6288, 
        N6287, N6286, N6285, N6284}) );
  hamming_N16000_CC16_DW01_add_34 add_367_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5928, N5927, N5926, N5925, N5924}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5938, N5937, N5936, N5935, N5934}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__95, SYNOPSYS_UNCONNECTED__96, 
        SYNOPSYS_UNCONNECTED__97, SYNOPSYS_UNCONNECTED__98, N6279, N6278, 
        N6277, N6276, N6275, N6274}) );
  hamming_N16000_CC16_DW01_add_35 add_368_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5908, N5907, N5906, N5905, N5904}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5918, N5917, N5916, N5915, N5914}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__99, SYNOPSYS_UNCONNECTED__100, 
        SYNOPSYS_UNCONNECTED__101, SYNOPSYS_UNCONNECTED__102, N6269, N6268, 
        N6267, N6266, N6265, N6264}) );
  hamming_N16000_CC16_DW01_add_36 add_369_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5888, N5887, N5886, N5885, N5884}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5898, N5897, N5896, N5895, N5894}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__103, SYNOPSYS_UNCONNECTED__104, 
        SYNOPSYS_UNCONNECTED__105, SYNOPSYS_UNCONNECTED__106, N6259, N6258, 
        N6257, N6256, N6255, N6254}) );
  hamming_N16000_CC16_DW01_add_37 add_370_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5868, N5867, N5866, N5865, N5864}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5878, N5877, N5876, N5875, N5874}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__107, SYNOPSYS_UNCONNECTED__108, 
        SYNOPSYS_UNCONNECTED__109, SYNOPSYS_UNCONNECTED__110, N6249, N6248, 
        N6247, N6246, N6245, N6244}) );
  hamming_N16000_CC16_DW01_add_38 add_371_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5848, N5847, N5846, N5845, N5844}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5858, N5857, N5856, N5855, N5854}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__111, SYNOPSYS_UNCONNECTED__112, 
        SYNOPSYS_UNCONNECTED__113, SYNOPSYS_UNCONNECTED__114, N6239, N6238, 
        N6237, N6236, N6235, N6234}) );
  hamming_N16000_CC16_DW01_add_39 add_372_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5828, N5827, N5826, N5825, N5824}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5838, N5837, N5836, N5835, N5834}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__115, SYNOPSYS_UNCONNECTED__116, 
        SYNOPSYS_UNCONNECTED__117, SYNOPSYS_UNCONNECTED__118, N6229, N6228, 
        N6227, N6226, N6225, N6224}) );
  hamming_N16000_CC16_DW01_add_40 add_373_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5808, N5807, N5806, N5805, N5804}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5818, N5817, N5816, N5815, N5814}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__119, SYNOPSYS_UNCONNECTED__120, 
        SYNOPSYS_UNCONNECTED__121, SYNOPSYS_UNCONNECTED__122, N6219, N6218, 
        N6217, N6216, N6215, N6214}) );
  hamming_N16000_CC16_DW01_add_41 add_374_root_add_47_I1000 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5788, N5787, N5786, N5785, N5784}), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, N5798, N5797, N5796, N5795, N5794}), .CI(1'b0), 
        .SUM({SYNOPSYS_UNCONNECTED__123, SYNOPSYS_UNCONNECTED__124, 
        SYNOPSYS_UNCONNECTED__125, SYNOPSYS_UNCONNECTED__126, N6209, N6208, 
        N6207, N6206, N6205, N6204}) );
  NAND U1686 ( .A(n687), .B(n688), .Z(N6198) );
  NANDN U1687 ( .A(n689), .B(n690), .Z(n688) );
  OR U1688 ( .A(n691), .B(n692), .Z(n690) );
  NAND U1689 ( .A(n691), .B(n692), .Z(n687) );
  XOR U1690 ( .A(n691), .B(n693), .Z(N6197) );
  XNOR U1691 ( .A(n689), .B(n692), .Z(n693) );
  AND U1692 ( .A(n694), .B(n695), .Z(n692) );
  NANDN U1693 ( .A(n696), .B(n697), .Z(n695) );
  NANDN U1694 ( .A(n698), .B(n699), .Z(n697) );
  NANDN U1695 ( .A(n699), .B(n698), .Z(n694) );
  NAND U1696 ( .A(n700), .B(n701), .Z(n689) );
  NANDN U1697 ( .A(n702), .B(n703), .Z(n701) );
  OR U1698 ( .A(n704), .B(n705), .Z(n703) );
  NAND U1699 ( .A(n705), .B(n704), .Z(n700) );
  AND U1700 ( .A(n706), .B(n707), .Z(n691) );
  NANDN U1701 ( .A(n708), .B(n709), .Z(n707) );
  NANDN U1702 ( .A(n710), .B(n711), .Z(n709) );
  NANDN U1703 ( .A(n711), .B(n710), .Z(n706) );
  XOR U1704 ( .A(n705), .B(n712), .Z(N6196) );
  XOR U1705 ( .A(n702), .B(n704), .Z(n712) );
  XNOR U1706 ( .A(n698), .B(n713), .Z(n704) );
  XNOR U1707 ( .A(n696), .B(n699), .Z(n713) );
  NAND U1708 ( .A(n714), .B(n715), .Z(n699) );
  NAND U1709 ( .A(n716), .B(n717), .Z(n715) );
  OR U1710 ( .A(n718), .B(n719), .Z(n716) );
  NANDN U1711 ( .A(n720), .B(n718), .Z(n714) );
  IV U1712 ( .A(n719), .Z(n720) );
  NAND U1713 ( .A(n721), .B(n722), .Z(n696) );
  NAND U1714 ( .A(n723), .B(n724), .Z(n722) );
  NANDN U1715 ( .A(n725), .B(n726), .Z(n723) );
  NANDN U1716 ( .A(n726), .B(n725), .Z(n721) );
  AND U1717 ( .A(n727), .B(n728), .Z(n698) );
  NAND U1718 ( .A(n729), .B(n730), .Z(n728) );
  OR U1719 ( .A(n731), .B(n732), .Z(n729) );
  NANDN U1720 ( .A(n733), .B(n731), .Z(n727) );
  NAND U1721 ( .A(n734), .B(n735), .Z(n702) );
  NANDN U1722 ( .A(n736), .B(n737), .Z(n735) );
  OR U1723 ( .A(n738), .B(n739), .Z(n737) );
  NANDN U1724 ( .A(n740), .B(n738), .Z(n734) );
  IV U1725 ( .A(n739), .Z(n740) );
  XNOR U1726 ( .A(n710), .B(n741), .Z(n705) );
  XNOR U1727 ( .A(n708), .B(n711), .Z(n741) );
  NAND U1728 ( .A(n742), .B(n743), .Z(n711) );
  NAND U1729 ( .A(n744), .B(n745), .Z(n743) );
  OR U1730 ( .A(n746), .B(n747), .Z(n744) );
  NANDN U1731 ( .A(n748), .B(n746), .Z(n742) );
  IV U1732 ( .A(n747), .Z(n748) );
  NAND U1733 ( .A(n749), .B(n750), .Z(n708) );
  NAND U1734 ( .A(n751), .B(n752), .Z(n750) );
  NANDN U1735 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U1736 ( .A(n754), .B(n753), .Z(n749) );
  AND U1737 ( .A(n755), .B(n756), .Z(n710) );
  NAND U1738 ( .A(n757), .B(n758), .Z(n756) );
  OR U1739 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U1740 ( .A(n761), .B(n759), .Z(n755) );
  XNOR U1741 ( .A(n736), .B(n762), .Z(N6195) );
  XOR U1742 ( .A(n738), .B(n739), .Z(n762) );
  XNOR U1743 ( .A(n752), .B(n763), .Z(n739) );
  XOR U1744 ( .A(n753), .B(n754), .Z(n763) );
  XOR U1745 ( .A(n759), .B(n764), .Z(n754) );
  XOR U1746 ( .A(n758), .B(n761), .Z(n764) );
  IV U1747 ( .A(n760), .Z(n761) );
  NAND U1748 ( .A(n765), .B(n766), .Z(n760) );
  OR U1749 ( .A(n767), .B(n768), .Z(n766) );
  OR U1750 ( .A(n769), .B(n770), .Z(n765) );
  NAND U1751 ( .A(n771), .B(n772), .Z(n758) );
  OR U1752 ( .A(n773), .B(n774), .Z(n772) );
  OR U1753 ( .A(n775), .B(n776), .Z(n771) );
  NOR U1754 ( .A(n777), .B(n778), .Z(n759) );
  ANDN U1755 ( .B(n779), .A(n780), .Z(n753) );
  XNOR U1756 ( .A(n746), .B(n781), .Z(n752) );
  XNOR U1757 ( .A(n745), .B(n747), .Z(n781) );
  NAND U1758 ( .A(n782), .B(n783), .Z(n747) );
  OR U1759 ( .A(n784), .B(n785), .Z(n783) );
  OR U1760 ( .A(n786), .B(n787), .Z(n782) );
  NAND U1761 ( .A(n788), .B(n789), .Z(n745) );
  OR U1762 ( .A(n790), .B(n791), .Z(n789) );
  OR U1763 ( .A(n792), .B(n793), .Z(n788) );
  ANDN U1764 ( .B(n794), .A(n795), .Z(n746) );
  IV U1765 ( .A(n796), .Z(n794) );
  ANDN U1766 ( .B(n797), .A(n798), .Z(n738) );
  XOR U1767 ( .A(n724), .B(n799), .Z(n736) );
  XOR U1768 ( .A(n725), .B(n726), .Z(n799) );
  XOR U1769 ( .A(n731), .B(n800), .Z(n726) );
  XOR U1770 ( .A(n730), .B(n733), .Z(n800) );
  IV U1771 ( .A(n732), .Z(n733) );
  NAND U1772 ( .A(n801), .B(n802), .Z(n732) );
  OR U1773 ( .A(n803), .B(n804), .Z(n802) );
  OR U1774 ( .A(n805), .B(n806), .Z(n801) );
  NAND U1775 ( .A(n807), .B(n808), .Z(n730) );
  OR U1776 ( .A(n809), .B(n810), .Z(n808) );
  OR U1777 ( .A(n811), .B(n812), .Z(n807) );
  NOR U1778 ( .A(n813), .B(n814), .Z(n731) );
  ANDN U1779 ( .B(n815), .A(n816), .Z(n725) );
  IV U1780 ( .A(n817), .Z(n815) );
  XNOR U1781 ( .A(n718), .B(n818), .Z(n724) );
  XNOR U1782 ( .A(n717), .B(n719), .Z(n818) );
  NAND U1783 ( .A(n819), .B(n820), .Z(n719) );
  OR U1784 ( .A(n821), .B(n822), .Z(n820) );
  OR U1785 ( .A(n823), .B(n824), .Z(n819) );
  NAND U1786 ( .A(n825), .B(n826), .Z(n717) );
  OR U1787 ( .A(n827), .B(n828), .Z(n826) );
  OR U1788 ( .A(n829), .B(n830), .Z(n825) );
  ANDN U1789 ( .B(n831), .A(n832), .Z(n718) );
  IV U1790 ( .A(n833), .Z(n831) );
  XNOR U1791 ( .A(n798), .B(n797), .Z(N6194) );
  XOR U1792 ( .A(n817), .B(n816), .Z(n797) );
  XNOR U1793 ( .A(n832), .B(n833), .Z(n816) );
  XNOR U1794 ( .A(n827), .B(n828), .Z(n833) );
  XNOR U1795 ( .A(n829), .B(n830), .Z(n828) );
  XNOR U1796 ( .A(y[988]), .B(x[988]), .Z(n830) );
  XNOR U1797 ( .A(y[989]), .B(x[989]), .Z(n829) );
  XNOR U1798 ( .A(y[987]), .B(x[987]), .Z(n827) );
  XNOR U1799 ( .A(n821), .B(n822), .Z(n832) );
  XNOR U1800 ( .A(y[984]), .B(x[984]), .Z(n822) );
  XNOR U1801 ( .A(n823), .B(n824), .Z(n821) );
  XNOR U1802 ( .A(y[985]), .B(x[985]), .Z(n824) );
  XNOR U1803 ( .A(y[986]), .B(x[986]), .Z(n823) );
  XNOR U1804 ( .A(n814), .B(n813), .Z(n817) );
  XNOR U1805 ( .A(n809), .B(n810), .Z(n813) );
  XNOR U1806 ( .A(y[981]), .B(x[981]), .Z(n810) );
  XNOR U1807 ( .A(n811), .B(n812), .Z(n809) );
  XNOR U1808 ( .A(y[982]), .B(x[982]), .Z(n812) );
  XNOR U1809 ( .A(y[983]), .B(x[983]), .Z(n811) );
  XNOR U1810 ( .A(n803), .B(n804), .Z(n814) );
  XNOR U1811 ( .A(y[978]), .B(x[978]), .Z(n804) );
  XNOR U1812 ( .A(n805), .B(n806), .Z(n803) );
  XNOR U1813 ( .A(y[979]), .B(x[979]), .Z(n806) );
  XNOR U1814 ( .A(y[980]), .B(x[980]), .Z(n805) );
  XOR U1815 ( .A(n779), .B(n780), .Z(n798) );
  XNOR U1816 ( .A(n795), .B(n796), .Z(n780) );
  XNOR U1817 ( .A(n790), .B(n791), .Z(n796) );
  XNOR U1818 ( .A(n792), .B(n793), .Z(n791) );
  XNOR U1819 ( .A(y[976]), .B(x[976]), .Z(n793) );
  XNOR U1820 ( .A(y[977]), .B(x[977]), .Z(n792) );
  XNOR U1821 ( .A(y[975]), .B(x[975]), .Z(n790) );
  XNOR U1822 ( .A(n784), .B(n785), .Z(n795) );
  XNOR U1823 ( .A(y[972]), .B(x[972]), .Z(n785) );
  XNOR U1824 ( .A(n786), .B(n787), .Z(n784) );
  XNOR U1825 ( .A(y[973]), .B(x[973]), .Z(n787) );
  XNOR U1826 ( .A(y[974]), .B(x[974]), .Z(n786) );
  XOR U1827 ( .A(n778), .B(n777), .Z(n779) );
  XNOR U1828 ( .A(n773), .B(n774), .Z(n777) );
  XNOR U1829 ( .A(y[969]), .B(x[969]), .Z(n774) );
  XNOR U1830 ( .A(n775), .B(n776), .Z(n773) );
  XNOR U1831 ( .A(y[970]), .B(x[970]), .Z(n776) );
  XNOR U1832 ( .A(y[971]), .B(x[971]), .Z(n775) );
  XNOR U1833 ( .A(n767), .B(n768), .Z(n778) );
  XNOR U1834 ( .A(y[966]), .B(x[966]), .Z(n768) );
  XNOR U1835 ( .A(n769), .B(n770), .Z(n767) );
  XNOR U1836 ( .A(y[967]), .B(x[967]), .Z(n770) );
  XNOR U1837 ( .A(y[968]), .B(x[968]), .Z(n769) );
  NAND U1838 ( .A(n834), .B(n835), .Z(N6188) );
  NANDN U1839 ( .A(n836), .B(n837), .Z(n835) );
  OR U1840 ( .A(n838), .B(n839), .Z(n837) );
  NAND U1841 ( .A(n838), .B(n839), .Z(n834) );
  XOR U1842 ( .A(n838), .B(n840), .Z(N6187) );
  XNOR U1843 ( .A(n836), .B(n839), .Z(n840) );
  AND U1844 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U1845 ( .A(n843), .B(n844), .Z(n842) );
  NANDN U1846 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U1847 ( .A(n846), .B(n845), .Z(n841) );
  NAND U1848 ( .A(n847), .B(n848), .Z(n836) );
  NANDN U1849 ( .A(n849), .B(n850), .Z(n848) );
  OR U1850 ( .A(n851), .B(n852), .Z(n850) );
  NAND U1851 ( .A(n852), .B(n851), .Z(n847) );
  AND U1852 ( .A(n853), .B(n854), .Z(n838) );
  NANDN U1853 ( .A(n855), .B(n856), .Z(n854) );
  NANDN U1854 ( .A(n857), .B(n858), .Z(n856) );
  NANDN U1855 ( .A(n858), .B(n857), .Z(n853) );
  XOR U1856 ( .A(n852), .B(n859), .Z(N6186) );
  XOR U1857 ( .A(n849), .B(n851), .Z(n859) );
  XNOR U1858 ( .A(n845), .B(n860), .Z(n851) );
  XNOR U1859 ( .A(n843), .B(n846), .Z(n860) );
  NAND U1860 ( .A(n861), .B(n862), .Z(n846) );
  NAND U1861 ( .A(n863), .B(n864), .Z(n862) );
  OR U1862 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U1863 ( .A(n867), .B(n865), .Z(n861) );
  IV U1864 ( .A(n866), .Z(n867) );
  NAND U1865 ( .A(n868), .B(n869), .Z(n843) );
  NAND U1866 ( .A(n870), .B(n871), .Z(n869) );
  NANDN U1867 ( .A(n872), .B(n873), .Z(n870) );
  NANDN U1868 ( .A(n873), .B(n872), .Z(n868) );
  AND U1869 ( .A(n874), .B(n875), .Z(n845) );
  NAND U1870 ( .A(n876), .B(n877), .Z(n875) );
  OR U1871 ( .A(n878), .B(n879), .Z(n876) );
  NANDN U1872 ( .A(n880), .B(n878), .Z(n874) );
  NAND U1873 ( .A(n881), .B(n882), .Z(n849) );
  NANDN U1874 ( .A(n883), .B(n884), .Z(n882) );
  OR U1875 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U1876 ( .A(n887), .B(n885), .Z(n881) );
  IV U1877 ( .A(n886), .Z(n887) );
  XNOR U1878 ( .A(n857), .B(n888), .Z(n852) );
  XNOR U1879 ( .A(n855), .B(n858), .Z(n888) );
  NAND U1880 ( .A(n889), .B(n890), .Z(n858) );
  NAND U1881 ( .A(n891), .B(n892), .Z(n890) );
  OR U1882 ( .A(n893), .B(n894), .Z(n891) );
  NANDN U1883 ( .A(n895), .B(n893), .Z(n889) );
  IV U1884 ( .A(n894), .Z(n895) );
  NAND U1885 ( .A(n896), .B(n897), .Z(n855) );
  NAND U1886 ( .A(n898), .B(n899), .Z(n897) );
  NANDN U1887 ( .A(n900), .B(n901), .Z(n898) );
  NANDN U1888 ( .A(n901), .B(n900), .Z(n896) );
  AND U1889 ( .A(n902), .B(n903), .Z(n857) );
  NAND U1890 ( .A(n904), .B(n905), .Z(n903) );
  OR U1891 ( .A(n906), .B(n907), .Z(n904) );
  NANDN U1892 ( .A(n908), .B(n906), .Z(n902) );
  XNOR U1893 ( .A(n883), .B(n909), .Z(N6185) );
  XOR U1894 ( .A(n885), .B(n886), .Z(n909) );
  XNOR U1895 ( .A(n899), .B(n910), .Z(n886) );
  XOR U1896 ( .A(n900), .B(n901), .Z(n910) );
  XOR U1897 ( .A(n906), .B(n911), .Z(n901) );
  XOR U1898 ( .A(n905), .B(n908), .Z(n911) );
  IV U1899 ( .A(n907), .Z(n908) );
  NAND U1900 ( .A(n912), .B(n913), .Z(n907) );
  OR U1901 ( .A(n914), .B(n915), .Z(n913) );
  OR U1902 ( .A(n916), .B(n917), .Z(n912) );
  NAND U1903 ( .A(n918), .B(n919), .Z(n905) );
  OR U1904 ( .A(n920), .B(n921), .Z(n919) );
  OR U1905 ( .A(n922), .B(n923), .Z(n918) );
  NOR U1906 ( .A(n924), .B(n925), .Z(n906) );
  ANDN U1907 ( .B(n926), .A(n927), .Z(n900) );
  XNOR U1908 ( .A(n893), .B(n928), .Z(n899) );
  XNOR U1909 ( .A(n892), .B(n894), .Z(n928) );
  NAND U1910 ( .A(n929), .B(n930), .Z(n894) );
  OR U1911 ( .A(n931), .B(n932), .Z(n930) );
  OR U1912 ( .A(n933), .B(n934), .Z(n929) );
  NAND U1913 ( .A(n935), .B(n936), .Z(n892) );
  OR U1914 ( .A(n937), .B(n938), .Z(n936) );
  OR U1915 ( .A(n939), .B(n940), .Z(n935) );
  ANDN U1916 ( .B(n941), .A(n942), .Z(n893) );
  IV U1917 ( .A(n943), .Z(n941) );
  ANDN U1918 ( .B(n944), .A(n945), .Z(n885) );
  XOR U1919 ( .A(n871), .B(n946), .Z(n883) );
  XOR U1920 ( .A(n872), .B(n873), .Z(n946) );
  XOR U1921 ( .A(n878), .B(n947), .Z(n873) );
  XOR U1922 ( .A(n877), .B(n880), .Z(n947) );
  IV U1923 ( .A(n879), .Z(n880) );
  NAND U1924 ( .A(n948), .B(n949), .Z(n879) );
  OR U1925 ( .A(n950), .B(n951), .Z(n949) );
  OR U1926 ( .A(n952), .B(n953), .Z(n948) );
  NAND U1927 ( .A(n954), .B(n955), .Z(n877) );
  OR U1928 ( .A(n956), .B(n957), .Z(n955) );
  OR U1929 ( .A(n958), .B(n959), .Z(n954) );
  NOR U1930 ( .A(n960), .B(n961), .Z(n878) );
  ANDN U1931 ( .B(n962), .A(n963), .Z(n872) );
  IV U1932 ( .A(n964), .Z(n962) );
  XNOR U1933 ( .A(n865), .B(n965), .Z(n871) );
  XNOR U1934 ( .A(n864), .B(n866), .Z(n965) );
  NAND U1935 ( .A(n966), .B(n967), .Z(n866) );
  OR U1936 ( .A(n968), .B(n969), .Z(n967) );
  OR U1937 ( .A(n970), .B(n971), .Z(n966) );
  NAND U1938 ( .A(n972), .B(n973), .Z(n864) );
  OR U1939 ( .A(n974), .B(n975), .Z(n973) );
  OR U1940 ( .A(n976), .B(n977), .Z(n972) );
  ANDN U1941 ( .B(n978), .A(n979), .Z(n865) );
  IV U1942 ( .A(n980), .Z(n978) );
  XNOR U1943 ( .A(n945), .B(n944), .Z(N6184) );
  XOR U1944 ( .A(n964), .B(n963), .Z(n944) );
  XNOR U1945 ( .A(n979), .B(n980), .Z(n963) );
  XNOR U1946 ( .A(n974), .B(n975), .Z(n980) );
  XNOR U1947 ( .A(n976), .B(n977), .Z(n975) );
  XNOR U1948 ( .A(y[964]), .B(x[964]), .Z(n977) );
  XNOR U1949 ( .A(y[965]), .B(x[965]), .Z(n976) );
  XNOR U1950 ( .A(y[963]), .B(x[963]), .Z(n974) );
  XNOR U1951 ( .A(n968), .B(n969), .Z(n979) );
  XNOR U1952 ( .A(y[960]), .B(x[960]), .Z(n969) );
  XNOR U1953 ( .A(n970), .B(n971), .Z(n968) );
  XNOR U1954 ( .A(y[961]), .B(x[961]), .Z(n971) );
  XNOR U1955 ( .A(y[962]), .B(x[962]), .Z(n970) );
  XNOR U1956 ( .A(n961), .B(n960), .Z(n964) );
  XNOR U1957 ( .A(n956), .B(n957), .Z(n960) );
  XNOR U1958 ( .A(y[957]), .B(x[957]), .Z(n957) );
  XNOR U1959 ( .A(n958), .B(n959), .Z(n956) );
  XNOR U1960 ( .A(y[958]), .B(x[958]), .Z(n959) );
  XNOR U1961 ( .A(y[959]), .B(x[959]), .Z(n958) );
  XNOR U1962 ( .A(n950), .B(n951), .Z(n961) );
  XNOR U1963 ( .A(y[954]), .B(x[954]), .Z(n951) );
  XNOR U1964 ( .A(n952), .B(n953), .Z(n950) );
  XNOR U1965 ( .A(y[955]), .B(x[955]), .Z(n953) );
  XNOR U1966 ( .A(y[956]), .B(x[956]), .Z(n952) );
  XOR U1967 ( .A(n926), .B(n927), .Z(n945) );
  XNOR U1968 ( .A(n942), .B(n943), .Z(n927) );
  XNOR U1969 ( .A(n937), .B(n938), .Z(n943) );
  XNOR U1970 ( .A(n939), .B(n940), .Z(n938) );
  XNOR U1971 ( .A(y[952]), .B(x[952]), .Z(n940) );
  XNOR U1972 ( .A(y[953]), .B(x[953]), .Z(n939) );
  XNOR U1973 ( .A(y[951]), .B(x[951]), .Z(n937) );
  XNOR U1974 ( .A(n931), .B(n932), .Z(n942) );
  XNOR U1975 ( .A(y[948]), .B(x[948]), .Z(n932) );
  XNOR U1976 ( .A(n933), .B(n934), .Z(n931) );
  XNOR U1977 ( .A(y[949]), .B(x[949]), .Z(n934) );
  XNOR U1978 ( .A(y[950]), .B(x[950]), .Z(n933) );
  XOR U1979 ( .A(n925), .B(n924), .Z(n926) );
  XNOR U1980 ( .A(n920), .B(n921), .Z(n924) );
  XNOR U1981 ( .A(y[945]), .B(x[945]), .Z(n921) );
  XNOR U1982 ( .A(n922), .B(n923), .Z(n920) );
  XNOR U1983 ( .A(y[946]), .B(x[946]), .Z(n923) );
  XNOR U1984 ( .A(y[947]), .B(x[947]), .Z(n922) );
  XNOR U1985 ( .A(n914), .B(n915), .Z(n925) );
  XNOR U1986 ( .A(y[942]), .B(x[942]), .Z(n915) );
  XNOR U1987 ( .A(n916), .B(n917), .Z(n914) );
  XNOR U1988 ( .A(y[943]), .B(x[943]), .Z(n917) );
  XNOR U1989 ( .A(y[944]), .B(x[944]), .Z(n916) );
  NAND U1990 ( .A(n981), .B(n982), .Z(N6178) );
  NANDN U1991 ( .A(n983), .B(n984), .Z(n982) );
  OR U1992 ( .A(n985), .B(n986), .Z(n984) );
  NAND U1993 ( .A(n985), .B(n986), .Z(n981) );
  XOR U1994 ( .A(n985), .B(n987), .Z(N6177) );
  XNOR U1995 ( .A(n983), .B(n986), .Z(n987) );
  AND U1996 ( .A(n988), .B(n989), .Z(n986) );
  NANDN U1997 ( .A(n990), .B(n991), .Z(n989) );
  NANDN U1998 ( .A(n992), .B(n993), .Z(n991) );
  NANDN U1999 ( .A(n993), .B(n992), .Z(n988) );
  NAND U2000 ( .A(n994), .B(n995), .Z(n983) );
  NANDN U2001 ( .A(n996), .B(n997), .Z(n995) );
  OR U2002 ( .A(n998), .B(n999), .Z(n997) );
  NAND U2003 ( .A(n999), .B(n998), .Z(n994) );
  AND U2004 ( .A(n1000), .B(n1001), .Z(n985) );
  NANDN U2005 ( .A(n1002), .B(n1003), .Z(n1001) );
  NANDN U2006 ( .A(n1004), .B(n1005), .Z(n1003) );
  NANDN U2007 ( .A(n1005), .B(n1004), .Z(n1000) );
  XOR U2008 ( .A(n999), .B(n1006), .Z(N6176) );
  XOR U2009 ( .A(n996), .B(n998), .Z(n1006) );
  XNOR U2010 ( .A(n992), .B(n1007), .Z(n998) );
  XNOR U2011 ( .A(n990), .B(n993), .Z(n1007) );
  NAND U2012 ( .A(n1008), .B(n1009), .Z(n993) );
  NAND U2013 ( .A(n1010), .B(n1011), .Z(n1009) );
  OR U2014 ( .A(n1012), .B(n1013), .Z(n1010) );
  NANDN U2015 ( .A(n1014), .B(n1012), .Z(n1008) );
  IV U2016 ( .A(n1013), .Z(n1014) );
  NAND U2017 ( .A(n1015), .B(n1016), .Z(n990) );
  NAND U2018 ( .A(n1017), .B(n1018), .Z(n1016) );
  NANDN U2019 ( .A(n1019), .B(n1020), .Z(n1017) );
  NANDN U2020 ( .A(n1020), .B(n1019), .Z(n1015) );
  AND U2021 ( .A(n1021), .B(n1022), .Z(n992) );
  NAND U2022 ( .A(n1023), .B(n1024), .Z(n1022) );
  OR U2023 ( .A(n1025), .B(n1026), .Z(n1023) );
  NANDN U2024 ( .A(n1027), .B(n1025), .Z(n1021) );
  NAND U2025 ( .A(n1028), .B(n1029), .Z(n996) );
  NANDN U2026 ( .A(n1030), .B(n1031), .Z(n1029) );
  OR U2027 ( .A(n1032), .B(n1033), .Z(n1031) );
  NANDN U2028 ( .A(n1034), .B(n1032), .Z(n1028) );
  IV U2029 ( .A(n1033), .Z(n1034) );
  XNOR U2030 ( .A(n1004), .B(n1035), .Z(n999) );
  XNOR U2031 ( .A(n1002), .B(n1005), .Z(n1035) );
  NAND U2032 ( .A(n1036), .B(n1037), .Z(n1005) );
  NAND U2033 ( .A(n1038), .B(n1039), .Z(n1037) );
  OR U2034 ( .A(n1040), .B(n1041), .Z(n1038) );
  NANDN U2035 ( .A(n1042), .B(n1040), .Z(n1036) );
  IV U2036 ( .A(n1041), .Z(n1042) );
  NAND U2037 ( .A(n1043), .B(n1044), .Z(n1002) );
  NAND U2038 ( .A(n1045), .B(n1046), .Z(n1044) );
  NANDN U2039 ( .A(n1047), .B(n1048), .Z(n1045) );
  NANDN U2040 ( .A(n1048), .B(n1047), .Z(n1043) );
  AND U2041 ( .A(n1049), .B(n1050), .Z(n1004) );
  NAND U2042 ( .A(n1051), .B(n1052), .Z(n1050) );
  OR U2043 ( .A(n1053), .B(n1054), .Z(n1051) );
  NANDN U2044 ( .A(n1055), .B(n1053), .Z(n1049) );
  XNOR U2045 ( .A(n1030), .B(n1056), .Z(N6175) );
  XOR U2046 ( .A(n1032), .B(n1033), .Z(n1056) );
  XNOR U2047 ( .A(n1046), .B(n1057), .Z(n1033) );
  XOR U2048 ( .A(n1047), .B(n1048), .Z(n1057) );
  XOR U2049 ( .A(n1053), .B(n1058), .Z(n1048) );
  XOR U2050 ( .A(n1052), .B(n1055), .Z(n1058) );
  IV U2051 ( .A(n1054), .Z(n1055) );
  NAND U2052 ( .A(n1059), .B(n1060), .Z(n1054) );
  OR U2053 ( .A(n1061), .B(n1062), .Z(n1060) );
  OR U2054 ( .A(n1063), .B(n1064), .Z(n1059) );
  NAND U2055 ( .A(n1065), .B(n1066), .Z(n1052) );
  OR U2056 ( .A(n1067), .B(n1068), .Z(n1066) );
  OR U2057 ( .A(n1069), .B(n1070), .Z(n1065) );
  NOR U2058 ( .A(n1071), .B(n1072), .Z(n1053) );
  ANDN U2059 ( .B(n1073), .A(n1074), .Z(n1047) );
  XNOR U2060 ( .A(n1040), .B(n1075), .Z(n1046) );
  XNOR U2061 ( .A(n1039), .B(n1041), .Z(n1075) );
  NAND U2062 ( .A(n1076), .B(n1077), .Z(n1041) );
  OR U2063 ( .A(n1078), .B(n1079), .Z(n1077) );
  OR U2064 ( .A(n1080), .B(n1081), .Z(n1076) );
  NAND U2065 ( .A(n1082), .B(n1083), .Z(n1039) );
  OR U2066 ( .A(n1084), .B(n1085), .Z(n1083) );
  OR U2067 ( .A(n1086), .B(n1087), .Z(n1082) );
  ANDN U2068 ( .B(n1088), .A(n1089), .Z(n1040) );
  IV U2069 ( .A(n1090), .Z(n1088) );
  ANDN U2070 ( .B(n1091), .A(n1092), .Z(n1032) );
  XOR U2071 ( .A(n1018), .B(n1093), .Z(n1030) );
  XOR U2072 ( .A(n1019), .B(n1020), .Z(n1093) );
  XOR U2073 ( .A(n1025), .B(n1094), .Z(n1020) );
  XOR U2074 ( .A(n1024), .B(n1027), .Z(n1094) );
  IV U2075 ( .A(n1026), .Z(n1027) );
  NAND U2076 ( .A(n1095), .B(n1096), .Z(n1026) );
  OR U2077 ( .A(n1097), .B(n1098), .Z(n1096) );
  OR U2078 ( .A(n1099), .B(n1100), .Z(n1095) );
  NAND U2079 ( .A(n1101), .B(n1102), .Z(n1024) );
  OR U2080 ( .A(n1103), .B(n1104), .Z(n1102) );
  OR U2081 ( .A(n1105), .B(n1106), .Z(n1101) );
  NOR U2082 ( .A(n1107), .B(n1108), .Z(n1025) );
  ANDN U2083 ( .B(n1109), .A(n1110), .Z(n1019) );
  IV U2084 ( .A(n1111), .Z(n1109) );
  XNOR U2085 ( .A(n1012), .B(n1112), .Z(n1018) );
  XNOR U2086 ( .A(n1011), .B(n1013), .Z(n1112) );
  NAND U2087 ( .A(n1113), .B(n1114), .Z(n1013) );
  OR U2088 ( .A(n1115), .B(n1116), .Z(n1114) );
  OR U2089 ( .A(n1117), .B(n1118), .Z(n1113) );
  NAND U2090 ( .A(n1119), .B(n1120), .Z(n1011) );
  OR U2091 ( .A(n1121), .B(n1122), .Z(n1120) );
  OR U2092 ( .A(n1123), .B(n1124), .Z(n1119) );
  ANDN U2093 ( .B(n1125), .A(n1126), .Z(n1012) );
  IV U2094 ( .A(n1127), .Z(n1125) );
  XNOR U2095 ( .A(n1092), .B(n1091), .Z(N6174) );
  XOR U2096 ( .A(n1111), .B(n1110), .Z(n1091) );
  XNOR U2097 ( .A(n1126), .B(n1127), .Z(n1110) );
  XNOR U2098 ( .A(n1121), .B(n1122), .Z(n1127) );
  XNOR U2099 ( .A(n1123), .B(n1124), .Z(n1122) );
  XNOR U2100 ( .A(y[940]), .B(x[940]), .Z(n1124) );
  XNOR U2101 ( .A(y[941]), .B(x[941]), .Z(n1123) );
  XNOR U2102 ( .A(y[939]), .B(x[939]), .Z(n1121) );
  XNOR U2103 ( .A(n1115), .B(n1116), .Z(n1126) );
  XNOR U2104 ( .A(y[936]), .B(x[936]), .Z(n1116) );
  XNOR U2105 ( .A(n1117), .B(n1118), .Z(n1115) );
  XNOR U2106 ( .A(y[937]), .B(x[937]), .Z(n1118) );
  XNOR U2107 ( .A(y[938]), .B(x[938]), .Z(n1117) );
  XNOR U2108 ( .A(n1108), .B(n1107), .Z(n1111) );
  XNOR U2109 ( .A(n1103), .B(n1104), .Z(n1107) );
  XNOR U2110 ( .A(y[933]), .B(x[933]), .Z(n1104) );
  XNOR U2111 ( .A(n1105), .B(n1106), .Z(n1103) );
  XNOR U2112 ( .A(y[934]), .B(x[934]), .Z(n1106) );
  XNOR U2113 ( .A(y[935]), .B(x[935]), .Z(n1105) );
  XNOR U2114 ( .A(n1097), .B(n1098), .Z(n1108) );
  XNOR U2115 ( .A(y[930]), .B(x[930]), .Z(n1098) );
  XNOR U2116 ( .A(n1099), .B(n1100), .Z(n1097) );
  XNOR U2117 ( .A(y[931]), .B(x[931]), .Z(n1100) );
  XNOR U2118 ( .A(y[932]), .B(x[932]), .Z(n1099) );
  XOR U2119 ( .A(n1073), .B(n1074), .Z(n1092) );
  XNOR U2120 ( .A(n1089), .B(n1090), .Z(n1074) );
  XNOR U2121 ( .A(n1084), .B(n1085), .Z(n1090) );
  XNOR U2122 ( .A(n1086), .B(n1087), .Z(n1085) );
  XNOR U2123 ( .A(y[928]), .B(x[928]), .Z(n1087) );
  XNOR U2124 ( .A(y[929]), .B(x[929]), .Z(n1086) );
  XNOR U2125 ( .A(y[927]), .B(x[927]), .Z(n1084) );
  XNOR U2126 ( .A(n1078), .B(n1079), .Z(n1089) );
  XNOR U2127 ( .A(y[924]), .B(x[924]), .Z(n1079) );
  XNOR U2128 ( .A(n1080), .B(n1081), .Z(n1078) );
  XNOR U2129 ( .A(y[925]), .B(x[925]), .Z(n1081) );
  XNOR U2130 ( .A(y[926]), .B(x[926]), .Z(n1080) );
  XOR U2131 ( .A(n1072), .B(n1071), .Z(n1073) );
  XNOR U2132 ( .A(n1067), .B(n1068), .Z(n1071) );
  XNOR U2133 ( .A(y[921]), .B(x[921]), .Z(n1068) );
  XNOR U2134 ( .A(n1069), .B(n1070), .Z(n1067) );
  XNOR U2135 ( .A(y[922]), .B(x[922]), .Z(n1070) );
  XNOR U2136 ( .A(y[923]), .B(x[923]), .Z(n1069) );
  XNOR U2137 ( .A(n1061), .B(n1062), .Z(n1072) );
  XNOR U2138 ( .A(y[918]), .B(x[918]), .Z(n1062) );
  XNOR U2139 ( .A(n1063), .B(n1064), .Z(n1061) );
  XNOR U2140 ( .A(y[919]), .B(x[919]), .Z(n1064) );
  XNOR U2141 ( .A(y[920]), .B(x[920]), .Z(n1063) );
  NAND U2142 ( .A(n1128), .B(n1129), .Z(N6168) );
  NANDN U2143 ( .A(n1130), .B(n1131), .Z(n1129) );
  OR U2144 ( .A(n1132), .B(n1133), .Z(n1131) );
  NAND U2145 ( .A(n1132), .B(n1133), .Z(n1128) );
  XOR U2146 ( .A(n1132), .B(n1134), .Z(N6167) );
  XNOR U2147 ( .A(n1130), .B(n1133), .Z(n1134) );
  AND U2148 ( .A(n1135), .B(n1136), .Z(n1133) );
  NANDN U2149 ( .A(n1137), .B(n1138), .Z(n1136) );
  NANDN U2150 ( .A(n1139), .B(n1140), .Z(n1138) );
  NANDN U2151 ( .A(n1140), .B(n1139), .Z(n1135) );
  NAND U2152 ( .A(n1141), .B(n1142), .Z(n1130) );
  NANDN U2153 ( .A(n1143), .B(n1144), .Z(n1142) );
  OR U2154 ( .A(n1145), .B(n1146), .Z(n1144) );
  NAND U2155 ( .A(n1146), .B(n1145), .Z(n1141) );
  AND U2156 ( .A(n1147), .B(n1148), .Z(n1132) );
  NANDN U2157 ( .A(n1149), .B(n1150), .Z(n1148) );
  NANDN U2158 ( .A(n1151), .B(n1152), .Z(n1150) );
  NANDN U2159 ( .A(n1152), .B(n1151), .Z(n1147) );
  XOR U2160 ( .A(n1146), .B(n1153), .Z(N6166) );
  XOR U2161 ( .A(n1143), .B(n1145), .Z(n1153) );
  XNOR U2162 ( .A(n1139), .B(n1154), .Z(n1145) );
  XNOR U2163 ( .A(n1137), .B(n1140), .Z(n1154) );
  NAND U2164 ( .A(n1155), .B(n1156), .Z(n1140) );
  NAND U2165 ( .A(n1157), .B(n1158), .Z(n1156) );
  OR U2166 ( .A(n1159), .B(n1160), .Z(n1157) );
  NANDN U2167 ( .A(n1161), .B(n1159), .Z(n1155) );
  IV U2168 ( .A(n1160), .Z(n1161) );
  NAND U2169 ( .A(n1162), .B(n1163), .Z(n1137) );
  NAND U2170 ( .A(n1164), .B(n1165), .Z(n1163) );
  NANDN U2171 ( .A(n1166), .B(n1167), .Z(n1164) );
  NANDN U2172 ( .A(n1167), .B(n1166), .Z(n1162) );
  AND U2173 ( .A(n1168), .B(n1169), .Z(n1139) );
  NAND U2174 ( .A(n1170), .B(n1171), .Z(n1169) );
  OR U2175 ( .A(n1172), .B(n1173), .Z(n1170) );
  NANDN U2176 ( .A(n1174), .B(n1172), .Z(n1168) );
  NAND U2177 ( .A(n1175), .B(n1176), .Z(n1143) );
  NANDN U2178 ( .A(n1177), .B(n1178), .Z(n1176) );
  OR U2179 ( .A(n1179), .B(n1180), .Z(n1178) );
  NANDN U2180 ( .A(n1181), .B(n1179), .Z(n1175) );
  IV U2181 ( .A(n1180), .Z(n1181) );
  XNOR U2182 ( .A(n1151), .B(n1182), .Z(n1146) );
  XNOR U2183 ( .A(n1149), .B(n1152), .Z(n1182) );
  NAND U2184 ( .A(n1183), .B(n1184), .Z(n1152) );
  NAND U2185 ( .A(n1185), .B(n1186), .Z(n1184) );
  OR U2186 ( .A(n1187), .B(n1188), .Z(n1185) );
  NANDN U2187 ( .A(n1189), .B(n1187), .Z(n1183) );
  IV U2188 ( .A(n1188), .Z(n1189) );
  NAND U2189 ( .A(n1190), .B(n1191), .Z(n1149) );
  NAND U2190 ( .A(n1192), .B(n1193), .Z(n1191) );
  NANDN U2191 ( .A(n1194), .B(n1195), .Z(n1192) );
  NANDN U2192 ( .A(n1195), .B(n1194), .Z(n1190) );
  AND U2193 ( .A(n1196), .B(n1197), .Z(n1151) );
  NAND U2194 ( .A(n1198), .B(n1199), .Z(n1197) );
  OR U2195 ( .A(n1200), .B(n1201), .Z(n1198) );
  NANDN U2196 ( .A(n1202), .B(n1200), .Z(n1196) );
  XNOR U2197 ( .A(n1177), .B(n1203), .Z(N6165) );
  XOR U2198 ( .A(n1179), .B(n1180), .Z(n1203) );
  XNOR U2199 ( .A(n1193), .B(n1204), .Z(n1180) );
  XOR U2200 ( .A(n1194), .B(n1195), .Z(n1204) );
  XOR U2201 ( .A(n1200), .B(n1205), .Z(n1195) );
  XOR U2202 ( .A(n1199), .B(n1202), .Z(n1205) );
  IV U2203 ( .A(n1201), .Z(n1202) );
  NAND U2204 ( .A(n1206), .B(n1207), .Z(n1201) );
  OR U2205 ( .A(n1208), .B(n1209), .Z(n1207) );
  OR U2206 ( .A(n1210), .B(n1211), .Z(n1206) );
  NAND U2207 ( .A(n1212), .B(n1213), .Z(n1199) );
  OR U2208 ( .A(n1214), .B(n1215), .Z(n1213) );
  OR U2209 ( .A(n1216), .B(n1217), .Z(n1212) );
  NOR U2210 ( .A(n1218), .B(n1219), .Z(n1200) );
  ANDN U2211 ( .B(n1220), .A(n1221), .Z(n1194) );
  XNOR U2212 ( .A(n1187), .B(n1222), .Z(n1193) );
  XNOR U2213 ( .A(n1186), .B(n1188), .Z(n1222) );
  NAND U2214 ( .A(n1223), .B(n1224), .Z(n1188) );
  OR U2215 ( .A(n1225), .B(n1226), .Z(n1224) );
  OR U2216 ( .A(n1227), .B(n1228), .Z(n1223) );
  NAND U2217 ( .A(n1229), .B(n1230), .Z(n1186) );
  OR U2218 ( .A(n1231), .B(n1232), .Z(n1230) );
  OR U2219 ( .A(n1233), .B(n1234), .Z(n1229) );
  ANDN U2220 ( .B(n1235), .A(n1236), .Z(n1187) );
  IV U2221 ( .A(n1237), .Z(n1235) );
  ANDN U2222 ( .B(n1238), .A(n1239), .Z(n1179) );
  XOR U2223 ( .A(n1165), .B(n1240), .Z(n1177) );
  XOR U2224 ( .A(n1166), .B(n1167), .Z(n1240) );
  XOR U2225 ( .A(n1172), .B(n1241), .Z(n1167) );
  XOR U2226 ( .A(n1171), .B(n1174), .Z(n1241) );
  IV U2227 ( .A(n1173), .Z(n1174) );
  NAND U2228 ( .A(n1242), .B(n1243), .Z(n1173) );
  OR U2229 ( .A(n1244), .B(n1245), .Z(n1243) );
  OR U2230 ( .A(n1246), .B(n1247), .Z(n1242) );
  NAND U2231 ( .A(n1248), .B(n1249), .Z(n1171) );
  OR U2232 ( .A(n1250), .B(n1251), .Z(n1249) );
  OR U2233 ( .A(n1252), .B(n1253), .Z(n1248) );
  NOR U2234 ( .A(n1254), .B(n1255), .Z(n1172) );
  ANDN U2235 ( .B(n1256), .A(n1257), .Z(n1166) );
  IV U2236 ( .A(n1258), .Z(n1256) );
  XNOR U2237 ( .A(n1159), .B(n1259), .Z(n1165) );
  XNOR U2238 ( .A(n1158), .B(n1160), .Z(n1259) );
  NAND U2239 ( .A(n1260), .B(n1261), .Z(n1160) );
  OR U2240 ( .A(n1262), .B(n1263), .Z(n1261) );
  OR U2241 ( .A(n1264), .B(n1265), .Z(n1260) );
  NAND U2242 ( .A(n1266), .B(n1267), .Z(n1158) );
  OR U2243 ( .A(n1268), .B(n1269), .Z(n1267) );
  OR U2244 ( .A(n1270), .B(n1271), .Z(n1266) );
  ANDN U2245 ( .B(n1272), .A(n1273), .Z(n1159) );
  IV U2246 ( .A(n1274), .Z(n1272) );
  XNOR U2247 ( .A(n1239), .B(n1238), .Z(N6164) );
  XOR U2248 ( .A(n1258), .B(n1257), .Z(n1238) );
  XNOR U2249 ( .A(n1273), .B(n1274), .Z(n1257) );
  XNOR U2250 ( .A(n1268), .B(n1269), .Z(n1274) );
  XNOR U2251 ( .A(n1270), .B(n1271), .Z(n1269) );
  XNOR U2252 ( .A(y[916]), .B(x[916]), .Z(n1271) );
  XNOR U2253 ( .A(y[917]), .B(x[917]), .Z(n1270) );
  XNOR U2254 ( .A(y[915]), .B(x[915]), .Z(n1268) );
  XNOR U2255 ( .A(n1262), .B(n1263), .Z(n1273) );
  XNOR U2256 ( .A(y[912]), .B(x[912]), .Z(n1263) );
  XNOR U2257 ( .A(n1264), .B(n1265), .Z(n1262) );
  XNOR U2258 ( .A(y[913]), .B(x[913]), .Z(n1265) );
  XNOR U2259 ( .A(y[914]), .B(x[914]), .Z(n1264) );
  XNOR U2260 ( .A(n1255), .B(n1254), .Z(n1258) );
  XNOR U2261 ( .A(n1250), .B(n1251), .Z(n1254) );
  XNOR U2262 ( .A(y[909]), .B(x[909]), .Z(n1251) );
  XNOR U2263 ( .A(n1252), .B(n1253), .Z(n1250) );
  XNOR U2264 ( .A(y[910]), .B(x[910]), .Z(n1253) );
  XNOR U2265 ( .A(y[911]), .B(x[911]), .Z(n1252) );
  XNOR U2266 ( .A(n1244), .B(n1245), .Z(n1255) );
  XNOR U2267 ( .A(y[906]), .B(x[906]), .Z(n1245) );
  XNOR U2268 ( .A(n1246), .B(n1247), .Z(n1244) );
  XNOR U2269 ( .A(y[907]), .B(x[907]), .Z(n1247) );
  XNOR U2270 ( .A(y[908]), .B(x[908]), .Z(n1246) );
  XOR U2271 ( .A(n1220), .B(n1221), .Z(n1239) );
  XNOR U2272 ( .A(n1236), .B(n1237), .Z(n1221) );
  XNOR U2273 ( .A(n1231), .B(n1232), .Z(n1237) );
  XNOR U2274 ( .A(n1233), .B(n1234), .Z(n1232) );
  XNOR U2275 ( .A(y[904]), .B(x[904]), .Z(n1234) );
  XNOR U2276 ( .A(y[905]), .B(x[905]), .Z(n1233) );
  XNOR U2277 ( .A(y[903]), .B(x[903]), .Z(n1231) );
  XNOR U2278 ( .A(n1225), .B(n1226), .Z(n1236) );
  XNOR U2279 ( .A(y[900]), .B(x[900]), .Z(n1226) );
  XNOR U2280 ( .A(n1227), .B(n1228), .Z(n1225) );
  XNOR U2281 ( .A(y[901]), .B(x[901]), .Z(n1228) );
  XNOR U2282 ( .A(y[902]), .B(x[902]), .Z(n1227) );
  XOR U2283 ( .A(n1219), .B(n1218), .Z(n1220) );
  XNOR U2284 ( .A(n1214), .B(n1215), .Z(n1218) );
  XNOR U2285 ( .A(y[897]), .B(x[897]), .Z(n1215) );
  XNOR U2286 ( .A(n1216), .B(n1217), .Z(n1214) );
  XNOR U2287 ( .A(y[898]), .B(x[898]), .Z(n1217) );
  XNOR U2288 ( .A(y[899]), .B(x[899]), .Z(n1216) );
  XNOR U2289 ( .A(n1208), .B(n1209), .Z(n1219) );
  XNOR U2290 ( .A(y[894]), .B(x[894]), .Z(n1209) );
  XNOR U2291 ( .A(n1210), .B(n1211), .Z(n1208) );
  XNOR U2292 ( .A(y[895]), .B(x[895]), .Z(n1211) );
  XNOR U2293 ( .A(y[896]), .B(x[896]), .Z(n1210) );
  NAND U2294 ( .A(n1275), .B(n1276), .Z(N6158) );
  NANDN U2295 ( .A(n1277), .B(n1278), .Z(n1276) );
  OR U2296 ( .A(n1279), .B(n1280), .Z(n1278) );
  NAND U2297 ( .A(n1279), .B(n1280), .Z(n1275) );
  XOR U2298 ( .A(n1279), .B(n1281), .Z(N6157) );
  XNOR U2299 ( .A(n1277), .B(n1280), .Z(n1281) );
  AND U2300 ( .A(n1282), .B(n1283), .Z(n1280) );
  NANDN U2301 ( .A(n1284), .B(n1285), .Z(n1283) );
  NANDN U2302 ( .A(n1286), .B(n1287), .Z(n1285) );
  NANDN U2303 ( .A(n1287), .B(n1286), .Z(n1282) );
  NAND U2304 ( .A(n1288), .B(n1289), .Z(n1277) );
  NANDN U2305 ( .A(n1290), .B(n1291), .Z(n1289) );
  OR U2306 ( .A(n1292), .B(n1293), .Z(n1291) );
  NAND U2307 ( .A(n1293), .B(n1292), .Z(n1288) );
  AND U2308 ( .A(n1294), .B(n1295), .Z(n1279) );
  NANDN U2309 ( .A(n1296), .B(n1297), .Z(n1295) );
  NANDN U2310 ( .A(n1298), .B(n1299), .Z(n1297) );
  NANDN U2311 ( .A(n1299), .B(n1298), .Z(n1294) );
  XOR U2312 ( .A(n1293), .B(n1300), .Z(N6156) );
  XOR U2313 ( .A(n1290), .B(n1292), .Z(n1300) );
  XNOR U2314 ( .A(n1286), .B(n1301), .Z(n1292) );
  XNOR U2315 ( .A(n1284), .B(n1287), .Z(n1301) );
  NAND U2316 ( .A(n1302), .B(n1303), .Z(n1287) );
  NAND U2317 ( .A(n1304), .B(n1305), .Z(n1303) );
  OR U2318 ( .A(n1306), .B(n1307), .Z(n1304) );
  NANDN U2319 ( .A(n1308), .B(n1306), .Z(n1302) );
  IV U2320 ( .A(n1307), .Z(n1308) );
  NAND U2321 ( .A(n1309), .B(n1310), .Z(n1284) );
  NAND U2322 ( .A(n1311), .B(n1312), .Z(n1310) );
  NANDN U2323 ( .A(n1313), .B(n1314), .Z(n1311) );
  NANDN U2324 ( .A(n1314), .B(n1313), .Z(n1309) );
  AND U2325 ( .A(n1315), .B(n1316), .Z(n1286) );
  NAND U2326 ( .A(n1317), .B(n1318), .Z(n1316) );
  OR U2327 ( .A(n1319), .B(n1320), .Z(n1317) );
  NANDN U2328 ( .A(n1321), .B(n1319), .Z(n1315) );
  NAND U2329 ( .A(n1322), .B(n1323), .Z(n1290) );
  NANDN U2330 ( .A(n1324), .B(n1325), .Z(n1323) );
  OR U2331 ( .A(n1326), .B(n1327), .Z(n1325) );
  NANDN U2332 ( .A(n1328), .B(n1326), .Z(n1322) );
  IV U2333 ( .A(n1327), .Z(n1328) );
  XNOR U2334 ( .A(n1298), .B(n1329), .Z(n1293) );
  XNOR U2335 ( .A(n1296), .B(n1299), .Z(n1329) );
  NAND U2336 ( .A(n1330), .B(n1331), .Z(n1299) );
  NAND U2337 ( .A(n1332), .B(n1333), .Z(n1331) );
  OR U2338 ( .A(n1334), .B(n1335), .Z(n1332) );
  NANDN U2339 ( .A(n1336), .B(n1334), .Z(n1330) );
  IV U2340 ( .A(n1335), .Z(n1336) );
  NAND U2341 ( .A(n1337), .B(n1338), .Z(n1296) );
  NAND U2342 ( .A(n1339), .B(n1340), .Z(n1338) );
  NANDN U2343 ( .A(n1341), .B(n1342), .Z(n1339) );
  NANDN U2344 ( .A(n1342), .B(n1341), .Z(n1337) );
  AND U2345 ( .A(n1343), .B(n1344), .Z(n1298) );
  NAND U2346 ( .A(n1345), .B(n1346), .Z(n1344) );
  OR U2347 ( .A(n1347), .B(n1348), .Z(n1345) );
  NANDN U2348 ( .A(n1349), .B(n1347), .Z(n1343) );
  XNOR U2349 ( .A(n1324), .B(n1350), .Z(N6155) );
  XOR U2350 ( .A(n1326), .B(n1327), .Z(n1350) );
  XNOR U2351 ( .A(n1340), .B(n1351), .Z(n1327) );
  XOR U2352 ( .A(n1341), .B(n1342), .Z(n1351) );
  XOR U2353 ( .A(n1347), .B(n1352), .Z(n1342) );
  XOR U2354 ( .A(n1346), .B(n1349), .Z(n1352) );
  IV U2355 ( .A(n1348), .Z(n1349) );
  NAND U2356 ( .A(n1353), .B(n1354), .Z(n1348) );
  OR U2357 ( .A(n1355), .B(n1356), .Z(n1354) );
  OR U2358 ( .A(n1357), .B(n1358), .Z(n1353) );
  NAND U2359 ( .A(n1359), .B(n1360), .Z(n1346) );
  OR U2360 ( .A(n1361), .B(n1362), .Z(n1360) );
  OR U2361 ( .A(n1363), .B(n1364), .Z(n1359) );
  NOR U2362 ( .A(n1365), .B(n1366), .Z(n1347) );
  ANDN U2363 ( .B(n1367), .A(n1368), .Z(n1341) );
  XNOR U2364 ( .A(n1334), .B(n1369), .Z(n1340) );
  XNOR U2365 ( .A(n1333), .B(n1335), .Z(n1369) );
  NAND U2366 ( .A(n1370), .B(n1371), .Z(n1335) );
  OR U2367 ( .A(n1372), .B(n1373), .Z(n1371) );
  OR U2368 ( .A(n1374), .B(n1375), .Z(n1370) );
  NAND U2369 ( .A(n1376), .B(n1377), .Z(n1333) );
  OR U2370 ( .A(n1378), .B(n1379), .Z(n1377) );
  OR U2371 ( .A(n1380), .B(n1381), .Z(n1376) );
  ANDN U2372 ( .B(n1382), .A(n1383), .Z(n1334) );
  IV U2373 ( .A(n1384), .Z(n1382) );
  ANDN U2374 ( .B(n1385), .A(n1386), .Z(n1326) );
  XOR U2375 ( .A(n1312), .B(n1387), .Z(n1324) );
  XOR U2376 ( .A(n1313), .B(n1314), .Z(n1387) );
  XOR U2377 ( .A(n1319), .B(n1388), .Z(n1314) );
  XOR U2378 ( .A(n1318), .B(n1321), .Z(n1388) );
  IV U2379 ( .A(n1320), .Z(n1321) );
  NAND U2380 ( .A(n1389), .B(n1390), .Z(n1320) );
  OR U2381 ( .A(n1391), .B(n1392), .Z(n1390) );
  OR U2382 ( .A(n1393), .B(n1394), .Z(n1389) );
  NAND U2383 ( .A(n1395), .B(n1396), .Z(n1318) );
  OR U2384 ( .A(n1397), .B(n1398), .Z(n1396) );
  OR U2385 ( .A(n1399), .B(n1400), .Z(n1395) );
  NOR U2386 ( .A(n1401), .B(n1402), .Z(n1319) );
  ANDN U2387 ( .B(n1403), .A(n1404), .Z(n1313) );
  IV U2388 ( .A(n1405), .Z(n1403) );
  XNOR U2389 ( .A(n1306), .B(n1406), .Z(n1312) );
  XNOR U2390 ( .A(n1305), .B(n1307), .Z(n1406) );
  NAND U2391 ( .A(n1407), .B(n1408), .Z(n1307) );
  OR U2392 ( .A(n1409), .B(n1410), .Z(n1408) );
  OR U2393 ( .A(n1411), .B(n1412), .Z(n1407) );
  NAND U2394 ( .A(n1413), .B(n1414), .Z(n1305) );
  OR U2395 ( .A(n1415), .B(n1416), .Z(n1414) );
  OR U2396 ( .A(n1417), .B(n1418), .Z(n1413) );
  ANDN U2397 ( .B(n1419), .A(n1420), .Z(n1306) );
  IV U2398 ( .A(n1421), .Z(n1419) );
  XNOR U2399 ( .A(n1386), .B(n1385), .Z(N6154) );
  XOR U2400 ( .A(n1405), .B(n1404), .Z(n1385) );
  XNOR U2401 ( .A(n1420), .B(n1421), .Z(n1404) );
  XNOR U2402 ( .A(n1415), .B(n1416), .Z(n1421) );
  XNOR U2403 ( .A(n1417), .B(n1418), .Z(n1416) );
  XNOR U2404 ( .A(y[892]), .B(x[892]), .Z(n1418) );
  XNOR U2405 ( .A(y[893]), .B(x[893]), .Z(n1417) );
  XNOR U2406 ( .A(y[891]), .B(x[891]), .Z(n1415) );
  XNOR U2407 ( .A(n1409), .B(n1410), .Z(n1420) );
  XNOR U2408 ( .A(y[888]), .B(x[888]), .Z(n1410) );
  XNOR U2409 ( .A(n1411), .B(n1412), .Z(n1409) );
  XNOR U2410 ( .A(y[889]), .B(x[889]), .Z(n1412) );
  XNOR U2411 ( .A(y[890]), .B(x[890]), .Z(n1411) );
  XNOR U2412 ( .A(n1402), .B(n1401), .Z(n1405) );
  XNOR U2413 ( .A(n1397), .B(n1398), .Z(n1401) );
  XNOR U2414 ( .A(y[885]), .B(x[885]), .Z(n1398) );
  XNOR U2415 ( .A(n1399), .B(n1400), .Z(n1397) );
  XNOR U2416 ( .A(y[886]), .B(x[886]), .Z(n1400) );
  XNOR U2417 ( .A(y[887]), .B(x[887]), .Z(n1399) );
  XNOR U2418 ( .A(n1391), .B(n1392), .Z(n1402) );
  XNOR U2419 ( .A(y[882]), .B(x[882]), .Z(n1392) );
  XNOR U2420 ( .A(n1393), .B(n1394), .Z(n1391) );
  XNOR U2421 ( .A(y[883]), .B(x[883]), .Z(n1394) );
  XNOR U2422 ( .A(y[884]), .B(x[884]), .Z(n1393) );
  XOR U2423 ( .A(n1367), .B(n1368), .Z(n1386) );
  XNOR U2424 ( .A(n1383), .B(n1384), .Z(n1368) );
  XNOR U2425 ( .A(n1378), .B(n1379), .Z(n1384) );
  XNOR U2426 ( .A(n1380), .B(n1381), .Z(n1379) );
  XNOR U2427 ( .A(y[880]), .B(x[880]), .Z(n1381) );
  XNOR U2428 ( .A(y[881]), .B(x[881]), .Z(n1380) );
  XNOR U2429 ( .A(y[879]), .B(x[879]), .Z(n1378) );
  XNOR U2430 ( .A(n1372), .B(n1373), .Z(n1383) );
  XNOR U2431 ( .A(y[876]), .B(x[876]), .Z(n1373) );
  XNOR U2432 ( .A(n1374), .B(n1375), .Z(n1372) );
  XNOR U2433 ( .A(y[877]), .B(x[877]), .Z(n1375) );
  XNOR U2434 ( .A(y[878]), .B(x[878]), .Z(n1374) );
  XOR U2435 ( .A(n1366), .B(n1365), .Z(n1367) );
  XNOR U2436 ( .A(n1361), .B(n1362), .Z(n1365) );
  XNOR U2437 ( .A(y[873]), .B(x[873]), .Z(n1362) );
  XNOR U2438 ( .A(n1363), .B(n1364), .Z(n1361) );
  XNOR U2439 ( .A(y[874]), .B(x[874]), .Z(n1364) );
  XNOR U2440 ( .A(y[875]), .B(x[875]), .Z(n1363) );
  XNOR U2441 ( .A(n1355), .B(n1356), .Z(n1366) );
  XNOR U2442 ( .A(y[870]), .B(x[870]), .Z(n1356) );
  XNOR U2443 ( .A(n1357), .B(n1358), .Z(n1355) );
  XNOR U2444 ( .A(y[871]), .B(x[871]), .Z(n1358) );
  XNOR U2445 ( .A(y[872]), .B(x[872]), .Z(n1357) );
  NAND U2446 ( .A(n1422), .B(n1423), .Z(N6148) );
  NANDN U2447 ( .A(n1424), .B(n1425), .Z(n1423) );
  OR U2448 ( .A(n1426), .B(n1427), .Z(n1425) );
  NAND U2449 ( .A(n1426), .B(n1427), .Z(n1422) );
  XOR U2450 ( .A(n1426), .B(n1428), .Z(N6147) );
  XNOR U2451 ( .A(n1424), .B(n1427), .Z(n1428) );
  AND U2452 ( .A(n1429), .B(n1430), .Z(n1427) );
  NANDN U2453 ( .A(n1431), .B(n1432), .Z(n1430) );
  NANDN U2454 ( .A(n1433), .B(n1434), .Z(n1432) );
  NANDN U2455 ( .A(n1434), .B(n1433), .Z(n1429) );
  NAND U2456 ( .A(n1435), .B(n1436), .Z(n1424) );
  NANDN U2457 ( .A(n1437), .B(n1438), .Z(n1436) );
  OR U2458 ( .A(n1439), .B(n1440), .Z(n1438) );
  NAND U2459 ( .A(n1440), .B(n1439), .Z(n1435) );
  AND U2460 ( .A(n1441), .B(n1442), .Z(n1426) );
  NANDN U2461 ( .A(n1443), .B(n1444), .Z(n1442) );
  NANDN U2462 ( .A(n1445), .B(n1446), .Z(n1444) );
  NANDN U2463 ( .A(n1446), .B(n1445), .Z(n1441) );
  XOR U2464 ( .A(n1440), .B(n1447), .Z(N6146) );
  XOR U2465 ( .A(n1437), .B(n1439), .Z(n1447) );
  XNOR U2466 ( .A(n1433), .B(n1448), .Z(n1439) );
  XNOR U2467 ( .A(n1431), .B(n1434), .Z(n1448) );
  NAND U2468 ( .A(n1449), .B(n1450), .Z(n1434) );
  NAND U2469 ( .A(n1451), .B(n1452), .Z(n1450) );
  OR U2470 ( .A(n1453), .B(n1454), .Z(n1451) );
  NANDN U2471 ( .A(n1455), .B(n1453), .Z(n1449) );
  IV U2472 ( .A(n1454), .Z(n1455) );
  NAND U2473 ( .A(n1456), .B(n1457), .Z(n1431) );
  NAND U2474 ( .A(n1458), .B(n1459), .Z(n1457) );
  NANDN U2475 ( .A(n1460), .B(n1461), .Z(n1458) );
  NANDN U2476 ( .A(n1461), .B(n1460), .Z(n1456) );
  AND U2477 ( .A(n1462), .B(n1463), .Z(n1433) );
  NAND U2478 ( .A(n1464), .B(n1465), .Z(n1463) );
  OR U2479 ( .A(n1466), .B(n1467), .Z(n1464) );
  NANDN U2480 ( .A(n1468), .B(n1466), .Z(n1462) );
  NAND U2481 ( .A(n1469), .B(n1470), .Z(n1437) );
  NANDN U2482 ( .A(n1471), .B(n1472), .Z(n1470) );
  OR U2483 ( .A(n1473), .B(n1474), .Z(n1472) );
  NANDN U2484 ( .A(n1475), .B(n1473), .Z(n1469) );
  IV U2485 ( .A(n1474), .Z(n1475) );
  XNOR U2486 ( .A(n1445), .B(n1476), .Z(n1440) );
  XNOR U2487 ( .A(n1443), .B(n1446), .Z(n1476) );
  NAND U2488 ( .A(n1477), .B(n1478), .Z(n1446) );
  NAND U2489 ( .A(n1479), .B(n1480), .Z(n1478) );
  OR U2490 ( .A(n1481), .B(n1482), .Z(n1479) );
  NANDN U2491 ( .A(n1483), .B(n1481), .Z(n1477) );
  IV U2492 ( .A(n1482), .Z(n1483) );
  NAND U2493 ( .A(n1484), .B(n1485), .Z(n1443) );
  NAND U2494 ( .A(n1486), .B(n1487), .Z(n1485) );
  NANDN U2495 ( .A(n1488), .B(n1489), .Z(n1486) );
  NANDN U2496 ( .A(n1489), .B(n1488), .Z(n1484) );
  AND U2497 ( .A(n1490), .B(n1491), .Z(n1445) );
  NAND U2498 ( .A(n1492), .B(n1493), .Z(n1491) );
  OR U2499 ( .A(n1494), .B(n1495), .Z(n1492) );
  NANDN U2500 ( .A(n1496), .B(n1494), .Z(n1490) );
  XNOR U2501 ( .A(n1471), .B(n1497), .Z(N6145) );
  XOR U2502 ( .A(n1473), .B(n1474), .Z(n1497) );
  XNOR U2503 ( .A(n1487), .B(n1498), .Z(n1474) );
  XOR U2504 ( .A(n1488), .B(n1489), .Z(n1498) );
  XOR U2505 ( .A(n1494), .B(n1499), .Z(n1489) );
  XOR U2506 ( .A(n1493), .B(n1496), .Z(n1499) );
  IV U2507 ( .A(n1495), .Z(n1496) );
  NAND U2508 ( .A(n1500), .B(n1501), .Z(n1495) );
  OR U2509 ( .A(n1502), .B(n1503), .Z(n1501) );
  OR U2510 ( .A(n1504), .B(n1505), .Z(n1500) );
  NAND U2511 ( .A(n1506), .B(n1507), .Z(n1493) );
  OR U2512 ( .A(n1508), .B(n1509), .Z(n1507) );
  OR U2513 ( .A(n1510), .B(n1511), .Z(n1506) );
  NOR U2514 ( .A(n1512), .B(n1513), .Z(n1494) );
  ANDN U2515 ( .B(n1514), .A(n1515), .Z(n1488) );
  XNOR U2516 ( .A(n1481), .B(n1516), .Z(n1487) );
  XNOR U2517 ( .A(n1480), .B(n1482), .Z(n1516) );
  NAND U2518 ( .A(n1517), .B(n1518), .Z(n1482) );
  OR U2519 ( .A(n1519), .B(n1520), .Z(n1518) );
  OR U2520 ( .A(n1521), .B(n1522), .Z(n1517) );
  NAND U2521 ( .A(n1523), .B(n1524), .Z(n1480) );
  OR U2522 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U2523 ( .A(n1527), .B(n1528), .Z(n1523) );
  ANDN U2524 ( .B(n1529), .A(n1530), .Z(n1481) );
  IV U2525 ( .A(n1531), .Z(n1529) );
  ANDN U2526 ( .B(n1532), .A(n1533), .Z(n1473) );
  XOR U2527 ( .A(n1459), .B(n1534), .Z(n1471) );
  XOR U2528 ( .A(n1460), .B(n1461), .Z(n1534) );
  XOR U2529 ( .A(n1466), .B(n1535), .Z(n1461) );
  XOR U2530 ( .A(n1465), .B(n1468), .Z(n1535) );
  IV U2531 ( .A(n1467), .Z(n1468) );
  NAND U2532 ( .A(n1536), .B(n1537), .Z(n1467) );
  OR U2533 ( .A(n1538), .B(n1539), .Z(n1537) );
  OR U2534 ( .A(n1540), .B(n1541), .Z(n1536) );
  NAND U2535 ( .A(n1542), .B(n1543), .Z(n1465) );
  OR U2536 ( .A(n1544), .B(n1545), .Z(n1543) );
  OR U2537 ( .A(n1546), .B(n1547), .Z(n1542) );
  NOR U2538 ( .A(n1548), .B(n1549), .Z(n1466) );
  ANDN U2539 ( .B(n1550), .A(n1551), .Z(n1460) );
  IV U2540 ( .A(n1552), .Z(n1550) );
  XNOR U2541 ( .A(n1453), .B(n1553), .Z(n1459) );
  XNOR U2542 ( .A(n1452), .B(n1454), .Z(n1553) );
  NAND U2543 ( .A(n1554), .B(n1555), .Z(n1454) );
  OR U2544 ( .A(n1556), .B(n1557), .Z(n1555) );
  OR U2545 ( .A(n1558), .B(n1559), .Z(n1554) );
  NAND U2546 ( .A(n1560), .B(n1561), .Z(n1452) );
  OR U2547 ( .A(n1562), .B(n1563), .Z(n1561) );
  OR U2548 ( .A(n1564), .B(n1565), .Z(n1560) );
  ANDN U2549 ( .B(n1566), .A(n1567), .Z(n1453) );
  IV U2550 ( .A(n1568), .Z(n1566) );
  XNOR U2551 ( .A(n1533), .B(n1532), .Z(N6144) );
  XOR U2552 ( .A(n1552), .B(n1551), .Z(n1532) );
  XNOR U2553 ( .A(n1567), .B(n1568), .Z(n1551) );
  XNOR U2554 ( .A(n1562), .B(n1563), .Z(n1568) );
  XNOR U2555 ( .A(n1564), .B(n1565), .Z(n1563) );
  XNOR U2556 ( .A(y[868]), .B(x[868]), .Z(n1565) );
  XNOR U2557 ( .A(y[869]), .B(x[869]), .Z(n1564) );
  XNOR U2558 ( .A(y[867]), .B(x[867]), .Z(n1562) );
  XNOR U2559 ( .A(n1556), .B(n1557), .Z(n1567) );
  XNOR U2560 ( .A(y[864]), .B(x[864]), .Z(n1557) );
  XNOR U2561 ( .A(n1558), .B(n1559), .Z(n1556) );
  XNOR U2562 ( .A(y[865]), .B(x[865]), .Z(n1559) );
  XNOR U2563 ( .A(y[866]), .B(x[866]), .Z(n1558) );
  XNOR U2564 ( .A(n1549), .B(n1548), .Z(n1552) );
  XNOR U2565 ( .A(n1544), .B(n1545), .Z(n1548) );
  XNOR U2566 ( .A(y[861]), .B(x[861]), .Z(n1545) );
  XNOR U2567 ( .A(n1546), .B(n1547), .Z(n1544) );
  XNOR U2568 ( .A(y[862]), .B(x[862]), .Z(n1547) );
  XNOR U2569 ( .A(y[863]), .B(x[863]), .Z(n1546) );
  XNOR U2570 ( .A(n1538), .B(n1539), .Z(n1549) );
  XNOR U2571 ( .A(y[858]), .B(x[858]), .Z(n1539) );
  XNOR U2572 ( .A(n1540), .B(n1541), .Z(n1538) );
  XNOR U2573 ( .A(y[859]), .B(x[859]), .Z(n1541) );
  XNOR U2574 ( .A(y[860]), .B(x[860]), .Z(n1540) );
  XOR U2575 ( .A(n1514), .B(n1515), .Z(n1533) );
  XNOR U2576 ( .A(n1530), .B(n1531), .Z(n1515) );
  XNOR U2577 ( .A(n1525), .B(n1526), .Z(n1531) );
  XNOR U2578 ( .A(n1527), .B(n1528), .Z(n1526) );
  XNOR U2579 ( .A(y[856]), .B(x[856]), .Z(n1528) );
  XNOR U2580 ( .A(y[857]), .B(x[857]), .Z(n1527) );
  XNOR U2581 ( .A(y[855]), .B(x[855]), .Z(n1525) );
  XNOR U2582 ( .A(n1519), .B(n1520), .Z(n1530) );
  XNOR U2583 ( .A(y[852]), .B(x[852]), .Z(n1520) );
  XNOR U2584 ( .A(n1521), .B(n1522), .Z(n1519) );
  XNOR U2585 ( .A(y[853]), .B(x[853]), .Z(n1522) );
  XNOR U2586 ( .A(y[854]), .B(x[854]), .Z(n1521) );
  XOR U2587 ( .A(n1513), .B(n1512), .Z(n1514) );
  XNOR U2588 ( .A(n1508), .B(n1509), .Z(n1512) );
  XNOR U2589 ( .A(y[849]), .B(x[849]), .Z(n1509) );
  XNOR U2590 ( .A(n1510), .B(n1511), .Z(n1508) );
  XNOR U2591 ( .A(y[850]), .B(x[850]), .Z(n1511) );
  XNOR U2592 ( .A(y[851]), .B(x[851]), .Z(n1510) );
  XNOR U2593 ( .A(n1502), .B(n1503), .Z(n1513) );
  XNOR U2594 ( .A(y[846]), .B(x[846]), .Z(n1503) );
  XNOR U2595 ( .A(n1504), .B(n1505), .Z(n1502) );
  XNOR U2596 ( .A(y[847]), .B(x[847]), .Z(n1505) );
  XNOR U2597 ( .A(y[848]), .B(x[848]), .Z(n1504) );
  NAND U2598 ( .A(n1569), .B(n1570), .Z(N6138) );
  NANDN U2599 ( .A(n1571), .B(n1572), .Z(n1570) );
  OR U2600 ( .A(n1573), .B(n1574), .Z(n1572) );
  NAND U2601 ( .A(n1573), .B(n1574), .Z(n1569) );
  XOR U2602 ( .A(n1573), .B(n1575), .Z(N6137) );
  XNOR U2603 ( .A(n1571), .B(n1574), .Z(n1575) );
  AND U2604 ( .A(n1576), .B(n1577), .Z(n1574) );
  NANDN U2605 ( .A(n1578), .B(n1579), .Z(n1577) );
  NANDN U2606 ( .A(n1580), .B(n1581), .Z(n1579) );
  NANDN U2607 ( .A(n1581), .B(n1580), .Z(n1576) );
  NAND U2608 ( .A(n1582), .B(n1583), .Z(n1571) );
  NANDN U2609 ( .A(n1584), .B(n1585), .Z(n1583) );
  OR U2610 ( .A(n1586), .B(n1587), .Z(n1585) );
  NAND U2611 ( .A(n1587), .B(n1586), .Z(n1582) );
  AND U2612 ( .A(n1588), .B(n1589), .Z(n1573) );
  NANDN U2613 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U2614 ( .A(n1592), .B(n1593), .Z(n1591) );
  NANDN U2615 ( .A(n1593), .B(n1592), .Z(n1588) );
  XOR U2616 ( .A(n1587), .B(n1594), .Z(N6136) );
  XOR U2617 ( .A(n1584), .B(n1586), .Z(n1594) );
  XNOR U2618 ( .A(n1580), .B(n1595), .Z(n1586) );
  XNOR U2619 ( .A(n1578), .B(n1581), .Z(n1595) );
  NAND U2620 ( .A(n1596), .B(n1597), .Z(n1581) );
  NAND U2621 ( .A(n1598), .B(n1599), .Z(n1597) );
  OR U2622 ( .A(n1600), .B(n1601), .Z(n1598) );
  NANDN U2623 ( .A(n1602), .B(n1600), .Z(n1596) );
  IV U2624 ( .A(n1601), .Z(n1602) );
  NAND U2625 ( .A(n1603), .B(n1604), .Z(n1578) );
  NAND U2626 ( .A(n1605), .B(n1606), .Z(n1604) );
  NANDN U2627 ( .A(n1607), .B(n1608), .Z(n1605) );
  NANDN U2628 ( .A(n1608), .B(n1607), .Z(n1603) );
  AND U2629 ( .A(n1609), .B(n1610), .Z(n1580) );
  NAND U2630 ( .A(n1611), .B(n1612), .Z(n1610) );
  OR U2631 ( .A(n1613), .B(n1614), .Z(n1611) );
  NANDN U2632 ( .A(n1615), .B(n1613), .Z(n1609) );
  NAND U2633 ( .A(n1616), .B(n1617), .Z(n1584) );
  NANDN U2634 ( .A(n1618), .B(n1619), .Z(n1617) );
  OR U2635 ( .A(n1620), .B(n1621), .Z(n1619) );
  NANDN U2636 ( .A(n1622), .B(n1620), .Z(n1616) );
  IV U2637 ( .A(n1621), .Z(n1622) );
  XNOR U2638 ( .A(n1592), .B(n1623), .Z(n1587) );
  XNOR U2639 ( .A(n1590), .B(n1593), .Z(n1623) );
  NAND U2640 ( .A(n1624), .B(n1625), .Z(n1593) );
  NAND U2641 ( .A(n1626), .B(n1627), .Z(n1625) );
  OR U2642 ( .A(n1628), .B(n1629), .Z(n1626) );
  NANDN U2643 ( .A(n1630), .B(n1628), .Z(n1624) );
  IV U2644 ( .A(n1629), .Z(n1630) );
  NAND U2645 ( .A(n1631), .B(n1632), .Z(n1590) );
  NAND U2646 ( .A(n1633), .B(n1634), .Z(n1632) );
  NANDN U2647 ( .A(n1635), .B(n1636), .Z(n1633) );
  NANDN U2648 ( .A(n1636), .B(n1635), .Z(n1631) );
  AND U2649 ( .A(n1637), .B(n1638), .Z(n1592) );
  NAND U2650 ( .A(n1639), .B(n1640), .Z(n1638) );
  OR U2651 ( .A(n1641), .B(n1642), .Z(n1639) );
  NANDN U2652 ( .A(n1643), .B(n1641), .Z(n1637) );
  XNOR U2653 ( .A(n1618), .B(n1644), .Z(N6135) );
  XOR U2654 ( .A(n1620), .B(n1621), .Z(n1644) );
  XNOR U2655 ( .A(n1634), .B(n1645), .Z(n1621) );
  XOR U2656 ( .A(n1635), .B(n1636), .Z(n1645) );
  XOR U2657 ( .A(n1641), .B(n1646), .Z(n1636) );
  XOR U2658 ( .A(n1640), .B(n1643), .Z(n1646) );
  IV U2659 ( .A(n1642), .Z(n1643) );
  NAND U2660 ( .A(n1647), .B(n1648), .Z(n1642) );
  OR U2661 ( .A(n1649), .B(n1650), .Z(n1648) );
  OR U2662 ( .A(n1651), .B(n1652), .Z(n1647) );
  NAND U2663 ( .A(n1653), .B(n1654), .Z(n1640) );
  OR U2664 ( .A(n1655), .B(n1656), .Z(n1654) );
  OR U2665 ( .A(n1657), .B(n1658), .Z(n1653) );
  NOR U2666 ( .A(n1659), .B(n1660), .Z(n1641) );
  ANDN U2667 ( .B(n1661), .A(n1662), .Z(n1635) );
  XNOR U2668 ( .A(n1628), .B(n1663), .Z(n1634) );
  XNOR U2669 ( .A(n1627), .B(n1629), .Z(n1663) );
  NAND U2670 ( .A(n1664), .B(n1665), .Z(n1629) );
  OR U2671 ( .A(n1666), .B(n1667), .Z(n1665) );
  OR U2672 ( .A(n1668), .B(n1669), .Z(n1664) );
  NAND U2673 ( .A(n1670), .B(n1671), .Z(n1627) );
  OR U2674 ( .A(n1672), .B(n1673), .Z(n1671) );
  OR U2675 ( .A(n1674), .B(n1675), .Z(n1670) );
  ANDN U2676 ( .B(n1676), .A(n1677), .Z(n1628) );
  IV U2677 ( .A(n1678), .Z(n1676) );
  ANDN U2678 ( .B(n1679), .A(n1680), .Z(n1620) );
  XOR U2679 ( .A(n1606), .B(n1681), .Z(n1618) );
  XOR U2680 ( .A(n1607), .B(n1608), .Z(n1681) );
  XOR U2681 ( .A(n1613), .B(n1682), .Z(n1608) );
  XOR U2682 ( .A(n1612), .B(n1615), .Z(n1682) );
  IV U2683 ( .A(n1614), .Z(n1615) );
  NAND U2684 ( .A(n1683), .B(n1684), .Z(n1614) );
  OR U2685 ( .A(n1685), .B(n1686), .Z(n1684) );
  OR U2686 ( .A(n1687), .B(n1688), .Z(n1683) );
  NAND U2687 ( .A(n1689), .B(n1690), .Z(n1612) );
  OR U2688 ( .A(n1691), .B(n1692), .Z(n1690) );
  OR U2689 ( .A(n1693), .B(n1694), .Z(n1689) );
  NOR U2690 ( .A(n1695), .B(n1696), .Z(n1613) );
  ANDN U2691 ( .B(n1697), .A(n1698), .Z(n1607) );
  IV U2692 ( .A(n1699), .Z(n1697) );
  XNOR U2693 ( .A(n1600), .B(n1700), .Z(n1606) );
  XNOR U2694 ( .A(n1599), .B(n1601), .Z(n1700) );
  NAND U2695 ( .A(n1701), .B(n1702), .Z(n1601) );
  OR U2696 ( .A(n1703), .B(n1704), .Z(n1702) );
  OR U2697 ( .A(n1705), .B(n1706), .Z(n1701) );
  NAND U2698 ( .A(n1707), .B(n1708), .Z(n1599) );
  OR U2699 ( .A(n1709), .B(n1710), .Z(n1708) );
  OR U2700 ( .A(n1711), .B(n1712), .Z(n1707) );
  ANDN U2701 ( .B(n1713), .A(n1714), .Z(n1600) );
  IV U2702 ( .A(n1715), .Z(n1713) );
  XNOR U2703 ( .A(n1680), .B(n1679), .Z(N6134) );
  XOR U2704 ( .A(n1699), .B(n1698), .Z(n1679) );
  XNOR U2705 ( .A(n1714), .B(n1715), .Z(n1698) );
  XNOR U2706 ( .A(n1709), .B(n1710), .Z(n1715) );
  XNOR U2707 ( .A(n1711), .B(n1712), .Z(n1710) );
  XNOR U2708 ( .A(y[844]), .B(x[844]), .Z(n1712) );
  XNOR U2709 ( .A(y[845]), .B(x[845]), .Z(n1711) );
  XNOR U2710 ( .A(y[843]), .B(x[843]), .Z(n1709) );
  XNOR U2711 ( .A(n1703), .B(n1704), .Z(n1714) );
  XNOR U2712 ( .A(y[840]), .B(x[840]), .Z(n1704) );
  XNOR U2713 ( .A(n1705), .B(n1706), .Z(n1703) );
  XNOR U2714 ( .A(y[841]), .B(x[841]), .Z(n1706) );
  XNOR U2715 ( .A(y[842]), .B(x[842]), .Z(n1705) );
  XNOR U2716 ( .A(n1696), .B(n1695), .Z(n1699) );
  XNOR U2717 ( .A(n1691), .B(n1692), .Z(n1695) );
  XNOR U2718 ( .A(y[837]), .B(x[837]), .Z(n1692) );
  XNOR U2719 ( .A(n1693), .B(n1694), .Z(n1691) );
  XNOR U2720 ( .A(y[838]), .B(x[838]), .Z(n1694) );
  XNOR U2721 ( .A(y[839]), .B(x[839]), .Z(n1693) );
  XNOR U2722 ( .A(n1685), .B(n1686), .Z(n1696) );
  XNOR U2723 ( .A(y[834]), .B(x[834]), .Z(n1686) );
  XNOR U2724 ( .A(n1687), .B(n1688), .Z(n1685) );
  XNOR U2725 ( .A(y[835]), .B(x[835]), .Z(n1688) );
  XNOR U2726 ( .A(y[836]), .B(x[836]), .Z(n1687) );
  XOR U2727 ( .A(n1661), .B(n1662), .Z(n1680) );
  XNOR U2728 ( .A(n1677), .B(n1678), .Z(n1662) );
  XNOR U2729 ( .A(n1672), .B(n1673), .Z(n1678) );
  XNOR U2730 ( .A(n1674), .B(n1675), .Z(n1673) );
  XNOR U2731 ( .A(y[832]), .B(x[832]), .Z(n1675) );
  XNOR U2732 ( .A(y[833]), .B(x[833]), .Z(n1674) );
  XNOR U2733 ( .A(y[831]), .B(x[831]), .Z(n1672) );
  XNOR U2734 ( .A(n1666), .B(n1667), .Z(n1677) );
  XNOR U2735 ( .A(y[828]), .B(x[828]), .Z(n1667) );
  XNOR U2736 ( .A(n1668), .B(n1669), .Z(n1666) );
  XNOR U2737 ( .A(y[829]), .B(x[829]), .Z(n1669) );
  XNOR U2738 ( .A(y[830]), .B(x[830]), .Z(n1668) );
  XOR U2739 ( .A(n1660), .B(n1659), .Z(n1661) );
  XNOR U2740 ( .A(n1655), .B(n1656), .Z(n1659) );
  XNOR U2741 ( .A(y[825]), .B(x[825]), .Z(n1656) );
  XNOR U2742 ( .A(n1657), .B(n1658), .Z(n1655) );
  XNOR U2743 ( .A(y[826]), .B(x[826]), .Z(n1658) );
  XNOR U2744 ( .A(y[827]), .B(x[827]), .Z(n1657) );
  XNOR U2745 ( .A(n1649), .B(n1650), .Z(n1660) );
  XNOR U2746 ( .A(y[822]), .B(x[822]), .Z(n1650) );
  XNOR U2747 ( .A(n1651), .B(n1652), .Z(n1649) );
  XNOR U2748 ( .A(y[823]), .B(x[823]), .Z(n1652) );
  XNOR U2749 ( .A(y[824]), .B(x[824]), .Z(n1651) );
  NAND U2750 ( .A(n1716), .B(n1717), .Z(N6128) );
  NANDN U2751 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U2752 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U2753 ( .A(n1720), .B(n1721), .Z(n1716) );
  XOR U2754 ( .A(n1720), .B(n1722), .Z(N6127) );
  XNOR U2755 ( .A(n1718), .B(n1721), .Z(n1722) );
  AND U2756 ( .A(n1723), .B(n1724), .Z(n1721) );
  NANDN U2757 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U2758 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U2759 ( .A(n1728), .B(n1727), .Z(n1723) );
  NAND U2760 ( .A(n1729), .B(n1730), .Z(n1718) );
  NANDN U2761 ( .A(n1731), .B(n1732), .Z(n1730) );
  OR U2762 ( .A(n1733), .B(n1734), .Z(n1732) );
  NAND U2763 ( .A(n1734), .B(n1733), .Z(n1729) );
  AND U2764 ( .A(n1735), .B(n1736), .Z(n1720) );
  NANDN U2765 ( .A(n1737), .B(n1738), .Z(n1736) );
  NANDN U2766 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U2767 ( .A(n1740), .B(n1739), .Z(n1735) );
  XOR U2768 ( .A(n1734), .B(n1741), .Z(N6126) );
  XOR U2769 ( .A(n1731), .B(n1733), .Z(n1741) );
  XNOR U2770 ( .A(n1727), .B(n1742), .Z(n1733) );
  XNOR U2771 ( .A(n1725), .B(n1728), .Z(n1742) );
  NAND U2772 ( .A(n1743), .B(n1744), .Z(n1728) );
  NAND U2773 ( .A(n1745), .B(n1746), .Z(n1744) );
  OR U2774 ( .A(n1747), .B(n1748), .Z(n1745) );
  NANDN U2775 ( .A(n1749), .B(n1747), .Z(n1743) );
  IV U2776 ( .A(n1748), .Z(n1749) );
  NAND U2777 ( .A(n1750), .B(n1751), .Z(n1725) );
  NAND U2778 ( .A(n1752), .B(n1753), .Z(n1751) );
  NANDN U2779 ( .A(n1754), .B(n1755), .Z(n1752) );
  NANDN U2780 ( .A(n1755), .B(n1754), .Z(n1750) );
  AND U2781 ( .A(n1756), .B(n1757), .Z(n1727) );
  NAND U2782 ( .A(n1758), .B(n1759), .Z(n1757) );
  OR U2783 ( .A(n1760), .B(n1761), .Z(n1758) );
  NANDN U2784 ( .A(n1762), .B(n1760), .Z(n1756) );
  NAND U2785 ( .A(n1763), .B(n1764), .Z(n1731) );
  NANDN U2786 ( .A(n1765), .B(n1766), .Z(n1764) );
  OR U2787 ( .A(n1767), .B(n1768), .Z(n1766) );
  NANDN U2788 ( .A(n1769), .B(n1767), .Z(n1763) );
  IV U2789 ( .A(n1768), .Z(n1769) );
  XNOR U2790 ( .A(n1739), .B(n1770), .Z(n1734) );
  XNOR U2791 ( .A(n1737), .B(n1740), .Z(n1770) );
  NAND U2792 ( .A(n1771), .B(n1772), .Z(n1740) );
  NAND U2793 ( .A(n1773), .B(n1774), .Z(n1772) );
  OR U2794 ( .A(n1775), .B(n1776), .Z(n1773) );
  NANDN U2795 ( .A(n1777), .B(n1775), .Z(n1771) );
  IV U2796 ( .A(n1776), .Z(n1777) );
  NAND U2797 ( .A(n1778), .B(n1779), .Z(n1737) );
  NAND U2798 ( .A(n1780), .B(n1781), .Z(n1779) );
  NANDN U2799 ( .A(n1782), .B(n1783), .Z(n1780) );
  NANDN U2800 ( .A(n1783), .B(n1782), .Z(n1778) );
  AND U2801 ( .A(n1784), .B(n1785), .Z(n1739) );
  NAND U2802 ( .A(n1786), .B(n1787), .Z(n1785) );
  OR U2803 ( .A(n1788), .B(n1789), .Z(n1786) );
  NANDN U2804 ( .A(n1790), .B(n1788), .Z(n1784) );
  XNOR U2805 ( .A(n1765), .B(n1791), .Z(N6125) );
  XOR U2806 ( .A(n1767), .B(n1768), .Z(n1791) );
  XNOR U2807 ( .A(n1781), .B(n1792), .Z(n1768) );
  XOR U2808 ( .A(n1782), .B(n1783), .Z(n1792) );
  XOR U2809 ( .A(n1788), .B(n1793), .Z(n1783) );
  XOR U2810 ( .A(n1787), .B(n1790), .Z(n1793) );
  IV U2811 ( .A(n1789), .Z(n1790) );
  NAND U2812 ( .A(n1794), .B(n1795), .Z(n1789) );
  OR U2813 ( .A(n1796), .B(n1797), .Z(n1795) );
  OR U2814 ( .A(n1798), .B(n1799), .Z(n1794) );
  NAND U2815 ( .A(n1800), .B(n1801), .Z(n1787) );
  OR U2816 ( .A(n1802), .B(n1803), .Z(n1801) );
  OR U2817 ( .A(n1804), .B(n1805), .Z(n1800) );
  NOR U2818 ( .A(n1806), .B(n1807), .Z(n1788) );
  ANDN U2819 ( .B(n1808), .A(n1809), .Z(n1782) );
  XNOR U2820 ( .A(n1775), .B(n1810), .Z(n1781) );
  XNOR U2821 ( .A(n1774), .B(n1776), .Z(n1810) );
  NAND U2822 ( .A(n1811), .B(n1812), .Z(n1776) );
  OR U2823 ( .A(n1813), .B(n1814), .Z(n1812) );
  OR U2824 ( .A(n1815), .B(n1816), .Z(n1811) );
  NAND U2825 ( .A(n1817), .B(n1818), .Z(n1774) );
  OR U2826 ( .A(n1819), .B(n1820), .Z(n1818) );
  OR U2827 ( .A(n1821), .B(n1822), .Z(n1817) );
  ANDN U2828 ( .B(n1823), .A(n1824), .Z(n1775) );
  IV U2829 ( .A(n1825), .Z(n1823) );
  ANDN U2830 ( .B(n1826), .A(n1827), .Z(n1767) );
  XOR U2831 ( .A(n1753), .B(n1828), .Z(n1765) );
  XOR U2832 ( .A(n1754), .B(n1755), .Z(n1828) );
  XOR U2833 ( .A(n1760), .B(n1829), .Z(n1755) );
  XOR U2834 ( .A(n1759), .B(n1762), .Z(n1829) );
  IV U2835 ( .A(n1761), .Z(n1762) );
  NAND U2836 ( .A(n1830), .B(n1831), .Z(n1761) );
  OR U2837 ( .A(n1832), .B(n1833), .Z(n1831) );
  OR U2838 ( .A(n1834), .B(n1835), .Z(n1830) );
  NAND U2839 ( .A(n1836), .B(n1837), .Z(n1759) );
  OR U2840 ( .A(n1838), .B(n1839), .Z(n1837) );
  OR U2841 ( .A(n1840), .B(n1841), .Z(n1836) );
  NOR U2842 ( .A(n1842), .B(n1843), .Z(n1760) );
  ANDN U2843 ( .B(n1844), .A(n1845), .Z(n1754) );
  IV U2844 ( .A(n1846), .Z(n1844) );
  XNOR U2845 ( .A(n1747), .B(n1847), .Z(n1753) );
  XNOR U2846 ( .A(n1746), .B(n1748), .Z(n1847) );
  NAND U2847 ( .A(n1848), .B(n1849), .Z(n1748) );
  OR U2848 ( .A(n1850), .B(n1851), .Z(n1849) );
  OR U2849 ( .A(n1852), .B(n1853), .Z(n1848) );
  NAND U2850 ( .A(n1854), .B(n1855), .Z(n1746) );
  OR U2851 ( .A(n1856), .B(n1857), .Z(n1855) );
  OR U2852 ( .A(n1858), .B(n1859), .Z(n1854) );
  ANDN U2853 ( .B(n1860), .A(n1861), .Z(n1747) );
  IV U2854 ( .A(n1862), .Z(n1860) );
  XNOR U2855 ( .A(n1827), .B(n1826), .Z(N6124) );
  XOR U2856 ( .A(n1846), .B(n1845), .Z(n1826) );
  XNOR U2857 ( .A(n1861), .B(n1862), .Z(n1845) );
  XNOR U2858 ( .A(n1856), .B(n1857), .Z(n1862) );
  XNOR U2859 ( .A(n1858), .B(n1859), .Z(n1857) );
  XNOR U2860 ( .A(y[820]), .B(x[820]), .Z(n1859) );
  XNOR U2861 ( .A(y[821]), .B(x[821]), .Z(n1858) );
  XNOR U2862 ( .A(y[819]), .B(x[819]), .Z(n1856) );
  XNOR U2863 ( .A(n1850), .B(n1851), .Z(n1861) );
  XNOR U2864 ( .A(y[816]), .B(x[816]), .Z(n1851) );
  XNOR U2865 ( .A(n1852), .B(n1853), .Z(n1850) );
  XNOR U2866 ( .A(y[817]), .B(x[817]), .Z(n1853) );
  XNOR U2867 ( .A(y[818]), .B(x[818]), .Z(n1852) );
  XNOR U2868 ( .A(n1843), .B(n1842), .Z(n1846) );
  XNOR U2869 ( .A(n1838), .B(n1839), .Z(n1842) );
  XNOR U2870 ( .A(y[813]), .B(x[813]), .Z(n1839) );
  XNOR U2871 ( .A(n1840), .B(n1841), .Z(n1838) );
  XNOR U2872 ( .A(y[814]), .B(x[814]), .Z(n1841) );
  XNOR U2873 ( .A(y[815]), .B(x[815]), .Z(n1840) );
  XNOR U2874 ( .A(n1832), .B(n1833), .Z(n1843) );
  XNOR U2875 ( .A(y[810]), .B(x[810]), .Z(n1833) );
  XNOR U2876 ( .A(n1834), .B(n1835), .Z(n1832) );
  XNOR U2877 ( .A(y[811]), .B(x[811]), .Z(n1835) );
  XNOR U2878 ( .A(y[812]), .B(x[812]), .Z(n1834) );
  XOR U2879 ( .A(n1808), .B(n1809), .Z(n1827) );
  XNOR U2880 ( .A(n1824), .B(n1825), .Z(n1809) );
  XNOR U2881 ( .A(n1819), .B(n1820), .Z(n1825) );
  XNOR U2882 ( .A(n1821), .B(n1822), .Z(n1820) );
  XNOR U2883 ( .A(y[808]), .B(x[808]), .Z(n1822) );
  XNOR U2884 ( .A(y[809]), .B(x[809]), .Z(n1821) );
  XNOR U2885 ( .A(y[807]), .B(x[807]), .Z(n1819) );
  XNOR U2886 ( .A(n1813), .B(n1814), .Z(n1824) );
  XNOR U2887 ( .A(y[804]), .B(x[804]), .Z(n1814) );
  XNOR U2888 ( .A(n1815), .B(n1816), .Z(n1813) );
  XNOR U2889 ( .A(y[805]), .B(x[805]), .Z(n1816) );
  XNOR U2890 ( .A(y[806]), .B(x[806]), .Z(n1815) );
  XOR U2891 ( .A(n1807), .B(n1806), .Z(n1808) );
  XNOR U2892 ( .A(n1802), .B(n1803), .Z(n1806) );
  XNOR U2893 ( .A(y[801]), .B(x[801]), .Z(n1803) );
  XNOR U2894 ( .A(n1804), .B(n1805), .Z(n1802) );
  XNOR U2895 ( .A(y[802]), .B(x[802]), .Z(n1805) );
  XNOR U2896 ( .A(y[803]), .B(x[803]), .Z(n1804) );
  XNOR U2897 ( .A(n1796), .B(n1797), .Z(n1807) );
  XNOR U2898 ( .A(y[798]), .B(x[798]), .Z(n1797) );
  XNOR U2899 ( .A(n1798), .B(n1799), .Z(n1796) );
  XNOR U2900 ( .A(y[799]), .B(x[799]), .Z(n1799) );
  XNOR U2901 ( .A(y[800]), .B(x[800]), .Z(n1798) );
  NAND U2902 ( .A(n1863), .B(n1864), .Z(N6118) );
  NANDN U2903 ( .A(n1865), .B(n1866), .Z(n1864) );
  OR U2904 ( .A(n1867), .B(n1868), .Z(n1866) );
  NAND U2905 ( .A(n1867), .B(n1868), .Z(n1863) );
  XOR U2906 ( .A(n1867), .B(n1869), .Z(N6117) );
  XNOR U2907 ( .A(n1865), .B(n1868), .Z(n1869) );
  AND U2908 ( .A(n1870), .B(n1871), .Z(n1868) );
  NANDN U2909 ( .A(n1872), .B(n1873), .Z(n1871) );
  NANDN U2910 ( .A(n1874), .B(n1875), .Z(n1873) );
  NANDN U2911 ( .A(n1875), .B(n1874), .Z(n1870) );
  NAND U2912 ( .A(n1876), .B(n1877), .Z(n1865) );
  NANDN U2913 ( .A(n1878), .B(n1879), .Z(n1877) );
  OR U2914 ( .A(n1880), .B(n1881), .Z(n1879) );
  NAND U2915 ( .A(n1881), .B(n1880), .Z(n1876) );
  AND U2916 ( .A(n1882), .B(n1883), .Z(n1867) );
  NANDN U2917 ( .A(n1884), .B(n1885), .Z(n1883) );
  NANDN U2918 ( .A(n1886), .B(n1887), .Z(n1885) );
  NANDN U2919 ( .A(n1887), .B(n1886), .Z(n1882) );
  XOR U2920 ( .A(n1881), .B(n1888), .Z(N6116) );
  XOR U2921 ( .A(n1878), .B(n1880), .Z(n1888) );
  XNOR U2922 ( .A(n1874), .B(n1889), .Z(n1880) );
  XNOR U2923 ( .A(n1872), .B(n1875), .Z(n1889) );
  NAND U2924 ( .A(n1890), .B(n1891), .Z(n1875) );
  NAND U2925 ( .A(n1892), .B(n1893), .Z(n1891) );
  OR U2926 ( .A(n1894), .B(n1895), .Z(n1892) );
  NANDN U2927 ( .A(n1896), .B(n1894), .Z(n1890) );
  IV U2928 ( .A(n1895), .Z(n1896) );
  NAND U2929 ( .A(n1897), .B(n1898), .Z(n1872) );
  NAND U2930 ( .A(n1899), .B(n1900), .Z(n1898) );
  NANDN U2931 ( .A(n1901), .B(n1902), .Z(n1899) );
  NANDN U2932 ( .A(n1902), .B(n1901), .Z(n1897) );
  AND U2933 ( .A(n1903), .B(n1904), .Z(n1874) );
  NAND U2934 ( .A(n1905), .B(n1906), .Z(n1904) );
  OR U2935 ( .A(n1907), .B(n1908), .Z(n1905) );
  NANDN U2936 ( .A(n1909), .B(n1907), .Z(n1903) );
  NAND U2937 ( .A(n1910), .B(n1911), .Z(n1878) );
  NANDN U2938 ( .A(n1912), .B(n1913), .Z(n1911) );
  OR U2939 ( .A(n1914), .B(n1915), .Z(n1913) );
  NANDN U2940 ( .A(n1916), .B(n1914), .Z(n1910) );
  IV U2941 ( .A(n1915), .Z(n1916) );
  XNOR U2942 ( .A(n1886), .B(n1917), .Z(n1881) );
  XNOR U2943 ( .A(n1884), .B(n1887), .Z(n1917) );
  NAND U2944 ( .A(n1918), .B(n1919), .Z(n1887) );
  NAND U2945 ( .A(n1920), .B(n1921), .Z(n1919) );
  OR U2946 ( .A(n1922), .B(n1923), .Z(n1920) );
  NANDN U2947 ( .A(n1924), .B(n1922), .Z(n1918) );
  IV U2948 ( .A(n1923), .Z(n1924) );
  NAND U2949 ( .A(n1925), .B(n1926), .Z(n1884) );
  NAND U2950 ( .A(n1927), .B(n1928), .Z(n1926) );
  NANDN U2951 ( .A(n1929), .B(n1930), .Z(n1927) );
  NANDN U2952 ( .A(n1930), .B(n1929), .Z(n1925) );
  AND U2953 ( .A(n1931), .B(n1932), .Z(n1886) );
  NAND U2954 ( .A(n1933), .B(n1934), .Z(n1932) );
  OR U2955 ( .A(n1935), .B(n1936), .Z(n1933) );
  NANDN U2956 ( .A(n1937), .B(n1935), .Z(n1931) );
  XNOR U2957 ( .A(n1912), .B(n1938), .Z(N6115) );
  XOR U2958 ( .A(n1914), .B(n1915), .Z(n1938) );
  XNOR U2959 ( .A(n1928), .B(n1939), .Z(n1915) );
  XOR U2960 ( .A(n1929), .B(n1930), .Z(n1939) );
  XOR U2961 ( .A(n1935), .B(n1940), .Z(n1930) );
  XOR U2962 ( .A(n1934), .B(n1937), .Z(n1940) );
  IV U2963 ( .A(n1936), .Z(n1937) );
  NAND U2964 ( .A(n1941), .B(n1942), .Z(n1936) );
  OR U2965 ( .A(n1943), .B(n1944), .Z(n1942) );
  OR U2966 ( .A(n1945), .B(n1946), .Z(n1941) );
  NAND U2967 ( .A(n1947), .B(n1948), .Z(n1934) );
  OR U2968 ( .A(n1949), .B(n1950), .Z(n1948) );
  OR U2969 ( .A(n1951), .B(n1952), .Z(n1947) );
  NOR U2970 ( .A(n1953), .B(n1954), .Z(n1935) );
  ANDN U2971 ( .B(n1955), .A(n1956), .Z(n1929) );
  XNOR U2972 ( .A(n1922), .B(n1957), .Z(n1928) );
  XNOR U2973 ( .A(n1921), .B(n1923), .Z(n1957) );
  NAND U2974 ( .A(n1958), .B(n1959), .Z(n1923) );
  OR U2975 ( .A(n1960), .B(n1961), .Z(n1959) );
  OR U2976 ( .A(n1962), .B(n1963), .Z(n1958) );
  NAND U2977 ( .A(n1964), .B(n1965), .Z(n1921) );
  OR U2978 ( .A(n1966), .B(n1967), .Z(n1965) );
  OR U2979 ( .A(n1968), .B(n1969), .Z(n1964) );
  ANDN U2980 ( .B(n1970), .A(n1971), .Z(n1922) );
  IV U2981 ( .A(n1972), .Z(n1970) );
  ANDN U2982 ( .B(n1973), .A(n1974), .Z(n1914) );
  XOR U2983 ( .A(n1900), .B(n1975), .Z(n1912) );
  XOR U2984 ( .A(n1901), .B(n1902), .Z(n1975) );
  XOR U2985 ( .A(n1907), .B(n1976), .Z(n1902) );
  XOR U2986 ( .A(n1906), .B(n1909), .Z(n1976) );
  IV U2987 ( .A(n1908), .Z(n1909) );
  NAND U2988 ( .A(n1977), .B(n1978), .Z(n1908) );
  OR U2989 ( .A(n1979), .B(n1980), .Z(n1978) );
  OR U2990 ( .A(n1981), .B(n1982), .Z(n1977) );
  NAND U2991 ( .A(n1983), .B(n1984), .Z(n1906) );
  OR U2992 ( .A(n1985), .B(n1986), .Z(n1984) );
  OR U2993 ( .A(n1987), .B(n1988), .Z(n1983) );
  NOR U2994 ( .A(n1989), .B(n1990), .Z(n1907) );
  ANDN U2995 ( .B(n1991), .A(n1992), .Z(n1901) );
  IV U2996 ( .A(n1993), .Z(n1991) );
  XNOR U2997 ( .A(n1894), .B(n1994), .Z(n1900) );
  XNOR U2998 ( .A(n1893), .B(n1895), .Z(n1994) );
  NAND U2999 ( .A(n1995), .B(n1996), .Z(n1895) );
  OR U3000 ( .A(n1997), .B(n1998), .Z(n1996) );
  OR U3001 ( .A(n1999), .B(n2000), .Z(n1995) );
  NAND U3002 ( .A(n2001), .B(n2002), .Z(n1893) );
  OR U3003 ( .A(n2003), .B(n2004), .Z(n2002) );
  OR U3004 ( .A(n2005), .B(n2006), .Z(n2001) );
  ANDN U3005 ( .B(n2007), .A(n2008), .Z(n1894) );
  IV U3006 ( .A(n2009), .Z(n2007) );
  XNOR U3007 ( .A(n1974), .B(n1973), .Z(N6114) );
  XOR U3008 ( .A(n1993), .B(n1992), .Z(n1973) );
  XNOR U3009 ( .A(n2008), .B(n2009), .Z(n1992) );
  XNOR U3010 ( .A(n2003), .B(n2004), .Z(n2009) );
  XNOR U3011 ( .A(n2005), .B(n2006), .Z(n2004) );
  XNOR U3012 ( .A(y[796]), .B(x[796]), .Z(n2006) );
  XNOR U3013 ( .A(y[797]), .B(x[797]), .Z(n2005) );
  XNOR U3014 ( .A(y[795]), .B(x[795]), .Z(n2003) );
  XNOR U3015 ( .A(n1997), .B(n1998), .Z(n2008) );
  XNOR U3016 ( .A(y[792]), .B(x[792]), .Z(n1998) );
  XNOR U3017 ( .A(n1999), .B(n2000), .Z(n1997) );
  XNOR U3018 ( .A(y[793]), .B(x[793]), .Z(n2000) );
  XNOR U3019 ( .A(y[794]), .B(x[794]), .Z(n1999) );
  XNOR U3020 ( .A(n1990), .B(n1989), .Z(n1993) );
  XNOR U3021 ( .A(n1985), .B(n1986), .Z(n1989) );
  XNOR U3022 ( .A(y[789]), .B(x[789]), .Z(n1986) );
  XNOR U3023 ( .A(n1987), .B(n1988), .Z(n1985) );
  XNOR U3024 ( .A(y[790]), .B(x[790]), .Z(n1988) );
  XNOR U3025 ( .A(y[791]), .B(x[791]), .Z(n1987) );
  XNOR U3026 ( .A(n1979), .B(n1980), .Z(n1990) );
  XNOR U3027 ( .A(y[786]), .B(x[786]), .Z(n1980) );
  XNOR U3028 ( .A(n1981), .B(n1982), .Z(n1979) );
  XNOR U3029 ( .A(y[787]), .B(x[787]), .Z(n1982) );
  XNOR U3030 ( .A(y[788]), .B(x[788]), .Z(n1981) );
  XOR U3031 ( .A(n1955), .B(n1956), .Z(n1974) );
  XNOR U3032 ( .A(n1971), .B(n1972), .Z(n1956) );
  XNOR U3033 ( .A(n1966), .B(n1967), .Z(n1972) );
  XNOR U3034 ( .A(n1968), .B(n1969), .Z(n1967) );
  XNOR U3035 ( .A(y[784]), .B(x[784]), .Z(n1969) );
  XNOR U3036 ( .A(y[785]), .B(x[785]), .Z(n1968) );
  XNOR U3037 ( .A(y[783]), .B(x[783]), .Z(n1966) );
  XNOR U3038 ( .A(n1960), .B(n1961), .Z(n1971) );
  XNOR U3039 ( .A(y[780]), .B(x[780]), .Z(n1961) );
  XNOR U3040 ( .A(n1962), .B(n1963), .Z(n1960) );
  XNOR U3041 ( .A(y[781]), .B(x[781]), .Z(n1963) );
  XNOR U3042 ( .A(y[782]), .B(x[782]), .Z(n1962) );
  XOR U3043 ( .A(n1954), .B(n1953), .Z(n1955) );
  XNOR U3044 ( .A(n1949), .B(n1950), .Z(n1953) );
  XNOR U3045 ( .A(y[777]), .B(x[777]), .Z(n1950) );
  XNOR U3046 ( .A(n1951), .B(n1952), .Z(n1949) );
  XNOR U3047 ( .A(y[778]), .B(x[778]), .Z(n1952) );
  XNOR U3048 ( .A(y[779]), .B(x[779]), .Z(n1951) );
  XNOR U3049 ( .A(n1943), .B(n1944), .Z(n1954) );
  XNOR U3050 ( .A(y[774]), .B(x[774]), .Z(n1944) );
  XNOR U3051 ( .A(n1945), .B(n1946), .Z(n1943) );
  XNOR U3052 ( .A(y[775]), .B(x[775]), .Z(n1946) );
  XNOR U3053 ( .A(y[776]), .B(x[776]), .Z(n1945) );
  NAND U3054 ( .A(n2010), .B(n2011), .Z(N6108) );
  NANDN U3055 ( .A(n2012), .B(n2013), .Z(n2011) );
  OR U3056 ( .A(n2014), .B(n2015), .Z(n2013) );
  NAND U3057 ( .A(n2014), .B(n2015), .Z(n2010) );
  XOR U3058 ( .A(n2014), .B(n2016), .Z(N6107) );
  XNOR U3059 ( .A(n2012), .B(n2015), .Z(n2016) );
  AND U3060 ( .A(n2017), .B(n2018), .Z(n2015) );
  NANDN U3061 ( .A(n2019), .B(n2020), .Z(n2018) );
  NANDN U3062 ( .A(n2021), .B(n2022), .Z(n2020) );
  NANDN U3063 ( .A(n2022), .B(n2021), .Z(n2017) );
  NAND U3064 ( .A(n2023), .B(n2024), .Z(n2012) );
  NANDN U3065 ( .A(n2025), .B(n2026), .Z(n2024) );
  OR U3066 ( .A(n2027), .B(n2028), .Z(n2026) );
  NAND U3067 ( .A(n2028), .B(n2027), .Z(n2023) );
  AND U3068 ( .A(n2029), .B(n2030), .Z(n2014) );
  NANDN U3069 ( .A(n2031), .B(n2032), .Z(n2030) );
  NANDN U3070 ( .A(n2033), .B(n2034), .Z(n2032) );
  NANDN U3071 ( .A(n2034), .B(n2033), .Z(n2029) );
  XOR U3072 ( .A(n2028), .B(n2035), .Z(N6106) );
  XOR U3073 ( .A(n2025), .B(n2027), .Z(n2035) );
  XNOR U3074 ( .A(n2021), .B(n2036), .Z(n2027) );
  XNOR U3075 ( .A(n2019), .B(n2022), .Z(n2036) );
  NAND U3076 ( .A(n2037), .B(n2038), .Z(n2022) );
  NAND U3077 ( .A(n2039), .B(n2040), .Z(n2038) );
  OR U3078 ( .A(n2041), .B(n2042), .Z(n2039) );
  NANDN U3079 ( .A(n2043), .B(n2041), .Z(n2037) );
  IV U3080 ( .A(n2042), .Z(n2043) );
  NAND U3081 ( .A(n2044), .B(n2045), .Z(n2019) );
  NAND U3082 ( .A(n2046), .B(n2047), .Z(n2045) );
  NANDN U3083 ( .A(n2048), .B(n2049), .Z(n2046) );
  NANDN U3084 ( .A(n2049), .B(n2048), .Z(n2044) );
  AND U3085 ( .A(n2050), .B(n2051), .Z(n2021) );
  NAND U3086 ( .A(n2052), .B(n2053), .Z(n2051) );
  OR U3087 ( .A(n2054), .B(n2055), .Z(n2052) );
  NANDN U3088 ( .A(n2056), .B(n2054), .Z(n2050) );
  NAND U3089 ( .A(n2057), .B(n2058), .Z(n2025) );
  NANDN U3090 ( .A(n2059), .B(n2060), .Z(n2058) );
  OR U3091 ( .A(n2061), .B(n2062), .Z(n2060) );
  NANDN U3092 ( .A(n2063), .B(n2061), .Z(n2057) );
  IV U3093 ( .A(n2062), .Z(n2063) );
  XNOR U3094 ( .A(n2033), .B(n2064), .Z(n2028) );
  XNOR U3095 ( .A(n2031), .B(n2034), .Z(n2064) );
  NAND U3096 ( .A(n2065), .B(n2066), .Z(n2034) );
  NAND U3097 ( .A(n2067), .B(n2068), .Z(n2066) );
  OR U3098 ( .A(n2069), .B(n2070), .Z(n2067) );
  NANDN U3099 ( .A(n2071), .B(n2069), .Z(n2065) );
  IV U3100 ( .A(n2070), .Z(n2071) );
  NAND U3101 ( .A(n2072), .B(n2073), .Z(n2031) );
  NAND U3102 ( .A(n2074), .B(n2075), .Z(n2073) );
  NANDN U3103 ( .A(n2076), .B(n2077), .Z(n2074) );
  NANDN U3104 ( .A(n2077), .B(n2076), .Z(n2072) );
  AND U3105 ( .A(n2078), .B(n2079), .Z(n2033) );
  NAND U3106 ( .A(n2080), .B(n2081), .Z(n2079) );
  OR U3107 ( .A(n2082), .B(n2083), .Z(n2080) );
  NANDN U3108 ( .A(n2084), .B(n2082), .Z(n2078) );
  XNOR U3109 ( .A(n2059), .B(n2085), .Z(N6105) );
  XOR U3110 ( .A(n2061), .B(n2062), .Z(n2085) );
  XNOR U3111 ( .A(n2075), .B(n2086), .Z(n2062) );
  XOR U3112 ( .A(n2076), .B(n2077), .Z(n2086) );
  XOR U3113 ( .A(n2082), .B(n2087), .Z(n2077) );
  XOR U3114 ( .A(n2081), .B(n2084), .Z(n2087) );
  IV U3115 ( .A(n2083), .Z(n2084) );
  NAND U3116 ( .A(n2088), .B(n2089), .Z(n2083) );
  OR U3117 ( .A(n2090), .B(n2091), .Z(n2089) );
  OR U3118 ( .A(n2092), .B(n2093), .Z(n2088) );
  NAND U3119 ( .A(n2094), .B(n2095), .Z(n2081) );
  OR U3120 ( .A(n2096), .B(n2097), .Z(n2095) );
  OR U3121 ( .A(n2098), .B(n2099), .Z(n2094) );
  NOR U3122 ( .A(n2100), .B(n2101), .Z(n2082) );
  ANDN U3123 ( .B(n2102), .A(n2103), .Z(n2076) );
  XNOR U3124 ( .A(n2069), .B(n2104), .Z(n2075) );
  XNOR U3125 ( .A(n2068), .B(n2070), .Z(n2104) );
  NAND U3126 ( .A(n2105), .B(n2106), .Z(n2070) );
  OR U3127 ( .A(n2107), .B(n2108), .Z(n2106) );
  OR U3128 ( .A(n2109), .B(n2110), .Z(n2105) );
  NAND U3129 ( .A(n2111), .B(n2112), .Z(n2068) );
  OR U3130 ( .A(n2113), .B(n2114), .Z(n2112) );
  OR U3131 ( .A(n2115), .B(n2116), .Z(n2111) );
  ANDN U3132 ( .B(n2117), .A(n2118), .Z(n2069) );
  IV U3133 ( .A(n2119), .Z(n2117) );
  ANDN U3134 ( .B(n2120), .A(n2121), .Z(n2061) );
  XOR U3135 ( .A(n2047), .B(n2122), .Z(n2059) );
  XOR U3136 ( .A(n2048), .B(n2049), .Z(n2122) );
  XOR U3137 ( .A(n2054), .B(n2123), .Z(n2049) );
  XOR U3138 ( .A(n2053), .B(n2056), .Z(n2123) );
  IV U3139 ( .A(n2055), .Z(n2056) );
  NAND U3140 ( .A(n2124), .B(n2125), .Z(n2055) );
  OR U3141 ( .A(n2126), .B(n2127), .Z(n2125) );
  OR U3142 ( .A(n2128), .B(n2129), .Z(n2124) );
  NAND U3143 ( .A(n2130), .B(n2131), .Z(n2053) );
  OR U3144 ( .A(n2132), .B(n2133), .Z(n2131) );
  OR U3145 ( .A(n2134), .B(n2135), .Z(n2130) );
  NOR U3146 ( .A(n2136), .B(n2137), .Z(n2054) );
  ANDN U3147 ( .B(n2138), .A(n2139), .Z(n2048) );
  IV U3148 ( .A(n2140), .Z(n2138) );
  XNOR U3149 ( .A(n2041), .B(n2141), .Z(n2047) );
  XNOR U3150 ( .A(n2040), .B(n2042), .Z(n2141) );
  NAND U3151 ( .A(n2142), .B(n2143), .Z(n2042) );
  OR U3152 ( .A(n2144), .B(n2145), .Z(n2143) );
  OR U3153 ( .A(n2146), .B(n2147), .Z(n2142) );
  NAND U3154 ( .A(n2148), .B(n2149), .Z(n2040) );
  OR U3155 ( .A(n2150), .B(n2151), .Z(n2149) );
  OR U3156 ( .A(n2152), .B(n2153), .Z(n2148) );
  ANDN U3157 ( .B(n2154), .A(n2155), .Z(n2041) );
  IV U3158 ( .A(n2156), .Z(n2154) );
  XNOR U3159 ( .A(n2121), .B(n2120), .Z(N6104) );
  XOR U3160 ( .A(n2140), .B(n2139), .Z(n2120) );
  XNOR U3161 ( .A(n2155), .B(n2156), .Z(n2139) );
  XNOR U3162 ( .A(n2150), .B(n2151), .Z(n2156) );
  XNOR U3163 ( .A(n2152), .B(n2153), .Z(n2151) );
  XNOR U3164 ( .A(y[772]), .B(x[772]), .Z(n2153) );
  XNOR U3165 ( .A(y[773]), .B(x[773]), .Z(n2152) );
  XNOR U3166 ( .A(y[771]), .B(x[771]), .Z(n2150) );
  XNOR U3167 ( .A(n2144), .B(n2145), .Z(n2155) );
  XNOR U3168 ( .A(y[768]), .B(x[768]), .Z(n2145) );
  XNOR U3169 ( .A(n2146), .B(n2147), .Z(n2144) );
  XNOR U3170 ( .A(y[769]), .B(x[769]), .Z(n2147) );
  XNOR U3171 ( .A(y[770]), .B(x[770]), .Z(n2146) );
  XNOR U3172 ( .A(n2137), .B(n2136), .Z(n2140) );
  XNOR U3173 ( .A(n2132), .B(n2133), .Z(n2136) );
  XNOR U3174 ( .A(y[765]), .B(x[765]), .Z(n2133) );
  XNOR U3175 ( .A(n2134), .B(n2135), .Z(n2132) );
  XNOR U3176 ( .A(y[766]), .B(x[766]), .Z(n2135) );
  XNOR U3177 ( .A(y[767]), .B(x[767]), .Z(n2134) );
  XNOR U3178 ( .A(n2126), .B(n2127), .Z(n2137) );
  XNOR U3179 ( .A(y[762]), .B(x[762]), .Z(n2127) );
  XNOR U3180 ( .A(n2128), .B(n2129), .Z(n2126) );
  XNOR U3181 ( .A(y[763]), .B(x[763]), .Z(n2129) );
  XNOR U3182 ( .A(y[764]), .B(x[764]), .Z(n2128) );
  XOR U3183 ( .A(n2102), .B(n2103), .Z(n2121) );
  XNOR U3184 ( .A(n2118), .B(n2119), .Z(n2103) );
  XNOR U3185 ( .A(n2113), .B(n2114), .Z(n2119) );
  XNOR U3186 ( .A(n2115), .B(n2116), .Z(n2114) );
  XNOR U3187 ( .A(y[760]), .B(x[760]), .Z(n2116) );
  XNOR U3188 ( .A(y[761]), .B(x[761]), .Z(n2115) );
  XNOR U3189 ( .A(y[759]), .B(x[759]), .Z(n2113) );
  XNOR U3190 ( .A(n2107), .B(n2108), .Z(n2118) );
  XNOR U3191 ( .A(y[756]), .B(x[756]), .Z(n2108) );
  XNOR U3192 ( .A(n2109), .B(n2110), .Z(n2107) );
  XNOR U3193 ( .A(y[757]), .B(x[757]), .Z(n2110) );
  XNOR U3194 ( .A(y[758]), .B(x[758]), .Z(n2109) );
  XOR U3195 ( .A(n2101), .B(n2100), .Z(n2102) );
  XNOR U3196 ( .A(n2096), .B(n2097), .Z(n2100) );
  XNOR U3197 ( .A(y[753]), .B(x[753]), .Z(n2097) );
  XNOR U3198 ( .A(n2098), .B(n2099), .Z(n2096) );
  XNOR U3199 ( .A(y[754]), .B(x[754]), .Z(n2099) );
  XNOR U3200 ( .A(y[755]), .B(x[755]), .Z(n2098) );
  XNOR U3201 ( .A(n2090), .B(n2091), .Z(n2101) );
  XNOR U3202 ( .A(y[750]), .B(x[750]), .Z(n2091) );
  XNOR U3203 ( .A(n2092), .B(n2093), .Z(n2090) );
  XNOR U3204 ( .A(y[751]), .B(x[751]), .Z(n2093) );
  XNOR U3205 ( .A(y[752]), .B(x[752]), .Z(n2092) );
  NAND U3206 ( .A(n2157), .B(n2158), .Z(N6098) );
  NANDN U3207 ( .A(n2159), .B(n2160), .Z(n2158) );
  OR U3208 ( .A(n2161), .B(n2162), .Z(n2160) );
  NAND U3209 ( .A(n2161), .B(n2162), .Z(n2157) );
  XOR U3210 ( .A(n2161), .B(n2163), .Z(N6097) );
  XNOR U3211 ( .A(n2159), .B(n2162), .Z(n2163) );
  AND U3212 ( .A(n2164), .B(n2165), .Z(n2162) );
  NANDN U3213 ( .A(n2166), .B(n2167), .Z(n2165) );
  NANDN U3214 ( .A(n2168), .B(n2169), .Z(n2167) );
  NANDN U3215 ( .A(n2169), .B(n2168), .Z(n2164) );
  NAND U3216 ( .A(n2170), .B(n2171), .Z(n2159) );
  NANDN U3217 ( .A(n2172), .B(n2173), .Z(n2171) );
  OR U3218 ( .A(n2174), .B(n2175), .Z(n2173) );
  NAND U3219 ( .A(n2175), .B(n2174), .Z(n2170) );
  AND U3220 ( .A(n2176), .B(n2177), .Z(n2161) );
  NANDN U3221 ( .A(n2178), .B(n2179), .Z(n2177) );
  NANDN U3222 ( .A(n2180), .B(n2181), .Z(n2179) );
  NANDN U3223 ( .A(n2181), .B(n2180), .Z(n2176) );
  XOR U3224 ( .A(n2175), .B(n2182), .Z(N6096) );
  XOR U3225 ( .A(n2172), .B(n2174), .Z(n2182) );
  XNOR U3226 ( .A(n2168), .B(n2183), .Z(n2174) );
  XNOR U3227 ( .A(n2166), .B(n2169), .Z(n2183) );
  NAND U3228 ( .A(n2184), .B(n2185), .Z(n2169) );
  NAND U3229 ( .A(n2186), .B(n2187), .Z(n2185) );
  OR U3230 ( .A(n2188), .B(n2189), .Z(n2186) );
  NANDN U3231 ( .A(n2190), .B(n2188), .Z(n2184) );
  IV U3232 ( .A(n2189), .Z(n2190) );
  NAND U3233 ( .A(n2191), .B(n2192), .Z(n2166) );
  NAND U3234 ( .A(n2193), .B(n2194), .Z(n2192) );
  NANDN U3235 ( .A(n2195), .B(n2196), .Z(n2193) );
  NANDN U3236 ( .A(n2196), .B(n2195), .Z(n2191) );
  AND U3237 ( .A(n2197), .B(n2198), .Z(n2168) );
  NAND U3238 ( .A(n2199), .B(n2200), .Z(n2198) );
  OR U3239 ( .A(n2201), .B(n2202), .Z(n2199) );
  NANDN U3240 ( .A(n2203), .B(n2201), .Z(n2197) );
  NAND U3241 ( .A(n2204), .B(n2205), .Z(n2172) );
  NANDN U3242 ( .A(n2206), .B(n2207), .Z(n2205) );
  OR U3243 ( .A(n2208), .B(n2209), .Z(n2207) );
  NANDN U3244 ( .A(n2210), .B(n2208), .Z(n2204) );
  IV U3245 ( .A(n2209), .Z(n2210) );
  XNOR U3246 ( .A(n2180), .B(n2211), .Z(n2175) );
  XNOR U3247 ( .A(n2178), .B(n2181), .Z(n2211) );
  NAND U3248 ( .A(n2212), .B(n2213), .Z(n2181) );
  NAND U3249 ( .A(n2214), .B(n2215), .Z(n2213) );
  OR U3250 ( .A(n2216), .B(n2217), .Z(n2214) );
  NANDN U3251 ( .A(n2218), .B(n2216), .Z(n2212) );
  IV U3252 ( .A(n2217), .Z(n2218) );
  NAND U3253 ( .A(n2219), .B(n2220), .Z(n2178) );
  NAND U3254 ( .A(n2221), .B(n2222), .Z(n2220) );
  NANDN U3255 ( .A(n2223), .B(n2224), .Z(n2221) );
  NANDN U3256 ( .A(n2224), .B(n2223), .Z(n2219) );
  AND U3257 ( .A(n2225), .B(n2226), .Z(n2180) );
  NAND U3258 ( .A(n2227), .B(n2228), .Z(n2226) );
  OR U3259 ( .A(n2229), .B(n2230), .Z(n2227) );
  NANDN U3260 ( .A(n2231), .B(n2229), .Z(n2225) );
  XNOR U3261 ( .A(n2206), .B(n2232), .Z(N6095) );
  XOR U3262 ( .A(n2208), .B(n2209), .Z(n2232) );
  XNOR U3263 ( .A(n2222), .B(n2233), .Z(n2209) );
  XOR U3264 ( .A(n2223), .B(n2224), .Z(n2233) );
  XOR U3265 ( .A(n2229), .B(n2234), .Z(n2224) );
  XOR U3266 ( .A(n2228), .B(n2231), .Z(n2234) );
  IV U3267 ( .A(n2230), .Z(n2231) );
  NAND U3268 ( .A(n2235), .B(n2236), .Z(n2230) );
  OR U3269 ( .A(n2237), .B(n2238), .Z(n2236) );
  OR U3270 ( .A(n2239), .B(n2240), .Z(n2235) );
  NAND U3271 ( .A(n2241), .B(n2242), .Z(n2228) );
  OR U3272 ( .A(n2243), .B(n2244), .Z(n2242) );
  OR U3273 ( .A(n2245), .B(n2246), .Z(n2241) );
  NOR U3274 ( .A(n2247), .B(n2248), .Z(n2229) );
  ANDN U3275 ( .B(n2249), .A(n2250), .Z(n2223) );
  XNOR U3276 ( .A(n2216), .B(n2251), .Z(n2222) );
  XNOR U3277 ( .A(n2215), .B(n2217), .Z(n2251) );
  NAND U3278 ( .A(n2252), .B(n2253), .Z(n2217) );
  OR U3279 ( .A(n2254), .B(n2255), .Z(n2253) );
  OR U3280 ( .A(n2256), .B(n2257), .Z(n2252) );
  NAND U3281 ( .A(n2258), .B(n2259), .Z(n2215) );
  OR U3282 ( .A(n2260), .B(n2261), .Z(n2259) );
  OR U3283 ( .A(n2262), .B(n2263), .Z(n2258) );
  ANDN U3284 ( .B(n2264), .A(n2265), .Z(n2216) );
  IV U3285 ( .A(n2266), .Z(n2264) );
  ANDN U3286 ( .B(n2267), .A(n2268), .Z(n2208) );
  XOR U3287 ( .A(n2194), .B(n2269), .Z(n2206) );
  XOR U3288 ( .A(n2195), .B(n2196), .Z(n2269) );
  XOR U3289 ( .A(n2201), .B(n2270), .Z(n2196) );
  XOR U3290 ( .A(n2200), .B(n2203), .Z(n2270) );
  IV U3291 ( .A(n2202), .Z(n2203) );
  NAND U3292 ( .A(n2271), .B(n2272), .Z(n2202) );
  OR U3293 ( .A(n2273), .B(n2274), .Z(n2272) );
  OR U3294 ( .A(n2275), .B(n2276), .Z(n2271) );
  NAND U3295 ( .A(n2277), .B(n2278), .Z(n2200) );
  OR U3296 ( .A(n2279), .B(n2280), .Z(n2278) );
  OR U3297 ( .A(n2281), .B(n2282), .Z(n2277) );
  NOR U3298 ( .A(n2283), .B(n2284), .Z(n2201) );
  ANDN U3299 ( .B(n2285), .A(n2286), .Z(n2195) );
  IV U3300 ( .A(n2287), .Z(n2285) );
  XNOR U3301 ( .A(n2188), .B(n2288), .Z(n2194) );
  XNOR U3302 ( .A(n2187), .B(n2189), .Z(n2288) );
  NAND U3303 ( .A(n2289), .B(n2290), .Z(n2189) );
  OR U3304 ( .A(n2291), .B(n2292), .Z(n2290) );
  OR U3305 ( .A(n2293), .B(n2294), .Z(n2289) );
  NAND U3306 ( .A(n2295), .B(n2296), .Z(n2187) );
  OR U3307 ( .A(n2297), .B(n2298), .Z(n2296) );
  OR U3308 ( .A(n2299), .B(n2300), .Z(n2295) );
  ANDN U3309 ( .B(n2301), .A(n2302), .Z(n2188) );
  IV U3310 ( .A(n2303), .Z(n2301) );
  XNOR U3311 ( .A(n2268), .B(n2267), .Z(N6094) );
  XOR U3312 ( .A(n2287), .B(n2286), .Z(n2267) );
  XNOR U3313 ( .A(n2302), .B(n2303), .Z(n2286) );
  XNOR U3314 ( .A(n2297), .B(n2298), .Z(n2303) );
  XNOR U3315 ( .A(n2299), .B(n2300), .Z(n2298) );
  XNOR U3316 ( .A(y[748]), .B(x[748]), .Z(n2300) );
  XNOR U3317 ( .A(y[749]), .B(x[749]), .Z(n2299) );
  XNOR U3318 ( .A(y[747]), .B(x[747]), .Z(n2297) );
  XNOR U3319 ( .A(n2291), .B(n2292), .Z(n2302) );
  XNOR U3320 ( .A(y[744]), .B(x[744]), .Z(n2292) );
  XNOR U3321 ( .A(n2293), .B(n2294), .Z(n2291) );
  XNOR U3322 ( .A(y[745]), .B(x[745]), .Z(n2294) );
  XNOR U3323 ( .A(y[746]), .B(x[746]), .Z(n2293) );
  XNOR U3324 ( .A(n2284), .B(n2283), .Z(n2287) );
  XNOR U3325 ( .A(n2279), .B(n2280), .Z(n2283) );
  XNOR U3326 ( .A(y[741]), .B(x[741]), .Z(n2280) );
  XNOR U3327 ( .A(n2281), .B(n2282), .Z(n2279) );
  XNOR U3328 ( .A(y[742]), .B(x[742]), .Z(n2282) );
  XNOR U3329 ( .A(y[743]), .B(x[743]), .Z(n2281) );
  XNOR U3330 ( .A(n2273), .B(n2274), .Z(n2284) );
  XNOR U3331 ( .A(y[738]), .B(x[738]), .Z(n2274) );
  XNOR U3332 ( .A(n2275), .B(n2276), .Z(n2273) );
  XNOR U3333 ( .A(y[739]), .B(x[739]), .Z(n2276) );
  XNOR U3334 ( .A(y[740]), .B(x[740]), .Z(n2275) );
  XOR U3335 ( .A(n2249), .B(n2250), .Z(n2268) );
  XNOR U3336 ( .A(n2265), .B(n2266), .Z(n2250) );
  XNOR U3337 ( .A(n2260), .B(n2261), .Z(n2266) );
  XNOR U3338 ( .A(n2262), .B(n2263), .Z(n2261) );
  XNOR U3339 ( .A(y[736]), .B(x[736]), .Z(n2263) );
  XNOR U3340 ( .A(y[737]), .B(x[737]), .Z(n2262) );
  XNOR U3341 ( .A(y[735]), .B(x[735]), .Z(n2260) );
  XNOR U3342 ( .A(n2254), .B(n2255), .Z(n2265) );
  XNOR U3343 ( .A(y[732]), .B(x[732]), .Z(n2255) );
  XNOR U3344 ( .A(n2256), .B(n2257), .Z(n2254) );
  XNOR U3345 ( .A(y[733]), .B(x[733]), .Z(n2257) );
  XNOR U3346 ( .A(y[734]), .B(x[734]), .Z(n2256) );
  XOR U3347 ( .A(n2248), .B(n2247), .Z(n2249) );
  XNOR U3348 ( .A(n2243), .B(n2244), .Z(n2247) );
  XNOR U3349 ( .A(y[729]), .B(x[729]), .Z(n2244) );
  XNOR U3350 ( .A(n2245), .B(n2246), .Z(n2243) );
  XNOR U3351 ( .A(y[730]), .B(x[730]), .Z(n2246) );
  XNOR U3352 ( .A(y[731]), .B(x[731]), .Z(n2245) );
  XNOR U3353 ( .A(n2237), .B(n2238), .Z(n2248) );
  XNOR U3354 ( .A(y[726]), .B(x[726]), .Z(n2238) );
  XNOR U3355 ( .A(n2239), .B(n2240), .Z(n2237) );
  XNOR U3356 ( .A(y[727]), .B(x[727]), .Z(n2240) );
  XNOR U3357 ( .A(y[728]), .B(x[728]), .Z(n2239) );
  NAND U3358 ( .A(n2304), .B(n2305), .Z(N6088) );
  NANDN U3359 ( .A(n2306), .B(n2307), .Z(n2305) );
  OR U3360 ( .A(n2308), .B(n2309), .Z(n2307) );
  NAND U3361 ( .A(n2308), .B(n2309), .Z(n2304) );
  XOR U3362 ( .A(n2308), .B(n2310), .Z(N6087) );
  XNOR U3363 ( .A(n2306), .B(n2309), .Z(n2310) );
  AND U3364 ( .A(n2311), .B(n2312), .Z(n2309) );
  NANDN U3365 ( .A(n2313), .B(n2314), .Z(n2312) );
  NANDN U3366 ( .A(n2315), .B(n2316), .Z(n2314) );
  NANDN U3367 ( .A(n2316), .B(n2315), .Z(n2311) );
  NAND U3368 ( .A(n2317), .B(n2318), .Z(n2306) );
  NANDN U3369 ( .A(n2319), .B(n2320), .Z(n2318) );
  OR U3370 ( .A(n2321), .B(n2322), .Z(n2320) );
  NAND U3371 ( .A(n2322), .B(n2321), .Z(n2317) );
  AND U3372 ( .A(n2323), .B(n2324), .Z(n2308) );
  NANDN U3373 ( .A(n2325), .B(n2326), .Z(n2324) );
  NANDN U3374 ( .A(n2327), .B(n2328), .Z(n2326) );
  NANDN U3375 ( .A(n2328), .B(n2327), .Z(n2323) );
  XOR U3376 ( .A(n2322), .B(n2329), .Z(N6086) );
  XOR U3377 ( .A(n2319), .B(n2321), .Z(n2329) );
  XNOR U3378 ( .A(n2315), .B(n2330), .Z(n2321) );
  XNOR U3379 ( .A(n2313), .B(n2316), .Z(n2330) );
  NAND U3380 ( .A(n2331), .B(n2332), .Z(n2316) );
  NAND U3381 ( .A(n2333), .B(n2334), .Z(n2332) );
  OR U3382 ( .A(n2335), .B(n2336), .Z(n2333) );
  NANDN U3383 ( .A(n2337), .B(n2335), .Z(n2331) );
  IV U3384 ( .A(n2336), .Z(n2337) );
  NAND U3385 ( .A(n2338), .B(n2339), .Z(n2313) );
  NAND U3386 ( .A(n2340), .B(n2341), .Z(n2339) );
  NANDN U3387 ( .A(n2342), .B(n2343), .Z(n2340) );
  NANDN U3388 ( .A(n2343), .B(n2342), .Z(n2338) );
  AND U3389 ( .A(n2344), .B(n2345), .Z(n2315) );
  NAND U3390 ( .A(n2346), .B(n2347), .Z(n2345) );
  OR U3391 ( .A(n2348), .B(n2349), .Z(n2346) );
  NANDN U3392 ( .A(n2350), .B(n2348), .Z(n2344) );
  NAND U3393 ( .A(n2351), .B(n2352), .Z(n2319) );
  NANDN U3394 ( .A(n2353), .B(n2354), .Z(n2352) );
  OR U3395 ( .A(n2355), .B(n2356), .Z(n2354) );
  NANDN U3396 ( .A(n2357), .B(n2355), .Z(n2351) );
  IV U3397 ( .A(n2356), .Z(n2357) );
  XNOR U3398 ( .A(n2327), .B(n2358), .Z(n2322) );
  XNOR U3399 ( .A(n2325), .B(n2328), .Z(n2358) );
  NAND U3400 ( .A(n2359), .B(n2360), .Z(n2328) );
  NAND U3401 ( .A(n2361), .B(n2362), .Z(n2360) );
  OR U3402 ( .A(n2363), .B(n2364), .Z(n2361) );
  NANDN U3403 ( .A(n2365), .B(n2363), .Z(n2359) );
  IV U3404 ( .A(n2364), .Z(n2365) );
  NAND U3405 ( .A(n2366), .B(n2367), .Z(n2325) );
  NAND U3406 ( .A(n2368), .B(n2369), .Z(n2367) );
  NANDN U3407 ( .A(n2370), .B(n2371), .Z(n2368) );
  NANDN U3408 ( .A(n2371), .B(n2370), .Z(n2366) );
  AND U3409 ( .A(n2372), .B(n2373), .Z(n2327) );
  NAND U3410 ( .A(n2374), .B(n2375), .Z(n2373) );
  OR U3411 ( .A(n2376), .B(n2377), .Z(n2374) );
  NANDN U3412 ( .A(n2378), .B(n2376), .Z(n2372) );
  XNOR U3413 ( .A(n2353), .B(n2379), .Z(N6085) );
  XOR U3414 ( .A(n2355), .B(n2356), .Z(n2379) );
  XNOR U3415 ( .A(n2369), .B(n2380), .Z(n2356) );
  XOR U3416 ( .A(n2370), .B(n2371), .Z(n2380) );
  XOR U3417 ( .A(n2376), .B(n2381), .Z(n2371) );
  XOR U3418 ( .A(n2375), .B(n2378), .Z(n2381) );
  IV U3419 ( .A(n2377), .Z(n2378) );
  NAND U3420 ( .A(n2382), .B(n2383), .Z(n2377) );
  OR U3421 ( .A(n2384), .B(n2385), .Z(n2383) );
  OR U3422 ( .A(n2386), .B(n2387), .Z(n2382) );
  NAND U3423 ( .A(n2388), .B(n2389), .Z(n2375) );
  OR U3424 ( .A(n2390), .B(n2391), .Z(n2389) );
  OR U3425 ( .A(n2392), .B(n2393), .Z(n2388) );
  NOR U3426 ( .A(n2394), .B(n2395), .Z(n2376) );
  ANDN U3427 ( .B(n2396), .A(n2397), .Z(n2370) );
  XNOR U3428 ( .A(n2363), .B(n2398), .Z(n2369) );
  XNOR U3429 ( .A(n2362), .B(n2364), .Z(n2398) );
  NAND U3430 ( .A(n2399), .B(n2400), .Z(n2364) );
  OR U3431 ( .A(n2401), .B(n2402), .Z(n2400) );
  OR U3432 ( .A(n2403), .B(n2404), .Z(n2399) );
  NAND U3433 ( .A(n2405), .B(n2406), .Z(n2362) );
  OR U3434 ( .A(n2407), .B(n2408), .Z(n2406) );
  OR U3435 ( .A(n2409), .B(n2410), .Z(n2405) );
  ANDN U3436 ( .B(n2411), .A(n2412), .Z(n2363) );
  IV U3437 ( .A(n2413), .Z(n2411) );
  ANDN U3438 ( .B(n2414), .A(n2415), .Z(n2355) );
  XOR U3439 ( .A(n2341), .B(n2416), .Z(n2353) );
  XOR U3440 ( .A(n2342), .B(n2343), .Z(n2416) );
  XOR U3441 ( .A(n2348), .B(n2417), .Z(n2343) );
  XOR U3442 ( .A(n2347), .B(n2350), .Z(n2417) );
  IV U3443 ( .A(n2349), .Z(n2350) );
  NAND U3444 ( .A(n2418), .B(n2419), .Z(n2349) );
  OR U3445 ( .A(n2420), .B(n2421), .Z(n2419) );
  OR U3446 ( .A(n2422), .B(n2423), .Z(n2418) );
  NAND U3447 ( .A(n2424), .B(n2425), .Z(n2347) );
  OR U3448 ( .A(n2426), .B(n2427), .Z(n2425) );
  OR U3449 ( .A(n2428), .B(n2429), .Z(n2424) );
  NOR U3450 ( .A(n2430), .B(n2431), .Z(n2348) );
  ANDN U3451 ( .B(n2432), .A(n2433), .Z(n2342) );
  IV U3452 ( .A(n2434), .Z(n2432) );
  XNOR U3453 ( .A(n2335), .B(n2435), .Z(n2341) );
  XNOR U3454 ( .A(n2334), .B(n2336), .Z(n2435) );
  NAND U3455 ( .A(n2436), .B(n2437), .Z(n2336) );
  OR U3456 ( .A(n2438), .B(n2439), .Z(n2437) );
  OR U3457 ( .A(n2440), .B(n2441), .Z(n2436) );
  NAND U3458 ( .A(n2442), .B(n2443), .Z(n2334) );
  OR U3459 ( .A(n2444), .B(n2445), .Z(n2443) );
  OR U3460 ( .A(n2446), .B(n2447), .Z(n2442) );
  ANDN U3461 ( .B(n2448), .A(n2449), .Z(n2335) );
  IV U3462 ( .A(n2450), .Z(n2448) );
  XNOR U3463 ( .A(n2415), .B(n2414), .Z(N6084) );
  XOR U3464 ( .A(n2434), .B(n2433), .Z(n2414) );
  XNOR U3465 ( .A(n2449), .B(n2450), .Z(n2433) );
  XNOR U3466 ( .A(n2444), .B(n2445), .Z(n2450) );
  XNOR U3467 ( .A(n2446), .B(n2447), .Z(n2445) );
  XNOR U3468 ( .A(y[724]), .B(x[724]), .Z(n2447) );
  XNOR U3469 ( .A(y[725]), .B(x[725]), .Z(n2446) );
  XNOR U3470 ( .A(y[723]), .B(x[723]), .Z(n2444) );
  XNOR U3471 ( .A(n2438), .B(n2439), .Z(n2449) );
  XNOR U3472 ( .A(y[720]), .B(x[720]), .Z(n2439) );
  XNOR U3473 ( .A(n2440), .B(n2441), .Z(n2438) );
  XNOR U3474 ( .A(y[721]), .B(x[721]), .Z(n2441) );
  XNOR U3475 ( .A(y[722]), .B(x[722]), .Z(n2440) );
  XNOR U3476 ( .A(n2431), .B(n2430), .Z(n2434) );
  XNOR U3477 ( .A(n2426), .B(n2427), .Z(n2430) );
  XNOR U3478 ( .A(y[717]), .B(x[717]), .Z(n2427) );
  XNOR U3479 ( .A(n2428), .B(n2429), .Z(n2426) );
  XNOR U3480 ( .A(y[718]), .B(x[718]), .Z(n2429) );
  XNOR U3481 ( .A(y[719]), .B(x[719]), .Z(n2428) );
  XNOR U3482 ( .A(n2420), .B(n2421), .Z(n2431) );
  XNOR U3483 ( .A(y[714]), .B(x[714]), .Z(n2421) );
  XNOR U3484 ( .A(n2422), .B(n2423), .Z(n2420) );
  XNOR U3485 ( .A(y[715]), .B(x[715]), .Z(n2423) );
  XNOR U3486 ( .A(y[716]), .B(x[716]), .Z(n2422) );
  XOR U3487 ( .A(n2396), .B(n2397), .Z(n2415) );
  XNOR U3488 ( .A(n2412), .B(n2413), .Z(n2397) );
  XNOR U3489 ( .A(n2407), .B(n2408), .Z(n2413) );
  XNOR U3490 ( .A(n2409), .B(n2410), .Z(n2408) );
  XNOR U3491 ( .A(y[712]), .B(x[712]), .Z(n2410) );
  XNOR U3492 ( .A(y[713]), .B(x[713]), .Z(n2409) );
  XNOR U3493 ( .A(y[711]), .B(x[711]), .Z(n2407) );
  XNOR U3494 ( .A(n2401), .B(n2402), .Z(n2412) );
  XNOR U3495 ( .A(y[708]), .B(x[708]), .Z(n2402) );
  XNOR U3496 ( .A(n2403), .B(n2404), .Z(n2401) );
  XNOR U3497 ( .A(y[709]), .B(x[709]), .Z(n2404) );
  XNOR U3498 ( .A(y[710]), .B(x[710]), .Z(n2403) );
  XOR U3499 ( .A(n2395), .B(n2394), .Z(n2396) );
  XNOR U3500 ( .A(n2390), .B(n2391), .Z(n2394) );
  XNOR U3501 ( .A(y[705]), .B(x[705]), .Z(n2391) );
  XNOR U3502 ( .A(n2392), .B(n2393), .Z(n2390) );
  XNOR U3503 ( .A(y[706]), .B(x[706]), .Z(n2393) );
  XNOR U3504 ( .A(y[707]), .B(x[707]), .Z(n2392) );
  XNOR U3505 ( .A(n2384), .B(n2385), .Z(n2395) );
  XNOR U3506 ( .A(y[702]), .B(x[702]), .Z(n2385) );
  XNOR U3507 ( .A(n2386), .B(n2387), .Z(n2384) );
  XNOR U3508 ( .A(y[703]), .B(x[703]), .Z(n2387) );
  XNOR U3509 ( .A(y[704]), .B(x[704]), .Z(n2386) );
  NAND U3510 ( .A(n2451), .B(n2452), .Z(N6078) );
  NANDN U3511 ( .A(n2453), .B(n2454), .Z(n2452) );
  OR U3512 ( .A(n2455), .B(n2456), .Z(n2454) );
  NAND U3513 ( .A(n2455), .B(n2456), .Z(n2451) );
  XOR U3514 ( .A(n2455), .B(n2457), .Z(N6077) );
  XNOR U3515 ( .A(n2453), .B(n2456), .Z(n2457) );
  AND U3516 ( .A(n2458), .B(n2459), .Z(n2456) );
  NANDN U3517 ( .A(n2460), .B(n2461), .Z(n2459) );
  NANDN U3518 ( .A(n2462), .B(n2463), .Z(n2461) );
  NANDN U3519 ( .A(n2463), .B(n2462), .Z(n2458) );
  NAND U3520 ( .A(n2464), .B(n2465), .Z(n2453) );
  NANDN U3521 ( .A(n2466), .B(n2467), .Z(n2465) );
  OR U3522 ( .A(n2468), .B(n2469), .Z(n2467) );
  NAND U3523 ( .A(n2469), .B(n2468), .Z(n2464) );
  AND U3524 ( .A(n2470), .B(n2471), .Z(n2455) );
  NANDN U3525 ( .A(n2472), .B(n2473), .Z(n2471) );
  NANDN U3526 ( .A(n2474), .B(n2475), .Z(n2473) );
  NANDN U3527 ( .A(n2475), .B(n2474), .Z(n2470) );
  XOR U3528 ( .A(n2469), .B(n2476), .Z(N6076) );
  XOR U3529 ( .A(n2466), .B(n2468), .Z(n2476) );
  XNOR U3530 ( .A(n2462), .B(n2477), .Z(n2468) );
  XNOR U3531 ( .A(n2460), .B(n2463), .Z(n2477) );
  NAND U3532 ( .A(n2478), .B(n2479), .Z(n2463) );
  NAND U3533 ( .A(n2480), .B(n2481), .Z(n2479) );
  OR U3534 ( .A(n2482), .B(n2483), .Z(n2480) );
  NANDN U3535 ( .A(n2484), .B(n2482), .Z(n2478) );
  IV U3536 ( .A(n2483), .Z(n2484) );
  NAND U3537 ( .A(n2485), .B(n2486), .Z(n2460) );
  NAND U3538 ( .A(n2487), .B(n2488), .Z(n2486) );
  NANDN U3539 ( .A(n2489), .B(n2490), .Z(n2487) );
  NANDN U3540 ( .A(n2490), .B(n2489), .Z(n2485) );
  AND U3541 ( .A(n2491), .B(n2492), .Z(n2462) );
  NAND U3542 ( .A(n2493), .B(n2494), .Z(n2492) );
  OR U3543 ( .A(n2495), .B(n2496), .Z(n2493) );
  NANDN U3544 ( .A(n2497), .B(n2495), .Z(n2491) );
  NAND U3545 ( .A(n2498), .B(n2499), .Z(n2466) );
  NANDN U3546 ( .A(n2500), .B(n2501), .Z(n2499) );
  OR U3547 ( .A(n2502), .B(n2503), .Z(n2501) );
  NANDN U3548 ( .A(n2504), .B(n2502), .Z(n2498) );
  IV U3549 ( .A(n2503), .Z(n2504) );
  XNOR U3550 ( .A(n2474), .B(n2505), .Z(n2469) );
  XNOR U3551 ( .A(n2472), .B(n2475), .Z(n2505) );
  NAND U3552 ( .A(n2506), .B(n2507), .Z(n2475) );
  NAND U3553 ( .A(n2508), .B(n2509), .Z(n2507) );
  OR U3554 ( .A(n2510), .B(n2511), .Z(n2508) );
  NANDN U3555 ( .A(n2512), .B(n2510), .Z(n2506) );
  IV U3556 ( .A(n2511), .Z(n2512) );
  NAND U3557 ( .A(n2513), .B(n2514), .Z(n2472) );
  NAND U3558 ( .A(n2515), .B(n2516), .Z(n2514) );
  NANDN U3559 ( .A(n2517), .B(n2518), .Z(n2515) );
  NANDN U3560 ( .A(n2518), .B(n2517), .Z(n2513) );
  AND U3561 ( .A(n2519), .B(n2520), .Z(n2474) );
  NAND U3562 ( .A(n2521), .B(n2522), .Z(n2520) );
  OR U3563 ( .A(n2523), .B(n2524), .Z(n2521) );
  NANDN U3564 ( .A(n2525), .B(n2523), .Z(n2519) );
  XNOR U3565 ( .A(n2500), .B(n2526), .Z(N6075) );
  XOR U3566 ( .A(n2502), .B(n2503), .Z(n2526) );
  XNOR U3567 ( .A(n2516), .B(n2527), .Z(n2503) );
  XOR U3568 ( .A(n2517), .B(n2518), .Z(n2527) );
  XOR U3569 ( .A(n2523), .B(n2528), .Z(n2518) );
  XOR U3570 ( .A(n2522), .B(n2525), .Z(n2528) );
  IV U3571 ( .A(n2524), .Z(n2525) );
  NAND U3572 ( .A(n2529), .B(n2530), .Z(n2524) );
  OR U3573 ( .A(n2531), .B(n2532), .Z(n2530) );
  OR U3574 ( .A(n2533), .B(n2534), .Z(n2529) );
  NAND U3575 ( .A(n2535), .B(n2536), .Z(n2522) );
  OR U3576 ( .A(n2537), .B(n2538), .Z(n2536) );
  OR U3577 ( .A(n2539), .B(n2540), .Z(n2535) );
  NOR U3578 ( .A(n2541), .B(n2542), .Z(n2523) );
  ANDN U3579 ( .B(n2543), .A(n2544), .Z(n2517) );
  XNOR U3580 ( .A(n2510), .B(n2545), .Z(n2516) );
  XNOR U3581 ( .A(n2509), .B(n2511), .Z(n2545) );
  NAND U3582 ( .A(n2546), .B(n2547), .Z(n2511) );
  OR U3583 ( .A(n2548), .B(n2549), .Z(n2547) );
  OR U3584 ( .A(n2550), .B(n2551), .Z(n2546) );
  NAND U3585 ( .A(n2552), .B(n2553), .Z(n2509) );
  OR U3586 ( .A(n2554), .B(n2555), .Z(n2553) );
  OR U3587 ( .A(n2556), .B(n2557), .Z(n2552) );
  ANDN U3588 ( .B(n2558), .A(n2559), .Z(n2510) );
  IV U3589 ( .A(n2560), .Z(n2558) );
  ANDN U3590 ( .B(n2561), .A(n2562), .Z(n2502) );
  XOR U3591 ( .A(n2488), .B(n2563), .Z(n2500) );
  XOR U3592 ( .A(n2489), .B(n2490), .Z(n2563) );
  XOR U3593 ( .A(n2495), .B(n2564), .Z(n2490) );
  XOR U3594 ( .A(n2494), .B(n2497), .Z(n2564) );
  IV U3595 ( .A(n2496), .Z(n2497) );
  NAND U3596 ( .A(n2565), .B(n2566), .Z(n2496) );
  OR U3597 ( .A(n2567), .B(n2568), .Z(n2566) );
  OR U3598 ( .A(n2569), .B(n2570), .Z(n2565) );
  NAND U3599 ( .A(n2571), .B(n2572), .Z(n2494) );
  OR U3600 ( .A(n2573), .B(n2574), .Z(n2572) );
  OR U3601 ( .A(n2575), .B(n2576), .Z(n2571) );
  NOR U3602 ( .A(n2577), .B(n2578), .Z(n2495) );
  ANDN U3603 ( .B(n2579), .A(n2580), .Z(n2489) );
  IV U3604 ( .A(n2581), .Z(n2579) );
  XNOR U3605 ( .A(n2482), .B(n2582), .Z(n2488) );
  XNOR U3606 ( .A(n2481), .B(n2483), .Z(n2582) );
  NAND U3607 ( .A(n2583), .B(n2584), .Z(n2483) );
  OR U3608 ( .A(n2585), .B(n2586), .Z(n2584) );
  OR U3609 ( .A(n2587), .B(n2588), .Z(n2583) );
  NAND U3610 ( .A(n2589), .B(n2590), .Z(n2481) );
  OR U3611 ( .A(n2591), .B(n2592), .Z(n2590) );
  OR U3612 ( .A(n2593), .B(n2594), .Z(n2589) );
  ANDN U3613 ( .B(n2595), .A(n2596), .Z(n2482) );
  IV U3614 ( .A(n2597), .Z(n2595) );
  XNOR U3615 ( .A(n2562), .B(n2561), .Z(N6074) );
  XOR U3616 ( .A(n2581), .B(n2580), .Z(n2561) );
  XNOR U3617 ( .A(n2596), .B(n2597), .Z(n2580) );
  XNOR U3618 ( .A(n2591), .B(n2592), .Z(n2597) );
  XNOR U3619 ( .A(n2593), .B(n2594), .Z(n2592) );
  XNOR U3620 ( .A(y[700]), .B(x[700]), .Z(n2594) );
  XNOR U3621 ( .A(y[701]), .B(x[701]), .Z(n2593) );
  XNOR U3622 ( .A(y[699]), .B(x[699]), .Z(n2591) );
  XNOR U3623 ( .A(n2585), .B(n2586), .Z(n2596) );
  XNOR U3624 ( .A(y[696]), .B(x[696]), .Z(n2586) );
  XNOR U3625 ( .A(n2587), .B(n2588), .Z(n2585) );
  XNOR U3626 ( .A(y[697]), .B(x[697]), .Z(n2588) );
  XNOR U3627 ( .A(y[698]), .B(x[698]), .Z(n2587) );
  XNOR U3628 ( .A(n2578), .B(n2577), .Z(n2581) );
  XNOR U3629 ( .A(n2573), .B(n2574), .Z(n2577) );
  XNOR U3630 ( .A(y[693]), .B(x[693]), .Z(n2574) );
  XNOR U3631 ( .A(n2575), .B(n2576), .Z(n2573) );
  XNOR U3632 ( .A(y[694]), .B(x[694]), .Z(n2576) );
  XNOR U3633 ( .A(y[695]), .B(x[695]), .Z(n2575) );
  XNOR U3634 ( .A(n2567), .B(n2568), .Z(n2578) );
  XNOR U3635 ( .A(y[690]), .B(x[690]), .Z(n2568) );
  XNOR U3636 ( .A(n2569), .B(n2570), .Z(n2567) );
  XNOR U3637 ( .A(y[691]), .B(x[691]), .Z(n2570) );
  XNOR U3638 ( .A(y[692]), .B(x[692]), .Z(n2569) );
  XOR U3639 ( .A(n2543), .B(n2544), .Z(n2562) );
  XNOR U3640 ( .A(n2559), .B(n2560), .Z(n2544) );
  XNOR U3641 ( .A(n2554), .B(n2555), .Z(n2560) );
  XNOR U3642 ( .A(n2556), .B(n2557), .Z(n2555) );
  XNOR U3643 ( .A(y[688]), .B(x[688]), .Z(n2557) );
  XNOR U3644 ( .A(y[689]), .B(x[689]), .Z(n2556) );
  XNOR U3645 ( .A(y[687]), .B(x[687]), .Z(n2554) );
  XNOR U3646 ( .A(n2548), .B(n2549), .Z(n2559) );
  XNOR U3647 ( .A(y[684]), .B(x[684]), .Z(n2549) );
  XNOR U3648 ( .A(n2550), .B(n2551), .Z(n2548) );
  XNOR U3649 ( .A(y[685]), .B(x[685]), .Z(n2551) );
  XNOR U3650 ( .A(y[686]), .B(x[686]), .Z(n2550) );
  XOR U3651 ( .A(n2542), .B(n2541), .Z(n2543) );
  XNOR U3652 ( .A(n2537), .B(n2538), .Z(n2541) );
  XNOR U3653 ( .A(y[681]), .B(x[681]), .Z(n2538) );
  XNOR U3654 ( .A(n2539), .B(n2540), .Z(n2537) );
  XNOR U3655 ( .A(y[682]), .B(x[682]), .Z(n2540) );
  XNOR U3656 ( .A(y[683]), .B(x[683]), .Z(n2539) );
  XNOR U3657 ( .A(n2531), .B(n2532), .Z(n2542) );
  XNOR U3658 ( .A(y[678]), .B(x[678]), .Z(n2532) );
  XNOR U3659 ( .A(n2533), .B(n2534), .Z(n2531) );
  XNOR U3660 ( .A(y[679]), .B(x[679]), .Z(n2534) );
  XNOR U3661 ( .A(y[680]), .B(x[680]), .Z(n2533) );
  NAND U3662 ( .A(n2598), .B(n2599), .Z(N6068) );
  NANDN U3663 ( .A(n2600), .B(n2601), .Z(n2599) );
  OR U3664 ( .A(n2602), .B(n2603), .Z(n2601) );
  NAND U3665 ( .A(n2602), .B(n2603), .Z(n2598) );
  XOR U3666 ( .A(n2602), .B(n2604), .Z(N6067) );
  XNOR U3667 ( .A(n2600), .B(n2603), .Z(n2604) );
  AND U3668 ( .A(n2605), .B(n2606), .Z(n2603) );
  NANDN U3669 ( .A(n2607), .B(n2608), .Z(n2606) );
  NANDN U3670 ( .A(n2609), .B(n2610), .Z(n2608) );
  NANDN U3671 ( .A(n2610), .B(n2609), .Z(n2605) );
  NAND U3672 ( .A(n2611), .B(n2612), .Z(n2600) );
  NANDN U3673 ( .A(n2613), .B(n2614), .Z(n2612) );
  OR U3674 ( .A(n2615), .B(n2616), .Z(n2614) );
  NAND U3675 ( .A(n2616), .B(n2615), .Z(n2611) );
  AND U3676 ( .A(n2617), .B(n2618), .Z(n2602) );
  NANDN U3677 ( .A(n2619), .B(n2620), .Z(n2618) );
  NANDN U3678 ( .A(n2621), .B(n2622), .Z(n2620) );
  NANDN U3679 ( .A(n2622), .B(n2621), .Z(n2617) );
  XOR U3680 ( .A(n2616), .B(n2623), .Z(N6066) );
  XOR U3681 ( .A(n2613), .B(n2615), .Z(n2623) );
  XNOR U3682 ( .A(n2609), .B(n2624), .Z(n2615) );
  XNOR U3683 ( .A(n2607), .B(n2610), .Z(n2624) );
  NAND U3684 ( .A(n2625), .B(n2626), .Z(n2610) );
  NAND U3685 ( .A(n2627), .B(n2628), .Z(n2626) );
  OR U3686 ( .A(n2629), .B(n2630), .Z(n2627) );
  NANDN U3687 ( .A(n2631), .B(n2629), .Z(n2625) );
  IV U3688 ( .A(n2630), .Z(n2631) );
  NAND U3689 ( .A(n2632), .B(n2633), .Z(n2607) );
  NAND U3690 ( .A(n2634), .B(n2635), .Z(n2633) );
  NANDN U3691 ( .A(n2636), .B(n2637), .Z(n2634) );
  NANDN U3692 ( .A(n2637), .B(n2636), .Z(n2632) );
  AND U3693 ( .A(n2638), .B(n2639), .Z(n2609) );
  NAND U3694 ( .A(n2640), .B(n2641), .Z(n2639) );
  OR U3695 ( .A(n2642), .B(n2643), .Z(n2640) );
  NANDN U3696 ( .A(n2644), .B(n2642), .Z(n2638) );
  NAND U3697 ( .A(n2645), .B(n2646), .Z(n2613) );
  NANDN U3698 ( .A(n2647), .B(n2648), .Z(n2646) );
  OR U3699 ( .A(n2649), .B(n2650), .Z(n2648) );
  NANDN U3700 ( .A(n2651), .B(n2649), .Z(n2645) );
  IV U3701 ( .A(n2650), .Z(n2651) );
  XNOR U3702 ( .A(n2621), .B(n2652), .Z(n2616) );
  XNOR U3703 ( .A(n2619), .B(n2622), .Z(n2652) );
  NAND U3704 ( .A(n2653), .B(n2654), .Z(n2622) );
  NAND U3705 ( .A(n2655), .B(n2656), .Z(n2654) );
  OR U3706 ( .A(n2657), .B(n2658), .Z(n2655) );
  NANDN U3707 ( .A(n2659), .B(n2657), .Z(n2653) );
  IV U3708 ( .A(n2658), .Z(n2659) );
  NAND U3709 ( .A(n2660), .B(n2661), .Z(n2619) );
  NAND U3710 ( .A(n2662), .B(n2663), .Z(n2661) );
  NANDN U3711 ( .A(n2664), .B(n2665), .Z(n2662) );
  NANDN U3712 ( .A(n2665), .B(n2664), .Z(n2660) );
  AND U3713 ( .A(n2666), .B(n2667), .Z(n2621) );
  NAND U3714 ( .A(n2668), .B(n2669), .Z(n2667) );
  OR U3715 ( .A(n2670), .B(n2671), .Z(n2668) );
  NANDN U3716 ( .A(n2672), .B(n2670), .Z(n2666) );
  XNOR U3717 ( .A(n2647), .B(n2673), .Z(N6065) );
  XOR U3718 ( .A(n2649), .B(n2650), .Z(n2673) );
  XNOR U3719 ( .A(n2663), .B(n2674), .Z(n2650) );
  XOR U3720 ( .A(n2664), .B(n2665), .Z(n2674) );
  XOR U3721 ( .A(n2670), .B(n2675), .Z(n2665) );
  XOR U3722 ( .A(n2669), .B(n2672), .Z(n2675) );
  IV U3723 ( .A(n2671), .Z(n2672) );
  NAND U3724 ( .A(n2676), .B(n2677), .Z(n2671) );
  OR U3725 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U3726 ( .A(n2680), .B(n2681), .Z(n2676) );
  NAND U3727 ( .A(n2682), .B(n2683), .Z(n2669) );
  OR U3728 ( .A(n2684), .B(n2685), .Z(n2683) );
  OR U3729 ( .A(n2686), .B(n2687), .Z(n2682) );
  NOR U3730 ( .A(n2688), .B(n2689), .Z(n2670) );
  ANDN U3731 ( .B(n2690), .A(n2691), .Z(n2664) );
  XNOR U3732 ( .A(n2657), .B(n2692), .Z(n2663) );
  XNOR U3733 ( .A(n2656), .B(n2658), .Z(n2692) );
  NAND U3734 ( .A(n2693), .B(n2694), .Z(n2658) );
  OR U3735 ( .A(n2695), .B(n2696), .Z(n2694) );
  OR U3736 ( .A(n2697), .B(n2698), .Z(n2693) );
  NAND U3737 ( .A(n2699), .B(n2700), .Z(n2656) );
  OR U3738 ( .A(n2701), .B(n2702), .Z(n2700) );
  OR U3739 ( .A(n2703), .B(n2704), .Z(n2699) );
  ANDN U3740 ( .B(n2705), .A(n2706), .Z(n2657) );
  IV U3741 ( .A(n2707), .Z(n2705) );
  ANDN U3742 ( .B(n2708), .A(n2709), .Z(n2649) );
  XOR U3743 ( .A(n2635), .B(n2710), .Z(n2647) );
  XOR U3744 ( .A(n2636), .B(n2637), .Z(n2710) );
  XOR U3745 ( .A(n2642), .B(n2711), .Z(n2637) );
  XOR U3746 ( .A(n2641), .B(n2644), .Z(n2711) );
  IV U3747 ( .A(n2643), .Z(n2644) );
  NAND U3748 ( .A(n2712), .B(n2713), .Z(n2643) );
  OR U3749 ( .A(n2714), .B(n2715), .Z(n2713) );
  OR U3750 ( .A(n2716), .B(n2717), .Z(n2712) );
  NAND U3751 ( .A(n2718), .B(n2719), .Z(n2641) );
  OR U3752 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U3753 ( .A(n2722), .B(n2723), .Z(n2718) );
  NOR U3754 ( .A(n2724), .B(n2725), .Z(n2642) );
  ANDN U3755 ( .B(n2726), .A(n2727), .Z(n2636) );
  IV U3756 ( .A(n2728), .Z(n2726) );
  XNOR U3757 ( .A(n2629), .B(n2729), .Z(n2635) );
  XNOR U3758 ( .A(n2628), .B(n2630), .Z(n2729) );
  NAND U3759 ( .A(n2730), .B(n2731), .Z(n2630) );
  OR U3760 ( .A(n2732), .B(n2733), .Z(n2731) );
  OR U3761 ( .A(n2734), .B(n2735), .Z(n2730) );
  NAND U3762 ( .A(n2736), .B(n2737), .Z(n2628) );
  OR U3763 ( .A(n2738), .B(n2739), .Z(n2737) );
  OR U3764 ( .A(n2740), .B(n2741), .Z(n2736) );
  ANDN U3765 ( .B(n2742), .A(n2743), .Z(n2629) );
  IV U3766 ( .A(n2744), .Z(n2742) );
  XNOR U3767 ( .A(n2709), .B(n2708), .Z(N6064) );
  XOR U3768 ( .A(n2728), .B(n2727), .Z(n2708) );
  XNOR U3769 ( .A(n2743), .B(n2744), .Z(n2727) );
  XNOR U3770 ( .A(n2738), .B(n2739), .Z(n2744) );
  XNOR U3771 ( .A(n2740), .B(n2741), .Z(n2739) );
  XNOR U3772 ( .A(y[676]), .B(x[676]), .Z(n2741) );
  XNOR U3773 ( .A(y[677]), .B(x[677]), .Z(n2740) );
  XNOR U3774 ( .A(y[675]), .B(x[675]), .Z(n2738) );
  XNOR U3775 ( .A(n2732), .B(n2733), .Z(n2743) );
  XNOR U3776 ( .A(y[672]), .B(x[672]), .Z(n2733) );
  XNOR U3777 ( .A(n2734), .B(n2735), .Z(n2732) );
  XNOR U3778 ( .A(y[673]), .B(x[673]), .Z(n2735) );
  XNOR U3779 ( .A(y[674]), .B(x[674]), .Z(n2734) );
  XNOR U3780 ( .A(n2725), .B(n2724), .Z(n2728) );
  XNOR U3781 ( .A(n2720), .B(n2721), .Z(n2724) );
  XNOR U3782 ( .A(y[669]), .B(x[669]), .Z(n2721) );
  XNOR U3783 ( .A(n2722), .B(n2723), .Z(n2720) );
  XNOR U3784 ( .A(y[670]), .B(x[670]), .Z(n2723) );
  XNOR U3785 ( .A(y[671]), .B(x[671]), .Z(n2722) );
  XNOR U3786 ( .A(n2714), .B(n2715), .Z(n2725) );
  XNOR U3787 ( .A(y[666]), .B(x[666]), .Z(n2715) );
  XNOR U3788 ( .A(n2716), .B(n2717), .Z(n2714) );
  XNOR U3789 ( .A(y[667]), .B(x[667]), .Z(n2717) );
  XNOR U3790 ( .A(y[668]), .B(x[668]), .Z(n2716) );
  XOR U3791 ( .A(n2690), .B(n2691), .Z(n2709) );
  XNOR U3792 ( .A(n2706), .B(n2707), .Z(n2691) );
  XNOR U3793 ( .A(n2701), .B(n2702), .Z(n2707) );
  XNOR U3794 ( .A(n2703), .B(n2704), .Z(n2702) );
  XNOR U3795 ( .A(y[664]), .B(x[664]), .Z(n2704) );
  XNOR U3796 ( .A(y[665]), .B(x[665]), .Z(n2703) );
  XNOR U3797 ( .A(y[663]), .B(x[663]), .Z(n2701) );
  XNOR U3798 ( .A(n2695), .B(n2696), .Z(n2706) );
  XNOR U3799 ( .A(y[660]), .B(x[660]), .Z(n2696) );
  XNOR U3800 ( .A(n2697), .B(n2698), .Z(n2695) );
  XNOR U3801 ( .A(y[661]), .B(x[661]), .Z(n2698) );
  XNOR U3802 ( .A(y[662]), .B(x[662]), .Z(n2697) );
  XOR U3803 ( .A(n2689), .B(n2688), .Z(n2690) );
  XNOR U3804 ( .A(n2684), .B(n2685), .Z(n2688) );
  XNOR U3805 ( .A(y[657]), .B(x[657]), .Z(n2685) );
  XNOR U3806 ( .A(n2686), .B(n2687), .Z(n2684) );
  XNOR U3807 ( .A(y[658]), .B(x[658]), .Z(n2687) );
  XNOR U3808 ( .A(y[659]), .B(x[659]), .Z(n2686) );
  XNOR U3809 ( .A(n2678), .B(n2679), .Z(n2689) );
  XNOR U3810 ( .A(y[654]), .B(x[654]), .Z(n2679) );
  XNOR U3811 ( .A(n2680), .B(n2681), .Z(n2678) );
  XNOR U3812 ( .A(y[655]), .B(x[655]), .Z(n2681) );
  XNOR U3813 ( .A(y[656]), .B(x[656]), .Z(n2680) );
  NAND U3814 ( .A(n2745), .B(n2746), .Z(N6058) );
  NANDN U3815 ( .A(n2747), .B(n2748), .Z(n2746) );
  OR U3816 ( .A(n2749), .B(n2750), .Z(n2748) );
  NAND U3817 ( .A(n2749), .B(n2750), .Z(n2745) );
  XOR U3818 ( .A(n2749), .B(n2751), .Z(N6057) );
  XNOR U3819 ( .A(n2747), .B(n2750), .Z(n2751) );
  AND U3820 ( .A(n2752), .B(n2753), .Z(n2750) );
  NANDN U3821 ( .A(n2754), .B(n2755), .Z(n2753) );
  NANDN U3822 ( .A(n2756), .B(n2757), .Z(n2755) );
  NANDN U3823 ( .A(n2757), .B(n2756), .Z(n2752) );
  NAND U3824 ( .A(n2758), .B(n2759), .Z(n2747) );
  NANDN U3825 ( .A(n2760), .B(n2761), .Z(n2759) );
  OR U3826 ( .A(n2762), .B(n2763), .Z(n2761) );
  NAND U3827 ( .A(n2763), .B(n2762), .Z(n2758) );
  AND U3828 ( .A(n2764), .B(n2765), .Z(n2749) );
  NANDN U3829 ( .A(n2766), .B(n2767), .Z(n2765) );
  NANDN U3830 ( .A(n2768), .B(n2769), .Z(n2767) );
  NANDN U3831 ( .A(n2769), .B(n2768), .Z(n2764) );
  XOR U3832 ( .A(n2763), .B(n2770), .Z(N6056) );
  XOR U3833 ( .A(n2760), .B(n2762), .Z(n2770) );
  XNOR U3834 ( .A(n2756), .B(n2771), .Z(n2762) );
  XNOR U3835 ( .A(n2754), .B(n2757), .Z(n2771) );
  NAND U3836 ( .A(n2772), .B(n2773), .Z(n2757) );
  NAND U3837 ( .A(n2774), .B(n2775), .Z(n2773) );
  OR U3838 ( .A(n2776), .B(n2777), .Z(n2774) );
  NANDN U3839 ( .A(n2778), .B(n2776), .Z(n2772) );
  IV U3840 ( .A(n2777), .Z(n2778) );
  NAND U3841 ( .A(n2779), .B(n2780), .Z(n2754) );
  NAND U3842 ( .A(n2781), .B(n2782), .Z(n2780) );
  NANDN U3843 ( .A(n2783), .B(n2784), .Z(n2781) );
  NANDN U3844 ( .A(n2784), .B(n2783), .Z(n2779) );
  AND U3845 ( .A(n2785), .B(n2786), .Z(n2756) );
  NAND U3846 ( .A(n2787), .B(n2788), .Z(n2786) );
  OR U3847 ( .A(n2789), .B(n2790), .Z(n2787) );
  NANDN U3848 ( .A(n2791), .B(n2789), .Z(n2785) );
  NAND U3849 ( .A(n2792), .B(n2793), .Z(n2760) );
  NANDN U3850 ( .A(n2794), .B(n2795), .Z(n2793) );
  OR U3851 ( .A(n2796), .B(n2797), .Z(n2795) );
  NANDN U3852 ( .A(n2798), .B(n2796), .Z(n2792) );
  IV U3853 ( .A(n2797), .Z(n2798) );
  XNOR U3854 ( .A(n2768), .B(n2799), .Z(n2763) );
  XNOR U3855 ( .A(n2766), .B(n2769), .Z(n2799) );
  NAND U3856 ( .A(n2800), .B(n2801), .Z(n2769) );
  NAND U3857 ( .A(n2802), .B(n2803), .Z(n2801) );
  OR U3858 ( .A(n2804), .B(n2805), .Z(n2802) );
  NANDN U3859 ( .A(n2806), .B(n2804), .Z(n2800) );
  IV U3860 ( .A(n2805), .Z(n2806) );
  NAND U3861 ( .A(n2807), .B(n2808), .Z(n2766) );
  NAND U3862 ( .A(n2809), .B(n2810), .Z(n2808) );
  NANDN U3863 ( .A(n2811), .B(n2812), .Z(n2809) );
  NANDN U3864 ( .A(n2812), .B(n2811), .Z(n2807) );
  AND U3865 ( .A(n2813), .B(n2814), .Z(n2768) );
  NAND U3866 ( .A(n2815), .B(n2816), .Z(n2814) );
  OR U3867 ( .A(n2817), .B(n2818), .Z(n2815) );
  NANDN U3868 ( .A(n2819), .B(n2817), .Z(n2813) );
  XNOR U3869 ( .A(n2794), .B(n2820), .Z(N6055) );
  XOR U3870 ( .A(n2796), .B(n2797), .Z(n2820) );
  XNOR U3871 ( .A(n2810), .B(n2821), .Z(n2797) );
  XOR U3872 ( .A(n2811), .B(n2812), .Z(n2821) );
  XOR U3873 ( .A(n2817), .B(n2822), .Z(n2812) );
  XOR U3874 ( .A(n2816), .B(n2819), .Z(n2822) );
  IV U3875 ( .A(n2818), .Z(n2819) );
  NAND U3876 ( .A(n2823), .B(n2824), .Z(n2818) );
  OR U3877 ( .A(n2825), .B(n2826), .Z(n2824) );
  OR U3878 ( .A(n2827), .B(n2828), .Z(n2823) );
  NAND U3879 ( .A(n2829), .B(n2830), .Z(n2816) );
  OR U3880 ( .A(n2831), .B(n2832), .Z(n2830) );
  OR U3881 ( .A(n2833), .B(n2834), .Z(n2829) );
  NOR U3882 ( .A(n2835), .B(n2836), .Z(n2817) );
  ANDN U3883 ( .B(n2837), .A(n2838), .Z(n2811) );
  XNOR U3884 ( .A(n2804), .B(n2839), .Z(n2810) );
  XNOR U3885 ( .A(n2803), .B(n2805), .Z(n2839) );
  NAND U3886 ( .A(n2840), .B(n2841), .Z(n2805) );
  OR U3887 ( .A(n2842), .B(n2843), .Z(n2841) );
  OR U3888 ( .A(n2844), .B(n2845), .Z(n2840) );
  NAND U3889 ( .A(n2846), .B(n2847), .Z(n2803) );
  OR U3890 ( .A(n2848), .B(n2849), .Z(n2847) );
  OR U3891 ( .A(n2850), .B(n2851), .Z(n2846) );
  ANDN U3892 ( .B(n2852), .A(n2853), .Z(n2804) );
  IV U3893 ( .A(n2854), .Z(n2852) );
  ANDN U3894 ( .B(n2855), .A(n2856), .Z(n2796) );
  XOR U3895 ( .A(n2782), .B(n2857), .Z(n2794) );
  XOR U3896 ( .A(n2783), .B(n2784), .Z(n2857) );
  XOR U3897 ( .A(n2789), .B(n2858), .Z(n2784) );
  XOR U3898 ( .A(n2788), .B(n2791), .Z(n2858) );
  IV U3899 ( .A(n2790), .Z(n2791) );
  NAND U3900 ( .A(n2859), .B(n2860), .Z(n2790) );
  OR U3901 ( .A(n2861), .B(n2862), .Z(n2860) );
  OR U3902 ( .A(n2863), .B(n2864), .Z(n2859) );
  NAND U3903 ( .A(n2865), .B(n2866), .Z(n2788) );
  OR U3904 ( .A(n2867), .B(n2868), .Z(n2866) );
  OR U3905 ( .A(n2869), .B(n2870), .Z(n2865) );
  NOR U3906 ( .A(n2871), .B(n2872), .Z(n2789) );
  ANDN U3907 ( .B(n2873), .A(n2874), .Z(n2783) );
  IV U3908 ( .A(n2875), .Z(n2873) );
  XNOR U3909 ( .A(n2776), .B(n2876), .Z(n2782) );
  XNOR U3910 ( .A(n2775), .B(n2777), .Z(n2876) );
  NAND U3911 ( .A(n2877), .B(n2878), .Z(n2777) );
  OR U3912 ( .A(n2879), .B(n2880), .Z(n2878) );
  OR U3913 ( .A(n2881), .B(n2882), .Z(n2877) );
  NAND U3914 ( .A(n2883), .B(n2884), .Z(n2775) );
  OR U3915 ( .A(n2885), .B(n2886), .Z(n2884) );
  OR U3916 ( .A(n2887), .B(n2888), .Z(n2883) );
  ANDN U3917 ( .B(n2889), .A(n2890), .Z(n2776) );
  IV U3918 ( .A(n2891), .Z(n2889) );
  XNOR U3919 ( .A(n2856), .B(n2855), .Z(N6054) );
  XOR U3920 ( .A(n2875), .B(n2874), .Z(n2855) );
  XNOR U3921 ( .A(n2890), .B(n2891), .Z(n2874) );
  XNOR U3922 ( .A(n2885), .B(n2886), .Z(n2891) );
  XNOR U3923 ( .A(n2887), .B(n2888), .Z(n2886) );
  XNOR U3924 ( .A(y[652]), .B(x[652]), .Z(n2888) );
  XNOR U3925 ( .A(y[653]), .B(x[653]), .Z(n2887) );
  XNOR U3926 ( .A(y[651]), .B(x[651]), .Z(n2885) );
  XNOR U3927 ( .A(n2879), .B(n2880), .Z(n2890) );
  XNOR U3928 ( .A(y[648]), .B(x[648]), .Z(n2880) );
  XNOR U3929 ( .A(n2881), .B(n2882), .Z(n2879) );
  XNOR U3930 ( .A(y[649]), .B(x[649]), .Z(n2882) );
  XNOR U3931 ( .A(y[650]), .B(x[650]), .Z(n2881) );
  XNOR U3932 ( .A(n2872), .B(n2871), .Z(n2875) );
  XNOR U3933 ( .A(n2867), .B(n2868), .Z(n2871) );
  XNOR U3934 ( .A(y[645]), .B(x[645]), .Z(n2868) );
  XNOR U3935 ( .A(n2869), .B(n2870), .Z(n2867) );
  XNOR U3936 ( .A(y[646]), .B(x[646]), .Z(n2870) );
  XNOR U3937 ( .A(y[647]), .B(x[647]), .Z(n2869) );
  XNOR U3938 ( .A(n2861), .B(n2862), .Z(n2872) );
  XNOR U3939 ( .A(y[642]), .B(x[642]), .Z(n2862) );
  XNOR U3940 ( .A(n2863), .B(n2864), .Z(n2861) );
  XNOR U3941 ( .A(y[643]), .B(x[643]), .Z(n2864) );
  XNOR U3942 ( .A(y[644]), .B(x[644]), .Z(n2863) );
  XOR U3943 ( .A(n2837), .B(n2838), .Z(n2856) );
  XNOR U3944 ( .A(n2853), .B(n2854), .Z(n2838) );
  XNOR U3945 ( .A(n2848), .B(n2849), .Z(n2854) );
  XNOR U3946 ( .A(n2850), .B(n2851), .Z(n2849) );
  XNOR U3947 ( .A(y[640]), .B(x[640]), .Z(n2851) );
  XNOR U3948 ( .A(y[641]), .B(x[641]), .Z(n2850) );
  XNOR U3949 ( .A(y[639]), .B(x[639]), .Z(n2848) );
  XNOR U3950 ( .A(n2842), .B(n2843), .Z(n2853) );
  XNOR U3951 ( .A(y[636]), .B(x[636]), .Z(n2843) );
  XNOR U3952 ( .A(n2844), .B(n2845), .Z(n2842) );
  XNOR U3953 ( .A(y[637]), .B(x[637]), .Z(n2845) );
  XNOR U3954 ( .A(y[638]), .B(x[638]), .Z(n2844) );
  XOR U3955 ( .A(n2836), .B(n2835), .Z(n2837) );
  XNOR U3956 ( .A(n2831), .B(n2832), .Z(n2835) );
  XNOR U3957 ( .A(y[633]), .B(x[633]), .Z(n2832) );
  XNOR U3958 ( .A(n2833), .B(n2834), .Z(n2831) );
  XNOR U3959 ( .A(y[634]), .B(x[634]), .Z(n2834) );
  XNOR U3960 ( .A(y[635]), .B(x[635]), .Z(n2833) );
  XNOR U3961 ( .A(n2825), .B(n2826), .Z(n2836) );
  XNOR U3962 ( .A(y[630]), .B(x[630]), .Z(n2826) );
  XNOR U3963 ( .A(n2827), .B(n2828), .Z(n2825) );
  XNOR U3964 ( .A(y[631]), .B(x[631]), .Z(n2828) );
  XNOR U3965 ( .A(y[632]), .B(x[632]), .Z(n2827) );
  NAND U3966 ( .A(n2892), .B(n2893), .Z(N6048) );
  NANDN U3967 ( .A(n2894), .B(n2895), .Z(n2893) );
  OR U3968 ( .A(n2896), .B(n2897), .Z(n2895) );
  NAND U3969 ( .A(n2896), .B(n2897), .Z(n2892) );
  XOR U3970 ( .A(n2896), .B(n2898), .Z(N6047) );
  XNOR U3971 ( .A(n2894), .B(n2897), .Z(n2898) );
  AND U3972 ( .A(n2899), .B(n2900), .Z(n2897) );
  NANDN U3973 ( .A(n2901), .B(n2902), .Z(n2900) );
  NANDN U3974 ( .A(n2903), .B(n2904), .Z(n2902) );
  NANDN U3975 ( .A(n2904), .B(n2903), .Z(n2899) );
  NAND U3976 ( .A(n2905), .B(n2906), .Z(n2894) );
  NANDN U3977 ( .A(n2907), .B(n2908), .Z(n2906) );
  OR U3978 ( .A(n2909), .B(n2910), .Z(n2908) );
  NAND U3979 ( .A(n2910), .B(n2909), .Z(n2905) );
  AND U3980 ( .A(n2911), .B(n2912), .Z(n2896) );
  NANDN U3981 ( .A(n2913), .B(n2914), .Z(n2912) );
  NANDN U3982 ( .A(n2915), .B(n2916), .Z(n2914) );
  NANDN U3983 ( .A(n2916), .B(n2915), .Z(n2911) );
  XOR U3984 ( .A(n2910), .B(n2917), .Z(N6046) );
  XOR U3985 ( .A(n2907), .B(n2909), .Z(n2917) );
  XNOR U3986 ( .A(n2903), .B(n2918), .Z(n2909) );
  XNOR U3987 ( .A(n2901), .B(n2904), .Z(n2918) );
  NAND U3988 ( .A(n2919), .B(n2920), .Z(n2904) );
  NAND U3989 ( .A(n2921), .B(n2922), .Z(n2920) );
  OR U3990 ( .A(n2923), .B(n2924), .Z(n2921) );
  NANDN U3991 ( .A(n2925), .B(n2923), .Z(n2919) );
  IV U3992 ( .A(n2924), .Z(n2925) );
  NAND U3993 ( .A(n2926), .B(n2927), .Z(n2901) );
  NAND U3994 ( .A(n2928), .B(n2929), .Z(n2927) );
  NANDN U3995 ( .A(n2930), .B(n2931), .Z(n2928) );
  NANDN U3996 ( .A(n2931), .B(n2930), .Z(n2926) );
  AND U3997 ( .A(n2932), .B(n2933), .Z(n2903) );
  NAND U3998 ( .A(n2934), .B(n2935), .Z(n2933) );
  OR U3999 ( .A(n2936), .B(n2937), .Z(n2934) );
  NANDN U4000 ( .A(n2938), .B(n2936), .Z(n2932) );
  NAND U4001 ( .A(n2939), .B(n2940), .Z(n2907) );
  NANDN U4002 ( .A(n2941), .B(n2942), .Z(n2940) );
  OR U4003 ( .A(n2943), .B(n2944), .Z(n2942) );
  NANDN U4004 ( .A(n2945), .B(n2943), .Z(n2939) );
  IV U4005 ( .A(n2944), .Z(n2945) );
  XNOR U4006 ( .A(n2915), .B(n2946), .Z(n2910) );
  XNOR U4007 ( .A(n2913), .B(n2916), .Z(n2946) );
  NAND U4008 ( .A(n2947), .B(n2948), .Z(n2916) );
  NAND U4009 ( .A(n2949), .B(n2950), .Z(n2948) );
  OR U4010 ( .A(n2951), .B(n2952), .Z(n2949) );
  NANDN U4011 ( .A(n2953), .B(n2951), .Z(n2947) );
  IV U4012 ( .A(n2952), .Z(n2953) );
  NAND U4013 ( .A(n2954), .B(n2955), .Z(n2913) );
  NAND U4014 ( .A(n2956), .B(n2957), .Z(n2955) );
  NANDN U4015 ( .A(n2958), .B(n2959), .Z(n2956) );
  NANDN U4016 ( .A(n2959), .B(n2958), .Z(n2954) );
  AND U4017 ( .A(n2960), .B(n2961), .Z(n2915) );
  NAND U4018 ( .A(n2962), .B(n2963), .Z(n2961) );
  OR U4019 ( .A(n2964), .B(n2965), .Z(n2962) );
  NANDN U4020 ( .A(n2966), .B(n2964), .Z(n2960) );
  XNOR U4021 ( .A(n2941), .B(n2967), .Z(N6045) );
  XOR U4022 ( .A(n2943), .B(n2944), .Z(n2967) );
  XNOR U4023 ( .A(n2957), .B(n2968), .Z(n2944) );
  XOR U4024 ( .A(n2958), .B(n2959), .Z(n2968) );
  XOR U4025 ( .A(n2964), .B(n2969), .Z(n2959) );
  XOR U4026 ( .A(n2963), .B(n2966), .Z(n2969) );
  IV U4027 ( .A(n2965), .Z(n2966) );
  NAND U4028 ( .A(n2970), .B(n2971), .Z(n2965) );
  OR U4029 ( .A(n2972), .B(n2973), .Z(n2971) );
  OR U4030 ( .A(n2974), .B(n2975), .Z(n2970) );
  NAND U4031 ( .A(n2976), .B(n2977), .Z(n2963) );
  OR U4032 ( .A(n2978), .B(n2979), .Z(n2977) );
  OR U4033 ( .A(n2980), .B(n2981), .Z(n2976) );
  NOR U4034 ( .A(n2982), .B(n2983), .Z(n2964) );
  ANDN U4035 ( .B(n2984), .A(n2985), .Z(n2958) );
  XNOR U4036 ( .A(n2951), .B(n2986), .Z(n2957) );
  XNOR U4037 ( .A(n2950), .B(n2952), .Z(n2986) );
  NAND U4038 ( .A(n2987), .B(n2988), .Z(n2952) );
  OR U4039 ( .A(n2989), .B(n2990), .Z(n2988) );
  OR U4040 ( .A(n2991), .B(n2992), .Z(n2987) );
  NAND U4041 ( .A(n2993), .B(n2994), .Z(n2950) );
  OR U4042 ( .A(n2995), .B(n2996), .Z(n2994) );
  OR U4043 ( .A(n2997), .B(n2998), .Z(n2993) );
  ANDN U4044 ( .B(n2999), .A(n3000), .Z(n2951) );
  IV U4045 ( .A(n3001), .Z(n2999) );
  ANDN U4046 ( .B(n3002), .A(n3003), .Z(n2943) );
  XOR U4047 ( .A(n2929), .B(n3004), .Z(n2941) );
  XOR U4048 ( .A(n2930), .B(n2931), .Z(n3004) );
  XOR U4049 ( .A(n2936), .B(n3005), .Z(n2931) );
  XOR U4050 ( .A(n2935), .B(n2938), .Z(n3005) );
  IV U4051 ( .A(n2937), .Z(n2938) );
  NAND U4052 ( .A(n3006), .B(n3007), .Z(n2937) );
  OR U4053 ( .A(n3008), .B(n3009), .Z(n3007) );
  OR U4054 ( .A(n3010), .B(n3011), .Z(n3006) );
  NAND U4055 ( .A(n3012), .B(n3013), .Z(n2935) );
  OR U4056 ( .A(n3014), .B(n3015), .Z(n3013) );
  OR U4057 ( .A(n3016), .B(n3017), .Z(n3012) );
  NOR U4058 ( .A(n3018), .B(n3019), .Z(n2936) );
  ANDN U4059 ( .B(n3020), .A(n3021), .Z(n2930) );
  IV U4060 ( .A(n3022), .Z(n3020) );
  XNOR U4061 ( .A(n2923), .B(n3023), .Z(n2929) );
  XNOR U4062 ( .A(n2922), .B(n2924), .Z(n3023) );
  NAND U4063 ( .A(n3024), .B(n3025), .Z(n2924) );
  OR U4064 ( .A(n3026), .B(n3027), .Z(n3025) );
  OR U4065 ( .A(n3028), .B(n3029), .Z(n3024) );
  NAND U4066 ( .A(n3030), .B(n3031), .Z(n2922) );
  OR U4067 ( .A(n3032), .B(n3033), .Z(n3031) );
  OR U4068 ( .A(n3034), .B(n3035), .Z(n3030) );
  ANDN U4069 ( .B(n3036), .A(n3037), .Z(n2923) );
  IV U4070 ( .A(n3038), .Z(n3036) );
  XNOR U4071 ( .A(n3003), .B(n3002), .Z(N6044) );
  XOR U4072 ( .A(n3022), .B(n3021), .Z(n3002) );
  XNOR U4073 ( .A(n3037), .B(n3038), .Z(n3021) );
  XNOR U4074 ( .A(n3032), .B(n3033), .Z(n3038) );
  XNOR U4075 ( .A(n3034), .B(n3035), .Z(n3033) );
  XNOR U4076 ( .A(y[628]), .B(x[628]), .Z(n3035) );
  XNOR U4077 ( .A(y[629]), .B(x[629]), .Z(n3034) );
  XNOR U4078 ( .A(y[627]), .B(x[627]), .Z(n3032) );
  XNOR U4079 ( .A(n3026), .B(n3027), .Z(n3037) );
  XNOR U4080 ( .A(y[624]), .B(x[624]), .Z(n3027) );
  XNOR U4081 ( .A(n3028), .B(n3029), .Z(n3026) );
  XNOR U4082 ( .A(y[625]), .B(x[625]), .Z(n3029) );
  XNOR U4083 ( .A(y[626]), .B(x[626]), .Z(n3028) );
  XNOR U4084 ( .A(n3019), .B(n3018), .Z(n3022) );
  XNOR U4085 ( .A(n3014), .B(n3015), .Z(n3018) );
  XNOR U4086 ( .A(y[621]), .B(x[621]), .Z(n3015) );
  XNOR U4087 ( .A(n3016), .B(n3017), .Z(n3014) );
  XNOR U4088 ( .A(y[622]), .B(x[622]), .Z(n3017) );
  XNOR U4089 ( .A(y[623]), .B(x[623]), .Z(n3016) );
  XNOR U4090 ( .A(n3008), .B(n3009), .Z(n3019) );
  XNOR U4091 ( .A(y[618]), .B(x[618]), .Z(n3009) );
  XNOR U4092 ( .A(n3010), .B(n3011), .Z(n3008) );
  XNOR U4093 ( .A(y[619]), .B(x[619]), .Z(n3011) );
  XNOR U4094 ( .A(y[620]), .B(x[620]), .Z(n3010) );
  XOR U4095 ( .A(n2984), .B(n2985), .Z(n3003) );
  XNOR U4096 ( .A(n3000), .B(n3001), .Z(n2985) );
  XNOR U4097 ( .A(n2995), .B(n2996), .Z(n3001) );
  XNOR U4098 ( .A(n2997), .B(n2998), .Z(n2996) );
  XNOR U4099 ( .A(y[616]), .B(x[616]), .Z(n2998) );
  XNOR U4100 ( .A(y[617]), .B(x[617]), .Z(n2997) );
  XNOR U4101 ( .A(y[615]), .B(x[615]), .Z(n2995) );
  XNOR U4102 ( .A(n2989), .B(n2990), .Z(n3000) );
  XNOR U4103 ( .A(y[612]), .B(x[612]), .Z(n2990) );
  XNOR U4104 ( .A(n2991), .B(n2992), .Z(n2989) );
  XNOR U4105 ( .A(y[613]), .B(x[613]), .Z(n2992) );
  XNOR U4106 ( .A(y[614]), .B(x[614]), .Z(n2991) );
  XOR U4107 ( .A(n2983), .B(n2982), .Z(n2984) );
  XNOR U4108 ( .A(n2978), .B(n2979), .Z(n2982) );
  XNOR U4109 ( .A(y[609]), .B(x[609]), .Z(n2979) );
  XNOR U4110 ( .A(n2980), .B(n2981), .Z(n2978) );
  XNOR U4111 ( .A(y[610]), .B(x[610]), .Z(n2981) );
  XNOR U4112 ( .A(y[611]), .B(x[611]), .Z(n2980) );
  XNOR U4113 ( .A(n2972), .B(n2973), .Z(n2983) );
  XNOR U4114 ( .A(y[606]), .B(x[606]), .Z(n2973) );
  XNOR U4115 ( .A(n2974), .B(n2975), .Z(n2972) );
  XNOR U4116 ( .A(y[607]), .B(x[607]), .Z(n2975) );
  XNOR U4117 ( .A(y[608]), .B(x[608]), .Z(n2974) );
  NAND U4118 ( .A(n3039), .B(n3040), .Z(N6038) );
  NANDN U4119 ( .A(n3041), .B(n3042), .Z(n3040) );
  OR U4120 ( .A(n3043), .B(n3044), .Z(n3042) );
  NAND U4121 ( .A(n3043), .B(n3044), .Z(n3039) );
  XOR U4122 ( .A(n3043), .B(n3045), .Z(N6037) );
  XNOR U4123 ( .A(n3041), .B(n3044), .Z(n3045) );
  AND U4124 ( .A(n3046), .B(n3047), .Z(n3044) );
  NANDN U4125 ( .A(n3048), .B(n3049), .Z(n3047) );
  NANDN U4126 ( .A(n3050), .B(n3051), .Z(n3049) );
  NANDN U4127 ( .A(n3051), .B(n3050), .Z(n3046) );
  NAND U4128 ( .A(n3052), .B(n3053), .Z(n3041) );
  NANDN U4129 ( .A(n3054), .B(n3055), .Z(n3053) );
  OR U4130 ( .A(n3056), .B(n3057), .Z(n3055) );
  NAND U4131 ( .A(n3057), .B(n3056), .Z(n3052) );
  AND U4132 ( .A(n3058), .B(n3059), .Z(n3043) );
  NANDN U4133 ( .A(n3060), .B(n3061), .Z(n3059) );
  NANDN U4134 ( .A(n3062), .B(n3063), .Z(n3061) );
  NANDN U4135 ( .A(n3063), .B(n3062), .Z(n3058) );
  XOR U4136 ( .A(n3057), .B(n3064), .Z(N6036) );
  XOR U4137 ( .A(n3054), .B(n3056), .Z(n3064) );
  XNOR U4138 ( .A(n3050), .B(n3065), .Z(n3056) );
  XNOR U4139 ( .A(n3048), .B(n3051), .Z(n3065) );
  NAND U4140 ( .A(n3066), .B(n3067), .Z(n3051) );
  NAND U4141 ( .A(n3068), .B(n3069), .Z(n3067) );
  OR U4142 ( .A(n3070), .B(n3071), .Z(n3068) );
  NANDN U4143 ( .A(n3072), .B(n3070), .Z(n3066) );
  IV U4144 ( .A(n3071), .Z(n3072) );
  NAND U4145 ( .A(n3073), .B(n3074), .Z(n3048) );
  NAND U4146 ( .A(n3075), .B(n3076), .Z(n3074) );
  NANDN U4147 ( .A(n3077), .B(n3078), .Z(n3075) );
  NANDN U4148 ( .A(n3078), .B(n3077), .Z(n3073) );
  AND U4149 ( .A(n3079), .B(n3080), .Z(n3050) );
  NAND U4150 ( .A(n3081), .B(n3082), .Z(n3080) );
  OR U4151 ( .A(n3083), .B(n3084), .Z(n3081) );
  NANDN U4152 ( .A(n3085), .B(n3083), .Z(n3079) );
  NAND U4153 ( .A(n3086), .B(n3087), .Z(n3054) );
  NANDN U4154 ( .A(n3088), .B(n3089), .Z(n3087) );
  OR U4155 ( .A(n3090), .B(n3091), .Z(n3089) );
  NANDN U4156 ( .A(n3092), .B(n3090), .Z(n3086) );
  IV U4157 ( .A(n3091), .Z(n3092) );
  XNOR U4158 ( .A(n3062), .B(n3093), .Z(n3057) );
  XNOR U4159 ( .A(n3060), .B(n3063), .Z(n3093) );
  NAND U4160 ( .A(n3094), .B(n3095), .Z(n3063) );
  NAND U4161 ( .A(n3096), .B(n3097), .Z(n3095) );
  OR U4162 ( .A(n3098), .B(n3099), .Z(n3096) );
  NANDN U4163 ( .A(n3100), .B(n3098), .Z(n3094) );
  IV U4164 ( .A(n3099), .Z(n3100) );
  NAND U4165 ( .A(n3101), .B(n3102), .Z(n3060) );
  NAND U4166 ( .A(n3103), .B(n3104), .Z(n3102) );
  NANDN U4167 ( .A(n3105), .B(n3106), .Z(n3103) );
  NANDN U4168 ( .A(n3106), .B(n3105), .Z(n3101) );
  AND U4169 ( .A(n3107), .B(n3108), .Z(n3062) );
  NAND U4170 ( .A(n3109), .B(n3110), .Z(n3108) );
  OR U4171 ( .A(n3111), .B(n3112), .Z(n3109) );
  NANDN U4172 ( .A(n3113), .B(n3111), .Z(n3107) );
  XNOR U4173 ( .A(n3088), .B(n3114), .Z(N6035) );
  XOR U4174 ( .A(n3090), .B(n3091), .Z(n3114) );
  XNOR U4175 ( .A(n3104), .B(n3115), .Z(n3091) );
  XOR U4176 ( .A(n3105), .B(n3106), .Z(n3115) );
  XOR U4177 ( .A(n3111), .B(n3116), .Z(n3106) );
  XOR U4178 ( .A(n3110), .B(n3113), .Z(n3116) );
  IV U4179 ( .A(n3112), .Z(n3113) );
  NAND U4180 ( .A(n3117), .B(n3118), .Z(n3112) );
  OR U4181 ( .A(n3119), .B(n3120), .Z(n3118) );
  OR U4182 ( .A(n3121), .B(n3122), .Z(n3117) );
  NAND U4183 ( .A(n3123), .B(n3124), .Z(n3110) );
  OR U4184 ( .A(n3125), .B(n3126), .Z(n3124) );
  OR U4185 ( .A(n3127), .B(n3128), .Z(n3123) );
  NOR U4186 ( .A(n3129), .B(n3130), .Z(n3111) );
  ANDN U4187 ( .B(n3131), .A(n3132), .Z(n3105) );
  XNOR U4188 ( .A(n3098), .B(n3133), .Z(n3104) );
  XNOR U4189 ( .A(n3097), .B(n3099), .Z(n3133) );
  NAND U4190 ( .A(n3134), .B(n3135), .Z(n3099) );
  OR U4191 ( .A(n3136), .B(n3137), .Z(n3135) );
  OR U4192 ( .A(n3138), .B(n3139), .Z(n3134) );
  NAND U4193 ( .A(n3140), .B(n3141), .Z(n3097) );
  OR U4194 ( .A(n3142), .B(n3143), .Z(n3141) );
  OR U4195 ( .A(n3144), .B(n3145), .Z(n3140) );
  ANDN U4196 ( .B(n3146), .A(n3147), .Z(n3098) );
  IV U4197 ( .A(n3148), .Z(n3146) );
  ANDN U4198 ( .B(n3149), .A(n3150), .Z(n3090) );
  XOR U4199 ( .A(n3076), .B(n3151), .Z(n3088) );
  XOR U4200 ( .A(n3077), .B(n3078), .Z(n3151) );
  XOR U4201 ( .A(n3083), .B(n3152), .Z(n3078) );
  XOR U4202 ( .A(n3082), .B(n3085), .Z(n3152) );
  IV U4203 ( .A(n3084), .Z(n3085) );
  NAND U4204 ( .A(n3153), .B(n3154), .Z(n3084) );
  OR U4205 ( .A(n3155), .B(n3156), .Z(n3154) );
  OR U4206 ( .A(n3157), .B(n3158), .Z(n3153) );
  NAND U4207 ( .A(n3159), .B(n3160), .Z(n3082) );
  OR U4208 ( .A(n3161), .B(n3162), .Z(n3160) );
  OR U4209 ( .A(n3163), .B(n3164), .Z(n3159) );
  NOR U4210 ( .A(n3165), .B(n3166), .Z(n3083) );
  ANDN U4211 ( .B(n3167), .A(n3168), .Z(n3077) );
  IV U4212 ( .A(n3169), .Z(n3167) );
  XNOR U4213 ( .A(n3070), .B(n3170), .Z(n3076) );
  XNOR U4214 ( .A(n3069), .B(n3071), .Z(n3170) );
  NAND U4215 ( .A(n3171), .B(n3172), .Z(n3071) );
  OR U4216 ( .A(n3173), .B(n3174), .Z(n3172) );
  OR U4217 ( .A(n3175), .B(n3176), .Z(n3171) );
  NAND U4218 ( .A(n3177), .B(n3178), .Z(n3069) );
  OR U4219 ( .A(n3179), .B(n3180), .Z(n3178) );
  OR U4220 ( .A(n3181), .B(n3182), .Z(n3177) );
  ANDN U4221 ( .B(n3183), .A(n3184), .Z(n3070) );
  IV U4222 ( .A(n3185), .Z(n3183) );
  XNOR U4223 ( .A(n3150), .B(n3149), .Z(N6034) );
  XOR U4224 ( .A(n3169), .B(n3168), .Z(n3149) );
  XNOR U4225 ( .A(n3184), .B(n3185), .Z(n3168) );
  XNOR U4226 ( .A(n3179), .B(n3180), .Z(n3185) );
  XNOR U4227 ( .A(n3181), .B(n3182), .Z(n3180) );
  XNOR U4228 ( .A(y[604]), .B(x[604]), .Z(n3182) );
  XNOR U4229 ( .A(y[605]), .B(x[605]), .Z(n3181) );
  XNOR U4230 ( .A(y[603]), .B(x[603]), .Z(n3179) );
  XNOR U4231 ( .A(n3173), .B(n3174), .Z(n3184) );
  XNOR U4232 ( .A(y[600]), .B(x[600]), .Z(n3174) );
  XNOR U4233 ( .A(n3175), .B(n3176), .Z(n3173) );
  XNOR U4234 ( .A(y[601]), .B(x[601]), .Z(n3176) );
  XNOR U4235 ( .A(y[602]), .B(x[602]), .Z(n3175) );
  XNOR U4236 ( .A(n3166), .B(n3165), .Z(n3169) );
  XNOR U4237 ( .A(n3161), .B(n3162), .Z(n3165) );
  XNOR U4238 ( .A(y[597]), .B(x[597]), .Z(n3162) );
  XNOR U4239 ( .A(n3163), .B(n3164), .Z(n3161) );
  XNOR U4240 ( .A(y[598]), .B(x[598]), .Z(n3164) );
  XNOR U4241 ( .A(y[599]), .B(x[599]), .Z(n3163) );
  XNOR U4242 ( .A(n3155), .B(n3156), .Z(n3166) );
  XNOR U4243 ( .A(y[594]), .B(x[594]), .Z(n3156) );
  XNOR U4244 ( .A(n3157), .B(n3158), .Z(n3155) );
  XNOR U4245 ( .A(y[595]), .B(x[595]), .Z(n3158) );
  XNOR U4246 ( .A(y[596]), .B(x[596]), .Z(n3157) );
  XOR U4247 ( .A(n3131), .B(n3132), .Z(n3150) );
  XNOR U4248 ( .A(n3147), .B(n3148), .Z(n3132) );
  XNOR U4249 ( .A(n3142), .B(n3143), .Z(n3148) );
  XNOR U4250 ( .A(n3144), .B(n3145), .Z(n3143) );
  XNOR U4251 ( .A(y[592]), .B(x[592]), .Z(n3145) );
  XNOR U4252 ( .A(y[593]), .B(x[593]), .Z(n3144) );
  XNOR U4253 ( .A(y[591]), .B(x[591]), .Z(n3142) );
  XNOR U4254 ( .A(n3136), .B(n3137), .Z(n3147) );
  XNOR U4255 ( .A(y[588]), .B(x[588]), .Z(n3137) );
  XNOR U4256 ( .A(n3138), .B(n3139), .Z(n3136) );
  XNOR U4257 ( .A(y[589]), .B(x[589]), .Z(n3139) );
  XNOR U4258 ( .A(y[590]), .B(x[590]), .Z(n3138) );
  XOR U4259 ( .A(n3130), .B(n3129), .Z(n3131) );
  XNOR U4260 ( .A(n3125), .B(n3126), .Z(n3129) );
  XNOR U4261 ( .A(y[585]), .B(x[585]), .Z(n3126) );
  XNOR U4262 ( .A(n3127), .B(n3128), .Z(n3125) );
  XNOR U4263 ( .A(y[586]), .B(x[586]), .Z(n3128) );
  XNOR U4264 ( .A(y[587]), .B(x[587]), .Z(n3127) );
  XNOR U4265 ( .A(n3119), .B(n3120), .Z(n3130) );
  XNOR U4266 ( .A(y[582]), .B(x[582]), .Z(n3120) );
  XNOR U4267 ( .A(n3121), .B(n3122), .Z(n3119) );
  XNOR U4268 ( .A(y[583]), .B(x[583]), .Z(n3122) );
  XNOR U4269 ( .A(y[584]), .B(x[584]), .Z(n3121) );
  NAND U4270 ( .A(n3186), .B(n3187), .Z(N6028) );
  NANDN U4271 ( .A(n3188), .B(n3189), .Z(n3187) );
  OR U4272 ( .A(n3190), .B(n3191), .Z(n3189) );
  NAND U4273 ( .A(n3190), .B(n3191), .Z(n3186) );
  XOR U4274 ( .A(n3190), .B(n3192), .Z(N6027) );
  XNOR U4275 ( .A(n3188), .B(n3191), .Z(n3192) );
  AND U4276 ( .A(n3193), .B(n3194), .Z(n3191) );
  NANDN U4277 ( .A(n3195), .B(n3196), .Z(n3194) );
  NANDN U4278 ( .A(n3197), .B(n3198), .Z(n3196) );
  NANDN U4279 ( .A(n3198), .B(n3197), .Z(n3193) );
  NAND U4280 ( .A(n3199), .B(n3200), .Z(n3188) );
  NANDN U4281 ( .A(n3201), .B(n3202), .Z(n3200) );
  OR U4282 ( .A(n3203), .B(n3204), .Z(n3202) );
  NAND U4283 ( .A(n3204), .B(n3203), .Z(n3199) );
  AND U4284 ( .A(n3205), .B(n3206), .Z(n3190) );
  NANDN U4285 ( .A(n3207), .B(n3208), .Z(n3206) );
  NANDN U4286 ( .A(n3209), .B(n3210), .Z(n3208) );
  NANDN U4287 ( .A(n3210), .B(n3209), .Z(n3205) );
  XOR U4288 ( .A(n3204), .B(n3211), .Z(N6026) );
  XOR U4289 ( .A(n3201), .B(n3203), .Z(n3211) );
  XNOR U4290 ( .A(n3197), .B(n3212), .Z(n3203) );
  XNOR U4291 ( .A(n3195), .B(n3198), .Z(n3212) );
  NAND U4292 ( .A(n3213), .B(n3214), .Z(n3198) );
  NAND U4293 ( .A(n3215), .B(n3216), .Z(n3214) );
  OR U4294 ( .A(n3217), .B(n3218), .Z(n3215) );
  NANDN U4295 ( .A(n3219), .B(n3217), .Z(n3213) );
  IV U4296 ( .A(n3218), .Z(n3219) );
  NAND U4297 ( .A(n3220), .B(n3221), .Z(n3195) );
  NAND U4298 ( .A(n3222), .B(n3223), .Z(n3221) );
  NANDN U4299 ( .A(n3224), .B(n3225), .Z(n3222) );
  NANDN U4300 ( .A(n3225), .B(n3224), .Z(n3220) );
  AND U4301 ( .A(n3226), .B(n3227), .Z(n3197) );
  NAND U4302 ( .A(n3228), .B(n3229), .Z(n3227) );
  OR U4303 ( .A(n3230), .B(n3231), .Z(n3228) );
  NANDN U4304 ( .A(n3232), .B(n3230), .Z(n3226) );
  NAND U4305 ( .A(n3233), .B(n3234), .Z(n3201) );
  NANDN U4306 ( .A(n3235), .B(n3236), .Z(n3234) );
  OR U4307 ( .A(n3237), .B(n3238), .Z(n3236) );
  NANDN U4308 ( .A(n3239), .B(n3237), .Z(n3233) );
  IV U4309 ( .A(n3238), .Z(n3239) );
  XNOR U4310 ( .A(n3209), .B(n3240), .Z(n3204) );
  XNOR U4311 ( .A(n3207), .B(n3210), .Z(n3240) );
  NAND U4312 ( .A(n3241), .B(n3242), .Z(n3210) );
  NAND U4313 ( .A(n3243), .B(n3244), .Z(n3242) );
  OR U4314 ( .A(n3245), .B(n3246), .Z(n3243) );
  NANDN U4315 ( .A(n3247), .B(n3245), .Z(n3241) );
  IV U4316 ( .A(n3246), .Z(n3247) );
  NAND U4317 ( .A(n3248), .B(n3249), .Z(n3207) );
  NAND U4318 ( .A(n3250), .B(n3251), .Z(n3249) );
  NANDN U4319 ( .A(n3252), .B(n3253), .Z(n3250) );
  NANDN U4320 ( .A(n3253), .B(n3252), .Z(n3248) );
  AND U4321 ( .A(n3254), .B(n3255), .Z(n3209) );
  NAND U4322 ( .A(n3256), .B(n3257), .Z(n3255) );
  OR U4323 ( .A(n3258), .B(n3259), .Z(n3256) );
  NANDN U4324 ( .A(n3260), .B(n3258), .Z(n3254) );
  XNOR U4325 ( .A(n3235), .B(n3261), .Z(N6025) );
  XOR U4326 ( .A(n3237), .B(n3238), .Z(n3261) );
  XNOR U4327 ( .A(n3251), .B(n3262), .Z(n3238) );
  XOR U4328 ( .A(n3252), .B(n3253), .Z(n3262) );
  XOR U4329 ( .A(n3258), .B(n3263), .Z(n3253) );
  XOR U4330 ( .A(n3257), .B(n3260), .Z(n3263) );
  IV U4331 ( .A(n3259), .Z(n3260) );
  NAND U4332 ( .A(n3264), .B(n3265), .Z(n3259) );
  OR U4333 ( .A(n3266), .B(n3267), .Z(n3265) );
  OR U4334 ( .A(n3268), .B(n3269), .Z(n3264) );
  NAND U4335 ( .A(n3270), .B(n3271), .Z(n3257) );
  OR U4336 ( .A(n3272), .B(n3273), .Z(n3271) );
  OR U4337 ( .A(n3274), .B(n3275), .Z(n3270) );
  NOR U4338 ( .A(n3276), .B(n3277), .Z(n3258) );
  ANDN U4339 ( .B(n3278), .A(n3279), .Z(n3252) );
  XNOR U4340 ( .A(n3245), .B(n3280), .Z(n3251) );
  XNOR U4341 ( .A(n3244), .B(n3246), .Z(n3280) );
  NAND U4342 ( .A(n3281), .B(n3282), .Z(n3246) );
  OR U4343 ( .A(n3283), .B(n3284), .Z(n3282) );
  OR U4344 ( .A(n3285), .B(n3286), .Z(n3281) );
  NAND U4345 ( .A(n3287), .B(n3288), .Z(n3244) );
  OR U4346 ( .A(n3289), .B(n3290), .Z(n3288) );
  OR U4347 ( .A(n3291), .B(n3292), .Z(n3287) );
  ANDN U4348 ( .B(n3293), .A(n3294), .Z(n3245) );
  IV U4349 ( .A(n3295), .Z(n3293) );
  ANDN U4350 ( .B(n3296), .A(n3297), .Z(n3237) );
  XOR U4351 ( .A(n3223), .B(n3298), .Z(n3235) );
  XOR U4352 ( .A(n3224), .B(n3225), .Z(n3298) );
  XOR U4353 ( .A(n3230), .B(n3299), .Z(n3225) );
  XOR U4354 ( .A(n3229), .B(n3232), .Z(n3299) );
  IV U4355 ( .A(n3231), .Z(n3232) );
  NAND U4356 ( .A(n3300), .B(n3301), .Z(n3231) );
  OR U4357 ( .A(n3302), .B(n3303), .Z(n3301) );
  OR U4358 ( .A(n3304), .B(n3305), .Z(n3300) );
  NAND U4359 ( .A(n3306), .B(n3307), .Z(n3229) );
  OR U4360 ( .A(n3308), .B(n3309), .Z(n3307) );
  OR U4361 ( .A(n3310), .B(n3311), .Z(n3306) );
  NOR U4362 ( .A(n3312), .B(n3313), .Z(n3230) );
  ANDN U4363 ( .B(n3314), .A(n3315), .Z(n3224) );
  IV U4364 ( .A(n3316), .Z(n3314) );
  XNOR U4365 ( .A(n3217), .B(n3317), .Z(n3223) );
  XNOR U4366 ( .A(n3216), .B(n3218), .Z(n3317) );
  NAND U4367 ( .A(n3318), .B(n3319), .Z(n3218) );
  OR U4368 ( .A(n3320), .B(n3321), .Z(n3319) );
  OR U4369 ( .A(n3322), .B(n3323), .Z(n3318) );
  NAND U4370 ( .A(n3324), .B(n3325), .Z(n3216) );
  OR U4371 ( .A(n3326), .B(n3327), .Z(n3325) );
  OR U4372 ( .A(n3328), .B(n3329), .Z(n3324) );
  ANDN U4373 ( .B(n3330), .A(n3331), .Z(n3217) );
  IV U4374 ( .A(n3332), .Z(n3330) );
  XNOR U4375 ( .A(n3297), .B(n3296), .Z(N6024) );
  XOR U4376 ( .A(n3316), .B(n3315), .Z(n3296) );
  XNOR U4377 ( .A(n3331), .B(n3332), .Z(n3315) );
  XNOR U4378 ( .A(n3326), .B(n3327), .Z(n3332) );
  XNOR U4379 ( .A(n3328), .B(n3329), .Z(n3327) );
  XNOR U4380 ( .A(y[580]), .B(x[580]), .Z(n3329) );
  XNOR U4381 ( .A(y[581]), .B(x[581]), .Z(n3328) );
  XNOR U4382 ( .A(y[579]), .B(x[579]), .Z(n3326) );
  XNOR U4383 ( .A(n3320), .B(n3321), .Z(n3331) );
  XNOR U4384 ( .A(y[576]), .B(x[576]), .Z(n3321) );
  XNOR U4385 ( .A(n3322), .B(n3323), .Z(n3320) );
  XNOR U4386 ( .A(y[577]), .B(x[577]), .Z(n3323) );
  XNOR U4387 ( .A(y[578]), .B(x[578]), .Z(n3322) );
  XNOR U4388 ( .A(n3313), .B(n3312), .Z(n3316) );
  XNOR U4389 ( .A(n3308), .B(n3309), .Z(n3312) );
  XNOR U4390 ( .A(y[573]), .B(x[573]), .Z(n3309) );
  XNOR U4391 ( .A(n3310), .B(n3311), .Z(n3308) );
  XNOR U4392 ( .A(y[574]), .B(x[574]), .Z(n3311) );
  XNOR U4393 ( .A(y[575]), .B(x[575]), .Z(n3310) );
  XNOR U4394 ( .A(n3302), .B(n3303), .Z(n3313) );
  XNOR U4395 ( .A(y[570]), .B(x[570]), .Z(n3303) );
  XNOR U4396 ( .A(n3304), .B(n3305), .Z(n3302) );
  XNOR U4397 ( .A(y[571]), .B(x[571]), .Z(n3305) );
  XNOR U4398 ( .A(y[572]), .B(x[572]), .Z(n3304) );
  XOR U4399 ( .A(n3278), .B(n3279), .Z(n3297) );
  XNOR U4400 ( .A(n3294), .B(n3295), .Z(n3279) );
  XNOR U4401 ( .A(n3289), .B(n3290), .Z(n3295) );
  XNOR U4402 ( .A(n3291), .B(n3292), .Z(n3290) );
  XNOR U4403 ( .A(y[568]), .B(x[568]), .Z(n3292) );
  XNOR U4404 ( .A(y[569]), .B(x[569]), .Z(n3291) );
  XNOR U4405 ( .A(y[567]), .B(x[567]), .Z(n3289) );
  XNOR U4406 ( .A(n3283), .B(n3284), .Z(n3294) );
  XNOR U4407 ( .A(y[564]), .B(x[564]), .Z(n3284) );
  XNOR U4408 ( .A(n3285), .B(n3286), .Z(n3283) );
  XNOR U4409 ( .A(y[565]), .B(x[565]), .Z(n3286) );
  XNOR U4410 ( .A(y[566]), .B(x[566]), .Z(n3285) );
  XOR U4411 ( .A(n3277), .B(n3276), .Z(n3278) );
  XNOR U4412 ( .A(n3272), .B(n3273), .Z(n3276) );
  XNOR U4413 ( .A(y[561]), .B(x[561]), .Z(n3273) );
  XNOR U4414 ( .A(n3274), .B(n3275), .Z(n3272) );
  XNOR U4415 ( .A(y[562]), .B(x[562]), .Z(n3275) );
  XNOR U4416 ( .A(y[563]), .B(x[563]), .Z(n3274) );
  XNOR U4417 ( .A(n3266), .B(n3267), .Z(n3277) );
  XNOR U4418 ( .A(y[558]), .B(x[558]), .Z(n3267) );
  XNOR U4419 ( .A(n3268), .B(n3269), .Z(n3266) );
  XNOR U4420 ( .A(y[559]), .B(x[559]), .Z(n3269) );
  XNOR U4421 ( .A(y[560]), .B(x[560]), .Z(n3268) );
  NAND U4422 ( .A(n3333), .B(n3334), .Z(N6018) );
  NANDN U4423 ( .A(n3335), .B(n3336), .Z(n3334) );
  OR U4424 ( .A(n3337), .B(n3338), .Z(n3336) );
  NAND U4425 ( .A(n3337), .B(n3338), .Z(n3333) );
  XOR U4426 ( .A(n3337), .B(n3339), .Z(N6017) );
  XNOR U4427 ( .A(n3335), .B(n3338), .Z(n3339) );
  AND U4428 ( .A(n3340), .B(n3341), .Z(n3338) );
  NANDN U4429 ( .A(n3342), .B(n3343), .Z(n3341) );
  NANDN U4430 ( .A(n3344), .B(n3345), .Z(n3343) );
  NANDN U4431 ( .A(n3345), .B(n3344), .Z(n3340) );
  NAND U4432 ( .A(n3346), .B(n3347), .Z(n3335) );
  NANDN U4433 ( .A(n3348), .B(n3349), .Z(n3347) );
  OR U4434 ( .A(n3350), .B(n3351), .Z(n3349) );
  NAND U4435 ( .A(n3351), .B(n3350), .Z(n3346) );
  AND U4436 ( .A(n3352), .B(n3353), .Z(n3337) );
  NANDN U4437 ( .A(n3354), .B(n3355), .Z(n3353) );
  NANDN U4438 ( .A(n3356), .B(n3357), .Z(n3355) );
  NANDN U4439 ( .A(n3357), .B(n3356), .Z(n3352) );
  XOR U4440 ( .A(n3351), .B(n3358), .Z(N6016) );
  XOR U4441 ( .A(n3348), .B(n3350), .Z(n3358) );
  XNOR U4442 ( .A(n3344), .B(n3359), .Z(n3350) );
  XNOR U4443 ( .A(n3342), .B(n3345), .Z(n3359) );
  NAND U4444 ( .A(n3360), .B(n3361), .Z(n3345) );
  NAND U4445 ( .A(n3362), .B(n3363), .Z(n3361) );
  OR U4446 ( .A(n3364), .B(n3365), .Z(n3362) );
  NANDN U4447 ( .A(n3366), .B(n3364), .Z(n3360) );
  IV U4448 ( .A(n3365), .Z(n3366) );
  NAND U4449 ( .A(n3367), .B(n3368), .Z(n3342) );
  NAND U4450 ( .A(n3369), .B(n3370), .Z(n3368) );
  NANDN U4451 ( .A(n3371), .B(n3372), .Z(n3369) );
  NANDN U4452 ( .A(n3372), .B(n3371), .Z(n3367) );
  AND U4453 ( .A(n3373), .B(n3374), .Z(n3344) );
  NAND U4454 ( .A(n3375), .B(n3376), .Z(n3374) );
  OR U4455 ( .A(n3377), .B(n3378), .Z(n3375) );
  NANDN U4456 ( .A(n3379), .B(n3377), .Z(n3373) );
  NAND U4457 ( .A(n3380), .B(n3381), .Z(n3348) );
  NANDN U4458 ( .A(n3382), .B(n3383), .Z(n3381) );
  OR U4459 ( .A(n3384), .B(n3385), .Z(n3383) );
  NANDN U4460 ( .A(n3386), .B(n3384), .Z(n3380) );
  IV U4461 ( .A(n3385), .Z(n3386) );
  XNOR U4462 ( .A(n3356), .B(n3387), .Z(n3351) );
  XNOR U4463 ( .A(n3354), .B(n3357), .Z(n3387) );
  NAND U4464 ( .A(n3388), .B(n3389), .Z(n3357) );
  NAND U4465 ( .A(n3390), .B(n3391), .Z(n3389) );
  OR U4466 ( .A(n3392), .B(n3393), .Z(n3390) );
  NANDN U4467 ( .A(n3394), .B(n3392), .Z(n3388) );
  IV U4468 ( .A(n3393), .Z(n3394) );
  NAND U4469 ( .A(n3395), .B(n3396), .Z(n3354) );
  NAND U4470 ( .A(n3397), .B(n3398), .Z(n3396) );
  NANDN U4471 ( .A(n3399), .B(n3400), .Z(n3397) );
  NANDN U4472 ( .A(n3400), .B(n3399), .Z(n3395) );
  AND U4473 ( .A(n3401), .B(n3402), .Z(n3356) );
  NAND U4474 ( .A(n3403), .B(n3404), .Z(n3402) );
  OR U4475 ( .A(n3405), .B(n3406), .Z(n3403) );
  NANDN U4476 ( .A(n3407), .B(n3405), .Z(n3401) );
  XNOR U4477 ( .A(n3382), .B(n3408), .Z(N6015) );
  XOR U4478 ( .A(n3384), .B(n3385), .Z(n3408) );
  XNOR U4479 ( .A(n3398), .B(n3409), .Z(n3385) );
  XOR U4480 ( .A(n3399), .B(n3400), .Z(n3409) );
  XOR U4481 ( .A(n3405), .B(n3410), .Z(n3400) );
  XOR U4482 ( .A(n3404), .B(n3407), .Z(n3410) );
  IV U4483 ( .A(n3406), .Z(n3407) );
  NAND U4484 ( .A(n3411), .B(n3412), .Z(n3406) );
  OR U4485 ( .A(n3413), .B(n3414), .Z(n3412) );
  OR U4486 ( .A(n3415), .B(n3416), .Z(n3411) );
  NAND U4487 ( .A(n3417), .B(n3418), .Z(n3404) );
  OR U4488 ( .A(n3419), .B(n3420), .Z(n3418) );
  OR U4489 ( .A(n3421), .B(n3422), .Z(n3417) );
  NOR U4490 ( .A(n3423), .B(n3424), .Z(n3405) );
  ANDN U4491 ( .B(n3425), .A(n3426), .Z(n3399) );
  XNOR U4492 ( .A(n3392), .B(n3427), .Z(n3398) );
  XNOR U4493 ( .A(n3391), .B(n3393), .Z(n3427) );
  NAND U4494 ( .A(n3428), .B(n3429), .Z(n3393) );
  OR U4495 ( .A(n3430), .B(n3431), .Z(n3429) );
  OR U4496 ( .A(n3432), .B(n3433), .Z(n3428) );
  NAND U4497 ( .A(n3434), .B(n3435), .Z(n3391) );
  OR U4498 ( .A(n3436), .B(n3437), .Z(n3435) );
  OR U4499 ( .A(n3438), .B(n3439), .Z(n3434) );
  ANDN U4500 ( .B(n3440), .A(n3441), .Z(n3392) );
  IV U4501 ( .A(n3442), .Z(n3440) );
  ANDN U4502 ( .B(n3443), .A(n3444), .Z(n3384) );
  XOR U4503 ( .A(n3370), .B(n3445), .Z(n3382) );
  XOR U4504 ( .A(n3371), .B(n3372), .Z(n3445) );
  XOR U4505 ( .A(n3377), .B(n3446), .Z(n3372) );
  XOR U4506 ( .A(n3376), .B(n3379), .Z(n3446) );
  IV U4507 ( .A(n3378), .Z(n3379) );
  NAND U4508 ( .A(n3447), .B(n3448), .Z(n3378) );
  OR U4509 ( .A(n3449), .B(n3450), .Z(n3448) );
  OR U4510 ( .A(n3451), .B(n3452), .Z(n3447) );
  NAND U4511 ( .A(n3453), .B(n3454), .Z(n3376) );
  OR U4512 ( .A(n3455), .B(n3456), .Z(n3454) );
  OR U4513 ( .A(n3457), .B(n3458), .Z(n3453) );
  NOR U4514 ( .A(n3459), .B(n3460), .Z(n3377) );
  ANDN U4515 ( .B(n3461), .A(n3462), .Z(n3371) );
  IV U4516 ( .A(n3463), .Z(n3461) );
  XNOR U4517 ( .A(n3364), .B(n3464), .Z(n3370) );
  XNOR U4518 ( .A(n3363), .B(n3365), .Z(n3464) );
  NAND U4519 ( .A(n3465), .B(n3466), .Z(n3365) );
  OR U4520 ( .A(n3467), .B(n3468), .Z(n3466) );
  OR U4521 ( .A(n3469), .B(n3470), .Z(n3465) );
  NAND U4522 ( .A(n3471), .B(n3472), .Z(n3363) );
  OR U4523 ( .A(n3473), .B(n3474), .Z(n3472) );
  OR U4524 ( .A(n3475), .B(n3476), .Z(n3471) );
  ANDN U4525 ( .B(n3477), .A(n3478), .Z(n3364) );
  IV U4526 ( .A(n3479), .Z(n3477) );
  XNOR U4527 ( .A(n3444), .B(n3443), .Z(N6014) );
  XOR U4528 ( .A(n3463), .B(n3462), .Z(n3443) );
  XNOR U4529 ( .A(n3478), .B(n3479), .Z(n3462) );
  XNOR U4530 ( .A(n3473), .B(n3474), .Z(n3479) );
  XNOR U4531 ( .A(n3475), .B(n3476), .Z(n3474) );
  XNOR U4532 ( .A(y[556]), .B(x[556]), .Z(n3476) );
  XNOR U4533 ( .A(y[557]), .B(x[557]), .Z(n3475) );
  XNOR U4534 ( .A(y[555]), .B(x[555]), .Z(n3473) );
  XNOR U4535 ( .A(n3467), .B(n3468), .Z(n3478) );
  XNOR U4536 ( .A(y[552]), .B(x[552]), .Z(n3468) );
  XNOR U4537 ( .A(n3469), .B(n3470), .Z(n3467) );
  XNOR U4538 ( .A(y[553]), .B(x[553]), .Z(n3470) );
  XNOR U4539 ( .A(y[554]), .B(x[554]), .Z(n3469) );
  XNOR U4540 ( .A(n3460), .B(n3459), .Z(n3463) );
  XNOR U4541 ( .A(n3455), .B(n3456), .Z(n3459) );
  XNOR U4542 ( .A(y[549]), .B(x[549]), .Z(n3456) );
  XNOR U4543 ( .A(n3457), .B(n3458), .Z(n3455) );
  XNOR U4544 ( .A(y[550]), .B(x[550]), .Z(n3458) );
  XNOR U4545 ( .A(y[551]), .B(x[551]), .Z(n3457) );
  XNOR U4546 ( .A(n3449), .B(n3450), .Z(n3460) );
  XNOR U4547 ( .A(y[546]), .B(x[546]), .Z(n3450) );
  XNOR U4548 ( .A(n3451), .B(n3452), .Z(n3449) );
  XNOR U4549 ( .A(y[547]), .B(x[547]), .Z(n3452) );
  XNOR U4550 ( .A(y[548]), .B(x[548]), .Z(n3451) );
  XOR U4551 ( .A(n3425), .B(n3426), .Z(n3444) );
  XNOR U4552 ( .A(n3441), .B(n3442), .Z(n3426) );
  XNOR U4553 ( .A(n3436), .B(n3437), .Z(n3442) );
  XNOR U4554 ( .A(n3438), .B(n3439), .Z(n3437) );
  XNOR U4555 ( .A(y[544]), .B(x[544]), .Z(n3439) );
  XNOR U4556 ( .A(y[545]), .B(x[545]), .Z(n3438) );
  XNOR U4557 ( .A(y[543]), .B(x[543]), .Z(n3436) );
  XNOR U4558 ( .A(n3430), .B(n3431), .Z(n3441) );
  XNOR U4559 ( .A(y[540]), .B(x[540]), .Z(n3431) );
  XNOR U4560 ( .A(n3432), .B(n3433), .Z(n3430) );
  XNOR U4561 ( .A(y[541]), .B(x[541]), .Z(n3433) );
  XNOR U4562 ( .A(y[542]), .B(x[542]), .Z(n3432) );
  XOR U4563 ( .A(n3424), .B(n3423), .Z(n3425) );
  XNOR U4564 ( .A(n3419), .B(n3420), .Z(n3423) );
  XNOR U4565 ( .A(y[537]), .B(x[537]), .Z(n3420) );
  XNOR U4566 ( .A(n3421), .B(n3422), .Z(n3419) );
  XNOR U4567 ( .A(y[538]), .B(x[538]), .Z(n3422) );
  XNOR U4568 ( .A(y[539]), .B(x[539]), .Z(n3421) );
  XNOR U4569 ( .A(n3413), .B(n3414), .Z(n3424) );
  XNOR U4570 ( .A(y[534]), .B(x[534]), .Z(n3414) );
  XNOR U4571 ( .A(n3415), .B(n3416), .Z(n3413) );
  XNOR U4572 ( .A(y[535]), .B(x[535]), .Z(n3416) );
  XNOR U4573 ( .A(y[536]), .B(x[536]), .Z(n3415) );
  NAND U4574 ( .A(n3480), .B(n3481), .Z(N6008) );
  NANDN U4575 ( .A(n3482), .B(n3483), .Z(n3481) );
  OR U4576 ( .A(n3484), .B(n3485), .Z(n3483) );
  NAND U4577 ( .A(n3484), .B(n3485), .Z(n3480) );
  XOR U4578 ( .A(n3484), .B(n3486), .Z(N6007) );
  XNOR U4579 ( .A(n3482), .B(n3485), .Z(n3486) );
  AND U4580 ( .A(n3487), .B(n3488), .Z(n3485) );
  NANDN U4581 ( .A(n3489), .B(n3490), .Z(n3488) );
  NANDN U4582 ( .A(n3491), .B(n3492), .Z(n3490) );
  NANDN U4583 ( .A(n3492), .B(n3491), .Z(n3487) );
  NAND U4584 ( .A(n3493), .B(n3494), .Z(n3482) );
  NANDN U4585 ( .A(n3495), .B(n3496), .Z(n3494) );
  OR U4586 ( .A(n3497), .B(n3498), .Z(n3496) );
  NAND U4587 ( .A(n3498), .B(n3497), .Z(n3493) );
  AND U4588 ( .A(n3499), .B(n3500), .Z(n3484) );
  NANDN U4589 ( .A(n3501), .B(n3502), .Z(n3500) );
  NANDN U4590 ( .A(n3503), .B(n3504), .Z(n3502) );
  NANDN U4591 ( .A(n3504), .B(n3503), .Z(n3499) );
  XOR U4592 ( .A(n3498), .B(n3505), .Z(N6006) );
  XOR U4593 ( .A(n3495), .B(n3497), .Z(n3505) );
  XNOR U4594 ( .A(n3491), .B(n3506), .Z(n3497) );
  XNOR U4595 ( .A(n3489), .B(n3492), .Z(n3506) );
  NAND U4596 ( .A(n3507), .B(n3508), .Z(n3492) );
  NAND U4597 ( .A(n3509), .B(n3510), .Z(n3508) );
  OR U4598 ( .A(n3511), .B(n3512), .Z(n3509) );
  NANDN U4599 ( .A(n3513), .B(n3511), .Z(n3507) );
  IV U4600 ( .A(n3512), .Z(n3513) );
  NAND U4601 ( .A(n3514), .B(n3515), .Z(n3489) );
  NAND U4602 ( .A(n3516), .B(n3517), .Z(n3515) );
  NANDN U4603 ( .A(n3518), .B(n3519), .Z(n3516) );
  NANDN U4604 ( .A(n3519), .B(n3518), .Z(n3514) );
  AND U4605 ( .A(n3520), .B(n3521), .Z(n3491) );
  NAND U4606 ( .A(n3522), .B(n3523), .Z(n3521) );
  OR U4607 ( .A(n3524), .B(n3525), .Z(n3522) );
  NANDN U4608 ( .A(n3526), .B(n3524), .Z(n3520) );
  NAND U4609 ( .A(n3527), .B(n3528), .Z(n3495) );
  NANDN U4610 ( .A(n3529), .B(n3530), .Z(n3528) );
  OR U4611 ( .A(n3531), .B(n3532), .Z(n3530) );
  NANDN U4612 ( .A(n3533), .B(n3531), .Z(n3527) );
  IV U4613 ( .A(n3532), .Z(n3533) );
  XNOR U4614 ( .A(n3503), .B(n3534), .Z(n3498) );
  XNOR U4615 ( .A(n3501), .B(n3504), .Z(n3534) );
  NAND U4616 ( .A(n3535), .B(n3536), .Z(n3504) );
  NAND U4617 ( .A(n3537), .B(n3538), .Z(n3536) );
  OR U4618 ( .A(n3539), .B(n3540), .Z(n3537) );
  NANDN U4619 ( .A(n3541), .B(n3539), .Z(n3535) );
  IV U4620 ( .A(n3540), .Z(n3541) );
  NAND U4621 ( .A(n3542), .B(n3543), .Z(n3501) );
  NAND U4622 ( .A(n3544), .B(n3545), .Z(n3543) );
  NANDN U4623 ( .A(n3546), .B(n3547), .Z(n3544) );
  NANDN U4624 ( .A(n3547), .B(n3546), .Z(n3542) );
  AND U4625 ( .A(n3548), .B(n3549), .Z(n3503) );
  NAND U4626 ( .A(n3550), .B(n3551), .Z(n3549) );
  OR U4627 ( .A(n3552), .B(n3553), .Z(n3550) );
  NANDN U4628 ( .A(n3554), .B(n3552), .Z(n3548) );
  XNOR U4629 ( .A(n3529), .B(n3555), .Z(N6005) );
  XOR U4630 ( .A(n3531), .B(n3532), .Z(n3555) );
  XNOR U4631 ( .A(n3545), .B(n3556), .Z(n3532) );
  XOR U4632 ( .A(n3546), .B(n3547), .Z(n3556) );
  XOR U4633 ( .A(n3552), .B(n3557), .Z(n3547) );
  XOR U4634 ( .A(n3551), .B(n3554), .Z(n3557) );
  IV U4635 ( .A(n3553), .Z(n3554) );
  NAND U4636 ( .A(n3558), .B(n3559), .Z(n3553) );
  OR U4637 ( .A(n3560), .B(n3561), .Z(n3559) );
  OR U4638 ( .A(n3562), .B(n3563), .Z(n3558) );
  NAND U4639 ( .A(n3564), .B(n3565), .Z(n3551) );
  OR U4640 ( .A(n3566), .B(n3567), .Z(n3565) );
  OR U4641 ( .A(n3568), .B(n3569), .Z(n3564) );
  NOR U4642 ( .A(n3570), .B(n3571), .Z(n3552) );
  ANDN U4643 ( .B(n3572), .A(n3573), .Z(n3546) );
  XNOR U4644 ( .A(n3539), .B(n3574), .Z(n3545) );
  XNOR U4645 ( .A(n3538), .B(n3540), .Z(n3574) );
  NAND U4646 ( .A(n3575), .B(n3576), .Z(n3540) );
  OR U4647 ( .A(n3577), .B(n3578), .Z(n3576) );
  OR U4648 ( .A(n3579), .B(n3580), .Z(n3575) );
  NAND U4649 ( .A(n3581), .B(n3582), .Z(n3538) );
  OR U4650 ( .A(n3583), .B(n3584), .Z(n3582) );
  OR U4651 ( .A(n3585), .B(n3586), .Z(n3581) );
  ANDN U4652 ( .B(n3587), .A(n3588), .Z(n3539) );
  IV U4653 ( .A(n3589), .Z(n3587) );
  ANDN U4654 ( .B(n3590), .A(n3591), .Z(n3531) );
  XOR U4655 ( .A(n3517), .B(n3592), .Z(n3529) );
  XOR U4656 ( .A(n3518), .B(n3519), .Z(n3592) );
  XOR U4657 ( .A(n3524), .B(n3593), .Z(n3519) );
  XOR U4658 ( .A(n3523), .B(n3526), .Z(n3593) );
  IV U4659 ( .A(n3525), .Z(n3526) );
  NAND U4660 ( .A(n3594), .B(n3595), .Z(n3525) );
  OR U4661 ( .A(n3596), .B(n3597), .Z(n3595) );
  OR U4662 ( .A(n3598), .B(n3599), .Z(n3594) );
  NAND U4663 ( .A(n3600), .B(n3601), .Z(n3523) );
  OR U4664 ( .A(n3602), .B(n3603), .Z(n3601) );
  OR U4665 ( .A(n3604), .B(n3605), .Z(n3600) );
  NOR U4666 ( .A(n3606), .B(n3607), .Z(n3524) );
  ANDN U4667 ( .B(n3608), .A(n3609), .Z(n3518) );
  IV U4668 ( .A(n3610), .Z(n3608) );
  XNOR U4669 ( .A(n3511), .B(n3611), .Z(n3517) );
  XNOR U4670 ( .A(n3510), .B(n3512), .Z(n3611) );
  NAND U4671 ( .A(n3612), .B(n3613), .Z(n3512) );
  OR U4672 ( .A(n3614), .B(n3615), .Z(n3613) );
  OR U4673 ( .A(n3616), .B(n3617), .Z(n3612) );
  NAND U4674 ( .A(n3618), .B(n3619), .Z(n3510) );
  OR U4675 ( .A(n3620), .B(n3621), .Z(n3619) );
  OR U4676 ( .A(n3622), .B(n3623), .Z(n3618) );
  ANDN U4677 ( .B(n3624), .A(n3625), .Z(n3511) );
  IV U4678 ( .A(n3626), .Z(n3624) );
  XNOR U4679 ( .A(n3591), .B(n3590), .Z(N6004) );
  XOR U4680 ( .A(n3610), .B(n3609), .Z(n3590) );
  XNOR U4681 ( .A(n3625), .B(n3626), .Z(n3609) );
  XNOR U4682 ( .A(n3620), .B(n3621), .Z(n3626) );
  XNOR U4683 ( .A(n3622), .B(n3623), .Z(n3621) );
  XNOR U4684 ( .A(y[532]), .B(x[532]), .Z(n3623) );
  XNOR U4685 ( .A(y[533]), .B(x[533]), .Z(n3622) );
  XNOR U4686 ( .A(y[531]), .B(x[531]), .Z(n3620) );
  XNOR U4687 ( .A(n3614), .B(n3615), .Z(n3625) );
  XNOR U4688 ( .A(y[528]), .B(x[528]), .Z(n3615) );
  XNOR U4689 ( .A(n3616), .B(n3617), .Z(n3614) );
  XNOR U4690 ( .A(y[529]), .B(x[529]), .Z(n3617) );
  XNOR U4691 ( .A(y[530]), .B(x[530]), .Z(n3616) );
  XNOR U4692 ( .A(n3607), .B(n3606), .Z(n3610) );
  XNOR U4693 ( .A(n3602), .B(n3603), .Z(n3606) );
  XNOR U4694 ( .A(y[525]), .B(x[525]), .Z(n3603) );
  XNOR U4695 ( .A(n3604), .B(n3605), .Z(n3602) );
  XNOR U4696 ( .A(y[526]), .B(x[526]), .Z(n3605) );
  XNOR U4697 ( .A(y[527]), .B(x[527]), .Z(n3604) );
  XNOR U4698 ( .A(n3596), .B(n3597), .Z(n3607) );
  XNOR U4699 ( .A(y[522]), .B(x[522]), .Z(n3597) );
  XNOR U4700 ( .A(n3598), .B(n3599), .Z(n3596) );
  XNOR U4701 ( .A(y[523]), .B(x[523]), .Z(n3599) );
  XNOR U4702 ( .A(y[524]), .B(x[524]), .Z(n3598) );
  XOR U4703 ( .A(n3572), .B(n3573), .Z(n3591) );
  XNOR U4704 ( .A(n3588), .B(n3589), .Z(n3573) );
  XNOR U4705 ( .A(n3583), .B(n3584), .Z(n3589) );
  XNOR U4706 ( .A(n3585), .B(n3586), .Z(n3584) );
  XNOR U4707 ( .A(y[520]), .B(x[520]), .Z(n3586) );
  XNOR U4708 ( .A(y[521]), .B(x[521]), .Z(n3585) );
  XNOR U4709 ( .A(y[519]), .B(x[519]), .Z(n3583) );
  XNOR U4710 ( .A(n3577), .B(n3578), .Z(n3588) );
  XNOR U4711 ( .A(y[516]), .B(x[516]), .Z(n3578) );
  XNOR U4712 ( .A(n3579), .B(n3580), .Z(n3577) );
  XNOR U4713 ( .A(y[517]), .B(x[517]), .Z(n3580) );
  XNOR U4714 ( .A(y[518]), .B(x[518]), .Z(n3579) );
  XOR U4715 ( .A(n3571), .B(n3570), .Z(n3572) );
  XNOR U4716 ( .A(n3566), .B(n3567), .Z(n3570) );
  XNOR U4717 ( .A(y[513]), .B(x[513]), .Z(n3567) );
  XNOR U4718 ( .A(n3568), .B(n3569), .Z(n3566) );
  XNOR U4719 ( .A(y[514]), .B(x[514]), .Z(n3569) );
  XNOR U4720 ( .A(y[515]), .B(x[515]), .Z(n3568) );
  XNOR U4721 ( .A(n3560), .B(n3561), .Z(n3571) );
  XNOR U4722 ( .A(y[510]), .B(x[510]), .Z(n3561) );
  XNOR U4723 ( .A(n3562), .B(n3563), .Z(n3560) );
  XNOR U4724 ( .A(y[511]), .B(x[511]), .Z(n3563) );
  XNOR U4725 ( .A(y[512]), .B(x[512]), .Z(n3562) );
  NAND U4726 ( .A(n3627), .B(n3628), .Z(N5998) );
  NANDN U4727 ( .A(n3629), .B(n3630), .Z(n3628) );
  OR U4728 ( .A(n3631), .B(n3632), .Z(n3630) );
  NAND U4729 ( .A(n3631), .B(n3632), .Z(n3627) );
  XOR U4730 ( .A(n3631), .B(n3633), .Z(N5997) );
  XNOR U4731 ( .A(n3629), .B(n3632), .Z(n3633) );
  AND U4732 ( .A(n3634), .B(n3635), .Z(n3632) );
  NANDN U4733 ( .A(n3636), .B(n3637), .Z(n3635) );
  NANDN U4734 ( .A(n3638), .B(n3639), .Z(n3637) );
  NANDN U4735 ( .A(n3639), .B(n3638), .Z(n3634) );
  NAND U4736 ( .A(n3640), .B(n3641), .Z(n3629) );
  NANDN U4737 ( .A(n3642), .B(n3643), .Z(n3641) );
  OR U4738 ( .A(n3644), .B(n3645), .Z(n3643) );
  NAND U4739 ( .A(n3645), .B(n3644), .Z(n3640) );
  AND U4740 ( .A(n3646), .B(n3647), .Z(n3631) );
  NANDN U4741 ( .A(n3648), .B(n3649), .Z(n3647) );
  NANDN U4742 ( .A(n3650), .B(n3651), .Z(n3649) );
  NANDN U4743 ( .A(n3651), .B(n3650), .Z(n3646) );
  XOR U4744 ( .A(n3645), .B(n3652), .Z(N5996) );
  XOR U4745 ( .A(n3642), .B(n3644), .Z(n3652) );
  XNOR U4746 ( .A(n3638), .B(n3653), .Z(n3644) );
  XNOR U4747 ( .A(n3636), .B(n3639), .Z(n3653) );
  NAND U4748 ( .A(n3654), .B(n3655), .Z(n3639) );
  NAND U4749 ( .A(n3656), .B(n3657), .Z(n3655) );
  OR U4750 ( .A(n3658), .B(n3659), .Z(n3656) );
  NANDN U4751 ( .A(n3660), .B(n3658), .Z(n3654) );
  IV U4752 ( .A(n3659), .Z(n3660) );
  NAND U4753 ( .A(n3661), .B(n3662), .Z(n3636) );
  NAND U4754 ( .A(n3663), .B(n3664), .Z(n3662) );
  NANDN U4755 ( .A(n3665), .B(n3666), .Z(n3663) );
  NANDN U4756 ( .A(n3666), .B(n3665), .Z(n3661) );
  AND U4757 ( .A(n3667), .B(n3668), .Z(n3638) );
  NAND U4758 ( .A(n3669), .B(n3670), .Z(n3668) );
  OR U4759 ( .A(n3671), .B(n3672), .Z(n3669) );
  NANDN U4760 ( .A(n3673), .B(n3671), .Z(n3667) );
  NAND U4761 ( .A(n3674), .B(n3675), .Z(n3642) );
  NANDN U4762 ( .A(n3676), .B(n3677), .Z(n3675) );
  OR U4763 ( .A(n3678), .B(n3679), .Z(n3677) );
  NANDN U4764 ( .A(n3680), .B(n3678), .Z(n3674) );
  IV U4765 ( .A(n3679), .Z(n3680) );
  XNOR U4766 ( .A(n3650), .B(n3681), .Z(n3645) );
  XNOR U4767 ( .A(n3648), .B(n3651), .Z(n3681) );
  NAND U4768 ( .A(n3682), .B(n3683), .Z(n3651) );
  NAND U4769 ( .A(n3684), .B(n3685), .Z(n3683) );
  OR U4770 ( .A(n3686), .B(n3687), .Z(n3684) );
  NANDN U4771 ( .A(n3688), .B(n3686), .Z(n3682) );
  IV U4772 ( .A(n3687), .Z(n3688) );
  NAND U4773 ( .A(n3689), .B(n3690), .Z(n3648) );
  NAND U4774 ( .A(n3691), .B(n3692), .Z(n3690) );
  NANDN U4775 ( .A(n3693), .B(n3694), .Z(n3691) );
  NANDN U4776 ( .A(n3694), .B(n3693), .Z(n3689) );
  AND U4777 ( .A(n3695), .B(n3696), .Z(n3650) );
  NAND U4778 ( .A(n3697), .B(n3698), .Z(n3696) );
  OR U4779 ( .A(n3699), .B(n3700), .Z(n3697) );
  NANDN U4780 ( .A(n3701), .B(n3699), .Z(n3695) );
  XNOR U4781 ( .A(n3676), .B(n3702), .Z(N5995) );
  XOR U4782 ( .A(n3678), .B(n3679), .Z(n3702) );
  XNOR U4783 ( .A(n3692), .B(n3703), .Z(n3679) );
  XOR U4784 ( .A(n3693), .B(n3694), .Z(n3703) );
  XOR U4785 ( .A(n3699), .B(n3704), .Z(n3694) );
  XOR U4786 ( .A(n3698), .B(n3701), .Z(n3704) );
  IV U4787 ( .A(n3700), .Z(n3701) );
  NAND U4788 ( .A(n3705), .B(n3706), .Z(n3700) );
  OR U4789 ( .A(n3707), .B(n3708), .Z(n3706) );
  OR U4790 ( .A(n3709), .B(n3710), .Z(n3705) );
  NAND U4791 ( .A(n3711), .B(n3712), .Z(n3698) );
  OR U4792 ( .A(n3713), .B(n3714), .Z(n3712) );
  OR U4793 ( .A(n3715), .B(n3716), .Z(n3711) );
  NOR U4794 ( .A(n3717), .B(n3718), .Z(n3699) );
  ANDN U4795 ( .B(n3719), .A(n3720), .Z(n3693) );
  XNOR U4796 ( .A(n3686), .B(n3721), .Z(n3692) );
  XNOR U4797 ( .A(n3685), .B(n3687), .Z(n3721) );
  NAND U4798 ( .A(n3722), .B(n3723), .Z(n3687) );
  OR U4799 ( .A(n3724), .B(n3725), .Z(n3723) );
  OR U4800 ( .A(n3726), .B(n3727), .Z(n3722) );
  NAND U4801 ( .A(n3728), .B(n3729), .Z(n3685) );
  OR U4802 ( .A(n3730), .B(n3731), .Z(n3729) );
  OR U4803 ( .A(n3732), .B(n3733), .Z(n3728) );
  ANDN U4804 ( .B(n3734), .A(n3735), .Z(n3686) );
  IV U4805 ( .A(n3736), .Z(n3734) );
  ANDN U4806 ( .B(n3737), .A(n3738), .Z(n3678) );
  XOR U4807 ( .A(n3664), .B(n3739), .Z(n3676) );
  XOR U4808 ( .A(n3665), .B(n3666), .Z(n3739) );
  XOR U4809 ( .A(n3671), .B(n3740), .Z(n3666) );
  XOR U4810 ( .A(n3670), .B(n3673), .Z(n3740) );
  IV U4811 ( .A(n3672), .Z(n3673) );
  NAND U4812 ( .A(n3741), .B(n3742), .Z(n3672) );
  OR U4813 ( .A(n3743), .B(n3744), .Z(n3742) );
  OR U4814 ( .A(n3745), .B(n3746), .Z(n3741) );
  NAND U4815 ( .A(n3747), .B(n3748), .Z(n3670) );
  OR U4816 ( .A(n3749), .B(n3750), .Z(n3748) );
  OR U4817 ( .A(n3751), .B(n3752), .Z(n3747) );
  NOR U4818 ( .A(n3753), .B(n3754), .Z(n3671) );
  ANDN U4819 ( .B(n3755), .A(n3756), .Z(n3665) );
  IV U4820 ( .A(n3757), .Z(n3755) );
  XNOR U4821 ( .A(n3658), .B(n3758), .Z(n3664) );
  XNOR U4822 ( .A(n3657), .B(n3659), .Z(n3758) );
  NAND U4823 ( .A(n3759), .B(n3760), .Z(n3659) );
  OR U4824 ( .A(n3761), .B(n3762), .Z(n3760) );
  OR U4825 ( .A(n3763), .B(n3764), .Z(n3759) );
  NAND U4826 ( .A(n3765), .B(n3766), .Z(n3657) );
  OR U4827 ( .A(n3767), .B(n3768), .Z(n3766) );
  OR U4828 ( .A(n3769), .B(n3770), .Z(n3765) );
  ANDN U4829 ( .B(n3771), .A(n3772), .Z(n3658) );
  IV U4830 ( .A(n3773), .Z(n3771) );
  XNOR U4831 ( .A(n3738), .B(n3737), .Z(N5994) );
  XOR U4832 ( .A(n3757), .B(n3756), .Z(n3737) );
  XNOR U4833 ( .A(n3772), .B(n3773), .Z(n3756) );
  XNOR U4834 ( .A(n3767), .B(n3768), .Z(n3773) );
  XNOR U4835 ( .A(n3769), .B(n3770), .Z(n3768) );
  XNOR U4836 ( .A(y[508]), .B(x[508]), .Z(n3770) );
  XNOR U4837 ( .A(y[509]), .B(x[509]), .Z(n3769) );
  XNOR U4838 ( .A(y[507]), .B(x[507]), .Z(n3767) );
  XNOR U4839 ( .A(n3761), .B(n3762), .Z(n3772) );
  XNOR U4840 ( .A(y[504]), .B(x[504]), .Z(n3762) );
  XNOR U4841 ( .A(n3763), .B(n3764), .Z(n3761) );
  XNOR U4842 ( .A(y[505]), .B(x[505]), .Z(n3764) );
  XNOR U4843 ( .A(y[506]), .B(x[506]), .Z(n3763) );
  XNOR U4844 ( .A(n3754), .B(n3753), .Z(n3757) );
  XNOR U4845 ( .A(n3749), .B(n3750), .Z(n3753) );
  XNOR U4846 ( .A(y[501]), .B(x[501]), .Z(n3750) );
  XNOR U4847 ( .A(n3751), .B(n3752), .Z(n3749) );
  XNOR U4848 ( .A(y[502]), .B(x[502]), .Z(n3752) );
  XNOR U4849 ( .A(y[503]), .B(x[503]), .Z(n3751) );
  XNOR U4850 ( .A(n3743), .B(n3744), .Z(n3754) );
  XNOR U4851 ( .A(y[498]), .B(x[498]), .Z(n3744) );
  XNOR U4852 ( .A(n3745), .B(n3746), .Z(n3743) );
  XNOR U4853 ( .A(y[499]), .B(x[499]), .Z(n3746) );
  XNOR U4854 ( .A(y[500]), .B(x[500]), .Z(n3745) );
  XOR U4855 ( .A(n3719), .B(n3720), .Z(n3738) );
  XNOR U4856 ( .A(n3735), .B(n3736), .Z(n3720) );
  XNOR U4857 ( .A(n3730), .B(n3731), .Z(n3736) );
  XNOR U4858 ( .A(n3732), .B(n3733), .Z(n3731) );
  XNOR U4859 ( .A(y[496]), .B(x[496]), .Z(n3733) );
  XNOR U4860 ( .A(y[497]), .B(x[497]), .Z(n3732) );
  XNOR U4861 ( .A(y[495]), .B(x[495]), .Z(n3730) );
  XNOR U4862 ( .A(n3724), .B(n3725), .Z(n3735) );
  XNOR U4863 ( .A(y[492]), .B(x[492]), .Z(n3725) );
  XNOR U4864 ( .A(n3726), .B(n3727), .Z(n3724) );
  XNOR U4865 ( .A(y[493]), .B(x[493]), .Z(n3727) );
  XNOR U4866 ( .A(y[494]), .B(x[494]), .Z(n3726) );
  XOR U4867 ( .A(n3718), .B(n3717), .Z(n3719) );
  XNOR U4868 ( .A(n3713), .B(n3714), .Z(n3717) );
  XNOR U4869 ( .A(y[489]), .B(x[489]), .Z(n3714) );
  XNOR U4870 ( .A(n3715), .B(n3716), .Z(n3713) );
  XNOR U4871 ( .A(y[490]), .B(x[490]), .Z(n3716) );
  XNOR U4872 ( .A(y[491]), .B(x[491]), .Z(n3715) );
  XNOR U4873 ( .A(n3707), .B(n3708), .Z(n3718) );
  XNOR U4874 ( .A(y[486]), .B(x[486]), .Z(n3708) );
  XNOR U4875 ( .A(n3709), .B(n3710), .Z(n3707) );
  XNOR U4876 ( .A(y[487]), .B(x[487]), .Z(n3710) );
  XNOR U4877 ( .A(y[488]), .B(x[488]), .Z(n3709) );
  NAND U4878 ( .A(n3774), .B(n3775), .Z(N5988) );
  NANDN U4879 ( .A(n3776), .B(n3777), .Z(n3775) );
  OR U4880 ( .A(n3778), .B(n3779), .Z(n3777) );
  NAND U4881 ( .A(n3778), .B(n3779), .Z(n3774) );
  XOR U4882 ( .A(n3778), .B(n3780), .Z(N5987) );
  XNOR U4883 ( .A(n3776), .B(n3779), .Z(n3780) );
  AND U4884 ( .A(n3781), .B(n3782), .Z(n3779) );
  NANDN U4885 ( .A(n3783), .B(n3784), .Z(n3782) );
  NANDN U4886 ( .A(n3785), .B(n3786), .Z(n3784) );
  NANDN U4887 ( .A(n3786), .B(n3785), .Z(n3781) );
  NAND U4888 ( .A(n3787), .B(n3788), .Z(n3776) );
  NANDN U4889 ( .A(n3789), .B(n3790), .Z(n3788) );
  OR U4890 ( .A(n3791), .B(n3792), .Z(n3790) );
  NAND U4891 ( .A(n3792), .B(n3791), .Z(n3787) );
  AND U4892 ( .A(n3793), .B(n3794), .Z(n3778) );
  NANDN U4893 ( .A(n3795), .B(n3796), .Z(n3794) );
  NANDN U4894 ( .A(n3797), .B(n3798), .Z(n3796) );
  NANDN U4895 ( .A(n3798), .B(n3797), .Z(n3793) );
  XOR U4896 ( .A(n3792), .B(n3799), .Z(N5986) );
  XOR U4897 ( .A(n3789), .B(n3791), .Z(n3799) );
  XNOR U4898 ( .A(n3785), .B(n3800), .Z(n3791) );
  XNOR U4899 ( .A(n3783), .B(n3786), .Z(n3800) );
  NAND U4900 ( .A(n3801), .B(n3802), .Z(n3786) );
  NAND U4901 ( .A(n3803), .B(n3804), .Z(n3802) );
  OR U4902 ( .A(n3805), .B(n3806), .Z(n3803) );
  NANDN U4903 ( .A(n3807), .B(n3805), .Z(n3801) );
  IV U4904 ( .A(n3806), .Z(n3807) );
  NAND U4905 ( .A(n3808), .B(n3809), .Z(n3783) );
  NAND U4906 ( .A(n3810), .B(n3811), .Z(n3809) );
  NANDN U4907 ( .A(n3812), .B(n3813), .Z(n3810) );
  NANDN U4908 ( .A(n3813), .B(n3812), .Z(n3808) );
  AND U4909 ( .A(n3814), .B(n3815), .Z(n3785) );
  NAND U4910 ( .A(n3816), .B(n3817), .Z(n3815) );
  OR U4911 ( .A(n3818), .B(n3819), .Z(n3816) );
  NANDN U4912 ( .A(n3820), .B(n3818), .Z(n3814) );
  NAND U4913 ( .A(n3821), .B(n3822), .Z(n3789) );
  NANDN U4914 ( .A(n3823), .B(n3824), .Z(n3822) );
  OR U4915 ( .A(n3825), .B(n3826), .Z(n3824) );
  NANDN U4916 ( .A(n3827), .B(n3825), .Z(n3821) );
  IV U4917 ( .A(n3826), .Z(n3827) );
  XNOR U4918 ( .A(n3797), .B(n3828), .Z(n3792) );
  XNOR U4919 ( .A(n3795), .B(n3798), .Z(n3828) );
  NAND U4920 ( .A(n3829), .B(n3830), .Z(n3798) );
  NAND U4921 ( .A(n3831), .B(n3832), .Z(n3830) );
  OR U4922 ( .A(n3833), .B(n3834), .Z(n3831) );
  NANDN U4923 ( .A(n3835), .B(n3833), .Z(n3829) );
  IV U4924 ( .A(n3834), .Z(n3835) );
  NAND U4925 ( .A(n3836), .B(n3837), .Z(n3795) );
  NAND U4926 ( .A(n3838), .B(n3839), .Z(n3837) );
  NANDN U4927 ( .A(n3840), .B(n3841), .Z(n3838) );
  NANDN U4928 ( .A(n3841), .B(n3840), .Z(n3836) );
  AND U4929 ( .A(n3842), .B(n3843), .Z(n3797) );
  NAND U4930 ( .A(n3844), .B(n3845), .Z(n3843) );
  OR U4931 ( .A(n3846), .B(n3847), .Z(n3844) );
  NANDN U4932 ( .A(n3848), .B(n3846), .Z(n3842) );
  XNOR U4933 ( .A(n3823), .B(n3849), .Z(N5985) );
  XOR U4934 ( .A(n3825), .B(n3826), .Z(n3849) );
  XNOR U4935 ( .A(n3839), .B(n3850), .Z(n3826) );
  XOR U4936 ( .A(n3840), .B(n3841), .Z(n3850) );
  XOR U4937 ( .A(n3846), .B(n3851), .Z(n3841) );
  XOR U4938 ( .A(n3845), .B(n3848), .Z(n3851) );
  IV U4939 ( .A(n3847), .Z(n3848) );
  NAND U4940 ( .A(n3852), .B(n3853), .Z(n3847) );
  OR U4941 ( .A(n3854), .B(n3855), .Z(n3853) );
  OR U4942 ( .A(n3856), .B(n3857), .Z(n3852) );
  NAND U4943 ( .A(n3858), .B(n3859), .Z(n3845) );
  OR U4944 ( .A(n3860), .B(n3861), .Z(n3859) );
  OR U4945 ( .A(n3862), .B(n3863), .Z(n3858) );
  NOR U4946 ( .A(n3864), .B(n3865), .Z(n3846) );
  ANDN U4947 ( .B(n3866), .A(n3867), .Z(n3840) );
  XNOR U4948 ( .A(n3833), .B(n3868), .Z(n3839) );
  XNOR U4949 ( .A(n3832), .B(n3834), .Z(n3868) );
  NAND U4950 ( .A(n3869), .B(n3870), .Z(n3834) );
  OR U4951 ( .A(n3871), .B(n3872), .Z(n3870) );
  OR U4952 ( .A(n3873), .B(n3874), .Z(n3869) );
  NAND U4953 ( .A(n3875), .B(n3876), .Z(n3832) );
  OR U4954 ( .A(n3877), .B(n3878), .Z(n3876) );
  OR U4955 ( .A(n3879), .B(n3880), .Z(n3875) );
  ANDN U4956 ( .B(n3881), .A(n3882), .Z(n3833) );
  IV U4957 ( .A(n3883), .Z(n3881) );
  ANDN U4958 ( .B(n3884), .A(n3885), .Z(n3825) );
  XOR U4959 ( .A(n3811), .B(n3886), .Z(n3823) );
  XOR U4960 ( .A(n3812), .B(n3813), .Z(n3886) );
  XOR U4961 ( .A(n3818), .B(n3887), .Z(n3813) );
  XOR U4962 ( .A(n3817), .B(n3820), .Z(n3887) );
  IV U4963 ( .A(n3819), .Z(n3820) );
  NAND U4964 ( .A(n3888), .B(n3889), .Z(n3819) );
  OR U4965 ( .A(n3890), .B(n3891), .Z(n3889) );
  OR U4966 ( .A(n3892), .B(n3893), .Z(n3888) );
  NAND U4967 ( .A(n3894), .B(n3895), .Z(n3817) );
  OR U4968 ( .A(n3896), .B(n3897), .Z(n3895) );
  OR U4969 ( .A(n3898), .B(n3899), .Z(n3894) );
  NOR U4970 ( .A(n3900), .B(n3901), .Z(n3818) );
  ANDN U4971 ( .B(n3902), .A(n3903), .Z(n3812) );
  IV U4972 ( .A(n3904), .Z(n3902) );
  XNOR U4973 ( .A(n3805), .B(n3905), .Z(n3811) );
  XNOR U4974 ( .A(n3804), .B(n3806), .Z(n3905) );
  NAND U4975 ( .A(n3906), .B(n3907), .Z(n3806) );
  OR U4976 ( .A(n3908), .B(n3909), .Z(n3907) );
  OR U4977 ( .A(n3910), .B(n3911), .Z(n3906) );
  NAND U4978 ( .A(n3912), .B(n3913), .Z(n3804) );
  OR U4979 ( .A(n3914), .B(n3915), .Z(n3913) );
  OR U4980 ( .A(n3916), .B(n3917), .Z(n3912) );
  ANDN U4981 ( .B(n3918), .A(n3919), .Z(n3805) );
  IV U4982 ( .A(n3920), .Z(n3918) );
  XNOR U4983 ( .A(n3885), .B(n3884), .Z(N5984) );
  XOR U4984 ( .A(n3904), .B(n3903), .Z(n3884) );
  XNOR U4985 ( .A(n3919), .B(n3920), .Z(n3903) );
  XNOR U4986 ( .A(n3914), .B(n3915), .Z(n3920) );
  XNOR U4987 ( .A(n3916), .B(n3917), .Z(n3915) );
  XNOR U4988 ( .A(y[484]), .B(x[484]), .Z(n3917) );
  XNOR U4989 ( .A(y[485]), .B(x[485]), .Z(n3916) );
  XNOR U4990 ( .A(y[483]), .B(x[483]), .Z(n3914) );
  XNOR U4991 ( .A(n3908), .B(n3909), .Z(n3919) );
  XNOR U4992 ( .A(y[480]), .B(x[480]), .Z(n3909) );
  XNOR U4993 ( .A(n3910), .B(n3911), .Z(n3908) );
  XNOR U4994 ( .A(y[481]), .B(x[481]), .Z(n3911) );
  XNOR U4995 ( .A(y[482]), .B(x[482]), .Z(n3910) );
  XNOR U4996 ( .A(n3901), .B(n3900), .Z(n3904) );
  XNOR U4997 ( .A(n3896), .B(n3897), .Z(n3900) );
  XNOR U4998 ( .A(y[477]), .B(x[477]), .Z(n3897) );
  XNOR U4999 ( .A(n3898), .B(n3899), .Z(n3896) );
  XNOR U5000 ( .A(y[478]), .B(x[478]), .Z(n3899) );
  XNOR U5001 ( .A(y[479]), .B(x[479]), .Z(n3898) );
  XNOR U5002 ( .A(n3890), .B(n3891), .Z(n3901) );
  XNOR U5003 ( .A(y[474]), .B(x[474]), .Z(n3891) );
  XNOR U5004 ( .A(n3892), .B(n3893), .Z(n3890) );
  XNOR U5005 ( .A(y[475]), .B(x[475]), .Z(n3893) );
  XNOR U5006 ( .A(y[476]), .B(x[476]), .Z(n3892) );
  XOR U5007 ( .A(n3866), .B(n3867), .Z(n3885) );
  XNOR U5008 ( .A(n3882), .B(n3883), .Z(n3867) );
  XNOR U5009 ( .A(n3877), .B(n3878), .Z(n3883) );
  XNOR U5010 ( .A(n3879), .B(n3880), .Z(n3878) );
  XNOR U5011 ( .A(y[472]), .B(x[472]), .Z(n3880) );
  XNOR U5012 ( .A(y[473]), .B(x[473]), .Z(n3879) );
  XNOR U5013 ( .A(y[471]), .B(x[471]), .Z(n3877) );
  XNOR U5014 ( .A(n3871), .B(n3872), .Z(n3882) );
  XNOR U5015 ( .A(y[468]), .B(x[468]), .Z(n3872) );
  XNOR U5016 ( .A(n3873), .B(n3874), .Z(n3871) );
  XNOR U5017 ( .A(y[469]), .B(x[469]), .Z(n3874) );
  XNOR U5018 ( .A(y[470]), .B(x[470]), .Z(n3873) );
  XOR U5019 ( .A(n3865), .B(n3864), .Z(n3866) );
  XNOR U5020 ( .A(n3860), .B(n3861), .Z(n3864) );
  XNOR U5021 ( .A(y[465]), .B(x[465]), .Z(n3861) );
  XNOR U5022 ( .A(n3862), .B(n3863), .Z(n3860) );
  XNOR U5023 ( .A(y[466]), .B(x[466]), .Z(n3863) );
  XNOR U5024 ( .A(y[467]), .B(x[467]), .Z(n3862) );
  XNOR U5025 ( .A(n3854), .B(n3855), .Z(n3865) );
  XNOR U5026 ( .A(y[462]), .B(x[462]), .Z(n3855) );
  XNOR U5027 ( .A(n3856), .B(n3857), .Z(n3854) );
  XNOR U5028 ( .A(y[463]), .B(x[463]), .Z(n3857) );
  XNOR U5029 ( .A(y[464]), .B(x[464]), .Z(n3856) );
  NAND U5030 ( .A(n3921), .B(n3922), .Z(N5978) );
  NANDN U5031 ( .A(n3923), .B(n3924), .Z(n3922) );
  OR U5032 ( .A(n3925), .B(n3926), .Z(n3924) );
  NAND U5033 ( .A(n3925), .B(n3926), .Z(n3921) );
  XOR U5034 ( .A(n3925), .B(n3927), .Z(N5977) );
  XNOR U5035 ( .A(n3923), .B(n3926), .Z(n3927) );
  AND U5036 ( .A(n3928), .B(n3929), .Z(n3926) );
  NANDN U5037 ( .A(n3930), .B(n3931), .Z(n3929) );
  NANDN U5038 ( .A(n3932), .B(n3933), .Z(n3931) );
  NANDN U5039 ( .A(n3933), .B(n3932), .Z(n3928) );
  NAND U5040 ( .A(n3934), .B(n3935), .Z(n3923) );
  NANDN U5041 ( .A(n3936), .B(n3937), .Z(n3935) );
  OR U5042 ( .A(n3938), .B(n3939), .Z(n3937) );
  NAND U5043 ( .A(n3939), .B(n3938), .Z(n3934) );
  AND U5044 ( .A(n3940), .B(n3941), .Z(n3925) );
  NANDN U5045 ( .A(n3942), .B(n3943), .Z(n3941) );
  NANDN U5046 ( .A(n3944), .B(n3945), .Z(n3943) );
  NANDN U5047 ( .A(n3945), .B(n3944), .Z(n3940) );
  XOR U5048 ( .A(n3939), .B(n3946), .Z(N5976) );
  XOR U5049 ( .A(n3936), .B(n3938), .Z(n3946) );
  XNOR U5050 ( .A(n3932), .B(n3947), .Z(n3938) );
  XNOR U5051 ( .A(n3930), .B(n3933), .Z(n3947) );
  NAND U5052 ( .A(n3948), .B(n3949), .Z(n3933) );
  NAND U5053 ( .A(n3950), .B(n3951), .Z(n3949) );
  OR U5054 ( .A(n3952), .B(n3953), .Z(n3950) );
  NANDN U5055 ( .A(n3954), .B(n3952), .Z(n3948) );
  IV U5056 ( .A(n3953), .Z(n3954) );
  NAND U5057 ( .A(n3955), .B(n3956), .Z(n3930) );
  NAND U5058 ( .A(n3957), .B(n3958), .Z(n3956) );
  NANDN U5059 ( .A(n3959), .B(n3960), .Z(n3957) );
  NANDN U5060 ( .A(n3960), .B(n3959), .Z(n3955) );
  AND U5061 ( .A(n3961), .B(n3962), .Z(n3932) );
  NAND U5062 ( .A(n3963), .B(n3964), .Z(n3962) );
  OR U5063 ( .A(n3965), .B(n3966), .Z(n3963) );
  NANDN U5064 ( .A(n3967), .B(n3965), .Z(n3961) );
  NAND U5065 ( .A(n3968), .B(n3969), .Z(n3936) );
  NANDN U5066 ( .A(n3970), .B(n3971), .Z(n3969) );
  OR U5067 ( .A(n3972), .B(n3973), .Z(n3971) );
  NANDN U5068 ( .A(n3974), .B(n3972), .Z(n3968) );
  IV U5069 ( .A(n3973), .Z(n3974) );
  XNOR U5070 ( .A(n3944), .B(n3975), .Z(n3939) );
  XNOR U5071 ( .A(n3942), .B(n3945), .Z(n3975) );
  NAND U5072 ( .A(n3976), .B(n3977), .Z(n3945) );
  NAND U5073 ( .A(n3978), .B(n3979), .Z(n3977) );
  OR U5074 ( .A(n3980), .B(n3981), .Z(n3978) );
  NANDN U5075 ( .A(n3982), .B(n3980), .Z(n3976) );
  IV U5076 ( .A(n3981), .Z(n3982) );
  NAND U5077 ( .A(n3983), .B(n3984), .Z(n3942) );
  NAND U5078 ( .A(n3985), .B(n3986), .Z(n3984) );
  NANDN U5079 ( .A(n3987), .B(n3988), .Z(n3985) );
  NANDN U5080 ( .A(n3988), .B(n3987), .Z(n3983) );
  AND U5081 ( .A(n3989), .B(n3990), .Z(n3944) );
  NAND U5082 ( .A(n3991), .B(n3992), .Z(n3990) );
  OR U5083 ( .A(n3993), .B(n3994), .Z(n3991) );
  NANDN U5084 ( .A(n3995), .B(n3993), .Z(n3989) );
  XNOR U5085 ( .A(n3970), .B(n3996), .Z(N5975) );
  XOR U5086 ( .A(n3972), .B(n3973), .Z(n3996) );
  XNOR U5087 ( .A(n3986), .B(n3997), .Z(n3973) );
  XOR U5088 ( .A(n3987), .B(n3988), .Z(n3997) );
  XOR U5089 ( .A(n3993), .B(n3998), .Z(n3988) );
  XOR U5090 ( .A(n3992), .B(n3995), .Z(n3998) );
  IV U5091 ( .A(n3994), .Z(n3995) );
  NAND U5092 ( .A(n3999), .B(n4000), .Z(n3994) );
  OR U5093 ( .A(n4001), .B(n4002), .Z(n4000) );
  OR U5094 ( .A(n4003), .B(n4004), .Z(n3999) );
  NAND U5095 ( .A(n4005), .B(n4006), .Z(n3992) );
  OR U5096 ( .A(n4007), .B(n4008), .Z(n4006) );
  OR U5097 ( .A(n4009), .B(n4010), .Z(n4005) );
  NOR U5098 ( .A(n4011), .B(n4012), .Z(n3993) );
  ANDN U5099 ( .B(n4013), .A(n4014), .Z(n3987) );
  XNOR U5100 ( .A(n3980), .B(n4015), .Z(n3986) );
  XNOR U5101 ( .A(n3979), .B(n3981), .Z(n4015) );
  NAND U5102 ( .A(n4016), .B(n4017), .Z(n3981) );
  OR U5103 ( .A(n4018), .B(n4019), .Z(n4017) );
  OR U5104 ( .A(n4020), .B(n4021), .Z(n4016) );
  NAND U5105 ( .A(n4022), .B(n4023), .Z(n3979) );
  OR U5106 ( .A(n4024), .B(n4025), .Z(n4023) );
  OR U5107 ( .A(n4026), .B(n4027), .Z(n4022) );
  ANDN U5108 ( .B(n4028), .A(n4029), .Z(n3980) );
  IV U5109 ( .A(n4030), .Z(n4028) );
  ANDN U5110 ( .B(n4031), .A(n4032), .Z(n3972) );
  XOR U5111 ( .A(n3958), .B(n4033), .Z(n3970) );
  XOR U5112 ( .A(n3959), .B(n3960), .Z(n4033) );
  XOR U5113 ( .A(n3965), .B(n4034), .Z(n3960) );
  XOR U5114 ( .A(n3964), .B(n3967), .Z(n4034) );
  IV U5115 ( .A(n3966), .Z(n3967) );
  NAND U5116 ( .A(n4035), .B(n4036), .Z(n3966) );
  OR U5117 ( .A(n4037), .B(n4038), .Z(n4036) );
  OR U5118 ( .A(n4039), .B(n4040), .Z(n4035) );
  NAND U5119 ( .A(n4041), .B(n4042), .Z(n3964) );
  OR U5120 ( .A(n4043), .B(n4044), .Z(n4042) );
  OR U5121 ( .A(n4045), .B(n4046), .Z(n4041) );
  NOR U5122 ( .A(n4047), .B(n4048), .Z(n3965) );
  ANDN U5123 ( .B(n4049), .A(n4050), .Z(n3959) );
  IV U5124 ( .A(n4051), .Z(n4049) );
  XNOR U5125 ( .A(n3952), .B(n4052), .Z(n3958) );
  XNOR U5126 ( .A(n3951), .B(n3953), .Z(n4052) );
  NAND U5127 ( .A(n4053), .B(n4054), .Z(n3953) );
  OR U5128 ( .A(n4055), .B(n4056), .Z(n4054) );
  OR U5129 ( .A(n4057), .B(n4058), .Z(n4053) );
  NAND U5130 ( .A(n4059), .B(n4060), .Z(n3951) );
  OR U5131 ( .A(n4061), .B(n4062), .Z(n4060) );
  OR U5132 ( .A(n4063), .B(n4064), .Z(n4059) );
  ANDN U5133 ( .B(n4065), .A(n4066), .Z(n3952) );
  IV U5134 ( .A(n4067), .Z(n4065) );
  XNOR U5135 ( .A(n4032), .B(n4031), .Z(N5974) );
  XOR U5136 ( .A(n4051), .B(n4050), .Z(n4031) );
  XNOR U5137 ( .A(n4066), .B(n4067), .Z(n4050) );
  XNOR U5138 ( .A(n4061), .B(n4062), .Z(n4067) );
  XNOR U5139 ( .A(n4063), .B(n4064), .Z(n4062) );
  XNOR U5140 ( .A(y[460]), .B(x[460]), .Z(n4064) );
  XNOR U5141 ( .A(y[461]), .B(x[461]), .Z(n4063) );
  XNOR U5142 ( .A(y[459]), .B(x[459]), .Z(n4061) );
  XNOR U5143 ( .A(n4055), .B(n4056), .Z(n4066) );
  XNOR U5144 ( .A(y[456]), .B(x[456]), .Z(n4056) );
  XNOR U5145 ( .A(n4057), .B(n4058), .Z(n4055) );
  XNOR U5146 ( .A(y[457]), .B(x[457]), .Z(n4058) );
  XNOR U5147 ( .A(y[458]), .B(x[458]), .Z(n4057) );
  XNOR U5148 ( .A(n4048), .B(n4047), .Z(n4051) );
  XNOR U5149 ( .A(n4043), .B(n4044), .Z(n4047) );
  XNOR U5150 ( .A(y[453]), .B(x[453]), .Z(n4044) );
  XNOR U5151 ( .A(n4045), .B(n4046), .Z(n4043) );
  XNOR U5152 ( .A(y[454]), .B(x[454]), .Z(n4046) );
  XNOR U5153 ( .A(y[455]), .B(x[455]), .Z(n4045) );
  XNOR U5154 ( .A(n4037), .B(n4038), .Z(n4048) );
  XNOR U5155 ( .A(y[450]), .B(x[450]), .Z(n4038) );
  XNOR U5156 ( .A(n4039), .B(n4040), .Z(n4037) );
  XNOR U5157 ( .A(y[451]), .B(x[451]), .Z(n4040) );
  XNOR U5158 ( .A(y[452]), .B(x[452]), .Z(n4039) );
  XOR U5159 ( .A(n4013), .B(n4014), .Z(n4032) );
  XNOR U5160 ( .A(n4029), .B(n4030), .Z(n4014) );
  XNOR U5161 ( .A(n4024), .B(n4025), .Z(n4030) );
  XNOR U5162 ( .A(n4026), .B(n4027), .Z(n4025) );
  XNOR U5163 ( .A(y[448]), .B(x[448]), .Z(n4027) );
  XNOR U5164 ( .A(y[449]), .B(x[449]), .Z(n4026) );
  XNOR U5165 ( .A(y[447]), .B(x[447]), .Z(n4024) );
  XNOR U5166 ( .A(n4018), .B(n4019), .Z(n4029) );
  XNOR U5167 ( .A(y[444]), .B(x[444]), .Z(n4019) );
  XNOR U5168 ( .A(n4020), .B(n4021), .Z(n4018) );
  XNOR U5169 ( .A(y[445]), .B(x[445]), .Z(n4021) );
  XNOR U5170 ( .A(y[446]), .B(x[446]), .Z(n4020) );
  XOR U5171 ( .A(n4012), .B(n4011), .Z(n4013) );
  XNOR U5172 ( .A(n4007), .B(n4008), .Z(n4011) );
  XNOR U5173 ( .A(y[441]), .B(x[441]), .Z(n4008) );
  XNOR U5174 ( .A(n4009), .B(n4010), .Z(n4007) );
  XNOR U5175 ( .A(y[442]), .B(x[442]), .Z(n4010) );
  XNOR U5176 ( .A(y[443]), .B(x[443]), .Z(n4009) );
  XNOR U5177 ( .A(n4001), .B(n4002), .Z(n4012) );
  XNOR U5178 ( .A(y[438]), .B(x[438]), .Z(n4002) );
  XNOR U5179 ( .A(n4003), .B(n4004), .Z(n4001) );
  XNOR U5180 ( .A(y[439]), .B(x[439]), .Z(n4004) );
  XNOR U5181 ( .A(y[440]), .B(x[440]), .Z(n4003) );
  NAND U5182 ( .A(n4068), .B(n4069), .Z(N5968) );
  NANDN U5183 ( .A(n4070), .B(n4071), .Z(n4069) );
  OR U5184 ( .A(n4072), .B(n4073), .Z(n4071) );
  NAND U5185 ( .A(n4072), .B(n4073), .Z(n4068) );
  XOR U5186 ( .A(n4072), .B(n4074), .Z(N5967) );
  XNOR U5187 ( .A(n4070), .B(n4073), .Z(n4074) );
  AND U5188 ( .A(n4075), .B(n4076), .Z(n4073) );
  NANDN U5189 ( .A(n4077), .B(n4078), .Z(n4076) );
  NANDN U5190 ( .A(n4079), .B(n4080), .Z(n4078) );
  NANDN U5191 ( .A(n4080), .B(n4079), .Z(n4075) );
  NAND U5192 ( .A(n4081), .B(n4082), .Z(n4070) );
  NANDN U5193 ( .A(n4083), .B(n4084), .Z(n4082) );
  OR U5194 ( .A(n4085), .B(n4086), .Z(n4084) );
  NAND U5195 ( .A(n4086), .B(n4085), .Z(n4081) );
  AND U5196 ( .A(n4087), .B(n4088), .Z(n4072) );
  NANDN U5197 ( .A(n4089), .B(n4090), .Z(n4088) );
  NANDN U5198 ( .A(n4091), .B(n4092), .Z(n4090) );
  NANDN U5199 ( .A(n4092), .B(n4091), .Z(n4087) );
  XOR U5200 ( .A(n4086), .B(n4093), .Z(N5966) );
  XOR U5201 ( .A(n4083), .B(n4085), .Z(n4093) );
  XNOR U5202 ( .A(n4079), .B(n4094), .Z(n4085) );
  XNOR U5203 ( .A(n4077), .B(n4080), .Z(n4094) );
  NAND U5204 ( .A(n4095), .B(n4096), .Z(n4080) );
  NAND U5205 ( .A(n4097), .B(n4098), .Z(n4096) );
  OR U5206 ( .A(n4099), .B(n4100), .Z(n4097) );
  NANDN U5207 ( .A(n4101), .B(n4099), .Z(n4095) );
  IV U5208 ( .A(n4100), .Z(n4101) );
  NAND U5209 ( .A(n4102), .B(n4103), .Z(n4077) );
  NAND U5210 ( .A(n4104), .B(n4105), .Z(n4103) );
  NANDN U5211 ( .A(n4106), .B(n4107), .Z(n4104) );
  NANDN U5212 ( .A(n4107), .B(n4106), .Z(n4102) );
  AND U5213 ( .A(n4108), .B(n4109), .Z(n4079) );
  NAND U5214 ( .A(n4110), .B(n4111), .Z(n4109) );
  OR U5215 ( .A(n4112), .B(n4113), .Z(n4110) );
  NANDN U5216 ( .A(n4114), .B(n4112), .Z(n4108) );
  NAND U5217 ( .A(n4115), .B(n4116), .Z(n4083) );
  NANDN U5218 ( .A(n4117), .B(n4118), .Z(n4116) );
  OR U5219 ( .A(n4119), .B(n4120), .Z(n4118) );
  NANDN U5220 ( .A(n4121), .B(n4119), .Z(n4115) );
  IV U5221 ( .A(n4120), .Z(n4121) );
  XNOR U5222 ( .A(n4091), .B(n4122), .Z(n4086) );
  XNOR U5223 ( .A(n4089), .B(n4092), .Z(n4122) );
  NAND U5224 ( .A(n4123), .B(n4124), .Z(n4092) );
  NAND U5225 ( .A(n4125), .B(n4126), .Z(n4124) );
  OR U5226 ( .A(n4127), .B(n4128), .Z(n4125) );
  NANDN U5227 ( .A(n4129), .B(n4127), .Z(n4123) );
  IV U5228 ( .A(n4128), .Z(n4129) );
  NAND U5229 ( .A(n4130), .B(n4131), .Z(n4089) );
  NAND U5230 ( .A(n4132), .B(n4133), .Z(n4131) );
  NANDN U5231 ( .A(n4134), .B(n4135), .Z(n4132) );
  NANDN U5232 ( .A(n4135), .B(n4134), .Z(n4130) );
  AND U5233 ( .A(n4136), .B(n4137), .Z(n4091) );
  NAND U5234 ( .A(n4138), .B(n4139), .Z(n4137) );
  OR U5235 ( .A(n4140), .B(n4141), .Z(n4138) );
  NANDN U5236 ( .A(n4142), .B(n4140), .Z(n4136) );
  XNOR U5237 ( .A(n4117), .B(n4143), .Z(N5965) );
  XOR U5238 ( .A(n4119), .B(n4120), .Z(n4143) );
  XNOR U5239 ( .A(n4133), .B(n4144), .Z(n4120) );
  XOR U5240 ( .A(n4134), .B(n4135), .Z(n4144) );
  XOR U5241 ( .A(n4140), .B(n4145), .Z(n4135) );
  XOR U5242 ( .A(n4139), .B(n4142), .Z(n4145) );
  IV U5243 ( .A(n4141), .Z(n4142) );
  NAND U5244 ( .A(n4146), .B(n4147), .Z(n4141) );
  OR U5245 ( .A(n4148), .B(n4149), .Z(n4147) );
  OR U5246 ( .A(n4150), .B(n4151), .Z(n4146) );
  NAND U5247 ( .A(n4152), .B(n4153), .Z(n4139) );
  OR U5248 ( .A(n4154), .B(n4155), .Z(n4153) );
  OR U5249 ( .A(n4156), .B(n4157), .Z(n4152) );
  NOR U5250 ( .A(n4158), .B(n4159), .Z(n4140) );
  ANDN U5251 ( .B(n4160), .A(n4161), .Z(n4134) );
  XNOR U5252 ( .A(n4127), .B(n4162), .Z(n4133) );
  XNOR U5253 ( .A(n4126), .B(n4128), .Z(n4162) );
  NAND U5254 ( .A(n4163), .B(n4164), .Z(n4128) );
  OR U5255 ( .A(n4165), .B(n4166), .Z(n4164) );
  OR U5256 ( .A(n4167), .B(n4168), .Z(n4163) );
  NAND U5257 ( .A(n4169), .B(n4170), .Z(n4126) );
  OR U5258 ( .A(n4171), .B(n4172), .Z(n4170) );
  OR U5259 ( .A(n4173), .B(n4174), .Z(n4169) );
  ANDN U5260 ( .B(n4175), .A(n4176), .Z(n4127) );
  IV U5261 ( .A(n4177), .Z(n4175) );
  ANDN U5262 ( .B(n4178), .A(n4179), .Z(n4119) );
  XOR U5263 ( .A(n4105), .B(n4180), .Z(n4117) );
  XOR U5264 ( .A(n4106), .B(n4107), .Z(n4180) );
  XOR U5265 ( .A(n4112), .B(n4181), .Z(n4107) );
  XOR U5266 ( .A(n4111), .B(n4114), .Z(n4181) );
  IV U5267 ( .A(n4113), .Z(n4114) );
  NAND U5268 ( .A(n4182), .B(n4183), .Z(n4113) );
  OR U5269 ( .A(n4184), .B(n4185), .Z(n4183) );
  OR U5270 ( .A(n4186), .B(n4187), .Z(n4182) );
  NAND U5271 ( .A(n4188), .B(n4189), .Z(n4111) );
  OR U5272 ( .A(n4190), .B(n4191), .Z(n4189) );
  OR U5273 ( .A(n4192), .B(n4193), .Z(n4188) );
  NOR U5274 ( .A(n4194), .B(n4195), .Z(n4112) );
  ANDN U5275 ( .B(n4196), .A(n4197), .Z(n4106) );
  IV U5276 ( .A(n4198), .Z(n4196) );
  XNOR U5277 ( .A(n4099), .B(n4199), .Z(n4105) );
  XNOR U5278 ( .A(n4098), .B(n4100), .Z(n4199) );
  NAND U5279 ( .A(n4200), .B(n4201), .Z(n4100) );
  OR U5280 ( .A(n4202), .B(n4203), .Z(n4201) );
  OR U5281 ( .A(n4204), .B(n4205), .Z(n4200) );
  NAND U5282 ( .A(n4206), .B(n4207), .Z(n4098) );
  OR U5283 ( .A(n4208), .B(n4209), .Z(n4207) );
  OR U5284 ( .A(n4210), .B(n4211), .Z(n4206) );
  ANDN U5285 ( .B(n4212), .A(n4213), .Z(n4099) );
  IV U5286 ( .A(n4214), .Z(n4212) );
  XNOR U5287 ( .A(n4179), .B(n4178), .Z(N5964) );
  XOR U5288 ( .A(n4198), .B(n4197), .Z(n4178) );
  XNOR U5289 ( .A(n4213), .B(n4214), .Z(n4197) );
  XNOR U5290 ( .A(n4208), .B(n4209), .Z(n4214) );
  XNOR U5291 ( .A(n4210), .B(n4211), .Z(n4209) );
  XNOR U5292 ( .A(y[436]), .B(x[436]), .Z(n4211) );
  XNOR U5293 ( .A(y[437]), .B(x[437]), .Z(n4210) );
  XNOR U5294 ( .A(y[435]), .B(x[435]), .Z(n4208) );
  XNOR U5295 ( .A(n4202), .B(n4203), .Z(n4213) );
  XNOR U5296 ( .A(y[432]), .B(x[432]), .Z(n4203) );
  XNOR U5297 ( .A(n4204), .B(n4205), .Z(n4202) );
  XNOR U5298 ( .A(y[433]), .B(x[433]), .Z(n4205) );
  XNOR U5299 ( .A(y[434]), .B(x[434]), .Z(n4204) );
  XNOR U5300 ( .A(n4195), .B(n4194), .Z(n4198) );
  XNOR U5301 ( .A(n4190), .B(n4191), .Z(n4194) );
  XNOR U5302 ( .A(y[429]), .B(x[429]), .Z(n4191) );
  XNOR U5303 ( .A(n4192), .B(n4193), .Z(n4190) );
  XNOR U5304 ( .A(y[430]), .B(x[430]), .Z(n4193) );
  XNOR U5305 ( .A(y[431]), .B(x[431]), .Z(n4192) );
  XNOR U5306 ( .A(n4184), .B(n4185), .Z(n4195) );
  XNOR U5307 ( .A(y[426]), .B(x[426]), .Z(n4185) );
  XNOR U5308 ( .A(n4186), .B(n4187), .Z(n4184) );
  XNOR U5309 ( .A(y[427]), .B(x[427]), .Z(n4187) );
  XNOR U5310 ( .A(y[428]), .B(x[428]), .Z(n4186) );
  XOR U5311 ( .A(n4160), .B(n4161), .Z(n4179) );
  XNOR U5312 ( .A(n4176), .B(n4177), .Z(n4161) );
  XNOR U5313 ( .A(n4171), .B(n4172), .Z(n4177) );
  XNOR U5314 ( .A(n4173), .B(n4174), .Z(n4172) );
  XNOR U5315 ( .A(y[424]), .B(x[424]), .Z(n4174) );
  XNOR U5316 ( .A(y[425]), .B(x[425]), .Z(n4173) );
  XNOR U5317 ( .A(y[423]), .B(x[423]), .Z(n4171) );
  XNOR U5318 ( .A(n4165), .B(n4166), .Z(n4176) );
  XNOR U5319 ( .A(y[420]), .B(x[420]), .Z(n4166) );
  XNOR U5320 ( .A(n4167), .B(n4168), .Z(n4165) );
  XNOR U5321 ( .A(y[421]), .B(x[421]), .Z(n4168) );
  XNOR U5322 ( .A(y[422]), .B(x[422]), .Z(n4167) );
  XOR U5323 ( .A(n4159), .B(n4158), .Z(n4160) );
  XNOR U5324 ( .A(n4154), .B(n4155), .Z(n4158) );
  XNOR U5325 ( .A(y[417]), .B(x[417]), .Z(n4155) );
  XNOR U5326 ( .A(n4156), .B(n4157), .Z(n4154) );
  XNOR U5327 ( .A(y[418]), .B(x[418]), .Z(n4157) );
  XNOR U5328 ( .A(y[419]), .B(x[419]), .Z(n4156) );
  XNOR U5329 ( .A(n4148), .B(n4149), .Z(n4159) );
  XNOR U5330 ( .A(y[414]), .B(x[414]), .Z(n4149) );
  XNOR U5331 ( .A(n4150), .B(n4151), .Z(n4148) );
  XNOR U5332 ( .A(y[415]), .B(x[415]), .Z(n4151) );
  XNOR U5333 ( .A(y[416]), .B(x[416]), .Z(n4150) );
  NAND U5334 ( .A(n4215), .B(n4216), .Z(N5958) );
  NANDN U5335 ( .A(n4217), .B(n4218), .Z(n4216) );
  OR U5336 ( .A(n4219), .B(n4220), .Z(n4218) );
  NAND U5337 ( .A(n4219), .B(n4220), .Z(n4215) );
  XOR U5338 ( .A(n4219), .B(n4221), .Z(N5957) );
  XNOR U5339 ( .A(n4217), .B(n4220), .Z(n4221) );
  AND U5340 ( .A(n4222), .B(n4223), .Z(n4220) );
  NANDN U5341 ( .A(n4224), .B(n4225), .Z(n4223) );
  NANDN U5342 ( .A(n4226), .B(n4227), .Z(n4225) );
  NANDN U5343 ( .A(n4227), .B(n4226), .Z(n4222) );
  NAND U5344 ( .A(n4228), .B(n4229), .Z(n4217) );
  NANDN U5345 ( .A(n4230), .B(n4231), .Z(n4229) );
  OR U5346 ( .A(n4232), .B(n4233), .Z(n4231) );
  NAND U5347 ( .A(n4233), .B(n4232), .Z(n4228) );
  AND U5348 ( .A(n4234), .B(n4235), .Z(n4219) );
  NANDN U5349 ( .A(n4236), .B(n4237), .Z(n4235) );
  NANDN U5350 ( .A(n4238), .B(n4239), .Z(n4237) );
  NANDN U5351 ( .A(n4239), .B(n4238), .Z(n4234) );
  XOR U5352 ( .A(n4233), .B(n4240), .Z(N5956) );
  XOR U5353 ( .A(n4230), .B(n4232), .Z(n4240) );
  XNOR U5354 ( .A(n4226), .B(n4241), .Z(n4232) );
  XNOR U5355 ( .A(n4224), .B(n4227), .Z(n4241) );
  NAND U5356 ( .A(n4242), .B(n4243), .Z(n4227) );
  NAND U5357 ( .A(n4244), .B(n4245), .Z(n4243) );
  OR U5358 ( .A(n4246), .B(n4247), .Z(n4244) );
  NANDN U5359 ( .A(n4248), .B(n4246), .Z(n4242) );
  IV U5360 ( .A(n4247), .Z(n4248) );
  NAND U5361 ( .A(n4249), .B(n4250), .Z(n4224) );
  NAND U5362 ( .A(n4251), .B(n4252), .Z(n4250) );
  NANDN U5363 ( .A(n4253), .B(n4254), .Z(n4251) );
  NANDN U5364 ( .A(n4254), .B(n4253), .Z(n4249) );
  AND U5365 ( .A(n4255), .B(n4256), .Z(n4226) );
  NAND U5366 ( .A(n4257), .B(n4258), .Z(n4256) );
  OR U5367 ( .A(n4259), .B(n4260), .Z(n4257) );
  NANDN U5368 ( .A(n4261), .B(n4259), .Z(n4255) );
  NAND U5369 ( .A(n4262), .B(n4263), .Z(n4230) );
  NANDN U5370 ( .A(n4264), .B(n4265), .Z(n4263) );
  OR U5371 ( .A(n4266), .B(n4267), .Z(n4265) );
  NANDN U5372 ( .A(n4268), .B(n4266), .Z(n4262) );
  IV U5373 ( .A(n4267), .Z(n4268) );
  XNOR U5374 ( .A(n4238), .B(n4269), .Z(n4233) );
  XNOR U5375 ( .A(n4236), .B(n4239), .Z(n4269) );
  NAND U5376 ( .A(n4270), .B(n4271), .Z(n4239) );
  NAND U5377 ( .A(n4272), .B(n4273), .Z(n4271) );
  OR U5378 ( .A(n4274), .B(n4275), .Z(n4272) );
  NANDN U5379 ( .A(n4276), .B(n4274), .Z(n4270) );
  IV U5380 ( .A(n4275), .Z(n4276) );
  NAND U5381 ( .A(n4277), .B(n4278), .Z(n4236) );
  NAND U5382 ( .A(n4279), .B(n4280), .Z(n4278) );
  NANDN U5383 ( .A(n4281), .B(n4282), .Z(n4279) );
  NANDN U5384 ( .A(n4282), .B(n4281), .Z(n4277) );
  AND U5385 ( .A(n4283), .B(n4284), .Z(n4238) );
  NAND U5386 ( .A(n4285), .B(n4286), .Z(n4284) );
  OR U5387 ( .A(n4287), .B(n4288), .Z(n4285) );
  NANDN U5388 ( .A(n4289), .B(n4287), .Z(n4283) );
  XNOR U5389 ( .A(n4264), .B(n4290), .Z(N5955) );
  XOR U5390 ( .A(n4266), .B(n4267), .Z(n4290) );
  XNOR U5391 ( .A(n4280), .B(n4291), .Z(n4267) );
  XOR U5392 ( .A(n4281), .B(n4282), .Z(n4291) );
  XOR U5393 ( .A(n4287), .B(n4292), .Z(n4282) );
  XOR U5394 ( .A(n4286), .B(n4289), .Z(n4292) );
  IV U5395 ( .A(n4288), .Z(n4289) );
  NAND U5396 ( .A(n4293), .B(n4294), .Z(n4288) );
  OR U5397 ( .A(n4295), .B(n4296), .Z(n4294) );
  OR U5398 ( .A(n4297), .B(n4298), .Z(n4293) );
  NAND U5399 ( .A(n4299), .B(n4300), .Z(n4286) );
  OR U5400 ( .A(n4301), .B(n4302), .Z(n4300) );
  OR U5401 ( .A(n4303), .B(n4304), .Z(n4299) );
  NOR U5402 ( .A(n4305), .B(n4306), .Z(n4287) );
  ANDN U5403 ( .B(n4307), .A(n4308), .Z(n4281) );
  XNOR U5404 ( .A(n4274), .B(n4309), .Z(n4280) );
  XNOR U5405 ( .A(n4273), .B(n4275), .Z(n4309) );
  NAND U5406 ( .A(n4310), .B(n4311), .Z(n4275) );
  OR U5407 ( .A(n4312), .B(n4313), .Z(n4311) );
  OR U5408 ( .A(n4314), .B(n4315), .Z(n4310) );
  NAND U5409 ( .A(n4316), .B(n4317), .Z(n4273) );
  OR U5410 ( .A(n4318), .B(n4319), .Z(n4317) );
  OR U5411 ( .A(n4320), .B(n4321), .Z(n4316) );
  ANDN U5412 ( .B(n4322), .A(n4323), .Z(n4274) );
  IV U5413 ( .A(n4324), .Z(n4322) );
  ANDN U5414 ( .B(n4325), .A(n4326), .Z(n4266) );
  XOR U5415 ( .A(n4252), .B(n4327), .Z(n4264) );
  XOR U5416 ( .A(n4253), .B(n4254), .Z(n4327) );
  XOR U5417 ( .A(n4259), .B(n4328), .Z(n4254) );
  XOR U5418 ( .A(n4258), .B(n4261), .Z(n4328) );
  IV U5419 ( .A(n4260), .Z(n4261) );
  NAND U5420 ( .A(n4329), .B(n4330), .Z(n4260) );
  OR U5421 ( .A(n4331), .B(n4332), .Z(n4330) );
  OR U5422 ( .A(n4333), .B(n4334), .Z(n4329) );
  NAND U5423 ( .A(n4335), .B(n4336), .Z(n4258) );
  OR U5424 ( .A(n4337), .B(n4338), .Z(n4336) );
  OR U5425 ( .A(n4339), .B(n4340), .Z(n4335) );
  NOR U5426 ( .A(n4341), .B(n4342), .Z(n4259) );
  ANDN U5427 ( .B(n4343), .A(n4344), .Z(n4253) );
  IV U5428 ( .A(n4345), .Z(n4343) );
  XNOR U5429 ( .A(n4246), .B(n4346), .Z(n4252) );
  XNOR U5430 ( .A(n4245), .B(n4247), .Z(n4346) );
  NAND U5431 ( .A(n4347), .B(n4348), .Z(n4247) );
  OR U5432 ( .A(n4349), .B(n4350), .Z(n4348) );
  OR U5433 ( .A(n4351), .B(n4352), .Z(n4347) );
  NAND U5434 ( .A(n4353), .B(n4354), .Z(n4245) );
  OR U5435 ( .A(n4355), .B(n4356), .Z(n4354) );
  OR U5436 ( .A(n4357), .B(n4358), .Z(n4353) );
  ANDN U5437 ( .B(n4359), .A(n4360), .Z(n4246) );
  IV U5438 ( .A(n4361), .Z(n4359) );
  XNOR U5439 ( .A(n4326), .B(n4325), .Z(N5954) );
  XOR U5440 ( .A(n4345), .B(n4344), .Z(n4325) );
  XNOR U5441 ( .A(n4360), .B(n4361), .Z(n4344) );
  XNOR U5442 ( .A(n4355), .B(n4356), .Z(n4361) );
  XNOR U5443 ( .A(n4357), .B(n4358), .Z(n4356) );
  XNOR U5444 ( .A(y[412]), .B(x[412]), .Z(n4358) );
  XNOR U5445 ( .A(y[413]), .B(x[413]), .Z(n4357) );
  XNOR U5446 ( .A(y[411]), .B(x[411]), .Z(n4355) );
  XNOR U5447 ( .A(n4349), .B(n4350), .Z(n4360) );
  XNOR U5448 ( .A(y[408]), .B(x[408]), .Z(n4350) );
  XNOR U5449 ( .A(n4351), .B(n4352), .Z(n4349) );
  XNOR U5450 ( .A(y[409]), .B(x[409]), .Z(n4352) );
  XNOR U5451 ( .A(y[410]), .B(x[410]), .Z(n4351) );
  XNOR U5452 ( .A(n4342), .B(n4341), .Z(n4345) );
  XNOR U5453 ( .A(n4337), .B(n4338), .Z(n4341) );
  XNOR U5454 ( .A(y[405]), .B(x[405]), .Z(n4338) );
  XNOR U5455 ( .A(n4339), .B(n4340), .Z(n4337) );
  XNOR U5456 ( .A(y[406]), .B(x[406]), .Z(n4340) );
  XNOR U5457 ( .A(y[407]), .B(x[407]), .Z(n4339) );
  XNOR U5458 ( .A(n4331), .B(n4332), .Z(n4342) );
  XNOR U5459 ( .A(y[402]), .B(x[402]), .Z(n4332) );
  XNOR U5460 ( .A(n4333), .B(n4334), .Z(n4331) );
  XNOR U5461 ( .A(y[403]), .B(x[403]), .Z(n4334) );
  XNOR U5462 ( .A(y[404]), .B(x[404]), .Z(n4333) );
  XOR U5463 ( .A(n4307), .B(n4308), .Z(n4326) );
  XNOR U5464 ( .A(n4323), .B(n4324), .Z(n4308) );
  XNOR U5465 ( .A(n4318), .B(n4319), .Z(n4324) );
  XNOR U5466 ( .A(n4320), .B(n4321), .Z(n4319) );
  XNOR U5467 ( .A(y[400]), .B(x[400]), .Z(n4321) );
  XNOR U5468 ( .A(y[401]), .B(x[401]), .Z(n4320) );
  XNOR U5469 ( .A(y[399]), .B(x[399]), .Z(n4318) );
  XNOR U5470 ( .A(n4312), .B(n4313), .Z(n4323) );
  XNOR U5471 ( .A(y[396]), .B(x[396]), .Z(n4313) );
  XNOR U5472 ( .A(n4314), .B(n4315), .Z(n4312) );
  XNOR U5473 ( .A(y[397]), .B(x[397]), .Z(n4315) );
  XNOR U5474 ( .A(y[398]), .B(x[398]), .Z(n4314) );
  XOR U5475 ( .A(n4306), .B(n4305), .Z(n4307) );
  XNOR U5476 ( .A(n4301), .B(n4302), .Z(n4305) );
  XNOR U5477 ( .A(y[393]), .B(x[393]), .Z(n4302) );
  XNOR U5478 ( .A(n4303), .B(n4304), .Z(n4301) );
  XNOR U5479 ( .A(y[394]), .B(x[394]), .Z(n4304) );
  XNOR U5480 ( .A(y[395]), .B(x[395]), .Z(n4303) );
  XNOR U5481 ( .A(n4295), .B(n4296), .Z(n4306) );
  XNOR U5482 ( .A(y[390]), .B(x[390]), .Z(n4296) );
  XNOR U5483 ( .A(n4297), .B(n4298), .Z(n4295) );
  XNOR U5484 ( .A(y[391]), .B(x[391]), .Z(n4298) );
  XNOR U5485 ( .A(y[392]), .B(x[392]), .Z(n4297) );
  NAND U5486 ( .A(n4362), .B(n4363), .Z(N5948) );
  NANDN U5487 ( .A(n4364), .B(n4365), .Z(n4363) );
  OR U5488 ( .A(n4366), .B(n4367), .Z(n4365) );
  NAND U5489 ( .A(n4366), .B(n4367), .Z(n4362) );
  XOR U5490 ( .A(n4366), .B(n4368), .Z(N5947) );
  XNOR U5491 ( .A(n4364), .B(n4367), .Z(n4368) );
  AND U5492 ( .A(n4369), .B(n4370), .Z(n4367) );
  NANDN U5493 ( .A(n4371), .B(n4372), .Z(n4370) );
  NANDN U5494 ( .A(n4373), .B(n4374), .Z(n4372) );
  NANDN U5495 ( .A(n4374), .B(n4373), .Z(n4369) );
  NAND U5496 ( .A(n4375), .B(n4376), .Z(n4364) );
  NANDN U5497 ( .A(n4377), .B(n4378), .Z(n4376) );
  OR U5498 ( .A(n4379), .B(n4380), .Z(n4378) );
  NAND U5499 ( .A(n4380), .B(n4379), .Z(n4375) );
  AND U5500 ( .A(n4381), .B(n4382), .Z(n4366) );
  NANDN U5501 ( .A(n4383), .B(n4384), .Z(n4382) );
  NANDN U5502 ( .A(n4385), .B(n4386), .Z(n4384) );
  NANDN U5503 ( .A(n4386), .B(n4385), .Z(n4381) );
  XOR U5504 ( .A(n4380), .B(n4387), .Z(N5946) );
  XOR U5505 ( .A(n4377), .B(n4379), .Z(n4387) );
  XNOR U5506 ( .A(n4373), .B(n4388), .Z(n4379) );
  XNOR U5507 ( .A(n4371), .B(n4374), .Z(n4388) );
  NAND U5508 ( .A(n4389), .B(n4390), .Z(n4374) );
  NAND U5509 ( .A(n4391), .B(n4392), .Z(n4390) );
  OR U5510 ( .A(n4393), .B(n4394), .Z(n4391) );
  NANDN U5511 ( .A(n4395), .B(n4393), .Z(n4389) );
  IV U5512 ( .A(n4394), .Z(n4395) );
  NAND U5513 ( .A(n4396), .B(n4397), .Z(n4371) );
  NAND U5514 ( .A(n4398), .B(n4399), .Z(n4397) );
  NANDN U5515 ( .A(n4400), .B(n4401), .Z(n4398) );
  NANDN U5516 ( .A(n4401), .B(n4400), .Z(n4396) );
  AND U5517 ( .A(n4402), .B(n4403), .Z(n4373) );
  NAND U5518 ( .A(n4404), .B(n4405), .Z(n4403) );
  OR U5519 ( .A(n4406), .B(n4407), .Z(n4404) );
  NANDN U5520 ( .A(n4408), .B(n4406), .Z(n4402) );
  NAND U5521 ( .A(n4409), .B(n4410), .Z(n4377) );
  NANDN U5522 ( .A(n4411), .B(n4412), .Z(n4410) );
  OR U5523 ( .A(n4413), .B(n4414), .Z(n4412) );
  NANDN U5524 ( .A(n4415), .B(n4413), .Z(n4409) );
  IV U5525 ( .A(n4414), .Z(n4415) );
  XNOR U5526 ( .A(n4385), .B(n4416), .Z(n4380) );
  XNOR U5527 ( .A(n4383), .B(n4386), .Z(n4416) );
  NAND U5528 ( .A(n4417), .B(n4418), .Z(n4386) );
  NAND U5529 ( .A(n4419), .B(n4420), .Z(n4418) );
  OR U5530 ( .A(n4421), .B(n4422), .Z(n4419) );
  NANDN U5531 ( .A(n4423), .B(n4421), .Z(n4417) );
  IV U5532 ( .A(n4422), .Z(n4423) );
  NAND U5533 ( .A(n4424), .B(n4425), .Z(n4383) );
  NAND U5534 ( .A(n4426), .B(n4427), .Z(n4425) );
  NANDN U5535 ( .A(n4428), .B(n4429), .Z(n4426) );
  NANDN U5536 ( .A(n4429), .B(n4428), .Z(n4424) );
  AND U5537 ( .A(n4430), .B(n4431), .Z(n4385) );
  NAND U5538 ( .A(n4432), .B(n4433), .Z(n4431) );
  OR U5539 ( .A(n4434), .B(n4435), .Z(n4432) );
  NANDN U5540 ( .A(n4436), .B(n4434), .Z(n4430) );
  XNOR U5541 ( .A(n4411), .B(n4437), .Z(N5945) );
  XOR U5542 ( .A(n4413), .B(n4414), .Z(n4437) );
  XNOR U5543 ( .A(n4427), .B(n4438), .Z(n4414) );
  XOR U5544 ( .A(n4428), .B(n4429), .Z(n4438) );
  XOR U5545 ( .A(n4434), .B(n4439), .Z(n4429) );
  XOR U5546 ( .A(n4433), .B(n4436), .Z(n4439) );
  IV U5547 ( .A(n4435), .Z(n4436) );
  NAND U5548 ( .A(n4440), .B(n4441), .Z(n4435) );
  OR U5549 ( .A(n4442), .B(n4443), .Z(n4441) );
  OR U5550 ( .A(n4444), .B(n4445), .Z(n4440) );
  NAND U5551 ( .A(n4446), .B(n4447), .Z(n4433) );
  OR U5552 ( .A(n4448), .B(n4449), .Z(n4447) );
  OR U5553 ( .A(n4450), .B(n4451), .Z(n4446) );
  NOR U5554 ( .A(n4452), .B(n4453), .Z(n4434) );
  ANDN U5555 ( .B(n4454), .A(n4455), .Z(n4428) );
  XNOR U5556 ( .A(n4421), .B(n4456), .Z(n4427) );
  XNOR U5557 ( .A(n4420), .B(n4422), .Z(n4456) );
  NAND U5558 ( .A(n4457), .B(n4458), .Z(n4422) );
  OR U5559 ( .A(n4459), .B(n4460), .Z(n4458) );
  OR U5560 ( .A(n4461), .B(n4462), .Z(n4457) );
  NAND U5561 ( .A(n4463), .B(n4464), .Z(n4420) );
  OR U5562 ( .A(n4465), .B(n4466), .Z(n4464) );
  OR U5563 ( .A(n4467), .B(n4468), .Z(n4463) );
  ANDN U5564 ( .B(n4469), .A(n4470), .Z(n4421) );
  IV U5565 ( .A(n4471), .Z(n4469) );
  ANDN U5566 ( .B(n4472), .A(n4473), .Z(n4413) );
  XOR U5567 ( .A(n4399), .B(n4474), .Z(n4411) );
  XOR U5568 ( .A(n4400), .B(n4401), .Z(n4474) );
  XOR U5569 ( .A(n4406), .B(n4475), .Z(n4401) );
  XOR U5570 ( .A(n4405), .B(n4408), .Z(n4475) );
  IV U5571 ( .A(n4407), .Z(n4408) );
  NAND U5572 ( .A(n4476), .B(n4477), .Z(n4407) );
  OR U5573 ( .A(n4478), .B(n4479), .Z(n4477) );
  OR U5574 ( .A(n4480), .B(n4481), .Z(n4476) );
  NAND U5575 ( .A(n4482), .B(n4483), .Z(n4405) );
  OR U5576 ( .A(n4484), .B(n4485), .Z(n4483) );
  OR U5577 ( .A(n4486), .B(n4487), .Z(n4482) );
  NOR U5578 ( .A(n4488), .B(n4489), .Z(n4406) );
  ANDN U5579 ( .B(n4490), .A(n4491), .Z(n4400) );
  IV U5580 ( .A(n4492), .Z(n4490) );
  XNOR U5581 ( .A(n4393), .B(n4493), .Z(n4399) );
  XNOR U5582 ( .A(n4392), .B(n4394), .Z(n4493) );
  NAND U5583 ( .A(n4494), .B(n4495), .Z(n4394) );
  OR U5584 ( .A(n4496), .B(n4497), .Z(n4495) );
  OR U5585 ( .A(n4498), .B(n4499), .Z(n4494) );
  NAND U5586 ( .A(n4500), .B(n4501), .Z(n4392) );
  OR U5587 ( .A(n4502), .B(n4503), .Z(n4501) );
  OR U5588 ( .A(n4504), .B(n4505), .Z(n4500) );
  ANDN U5589 ( .B(n4506), .A(n4507), .Z(n4393) );
  IV U5590 ( .A(n4508), .Z(n4506) );
  XNOR U5591 ( .A(n4473), .B(n4472), .Z(N5944) );
  XOR U5592 ( .A(n4492), .B(n4491), .Z(n4472) );
  XNOR U5593 ( .A(n4507), .B(n4508), .Z(n4491) );
  XNOR U5594 ( .A(n4502), .B(n4503), .Z(n4508) );
  XNOR U5595 ( .A(n4504), .B(n4505), .Z(n4503) );
  XNOR U5596 ( .A(y[388]), .B(x[388]), .Z(n4505) );
  XNOR U5597 ( .A(y[389]), .B(x[389]), .Z(n4504) );
  XNOR U5598 ( .A(y[387]), .B(x[387]), .Z(n4502) );
  XNOR U5599 ( .A(n4496), .B(n4497), .Z(n4507) );
  XNOR U5600 ( .A(y[384]), .B(x[384]), .Z(n4497) );
  XNOR U5601 ( .A(n4498), .B(n4499), .Z(n4496) );
  XNOR U5602 ( .A(y[385]), .B(x[385]), .Z(n4499) );
  XNOR U5603 ( .A(y[386]), .B(x[386]), .Z(n4498) );
  XNOR U5604 ( .A(n4489), .B(n4488), .Z(n4492) );
  XNOR U5605 ( .A(n4484), .B(n4485), .Z(n4488) );
  XNOR U5606 ( .A(y[381]), .B(x[381]), .Z(n4485) );
  XNOR U5607 ( .A(n4486), .B(n4487), .Z(n4484) );
  XNOR U5608 ( .A(y[382]), .B(x[382]), .Z(n4487) );
  XNOR U5609 ( .A(y[383]), .B(x[383]), .Z(n4486) );
  XNOR U5610 ( .A(n4478), .B(n4479), .Z(n4489) );
  XNOR U5611 ( .A(y[378]), .B(x[378]), .Z(n4479) );
  XNOR U5612 ( .A(n4480), .B(n4481), .Z(n4478) );
  XNOR U5613 ( .A(y[379]), .B(x[379]), .Z(n4481) );
  XNOR U5614 ( .A(y[380]), .B(x[380]), .Z(n4480) );
  XOR U5615 ( .A(n4454), .B(n4455), .Z(n4473) );
  XNOR U5616 ( .A(n4470), .B(n4471), .Z(n4455) );
  XNOR U5617 ( .A(n4465), .B(n4466), .Z(n4471) );
  XNOR U5618 ( .A(n4467), .B(n4468), .Z(n4466) );
  XNOR U5619 ( .A(y[376]), .B(x[376]), .Z(n4468) );
  XNOR U5620 ( .A(y[377]), .B(x[377]), .Z(n4467) );
  XNOR U5621 ( .A(y[375]), .B(x[375]), .Z(n4465) );
  XNOR U5622 ( .A(n4459), .B(n4460), .Z(n4470) );
  XNOR U5623 ( .A(y[372]), .B(x[372]), .Z(n4460) );
  XNOR U5624 ( .A(n4461), .B(n4462), .Z(n4459) );
  XNOR U5625 ( .A(y[373]), .B(x[373]), .Z(n4462) );
  XNOR U5626 ( .A(y[374]), .B(x[374]), .Z(n4461) );
  XOR U5627 ( .A(n4453), .B(n4452), .Z(n4454) );
  XNOR U5628 ( .A(n4448), .B(n4449), .Z(n4452) );
  XNOR U5629 ( .A(y[369]), .B(x[369]), .Z(n4449) );
  XNOR U5630 ( .A(n4450), .B(n4451), .Z(n4448) );
  XNOR U5631 ( .A(y[370]), .B(x[370]), .Z(n4451) );
  XNOR U5632 ( .A(y[371]), .B(x[371]), .Z(n4450) );
  XNOR U5633 ( .A(n4442), .B(n4443), .Z(n4453) );
  XNOR U5634 ( .A(y[366]), .B(x[366]), .Z(n4443) );
  XNOR U5635 ( .A(n4444), .B(n4445), .Z(n4442) );
  XNOR U5636 ( .A(y[367]), .B(x[367]), .Z(n4445) );
  XNOR U5637 ( .A(y[368]), .B(x[368]), .Z(n4444) );
  NAND U5638 ( .A(n4509), .B(n4510), .Z(N5938) );
  NANDN U5639 ( .A(n4511), .B(n4512), .Z(n4510) );
  OR U5640 ( .A(n4513), .B(n4514), .Z(n4512) );
  NAND U5641 ( .A(n4513), .B(n4514), .Z(n4509) );
  XOR U5642 ( .A(n4513), .B(n4515), .Z(N5937) );
  XNOR U5643 ( .A(n4511), .B(n4514), .Z(n4515) );
  AND U5644 ( .A(n4516), .B(n4517), .Z(n4514) );
  NANDN U5645 ( .A(n4518), .B(n4519), .Z(n4517) );
  NANDN U5646 ( .A(n4520), .B(n4521), .Z(n4519) );
  NANDN U5647 ( .A(n4521), .B(n4520), .Z(n4516) );
  NAND U5648 ( .A(n4522), .B(n4523), .Z(n4511) );
  NANDN U5649 ( .A(n4524), .B(n4525), .Z(n4523) );
  OR U5650 ( .A(n4526), .B(n4527), .Z(n4525) );
  NAND U5651 ( .A(n4527), .B(n4526), .Z(n4522) );
  AND U5652 ( .A(n4528), .B(n4529), .Z(n4513) );
  NANDN U5653 ( .A(n4530), .B(n4531), .Z(n4529) );
  NANDN U5654 ( .A(n4532), .B(n4533), .Z(n4531) );
  NANDN U5655 ( .A(n4533), .B(n4532), .Z(n4528) );
  XOR U5656 ( .A(n4527), .B(n4534), .Z(N5936) );
  XOR U5657 ( .A(n4524), .B(n4526), .Z(n4534) );
  XNOR U5658 ( .A(n4520), .B(n4535), .Z(n4526) );
  XNOR U5659 ( .A(n4518), .B(n4521), .Z(n4535) );
  NAND U5660 ( .A(n4536), .B(n4537), .Z(n4521) );
  NAND U5661 ( .A(n4538), .B(n4539), .Z(n4537) );
  OR U5662 ( .A(n4540), .B(n4541), .Z(n4538) );
  NANDN U5663 ( .A(n4542), .B(n4540), .Z(n4536) );
  IV U5664 ( .A(n4541), .Z(n4542) );
  NAND U5665 ( .A(n4543), .B(n4544), .Z(n4518) );
  NAND U5666 ( .A(n4545), .B(n4546), .Z(n4544) );
  NANDN U5667 ( .A(n4547), .B(n4548), .Z(n4545) );
  NANDN U5668 ( .A(n4548), .B(n4547), .Z(n4543) );
  AND U5669 ( .A(n4549), .B(n4550), .Z(n4520) );
  NAND U5670 ( .A(n4551), .B(n4552), .Z(n4550) );
  OR U5671 ( .A(n4553), .B(n4554), .Z(n4551) );
  NANDN U5672 ( .A(n4555), .B(n4553), .Z(n4549) );
  NAND U5673 ( .A(n4556), .B(n4557), .Z(n4524) );
  NANDN U5674 ( .A(n4558), .B(n4559), .Z(n4557) );
  OR U5675 ( .A(n4560), .B(n4561), .Z(n4559) );
  NANDN U5676 ( .A(n4562), .B(n4560), .Z(n4556) );
  IV U5677 ( .A(n4561), .Z(n4562) );
  XNOR U5678 ( .A(n4532), .B(n4563), .Z(n4527) );
  XNOR U5679 ( .A(n4530), .B(n4533), .Z(n4563) );
  NAND U5680 ( .A(n4564), .B(n4565), .Z(n4533) );
  NAND U5681 ( .A(n4566), .B(n4567), .Z(n4565) );
  OR U5682 ( .A(n4568), .B(n4569), .Z(n4566) );
  NANDN U5683 ( .A(n4570), .B(n4568), .Z(n4564) );
  IV U5684 ( .A(n4569), .Z(n4570) );
  NAND U5685 ( .A(n4571), .B(n4572), .Z(n4530) );
  NAND U5686 ( .A(n4573), .B(n4574), .Z(n4572) );
  NANDN U5687 ( .A(n4575), .B(n4576), .Z(n4573) );
  NANDN U5688 ( .A(n4576), .B(n4575), .Z(n4571) );
  AND U5689 ( .A(n4577), .B(n4578), .Z(n4532) );
  NAND U5690 ( .A(n4579), .B(n4580), .Z(n4578) );
  OR U5691 ( .A(n4581), .B(n4582), .Z(n4579) );
  NANDN U5692 ( .A(n4583), .B(n4581), .Z(n4577) );
  XNOR U5693 ( .A(n4558), .B(n4584), .Z(N5935) );
  XOR U5694 ( .A(n4560), .B(n4561), .Z(n4584) );
  XNOR U5695 ( .A(n4574), .B(n4585), .Z(n4561) );
  XOR U5696 ( .A(n4575), .B(n4576), .Z(n4585) );
  XOR U5697 ( .A(n4581), .B(n4586), .Z(n4576) );
  XOR U5698 ( .A(n4580), .B(n4583), .Z(n4586) );
  IV U5699 ( .A(n4582), .Z(n4583) );
  NAND U5700 ( .A(n4587), .B(n4588), .Z(n4582) );
  OR U5701 ( .A(n4589), .B(n4590), .Z(n4588) );
  OR U5702 ( .A(n4591), .B(n4592), .Z(n4587) );
  NAND U5703 ( .A(n4593), .B(n4594), .Z(n4580) );
  OR U5704 ( .A(n4595), .B(n4596), .Z(n4594) );
  OR U5705 ( .A(n4597), .B(n4598), .Z(n4593) );
  NOR U5706 ( .A(n4599), .B(n4600), .Z(n4581) );
  ANDN U5707 ( .B(n4601), .A(n4602), .Z(n4575) );
  XNOR U5708 ( .A(n4568), .B(n4603), .Z(n4574) );
  XNOR U5709 ( .A(n4567), .B(n4569), .Z(n4603) );
  NAND U5710 ( .A(n4604), .B(n4605), .Z(n4569) );
  OR U5711 ( .A(n4606), .B(n4607), .Z(n4605) );
  OR U5712 ( .A(n4608), .B(n4609), .Z(n4604) );
  NAND U5713 ( .A(n4610), .B(n4611), .Z(n4567) );
  OR U5714 ( .A(n4612), .B(n4613), .Z(n4611) );
  OR U5715 ( .A(n4614), .B(n4615), .Z(n4610) );
  ANDN U5716 ( .B(n4616), .A(n4617), .Z(n4568) );
  IV U5717 ( .A(n4618), .Z(n4616) );
  ANDN U5718 ( .B(n4619), .A(n4620), .Z(n4560) );
  XOR U5719 ( .A(n4546), .B(n4621), .Z(n4558) );
  XOR U5720 ( .A(n4547), .B(n4548), .Z(n4621) );
  XOR U5721 ( .A(n4553), .B(n4622), .Z(n4548) );
  XOR U5722 ( .A(n4552), .B(n4555), .Z(n4622) );
  IV U5723 ( .A(n4554), .Z(n4555) );
  NAND U5724 ( .A(n4623), .B(n4624), .Z(n4554) );
  OR U5725 ( .A(n4625), .B(n4626), .Z(n4624) );
  OR U5726 ( .A(n4627), .B(n4628), .Z(n4623) );
  NAND U5727 ( .A(n4629), .B(n4630), .Z(n4552) );
  OR U5728 ( .A(n4631), .B(n4632), .Z(n4630) );
  OR U5729 ( .A(n4633), .B(n4634), .Z(n4629) );
  NOR U5730 ( .A(n4635), .B(n4636), .Z(n4553) );
  ANDN U5731 ( .B(n4637), .A(n4638), .Z(n4547) );
  IV U5732 ( .A(n4639), .Z(n4637) );
  XNOR U5733 ( .A(n4540), .B(n4640), .Z(n4546) );
  XNOR U5734 ( .A(n4539), .B(n4541), .Z(n4640) );
  NAND U5735 ( .A(n4641), .B(n4642), .Z(n4541) );
  OR U5736 ( .A(n4643), .B(n4644), .Z(n4642) );
  OR U5737 ( .A(n4645), .B(n4646), .Z(n4641) );
  NAND U5738 ( .A(n4647), .B(n4648), .Z(n4539) );
  OR U5739 ( .A(n4649), .B(n4650), .Z(n4648) );
  OR U5740 ( .A(n4651), .B(n4652), .Z(n4647) );
  ANDN U5741 ( .B(n4653), .A(n4654), .Z(n4540) );
  IV U5742 ( .A(n4655), .Z(n4653) );
  XNOR U5743 ( .A(n4620), .B(n4619), .Z(N5934) );
  XOR U5744 ( .A(n4639), .B(n4638), .Z(n4619) );
  XNOR U5745 ( .A(n4654), .B(n4655), .Z(n4638) );
  XNOR U5746 ( .A(n4649), .B(n4650), .Z(n4655) );
  XNOR U5747 ( .A(n4651), .B(n4652), .Z(n4650) );
  XNOR U5748 ( .A(y[364]), .B(x[364]), .Z(n4652) );
  XNOR U5749 ( .A(y[365]), .B(x[365]), .Z(n4651) );
  XNOR U5750 ( .A(y[363]), .B(x[363]), .Z(n4649) );
  XNOR U5751 ( .A(n4643), .B(n4644), .Z(n4654) );
  XNOR U5752 ( .A(y[360]), .B(x[360]), .Z(n4644) );
  XNOR U5753 ( .A(n4645), .B(n4646), .Z(n4643) );
  XNOR U5754 ( .A(y[361]), .B(x[361]), .Z(n4646) );
  XNOR U5755 ( .A(y[362]), .B(x[362]), .Z(n4645) );
  XNOR U5756 ( .A(n4636), .B(n4635), .Z(n4639) );
  XNOR U5757 ( .A(n4631), .B(n4632), .Z(n4635) );
  XNOR U5758 ( .A(y[357]), .B(x[357]), .Z(n4632) );
  XNOR U5759 ( .A(n4633), .B(n4634), .Z(n4631) );
  XNOR U5760 ( .A(y[358]), .B(x[358]), .Z(n4634) );
  XNOR U5761 ( .A(y[359]), .B(x[359]), .Z(n4633) );
  XNOR U5762 ( .A(n4625), .B(n4626), .Z(n4636) );
  XNOR U5763 ( .A(y[354]), .B(x[354]), .Z(n4626) );
  XNOR U5764 ( .A(n4627), .B(n4628), .Z(n4625) );
  XNOR U5765 ( .A(y[355]), .B(x[355]), .Z(n4628) );
  XNOR U5766 ( .A(y[356]), .B(x[356]), .Z(n4627) );
  XOR U5767 ( .A(n4601), .B(n4602), .Z(n4620) );
  XNOR U5768 ( .A(n4617), .B(n4618), .Z(n4602) );
  XNOR U5769 ( .A(n4612), .B(n4613), .Z(n4618) );
  XNOR U5770 ( .A(n4614), .B(n4615), .Z(n4613) );
  XNOR U5771 ( .A(y[352]), .B(x[352]), .Z(n4615) );
  XNOR U5772 ( .A(y[353]), .B(x[353]), .Z(n4614) );
  XNOR U5773 ( .A(y[351]), .B(x[351]), .Z(n4612) );
  XNOR U5774 ( .A(n4606), .B(n4607), .Z(n4617) );
  XNOR U5775 ( .A(y[348]), .B(x[348]), .Z(n4607) );
  XNOR U5776 ( .A(n4608), .B(n4609), .Z(n4606) );
  XNOR U5777 ( .A(y[349]), .B(x[349]), .Z(n4609) );
  XNOR U5778 ( .A(y[350]), .B(x[350]), .Z(n4608) );
  XOR U5779 ( .A(n4600), .B(n4599), .Z(n4601) );
  XNOR U5780 ( .A(n4595), .B(n4596), .Z(n4599) );
  XNOR U5781 ( .A(y[345]), .B(x[345]), .Z(n4596) );
  XNOR U5782 ( .A(n4597), .B(n4598), .Z(n4595) );
  XNOR U5783 ( .A(y[346]), .B(x[346]), .Z(n4598) );
  XNOR U5784 ( .A(y[347]), .B(x[347]), .Z(n4597) );
  XNOR U5785 ( .A(n4589), .B(n4590), .Z(n4600) );
  XNOR U5786 ( .A(y[342]), .B(x[342]), .Z(n4590) );
  XNOR U5787 ( .A(n4591), .B(n4592), .Z(n4589) );
  XNOR U5788 ( .A(y[343]), .B(x[343]), .Z(n4592) );
  XNOR U5789 ( .A(y[344]), .B(x[344]), .Z(n4591) );
  NAND U5790 ( .A(n4656), .B(n4657), .Z(N5928) );
  NANDN U5791 ( .A(n4658), .B(n4659), .Z(n4657) );
  OR U5792 ( .A(n4660), .B(n4661), .Z(n4659) );
  NAND U5793 ( .A(n4660), .B(n4661), .Z(n4656) );
  XOR U5794 ( .A(n4660), .B(n4662), .Z(N5927) );
  XNOR U5795 ( .A(n4658), .B(n4661), .Z(n4662) );
  AND U5796 ( .A(n4663), .B(n4664), .Z(n4661) );
  NANDN U5797 ( .A(n4665), .B(n4666), .Z(n4664) );
  NANDN U5798 ( .A(n4667), .B(n4668), .Z(n4666) );
  NANDN U5799 ( .A(n4668), .B(n4667), .Z(n4663) );
  NAND U5800 ( .A(n4669), .B(n4670), .Z(n4658) );
  NANDN U5801 ( .A(n4671), .B(n4672), .Z(n4670) );
  OR U5802 ( .A(n4673), .B(n4674), .Z(n4672) );
  NAND U5803 ( .A(n4674), .B(n4673), .Z(n4669) );
  AND U5804 ( .A(n4675), .B(n4676), .Z(n4660) );
  NANDN U5805 ( .A(n4677), .B(n4678), .Z(n4676) );
  NANDN U5806 ( .A(n4679), .B(n4680), .Z(n4678) );
  NANDN U5807 ( .A(n4680), .B(n4679), .Z(n4675) );
  XOR U5808 ( .A(n4674), .B(n4681), .Z(N5926) );
  XOR U5809 ( .A(n4671), .B(n4673), .Z(n4681) );
  XNOR U5810 ( .A(n4667), .B(n4682), .Z(n4673) );
  XNOR U5811 ( .A(n4665), .B(n4668), .Z(n4682) );
  NAND U5812 ( .A(n4683), .B(n4684), .Z(n4668) );
  NAND U5813 ( .A(n4685), .B(n4686), .Z(n4684) );
  OR U5814 ( .A(n4687), .B(n4688), .Z(n4685) );
  NANDN U5815 ( .A(n4689), .B(n4687), .Z(n4683) );
  IV U5816 ( .A(n4688), .Z(n4689) );
  NAND U5817 ( .A(n4690), .B(n4691), .Z(n4665) );
  NAND U5818 ( .A(n4692), .B(n4693), .Z(n4691) );
  NANDN U5819 ( .A(n4694), .B(n4695), .Z(n4692) );
  NANDN U5820 ( .A(n4695), .B(n4694), .Z(n4690) );
  AND U5821 ( .A(n4696), .B(n4697), .Z(n4667) );
  NAND U5822 ( .A(n4698), .B(n4699), .Z(n4697) );
  OR U5823 ( .A(n4700), .B(n4701), .Z(n4698) );
  NANDN U5824 ( .A(n4702), .B(n4700), .Z(n4696) );
  NAND U5825 ( .A(n4703), .B(n4704), .Z(n4671) );
  NANDN U5826 ( .A(n4705), .B(n4706), .Z(n4704) );
  OR U5827 ( .A(n4707), .B(n4708), .Z(n4706) );
  NANDN U5828 ( .A(n4709), .B(n4707), .Z(n4703) );
  IV U5829 ( .A(n4708), .Z(n4709) );
  XNOR U5830 ( .A(n4679), .B(n4710), .Z(n4674) );
  XNOR U5831 ( .A(n4677), .B(n4680), .Z(n4710) );
  NAND U5832 ( .A(n4711), .B(n4712), .Z(n4680) );
  NAND U5833 ( .A(n4713), .B(n4714), .Z(n4712) );
  OR U5834 ( .A(n4715), .B(n4716), .Z(n4713) );
  NANDN U5835 ( .A(n4717), .B(n4715), .Z(n4711) );
  IV U5836 ( .A(n4716), .Z(n4717) );
  NAND U5837 ( .A(n4718), .B(n4719), .Z(n4677) );
  NAND U5838 ( .A(n4720), .B(n4721), .Z(n4719) );
  NANDN U5839 ( .A(n4722), .B(n4723), .Z(n4720) );
  NANDN U5840 ( .A(n4723), .B(n4722), .Z(n4718) );
  AND U5841 ( .A(n4724), .B(n4725), .Z(n4679) );
  NAND U5842 ( .A(n4726), .B(n4727), .Z(n4725) );
  OR U5843 ( .A(n4728), .B(n4729), .Z(n4726) );
  NANDN U5844 ( .A(n4730), .B(n4728), .Z(n4724) );
  XNOR U5845 ( .A(n4705), .B(n4731), .Z(N5925) );
  XOR U5846 ( .A(n4707), .B(n4708), .Z(n4731) );
  XNOR U5847 ( .A(n4721), .B(n4732), .Z(n4708) );
  XOR U5848 ( .A(n4722), .B(n4723), .Z(n4732) );
  XOR U5849 ( .A(n4728), .B(n4733), .Z(n4723) );
  XOR U5850 ( .A(n4727), .B(n4730), .Z(n4733) );
  IV U5851 ( .A(n4729), .Z(n4730) );
  NAND U5852 ( .A(n4734), .B(n4735), .Z(n4729) );
  OR U5853 ( .A(n4736), .B(n4737), .Z(n4735) );
  OR U5854 ( .A(n4738), .B(n4739), .Z(n4734) );
  NAND U5855 ( .A(n4740), .B(n4741), .Z(n4727) );
  OR U5856 ( .A(n4742), .B(n4743), .Z(n4741) );
  OR U5857 ( .A(n4744), .B(n4745), .Z(n4740) );
  NOR U5858 ( .A(n4746), .B(n4747), .Z(n4728) );
  ANDN U5859 ( .B(n4748), .A(n4749), .Z(n4722) );
  XNOR U5860 ( .A(n4715), .B(n4750), .Z(n4721) );
  XNOR U5861 ( .A(n4714), .B(n4716), .Z(n4750) );
  NAND U5862 ( .A(n4751), .B(n4752), .Z(n4716) );
  OR U5863 ( .A(n4753), .B(n4754), .Z(n4752) );
  OR U5864 ( .A(n4755), .B(n4756), .Z(n4751) );
  NAND U5865 ( .A(n4757), .B(n4758), .Z(n4714) );
  OR U5866 ( .A(n4759), .B(n4760), .Z(n4758) );
  OR U5867 ( .A(n4761), .B(n4762), .Z(n4757) );
  ANDN U5868 ( .B(n4763), .A(n4764), .Z(n4715) );
  IV U5869 ( .A(n4765), .Z(n4763) );
  ANDN U5870 ( .B(n4766), .A(n4767), .Z(n4707) );
  XOR U5871 ( .A(n4693), .B(n4768), .Z(n4705) );
  XOR U5872 ( .A(n4694), .B(n4695), .Z(n4768) );
  XOR U5873 ( .A(n4700), .B(n4769), .Z(n4695) );
  XOR U5874 ( .A(n4699), .B(n4702), .Z(n4769) );
  IV U5875 ( .A(n4701), .Z(n4702) );
  NAND U5876 ( .A(n4770), .B(n4771), .Z(n4701) );
  OR U5877 ( .A(n4772), .B(n4773), .Z(n4771) );
  OR U5878 ( .A(n4774), .B(n4775), .Z(n4770) );
  NAND U5879 ( .A(n4776), .B(n4777), .Z(n4699) );
  OR U5880 ( .A(n4778), .B(n4779), .Z(n4777) );
  OR U5881 ( .A(n4780), .B(n4781), .Z(n4776) );
  NOR U5882 ( .A(n4782), .B(n4783), .Z(n4700) );
  ANDN U5883 ( .B(n4784), .A(n4785), .Z(n4694) );
  IV U5884 ( .A(n4786), .Z(n4784) );
  XNOR U5885 ( .A(n4687), .B(n4787), .Z(n4693) );
  XNOR U5886 ( .A(n4686), .B(n4688), .Z(n4787) );
  NAND U5887 ( .A(n4788), .B(n4789), .Z(n4688) );
  OR U5888 ( .A(n4790), .B(n4791), .Z(n4789) );
  OR U5889 ( .A(n4792), .B(n4793), .Z(n4788) );
  NAND U5890 ( .A(n4794), .B(n4795), .Z(n4686) );
  OR U5891 ( .A(n4796), .B(n4797), .Z(n4795) );
  OR U5892 ( .A(n4798), .B(n4799), .Z(n4794) );
  ANDN U5893 ( .B(n4800), .A(n4801), .Z(n4687) );
  IV U5894 ( .A(n4802), .Z(n4800) );
  XNOR U5895 ( .A(n4767), .B(n4766), .Z(N5924) );
  XOR U5896 ( .A(n4786), .B(n4785), .Z(n4766) );
  XNOR U5897 ( .A(n4801), .B(n4802), .Z(n4785) );
  XNOR U5898 ( .A(n4796), .B(n4797), .Z(n4802) );
  XNOR U5899 ( .A(n4798), .B(n4799), .Z(n4797) );
  XNOR U5900 ( .A(y[340]), .B(x[340]), .Z(n4799) );
  XNOR U5901 ( .A(y[341]), .B(x[341]), .Z(n4798) );
  XNOR U5902 ( .A(y[339]), .B(x[339]), .Z(n4796) );
  XNOR U5903 ( .A(n4790), .B(n4791), .Z(n4801) );
  XNOR U5904 ( .A(y[336]), .B(x[336]), .Z(n4791) );
  XNOR U5905 ( .A(n4792), .B(n4793), .Z(n4790) );
  XNOR U5906 ( .A(y[337]), .B(x[337]), .Z(n4793) );
  XNOR U5907 ( .A(y[338]), .B(x[338]), .Z(n4792) );
  XNOR U5908 ( .A(n4783), .B(n4782), .Z(n4786) );
  XNOR U5909 ( .A(n4778), .B(n4779), .Z(n4782) );
  XNOR U5910 ( .A(y[333]), .B(x[333]), .Z(n4779) );
  XNOR U5911 ( .A(n4780), .B(n4781), .Z(n4778) );
  XNOR U5912 ( .A(y[334]), .B(x[334]), .Z(n4781) );
  XNOR U5913 ( .A(y[335]), .B(x[335]), .Z(n4780) );
  XNOR U5914 ( .A(n4772), .B(n4773), .Z(n4783) );
  XNOR U5915 ( .A(y[330]), .B(x[330]), .Z(n4773) );
  XNOR U5916 ( .A(n4774), .B(n4775), .Z(n4772) );
  XNOR U5917 ( .A(y[331]), .B(x[331]), .Z(n4775) );
  XNOR U5918 ( .A(y[332]), .B(x[332]), .Z(n4774) );
  XOR U5919 ( .A(n4748), .B(n4749), .Z(n4767) );
  XNOR U5920 ( .A(n4764), .B(n4765), .Z(n4749) );
  XNOR U5921 ( .A(n4759), .B(n4760), .Z(n4765) );
  XNOR U5922 ( .A(n4761), .B(n4762), .Z(n4760) );
  XNOR U5923 ( .A(y[328]), .B(x[328]), .Z(n4762) );
  XNOR U5924 ( .A(y[329]), .B(x[329]), .Z(n4761) );
  XNOR U5925 ( .A(y[327]), .B(x[327]), .Z(n4759) );
  XNOR U5926 ( .A(n4753), .B(n4754), .Z(n4764) );
  XNOR U5927 ( .A(y[324]), .B(x[324]), .Z(n4754) );
  XNOR U5928 ( .A(n4755), .B(n4756), .Z(n4753) );
  XNOR U5929 ( .A(y[325]), .B(x[325]), .Z(n4756) );
  XNOR U5930 ( .A(y[326]), .B(x[326]), .Z(n4755) );
  XOR U5931 ( .A(n4747), .B(n4746), .Z(n4748) );
  XNOR U5932 ( .A(n4742), .B(n4743), .Z(n4746) );
  XNOR U5933 ( .A(y[321]), .B(x[321]), .Z(n4743) );
  XNOR U5934 ( .A(n4744), .B(n4745), .Z(n4742) );
  XNOR U5935 ( .A(y[322]), .B(x[322]), .Z(n4745) );
  XNOR U5936 ( .A(y[323]), .B(x[323]), .Z(n4744) );
  XNOR U5937 ( .A(n4736), .B(n4737), .Z(n4747) );
  XNOR U5938 ( .A(y[318]), .B(x[318]), .Z(n4737) );
  XNOR U5939 ( .A(n4738), .B(n4739), .Z(n4736) );
  XNOR U5940 ( .A(y[319]), .B(x[319]), .Z(n4739) );
  XNOR U5941 ( .A(y[320]), .B(x[320]), .Z(n4738) );
  NAND U5942 ( .A(n4803), .B(n4804), .Z(N5918) );
  NANDN U5943 ( .A(n4805), .B(n4806), .Z(n4804) );
  OR U5944 ( .A(n4807), .B(n4808), .Z(n4806) );
  NAND U5945 ( .A(n4807), .B(n4808), .Z(n4803) );
  XOR U5946 ( .A(n4807), .B(n4809), .Z(N5917) );
  XNOR U5947 ( .A(n4805), .B(n4808), .Z(n4809) );
  AND U5948 ( .A(n4810), .B(n4811), .Z(n4808) );
  NANDN U5949 ( .A(n4812), .B(n4813), .Z(n4811) );
  NANDN U5950 ( .A(n4814), .B(n4815), .Z(n4813) );
  NANDN U5951 ( .A(n4815), .B(n4814), .Z(n4810) );
  NAND U5952 ( .A(n4816), .B(n4817), .Z(n4805) );
  NANDN U5953 ( .A(n4818), .B(n4819), .Z(n4817) );
  OR U5954 ( .A(n4820), .B(n4821), .Z(n4819) );
  NAND U5955 ( .A(n4821), .B(n4820), .Z(n4816) );
  AND U5956 ( .A(n4822), .B(n4823), .Z(n4807) );
  NANDN U5957 ( .A(n4824), .B(n4825), .Z(n4823) );
  NANDN U5958 ( .A(n4826), .B(n4827), .Z(n4825) );
  NANDN U5959 ( .A(n4827), .B(n4826), .Z(n4822) );
  XOR U5960 ( .A(n4821), .B(n4828), .Z(N5916) );
  XOR U5961 ( .A(n4818), .B(n4820), .Z(n4828) );
  XNOR U5962 ( .A(n4814), .B(n4829), .Z(n4820) );
  XNOR U5963 ( .A(n4812), .B(n4815), .Z(n4829) );
  NAND U5964 ( .A(n4830), .B(n4831), .Z(n4815) );
  NAND U5965 ( .A(n4832), .B(n4833), .Z(n4831) );
  OR U5966 ( .A(n4834), .B(n4835), .Z(n4832) );
  NANDN U5967 ( .A(n4836), .B(n4834), .Z(n4830) );
  IV U5968 ( .A(n4835), .Z(n4836) );
  NAND U5969 ( .A(n4837), .B(n4838), .Z(n4812) );
  NAND U5970 ( .A(n4839), .B(n4840), .Z(n4838) );
  NANDN U5971 ( .A(n4841), .B(n4842), .Z(n4839) );
  NANDN U5972 ( .A(n4842), .B(n4841), .Z(n4837) );
  AND U5973 ( .A(n4843), .B(n4844), .Z(n4814) );
  NAND U5974 ( .A(n4845), .B(n4846), .Z(n4844) );
  OR U5975 ( .A(n4847), .B(n4848), .Z(n4845) );
  NANDN U5976 ( .A(n4849), .B(n4847), .Z(n4843) );
  NAND U5977 ( .A(n4850), .B(n4851), .Z(n4818) );
  NANDN U5978 ( .A(n4852), .B(n4853), .Z(n4851) );
  OR U5979 ( .A(n4854), .B(n4855), .Z(n4853) );
  NANDN U5980 ( .A(n4856), .B(n4854), .Z(n4850) );
  IV U5981 ( .A(n4855), .Z(n4856) );
  XNOR U5982 ( .A(n4826), .B(n4857), .Z(n4821) );
  XNOR U5983 ( .A(n4824), .B(n4827), .Z(n4857) );
  NAND U5984 ( .A(n4858), .B(n4859), .Z(n4827) );
  NAND U5985 ( .A(n4860), .B(n4861), .Z(n4859) );
  OR U5986 ( .A(n4862), .B(n4863), .Z(n4860) );
  NANDN U5987 ( .A(n4864), .B(n4862), .Z(n4858) );
  IV U5988 ( .A(n4863), .Z(n4864) );
  NAND U5989 ( .A(n4865), .B(n4866), .Z(n4824) );
  NAND U5990 ( .A(n4867), .B(n4868), .Z(n4866) );
  NANDN U5991 ( .A(n4869), .B(n4870), .Z(n4867) );
  NANDN U5992 ( .A(n4870), .B(n4869), .Z(n4865) );
  AND U5993 ( .A(n4871), .B(n4872), .Z(n4826) );
  NAND U5994 ( .A(n4873), .B(n4874), .Z(n4872) );
  OR U5995 ( .A(n4875), .B(n4876), .Z(n4873) );
  NANDN U5996 ( .A(n4877), .B(n4875), .Z(n4871) );
  XNOR U5997 ( .A(n4852), .B(n4878), .Z(N5915) );
  XOR U5998 ( .A(n4854), .B(n4855), .Z(n4878) );
  XNOR U5999 ( .A(n4868), .B(n4879), .Z(n4855) );
  XOR U6000 ( .A(n4869), .B(n4870), .Z(n4879) );
  XOR U6001 ( .A(n4875), .B(n4880), .Z(n4870) );
  XOR U6002 ( .A(n4874), .B(n4877), .Z(n4880) );
  IV U6003 ( .A(n4876), .Z(n4877) );
  NAND U6004 ( .A(n4881), .B(n4882), .Z(n4876) );
  OR U6005 ( .A(n4883), .B(n4884), .Z(n4882) );
  OR U6006 ( .A(n4885), .B(n4886), .Z(n4881) );
  NAND U6007 ( .A(n4887), .B(n4888), .Z(n4874) );
  OR U6008 ( .A(n4889), .B(n4890), .Z(n4888) );
  OR U6009 ( .A(n4891), .B(n4892), .Z(n4887) );
  NOR U6010 ( .A(n4893), .B(n4894), .Z(n4875) );
  ANDN U6011 ( .B(n4895), .A(n4896), .Z(n4869) );
  XNOR U6012 ( .A(n4862), .B(n4897), .Z(n4868) );
  XNOR U6013 ( .A(n4861), .B(n4863), .Z(n4897) );
  NAND U6014 ( .A(n4898), .B(n4899), .Z(n4863) );
  OR U6015 ( .A(n4900), .B(n4901), .Z(n4899) );
  OR U6016 ( .A(n4902), .B(n4903), .Z(n4898) );
  NAND U6017 ( .A(n4904), .B(n4905), .Z(n4861) );
  OR U6018 ( .A(n4906), .B(n4907), .Z(n4905) );
  OR U6019 ( .A(n4908), .B(n4909), .Z(n4904) );
  ANDN U6020 ( .B(n4910), .A(n4911), .Z(n4862) );
  IV U6021 ( .A(n4912), .Z(n4910) );
  ANDN U6022 ( .B(n4913), .A(n4914), .Z(n4854) );
  XOR U6023 ( .A(n4840), .B(n4915), .Z(n4852) );
  XOR U6024 ( .A(n4841), .B(n4842), .Z(n4915) );
  XOR U6025 ( .A(n4847), .B(n4916), .Z(n4842) );
  XOR U6026 ( .A(n4846), .B(n4849), .Z(n4916) );
  IV U6027 ( .A(n4848), .Z(n4849) );
  NAND U6028 ( .A(n4917), .B(n4918), .Z(n4848) );
  OR U6029 ( .A(n4919), .B(n4920), .Z(n4918) );
  OR U6030 ( .A(n4921), .B(n4922), .Z(n4917) );
  NAND U6031 ( .A(n4923), .B(n4924), .Z(n4846) );
  OR U6032 ( .A(n4925), .B(n4926), .Z(n4924) );
  OR U6033 ( .A(n4927), .B(n4928), .Z(n4923) );
  NOR U6034 ( .A(n4929), .B(n4930), .Z(n4847) );
  ANDN U6035 ( .B(n4931), .A(n4932), .Z(n4841) );
  IV U6036 ( .A(n4933), .Z(n4931) );
  XNOR U6037 ( .A(n4834), .B(n4934), .Z(n4840) );
  XNOR U6038 ( .A(n4833), .B(n4835), .Z(n4934) );
  NAND U6039 ( .A(n4935), .B(n4936), .Z(n4835) );
  OR U6040 ( .A(n4937), .B(n4938), .Z(n4936) );
  OR U6041 ( .A(n4939), .B(n4940), .Z(n4935) );
  NAND U6042 ( .A(n4941), .B(n4942), .Z(n4833) );
  OR U6043 ( .A(n4943), .B(n4944), .Z(n4942) );
  OR U6044 ( .A(n4945), .B(n4946), .Z(n4941) );
  ANDN U6045 ( .B(n4947), .A(n4948), .Z(n4834) );
  IV U6046 ( .A(n4949), .Z(n4947) );
  XNOR U6047 ( .A(n4914), .B(n4913), .Z(N5914) );
  XOR U6048 ( .A(n4933), .B(n4932), .Z(n4913) );
  XNOR U6049 ( .A(n4948), .B(n4949), .Z(n4932) );
  XNOR U6050 ( .A(n4943), .B(n4944), .Z(n4949) );
  XNOR U6051 ( .A(n4945), .B(n4946), .Z(n4944) );
  XNOR U6052 ( .A(y[316]), .B(x[316]), .Z(n4946) );
  XNOR U6053 ( .A(y[317]), .B(x[317]), .Z(n4945) );
  XNOR U6054 ( .A(y[315]), .B(x[315]), .Z(n4943) );
  XNOR U6055 ( .A(n4937), .B(n4938), .Z(n4948) );
  XNOR U6056 ( .A(y[312]), .B(x[312]), .Z(n4938) );
  XNOR U6057 ( .A(n4939), .B(n4940), .Z(n4937) );
  XNOR U6058 ( .A(y[313]), .B(x[313]), .Z(n4940) );
  XNOR U6059 ( .A(y[314]), .B(x[314]), .Z(n4939) );
  XNOR U6060 ( .A(n4930), .B(n4929), .Z(n4933) );
  XNOR U6061 ( .A(n4925), .B(n4926), .Z(n4929) );
  XNOR U6062 ( .A(y[309]), .B(x[309]), .Z(n4926) );
  XNOR U6063 ( .A(n4927), .B(n4928), .Z(n4925) );
  XNOR U6064 ( .A(y[310]), .B(x[310]), .Z(n4928) );
  XNOR U6065 ( .A(y[311]), .B(x[311]), .Z(n4927) );
  XNOR U6066 ( .A(n4919), .B(n4920), .Z(n4930) );
  XNOR U6067 ( .A(y[306]), .B(x[306]), .Z(n4920) );
  XNOR U6068 ( .A(n4921), .B(n4922), .Z(n4919) );
  XNOR U6069 ( .A(y[307]), .B(x[307]), .Z(n4922) );
  XNOR U6070 ( .A(y[308]), .B(x[308]), .Z(n4921) );
  XOR U6071 ( .A(n4895), .B(n4896), .Z(n4914) );
  XNOR U6072 ( .A(n4911), .B(n4912), .Z(n4896) );
  XNOR U6073 ( .A(n4906), .B(n4907), .Z(n4912) );
  XNOR U6074 ( .A(n4908), .B(n4909), .Z(n4907) );
  XNOR U6075 ( .A(y[304]), .B(x[304]), .Z(n4909) );
  XNOR U6076 ( .A(y[305]), .B(x[305]), .Z(n4908) );
  XNOR U6077 ( .A(y[303]), .B(x[303]), .Z(n4906) );
  XNOR U6078 ( .A(n4900), .B(n4901), .Z(n4911) );
  XNOR U6079 ( .A(y[300]), .B(x[300]), .Z(n4901) );
  XNOR U6080 ( .A(n4902), .B(n4903), .Z(n4900) );
  XNOR U6081 ( .A(y[301]), .B(x[301]), .Z(n4903) );
  XNOR U6082 ( .A(y[302]), .B(x[302]), .Z(n4902) );
  XOR U6083 ( .A(n4894), .B(n4893), .Z(n4895) );
  XNOR U6084 ( .A(n4889), .B(n4890), .Z(n4893) );
  XNOR U6085 ( .A(y[297]), .B(x[297]), .Z(n4890) );
  XNOR U6086 ( .A(n4891), .B(n4892), .Z(n4889) );
  XNOR U6087 ( .A(y[298]), .B(x[298]), .Z(n4892) );
  XNOR U6088 ( .A(y[299]), .B(x[299]), .Z(n4891) );
  XNOR U6089 ( .A(n4883), .B(n4884), .Z(n4894) );
  XNOR U6090 ( .A(y[294]), .B(x[294]), .Z(n4884) );
  XNOR U6091 ( .A(n4885), .B(n4886), .Z(n4883) );
  XNOR U6092 ( .A(y[295]), .B(x[295]), .Z(n4886) );
  XNOR U6093 ( .A(y[296]), .B(x[296]), .Z(n4885) );
  NAND U6094 ( .A(n4950), .B(n4951), .Z(N5908) );
  NANDN U6095 ( .A(n4952), .B(n4953), .Z(n4951) );
  OR U6096 ( .A(n4954), .B(n4955), .Z(n4953) );
  NAND U6097 ( .A(n4954), .B(n4955), .Z(n4950) );
  XOR U6098 ( .A(n4954), .B(n4956), .Z(N5907) );
  XNOR U6099 ( .A(n4952), .B(n4955), .Z(n4956) );
  AND U6100 ( .A(n4957), .B(n4958), .Z(n4955) );
  NANDN U6101 ( .A(n4959), .B(n4960), .Z(n4958) );
  NANDN U6102 ( .A(n4961), .B(n4962), .Z(n4960) );
  NANDN U6103 ( .A(n4962), .B(n4961), .Z(n4957) );
  NAND U6104 ( .A(n4963), .B(n4964), .Z(n4952) );
  NANDN U6105 ( .A(n4965), .B(n4966), .Z(n4964) );
  OR U6106 ( .A(n4967), .B(n4968), .Z(n4966) );
  NAND U6107 ( .A(n4968), .B(n4967), .Z(n4963) );
  AND U6108 ( .A(n4969), .B(n4970), .Z(n4954) );
  NANDN U6109 ( .A(n4971), .B(n4972), .Z(n4970) );
  NANDN U6110 ( .A(n4973), .B(n4974), .Z(n4972) );
  NANDN U6111 ( .A(n4974), .B(n4973), .Z(n4969) );
  XOR U6112 ( .A(n4968), .B(n4975), .Z(N5906) );
  XOR U6113 ( .A(n4965), .B(n4967), .Z(n4975) );
  XNOR U6114 ( .A(n4961), .B(n4976), .Z(n4967) );
  XNOR U6115 ( .A(n4959), .B(n4962), .Z(n4976) );
  NAND U6116 ( .A(n4977), .B(n4978), .Z(n4962) );
  NAND U6117 ( .A(n4979), .B(n4980), .Z(n4978) );
  OR U6118 ( .A(n4981), .B(n4982), .Z(n4979) );
  NANDN U6119 ( .A(n4983), .B(n4981), .Z(n4977) );
  IV U6120 ( .A(n4982), .Z(n4983) );
  NAND U6121 ( .A(n4984), .B(n4985), .Z(n4959) );
  NAND U6122 ( .A(n4986), .B(n4987), .Z(n4985) );
  NANDN U6123 ( .A(n4988), .B(n4989), .Z(n4986) );
  NANDN U6124 ( .A(n4989), .B(n4988), .Z(n4984) );
  AND U6125 ( .A(n4990), .B(n4991), .Z(n4961) );
  NAND U6126 ( .A(n4992), .B(n4993), .Z(n4991) );
  OR U6127 ( .A(n4994), .B(n4995), .Z(n4992) );
  NANDN U6128 ( .A(n4996), .B(n4994), .Z(n4990) );
  NAND U6129 ( .A(n4997), .B(n4998), .Z(n4965) );
  NANDN U6130 ( .A(n4999), .B(n5000), .Z(n4998) );
  OR U6131 ( .A(n5001), .B(n5002), .Z(n5000) );
  NANDN U6132 ( .A(n5003), .B(n5001), .Z(n4997) );
  IV U6133 ( .A(n5002), .Z(n5003) );
  XNOR U6134 ( .A(n4973), .B(n5004), .Z(n4968) );
  XNOR U6135 ( .A(n4971), .B(n4974), .Z(n5004) );
  NAND U6136 ( .A(n5005), .B(n5006), .Z(n4974) );
  NAND U6137 ( .A(n5007), .B(n5008), .Z(n5006) );
  OR U6138 ( .A(n5009), .B(n5010), .Z(n5007) );
  NANDN U6139 ( .A(n5011), .B(n5009), .Z(n5005) );
  IV U6140 ( .A(n5010), .Z(n5011) );
  NAND U6141 ( .A(n5012), .B(n5013), .Z(n4971) );
  NAND U6142 ( .A(n5014), .B(n5015), .Z(n5013) );
  NANDN U6143 ( .A(n5016), .B(n5017), .Z(n5014) );
  NANDN U6144 ( .A(n5017), .B(n5016), .Z(n5012) );
  AND U6145 ( .A(n5018), .B(n5019), .Z(n4973) );
  NAND U6146 ( .A(n5020), .B(n5021), .Z(n5019) );
  OR U6147 ( .A(n5022), .B(n5023), .Z(n5020) );
  NANDN U6148 ( .A(n5024), .B(n5022), .Z(n5018) );
  XNOR U6149 ( .A(n4999), .B(n5025), .Z(N5905) );
  XOR U6150 ( .A(n5001), .B(n5002), .Z(n5025) );
  XNOR U6151 ( .A(n5015), .B(n5026), .Z(n5002) );
  XOR U6152 ( .A(n5016), .B(n5017), .Z(n5026) );
  XOR U6153 ( .A(n5022), .B(n5027), .Z(n5017) );
  XOR U6154 ( .A(n5021), .B(n5024), .Z(n5027) );
  IV U6155 ( .A(n5023), .Z(n5024) );
  NAND U6156 ( .A(n5028), .B(n5029), .Z(n5023) );
  OR U6157 ( .A(n5030), .B(n5031), .Z(n5029) );
  OR U6158 ( .A(n5032), .B(n5033), .Z(n5028) );
  NAND U6159 ( .A(n5034), .B(n5035), .Z(n5021) );
  OR U6160 ( .A(n5036), .B(n5037), .Z(n5035) );
  OR U6161 ( .A(n5038), .B(n5039), .Z(n5034) );
  NOR U6162 ( .A(n5040), .B(n5041), .Z(n5022) );
  ANDN U6163 ( .B(n5042), .A(n5043), .Z(n5016) );
  XNOR U6164 ( .A(n5009), .B(n5044), .Z(n5015) );
  XNOR U6165 ( .A(n5008), .B(n5010), .Z(n5044) );
  NAND U6166 ( .A(n5045), .B(n5046), .Z(n5010) );
  OR U6167 ( .A(n5047), .B(n5048), .Z(n5046) );
  OR U6168 ( .A(n5049), .B(n5050), .Z(n5045) );
  NAND U6169 ( .A(n5051), .B(n5052), .Z(n5008) );
  OR U6170 ( .A(n5053), .B(n5054), .Z(n5052) );
  OR U6171 ( .A(n5055), .B(n5056), .Z(n5051) );
  ANDN U6172 ( .B(n5057), .A(n5058), .Z(n5009) );
  IV U6173 ( .A(n5059), .Z(n5057) );
  ANDN U6174 ( .B(n5060), .A(n5061), .Z(n5001) );
  XOR U6175 ( .A(n4987), .B(n5062), .Z(n4999) );
  XOR U6176 ( .A(n4988), .B(n4989), .Z(n5062) );
  XOR U6177 ( .A(n4994), .B(n5063), .Z(n4989) );
  XOR U6178 ( .A(n4993), .B(n4996), .Z(n5063) );
  IV U6179 ( .A(n4995), .Z(n4996) );
  NAND U6180 ( .A(n5064), .B(n5065), .Z(n4995) );
  OR U6181 ( .A(n5066), .B(n5067), .Z(n5065) );
  OR U6182 ( .A(n5068), .B(n5069), .Z(n5064) );
  NAND U6183 ( .A(n5070), .B(n5071), .Z(n4993) );
  OR U6184 ( .A(n5072), .B(n5073), .Z(n5071) );
  OR U6185 ( .A(n5074), .B(n5075), .Z(n5070) );
  NOR U6186 ( .A(n5076), .B(n5077), .Z(n4994) );
  ANDN U6187 ( .B(n5078), .A(n5079), .Z(n4988) );
  IV U6188 ( .A(n5080), .Z(n5078) );
  XNOR U6189 ( .A(n4981), .B(n5081), .Z(n4987) );
  XNOR U6190 ( .A(n4980), .B(n4982), .Z(n5081) );
  NAND U6191 ( .A(n5082), .B(n5083), .Z(n4982) );
  OR U6192 ( .A(n5084), .B(n5085), .Z(n5083) );
  OR U6193 ( .A(n5086), .B(n5087), .Z(n5082) );
  NAND U6194 ( .A(n5088), .B(n5089), .Z(n4980) );
  OR U6195 ( .A(n5090), .B(n5091), .Z(n5089) );
  OR U6196 ( .A(n5092), .B(n5093), .Z(n5088) );
  ANDN U6197 ( .B(n5094), .A(n5095), .Z(n4981) );
  IV U6198 ( .A(n5096), .Z(n5094) );
  XNOR U6199 ( .A(n5061), .B(n5060), .Z(N5904) );
  XOR U6200 ( .A(n5080), .B(n5079), .Z(n5060) );
  XNOR U6201 ( .A(n5095), .B(n5096), .Z(n5079) );
  XNOR U6202 ( .A(n5090), .B(n5091), .Z(n5096) );
  XNOR U6203 ( .A(n5092), .B(n5093), .Z(n5091) );
  XNOR U6204 ( .A(y[292]), .B(x[292]), .Z(n5093) );
  XNOR U6205 ( .A(y[293]), .B(x[293]), .Z(n5092) );
  XNOR U6206 ( .A(y[291]), .B(x[291]), .Z(n5090) );
  XNOR U6207 ( .A(n5084), .B(n5085), .Z(n5095) );
  XNOR U6208 ( .A(y[288]), .B(x[288]), .Z(n5085) );
  XNOR U6209 ( .A(n5086), .B(n5087), .Z(n5084) );
  XNOR U6210 ( .A(y[289]), .B(x[289]), .Z(n5087) );
  XNOR U6211 ( .A(y[290]), .B(x[290]), .Z(n5086) );
  XNOR U6212 ( .A(n5077), .B(n5076), .Z(n5080) );
  XNOR U6213 ( .A(n5072), .B(n5073), .Z(n5076) );
  XNOR U6214 ( .A(y[285]), .B(x[285]), .Z(n5073) );
  XNOR U6215 ( .A(n5074), .B(n5075), .Z(n5072) );
  XNOR U6216 ( .A(y[286]), .B(x[286]), .Z(n5075) );
  XNOR U6217 ( .A(y[287]), .B(x[287]), .Z(n5074) );
  XNOR U6218 ( .A(n5066), .B(n5067), .Z(n5077) );
  XNOR U6219 ( .A(y[282]), .B(x[282]), .Z(n5067) );
  XNOR U6220 ( .A(n5068), .B(n5069), .Z(n5066) );
  XNOR U6221 ( .A(y[283]), .B(x[283]), .Z(n5069) );
  XNOR U6222 ( .A(y[284]), .B(x[284]), .Z(n5068) );
  XOR U6223 ( .A(n5042), .B(n5043), .Z(n5061) );
  XNOR U6224 ( .A(n5058), .B(n5059), .Z(n5043) );
  XNOR U6225 ( .A(n5053), .B(n5054), .Z(n5059) );
  XNOR U6226 ( .A(n5055), .B(n5056), .Z(n5054) );
  XNOR U6227 ( .A(y[280]), .B(x[280]), .Z(n5056) );
  XNOR U6228 ( .A(y[281]), .B(x[281]), .Z(n5055) );
  XNOR U6229 ( .A(y[279]), .B(x[279]), .Z(n5053) );
  XNOR U6230 ( .A(n5047), .B(n5048), .Z(n5058) );
  XNOR U6231 ( .A(y[276]), .B(x[276]), .Z(n5048) );
  XNOR U6232 ( .A(n5049), .B(n5050), .Z(n5047) );
  XNOR U6233 ( .A(y[277]), .B(x[277]), .Z(n5050) );
  XNOR U6234 ( .A(y[278]), .B(x[278]), .Z(n5049) );
  XOR U6235 ( .A(n5041), .B(n5040), .Z(n5042) );
  XNOR U6236 ( .A(n5036), .B(n5037), .Z(n5040) );
  XNOR U6237 ( .A(y[273]), .B(x[273]), .Z(n5037) );
  XNOR U6238 ( .A(n5038), .B(n5039), .Z(n5036) );
  XNOR U6239 ( .A(y[274]), .B(x[274]), .Z(n5039) );
  XNOR U6240 ( .A(y[275]), .B(x[275]), .Z(n5038) );
  XNOR U6241 ( .A(n5030), .B(n5031), .Z(n5041) );
  XNOR U6242 ( .A(y[270]), .B(x[270]), .Z(n5031) );
  XNOR U6243 ( .A(n5032), .B(n5033), .Z(n5030) );
  XNOR U6244 ( .A(y[271]), .B(x[271]), .Z(n5033) );
  XNOR U6245 ( .A(y[272]), .B(x[272]), .Z(n5032) );
  NAND U6246 ( .A(n5097), .B(n5098), .Z(N5898) );
  NANDN U6247 ( .A(n5099), .B(n5100), .Z(n5098) );
  OR U6248 ( .A(n5101), .B(n5102), .Z(n5100) );
  NAND U6249 ( .A(n5101), .B(n5102), .Z(n5097) );
  XOR U6250 ( .A(n5101), .B(n5103), .Z(N5897) );
  XNOR U6251 ( .A(n5099), .B(n5102), .Z(n5103) );
  AND U6252 ( .A(n5104), .B(n5105), .Z(n5102) );
  NANDN U6253 ( .A(n5106), .B(n5107), .Z(n5105) );
  NANDN U6254 ( .A(n5108), .B(n5109), .Z(n5107) );
  NANDN U6255 ( .A(n5109), .B(n5108), .Z(n5104) );
  NAND U6256 ( .A(n5110), .B(n5111), .Z(n5099) );
  NANDN U6257 ( .A(n5112), .B(n5113), .Z(n5111) );
  OR U6258 ( .A(n5114), .B(n5115), .Z(n5113) );
  NAND U6259 ( .A(n5115), .B(n5114), .Z(n5110) );
  AND U6260 ( .A(n5116), .B(n5117), .Z(n5101) );
  NANDN U6261 ( .A(n5118), .B(n5119), .Z(n5117) );
  NANDN U6262 ( .A(n5120), .B(n5121), .Z(n5119) );
  NANDN U6263 ( .A(n5121), .B(n5120), .Z(n5116) );
  XOR U6264 ( .A(n5115), .B(n5122), .Z(N5896) );
  XOR U6265 ( .A(n5112), .B(n5114), .Z(n5122) );
  XNOR U6266 ( .A(n5108), .B(n5123), .Z(n5114) );
  XNOR U6267 ( .A(n5106), .B(n5109), .Z(n5123) );
  NAND U6268 ( .A(n5124), .B(n5125), .Z(n5109) );
  NAND U6269 ( .A(n5126), .B(n5127), .Z(n5125) );
  OR U6270 ( .A(n5128), .B(n5129), .Z(n5126) );
  NANDN U6271 ( .A(n5130), .B(n5128), .Z(n5124) );
  IV U6272 ( .A(n5129), .Z(n5130) );
  NAND U6273 ( .A(n5131), .B(n5132), .Z(n5106) );
  NAND U6274 ( .A(n5133), .B(n5134), .Z(n5132) );
  NANDN U6275 ( .A(n5135), .B(n5136), .Z(n5133) );
  NANDN U6276 ( .A(n5136), .B(n5135), .Z(n5131) );
  AND U6277 ( .A(n5137), .B(n5138), .Z(n5108) );
  NAND U6278 ( .A(n5139), .B(n5140), .Z(n5138) );
  OR U6279 ( .A(n5141), .B(n5142), .Z(n5139) );
  NANDN U6280 ( .A(n5143), .B(n5141), .Z(n5137) );
  NAND U6281 ( .A(n5144), .B(n5145), .Z(n5112) );
  NANDN U6282 ( .A(n5146), .B(n5147), .Z(n5145) );
  OR U6283 ( .A(n5148), .B(n5149), .Z(n5147) );
  NANDN U6284 ( .A(n5150), .B(n5148), .Z(n5144) );
  IV U6285 ( .A(n5149), .Z(n5150) );
  XNOR U6286 ( .A(n5120), .B(n5151), .Z(n5115) );
  XNOR U6287 ( .A(n5118), .B(n5121), .Z(n5151) );
  NAND U6288 ( .A(n5152), .B(n5153), .Z(n5121) );
  NAND U6289 ( .A(n5154), .B(n5155), .Z(n5153) );
  OR U6290 ( .A(n5156), .B(n5157), .Z(n5154) );
  NANDN U6291 ( .A(n5158), .B(n5156), .Z(n5152) );
  IV U6292 ( .A(n5157), .Z(n5158) );
  NAND U6293 ( .A(n5159), .B(n5160), .Z(n5118) );
  NAND U6294 ( .A(n5161), .B(n5162), .Z(n5160) );
  NANDN U6295 ( .A(n5163), .B(n5164), .Z(n5161) );
  NANDN U6296 ( .A(n5164), .B(n5163), .Z(n5159) );
  AND U6297 ( .A(n5165), .B(n5166), .Z(n5120) );
  NAND U6298 ( .A(n5167), .B(n5168), .Z(n5166) );
  OR U6299 ( .A(n5169), .B(n5170), .Z(n5167) );
  NANDN U6300 ( .A(n5171), .B(n5169), .Z(n5165) );
  XNOR U6301 ( .A(n5146), .B(n5172), .Z(N5895) );
  XOR U6302 ( .A(n5148), .B(n5149), .Z(n5172) );
  XNOR U6303 ( .A(n5162), .B(n5173), .Z(n5149) );
  XOR U6304 ( .A(n5163), .B(n5164), .Z(n5173) );
  XOR U6305 ( .A(n5169), .B(n5174), .Z(n5164) );
  XOR U6306 ( .A(n5168), .B(n5171), .Z(n5174) );
  IV U6307 ( .A(n5170), .Z(n5171) );
  NAND U6308 ( .A(n5175), .B(n5176), .Z(n5170) );
  OR U6309 ( .A(n5177), .B(n5178), .Z(n5176) );
  OR U6310 ( .A(n5179), .B(n5180), .Z(n5175) );
  NAND U6311 ( .A(n5181), .B(n5182), .Z(n5168) );
  OR U6312 ( .A(n5183), .B(n5184), .Z(n5182) );
  OR U6313 ( .A(n5185), .B(n5186), .Z(n5181) );
  NOR U6314 ( .A(n5187), .B(n5188), .Z(n5169) );
  ANDN U6315 ( .B(n5189), .A(n5190), .Z(n5163) );
  XNOR U6316 ( .A(n5156), .B(n5191), .Z(n5162) );
  XNOR U6317 ( .A(n5155), .B(n5157), .Z(n5191) );
  NAND U6318 ( .A(n5192), .B(n5193), .Z(n5157) );
  OR U6319 ( .A(n5194), .B(n5195), .Z(n5193) );
  OR U6320 ( .A(n5196), .B(n5197), .Z(n5192) );
  NAND U6321 ( .A(n5198), .B(n5199), .Z(n5155) );
  OR U6322 ( .A(n5200), .B(n5201), .Z(n5199) );
  OR U6323 ( .A(n5202), .B(n5203), .Z(n5198) );
  ANDN U6324 ( .B(n5204), .A(n5205), .Z(n5156) );
  IV U6325 ( .A(n5206), .Z(n5204) );
  ANDN U6326 ( .B(n5207), .A(n5208), .Z(n5148) );
  XOR U6327 ( .A(n5134), .B(n5209), .Z(n5146) );
  XOR U6328 ( .A(n5135), .B(n5136), .Z(n5209) );
  XOR U6329 ( .A(n5141), .B(n5210), .Z(n5136) );
  XOR U6330 ( .A(n5140), .B(n5143), .Z(n5210) );
  IV U6331 ( .A(n5142), .Z(n5143) );
  NAND U6332 ( .A(n5211), .B(n5212), .Z(n5142) );
  OR U6333 ( .A(n5213), .B(n5214), .Z(n5212) );
  OR U6334 ( .A(n5215), .B(n5216), .Z(n5211) );
  NAND U6335 ( .A(n5217), .B(n5218), .Z(n5140) );
  OR U6336 ( .A(n5219), .B(n5220), .Z(n5218) );
  OR U6337 ( .A(n5221), .B(n5222), .Z(n5217) );
  NOR U6338 ( .A(n5223), .B(n5224), .Z(n5141) );
  ANDN U6339 ( .B(n5225), .A(n5226), .Z(n5135) );
  IV U6340 ( .A(n5227), .Z(n5225) );
  XNOR U6341 ( .A(n5128), .B(n5228), .Z(n5134) );
  XNOR U6342 ( .A(n5127), .B(n5129), .Z(n5228) );
  NAND U6343 ( .A(n5229), .B(n5230), .Z(n5129) );
  OR U6344 ( .A(n5231), .B(n5232), .Z(n5230) );
  OR U6345 ( .A(n5233), .B(n5234), .Z(n5229) );
  NAND U6346 ( .A(n5235), .B(n5236), .Z(n5127) );
  OR U6347 ( .A(n5237), .B(n5238), .Z(n5236) );
  OR U6348 ( .A(n5239), .B(n5240), .Z(n5235) );
  ANDN U6349 ( .B(n5241), .A(n5242), .Z(n5128) );
  IV U6350 ( .A(n5243), .Z(n5241) );
  XNOR U6351 ( .A(n5208), .B(n5207), .Z(N5894) );
  XOR U6352 ( .A(n5227), .B(n5226), .Z(n5207) );
  XNOR U6353 ( .A(n5242), .B(n5243), .Z(n5226) );
  XNOR U6354 ( .A(n5237), .B(n5238), .Z(n5243) );
  XNOR U6355 ( .A(n5239), .B(n5240), .Z(n5238) );
  XNOR U6356 ( .A(y[268]), .B(x[268]), .Z(n5240) );
  XNOR U6357 ( .A(y[269]), .B(x[269]), .Z(n5239) );
  XNOR U6358 ( .A(y[267]), .B(x[267]), .Z(n5237) );
  XNOR U6359 ( .A(n5231), .B(n5232), .Z(n5242) );
  XNOR U6360 ( .A(y[264]), .B(x[264]), .Z(n5232) );
  XNOR U6361 ( .A(n5233), .B(n5234), .Z(n5231) );
  XNOR U6362 ( .A(y[265]), .B(x[265]), .Z(n5234) );
  XNOR U6363 ( .A(y[266]), .B(x[266]), .Z(n5233) );
  XNOR U6364 ( .A(n5224), .B(n5223), .Z(n5227) );
  XNOR U6365 ( .A(n5219), .B(n5220), .Z(n5223) );
  XNOR U6366 ( .A(y[261]), .B(x[261]), .Z(n5220) );
  XNOR U6367 ( .A(n5221), .B(n5222), .Z(n5219) );
  XNOR U6368 ( .A(y[262]), .B(x[262]), .Z(n5222) );
  XNOR U6369 ( .A(y[263]), .B(x[263]), .Z(n5221) );
  XNOR U6370 ( .A(n5213), .B(n5214), .Z(n5224) );
  XNOR U6371 ( .A(y[258]), .B(x[258]), .Z(n5214) );
  XNOR U6372 ( .A(n5215), .B(n5216), .Z(n5213) );
  XNOR U6373 ( .A(y[259]), .B(x[259]), .Z(n5216) );
  XNOR U6374 ( .A(y[260]), .B(x[260]), .Z(n5215) );
  XOR U6375 ( .A(n5189), .B(n5190), .Z(n5208) );
  XNOR U6376 ( .A(n5205), .B(n5206), .Z(n5190) );
  XNOR U6377 ( .A(n5200), .B(n5201), .Z(n5206) );
  XNOR U6378 ( .A(n5202), .B(n5203), .Z(n5201) );
  XNOR U6379 ( .A(y[256]), .B(x[256]), .Z(n5203) );
  XNOR U6380 ( .A(y[257]), .B(x[257]), .Z(n5202) );
  XNOR U6381 ( .A(y[255]), .B(x[255]), .Z(n5200) );
  XNOR U6382 ( .A(n5194), .B(n5195), .Z(n5205) );
  XNOR U6383 ( .A(y[252]), .B(x[252]), .Z(n5195) );
  XNOR U6384 ( .A(n5196), .B(n5197), .Z(n5194) );
  XNOR U6385 ( .A(y[253]), .B(x[253]), .Z(n5197) );
  XNOR U6386 ( .A(y[254]), .B(x[254]), .Z(n5196) );
  XOR U6387 ( .A(n5188), .B(n5187), .Z(n5189) );
  XNOR U6388 ( .A(n5183), .B(n5184), .Z(n5187) );
  XNOR U6389 ( .A(y[249]), .B(x[249]), .Z(n5184) );
  XNOR U6390 ( .A(n5185), .B(n5186), .Z(n5183) );
  XNOR U6391 ( .A(y[250]), .B(x[250]), .Z(n5186) );
  XNOR U6392 ( .A(y[251]), .B(x[251]), .Z(n5185) );
  XNOR U6393 ( .A(n5177), .B(n5178), .Z(n5188) );
  XNOR U6394 ( .A(y[246]), .B(x[246]), .Z(n5178) );
  XNOR U6395 ( .A(n5179), .B(n5180), .Z(n5177) );
  XNOR U6396 ( .A(y[247]), .B(x[247]), .Z(n5180) );
  XNOR U6397 ( .A(y[248]), .B(x[248]), .Z(n5179) );
  NAND U6398 ( .A(n5244), .B(n5245), .Z(N5888) );
  NANDN U6399 ( .A(n5246), .B(n5247), .Z(n5245) );
  OR U6400 ( .A(n5248), .B(n5249), .Z(n5247) );
  NAND U6401 ( .A(n5248), .B(n5249), .Z(n5244) );
  XOR U6402 ( .A(n5248), .B(n5250), .Z(N5887) );
  XNOR U6403 ( .A(n5246), .B(n5249), .Z(n5250) );
  AND U6404 ( .A(n5251), .B(n5252), .Z(n5249) );
  NANDN U6405 ( .A(n5253), .B(n5254), .Z(n5252) );
  NANDN U6406 ( .A(n5255), .B(n5256), .Z(n5254) );
  NANDN U6407 ( .A(n5256), .B(n5255), .Z(n5251) );
  NAND U6408 ( .A(n5257), .B(n5258), .Z(n5246) );
  NANDN U6409 ( .A(n5259), .B(n5260), .Z(n5258) );
  OR U6410 ( .A(n5261), .B(n5262), .Z(n5260) );
  NAND U6411 ( .A(n5262), .B(n5261), .Z(n5257) );
  AND U6412 ( .A(n5263), .B(n5264), .Z(n5248) );
  NANDN U6413 ( .A(n5265), .B(n5266), .Z(n5264) );
  NANDN U6414 ( .A(n5267), .B(n5268), .Z(n5266) );
  NANDN U6415 ( .A(n5268), .B(n5267), .Z(n5263) );
  XOR U6416 ( .A(n5262), .B(n5269), .Z(N5886) );
  XOR U6417 ( .A(n5259), .B(n5261), .Z(n5269) );
  XNOR U6418 ( .A(n5255), .B(n5270), .Z(n5261) );
  XNOR U6419 ( .A(n5253), .B(n5256), .Z(n5270) );
  NAND U6420 ( .A(n5271), .B(n5272), .Z(n5256) );
  NAND U6421 ( .A(n5273), .B(n5274), .Z(n5272) );
  OR U6422 ( .A(n5275), .B(n5276), .Z(n5273) );
  NANDN U6423 ( .A(n5277), .B(n5275), .Z(n5271) );
  IV U6424 ( .A(n5276), .Z(n5277) );
  NAND U6425 ( .A(n5278), .B(n5279), .Z(n5253) );
  NAND U6426 ( .A(n5280), .B(n5281), .Z(n5279) );
  NANDN U6427 ( .A(n5282), .B(n5283), .Z(n5280) );
  NANDN U6428 ( .A(n5283), .B(n5282), .Z(n5278) );
  AND U6429 ( .A(n5284), .B(n5285), .Z(n5255) );
  NAND U6430 ( .A(n5286), .B(n5287), .Z(n5285) );
  OR U6431 ( .A(n5288), .B(n5289), .Z(n5286) );
  NANDN U6432 ( .A(n5290), .B(n5288), .Z(n5284) );
  NAND U6433 ( .A(n5291), .B(n5292), .Z(n5259) );
  NANDN U6434 ( .A(n5293), .B(n5294), .Z(n5292) );
  OR U6435 ( .A(n5295), .B(n5296), .Z(n5294) );
  NANDN U6436 ( .A(n5297), .B(n5295), .Z(n5291) );
  IV U6437 ( .A(n5296), .Z(n5297) );
  XNOR U6438 ( .A(n5267), .B(n5298), .Z(n5262) );
  XNOR U6439 ( .A(n5265), .B(n5268), .Z(n5298) );
  NAND U6440 ( .A(n5299), .B(n5300), .Z(n5268) );
  NAND U6441 ( .A(n5301), .B(n5302), .Z(n5300) );
  OR U6442 ( .A(n5303), .B(n5304), .Z(n5301) );
  NANDN U6443 ( .A(n5305), .B(n5303), .Z(n5299) );
  IV U6444 ( .A(n5304), .Z(n5305) );
  NAND U6445 ( .A(n5306), .B(n5307), .Z(n5265) );
  NAND U6446 ( .A(n5308), .B(n5309), .Z(n5307) );
  NANDN U6447 ( .A(n5310), .B(n5311), .Z(n5308) );
  NANDN U6448 ( .A(n5311), .B(n5310), .Z(n5306) );
  AND U6449 ( .A(n5312), .B(n5313), .Z(n5267) );
  NAND U6450 ( .A(n5314), .B(n5315), .Z(n5313) );
  OR U6451 ( .A(n5316), .B(n5317), .Z(n5314) );
  NANDN U6452 ( .A(n5318), .B(n5316), .Z(n5312) );
  XNOR U6453 ( .A(n5293), .B(n5319), .Z(N5885) );
  XOR U6454 ( .A(n5295), .B(n5296), .Z(n5319) );
  XNOR U6455 ( .A(n5309), .B(n5320), .Z(n5296) );
  XOR U6456 ( .A(n5310), .B(n5311), .Z(n5320) );
  XOR U6457 ( .A(n5316), .B(n5321), .Z(n5311) );
  XOR U6458 ( .A(n5315), .B(n5318), .Z(n5321) );
  IV U6459 ( .A(n5317), .Z(n5318) );
  NAND U6460 ( .A(n5322), .B(n5323), .Z(n5317) );
  OR U6461 ( .A(n5324), .B(n5325), .Z(n5323) );
  OR U6462 ( .A(n5326), .B(n5327), .Z(n5322) );
  NAND U6463 ( .A(n5328), .B(n5329), .Z(n5315) );
  OR U6464 ( .A(n5330), .B(n5331), .Z(n5329) );
  OR U6465 ( .A(n5332), .B(n5333), .Z(n5328) );
  NOR U6466 ( .A(n5334), .B(n5335), .Z(n5316) );
  ANDN U6467 ( .B(n5336), .A(n5337), .Z(n5310) );
  XNOR U6468 ( .A(n5303), .B(n5338), .Z(n5309) );
  XNOR U6469 ( .A(n5302), .B(n5304), .Z(n5338) );
  NAND U6470 ( .A(n5339), .B(n5340), .Z(n5304) );
  OR U6471 ( .A(n5341), .B(n5342), .Z(n5340) );
  OR U6472 ( .A(n5343), .B(n5344), .Z(n5339) );
  NAND U6473 ( .A(n5345), .B(n5346), .Z(n5302) );
  OR U6474 ( .A(n5347), .B(n5348), .Z(n5346) );
  OR U6475 ( .A(n5349), .B(n5350), .Z(n5345) );
  ANDN U6476 ( .B(n5351), .A(n5352), .Z(n5303) );
  IV U6477 ( .A(n5353), .Z(n5351) );
  ANDN U6478 ( .B(n5354), .A(n5355), .Z(n5295) );
  XOR U6479 ( .A(n5281), .B(n5356), .Z(n5293) );
  XOR U6480 ( .A(n5282), .B(n5283), .Z(n5356) );
  XOR U6481 ( .A(n5288), .B(n5357), .Z(n5283) );
  XOR U6482 ( .A(n5287), .B(n5290), .Z(n5357) );
  IV U6483 ( .A(n5289), .Z(n5290) );
  NAND U6484 ( .A(n5358), .B(n5359), .Z(n5289) );
  OR U6485 ( .A(n5360), .B(n5361), .Z(n5359) );
  OR U6486 ( .A(n5362), .B(n5363), .Z(n5358) );
  NAND U6487 ( .A(n5364), .B(n5365), .Z(n5287) );
  OR U6488 ( .A(n5366), .B(n5367), .Z(n5365) );
  OR U6489 ( .A(n5368), .B(n5369), .Z(n5364) );
  NOR U6490 ( .A(n5370), .B(n5371), .Z(n5288) );
  ANDN U6491 ( .B(n5372), .A(n5373), .Z(n5282) );
  IV U6492 ( .A(n5374), .Z(n5372) );
  XNOR U6493 ( .A(n5275), .B(n5375), .Z(n5281) );
  XNOR U6494 ( .A(n5274), .B(n5276), .Z(n5375) );
  NAND U6495 ( .A(n5376), .B(n5377), .Z(n5276) );
  OR U6496 ( .A(n5378), .B(n5379), .Z(n5377) );
  OR U6497 ( .A(n5380), .B(n5381), .Z(n5376) );
  NAND U6498 ( .A(n5382), .B(n5383), .Z(n5274) );
  OR U6499 ( .A(n5384), .B(n5385), .Z(n5383) );
  OR U6500 ( .A(n5386), .B(n5387), .Z(n5382) );
  ANDN U6501 ( .B(n5388), .A(n5389), .Z(n5275) );
  IV U6502 ( .A(n5390), .Z(n5388) );
  XNOR U6503 ( .A(n5355), .B(n5354), .Z(N5884) );
  XOR U6504 ( .A(n5374), .B(n5373), .Z(n5354) );
  XNOR U6505 ( .A(n5389), .B(n5390), .Z(n5373) );
  XNOR U6506 ( .A(n5384), .B(n5385), .Z(n5390) );
  XNOR U6507 ( .A(n5386), .B(n5387), .Z(n5385) );
  XNOR U6508 ( .A(y[244]), .B(x[244]), .Z(n5387) );
  XNOR U6509 ( .A(y[245]), .B(x[245]), .Z(n5386) );
  XNOR U6510 ( .A(y[243]), .B(x[243]), .Z(n5384) );
  XNOR U6511 ( .A(n5378), .B(n5379), .Z(n5389) );
  XNOR U6512 ( .A(y[240]), .B(x[240]), .Z(n5379) );
  XNOR U6513 ( .A(n5380), .B(n5381), .Z(n5378) );
  XNOR U6514 ( .A(y[241]), .B(x[241]), .Z(n5381) );
  XNOR U6515 ( .A(y[242]), .B(x[242]), .Z(n5380) );
  XNOR U6516 ( .A(n5371), .B(n5370), .Z(n5374) );
  XNOR U6517 ( .A(n5366), .B(n5367), .Z(n5370) );
  XNOR U6518 ( .A(y[237]), .B(x[237]), .Z(n5367) );
  XNOR U6519 ( .A(n5368), .B(n5369), .Z(n5366) );
  XNOR U6520 ( .A(y[238]), .B(x[238]), .Z(n5369) );
  XNOR U6521 ( .A(y[239]), .B(x[239]), .Z(n5368) );
  XNOR U6522 ( .A(n5360), .B(n5361), .Z(n5371) );
  XNOR U6523 ( .A(y[234]), .B(x[234]), .Z(n5361) );
  XNOR U6524 ( .A(n5362), .B(n5363), .Z(n5360) );
  XNOR U6525 ( .A(y[235]), .B(x[235]), .Z(n5363) );
  XNOR U6526 ( .A(y[236]), .B(x[236]), .Z(n5362) );
  XOR U6527 ( .A(n5336), .B(n5337), .Z(n5355) );
  XNOR U6528 ( .A(n5352), .B(n5353), .Z(n5337) );
  XNOR U6529 ( .A(n5347), .B(n5348), .Z(n5353) );
  XNOR U6530 ( .A(n5349), .B(n5350), .Z(n5348) );
  XNOR U6531 ( .A(y[232]), .B(x[232]), .Z(n5350) );
  XNOR U6532 ( .A(y[233]), .B(x[233]), .Z(n5349) );
  XNOR U6533 ( .A(y[231]), .B(x[231]), .Z(n5347) );
  XNOR U6534 ( .A(n5341), .B(n5342), .Z(n5352) );
  XNOR U6535 ( .A(y[228]), .B(x[228]), .Z(n5342) );
  XNOR U6536 ( .A(n5343), .B(n5344), .Z(n5341) );
  XNOR U6537 ( .A(y[229]), .B(x[229]), .Z(n5344) );
  XNOR U6538 ( .A(y[230]), .B(x[230]), .Z(n5343) );
  XOR U6539 ( .A(n5335), .B(n5334), .Z(n5336) );
  XNOR U6540 ( .A(n5330), .B(n5331), .Z(n5334) );
  XNOR U6541 ( .A(y[225]), .B(x[225]), .Z(n5331) );
  XNOR U6542 ( .A(n5332), .B(n5333), .Z(n5330) );
  XNOR U6543 ( .A(y[226]), .B(x[226]), .Z(n5333) );
  XNOR U6544 ( .A(y[227]), .B(x[227]), .Z(n5332) );
  XNOR U6545 ( .A(n5324), .B(n5325), .Z(n5335) );
  XNOR U6546 ( .A(y[222]), .B(x[222]), .Z(n5325) );
  XNOR U6547 ( .A(n5326), .B(n5327), .Z(n5324) );
  XNOR U6548 ( .A(y[223]), .B(x[223]), .Z(n5327) );
  XNOR U6549 ( .A(y[224]), .B(x[224]), .Z(n5326) );
  NAND U6550 ( .A(n5391), .B(n5392), .Z(N5878) );
  NANDN U6551 ( .A(n5393), .B(n5394), .Z(n5392) );
  OR U6552 ( .A(n5395), .B(n5396), .Z(n5394) );
  NAND U6553 ( .A(n5395), .B(n5396), .Z(n5391) );
  XOR U6554 ( .A(n5395), .B(n5397), .Z(N5877) );
  XNOR U6555 ( .A(n5393), .B(n5396), .Z(n5397) );
  AND U6556 ( .A(n5398), .B(n5399), .Z(n5396) );
  NANDN U6557 ( .A(n5400), .B(n5401), .Z(n5399) );
  NANDN U6558 ( .A(n5402), .B(n5403), .Z(n5401) );
  NANDN U6559 ( .A(n5403), .B(n5402), .Z(n5398) );
  NAND U6560 ( .A(n5404), .B(n5405), .Z(n5393) );
  NANDN U6561 ( .A(n5406), .B(n5407), .Z(n5405) );
  OR U6562 ( .A(n5408), .B(n5409), .Z(n5407) );
  NAND U6563 ( .A(n5409), .B(n5408), .Z(n5404) );
  AND U6564 ( .A(n5410), .B(n5411), .Z(n5395) );
  NANDN U6565 ( .A(n5412), .B(n5413), .Z(n5411) );
  NANDN U6566 ( .A(n5414), .B(n5415), .Z(n5413) );
  NANDN U6567 ( .A(n5415), .B(n5414), .Z(n5410) );
  XOR U6568 ( .A(n5409), .B(n5416), .Z(N5876) );
  XOR U6569 ( .A(n5406), .B(n5408), .Z(n5416) );
  XNOR U6570 ( .A(n5402), .B(n5417), .Z(n5408) );
  XNOR U6571 ( .A(n5400), .B(n5403), .Z(n5417) );
  NAND U6572 ( .A(n5418), .B(n5419), .Z(n5403) );
  NAND U6573 ( .A(n5420), .B(n5421), .Z(n5419) );
  OR U6574 ( .A(n5422), .B(n5423), .Z(n5420) );
  NANDN U6575 ( .A(n5424), .B(n5422), .Z(n5418) );
  IV U6576 ( .A(n5423), .Z(n5424) );
  NAND U6577 ( .A(n5425), .B(n5426), .Z(n5400) );
  NAND U6578 ( .A(n5427), .B(n5428), .Z(n5426) );
  NANDN U6579 ( .A(n5429), .B(n5430), .Z(n5427) );
  NANDN U6580 ( .A(n5430), .B(n5429), .Z(n5425) );
  AND U6581 ( .A(n5431), .B(n5432), .Z(n5402) );
  NAND U6582 ( .A(n5433), .B(n5434), .Z(n5432) );
  OR U6583 ( .A(n5435), .B(n5436), .Z(n5433) );
  NANDN U6584 ( .A(n5437), .B(n5435), .Z(n5431) );
  NAND U6585 ( .A(n5438), .B(n5439), .Z(n5406) );
  NANDN U6586 ( .A(n5440), .B(n5441), .Z(n5439) );
  OR U6587 ( .A(n5442), .B(n5443), .Z(n5441) );
  NANDN U6588 ( .A(n5444), .B(n5442), .Z(n5438) );
  IV U6589 ( .A(n5443), .Z(n5444) );
  XNOR U6590 ( .A(n5414), .B(n5445), .Z(n5409) );
  XNOR U6591 ( .A(n5412), .B(n5415), .Z(n5445) );
  NAND U6592 ( .A(n5446), .B(n5447), .Z(n5415) );
  NAND U6593 ( .A(n5448), .B(n5449), .Z(n5447) );
  OR U6594 ( .A(n5450), .B(n5451), .Z(n5448) );
  NANDN U6595 ( .A(n5452), .B(n5450), .Z(n5446) );
  IV U6596 ( .A(n5451), .Z(n5452) );
  NAND U6597 ( .A(n5453), .B(n5454), .Z(n5412) );
  NAND U6598 ( .A(n5455), .B(n5456), .Z(n5454) );
  NANDN U6599 ( .A(n5457), .B(n5458), .Z(n5455) );
  NANDN U6600 ( .A(n5458), .B(n5457), .Z(n5453) );
  AND U6601 ( .A(n5459), .B(n5460), .Z(n5414) );
  NAND U6602 ( .A(n5461), .B(n5462), .Z(n5460) );
  OR U6603 ( .A(n5463), .B(n5464), .Z(n5461) );
  NANDN U6604 ( .A(n5465), .B(n5463), .Z(n5459) );
  XNOR U6605 ( .A(n5440), .B(n5466), .Z(N5875) );
  XOR U6606 ( .A(n5442), .B(n5443), .Z(n5466) );
  XNOR U6607 ( .A(n5456), .B(n5467), .Z(n5443) );
  XOR U6608 ( .A(n5457), .B(n5458), .Z(n5467) );
  XOR U6609 ( .A(n5463), .B(n5468), .Z(n5458) );
  XOR U6610 ( .A(n5462), .B(n5465), .Z(n5468) );
  IV U6611 ( .A(n5464), .Z(n5465) );
  NAND U6612 ( .A(n5469), .B(n5470), .Z(n5464) );
  OR U6613 ( .A(n5471), .B(n5472), .Z(n5470) );
  OR U6614 ( .A(n5473), .B(n5474), .Z(n5469) );
  NAND U6615 ( .A(n5475), .B(n5476), .Z(n5462) );
  OR U6616 ( .A(n5477), .B(n5478), .Z(n5476) );
  OR U6617 ( .A(n5479), .B(n5480), .Z(n5475) );
  NOR U6618 ( .A(n5481), .B(n5482), .Z(n5463) );
  ANDN U6619 ( .B(n5483), .A(n5484), .Z(n5457) );
  XNOR U6620 ( .A(n5450), .B(n5485), .Z(n5456) );
  XNOR U6621 ( .A(n5449), .B(n5451), .Z(n5485) );
  NAND U6622 ( .A(n5486), .B(n5487), .Z(n5451) );
  OR U6623 ( .A(n5488), .B(n5489), .Z(n5487) );
  OR U6624 ( .A(n5490), .B(n5491), .Z(n5486) );
  NAND U6625 ( .A(n5492), .B(n5493), .Z(n5449) );
  OR U6626 ( .A(n5494), .B(n5495), .Z(n5493) );
  OR U6627 ( .A(n5496), .B(n5497), .Z(n5492) );
  ANDN U6628 ( .B(n5498), .A(n5499), .Z(n5450) );
  IV U6629 ( .A(n5500), .Z(n5498) );
  ANDN U6630 ( .B(n5501), .A(n5502), .Z(n5442) );
  XOR U6631 ( .A(n5428), .B(n5503), .Z(n5440) );
  XOR U6632 ( .A(n5429), .B(n5430), .Z(n5503) );
  XOR U6633 ( .A(n5435), .B(n5504), .Z(n5430) );
  XOR U6634 ( .A(n5434), .B(n5437), .Z(n5504) );
  IV U6635 ( .A(n5436), .Z(n5437) );
  NAND U6636 ( .A(n5505), .B(n5506), .Z(n5436) );
  OR U6637 ( .A(n5507), .B(n5508), .Z(n5506) );
  OR U6638 ( .A(n5509), .B(n5510), .Z(n5505) );
  NAND U6639 ( .A(n5511), .B(n5512), .Z(n5434) );
  OR U6640 ( .A(n5513), .B(n5514), .Z(n5512) );
  OR U6641 ( .A(n5515), .B(n5516), .Z(n5511) );
  NOR U6642 ( .A(n5517), .B(n5518), .Z(n5435) );
  ANDN U6643 ( .B(n5519), .A(n5520), .Z(n5429) );
  IV U6644 ( .A(n5521), .Z(n5519) );
  XNOR U6645 ( .A(n5422), .B(n5522), .Z(n5428) );
  XNOR U6646 ( .A(n5421), .B(n5423), .Z(n5522) );
  NAND U6647 ( .A(n5523), .B(n5524), .Z(n5423) );
  OR U6648 ( .A(n5525), .B(n5526), .Z(n5524) );
  OR U6649 ( .A(n5527), .B(n5528), .Z(n5523) );
  NAND U6650 ( .A(n5529), .B(n5530), .Z(n5421) );
  OR U6651 ( .A(n5531), .B(n5532), .Z(n5530) );
  OR U6652 ( .A(n5533), .B(n5534), .Z(n5529) );
  ANDN U6653 ( .B(n5535), .A(n5536), .Z(n5422) );
  IV U6654 ( .A(n5537), .Z(n5535) );
  XNOR U6655 ( .A(n5502), .B(n5501), .Z(N5874) );
  XOR U6656 ( .A(n5521), .B(n5520), .Z(n5501) );
  XNOR U6657 ( .A(n5536), .B(n5537), .Z(n5520) );
  XNOR U6658 ( .A(n5531), .B(n5532), .Z(n5537) );
  XNOR U6659 ( .A(n5533), .B(n5534), .Z(n5532) );
  XNOR U6660 ( .A(y[220]), .B(x[220]), .Z(n5534) );
  XNOR U6661 ( .A(y[221]), .B(x[221]), .Z(n5533) );
  XNOR U6662 ( .A(y[219]), .B(x[219]), .Z(n5531) );
  XNOR U6663 ( .A(n5525), .B(n5526), .Z(n5536) );
  XNOR U6664 ( .A(y[216]), .B(x[216]), .Z(n5526) );
  XNOR U6665 ( .A(n5527), .B(n5528), .Z(n5525) );
  XNOR U6666 ( .A(y[217]), .B(x[217]), .Z(n5528) );
  XNOR U6667 ( .A(y[218]), .B(x[218]), .Z(n5527) );
  XNOR U6668 ( .A(n5518), .B(n5517), .Z(n5521) );
  XNOR U6669 ( .A(n5513), .B(n5514), .Z(n5517) );
  XNOR U6670 ( .A(y[213]), .B(x[213]), .Z(n5514) );
  XNOR U6671 ( .A(n5515), .B(n5516), .Z(n5513) );
  XNOR U6672 ( .A(y[214]), .B(x[214]), .Z(n5516) );
  XNOR U6673 ( .A(y[215]), .B(x[215]), .Z(n5515) );
  XNOR U6674 ( .A(n5507), .B(n5508), .Z(n5518) );
  XNOR U6675 ( .A(y[210]), .B(x[210]), .Z(n5508) );
  XNOR U6676 ( .A(n5509), .B(n5510), .Z(n5507) );
  XNOR U6677 ( .A(y[211]), .B(x[211]), .Z(n5510) );
  XNOR U6678 ( .A(y[212]), .B(x[212]), .Z(n5509) );
  XOR U6679 ( .A(n5483), .B(n5484), .Z(n5502) );
  XNOR U6680 ( .A(n5499), .B(n5500), .Z(n5484) );
  XNOR U6681 ( .A(n5494), .B(n5495), .Z(n5500) );
  XNOR U6682 ( .A(n5496), .B(n5497), .Z(n5495) );
  XNOR U6683 ( .A(y[208]), .B(x[208]), .Z(n5497) );
  XNOR U6684 ( .A(y[209]), .B(x[209]), .Z(n5496) );
  XNOR U6685 ( .A(y[207]), .B(x[207]), .Z(n5494) );
  XNOR U6686 ( .A(n5488), .B(n5489), .Z(n5499) );
  XNOR U6687 ( .A(y[204]), .B(x[204]), .Z(n5489) );
  XNOR U6688 ( .A(n5490), .B(n5491), .Z(n5488) );
  XNOR U6689 ( .A(y[205]), .B(x[205]), .Z(n5491) );
  XNOR U6690 ( .A(y[206]), .B(x[206]), .Z(n5490) );
  XOR U6691 ( .A(n5482), .B(n5481), .Z(n5483) );
  XNOR U6692 ( .A(n5477), .B(n5478), .Z(n5481) );
  XNOR U6693 ( .A(y[201]), .B(x[201]), .Z(n5478) );
  XNOR U6694 ( .A(n5479), .B(n5480), .Z(n5477) );
  XNOR U6695 ( .A(y[202]), .B(x[202]), .Z(n5480) );
  XNOR U6696 ( .A(y[203]), .B(x[203]), .Z(n5479) );
  XNOR U6697 ( .A(n5471), .B(n5472), .Z(n5482) );
  XNOR U6698 ( .A(y[198]), .B(x[198]), .Z(n5472) );
  XNOR U6699 ( .A(n5473), .B(n5474), .Z(n5471) );
  XNOR U6700 ( .A(y[199]), .B(x[199]), .Z(n5474) );
  XNOR U6701 ( .A(y[200]), .B(x[200]), .Z(n5473) );
  NAND U6702 ( .A(n5538), .B(n5539), .Z(N5868) );
  NANDN U6703 ( .A(n5540), .B(n5541), .Z(n5539) );
  OR U6704 ( .A(n5542), .B(n5543), .Z(n5541) );
  NAND U6705 ( .A(n5542), .B(n5543), .Z(n5538) );
  XOR U6706 ( .A(n5542), .B(n5544), .Z(N5867) );
  XNOR U6707 ( .A(n5540), .B(n5543), .Z(n5544) );
  AND U6708 ( .A(n5545), .B(n5546), .Z(n5543) );
  NANDN U6709 ( .A(n5547), .B(n5548), .Z(n5546) );
  NANDN U6710 ( .A(n5549), .B(n5550), .Z(n5548) );
  NANDN U6711 ( .A(n5550), .B(n5549), .Z(n5545) );
  NAND U6712 ( .A(n5551), .B(n5552), .Z(n5540) );
  NANDN U6713 ( .A(n5553), .B(n5554), .Z(n5552) );
  OR U6714 ( .A(n5555), .B(n5556), .Z(n5554) );
  NAND U6715 ( .A(n5556), .B(n5555), .Z(n5551) );
  AND U6716 ( .A(n5557), .B(n5558), .Z(n5542) );
  NANDN U6717 ( .A(n5559), .B(n5560), .Z(n5558) );
  NANDN U6718 ( .A(n5561), .B(n5562), .Z(n5560) );
  NANDN U6719 ( .A(n5562), .B(n5561), .Z(n5557) );
  XOR U6720 ( .A(n5556), .B(n5563), .Z(N5866) );
  XOR U6721 ( .A(n5553), .B(n5555), .Z(n5563) );
  XNOR U6722 ( .A(n5549), .B(n5564), .Z(n5555) );
  XNOR U6723 ( .A(n5547), .B(n5550), .Z(n5564) );
  NAND U6724 ( .A(n5565), .B(n5566), .Z(n5550) );
  NAND U6725 ( .A(n5567), .B(n5568), .Z(n5566) );
  OR U6726 ( .A(n5569), .B(n5570), .Z(n5567) );
  NANDN U6727 ( .A(n5571), .B(n5569), .Z(n5565) );
  IV U6728 ( .A(n5570), .Z(n5571) );
  NAND U6729 ( .A(n5572), .B(n5573), .Z(n5547) );
  NAND U6730 ( .A(n5574), .B(n5575), .Z(n5573) );
  NANDN U6731 ( .A(n5576), .B(n5577), .Z(n5574) );
  NANDN U6732 ( .A(n5577), .B(n5576), .Z(n5572) );
  AND U6733 ( .A(n5578), .B(n5579), .Z(n5549) );
  NAND U6734 ( .A(n5580), .B(n5581), .Z(n5579) );
  OR U6735 ( .A(n5582), .B(n5583), .Z(n5580) );
  NANDN U6736 ( .A(n5584), .B(n5582), .Z(n5578) );
  NAND U6737 ( .A(n5585), .B(n5586), .Z(n5553) );
  NANDN U6738 ( .A(n5587), .B(n5588), .Z(n5586) );
  OR U6739 ( .A(n5589), .B(n5590), .Z(n5588) );
  NANDN U6740 ( .A(n5591), .B(n5589), .Z(n5585) );
  IV U6741 ( .A(n5590), .Z(n5591) );
  XNOR U6742 ( .A(n5561), .B(n5592), .Z(n5556) );
  XNOR U6743 ( .A(n5559), .B(n5562), .Z(n5592) );
  NAND U6744 ( .A(n5593), .B(n5594), .Z(n5562) );
  NAND U6745 ( .A(n5595), .B(n5596), .Z(n5594) );
  OR U6746 ( .A(n5597), .B(n5598), .Z(n5595) );
  NANDN U6747 ( .A(n5599), .B(n5597), .Z(n5593) );
  IV U6748 ( .A(n5598), .Z(n5599) );
  NAND U6749 ( .A(n5600), .B(n5601), .Z(n5559) );
  NAND U6750 ( .A(n5602), .B(n5603), .Z(n5601) );
  NANDN U6751 ( .A(n5604), .B(n5605), .Z(n5602) );
  NANDN U6752 ( .A(n5605), .B(n5604), .Z(n5600) );
  AND U6753 ( .A(n5606), .B(n5607), .Z(n5561) );
  NAND U6754 ( .A(n5608), .B(n5609), .Z(n5607) );
  OR U6755 ( .A(n5610), .B(n5611), .Z(n5608) );
  NANDN U6756 ( .A(n5612), .B(n5610), .Z(n5606) );
  XNOR U6757 ( .A(n5587), .B(n5613), .Z(N5865) );
  XOR U6758 ( .A(n5589), .B(n5590), .Z(n5613) );
  XNOR U6759 ( .A(n5603), .B(n5614), .Z(n5590) );
  XOR U6760 ( .A(n5604), .B(n5605), .Z(n5614) );
  XOR U6761 ( .A(n5610), .B(n5615), .Z(n5605) );
  XOR U6762 ( .A(n5609), .B(n5612), .Z(n5615) );
  IV U6763 ( .A(n5611), .Z(n5612) );
  NAND U6764 ( .A(n5616), .B(n5617), .Z(n5611) );
  OR U6765 ( .A(n5618), .B(n5619), .Z(n5617) );
  OR U6766 ( .A(n5620), .B(n5621), .Z(n5616) );
  NAND U6767 ( .A(n5622), .B(n5623), .Z(n5609) );
  OR U6768 ( .A(n5624), .B(n5625), .Z(n5623) );
  OR U6769 ( .A(n5626), .B(n5627), .Z(n5622) );
  NOR U6770 ( .A(n5628), .B(n5629), .Z(n5610) );
  ANDN U6771 ( .B(n5630), .A(n5631), .Z(n5604) );
  XNOR U6772 ( .A(n5597), .B(n5632), .Z(n5603) );
  XNOR U6773 ( .A(n5596), .B(n5598), .Z(n5632) );
  NAND U6774 ( .A(n5633), .B(n5634), .Z(n5598) );
  OR U6775 ( .A(n5635), .B(n5636), .Z(n5634) );
  OR U6776 ( .A(n5637), .B(n5638), .Z(n5633) );
  NAND U6777 ( .A(n5639), .B(n5640), .Z(n5596) );
  OR U6778 ( .A(n5641), .B(n5642), .Z(n5640) );
  OR U6779 ( .A(n5643), .B(n5644), .Z(n5639) );
  ANDN U6780 ( .B(n5645), .A(n5646), .Z(n5597) );
  IV U6781 ( .A(n5647), .Z(n5645) );
  ANDN U6782 ( .B(n5648), .A(n5649), .Z(n5589) );
  XOR U6783 ( .A(n5575), .B(n5650), .Z(n5587) );
  XOR U6784 ( .A(n5576), .B(n5577), .Z(n5650) );
  XOR U6785 ( .A(n5582), .B(n5651), .Z(n5577) );
  XOR U6786 ( .A(n5581), .B(n5584), .Z(n5651) );
  IV U6787 ( .A(n5583), .Z(n5584) );
  NAND U6788 ( .A(n5652), .B(n5653), .Z(n5583) );
  OR U6789 ( .A(n5654), .B(n5655), .Z(n5653) );
  OR U6790 ( .A(n5656), .B(n5657), .Z(n5652) );
  NAND U6791 ( .A(n5658), .B(n5659), .Z(n5581) );
  OR U6792 ( .A(n5660), .B(n5661), .Z(n5659) );
  OR U6793 ( .A(n5662), .B(n5663), .Z(n5658) );
  NOR U6794 ( .A(n5664), .B(n5665), .Z(n5582) );
  ANDN U6795 ( .B(n5666), .A(n5667), .Z(n5576) );
  IV U6796 ( .A(n5668), .Z(n5666) );
  XNOR U6797 ( .A(n5569), .B(n5669), .Z(n5575) );
  XNOR U6798 ( .A(n5568), .B(n5570), .Z(n5669) );
  NAND U6799 ( .A(n5670), .B(n5671), .Z(n5570) );
  OR U6800 ( .A(n5672), .B(n5673), .Z(n5671) );
  OR U6801 ( .A(n5674), .B(n5675), .Z(n5670) );
  NAND U6802 ( .A(n5676), .B(n5677), .Z(n5568) );
  OR U6803 ( .A(n5678), .B(n5679), .Z(n5677) );
  OR U6804 ( .A(n5680), .B(n5681), .Z(n5676) );
  ANDN U6805 ( .B(n5682), .A(n5683), .Z(n5569) );
  IV U6806 ( .A(n5684), .Z(n5682) );
  XNOR U6807 ( .A(n5649), .B(n5648), .Z(N5864) );
  XOR U6808 ( .A(n5668), .B(n5667), .Z(n5648) );
  XNOR U6809 ( .A(n5683), .B(n5684), .Z(n5667) );
  XNOR U6810 ( .A(n5678), .B(n5679), .Z(n5684) );
  XNOR U6811 ( .A(n5680), .B(n5681), .Z(n5679) );
  XNOR U6812 ( .A(y[196]), .B(x[196]), .Z(n5681) );
  XNOR U6813 ( .A(y[197]), .B(x[197]), .Z(n5680) );
  XNOR U6814 ( .A(y[195]), .B(x[195]), .Z(n5678) );
  XNOR U6815 ( .A(n5672), .B(n5673), .Z(n5683) );
  XNOR U6816 ( .A(y[192]), .B(x[192]), .Z(n5673) );
  XNOR U6817 ( .A(n5674), .B(n5675), .Z(n5672) );
  XNOR U6818 ( .A(y[193]), .B(x[193]), .Z(n5675) );
  XNOR U6819 ( .A(y[194]), .B(x[194]), .Z(n5674) );
  XNOR U6820 ( .A(n5665), .B(n5664), .Z(n5668) );
  XNOR U6821 ( .A(n5660), .B(n5661), .Z(n5664) );
  XNOR U6822 ( .A(y[189]), .B(x[189]), .Z(n5661) );
  XNOR U6823 ( .A(n5662), .B(n5663), .Z(n5660) );
  XNOR U6824 ( .A(y[190]), .B(x[190]), .Z(n5663) );
  XNOR U6825 ( .A(y[191]), .B(x[191]), .Z(n5662) );
  XNOR U6826 ( .A(n5654), .B(n5655), .Z(n5665) );
  XNOR U6827 ( .A(y[186]), .B(x[186]), .Z(n5655) );
  XNOR U6828 ( .A(n5656), .B(n5657), .Z(n5654) );
  XNOR U6829 ( .A(y[187]), .B(x[187]), .Z(n5657) );
  XNOR U6830 ( .A(y[188]), .B(x[188]), .Z(n5656) );
  XOR U6831 ( .A(n5630), .B(n5631), .Z(n5649) );
  XNOR U6832 ( .A(n5646), .B(n5647), .Z(n5631) );
  XNOR U6833 ( .A(n5641), .B(n5642), .Z(n5647) );
  XNOR U6834 ( .A(n5643), .B(n5644), .Z(n5642) );
  XNOR U6835 ( .A(y[184]), .B(x[184]), .Z(n5644) );
  XNOR U6836 ( .A(y[185]), .B(x[185]), .Z(n5643) );
  XNOR U6837 ( .A(y[183]), .B(x[183]), .Z(n5641) );
  XNOR U6838 ( .A(n5635), .B(n5636), .Z(n5646) );
  XNOR U6839 ( .A(y[180]), .B(x[180]), .Z(n5636) );
  XNOR U6840 ( .A(n5637), .B(n5638), .Z(n5635) );
  XNOR U6841 ( .A(y[181]), .B(x[181]), .Z(n5638) );
  XNOR U6842 ( .A(y[182]), .B(x[182]), .Z(n5637) );
  XOR U6843 ( .A(n5629), .B(n5628), .Z(n5630) );
  XNOR U6844 ( .A(n5624), .B(n5625), .Z(n5628) );
  XNOR U6845 ( .A(y[177]), .B(x[177]), .Z(n5625) );
  XNOR U6846 ( .A(n5626), .B(n5627), .Z(n5624) );
  XNOR U6847 ( .A(y[178]), .B(x[178]), .Z(n5627) );
  XNOR U6848 ( .A(y[179]), .B(x[179]), .Z(n5626) );
  XNOR U6849 ( .A(n5618), .B(n5619), .Z(n5629) );
  XNOR U6850 ( .A(y[174]), .B(x[174]), .Z(n5619) );
  XNOR U6851 ( .A(n5620), .B(n5621), .Z(n5618) );
  XNOR U6852 ( .A(y[175]), .B(x[175]), .Z(n5621) );
  XNOR U6853 ( .A(y[176]), .B(x[176]), .Z(n5620) );
  NAND U6854 ( .A(n5685), .B(n5686), .Z(N5858) );
  NANDN U6855 ( .A(n5687), .B(n5688), .Z(n5686) );
  OR U6856 ( .A(n5689), .B(n5690), .Z(n5688) );
  NAND U6857 ( .A(n5689), .B(n5690), .Z(n5685) );
  XOR U6858 ( .A(n5689), .B(n5691), .Z(N5857) );
  XNOR U6859 ( .A(n5687), .B(n5690), .Z(n5691) );
  AND U6860 ( .A(n5692), .B(n5693), .Z(n5690) );
  NANDN U6861 ( .A(n5694), .B(n5695), .Z(n5693) );
  NANDN U6862 ( .A(n5696), .B(n5697), .Z(n5695) );
  NANDN U6863 ( .A(n5697), .B(n5696), .Z(n5692) );
  NAND U6864 ( .A(n5698), .B(n5699), .Z(n5687) );
  NANDN U6865 ( .A(n5700), .B(n5701), .Z(n5699) );
  OR U6866 ( .A(n5702), .B(n5703), .Z(n5701) );
  NAND U6867 ( .A(n5703), .B(n5702), .Z(n5698) );
  AND U6868 ( .A(n5704), .B(n5705), .Z(n5689) );
  NANDN U6869 ( .A(n5706), .B(n5707), .Z(n5705) );
  NANDN U6870 ( .A(n5708), .B(n5709), .Z(n5707) );
  NANDN U6871 ( .A(n5709), .B(n5708), .Z(n5704) );
  XOR U6872 ( .A(n5703), .B(n5710), .Z(N5856) );
  XOR U6873 ( .A(n5700), .B(n5702), .Z(n5710) );
  XNOR U6874 ( .A(n5696), .B(n5711), .Z(n5702) );
  XNOR U6875 ( .A(n5694), .B(n5697), .Z(n5711) );
  NAND U6876 ( .A(n5712), .B(n5713), .Z(n5697) );
  NAND U6877 ( .A(n5714), .B(n5715), .Z(n5713) );
  OR U6878 ( .A(n5716), .B(n5717), .Z(n5714) );
  NANDN U6879 ( .A(n5718), .B(n5716), .Z(n5712) );
  IV U6880 ( .A(n5717), .Z(n5718) );
  NAND U6881 ( .A(n5719), .B(n5720), .Z(n5694) );
  NAND U6882 ( .A(n5721), .B(n5722), .Z(n5720) );
  NANDN U6883 ( .A(n5723), .B(n5724), .Z(n5721) );
  NANDN U6884 ( .A(n5724), .B(n5723), .Z(n5719) );
  AND U6885 ( .A(n5725), .B(n5726), .Z(n5696) );
  NAND U6886 ( .A(n5727), .B(n5728), .Z(n5726) );
  OR U6887 ( .A(n5729), .B(n5730), .Z(n5727) );
  NANDN U6888 ( .A(n5731), .B(n5729), .Z(n5725) );
  NAND U6889 ( .A(n5732), .B(n5733), .Z(n5700) );
  NANDN U6890 ( .A(n5734), .B(n5735), .Z(n5733) );
  OR U6891 ( .A(n5736), .B(n5737), .Z(n5735) );
  NANDN U6892 ( .A(n5738), .B(n5736), .Z(n5732) );
  IV U6893 ( .A(n5737), .Z(n5738) );
  XNOR U6894 ( .A(n5708), .B(n5739), .Z(n5703) );
  XNOR U6895 ( .A(n5706), .B(n5709), .Z(n5739) );
  NAND U6896 ( .A(n5740), .B(n5741), .Z(n5709) );
  NAND U6897 ( .A(n5742), .B(n5743), .Z(n5741) );
  OR U6898 ( .A(n5744), .B(n5745), .Z(n5742) );
  NANDN U6899 ( .A(n5746), .B(n5744), .Z(n5740) );
  IV U6900 ( .A(n5745), .Z(n5746) );
  NAND U6901 ( .A(n5747), .B(n5748), .Z(n5706) );
  NAND U6902 ( .A(n5749), .B(n5750), .Z(n5748) );
  NANDN U6903 ( .A(n5751), .B(n5752), .Z(n5749) );
  NANDN U6904 ( .A(n5752), .B(n5751), .Z(n5747) );
  AND U6905 ( .A(n5753), .B(n5754), .Z(n5708) );
  NAND U6906 ( .A(n5755), .B(n5756), .Z(n5754) );
  OR U6907 ( .A(n5757), .B(n5758), .Z(n5755) );
  NANDN U6908 ( .A(n5759), .B(n5757), .Z(n5753) );
  XNOR U6909 ( .A(n5734), .B(n5760), .Z(N5855) );
  XOR U6910 ( .A(n5736), .B(n5737), .Z(n5760) );
  XNOR U6911 ( .A(n5750), .B(n5761), .Z(n5737) );
  XOR U6912 ( .A(n5751), .B(n5752), .Z(n5761) );
  XOR U6913 ( .A(n5757), .B(n5762), .Z(n5752) );
  XOR U6914 ( .A(n5756), .B(n5759), .Z(n5762) );
  IV U6915 ( .A(n5758), .Z(n5759) );
  NAND U6916 ( .A(n5763), .B(n5764), .Z(n5758) );
  OR U6917 ( .A(n5765), .B(n5766), .Z(n5764) );
  OR U6918 ( .A(n5767), .B(n5768), .Z(n5763) );
  NAND U6919 ( .A(n5769), .B(n5770), .Z(n5756) );
  OR U6920 ( .A(n5771), .B(n5772), .Z(n5770) );
  OR U6921 ( .A(n5773), .B(n5774), .Z(n5769) );
  NOR U6922 ( .A(n5775), .B(n5776), .Z(n5757) );
  ANDN U6923 ( .B(n5777), .A(n5778), .Z(n5751) );
  XNOR U6924 ( .A(n5744), .B(n5779), .Z(n5750) );
  XNOR U6925 ( .A(n5743), .B(n5745), .Z(n5779) );
  NAND U6926 ( .A(n5780), .B(n5781), .Z(n5745) );
  OR U6927 ( .A(n5782), .B(n5783), .Z(n5781) );
  OR U6928 ( .A(n5784), .B(n5785), .Z(n5780) );
  NAND U6929 ( .A(n5786), .B(n5787), .Z(n5743) );
  OR U6930 ( .A(n5788), .B(n5789), .Z(n5787) );
  OR U6931 ( .A(n5790), .B(n5791), .Z(n5786) );
  ANDN U6932 ( .B(n5792), .A(n5793), .Z(n5744) );
  IV U6933 ( .A(n5794), .Z(n5792) );
  ANDN U6934 ( .B(n5795), .A(n5796), .Z(n5736) );
  XOR U6935 ( .A(n5722), .B(n5797), .Z(n5734) );
  XOR U6936 ( .A(n5723), .B(n5724), .Z(n5797) );
  XOR U6937 ( .A(n5729), .B(n5798), .Z(n5724) );
  XOR U6938 ( .A(n5728), .B(n5731), .Z(n5798) );
  IV U6939 ( .A(n5730), .Z(n5731) );
  NAND U6940 ( .A(n5799), .B(n5800), .Z(n5730) );
  OR U6941 ( .A(n5801), .B(n5802), .Z(n5800) );
  OR U6942 ( .A(n5803), .B(n5804), .Z(n5799) );
  NAND U6943 ( .A(n5805), .B(n5806), .Z(n5728) );
  OR U6944 ( .A(n5807), .B(n5808), .Z(n5806) );
  OR U6945 ( .A(n5809), .B(n5810), .Z(n5805) );
  NOR U6946 ( .A(n5811), .B(n5812), .Z(n5729) );
  ANDN U6947 ( .B(n5813), .A(n5814), .Z(n5723) );
  IV U6948 ( .A(n5815), .Z(n5813) );
  XNOR U6949 ( .A(n5716), .B(n5816), .Z(n5722) );
  XNOR U6950 ( .A(n5715), .B(n5717), .Z(n5816) );
  NAND U6951 ( .A(n5817), .B(n5818), .Z(n5717) );
  OR U6952 ( .A(n5819), .B(n5820), .Z(n5818) );
  OR U6953 ( .A(n5821), .B(n5822), .Z(n5817) );
  NAND U6954 ( .A(n5823), .B(n5824), .Z(n5715) );
  OR U6955 ( .A(n5825), .B(n5826), .Z(n5824) );
  OR U6956 ( .A(n5827), .B(n5828), .Z(n5823) );
  ANDN U6957 ( .B(n5829), .A(n5830), .Z(n5716) );
  IV U6958 ( .A(n5831), .Z(n5829) );
  XNOR U6959 ( .A(n5796), .B(n5795), .Z(N5854) );
  XOR U6960 ( .A(n5815), .B(n5814), .Z(n5795) );
  XNOR U6961 ( .A(n5830), .B(n5831), .Z(n5814) );
  XNOR U6962 ( .A(n5825), .B(n5826), .Z(n5831) );
  XNOR U6963 ( .A(n5827), .B(n5828), .Z(n5826) );
  XNOR U6964 ( .A(y[172]), .B(x[172]), .Z(n5828) );
  XNOR U6965 ( .A(y[173]), .B(x[173]), .Z(n5827) );
  XNOR U6966 ( .A(y[171]), .B(x[171]), .Z(n5825) );
  XNOR U6967 ( .A(n5819), .B(n5820), .Z(n5830) );
  XNOR U6968 ( .A(y[168]), .B(x[168]), .Z(n5820) );
  XNOR U6969 ( .A(n5821), .B(n5822), .Z(n5819) );
  XNOR U6970 ( .A(y[169]), .B(x[169]), .Z(n5822) );
  XNOR U6971 ( .A(y[170]), .B(x[170]), .Z(n5821) );
  XNOR U6972 ( .A(n5812), .B(n5811), .Z(n5815) );
  XNOR U6973 ( .A(n5807), .B(n5808), .Z(n5811) );
  XNOR U6974 ( .A(y[165]), .B(x[165]), .Z(n5808) );
  XNOR U6975 ( .A(n5809), .B(n5810), .Z(n5807) );
  XNOR U6976 ( .A(y[166]), .B(x[166]), .Z(n5810) );
  XNOR U6977 ( .A(y[167]), .B(x[167]), .Z(n5809) );
  XNOR U6978 ( .A(n5801), .B(n5802), .Z(n5812) );
  XNOR U6979 ( .A(y[162]), .B(x[162]), .Z(n5802) );
  XNOR U6980 ( .A(n5803), .B(n5804), .Z(n5801) );
  XNOR U6981 ( .A(y[163]), .B(x[163]), .Z(n5804) );
  XNOR U6982 ( .A(y[164]), .B(x[164]), .Z(n5803) );
  XOR U6983 ( .A(n5777), .B(n5778), .Z(n5796) );
  XNOR U6984 ( .A(n5793), .B(n5794), .Z(n5778) );
  XNOR U6985 ( .A(n5788), .B(n5789), .Z(n5794) );
  XNOR U6986 ( .A(n5790), .B(n5791), .Z(n5789) );
  XNOR U6987 ( .A(y[160]), .B(x[160]), .Z(n5791) );
  XNOR U6988 ( .A(y[161]), .B(x[161]), .Z(n5790) );
  XNOR U6989 ( .A(y[159]), .B(x[159]), .Z(n5788) );
  XNOR U6990 ( .A(n5782), .B(n5783), .Z(n5793) );
  XNOR U6991 ( .A(y[156]), .B(x[156]), .Z(n5783) );
  XNOR U6992 ( .A(n5784), .B(n5785), .Z(n5782) );
  XNOR U6993 ( .A(y[157]), .B(x[157]), .Z(n5785) );
  XNOR U6994 ( .A(y[158]), .B(x[158]), .Z(n5784) );
  XOR U6995 ( .A(n5776), .B(n5775), .Z(n5777) );
  XNOR U6996 ( .A(n5771), .B(n5772), .Z(n5775) );
  XNOR U6997 ( .A(y[153]), .B(x[153]), .Z(n5772) );
  XNOR U6998 ( .A(n5773), .B(n5774), .Z(n5771) );
  XNOR U6999 ( .A(y[154]), .B(x[154]), .Z(n5774) );
  XNOR U7000 ( .A(y[155]), .B(x[155]), .Z(n5773) );
  XNOR U7001 ( .A(n5765), .B(n5766), .Z(n5776) );
  XNOR U7002 ( .A(y[150]), .B(x[150]), .Z(n5766) );
  XNOR U7003 ( .A(n5767), .B(n5768), .Z(n5765) );
  XNOR U7004 ( .A(y[151]), .B(x[151]), .Z(n5768) );
  XNOR U7005 ( .A(y[152]), .B(x[152]), .Z(n5767) );
  NAND U7006 ( .A(n5832), .B(n5833), .Z(N5848) );
  NANDN U7007 ( .A(n5834), .B(n5835), .Z(n5833) );
  OR U7008 ( .A(n5836), .B(n5837), .Z(n5835) );
  NAND U7009 ( .A(n5836), .B(n5837), .Z(n5832) );
  XOR U7010 ( .A(n5836), .B(n5838), .Z(N5847) );
  XNOR U7011 ( .A(n5834), .B(n5837), .Z(n5838) );
  AND U7012 ( .A(n5839), .B(n5840), .Z(n5837) );
  NANDN U7013 ( .A(n5841), .B(n5842), .Z(n5840) );
  NANDN U7014 ( .A(n5843), .B(n5844), .Z(n5842) );
  NANDN U7015 ( .A(n5844), .B(n5843), .Z(n5839) );
  NAND U7016 ( .A(n5845), .B(n5846), .Z(n5834) );
  NANDN U7017 ( .A(n5847), .B(n5848), .Z(n5846) );
  OR U7018 ( .A(n5849), .B(n5850), .Z(n5848) );
  NAND U7019 ( .A(n5850), .B(n5849), .Z(n5845) );
  AND U7020 ( .A(n5851), .B(n5852), .Z(n5836) );
  NANDN U7021 ( .A(n5853), .B(n5854), .Z(n5852) );
  NANDN U7022 ( .A(n5855), .B(n5856), .Z(n5854) );
  NANDN U7023 ( .A(n5856), .B(n5855), .Z(n5851) );
  XOR U7024 ( .A(n5850), .B(n5857), .Z(N5846) );
  XOR U7025 ( .A(n5847), .B(n5849), .Z(n5857) );
  XNOR U7026 ( .A(n5843), .B(n5858), .Z(n5849) );
  XNOR U7027 ( .A(n5841), .B(n5844), .Z(n5858) );
  NAND U7028 ( .A(n5859), .B(n5860), .Z(n5844) );
  NAND U7029 ( .A(n5861), .B(n5862), .Z(n5860) );
  OR U7030 ( .A(n5863), .B(n5864), .Z(n5861) );
  NANDN U7031 ( .A(n5865), .B(n5863), .Z(n5859) );
  IV U7032 ( .A(n5864), .Z(n5865) );
  NAND U7033 ( .A(n5866), .B(n5867), .Z(n5841) );
  NAND U7034 ( .A(n5868), .B(n5869), .Z(n5867) );
  NANDN U7035 ( .A(n5870), .B(n5871), .Z(n5868) );
  NANDN U7036 ( .A(n5871), .B(n5870), .Z(n5866) );
  AND U7037 ( .A(n5872), .B(n5873), .Z(n5843) );
  NAND U7038 ( .A(n5874), .B(n5875), .Z(n5873) );
  OR U7039 ( .A(n5876), .B(n5877), .Z(n5874) );
  NANDN U7040 ( .A(n5878), .B(n5876), .Z(n5872) );
  NAND U7041 ( .A(n5879), .B(n5880), .Z(n5847) );
  NANDN U7042 ( .A(n5881), .B(n5882), .Z(n5880) );
  OR U7043 ( .A(n5883), .B(n5884), .Z(n5882) );
  NANDN U7044 ( .A(n5885), .B(n5883), .Z(n5879) );
  IV U7045 ( .A(n5884), .Z(n5885) );
  XNOR U7046 ( .A(n5855), .B(n5886), .Z(n5850) );
  XNOR U7047 ( .A(n5853), .B(n5856), .Z(n5886) );
  NAND U7048 ( .A(n5887), .B(n5888), .Z(n5856) );
  NAND U7049 ( .A(n5889), .B(n5890), .Z(n5888) );
  OR U7050 ( .A(n5891), .B(n5892), .Z(n5889) );
  NANDN U7051 ( .A(n5893), .B(n5891), .Z(n5887) );
  IV U7052 ( .A(n5892), .Z(n5893) );
  NAND U7053 ( .A(n5894), .B(n5895), .Z(n5853) );
  NAND U7054 ( .A(n5896), .B(n5897), .Z(n5895) );
  NANDN U7055 ( .A(n5898), .B(n5899), .Z(n5896) );
  NANDN U7056 ( .A(n5899), .B(n5898), .Z(n5894) );
  AND U7057 ( .A(n5900), .B(n5901), .Z(n5855) );
  NAND U7058 ( .A(n5902), .B(n5903), .Z(n5901) );
  OR U7059 ( .A(n5904), .B(n5905), .Z(n5902) );
  NANDN U7060 ( .A(n5906), .B(n5904), .Z(n5900) );
  XNOR U7061 ( .A(n5881), .B(n5907), .Z(N5845) );
  XOR U7062 ( .A(n5883), .B(n5884), .Z(n5907) );
  XNOR U7063 ( .A(n5897), .B(n5908), .Z(n5884) );
  XOR U7064 ( .A(n5898), .B(n5899), .Z(n5908) );
  XOR U7065 ( .A(n5904), .B(n5909), .Z(n5899) );
  XOR U7066 ( .A(n5903), .B(n5906), .Z(n5909) );
  IV U7067 ( .A(n5905), .Z(n5906) );
  NAND U7068 ( .A(n5910), .B(n5911), .Z(n5905) );
  OR U7069 ( .A(n5912), .B(n5913), .Z(n5911) );
  OR U7070 ( .A(n5914), .B(n5915), .Z(n5910) );
  NAND U7071 ( .A(n5916), .B(n5917), .Z(n5903) );
  OR U7072 ( .A(n5918), .B(n5919), .Z(n5917) );
  OR U7073 ( .A(n5920), .B(n5921), .Z(n5916) );
  NOR U7074 ( .A(n5922), .B(n5923), .Z(n5904) );
  ANDN U7075 ( .B(n5924), .A(n5925), .Z(n5898) );
  XNOR U7076 ( .A(n5891), .B(n5926), .Z(n5897) );
  XNOR U7077 ( .A(n5890), .B(n5892), .Z(n5926) );
  NAND U7078 ( .A(n5927), .B(n5928), .Z(n5892) );
  OR U7079 ( .A(n5929), .B(n5930), .Z(n5928) );
  OR U7080 ( .A(n5931), .B(n5932), .Z(n5927) );
  NAND U7081 ( .A(n5933), .B(n5934), .Z(n5890) );
  OR U7082 ( .A(n5935), .B(n5936), .Z(n5934) );
  OR U7083 ( .A(n5937), .B(n5938), .Z(n5933) );
  ANDN U7084 ( .B(n5939), .A(n5940), .Z(n5891) );
  IV U7085 ( .A(n5941), .Z(n5939) );
  ANDN U7086 ( .B(n5942), .A(n5943), .Z(n5883) );
  XOR U7087 ( .A(n5869), .B(n5944), .Z(n5881) );
  XOR U7088 ( .A(n5870), .B(n5871), .Z(n5944) );
  XOR U7089 ( .A(n5876), .B(n5945), .Z(n5871) );
  XOR U7090 ( .A(n5875), .B(n5878), .Z(n5945) );
  IV U7091 ( .A(n5877), .Z(n5878) );
  NAND U7092 ( .A(n5946), .B(n5947), .Z(n5877) );
  OR U7093 ( .A(n5948), .B(n5949), .Z(n5947) );
  OR U7094 ( .A(n5950), .B(n5951), .Z(n5946) );
  NAND U7095 ( .A(n5952), .B(n5953), .Z(n5875) );
  OR U7096 ( .A(n5954), .B(n5955), .Z(n5953) );
  OR U7097 ( .A(n5956), .B(n5957), .Z(n5952) );
  NOR U7098 ( .A(n5958), .B(n5959), .Z(n5876) );
  ANDN U7099 ( .B(n5960), .A(n5961), .Z(n5870) );
  IV U7100 ( .A(n5962), .Z(n5960) );
  XNOR U7101 ( .A(n5863), .B(n5963), .Z(n5869) );
  XNOR U7102 ( .A(n5862), .B(n5864), .Z(n5963) );
  NAND U7103 ( .A(n5964), .B(n5965), .Z(n5864) );
  OR U7104 ( .A(n5966), .B(n5967), .Z(n5965) );
  OR U7105 ( .A(n5968), .B(n5969), .Z(n5964) );
  NAND U7106 ( .A(n5970), .B(n5971), .Z(n5862) );
  OR U7107 ( .A(n5972), .B(n5973), .Z(n5971) );
  OR U7108 ( .A(n5974), .B(n5975), .Z(n5970) );
  ANDN U7109 ( .B(n5976), .A(n5977), .Z(n5863) );
  IV U7110 ( .A(n5978), .Z(n5976) );
  XNOR U7111 ( .A(n5943), .B(n5942), .Z(N5844) );
  XOR U7112 ( .A(n5962), .B(n5961), .Z(n5942) );
  XNOR U7113 ( .A(n5977), .B(n5978), .Z(n5961) );
  XNOR U7114 ( .A(n5972), .B(n5973), .Z(n5978) );
  XNOR U7115 ( .A(n5974), .B(n5975), .Z(n5973) );
  XNOR U7116 ( .A(y[148]), .B(x[148]), .Z(n5975) );
  XNOR U7117 ( .A(y[149]), .B(x[149]), .Z(n5974) );
  XNOR U7118 ( .A(y[147]), .B(x[147]), .Z(n5972) );
  XNOR U7119 ( .A(n5966), .B(n5967), .Z(n5977) );
  XNOR U7120 ( .A(y[144]), .B(x[144]), .Z(n5967) );
  XNOR U7121 ( .A(n5968), .B(n5969), .Z(n5966) );
  XNOR U7122 ( .A(y[145]), .B(x[145]), .Z(n5969) );
  XNOR U7123 ( .A(y[146]), .B(x[146]), .Z(n5968) );
  XNOR U7124 ( .A(n5959), .B(n5958), .Z(n5962) );
  XNOR U7125 ( .A(n5954), .B(n5955), .Z(n5958) );
  XNOR U7126 ( .A(y[141]), .B(x[141]), .Z(n5955) );
  XNOR U7127 ( .A(n5956), .B(n5957), .Z(n5954) );
  XNOR U7128 ( .A(y[142]), .B(x[142]), .Z(n5957) );
  XNOR U7129 ( .A(y[143]), .B(x[143]), .Z(n5956) );
  XNOR U7130 ( .A(n5948), .B(n5949), .Z(n5959) );
  XNOR U7131 ( .A(y[138]), .B(x[138]), .Z(n5949) );
  XNOR U7132 ( .A(n5950), .B(n5951), .Z(n5948) );
  XNOR U7133 ( .A(y[139]), .B(x[139]), .Z(n5951) );
  XNOR U7134 ( .A(y[140]), .B(x[140]), .Z(n5950) );
  XOR U7135 ( .A(n5924), .B(n5925), .Z(n5943) );
  XNOR U7136 ( .A(n5940), .B(n5941), .Z(n5925) );
  XNOR U7137 ( .A(n5935), .B(n5936), .Z(n5941) );
  XNOR U7138 ( .A(n5937), .B(n5938), .Z(n5936) );
  XNOR U7139 ( .A(y[136]), .B(x[136]), .Z(n5938) );
  XNOR U7140 ( .A(y[137]), .B(x[137]), .Z(n5937) );
  XNOR U7141 ( .A(y[135]), .B(x[135]), .Z(n5935) );
  XNOR U7142 ( .A(n5929), .B(n5930), .Z(n5940) );
  XNOR U7143 ( .A(y[132]), .B(x[132]), .Z(n5930) );
  XNOR U7144 ( .A(n5931), .B(n5932), .Z(n5929) );
  XNOR U7145 ( .A(y[133]), .B(x[133]), .Z(n5932) );
  XNOR U7146 ( .A(y[134]), .B(x[134]), .Z(n5931) );
  XOR U7147 ( .A(n5923), .B(n5922), .Z(n5924) );
  XNOR U7148 ( .A(n5918), .B(n5919), .Z(n5922) );
  XNOR U7149 ( .A(y[129]), .B(x[129]), .Z(n5919) );
  XNOR U7150 ( .A(n5920), .B(n5921), .Z(n5918) );
  XNOR U7151 ( .A(y[130]), .B(x[130]), .Z(n5921) );
  XNOR U7152 ( .A(y[131]), .B(x[131]), .Z(n5920) );
  XNOR U7153 ( .A(n5912), .B(n5913), .Z(n5923) );
  XNOR U7154 ( .A(y[126]), .B(x[126]), .Z(n5913) );
  XNOR U7155 ( .A(n5914), .B(n5915), .Z(n5912) );
  XNOR U7156 ( .A(y[127]), .B(x[127]), .Z(n5915) );
  XNOR U7157 ( .A(y[128]), .B(x[128]), .Z(n5914) );
  NAND U7158 ( .A(n5979), .B(n5980), .Z(N5838) );
  NANDN U7159 ( .A(n5981), .B(n5982), .Z(n5980) );
  OR U7160 ( .A(n5983), .B(n5984), .Z(n5982) );
  NAND U7161 ( .A(n5983), .B(n5984), .Z(n5979) );
  XOR U7162 ( .A(n5983), .B(n5985), .Z(N5837) );
  XNOR U7163 ( .A(n5981), .B(n5984), .Z(n5985) );
  AND U7164 ( .A(n5986), .B(n5987), .Z(n5984) );
  NANDN U7165 ( .A(n5988), .B(n5989), .Z(n5987) );
  NANDN U7166 ( .A(n5990), .B(n5991), .Z(n5989) );
  NANDN U7167 ( .A(n5991), .B(n5990), .Z(n5986) );
  NAND U7168 ( .A(n5992), .B(n5993), .Z(n5981) );
  NANDN U7169 ( .A(n5994), .B(n5995), .Z(n5993) );
  OR U7170 ( .A(n5996), .B(n5997), .Z(n5995) );
  NAND U7171 ( .A(n5997), .B(n5996), .Z(n5992) );
  AND U7172 ( .A(n5998), .B(n5999), .Z(n5983) );
  NANDN U7173 ( .A(n6000), .B(n6001), .Z(n5999) );
  NANDN U7174 ( .A(n6002), .B(n6003), .Z(n6001) );
  NANDN U7175 ( .A(n6003), .B(n6002), .Z(n5998) );
  XOR U7176 ( .A(n5997), .B(n6004), .Z(N5836) );
  XOR U7177 ( .A(n5994), .B(n5996), .Z(n6004) );
  XNOR U7178 ( .A(n5990), .B(n6005), .Z(n5996) );
  XNOR U7179 ( .A(n5988), .B(n5991), .Z(n6005) );
  NAND U7180 ( .A(n6006), .B(n6007), .Z(n5991) );
  NAND U7181 ( .A(n6008), .B(n6009), .Z(n6007) );
  OR U7182 ( .A(n6010), .B(n6011), .Z(n6008) );
  NANDN U7183 ( .A(n6012), .B(n6010), .Z(n6006) );
  IV U7184 ( .A(n6011), .Z(n6012) );
  NAND U7185 ( .A(n6013), .B(n6014), .Z(n5988) );
  NAND U7186 ( .A(n6015), .B(n6016), .Z(n6014) );
  NANDN U7187 ( .A(n6017), .B(n6018), .Z(n6015) );
  NANDN U7188 ( .A(n6018), .B(n6017), .Z(n6013) );
  AND U7189 ( .A(n6019), .B(n6020), .Z(n5990) );
  NAND U7190 ( .A(n6021), .B(n6022), .Z(n6020) );
  OR U7191 ( .A(n6023), .B(n6024), .Z(n6021) );
  NANDN U7192 ( .A(n6025), .B(n6023), .Z(n6019) );
  NAND U7193 ( .A(n6026), .B(n6027), .Z(n5994) );
  NANDN U7194 ( .A(n6028), .B(n6029), .Z(n6027) );
  OR U7195 ( .A(n6030), .B(n6031), .Z(n6029) );
  NANDN U7196 ( .A(n6032), .B(n6030), .Z(n6026) );
  IV U7197 ( .A(n6031), .Z(n6032) );
  XNOR U7198 ( .A(n6002), .B(n6033), .Z(n5997) );
  XNOR U7199 ( .A(n6000), .B(n6003), .Z(n6033) );
  NAND U7200 ( .A(n6034), .B(n6035), .Z(n6003) );
  NAND U7201 ( .A(n6036), .B(n6037), .Z(n6035) );
  OR U7202 ( .A(n6038), .B(n6039), .Z(n6036) );
  NANDN U7203 ( .A(n6040), .B(n6038), .Z(n6034) );
  IV U7204 ( .A(n6039), .Z(n6040) );
  NAND U7205 ( .A(n6041), .B(n6042), .Z(n6000) );
  NAND U7206 ( .A(n6043), .B(n6044), .Z(n6042) );
  NANDN U7207 ( .A(n6045), .B(n6046), .Z(n6043) );
  NANDN U7208 ( .A(n6046), .B(n6045), .Z(n6041) );
  AND U7209 ( .A(n6047), .B(n6048), .Z(n6002) );
  NAND U7210 ( .A(n6049), .B(n6050), .Z(n6048) );
  OR U7211 ( .A(n6051), .B(n6052), .Z(n6049) );
  NANDN U7212 ( .A(n6053), .B(n6051), .Z(n6047) );
  XNOR U7213 ( .A(n6028), .B(n6054), .Z(N5835) );
  XOR U7214 ( .A(n6030), .B(n6031), .Z(n6054) );
  XNOR U7215 ( .A(n6044), .B(n6055), .Z(n6031) );
  XOR U7216 ( .A(n6045), .B(n6046), .Z(n6055) );
  XOR U7217 ( .A(n6051), .B(n6056), .Z(n6046) );
  XOR U7218 ( .A(n6050), .B(n6053), .Z(n6056) );
  IV U7219 ( .A(n6052), .Z(n6053) );
  NAND U7220 ( .A(n6057), .B(n6058), .Z(n6052) );
  OR U7221 ( .A(n6059), .B(n6060), .Z(n6058) );
  OR U7222 ( .A(n6061), .B(n6062), .Z(n6057) );
  NAND U7223 ( .A(n6063), .B(n6064), .Z(n6050) );
  OR U7224 ( .A(n6065), .B(n6066), .Z(n6064) );
  OR U7225 ( .A(n6067), .B(n6068), .Z(n6063) );
  NOR U7226 ( .A(n6069), .B(n6070), .Z(n6051) );
  ANDN U7227 ( .B(n6071), .A(n6072), .Z(n6045) );
  XNOR U7228 ( .A(n6038), .B(n6073), .Z(n6044) );
  XNOR U7229 ( .A(n6037), .B(n6039), .Z(n6073) );
  NAND U7230 ( .A(n6074), .B(n6075), .Z(n6039) );
  OR U7231 ( .A(n6076), .B(n6077), .Z(n6075) );
  OR U7232 ( .A(n6078), .B(n6079), .Z(n6074) );
  NAND U7233 ( .A(n6080), .B(n6081), .Z(n6037) );
  OR U7234 ( .A(n6082), .B(n6083), .Z(n6081) );
  OR U7235 ( .A(n6084), .B(n6085), .Z(n6080) );
  ANDN U7236 ( .B(n6086), .A(n6087), .Z(n6038) );
  IV U7237 ( .A(n6088), .Z(n6086) );
  ANDN U7238 ( .B(n6089), .A(n6090), .Z(n6030) );
  XOR U7239 ( .A(n6016), .B(n6091), .Z(n6028) );
  XOR U7240 ( .A(n6017), .B(n6018), .Z(n6091) );
  XOR U7241 ( .A(n6023), .B(n6092), .Z(n6018) );
  XOR U7242 ( .A(n6022), .B(n6025), .Z(n6092) );
  IV U7243 ( .A(n6024), .Z(n6025) );
  NAND U7244 ( .A(n6093), .B(n6094), .Z(n6024) );
  OR U7245 ( .A(n6095), .B(n6096), .Z(n6094) );
  OR U7246 ( .A(n6097), .B(n6098), .Z(n6093) );
  NAND U7247 ( .A(n6099), .B(n6100), .Z(n6022) );
  OR U7248 ( .A(n6101), .B(n6102), .Z(n6100) );
  OR U7249 ( .A(n6103), .B(n6104), .Z(n6099) );
  NOR U7250 ( .A(n6105), .B(n6106), .Z(n6023) );
  ANDN U7251 ( .B(n6107), .A(n6108), .Z(n6017) );
  IV U7252 ( .A(n6109), .Z(n6107) );
  XNOR U7253 ( .A(n6010), .B(n6110), .Z(n6016) );
  XNOR U7254 ( .A(n6009), .B(n6011), .Z(n6110) );
  NAND U7255 ( .A(n6111), .B(n6112), .Z(n6011) );
  OR U7256 ( .A(n6113), .B(n6114), .Z(n6112) );
  OR U7257 ( .A(n6115), .B(n6116), .Z(n6111) );
  NAND U7258 ( .A(n6117), .B(n6118), .Z(n6009) );
  OR U7259 ( .A(n6119), .B(n6120), .Z(n6118) );
  OR U7260 ( .A(n6121), .B(n6122), .Z(n6117) );
  ANDN U7261 ( .B(n6123), .A(n6124), .Z(n6010) );
  IV U7262 ( .A(n6125), .Z(n6123) );
  XNOR U7263 ( .A(n6090), .B(n6089), .Z(N5834) );
  XOR U7264 ( .A(n6109), .B(n6108), .Z(n6089) );
  XNOR U7265 ( .A(n6124), .B(n6125), .Z(n6108) );
  XNOR U7266 ( .A(n6119), .B(n6120), .Z(n6125) );
  XNOR U7267 ( .A(n6121), .B(n6122), .Z(n6120) );
  XNOR U7268 ( .A(y[124]), .B(x[124]), .Z(n6122) );
  XNOR U7269 ( .A(y[125]), .B(x[125]), .Z(n6121) );
  XNOR U7270 ( .A(y[123]), .B(x[123]), .Z(n6119) );
  XNOR U7271 ( .A(n6113), .B(n6114), .Z(n6124) );
  XNOR U7272 ( .A(y[120]), .B(x[120]), .Z(n6114) );
  XNOR U7273 ( .A(n6115), .B(n6116), .Z(n6113) );
  XNOR U7274 ( .A(y[121]), .B(x[121]), .Z(n6116) );
  XNOR U7275 ( .A(y[122]), .B(x[122]), .Z(n6115) );
  XNOR U7276 ( .A(n6106), .B(n6105), .Z(n6109) );
  XNOR U7277 ( .A(n6101), .B(n6102), .Z(n6105) );
  XNOR U7278 ( .A(y[117]), .B(x[117]), .Z(n6102) );
  XNOR U7279 ( .A(n6103), .B(n6104), .Z(n6101) );
  XNOR U7280 ( .A(y[118]), .B(x[118]), .Z(n6104) );
  XNOR U7281 ( .A(y[119]), .B(x[119]), .Z(n6103) );
  XNOR U7282 ( .A(n6095), .B(n6096), .Z(n6106) );
  XNOR U7283 ( .A(y[114]), .B(x[114]), .Z(n6096) );
  XNOR U7284 ( .A(n6097), .B(n6098), .Z(n6095) );
  XNOR U7285 ( .A(y[115]), .B(x[115]), .Z(n6098) );
  XNOR U7286 ( .A(y[116]), .B(x[116]), .Z(n6097) );
  XOR U7287 ( .A(n6071), .B(n6072), .Z(n6090) );
  XNOR U7288 ( .A(n6087), .B(n6088), .Z(n6072) );
  XNOR U7289 ( .A(n6082), .B(n6083), .Z(n6088) );
  XNOR U7290 ( .A(n6084), .B(n6085), .Z(n6083) );
  XNOR U7291 ( .A(y[112]), .B(x[112]), .Z(n6085) );
  XNOR U7292 ( .A(y[113]), .B(x[113]), .Z(n6084) );
  XNOR U7293 ( .A(y[111]), .B(x[111]), .Z(n6082) );
  XNOR U7294 ( .A(n6076), .B(n6077), .Z(n6087) );
  XNOR U7295 ( .A(y[108]), .B(x[108]), .Z(n6077) );
  XNOR U7296 ( .A(n6078), .B(n6079), .Z(n6076) );
  XNOR U7297 ( .A(y[109]), .B(x[109]), .Z(n6079) );
  XNOR U7298 ( .A(y[110]), .B(x[110]), .Z(n6078) );
  XOR U7299 ( .A(n6070), .B(n6069), .Z(n6071) );
  XNOR U7300 ( .A(n6065), .B(n6066), .Z(n6069) );
  XNOR U7301 ( .A(y[105]), .B(x[105]), .Z(n6066) );
  XNOR U7302 ( .A(n6067), .B(n6068), .Z(n6065) );
  XNOR U7303 ( .A(y[106]), .B(x[106]), .Z(n6068) );
  XNOR U7304 ( .A(y[107]), .B(x[107]), .Z(n6067) );
  XNOR U7305 ( .A(n6059), .B(n6060), .Z(n6070) );
  XNOR U7306 ( .A(y[102]), .B(x[102]), .Z(n6060) );
  XNOR U7307 ( .A(n6061), .B(n6062), .Z(n6059) );
  XNOR U7308 ( .A(y[103]), .B(x[103]), .Z(n6062) );
  XNOR U7309 ( .A(y[104]), .B(x[104]), .Z(n6061) );
  NAND U7310 ( .A(n6126), .B(n6127), .Z(N5828) );
  NANDN U7311 ( .A(n6128), .B(n6129), .Z(n6127) );
  OR U7312 ( .A(n6130), .B(n6131), .Z(n6129) );
  NAND U7313 ( .A(n6130), .B(n6131), .Z(n6126) );
  XOR U7314 ( .A(n6130), .B(n6132), .Z(N5827) );
  XNOR U7315 ( .A(n6128), .B(n6131), .Z(n6132) );
  AND U7316 ( .A(n6133), .B(n6134), .Z(n6131) );
  NANDN U7317 ( .A(n6135), .B(n6136), .Z(n6134) );
  NANDN U7318 ( .A(n6137), .B(n6138), .Z(n6136) );
  NANDN U7319 ( .A(n6138), .B(n6137), .Z(n6133) );
  NAND U7320 ( .A(n6139), .B(n6140), .Z(n6128) );
  NANDN U7321 ( .A(n6141), .B(n6142), .Z(n6140) );
  OR U7322 ( .A(n6143), .B(n6144), .Z(n6142) );
  NAND U7323 ( .A(n6144), .B(n6143), .Z(n6139) );
  AND U7324 ( .A(n6145), .B(n6146), .Z(n6130) );
  NANDN U7325 ( .A(n6147), .B(n6148), .Z(n6146) );
  NANDN U7326 ( .A(n6149), .B(n6150), .Z(n6148) );
  NANDN U7327 ( .A(n6150), .B(n6149), .Z(n6145) );
  XOR U7328 ( .A(n6144), .B(n6151), .Z(N5826) );
  XOR U7329 ( .A(n6141), .B(n6143), .Z(n6151) );
  XNOR U7330 ( .A(n6137), .B(n6152), .Z(n6143) );
  XNOR U7331 ( .A(n6135), .B(n6138), .Z(n6152) );
  NAND U7332 ( .A(n6153), .B(n6154), .Z(n6138) );
  NAND U7333 ( .A(n6155), .B(n6156), .Z(n6154) );
  OR U7334 ( .A(n6157), .B(n6158), .Z(n6155) );
  NANDN U7335 ( .A(n6159), .B(n6157), .Z(n6153) );
  IV U7336 ( .A(n6158), .Z(n6159) );
  NAND U7337 ( .A(n6160), .B(n6161), .Z(n6135) );
  NAND U7338 ( .A(n6162), .B(n6163), .Z(n6161) );
  NANDN U7339 ( .A(n6164), .B(n6165), .Z(n6162) );
  NANDN U7340 ( .A(n6165), .B(n6164), .Z(n6160) );
  AND U7341 ( .A(n6166), .B(n6167), .Z(n6137) );
  NAND U7342 ( .A(n6168), .B(n6169), .Z(n6167) );
  OR U7343 ( .A(n6170), .B(n6171), .Z(n6168) );
  NANDN U7344 ( .A(n6172), .B(n6170), .Z(n6166) );
  NAND U7345 ( .A(n6173), .B(n6174), .Z(n6141) );
  NANDN U7346 ( .A(n6175), .B(n6176), .Z(n6174) );
  OR U7347 ( .A(n6177), .B(n6178), .Z(n6176) );
  NANDN U7348 ( .A(n6179), .B(n6177), .Z(n6173) );
  IV U7349 ( .A(n6178), .Z(n6179) );
  XNOR U7350 ( .A(n6149), .B(n6180), .Z(n6144) );
  XNOR U7351 ( .A(n6147), .B(n6150), .Z(n6180) );
  NAND U7352 ( .A(n6181), .B(n6182), .Z(n6150) );
  NAND U7353 ( .A(n6183), .B(n6184), .Z(n6182) );
  OR U7354 ( .A(n6185), .B(n6186), .Z(n6183) );
  NANDN U7355 ( .A(n6187), .B(n6185), .Z(n6181) );
  IV U7356 ( .A(n6186), .Z(n6187) );
  NAND U7357 ( .A(n6188), .B(n6189), .Z(n6147) );
  NAND U7358 ( .A(n6190), .B(n6191), .Z(n6189) );
  NANDN U7359 ( .A(n6192), .B(n6193), .Z(n6190) );
  NANDN U7360 ( .A(n6193), .B(n6192), .Z(n6188) );
  AND U7361 ( .A(n6194), .B(n6195), .Z(n6149) );
  NAND U7362 ( .A(n6196), .B(n6197), .Z(n6195) );
  OR U7363 ( .A(n6198), .B(n6199), .Z(n6196) );
  NANDN U7364 ( .A(n6200), .B(n6198), .Z(n6194) );
  XNOR U7365 ( .A(n6175), .B(n6201), .Z(N5825) );
  XOR U7366 ( .A(n6177), .B(n6178), .Z(n6201) );
  XNOR U7367 ( .A(n6191), .B(n6202), .Z(n6178) );
  XOR U7368 ( .A(n6192), .B(n6193), .Z(n6202) );
  XOR U7369 ( .A(n6198), .B(n6203), .Z(n6193) );
  XOR U7370 ( .A(n6197), .B(n6200), .Z(n6203) );
  IV U7371 ( .A(n6199), .Z(n6200) );
  NAND U7372 ( .A(n6204), .B(n6205), .Z(n6199) );
  OR U7373 ( .A(n6206), .B(n6207), .Z(n6205) );
  OR U7374 ( .A(n6208), .B(n6209), .Z(n6204) );
  NAND U7375 ( .A(n6210), .B(n6211), .Z(n6197) );
  OR U7376 ( .A(n6212), .B(n6213), .Z(n6211) );
  OR U7377 ( .A(n6214), .B(n6215), .Z(n6210) );
  NOR U7378 ( .A(n6216), .B(n6217), .Z(n6198) );
  ANDN U7379 ( .B(n6218), .A(n6219), .Z(n6192) );
  XNOR U7380 ( .A(n6185), .B(n6220), .Z(n6191) );
  XNOR U7381 ( .A(n6184), .B(n6186), .Z(n6220) );
  NAND U7382 ( .A(n6221), .B(n6222), .Z(n6186) );
  OR U7383 ( .A(n6223), .B(n6224), .Z(n6222) );
  OR U7384 ( .A(n6225), .B(n6226), .Z(n6221) );
  NAND U7385 ( .A(n6227), .B(n6228), .Z(n6184) );
  OR U7386 ( .A(n6229), .B(n6230), .Z(n6228) );
  OR U7387 ( .A(n6231), .B(n6232), .Z(n6227) );
  ANDN U7388 ( .B(n6233), .A(n6234), .Z(n6185) );
  IV U7389 ( .A(n6235), .Z(n6233) );
  ANDN U7390 ( .B(n6236), .A(n6237), .Z(n6177) );
  XOR U7391 ( .A(n6163), .B(n6238), .Z(n6175) );
  XOR U7392 ( .A(n6164), .B(n6165), .Z(n6238) );
  XOR U7393 ( .A(n6170), .B(n6239), .Z(n6165) );
  XOR U7394 ( .A(n6169), .B(n6172), .Z(n6239) );
  IV U7395 ( .A(n6171), .Z(n6172) );
  NAND U7396 ( .A(n6240), .B(n6241), .Z(n6171) );
  OR U7397 ( .A(n6242), .B(n6243), .Z(n6241) );
  OR U7398 ( .A(n6244), .B(n6245), .Z(n6240) );
  NAND U7399 ( .A(n6246), .B(n6247), .Z(n6169) );
  OR U7400 ( .A(n6248), .B(n6249), .Z(n6247) );
  OR U7401 ( .A(n6250), .B(n6251), .Z(n6246) );
  NOR U7402 ( .A(n6252), .B(n6253), .Z(n6170) );
  ANDN U7403 ( .B(n6254), .A(n6255), .Z(n6164) );
  IV U7404 ( .A(n6256), .Z(n6254) );
  XNOR U7405 ( .A(n6157), .B(n6257), .Z(n6163) );
  XNOR U7406 ( .A(n6156), .B(n6158), .Z(n6257) );
  NAND U7407 ( .A(n6258), .B(n6259), .Z(n6158) );
  OR U7408 ( .A(n6260), .B(n6261), .Z(n6259) );
  OR U7409 ( .A(n6262), .B(n6263), .Z(n6258) );
  NAND U7410 ( .A(n6264), .B(n6265), .Z(n6156) );
  OR U7411 ( .A(n6266), .B(n6267), .Z(n6265) );
  OR U7412 ( .A(n6268), .B(n6269), .Z(n6264) );
  ANDN U7413 ( .B(n6270), .A(n6271), .Z(n6157) );
  IV U7414 ( .A(n6272), .Z(n6270) );
  XNOR U7415 ( .A(n6237), .B(n6236), .Z(N5824) );
  XOR U7416 ( .A(n6256), .B(n6255), .Z(n6236) );
  XNOR U7417 ( .A(n6271), .B(n6272), .Z(n6255) );
  XNOR U7418 ( .A(n6266), .B(n6267), .Z(n6272) );
  XNOR U7419 ( .A(n6268), .B(n6269), .Z(n6267) );
  XNOR U7420 ( .A(y[100]), .B(x[100]), .Z(n6269) );
  XNOR U7421 ( .A(y[101]), .B(x[101]), .Z(n6268) );
  XNOR U7422 ( .A(y[99]), .B(x[99]), .Z(n6266) );
  XNOR U7423 ( .A(n6260), .B(n6261), .Z(n6271) );
  XNOR U7424 ( .A(y[96]), .B(x[96]), .Z(n6261) );
  XNOR U7425 ( .A(n6262), .B(n6263), .Z(n6260) );
  XNOR U7426 ( .A(y[97]), .B(x[97]), .Z(n6263) );
  XNOR U7427 ( .A(y[98]), .B(x[98]), .Z(n6262) );
  XNOR U7428 ( .A(n6253), .B(n6252), .Z(n6256) );
  XNOR U7429 ( .A(n6248), .B(n6249), .Z(n6252) );
  XNOR U7430 ( .A(y[93]), .B(x[93]), .Z(n6249) );
  XNOR U7431 ( .A(n6250), .B(n6251), .Z(n6248) );
  XNOR U7432 ( .A(y[94]), .B(x[94]), .Z(n6251) );
  XNOR U7433 ( .A(y[95]), .B(x[95]), .Z(n6250) );
  XNOR U7434 ( .A(n6242), .B(n6243), .Z(n6253) );
  XNOR U7435 ( .A(y[90]), .B(x[90]), .Z(n6243) );
  XNOR U7436 ( .A(n6244), .B(n6245), .Z(n6242) );
  XNOR U7437 ( .A(y[91]), .B(x[91]), .Z(n6245) );
  XNOR U7438 ( .A(y[92]), .B(x[92]), .Z(n6244) );
  XOR U7439 ( .A(n6218), .B(n6219), .Z(n6237) );
  XNOR U7440 ( .A(n6234), .B(n6235), .Z(n6219) );
  XNOR U7441 ( .A(n6229), .B(n6230), .Z(n6235) );
  XNOR U7442 ( .A(n6231), .B(n6232), .Z(n6230) );
  XNOR U7443 ( .A(y[88]), .B(x[88]), .Z(n6232) );
  XNOR U7444 ( .A(y[89]), .B(x[89]), .Z(n6231) );
  XNOR U7445 ( .A(y[87]), .B(x[87]), .Z(n6229) );
  XNOR U7446 ( .A(n6223), .B(n6224), .Z(n6234) );
  XNOR U7447 ( .A(y[84]), .B(x[84]), .Z(n6224) );
  XNOR U7448 ( .A(n6225), .B(n6226), .Z(n6223) );
  XNOR U7449 ( .A(y[85]), .B(x[85]), .Z(n6226) );
  XNOR U7450 ( .A(y[86]), .B(x[86]), .Z(n6225) );
  XOR U7451 ( .A(n6217), .B(n6216), .Z(n6218) );
  XNOR U7452 ( .A(n6212), .B(n6213), .Z(n6216) );
  XNOR U7453 ( .A(y[81]), .B(x[81]), .Z(n6213) );
  XNOR U7454 ( .A(n6214), .B(n6215), .Z(n6212) );
  XNOR U7455 ( .A(y[82]), .B(x[82]), .Z(n6215) );
  XNOR U7456 ( .A(y[83]), .B(x[83]), .Z(n6214) );
  XNOR U7457 ( .A(n6206), .B(n6207), .Z(n6217) );
  XNOR U7458 ( .A(y[78]), .B(x[78]), .Z(n6207) );
  XNOR U7459 ( .A(n6208), .B(n6209), .Z(n6206) );
  XNOR U7460 ( .A(y[79]), .B(x[79]), .Z(n6209) );
  XNOR U7461 ( .A(y[80]), .B(x[80]), .Z(n6208) );
  NAND U7462 ( .A(n6273), .B(n6274), .Z(N5818) );
  NANDN U7463 ( .A(n6275), .B(n6276), .Z(n6274) );
  OR U7464 ( .A(n6277), .B(n6278), .Z(n6276) );
  NAND U7465 ( .A(n6277), .B(n6278), .Z(n6273) );
  XOR U7466 ( .A(n6277), .B(n6279), .Z(N5817) );
  XNOR U7467 ( .A(n6275), .B(n6278), .Z(n6279) );
  AND U7468 ( .A(n6280), .B(n6281), .Z(n6278) );
  NANDN U7469 ( .A(n6282), .B(n6283), .Z(n6281) );
  NANDN U7470 ( .A(n6284), .B(n6285), .Z(n6283) );
  NANDN U7471 ( .A(n6285), .B(n6284), .Z(n6280) );
  NAND U7472 ( .A(n6286), .B(n6287), .Z(n6275) );
  NANDN U7473 ( .A(n6288), .B(n6289), .Z(n6287) );
  OR U7474 ( .A(n6290), .B(n6291), .Z(n6289) );
  NAND U7475 ( .A(n6291), .B(n6290), .Z(n6286) );
  AND U7476 ( .A(n6292), .B(n6293), .Z(n6277) );
  NANDN U7477 ( .A(n6294), .B(n6295), .Z(n6293) );
  NANDN U7478 ( .A(n6296), .B(n6297), .Z(n6295) );
  NANDN U7479 ( .A(n6297), .B(n6296), .Z(n6292) );
  XOR U7480 ( .A(n6291), .B(n6298), .Z(N5816) );
  XOR U7481 ( .A(n6288), .B(n6290), .Z(n6298) );
  XNOR U7482 ( .A(n6284), .B(n6299), .Z(n6290) );
  XNOR U7483 ( .A(n6282), .B(n6285), .Z(n6299) );
  NAND U7484 ( .A(n6300), .B(n6301), .Z(n6285) );
  NAND U7485 ( .A(n6302), .B(n6303), .Z(n6301) );
  OR U7486 ( .A(n6304), .B(n6305), .Z(n6302) );
  NANDN U7487 ( .A(n6306), .B(n6304), .Z(n6300) );
  IV U7488 ( .A(n6305), .Z(n6306) );
  NAND U7489 ( .A(n6307), .B(n6308), .Z(n6282) );
  NAND U7490 ( .A(n6309), .B(n6310), .Z(n6308) );
  NANDN U7491 ( .A(n6311), .B(n6312), .Z(n6309) );
  NANDN U7492 ( .A(n6312), .B(n6311), .Z(n6307) );
  AND U7493 ( .A(n6313), .B(n6314), .Z(n6284) );
  NAND U7494 ( .A(n6315), .B(n6316), .Z(n6314) );
  OR U7495 ( .A(n6317), .B(n6318), .Z(n6315) );
  NANDN U7496 ( .A(n6319), .B(n6317), .Z(n6313) );
  NAND U7497 ( .A(n6320), .B(n6321), .Z(n6288) );
  NANDN U7498 ( .A(n6322), .B(n6323), .Z(n6321) );
  OR U7499 ( .A(n6324), .B(n6325), .Z(n6323) );
  NANDN U7500 ( .A(n6326), .B(n6324), .Z(n6320) );
  IV U7501 ( .A(n6325), .Z(n6326) );
  XNOR U7502 ( .A(n6296), .B(n6327), .Z(n6291) );
  XNOR U7503 ( .A(n6294), .B(n6297), .Z(n6327) );
  NAND U7504 ( .A(n6328), .B(n6329), .Z(n6297) );
  NAND U7505 ( .A(n6330), .B(n6331), .Z(n6329) );
  OR U7506 ( .A(n6332), .B(n6333), .Z(n6330) );
  NANDN U7507 ( .A(n6334), .B(n6332), .Z(n6328) );
  IV U7508 ( .A(n6333), .Z(n6334) );
  NAND U7509 ( .A(n6335), .B(n6336), .Z(n6294) );
  NAND U7510 ( .A(n6337), .B(n6338), .Z(n6336) );
  NANDN U7511 ( .A(n6339), .B(n6340), .Z(n6337) );
  NANDN U7512 ( .A(n6340), .B(n6339), .Z(n6335) );
  AND U7513 ( .A(n6341), .B(n6342), .Z(n6296) );
  NAND U7514 ( .A(n6343), .B(n6344), .Z(n6342) );
  OR U7515 ( .A(n6345), .B(n6346), .Z(n6343) );
  NANDN U7516 ( .A(n6347), .B(n6345), .Z(n6341) );
  XNOR U7517 ( .A(n6322), .B(n6348), .Z(N5815) );
  XOR U7518 ( .A(n6324), .B(n6325), .Z(n6348) );
  XNOR U7519 ( .A(n6338), .B(n6349), .Z(n6325) );
  XOR U7520 ( .A(n6339), .B(n6340), .Z(n6349) );
  XOR U7521 ( .A(n6345), .B(n6350), .Z(n6340) );
  XOR U7522 ( .A(n6344), .B(n6347), .Z(n6350) );
  IV U7523 ( .A(n6346), .Z(n6347) );
  NAND U7524 ( .A(n6351), .B(n6352), .Z(n6346) );
  OR U7525 ( .A(n6353), .B(n6354), .Z(n6352) );
  OR U7526 ( .A(n6355), .B(n6356), .Z(n6351) );
  NAND U7527 ( .A(n6357), .B(n6358), .Z(n6344) );
  OR U7528 ( .A(n6359), .B(n6360), .Z(n6358) );
  OR U7529 ( .A(n6361), .B(n6362), .Z(n6357) );
  NOR U7530 ( .A(n6363), .B(n6364), .Z(n6345) );
  ANDN U7531 ( .B(n6365), .A(n6366), .Z(n6339) );
  XNOR U7532 ( .A(n6332), .B(n6367), .Z(n6338) );
  XNOR U7533 ( .A(n6331), .B(n6333), .Z(n6367) );
  NAND U7534 ( .A(n6368), .B(n6369), .Z(n6333) );
  OR U7535 ( .A(n6370), .B(n6371), .Z(n6369) );
  OR U7536 ( .A(n6372), .B(n6373), .Z(n6368) );
  NAND U7537 ( .A(n6374), .B(n6375), .Z(n6331) );
  OR U7538 ( .A(n6376), .B(n6377), .Z(n6375) );
  OR U7539 ( .A(n6378), .B(n6379), .Z(n6374) );
  ANDN U7540 ( .B(n6380), .A(n6381), .Z(n6332) );
  IV U7541 ( .A(n6382), .Z(n6380) );
  ANDN U7542 ( .B(n6383), .A(n6384), .Z(n6324) );
  XOR U7543 ( .A(n6310), .B(n6385), .Z(n6322) );
  XOR U7544 ( .A(n6311), .B(n6312), .Z(n6385) );
  XOR U7545 ( .A(n6317), .B(n6386), .Z(n6312) );
  XOR U7546 ( .A(n6316), .B(n6319), .Z(n6386) );
  IV U7547 ( .A(n6318), .Z(n6319) );
  NAND U7548 ( .A(n6387), .B(n6388), .Z(n6318) );
  OR U7549 ( .A(n6389), .B(n6390), .Z(n6388) );
  OR U7550 ( .A(n6391), .B(n6392), .Z(n6387) );
  NAND U7551 ( .A(n6393), .B(n6394), .Z(n6316) );
  OR U7552 ( .A(n6395), .B(n6396), .Z(n6394) );
  OR U7553 ( .A(n6397), .B(n6398), .Z(n6393) );
  NOR U7554 ( .A(n6399), .B(n6400), .Z(n6317) );
  ANDN U7555 ( .B(n6401), .A(n6402), .Z(n6311) );
  IV U7556 ( .A(n6403), .Z(n6401) );
  XNOR U7557 ( .A(n6304), .B(n6404), .Z(n6310) );
  XNOR U7558 ( .A(n6303), .B(n6305), .Z(n6404) );
  NAND U7559 ( .A(n6405), .B(n6406), .Z(n6305) );
  OR U7560 ( .A(n6407), .B(n6408), .Z(n6406) );
  OR U7561 ( .A(n6409), .B(n6410), .Z(n6405) );
  NAND U7562 ( .A(n6411), .B(n6412), .Z(n6303) );
  OR U7563 ( .A(n6413), .B(n6414), .Z(n6412) );
  OR U7564 ( .A(n6415), .B(n6416), .Z(n6411) );
  ANDN U7565 ( .B(n6417), .A(n6418), .Z(n6304) );
  IV U7566 ( .A(n6419), .Z(n6417) );
  XNOR U7567 ( .A(n6384), .B(n6383), .Z(N5814) );
  XOR U7568 ( .A(n6403), .B(n6402), .Z(n6383) );
  XNOR U7569 ( .A(n6418), .B(n6419), .Z(n6402) );
  XNOR U7570 ( .A(n6413), .B(n6414), .Z(n6419) );
  XNOR U7571 ( .A(n6415), .B(n6416), .Z(n6414) );
  XNOR U7572 ( .A(y[76]), .B(x[76]), .Z(n6416) );
  XNOR U7573 ( .A(y[77]), .B(x[77]), .Z(n6415) );
  XNOR U7574 ( .A(y[75]), .B(x[75]), .Z(n6413) );
  XNOR U7575 ( .A(n6407), .B(n6408), .Z(n6418) );
  XNOR U7576 ( .A(y[72]), .B(x[72]), .Z(n6408) );
  XNOR U7577 ( .A(n6409), .B(n6410), .Z(n6407) );
  XNOR U7578 ( .A(y[73]), .B(x[73]), .Z(n6410) );
  XNOR U7579 ( .A(y[74]), .B(x[74]), .Z(n6409) );
  XNOR U7580 ( .A(n6400), .B(n6399), .Z(n6403) );
  XNOR U7581 ( .A(n6395), .B(n6396), .Z(n6399) );
  XNOR U7582 ( .A(y[69]), .B(x[69]), .Z(n6396) );
  XNOR U7583 ( .A(n6397), .B(n6398), .Z(n6395) );
  XNOR U7584 ( .A(y[70]), .B(x[70]), .Z(n6398) );
  XNOR U7585 ( .A(y[71]), .B(x[71]), .Z(n6397) );
  XNOR U7586 ( .A(n6389), .B(n6390), .Z(n6400) );
  XNOR U7587 ( .A(y[66]), .B(x[66]), .Z(n6390) );
  XNOR U7588 ( .A(n6391), .B(n6392), .Z(n6389) );
  XNOR U7589 ( .A(y[67]), .B(x[67]), .Z(n6392) );
  XNOR U7590 ( .A(y[68]), .B(x[68]), .Z(n6391) );
  XOR U7591 ( .A(n6365), .B(n6366), .Z(n6384) );
  XNOR U7592 ( .A(n6381), .B(n6382), .Z(n6366) );
  XNOR U7593 ( .A(n6376), .B(n6377), .Z(n6382) );
  XNOR U7594 ( .A(n6378), .B(n6379), .Z(n6377) );
  XNOR U7595 ( .A(y[64]), .B(x[64]), .Z(n6379) );
  XNOR U7596 ( .A(y[65]), .B(x[65]), .Z(n6378) );
  XNOR U7597 ( .A(y[63]), .B(x[63]), .Z(n6376) );
  XNOR U7598 ( .A(n6370), .B(n6371), .Z(n6381) );
  XNOR U7599 ( .A(y[60]), .B(x[60]), .Z(n6371) );
  XNOR U7600 ( .A(n6372), .B(n6373), .Z(n6370) );
  XNOR U7601 ( .A(y[61]), .B(x[61]), .Z(n6373) );
  XNOR U7602 ( .A(y[62]), .B(x[62]), .Z(n6372) );
  XOR U7603 ( .A(n6364), .B(n6363), .Z(n6365) );
  XNOR U7604 ( .A(n6359), .B(n6360), .Z(n6363) );
  XNOR U7605 ( .A(y[57]), .B(x[57]), .Z(n6360) );
  XNOR U7606 ( .A(n6361), .B(n6362), .Z(n6359) );
  XNOR U7607 ( .A(y[58]), .B(x[58]), .Z(n6362) );
  XNOR U7608 ( .A(y[59]), .B(x[59]), .Z(n6361) );
  XNOR U7609 ( .A(n6353), .B(n6354), .Z(n6364) );
  XNOR U7610 ( .A(y[54]), .B(x[54]), .Z(n6354) );
  XNOR U7611 ( .A(n6355), .B(n6356), .Z(n6353) );
  XNOR U7612 ( .A(y[55]), .B(x[55]), .Z(n6356) );
  XNOR U7613 ( .A(y[56]), .B(x[56]), .Z(n6355) );
  NAND U7614 ( .A(n6420), .B(n6421), .Z(N5808) );
  NANDN U7615 ( .A(n6422), .B(n6423), .Z(n6421) );
  OR U7616 ( .A(n6424), .B(n6425), .Z(n6423) );
  NAND U7617 ( .A(n6424), .B(n6425), .Z(n6420) );
  XOR U7618 ( .A(n6424), .B(n6426), .Z(N5807) );
  XNOR U7619 ( .A(n6422), .B(n6425), .Z(n6426) );
  AND U7620 ( .A(n6427), .B(n6428), .Z(n6425) );
  NANDN U7621 ( .A(n6429), .B(n6430), .Z(n6428) );
  NANDN U7622 ( .A(n6431), .B(n6432), .Z(n6430) );
  NANDN U7623 ( .A(n6432), .B(n6431), .Z(n6427) );
  NAND U7624 ( .A(n6433), .B(n6434), .Z(n6422) );
  NANDN U7625 ( .A(n6435), .B(n6436), .Z(n6434) );
  OR U7626 ( .A(n6437), .B(n6438), .Z(n6436) );
  NAND U7627 ( .A(n6438), .B(n6437), .Z(n6433) );
  AND U7628 ( .A(n6439), .B(n6440), .Z(n6424) );
  NANDN U7629 ( .A(n6441), .B(n6442), .Z(n6440) );
  NANDN U7630 ( .A(n6443), .B(n6444), .Z(n6442) );
  NANDN U7631 ( .A(n6444), .B(n6443), .Z(n6439) );
  XOR U7632 ( .A(n6438), .B(n6445), .Z(N5806) );
  XOR U7633 ( .A(n6435), .B(n6437), .Z(n6445) );
  XNOR U7634 ( .A(n6431), .B(n6446), .Z(n6437) );
  XNOR U7635 ( .A(n6429), .B(n6432), .Z(n6446) );
  NAND U7636 ( .A(n6447), .B(n6448), .Z(n6432) );
  NAND U7637 ( .A(n6449), .B(n6450), .Z(n6448) );
  OR U7638 ( .A(n6451), .B(n6452), .Z(n6449) );
  NANDN U7639 ( .A(n6453), .B(n6451), .Z(n6447) );
  IV U7640 ( .A(n6452), .Z(n6453) );
  NAND U7641 ( .A(n6454), .B(n6455), .Z(n6429) );
  NAND U7642 ( .A(n6456), .B(n6457), .Z(n6455) );
  NANDN U7643 ( .A(n6458), .B(n6459), .Z(n6456) );
  NANDN U7644 ( .A(n6459), .B(n6458), .Z(n6454) );
  AND U7645 ( .A(n6460), .B(n6461), .Z(n6431) );
  NAND U7646 ( .A(n6462), .B(n6463), .Z(n6461) );
  OR U7647 ( .A(n6464), .B(n6465), .Z(n6462) );
  NANDN U7648 ( .A(n6466), .B(n6464), .Z(n6460) );
  NAND U7649 ( .A(n6467), .B(n6468), .Z(n6435) );
  NANDN U7650 ( .A(n6469), .B(n6470), .Z(n6468) );
  OR U7651 ( .A(n6471), .B(n6472), .Z(n6470) );
  NANDN U7652 ( .A(n6473), .B(n6471), .Z(n6467) );
  IV U7653 ( .A(n6472), .Z(n6473) );
  XNOR U7654 ( .A(n6443), .B(n6474), .Z(n6438) );
  XNOR U7655 ( .A(n6441), .B(n6444), .Z(n6474) );
  NAND U7656 ( .A(n6475), .B(n6476), .Z(n6444) );
  NAND U7657 ( .A(n6477), .B(n6478), .Z(n6476) );
  OR U7658 ( .A(n6479), .B(n6480), .Z(n6477) );
  NANDN U7659 ( .A(n6481), .B(n6479), .Z(n6475) );
  IV U7660 ( .A(n6480), .Z(n6481) );
  NAND U7661 ( .A(n6482), .B(n6483), .Z(n6441) );
  NAND U7662 ( .A(n6484), .B(n6485), .Z(n6483) );
  NANDN U7663 ( .A(n6486), .B(n6487), .Z(n6484) );
  NANDN U7664 ( .A(n6487), .B(n6486), .Z(n6482) );
  AND U7665 ( .A(n6488), .B(n6489), .Z(n6443) );
  NAND U7666 ( .A(n6490), .B(n6491), .Z(n6489) );
  OR U7667 ( .A(n6492), .B(n6493), .Z(n6490) );
  NANDN U7668 ( .A(n6494), .B(n6492), .Z(n6488) );
  XNOR U7669 ( .A(n6469), .B(n6495), .Z(N5805) );
  XOR U7670 ( .A(n6471), .B(n6472), .Z(n6495) );
  XNOR U7671 ( .A(n6485), .B(n6496), .Z(n6472) );
  XOR U7672 ( .A(n6486), .B(n6487), .Z(n6496) );
  XOR U7673 ( .A(n6492), .B(n6497), .Z(n6487) );
  XOR U7674 ( .A(n6491), .B(n6494), .Z(n6497) );
  IV U7675 ( .A(n6493), .Z(n6494) );
  NAND U7676 ( .A(n6498), .B(n6499), .Z(n6493) );
  OR U7677 ( .A(n6500), .B(n6501), .Z(n6499) );
  OR U7678 ( .A(n6502), .B(n6503), .Z(n6498) );
  NAND U7679 ( .A(n6504), .B(n6505), .Z(n6491) );
  OR U7680 ( .A(n6506), .B(n6507), .Z(n6505) );
  OR U7681 ( .A(n6508), .B(n6509), .Z(n6504) );
  NOR U7682 ( .A(n6510), .B(n6511), .Z(n6492) );
  ANDN U7683 ( .B(n6512), .A(n6513), .Z(n6486) );
  XNOR U7684 ( .A(n6479), .B(n6514), .Z(n6485) );
  XNOR U7685 ( .A(n6478), .B(n6480), .Z(n6514) );
  NAND U7686 ( .A(n6515), .B(n6516), .Z(n6480) );
  OR U7687 ( .A(n6517), .B(n6518), .Z(n6516) );
  OR U7688 ( .A(n6519), .B(n6520), .Z(n6515) );
  NAND U7689 ( .A(n6521), .B(n6522), .Z(n6478) );
  OR U7690 ( .A(n6523), .B(n6524), .Z(n6522) );
  OR U7691 ( .A(n6525), .B(n6526), .Z(n6521) );
  ANDN U7692 ( .B(n6527), .A(n6528), .Z(n6479) );
  IV U7693 ( .A(n6529), .Z(n6527) );
  ANDN U7694 ( .B(n6530), .A(n6531), .Z(n6471) );
  XOR U7695 ( .A(n6457), .B(n6532), .Z(n6469) );
  XOR U7696 ( .A(n6458), .B(n6459), .Z(n6532) );
  XOR U7697 ( .A(n6464), .B(n6533), .Z(n6459) );
  XOR U7698 ( .A(n6463), .B(n6466), .Z(n6533) );
  IV U7699 ( .A(n6465), .Z(n6466) );
  NAND U7700 ( .A(n6534), .B(n6535), .Z(n6465) );
  OR U7701 ( .A(n6536), .B(n6537), .Z(n6535) );
  OR U7702 ( .A(n6538), .B(n6539), .Z(n6534) );
  NAND U7703 ( .A(n6540), .B(n6541), .Z(n6463) );
  OR U7704 ( .A(n6542), .B(n6543), .Z(n6541) );
  OR U7705 ( .A(n6544), .B(n6545), .Z(n6540) );
  NOR U7706 ( .A(n6546), .B(n6547), .Z(n6464) );
  ANDN U7707 ( .B(n6548), .A(n6549), .Z(n6458) );
  IV U7708 ( .A(n6550), .Z(n6548) );
  XNOR U7709 ( .A(n6451), .B(n6551), .Z(n6457) );
  XNOR U7710 ( .A(n6450), .B(n6452), .Z(n6551) );
  NAND U7711 ( .A(n6552), .B(n6553), .Z(n6452) );
  OR U7712 ( .A(n6554), .B(n6555), .Z(n6553) );
  OR U7713 ( .A(n6556), .B(n6557), .Z(n6552) );
  NAND U7714 ( .A(n6558), .B(n6559), .Z(n6450) );
  OR U7715 ( .A(n6560), .B(n6561), .Z(n6559) );
  OR U7716 ( .A(n6562), .B(n6563), .Z(n6558) );
  ANDN U7717 ( .B(n6564), .A(n6565), .Z(n6451) );
  IV U7718 ( .A(n6566), .Z(n6564) );
  XNOR U7719 ( .A(n6531), .B(n6530), .Z(N5804) );
  XOR U7720 ( .A(n6550), .B(n6549), .Z(n6530) );
  XNOR U7721 ( .A(n6565), .B(n6566), .Z(n6549) );
  XNOR U7722 ( .A(n6560), .B(n6561), .Z(n6566) );
  XNOR U7723 ( .A(n6562), .B(n6563), .Z(n6561) );
  XNOR U7724 ( .A(y[52]), .B(x[52]), .Z(n6563) );
  XNOR U7725 ( .A(y[53]), .B(x[53]), .Z(n6562) );
  XNOR U7726 ( .A(y[51]), .B(x[51]), .Z(n6560) );
  XNOR U7727 ( .A(n6554), .B(n6555), .Z(n6565) );
  XNOR U7728 ( .A(y[48]), .B(x[48]), .Z(n6555) );
  XNOR U7729 ( .A(n6556), .B(n6557), .Z(n6554) );
  XNOR U7730 ( .A(y[49]), .B(x[49]), .Z(n6557) );
  XNOR U7731 ( .A(y[50]), .B(x[50]), .Z(n6556) );
  XNOR U7732 ( .A(n6547), .B(n6546), .Z(n6550) );
  XNOR U7733 ( .A(n6542), .B(n6543), .Z(n6546) );
  XNOR U7734 ( .A(y[45]), .B(x[45]), .Z(n6543) );
  XNOR U7735 ( .A(n6544), .B(n6545), .Z(n6542) );
  XNOR U7736 ( .A(y[46]), .B(x[46]), .Z(n6545) );
  XNOR U7737 ( .A(y[47]), .B(x[47]), .Z(n6544) );
  XNOR U7738 ( .A(n6536), .B(n6537), .Z(n6547) );
  XNOR U7739 ( .A(y[42]), .B(x[42]), .Z(n6537) );
  XNOR U7740 ( .A(n6538), .B(n6539), .Z(n6536) );
  XNOR U7741 ( .A(y[43]), .B(x[43]), .Z(n6539) );
  XNOR U7742 ( .A(y[44]), .B(x[44]), .Z(n6538) );
  XOR U7743 ( .A(n6512), .B(n6513), .Z(n6531) );
  XNOR U7744 ( .A(n6528), .B(n6529), .Z(n6513) );
  XNOR U7745 ( .A(n6523), .B(n6524), .Z(n6529) );
  XNOR U7746 ( .A(n6525), .B(n6526), .Z(n6524) );
  XNOR U7747 ( .A(y[40]), .B(x[40]), .Z(n6526) );
  XNOR U7748 ( .A(y[41]), .B(x[41]), .Z(n6525) );
  XNOR U7749 ( .A(y[39]), .B(x[39]), .Z(n6523) );
  XNOR U7750 ( .A(n6517), .B(n6518), .Z(n6528) );
  XNOR U7751 ( .A(y[36]), .B(x[36]), .Z(n6518) );
  XNOR U7752 ( .A(n6519), .B(n6520), .Z(n6517) );
  XNOR U7753 ( .A(y[37]), .B(x[37]), .Z(n6520) );
  XNOR U7754 ( .A(y[38]), .B(x[38]), .Z(n6519) );
  XOR U7755 ( .A(n6511), .B(n6510), .Z(n6512) );
  XNOR U7756 ( .A(n6506), .B(n6507), .Z(n6510) );
  XNOR U7757 ( .A(y[33]), .B(x[33]), .Z(n6507) );
  XNOR U7758 ( .A(n6508), .B(n6509), .Z(n6506) );
  XNOR U7759 ( .A(y[34]), .B(x[34]), .Z(n6509) );
  XNOR U7760 ( .A(y[35]), .B(x[35]), .Z(n6508) );
  XNOR U7761 ( .A(n6500), .B(n6501), .Z(n6511) );
  XNOR U7762 ( .A(y[30]), .B(x[30]), .Z(n6501) );
  XNOR U7763 ( .A(n6502), .B(n6503), .Z(n6500) );
  XNOR U7764 ( .A(y[31]), .B(x[31]), .Z(n6503) );
  XNOR U7765 ( .A(y[32]), .B(x[32]), .Z(n6502) );
  NAND U7766 ( .A(n6567), .B(n6568), .Z(N5798) );
  NANDN U7767 ( .A(n6569), .B(n6570), .Z(n6568) );
  OR U7768 ( .A(n6571), .B(n6572), .Z(n6570) );
  NAND U7769 ( .A(n6571), .B(n6572), .Z(n6567) );
  XOR U7770 ( .A(n6571), .B(n6573), .Z(N5797) );
  XNOR U7771 ( .A(n6569), .B(n6572), .Z(n6573) );
  AND U7772 ( .A(n6574), .B(n6575), .Z(n6572) );
  NANDN U7773 ( .A(n6576), .B(n6577), .Z(n6575) );
  NANDN U7774 ( .A(n6578), .B(n6579), .Z(n6577) );
  NANDN U7775 ( .A(n6579), .B(n6578), .Z(n6574) );
  NAND U7776 ( .A(n6580), .B(n6581), .Z(n6569) );
  NANDN U7777 ( .A(n6582), .B(n6583), .Z(n6581) );
  OR U7778 ( .A(n6584), .B(n6585), .Z(n6583) );
  NAND U7779 ( .A(n6585), .B(n6584), .Z(n6580) );
  AND U7780 ( .A(n6586), .B(n6587), .Z(n6571) );
  NANDN U7781 ( .A(n6588), .B(n6589), .Z(n6587) );
  NANDN U7782 ( .A(n6590), .B(n6591), .Z(n6589) );
  NANDN U7783 ( .A(n6591), .B(n6590), .Z(n6586) );
  XOR U7784 ( .A(n6585), .B(n6592), .Z(N5796) );
  XOR U7785 ( .A(n6582), .B(n6584), .Z(n6592) );
  XNOR U7786 ( .A(n6578), .B(n6593), .Z(n6584) );
  XNOR U7787 ( .A(n6576), .B(n6579), .Z(n6593) );
  NAND U7788 ( .A(n6594), .B(n6595), .Z(n6579) );
  NAND U7789 ( .A(n6596), .B(n6597), .Z(n6595) );
  OR U7790 ( .A(n6598), .B(n6599), .Z(n6596) );
  NANDN U7791 ( .A(n6600), .B(n6598), .Z(n6594) );
  IV U7792 ( .A(n6599), .Z(n6600) );
  NAND U7793 ( .A(n6601), .B(n6602), .Z(n6576) );
  NAND U7794 ( .A(n6603), .B(n6604), .Z(n6602) );
  NANDN U7795 ( .A(n6605), .B(n6606), .Z(n6603) );
  NANDN U7796 ( .A(n6606), .B(n6605), .Z(n6601) );
  AND U7797 ( .A(n6607), .B(n6608), .Z(n6578) );
  NAND U7798 ( .A(n6609), .B(n6610), .Z(n6608) );
  OR U7799 ( .A(n6611), .B(n6612), .Z(n6609) );
  NANDN U7800 ( .A(n6613), .B(n6611), .Z(n6607) );
  NAND U7801 ( .A(n6614), .B(n6615), .Z(n6582) );
  NANDN U7802 ( .A(n6616), .B(n6617), .Z(n6615) );
  OR U7803 ( .A(n6618), .B(n6619), .Z(n6617) );
  NANDN U7804 ( .A(n6620), .B(n6618), .Z(n6614) );
  IV U7805 ( .A(n6619), .Z(n6620) );
  XNOR U7806 ( .A(n6590), .B(n6621), .Z(n6585) );
  XNOR U7807 ( .A(n6588), .B(n6591), .Z(n6621) );
  NAND U7808 ( .A(n6622), .B(n6623), .Z(n6591) );
  NAND U7809 ( .A(n6624), .B(n6625), .Z(n6623) );
  OR U7810 ( .A(n6626), .B(n6627), .Z(n6624) );
  NANDN U7811 ( .A(n6628), .B(n6626), .Z(n6622) );
  IV U7812 ( .A(n6627), .Z(n6628) );
  NAND U7813 ( .A(n6629), .B(n6630), .Z(n6588) );
  NAND U7814 ( .A(n6631), .B(n6632), .Z(n6630) );
  NANDN U7815 ( .A(n6633), .B(n6634), .Z(n6631) );
  NANDN U7816 ( .A(n6634), .B(n6633), .Z(n6629) );
  AND U7817 ( .A(n6635), .B(n6636), .Z(n6590) );
  NAND U7818 ( .A(n6637), .B(n6638), .Z(n6636) );
  OR U7819 ( .A(n6639), .B(n6640), .Z(n6637) );
  NANDN U7820 ( .A(n6641), .B(n6639), .Z(n6635) );
  IV U7821 ( .A(n6640), .Z(n6641) );
  XNOR U7822 ( .A(n6616), .B(n6642), .Z(N5795) );
  XOR U7823 ( .A(n6618), .B(n6619), .Z(n6642) );
  XNOR U7824 ( .A(n6632), .B(n6643), .Z(n6619) );
  XOR U7825 ( .A(n6633), .B(n6634), .Z(n6643) );
  XOR U7826 ( .A(n6639), .B(n6644), .Z(n6634) );
  XNOR U7827 ( .A(n6638), .B(n6640), .Z(n6644) );
  NAND U7828 ( .A(n6645), .B(n6646), .Z(n6640) );
  OR U7829 ( .A(n6647), .B(n6648), .Z(n6646) );
  IV U7830 ( .A(n6649), .Z(n6648) );
  OR U7831 ( .A(n6650), .B(n6651), .Z(n6645) );
  NAND U7832 ( .A(n6652), .B(n6653), .Z(n6638) );
  OR U7833 ( .A(n6654), .B(n6655), .Z(n6653) );
  OR U7834 ( .A(n6656), .B(n6657), .Z(n6652) );
  ANDN U7835 ( .B(n6658), .A(n6659), .Z(n6639) );
  IV U7836 ( .A(n6660), .Z(n6658) );
  NOR U7837 ( .A(n6661), .B(n6662), .Z(n6633) );
  XNOR U7838 ( .A(n6626), .B(n6663), .Z(n6632) );
  XNOR U7839 ( .A(n6625), .B(n6627), .Z(n6663) );
  NAND U7840 ( .A(n6664), .B(n6665), .Z(n6627) );
  OR U7841 ( .A(n6666), .B(n6667), .Z(n6665) );
  OR U7842 ( .A(n6668), .B(n6669), .Z(n6664) );
  NAND U7843 ( .A(n6670), .B(n6671), .Z(n6625) );
  OR U7844 ( .A(n6672), .B(n6673), .Z(n6671) );
  OR U7845 ( .A(n6674), .B(n6675), .Z(n6670) );
  ANDN U7846 ( .B(n6676), .A(n6677), .Z(n6626) );
  IV U7847 ( .A(n6678), .Z(n6676) );
  ANDN U7848 ( .B(n6679), .A(n6680), .Z(n6618) );
  XOR U7849 ( .A(n6604), .B(n6681), .Z(n6616) );
  XOR U7850 ( .A(n6605), .B(n6606), .Z(n6681) );
  XOR U7851 ( .A(n6611), .B(n6682), .Z(n6606) );
  XOR U7852 ( .A(n6610), .B(n6613), .Z(n6682) );
  IV U7853 ( .A(n6612), .Z(n6613) );
  NAND U7854 ( .A(n6683), .B(n6684), .Z(n6612) );
  OR U7855 ( .A(n6685), .B(n6686), .Z(n6684) );
  OR U7856 ( .A(n6687), .B(n6688), .Z(n6683) );
  NAND U7857 ( .A(n6689), .B(n6690), .Z(n6610) );
  OR U7858 ( .A(n6691), .B(n6692), .Z(n6690) );
  OR U7859 ( .A(n6693), .B(n6694), .Z(n6689) );
  NOR U7860 ( .A(n6695), .B(n6696), .Z(n6611) );
  ANDN U7861 ( .B(n6697), .A(n6698), .Z(n6605) );
  IV U7862 ( .A(n6699), .Z(n6697) );
  XNOR U7863 ( .A(n6598), .B(n6700), .Z(n6604) );
  XNOR U7864 ( .A(n6597), .B(n6599), .Z(n6700) );
  NAND U7865 ( .A(n6701), .B(n6702), .Z(n6599) );
  OR U7866 ( .A(n6703), .B(n6704), .Z(n6702) );
  OR U7867 ( .A(n6705), .B(n6706), .Z(n6701) );
  NAND U7868 ( .A(n6707), .B(n6708), .Z(n6597) );
  OR U7869 ( .A(n6709), .B(n6710), .Z(n6708) );
  OR U7870 ( .A(n6711), .B(n6712), .Z(n6707) );
  ANDN U7871 ( .B(n6713), .A(n6714), .Z(n6598) );
  IV U7872 ( .A(n6715), .Z(n6713) );
  XNOR U7873 ( .A(n6680), .B(n6679), .Z(N5794) );
  XOR U7874 ( .A(n6699), .B(n6698), .Z(n6679) );
  XNOR U7875 ( .A(n6714), .B(n6715), .Z(n6698) );
  XNOR U7876 ( .A(n6709), .B(n6710), .Z(n6715) );
  XNOR U7877 ( .A(n6711), .B(n6712), .Z(n6710) );
  XNOR U7878 ( .A(y[28]), .B(x[28]), .Z(n6712) );
  XNOR U7879 ( .A(y[29]), .B(x[29]), .Z(n6711) );
  XNOR U7880 ( .A(y[27]), .B(x[27]), .Z(n6709) );
  XNOR U7881 ( .A(n6703), .B(n6704), .Z(n6714) );
  XNOR U7882 ( .A(y[24]), .B(x[24]), .Z(n6704) );
  XNOR U7883 ( .A(n6705), .B(n6706), .Z(n6703) );
  XNOR U7884 ( .A(y[25]), .B(x[25]), .Z(n6706) );
  XNOR U7885 ( .A(y[26]), .B(x[26]), .Z(n6705) );
  XNOR U7886 ( .A(n6696), .B(n6695), .Z(n6699) );
  XNOR U7887 ( .A(n6691), .B(n6692), .Z(n6695) );
  XNOR U7888 ( .A(y[21]), .B(x[21]), .Z(n6692) );
  XNOR U7889 ( .A(n6693), .B(n6694), .Z(n6691) );
  XNOR U7890 ( .A(y[22]), .B(x[22]), .Z(n6694) );
  XNOR U7891 ( .A(y[23]), .B(x[23]), .Z(n6693) );
  XNOR U7892 ( .A(n6685), .B(n6686), .Z(n6696) );
  XNOR U7893 ( .A(y[18]), .B(x[18]), .Z(n6686) );
  XNOR U7894 ( .A(n6687), .B(n6688), .Z(n6685) );
  XNOR U7895 ( .A(y[19]), .B(x[19]), .Z(n6688) );
  XNOR U7896 ( .A(y[20]), .B(x[20]), .Z(n6687) );
  XNOR U7897 ( .A(n6661), .B(n6662), .Z(n6680) );
  XNOR U7898 ( .A(n6677), .B(n6678), .Z(n6662) );
  XNOR U7899 ( .A(n6672), .B(n6673), .Z(n6678) );
  XNOR U7900 ( .A(n6674), .B(n6675), .Z(n6673) );
  XNOR U7901 ( .A(y[16]), .B(x[16]), .Z(n6675) );
  XNOR U7902 ( .A(y[17]), .B(x[17]), .Z(n6674) );
  XNOR U7903 ( .A(y[15]), .B(x[15]), .Z(n6672) );
  XNOR U7904 ( .A(n6666), .B(n6667), .Z(n6677) );
  XNOR U7905 ( .A(y[12]), .B(x[12]), .Z(n6667) );
  XNOR U7906 ( .A(n6668), .B(n6669), .Z(n6666) );
  XNOR U7907 ( .A(y[13]), .B(x[13]), .Z(n6669) );
  XNOR U7908 ( .A(y[14]), .B(x[14]), .Z(n6668) );
  XNOR U7909 ( .A(n6660), .B(n6659), .Z(n6661) );
  XNOR U7910 ( .A(n6654), .B(n6655), .Z(n6659) );
  XNOR U7911 ( .A(y[9]), .B(x[9]), .Z(n6655) );
  XNOR U7912 ( .A(n6656), .B(n6657), .Z(n6654) );
  XNOR U7913 ( .A(y[10]), .B(x[10]), .Z(n6657) );
  XNOR U7914 ( .A(y[11]), .B(x[11]), .Z(n6656) );
  XOR U7915 ( .A(n6647), .B(n6649), .Z(n6660) );
  XOR U7916 ( .A(n6650), .B(n6651), .Z(n6649) );
  XNOR U7917 ( .A(y[7]), .B(x[7]), .Z(n6651) );
  XNOR U7918 ( .A(y[8]), .B(x[8]), .Z(n6650) );
  XNOR U7919 ( .A(y[6]), .B(x[6]), .Z(n6647) );
  ANDN U7920 ( .B(n6716), .A(n6717), .Z(N5788) );
  XNOR U7921 ( .A(n6717), .B(n6716), .Z(N5787) );
  ANDN U7922 ( .B(n6718), .A(n6719), .Z(n6716) );
  NAND U7923 ( .A(n6720), .B(n6721), .Z(n6717) );
  NANDN U7924 ( .A(n6722), .B(n6723), .Z(n6721) );
  OR U7925 ( .A(n6724), .B(n6725), .Z(n6723) );
  NAND U7926 ( .A(n6724), .B(n6725), .Z(n6720) );
  XNOR U7927 ( .A(n6724), .B(n6726), .Z(N5786) );
  XNOR U7928 ( .A(n6722), .B(n6725), .Z(n6726) );
  AND U7929 ( .A(n6727), .B(n6728), .Z(n6725) );
  NAND U7930 ( .A(n6729), .B(n6730), .Z(n6728) );
  OR U7931 ( .A(n6731), .B(n6732), .Z(n6729) );
  NANDN U7932 ( .A(n6733), .B(n6731), .Z(n6727) );
  IV U7933 ( .A(n6732), .Z(n6733) );
  NAND U7934 ( .A(n6734), .B(n6735), .Z(n6722) );
  NANDN U7935 ( .A(n6736), .B(n6737), .Z(n6735) );
  OR U7936 ( .A(n6738), .B(n6739), .Z(n6737) );
  NAND U7937 ( .A(n6739), .B(n6738), .Z(n6734) );
  XOR U7938 ( .A(n6719), .B(n6718), .Z(n6724) );
  NAND U7939 ( .A(n6740), .B(n6741), .Z(n6718) );
  OR U7940 ( .A(n6742), .B(n6743), .Z(n6741) );
  OR U7941 ( .A(n6744), .B(n6745), .Z(n6740) );
  AND U7942 ( .A(n6746), .B(n6747), .Z(n6719) );
  NAND U7943 ( .A(n6748), .B(n6749), .Z(n6747) );
  NAND U7944 ( .A(n6750), .B(n6751), .Z(n6748) );
  OR U7945 ( .A(n6750), .B(n6751), .Z(n6746) );
  XNOR U7946 ( .A(n6736), .B(n6752), .Z(N5785) );
  XOR U7947 ( .A(n6738), .B(n6739), .Z(n6752) );
  XNOR U7948 ( .A(n6731), .B(n6753), .Z(n6739) );
  XNOR U7949 ( .A(n6730), .B(n6732), .Z(n6753) );
  NAND U7950 ( .A(n6754), .B(n6755), .Z(n6732) );
  OR U7951 ( .A(n6756), .B(n6757), .Z(n6755) );
  OR U7952 ( .A(n6758), .B(n6759), .Z(n6754) );
  NAND U7953 ( .A(n6760), .B(n6761), .Z(n6730) );
  OR U7954 ( .A(n6762), .B(n6763), .Z(n6761) );
  OR U7955 ( .A(n6764), .B(n6765), .Z(n6760) );
  ANDN U7956 ( .B(n6766), .A(n6767), .Z(n6731) );
  IV U7957 ( .A(n6768), .Z(n6766) );
  ANDN U7958 ( .B(n6769), .A(n6770), .Z(n6738) );
  XNOR U7959 ( .A(n6749), .B(n6771), .Z(n6736) );
  XOR U7960 ( .A(n6751), .B(n6750), .Z(n6771) );
  OR U7961 ( .A(n6772), .B(n6773), .Z(n6750) );
  AND U7962 ( .A(n6774), .B(n6775), .Z(n6751) );
  OR U7963 ( .A(n6776), .B(n6777), .Z(n6775) );
  OR U7964 ( .A(n6778), .B(n6779), .Z(n6774) );
  XOR U7965 ( .A(n6742), .B(n6743), .Z(n6749) );
  XOR U7966 ( .A(n6780), .B(n6744), .Z(n6743) );
  AND U7967 ( .A(n6781), .B(n6782), .Z(n6744) );
  OR U7968 ( .A(n6783), .B(n6784), .Z(n6782) );
  OR U7969 ( .A(n6785), .B(n6786), .Z(n6781) );
  IV U7970 ( .A(n6745), .Z(n6780) );
  AND U7971 ( .A(n6787), .B(n6788), .Z(n6745) );
  NANDN U7972 ( .A(n6789), .B(n6790), .Z(n6788) );
  OR U7973 ( .A(n6791), .B(n6792), .Z(n6787) );
  AND U7974 ( .A(n6793), .B(n6794), .Z(n6742) );
  NANDN U7975 ( .A(n6795), .B(n6796), .Z(n6794) );
  NANDN U7976 ( .A(n6797), .B(n6798), .Z(n6793) );
  XNOR U7977 ( .A(n6770), .B(n6769), .Z(N5784) );
  XOR U7978 ( .A(n6773), .B(n6772), .Z(n6769) );
  XOR U7979 ( .A(n6795), .B(n6796), .Z(n6772) );
  XNOR U7980 ( .A(n6797), .B(n6798), .Z(n6796) );
  XOR U7981 ( .A(n6784), .B(n6783), .Z(n6798) );
  XNOR U7982 ( .A(y[0]), .B(x[0]), .Z(n6783) );
  XNOR U7983 ( .A(n6786), .B(n6785), .Z(n6784) );
  XNOR U7984 ( .A(y[1]), .B(x[1]), .Z(n6785) );
  XNOR U7985 ( .A(y[2]), .B(x[2]), .Z(n6786) );
  XOR U7986 ( .A(n6790), .B(n6789), .Z(n6797) );
  XNOR U7987 ( .A(y[3]), .B(x[3]), .Z(n6789) );
  XOR U7988 ( .A(n6792), .B(n6791), .Z(n6790) );
  XNOR U7989 ( .A(y[4]), .B(x[4]), .Z(n6791) );
  XNOR U7990 ( .A(y[5]), .B(x[5]), .Z(n6792) );
  XNOR U7991 ( .A(y[999]), .B(x[999]), .Z(n6795) );
  XNOR U7992 ( .A(n6776), .B(n6777), .Z(n6773) );
  XNOR U7993 ( .A(y[996]), .B(x[996]), .Z(n6777) );
  XNOR U7994 ( .A(n6778), .B(n6779), .Z(n6776) );
  XNOR U7995 ( .A(y[997]), .B(x[997]), .Z(n6779) );
  XNOR U7996 ( .A(y[998]), .B(x[998]), .Z(n6778) );
  XNOR U7997 ( .A(n6767), .B(n6768), .Z(n6770) );
  XNOR U7998 ( .A(n6762), .B(n6763), .Z(n6768) );
  XNOR U7999 ( .A(n6764), .B(n6765), .Z(n6763) );
  XNOR U8000 ( .A(y[994]), .B(x[994]), .Z(n6765) );
  XNOR U8001 ( .A(y[995]), .B(x[995]), .Z(n6764) );
  XNOR U8002 ( .A(y[993]), .B(x[993]), .Z(n6762) );
  XNOR U8003 ( .A(n6756), .B(n6757), .Z(n6767) );
  XNOR U8004 ( .A(y[990]), .B(x[990]), .Z(n6757) );
  XNOR U8005 ( .A(n6758), .B(n6759), .Z(n6756) );
  XNOR U8006 ( .A(y[991]), .B(x[991]), .Z(n6759) );
  XNOR U8007 ( .A(y[992]), .B(x[992]), .Z(n6758) );
endmodule

