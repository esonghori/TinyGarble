
module modmult_N256_CC512 ( clk, rst, start, x, y, n, o );
  input [255:0] x;
  input [255:0] y;
  input [255:0] n;
  output [255:0] o;
  input clk, rst, start;


endmodule


module modexp_2N_NN_N256_CC262144 ( clk, rst, m, e, n, c );
  input [255:0] m;
  input [255:0] e;
  input [255:0] n;
  output [255:0] c;
  input clk, rst;
  wire   init, mul_pow, first_one, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012;
  wire   [511:0] start_in;
  wire   [511:0] start_reg;
  wire   [255:0] ereg;
  wire   [255:0] o;
  wire   [255:0] creg;
  wire   [255:0] x;
  wire   [255:0] y;

  modmult_N256_CC512 modmult_1 ( .clk(clk), .rst(rst), .start(start_in[0]), 
        .x(x), .y(y), .n(n), .o(o) );
  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \start_reg_reg[0]  ( .D(start_in[511]), .CLK(clk), .RST(rst), .Q(
        start_reg[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .Q(
        start_reg[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .Q(
        start_reg[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .Q(
        start_reg[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .Q(
        start_reg[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .Q(
        start_reg[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .Q(
        start_reg[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .Q(
        start_reg[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .Q(
        start_reg[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .Q(
        start_reg[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .Q(
        start_reg[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .Q(
        start_reg[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .Q(
        start_reg[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .Q(
        start_reg[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .Q(
        start_reg[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .Q(
        start_reg[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .Q(
        start_reg[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .Q(
        start_reg[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .Q(
        start_reg[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .Q(
        start_reg[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .Q(
        start_reg[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .Q(
        start_reg[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .Q(
        start_reg[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .Q(
        start_reg[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .Q(
        start_reg[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .Q(
        start_reg[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .Q(
        start_reg[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .Q(
        start_reg[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .Q(
        start_reg[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .Q(
        start_reg[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .Q(
        start_reg[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .Q(
        start_reg[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .Q(
        start_reg[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .Q(
        start_reg[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .Q(
        start_reg[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .Q(
        start_reg[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .Q(
        start_reg[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .Q(
        start_reg[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .Q(
        start_reg[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .Q(
        start_reg[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .Q(
        start_reg[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .Q(
        start_reg[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .Q(
        start_reg[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .Q(
        start_reg[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .Q(
        start_reg[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .Q(
        start_reg[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .Q(
        start_reg[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .Q(
        start_reg[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .Q(
        start_reg[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .Q(
        start_reg[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .Q(
        start_reg[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .Q(
        start_reg[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .Q(
        start_reg[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .Q(
        start_reg[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .Q(
        start_reg[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .Q(
        start_reg[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .Q(
        start_reg[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .Q(
        start_reg[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .Q(
        start_reg[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .Q(
        start_reg[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .Q(
        start_reg[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .Q(
        start_reg[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .Q(
        start_reg[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .Q(
        start_reg[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .Q(
        start_reg[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .Q(
        start_reg[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .Q(
        start_reg[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .Q(
        start_reg[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .Q(
        start_reg[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .Q(
        start_reg[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .Q(
        start_reg[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .Q(
        start_reg[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .Q(
        start_reg[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .Q(
        start_reg[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .Q(
        start_reg[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .Q(
        start_reg[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .Q(
        start_reg[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .Q(
        start_reg[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .Q(
        start_reg[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .Q(
        start_reg[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .Q(
        start_reg[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .Q(
        start_reg[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .Q(
        start_reg[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .Q(
        start_reg[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .Q(
        start_reg[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .Q(
        start_reg[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .Q(
        start_reg[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .Q(
        start_reg[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .Q(
        start_reg[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .Q(
        start_reg[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .Q(
        start_reg[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .Q(
        start_reg[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .Q(
        start_reg[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .Q(
        start_reg[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .Q(
        start_reg[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .Q(
        start_reg[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .Q(
        start_reg[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .Q(
        start_reg[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .Q(
        start_reg[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .Q(
        start_reg[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .Q(
        start_reg[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .Q(
        start_reg[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .Q(
        start_reg[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .Q(
        start_reg[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .Q(
        start_reg[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .Q(
        start_reg[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .Q(
        start_reg[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .Q(
        start_reg[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .Q(
        start_reg[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .Q(
        start_reg[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .Q(
        start_reg[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .Q(
        start_reg[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .Q(
        start_reg[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .Q(
        start_reg[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .Q(
        start_reg[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .Q(
        start_reg[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .Q(
        start_reg[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .Q(
        start_reg[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .Q(
        start_reg[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .Q(
        start_reg[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .Q(
        start_reg[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .Q(
        start_reg[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .Q(
        start_reg[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .Q(
        start_reg[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .Q(
        start_reg[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .Q(
        start_reg[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .Q(
        start_reg[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .Q(
        start_reg[127]) );
  DFF \start_reg_reg[128]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .Q(
        start_reg[128]) );
  DFF \start_reg_reg[129]  ( .D(start_in[128]), .CLK(clk), .RST(rst), .Q(
        start_reg[129]) );
  DFF \start_reg_reg[130]  ( .D(start_in[129]), .CLK(clk), .RST(rst), .Q(
        start_reg[130]) );
  DFF \start_reg_reg[131]  ( .D(start_in[130]), .CLK(clk), .RST(rst), .Q(
        start_reg[131]) );
  DFF \start_reg_reg[132]  ( .D(start_in[131]), .CLK(clk), .RST(rst), .Q(
        start_reg[132]) );
  DFF \start_reg_reg[133]  ( .D(start_in[132]), .CLK(clk), .RST(rst), .Q(
        start_reg[133]) );
  DFF \start_reg_reg[134]  ( .D(start_in[133]), .CLK(clk), .RST(rst), .Q(
        start_reg[134]) );
  DFF \start_reg_reg[135]  ( .D(start_in[134]), .CLK(clk), .RST(rst), .Q(
        start_reg[135]) );
  DFF \start_reg_reg[136]  ( .D(start_in[135]), .CLK(clk), .RST(rst), .Q(
        start_reg[136]) );
  DFF \start_reg_reg[137]  ( .D(start_in[136]), .CLK(clk), .RST(rst), .Q(
        start_reg[137]) );
  DFF \start_reg_reg[138]  ( .D(start_in[137]), .CLK(clk), .RST(rst), .Q(
        start_reg[138]) );
  DFF \start_reg_reg[139]  ( .D(start_in[138]), .CLK(clk), .RST(rst), .Q(
        start_reg[139]) );
  DFF \start_reg_reg[140]  ( .D(start_in[139]), .CLK(clk), .RST(rst), .Q(
        start_reg[140]) );
  DFF \start_reg_reg[141]  ( .D(start_in[140]), .CLK(clk), .RST(rst), .Q(
        start_reg[141]) );
  DFF \start_reg_reg[142]  ( .D(start_in[141]), .CLK(clk), .RST(rst), .Q(
        start_reg[142]) );
  DFF \start_reg_reg[143]  ( .D(start_in[142]), .CLK(clk), .RST(rst), .Q(
        start_reg[143]) );
  DFF \start_reg_reg[144]  ( .D(start_in[143]), .CLK(clk), .RST(rst), .Q(
        start_reg[144]) );
  DFF \start_reg_reg[145]  ( .D(start_in[144]), .CLK(clk), .RST(rst), .Q(
        start_reg[145]) );
  DFF \start_reg_reg[146]  ( .D(start_in[145]), .CLK(clk), .RST(rst), .Q(
        start_reg[146]) );
  DFF \start_reg_reg[147]  ( .D(start_in[146]), .CLK(clk), .RST(rst), .Q(
        start_reg[147]) );
  DFF \start_reg_reg[148]  ( .D(start_in[147]), .CLK(clk), .RST(rst), .Q(
        start_reg[148]) );
  DFF \start_reg_reg[149]  ( .D(start_in[148]), .CLK(clk), .RST(rst), .Q(
        start_reg[149]) );
  DFF \start_reg_reg[150]  ( .D(start_in[149]), .CLK(clk), .RST(rst), .Q(
        start_reg[150]) );
  DFF \start_reg_reg[151]  ( .D(start_in[150]), .CLK(clk), .RST(rst), .Q(
        start_reg[151]) );
  DFF \start_reg_reg[152]  ( .D(start_in[151]), .CLK(clk), .RST(rst), .Q(
        start_reg[152]) );
  DFF \start_reg_reg[153]  ( .D(start_in[152]), .CLK(clk), .RST(rst), .Q(
        start_reg[153]) );
  DFF \start_reg_reg[154]  ( .D(start_in[153]), .CLK(clk), .RST(rst), .Q(
        start_reg[154]) );
  DFF \start_reg_reg[155]  ( .D(start_in[154]), .CLK(clk), .RST(rst), .Q(
        start_reg[155]) );
  DFF \start_reg_reg[156]  ( .D(start_in[155]), .CLK(clk), .RST(rst), .Q(
        start_reg[156]) );
  DFF \start_reg_reg[157]  ( .D(start_in[156]), .CLK(clk), .RST(rst), .Q(
        start_reg[157]) );
  DFF \start_reg_reg[158]  ( .D(start_in[157]), .CLK(clk), .RST(rst), .Q(
        start_reg[158]) );
  DFF \start_reg_reg[159]  ( .D(start_in[158]), .CLK(clk), .RST(rst), .Q(
        start_reg[159]) );
  DFF \start_reg_reg[160]  ( .D(start_in[159]), .CLK(clk), .RST(rst), .Q(
        start_reg[160]) );
  DFF \start_reg_reg[161]  ( .D(start_in[160]), .CLK(clk), .RST(rst), .Q(
        start_reg[161]) );
  DFF \start_reg_reg[162]  ( .D(start_in[161]), .CLK(clk), .RST(rst), .Q(
        start_reg[162]) );
  DFF \start_reg_reg[163]  ( .D(start_in[162]), .CLK(clk), .RST(rst), .Q(
        start_reg[163]) );
  DFF \start_reg_reg[164]  ( .D(start_in[163]), .CLK(clk), .RST(rst), .Q(
        start_reg[164]) );
  DFF \start_reg_reg[165]  ( .D(start_in[164]), .CLK(clk), .RST(rst), .Q(
        start_reg[165]) );
  DFF \start_reg_reg[166]  ( .D(start_in[165]), .CLK(clk), .RST(rst), .Q(
        start_reg[166]) );
  DFF \start_reg_reg[167]  ( .D(start_in[166]), .CLK(clk), .RST(rst), .Q(
        start_reg[167]) );
  DFF \start_reg_reg[168]  ( .D(start_in[167]), .CLK(clk), .RST(rst), .Q(
        start_reg[168]) );
  DFF \start_reg_reg[169]  ( .D(start_in[168]), .CLK(clk), .RST(rst), .Q(
        start_reg[169]) );
  DFF \start_reg_reg[170]  ( .D(start_in[169]), .CLK(clk), .RST(rst), .Q(
        start_reg[170]) );
  DFF \start_reg_reg[171]  ( .D(start_in[170]), .CLK(clk), .RST(rst), .Q(
        start_reg[171]) );
  DFF \start_reg_reg[172]  ( .D(start_in[171]), .CLK(clk), .RST(rst), .Q(
        start_reg[172]) );
  DFF \start_reg_reg[173]  ( .D(start_in[172]), .CLK(clk), .RST(rst), .Q(
        start_reg[173]) );
  DFF \start_reg_reg[174]  ( .D(start_in[173]), .CLK(clk), .RST(rst), .Q(
        start_reg[174]) );
  DFF \start_reg_reg[175]  ( .D(start_in[174]), .CLK(clk), .RST(rst), .Q(
        start_reg[175]) );
  DFF \start_reg_reg[176]  ( .D(start_in[175]), .CLK(clk), .RST(rst), .Q(
        start_reg[176]) );
  DFF \start_reg_reg[177]  ( .D(start_in[176]), .CLK(clk), .RST(rst), .Q(
        start_reg[177]) );
  DFF \start_reg_reg[178]  ( .D(start_in[177]), .CLK(clk), .RST(rst), .Q(
        start_reg[178]) );
  DFF \start_reg_reg[179]  ( .D(start_in[178]), .CLK(clk), .RST(rst), .Q(
        start_reg[179]) );
  DFF \start_reg_reg[180]  ( .D(start_in[179]), .CLK(clk), .RST(rst), .Q(
        start_reg[180]) );
  DFF \start_reg_reg[181]  ( .D(start_in[180]), .CLK(clk), .RST(rst), .Q(
        start_reg[181]) );
  DFF \start_reg_reg[182]  ( .D(start_in[181]), .CLK(clk), .RST(rst), .Q(
        start_reg[182]) );
  DFF \start_reg_reg[183]  ( .D(start_in[182]), .CLK(clk), .RST(rst), .Q(
        start_reg[183]) );
  DFF \start_reg_reg[184]  ( .D(start_in[183]), .CLK(clk), .RST(rst), .Q(
        start_reg[184]) );
  DFF \start_reg_reg[185]  ( .D(start_in[184]), .CLK(clk), .RST(rst), .Q(
        start_reg[185]) );
  DFF \start_reg_reg[186]  ( .D(start_in[185]), .CLK(clk), .RST(rst), .Q(
        start_reg[186]) );
  DFF \start_reg_reg[187]  ( .D(start_in[186]), .CLK(clk), .RST(rst), .Q(
        start_reg[187]) );
  DFF \start_reg_reg[188]  ( .D(start_in[187]), .CLK(clk), .RST(rst), .Q(
        start_reg[188]) );
  DFF \start_reg_reg[189]  ( .D(start_in[188]), .CLK(clk), .RST(rst), .Q(
        start_reg[189]) );
  DFF \start_reg_reg[190]  ( .D(start_in[189]), .CLK(clk), .RST(rst), .Q(
        start_reg[190]) );
  DFF \start_reg_reg[191]  ( .D(start_in[190]), .CLK(clk), .RST(rst), .Q(
        start_reg[191]) );
  DFF \start_reg_reg[192]  ( .D(start_in[191]), .CLK(clk), .RST(rst), .Q(
        start_reg[192]) );
  DFF \start_reg_reg[193]  ( .D(start_in[192]), .CLK(clk), .RST(rst), .Q(
        start_reg[193]) );
  DFF \start_reg_reg[194]  ( .D(start_in[193]), .CLK(clk), .RST(rst), .Q(
        start_reg[194]) );
  DFF \start_reg_reg[195]  ( .D(start_in[194]), .CLK(clk), .RST(rst), .Q(
        start_reg[195]) );
  DFF \start_reg_reg[196]  ( .D(start_in[195]), .CLK(clk), .RST(rst), .Q(
        start_reg[196]) );
  DFF \start_reg_reg[197]  ( .D(start_in[196]), .CLK(clk), .RST(rst), .Q(
        start_reg[197]) );
  DFF \start_reg_reg[198]  ( .D(start_in[197]), .CLK(clk), .RST(rst), .Q(
        start_reg[198]) );
  DFF \start_reg_reg[199]  ( .D(start_in[198]), .CLK(clk), .RST(rst), .Q(
        start_reg[199]) );
  DFF \start_reg_reg[200]  ( .D(start_in[199]), .CLK(clk), .RST(rst), .Q(
        start_reg[200]) );
  DFF \start_reg_reg[201]  ( .D(start_in[200]), .CLK(clk), .RST(rst), .Q(
        start_reg[201]) );
  DFF \start_reg_reg[202]  ( .D(start_in[201]), .CLK(clk), .RST(rst), .Q(
        start_reg[202]) );
  DFF \start_reg_reg[203]  ( .D(start_in[202]), .CLK(clk), .RST(rst), .Q(
        start_reg[203]) );
  DFF \start_reg_reg[204]  ( .D(start_in[203]), .CLK(clk), .RST(rst), .Q(
        start_reg[204]) );
  DFF \start_reg_reg[205]  ( .D(start_in[204]), .CLK(clk), .RST(rst), .Q(
        start_reg[205]) );
  DFF \start_reg_reg[206]  ( .D(start_in[205]), .CLK(clk), .RST(rst), .Q(
        start_reg[206]) );
  DFF \start_reg_reg[207]  ( .D(start_in[206]), .CLK(clk), .RST(rst), .Q(
        start_reg[207]) );
  DFF \start_reg_reg[208]  ( .D(start_in[207]), .CLK(clk), .RST(rst), .Q(
        start_reg[208]) );
  DFF \start_reg_reg[209]  ( .D(start_in[208]), .CLK(clk), .RST(rst), .Q(
        start_reg[209]) );
  DFF \start_reg_reg[210]  ( .D(start_in[209]), .CLK(clk), .RST(rst), .Q(
        start_reg[210]) );
  DFF \start_reg_reg[211]  ( .D(start_in[210]), .CLK(clk), .RST(rst), .Q(
        start_reg[211]) );
  DFF \start_reg_reg[212]  ( .D(start_in[211]), .CLK(clk), .RST(rst), .Q(
        start_reg[212]) );
  DFF \start_reg_reg[213]  ( .D(start_in[212]), .CLK(clk), .RST(rst), .Q(
        start_reg[213]) );
  DFF \start_reg_reg[214]  ( .D(start_in[213]), .CLK(clk), .RST(rst), .Q(
        start_reg[214]) );
  DFF \start_reg_reg[215]  ( .D(start_in[214]), .CLK(clk), .RST(rst), .Q(
        start_reg[215]) );
  DFF \start_reg_reg[216]  ( .D(start_in[215]), .CLK(clk), .RST(rst), .Q(
        start_reg[216]) );
  DFF \start_reg_reg[217]  ( .D(start_in[216]), .CLK(clk), .RST(rst), .Q(
        start_reg[217]) );
  DFF \start_reg_reg[218]  ( .D(start_in[217]), .CLK(clk), .RST(rst), .Q(
        start_reg[218]) );
  DFF \start_reg_reg[219]  ( .D(start_in[218]), .CLK(clk), .RST(rst), .Q(
        start_reg[219]) );
  DFF \start_reg_reg[220]  ( .D(start_in[219]), .CLK(clk), .RST(rst), .Q(
        start_reg[220]) );
  DFF \start_reg_reg[221]  ( .D(start_in[220]), .CLK(clk), .RST(rst), .Q(
        start_reg[221]) );
  DFF \start_reg_reg[222]  ( .D(start_in[221]), .CLK(clk), .RST(rst), .Q(
        start_reg[222]) );
  DFF \start_reg_reg[223]  ( .D(start_in[222]), .CLK(clk), .RST(rst), .Q(
        start_reg[223]) );
  DFF \start_reg_reg[224]  ( .D(start_in[223]), .CLK(clk), .RST(rst), .Q(
        start_reg[224]) );
  DFF \start_reg_reg[225]  ( .D(start_in[224]), .CLK(clk), .RST(rst), .Q(
        start_reg[225]) );
  DFF \start_reg_reg[226]  ( .D(start_in[225]), .CLK(clk), .RST(rst), .Q(
        start_reg[226]) );
  DFF \start_reg_reg[227]  ( .D(start_in[226]), .CLK(clk), .RST(rst), .Q(
        start_reg[227]) );
  DFF \start_reg_reg[228]  ( .D(start_in[227]), .CLK(clk), .RST(rst), .Q(
        start_reg[228]) );
  DFF \start_reg_reg[229]  ( .D(start_in[228]), .CLK(clk), .RST(rst), .Q(
        start_reg[229]) );
  DFF \start_reg_reg[230]  ( .D(start_in[229]), .CLK(clk), .RST(rst), .Q(
        start_reg[230]) );
  DFF \start_reg_reg[231]  ( .D(start_in[230]), .CLK(clk), .RST(rst), .Q(
        start_reg[231]) );
  DFF \start_reg_reg[232]  ( .D(start_in[231]), .CLK(clk), .RST(rst), .Q(
        start_reg[232]) );
  DFF \start_reg_reg[233]  ( .D(start_in[232]), .CLK(clk), .RST(rst), .Q(
        start_reg[233]) );
  DFF \start_reg_reg[234]  ( .D(start_in[233]), .CLK(clk), .RST(rst), .Q(
        start_reg[234]) );
  DFF \start_reg_reg[235]  ( .D(start_in[234]), .CLK(clk), .RST(rst), .Q(
        start_reg[235]) );
  DFF \start_reg_reg[236]  ( .D(start_in[235]), .CLK(clk), .RST(rst), .Q(
        start_reg[236]) );
  DFF \start_reg_reg[237]  ( .D(start_in[236]), .CLK(clk), .RST(rst), .Q(
        start_reg[237]) );
  DFF \start_reg_reg[238]  ( .D(start_in[237]), .CLK(clk), .RST(rst), .Q(
        start_reg[238]) );
  DFF \start_reg_reg[239]  ( .D(start_in[238]), .CLK(clk), .RST(rst), .Q(
        start_reg[239]) );
  DFF \start_reg_reg[240]  ( .D(start_in[239]), .CLK(clk), .RST(rst), .Q(
        start_reg[240]) );
  DFF \start_reg_reg[241]  ( .D(start_in[240]), .CLK(clk), .RST(rst), .Q(
        start_reg[241]) );
  DFF \start_reg_reg[242]  ( .D(start_in[241]), .CLK(clk), .RST(rst), .Q(
        start_reg[242]) );
  DFF \start_reg_reg[243]  ( .D(start_in[242]), .CLK(clk), .RST(rst), .Q(
        start_reg[243]) );
  DFF \start_reg_reg[244]  ( .D(start_in[243]), .CLK(clk), .RST(rst), .Q(
        start_reg[244]) );
  DFF \start_reg_reg[245]  ( .D(start_in[244]), .CLK(clk), .RST(rst), .Q(
        start_reg[245]) );
  DFF \start_reg_reg[246]  ( .D(start_in[245]), .CLK(clk), .RST(rst), .Q(
        start_reg[246]) );
  DFF \start_reg_reg[247]  ( .D(start_in[246]), .CLK(clk), .RST(rst), .Q(
        start_reg[247]) );
  DFF \start_reg_reg[248]  ( .D(start_in[247]), .CLK(clk), .RST(rst), .Q(
        start_reg[248]) );
  DFF \start_reg_reg[249]  ( .D(start_in[248]), .CLK(clk), .RST(rst), .Q(
        start_reg[249]) );
  DFF \start_reg_reg[250]  ( .D(start_in[249]), .CLK(clk), .RST(rst), .Q(
        start_reg[250]) );
  DFF \start_reg_reg[251]  ( .D(start_in[250]), .CLK(clk), .RST(rst), .Q(
        start_reg[251]) );
  DFF \start_reg_reg[252]  ( .D(start_in[251]), .CLK(clk), .RST(rst), .Q(
        start_reg[252]) );
  DFF \start_reg_reg[253]  ( .D(start_in[252]), .CLK(clk), .RST(rst), .Q(
        start_reg[253]) );
  DFF \start_reg_reg[254]  ( .D(start_in[253]), .CLK(clk), .RST(rst), .Q(
        start_reg[254]) );
  DFF \start_reg_reg[255]  ( .D(start_in[254]), .CLK(clk), .RST(rst), .Q(
        start_reg[255]) );
  DFF \start_reg_reg[256]  ( .D(start_in[255]), .CLK(clk), .RST(rst), .Q(
        start_reg[256]) );
  DFF \start_reg_reg[257]  ( .D(start_in[256]), .CLK(clk), .RST(rst), .Q(
        start_reg[257]) );
  DFF \start_reg_reg[258]  ( .D(start_in[257]), .CLK(clk), .RST(rst), .Q(
        start_reg[258]) );
  DFF \start_reg_reg[259]  ( .D(start_in[258]), .CLK(clk), .RST(rst), .Q(
        start_reg[259]) );
  DFF \start_reg_reg[260]  ( .D(start_in[259]), .CLK(clk), .RST(rst), .Q(
        start_reg[260]) );
  DFF \start_reg_reg[261]  ( .D(start_in[260]), .CLK(clk), .RST(rst), .Q(
        start_reg[261]) );
  DFF \start_reg_reg[262]  ( .D(start_in[261]), .CLK(clk), .RST(rst), .Q(
        start_reg[262]) );
  DFF \start_reg_reg[263]  ( .D(start_in[262]), .CLK(clk), .RST(rst), .Q(
        start_reg[263]) );
  DFF \start_reg_reg[264]  ( .D(start_in[263]), .CLK(clk), .RST(rst), .Q(
        start_reg[264]) );
  DFF \start_reg_reg[265]  ( .D(start_in[264]), .CLK(clk), .RST(rst), .Q(
        start_reg[265]) );
  DFF \start_reg_reg[266]  ( .D(start_in[265]), .CLK(clk), .RST(rst), .Q(
        start_reg[266]) );
  DFF \start_reg_reg[267]  ( .D(start_in[266]), .CLK(clk), .RST(rst), .Q(
        start_reg[267]) );
  DFF \start_reg_reg[268]  ( .D(start_in[267]), .CLK(clk), .RST(rst), .Q(
        start_reg[268]) );
  DFF \start_reg_reg[269]  ( .D(start_in[268]), .CLK(clk), .RST(rst), .Q(
        start_reg[269]) );
  DFF \start_reg_reg[270]  ( .D(start_in[269]), .CLK(clk), .RST(rst), .Q(
        start_reg[270]) );
  DFF \start_reg_reg[271]  ( .D(start_in[270]), .CLK(clk), .RST(rst), .Q(
        start_reg[271]) );
  DFF \start_reg_reg[272]  ( .D(start_in[271]), .CLK(clk), .RST(rst), .Q(
        start_reg[272]) );
  DFF \start_reg_reg[273]  ( .D(start_in[272]), .CLK(clk), .RST(rst), .Q(
        start_reg[273]) );
  DFF \start_reg_reg[274]  ( .D(start_in[273]), .CLK(clk), .RST(rst), .Q(
        start_reg[274]) );
  DFF \start_reg_reg[275]  ( .D(start_in[274]), .CLK(clk), .RST(rst), .Q(
        start_reg[275]) );
  DFF \start_reg_reg[276]  ( .D(start_in[275]), .CLK(clk), .RST(rst), .Q(
        start_reg[276]) );
  DFF \start_reg_reg[277]  ( .D(start_in[276]), .CLK(clk), .RST(rst), .Q(
        start_reg[277]) );
  DFF \start_reg_reg[278]  ( .D(start_in[277]), .CLK(clk), .RST(rst), .Q(
        start_reg[278]) );
  DFF \start_reg_reg[279]  ( .D(start_in[278]), .CLK(clk), .RST(rst), .Q(
        start_reg[279]) );
  DFF \start_reg_reg[280]  ( .D(start_in[279]), .CLK(clk), .RST(rst), .Q(
        start_reg[280]) );
  DFF \start_reg_reg[281]  ( .D(start_in[280]), .CLK(clk), .RST(rst), .Q(
        start_reg[281]) );
  DFF \start_reg_reg[282]  ( .D(start_in[281]), .CLK(clk), .RST(rst), .Q(
        start_reg[282]) );
  DFF \start_reg_reg[283]  ( .D(start_in[282]), .CLK(clk), .RST(rst), .Q(
        start_reg[283]) );
  DFF \start_reg_reg[284]  ( .D(start_in[283]), .CLK(clk), .RST(rst), .Q(
        start_reg[284]) );
  DFF \start_reg_reg[285]  ( .D(start_in[284]), .CLK(clk), .RST(rst), .Q(
        start_reg[285]) );
  DFF \start_reg_reg[286]  ( .D(start_in[285]), .CLK(clk), .RST(rst), .Q(
        start_reg[286]) );
  DFF \start_reg_reg[287]  ( .D(start_in[286]), .CLK(clk), .RST(rst), .Q(
        start_reg[287]) );
  DFF \start_reg_reg[288]  ( .D(start_in[287]), .CLK(clk), .RST(rst), .Q(
        start_reg[288]) );
  DFF \start_reg_reg[289]  ( .D(start_in[288]), .CLK(clk), .RST(rst), .Q(
        start_reg[289]) );
  DFF \start_reg_reg[290]  ( .D(start_in[289]), .CLK(clk), .RST(rst), .Q(
        start_reg[290]) );
  DFF \start_reg_reg[291]  ( .D(start_in[290]), .CLK(clk), .RST(rst), .Q(
        start_reg[291]) );
  DFF \start_reg_reg[292]  ( .D(start_in[291]), .CLK(clk), .RST(rst), .Q(
        start_reg[292]) );
  DFF \start_reg_reg[293]  ( .D(start_in[292]), .CLK(clk), .RST(rst), .Q(
        start_reg[293]) );
  DFF \start_reg_reg[294]  ( .D(start_in[293]), .CLK(clk), .RST(rst), .Q(
        start_reg[294]) );
  DFF \start_reg_reg[295]  ( .D(start_in[294]), .CLK(clk), .RST(rst), .Q(
        start_reg[295]) );
  DFF \start_reg_reg[296]  ( .D(start_in[295]), .CLK(clk), .RST(rst), .Q(
        start_reg[296]) );
  DFF \start_reg_reg[297]  ( .D(start_in[296]), .CLK(clk), .RST(rst), .Q(
        start_reg[297]) );
  DFF \start_reg_reg[298]  ( .D(start_in[297]), .CLK(clk), .RST(rst), .Q(
        start_reg[298]) );
  DFF \start_reg_reg[299]  ( .D(start_in[298]), .CLK(clk), .RST(rst), .Q(
        start_reg[299]) );
  DFF \start_reg_reg[300]  ( .D(start_in[299]), .CLK(clk), .RST(rst), .Q(
        start_reg[300]) );
  DFF \start_reg_reg[301]  ( .D(start_in[300]), .CLK(clk), .RST(rst), .Q(
        start_reg[301]) );
  DFF \start_reg_reg[302]  ( .D(start_in[301]), .CLK(clk), .RST(rst), .Q(
        start_reg[302]) );
  DFF \start_reg_reg[303]  ( .D(start_in[302]), .CLK(clk), .RST(rst), .Q(
        start_reg[303]) );
  DFF \start_reg_reg[304]  ( .D(start_in[303]), .CLK(clk), .RST(rst), .Q(
        start_reg[304]) );
  DFF \start_reg_reg[305]  ( .D(start_in[304]), .CLK(clk), .RST(rst), .Q(
        start_reg[305]) );
  DFF \start_reg_reg[306]  ( .D(start_in[305]), .CLK(clk), .RST(rst), .Q(
        start_reg[306]) );
  DFF \start_reg_reg[307]  ( .D(start_in[306]), .CLK(clk), .RST(rst), .Q(
        start_reg[307]) );
  DFF \start_reg_reg[308]  ( .D(start_in[307]), .CLK(clk), .RST(rst), .Q(
        start_reg[308]) );
  DFF \start_reg_reg[309]  ( .D(start_in[308]), .CLK(clk), .RST(rst), .Q(
        start_reg[309]) );
  DFF \start_reg_reg[310]  ( .D(start_in[309]), .CLK(clk), .RST(rst), .Q(
        start_reg[310]) );
  DFF \start_reg_reg[311]  ( .D(start_in[310]), .CLK(clk), .RST(rst), .Q(
        start_reg[311]) );
  DFF \start_reg_reg[312]  ( .D(start_in[311]), .CLK(clk), .RST(rst), .Q(
        start_reg[312]) );
  DFF \start_reg_reg[313]  ( .D(start_in[312]), .CLK(clk), .RST(rst), .Q(
        start_reg[313]) );
  DFF \start_reg_reg[314]  ( .D(start_in[313]), .CLK(clk), .RST(rst), .Q(
        start_reg[314]) );
  DFF \start_reg_reg[315]  ( .D(start_in[314]), .CLK(clk), .RST(rst), .Q(
        start_reg[315]) );
  DFF \start_reg_reg[316]  ( .D(start_in[315]), .CLK(clk), .RST(rst), .Q(
        start_reg[316]) );
  DFF \start_reg_reg[317]  ( .D(start_in[316]), .CLK(clk), .RST(rst), .Q(
        start_reg[317]) );
  DFF \start_reg_reg[318]  ( .D(start_in[317]), .CLK(clk), .RST(rst), .Q(
        start_reg[318]) );
  DFF \start_reg_reg[319]  ( .D(start_in[318]), .CLK(clk), .RST(rst), .Q(
        start_reg[319]) );
  DFF \start_reg_reg[320]  ( .D(start_in[319]), .CLK(clk), .RST(rst), .Q(
        start_reg[320]) );
  DFF \start_reg_reg[321]  ( .D(start_in[320]), .CLK(clk), .RST(rst), .Q(
        start_reg[321]) );
  DFF \start_reg_reg[322]  ( .D(start_in[321]), .CLK(clk), .RST(rst), .Q(
        start_reg[322]) );
  DFF \start_reg_reg[323]  ( .D(start_in[322]), .CLK(clk), .RST(rst), .Q(
        start_reg[323]) );
  DFF \start_reg_reg[324]  ( .D(start_in[323]), .CLK(clk), .RST(rst), .Q(
        start_reg[324]) );
  DFF \start_reg_reg[325]  ( .D(start_in[324]), .CLK(clk), .RST(rst), .Q(
        start_reg[325]) );
  DFF \start_reg_reg[326]  ( .D(start_in[325]), .CLK(clk), .RST(rst), .Q(
        start_reg[326]) );
  DFF \start_reg_reg[327]  ( .D(start_in[326]), .CLK(clk), .RST(rst), .Q(
        start_reg[327]) );
  DFF \start_reg_reg[328]  ( .D(start_in[327]), .CLK(clk), .RST(rst), .Q(
        start_reg[328]) );
  DFF \start_reg_reg[329]  ( .D(start_in[328]), .CLK(clk), .RST(rst), .Q(
        start_reg[329]) );
  DFF \start_reg_reg[330]  ( .D(start_in[329]), .CLK(clk), .RST(rst), .Q(
        start_reg[330]) );
  DFF \start_reg_reg[331]  ( .D(start_in[330]), .CLK(clk), .RST(rst), .Q(
        start_reg[331]) );
  DFF \start_reg_reg[332]  ( .D(start_in[331]), .CLK(clk), .RST(rst), .Q(
        start_reg[332]) );
  DFF \start_reg_reg[333]  ( .D(start_in[332]), .CLK(clk), .RST(rst), .Q(
        start_reg[333]) );
  DFF \start_reg_reg[334]  ( .D(start_in[333]), .CLK(clk), .RST(rst), .Q(
        start_reg[334]) );
  DFF \start_reg_reg[335]  ( .D(start_in[334]), .CLK(clk), .RST(rst), .Q(
        start_reg[335]) );
  DFF \start_reg_reg[336]  ( .D(start_in[335]), .CLK(clk), .RST(rst), .Q(
        start_reg[336]) );
  DFF \start_reg_reg[337]  ( .D(start_in[336]), .CLK(clk), .RST(rst), .Q(
        start_reg[337]) );
  DFF \start_reg_reg[338]  ( .D(start_in[337]), .CLK(clk), .RST(rst), .Q(
        start_reg[338]) );
  DFF \start_reg_reg[339]  ( .D(start_in[338]), .CLK(clk), .RST(rst), .Q(
        start_reg[339]) );
  DFF \start_reg_reg[340]  ( .D(start_in[339]), .CLK(clk), .RST(rst), .Q(
        start_reg[340]) );
  DFF \start_reg_reg[341]  ( .D(start_in[340]), .CLK(clk), .RST(rst), .Q(
        start_reg[341]) );
  DFF \start_reg_reg[342]  ( .D(start_in[341]), .CLK(clk), .RST(rst), .Q(
        start_reg[342]) );
  DFF \start_reg_reg[343]  ( .D(start_in[342]), .CLK(clk), .RST(rst), .Q(
        start_reg[343]) );
  DFF \start_reg_reg[344]  ( .D(start_in[343]), .CLK(clk), .RST(rst), .Q(
        start_reg[344]) );
  DFF \start_reg_reg[345]  ( .D(start_in[344]), .CLK(clk), .RST(rst), .Q(
        start_reg[345]) );
  DFF \start_reg_reg[346]  ( .D(start_in[345]), .CLK(clk), .RST(rst), .Q(
        start_reg[346]) );
  DFF \start_reg_reg[347]  ( .D(start_in[346]), .CLK(clk), .RST(rst), .Q(
        start_reg[347]) );
  DFF \start_reg_reg[348]  ( .D(start_in[347]), .CLK(clk), .RST(rst), .Q(
        start_reg[348]) );
  DFF \start_reg_reg[349]  ( .D(start_in[348]), .CLK(clk), .RST(rst), .Q(
        start_reg[349]) );
  DFF \start_reg_reg[350]  ( .D(start_in[349]), .CLK(clk), .RST(rst), .Q(
        start_reg[350]) );
  DFF \start_reg_reg[351]  ( .D(start_in[350]), .CLK(clk), .RST(rst), .Q(
        start_reg[351]) );
  DFF \start_reg_reg[352]  ( .D(start_in[351]), .CLK(clk), .RST(rst), .Q(
        start_reg[352]) );
  DFF \start_reg_reg[353]  ( .D(start_in[352]), .CLK(clk), .RST(rst), .Q(
        start_reg[353]) );
  DFF \start_reg_reg[354]  ( .D(start_in[353]), .CLK(clk), .RST(rst), .Q(
        start_reg[354]) );
  DFF \start_reg_reg[355]  ( .D(start_in[354]), .CLK(clk), .RST(rst), .Q(
        start_reg[355]) );
  DFF \start_reg_reg[356]  ( .D(start_in[355]), .CLK(clk), .RST(rst), .Q(
        start_reg[356]) );
  DFF \start_reg_reg[357]  ( .D(start_in[356]), .CLK(clk), .RST(rst), .Q(
        start_reg[357]) );
  DFF \start_reg_reg[358]  ( .D(start_in[357]), .CLK(clk), .RST(rst), .Q(
        start_reg[358]) );
  DFF \start_reg_reg[359]  ( .D(start_in[358]), .CLK(clk), .RST(rst), .Q(
        start_reg[359]) );
  DFF \start_reg_reg[360]  ( .D(start_in[359]), .CLK(clk), .RST(rst), .Q(
        start_reg[360]) );
  DFF \start_reg_reg[361]  ( .D(start_in[360]), .CLK(clk), .RST(rst), .Q(
        start_reg[361]) );
  DFF \start_reg_reg[362]  ( .D(start_in[361]), .CLK(clk), .RST(rst), .Q(
        start_reg[362]) );
  DFF \start_reg_reg[363]  ( .D(start_in[362]), .CLK(clk), .RST(rst), .Q(
        start_reg[363]) );
  DFF \start_reg_reg[364]  ( .D(start_in[363]), .CLK(clk), .RST(rst), .Q(
        start_reg[364]) );
  DFF \start_reg_reg[365]  ( .D(start_in[364]), .CLK(clk), .RST(rst), .Q(
        start_reg[365]) );
  DFF \start_reg_reg[366]  ( .D(start_in[365]), .CLK(clk), .RST(rst), .Q(
        start_reg[366]) );
  DFF \start_reg_reg[367]  ( .D(start_in[366]), .CLK(clk), .RST(rst), .Q(
        start_reg[367]) );
  DFF \start_reg_reg[368]  ( .D(start_in[367]), .CLK(clk), .RST(rst), .Q(
        start_reg[368]) );
  DFF \start_reg_reg[369]  ( .D(start_in[368]), .CLK(clk), .RST(rst), .Q(
        start_reg[369]) );
  DFF \start_reg_reg[370]  ( .D(start_in[369]), .CLK(clk), .RST(rst), .Q(
        start_reg[370]) );
  DFF \start_reg_reg[371]  ( .D(start_in[370]), .CLK(clk), .RST(rst), .Q(
        start_reg[371]) );
  DFF \start_reg_reg[372]  ( .D(start_in[371]), .CLK(clk), .RST(rst), .Q(
        start_reg[372]) );
  DFF \start_reg_reg[373]  ( .D(start_in[372]), .CLK(clk), .RST(rst), .Q(
        start_reg[373]) );
  DFF \start_reg_reg[374]  ( .D(start_in[373]), .CLK(clk), .RST(rst), .Q(
        start_reg[374]) );
  DFF \start_reg_reg[375]  ( .D(start_in[374]), .CLK(clk), .RST(rst), .Q(
        start_reg[375]) );
  DFF \start_reg_reg[376]  ( .D(start_in[375]), .CLK(clk), .RST(rst), .Q(
        start_reg[376]) );
  DFF \start_reg_reg[377]  ( .D(start_in[376]), .CLK(clk), .RST(rst), .Q(
        start_reg[377]) );
  DFF \start_reg_reg[378]  ( .D(start_in[377]), .CLK(clk), .RST(rst), .Q(
        start_reg[378]) );
  DFF \start_reg_reg[379]  ( .D(start_in[378]), .CLK(clk), .RST(rst), .Q(
        start_reg[379]) );
  DFF \start_reg_reg[380]  ( .D(start_in[379]), .CLK(clk), .RST(rst), .Q(
        start_reg[380]) );
  DFF \start_reg_reg[381]  ( .D(start_in[380]), .CLK(clk), .RST(rst), .Q(
        start_reg[381]) );
  DFF \start_reg_reg[382]  ( .D(start_in[381]), .CLK(clk), .RST(rst), .Q(
        start_reg[382]) );
  DFF \start_reg_reg[383]  ( .D(start_in[382]), .CLK(clk), .RST(rst), .Q(
        start_reg[383]) );
  DFF \start_reg_reg[384]  ( .D(start_in[383]), .CLK(clk), .RST(rst), .Q(
        start_reg[384]) );
  DFF \start_reg_reg[385]  ( .D(start_in[384]), .CLK(clk), .RST(rst), .Q(
        start_reg[385]) );
  DFF \start_reg_reg[386]  ( .D(start_in[385]), .CLK(clk), .RST(rst), .Q(
        start_reg[386]) );
  DFF \start_reg_reg[387]  ( .D(start_in[386]), .CLK(clk), .RST(rst), .Q(
        start_reg[387]) );
  DFF \start_reg_reg[388]  ( .D(start_in[387]), .CLK(clk), .RST(rst), .Q(
        start_reg[388]) );
  DFF \start_reg_reg[389]  ( .D(start_in[388]), .CLK(clk), .RST(rst), .Q(
        start_reg[389]) );
  DFF \start_reg_reg[390]  ( .D(start_in[389]), .CLK(clk), .RST(rst), .Q(
        start_reg[390]) );
  DFF \start_reg_reg[391]  ( .D(start_in[390]), .CLK(clk), .RST(rst), .Q(
        start_reg[391]) );
  DFF \start_reg_reg[392]  ( .D(start_in[391]), .CLK(clk), .RST(rst), .Q(
        start_reg[392]) );
  DFF \start_reg_reg[393]  ( .D(start_in[392]), .CLK(clk), .RST(rst), .Q(
        start_reg[393]) );
  DFF \start_reg_reg[394]  ( .D(start_in[393]), .CLK(clk), .RST(rst), .Q(
        start_reg[394]) );
  DFF \start_reg_reg[395]  ( .D(start_in[394]), .CLK(clk), .RST(rst), .Q(
        start_reg[395]) );
  DFF \start_reg_reg[396]  ( .D(start_in[395]), .CLK(clk), .RST(rst), .Q(
        start_reg[396]) );
  DFF \start_reg_reg[397]  ( .D(start_in[396]), .CLK(clk), .RST(rst), .Q(
        start_reg[397]) );
  DFF \start_reg_reg[398]  ( .D(start_in[397]), .CLK(clk), .RST(rst), .Q(
        start_reg[398]) );
  DFF \start_reg_reg[399]  ( .D(start_in[398]), .CLK(clk), .RST(rst), .Q(
        start_reg[399]) );
  DFF \start_reg_reg[400]  ( .D(start_in[399]), .CLK(clk), .RST(rst), .Q(
        start_reg[400]) );
  DFF \start_reg_reg[401]  ( .D(start_in[400]), .CLK(clk), .RST(rst), .Q(
        start_reg[401]) );
  DFF \start_reg_reg[402]  ( .D(start_in[401]), .CLK(clk), .RST(rst), .Q(
        start_reg[402]) );
  DFF \start_reg_reg[403]  ( .D(start_in[402]), .CLK(clk), .RST(rst), .Q(
        start_reg[403]) );
  DFF \start_reg_reg[404]  ( .D(start_in[403]), .CLK(clk), .RST(rst), .Q(
        start_reg[404]) );
  DFF \start_reg_reg[405]  ( .D(start_in[404]), .CLK(clk), .RST(rst), .Q(
        start_reg[405]) );
  DFF \start_reg_reg[406]  ( .D(start_in[405]), .CLK(clk), .RST(rst), .Q(
        start_reg[406]) );
  DFF \start_reg_reg[407]  ( .D(start_in[406]), .CLK(clk), .RST(rst), .Q(
        start_reg[407]) );
  DFF \start_reg_reg[408]  ( .D(start_in[407]), .CLK(clk), .RST(rst), .Q(
        start_reg[408]) );
  DFF \start_reg_reg[409]  ( .D(start_in[408]), .CLK(clk), .RST(rst), .Q(
        start_reg[409]) );
  DFF \start_reg_reg[410]  ( .D(start_in[409]), .CLK(clk), .RST(rst), .Q(
        start_reg[410]) );
  DFF \start_reg_reg[411]  ( .D(start_in[410]), .CLK(clk), .RST(rst), .Q(
        start_reg[411]) );
  DFF \start_reg_reg[412]  ( .D(start_in[411]), .CLK(clk), .RST(rst), .Q(
        start_reg[412]) );
  DFF \start_reg_reg[413]  ( .D(start_in[412]), .CLK(clk), .RST(rst), .Q(
        start_reg[413]) );
  DFF \start_reg_reg[414]  ( .D(start_in[413]), .CLK(clk), .RST(rst), .Q(
        start_reg[414]) );
  DFF \start_reg_reg[415]  ( .D(start_in[414]), .CLK(clk), .RST(rst), .Q(
        start_reg[415]) );
  DFF \start_reg_reg[416]  ( .D(start_in[415]), .CLK(clk), .RST(rst), .Q(
        start_reg[416]) );
  DFF \start_reg_reg[417]  ( .D(start_in[416]), .CLK(clk), .RST(rst), .Q(
        start_reg[417]) );
  DFF \start_reg_reg[418]  ( .D(start_in[417]), .CLK(clk), .RST(rst), .Q(
        start_reg[418]) );
  DFF \start_reg_reg[419]  ( .D(start_in[418]), .CLK(clk), .RST(rst), .Q(
        start_reg[419]) );
  DFF \start_reg_reg[420]  ( .D(start_in[419]), .CLK(clk), .RST(rst), .Q(
        start_reg[420]) );
  DFF \start_reg_reg[421]  ( .D(start_in[420]), .CLK(clk), .RST(rst), .Q(
        start_reg[421]) );
  DFF \start_reg_reg[422]  ( .D(start_in[421]), .CLK(clk), .RST(rst), .Q(
        start_reg[422]) );
  DFF \start_reg_reg[423]  ( .D(start_in[422]), .CLK(clk), .RST(rst), .Q(
        start_reg[423]) );
  DFF \start_reg_reg[424]  ( .D(start_in[423]), .CLK(clk), .RST(rst), .Q(
        start_reg[424]) );
  DFF \start_reg_reg[425]  ( .D(start_in[424]), .CLK(clk), .RST(rst), .Q(
        start_reg[425]) );
  DFF \start_reg_reg[426]  ( .D(start_in[425]), .CLK(clk), .RST(rst), .Q(
        start_reg[426]) );
  DFF \start_reg_reg[427]  ( .D(start_in[426]), .CLK(clk), .RST(rst), .Q(
        start_reg[427]) );
  DFF \start_reg_reg[428]  ( .D(start_in[427]), .CLK(clk), .RST(rst), .Q(
        start_reg[428]) );
  DFF \start_reg_reg[429]  ( .D(start_in[428]), .CLK(clk), .RST(rst), .Q(
        start_reg[429]) );
  DFF \start_reg_reg[430]  ( .D(start_in[429]), .CLK(clk), .RST(rst), .Q(
        start_reg[430]) );
  DFF \start_reg_reg[431]  ( .D(start_in[430]), .CLK(clk), .RST(rst), .Q(
        start_reg[431]) );
  DFF \start_reg_reg[432]  ( .D(start_in[431]), .CLK(clk), .RST(rst), .Q(
        start_reg[432]) );
  DFF \start_reg_reg[433]  ( .D(start_in[432]), .CLK(clk), .RST(rst), .Q(
        start_reg[433]) );
  DFF \start_reg_reg[434]  ( .D(start_in[433]), .CLK(clk), .RST(rst), .Q(
        start_reg[434]) );
  DFF \start_reg_reg[435]  ( .D(start_in[434]), .CLK(clk), .RST(rst), .Q(
        start_reg[435]) );
  DFF \start_reg_reg[436]  ( .D(start_in[435]), .CLK(clk), .RST(rst), .Q(
        start_reg[436]) );
  DFF \start_reg_reg[437]  ( .D(start_in[436]), .CLK(clk), .RST(rst), .Q(
        start_reg[437]) );
  DFF \start_reg_reg[438]  ( .D(start_in[437]), .CLK(clk), .RST(rst), .Q(
        start_reg[438]) );
  DFF \start_reg_reg[439]  ( .D(start_in[438]), .CLK(clk), .RST(rst), .Q(
        start_reg[439]) );
  DFF \start_reg_reg[440]  ( .D(start_in[439]), .CLK(clk), .RST(rst), .Q(
        start_reg[440]) );
  DFF \start_reg_reg[441]  ( .D(start_in[440]), .CLK(clk), .RST(rst), .Q(
        start_reg[441]) );
  DFF \start_reg_reg[442]  ( .D(start_in[441]), .CLK(clk), .RST(rst), .Q(
        start_reg[442]) );
  DFF \start_reg_reg[443]  ( .D(start_in[442]), .CLK(clk), .RST(rst), .Q(
        start_reg[443]) );
  DFF \start_reg_reg[444]  ( .D(start_in[443]), .CLK(clk), .RST(rst), .Q(
        start_reg[444]) );
  DFF \start_reg_reg[445]  ( .D(start_in[444]), .CLK(clk), .RST(rst), .Q(
        start_reg[445]) );
  DFF \start_reg_reg[446]  ( .D(start_in[445]), .CLK(clk), .RST(rst), .Q(
        start_reg[446]) );
  DFF \start_reg_reg[447]  ( .D(start_in[446]), .CLK(clk), .RST(rst), .Q(
        start_reg[447]) );
  DFF \start_reg_reg[448]  ( .D(start_in[447]), .CLK(clk), .RST(rst), .Q(
        start_reg[448]) );
  DFF \start_reg_reg[449]  ( .D(start_in[448]), .CLK(clk), .RST(rst), .Q(
        start_reg[449]) );
  DFF \start_reg_reg[450]  ( .D(start_in[449]), .CLK(clk), .RST(rst), .Q(
        start_reg[450]) );
  DFF \start_reg_reg[451]  ( .D(start_in[450]), .CLK(clk), .RST(rst), .Q(
        start_reg[451]) );
  DFF \start_reg_reg[452]  ( .D(start_in[451]), .CLK(clk), .RST(rst), .Q(
        start_reg[452]) );
  DFF \start_reg_reg[453]  ( .D(start_in[452]), .CLK(clk), .RST(rst), .Q(
        start_reg[453]) );
  DFF \start_reg_reg[454]  ( .D(start_in[453]), .CLK(clk), .RST(rst), .Q(
        start_reg[454]) );
  DFF \start_reg_reg[455]  ( .D(start_in[454]), .CLK(clk), .RST(rst), .Q(
        start_reg[455]) );
  DFF \start_reg_reg[456]  ( .D(start_in[455]), .CLK(clk), .RST(rst), .Q(
        start_reg[456]) );
  DFF \start_reg_reg[457]  ( .D(start_in[456]), .CLK(clk), .RST(rst), .Q(
        start_reg[457]) );
  DFF \start_reg_reg[458]  ( .D(start_in[457]), .CLK(clk), .RST(rst), .Q(
        start_reg[458]) );
  DFF \start_reg_reg[459]  ( .D(start_in[458]), .CLK(clk), .RST(rst), .Q(
        start_reg[459]) );
  DFF \start_reg_reg[460]  ( .D(start_in[459]), .CLK(clk), .RST(rst), .Q(
        start_reg[460]) );
  DFF \start_reg_reg[461]  ( .D(start_in[460]), .CLK(clk), .RST(rst), .Q(
        start_reg[461]) );
  DFF \start_reg_reg[462]  ( .D(start_in[461]), .CLK(clk), .RST(rst), .Q(
        start_reg[462]) );
  DFF \start_reg_reg[463]  ( .D(start_in[462]), .CLK(clk), .RST(rst), .Q(
        start_reg[463]) );
  DFF \start_reg_reg[464]  ( .D(start_in[463]), .CLK(clk), .RST(rst), .Q(
        start_reg[464]) );
  DFF \start_reg_reg[465]  ( .D(start_in[464]), .CLK(clk), .RST(rst), .Q(
        start_reg[465]) );
  DFF \start_reg_reg[466]  ( .D(start_in[465]), .CLK(clk), .RST(rst), .Q(
        start_reg[466]) );
  DFF \start_reg_reg[467]  ( .D(start_in[466]), .CLK(clk), .RST(rst), .Q(
        start_reg[467]) );
  DFF \start_reg_reg[468]  ( .D(start_in[467]), .CLK(clk), .RST(rst), .Q(
        start_reg[468]) );
  DFF \start_reg_reg[469]  ( .D(start_in[468]), .CLK(clk), .RST(rst), .Q(
        start_reg[469]) );
  DFF \start_reg_reg[470]  ( .D(start_in[469]), .CLK(clk), .RST(rst), .Q(
        start_reg[470]) );
  DFF \start_reg_reg[471]  ( .D(start_in[470]), .CLK(clk), .RST(rst), .Q(
        start_reg[471]) );
  DFF \start_reg_reg[472]  ( .D(start_in[471]), .CLK(clk), .RST(rst), .Q(
        start_reg[472]) );
  DFF \start_reg_reg[473]  ( .D(start_in[472]), .CLK(clk), .RST(rst), .Q(
        start_reg[473]) );
  DFF \start_reg_reg[474]  ( .D(start_in[473]), .CLK(clk), .RST(rst), .Q(
        start_reg[474]) );
  DFF \start_reg_reg[475]  ( .D(start_in[474]), .CLK(clk), .RST(rst), .Q(
        start_reg[475]) );
  DFF \start_reg_reg[476]  ( .D(start_in[475]), .CLK(clk), .RST(rst), .Q(
        start_reg[476]) );
  DFF \start_reg_reg[477]  ( .D(start_in[476]), .CLK(clk), .RST(rst), .Q(
        start_reg[477]) );
  DFF \start_reg_reg[478]  ( .D(start_in[477]), .CLK(clk), .RST(rst), .Q(
        start_reg[478]) );
  DFF \start_reg_reg[479]  ( .D(start_in[478]), .CLK(clk), .RST(rst), .Q(
        start_reg[479]) );
  DFF \start_reg_reg[480]  ( .D(start_in[479]), .CLK(clk), .RST(rst), .Q(
        start_reg[480]) );
  DFF \start_reg_reg[481]  ( .D(start_in[480]), .CLK(clk), .RST(rst), .Q(
        start_reg[481]) );
  DFF \start_reg_reg[482]  ( .D(start_in[481]), .CLK(clk), .RST(rst), .Q(
        start_reg[482]) );
  DFF \start_reg_reg[483]  ( .D(start_in[482]), .CLK(clk), .RST(rst), .Q(
        start_reg[483]) );
  DFF \start_reg_reg[484]  ( .D(start_in[483]), .CLK(clk), .RST(rst), .Q(
        start_reg[484]) );
  DFF \start_reg_reg[485]  ( .D(start_in[484]), .CLK(clk), .RST(rst), .Q(
        start_reg[485]) );
  DFF \start_reg_reg[486]  ( .D(start_in[485]), .CLK(clk), .RST(rst), .Q(
        start_reg[486]) );
  DFF \start_reg_reg[487]  ( .D(start_in[486]), .CLK(clk), .RST(rst), .Q(
        start_reg[487]) );
  DFF \start_reg_reg[488]  ( .D(start_in[487]), .CLK(clk), .RST(rst), .Q(
        start_reg[488]) );
  DFF \start_reg_reg[489]  ( .D(start_in[488]), .CLK(clk), .RST(rst), .Q(
        start_reg[489]) );
  DFF \start_reg_reg[490]  ( .D(start_in[489]), .CLK(clk), .RST(rst), .Q(
        start_reg[490]) );
  DFF \start_reg_reg[491]  ( .D(start_in[490]), .CLK(clk), .RST(rst), .Q(
        start_reg[491]) );
  DFF \start_reg_reg[492]  ( .D(start_in[491]), .CLK(clk), .RST(rst), .Q(
        start_reg[492]) );
  DFF \start_reg_reg[493]  ( .D(start_in[492]), .CLK(clk), .RST(rst), .Q(
        start_reg[493]) );
  DFF \start_reg_reg[494]  ( .D(start_in[493]), .CLK(clk), .RST(rst), .Q(
        start_reg[494]) );
  DFF \start_reg_reg[495]  ( .D(start_in[494]), .CLK(clk), .RST(rst), .Q(
        start_reg[495]) );
  DFF \start_reg_reg[496]  ( .D(start_in[495]), .CLK(clk), .RST(rst), .Q(
        start_reg[496]) );
  DFF \start_reg_reg[497]  ( .D(start_in[496]), .CLK(clk), .RST(rst), .Q(
        start_reg[497]) );
  DFF \start_reg_reg[498]  ( .D(start_in[497]), .CLK(clk), .RST(rst), .Q(
        start_reg[498]) );
  DFF \start_reg_reg[499]  ( .D(start_in[498]), .CLK(clk), .RST(rst), .Q(
        start_reg[499]) );
  DFF \start_reg_reg[500]  ( .D(start_in[499]), .CLK(clk), .RST(rst), .Q(
        start_reg[500]) );
  DFF \start_reg_reg[501]  ( .D(start_in[500]), .CLK(clk), .RST(rst), .Q(
        start_reg[501]) );
  DFF \start_reg_reg[502]  ( .D(start_in[501]), .CLK(clk), .RST(rst), .Q(
        start_reg[502]) );
  DFF \start_reg_reg[503]  ( .D(start_in[502]), .CLK(clk), .RST(rst), .Q(
        start_reg[503]) );
  DFF \start_reg_reg[504]  ( .D(start_in[503]), .CLK(clk), .RST(rst), .Q(
        start_reg[504]) );
  DFF \start_reg_reg[505]  ( .D(start_in[504]), .CLK(clk), .RST(rst), .Q(
        start_reg[505]) );
  DFF \start_reg_reg[506]  ( .D(start_in[505]), .CLK(clk), .RST(rst), .Q(
        start_reg[506]) );
  DFF \start_reg_reg[507]  ( .D(start_in[506]), .CLK(clk), .RST(rst), .Q(
        start_reg[507]) );
  DFF \start_reg_reg[508]  ( .D(start_in[507]), .CLK(clk), .RST(rst), .Q(
        start_reg[508]) );
  DFF \start_reg_reg[509]  ( .D(start_in[508]), .CLK(clk), .RST(rst), .Q(
        start_reg[509]) );
  DFF \start_reg_reg[510]  ( .D(start_in[509]), .CLK(clk), .RST(rst), .Q(
        start_reg[510]) );
  DFF \start_reg_reg[511]  ( .D(start_in[510]), .CLK(clk), .RST(rst), .Q(
        start_reg[511]) );
  DFF mul_pow_reg ( .D(n2315), .CLK(clk), .RST(rst), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(n2314), .CLK(clk), .RST(rst), .Q(ereg[0]) );
  DFF \ereg_reg[1]  ( .D(n2313), .CLK(clk), .RST(rst), .Q(ereg[1]) );
  DFF \ereg_reg[2]  ( .D(n2312), .CLK(clk), .RST(rst), .Q(ereg[2]) );
  DFF \ereg_reg[3]  ( .D(n2311), .CLK(clk), .RST(rst), .Q(ereg[3]) );
  DFF \ereg_reg[4]  ( .D(n2310), .CLK(clk), .RST(rst), .Q(ereg[4]) );
  DFF \ereg_reg[5]  ( .D(n2309), .CLK(clk), .RST(rst), .Q(ereg[5]) );
  DFF \ereg_reg[6]  ( .D(n2308), .CLK(clk), .RST(rst), .Q(ereg[6]) );
  DFF \ereg_reg[7]  ( .D(n2307), .CLK(clk), .RST(rst), .Q(ereg[7]) );
  DFF \ereg_reg[8]  ( .D(n2306), .CLK(clk), .RST(rst), .Q(ereg[8]) );
  DFF \ereg_reg[9]  ( .D(n2305), .CLK(clk), .RST(rst), .Q(ereg[9]) );
  DFF \ereg_reg[10]  ( .D(n2304), .CLK(clk), .RST(rst), .Q(ereg[10]) );
  DFF \ereg_reg[11]  ( .D(n2303), .CLK(clk), .RST(rst), .Q(ereg[11]) );
  DFF \ereg_reg[12]  ( .D(n2302), .CLK(clk), .RST(rst), .Q(ereg[12]) );
  DFF \ereg_reg[13]  ( .D(n2301), .CLK(clk), .RST(rst), .Q(ereg[13]) );
  DFF \ereg_reg[14]  ( .D(n2300), .CLK(clk), .RST(rst), .Q(ereg[14]) );
  DFF \ereg_reg[15]  ( .D(n2299), .CLK(clk), .RST(rst), .Q(ereg[15]) );
  DFF \ereg_reg[16]  ( .D(n2298), .CLK(clk), .RST(rst), .Q(ereg[16]) );
  DFF \ereg_reg[17]  ( .D(n2297), .CLK(clk), .RST(rst), .Q(ereg[17]) );
  DFF \ereg_reg[18]  ( .D(n2296), .CLK(clk), .RST(rst), .Q(ereg[18]) );
  DFF \ereg_reg[19]  ( .D(n2295), .CLK(clk), .RST(rst), .Q(ereg[19]) );
  DFF \ereg_reg[20]  ( .D(n2294), .CLK(clk), .RST(rst), .Q(ereg[20]) );
  DFF \ereg_reg[21]  ( .D(n2293), .CLK(clk), .RST(rst), .Q(ereg[21]) );
  DFF \ereg_reg[22]  ( .D(n2292), .CLK(clk), .RST(rst), .Q(ereg[22]) );
  DFF \ereg_reg[23]  ( .D(n2291), .CLK(clk), .RST(rst), .Q(ereg[23]) );
  DFF \ereg_reg[24]  ( .D(n2290), .CLK(clk), .RST(rst), .Q(ereg[24]) );
  DFF \ereg_reg[25]  ( .D(n2289), .CLK(clk), .RST(rst), .Q(ereg[25]) );
  DFF \ereg_reg[26]  ( .D(n2288), .CLK(clk), .RST(rst), .Q(ereg[26]) );
  DFF \ereg_reg[27]  ( .D(n2287), .CLK(clk), .RST(rst), .Q(ereg[27]) );
  DFF \ereg_reg[28]  ( .D(n2286), .CLK(clk), .RST(rst), .Q(ereg[28]) );
  DFF \ereg_reg[29]  ( .D(n2285), .CLK(clk), .RST(rst), .Q(ereg[29]) );
  DFF \ereg_reg[30]  ( .D(n2284), .CLK(clk), .RST(rst), .Q(ereg[30]) );
  DFF \ereg_reg[31]  ( .D(n2283), .CLK(clk), .RST(rst), .Q(ereg[31]) );
  DFF \ereg_reg[32]  ( .D(n2282), .CLK(clk), .RST(rst), .Q(ereg[32]) );
  DFF \ereg_reg[33]  ( .D(n2281), .CLK(clk), .RST(rst), .Q(ereg[33]) );
  DFF \ereg_reg[34]  ( .D(n2280), .CLK(clk), .RST(rst), .Q(ereg[34]) );
  DFF \ereg_reg[35]  ( .D(n2279), .CLK(clk), .RST(rst), .Q(ereg[35]) );
  DFF \ereg_reg[36]  ( .D(n2278), .CLK(clk), .RST(rst), .Q(ereg[36]) );
  DFF \ereg_reg[37]  ( .D(n2277), .CLK(clk), .RST(rst), .Q(ereg[37]) );
  DFF \ereg_reg[38]  ( .D(n2276), .CLK(clk), .RST(rst), .Q(ereg[38]) );
  DFF \ereg_reg[39]  ( .D(n2275), .CLK(clk), .RST(rst), .Q(ereg[39]) );
  DFF \ereg_reg[40]  ( .D(n2274), .CLK(clk), .RST(rst), .Q(ereg[40]) );
  DFF \ereg_reg[41]  ( .D(n2273), .CLK(clk), .RST(rst), .Q(ereg[41]) );
  DFF \ereg_reg[42]  ( .D(n2272), .CLK(clk), .RST(rst), .Q(ereg[42]) );
  DFF \ereg_reg[43]  ( .D(n2271), .CLK(clk), .RST(rst), .Q(ereg[43]) );
  DFF \ereg_reg[44]  ( .D(n2270), .CLK(clk), .RST(rst), .Q(ereg[44]) );
  DFF \ereg_reg[45]  ( .D(n2269), .CLK(clk), .RST(rst), .Q(ereg[45]) );
  DFF \ereg_reg[46]  ( .D(n2268), .CLK(clk), .RST(rst), .Q(ereg[46]) );
  DFF \ereg_reg[47]  ( .D(n2267), .CLK(clk), .RST(rst), .Q(ereg[47]) );
  DFF \ereg_reg[48]  ( .D(n2266), .CLK(clk), .RST(rst), .Q(ereg[48]) );
  DFF \ereg_reg[49]  ( .D(n2265), .CLK(clk), .RST(rst), .Q(ereg[49]) );
  DFF \ereg_reg[50]  ( .D(n2264), .CLK(clk), .RST(rst), .Q(ereg[50]) );
  DFF \ereg_reg[51]  ( .D(n2263), .CLK(clk), .RST(rst), .Q(ereg[51]) );
  DFF \ereg_reg[52]  ( .D(n2262), .CLK(clk), .RST(rst), .Q(ereg[52]) );
  DFF \ereg_reg[53]  ( .D(n2261), .CLK(clk), .RST(rst), .Q(ereg[53]) );
  DFF \ereg_reg[54]  ( .D(n2260), .CLK(clk), .RST(rst), .Q(ereg[54]) );
  DFF \ereg_reg[55]  ( .D(n2259), .CLK(clk), .RST(rst), .Q(ereg[55]) );
  DFF \ereg_reg[56]  ( .D(n2258), .CLK(clk), .RST(rst), .Q(ereg[56]) );
  DFF \ereg_reg[57]  ( .D(n2257), .CLK(clk), .RST(rst), .Q(ereg[57]) );
  DFF \ereg_reg[58]  ( .D(n2256), .CLK(clk), .RST(rst), .Q(ereg[58]) );
  DFF \ereg_reg[59]  ( .D(n2255), .CLK(clk), .RST(rst), .Q(ereg[59]) );
  DFF \ereg_reg[60]  ( .D(n2254), .CLK(clk), .RST(rst), .Q(ereg[60]) );
  DFF \ereg_reg[61]  ( .D(n2253), .CLK(clk), .RST(rst), .Q(ereg[61]) );
  DFF \ereg_reg[62]  ( .D(n2252), .CLK(clk), .RST(rst), .Q(ereg[62]) );
  DFF \ereg_reg[63]  ( .D(n2251), .CLK(clk), .RST(rst), .Q(ereg[63]) );
  DFF \ereg_reg[64]  ( .D(n2250), .CLK(clk), .RST(rst), .Q(ereg[64]) );
  DFF \ereg_reg[65]  ( .D(n2249), .CLK(clk), .RST(rst), .Q(ereg[65]) );
  DFF \ereg_reg[66]  ( .D(n2248), .CLK(clk), .RST(rst), .Q(ereg[66]) );
  DFF \ereg_reg[67]  ( .D(n2247), .CLK(clk), .RST(rst), .Q(ereg[67]) );
  DFF \ereg_reg[68]  ( .D(n2246), .CLK(clk), .RST(rst), .Q(ereg[68]) );
  DFF \ereg_reg[69]  ( .D(n2245), .CLK(clk), .RST(rst), .Q(ereg[69]) );
  DFF \ereg_reg[70]  ( .D(n2244), .CLK(clk), .RST(rst), .Q(ereg[70]) );
  DFF \ereg_reg[71]  ( .D(n2243), .CLK(clk), .RST(rst), .Q(ereg[71]) );
  DFF \ereg_reg[72]  ( .D(n2242), .CLK(clk), .RST(rst), .Q(ereg[72]) );
  DFF \ereg_reg[73]  ( .D(n2241), .CLK(clk), .RST(rst), .Q(ereg[73]) );
  DFF \ereg_reg[74]  ( .D(n2240), .CLK(clk), .RST(rst), .Q(ereg[74]) );
  DFF \ereg_reg[75]  ( .D(n2239), .CLK(clk), .RST(rst), .Q(ereg[75]) );
  DFF \ereg_reg[76]  ( .D(n2238), .CLK(clk), .RST(rst), .Q(ereg[76]) );
  DFF \ereg_reg[77]  ( .D(n2237), .CLK(clk), .RST(rst), .Q(ereg[77]) );
  DFF \ereg_reg[78]  ( .D(n2236), .CLK(clk), .RST(rst), .Q(ereg[78]) );
  DFF \ereg_reg[79]  ( .D(n2235), .CLK(clk), .RST(rst), .Q(ereg[79]) );
  DFF \ereg_reg[80]  ( .D(n2234), .CLK(clk), .RST(rst), .Q(ereg[80]) );
  DFF \ereg_reg[81]  ( .D(n2233), .CLK(clk), .RST(rst), .Q(ereg[81]) );
  DFF \ereg_reg[82]  ( .D(n2232), .CLK(clk), .RST(rst), .Q(ereg[82]) );
  DFF \ereg_reg[83]  ( .D(n2231), .CLK(clk), .RST(rst), .Q(ereg[83]) );
  DFF \ereg_reg[84]  ( .D(n2230), .CLK(clk), .RST(rst), .Q(ereg[84]) );
  DFF \ereg_reg[85]  ( .D(n2229), .CLK(clk), .RST(rst), .Q(ereg[85]) );
  DFF \ereg_reg[86]  ( .D(n2228), .CLK(clk), .RST(rst), .Q(ereg[86]) );
  DFF \ereg_reg[87]  ( .D(n2227), .CLK(clk), .RST(rst), .Q(ereg[87]) );
  DFF \ereg_reg[88]  ( .D(n2226), .CLK(clk), .RST(rst), .Q(ereg[88]) );
  DFF \ereg_reg[89]  ( .D(n2225), .CLK(clk), .RST(rst), .Q(ereg[89]) );
  DFF \ereg_reg[90]  ( .D(n2224), .CLK(clk), .RST(rst), .Q(ereg[90]) );
  DFF \ereg_reg[91]  ( .D(n2223), .CLK(clk), .RST(rst), .Q(ereg[91]) );
  DFF \ereg_reg[92]  ( .D(n2222), .CLK(clk), .RST(rst), .Q(ereg[92]) );
  DFF \ereg_reg[93]  ( .D(n2221), .CLK(clk), .RST(rst), .Q(ereg[93]) );
  DFF \ereg_reg[94]  ( .D(n2220), .CLK(clk), .RST(rst), .Q(ereg[94]) );
  DFF \ereg_reg[95]  ( .D(n2219), .CLK(clk), .RST(rst), .Q(ereg[95]) );
  DFF \ereg_reg[96]  ( .D(n2218), .CLK(clk), .RST(rst), .Q(ereg[96]) );
  DFF \ereg_reg[97]  ( .D(n2217), .CLK(clk), .RST(rst), .Q(ereg[97]) );
  DFF \ereg_reg[98]  ( .D(n2216), .CLK(clk), .RST(rst), .Q(ereg[98]) );
  DFF \ereg_reg[99]  ( .D(n2215), .CLK(clk), .RST(rst), .Q(ereg[99]) );
  DFF \ereg_reg[100]  ( .D(n2214), .CLK(clk), .RST(rst), .Q(ereg[100]) );
  DFF \ereg_reg[101]  ( .D(n2213), .CLK(clk), .RST(rst), .Q(ereg[101]) );
  DFF \ereg_reg[102]  ( .D(n2212), .CLK(clk), .RST(rst), .Q(ereg[102]) );
  DFF \ereg_reg[103]  ( .D(n2211), .CLK(clk), .RST(rst), .Q(ereg[103]) );
  DFF \ereg_reg[104]  ( .D(n2210), .CLK(clk), .RST(rst), .Q(ereg[104]) );
  DFF \ereg_reg[105]  ( .D(n2209), .CLK(clk), .RST(rst), .Q(ereg[105]) );
  DFF \ereg_reg[106]  ( .D(n2208), .CLK(clk), .RST(rst), .Q(ereg[106]) );
  DFF \ereg_reg[107]  ( .D(n2207), .CLK(clk), .RST(rst), .Q(ereg[107]) );
  DFF \ereg_reg[108]  ( .D(n2206), .CLK(clk), .RST(rst), .Q(ereg[108]) );
  DFF \ereg_reg[109]  ( .D(n2205), .CLK(clk), .RST(rst), .Q(ereg[109]) );
  DFF \ereg_reg[110]  ( .D(n2204), .CLK(clk), .RST(rst), .Q(ereg[110]) );
  DFF \ereg_reg[111]  ( .D(n2203), .CLK(clk), .RST(rst), .Q(ereg[111]) );
  DFF \ereg_reg[112]  ( .D(n2202), .CLK(clk), .RST(rst), .Q(ereg[112]) );
  DFF \ereg_reg[113]  ( .D(n2201), .CLK(clk), .RST(rst), .Q(ereg[113]) );
  DFF \ereg_reg[114]  ( .D(n2200), .CLK(clk), .RST(rst), .Q(ereg[114]) );
  DFF \ereg_reg[115]  ( .D(n2199), .CLK(clk), .RST(rst), .Q(ereg[115]) );
  DFF \ereg_reg[116]  ( .D(n2198), .CLK(clk), .RST(rst), .Q(ereg[116]) );
  DFF \ereg_reg[117]  ( .D(n2197), .CLK(clk), .RST(rst), .Q(ereg[117]) );
  DFF \ereg_reg[118]  ( .D(n2196), .CLK(clk), .RST(rst), .Q(ereg[118]) );
  DFF \ereg_reg[119]  ( .D(n2195), .CLK(clk), .RST(rst), .Q(ereg[119]) );
  DFF \ereg_reg[120]  ( .D(n2194), .CLK(clk), .RST(rst), .Q(ereg[120]) );
  DFF \ereg_reg[121]  ( .D(n2193), .CLK(clk), .RST(rst), .Q(ereg[121]) );
  DFF \ereg_reg[122]  ( .D(n2192), .CLK(clk), .RST(rst), .Q(ereg[122]) );
  DFF \ereg_reg[123]  ( .D(n2191), .CLK(clk), .RST(rst), .Q(ereg[123]) );
  DFF \ereg_reg[124]  ( .D(n2190), .CLK(clk), .RST(rst), .Q(ereg[124]) );
  DFF \ereg_reg[125]  ( .D(n2189), .CLK(clk), .RST(rst), .Q(ereg[125]) );
  DFF \ereg_reg[126]  ( .D(n2188), .CLK(clk), .RST(rst), .Q(ereg[126]) );
  DFF \ereg_reg[127]  ( .D(n2187), .CLK(clk), .RST(rst), .Q(ereg[127]) );
  DFF \ereg_reg[128]  ( .D(n2186), .CLK(clk), .RST(rst), .Q(ereg[128]) );
  DFF \ereg_reg[129]  ( .D(n2185), .CLK(clk), .RST(rst), .Q(ereg[129]) );
  DFF \ereg_reg[130]  ( .D(n2184), .CLK(clk), .RST(rst), .Q(ereg[130]) );
  DFF \ereg_reg[131]  ( .D(n2183), .CLK(clk), .RST(rst), .Q(ereg[131]) );
  DFF \ereg_reg[132]  ( .D(n2182), .CLK(clk), .RST(rst), .Q(ereg[132]) );
  DFF \ereg_reg[133]  ( .D(n2181), .CLK(clk), .RST(rst), .Q(ereg[133]) );
  DFF \ereg_reg[134]  ( .D(n2180), .CLK(clk), .RST(rst), .Q(ereg[134]) );
  DFF \ereg_reg[135]  ( .D(n2179), .CLK(clk), .RST(rst), .Q(ereg[135]) );
  DFF \ereg_reg[136]  ( .D(n2178), .CLK(clk), .RST(rst), .Q(ereg[136]) );
  DFF \ereg_reg[137]  ( .D(n2177), .CLK(clk), .RST(rst), .Q(ereg[137]) );
  DFF \ereg_reg[138]  ( .D(n2176), .CLK(clk), .RST(rst), .Q(ereg[138]) );
  DFF \ereg_reg[139]  ( .D(n2175), .CLK(clk), .RST(rst), .Q(ereg[139]) );
  DFF \ereg_reg[140]  ( .D(n2174), .CLK(clk), .RST(rst), .Q(ereg[140]) );
  DFF \ereg_reg[141]  ( .D(n2173), .CLK(clk), .RST(rst), .Q(ereg[141]) );
  DFF \ereg_reg[142]  ( .D(n2172), .CLK(clk), .RST(rst), .Q(ereg[142]) );
  DFF \ereg_reg[143]  ( .D(n2171), .CLK(clk), .RST(rst), .Q(ereg[143]) );
  DFF \ereg_reg[144]  ( .D(n2170), .CLK(clk), .RST(rst), .Q(ereg[144]) );
  DFF \ereg_reg[145]  ( .D(n2169), .CLK(clk), .RST(rst), .Q(ereg[145]) );
  DFF \ereg_reg[146]  ( .D(n2168), .CLK(clk), .RST(rst), .Q(ereg[146]) );
  DFF \ereg_reg[147]  ( .D(n2167), .CLK(clk), .RST(rst), .Q(ereg[147]) );
  DFF \ereg_reg[148]  ( .D(n2166), .CLK(clk), .RST(rst), .Q(ereg[148]) );
  DFF \ereg_reg[149]  ( .D(n2165), .CLK(clk), .RST(rst), .Q(ereg[149]) );
  DFF \ereg_reg[150]  ( .D(n2164), .CLK(clk), .RST(rst), .Q(ereg[150]) );
  DFF \ereg_reg[151]  ( .D(n2163), .CLK(clk), .RST(rst), .Q(ereg[151]) );
  DFF \ereg_reg[152]  ( .D(n2162), .CLK(clk), .RST(rst), .Q(ereg[152]) );
  DFF \ereg_reg[153]  ( .D(n2161), .CLK(clk), .RST(rst), .Q(ereg[153]) );
  DFF \ereg_reg[154]  ( .D(n2160), .CLK(clk), .RST(rst), .Q(ereg[154]) );
  DFF \ereg_reg[155]  ( .D(n2159), .CLK(clk), .RST(rst), .Q(ereg[155]) );
  DFF \ereg_reg[156]  ( .D(n2158), .CLK(clk), .RST(rst), .Q(ereg[156]) );
  DFF \ereg_reg[157]  ( .D(n2157), .CLK(clk), .RST(rst), .Q(ereg[157]) );
  DFF \ereg_reg[158]  ( .D(n2156), .CLK(clk), .RST(rst), .Q(ereg[158]) );
  DFF \ereg_reg[159]  ( .D(n2155), .CLK(clk), .RST(rst), .Q(ereg[159]) );
  DFF \ereg_reg[160]  ( .D(n2154), .CLK(clk), .RST(rst), .Q(ereg[160]) );
  DFF \ereg_reg[161]  ( .D(n2153), .CLK(clk), .RST(rst), .Q(ereg[161]) );
  DFF \ereg_reg[162]  ( .D(n2152), .CLK(clk), .RST(rst), .Q(ereg[162]) );
  DFF \ereg_reg[163]  ( .D(n2151), .CLK(clk), .RST(rst), .Q(ereg[163]) );
  DFF \ereg_reg[164]  ( .D(n2150), .CLK(clk), .RST(rst), .Q(ereg[164]) );
  DFF \ereg_reg[165]  ( .D(n2149), .CLK(clk), .RST(rst), .Q(ereg[165]) );
  DFF \ereg_reg[166]  ( .D(n2148), .CLK(clk), .RST(rst), .Q(ereg[166]) );
  DFF \ereg_reg[167]  ( .D(n2147), .CLK(clk), .RST(rst), .Q(ereg[167]) );
  DFF \ereg_reg[168]  ( .D(n2146), .CLK(clk), .RST(rst), .Q(ereg[168]) );
  DFF \ereg_reg[169]  ( .D(n2145), .CLK(clk), .RST(rst), .Q(ereg[169]) );
  DFF \ereg_reg[170]  ( .D(n2144), .CLK(clk), .RST(rst), .Q(ereg[170]) );
  DFF \ereg_reg[171]  ( .D(n2143), .CLK(clk), .RST(rst), .Q(ereg[171]) );
  DFF \ereg_reg[172]  ( .D(n2142), .CLK(clk), .RST(rst), .Q(ereg[172]) );
  DFF \ereg_reg[173]  ( .D(n2141), .CLK(clk), .RST(rst), .Q(ereg[173]) );
  DFF \ereg_reg[174]  ( .D(n2140), .CLK(clk), .RST(rst), .Q(ereg[174]) );
  DFF \ereg_reg[175]  ( .D(n2139), .CLK(clk), .RST(rst), .Q(ereg[175]) );
  DFF \ereg_reg[176]  ( .D(n2138), .CLK(clk), .RST(rst), .Q(ereg[176]) );
  DFF \ereg_reg[177]  ( .D(n2137), .CLK(clk), .RST(rst), .Q(ereg[177]) );
  DFF \ereg_reg[178]  ( .D(n2136), .CLK(clk), .RST(rst), .Q(ereg[178]) );
  DFF \ereg_reg[179]  ( .D(n2135), .CLK(clk), .RST(rst), .Q(ereg[179]) );
  DFF \ereg_reg[180]  ( .D(n2134), .CLK(clk), .RST(rst), .Q(ereg[180]) );
  DFF \ereg_reg[181]  ( .D(n2133), .CLK(clk), .RST(rst), .Q(ereg[181]) );
  DFF \ereg_reg[182]  ( .D(n2132), .CLK(clk), .RST(rst), .Q(ereg[182]) );
  DFF \ereg_reg[183]  ( .D(n2131), .CLK(clk), .RST(rst), .Q(ereg[183]) );
  DFF \ereg_reg[184]  ( .D(n2130), .CLK(clk), .RST(rst), .Q(ereg[184]) );
  DFF \ereg_reg[185]  ( .D(n2129), .CLK(clk), .RST(rst), .Q(ereg[185]) );
  DFF \ereg_reg[186]  ( .D(n2128), .CLK(clk), .RST(rst), .Q(ereg[186]) );
  DFF \ereg_reg[187]  ( .D(n2127), .CLK(clk), .RST(rst), .Q(ereg[187]) );
  DFF \ereg_reg[188]  ( .D(n2126), .CLK(clk), .RST(rst), .Q(ereg[188]) );
  DFF \ereg_reg[189]  ( .D(n2125), .CLK(clk), .RST(rst), .Q(ereg[189]) );
  DFF \ereg_reg[190]  ( .D(n2124), .CLK(clk), .RST(rst), .Q(ereg[190]) );
  DFF \ereg_reg[191]  ( .D(n2123), .CLK(clk), .RST(rst), .Q(ereg[191]) );
  DFF \ereg_reg[192]  ( .D(n2122), .CLK(clk), .RST(rst), .Q(ereg[192]) );
  DFF \ereg_reg[193]  ( .D(n2121), .CLK(clk), .RST(rst), .Q(ereg[193]) );
  DFF \ereg_reg[194]  ( .D(n2120), .CLK(clk), .RST(rst), .Q(ereg[194]) );
  DFF \ereg_reg[195]  ( .D(n2119), .CLK(clk), .RST(rst), .Q(ereg[195]) );
  DFF \ereg_reg[196]  ( .D(n2118), .CLK(clk), .RST(rst), .Q(ereg[196]) );
  DFF \ereg_reg[197]  ( .D(n2117), .CLK(clk), .RST(rst), .Q(ereg[197]) );
  DFF \ereg_reg[198]  ( .D(n2116), .CLK(clk), .RST(rst), .Q(ereg[198]) );
  DFF \ereg_reg[199]  ( .D(n2115), .CLK(clk), .RST(rst), .Q(ereg[199]) );
  DFF \ereg_reg[200]  ( .D(n2114), .CLK(clk), .RST(rst), .Q(ereg[200]) );
  DFF \ereg_reg[201]  ( .D(n2113), .CLK(clk), .RST(rst), .Q(ereg[201]) );
  DFF \ereg_reg[202]  ( .D(n2112), .CLK(clk), .RST(rst), .Q(ereg[202]) );
  DFF \ereg_reg[203]  ( .D(n2111), .CLK(clk), .RST(rst), .Q(ereg[203]) );
  DFF \ereg_reg[204]  ( .D(n2110), .CLK(clk), .RST(rst), .Q(ereg[204]) );
  DFF \ereg_reg[205]  ( .D(n2109), .CLK(clk), .RST(rst), .Q(ereg[205]) );
  DFF \ereg_reg[206]  ( .D(n2108), .CLK(clk), .RST(rst), .Q(ereg[206]) );
  DFF \ereg_reg[207]  ( .D(n2107), .CLK(clk), .RST(rst), .Q(ereg[207]) );
  DFF \ereg_reg[208]  ( .D(n2106), .CLK(clk), .RST(rst), .Q(ereg[208]) );
  DFF \ereg_reg[209]  ( .D(n2105), .CLK(clk), .RST(rst), .Q(ereg[209]) );
  DFF \ereg_reg[210]  ( .D(n2104), .CLK(clk), .RST(rst), .Q(ereg[210]) );
  DFF \ereg_reg[211]  ( .D(n2103), .CLK(clk), .RST(rst), .Q(ereg[211]) );
  DFF \ereg_reg[212]  ( .D(n2102), .CLK(clk), .RST(rst), .Q(ereg[212]) );
  DFF \ereg_reg[213]  ( .D(n2101), .CLK(clk), .RST(rst), .Q(ereg[213]) );
  DFF \ereg_reg[214]  ( .D(n2100), .CLK(clk), .RST(rst), .Q(ereg[214]) );
  DFF \ereg_reg[215]  ( .D(n2099), .CLK(clk), .RST(rst), .Q(ereg[215]) );
  DFF \ereg_reg[216]  ( .D(n2098), .CLK(clk), .RST(rst), .Q(ereg[216]) );
  DFF \ereg_reg[217]  ( .D(n2097), .CLK(clk), .RST(rst), .Q(ereg[217]) );
  DFF \ereg_reg[218]  ( .D(n2096), .CLK(clk), .RST(rst), .Q(ereg[218]) );
  DFF \ereg_reg[219]  ( .D(n2095), .CLK(clk), .RST(rst), .Q(ereg[219]) );
  DFF \ereg_reg[220]  ( .D(n2094), .CLK(clk), .RST(rst), .Q(ereg[220]) );
  DFF \ereg_reg[221]  ( .D(n2093), .CLK(clk), .RST(rst), .Q(ereg[221]) );
  DFF \ereg_reg[222]  ( .D(n2092), .CLK(clk), .RST(rst), .Q(ereg[222]) );
  DFF \ereg_reg[223]  ( .D(n2091), .CLK(clk), .RST(rst), .Q(ereg[223]) );
  DFF \ereg_reg[224]  ( .D(n2090), .CLK(clk), .RST(rst), .Q(ereg[224]) );
  DFF \ereg_reg[225]  ( .D(n2089), .CLK(clk), .RST(rst), .Q(ereg[225]) );
  DFF \ereg_reg[226]  ( .D(n2088), .CLK(clk), .RST(rst), .Q(ereg[226]) );
  DFF \ereg_reg[227]  ( .D(n2087), .CLK(clk), .RST(rst), .Q(ereg[227]) );
  DFF \ereg_reg[228]  ( .D(n2086), .CLK(clk), .RST(rst), .Q(ereg[228]) );
  DFF \ereg_reg[229]  ( .D(n2085), .CLK(clk), .RST(rst), .Q(ereg[229]) );
  DFF \ereg_reg[230]  ( .D(n2084), .CLK(clk), .RST(rst), .Q(ereg[230]) );
  DFF \ereg_reg[231]  ( .D(n2083), .CLK(clk), .RST(rst), .Q(ereg[231]) );
  DFF \ereg_reg[232]  ( .D(n2082), .CLK(clk), .RST(rst), .Q(ereg[232]) );
  DFF \ereg_reg[233]  ( .D(n2081), .CLK(clk), .RST(rst), .Q(ereg[233]) );
  DFF \ereg_reg[234]  ( .D(n2080), .CLK(clk), .RST(rst), .Q(ereg[234]) );
  DFF \ereg_reg[235]  ( .D(n2079), .CLK(clk), .RST(rst), .Q(ereg[235]) );
  DFF \ereg_reg[236]  ( .D(n2078), .CLK(clk), .RST(rst), .Q(ereg[236]) );
  DFF \ereg_reg[237]  ( .D(n2077), .CLK(clk), .RST(rst), .Q(ereg[237]) );
  DFF \ereg_reg[238]  ( .D(n2076), .CLK(clk), .RST(rst), .Q(ereg[238]) );
  DFF \ereg_reg[239]  ( .D(n2075), .CLK(clk), .RST(rst), .Q(ereg[239]) );
  DFF \ereg_reg[240]  ( .D(n2074), .CLK(clk), .RST(rst), .Q(ereg[240]) );
  DFF \ereg_reg[241]  ( .D(n2073), .CLK(clk), .RST(rst), .Q(ereg[241]) );
  DFF \ereg_reg[242]  ( .D(n2072), .CLK(clk), .RST(rst), .Q(ereg[242]) );
  DFF \ereg_reg[243]  ( .D(n2071), .CLK(clk), .RST(rst), .Q(ereg[243]) );
  DFF \ereg_reg[244]  ( .D(n2070), .CLK(clk), .RST(rst), .Q(ereg[244]) );
  DFF \ereg_reg[245]  ( .D(n2069), .CLK(clk), .RST(rst), .Q(ereg[245]) );
  DFF \ereg_reg[246]  ( .D(n2068), .CLK(clk), .RST(rst), .Q(ereg[246]) );
  DFF \ereg_reg[247]  ( .D(n2067), .CLK(clk), .RST(rst), .Q(ereg[247]) );
  DFF \ereg_reg[248]  ( .D(n2066), .CLK(clk), .RST(rst), .Q(ereg[248]) );
  DFF \ereg_reg[249]  ( .D(n2065), .CLK(clk), .RST(rst), .Q(ereg[249]) );
  DFF \ereg_reg[250]  ( .D(n2064), .CLK(clk), .RST(rst), .Q(ereg[250]) );
  DFF \ereg_reg[251]  ( .D(n2063), .CLK(clk), .RST(rst), .Q(ereg[251]) );
  DFF \ereg_reg[252]  ( .D(n2062), .CLK(clk), .RST(rst), .Q(ereg[252]) );
  DFF \ereg_reg[253]  ( .D(n2061), .CLK(clk), .RST(rst), .Q(ereg[253]) );
  DFF \ereg_reg[254]  ( .D(n2060), .CLK(clk), .RST(rst), .Q(ereg[254]) );
  DFF \ereg_reg[255]  ( .D(n2059), .CLK(clk), .RST(rst), .Q(ereg[255]) );
  DFF first_one_reg ( .D(n2058), .CLK(clk), .RST(rst), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(n2057), .CLK(clk), .RST(rst), .Q(creg[0]) );
  DFF \creg_reg[1]  ( .D(n2056), .CLK(clk), .RST(rst), .Q(creg[1]) );
  DFF \creg_reg[2]  ( .D(n2055), .CLK(clk), .RST(rst), .Q(creg[2]) );
  DFF \creg_reg[3]  ( .D(n2054), .CLK(clk), .RST(rst), .Q(creg[3]) );
  DFF \creg_reg[4]  ( .D(n2053), .CLK(clk), .RST(rst), .Q(creg[4]) );
  DFF \creg_reg[5]  ( .D(n2052), .CLK(clk), .RST(rst), .Q(creg[5]) );
  DFF \creg_reg[6]  ( .D(n2051), .CLK(clk), .RST(rst), .Q(creg[6]) );
  DFF \creg_reg[7]  ( .D(n2050), .CLK(clk), .RST(rst), .Q(creg[7]) );
  DFF \creg_reg[8]  ( .D(n2049), .CLK(clk), .RST(rst), .Q(creg[8]) );
  DFF \creg_reg[9]  ( .D(n2048), .CLK(clk), .RST(rst), .Q(creg[9]) );
  DFF \creg_reg[10]  ( .D(n2047), .CLK(clk), .RST(rst), .Q(creg[10]) );
  DFF \creg_reg[11]  ( .D(n2046), .CLK(clk), .RST(rst), .Q(creg[11]) );
  DFF \creg_reg[12]  ( .D(n2045), .CLK(clk), .RST(rst), .Q(creg[12]) );
  DFF \creg_reg[13]  ( .D(n2044), .CLK(clk), .RST(rst), .Q(creg[13]) );
  DFF \creg_reg[14]  ( .D(n2043), .CLK(clk), .RST(rst), .Q(creg[14]) );
  DFF \creg_reg[15]  ( .D(n2042), .CLK(clk), .RST(rst), .Q(creg[15]) );
  DFF \creg_reg[16]  ( .D(n2041), .CLK(clk), .RST(rst), .Q(creg[16]) );
  DFF \creg_reg[17]  ( .D(n2040), .CLK(clk), .RST(rst), .Q(creg[17]) );
  DFF \creg_reg[18]  ( .D(n2039), .CLK(clk), .RST(rst), .Q(creg[18]) );
  DFF \creg_reg[19]  ( .D(n2038), .CLK(clk), .RST(rst), .Q(creg[19]) );
  DFF \creg_reg[20]  ( .D(n2037), .CLK(clk), .RST(rst), .Q(creg[20]) );
  DFF \creg_reg[21]  ( .D(n2036), .CLK(clk), .RST(rst), .Q(creg[21]) );
  DFF \creg_reg[22]  ( .D(n2035), .CLK(clk), .RST(rst), .Q(creg[22]) );
  DFF \creg_reg[23]  ( .D(n2034), .CLK(clk), .RST(rst), .Q(creg[23]) );
  DFF \creg_reg[24]  ( .D(n2033), .CLK(clk), .RST(rst), .Q(creg[24]) );
  DFF \creg_reg[25]  ( .D(n2032), .CLK(clk), .RST(rst), .Q(creg[25]) );
  DFF \creg_reg[26]  ( .D(n2031), .CLK(clk), .RST(rst), .Q(creg[26]) );
  DFF \creg_reg[27]  ( .D(n2030), .CLK(clk), .RST(rst), .Q(creg[27]) );
  DFF \creg_reg[28]  ( .D(n2029), .CLK(clk), .RST(rst), .Q(creg[28]) );
  DFF \creg_reg[29]  ( .D(n2028), .CLK(clk), .RST(rst), .Q(creg[29]) );
  DFF \creg_reg[30]  ( .D(n2027), .CLK(clk), .RST(rst), .Q(creg[30]) );
  DFF \creg_reg[31]  ( .D(n2026), .CLK(clk), .RST(rst), .Q(creg[31]) );
  DFF \creg_reg[32]  ( .D(n2025), .CLK(clk), .RST(rst), .Q(creg[32]) );
  DFF \creg_reg[33]  ( .D(n2024), .CLK(clk), .RST(rst), .Q(creg[33]) );
  DFF \creg_reg[34]  ( .D(n2023), .CLK(clk), .RST(rst), .Q(creg[34]) );
  DFF \creg_reg[35]  ( .D(n2022), .CLK(clk), .RST(rst), .Q(creg[35]) );
  DFF \creg_reg[36]  ( .D(n2021), .CLK(clk), .RST(rst), .Q(creg[36]) );
  DFF \creg_reg[37]  ( .D(n2020), .CLK(clk), .RST(rst), .Q(creg[37]) );
  DFF \creg_reg[38]  ( .D(n2019), .CLK(clk), .RST(rst), .Q(creg[38]) );
  DFF \creg_reg[39]  ( .D(n2018), .CLK(clk), .RST(rst), .Q(creg[39]) );
  DFF \creg_reg[40]  ( .D(n2017), .CLK(clk), .RST(rst), .Q(creg[40]) );
  DFF \creg_reg[41]  ( .D(n2016), .CLK(clk), .RST(rst), .Q(creg[41]) );
  DFF \creg_reg[42]  ( .D(n2015), .CLK(clk), .RST(rst), .Q(creg[42]) );
  DFF \creg_reg[43]  ( .D(n2014), .CLK(clk), .RST(rst), .Q(creg[43]) );
  DFF \creg_reg[44]  ( .D(n2013), .CLK(clk), .RST(rst), .Q(creg[44]) );
  DFF \creg_reg[45]  ( .D(n2012), .CLK(clk), .RST(rst), .Q(creg[45]) );
  DFF \creg_reg[46]  ( .D(n2011), .CLK(clk), .RST(rst), .Q(creg[46]) );
  DFF \creg_reg[47]  ( .D(n2010), .CLK(clk), .RST(rst), .Q(creg[47]) );
  DFF \creg_reg[48]  ( .D(n2009), .CLK(clk), .RST(rst), .Q(creg[48]) );
  DFF \creg_reg[49]  ( .D(n2008), .CLK(clk), .RST(rst), .Q(creg[49]) );
  DFF \creg_reg[50]  ( .D(n2007), .CLK(clk), .RST(rst), .Q(creg[50]) );
  DFF \creg_reg[51]  ( .D(n2006), .CLK(clk), .RST(rst), .Q(creg[51]) );
  DFF \creg_reg[52]  ( .D(n2005), .CLK(clk), .RST(rst), .Q(creg[52]) );
  DFF \creg_reg[53]  ( .D(n2004), .CLK(clk), .RST(rst), .Q(creg[53]) );
  DFF \creg_reg[54]  ( .D(n2003), .CLK(clk), .RST(rst), .Q(creg[54]) );
  DFF \creg_reg[55]  ( .D(n2002), .CLK(clk), .RST(rst), .Q(creg[55]) );
  DFF \creg_reg[56]  ( .D(n2001), .CLK(clk), .RST(rst), .Q(creg[56]) );
  DFF \creg_reg[57]  ( .D(n2000), .CLK(clk), .RST(rst), .Q(creg[57]) );
  DFF \creg_reg[58]  ( .D(n1999), .CLK(clk), .RST(rst), .Q(creg[58]) );
  DFF \creg_reg[59]  ( .D(n1998), .CLK(clk), .RST(rst), .Q(creg[59]) );
  DFF \creg_reg[60]  ( .D(n1997), .CLK(clk), .RST(rst), .Q(creg[60]) );
  DFF \creg_reg[61]  ( .D(n1996), .CLK(clk), .RST(rst), .Q(creg[61]) );
  DFF \creg_reg[62]  ( .D(n1995), .CLK(clk), .RST(rst), .Q(creg[62]) );
  DFF \creg_reg[63]  ( .D(n1994), .CLK(clk), .RST(rst), .Q(creg[63]) );
  DFF \creg_reg[64]  ( .D(n1993), .CLK(clk), .RST(rst), .Q(creg[64]) );
  DFF \creg_reg[65]  ( .D(n1992), .CLK(clk), .RST(rst), .Q(creg[65]) );
  DFF \creg_reg[66]  ( .D(n1991), .CLK(clk), .RST(rst), .Q(creg[66]) );
  DFF \creg_reg[67]  ( .D(n1990), .CLK(clk), .RST(rst), .Q(creg[67]) );
  DFF \creg_reg[68]  ( .D(n1989), .CLK(clk), .RST(rst), .Q(creg[68]) );
  DFF \creg_reg[69]  ( .D(n1988), .CLK(clk), .RST(rst), .Q(creg[69]) );
  DFF \creg_reg[70]  ( .D(n1987), .CLK(clk), .RST(rst), .Q(creg[70]) );
  DFF \creg_reg[71]  ( .D(n1986), .CLK(clk), .RST(rst), .Q(creg[71]) );
  DFF \creg_reg[72]  ( .D(n1985), .CLK(clk), .RST(rst), .Q(creg[72]) );
  DFF \creg_reg[73]  ( .D(n1984), .CLK(clk), .RST(rst), .Q(creg[73]) );
  DFF \creg_reg[74]  ( .D(n1983), .CLK(clk), .RST(rst), .Q(creg[74]) );
  DFF \creg_reg[75]  ( .D(n1982), .CLK(clk), .RST(rst), .Q(creg[75]) );
  DFF \creg_reg[76]  ( .D(n1981), .CLK(clk), .RST(rst), .Q(creg[76]) );
  DFF \creg_reg[77]  ( .D(n1980), .CLK(clk), .RST(rst), .Q(creg[77]) );
  DFF \creg_reg[78]  ( .D(n1979), .CLK(clk), .RST(rst), .Q(creg[78]) );
  DFF \creg_reg[79]  ( .D(n1978), .CLK(clk), .RST(rst), .Q(creg[79]) );
  DFF \creg_reg[80]  ( .D(n1977), .CLK(clk), .RST(rst), .Q(creg[80]) );
  DFF \creg_reg[81]  ( .D(n1976), .CLK(clk), .RST(rst), .Q(creg[81]) );
  DFF \creg_reg[82]  ( .D(n1975), .CLK(clk), .RST(rst), .Q(creg[82]) );
  DFF \creg_reg[83]  ( .D(n1974), .CLK(clk), .RST(rst), .Q(creg[83]) );
  DFF \creg_reg[84]  ( .D(n1973), .CLK(clk), .RST(rst), .Q(creg[84]) );
  DFF \creg_reg[85]  ( .D(n1972), .CLK(clk), .RST(rst), .Q(creg[85]) );
  DFF \creg_reg[86]  ( .D(n1971), .CLK(clk), .RST(rst), .Q(creg[86]) );
  DFF \creg_reg[87]  ( .D(n1970), .CLK(clk), .RST(rst), .Q(creg[87]) );
  DFF \creg_reg[88]  ( .D(n1969), .CLK(clk), .RST(rst), .Q(creg[88]) );
  DFF \creg_reg[89]  ( .D(n1968), .CLK(clk), .RST(rst), .Q(creg[89]) );
  DFF \creg_reg[90]  ( .D(n1967), .CLK(clk), .RST(rst), .Q(creg[90]) );
  DFF \creg_reg[91]  ( .D(n1966), .CLK(clk), .RST(rst), .Q(creg[91]) );
  DFF \creg_reg[92]  ( .D(n1965), .CLK(clk), .RST(rst), .Q(creg[92]) );
  DFF \creg_reg[93]  ( .D(n1964), .CLK(clk), .RST(rst), .Q(creg[93]) );
  DFF \creg_reg[94]  ( .D(n1963), .CLK(clk), .RST(rst), .Q(creg[94]) );
  DFF \creg_reg[95]  ( .D(n1962), .CLK(clk), .RST(rst), .Q(creg[95]) );
  DFF \creg_reg[96]  ( .D(n1961), .CLK(clk), .RST(rst), .Q(creg[96]) );
  DFF \creg_reg[97]  ( .D(n1960), .CLK(clk), .RST(rst), .Q(creg[97]) );
  DFF \creg_reg[98]  ( .D(n1959), .CLK(clk), .RST(rst), .Q(creg[98]) );
  DFF \creg_reg[99]  ( .D(n1958), .CLK(clk), .RST(rst), .Q(creg[99]) );
  DFF \creg_reg[100]  ( .D(n1957), .CLK(clk), .RST(rst), .Q(creg[100]) );
  DFF \creg_reg[101]  ( .D(n1956), .CLK(clk), .RST(rst), .Q(creg[101]) );
  DFF \creg_reg[102]  ( .D(n1955), .CLK(clk), .RST(rst), .Q(creg[102]) );
  DFF \creg_reg[103]  ( .D(n1954), .CLK(clk), .RST(rst), .Q(creg[103]) );
  DFF \creg_reg[104]  ( .D(n1953), .CLK(clk), .RST(rst), .Q(creg[104]) );
  DFF \creg_reg[105]  ( .D(n1952), .CLK(clk), .RST(rst), .Q(creg[105]) );
  DFF \creg_reg[106]  ( .D(n1951), .CLK(clk), .RST(rst), .Q(creg[106]) );
  DFF \creg_reg[107]  ( .D(n1950), .CLK(clk), .RST(rst), .Q(creg[107]) );
  DFF \creg_reg[108]  ( .D(n1949), .CLK(clk), .RST(rst), .Q(creg[108]) );
  DFF \creg_reg[109]  ( .D(n1948), .CLK(clk), .RST(rst), .Q(creg[109]) );
  DFF \creg_reg[110]  ( .D(n1947), .CLK(clk), .RST(rst), .Q(creg[110]) );
  DFF \creg_reg[111]  ( .D(n1946), .CLK(clk), .RST(rst), .Q(creg[111]) );
  DFF \creg_reg[112]  ( .D(n1945), .CLK(clk), .RST(rst), .Q(creg[112]) );
  DFF \creg_reg[113]  ( .D(n1944), .CLK(clk), .RST(rst), .Q(creg[113]) );
  DFF \creg_reg[114]  ( .D(n1943), .CLK(clk), .RST(rst), .Q(creg[114]) );
  DFF \creg_reg[115]  ( .D(n1942), .CLK(clk), .RST(rst), .Q(creg[115]) );
  DFF \creg_reg[116]  ( .D(n1941), .CLK(clk), .RST(rst), .Q(creg[116]) );
  DFF \creg_reg[117]  ( .D(n1940), .CLK(clk), .RST(rst), .Q(creg[117]) );
  DFF \creg_reg[118]  ( .D(n1939), .CLK(clk), .RST(rst), .Q(creg[118]) );
  DFF \creg_reg[119]  ( .D(n1938), .CLK(clk), .RST(rst), .Q(creg[119]) );
  DFF \creg_reg[120]  ( .D(n1937), .CLK(clk), .RST(rst), .Q(creg[120]) );
  DFF \creg_reg[121]  ( .D(n1936), .CLK(clk), .RST(rst), .Q(creg[121]) );
  DFF \creg_reg[122]  ( .D(n1935), .CLK(clk), .RST(rst), .Q(creg[122]) );
  DFF \creg_reg[123]  ( .D(n1934), .CLK(clk), .RST(rst), .Q(creg[123]) );
  DFF \creg_reg[124]  ( .D(n1933), .CLK(clk), .RST(rst), .Q(creg[124]) );
  DFF \creg_reg[125]  ( .D(n1932), .CLK(clk), .RST(rst), .Q(creg[125]) );
  DFF \creg_reg[126]  ( .D(n1931), .CLK(clk), .RST(rst), .Q(creg[126]) );
  DFF \creg_reg[127]  ( .D(n1930), .CLK(clk), .RST(rst), .Q(creg[127]) );
  DFF \creg_reg[128]  ( .D(n1929), .CLK(clk), .RST(rst), .Q(creg[128]) );
  DFF \creg_reg[129]  ( .D(n1928), .CLK(clk), .RST(rst), .Q(creg[129]) );
  DFF \creg_reg[130]  ( .D(n1927), .CLK(clk), .RST(rst), .Q(creg[130]) );
  DFF \creg_reg[131]  ( .D(n1926), .CLK(clk), .RST(rst), .Q(creg[131]) );
  DFF \creg_reg[132]  ( .D(n1925), .CLK(clk), .RST(rst), .Q(creg[132]) );
  DFF \creg_reg[133]  ( .D(n1924), .CLK(clk), .RST(rst), .Q(creg[133]) );
  DFF \creg_reg[134]  ( .D(n1923), .CLK(clk), .RST(rst), .Q(creg[134]) );
  DFF \creg_reg[135]  ( .D(n1922), .CLK(clk), .RST(rst), .Q(creg[135]) );
  DFF \creg_reg[136]  ( .D(n1921), .CLK(clk), .RST(rst), .Q(creg[136]) );
  DFF \creg_reg[137]  ( .D(n1920), .CLK(clk), .RST(rst), .Q(creg[137]) );
  DFF \creg_reg[138]  ( .D(n1919), .CLK(clk), .RST(rst), .Q(creg[138]) );
  DFF \creg_reg[139]  ( .D(n1918), .CLK(clk), .RST(rst), .Q(creg[139]) );
  DFF \creg_reg[140]  ( .D(n1917), .CLK(clk), .RST(rst), .Q(creg[140]) );
  DFF \creg_reg[141]  ( .D(n1916), .CLK(clk), .RST(rst), .Q(creg[141]) );
  DFF \creg_reg[142]  ( .D(n1915), .CLK(clk), .RST(rst), .Q(creg[142]) );
  DFF \creg_reg[143]  ( .D(n1914), .CLK(clk), .RST(rst), .Q(creg[143]) );
  DFF \creg_reg[144]  ( .D(n1913), .CLK(clk), .RST(rst), .Q(creg[144]) );
  DFF \creg_reg[145]  ( .D(n1912), .CLK(clk), .RST(rst), .Q(creg[145]) );
  DFF \creg_reg[146]  ( .D(n1911), .CLK(clk), .RST(rst), .Q(creg[146]) );
  DFF \creg_reg[147]  ( .D(n1910), .CLK(clk), .RST(rst), .Q(creg[147]) );
  DFF \creg_reg[148]  ( .D(n1909), .CLK(clk), .RST(rst), .Q(creg[148]) );
  DFF \creg_reg[149]  ( .D(n1908), .CLK(clk), .RST(rst), .Q(creg[149]) );
  DFF \creg_reg[150]  ( .D(n1907), .CLK(clk), .RST(rst), .Q(creg[150]) );
  DFF \creg_reg[151]  ( .D(n1906), .CLK(clk), .RST(rst), .Q(creg[151]) );
  DFF \creg_reg[152]  ( .D(n1905), .CLK(clk), .RST(rst), .Q(creg[152]) );
  DFF \creg_reg[153]  ( .D(n1904), .CLK(clk), .RST(rst), .Q(creg[153]) );
  DFF \creg_reg[154]  ( .D(n1903), .CLK(clk), .RST(rst), .Q(creg[154]) );
  DFF \creg_reg[155]  ( .D(n1902), .CLK(clk), .RST(rst), .Q(creg[155]) );
  DFF \creg_reg[156]  ( .D(n1901), .CLK(clk), .RST(rst), .Q(creg[156]) );
  DFF \creg_reg[157]  ( .D(n1900), .CLK(clk), .RST(rst), .Q(creg[157]) );
  DFF \creg_reg[158]  ( .D(n1899), .CLK(clk), .RST(rst), .Q(creg[158]) );
  DFF \creg_reg[159]  ( .D(n1898), .CLK(clk), .RST(rst), .Q(creg[159]) );
  DFF \creg_reg[160]  ( .D(n1897), .CLK(clk), .RST(rst), .Q(creg[160]) );
  DFF \creg_reg[161]  ( .D(n1896), .CLK(clk), .RST(rst), .Q(creg[161]) );
  DFF \creg_reg[162]  ( .D(n1895), .CLK(clk), .RST(rst), .Q(creg[162]) );
  DFF \creg_reg[163]  ( .D(n1894), .CLK(clk), .RST(rst), .Q(creg[163]) );
  DFF \creg_reg[164]  ( .D(n1893), .CLK(clk), .RST(rst), .Q(creg[164]) );
  DFF \creg_reg[165]  ( .D(n1892), .CLK(clk), .RST(rst), .Q(creg[165]) );
  DFF \creg_reg[166]  ( .D(n1891), .CLK(clk), .RST(rst), .Q(creg[166]) );
  DFF \creg_reg[167]  ( .D(n1890), .CLK(clk), .RST(rst), .Q(creg[167]) );
  DFF \creg_reg[168]  ( .D(n1889), .CLK(clk), .RST(rst), .Q(creg[168]) );
  DFF \creg_reg[169]  ( .D(n1888), .CLK(clk), .RST(rst), .Q(creg[169]) );
  DFF \creg_reg[170]  ( .D(n1887), .CLK(clk), .RST(rst), .Q(creg[170]) );
  DFF \creg_reg[171]  ( .D(n1886), .CLK(clk), .RST(rst), .Q(creg[171]) );
  DFF \creg_reg[172]  ( .D(n1885), .CLK(clk), .RST(rst), .Q(creg[172]) );
  DFF \creg_reg[173]  ( .D(n1884), .CLK(clk), .RST(rst), .Q(creg[173]) );
  DFF \creg_reg[174]  ( .D(n1883), .CLK(clk), .RST(rst), .Q(creg[174]) );
  DFF \creg_reg[175]  ( .D(n1882), .CLK(clk), .RST(rst), .Q(creg[175]) );
  DFF \creg_reg[176]  ( .D(n1881), .CLK(clk), .RST(rst), .Q(creg[176]) );
  DFF \creg_reg[177]  ( .D(n1880), .CLK(clk), .RST(rst), .Q(creg[177]) );
  DFF \creg_reg[178]  ( .D(n1879), .CLK(clk), .RST(rst), .Q(creg[178]) );
  DFF \creg_reg[179]  ( .D(n1878), .CLK(clk), .RST(rst), .Q(creg[179]) );
  DFF \creg_reg[180]  ( .D(n1877), .CLK(clk), .RST(rst), .Q(creg[180]) );
  DFF \creg_reg[181]  ( .D(n1876), .CLK(clk), .RST(rst), .Q(creg[181]) );
  DFF \creg_reg[182]  ( .D(n1875), .CLK(clk), .RST(rst), .Q(creg[182]) );
  DFF \creg_reg[183]  ( .D(n1874), .CLK(clk), .RST(rst), .Q(creg[183]) );
  DFF \creg_reg[184]  ( .D(n1873), .CLK(clk), .RST(rst), .Q(creg[184]) );
  DFF \creg_reg[185]  ( .D(n1872), .CLK(clk), .RST(rst), .Q(creg[185]) );
  DFF \creg_reg[186]  ( .D(n1871), .CLK(clk), .RST(rst), .Q(creg[186]) );
  DFF \creg_reg[187]  ( .D(n1870), .CLK(clk), .RST(rst), .Q(creg[187]) );
  DFF \creg_reg[188]  ( .D(n1869), .CLK(clk), .RST(rst), .Q(creg[188]) );
  DFF \creg_reg[189]  ( .D(n1868), .CLK(clk), .RST(rst), .Q(creg[189]) );
  DFF \creg_reg[190]  ( .D(n1867), .CLK(clk), .RST(rst), .Q(creg[190]) );
  DFF \creg_reg[191]  ( .D(n1866), .CLK(clk), .RST(rst), .Q(creg[191]) );
  DFF \creg_reg[192]  ( .D(n1865), .CLK(clk), .RST(rst), .Q(creg[192]) );
  DFF \creg_reg[193]  ( .D(n1864), .CLK(clk), .RST(rst), .Q(creg[193]) );
  DFF \creg_reg[194]  ( .D(n1863), .CLK(clk), .RST(rst), .Q(creg[194]) );
  DFF \creg_reg[195]  ( .D(n1862), .CLK(clk), .RST(rst), .Q(creg[195]) );
  DFF \creg_reg[196]  ( .D(n1861), .CLK(clk), .RST(rst), .Q(creg[196]) );
  DFF \creg_reg[197]  ( .D(n1860), .CLK(clk), .RST(rst), .Q(creg[197]) );
  DFF \creg_reg[198]  ( .D(n1859), .CLK(clk), .RST(rst), .Q(creg[198]) );
  DFF \creg_reg[199]  ( .D(n1858), .CLK(clk), .RST(rst), .Q(creg[199]) );
  DFF \creg_reg[200]  ( .D(n1857), .CLK(clk), .RST(rst), .Q(creg[200]) );
  DFF \creg_reg[201]  ( .D(n1856), .CLK(clk), .RST(rst), .Q(creg[201]) );
  DFF \creg_reg[202]  ( .D(n1855), .CLK(clk), .RST(rst), .Q(creg[202]) );
  DFF \creg_reg[203]  ( .D(n1854), .CLK(clk), .RST(rst), .Q(creg[203]) );
  DFF \creg_reg[204]  ( .D(n1853), .CLK(clk), .RST(rst), .Q(creg[204]) );
  DFF \creg_reg[205]  ( .D(n1852), .CLK(clk), .RST(rst), .Q(creg[205]) );
  DFF \creg_reg[206]  ( .D(n1851), .CLK(clk), .RST(rst), .Q(creg[206]) );
  DFF \creg_reg[207]  ( .D(n1850), .CLK(clk), .RST(rst), .Q(creg[207]) );
  DFF \creg_reg[208]  ( .D(n1849), .CLK(clk), .RST(rst), .Q(creg[208]) );
  DFF \creg_reg[209]  ( .D(n1848), .CLK(clk), .RST(rst), .Q(creg[209]) );
  DFF \creg_reg[210]  ( .D(n1847), .CLK(clk), .RST(rst), .Q(creg[210]) );
  DFF \creg_reg[211]  ( .D(n1846), .CLK(clk), .RST(rst), .Q(creg[211]) );
  DFF \creg_reg[212]  ( .D(n1845), .CLK(clk), .RST(rst), .Q(creg[212]) );
  DFF \creg_reg[213]  ( .D(n1844), .CLK(clk), .RST(rst), .Q(creg[213]) );
  DFF \creg_reg[214]  ( .D(n1843), .CLK(clk), .RST(rst), .Q(creg[214]) );
  DFF \creg_reg[215]  ( .D(n1842), .CLK(clk), .RST(rst), .Q(creg[215]) );
  DFF \creg_reg[216]  ( .D(n1841), .CLK(clk), .RST(rst), .Q(creg[216]) );
  DFF \creg_reg[217]  ( .D(n1840), .CLK(clk), .RST(rst), .Q(creg[217]) );
  DFF \creg_reg[218]  ( .D(n1839), .CLK(clk), .RST(rst), .Q(creg[218]) );
  DFF \creg_reg[219]  ( .D(n1838), .CLK(clk), .RST(rst), .Q(creg[219]) );
  DFF \creg_reg[220]  ( .D(n1837), .CLK(clk), .RST(rst), .Q(creg[220]) );
  DFF \creg_reg[221]  ( .D(n1836), .CLK(clk), .RST(rst), .Q(creg[221]) );
  DFF \creg_reg[222]  ( .D(n1835), .CLK(clk), .RST(rst), .Q(creg[222]) );
  DFF \creg_reg[223]  ( .D(n1834), .CLK(clk), .RST(rst), .Q(creg[223]) );
  DFF \creg_reg[224]  ( .D(n1833), .CLK(clk), .RST(rst), .Q(creg[224]) );
  DFF \creg_reg[225]  ( .D(n1832), .CLK(clk), .RST(rst), .Q(creg[225]) );
  DFF \creg_reg[226]  ( .D(n1831), .CLK(clk), .RST(rst), .Q(creg[226]) );
  DFF \creg_reg[227]  ( .D(n1830), .CLK(clk), .RST(rst), .Q(creg[227]) );
  DFF \creg_reg[228]  ( .D(n1829), .CLK(clk), .RST(rst), .Q(creg[228]) );
  DFF \creg_reg[229]  ( .D(n1828), .CLK(clk), .RST(rst), .Q(creg[229]) );
  DFF \creg_reg[230]  ( .D(n1827), .CLK(clk), .RST(rst), .Q(creg[230]) );
  DFF \creg_reg[231]  ( .D(n1826), .CLK(clk), .RST(rst), .Q(creg[231]) );
  DFF \creg_reg[232]  ( .D(n1825), .CLK(clk), .RST(rst), .Q(creg[232]) );
  DFF \creg_reg[233]  ( .D(n1824), .CLK(clk), .RST(rst), .Q(creg[233]) );
  DFF \creg_reg[234]  ( .D(n1823), .CLK(clk), .RST(rst), .Q(creg[234]) );
  DFF \creg_reg[235]  ( .D(n1822), .CLK(clk), .RST(rst), .Q(creg[235]) );
  DFF \creg_reg[236]  ( .D(n1821), .CLK(clk), .RST(rst), .Q(creg[236]) );
  DFF \creg_reg[237]  ( .D(n1820), .CLK(clk), .RST(rst), .Q(creg[237]) );
  DFF \creg_reg[238]  ( .D(n1819), .CLK(clk), .RST(rst), .Q(creg[238]) );
  DFF \creg_reg[239]  ( .D(n1818), .CLK(clk), .RST(rst), .Q(creg[239]) );
  DFF \creg_reg[240]  ( .D(n1817), .CLK(clk), .RST(rst), .Q(creg[240]) );
  DFF \creg_reg[241]  ( .D(n1816), .CLK(clk), .RST(rst), .Q(creg[241]) );
  DFF \creg_reg[242]  ( .D(n1815), .CLK(clk), .RST(rst), .Q(creg[242]) );
  DFF \creg_reg[243]  ( .D(n1814), .CLK(clk), .RST(rst), .Q(creg[243]) );
  DFF \creg_reg[244]  ( .D(n1813), .CLK(clk), .RST(rst), .Q(creg[244]) );
  DFF \creg_reg[245]  ( .D(n1812), .CLK(clk), .RST(rst), .Q(creg[245]) );
  DFF \creg_reg[246]  ( .D(n1811), .CLK(clk), .RST(rst), .Q(creg[246]) );
  DFF \creg_reg[247]  ( .D(n1810), .CLK(clk), .RST(rst), .Q(creg[247]) );
  DFF \creg_reg[248]  ( .D(n1809), .CLK(clk), .RST(rst), .Q(creg[248]) );
  DFF \creg_reg[249]  ( .D(n1808), .CLK(clk), .RST(rst), .Q(creg[249]) );
  DFF \creg_reg[250]  ( .D(n1807), .CLK(clk), .RST(rst), .Q(creg[250]) );
  DFF \creg_reg[251]  ( .D(n1806), .CLK(clk), .RST(rst), .Q(creg[251]) );
  DFF \creg_reg[252]  ( .D(n1805), .CLK(clk), .RST(rst), .Q(creg[252]) );
  DFF \creg_reg[253]  ( .D(n1804), .CLK(clk), .RST(rst), .Q(creg[253]) );
  DFF \creg_reg[254]  ( .D(n1803), .CLK(clk), .RST(rst), .Q(creg[254]) );
  DFF \creg_reg[255]  ( .D(n1802), .CLK(clk), .RST(rst), .Q(creg[255]) );
  IV U5139 ( .A(n5983), .Z(n3857) );
  IV U5140 ( .A(n5987), .Z(n3858) );
  IV U5141 ( .A(init), .Z(n3859) );
  IV U5142 ( .A(init), .Z(n3860) );
  IV U5143 ( .A(init), .Z(n3861) );
  IV U5144 ( .A(init), .Z(n3862) );
  IV U5145 ( .A(init), .Z(n3863) );
  IV U5146 ( .A(init), .Z(n3864) );
  IV U5147 ( .A(init), .Z(n3865) );
  IV U5148 ( .A(init), .Z(n3866) );
  IV U5149 ( .A(init), .Z(n3867) );
  IV U5150 ( .A(init), .Z(n3868) );
  IV U5151 ( .A(init), .Z(n3869) );
  IV U5152 ( .A(init), .Z(n3870) );
  IV U5153 ( .A(init), .Z(n3871) );
  IV U5154 ( .A(init), .Z(n3872) );
  IV U5155 ( .A(init), .Z(n3873) );
  IV U5156 ( .A(init), .Z(n3874) );
  IV U5157 ( .A(init), .Z(n3875) );
  IV U5158 ( .A(init), .Z(n3876) );
  IV U5159 ( .A(init), .Z(n3877) );
  IV U5160 ( .A(init), .Z(n3878) );
  IV U5161 ( .A(init), .Z(n3879) );
  IV U5162 ( .A(init), .Z(n3880) );
  IV U5163 ( .A(init), .Z(n3881) );
  IV U5164 ( .A(init), .Z(n3882) );
  IV U5165 ( .A(init), .Z(n3883) );
  IV U5166 ( .A(init), .Z(n3884) );
  IV U5167 ( .A(init), .Z(n3885) );
  IV U5168 ( .A(init), .Z(n3886) );
  IV U5169 ( .A(init), .Z(n3887) );
  IV U5170 ( .A(init), .Z(n3888) );
  IV U5171 ( .A(init), .Z(n3889) );
  IV U5172 ( .A(init), .Z(n3890) );
  IV U5173 ( .A(init), .Z(n3891) );
  IV U5174 ( .A(init), .Z(n3892) );
  IV U5175 ( .A(init), .Z(n3893) );
  IV U5176 ( .A(init), .Z(n3894) );
  IV U5177 ( .A(init), .Z(n3895) );
  IV U5178 ( .A(init), .Z(n3896) );
  IV U5179 ( .A(init), .Z(n3897) );
  IV U5180 ( .A(init), .Z(n3898) );
  IV U5181 ( .A(init), .Z(n3899) );
  IV U5182 ( .A(init), .Z(n3900) );
  IV U5183 ( .A(init), .Z(n3901) );
  IV U5184 ( .A(init), .Z(n3902) );
  IV U5185 ( .A(init), .Z(n3903) );
  IV U5186 ( .A(init), .Z(n3904) );
  IV U5187 ( .A(init), .Z(n3905) );
  IV U5188 ( .A(init), .Z(n3906) );
  IV U5189 ( .A(init), .Z(n3907) );
  IV U5190 ( .A(init), .Z(n3908) );
  IV U5191 ( .A(init), .Z(n3909) );
  IV U5192 ( .A(init), .Z(n3910) );
  IV U5193 ( .A(init), .Z(n3911) );
  IV U5194 ( .A(init), .Z(n3912) );
  IV U5195 ( .A(init), .Z(n3913) );
  IV U5196 ( .A(init), .Z(n3914) );
  IV U5197 ( .A(init), .Z(n3915) );
  IV U5198 ( .A(init), .Z(n3916) );
  IV U5199 ( .A(init), .Z(n3917) );
  IV U5200 ( .A(init), .Z(n3918) );
  IV U5201 ( .A(init), .Z(n3919) );
  IV U5202 ( .A(init), .Z(n3920) );
  IV U5203 ( .A(init), .Z(n3921) );
  IV U5204 ( .A(init), .Z(n3922) );
  IV U5205 ( .A(init), .Z(n3923) );
  IV U5206 ( .A(init), .Z(n3924) );
  IV U5207 ( .A(init), .Z(n3925) );
  IV U5208 ( .A(init), .Z(n3926) );
  IV U5209 ( .A(init), .Z(n3927) );
  IV U5210 ( .A(init), .Z(n3928) );
  IV U5211 ( .A(init), .Z(n3929) );
  IV U5212 ( .A(init), .Z(n3930) );
  IV U5213 ( .A(init), .Z(n3931) );
  IV U5214 ( .A(init), .Z(n3932) );
  ANDN U5215 ( .B(e[255]), .A(init), .Z(n5992) );
  NAND U5216 ( .A(init), .B(ereg[255]), .Z(n3933) );
  NANDN U5217 ( .A(n5992), .B(n3933), .Z(n5987) );
  NAND U5218 ( .A(n3858), .B(creg[0]), .Z(n3935) );
  NAND U5219 ( .A(n5987), .B(o[0]), .Z(n3934) );
  NAND U5220 ( .A(n3935), .B(n3934), .Z(c[0]) );
  NAND U5221 ( .A(n3858), .B(creg[100]), .Z(n3937) );
  NAND U5222 ( .A(n5987), .B(o[100]), .Z(n3936) );
  NAND U5223 ( .A(n3937), .B(n3936), .Z(c[100]) );
  NAND U5224 ( .A(n3858), .B(creg[101]), .Z(n3939) );
  NAND U5225 ( .A(n5987), .B(o[101]), .Z(n3938) );
  NAND U5226 ( .A(n3939), .B(n3938), .Z(c[101]) );
  NAND U5227 ( .A(n3858), .B(creg[102]), .Z(n3941) );
  NAND U5228 ( .A(n5987), .B(o[102]), .Z(n3940) );
  NAND U5229 ( .A(n3941), .B(n3940), .Z(c[102]) );
  NAND U5230 ( .A(n3858), .B(creg[103]), .Z(n3943) );
  NAND U5231 ( .A(n5987), .B(o[103]), .Z(n3942) );
  NAND U5232 ( .A(n3943), .B(n3942), .Z(c[103]) );
  NAND U5233 ( .A(n3858), .B(creg[104]), .Z(n3945) );
  NAND U5234 ( .A(n5987), .B(o[104]), .Z(n3944) );
  NAND U5235 ( .A(n3945), .B(n3944), .Z(c[104]) );
  NAND U5236 ( .A(n3858), .B(creg[105]), .Z(n3947) );
  NAND U5237 ( .A(n5987), .B(o[105]), .Z(n3946) );
  NAND U5238 ( .A(n3947), .B(n3946), .Z(c[105]) );
  NAND U5239 ( .A(n3858), .B(creg[106]), .Z(n3949) );
  NAND U5240 ( .A(n5987), .B(o[106]), .Z(n3948) );
  NAND U5241 ( .A(n3949), .B(n3948), .Z(c[106]) );
  NAND U5242 ( .A(n3858), .B(creg[107]), .Z(n3951) );
  NAND U5243 ( .A(n5987), .B(o[107]), .Z(n3950) );
  NAND U5244 ( .A(n3951), .B(n3950), .Z(c[107]) );
  NAND U5245 ( .A(n3858), .B(creg[108]), .Z(n3953) );
  NAND U5246 ( .A(n5987), .B(o[108]), .Z(n3952) );
  NAND U5247 ( .A(n3953), .B(n3952), .Z(c[108]) );
  NAND U5248 ( .A(n3858), .B(creg[109]), .Z(n3955) );
  NAND U5249 ( .A(n5987), .B(o[109]), .Z(n3954) );
  NAND U5250 ( .A(n3955), .B(n3954), .Z(c[109]) );
  NAND U5251 ( .A(n3858), .B(creg[10]), .Z(n3957) );
  NAND U5252 ( .A(n5987), .B(o[10]), .Z(n3956) );
  NAND U5253 ( .A(n3957), .B(n3956), .Z(c[10]) );
  NAND U5254 ( .A(n3858), .B(creg[110]), .Z(n3959) );
  NAND U5255 ( .A(n5987), .B(o[110]), .Z(n3958) );
  NAND U5256 ( .A(n3959), .B(n3958), .Z(c[110]) );
  NAND U5257 ( .A(n3858), .B(creg[111]), .Z(n3961) );
  NAND U5258 ( .A(n5987), .B(o[111]), .Z(n3960) );
  NAND U5259 ( .A(n3961), .B(n3960), .Z(c[111]) );
  NAND U5260 ( .A(n3858), .B(creg[112]), .Z(n3963) );
  NAND U5261 ( .A(n5987), .B(o[112]), .Z(n3962) );
  NAND U5262 ( .A(n3963), .B(n3962), .Z(c[112]) );
  NAND U5263 ( .A(n3858), .B(creg[113]), .Z(n3965) );
  NAND U5264 ( .A(n5987), .B(o[113]), .Z(n3964) );
  NAND U5265 ( .A(n3965), .B(n3964), .Z(c[113]) );
  NAND U5266 ( .A(n3858), .B(creg[114]), .Z(n3967) );
  NAND U5267 ( .A(n5987), .B(o[114]), .Z(n3966) );
  NAND U5268 ( .A(n3967), .B(n3966), .Z(c[114]) );
  NAND U5269 ( .A(n3858), .B(creg[115]), .Z(n3969) );
  NAND U5270 ( .A(n5987), .B(o[115]), .Z(n3968) );
  NAND U5271 ( .A(n3969), .B(n3968), .Z(c[115]) );
  NAND U5272 ( .A(n3858), .B(creg[116]), .Z(n3971) );
  NAND U5273 ( .A(n5987), .B(o[116]), .Z(n3970) );
  NAND U5274 ( .A(n3971), .B(n3970), .Z(c[116]) );
  NAND U5275 ( .A(n3858), .B(creg[117]), .Z(n3973) );
  NAND U5276 ( .A(n5987), .B(o[117]), .Z(n3972) );
  NAND U5277 ( .A(n3973), .B(n3972), .Z(c[117]) );
  NAND U5278 ( .A(n3858), .B(creg[118]), .Z(n3975) );
  NAND U5279 ( .A(n5987), .B(o[118]), .Z(n3974) );
  NAND U5280 ( .A(n3975), .B(n3974), .Z(c[118]) );
  NAND U5281 ( .A(n3858), .B(creg[119]), .Z(n3977) );
  NAND U5282 ( .A(n5987), .B(o[119]), .Z(n3976) );
  NAND U5283 ( .A(n3977), .B(n3976), .Z(c[119]) );
  NAND U5284 ( .A(n3858), .B(creg[11]), .Z(n3979) );
  NAND U5285 ( .A(n5987), .B(o[11]), .Z(n3978) );
  NAND U5286 ( .A(n3979), .B(n3978), .Z(c[11]) );
  NAND U5287 ( .A(n3858), .B(creg[120]), .Z(n3981) );
  NAND U5288 ( .A(n5987), .B(o[120]), .Z(n3980) );
  NAND U5289 ( .A(n3981), .B(n3980), .Z(c[120]) );
  NAND U5290 ( .A(n3858), .B(creg[121]), .Z(n3983) );
  NAND U5291 ( .A(n5987), .B(o[121]), .Z(n3982) );
  NAND U5292 ( .A(n3983), .B(n3982), .Z(c[121]) );
  NAND U5293 ( .A(n3858), .B(creg[122]), .Z(n3985) );
  NAND U5294 ( .A(n5987), .B(o[122]), .Z(n3984) );
  NAND U5295 ( .A(n3985), .B(n3984), .Z(c[122]) );
  NAND U5296 ( .A(n3858), .B(creg[123]), .Z(n3987) );
  NAND U5297 ( .A(n5987), .B(o[123]), .Z(n3986) );
  NAND U5298 ( .A(n3987), .B(n3986), .Z(c[123]) );
  NAND U5299 ( .A(n3858), .B(creg[124]), .Z(n3989) );
  NAND U5300 ( .A(n5987), .B(o[124]), .Z(n3988) );
  NAND U5301 ( .A(n3989), .B(n3988), .Z(c[124]) );
  NAND U5302 ( .A(n3858), .B(creg[125]), .Z(n3991) );
  NAND U5303 ( .A(n5987), .B(o[125]), .Z(n3990) );
  NAND U5304 ( .A(n3991), .B(n3990), .Z(c[125]) );
  NAND U5305 ( .A(n3858), .B(creg[126]), .Z(n3993) );
  NAND U5306 ( .A(n5987), .B(o[126]), .Z(n3992) );
  NAND U5307 ( .A(n3993), .B(n3992), .Z(c[126]) );
  NAND U5308 ( .A(n3858), .B(creg[127]), .Z(n3995) );
  NAND U5309 ( .A(n5987), .B(o[127]), .Z(n3994) );
  NAND U5310 ( .A(n3995), .B(n3994), .Z(c[127]) );
  NAND U5311 ( .A(n3858), .B(creg[128]), .Z(n3997) );
  NAND U5312 ( .A(n5987), .B(o[128]), .Z(n3996) );
  NAND U5313 ( .A(n3997), .B(n3996), .Z(c[128]) );
  NAND U5314 ( .A(n3858), .B(creg[129]), .Z(n3999) );
  NAND U5315 ( .A(n5987), .B(o[129]), .Z(n3998) );
  NAND U5316 ( .A(n3999), .B(n3998), .Z(c[129]) );
  NAND U5317 ( .A(n3858), .B(creg[12]), .Z(n4001) );
  NAND U5318 ( .A(n5987), .B(o[12]), .Z(n4000) );
  NAND U5319 ( .A(n4001), .B(n4000), .Z(c[12]) );
  NAND U5320 ( .A(n3858), .B(creg[130]), .Z(n4003) );
  NAND U5321 ( .A(n5987), .B(o[130]), .Z(n4002) );
  NAND U5322 ( .A(n4003), .B(n4002), .Z(c[130]) );
  NAND U5323 ( .A(n3858), .B(creg[131]), .Z(n4005) );
  NAND U5324 ( .A(n5987), .B(o[131]), .Z(n4004) );
  NAND U5325 ( .A(n4005), .B(n4004), .Z(c[131]) );
  NAND U5326 ( .A(n3858), .B(creg[132]), .Z(n4007) );
  NAND U5327 ( .A(n5987), .B(o[132]), .Z(n4006) );
  NAND U5328 ( .A(n4007), .B(n4006), .Z(c[132]) );
  NAND U5329 ( .A(n3858), .B(creg[133]), .Z(n4009) );
  NAND U5330 ( .A(n5987), .B(o[133]), .Z(n4008) );
  NAND U5331 ( .A(n4009), .B(n4008), .Z(c[133]) );
  NAND U5332 ( .A(n3858), .B(creg[134]), .Z(n4011) );
  NAND U5333 ( .A(n5987), .B(o[134]), .Z(n4010) );
  NAND U5334 ( .A(n4011), .B(n4010), .Z(c[134]) );
  NAND U5335 ( .A(n3858), .B(creg[135]), .Z(n4013) );
  NAND U5336 ( .A(n5987), .B(o[135]), .Z(n4012) );
  NAND U5337 ( .A(n4013), .B(n4012), .Z(c[135]) );
  NAND U5338 ( .A(n3858), .B(creg[136]), .Z(n4015) );
  NAND U5339 ( .A(n5987), .B(o[136]), .Z(n4014) );
  NAND U5340 ( .A(n4015), .B(n4014), .Z(c[136]) );
  NAND U5341 ( .A(n3858), .B(creg[137]), .Z(n4017) );
  NAND U5342 ( .A(n5987), .B(o[137]), .Z(n4016) );
  NAND U5343 ( .A(n4017), .B(n4016), .Z(c[137]) );
  NAND U5344 ( .A(n3858), .B(creg[138]), .Z(n4019) );
  NAND U5345 ( .A(n5987), .B(o[138]), .Z(n4018) );
  NAND U5346 ( .A(n4019), .B(n4018), .Z(c[138]) );
  NAND U5347 ( .A(n3858), .B(creg[139]), .Z(n4021) );
  NAND U5348 ( .A(n5987), .B(o[139]), .Z(n4020) );
  NAND U5349 ( .A(n4021), .B(n4020), .Z(c[139]) );
  NAND U5350 ( .A(n3858), .B(creg[13]), .Z(n4023) );
  NAND U5351 ( .A(n5987), .B(o[13]), .Z(n4022) );
  NAND U5352 ( .A(n4023), .B(n4022), .Z(c[13]) );
  NAND U5353 ( .A(n3858), .B(creg[140]), .Z(n4025) );
  NAND U5354 ( .A(n5987), .B(o[140]), .Z(n4024) );
  NAND U5355 ( .A(n4025), .B(n4024), .Z(c[140]) );
  NAND U5356 ( .A(n3858), .B(creg[141]), .Z(n4027) );
  NAND U5357 ( .A(n5987), .B(o[141]), .Z(n4026) );
  NAND U5358 ( .A(n4027), .B(n4026), .Z(c[141]) );
  NAND U5359 ( .A(n3858), .B(creg[142]), .Z(n4029) );
  NAND U5360 ( .A(n5987), .B(o[142]), .Z(n4028) );
  NAND U5361 ( .A(n4029), .B(n4028), .Z(c[142]) );
  NAND U5362 ( .A(n3858), .B(creg[143]), .Z(n4031) );
  NAND U5363 ( .A(n5987), .B(o[143]), .Z(n4030) );
  NAND U5364 ( .A(n4031), .B(n4030), .Z(c[143]) );
  NAND U5365 ( .A(n3858), .B(creg[144]), .Z(n4033) );
  NAND U5366 ( .A(n5987), .B(o[144]), .Z(n4032) );
  NAND U5367 ( .A(n4033), .B(n4032), .Z(c[144]) );
  NAND U5368 ( .A(n3858), .B(creg[145]), .Z(n4035) );
  NAND U5369 ( .A(n5987), .B(o[145]), .Z(n4034) );
  NAND U5370 ( .A(n4035), .B(n4034), .Z(c[145]) );
  NAND U5371 ( .A(n3858), .B(creg[146]), .Z(n4037) );
  NAND U5372 ( .A(n5987), .B(o[146]), .Z(n4036) );
  NAND U5373 ( .A(n4037), .B(n4036), .Z(c[146]) );
  NAND U5374 ( .A(n3858), .B(creg[147]), .Z(n4039) );
  NAND U5375 ( .A(n5987), .B(o[147]), .Z(n4038) );
  NAND U5376 ( .A(n4039), .B(n4038), .Z(c[147]) );
  NAND U5377 ( .A(n3858), .B(creg[148]), .Z(n4041) );
  NAND U5378 ( .A(n5987), .B(o[148]), .Z(n4040) );
  NAND U5379 ( .A(n4041), .B(n4040), .Z(c[148]) );
  NAND U5380 ( .A(n3858), .B(creg[149]), .Z(n4043) );
  NAND U5381 ( .A(n5987), .B(o[149]), .Z(n4042) );
  NAND U5382 ( .A(n4043), .B(n4042), .Z(c[149]) );
  NAND U5383 ( .A(n3858), .B(creg[14]), .Z(n4045) );
  NAND U5384 ( .A(n5987), .B(o[14]), .Z(n4044) );
  NAND U5385 ( .A(n4045), .B(n4044), .Z(c[14]) );
  NAND U5386 ( .A(n3858), .B(creg[150]), .Z(n4047) );
  NAND U5387 ( .A(n5987), .B(o[150]), .Z(n4046) );
  NAND U5388 ( .A(n4047), .B(n4046), .Z(c[150]) );
  NAND U5389 ( .A(n3858), .B(creg[151]), .Z(n4049) );
  NAND U5390 ( .A(n5987), .B(o[151]), .Z(n4048) );
  NAND U5391 ( .A(n4049), .B(n4048), .Z(c[151]) );
  NAND U5392 ( .A(n3858), .B(creg[152]), .Z(n4051) );
  NAND U5393 ( .A(n5987), .B(o[152]), .Z(n4050) );
  NAND U5394 ( .A(n4051), .B(n4050), .Z(c[152]) );
  NAND U5395 ( .A(n3858), .B(creg[153]), .Z(n4053) );
  NAND U5396 ( .A(n5987), .B(o[153]), .Z(n4052) );
  NAND U5397 ( .A(n4053), .B(n4052), .Z(c[153]) );
  NAND U5398 ( .A(n3858), .B(creg[154]), .Z(n4055) );
  NAND U5399 ( .A(n5987), .B(o[154]), .Z(n4054) );
  NAND U5400 ( .A(n4055), .B(n4054), .Z(c[154]) );
  NAND U5401 ( .A(n3858), .B(creg[155]), .Z(n4057) );
  NAND U5402 ( .A(n5987), .B(o[155]), .Z(n4056) );
  NAND U5403 ( .A(n4057), .B(n4056), .Z(c[155]) );
  NAND U5404 ( .A(n3858), .B(creg[156]), .Z(n4059) );
  NAND U5405 ( .A(n5987), .B(o[156]), .Z(n4058) );
  NAND U5406 ( .A(n4059), .B(n4058), .Z(c[156]) );
  NAND U5407 ( .A(n3858), .B(creg[157]), .Z(n4061) );
  NAND U5408 ( .A(n5987), .B(o[157]), .Z(n4060) );
  NAND U5409 ( .A(n4061), .B(n4060), .Z(c[157]) );
  NAND U5410 ( .A(n3858), .B(creg[158]), .Z(n4063) );
  NAND U5411 ( .A(n5987), .B(o[158]), .Z(n4062) );
  NAND U5412 ( .A(n4063), .B(n4062), .Z(c[158]) );
  NAND U5413 ( .A(n3858), .B(creg[159]), .Z(n4065) );
  NAND U5414 ( .A(n5987), .B(o[159]), .Z(n4064) );
  NAND U5415 ( .A(n4065), .B(n4064), .Z(c[159]) );
  NAND U5416 ( .A(n3858), .B(creg[15]), .Z(n4067) );
  NAND U5417 ( .A(n5987), .B(o[15]), .Z(n4066) );
  NAND U5418 ( .A(n4067), .B(n4066), .Z(c[15]) );
  NAND U5419 ( .A(n3858), .B(creg[160]), .Z(n4069) );
  NAND U5420 ( .A(n5987), .B(o[160]), .Z(n4068) );
  NAND U5421 ( .A(n4069), .B(n4068), .Z(c[160]) );
  NAND U5422 ( .A(n3858), .B(creg[161]), .Z(n4071) );
  NAND U5423 ( .A(n5987), .B(o[161]), .Z(n4070) );
  NAND U5424 ( .A(n4071), .B(n4070), .Z(c[161]) );
  NAND U5425 ( .A(n3858), .B(creg[162]), .Z(n4073) );
  NAND U5426 ( .A(n5987), .B(o[162]), .Z(n4072) );
  NAND U5427 ( .A(n4073), .B(n4072), .Z(c[162]) );
  NAND U5428 ( .A(n3858), .B(creg[163]), .Z(n4075) );
  NAND U5429 ( .A(n5987), .B(o[163]), .Z(n4074) );
  NAND U5430 ( .A(n4075), .B(n4074), .Z(c[163]) );
  NAND U5431 ( .A(n3858), .B(creg[164]), .Z(n4077) );
  NAND U5432 ( .A(n5987), .B(o[164]), .Z(n4076) );
  NAND U5433 ( .A(n4077), .B(n4076), .Z(c[164]) );
  NAND U5434 ( .A(n3858), .B(creg[165]), .Z(n4079) );
  NAND U5435 ( .A(n5987), .B(o[165]), .Z(n4078) );
  NAND U5436 ( .A(n4079), .B(n4078), .Z(c[165]) );
  NAND U5437 ( .A(n3858), .B(creg[166]), .Z(n4081) );
  NAND U5438 ( .A(n5987), .B(o[166]), .Z(n4080) );
  NAND U5439 ( .A(n4081), .B(n4080), .Z(c[166]) );
  NAND U5440 ( .A(n3858), .B(creg[167]), .Z(n4083) );
  NAND U5441 ( .A(n5987), .B(o[167]), .Z(n4082) );
  NAND U5442 ( .A(n4083), .B(n4082), .Z(c[167]) );
  NAND U5443 ( .A(n3858), .B(creg[168]), .Z(n4085) );
  NAND U5444 ( .A(n5987), .B(o[168]), .Z(n4084) );
  NAND U5445 ( .A(n4085), .B(n4084), .Z(c[168]) );
  NAND U5446 ( .A(n3858), .B(creg[169]), .Z(n4087) );
  NAND U5447 ( .A(n5987), .B(o[169]), .Z(n4086) );
  NAND U5448 ( .A(n4087), .B(n4086), .Z(c[169]) );
  NAND U5449 ( .A(n3858), .B(creg[16]), .Z(n4089) );
  NAND U5450 ( .A(n5987), .B(o[16]), .Z(n4088) );
  NAND U5451 ( .A(n4089), .B(n4088), .Z(c[16]) );
  NAND U5452 ( .A(n3858), .B(creg[170]), .Z(n4091) );
  NAND U5453 ( .A(n5987), .B(o[170]), .Z(n4090) );
  NAND U5454 ( .A(n4091), .B(n4090), .Z(c[170]) );
  NAND U5455 ( .A(n3858), .B(creg[171]), .Z(n4093) );
  NAND U5456 ( .A(n5987), .B(o[171]), .Z(n4092) );
  NAND U5457 ( .A(n4093), .B(n4092), .Z(c[171]) );
  NAND U5458 ( .A(n3858), .B(creg[172]), .Z(n4095) );
  NAND U5459 ( .A(n5987), .B(o[172]), .Z(n4094) );
  NAND U5460 ( .A(n4095), .B(n4094), .Z(c[172]) );
  NAND U5461 ( .A(n3858), .B(creg[173]), .Z(n4097) );
  NAND U5462 ( .A(n5987), .B(o[173]), .Z(n4096) );
  NAND U5463 ( .A(n4097), .B(n4096), .Z(c[173]) );
  NAND U5464 ( .A(n3858), .B(creg[174]), .Z(n4099) );
  NAND U5465 ( .A(n5987), .B(o[174]), .Z(n4098) );
  NAND U5466 ( .A(n4099), .B(n4098), .Z(c[174]) );
  NAND U5467 ( .A(n3858), .B(creg[175]), .Z(n4101) );
  NAND U5468 ( .A(n5987), .B(o[175]), .Z(n4100) );
  NAND U5469 ( .A(n4101), .B(n4100), .Z(c[175]) );
  NAND U5470 ( .A(n3858), .B(creg[176]), .Z(n4103) );
  NAND U5471 ( .A(n5987), .B(o[176]), .Z(n4102) );
  NAND U5472 ( .A(n4103), .B(n4102), .Z(c[176]) );
  NAND U5473 ( .A(n3858), .B(creg[177]), .Z(n4105) );
  NAND U5474 ( .A(n5987), .B(o[177]), .Z(n4104) );
  NAND U5475 ( .A(n4105), .B(n4104), .Z(c[177]) );
  NAND U5476 ( .A(n3858), .B(creg[178]), .Z(n4107) );
  NAND U5477 ( .A(n5987), .B(o[178]), .Z(n4106) );
  NAND U5478 ( .A(n4107), .B(n4106), .Z(c[178]) );
  NAND U5479 ( .A(n3858), .B(creg[179]), .Z(n4109) );
  NAND U5480 ( .A(n5987), .B(o[179]), .Z(n4108) );
  NAND U5481 ( .A(n4109), .B(n4108), .Z(c[179]) );
  NAND U5482 ( .A(n3858), .B(creg[17]), .Z(n4111) );
  NAND U5483 ( .A(n5987), .B(o[17]), .Z(n4110) );
  NAND U5484 ( .A(n4111), .B(n4110), .Z(c[17]) );
  NAND U5485 ( .A(n3858), .B(creg[180]), .Z(n4113) );
  NAND U5486 ( .A(n5987), .B(o[180]), .Z(n4112) );
  NAND U5487 ( .A(n4113), .B(n4112), .Z(c[180]) );
  NAND U5488 ( .A(n3858), .B(creg[181]), .Z(n4115) );
  NAND U5489 ( .A(n5987), .B(o[181]), .Z(n4114) );
  NAND U5490 ( .A(n4115), .B(n4114), .Z(c[181]) );
  NAND U5491 ( .A(n3858), .B(creg[182]), .Z(n4117) );
  NAND U5492 ( .A(n5987), .B(o[182]), .Z(n4116) );
  NAND U5493 ( .A(n4117), .B(n4116), .Z(c[182]) );
  NAND U5494 ( .A(n3858), .B(creg[183]), .Z(n4119) );
  NAND U5495 ( .A(n5987), .B(o[183]), .Z(n4118) );
  NAND U5496 ( .A(n4119), .B(n4118), .Z(c[183]) );
  NAND U5497 ( .A(n3858), .B(creg[184]), .Z(n4121) );
  NAND U5498 ( .A(n5987), .B(o[184]), .Z(n4120) );
  NAND U5499 ( .A(n4121), .B(n4120), .Z(c[184]) );
  NAND U5500 ( .A(n3858), .B(creg[185]), .Z(n4123) );
  NAND U5501 ( .A(n5987), .B(o[185]), .Z(n4122) );
  NAND U5502 ( .A(n4123), .B(n4122), .Z(c[185]) );
  NAND U5503 ( .A(n3858), .B(creg[186]), .Z(n4125) );
  NAND U5504 ( .A(n5987), .B(o[186]), .Z(n4124) );
  NAND U5505 ( .A(n4125), .B(n4124), .Z(c[186]) );
  NAND U5506 ( .A(n3858), .B(creg[187]), .Z(n4127) );
  NAND U5507 ( .A(n5987), .B(o[187]), .Z(n4126) );
  NAND U5508 ( .A(n4127), .B(n4126), .Z(c[187]) );
  NAND U5509 ( .A(n3858), .B(creg[188]), .Z(n4129) );
  NAND U5510 ( .A(n5987), .B(o[188]), .Z(n4128) );
  NAND U5511 ( .A(n4129), .B(n4128), .Z(c[188]) );
  NAND U5512 ( .A(n3858), .B(creg[189]), .Z(n4131) );
  NAND U5513 ( .A(n5987), .B(o[189]), .Z(n4130) );
  NAND U5514 ( .A(n4131), .B(n4130), .Z(c[189]) );
  NAND U5515 ( .A(n3858), .B(creg[18]), .Z(n4133) );
  NAND U5516 ( .A(n5987), .B(o[18]), .Z(n4132) );
  NAND U5517 ( .A(n4133), .B(n4132), .Z(c[18]) );
  NAND U5518 ( .A(n3858), .B(creg[190]), .Z(n4135) );
  NAND U5519 ( .A(n5987), .B(o[190]), .Z(n4134) );
  NAND U5520 ( .A(n4135), .B(n4134), .Z(c[190]) );
  NAND U5521 ( .A(n3858), .B(creg[191]), .Z(n4137) );
  NAND U5522 ( .A(n5987), .B(o[191]), .Z(n4136) );
  NAND U5523 ( .A(n4137), .B(n4136), .Z(c[191]) );
  NAND U5524 ( .A(n3858), .B(creg[192]), .Z(n4139) );
  NAND U5525 ( .A(n5987), .B(o[192]), .Z(n4138) );
  NAND U5526 ( .A(n4139), .B(n4138), .Z(c[192]) );
  NAND U5527 ( .A(n3858), .B(creg[193]), .Z(n4141) );
  NAND U5528 ( .A(n5987), .B(o[193]), .Z(n4140) );
  NAND U5529 ( .A(n4141), .B(n4140), .Z(c[193]) );
  NAND U5530 ( .A(n3858), .B(creg[194]), .Z(n4143) );
  NAND U5531 ( .A(n5987), .B(o[194]), .Z(n4142) );
  NAND U5532 ( .A(n4143), .B(n4142), .Z(c[194]) );
  NAND U5533 ( .A(n3858), .B(creg[195]), .Z(n4145) );
  NAND U5534 ( .A(n5987), .B(o[195]), .Z(n4144) );
  NAND U5535 ( .A(n4145), .B(n4144), .Z(c[195]) );
  NAND U5536 ( .A(n3858), .B(creg[196]), .Z(n4147) );
  NAND U5537 ( .A(n5987), .B(o[196]), .Z(n4146) );
  NAND U5538 ( .A(n4147), .B(n4146), .Z(c[196]) );
  NAND U5539 ( .A(n3858), .B(creg[197]), .Z(n4149) );
  NAND U5540 ( .A(n5987), .B(o[197]), .Z(n4148) );
  NAND U5541 ( .A(n4149), .B(n4148), .Z(c[197]) );
  NAND U5542 ( .A(n3858), .B(creg[198]), .Z(n4151) );
  NAND U5543 ( .A(n5987), .B(o[198]), .Z(n4150) );
  NAND U5544 ( .A(n4151), .B(n4150), .Z(c[198]) );
  NAND U5545 ( .A(n3858), .B(creg[199]), .Z(n4153) );
  NAND U5546 ( .A(n5987), .B(o[199]), .Z(n4152) );
  NAND U5547 ( .A(n4153), .B(n4152), .Z(c[199]) );
  NAND U5548 ( .A(n3858), .B(creg[19]), .Z(n4155) );
  NAND U5549 ( .A(n5987), .B(o[19]), .Z(n4154) );
  NAND U5550 ( .A(n4155), .B(n4154), .Z(c[19]) );
  NAND U5551 ( .A(n3858), .B(creg[1]), .Z(n4157) );
  NAND U5552 ( .A(n5987), .B(o[1]), .Z(n4156) );
  NAND U5553 ( .A(n4157), .B(n4156), .Z(c[1]) );
  NAND U5554 ( .A(n3858), .B(creg[200]), .Z(n4159) );
  NAND U5555 ( .A(n5987), .B(o[200]), .Z(n4158) );
  NAND U5556 ( .A(n4159), .B(n4158), .Z(c[200]) );
  NAND U5557 ( .A(n3858), .B(creg[201]), .Z(n4161) );
  NAND U5558 ( .A(n5987), .B(o[201]), .Z(n4160) );
  NAND U5559 ( .A(n4161), .B(n4160), .Z(c[201]) );
  NAND U5560 ( .A(n3858), .B(creg[202]), .Z(n4163) );
  NAND U5561 ( .A(n5987), .B(o[202]), .Z(n4162) );
  NAND U5562 ( .A(n4163), .B(n4162), .Z(c[202]) );
  NAND U5563 ( .A(n3858), .B(creg[203]), .Z(n4165) );
  NAND U5564 ( .A(n5987), .B(o[203]), .Z(n4164) );
  NAND U5565 ( .A(n4165), .B(n4164), .Z(c[203]) );
  NAND U5566 ( .A(n3858), .B(creg[204]), .Z(n4167) );
  NAND U5567 ( .A(n5987), .B(o[204]), .Z(n4166) );
  NAND U5568 ( .A(n4167), .B(n4166), .Z(c[204]) );
  NAND U5569 ( .A(n3858), .B(creg[205]), .Z(n4169) );
  NAND U5570 ( .A(n5987), .B(o[205]), .Z(n4168) );
  NAND U5571 ( .A(n4169), .B(n4168), .Z(c[205]) );
  NAND U5572 ( .A(n3858), .B(creg[206]), .Z(n4171) );
  NAND U5573 ( .A(n5987), .B(o[206]), .Z(n4170) );
  NAND U5574 ( .A(n4171), .B(n4170), .Z(c[206]) );
  NAND U5575 ( .A(n3858), .B(creg[207]), .Z(n4173) );
  NAND U5576 ( .A(n5987), .B(o[207]), .Z(n4172) );
  NAND U5577 ( .A(n4173), .B(n4172), .Z(c[207]) );
  NAND U5578 ( .A(n3858), .B(creg[208]), .Z(n4175) );
  NAND U5579 ( .A(n5987), .B(o[208]), .Z(n4174) );
  NAND U5580 ( .A(n4175), .B(n4174), .Z(c[208]) );
  NAND U5581 ( .A(n3858), .B(creg[209]), .Z(n4177) );
  NAND U5582 ( .A(n5987), .B(o[209]), .Z(n4176) );
  NAND U5583 ( .A(n4177), .B(n4176), .Z(c[209]) );
  NAND U5584 ( .A(n3858), .B(creg[20]), .Z(n4179) );
  NAND U5585 ( .A(n5987), .B(o[20]), .Z(n4178) );
  NAND U5586 ( .A(n4179), .B(n4178), .Z(c[20]) );
  NAND U5587 ( .A(n3858), .B(creg[210]), .Z(n4181) );
  NAND U5588 ( .A(n5987), .B(o[210]), .Z(n4180) );
  NAND U5589 ( .A(n4181), .B(n4180), .Z(c[210]) );
  NAND U5590 ( .A(n3858), .B(creg[211]), .Z(n4183) );
  NAND U5591 ( .A(n5987), .B(o[211]), .Z(n4182) );
  NAND U5592 ( .A(n4183), .B(n4182), .Z(c[211]) );
  NAND U5593 ( .A(n3858), .B(creg[212]), .Z(n4185) );
  NAND U5594 ( .A(n5987), .B(o[212]), .Z(n4184) );
  NAND U5595 ( .A(n4185), .B(n4184), .Z(c[212]) );
  NAND U5596 ( .A(n3858), .B(creg[213]), .Z(n4187) );
  NAND U5597 ( .A(n5987), .B(o[213]), .Z(n4186) );
  NAND U5598 ( .A(n4187), .B(n4186), .Z(c[213]) );
  NAND U5599 ( .A(n3858), .B(creg[214]), .Z(n4189) );
  NAND U5600 ( .A(n5987), .B(o[214]), .Z(n4188) );
  NAND U5601 ( .A(n4189), .B(n4188), .Z(c[214]) );
  NAND U5602 ( .A(n3858), .B(creg[215]), .Z(n4191) );
  NAND U5603 ( .A(n5987), .B(o[215]), .Z(n4190) );
  NAND U5604 ( .A(n4191), .B(n4190), .Z(c[215]) );
  NAND U5605 ( .A(n3858), .B(creg[216]), .Z(n4193) );
  NAND U5606 ( .A(n5987), .B(o[216]), .Z(n4192) );
  NAND U5607 ( .A(n4193), .B(n4192), .Z(c[216]) );
  NAND U5608 ( .A(n3858), .B(creg[217]), .Z(n4195) );
  NAND U5609 ( .A(n5987), .B(o[217]), .Z(n4194) );
  NAND U5610 ( .A(n4195), .B(n4194), .Z(c[217]) );
  NAND U5611 ( .A(n3858), .B(creg[218]), .Z(n4197) );
  NAND U5612 ( .A(n5987), .B(o[218]), .Z(n4196) );
  NAND U5613 ( .A(n4197), .B(n4196), .Z(c[218]) );
  NAND U5614 ( .A(n3858), .B(creg[219]), .Z(n4199) );
  NAND U5615 ( .A(n5987), .B(o[219]), .Z(n4198) );
  NAND U5616 ( .A(n4199), .B(n4198), .Z(c[219]) );
  NAND U5617 ( .A(n3858), .B(creg[21]), .Z(n4201) );
  NAND U5618 ( .A(n5987), .B(o[21]), .Z(n4200) );
  NAND U5619 ( .A(n4201), .B(n4200), .Z(c[21]) );
  NAND U5620 ( .A(n3858), .B(creg[220]), .Z(n4203) );
  NAND U5621 ( .A(n5987), .B(o[220]), .Z(n4202) );
  NAND U5622 ( .A(n4203), .B(n4202), .Z(c[220]) );
  NAND U5623 ( .A(n3858), .B(creg[221]), .Z(n4205) );
  NAND U5624 ( .A(n5987), .B(o[221]), .Z(n4204) );
  NAND U5625 ( .A(n4205), .B(n4204), .Z(c[221]) );
  NAND U5626 ( .A(n3858), .B(creg[222]), .Z(n4207) );
  NAND U5627 ( .A(n5987), .B(o[222]), .Z(n4206) );
  NAND U5628 ( .A(n4207), .B(n4206), .Z(c[222]) );
  NAND U5629 ( .A(n3858), .B(creg[223]), .Z(n4209) );
  NAND U5630 ( .A(n5987), .B(o[223]), .Z(n4208) );
  NAND U5631 ( .A(n4209), .B(n4208), .Z(c[223]) );
  NAND U5632 ( .A(n3858), .B(creg[224]), .Z(n4211) );
  NAND U5633 ( .A(n5987), .B(o[224]), .Z(n4210) );
  NAND U5634 ( .A(n4211), .B(n4210), .Z(c[224]) );
  NAND U5635 ( .A(n3858), .B(creg[225]), .Z(n4213) );
  NAND U5636 ( .A(n5987), .B(o[225]), .Z(n4212) );
  NAND U5637 ( .A(n4213), .B(n4212), .Z(c[225]) );
  NAND U5638 ( .A(n3858), .B(creg[226]), .Z(n4215) );
  NAND U5639 ( .A(n5987), .B(o[226]), .Z(n4214) );
  NAND U5640 ( .A(n4215), .B(n4214), .Z(c[226]) );
  NAND U5641 ( .A(n3858), .B(creg[227]), .Z(n4217) );
  NAND U5642 ( .A(n5987), .B(o[227]), .Z(n4216) );
  NAND U5643 ( .A(n4217), .B(n4216), .Z(c[227]) );
  NAND U5644 ( .A(n3858), .B(creg[228]), .Z(n4219) );
  NAND U5645 ( .A(n5987), .B(o[228]), .Z(n4218) );
  NAND U5646 ( .A(n4219), .B(n4218), .Z(c[228]) );
  NAND U5647 ( .A(n3858), .B(creg[229]), .Z(n4221) );
  NAND U5648 ( .A(n5987), .B(o[229]), .Z(n4220) );
  NAND U5649 ( .A(n4221), .B(n4220), .Z(c[229]) );
  NAND U5650 ( .A(n3858), .B(creg[22]), .Z(n4223) );
  NAND U5651 ( .A(n5987), .B(o[22]), .Z(n4222) );
  NAND U5652 ( .A(n4223), .B(n4222), .Z(c[22]) );
  NAND U5653 ( .A(n3858), .B(creg[230]), .Z(n4225) );
  NAND U5654 ( .A(n5987), .B(o[230]), .Z(n4224) );
  NAND U5655 ( .A(n4225), .B(n4224), .Z(c[230]) );
  NAND U5656 ( .A(n3858), .B(creg[231]), .Z(n4227) );
  NAND U5657 ( .A(n5987), .B(o[231]), .Z(n4226) );
  NAND U5658 ( .A(n4227), .B(n4226), .Z(c[231]) );
  NAND U5659 ( .A(n3858), .B(creg[232]), .Z(n4229) );
  NAND U5660 ( .A(n5987), .B(o[232]), .Z(n4228) );
  NAND U5661 ( .A(n4229), .B(n4228), .Z(c[232]) );
  NAND U5662 ( .A(n3858), .B(creg[233]), .Z(n4231) );
  NAND U5663 ( .A(n5987), .B(o[233]), .Z(n4230) );
  NAND U5664 ( .A(n4231), .B(n4230), .Z(c[233]) );
  NAND U5665 ( .A(n3858), .B(creg[234]), .Z(n4233) );
  NAND U5666 ( .A(n5987), .B(o[234]), .Z(n4232) );
  NAND U5667 ( .A(n4233), .B(n4232), .Z(c[234]) );
  NAND U5668 ( .A(n3858), .B(creg[235]), .Z(n4235) );
  NAND U5669 ( .A(n5987), .B(o[235]), .Z(n4234) );
  NAND U5670 ( .A(n4235), .B(n4234), .Z(c[235]) );
  NAND U5671 ( .A(n3858), .B(creg[236]), .Z(n4237) );
  NAND U5672 ( .A(n5987), .B(o[236]), .Z(n4236) );
  NAND U5673 ( .A(n4237), .B(n4236), .Z(c[236]) );
  NAND U5674 ( .A(n3858), .B(creg[237]), .Z(n4239) );
  NAND U5675 ( .A(n5987), .B(o[237]), .Z(n4238) );
  NAND U5676 ( .A(n4239), .B(n4238), .Z(c[237]) );
  NAND U5677 ( .A(n3858), .B(creg[238]), .Z(n4241) );
  NAND U5678 ( .A(n5987), .B(o[238]), .Z(n4240) );
  NAND U5679 ( .A(n4241), .B(n4240), .Z(c[238]) );
  NAND U5680 ( .A(n3858), .B(creg[239]), .Z(n4243) );
  NAND U5681 ( .A(n5987), .B(o[239]), .Z(n4242) );
  NAND U5682 ( .A(n4243), .B(n4242), .Z(c[239]) );
  NAND U5683 ( .A(n3858), .B(creg[23]), .Z(n4245) );
  NAND U5684 ( .A(n5987), .B(o[23]), .Z(n4244) );
  NAND U5685 ( .A(n4245), .B(n4244), .Z(c[23]) );
  NAND U5686 ( .A(n3858), .B(creg[240]), .Z(n4247) );
  NAND U5687 ( .A(n5987), .B(o[240]), .Z(n4246) );
  NAND U5688 ( .A(n4247), .B(n4246), .Z(c[240]) );
  NAND U5689 ( .A(n3858), .B(creg[241]), .Z(n4249) );
  NAND U5690 ( .A(n5987), .B(o[241]), .Z(n4248) );
  NAND U5691 ( .A(n4249), .B(n4248), .Z(c[241]) );
  NAND U5692 ( .A(n3858), .B(creg[242]), .Z(n4251) );
  NAND U5693 ( .A(n5987), .B(o[242]), .Z(n4250) );
  NAND U5694 ( .A(n4251), .B(n4250), .Z(c[242]) );
  NAND U5695 ( .A(n3858), .B(creg[243]), .Z(n4253) );
  NAND U5696 ( .A(n5987), .B(o[243]), .Z(n4252) );
  NAND U5697 ( .A(n4253), .B(n4252), .Z(c[243]) );
  NAND U5698 ( .A(n3858), .B(creg[244]), .Z(n4255) );
  NAND U5699 ( .A(n5987), .B(o[244]), .Z(n4254) );
  NAND U5700 ( .A(n4255), .B(n4254), .Z(c[244]) );
  NAND U5701 ( .A(n3858), .B(creg[245]), .Z(n4257) );
  NAND U5702 ( .A(n5987), .B(o[245]), .Z(n4256) );
  NAND U5703 ( .A(n4257), .B(n4256), .Z(c[245]) );
  NAND U5704 ( .A(n3858), .B(creg[246]), .Z(n4259) );
  NAND U5705 ( .A(n5987), .B(o[246]), .Z(n4258) );
  NAND U5706 ( .A(n4259), .B(n4258), .Z(c[246]) );
  NAND U5707 ( .A(n3858), .B(creg[247]), .Z(n4261) );
  NAND U5708 ( .A(n5987), .B(o[247]), .Z(n4260) );
  NAND U5709 ( .A(n4261), .B(n4260), .Z(c[247]) );
  NAND U5710 ( .A(n3858), .B(creg[248]), .Z(n4263) );
  NAND U5711 ( .A(n5987), .B(o[248]), .Z(n4262) );
  NAND U5712 ( .A(n4263), .B(n4262), .Z(c[248]) );
  NAND U5713 ( .A(n3858), .B(creg[249]), .Z(n4265) );
  NAND U5714 ( .A(n5987), .B(o[249]), .Z(n4264) );
  NAND U5715 ( .A(n4265), .B(n4264), .Z(c[249]) );
  NAND U5716 ( .A(n3858), .B(creg[24]), .Z(n4267) );
  NAND U5717 ( .A(n5987), .B(o[24]), .Z(n4266) );
  NAND U5718 ( .A(n4267), .B(n4266), .Z(c[24]) );
  NAND U5719 ( .A(n3858), .B(creg[250]), .Z(n4269) );
  NAND U5720 ( .A(n5987), .B(o[250]), .Z(n4268) );
  NAND U5721 ( .A(n4269), .B(n4268), .Z(c[250]) );
  NAND U5722 ( .A(n3858), .B(creg[251]), .Z(n4271) );
  NAND U5723 ( .A(n5987), .B(o[251]), .Z(n4270) );
  NAND U5724 ( .A(n4271), .B(n4270), .Z(c[251]) );
  NAND U5725 ( .A(n3858), .B(creg[252]), .Z(n4273) );
  NAND U5726 ( .A(n5987), .B(o[252]), .Z(n4272) );
  NAND U5727 ( .A(n4273), .B(n4272), .Z(c[252]) );
  NAND U5728 ( .A(n3858), .B(creg[253]), .Z(n4275) );
  NAND U5729 ( .A(n5987), .B(o[253]), .Z(n4274) );
  NAND U5730 ( .A(n4275), .B(n4274), .Z(c[253]) );
  NAND U5731 ( .A(n3858), .B(creg[254]), .Z(n4277) );
  NAND U5732 ( .A(n5987), .B(o[254]), .Z(n4276) );
  NAND U5733 ( .A(n4277), .B(n4276), .Z(c[254]) );
  NAND U5734 ( .A(n3858), .B(creg[255]), .Z(n4279) );
  NAND U5735 ( .A(n5987), .B(o[255]), .Z(n4278) );
  NAND U5736 ( .A(n4279), .B(n4278), .Z(c[255]) );
  NAND U5737 ( .A(n3858), .B(creg[25]), .Z(n4281) );
  NAND U5738 ( .A(n5987), .B(o[25]), .Z(n4280) );
  NAND U5739 ( .A(n4281), .B(n4280), .Z(c[25]) );
  NAND U5740 ( .A(n3858), .B(creg[26]), .Z(n4283) );
  NAND U5741 ( .A(n5987), .B(o[26]), .Z(n4282) );
  NAND U5742 ( .A(n4283), .B(n4282), .Z(c[26]) );
  NAND U5743 ( .A(n3858), .B(creg[27]), .Z(n4285) );
  NAND U5744 ( .A(n5987), .B(o[27]), .Z(n4284) );
  NAND U5745 ( .A(n4285), .B(n4284), .Z(c[27]) );
  NAND U5746 ( .A(n3858), .B(creg[28]), .Z(n4287) );
  NAND U5747 ( .A(n5987), .B(o[28]), .Z(n4286) );
  NAND U5748 ( .A(n4287), .B(n4286), .Z(c[28]) );
  NAND U5749 ( .A(n3858), .B(creg[29]), .Z(n4289) );
  NAND U5750 ( .A(n5987), .B(o[29]), .Z(n4288) );
  NAND U5751 ( .A(n4289), .B(n4288), .Z(c[29]) );
  NAND U5752 ( .A(n3858), .B(creg[2]), .Z(n4291) );
  NAND U5753 ( .A(n5987), .B(o[2]), .Z(n4290) );
  NAND U5754 ( .A(n4291), .B(n4290), .Z(c[2]) );
  NAND U5755 ( .A(n3858), .B(creg[30]), .Z(n4293) );
  NAND U5756 ( .A(n5987), .B(o[30]), .Z(n4292) );
  NAND U5757 ( .A(n4293), .B(n4292), .Z(c[30]) );
  NAND U5758 ( .A(n3858), .B(creg[31]), .Z(n4295) );
  NAND U5759 ( .A(n5987), .B(o[31]), .Z(n4294) );
  NAND U5760 ( .A(n4295), .B(n4294), .Z(c[31]) );
  NAND U5761 ( .A(n3858), .B(creg[32]), .Z(n4297) );
  NAND U5762 ( .A(n5987), .B(o[32]), .Z(n4296) );
  NAND U5763 ( .A(n4297), .B(n4296), .Z(c[32]) );
  NAND U5764 ( .A(n3858), .B(creg[33]), .Z(n4299) );
  NAND U5765 ( .A(n5987), .B(o[33]), .Z(n4298) );
  NAND U5766 ( .A(n4299), .B(n4298), .Z(c[33]) );
  NAND U5767 ( .A(n3858), .B(creg[34]), .Z(n4301) );
  NAND U5768 ( .A(n5987), .B(o[34]), .Z(n4300) );
  NAND U5769 ( .A(n4301), .B(n4300), .Z(c[34]) );
  NAND U5770 ( .A(n3858), .B(creg[35]), .Z(n4303) );
  NAND U5771 ( .A(n5987), .B(o[35]), .Z(n4302) );
  NAND U5772 ( .A(n4303), .B(n4302), .Z(c[35]) );
  NAND U5773 ( .A(n3858), .B(creg[36]), .Z(n4305) );
  NAND U5774 ( .A(n5987), .B(o[36]), .Z(n4304) );
  NAND U5775 ( .A(n4305), .B(n4304), .Z(c[36]) );
  NAND U5776 ( .A(n3858), .B(creg[37]), .Z(n4307) );
  NAND U5777 ( .A(n5987), .B(o[37]), .Z(n4306) );
  NAND U5778 ( .A(n4307), .B(n4306), .Z(c[37]) );
  NAND U5779 ( .A(n3858), .B(creg[38]), .Z(n4309) );
  NAND U5780 ( .A(n5987), .B(o[38]), .Z(n4308) );
  NAND U5781 ( .A(n4309), .B(n4308), .Z(c[38]) );
  NAND U5782 ( .A(n3858), .B(creg[39]), .Z(n4311) );
  NAND U5783 ( .A(n5987), .B(o[39]), .Z(n4310) );
  NAND U5784 ( .A(n4311), .B(n4310), .Z(c[39]) );
  NAND U5785 ( .A(n3858), .B(creg[3]), .Z(n4313) );
  NAND U5786 ( .A(n5987), .B(o[3]), .Z(n4312) );
  NAND U5787 ( .A(n4313), .B(n4312), .Z(c[3]) );
  NAND U5788 ( .A(n3858), .B(creg[40]), .Z(n4315) );
  NAND U5789 ( .A(n5987), .B(o[40]), .Z(n4314) );
  NAND U5790 ( .A(n4315), .B(n4314), .Z(c[40]) );
  NAND U5791 ( .A(n3858), .B(creg[41]), .Z(n4317) );
  NAND U5792 ( .A(n5987), .B(o[41]), .Z(n4316) );
  NAND U5793 ( .A(n4317), .B(n4316), .Z(c[41]) );
  NAND U5794 ( .A(n3858), .B(creg[42]), .Z(n4319) );
  NAND U5795 ( .A(n5987), .B(o[42]), .Z(n4318) );
  NAND U5796 ( .A(n4319), .B(n4318), .Z(c[42]) );
  NAND U5797 ( .A(n3858), .B(creg[43]), .Z(n4321) );
  NAND U5798 ( .A(n5987), .B(o[43]), .Z(n4320) );
  NAND U5799 ( .A(n4321), .B(n4320), .Z(c[43]) );
  NAND U5800 ( .A(n3858), .B(creg[44]), .Z(n4323) );
  NAND U5801 ( .A(n5987), .B(o[44]), .Z(n4322) );
  NAND U5802 ( .A(n4323), .B(n4322), .Z(c[44]) );
  NAND U5803 ( .A(n3858), .B(creg[45]), .Z(n4325) );
  NAND U5804 ( .A(n5987), .B(o[45]), .Z(n4324) );
  NAND U5805 ( .A(n4325), .B(n4324), .Z(c[45]) );
  NAND U5806 ( .A(n3858), .B(creg[46]), .Z(n4327) );
  NAND U5807 ( .A(n5987), .B(o[46]), .Z(n4326) );
  NAND U5808 ( .A(n4327), .B(n4326), .Z(c[46]) );
  NAND U5809 ( .A(n3858), .B(creg[47]), .Z(n4329) );
  NAND U5810 ( .A(n5987), .B(o[47]), .Z(n4328) );
  NAND U5811 ( .A(n4329), .B(n4328), .Z(c[47]) );
  NAND U5812 ( .A(n3858), .B(creg[48]), .Z(n4331) );
  NAND U5813 ( .A(n5987), .B(o[48]), .Z(n4330) );
  NAND U5814 ( .A(n4331), .B(n4330), .Z(c[48]) );
  NAND U5815 ( .A(n3858), .B(creg[49]), .Z(n4333) );
  NAND U5816 ( .A(n5987), .B(o[49]), .Z(n4332) );
  NAND U5817 ( .A(n4333), .B(n4332), .Z(c[49]) );
  NAND U5818 ( .A(n3858), .B(creg[4]), .Z(n4335) );
  NAND U5819 ( .A(n5987), .B(o[4]), .Z(n4334) );
  NAND U5820 ( .A(n4335), .B(n4334), .Z(c[4]) );
  NAND U5821 ( .A(n3858), .B(creg[50]), .Z(n4337) );
  NAND U5822 ( .A(n5987), .B(o[50]), .Z(n4336) );
  NAND U5823 ( .A(n4337), .B(n4336), .Z(c[50]) );
  NAND U5824 ( .A(n3858), .B(creg[51]), .Z(n4339) );
  NAND U5825 ( .A(n5987), .B(o[51]), .Z(n4338) );
  NAND U5826 ( .A(n4339), .B(n4338), .Z(c[51]) );
  NAND U5827 ( .A(n3858), .B(creg[52]), .Z(n4341) );
  NAND U5828 ( .A(n5987), .B(o[52]), .Z(n4340) );
  NAND U5829 ( .A(n4341), .B(n4340), .Z(c[52]) );
  NAND U5830 ( .A(n3858), .B(creg[53]), .Z(n4343) );
  NAND U5831 ( .A(n5987), .B(o[53]), .Z(n4342) );
  NAND U5832 ( .A(n4343), .B(n4342), .Z(c[53]) );
  NAND U5833 ( .A(n3858), .B(creg[54]), .Z(n4345) );
  NAND U5834 ( .A(n5987), .B(o[54]), .Z(n4344) );
  NAND U5835 ( .A(n4345), .B(n4344), .Z(c[54]) );
  NAND U5836 ( .A(n3858), .B(creg[55]), .Z(n4347) );
  NAND U5837 ( .A(n5987), .B(o[55]), .Z(n4346) );
  NAND U5838 ( .A(n4347), .B(n4346), .Z(c[55]) );
  NAND U5839 ( .A(n3858), .B(creg[56]), .Z(n4349) );
  NAND U5840 ( .A(n5987), .B(o[56]), .Z(n4348) );
  NAND U5841 ( .A(n4349), .B(n4348), .Z(c[56]) );
  NAND U5842 ( .A(n3858), .B(creg[57]), .Z(n4351) );
  NAND U5843 ( .A(n5987), .B(o[57]), .Z(n4350) );
  NAND U5844 ( .A(n4351), .B(n4350), .Z(c[57]) );
  NAND U5845 ( .A(n3858), .B(creg[58]), .Z(n4353) );
  NAND U5846 ( .A(n5987), .B(o[58]), .Z(n4352) );
  NAND U5847 ( .A(n4353), .B(n4352), .Z(c[58]) );
  NAND U5848 ( .A(n3858), .B(creg[59]), .Z(n4355) );
  NAND U5849 ( .A(n5987), .B(o[59]), .Z(n4354) );
  NAND U5850 ( .A(n4355), .B(n4354), .Z(c[59]) );
  NAND U5851 ( .A(n3858), .B(creg[5]), .Z(n4357) );
  NAND U5852 ( .A(n5987), .B(o[5]), .Z(n4356) );
  NAND U5853 ( .A(n4357), .B(n4356), .Z(c[5]) );
  NAND U5854 ( .A(n3858), .B(creg[60]), .Z(n4359) );
  NAND U5855 ( .A(n5987), .B(o[60]), .Z(n4358) );
  NAND U5856 ( .A(n4359), .B(n4358), .Z(c[60]) );
  NAND U5857 ( .A(n3858), .B(creg[61]), .Z(n4361) );
  NAND U5858 ( .A(n5987), .B(o[61]), .Z(n4360) );
  NAND U5859 ( .A(n4361), .B(n4360), .Z(c[61]) );
  NAND U5860 ( .A(n3858), .B(creg[62]), .Z(n4363) );
  NAND U5861 ( .A(n5987), .B(o[62]), .Z(n4362) );
  NAND U5862 ( .A(n4363), .B(n4362), .Z(c[62]) );
  NAND U5863 ( .A(n3858), .B(creg[63]), .Z(n4365) );
  NAND U5864 ( .A(n5987), .B(o[63]), .Z(n4364) );
  NAND U5865 ( .A(n4365), .B(n4364), .Z(c[63]) );
  NAND U5866 ( .A(n3858), .B(creg[64]), .Z(n4367) );
  NAND U5867 ( .A(n5987), .B(o[64]), .Z(n4366) );
  NAND U5868 ( .A(n4367), .B(n4366), .Z(c[64]) );
  NAND U5869 ( .A(n3858), .B(creg[65]), .Z(n4369) );
  NAND U5870 ( .A(n5987), .B(o[65]), .Z(n4368) );
  NAND U5871 ( .A(n4369), .B(n4368), .Z(c[65]) );
  NAND U5872 ( .A(n3858), .B(creg[66]), .Z(n4371) );
  NAND U5873 ( .A(n5987), .B(o[66]), .Z(n4370) );
  NAND U5874 ( .A(n4371), .B(n4370), .Z(c[66]) );
  NAND U5875 ( .A(n3858), .B(creg[67]), .Z(n4373) );
  NAND U5876 ( .A(n5987), .B(o[67]), .Z(n4372) );
  NAND U5877 ( .A(n4373), .B(n4372), .Z(c[67]) );
  NAND U5878 ( .A(n3858), .B(creg[68]), .Z(n4375) );
  NAND U5879 ( .A(n5987), .B(o[68]), .Z(n4374) );
  NAND U5880 ( .A(n4375), .B(n4374), .Z(c[68]) );
  NAND U5881 ( .A(n3858), .B(creg[69]), .Z(n4377) );
  NAND U5882 ( .A(n5987), .B(o[69]), .Z(n4376) );
  NAND U5883 ( .A(n4377), .B(n4376), .Z(c[69]) );
  NAND U5884 ( .A(n3858), .B(creg[6]), .Z(n4379) );
  NAND U5885 ( .A(n5987), .B(o[6]), .Z(n4378) );
  NAND U5886 ( .A(n4379), .B(n4378), .Z(c[6]) );
  NAND U5887 ( .A(n3858), .B(creg[70]), .Z(n4381) );
  NAND U5888 ( .A(n5987), .B(o[70]), .Z(n4380) );
  NAND U5889 ( .A(n4381), .B(n4380), .Z(c[70]) );
  NAND U5890 ( .A(n3858), .B(creg[71]), .Z(n4383) );
  NAND U5891 ( .A(n5987), .B(o[71]), .Z(n4382) );
  NAND U5892 ( .A(n4383), .B(n4382), .Z(c[71]) );
  NAND U5893 ( .A(n3858), .B(creg[72]), .Z(n4385) );
  NAND U5894 ( .A(n5987), .B(o[72]), .Z(n4384) );
  NAND U5895 ( .A(n4385), .B(n4384), .Z(c[72]) );
  NAND U5896 ( .A(n3858), .B(creg[73]), .Z(n4387) );
  NAND U5897 ( .A(n5987), .B(o[73]), .Z(n4386) );
  NAND U5898 ( .A(n4387), .B(n4386), .Z(c[73]) );
  NAND U5899 ( .A(n3858), .B(creg[74]), .Z(n4389) );
  NAND U5900 ( .A(n5987), .B(o[74]), .Z(n4388) );
  NAND U5901 ( .A(n4389), .B(n4388), .Z(c[74]) );
  NAND U5902 ( .A(n3858), .B(creg[75]), .Z(n4391) );
  NAND U5903 ( .A(n5987), .B(o[75]), .Z(n4390) );
  NAND U5904 ( .A(n4391), .B(n4390), .Z(c[75]) );
  NAND U5905 ( .A(n3858), .B(creg[76]), .Z(n4393) );
  NAND U5906 ( .A(n5987), .B(o[76]), .Z(n4392) );
  NAND U5907 ( .A(n4393), .B(n4392), .Z(c[76]) );
  NAND U5908 ( .A(n3858), .B(creg[77]), .Z(n4395) );
  NAND U5909 ( .A(n5987), .B(o[77]), .Z(n4394) );
  NAND U5910 ( .A(n4395), .B(n4394), .Z(c[77]) );
  NAND U5911 ( .A(n3858), .B(creg[78]), .Z(n4397) );
  NAND U5912 ( .A(n5987), .B(o[78]), .Z(n4396) );
  NAND U5913 ( .A(n4397), .B(n4396), .Z(c[78]) );
  NAND U5914 ( .A(n3858), .B(creg[79]), .Z(n4399) );
  NAND U5915 ( .A(n5987), .B(o[79]), .Z(n4398) );
  NAND U5916 ( .A(n4399), .B(n4398), .Z(c[79]) );
  NAND U5917 ( .A(n3858), .B(creg[7]), .Z(n4401) );
  NAND U5918 ( .A(n5987), .B(o[7]), .Z(n4400) );
  NAND U5919 ( .A(n4401), .B(n4400), .Z(c[7]) );
  NAND U5920 ( .A(n3858), .B(creg[80]), .Z(n4403) );
  NAND U5921 ( .A(n5987), .B(o[80]), .Z(n4402) );
  NAND U5922 ( .A(n4403), .B(n4402), .Z(c[80]) );
  NAND U5923 ( .A(n3858), .B(creg[81]), .Z(n4405) );
  NAND U5924 ( .A(n5987), .B(o[81]), .Z(n4404) );
  NAND U5925 ( .A(n4405), .B(n4404), .Z(c[81]) );
  NAND U5926 ( .A(n3858), .B(creg[82]), .Z(n4407) );
  NAND U5927 ( .A(n5987), .B(o[82]), .Z(n4406) );
  NAND U5928 ( .A(n4407), .B(n4406), .Z(c[82]) );
  NAND U5929 ( .A(n3858), .B(creg[83]), .Z(n4409) );
  NAND U5930 ( .A(n5987), .B(o[83]), .Z(n4408) );
  NAND U5931 ( .A(n4409), .B(n4408), .Z(c[83]) );
  NAND U5932 ( .A(n3858), .B(creg[84]), .Z(n4411) );
  NAND U5933 ( .A(n5987), .B(o[84]), .Z(n4410) );
  NAND U5934 ( .A(n4411), .B(n4410), .Z(c[84]) );
  NAND U5935 ( .A(n3858), .B(creg[85]), .Z(n4413) );
  NAND U5936 ( .A(n5987), .B(o[85]), .Z(n4412) );
  NAND U5937 ( .A(n4413), .B(n4412), .Z(c[85]) );
  NAND U5938 ( .A(n3858), .B(creg[86]), .Z(n4415) );
  NAND U5939 ( .A(n5987), .B(o[86]), .Z(n4414) );
  NAND U5940 ( .A(n4415), .B(n4414), .Z(c[86]) );
  NAND U5941 ( .A(n3858), .B(creg[87]), .Z(n4417) );
  NAND U5942 ( .A(n5987), .B(o[87]), .Z(n4416) );
  NAND U5943 ( .A(n4417), .B(n4416), .Z(c[87]) );
  NAND U5944 ( .A(n3858), .B(creg[88]), .Z(n4419) );
  NAND U5945 ( .A(n5987), .B(o[88]), .Z(n4418) );
  NAND U5946 ( .A(n4419), .B(n4418), .Z(c[88]) );
  NAND U5947 ( .A(n3858), .B(creg[89]), .Z(n4421) );
  NAND U5948 ( .A(n5987), .B(o[89]), .Z(n4420) );
  NAND U5949 ( .A(n4421), .B(n4420), .Z(c[89]) );
  NAND U5950 ( .A(n3858), .B(creg[8]), .Z(n4423) );
  NAND U5951 ( .A(n5987), .B(o[8]), .Z(n4422) );
  NAND U5952 ( .A(n4423), .B(n4422), .Z(c[8]) );
  NAND U5953 ( .A(n3858), .B(creg[90]), .Z(n4425) );
  NAND U5954 ( .A(n5987), .B(o[90]), .Z(n4424) );
  NAND U5955 ( .A(n4425), .B(n4424), .Z(c[90]) );
  NAND U5956 ( .A(n3858), .B(creg[91]), .Z(n4427) );
  NAND U5957 ( .A(n5987), .B(o[91]), .Z(n4426) );
  NAND U5958 ( .A(n4427), .B(n4426), .Z(c[91]) );
  NAND U5959 ( .A(n3858), .B(creg[92]), .Z(n4429) );
  NAND U5960 ( .A(n5987), .B(o[92]), .Z(n4428) );
  NAND U5961 ( .A(n4429), .B(n4428), .Z(c[92]) );
  NAND U5962 ( .A(n3858), .B(creg[93]), .Z(n4431) );
  NAND U5963 ( .A(n5987), .B(o[93]), .Z(n4430) );
  NAND U5964 ( .A(n4431), .B(n4430), .Z(c[93]) );
  NAND U5965 ( .A(n3858), .B(creg[94]), .Z(n4433) );
  NAND U5966 ( .A(n5987), .B(o[94]), .Z(n4432) );
  NAND U5967 ( .A(n4433), .B(n4432), .Z(c[94]) );
  NAND U5968 ( .A(n3858), .B(creg[95]), .Z(n4435) );
  NAND U5969 ( .A(n5987), .B(o[95]), .Z(n4434) );
  NAND U5970 ( .A(n4435), .B(n4434), .Z(c[95]) );
  NAND U5971 ( .A(n3858), .B(creg[96]), .Z(n4437) );
  NAND U5972 ( .A(n5987), .B(o[96]), .Z(n4436) );
  NAND U5973 ( .A(n4437), .B(n4436), .Z(c[96]) );
  NAND U5974 ( .A(n3858), .B(creg[97]), .Z(n4439) );
  NAND U5975 ( .A(n5987), .B(o[97]), .Z(n4438) );
  NAND U5976 ( .A(n4439), .B(n4438), .Z(c[97]) );
  NAND U5977 ( .A(n3858), .B(creg[98]), .Z(n4441) );
  NAND U5978 ( .A(n5987), .B(o[98]), .Z(n4440) );
  NAND U5979 ( .A(n4441), .B(n4440), .Z(c[98]) );
  NAND U5980 ( .A(n3858), .B(creg[99]), .Z(n4443) );
  NAND U5981 ( .A(n5987), .B(o[99]), .Z(n4442) );
  NAND U5982 ( .A(n4443), .B(n4442), .Z(c[99]) );
  NAND U5983 ( .A(n3858), .B(creg[9]), .Z(n4445) );
  NAND U5984 ( .A(n5987), .B(o[9]), .Z(n4444) );
  NAND U5985 ( .A(n4445), .B(n4444), .Z(c[9]) );
  NANDN U5986 ( .A(start_reg[0]), .B(init), .Z(start_in[0]) );
  AND U5987 ( .A(start_reg[100]), .B(init), .Z(start_in[100]) );
  AND U5988 ( .A(start_reg[101]), .B(init), .Z(start_in[101]) );
  AND U5989 ( .A(start_reg[102]), .B(init), .Z(start_in[102]) );
  AND U5990 ( .A(start_reg[103]), .B(init), .Z(start_in[103]) );
  AND U5991 ( .A(start_reg[104]), .B(init), .Z(start_in[104]) );
  AND U5992 ( .A(start_reg[105]), .B(init), .Z(start_in[105]) );
  AND U5993 ( .A(start_reg[106]), .B(init), .Z(start_in[106]) );
  AND U5994 ( .A(start_reg[107]), .B(init), .Z(start_in[107]) );
  AND U5995 ( .A(start_reg[108]), .B(init), .Z(start_in[108]) );
  AND U5996 ( .A(start_reg[109]), .B(init), .Z(start_in[109]) );
  AND U5997 ( .A(start_reg[10]), .B(init), .Z(start_in[10]) );
  AND U5998 ( .A(start_reg[110]), .B(init), .Z(start_in[110]) );
  AND U5999 ( .A(start_reg[111]), .B(init), .Z(start_in[111]) );
  AND U6000 ( .A(start_reg[112]), .B(init), .Z(start_in[112]) );
  AND U6001 ( .A(start_reg[113]), .B(init), .Z(start_in[113]) );
  AND U6002 ( .A(start_reg[114]), .B(init), .Z(start_in[114]) );
  AND U6003 ( .A(start_reg[115]), .B(init), .Z(start_in[115]) );
  AND U6004 ( .A(start_reg[116]), .B(init), .Z(start_in[116]) );
  AND U6005 ( .A(start_reg[117]), .B(init), .Z(start_in[117]) );
  AND U6006 ( .A(start_reg[118]), .B(init), .Z(start_in[118]) );
  AND U6007 ( .A(start_reg[119]), .B(init), .Z(start_in[119]) );
  AND U6008 ( .A(start_reg[11]), .B(init), .Z(start_in[11]) );
  AND U6009 ( .A(start_reg[120]), .B(init), .Z(start_in[120]) );
  AND U6010 ( .A(start_reg[121]), .B(init), .Z(start_in[121]) );
  AND U6011 ( .A(start_reg[122]), .B(init), .Z(start_in[122]) );
  AND U6012 ( .A(start_reg[123]), .B(init), .Z(start_in[123]) );
  AND U6013 ( .A(start_reg[124]), .B(init), .Z(start_in[124]) );
  AND U6014 ( .A(start_reg[125]), .B(init), .Z(start_in[125]) );
  AND U6015 ( .A(start_reg[126]), .B(init), .Z(start_in[126]) );
  AND U6016 ( .A(start_reg[127]), .B(init), .Z(start_in[127]) );
  AND U6017 ( .A(start_reg[128]), .B(init), .Z(start_in[128]) );
  AND U6018 ( .A(start_reg[129]), .B(init), .Z(start_in[129]) );
  AND U6019 ( .A(start_reg[12]), .B(init), .Z(start_in[12]) );
  AND U6020 ( .A(start_reg[130]), .B(init), .Z(start_in[130]) );
  AND U6021 ( .A(start_reg[131]), .B(init), .Z(start_in[131]) );
  AND U6022 ( .A(start_reg[132]), .B(init), .Z(start_in[132]) );
  AND U6023 ( .A(start_reg[133]), .B(init), .Z(start_in[133]) );
  AND U6024 ( .A(start_reg[134]), .B(init), .Z(start_in[134]) );
  AND U6025 ( .A(start_reg[135]), .B(init), .Z(start_in[135]) );
  AND U6026 ( .A(start_reg[136]), .B(init), .Z(start_in[136]) );
  AND U6027 ( .A(start_reg[137]), .B(init), .Z(start_in[137]) );
  AND U6028 ( .A(start_reg[138]), .B(init), .Z(start_in[138]) );
  AND U6029 ( .A(start_reg[139]), .B(init), .Z(start_in[139]) );
  AND U6030 ( .A(start_reg[13]), .B(init), .Z(start_in[13]) );
  AND U6031 ( .A(start_reg[140]), .B(init), .Z(start_in[140]) );
  AND U6032 ( .A(start_reg[141]), .B(init), .Z(start_in[141]) );
  AND U6033 ( .A(start_reg[142]), .B(init), .Z(start_in[142]) );
  AND U6034 ( .A(start_reg[143]), .B(init), .Z(start_in[143]) );
  AND U6035 ( .A(start_reg[144]), .B(init), .Z(start_in[144]) );
  AND U6036 ( .A(start_reg[145]), .B(init), .Z(start_in[145]) );
  AND U6037 ( .A(start_reg[146]), .B(init), .Z(start_in[146]) );
  AND U6038 ( .A(start_reg[147]), .B(init), .Z(start_in[147]) );
  AND U6039 ( .A(start_reg[148]), .B(init), .Z(start_in[148]) );
  AND U6040 ( .A(start_reg[149]), .B(init), .Z(start_in[149]) );
  AND U6041 ( .A(start_reg[14]), .B(init), .Z(start_in[14]) );
  AND U6042 ( .A(start_reg[150]), .B(init), .Z(start_in[150]) );
  AND U6043 ( .A(start_reg[151]), .B(init), .Z(start_in[151]) );
  AND U6044 ( .A(start_reg[152]), .B(init), .Z(start_in[152]) );
  AND U6045 ( .A(start_reg[153]), .B(init), .Z(start_in[153]) );
  AND U6046 ( .A(start_reg[154]), .B(init), .Z(start_in[154]) );
  AND U6047 ( .A(start_reg[155]), .B(init), .Z(start_in[155]) );
  AND U6048 ( .A(start_reg[156]), .B(init), .Z(start_in[156]) );
  AND U6049 ( .A(start_reg[157]), .B(init), .Z(start_in[157]) );
  AND U6050 ( .A(start_reg[158]), .B(init), .Z(start_in[158]) );
  AND U6051 ( .A(start_reg[159]), .B(init), .Z(start_in[159]) );
  AND U6052 ( .A(start_reg[15]), .B(init), .Z(start_in[15]) );
  AND U6053 ( .A(start_reg[160]), .B(init), .Z(start_in[160]) );
  AND U6054 ( .A(start_reg[161]), .B(init), .Z(start_in[161]) );
  AND U6055 ( .A(start_reg[162]), .B(init), .Z(start_in[162]) );
  AND U6056 ( .A(start_reg[163]), .B(init), .Z(start_in[163]) );
  AND U6057 ( .A(start_reg[164]), .B(init), .Z(start_in[164]) );
  AND U6058 ( .A(start_reg[165]), .B(init), .Z(start_in[165]) );
  AND U6059 ( .A(start_reg[166]), .B(init), .Z(start_in[166]) );
  AND U6060 ( .A(start_reg[167]), .B(init), .Z(start_in[167]) );
  AND U6061 ( .A(start_reg[168]), .B(init), .Z(start_in[168]) );
  AND U6062 ( .A(start_reg[169]), .B(init), .Z(start_in[169]) );
  AND U6063 ( .A(start_reg[16]), .B(init), .Z(start_in[16]) );
  AND U6064 ( .A(start_reg[170]), .B(init), .Z(start_in[170]) );
  AND U6065 ( .A(start_reg[171]), .B(init), .Z(start_in[171]) );
  AND U6066 ( .A(start_reg[172]), .B(init), .Z(start_in[172]) );
  AND U6067 ( .A(start_reg[173]), .B(init), .Z(start_in[173]) );
  AND U6068 ( .A(start_reg[174]), .B(init), .Z(start_in[174]) );
  AND U6069 ( .A(start_reg[175]), .B(init), .Z(start_in[175]) );
  AND U6070 ( .A(start_reg[176]), .B(init), .Z(start_in[176]) );
  AND U6071 ( .A(start_reg[177]), .B(init), .Z(start_in[177]) );
  AND U6072 ( .A(start_reg[178]), .B(init), .Z(start_in[178]) );
  AND U6073 ( .A(start_reg[179]), .B(init), .Z(start_in[179]) );
  AND U6074 ( .A(start_reg[17]), .B(init), .Z(start_in[17]) );
  AND U6075 ( .A(start_reg[180]), .B(init), .Z(start_in[180]) );
  AND U6076 ( .A(start_reg[181]), .B(init), .Z(start_in[181]) );
  AND U6077 ( .A(start_reg[182]), .B(init), .Z(start_in[182]) );
  AND U6078 ( .A(start_reg[183]), .B(init), .Z(start_in[183]) );
  AND U6079 ( .A(start_reg[184]), .B(init), .Z(start_in[184]) );
  AND U6080 ( .A(start_reg[185]), .B(init), .Z(start_in[185]) );
  AND U6081 ( .A(start_reg[186]), .B(init), .Z(start_in[186]) );
  AND U6082 ( .A(start_reg[187]), .B(init), .Z(start_in[187]) );
  AND U6083 ( .A(start_reg[188]), .B(init), .Z(start_in[188]) );
  AND U6084 ( .A(start_reg[189]), .B(init), .Z(start_in[189]) );
  AND U6085 ( .A(start_reg[18]), .B(init), .Z(start_in[18]) );
  AND U6086 ( .A(start_reg[190]), .B(init), .Z(start_in[190]) );
  AND U6087 ( .A(start_reg[191]), .B(init), .Z(start_in[191]) );
  AND U6088 ( .A(start_reg[192]), .B(init), .Z(start_in[192]) );
  AND U6089 ( .A(start_reg[193]), .B(init), .Z(start_in[193]) );
  AND U6090 ( .A(start_reg[194]), .B(init), .Z(start_in[194]) );
  AND U6091 ( .A(start_reg[195]), .B(init), .Z(start_in[195]) );
  AND U6092 ( .A(start_reg[196]), .B(init), .Z(start_in[196]) );
  AND U6093 ( .A(start_reg[197]), .B(init), .Z(start_in[197]) );
  AND U6094 ( .A(start_reg[198]), .B(init), .Z(start_in[198]) );
  AND U6095 ( .A(start_reg[199]), .B(init), .Z(start_in[199]) );
  AND U6096 ( .A(start_reg[19]), .B(init), .Z(start_in[19]) );
  AND U6097 ( .A(start_reg[1]), .B(init), .Z(start_in[1]) );
  AND U6098 ( .A(start_reg[200]), .B(init), .Z(start_in[200]) );
  AND U6099 ( .A(start_reg[201]), .B(init), .Z(start_in[201]) );
  AND U6100 ( .A(start_reg[202]), .B(init), .Z(start_in[202]) );
  AND U6101 ( .A(start_reg[203]), .B(init), .Z(start_in[203]) );
  AND U6102 ( .A(start_reg[204]), .B(init), .Z(start_in[204]) );
  AND U6103 ( .A(start_reg[205]), .B(init), .Z(start_in[205]) );
  AND U6104 ( .A(start_reg[206]), .B(init), .Z(start_in[206]) );
  AND U6105 ( .A(start_reg[207]), .B(init), .Z(start_in[207]) );
  AND U6106 ( .A(start_reg[208]), .B(init), .Z(start_in[208]) );
  AND U6107 ( .A(start_reg[209]), .B(init), .Z(start_in[209]) );
  AND U6108 ( .A(start_reg[20]), .B(init), .Z(start_in[20]) );
  AND U6109 ( .A(start_reg[210]), .B(init), .Z(start_in[210]) );
  AND U6110 ( .A(start_reg[211]), .B(init), .Z(start_in[211]) );
  AND U6111 ( .A(start_reg[212]), .B(init), .Z(start_in[212]) );
  AND U6112 ( .A(start_reg[213]), .B(init), .Z(start_in[213]) );
  AND U6113 ( .A(start_reg[214]), .B(init), .Z(start_in[214]) );
  AND U6114 ( .A(start_reg[215]), .B(init), .Z(start_in[215]) );
  AND U6115 ( .A(start_reg[216]), .B(init), .Z(start_in[216]) );
  AND U6116 ( .A(start_reg[217]), .B(init), .Z(start_in[217]) );
  AND U6117 ( .A(start_reg[218]), .B(init), .Z(start_in[218]) );
  AND U6118 ( .A(start_reg[219]), .B(init), .Z(start_in[219]) );
  AND U6119 ( .A(start_reg[21]), .B(init), .Z(start_in[21]) );
  AND U6120 ( .A(start_reg[220]), .B(init), .Z(start_in[220]) );
  AND U6121 ( .A(start_reg[221]), .B(init), .Z(start_in[221]) );
  AND U6122 ( .A(start_reg[222]), .B(init), .Z(start_in[222]) );
  AND U6123 ( .A(start_reg[223]), .B(init), .Z(start_in[223]) );
  AND U6124 ( .A(start_reg[224]), .B(init), .Z(start_in[224]) );
  AND U6125 ( .A(start_reg[225]), .B(init), .Z(start_in[225]) );
  AND U6126 ( .A(start_reg[226]), .B(init), .Z(start_in[226]) );
  AND U6127 ( .A(start_reg[227]), .B(init), .Z(start_in[227]) );
  AND U6128 ( .A(start_reg[228]), .B(init), .Z(start_in[228]) );
  AND U6129 ( .A(start_reg[229]), .B(init), .Z(start_in[229]) );
  AND U6130 ( .A(start_reg[22]), .B(init), .Z(start_in[22]) );
  AND U6131 ( .A(start_reg[230]), .B(init), .Z(start_in[230]) );
  AND U6132 ( .A(start_reg[231]), .B(init), .Z(start_in[231]) );
  AND U6133 ( .A(start_reg[232]), .B(init), .Z(start_in[232]) );
  AND U6134 ( .A(start_reg[233]), .B(init), .Z(start_in[233]) );
  AND U6135 ( .A(start_reg[234]), .B(init), .Z(start_in[234]) );
  AND U6136 ( .A(start_reg[235]), .B(init), .Z(start_in[235]) );
  AND U6137 ( .A(start_reg[236]), .B(init), .Z(start_in[236]) );
  AND U6138 ( .A(start_reg[237]), .B(init), .Z(start_in[237]) );
  AND U6139 ( .A(start_reg[238]), .B(init), .Z(start_in[238]) );
  AND U6140 ( .A(start_reg[239]), .B(init), .Z(start_in[239]) );
  AND U6141 ( .A(start_reg[23]), .B(init), .Z(start_in[23]) );
  AND U6142 ( .A(start_reg[240]), .B(init), .Z(start_in[240]) );
  AND U6143 ( .A(start_reg[241]), .B(init), .Z(start_in[241]) );
  AND U6144 ( .A(start_reg[242]), .B(init), .Z(start_in[242]) );
  AND U6145 ( .A(start_reg[243]), .B(init), .Z(start_in[243]) );
  AND U6146 ( .A(start_reg[244]), .B(init), .Z(start_in[244]) );
  AND U6147 ( .A(start_reg[245]), .B(init), .Z(start_in[245]) );
  AND U6148 ( .A(start_reg[246]), .B(init), .Z(start_in[246]) );
  AND U6149 ( .A(start_reg[247]), .B(init), .Z(start_in[247]) );
  AND U6150 ( .A(start_reg[248]), .B(init), .Z(start_in[248]) );
  AND U6151 ( .A(start_reg[249]), .B(init), .Z(start_in[249]) );
  AND U6152 ( .A(start_reg[24]), .B(init), .Z(start_in[24]) );
  AND U6153 ( .A(start_reg[250]), .B(init), .Z(start_in[250]) );
  AND U6154 ( .A(start_reg[251]), .B(init), .Z(start_in[251]) );
  AND U6155 ( .A(start_reg[252]), .B(init), .Z(start_in[252]) );
  AND U6156 ( .A(start_reg[253]), .B(init), .Z(start_in[253]) );
  AND U6157 ( .A(start_reg[254]), .B(init), .Z(start_in[254]) );
  AND U6158 ( .A(start_reg[255]), .B(init), .Z(start_in[255]) );
  AND U6159 ( .A(start_reg[256]), .B(init), .Z(start_in[256]) );
  AND U6160 ( .A(start_reg[257]), .B(init), .Z(start_in[257]) );
  AND U6161 ( .A(start_reg[258]), .B(init), .Z(start_in[258]) );
  AND U6162 ( .A(start_reg[259]), .B(init), .Z(start_in[259]) );
  AND U6163 ( .A(start_reg[25]), .B(init), .Z(start_in[25]) );
  AND U6164 ( .A(start_reg[260]), .B(init), .Z(start_in[260]) );
  AND U6165 ( .A(start_reg[261]), .B(init), .Z(start_in[261]) );
  AND U6166 ( .A(start_reg[262]), .B(init), .Z(start_in[262]) );
  AND U6167 ( .A(start_reg[263]), .B(init), .Z(start_in[263]) );
  AND U6168 ( .A(start_reg[264]), .B(init), .Z(start_in[264]) );
  AND U6169 ( .A(start_reg[265]), .B(init), .Z(start_in[265]) );
  AND U6170 ( .A(start_reg[266]), .B(init), .Z(start_in[266]) );
  AND U6171 ( .A(start_reg[267]), .B(init), .Z(start_in[267]) );
  AND U6172 ( .A(start_reg[268]), .B(init), .Z(start_in[268]) );
  AND U6173 ( .A(start_reg[269]), .B(init), .Z(start_in[269]) );
  AND U6174 ( .A(start_reg[26]), .B(init), .Z(start_in[26]) );
  AND U6175 ( .A(start_reg[270]), .B(init), .Z(start_in[270]) );
  AND U6176 ( .A(start_reg[271]), .B(init), .Z(start_in[271]) );
  AND U6177 ( .A(start_reg[272]), .B(init), .Z(start_in[272]) );
  AND U6178 ( .A(start_reg[273]), .B(init), .Z(start_in[273]) );
  AND U6179 ( .A(start_reg[274]), .B(init), .Z(start_in[274]) );
  AND U6180 ( .A(start_reg[275]), .B(init), .Z(start_in[275]) );
  AND U6181 ( .A(start_reg[276]), .B(init), .Z(start_in[276]) );
  AND U6182 ( .A(start_reg[277]), .B(init), .Z(start_in[277]) );
  AND U6183 ( .A(start_reg[278]), .B(init), .Z(start_in[278]) );
  AND U6184 ( .A(start_reg[279]), .B(init), .Z(start_in[279]) );
  AND U6185 ( .A(start_reg[27]), .B(init), .Z(start_in[27]) );
  AND U6186 ( .A(start_reg[280]), .B(init), .Z(start_in[280]) );
  AND U6187 ( .A(start_reg[281]), .B(init), .Z(start_in[281]) );
  AND U6188 ( .A(start_reg[282]), .B(init), .Z(start_in[282]) );
  AND U6189 ( .A(start_reg[283]), .B(init), .Z(start_in[283]) );
  AND U6190 ( .A(start_reg[284]), .B(init), .Z(start_in[284]) );
  AND U6191 ( .A(start_reg[285]), .B(init), .Z(start_in[285]) );
  AND U6192 ( .A(start_reg[286]), .B(init), .Z(start_in[286]) );
  AND U6193 ( .A(start_reg[287]), .B(init), .Z(start_in[287]) );
  AND U6194 ( .A(start_reg[288]), .B(init), .Z(start_in[288]) );
  AND U6195 ( .A(start_reg[289]), .B(init), .Z(start_in[289]) );
  AND U6196 ( .A(start_reg[28]), .B(init), .Z(start_in[28]) );
  AND U6197 ( .A(start_reg[290]), .B(init), .Z(start_in[290]) );
  AND U6198 ( .A(start_reg[291]), .B(init), .Z(start_in[291]) );
  AND U6199 ( .A(start_reg[292]), .B(init), .Z(start_in[292]) );
  AND U6200 ( .A(start_reg[293]), .B(init), .Z(start_in[293]) );
  AND U6201 ( .A(start_reg[294]), .B(init), .Z(start_in[294]) );
  AND U6202 ( .A(start_reg[295]), .B(init), .Z(start_in[295]) );
  AND U6203 ( .A(start_reg[296]), .B(init), .Z(start_in[296]) );
  AND U6204 ( .A(start_reg[297]), .B(init), .Z(start_in[297]) );
  AND U6205 ( .A(start_reg[298]), .B(init), .Z(start_in[298]) );
  AND U6206 ( .A(start_reg[299]), .B(init), .Z(start_in[299]) );
  AND U6207 ( .A(start_reg[29]), .B(init), .Z(start_in[29]) );
  AND U6208 ( .A(start_reg[2]), .B(init), .Z(start_in[2]) );
  AND U6209 ( .A(start_reg[300]), .B(init), .Z(start_in[300]) );
  AND U6210 ( .A(start_reg[301]), .B(init), .Z(start_in[301]) );
  AND U6211 ( .A(start_reg[302]), .B(init), .Z(start_in[302]) );
  AND U6212 ( .A(start_reg[303]), .B(init), .Z(start_in[303]) );
  AND U6213 ( .A(start_reg[304]), .B(init), .Z(start_in[304]) );
  AND U6214 ( .A(start_reg[305]), .B(init), .Z(start_in[305]) );
  AND U6215 ( .A(start_reg[306]), .B(init), .Z(start_in[306]) );
  AND U6216 ( .A(start_reg[307]), .B(init), .Z(start_in[307]) );
  AND U6217 ( .A(start_reg[308]), .B(init), .Z(start_in[308]) );
  AND U6218 ( .A(start_reg[309]), .B(init), .Z(start_in[309]) );
  AND U6219 ( .A(start_reg[30]), .B(init), .Z(start_in[30]) );
  AND U6220 ( .A(start_reg[310]), .B(init), .Z(start_in[310]) );
  AND U6221 ( .A(start_reg[311]), .B(init), .Z(start_in[311]) );
  AND U6222 ( .A(start_reg[312]), .B(init), .Z(start_in[312]) );
  AND U6223 ( .A(start_reg[313]), .B(init), .Z(start_in[313]) );
  AND U6224 ( .A(start_reg[314]), .B(init), .Z(start_in[314]) );
  AND U6225 ( .A(start_reg[315]), .B(init), .Z(start_in[315]) );
  AND U6226 ( .A(start_reg[316]), .B(init), .Z(start_in[316]) );
  AND U6227 ( .A(start_reg[317]), .B(init), .Z(start_in[317]) );
  AND U6228 ( .A(start_reg[318]), .B(init), .Z(start_in[318]) );
  AND U6229 ( .A(start_reg[319]), .B(init), .Z(start_in[319]) );
  AND U6230 ( .A(start_reg[31]), .B(init), .Z(start_in[31]) );
  AND U6231 ( .A(start_reg[320]), .B(init), .Z(start_in[320]) );
  AND U6232 ( .A(start_reg[321]), .B(init), .Z(start_in[321]) );
  AND U6233 ( .A(start_reg[322]), .B(init), .Z(start_in[322]) );
  AND U6234 ( .A(start_reg[323]), .B(init), .Z(start_in[323]) );
  AND U6235 ( .A(start_reg[324]), .B(init), .Z(start_in[324]) );
  AND U6236 ( .A(start_reg[325]), .B(init), .Z(start_in[325]) );
  AND U6237 ( .A(start_reg[326]), .B(init), .Z(start_in[326]) );
  AND U6238 ( .A(start_reg[327]), .B(init), .Z(start_in[327]) );
  AND U6239 ( .A(start_reg[328]), .B(init), .Z(start_in[328]) );
  AND U6240 ( .A(start_reg[329]), .B(init), .Z(start_in[329]) );
  AND U6241 ( .A(start_reg[32]), .B(init), .Z(start_in[32]) );
  AND U6242 ( .A(start_reg[330]), .B(init), .Z(start_in[330]) );
  AND U6243 ( .A(start_reg[331]), .B(init), .Z(start_in[331]) );
  AND U6244 ( .A(start_reg[332]), .B(init), .Z(start_in[332]) );
  AND U6245 ( .A(start_reg[333]), .B(init), .Z(start_in[333]) );
  AND U6246 ( .A(start_reg[334]), .B(init), .Z(start_in[334]) );
  AND U6247 ( .A(start_reg[335]), .B(init), .Z(start_in[335]) );
  AND U6248 ( .A(start_reg[336]), .B(init), .Z(start_in[336]) );
  AND U6249 ( .A(start_reg[337]), .B(init), .Z(start_in[337]) );
  AND U6250 ( .A(start_reg[338]), .B(init), .Z(start_in[338]) );
  AND U6251 ( .A(start_reg[339]), .B(init), .Z(start_in[339]) );
  AND U6252 ( .A(start_reg[33]), .B(init), .Z(start_in[33]) );
  AND U6253 ( .A(start_reg[340]), .B(init), .Z(start_in[340]) );
  AND U6254 ( .A(start_reg[341]), .B(init), .Z(start_in[341]) );
  AND U6255 ( .A(start_reg[342]), .B(init), .Z(start_in[342]) );
  AND U6256 ( .A(start_reg[343]), .B(init), .Z(start_in[343]) );
  AND U6257 ( .A(start_reg[344]), .B(init), .Z(start_in[344]) );
  AND U6258 ( .A(start_reg[345]), .B(init), .Z(start_in[345]) );
  AND U6259 ( .A(start_reg[346]), .B(init), .Z(start_in[346]) );
  AND U6260 ( .A(start_reg[347]), .B(init), .Z(start_in[347]) );
  AND U6261 ( .A(start_reg[348]), .B(init), .Z(start_in[348]) );
  AND U6262 ( .A(start_reg[349]), .B(init), .Z(start_in[349]) );
  AND U6263 ( .A(start_reg[34]), .B(init), .Z(start_in[34]) );
  AND U6264 ( .A(start_reg[350]), .B(init), .Z(start_in[350]) );
  AND U6265 ( .A(start_reg[351]), .B(init), .Z(start_in[351]) );
  AND U6266 ( .A(start_reg[352]), .B(init), .Z(start_in[352]) );
  AND U6267 ( .A(start_reg[353]), .B(init), .Z(start_in[353]) );
  AND U6268 ( .A(start_reg[354]), .B(init), .Z(start_in[354]) );
  AND U6269 ( .A(start_reg[355]), .B(init), .Z(start_in[355]) );
  AND U6270 ( .A(start_reg[356]), .B(init), .Z(start_in[356]) );
  AND U6271 ( .A(start_reg[357]), .B(init), .Z(start_in[357]) );
  AND U6272 ( .A(start_reg[358]), .B(init), .Z(start_in[358]) );
  AND U6273 ( .A(start_reg[359]), .B(init), .Z(start_in[359]) );
  AND U6274 ( .A(start_reg[35]), .B(init), .Z(start_in[35]) );
  AND U6275 ( .A(start_reg[360]), .B(init), .Z(start_in[360]) );
  AND U6276 ( .A(start_reg[361]), .B(init), .Z(start_in[361]) );
  AND U6277 ( .A(start_reg[362]), .B(init), .Z(start_in[362]) );
  AND U6278 ( .A(start_reg[363]), .B(init), .Z(start_in[363]) );
  AND U6279 ( .A(start_reg[364]), .B(init), .Z(start_in[364]) );
  AND U6280 ( .A(start_reg[365]), .B(init), .Z(start_in[365]) );
  AND U6281 ( .A(start_reg[366]), .B(init), .Z(start_in[366]) );
  AND U6282 ( .A(start_reg[367]), .B(init), .Z(start_in[367]) );
  AND U6283 ( .A(start_reg[368]), .B(init), .Z(start_in[368]) );
  AND U6284 ( .A(start_reg[369]), .B(init), .Z(start_in[369]) );
  AND U6285 ( .A(start_reg[36]), .B(init), .Z(start_in[36]) );
  AND U6286 ( .A(start_reg[370]), .B(init), .Z(start_in[370]) );
  AND U6287 ( .A(start_reg[371]), .B(init), .Z(start_in[371]) );
  AND U6288 ( .A(start_reg[372]), .B(init), .Z(start_in[372]) );
  AND U6289 ( .A(start_reg[373]), .B(init), .Z(start_in[373]) );
  AND U6290 ( .A(start_reg[374]), .B(init), .Z(start_in[374]) );
  AND U6291 ( .A(start_reg[375]), .B(init), .Z(start_in[375]) );
  AND U6292 ( .A(start_reg[376]), .B(init), .Z(start_in[376]) );
  AND U6293 ( .A(start_reg[377]), .B(init), .Z(start_in[377]) );
  AND U6294 ( .A(start_reg[378]), .B(init), .Z(start_in[378]) );
  AND U6295 ( .A(start_reg[379]), .B(init), .Z(start_in[379]) );
  AND U6296 ( .A(start_reg[37]), .B(init), .Z(start_in[37]) );
  AND U6297 ( .A(start_reg[380]), .B(init), .Z(start_in[380]) );
  AND U6298 ( .A(start_reg[381]), .B(init), .Z(start_in[381]) );
  AND U6299 ( .A(start_reg[382]), .B(init), .Z(start_in[382]) );
  AND U6300 ( .A(start_reg[383]), .B(init), .Z(start_in[383]) );
  AND U6301 ( .A(start_reg[384]), .B(init), .Z(start_in[384]) );
  AND U6302 ( .A(start_reg[385]), .B(init), .Z(start_in[385]) );
  AND U6303 ( .A(start_reg[386]), .B(init), .Z(start_in[386]) );
  AND U6304 ( .A(start_reg[387]), .B(init), .Z(start_in[387]) );
  AND U6305 ( .A(start_reg[388]), .B(init), .Z(start_in[388]) );
  AND U6306 ( .A(start_reg[389]), .B(init), .Z(start_in[389]) );
  AND U6307 ( .A(start_reg[38]), .B(init), .Z(start_in[38]) );
  AND U6308 ( .A(start_reg[390]), .B(init), .Z(start_in[390]) );
  AND U6309 ( .A(start_reg[391]), .B(init), .Z(start_in[391]) );
  AND U6310 ( .A(start_reg[392]), .B(init), .Z(start_in[392]) );
  AND U6311 ( .A(start_reg[393]), .B(init), .Z(start_in[393]) );
  AND U6312 ( .A(start_reg[394]), .B(init), .Z(start_in[394]) );
  AND U6313 ( .A(start_reg[395]), .B(init), .Z(start_in[395]) );
  AND U6314 ( .A(start_reg[396]), .B(init), .Z(start_in[396]) );
  AND U6315 ( .A(start_reg[397]), .B(init), .Z(start_in[397]) );
  AND U6316 ( .A(start_reg[398]), .B(init), .Z(start_in[398]) );
  AND U6317 ( .A(start_reg[399]), .B(init), .Z(start_in[399]) );
  AND U6318 ( .A(start_reg[39]), .B(init), .Z(start_in[39]) );
  AND U6319 ( .A(start_reg[3]), .B(init), .Z(start_in[3]) );
  AND U6320 ( .A(start_reg[400]), .B(init), .Z(start_in[400]) );
  AND U6321 ( .A(start_reg[401]), .B(init), .Z(start_in[401]) );
  AND U6322 ( .A(start_reg[402]), .B(init), .Z(start_in[402]) );
  AND U6323 ( .A(start_reg[403]), .B(init), .Z(start_in[403]) );
  AND U6324 ( .A(start_reg[404]), .B(init), .Z(start_in[404]) );
  AND U6325 ( .A(start_reg[405]), .B(init), .Z(start_in[405]) );
  AND U6326 ( .A(start_reg[406]), .B(init), .Z(start_in[406]) );
  AND U6327 ( .A(start_reg[407]), .B(init), .Z(start_in[407]) );
  AND U6328 ( .A(start_reg[408]), .B(init), .Z(start_in[408]) );
  AND U6329 ( .A(start_reg[409]), .B(init), .Z(start_in[409]) );
  AND U6330 ( .A(start_reg[40]), .B(init), .Z(start_in[40]) );
  AND U6331 ( .A(start_reg[410]), .B(init), .Z(start_in[410]) );
  AND U6332 ( .A(start_reg[411]), .B(init), .Z(start_in[411]) );
  AND U6333 ( .A(start_reg[412]), .B(init), .Z(start_in[412]) );
  AND U6334 ( .A(start_reg[413]), .B(init), .Z(start_in[413]) );
  AND U6335 ( .A(start_reg[414]), .B(init), .Z(start_in[414]) );
  AND U6336 ( .A(start_reg[415]), .B(init), .Z(start_in[415]) );
  AND U6337 ( .A(start_reg[416]), .B(init), .Z(start_in[416]) );
  AND U6338 ( .A(start_reg[417]), .B(init), .Z(start_in[417]) );
  AND U6339 ( .A(start_reg[418]), .B(init), .Z(start_in[418]) );
  AND U6340 ( .A(start_reg[419]), .B(init), .Z(start_in[419]) );
  AND U6341 ( .A(start_reg[41]), .B(init), .Z(start_in[41]) );
  AND U6342 ( .A(start_reg[420]), .B(init), .Z(start_in[420]) );
  AND U6343 ( .A(start_reg[421]), .B(init), .Z(start_in[421]) );
  AND U6344 ( .A(start_reg[422]), .B(init), .Z(start_in[422]) );
  AND U6345 ( .A(start_reg[423]), .B(init), .Z(start_in[423]) );
  AND U6346 ( .A(start_reg[424]), .B(init), .Z(start_in[424]) );
  AND U6347 ( .A(start_reg[425]), .B(init), .Z(start_in[425]) );
  AND U6348 ( .A(start_reg[426]), .B(init), .Z(start_in[426]) );
  AND U6349 ( .A(start_reg[427]), .B(init), .Z(start_in[427]) );
  AND U6350 ( .A(start_reg[428]), .B(init), .Z(start_in[428]) );
  AND U6351 ( .A(start_reg[429]), .B(init), .Z(start_in[429]) );
  AND U6352 ( .A(start_reg[42]), .B(init), .Z(start_in[42]) );
  AND U6353 ( .A(start_reg[430]), .B(init), .Z(start_in[430]) );
  AND U6354 ( .A(start_reg[431]), .B(init), .Z(start_in[431]) );
  AND U6355 ( .A(start_reg[432]), .B(init), .Z(start_in[432]) );
  AND U6356 ( .A(start_reg[433]), .B(init), .Z(start_in[433]) );
  AND U6357 ( .A(start_reg[434]), .B(init), .Z(start_in[434]) );
  AND U6358 ( .A(start_reg[435]), .B(init), .Z(start_in[435]) );
  AND U6359 ( .A(start_reg[436]), .B(init), .Z(start_in[436]) );
  AND U6360 ( .A(start_reg[437]), .B(init), .Z(start_in[437]) );
  AND U6361 ( .A(start_reg[438]), .B(init), .Z(start_in[438]) );
  AND U6362 ( .A(start_reg[439]), .B(init), .Z(start_in[439]) );
  AND U6363 ( .A(start_reg[43]), .B(init), .Z(start_in[43]) );
  AND U6364 ( .A(start_reg[440]), .B(init), .Z(start_in[440]) );
  AND U6365 ( .A(start_reg[441]), .B(init), .Z(start_in[441]) );
  AND U6366 ( .A(start_reg[442]), .B(init), .Z(start_in[442]) );
  AND U6367 ( .A(start_reg[443]), .B(init), .Z(start_in[443]) );
  AND U6368 ( .A(start_reg[444]), .B(init), .Z(start_in[444]) );
  AND U6369 ( .A(start_reg[445]), .B(init), .Z(start_in[445]) );
  AND U6370 ( .A(start_reg[446]), .B(init), .Z(start_in[446]) );
  AND U6371 ( .A(start_reg[447]), .B(init), .Z(start_in[447]) );
  AND U6372 ( .A(start_reg[448]), .B(init), .Z(start_in[448]) );
  AND U6373 ( .A(start_reg[449]), .B(init), .Z(start_in[449]) );
  AND U6374 ( .A(start_reg[44]), .B(init), .Z(start_in[44]) );
  AND U6375 ( .A(start_reg[450]), .B(init), .Z(start_in[450]) );
  AND U6376 ( .A(start_reg[451]), .B(init), .Z(start_in[451]) );
  AND U6377 ( .A(start_reg[452]), .B(init), .Z(start_in[452]) );
  AND U6378 ( .A(start_reg[453]), .B(init), .Z(start_in[453]) );
  AND U6379 ( .A(start_reg[454]), .B(init), .Z(start_in[454]) );
  AND U6380 ( .A(start_reg[455]), .B(init), .Z(start_in[455]) );
  AND U6381 ( .A(start_reg[456]), .B(init), .Z(start_in[456]) );
  AND U6382 ( .A(start_reg[457]), .B(init), .Z(start_in[457]) );
  AND U6383 ( .A(start_reg[458]), .B(init), .Z(start_in[458]) );
  AND U6384 ( .A(start_reg[459]), .B(init), .Z(start_in[459]) );
  AND U6385 ( .A(start_reg[45]), .B(init), .Z(start_in[45]) );
  AND U6386 ( .A(start_reg[460]), .B(init), .Z(start_in[460]) );
  AND U6387 ( .A(start_reg[461]), .B(init), .Z(start_in[461]) );
  AND U6388 ( .A(start_reg[462]), .B(init), .Z(start_in[462]) );
  AND U6389 ( .A(start_reg[463]), .B(init), .Z(start_in[463]) );
  AND U6390 ( .A(start_reg[464]), .B(init), .Z(start_in[464]) );
  AND U6391 ( .A(start_reg[465]), .B(init), .Z(start_in[465]) );
  AND U6392 ( .A(start_reg[466]), .B(init), .Z(start_in[466]) );
  AND U6393 ( .A(start_reg[467]), .B(init), .Z(start_in[467]) );
  AND U6394 ( .A(start_reg[468]), .B(init), .Z(start_in[468]) );
  AND U6395 ( .A(start_reg[469]), .B(init), .Z(start_in[469]) );
  AND U6396 ( .A(start_reg[46]), .B(init), .Z(start_in[46]) );
  AND U6397 ( .A(start_reg[470]), .B(init), .Z(start_in[470]) );
  AND U6398 ( .A(start_reg[471]), .B(init), .Z(start_in[471]) );
  AND U6399 ( .A(start_reg[472]), .B(init), .Z(start_in[472]) );
  AND U6400 ( .A(start_reg[473]), .B(init), .Z(start_in[473]) );
  AND U6401 ( .A(start_reg[474]), .B(init), .Z(start_in[474]) );
  AND U6402 ( .A(start_reg[475]), .B(init), .Z(start_in[475]) );
  AND U6403 ( .A(start_reg[476]), .B(init), .Z(start_in[476]) );
  AND U6404 ( .A(start_reg[477]), .B(init), .Z(start_in[477]) );
  AND U6405 ( .A(start_reg[478]), .B(init), .Z(start_in[478]) );
  AND U6406 ( .A(start_reg[479]), .B(init), .Z(start_in[479]) );
  AND U6407 ( .A(start_reg[47]), .B(init), .Z(start_in[47]) );
  AND U6408 ( .A(start_reg[480]), .B(init), .Z(start_in[480]) );
  AND U6409 ( .A(start_reg[481]), .B(init), .Z(start_in[481]) );
  AND U6410 ( .A(start_reg[482]), .B(init), .Z(start_in[482]) );
  AND U6411 ( .A(start_reg[483]), .B(init), .Z(start_in[483]) );
  AND U6412 ( .A(start_reg[484]), .B(init), .Z(start_in[484]) );
  AND U6413 ( .A(start_reg[485]), .B(init), .Z(start_in[485]) );
  AND U6414 ( .A(start_reg[486]), .B(init), .Z(start_in[486]) );
  AND U6415 ( .A(start_reg[487]), .B(init), .Z(start_in[487]) );
  AND U6416 ( .A(start_reg[488]), .B(init), .Z(start_in[488]) );
  AND U6417 ( .A(start_reg[489]), .B(init), .Z(start_in[489]) );
  AND U6418 ( .A(start_reg[48]), .B(init), .Z(start_in[48]) );
  AND U6419 ( .A(start_reg[490]), .B(init), .Z(start_in[490]) );
  AND U6420 ( .A(start_reg[491]), .B(init), .Z(start_in[491]) );
  AND U6421 ( .A(start_reg[492]), .B(init), .Z(start_in[492]) );
  AND U6422 ( .A(start_reg[493]), .B(init), .Z(start_in[493]) );
  AND U6423 ( .A(start_reg[494]), .B(init), .Z(start_in[494]) );
  AND U6424 ( .A(start_reg[495]), .B(init), .Z(start_in[495]) );
  AND U6425 ( .A(start_reg[496]), .B(init), .Z(start_in[496]) );
  AND U6426 ( .A(start_reg[497]), .B(init), .Z(start_in[497]) );
  AND U6427 ( .A(start_reg[498]), .B(init), .Z(start_in[498]) );
  AND U6428 ( .A(start_reg[499]), .B(init), .Z(start_in[499]) );
  AND U6429 ( .A(start_reg[49]), .B(init), .Z(start_in[49]) );
  AND U6430 ( .A(start_reg[4]), .B(init), .Z(start_in[4]) );
  AND U6431 ( .A(start_reg[500]), .B(init), .Z(start_in[500]) );
  AND U6432 ( .A(start_reg[501]), .B(init), .Z(start_in[501]) );
  AND U6433 ( .A(start_reg[502]), .B(init), .Z(start_in[502]) );
  AND U6434 ( .A(start_reg[503]), .B(init), .Z(start_in[503]) );
  AND U6435 ( .A(start_reg[504]), .B(init), .Z(start_in[504]) );
  AND U6436 ( .A(start_reg[505]), .B(init), .Z(start_in[505]) );
  AND U6437 ( .A(start_reg[506]), .B(init), .Z(start_in[506]) );
  AND U6438 ( .A(start_reg[507]), .B(init), .Z(start_in[507]) );
  AND U6439 ( .A(start_reg[508]), .B(init), .Z(start_in[508]) );
  AND U6440 ( .A(start_reg[509]), .B(init), .Z(start_in[509]) );
  AND U6441 ( .A(start_reg[50]), .B(init), .Z(start_in[50]) );
  AND U6442 ( .A(start_reg[510]), .B(init), .Z(start_in[510]) );
  AND U6443 ( .A(start_reg[51]), .B(init), .Z(start_in[51]) );
  AND U6444 ( .A(start_reg[52]), .B(init), .Z(start_in[52]) );
  AND U6445 ( .A(start_reg[53]), .B(init), .Z(start_in[53]) );
  AND U6446 ( .A(start_reg[54]), .B(init), .Z(start_in[54]) );
  AND U6447 ( .A(start_reg[55]), .B(init), .Z(start_in[55]) );
  AND U6448 ( .A(start_reg[56]), .B(init), .Z(start_in[56]) );
  AND U6449 ( .A(start_reg[57]), .B(init), .Z(start_in[57]) );
  AND U6450 ( .A(start_reg[58]), .B(init), .Z(start_in[58]) );
  AND U6451 ( .A(start_reg[59]), .B(init), .Z(start_in[59]) );
  AND U6452 ( .A(start_reg[5]), .B(init), .Z(start_in[5]) );
  AND U6453 ( .A(start_reg[60]), .B(init), .Z(start_in[60]) );
  AND U6454 ( .A(start_reg[61]), .B(init), .Z(start_in[61]) );
  AND U6455 ( .A(start_reg[62]), .B(init), .Z(start_in[62]) );
  AND U6456 ( .A(start_reg[63]), .B(init), .Z(start_in[63]) );
  AND U6457 ( .A(start_reg[64]), .B(init), .Z(start_in[64]) );
  AND U6458 ( .A(start_reg[65]), .B(init), .Z(start_in[65]) );
  AND U6459 ( .A(start_reg[66]), .B(init), .Z(start_in[66]) );
  AND U6460 ( .A(start_reg[67]), .B(init), .Z(start_in[67]) );
  AND U6461 ( .A(start_reg[68]), .B(init), .Z(start_in[68]) );
  AND U6462 ( .A(start_reg[69]), .B(init), .Z(start_in[69]) );
  AND U6463 ( .A(start_reg[6]), .B(init), .Z(start_in[6]) );
  AND U6464 ( .A(start_reg[70]), .B(init), .Z(start_in[70]) );
  AND U6465 ( .A(start_reg[71]), .B(init), .Z(start_in[71]) );
  AND U6466 ( .A(start_reg[72]), .B(init), .Z(start_in[72]) );
  AND U6467 ( .A(start_reg[73]), .B(init), .Z(start_in[73]) );
  AND U6468 ( .A(start_reg[74]), .B(init), .Z(start_in[74]) );
  AND U6469 ( .A(start_reg[75]), .B(init), .Z(start_in[75]) );
  AND U6470 ( .A(start_reg[76]), .B(init), .Z(start_in[76]) );
  AND U6471 ( .A(start_reg[77]), .B(init), .Z(start_in[77]) );
  AND U6472 ( .A(start_reg[78]), .B(init), .Z(start_in[78]) );
  AND U6473 ( .A(start_reg[79]), .B(init), .Z(start_in[79]) );
  AND U6474 ( .A(start_reg[7]), .B(init), .Z(start_in[7]) );
  AND U6475 ( .A(start_reg[80]), .B(init), .Z(start_in[80]) );
  AND U6476 ( .A(start_reg[81]), .B(init), .Z(start_in[81]) );
  AND U6477 ( .A(start_reg[82]), .B(init), .Z(start_in[82]) );
  AND U6478 ( .A(start_reg[83]), .B(init), .Z(start_in[83]) );
  AND U6479 ( .A(start_reg[84]), .B(init), .Z(start_in[84]) );
  AND U6480 ( .A(start_reg[85]), .B(init), .Z(start_in[85]) );
  AND U6481 ( .A(start_reg[86]), .B(init), .Z(start_in[86]) );
  AND U6482 ( .A(start_reg[87]), .B(init), .Z(start_in[87]) );
  AND U6483 ( .A(start_reg[88]), .B(init), .Z(start_in[88]) );
  AND U6484 ( .A(start_reg[89]), .B(init), .Z(start_in[89]) );
  AND U6485 ( .A(start_reg[8]), .B(init), .Z(start_in[8]) );
  AND U6486 ( .A(start_reg[90]), .B(init), .Z(start_in[90]) );
  AND U6487 ( .A(start_reg[91]), .B(init), .Z(start_in[91]) );
  AND U6488 ( .A(start_reg[92]), .B(init), .Z(start_in[92]) );
  AND U6489 ( .A(start_reg[93]), .B(init), .Z(start_in[93]) );
  AND U6490 ( .A(start_reg[94]), .B(init), .Z(start_in[94]) );
  AND U6491 ( .A(start_reg[95]), .B(init), .Z(start_in[95]) );
  AND U6492 ( .A(start_reg[96]), .B(init), .Z(start_in[96]) );
  AND U6493 ( .A(start_reg[97]), .B(init), .Z(start_in[97]) );
  AND U6494 ( .A(start_reg[98]), .B(init), .Z(start_in[98]) );
  AND U6495 ( .A(start_reg[99]), .B(init), .Z(start_in[99]) );
  AND U6496 ( .A(start_reg[9]), .B(init), .Z(start_in[9]) );
  NAND U6497 ( .A(n3859), .B(m[0]), .Z(n4446) );
  NAND U6498 ( .A(init), .B(creg[0]), .Z(n4838) );
  NAND U6499 ( .A(n4446), .B(n4838), .Z(x[0]) );
  NAND U6500 ( .A(n3859), .B(m[100]), .Z(n4447) );
  NAND U6501 ( .A(init), .B(creg[100]), .Z(n4841) );
  NAND U6502 ( .A(n4447), .B(n4841), .Z(x[100]) );
  NAND U6503 ( .A(n3859), .B(m[101]), .Z(n4448) );
  NAND U6504 ( .A(init), .B(creg[101]), .Z(n4844) );
  NAND U6505 ( .A(n4448), .B(n4844), .Z(x[101]) );
  NAND U6506 ( .A(n3859), .B(m[102]), .Z(n4449) );
  NAND U6507 ( .A(init), .B(creg[102]), .Z(n4847) );
  NAND U6508 ( .A(n4449), .B(n4847), .Z(x[102]) );
  NAND U6509 ( .A(n3859), .B(m[103]), .Z(n4450) );
  NAND U6510 ( .A(init), .B(creg[103]), .Z(n4850) );
  NAND U6511 ( .A(n4450), .B(n4850), .Z(x[103]) );
  NAND U6512 ( .A(n3860), .B(m[104]), .Z(n4451) );
  NAND U6513 ( .A(init), .B(creg[104]), .Z(n4853) );
  NAND U6514 ( .A(n4451), .B(n4853), .Z(x[104]) );
  NAND U6515 ( .A(init), .B(creg[105]), .Z(n4453) );
  NAND U6516 ( .A(n3860), .B(m[105]), .Z(n4452) );
  NAND U6517 ( .A(n4453), .B(n4452), .Z(x[105]) );
  NAND U6518 ( .A(init), .B(creg[106]), .Z(n4455) );
  NAND U6519 ( .A(n3860), .B(m[106]), .Z(n4454) );
  NAND U6520 ( .A(n4455), .B(n4454), .Z(x[106]) );
  NAND U6521 ( .A(init), .B(creg[107]), .Z(n4457) );
  NAND U6522 ( .A(n3860), .B(m[107]), .Z(n4456) );
  NAND U6523 ( .A(n4457), .B(n4456), .Z(x[107]) );
  NAND U6524 ( .A(n3860), .B(m[108]), .Z(n4458) );
  NAND U6525 ( .A(init), .B(creg[108]), .Z(n4862) );
  NAND U6526 ( .A(n4458), .B(n4862), .Z(x[108]) );
  NAND U6527 ( .A(n3860), .B(m[109]), .Z(n4459) );
  NAND U6528 ( .A(init), .B(creg[109]), .Z(n4865) );
  NAND U6529 ( .A(n4459), .B(n4865), .Z(x[109]) );
  NAND U6530 ( .A(n3860), .B(m[10]), .Z(n4460) );
  NAND U6531 ( .A(init), .B(creg[10]), .Z(n4868) );
  NAND U6532 ( .A(n4460), .B(n4868), .Z(x[10]) );
  NAND U6533 ( .A(init), .B(creg[110]), .Z(n4462) );
  NAND U6534 ( .A(n3861), .B(m[110]), .Z(n4461) );
  NAND U6535 ( .A(n4462), .B(n4461), .Z(x[110]) );
  NAND U6536 ( .A(init), .B(creg[111]), .Z(n4464) );
  NAND U6537 ( .A(n3861), .B(m[111]), .Z(n4463) );
  NAND U6538 ( .A(n4464), .B(n4463), .Z(x[111]) );
  NAND U6539 ( .A(init), .B(creg[112]), .Z(n4466) );
  NAND U6540 ( .A(n3861), .B(m[112]), .Z(n4465) );
  NAND U6541 ( .A(n4466), .B(n4465), .Z(x[112]) );
  NAND U6542 ( .A(n3861), .B(m[113]), .Z(n4467) );
  NAND U6543 ( .A(init), .B(creg[113]), .Z(n4877) );
  NAND U6544 ( .A(n4467), .B(n4877), .Z(x[113]) );
  NAND U6545 ( .A(init), .B(creg[114]), .Z(n4469) );
  NAND U6546 ( .A(n3861), .B(m[114]), .Z(n4468) );
  NAND U6547 ( .A(n4469), .B(n4468), .Z(x[114]) );
  NAND U6548 ( .A(init), .B(creg[115]), .Z(n4471) );
  NAND U6549 ( .A(n3861), .B(m[115]), .Z(n4470) );
  NAND U6550 ( .A(n4471), .B(n4470), .Z(x[115]) );
  NAND U6551 ( .A(n3861), .B(m[116]), .Z(n4472) );
  NAND U6552 ( .A(init), .B(creg[116]), .Z(n4884) );
  NAND U6553 ( .A(n4472), .B(n4884), .Z(x[116]) );
  NAND U6554 ( .A(n3862), .B(m[117]), .Z(n4473) );
  NAND U6555 ( .A(init), .B(creg[117]), .Z(n4887) );
  NAND U6556 ( .A(n4473), .B(n4887), .Z(x[117]) );
  NAND U6557 ( .A(n3862), .B(m[118]), .Z(n4474) );
  NAND U6558 ( .A(init), .B(creg[118]), .Z(n4890) );
  NAND U6559 ( .A(n4474), .B(n4890), .Z(x[118]) );
  NAND U6560 ( .A(n3862), .B(m[119]), .Z(n4475) );
  NAND U6561 ( .A(init), .B(creg[119]), .Z(n4893) );
  NAND U6562 ( .A(n4475), .B(n4893), .Z(x[119]) );
  NAND U6563 ( .A(n3862), .B(m[11]), .Z(n4476) );
  NAND U6564 ( .A(init), .B(creg[11]), .Z(n4896) );
  NAND U6565 ( .A(n4476), .B(n4896), .Z(x[11]) );
  NAND U6566 ( .A(init), .B(creg[120]), .Z(n4478) );
  NAND U6567 ( .A(n3862), .B(m[120]), .Z(n4477) );
  NAND U6568 ( .A(n4478), .B(n4477), .Z(x[120]) );
  NAND U6569 ( .A(init), .B(creg[121]), .Z(n4480) );
  NAND U6570 ( .A(n3862), .B(m[121]), .Z(n4479) );
  NAND U6571 ( .A(n4480), .B(n4479), .Z(x[121]) );
  NAND U6572 ( .A(n3862), .B(m[122]), .Z(n4481) );
  NAND U6573 ( .A(init), .B(creg[122]), .Z(n4903) );
  NAND U6574 ( .A(n4481), .B(n4903), .Z(x[122]) );
  NAND U6575 ( .A(init), .B(creg[123]), .Z(n4483) );
  NAND U6576 ( .A(n3863), .B(m[123]), .Z(n4482) );
  NAND U6577 ( .A(n4483), .B(n4482), .Z(x[123]) );
  NAND U6578 ( .A(init), .B(creg[124]), .Z(n4485) );
  NAND U6579 ( .A(n3863), .B(m[124]), .Z(n4484) );
  NAND U6580 ( .A(n4485), .B(n4484), .Z(x[124]) );
  NAND U6581 ( .A(n3863), .B(m[125]), .Z(n4486) );
  NAND U6582 ( .A(init), .B(creg[125]), .Z(n4910) );
  NAND U6583 ( .A(n4486), .B(n4910), .Z(x[125]) );
  NAND U6584 ( .A(init), .B(creg[126]), .Z(n4488) );
  NAND U6585 ( .A(n3863), .B(m[126]), .Z(n4487) );
  NAND U6586 ( .A(n4488), .B(n4487), .Z(x[126]) );
  NAND U6587 ( .A(init), .B(creg[127]), .Z(n4490) );
  NAND U6588 ( .A(n3863), .B(m[127]), .Z(n4489) );
  NAND U6589 ( .A(n4490), .B(n4489), .Z(x[127]) );
  NAND U6590 ( .A(init), .B(creg[128]), .Z(n4492) );
  NAND U6591 ( .A(n3863), .B(m[128]), .Z(n4491) );
  NAND U6592 ( .A(n4492), .B(n4491), .Z(x[128]) );
  NAND U6593 ( .A(init), .B(creg[129]), .Z(n4494) );
  NAND U6594 ( .A(n3863), .B(m[129]), .Z(n4493) );
  NAND U6595 ( .A(n4494), .B(n4493), .Z(x[129]) );
  NAND U6596 ( .A(n3864), .B(m[12]), .Z(n4495) );
  NAND U6597 ( .A(init), .B(creg[12]), .Z(n4921) );
  NAND U6598 ( .A(n4495), .B(n4921), .Z(x[12]) );
  NAND U6599 ( .A(init), .B(creg[130]), .Z(n4497) );
  NAND U6600 ( .A(n3864), .B(m[130]), .Z(n4496) );
  NAND U6601 ( .A(n4497), .B(n4496), .Z(x[130]) );
  NAND U6602 ( .A(init), .B(creg[131]), .Z(n4499) );
  NAND U6603 ( .A(n3864), .B(m[131]), .Z(n4498) );
  NAND U6604 ( .A(n4499), .B(n4498), .Z(x[131]) );
  NAND U6605 ( .A(init), .B(creg[132]), .Z(n4501) );
  NAND U6606 ( .A(n3864), .B(m[132]), .Z(n4500) );
  NAND U6607 ( .A(n4501), .B(n4500), .Z(x[132]) );
  NAND U6608 ( .A(n3864), .B(m[133]), .Z(n4502) );
  NAND U6609 ( .A(init), .B(creg[133]), .Z(n4930) );
  NAND U6610 ( .A(n4502), .B(n4930), .Z(x[133]) );
  NAND U6611 ( .A(init), .B(creg[134]), .Z(n4504) );
  NAND U6612 ( .A(n3864), .B(m[134]), .Z(n4503) );
  NAND U6613 ( .A(n4504), .B(n4503), .Z(x[134]) );
  NAND U6614 ( .A(init), .B(creg[135]), .Z(n4506) );
  NAND U6615 ( .A(n3864), .B(m[135]), .Z(n4505) );
  NAND U6616 ( .A(n4506), .B(n4505), .Z(x[135]) );
  NAND U6617 ( .A(init), .B(creg[136]), .Z(n4508) );
  NAND U6618 ( .A(n3865), .B(m[136]), .Z(n4507) );
  NAND U6619 ( .A(n4508), .B(n4507), .Z(x[136]) );
  NAND U6620 ( .A(n3865), .B(m[137]), .Z(n4509) );
  NAND U6621 ( .A(init), .B(creg[137]), .Z(n4939) );
  NAND U6622 ( .A(n4509), .B(n4939), .Z(x[137]) );
  NAND U6623 ( .A(n3865), .B(m[138]), .Z(n4510) );
  NAND U6624 ( .A(init), .B(creg[138]), .Z(n4942) );
  NAND U6625 ( .A(n4510), .B(n4942), .Z(x[138]) );
  NAND U6626 ( .A(init), .B(creg[139]), .Z(n4512) );
  NAND U6627 ( .A(n3865), .B(m[139]), .Z(n4511) );
  NAND U6628 ( .A(n4512), .B(n4511), .Z(x[139]) );
  NAND U6629 ( .A(init), .B(creg[13]), .Z(n4514) );
  NAND U6630 ( .A(n3865), .B(m[13]), .Z(n4513) );
  NAND U6631 ( .A(n4514), .B(n4513), .Z(x[13]) );
  NAND U6632 ( .A(n3865), .B(m[140]), .Z(n4515) );
  NAND U6633 ( .A(init), .B(creg[140]), .Z(n4949) );
  NAND U6634 ( .A(n4515), .B(n4949), .Z(x[140]) );
  NAND U6635 ( .A(n3865), .B(m[141]), .Z(n4516) );
  NAND U6636 ( .A(init), .B(creg[141]), .Z(n4952) );
  NAND U6637 ( .A(n4516), .B(n4952), .Z(x[141]) );
  NAND U6638 ( .A(init), .B(creg[142]), .Z(n4518) );
  NAND U6639 ( .A(n3866), .B(m[142]), .Z(n4517) );
  NAND U6640 ( .A(n4518), .B(n4517), .Z(x[142]) );
  NAND U6641 ( .A(init), .B(creg[143]), .Z(n4520) );
  NAND U6642 ( .A(n3866), .B(m[143]), .Z(n4519) );
  NAND U6643 ( .A(n4520), .B(n4519), .Z(x[143]) );
  NAND U6644 ( .A(init), .B(creg[144]), .Z(n4522) );
  NAND U6645 ( .A(n3866), .B(m[144]), .Z(n4521) );
  NAND U6646 ( .A(n4522), .B(n4521), .Z(x[144]) );
  NAND U6647 ( .A(init), .B(creg[145]), .Z(n4524) );
  NAND U6648 ( .A(n3866), .B(m[145]), .Z(n4523) );
  NAND U6649 ( .A(n4524), .B(n4523), .Z(x[145]) );
  NAND U6650 ( .A(init), .B(creg[146]), .Z(n4526) );
  NAND U6651 ( .A(n3866), .B(m[146]), .Z(n4525) );
  NAND U6652 ( .A(n4526), .B(n4525), .Z(x[146]) );
  NAND U6653 ( .A(init), .B(creg[147]), .Z(n4528) );
  NAND U6654 ( .A(n3866), .B(m[147]), .Z(n4527) );
  NAND U6655 ( .A(n4528), .B(n4527), .Z(x[147]) );
  NAND U6656 ( .A(init), .B(creg[148]), .Z(n4530) );
  NAND U6657 ( .A(n3866), .B(m[148]), .Z(n4529) );
  NAND U6658 ( .A(n4530), .B(n4529), .Z(x[148]) );
  NAND U6659 ( .A(n3867), .B(m[149]), .Z(n4531) );
  NAND U6660 ( .A(init), .B(creg[149]), .Z(n4969) );
  NAND U6661 ( .A(n4531), .B(n4969), .Z(x[149]) );
  NAND U6662 ( .A(n3867), .B(m[14]), .Z(n4532) );
  NAND U6663 ( .A(init), .B(creg[14]), .Z(n4972) );
  NAND U6664 ( .A(n4532), .B(n4972), .Z(x[14]) );
  NAND U6665 ( .A(n3867), .B(m[150]), .Z(n4533) );
  NAND U6666 ( .A(init), .B(creg[150]), .Z(n4975) );
  NAND U6667 ( .A(n4533), .B(n4975), .Z(x[150]) );
  NAND U6668 ( .A(n3867), .B(m[151]), .Z(n4534) );
  NAND U6669 ( .A(init), .B(creg[151]), .Z(n4978) );
  NAND U6670 ( .A(n4534), .B(n4978), .Z(x[151]) );
  NAND U6671 ( .A(init), .B(creg[152]), .Z(n4536) );
  NAND U6672 ( .A(n3867), .B(m[152]), .Z(n4535) );
  NAND U6673 ( .A(n4536), .B(n4535), .Z(x[152]) );
  NAND U6674 ( .A(n3867), .B(m[153]), .Z(n4537) );
  NAND U6675 ( .A(init), .B(creg[153]), .Z(n4983) );
  NAND U6676 ( .A(n4537), .B(n4983), .Z(x[153]) );
  NAND U6677 ( .A(init), .B(creg[154]), .Z(n4539) );
  NAND U6678 ( .A(n3867), .B(m[154]), .Z(n4538) );
  NAND U6679 ( .A(n4539), .B(n4538), .Z(x[154]) );
  NAND U6680 ( .A(n3868), .B(m[155]), .Z(n4540) );
  NAND U6681 ( .A(init), .B(creg[155]), .Z(n4988) );
  NAND U6682 ( .A(n4540), .B(n4988), .Z(x[155]) );
  NAND U6683 ( .A(init), .B(creg[156]), .Z(n4542) );
  NAND U6684 ( .A(n3868), .B(m[156]), .Z(n4541) );
  NAND U6685 ( .A(n4542), .B(n4541), .Z(x[156]) );
  NAND U6686 ( .A(n3868), .B(m[157]), .Z(n4543) );
  NAND U6687 ( .A(init), .B(creg[157]), .Z(n4993) );
  NAND U6688 ( .A(n4543), .B(n4993), .Z(x[157]) );
  NAND U6689 ( .A(init), .B(creg[158]), .Z(n4545) );
  NAND U6690 ( .A(n3868), .B(m[158]), .Z(n4544) );
  NAND U6691 ( .A(n4545), .B(n4544), .Z(x[158]) );
  NAND U6692 ( .A(init), .B(creg[159]), .Z(n4547) );
  NAND U6693 ( .A(n3868), .B(m[159]), .Z(n4546) );
  NAND U6694 ( .A(n4547), .B(n4546), .Z(x[159]) );
  NAND U6695 ( .A(n3868), .B(m[15]), .Z(n4548) );
  NAND U6696 ( .A(init), .B(creg[15]), .Z(n5000) );
  NAND U6697 ( .A(n4548), .B(n5000), .Z(x[15]) );
  NAND U6698 ( .A(n3868), .B(m[160]), .Z(n4549) );
  NAND U6699 ( .A(init), .B(creg[160]), .Z(n5003) );
  NAND U6700 ( .A(n4549), .B(n5003), .Z(x[160]) );
  NAND U6701 ( .A(n3869), .B(m[161]), .Z(n4550) );
  NAND U6702 ( .A(init), .B(creg[161]), .Z(n5006) );
  NAND U6703 ( .A(n4550), .B(n5006), .Z(x[161]) );
  NAND U6704 ( .A(n3869), .B(m[162]), .Z(n4551) );
  NAND U6705 ( .A(init), .B(creg[162]), .Z(n5009) );
  NAND U6706 ( .A(n4551), .B(n5009), .Z(x[162]) );
  NAND U6707 ( .A(init), .B(creg[163]), .Z(n4553) );
  NAND U6708 ( .A(n3869), .B(m[163]), .Z(n4552) );
  NAND U6709 ( .A(n4553), .B(n4552), .Z(x[163]) );
  NAND U6710 ( .A(init), .B(creg[164]), .Z(n4555) );
  NAND U6711 ( .A(n3869), .B(m[164]), .Z(n4554) );
  NAND U6712 ( .A(n4555), .B(n4554), .Z(x[164]) );
  NAND U6713 ( .A(init), .B(creg[165]), .Z(n4557) );
  NAND U6714 ( .A(n3869), .B(m[165]), .Z(n4556) );
  NAND U6715 ( .A(n4557), .B(n4556), .Z(x[165]) );
  NAND U6716 ( .A(n3869), .B(m[166]), .Z(n4558) );
  NAND U6717 ( .A(init), .B(creg[166]), .Z(n5018) );
  NAND U6718 ( .A(n4558), .B(n5018), .Z(x[166]) );
  NAND U6719 ( .A(n3869), .B(m[167]), .Z(n4559) );
  NAND U6720 ( .A(init), .B(creg[167]), .Z(n5021) );
  NAND U6721 ( .A(n4559), .B(n5021), .Z(x[167]) );
  NAND U6722 ( .A(init), .B(creg[168]), .Z(n4561) );
  NAND U6723 ( .A(n3870), .B(m[168]), .Z(n4560) );
  NAND U6724 ( .A(n4561), .B(n4560), .Z(x[168]) );
  NAND U6725 ( .A(n3870), .B(m[169]), .Z(n4562) );
  NAND U6726 ( .A(init), .B(creg[169]), .Z(n5026) );
  NAND U6727 ( .A(n4562), .B(n5026), .Z(x[169]) );
  NAND U6728 ( .A(n3870), .B(m[16]), .Z(n4563) );
  NAND U6729 ( .A(init), .B(creg[16]), .Z(n5029) );
  NAND U6730 ( .A(n4563), .B(n5029), .Z(x[16]) );
  NAND U6731 ( .A(init), .B(creg[170]), .Z(n4565) );
  NAND U6732 ( .A(n3870), .B(m[170]), .Z(n4564) );
  NAND U6733 ( .A(n4565), .B(n4564), .Z(x[170]) );
  NAND U6734 ( .A(init), .B(creg[171]), .Z(n4567) );
  NAND U6735 ( .A(n3870), .B(m[171]), .Z(n4566) );
  NAND U6736 ( .A(n4567), .B(n4566), .Z(x[171]) );
  NAND U6737 ( .A(init), .B(creg[172]), .Z(n4569) );
  NAND U6738 ( .A(n3870), .B(m[172]), .Z(n4568) );
  NAND U6739 ( .A(n4569), .B(n4568), .Z(x[172]) );
  NAND U6740 ( .A(n3870), .B(m[173]), .Z(n4570) );
  NAND U6741 ( .A(init), .B(creg[173]), .Z(n5038) );
  NAND U6742 ( .A(n4570), .B(n5038), .Z(x[173]) );
  NAND U6743 ( .A(n3871), .B(m[174]), .Z(n4571) );
  NAND U6744 ( .A(init), .B(creg[174]), .Z(n5041) );
  NAND U6745 ( .A(n4571), .B(n5041), .Z(x[174]) );
  NAND U6746 ( .A(n3871), .B(m[175]), .Z(n4572) );
  NAND U6747 ( .A(init), .B(creg[175]), .Z(n5044) );
  NAND U6748 ( .A(n4572), .B(n5044), .Z(x[175]) );
  NAND U6749 ( .A(init), .B(creg[176]), .Z(n4574) );
  NAND U6750 ( .A(n3871), .B(m[176]), .Z(n4573) );
  NAND U6751 ( .A(n4574), .B(n4573), .Z(x[176]) );
  NAND U6752 ( .A(init), .B(creg[177]), .Z(n4576) );
  NAND U6753 ( .A(n3871), .B(m[177]), .Z(n4575) );
  NAND U6754 ( .A(n4576), .B(n4575), .Z(x[177]) );
  NAND U6755 ( .A(n3871), .B(m[178]), .Z(n4577) );
  NAND U6756 ( .A(init), .B(creg[178]), .Z(n5051) );
  NAND U6757 ( .A(n4577), .B(n5051), .Z(x[178]) );
  NAND U6758 ( .A(n3871), .B(m[179]), .Z(n4578) );
  NAND U6759 ( .A(init), .B(creg[179]), .Z(n5054) );
  NAND U6760 ( .A(n4578), .B(n5054), .Z(x[179]) );
  NAND U6761 ( .A(init), .B(creg[17]), .Z(n4580) );
  NAND U6762 ( .A(n3871), .B(m[17]), .Z(n4579) );
  NAND U6763 ( .A(n4580), .B(n4579), .Z(x[17]) );
  NAND U6764 ( .A(init), .B(creg[180]), .Z(n4582) );
  NAND U6765 ( .A(n3872), .B(m[180]), .Z(n4581) );
  NAND U6766 ( .A(n4582), .B(n4581), .Z(x[180]) );
  NAND U6767 ( .A(init), .B(creg[181]), .Z(n4584) );
  NAND U6768 ( .A(n3872), .B(m[181]), .Z(n4583) );
  NAND U6769 ( .A(n4584), .B(n4583), .Z(x[181]) );
  NAND U6770 ( .A(n3872), .B(m[182]), .Z(n4585) );
  NAND U6771 ( .A(init), .B(creg[182]), .Z(n5063) );
  NAND U6772 ( .A(n4585), .B(n5063), .Z(x[182]) );
  NAND U6773 ( .A(init), .B(creg[183]), .Z(n4587) );
  NAND U6774 ( .A(n3872), .B(m[183]), .Z(n4586) );
  NAND U6775 ( .A(n4587), .B(n4586), .Z(x[183]) );
  NAND U6776 ( .A(n3872), .B(m[184]), .Z(n4588) );
  NAND U6777 ( .A(init), .B(creg[184]), .Z(n5068) );
  NAND U6778 ( .A(n4588), .B(n5068), .Z(x[184]) );
  NAND U6779 ( .A(init), .B(creg[185]), .Z(n4590) );
  NAND U6780 ( .A(n3872), .B(m[185]), .Z(n4589) );
  NAND U6781 ( .A(n4590), .B(n4589), .Z(x[185]) );
  NAND U6782 ( .A(init), .B(creg[186]), .Z(n4592) );
  NAND U6783 ( .A(n3872), .B(m[186]), .Z(n4591) );
  NAND U6784 ( .A(n4592), .B(n4591), .Z(x[186]) );
  NAND U6785 ( .A(init), .B(creg[187]), .Z(n4594) );
  NAND U6786 ( .A(n3873), .B(m[187]), .Z(n4593) );
  NAND U6787 ( .A(n4594), .B(n4593), .Z(x[187]) );
  NAND U6788 ( .A(init), .B(creg[188]), .Z(n4596) );
  NAND U6789 ( .A(n3873), .B(m[188]), .Z(n4595) );
  NAND U6790 ( .A(n4596), .B(n4595), .Z(x[188]) );
  NAND U6791 ( .A(init), .B(creg[189]), .Z(n4598) );
  NAND U6792 ( .A(n3873), .B(m[189]), .Z(n4597) );
  NAND U6793 ( .A(n4598), .B(n4597), .Z(x[189]) );
  NAND U6794 ( .A(init), .B(creg[18]), .Z(n4600) );
  NAND U6795 ( .A(n3873), .B(m[18]), .Z(n4599) );
  NAND U6796 ( .A(n4600), .B(n4599), .Z(x[18]) );
  NAND U6797 ( .A(n3873), .B(m[190]), .Z(n4601) );
  NAND U6798 ( .A(init), .B(creg[190]), .Z(n5083) );
  NAND U6799 ( .A(n4601), .B(n5083), .Z(x[190]) );
  NAND U6800 ( .A(init), .B(creg[191]), .Z(n4603) );
  NAND U6801 ( .A(n3873), .B(m[191]), .Z(n4602) );
  NAND U6802 ( .A(n4603), .B(n4602), .Z(x[191]) );
  NAND U6803 ( .A(n3873), .B(m[192]), .Z(n4604) );
  NAND U6804 ( .A(init), .B(creg[192]), .Z(n5088) );
  NAND U6805 ( .A(n4604), .B(n5088), .Z(x[192]) );
  NAND U6806 ( .A(init), .B(creg[193]), .Z(n4606) );
  NAND U6807 ( .A(n3874), .B(m[193]), .Z(n4605) );
  NAND U6808 ( .A(n4606), .B(n4605), .Z(x[193]) );
  NAND U6809 ( .A(init), .B(creg[194]), .Z(n4608) );
  NAND U6810 ( .A(n3874), .B(m[194]), .Z(n4607) );
  NAND U6811 ( .A(n4608), .B(n4607), .Z(x[194]) );
  NAND U6812 ( .A(n3874), .B(m[195]), .Z(n4609) );
  NAND U6813 ( .A(init), .B(creg[195]), .Z(n5095) );
  NAND U6814 ( .A(n4609), .B(n5095), .Z(x[195]) );
  NAND U6815 ( .A(init), .B(creg[196]), .Z(n4611) );
  NAND U6816 ( .A(n3874), .B(m[196]), .Z(n4610) );
  NAND U6817 ( .A(n4611), .B(n4610), .Z(x[196]) );
  NAND U6818 ( .A(n3874), .B(m[197]), .Z(n4612) );
  NAND U6819 ( .A(init), .B(creg[197]), .Z(n5100) );
  NAND U6820 ( .A(n4612), .B(n5100), .Z(x[197]) );
  NAND U6821 ( .A(n3874), .B(m[198]), .Z(n4613) );
  NAND U6822 ( .A(init), .B(creg[198]), .Z(n5103) );
  NAND U6823 ( .A(n4613), .B(n5103), .Z(x[198]) );
  NAND U6824 ( .A(n3874), .B(m[199]), .Z(n4614) );
  NAND U6825 ( .A(init), .B(creg[199]), .Z(n5106) );
  NAND U6826 ( .A(n4614), .B(n5106), .Z(x[199]) );
  NAND U6827 ( .A(n3875), .B(m[19]), .Z(n4615) );
  NAND U6828 ( .A(init), .B(creg[19]), .Z(n5109) );
  NAND U6829 ( .A(n4615), .B(n5109), .Z(x[19]) );
  NAND U6830 ( .A(n3875), .B(m[1]), .Z(n4616) );
  NAND U6831 ( .A(init), .B(creg[1]), .Z(n5112) );
  NAND U6832 ( .A(n4616), .B(n5112), .Z(x[1]) );
  NAND U6833 ( .A(init), .B(creg[200]), .Z(n4618) );
  NAND U6834 ( .A(n3875), .B(m[200]), .Z(n4617) );
  NAND U6835 ( .A(n4618), .B(n4617), .Z(x[200]) );
  NAND U6836 ( .A(init), .B(creg[201]), .Z(n4620) );
  NAND U6837 ( .A(n3875), .B(m[201]), .Z(n4619) );
  NAND U6838 ( .A(n4620), .B(n4619), .Z(x[201]) );
  NAND U6839 ( .A(n3875), .B(m[202]), .Z(n4621) );
  NAND U6840 ( .A(init), .B(creg[202]), .Z(n5119) );
  NAND U6841 ( .A(n4621), .B(n5119), .Z(x[202]) );
  NAND U6842 ( .A(n3875), .B(m[203]), .Z(n4622) );
  NAND U6843 ( .A(init), .B(creg[203]), .Z(n5122) );
  NAND U6844 ( .A(n4622), .B(n5122), .Z(x[203]) );
  NAND U6845 ( .A(init), .B(creg[204]), .Z(n4624) );
  NAND U6846 ( .A(n3875), .B(m[204]), .Z(n4623) );
  NAND U6847 ( .A(n4624), .B(n4623), .Z(x[204]) );
  NAND U6848 ( .A(n3876), .B(m[205]), .Z(n4625) );
  NAND U6849 ( .A(init), .B(creg[205]), .Z(n5127) );
  NAND U6850 ( .A(n4625), .B(n5127), .Z(x[205]) );
  NAND U6851 ( .A(n3876), .B(m[206]), .Z(n4626) );
  NAND U6852 ( .A(init), .B(creg[206]), .Z(n5130) );
  NAND U6853 ( .A(n4626), .B(n5130), .Z(x[206]) );
  NAND U6854 ( .A(n3876), .B(m[207]), .Z(n4627) );
  NAND U6855 ( .A(init), .B(creg[207]), .Z(n5133) );
  NAND U6856 ( .A(n4627), .B(n5133), .Z(x[207]) );
  NAND U6857 ( .A(init), .B(creg[208]), .Z(n4629) );
  NAND U6858 ( .A(n3876), .B(m[208]), .Z(n4628) );
  NAND U6859 ( .A(n4629), .B(n4628), .Z(x[208]) );
  NAND U6860 ( .A(n3876), .B(m[209]), .Z(n4630) );
  NAND U6861 ( .A(init), .B(creg[209]), .Z(n5138) );
  NAND U6862 ( .A(n4630), .B(n5138), .Z(x[209]) );
  NAND U6863 ( .A(init), .B(creg[20]), .Z(n4632) );
  NAND U6864 ( .A(n3876), .B(m[20]), .Z(n4631) );
  NAND U6865 ( .A(n4632), .B(n4631), .Z(x[20]) );
  NAND U6866 ( .A(init), .B(creg[210]), .Z(n4634) );
  NAND U6867 ( .A(n3876), .B(m[210]), .Z(n4633) );
  NAND U6868 ( .A(n4634), .B(n4633), .Z(x[210]) );
  NAND U6869 ( .A(init), .B(creg[211]), .Z(n4636) );
  NAND U6870 ( .A(n3877), .B(m[211]), .Z(n4635) );
  NAND U6871 ( .A(n4636), .B(n4635), .Z(x[211]) );
  NAND U6872 ( .A(init), .B(creg[212]), .Z(n4638) );
  NAND U6873 ( .A(n3877), .B(m[212]), .Z(n4637) );
  NAND U6874 ( .A(n4638), .B(n4637), .Z(x[212]) );
  NAND U6875 ( .A(n3877), .B(m[213]), .Z(n4639) );
  NAND U6876 ( .A(init), .B(creg[213]), .Z(n5149) );
  NAND U6877 ( .A(n4639), .B(n5149), .Z(x[213]) );
  NAND U6878 ( .A(init), .B(creg[214]), .Z(n4641) );
  NAND U6879 ( .A(n3877), .B(m[214]), .Z(n4640) );
  NAND U6880 ( .A(n4641), .B(n4640), .Z(x[214]) );
  NAND U6881 ( .A(n3877), .B(m[215]), .Z(n4642) );
  NAND U6882 ( .A(init), .B(creg[215]), .Z(n5154) );
  NAND U6883 ( .A(n4642), .B(n5154), .Z(x[215]) );
  NAND U6884 ( .A(n3877), .B(m[216]), .Z(n4643) );
  NAND U6885 ( .A(init), .B(creg[216]), .Z(n5157) );
  NAND U6886 ( .A(n4643), .B(n5157), .Z(x[216]) );
  NAND U6887 ( .A(init), .B(creg[217]), .Z(n4645) );
  NAND U6888 ( .A(n3877), .B(m[217]), .Z(n4644) );
  NAND U6889 ( .A(n4645), .B(n4644), .Z(x[217]) );
  NAND U6890 ( .A(init), .B(creg[218]), .Z(n4647) );
  NAND U6891 ( .A(n3878), .B(m[218]), .Z(n4646) );
  NAND U6892 ( .A(n4647), .B(n4646), .Z(x[218]) );
  NAND U6893 ( .A(init), .B(creg[219]), .Z(n4649) );
  NAND U6894 ( .A(n3878), .B(m[219]), .Z(n4648) );
  NAND U6895 ( .A(n4649), .B(n4648), .Z(x[219]) );
  NAND U6896 ( .A(init), .B(creg[21]), .Z(n4651) );
  NAND U6897 ( .A(n3878), .B(m[21]), .Z(n4650) );
  NAND U6898 ( .A(n4651), .B(n4650), .Z(x[21]) );
  NAND U6899 ( .A(n3878), .B(m[220]), .Z(n4652) );
  NAND U6900 ( .A(init), .B(creg[220]), .Z(n5168) );
  NAND U6901 ( .A(n4652), .B(n5168), .Z(x[220]) );
  NAND U6902 ( .A(n3878), .B(m[221]), .Z(n4653) );
  NAND U6903 ( .A(init), .B(creg[221]), .Z(n5171) );
  NAND U6904 ( .A(n4653), .B(n5171), .Z(x[221]) );
  NAND U6905 ( .A(init), .B(creg[222]), .Z(n4655) );
  NAND U6906 ( .A(n3878), .B(m[222]), .Z(n4654) );
  NAND U6907 ( .A(n4655), .B(n4654), .Z(x[222]) );
  NAND U6908 ( .A(init), .B(creg[223]), .Z(n4657) );
  NAND U6909 ( .A(n3878), .B(m[223]), .Z(n4656) );
  NAND U6910 ( .A(n4657), .B(n4656), .Z(x[223]) );
  NAND U6911 ( .A(init), .B(creg[224]), .Z(n4659) );
  NAND U6912 ( .A(n3879), .B(m[224]), .Z(n4658) );
  NAND U6913 ( .A(n4659), .B(n4658), .Z(x[224]) );
  NAND U6914 ( .A(init), .B(creg[225]), .Z(n4661) );
  NAND U6915 ( .A(n3879), .B(m[225]), .Z(n4660) );
  NAND U6916 ( .A(n4661), .B(n4660), .Z(x[225]) );
  NAND U6917 ( .A(n3879), .B(m[226]), .Z(n4662) );
  NAND U6918 ( .A(init), .B(creg[226]), .Z(n5182) );
  NAND U6919 ( .A(n4662), .B(n5182), .Z(x[226]) );
  NAND U6920 ( .A(init), .B(creg[227]), .Z(n4664) );
  NAND U6921 ( .A(n3879), .B(m[227]), .Z(n4663) );
  NAND U6922 ( .A(n4664), .B(n4663), .Z(x[227]) );
  NAND U6923 ( .A(init), .B(creg[228]), .Z(n4666) );
  NAND U6924 ( .A(n3879), .B(m[228]), .Z(n4665) );
  NAND U6925 ( .A(n4666), .B(n4665), .Z(x[228]) );
  NAND U6926 ( .A(init), .B(creg[229]), .Z(n4668) );
  NAND U6927 ( .A(n3879), .B(m[229]), .Z(n4667) );
  NAND U6928 ( .A(n4668), .B(n4667), .Z(x[229]) );
  NAND U6929 ( .A(n3879), .B(m[22]), .Z(n4669) );
  NAND U6930 ( .A(init), .B(creg[22]), .Z(n5191) );
  NAND U6931 ( .A(n4669), .B(n5191), .Z(x[22]) );
  NAND U6932 ( .A(init), .B(creg[230]), .Z(n4671) );
  NAND U6933 ( .A(n3880), .B(m[230]), .Z(n4670) );
  NAND U6934 ( .A(n4671), .B(n4670), .Z(x[230]) );
  NAND U6935 ( .A(init), .B(creg[231]), .Z(n4673) );
  NAND U6936 ( .A(n3880), .B(m[231]), .Z(n4672) );
  NAND U6937 ( .A(n4673), .B(n4672), .Z(x[231]) );
  NAND U6938 ( .A(init), .B(creg[232]), .Z(n4675) );
  NAND U6939 ( .A(n3880), .B(m[232]), .Z(n4674) );
  NAND U6940 ( .A(n4675), .B(n4674), .Z(x[232]) );
  NAND U6941 ( .A(init), .B(creg[233]), .Z(n4677) );
  NAND U6942 ( .A(n3880), .B(m[233]), .Z(n4676) );
  NAND U6943 ( .A(n4677), .B(n4676), .Z(x[233]) );
  NAND U6944 ( .A(n3880), .B(m[234]), .Z(n4678) );
  NAND U6945 ( .A(init), .B(creg[234]), .Z(n5202) );
  NAND U6946 ( .A(n4678), .B(n5202), .Z(x[234]) );
  NAND U6947 ( .A(init), .B(creg[235]), .Z(n4680) );
  NAND U6948 ( .A(n3880), .B(m[235]), .Z(n4679) );
  NAND U6949 ( .A(n4680), .B(n4679), .Z(x[235]) );
  NAND U6950 ( .A(init), .B(creg[236]), .Z(n4682) );
  NAND U6951 ( .A(n3880), .B(m[236]), .Z(n4681) );
  NAND U6952 ( .A(n4682), .B(n4681), .Z(x[236]) );
  NAND U6953 ( .A(n3881), .B(m[237]), .Z(n4683) );
  NAND U6954 ( .A(init), .B(creg[237]), .Z(n5209) );
  NAND U6955 ( .A(n4683), .B(n5209), .Z(x[237]) );
  NAND U6956 ( .A(n3881), .B(m[238]), .Z(n4684) );
  NAND U6957 ( .A(init), .B(creg[238]), .Z(n5212) );
  NAND U6958 ( .A(n4684), .B(n5212), .Z(x[238]) );
  NAND U6959 ( .A(init), .B(creg[239]), .Z(n4686) );
  NAND U6960 ( .A(n3881), .B(m[239]), .Z(n4685) );
  NAND U6961 ( .A(n4686), .B(n4685), .Z(x[239]) );
  NAND U6962 ( .A(init), .B(creg[23]), .Z(n4688) );
  NAND U6963 ( .A(n3881), .B(m[23]), .Z(n4687) );
  NAND U6964 ( .A(n4688), .B(n4687), .Z(x[23]) );
  NAND U6965 ( .A(init), .B(creg[240]), .Z(n4690) );
  NAND U6966 ( .A(n3881), .B(m[240]), .Z(n4689) );
  NAND U6967 ( .A(n4690), .B(n4689), .Z(x[240]) );
  NAND U6968 ( .A(n3881), .B(m[241]), .Z(n4691) );
  NAND U6969 ( .A(init), .B(creg[241]), .Z(n5221) );
  NAND U6970 ( .A(n4691), .B(n5221), .Z(x[241]) );
  NAND U6971 ( .A(init), .B(creg[242]), .Z(n4693) );
  NAND U6972 ( .A(n3881), .B(m[242]), .Z(n4692) );
  NAND U6973 ( .A(n4693), .B(n4692), .Z(x[242]) );
  NAND U6974 ( .A(n3882), .B(m[243]), .Z(n4694) );
  NAND U6975 ( .A(init), .B(creg[243]), .Z(n5226) );
  NAND U6976 ( .A(n4694), .B(n5226), .Z(x[243]) );
  NAND U6977 ( .A(n3882), .B(m[244]), .Z(n4695) );
  NAND U6978 ( .A(init), .B(creg[244]), .Z(n5229) );
  NAND U6979 ( .A(n4695), .B(n5229), .Z(x[244]) );
  NAND U6980 ( .A(init), .B(creg[245]), .Z(n4697) );
  NAND U6981 ( .A(n3882), .B(m[245]), .Z(n4696) );
  NAND U6982 ( .A(n4697), .B(n4696), .Z(x[245]) );
  NAND U6983 ( .A(n3882), .B(m[246]), .Z(n4698) );
  NAND U6984 ( .A(init), .B(creg[246]), .Z(n5234) );
  NAND U6985 ( .A(n4698), .B(n5234), .Z(x[246]) );
  NAND U6986 ( .A(init), .B(creg[247]), .Z(n4700) );
  NAND U6987 ( .A(n3882), .B(m[247]), .Z(n4699) );
  NAND U6988 ( .A(n4700), .B(n4699), .Z(x[247]) );
  NAND U6989 ( .A(init), .B(creg[248]), .Z(n4702) );
  NAND U6990 ( .A(n3882), .B(m[248]), .Z(n4701) );
  NAND U6991 ( .A(n4702), .B(n4701), .Z(x[248]) );
  NAND U6992 ( .A(n3882), .B(m[249]), .Z(n4703) );
  NAND U6993 ( .A(init), .B(creg[249]), .Z(n5241) );
  NAND U6994 ( .A(n4703), .B(n5241), .Z(x[249]) );
  NAND U6995 ( .A(init), .B(creg[24]), .Z(n4705) );
  NAND U6996 ( .A(n3883), .B(m[24]), .Z(n4704) );
  NAND U6997 ( .A(n4705), .B(n4704), .Z(x[24]) );
  NAND U6998 ( .A(n3883), .B(m[250]), .Z(n4706) );
  NAND U6999 ( .A(init), .B(creg[250]), .Z(n5246) );
  NAND U7000 ( .A(n4706), .B(n5246), .Z(x[250]) );
  NAND U7001 ( .A(init), .B(creg[251]), .Z(n4708) );
  NAND U7002 ( .A(n3883), .B(m[251]), .Z(n4707) );
  NAND U7003 ( .A(n4708), .B(n4707), .Z(x[251]) );
  NAND U7004 ( .A(init), .B(creg[252]), .Z(n4710) );
  NAND U7005 ( .A(n3883), .B(m[252]), .Z(n4709) );
  NAND U7006 ( .A(n4710), .B(n4709), .Z(x[252]) );
  NAND U7007 ( .A(init), .B(creg[253]), .Z(n4712) );
  NAND U7008 ( .A(n3883), .B(m[253]), .Z(n4711) );
  NAND U7009 ( .A(n4712), .B(n4711), .Z(x[253]) );
  NAND U7010 ( .A(init), .B(creg[254]), .Z(n4714) );
  NAND U7011 ( .A(n3883), .B(m[254]), .Z(n4713) );
  NAND U7012 ( .A(n4714), .B(n4713), .Z(x[254]) );
  NAND U7013 ( .A(init), .B(creg[255]), .Z(n4716) );
  NAND U7014 ( .A(n3883), .B(m[255]), .Z(n4715) );
  NAND U7015 ( .A(n4716), .B(n4715), .Z(x[255]) );
  NAND U7016 ( .A(init), .B(creg[25]), .Z(n4718) );
  NAND U7017 ( .A(n3884), .B(m[25]), .Z(n4717) );
  NAND U7018 ( .A(n4718), .B(n4717), .Z(x[25]) );
  NAND U7019 ( .A(n3884), .B(m[26]), .Z(n4719) );
  NAND U7020 ( .A(init), .B(creg[26]), .Z(n5261) );
  NAND U7021 ( .A(n4719), .B(n5261), .Z(x[26]) );
  NAND U7022 ( .A(n3884), .B(m[27]), .Z(n4720) );
  NAND U7023 ( .A(init), .B(creg[27]), .Z(n5264) );
  NAND U7024 ( .A(n4720), .B(n5264), .Z(x[27]) );
  NAND U7025 ( .A(init), .B(creg[28]), .Z(n4722) );
  NAND U7026 ( .A(n3884), .B(m[28]), .Z(n4721) );
  NAND U7027 ( .A(n4722), .B(n4721), .Z(x[28]) );
  NAND U7028 ( .A(n3884), .B(m[29]), .Z(n4723) );
  NAND U7029 ( .A(init), .B(creg[29]), .Z(n5269) );
  NAND U7030 ( .A(n4723), .B(n5269), .Z(x[29]) );
  NAND U7031 ( .A(n3884), .B(m[2]), .Z(n4724) );
  NAND U7032 ( .A(init), .B(creg[2]), .Z(n5272) );
  NAND U7033 ( .A(n4724), .B(n5272), .Z(x[2]) );
  NAND U7034 ( .A(init), .B(creg[30]), .Z(n4726) );
  NAND U7035 ( .A(n3884), .B(m[30]), .Z(n4725) );
  NAND U7036 ( .A(n4726), .B(n4725), .Z(x[30]) );
  NAND U7037 ( .A(n3885), .B(m[31]), .Z(n4727) );
  NAND U7038 ( .A(init), .B(creg[31]), .Z(n5277) );
  NAND U7039 ( .A(n4727), .B(n5277), .Z(x[31]) );
  NAND U7040 ( .A(n3885), .B(m[32]), .Z(n4728) );
  NAND U7041 ( .A(init), .B(creg[32]), .Z(n5280) );
  NAND U7042 ( .A(n4728), .B(n5280), .Z(x[32]) );
  NAND U7043 ( .A(init), .B(creg[33]), .Z(n4730) );
  NAND U7044 ( .A(n3885), .B(m[33]), .Z(n4729) );
  NAND U7045 ( .A(n4730), .B(n4729), .Z(x[33]) );
  NAND U7046 ( .A(n3885), .B(m[34]), .Z(n4731) );
  NAND U7047 ( .A(init), .B(creg[34]), .Z(n5285) );
  NAND U7048 ( .A(n4731), .B(n5285), .Z(x[34]) );
  NAND U7049 ( .A(init), .B(creg[35]), .Z(n4733) );
  NAND U7050 ( .A(n3885), .B(m[35]), .Z(n4732) );
  NAND U7051 ( .A(n4733), .B(n4732), .Z(x[35]) );
  NAND U7052 ( .A(n3885), .B(m[36]), .Z(n4734) );
  NAND U7053 ( .A(init), .B(creg[36]), .Z(n5290) );
  NAND U7054 ( .A(n4734), .B(n5290), .Z(x[36]) );
  NAND U7055 ( .A(n3885), .B(m[37]), .Z(n4735) );
  NAND U7056 ( .A(init), .B(creg[37]), .Z(n5293) );
  NAND U7057 ( .A(n4735), .B(n5293), .Z(x[37]) );
  NAND U7058 ( .A(init), .B(creg[38]), .Z(n4737) );
  NAND U7059 ( .A(n3886), .B(m[38]), .Z(n4736) );
  NAND U7060 ( .A(n4737), .B(n4736), .Z(x[38]) );
  NAND U7061 ( .A(init), .B(creg[39]), .Z(n4739) );
  NAND U7062 ( .A(n3886), .B(m[39]), .Z(n4738) );
  NAND U7063 ( .A(n4739), .B(n4738), .Z(x[39]) );
  NAND U7064 ( .A(n3886), .B(m[3]), .Z(n4740) );
  NAND U7065 ( .A(init), .B(creg[3]), .Z(n5300) );
  NAND U7066 ( .A(n4740), .B(n5300), .Z(x[3]) );
  NAND U7067 ( .A(init), .B(creg[40]), .Z(n4742) );
  NAND U7068 ( .A(n3886), .B(m[40]), .Z(n4741) );
  NAND U7069 ( .A(n4742), .B(n4741), .Z(x[40]) );
  NAND U7070 ( .A(n3886), .B(m[41]), .Z(n4743) );
  NAND U7071 ( .A(init), .B(creg[41]), .Z(n5305) );
  NAND U7072 ( .A(n4743), .B(n5305), .Z(x[41]) );
  NAND U7073 ( .A(n3886), .B(m[42]), .Z(n4744) );
  NAND U7074 ( .A(init), .B(creg[42]), .Z(n5308) );
  NAND U7075 ( .A(n4744), .B(n5308), .Z(x[42]) );
  NAND U7076 ( .A(init), .B(creg[43]), .Z(n4746) );
  NAND U7077 ( .A(n3886), .B(m[43]), .Z(n4745) );
  NAND U7078 ( .A(n4746), .B(n4745), .Z(x[43]) );
  NAND U7079 ( .A(init), .B(creg[44]), .Z(n4748) );
  NAND U7080 ( .A(n3887), .B(m[44]), .Z(n4747) );
  NAND U7081 ( .A(n4748), .B(n4747), .Z(x[44]) );
  NAND U7082 ( .A(n3887), .B(m[45]), .Z(n4749) );
  NAND U7083 ( .A(init), .B(creg[45]), .Z(n5315) );
  NAND U7084 ( .A(n4749), .B(n5315), .Z(x[45]) );
  NAND U7085 ( .A(init), .B(creg[46]), .Z(n4751) );
  NAND U7086 ( .A(n3887), .B(m[46]), .Z(n4750) );
  NAND U7087 ( .A(n4751), .B(n4750), .Z(x[46]) );
  NAND U7088 ( .A(n3887), .B(m[47]), .Z(n4752) );
  NAND U7089 ( .A(init), .B(creg[47]), .Z(n5320) );
  NAND U7090 ( .A(n4752), .B(n5320), .Z(x[47]) );
  NAND U7091 ( .A(init), .B(creg[48]), .Z(n4754) );
  NAND U7092 ( .A(n3887), .B(m[48]), .Z(n4753) );
  NAND U7093 ( .A(n4754), .B(n4753), .Z(x[48]) );
  NAND U7094 ( .A(n3887), .B(m[49]), .Z(n4755) );
  NAND U7095 ( .A(init), .B(creg[49]), .Z(n5325) );
  NAND U7096 ( .A(n4755), .B(n5325), .Z(x[49]) );
  NAND U7097 ( .A(n3887), .B(m[4]), .Z(n4756) );
  NAND U7098 ( .A(init), .B(creg[4]), .Z(n5328) );
  NAND U7099 ( .A(n4756), .B(n5328), .Z(x[4]) );
  NAND U7100 ( .A(init), .B(creg[50]), .Z(n4758) );
  NAND U7101 ( .A(n3888), .B(m[50]), .Z(n4757) );
  NAND U7102 ( .A(n4758), .B(n4757), .Z(x[50]) );
  NAND U7103 ( .A(n3888), .B(m[51]), .Z(n4759) );
  NAND U7104 ( .A(init), .B(creg[51]), .Z(n5333) );
  NAND U7105 ( .A(n4759), .B(n5333), .Z(x[51]) );
  NAND U7106 ( .A(init), .B(creg[52]), .Z(n4761) );
  NAND U7107 ( .A(n3888), .B(m[52]), .Z(n4760) );
  NAND U7108 ( .A(n4761), .B(n4760), .Z(x[52]) );
  NAND U7109 ( .A(init), .B(creg[53]), .Z(n4763) );
  NAND U7110 ( .A(n3888), .B(m[53]), .Z(n4762) );
  NAND U7111 ( .A(n4763), .B(n4762), .Z(x[53]) );
  NAND U7112 ( .A(n3888), .B(m[54]), .Z(n4764) );
  NAND U7113 ( .A(init), .B(creg[54]), .Z(n5340) );
  NAND U7114 ( .A(n4764), .B(n5340), .Z(x[54]) );
  NAND U7115 ( .A(n3888), .B(m[55]), .Z(n4765) );
  NAND U7116 ( .A(init), .B(creg[55]), .Z(n5343) );
  NAND U7117 ( .A(n4765), .B(n5343), .Z(x[55]) );
  NAND U7118 ( .A(n3888), .B(m[56]), .Z(n4766) );
  NAND U7119 ( .A(init), .B(creg[56]), .Z(n5346) );
  NAND U7120 ( .A(n4766), .B(n5346), .Z(x[56]) );
  NAND U7121 ( .A(init), .B(creg[57]), .Z(n4768) );
  NAND U7122 ( .A(n3889), .B(m[57]), .Z(n4767) );
  NAND U7123 ( .A(n4768), .B(n4767), .Z(x[57]) );
  NAND U7124 ( .A(n3889), .B(m[58]), .Z(n4769) );
  NAND U7125 ( .A(init), .B(creg[58]), .Z(n5351) );
  NAND U7126 ( .A(n4769), .B(n5351), .Z(x[58]) );
  NAND U7127 ( .A(init), .B(creg[59]), .Z(n4771) );
  NAND U7128 ( .A(n3889), .B(m[59]), .Z(n4770) );
  NAND U7129 ( .A(n4771), .B(n4770), .Z(x[59]) );
  NAND U7130 ( .A(init), .B(creg[5]), .Z(n4773) );
  NAND U7131 ( .A(n3889), .B(m[5]), .Z(n4772) );
  NAND U7132 ( .A(n4773), .B(n4772), .Z(x[5]) );
  NAND U7133 ( .A(n3889), .B(m[60]), .Z(n4774) );
  NAND U7134 ( .A(init), .B(creg[60]), .Z(n5358) );
  NAND U7135 ( .A(n4774), .B(n5358), .Z(x[60]) );
  NAND U7136 ( .A(init), .B(creg[61]), .Z(n4776) );
  NAND U7137 ( .A(n3889), .B(m[61]), .Z(n4775) );
  NAND U7138 ( .A(n4776), .B(n4775), .Z(x[61]) );
  NAND U7139 ( .A(n3889), .B(m[62]), .Z(n4777) );
  NAND U7140 ( .A(init), .B(creg[62]), .Z(n5363) );
  NAND U7141 ( .A(n4777), .B(n5363), .Z(x[62]) );
  NAND U7142 ( .A(init), .B(creg[63]), .Z(n4779) );
  NAND U7143 ( .A(n3890), .B(m[63]), .Z(n4778) );
  NAND U7144 ( .A(n4779), .B(n4778), .Z(x[63]) );
  NAND U7145 ( .A(init), .B(creg[64]), .Z(n4781) );
  NAND U7146 ( .A(n3890), .B(m[64]), .Z(n4780) );
  NAND U7147 ( .A(n4781), .B(n4780), .Z(x[64]) );
  NAND U7148 ( .A(init), .B(creg[65]), .Z(n4783) );
  NAND U7149 ( .A(n3890), .B(m[65]), .Z(n4782) );
  NAND U7150 ( .A(n4783), .B(n4782), .Z(x[65]) );
  NAND U7151 ( .A(n3890), .B(m[66]), .Z(n4784) );
  NAND U7152 ( .A(init), .B(creg[66]), .Z(n5372) );
  NAND U7153 ( .A(n4784), .B(n5372), .Z(x[66]) );
  NAND U7154 ( .A(init), .B(creg[67]), .Z(n4786) );
  NAND U7155 ( .A(n3890), .B(m[67]), .Z(n4785) );
  NAND U7156 ( .A(n4786), .B(n4785), .Z(x[67]) );
  NAND U7157 ( .A(n3890), .B(m[68]), .Z(n4787) );
  NAND U7158 ( .A(init), .B(creg[68]), .Z(n5377) );
  NAND U7159 ( .A(n4787), .B(n5377), .Z(x[68]) );
  NAND U7160 ( .A(init), .B(creg[69]), .Z(n4789) );
  NAND U7161 ( .A(n3890), .B(m[69]), .Z(n4788) );
  NAND U7162 ( .A(n4789), .B(n4788), .Z(x[69]) );
  NAND U7163 ( .A(init), .B(creg[6]), .Z(n4791) );
  NAND U7164 ( .A(n3891), .B(m[6]), .Z(n4790) );
  NAND U7165 ( .A(n4791), .B(n4790), .Z(x[6]) );
  NAND U7166 ( .A(n3891), .B(m[70]), .Z(n4792) );
  NAND U7167 ( .A(init), .B(creg[70]), .Z(n5384) );
  NAND U7168 ( .A(n4792), .B(n5384), .Z(x[70]) );
  NAND U7169 ( .A(init), .B(creg[71]), .Z(n4794) );
  NAND U7170 ( .A(n3891), .B(m[71]), .Z(n4793) );
  NAND U7171 ( .A(n4794), .B(n4793), .Z(x[71]) );
  NAND U7172 ( .A(n3891), .B(m[72]), .Z(n4795) );
  NAND U7173 ( .A(init), .B(creg[72]), .Z(n5389) );
  NAND U7174 ( .A(n4795), .B(n5389), .Z(x[72]) );
  NAND U7175 ( .A(init), .B(creg[73]), .Z(n4797) );
  NAND U7176 ( .A(n3891), .B(m[73]), .Z(n4796) );
  NAND U7177 ( .A(n4797), .B(n4796), .Z(x[73]) );
  NAND U7178 ( .A(n3891), .B(m[74]), .Z(n4798) );
  NAND U7179 ( .A(init), .B(creg[74]), .Z(n5394) );
  NAND U7180 ( .A(n4798), .B(n5394), .Z(x[74]) );
  NAND U7181 ( .A(n3891), .B(m[75]), .Z(n4799) );
  NAND U7182 ( .A(init), .B(creg[75]), .Z(n5397) );
  NAND U7183 ( .A(n4799), .B(n5397), .Z(x[75]) );
  NAND U7184 ( .A(n3892), .B(m[76]), .Z(n4800) );
  NAND U7185 ( .A(init), .B(creg[76]), .Z(n5400) );
  NAND U7186 ( .A(n4800), .B(n5400), .Z(x[76]) );
  NAND U7187 ( .A(n3892), .B(m[77]), .Z(n4801) );
  NAND U7188 ( .A(init), .B(creg[77]), .Z(n5403) );
  NAND U7189 ( .A(n4801), .B(n5403), .Z(x[77]) );
  NAND U7190 ( .A(init), .B(creg[78]), .Z(n4803) );
  NAND U7191 ( .A(n3892), .B(m[78]), .Z(n4802) );
  NAND U7192 ( .A(n4803), .B(n4802), .Z(x[78]) );
  NAND U7193 ( .A(init), .B(creg[79]), .Z(n4805) );
  NAND U7194 ( .A(n3892), .B(m[79]), .Z(n4804) );
  NAND U7195 ( .A(n4805), .B(n4804), .Z(x[79]) );
  NAND U7196 ( .A(init), .B(creg[7]), .Z(n4807) );
  NAND U7197 ( .A(n3892), .B(m[7]), .Z(n4806) );
  NAND U7198 ( .A(n4807), .B(n4806), .Z(x[7]) );
  NAND U7199 ( .A(n3892), .B(m[80]), .Z(n4808) );
  NAND U7200 ( .A(init), .B(creg[80]), .Z(n5412) );
  NAND U7201 ( .A(n4808), .B(n5412), .Z(x[80]) );
  NAND U7202 ( .A(n3892), .B(m[81]), .Z(n4809) );
  NAND U7203 ( .A(init), .B(creg[81]), .Z(n5415) );
  NAND U7204 ( .A(n4809), .B(n5415), .Z(x[81]) );
  NAND U7205 ( .A(n3893), .B(m[82]), .Z(n4810) );
  NAND U7206 ( .A(init), .B(creg[82]), .Z(n5418) );
  NAND U7207 ( .A(n4810), .B(n5418), .Z(x[82]) );
  NAND U7208 ( .A(n3893), .B(m[83]), .Z(n4811) );
  NAND U7209 ( .A(init), .B(creg[83]), .Z(n5421) );
  NAND U7210 ( .A(n4811), .B(n5421), .Z(x[83]) );
  NAND U7211 ( .A(init), .B(creg[84]), .Z(n4813) );
  NAND U7212 ( .A(n3893), .B(m[84]), .Z(n4812) );
  NAND U7213 ( .A(n4813), .B(n4812), .Z(x[84]) );
  NAND U7214 ( .A(n3893), .B(m[85]), .Z(n4814) );
  NAND U7215 ( .A(init), .B(creg[85]), .Z(n5426) );
  NAND U7216 ( .A(n4814), .B(n5426), .Z(x[85]) );
  NAND U7217 ( .A(n3893), .B(m[86]), .Z(n4815) );
  NAND U7218 ( .A(init), .B(creg[86]), .Z(n5429) );
  NAND U7219 ( .A(n4815), .B(n5429), .Z(x[86]) );
  NAND U7220 ( .A(init), .B(creg[87]), .Z(n4817) );
  NAND U7221 ( .A(n3893), .B(m[87]), .Z(n4816) );
  NAND U7222 ( .A(n4817), .B(n4816), .Z(x[87]) );
  NAND U7223 ( .A(init), .B(creg[88]), .Z(n4819) );
  NAND U7224 ( .A(n3893), .B(m[88]), .Z(n4818) );
  NAND U7225 ( .A(n4819), .B(n4818), .Z(x[88]) );
  NAND U7226 ( .A(init), .B(creg[89]), .Z(n4821) );
  NAND U7227 ( .A(n3894), .B(m[89]), .Z(n4820) );
  NAND U7228 ( .A(n4821), .B(n4820), .Z(x[89]) );
  NAND U7229 ( .A(init), .B(creg[8]), .Z(n4823) );
  NAND U7230 ( .A(n3894), .B(m[8]), .Z(n4822) );
  NAND U7231 ( .A(n4823), .B(n4822), .Z(x[8]) );
  NAND U7232 ( .A(n3894), .B(m[90]), .Z(n4824) );
  NAND U7233 ( .A(init), .B(creg[90]), .Z(n5440) );
  NAND U7234 ( .A(n4824), .B(n5440), .Z(x[90]) );
  NAND U7235 ( .A(n3894), .B(m[91]), .Z(n4825) );
  NAND U7236 ( .A(init), .B(creg[91]), .Z(n5443) );
  NAND U7237 ( .A(n4825), .B(n5443), .Z(x[91]) );
  NAND U7238 ( .A(n3894), .B(m[92]), .Z(n4826) );
  NAND U7239 ( .A(init), .B(creg[92]), .Z(n5446) );
  NAND U7240 ( .A(n4826), .B(n5446), .Z(x[92]) );
  NAND U7241 ( .A(init), .B(creg[93]), .Z(n4828) );
  NAND U7242 ( .A(n3894), .B(m[93]), .Z(n4827) );
  NAND U7243 ( .A(n4828), .B(n4827), .Z(x[93]) );
  NAND U7244 ( .A(n3894), .B(m[94]), .Z(n4829) );
  NAND U7245 ( .A(init), .B(creg[94]), .Z(n5451) );
  NAND U7246 ( .A(n4829), .B(n5451), .Z(x[94]) );
  NAND U7247 ( .A(n3895), .B(m[95]), .Z(n4830) );
  NAND U7248 ( .A(init), .B(creg[95]), .Z(n5454) );
  NAND U7249 ( .A(n4830), .B(n5454), .Z(x[95]) );
  NAND U7250 ( .A(n3895), .B(m[96]), .Z(n4831) );
  NAND U7251 ( .A(init), .B(creg[96]), .Z(n5457) );
  NAND U7252 ( .A(n4831), .B(n5457), .Z(x[96]) );
  NAND U7253 ( .A(n3895), .B(m[97]), .Z(n4832) );
  NAND U7254 ( .A(init), .B(creg[97]), .Z(n5460) );
  NAND U7255 ( .A(n4832), .B(n5460), .Z(x[97]) );
  NAND U7256 ( .A(n3895), .B(m[98]), .Z(n4833) );
  NAND U7257 ( .A(init), .B(creg[98]), .Z(n5463) );
  NAND U7258 ( .A(n4833), .B(n5463), .Z(x[98]) );
  NAND U7259 ( .A(init), .B(creg[99]), .Z(n4835) );
  NAND U7260 ( .A(n3895), .B(m[99]), .Z(n4834) );
  NAND U7261 ( .A(n4835), .B(n4834), .Z(x[99]) );
  NAND U7262 ( .A(init), .B(creg[9]), .Z(n4837) );
  NAND U7263 ( .A(n3895), .B(m[9]), .Z(n4836) );
  NAND U7264 ( .A(n4837), .B(n4836), .Z(x[9]) );
  IV U7265 ( .A(mul_pow), .Z(n5986) );
  NANDN U7266 ( .A(n4838), .B(n5986), .Z(n4840) );
  NAND U7267 ( .A(init), .B(n5986), .Z(n5468) );
  NAND U7268 ( .A(n5468), .B(m[0]), .Z(n4839) );
  NAND U7269 ( .A(n4840), .B(n4839), .Z(y[0]) );
  NANDN U7270 ( .A(n4841), .B(n5986), .Z(n4843) );
  NAND U7271 ( .A(n5468), .B(m[100]), .Z(n4842) );
  NAND U7272 ( .A(n4843), .B(n4842), .Z(y[100]) );
  NANDN U7273 ( .A(n4844), .B(n5986), .Z(n4846) );
  NAND U7274 ( .A(n5468), .B(m[101]), .Z(n4845) );
  NAND U7275 ( .A(n4846), .B(n4845), .Z(y[101]) );
  NANDN U7276 ( .A(n4847), .B(n5986), .Z(n4849) );
  NAND U7277 ( .A(n5468), .B(m[102]), .Z(n4848) );
  NAND U7278 ( .A(n4849), .B(n4848), .Z(y[102]) );
  NANDN U7279 ( .A(n4850), .B(n5986), .Z(n4852) );
  NAND U7280 ( .A(n5468), .B(m[103]), .Z(n4851) );
  NAND U7281 ( .A(n4852), .B(n4851), .Z(y[103]) );
  NANDN U7282 ( .A(n4853), .B(n5986), .Z(n4855) );
  NAND U7283 ( .A(n5468), .B(m[104]), .Z(n4854) );
  NAND U7284 ( .A(n4855), .B(n4854), .Z(y[104]) );
  NAND U7285 ( .A(n5468), .B(m[105]), .Z(n4857) );
  NANDN U7286 ( .A(n5468), .B(creg[105]), .Z(n4856) );
  NAND U7287 ( .A(n4857), .B(n4856), .Z(y[105]) );
  NAND U7288 ( .A(n5468), .B(m[106]), .Z(n4859) );
  NANDN U7289 ( .A(n5468), .B(creg[106]), .Z(n4858) );
  NAND U7290 ( .A(n4859), .B(n4858), .Z(y[106]) );
  NAND U7291 ( .A(n5468), .B(m[107]), .Z(n4861) );
  NANDN U7292 ( .A(n5468), .B(creg[107]), .Z(n4860) );
  NAND U7293 ( .A(n4861), .B(n4860), .Z(y[107]) );
  NANDN U7294 ( .A(n4862), .B(n5986), .Z(n4864) );
  NAND U7295 ( .A(n5468), .B(m[108]), .Z(n4863) );
  NAND U7296 ( .A(n4864), .B(n4863), .Z(y[108]) );
  NANDN U7297 ( .A(n4865), .B(n5986), .Z(n4867) );
  NAND U7298 ( .A(n5468), .B(m[109]), .Z(n4866) );
  NAND U7299 ( .A(n4867), .B(n4866), .Z(y[109]) );
  NANDN U7300 ( .A(n4868), .B(n5986), .Z(n4870) );
  NAND U7301 ( .A(n5468), .B(m[10]), .Z(n4869) );
  NAND U7302 ( .A(n4870), .B(n4869), .Z(y[10]) );
  NAND U7303 ( .A(n5468), .B(m[110]), .Z(n4872) );
  NANDN U7304 ( .A(n5468), .B(creg[110]), .Z(n4871) );
  NAND U7305 ( .A(n4872), .B(n4871), .Z(y[110]) );
  NAND U7306 ( .A(n5468), .B(m[111]), .Z(n4874) );
  NANDN U7307 ( .A(n5468), .B(creg[111]), .Z(n4873) );
  NAND U7308 ( .A(n4874), .B(n4873), .Z(y[111]) );
  NAND U7309 ( .A(n5468), .B(m[112]), .Z(n4876) );
  NANDN U7310 ( .A(n5468), .B(creg[112]), .Z(n4875) );
  NAND U7311 ( .A(n4876), .B(n4875), .Z(y[112]) );
  NANDN U7312 ( .A(n4877), .B(n5986), .Z(n4879) );
  NAND U7313 ( .A(n5468), .B(m[113]), .Z(n4878) );
  NAND U7314 ( .A(n4879), .B(n4878), .Z(y[113]) );
  NAND U7315 ( .A(n5468), .B(m[114]), .Z(n4881) );
  NANDN U7316 ( .A(n5468), .B(creg[114]), .Z(n4880) );
  NAND U7317 ( .A(n4881), .B(n4880), .Z(y[114]) );
  NAND U7318 ( .A(n5468), .B(m[115]), .Z(n4883) );
  NANDN U7319 ( .A(n5468), .B(creg[115]), .Z(n4882) );
  NAND U7320 ( .A(n4883), .B(n4882), .Z(y[115]) );
  NANDN U7321 ( .A(n4884), .B(n5986), .Z(n4886) );
  NAND U7322 ( .A(n5468), .B(m[116]), .Z(n4885) );
  NAND U7323 ( .A(n4886), .B(n4885), .Z(y[116]) );
  NANDN U7324 ( .A(n4887), .B(n5986), .Z(n4889) );
  NAND U7325 ( .A(n5468), .B(m[117]), .Z(n4888) );
  NAND U7326 ( .A(n4889), .B(n4888), .Z(y[117]) );
  NANDN U7327 ( .A(n4890), .B(n5986), .Z(n4892) );
  NAND U7328 ( .A(n5468), .B(m[118]), .Z(n4891) );
  NAND U7329 ( .A(n4892), .B(n4891), .Z(y[118]) );
  NANDN U7330 ( .A(n4893), .B(n5986), .Z(n4895) );
  NAND U7331 ( .A(n5468), .B(m[119]), .Z(n4894) );
  NAND U7332 ( .A(n4895), .B(n4894), .Z(y[119]) );
  NANDN U7333 ( .A(n4896), .B(n5986), .Z(n4898) );
  NAND U7334 ( .A(n5468), .B(m[11]), .Z(n4897) );
  NAND U7335 ( .A(n4898), .B(n4897), .Z(y[11]) );
  NAND U7336 ( .A(n5468), .B(m[120]), .Z(n4900) );
  NANDN U7337 ( .A(n5468), .B(creg[120]), .Z(n4899) );
  NAND U7338 ( .A(n4900), .B(n4899), .Z(y[120]) );
  NAND U7339 ( .A(n5468), .B(m[121]), .Z(n4902) );
  NANDN U7340 ( .A(n5468), .B(creg[121]), .Z(n4901) );
  NAND U7341 ( .A(n4902), .B(n4901), .Z(y[121]) );
  NANDN U7342 ( .A(n4903), .B(n5986), .Z(n4905) );
  NAND U7343 ( .A(n5468), .B(m[122]), .Z(n4904) );
  NAND U7344 ( .A(n4905), .B(n4904), .Z(y[122]) );
  NAND U7345 ( .A(n5468), .B(m[123]), .Z(n4907) );
  NANDN U7346 ( .A(n5468), .B(creg[123]), .Z(n4906) );
  NAND U7347 ( .A(n4907), .B(n4906), .Z(y[123]) );
  NAND U7348 ( .A(n5468), .B(m[124]), .Z(n4909) );
  NANDN U7349 ( .A(n5468), .B(creg[124]), .Z(n4908) );
  NAND U7350 ( .A(n4909), .B(n4908), .Z(y[124]) );
  NANDN U7351 ( .A(n4910), .B(n5986), .Z(n4912) );
  NAND U7352 ( .A(n5468), .B(m[125]), .Z(n4911) );
  NAND U7353 ( .A(n4912), .B(n4911), .Z(y[125]) );
  NAND U7354 ( .A(n5468), .B(m[126]), .Z(n4914) );
  NANDN U7355 ( .A(n5468), .B(creg[126]), .Z(n4913) );
  NAND U7356 ( .A(n4914), .B(n4913), .Z(y[126]) );
  NAND U7357 ( .A(n5468), .B(m[127]), .Z(n4916) );
  NANDN U7358 ( .A(n5468), .B(creg[127]), .Z(n4915) );
  NAND U7359 ( .A(n4916), .B(n4915), .Z(y[127]) );
  NAND U7360 ( .A(n5468), .B(m[128]), .Z(n4918) );
  NANDN U7361 ( .A(n5468), .B(creg[128]), .Z(n4917) );
  NAND U7362 ( .A(n4918), .B(n4917), .Z(y[128]) );
  NAND U7363 ( .A(n5468), .B(m[129]), .Z(n4920) );
  NANDN U7364 ( .A(n5468), .B(creg[129]), .Z(n4919) );
  NAND U7365 ( .A(n4920), .B(n4919), .Z(y[129]) );
  NANDN U7366 ( .A(n4921), .B(n5986), .Z(n4923) );
  NAND U7367 ( .A(n5468), .B(m[12]), .Z(n4922) );
  NAND U7368 ( .A(n4923), .B(n4922), .Z(y[12]) );
  NAND U7369 ( .A(n5468), .B(m[130]), .Z(n4925) );
  NANDN U7370 ( .A(n5468), .B(creg[130]), .Z(n4924) );
  NAND U7371 ( .A(n4925), .B(n4924), .Z(y[130]) );
  NAND U7372 ( .A(n5468), .B(m[131]), .Z(n4927) );
  NANDN U7373 ( .A(n5468), .B(creg[131]), .Z(n4926) );
  NAND U7374 ( .A(n4927), .B(n4926), .Z(y[131]) );
  NAND U7375 ( .A(n5468), .B(m[132]), .Z(n4929) );
  NANDN U7376 ( .A(n5468), .B(creg[132]), .Z(n4928) );
  NAND U7377 ( .A(n4929), .B(n4928), .Z(y[132]) );
  NANDN U7378 ( .A(n4930), .B(n5986), .Z(n4932) );
  NAND U7379 ( .A(n5468), .B(m[133]), .Z(n4931) );
  NAND U7380 ( .A(n4932), .B(n4931), .Z(y[133]) );
  NAND U7381 ( .A(n5468), .B(m[134]), .Z(n4934) );
  NANDN U7382 ( .A(n5468), .B(creg[134]), .Z(n4933) );
  NAND U7383 ( .A(n4934), .B(n4933), .Z(y[134]) );
  NAND U7384 ( .A(n5468), .B(m[135]), .Z(n4936) );
  NANDN U7385 ( .A(n5468), .B(creg[135]), .Z(n4935) );
  NAND U7386 ( .A(n4936), .B(n4935), .Z(y[135]) );
  NAND U7387 ( .A(n5468), .B(m[136]), .Z(n4938) );
  NANDN U7388 ( .A(n5468), .B(creg[136]), .Z(n4937) );
  NAND U7389 ( .A(n4938), .B(n4937), .Z(y[136]) );
  NANDN U7390 ( .A(n4939), .B(n5986), .Z(n4941) );
  NAND U7391 ( .A(n5468), .B(m[137]), .Z(n4940) );
  NAND U7392 ( .A(n4941), .B(n4940), .Z(y[137]) );
  NANDN U7393 ( .A(n4942), .B(n5986), .Z(n4944) );
  NAND U7394 ( .A(n5468), .B(m[138]), .Z(n4943) );
  NAND U7395 ( .A(n4944), .B(n4943), .Z(y[138]) );
  NAND U7396 ( .A(n5468), .B(m[139]), .Z(n4946) );
  NANDN U7397 ( .A(n5468), .B(creg[139]), .Z(n4945) );
  NAND U7398 ( .A(n4946), .B(n4945), .Z(y[139]) );
  NAND U7399 ( .A(n5468), .B(m[13]), .Z(n4948) );
  NANDN U7400 ( .A(n5468), .B(creg[13]), .Z(n4947) );
  NAND U7401 ( .A(n4948), .B(n4947), .Z(y[13]) );
  NANDN U7402 ( .A(n4949), .B(n5986), .Z(n4951) );
  NAND U7403 ( .A(n5468), .B(m[140]), .Z(n4950) );
  NAND U7404 ( .A(n4951), .B(n4950), .Z(y[140]) );
  NANDN U7405 ( .A(n4952), .B(n5986), .Z(n4954) );
  NAND U7406 ( .A(n5468), .B(m[141]), .Z(n4953) );
  NAND U7407 ( .A(n4954), .B(n4953), .Z(y[141]) );
  NAND U7408 ( .A(n5468), .B(m[142]), .Z(n4956) );
  NANDN U7409 ( .A(n5468), .B(creg[142]), .Z(n4955) );
  NAND U7410 ( .A(n4956), .B(n4955), .Z(y[142]) );
  NAND U7411 ( .A(n5468), .B(m[143]), .Z(n4958) );
  NANDN U7412 ( .A(n5468), .B(creg[143]), .Z(n4957) );
  NAND U7413 ( .A(n4958), .B(n4957), .Z(y[143]) );
  NAND U7414 ( .A(n5468), .B(m[144]), .Z(n4960) );
  NANDN U7415 ( .A(n5468), .B(creg[144]), .Z(n4959) );
  NAND U7416 ( .A(n4960), .B(n4959), .Z(y[144]) );
  NAND U7417 ( .A(n5468), .B(m[145]), .Z(n4962) );
  NANDN U7418 ( .A(n5468), .B(creg[145]), .Z(n4961) );
  NAND U7419 ( .A(n4962), .B(n4961), .Z(y[145]) );
  NAND U7420 ( .A(n5468), .B(m[146]), .Z(n4964) );
  NANDN U7421 ( .A(n5468), .B(creg[146]), .Z(n4963) );
  NAND U7422 ( .A(n4964), .B(n4963), .Z(y[146]) );
  NAND U7423 ( .A(n5468), .B(m[147]), .Z(n4966) );
  NANDN U7424 ( .A(n5468), .B(creg[147]), .Z(n4965) );
  NAND U7425 ( .A(n4966), .B(n4965), .Z(y[147]) );
  NAND U7426 ( .A(n5468), .B(m[148]), .Z(n4968) );
  NANDN U7427 ( .A(n5468), .B(creg[148]), .Z(n4967) );
  NAND U7428 ( .A(n4968), .B(n4967), .Z(y[148]) );
  NANDN U7429 ( .A(n4969), .B(n5986), .Z(n4971) );
  NAND U7430 ( .A(n5468), .B(m[149]), .Z(n4970) );
  NAND U7431 ( .A(n4971), .B(n4970), .Z(y[149]) );
  NANDN U7432 ( .A(n4972), .B(n5986), .Z(n4974) );
  NAND U7433 ( .A(n5468), .B(m[14]), .Z(n4973) );
  NAND U7434 ( .A(n4974), .B(n4973), .Z(y[14]) );
  NANDN U7435 ( .A(n4975), .B(n5986), .Z(n4977) );
  NAND U7436 ( .A(n5468), .B(m[150]), .Z(n4976) );
  NAND U7437 ( .A(n4977), .B(n4976), .Z(y[150]) );
  NANDN U7438 ( .A(n4978), .B(n5986), .Z(n4980) );
  NAND U7439 ( .A(n5468), .B(m[151]), .Z(n4979) );
  NAND U7440 ( .A(n4980), .B(n4979), .Z(y[151]) );
  NAND U7441 ( .A(n5468), .B(m[152]), .Z(n4982) );
  NANDN U7442 ( .A(n5468), .B(creg[152]), .Z(n4981) );
  NAND U7443 ( .A(n4982), .B(n4981), .Z(y[152]) );
  NANDN U7444 ( .A(n4983), .B(n5986), .Z(n4985) );
  NAND U7445 ( .A(n5468), .B(m[153]), .Z(n4984) );
  NAND U7446 ( .A(n4985), .B(n4984), .Z(y[153]) );
  NAND U7447 ( .A(n5468), .B(m[154]), .Z(n4987) );
  NANDN U7448 ( .A(n5468), .B(creg[154]), .Z(n4986) );
  NAND U7449 ( .A(n4987), .B(n4986), .Z(y[154]) );
  NANDN U7450 ( .A(n4988), .B(n5986), .Z(n4990) );
  NAND U7451 ( .A(n5468), .B(m[155]), .Z(n4989) );
  NAND U7452 ( .A(n4990), .B(n4989), .Z(y[155]) );
  NAND U7453 ( .A(n5468), .B(m[156]), .Z(n4992) );
  NANDN U7454 ( .A(n5468), .B(creg[156]), .Z(n4991) );
  NAND U7455 ( .A(n4992), .B(n4991), .Z(y[156]) );
  NANDN U7456 ( .A(n4993), .B(n5986), .Z(n4995) );
  NAND U7457 ( .A(n5468), .B(m[157]), .Z(n4994) );
  NAND U7458 ( .A(n4995), .B(n4994), .Z(y[157]) );
  NAND U7459 ( .A(n5468), .B(m[158]), .Z(n4997) );
  NANDN U7460 ( .A(n5468), .B(creg[158]), .Z(n4996) );
  NAND U7461 ( .A(n4997), .B(n4996), .Z(y[158]) );
  NAND U7462 ( .A(n5468), .B(m[159]), .Z(n4999) );
  NANDN U7463 ( .A(n5468), .B(creg[159]), .Z(n4998) );
  NAND U7464 ( .A(n4999), .B(n4998), .Z(y[159]) );
  NANDN U7465 ( .A(n5000), .B(n5986), .Z(n5002) );
  NAND U7466 ( .A(n5468), .B(m[15]), .Z(n5001) );
  NAND U7467 ( .A(n5002), .B(n5001), .Z(y[15]) );
  NANDN U7468 ( .A(n5003), .B(n5986), .Z(n5005) );
  NAND U7469 ( .A(n5468), .B(m[160]), .Z(n5004) );
  NAND U7470 ( .A(n5005), .B(n5004), .Z(y[160]) );
  NANDN U7471 ( .A(n5006), .B(n5986), .Z(n5008) );
  NAND U7472 ( .A(n5468), .B(m[161]), .Z(n5007) );
  NAND U7473 ( .A(n5008), .B(n5007), .Z(y[161]) );
  NANDN U7474 ( .A(n5009), .B(n5986), .Z(n5011) );
  NAND U7475 ( .A(n5468), .B(m[162]), .Z(n5010) );
  NAND U7476 ( .A(n5011), .B(n5010), .Z(y[162]) );
  NAND U7477 ( .A(n5468), .B(m[163]), .Z(n5013) );
  NANDN U7478 ( .A(n5468), .B(creg[163]), .Z(n5012) );
  NAND U7479 ( .A(n5013), .B(n5012), .Z(y[163]) );
  NAND U7480 ( .A(n5468), .B(m[164]), .Z(n5015) );
  NANDN U7481 ( .A(n5468), .B(creg[164]), .Z(n5014) );
  NAND U7482 ( .A(n5015), .B(n5014), .Z(y[164]) );
  NAND U7483 ( .A(n5468), .B(m[165]), .Z(n5017) );
  NANDN U7484 ( .A(n5468), .B(creg[165]), .Z(n5016) );
  NAND U7485 ( .A(n5017), .B(n5016), .Z(y[165]) );
  NANDN U7486 ( .A(n5018), .B(n5986), .Z(n5020) );
  NAND U7487 ( .A(n5468), .B(m[166]), .Z(n5019) );
  NAND U7488 ( .A(n5020), .B(n5019), .Z(y[166]) );
  NANDN U7489 ( .A(n5021), .B(n5986), .Z(n5023) );
  NAND U7490 ( .A(n5468), .B(m[167]), .Z(n5022) );
  NAND U7491 ( .A(n5023), .B(n5022), .Z(y[167]) );
  NAND U7492 ( .A(n5468), .B(m[168]), .Z(n5025) );
  NANDN U7493 ( .A(n5468), .B(creg[168]), .Z(n5024) );
  NAND U7494 ( .A(n5025), .B(n5024), .Z(y[168]) );
  NANDN U7495 ( .A(n5026), .B(n5986), .Z(n5028) );
  NAND U7496 ( .A(n5468), .B(m[169]), .Z(n5027) );
  NAND U7497 ( .A(n5028), .B(n5027), .Z(y[169]) );
  NANDN U7498 ( .A(n5029), .B(n5986), .Z(n5031) );
  NAND U7499 ( .A(n5468), .B(m[16]), .Z(n5030) );
  NAND U7500 ( .A(n5031), .B(n5030), .Z(y[16]) );
  NAND U7501 ( .A(n5468), .B(m[170]), .Z(n5033) );
  NANDN U7502 ( .A(n5468), .B(creg[170]), .Z(n5032) );
  NAND U7503 ( .A(n5033), .B(n5032), .Z(y[170]) );
  NAND U7504 ( .A(n5468), .B(m[171]), .Z(n5035) );
  NANDN U7505 ( .A(n5468), .B(creg[171]), .Z(n5034) );
  NAND U7506 ( .A(n5035), .B(n5034), .Z(y[171]) );
  NAND U7507 ( .A(n5468), .B(m[172]), .Z(n5037) );
  NANDN U7508 ( .A(n5468), .B(creg[172]), .Z(n5036) );
  NAND U7509 ( .A(n5037), .B(n5036), .Z(y[172]) );
  NANDN U7510 ( .A(n5038), .B(n5986), .Z(n5040) );
  NAND U7511 ( .A(n5468), .B(m[173]), .Z(n5039) );
  NAND U7512 ( .A(n5040), .B(n5039), .Z(y[173]) );
  NANDN U7513 ( .A(n5041), .B(n5986), .Z(n5043) );
  NAND U7514 ( .A(n5468), .B(m[174]), .Z(n5042) );
  NAND U7515 ( .A(n5043), .B(n5042), .Z(y[174]) );
  NANDN U7516 ( .A(n5044), .B(n5986), .Z(n5046) );
  NAND U7517 ( .A(n5468), .B(m[175]), .Z(n5045) );
  NAND U7518 ( .A(n5046), .B(n5045), .Z(y[175]) );
  NAND U7519 ( .A(n5468), .B(m[176]), .Z(n5048) );
  NANDN U7520 ( .A(n5468), .B(creg[176]), .Z(n5047) );
  NAND U7521 ( .A(n5048), .B(n5047), .Z(y[176]) );
  NAND U7522 ( .A(n5468), .B(m[177]), .Z(n5050) );
  NANDN U7523 ( .A(n5468), .B(creg[177]), .Z(n5049) );
  NAND U7524 ( .A(n5050), .B(n5049), .Z(y[177]) );
  NANDN U7525 ( .A(n5051), .B(n5986), .Z(n5053) );
  NAND U7526 ( .A(n5468), .B(m[178]), .Z(n5052) );
  NAND U7527 ( .A(n5053), .B(n5052), .Z(y[178]) );
  NANDN U7528 ( .A(n5054), .B(n5986), .Z(n5056) );
  NAND U7529 ( .A(n5468), .B(m[179]), .Z(n5055) );
  NAND U7530 ( .A(n5056), .B(n5055), .Z(y[179]) );
  NAND U7531 ( .A(n5468), .B(m[17]), .Z(n5058) );
  NANDN U7532 ( .A(n5468), .B(creg[17]), .Z(n5057) );
  NAND U7533 ( .A(n5058), .B(n5057), .Z(y[17]) );
  NAND U7534 ( .A(n5468), .B(m[180]), .Z(n5060) );
  NANDN U7535 ( .A(n5468), .B(creg[180]), .Z(n5059) );
  NAND U7536 ( .A(n5060), .B(n5059), .Z(y[180]) );
  NAND U7537 ( .A(n5468), .B(m[181]), .Z(n5062) );
  NANDN U7538 ( .A(n5468), .B(creg[181]), .Z(n5061) );
  NAND U7539 ( .A(n5062), .B(n5061), .Z(y[181]) );
  NANDN U7540 ( .A(n5063), .B(n5986), .Z(n5065) );
  NAND U7541 ( .A(n5468), .B(m[182]), .Z(n5064) );
  NAND U7542 ( .A(n5065), .B(n5064), .Z(y[182]) );
  NAND U7543 ( .A(n5468), .B(m[183]), .Z(n5067) );
  NANDN U7544 ( .A(n5468), .B(creg[183]), .Z(n5066) );
  NAND U7545 ( .A(n5067), .B(n5066), .Z(y[183]) );
  NANDN U7546 ( .A(n5068), .B(n5986), .Z(n5070) );
  NAND U7547 ( .A(n5468), .B(m[184]), .Z(n5069) );
  NAND U7548 ( .A(n5070), .B(n5069), .Z(y[184]) );
  NAND U7549 ( .A(n5468), .B(m[185]), .Z(n5072) );
  NANDN U7550 ( .A(n5468), .B(creg[185]), .Z(n5071) );
  NAND U7551 ( .A(n5072), .B(n5071), .Z(y[185]) );
  NAND U7552 ( .A(n5468), .B(m[186]), .Z(n5074) );
  NANDN U7553 ( .A(n5468), .B(creg[186]), .Z(n5073) );
  NAND U7554 ( .A(n5074), .B(n5073), .Z(y[186]) );
  NAND U7555 ( .A(n5468), .B(m[187]), .Z(n5076) );
  NANDN U7556 ( .A(n5468), .B(creg[187]), .Z(n5075) );
  NAND U7557 ( .A(n5076), .B(n5075), .Z(y[187]) );
  NAND U7558 ( .A(n5468), .B(m[188]), .Z(n5078) );
  NANDN U7559 ( .A(n5468), .B(creg[188]), .Z(n5077) );
  NAND U7560 ( .A(n5078), .B(n5077), .Z(y[188]) );
  NAND U7561 ( .A(n5468), .B(m[189]), .Z(n5080) );
  NANDN U7562 ( .A(n5468), .B(creg[189]), .Z(n5079) );
  NAND U7563 ( .A(n5080), .B(n5079), .Z(y[189]) );
  NAND U7564 ( .A(n5468), .B(m[18]), .Z(n5082) );
  NANDN U7565 ( .A(n5468), .B(creg[18]), .Z(n5081) );
  NAND U7566 ( .A(n5082), .B(n5081), .Z(y[18]) );
  NANDN U7567 ( .A(n5083), .B(n5986), .Z(n5085) );
  NAND U7568 ( .A(n5468), .B(m[190]), .Z(n5084) );
  NAND U7569 ( .A(n5085), .B(n5084), .Z(y[190]) );
  NAND U7570 ( .A(n5468), .B(m[191]), .Z(n5087) );
  NANDN U7571 ( .A(n5468), .B(creg[191]), .Z(n5086) );
  NAND U7572 ( .A(n5087), .B(n5086), .Z(y[191]) );
  NANDN U7573 ( .A(n5088), .B(n5986), .Z(n5090) );
  NAND U7574 ( .A(n5468), .B(m[192]), .Z(n5089) );
  NAND U7575 ( .A(n5090), .B(n5089), .Z(y[192]) );
  NAND U7576 ( .A(n5468), .B(m[193]), .Z(n5092) );
  NANDN U7577 ( .A(n5468), .B(creg[193]), .Z(n5091) );
  NAND U7578 ( .A(n5092), .B(n5091), .Z(y[193]) );
  NAND U7579 ( .A(n5468), .B(m[194]), .Z(n5094) );
  NANDN U7580 ( .A(n5468), .B(creg[194]), .Z(n5093) );
  NAND U7581 ( .A(n5094), .B(n5093), .Z(y[194]) );
  NANDN U7582 ( .A(n5095), .B(n5986), .Z(n5097) );
  NAND U7583 ( .A(n5468), .B(m[195]), .Z(n5096) );
  NAND U7584 ( .A(n5097), .B(n5096), .Z(y[195]) );
  NAND U7585 ( .A(n5468), .B(m[196]), .Z(n5099) );
  NANDN U7586 ( .A(n5468), .B(creg[196]), .Z(n5098) );
  NAND U7587 ( .A(n5099), .B(n5098), .Z(y[196]) );
  NANDN U7588 ( .A(n5100), .B(n5986), .Z(n5102) );
  NAND U7589 ( .A(n5468), .B(m[197]), .Z(n5101) );
  NAND U7590 ( .A(n5102), .B(n5101), .Z(y[197]) );
  NANDN U7591 ( .A(n5103), .B(n5986), .Z(n5105) );
  NAND U7592 ( .A(n5468), .B(m[198]), .Z(n5104) );
  NAND U7593 ( .A(n5105), .B(n5104), .Z(y[198]) );
  NANDN U7594 ( .A(n5106), .B(n5986), .Z(n5108) );
  NAND U7595 ( .A(n5468), .B(m[199]), .Z(n5107) );
  NAND U7596 ( .A(n5108), .B(n5107), .Z(y[199]) );
  NANDN U7597 ( .A(n5109), .B(n5986), .Z(n5111) );
  NAND U7598 ( .A(n5468), .B(m[19]), .Z(n5110) );
  NAND U7599 ( .A(n5111), .B(n5110), .Z(y[19]) );
  NANDN U7600 ( .A(n5112), .B(n5986), .Z(n5114) );
  NAND U7601 ( .A(n5468), .B(m[1]), .Z(n5113) );
  NAND U7602 ( .A(n5114), .B(n5113), .Z(y[1]) );
  NAND U7603 ( .A(n5468), .B(m[200]), .Z(n5116) );
  NANDN U7604 ( .A(n5468), .B(creg[200]), .Z(n5115) );
  NAND U7605 ( .A(n5116), .B(n5115), .Z(y[200]) );
  NAND U7606 ( .A(n5468), .B(m[201]), .Z(n5118) );
  NANDN U7607 ( .A(n5468), .B(creg[201]), .Z(n5117) );
  NAND U7608 ( .A(n5118), .B(n5117), .Z(y[201]) );
  NANDN U7609 ( .A(n5119), .B(n5986), .Z(n5121) );
  NAND U7610 ( .A(n5468), .B(m[202]), .Z(n5120) );
  NAND U7611 ( .A(n5121), .B(n5120), .Z(y[202]) );
  NANDN U7612 ( .A(n5122), .B(n5986), .Z(n5124) );
  NAND U7613 ( .A(n5468), .B(m[203]), .Z(n5123) );
  NAND U7614 ( .A(n5124), .B(n5123), .Z(y[203]) );
  NAND U7615 ( .A(n5468), .B(m[204]), .Z(n5126) );
  NANDN U7616 ( .A(n5468), .B(creg[204]), .Z(n5125) );
  NAND U7617 ( .A(n5126), .B(n5125), .Z(y[204]) );
  NANDN U7618 ( .A(n5127), .B(n5986), .Z(n5129) );
  NAND U7619 ( .A(n5468), .B(m[205]), .Z(n5128) );
  NAND U7620 ( .A(n5129), .B(n5128), .Z(y[205]) );
  NANDN U7621 ( .A(n5130), .B(n5986), .Z(n5132) );
  NAND U7622 ( .A(n5468), .B(m[206]), .Z(n5131) );
  NAND U7623 ( .A(n5132), .B(n5131), .Z(y[206]) );
  NANDN U7624 ( .A(n5133), .B(n5986), .Z(n5135) );
  NAND U7625 ( .A(n5468), .B(m[207]), .Z(n5134) );
  NAND U7626 ( .A(n5135), .B(n5134), .Z(y[207]) );
  NAND U7627 ( .A(n5468), .B(m[208]), .Z(n5137) );
  NANDN U7628 ( .A(n5468), .B(creg[208]), .Z(n5136) );
  NAND U7629 ( .A(n5137), .B(n5136), .Z(y[208]) );
  NANDN U7630 ( .A(n5138), .B(n5986), .Z(n5140) );
  NAND U7631 ( .A(n5468), .B(m[209]), .Z(n5139) );
  NAND U7632 ( .A(n5140), .B(n5139), .Z(y[209]) );
  NAND U7633 ( .A(n5468), .B(m[20]), .Z(n5142) );
  NANDN U7634 ( .A(n5468), .B(creg[20]), .Z(n5141) );
  NAND U7635 ( .A(n5142), .B(n5141), .Z(y[20]) );
  NAND U7636 ( .A(n5468), .B(m[210]), .Z(n5144) );
  NANDN U7637 ( .A(n5468), .B(creg[210]), .Z(n5143) );
  NAND U7638 ( .A(n5144), .B(n5143), .Z(y[210]) );
  NAND U7639 ( .A(n5468), .B(m[211]), .Z(n5146) );
  NANDN U7640 ( .A(n5468), .B(creg[211]), .Z(n5145) );
  NAND U7641 ( .A(n5146), .B(n5145), .Z(y[211]) );
  NAND U7642 ( .A(n5468), .B(m[212]), .Z(n5148) );
  NANDN U7643 ( .A(n5468), .B(creg[212]), .Z(n5147) );
  NAND U7644 ( .A(n5148), .B(n5147), .Z(y[212]) );
  NANDN U7645 ( .A(n5149), .B(n5986), .Z(n5151) );
  NAND U7646 ( .A(n5468), .B(m[213]), .Z(n5150) );
  NAND U7647 ( .A(n5151), .B(n5150), .Z(y[213]) );
  NAND U7648 ( .A(n5468), .B(m[214]), .Z(n5153) );
  NANDN U7649 ( .A(n5468), .B(creg[214]), .Z(n5152) );
  NAND U7650 ( .A(n5153), .B(n5152), .Z(y[214]) );
  NANDN U7651 ( .A(n5154), .B(n5986), .Z(n5156) );
  NAND U7652 ( .A(n5468), .B(m[215]), .Z(n5155) );
  NAND U7653 ( .A(n5156), .B(n5155), .Z(y[215]) );
  NANDN U7654 ( .A(n5157), .B(n5986), .Z(n5159) );
  NAND U7655 ( .A(n5468), .B(m[216]), .Z(n5158) );
  NAND U7656 ( .A(n5159), .B(n5158), .Z(y[216]) );
  NAND U7657 ( .A(n5468), .B(m[217]), .Z(n5161) );
  NANDN U7658 ( .A(n5468), .B(creg[217]), .Z(n5160) );
  NAND U7659 ( .A(n5161), .B(n5160), .Z(y[217]) );
  NAND U7660 ( .A(n5468), .B(m[218]), .Z(n5163) );
  NANDN U7661 ( .A(n5468), .B(creg[218]), .Z(n5162) );
  NAND U7662 ( .A(n5163), .B(n5162), .Z(y[218]) );
  NAND U7663 ( .A(n5468), .B(m[219]), .Z(n5165) );
  NANDN U7664 ( .A(n5468), .B(creg[219]), .Z(n5164) );
  NAND U7665 ( .A(n5165), .B(n5164), .Z(y[219]) );
  NAND U7666 ( .A(n5468), .B(m[21]), .Z(n5167) );
  NANDN U7667 ( .A(n5468), .B(creg[21]), .Z(n5166) );
  NAND U7668 ( .A(n5167), .B(n5166), .Z(y[21]) );
  NANDN U7669 ( .A(n5168), .B(n5986), .Z(n5170) );
  NAND U7670 ( .A(n5468), .B(m[220]), .Z(n5169) );
  NAND U7671 ( .A(n5170), .B(n5169), .Z(y[220]) );
  NANDN U7672 ( .A(n5171), .B(n5986), .Z(n5173) );
  NAND U7673 ( .A(n5468), .B(m[221]), .Z(n5172) );
  NAND U7674 ( .A(n5173), .B(n5172), .Z(y[221]) );
  NAND U7675 ( .A(n5468), .B(m[222]), .Z(n5175) );
  NANDN U7676 ( .A(n5468), .B(creg[222]), .Z(n5174) );
  NAND U7677 ( .A(n5175), .B(n5174), .Z(y[222]) );
  NAND U7678 ( .A(n5468), .B(m[223]), .Z(n5177) );
  NANDN U7679 ( .A(n5468), .B(creg[223]), .Z(n5176) );
  NAND U7680 ( .A(n5177), .B(n5176), .Z(y[223]) );
  NAND U7681 ( .A(n5468), .B(m[224]), .Z(n5179) );
  NANDN U7682 ( .A(n5468), .B(creg[224]), .Z(n5178) );
  NAND U7683 ( .A(n5179), .B(n5178), .Z(y[224]) );
  NAND U7684 ( .A(n5468), .B(m[225]), .Z(n5181) );
  NANDN U7685 ( .A(n5468), .B(creg[225]), .Z(n5180) );
  NAND U7686 ( .A(n5181), .B(n5180), .Z(y[225]) );
  NANDN U7687 ( .A(n5182), .B(n5986), .Z(n5184) );
  NAND U7688 ( .A(n5468), .B(m[226]), .Z(n5183) );
  NAND U7689 ( .A(n5184), .B(n5183), .Z(y[226]) );
  NAND U7690 ( .A(n5468), .B(m[227]), .Z(n5186) );
  NANDN U7691 ( .A(n5468), .B(creg[227]), .Z(n5185) );
  NAND U7692 ( .A(n5186), .B(n5185), .Z(y[227]) );
  NAND U7693 ( .A(n5468), .B(m[228]), .Z(n5188) );
  NANDN U7694 ( .A(n5468), .B(creg[228]), .Z(n5187) );
  NAND U7695 ( .A(n5188), .B(n5187), .Z(y[228]) );
  NAND U7696 ( .A(n5468), .B(m[229]), .Z(n5190) );
  NANDN U7697 ( .A(n5468), .B(creg[229]), .Z(n5189) );
  NAND U7698 ( .A(n5190), .B(n5189), .Z(y[229]) );
  NANDN U7699 ( .A(n5191), .B(n5986), .Z(n5193) );
  NAND U7700 ( .A(n5468), .B(m[22]), .Z(n5192) );
  NAND U7701 ( .A(n5193), .B(n5192), .Z(y[22]) );
  NAND U7702 ( .A(n5468), .B(m[230]), .Z(n5195) );
  NANDN U7703 ( .A(n5468), .B(creg[230]), .Z(n5194) );
  NAND U7704 ( .A(n5195), .B(n5194), .Z(y[230]) );
  NAND U7705 ( .A(n5468), .B(m[231]), .Z(n5197) );
  NANDN U7706 ( .A(n5468), .B(creg[231]), .Z(n5196) );
  NAND U7707 ( .A(n5197), .B(n5196), .Z(y[231]) );
  NAND U7708 ( .A(n5468), .B(m[232]), .Z(n5199) );
  NANDN U7709 ( .A(n5468), .B(creg[232]), .Z(n5198) );
  NAND U7710 ( .A(n5199), .B(n5198), .Z(y[232]) );
  NAND U7711 ( .A(n5468), .B(m[233]), .Z(n5201) );
  NANDN U7712 ( .A(n5468), .B(creg[233]), .Z(n5200) );
  NAND U7713 ( .A(n5201), .B(n5200), .Z(y[233]) );
  NANDN U7714 ( .A(n5202), .B(n5986), .Z(n5204) );
  NAND U7715 ( .A(n5468), .B(m[234]), .Z(n5203) );
  NAND U7716 ( .A(n5204), .B(n5203), .Z(y[234]) );
  NAND U7717 ( .A(n5468), .B(m[235]), .Z(n5206) );
  NANDN U7718 ( .A(n5468), .B(creg[235]), .Z(n5205) );
  NAND U7719 ( .A(n5206), .B(n5205), .Z(y[235]) );
  NAND U7720 ( .A(n5468), .B(m[236]), .Z(n5208) );
  NANDN U7721 ( .A(n5468), .B(creg[236]), .Z(n5207) );
  NAND U7722 ( .A(n5208), .B(n5207), .Z(y[236]) );
  NANDN U7723 ( .A(n5209), .B(n5986), .Z(n5211) );
  NAND U7724 ( .A(n5468), .B(m[237]), .Z(n5210) );
  NAND U7725 ( .A(n5211), .B(n5210), .Z(y[237]) );
  NANDN U7726 ( .A(n5212), .B(n5986), .Z(n5214) );
  NAND U7727 ( .A(n5468), .B(m[238]), .Z(n5213) );
  NAND U7728 ( .A(n5214), .B(n5213), .Z(y[238]) );
  NAND U7729 ( .A(n5468), .B(m[239]), .Z(n5216) );
  NANDN U7730 ( .A(n5468), .B(creg[239]), .Z(n5215) );
  NAND U7731 ( .A(n5216), .B(n5215), .Z(y[239]) );
  NAND U7732 ( .A(n5468), .B(m[23]), .Z(n5218) );
  NANDN U7733 ( .A(n5468), .B(creg[23]), .Z(n5217) );
  NAND U7734 ( .A(n5218), .B(n5217), .Z(y[23]) );
  NAND U7735 ( .A(n5468), .B(m[240]), .Z(n5220) );
  NANDN U7736 ( .A(n5468), .B(creg[240]), .Z(n5219) );
  NAND U7737 ( .A(n5220), .B(n5219), .Z(y[240]) );
  NANDN U7738 ( .A(n5221), .B(n5986), .Z(n5223) );
  NAND U7739 ( .A(n5468), .B(m[241]), .Z(n5222) );
  NAND U7740 ( .A(n5223), .B(n5222), .Z(y[241]) );
  NAND U7741 ( .A(n5468), .B(m[242]), .Z(n5225) );
  NANDN U7742 ( .A(n5468), .B(creg[242]), .Z(n5224) );
  NAND U7743 ( .A(n5225), .B(n5224), .Z(y[242]) );
  NANDN U7744 ( .A(n5226), .B(n5986), .Z(n5228) );
  NAND U7745 ( .A(n5468), .B(m[243]), .Z(n5227) );
  NAND U7746 ( .A(n5228), .B(n5227), .Z(y[243]) );
  NANDN U7747 ( .A(n5229), .B(n5986), .Z(n5231) );
  NAND U7748 ( .A(n5468), .B(m[244]), .Z(n5230) );
  NAND U7749 ( .A(n5231), .B(n5230), .Z(y[244]) );
  NAND U7750 ( .A(n5468), .B(m[245]), .Z(n5233) );
  NANDN U7751 ( .A(n5468), .B(creg[245]), .Z(n5232) );
  NAND U7752 ( .A(n5233), .B(n5232), .Z(y[245]) );
  NANDN U7753 ( .A(n5234), .B(n5986), .Z(n5236) );
  NAND U7754 ( .A(n5468), .B(m[246]), .Z(n5235) );
  NAND U7755 ( .A(n5236), .B(n5235), .Z(y[246]) );
  NAND U7756 ( .A(n5468), .B(m[247]), .Z(n5238) );
  NANDN U7757 ( .A(n5468), .B(creg[247]), .Z(n5237) );
  NAND U7758 ( .A(n5238), .B(n5237), .Z(y[247]) );
  NAND U7759 ( .A(n5468), .B(m[248]), .Z(n5240) );
  NANDN U7760 ( .A(n5468), .B(creg[248]), .Z(n5239) );
  NAND U7761 ( .A(n5240), .B(n5239), .Z(y[248]) );
  NANDN U7762 ( .A(n5241), .B(n5986), .Z(n5243) );
  NAND U7763 ( .A(n5468), .B(m[249]), .Z(n5242) );
  NAND U7764 ( .A(n5243), .B(n5242), .Z(y[249]) );
  NAND U7765 ( .A(n5468), .B(m[24]), .Z(n5245) );
  NANDN U7766 ( .A(n5468), .B(creg[24]), .Z(n5244) );
  NAND U7767 ( .A(n5245), .B(n5244), .Z(y[24]) );
  NANDN U7768 ( .A(n5246), .B(n5986), .Z(n5248) );
  NAND U7769 ( .A(n5468), .B(m[250]), .Z(n5247) );
  NAND U7770 ( .A(n5248), .B(n5247), .Z(y[250]) );
  NAND U7771 ( .A(n5468), .B(m[251]), .Z(n5250) );
  NANDN U7772 ( .A(n5468), .B(creg[251]), .Z(n5249) );
  NAND U7773 ( .A(n5250), .B(n5249), .Z(y[251]) );
  NAND U7774 ( .A(n5468), .B(m[252]), .Z(n5252) );
  NANDN U7775 ( .A(n5468), .B(creg[252]), .Z(n5251) );
  NAND U7776 ( .A(n5252), .B(n5251), .Z(y[252]) );
  NAND U7777 ( .A(n5468), .B(m[253]), .Z(n5254) );
  NANDN U7778 ( .A(n5468), .B(creg[253]), .Z(n5253) );
  NAND U7779 ( .A(n5254), .B(n5253), .Z(y[253]) );
  NAND U7780 ( .A(n5468), .B(m[254]), .Z(n5256) );
  NANDN U7781 ( .A(n5468), .B(creg[254]), .Z(n5255) );
  NAND U7782 ( .A(n5256), .B(n5255), .Z(y[254]) );
  NAND U7783 ( .A(n5468), .B(m[255]), .Z(n5258) );
  NANDN U7784 ( .A(n5468), .B(creg[255]), .Z(n5257) );
  NAND U7785 ( .A(n5258), .B(n5257), .Z(y[255]) );
  NAND U7786 ( .A(n5468), .B(m[25]), .Z(n5260) );
  NANDN U7787 ( .A(n5468), .B(creg[25]), .Z(n5259) );
  NAND U7788 ( .A(n5260), .B(n5259), .Z(y[25]) );
  NANDN U7789 ( .A(n5261), .B(n5986), .Z(n5263) );
  NAND U7790 ( .A(n5468), .B(m[26]), .Z(n5262) );
  NAND U7791 ( .A(n5263), .B(n5262), .Z(y[26]) );
  NANDN U7792 ( .A(n5264), .B(n5986), .Z(n5266) );
  NAND U7793 ( .A(n5468), .B(m[27]), .Z(n5265) );
  NAND U7794 ( .A(n5266), .B(n5265), .Z(y[27]) );
  NAND U7795 ( .A(n5468), .B(m[28]), .Z(n5268) );
  NANDN U7796 ( .A(n5468), .B(creg[28]), .Z(n5267) );
  NAND U7797 ( .A(n5268), .B(n5267), .Z(y[28]) );
  NANDN U7798 ( .A(n5269), .B(n5986), .Z(n5271) );
  NAND U7799 ( .A(n5468), .B(m[29]), .Z(n5270) );
  NAND U7800 ( .A(n5271), .B(n5270), .Z(y[29]) );
  NANDN U7801 ( .A(n5272), .B(n5986), .Z(n5274) );
  NAND U7802 ( .A(n5468), .B(m[2]), .Z(n5273) );
  NAND U7803 ( .A(n5274), .B(n5273), .Z(y[2]) );
  NAND U7804 ( .A(n5468), .B(m[30]), .Z(n5276) );
  NANDN U7805 ( .A(n5468), .B(creg[30]), .Z(n5275) );
  NAND U7806 ( .A(n5276), .B(n5275), .Z(y[30]) );
  NANDN U7807 ( .A(n5277), .B(n5986), .Z(n5279) );
  NAND U7808 ( .A(n5468), .B(m[31]), .Z(n5278) );
  NAND U7809 ( .A(n5279), .B(n5278), .Z(y[31]) );
  NANDN U7810 ( .A(n5280), .B(n5986), .Z(n5282) );
  NAND U7811 ( .A(n5468), .B(m[32]), .Z(n5281) );
  NAND U7812 ( .A(n5282), .B(n5281), .Z(y[32]) );
  NAND U7813 ( .A(n5468), .B(m[33]), .Z(n5284) );
  NANDN U7814 ( .A(n5468), .B(creg[33]), .Z(n5283) );
  NAND U7815 ( .A(n5284), .B(n5283), .Z(y[33]) );
  NANDN U7816 ( .A(n5285), .B(n5986), .Z(n5287) );
  NAND U7817 ( .A(n5468), .B(m[34]), .Z(n5286) );
  NAND U7818 ( .A(n5287), .B(n5286), .Z(y[34]) );
  NAND U7819 ( .A(n5468), .B(m[35]), .Z(n5289) );
  NANDN U7820 ( .A(n5468), .B(creg[35]), .Z(n5288) );
  NAND U7821 ( .A(n5289), .B(n5288), .Z(y[35]) );
  NANDN U7822 ( .A(n5290), .B(n5986), .Z(n5292) );
  NAND U7823 ( .A(n5468), .B(m[36]), .Z(n5291) );
  NAND U7824 ( .A(n5292), .B(n5291), .Z(y[36]) );
  NANDN U7825 ( .A(n5293), .B(n5986), .Z(n5295) );
  NAND U7826 ( .A(n5468), .B(m[37]), .Z(n5294) );
  NAND U7827 ( .A(n5295), .B(n5294), .Z(y[37]) );
  NAND U7828 ( .A(n5468), .B(m[38]), .Z(n5297) );
  NANDN U7829 ( .A(n5468), .B(creg[38]), .Z(n5296) );
  NAND U7830 ( .A(n5297), .B(n5296), .Z(y[38]) );
  NAND U7831 ( .A(n5468), .B(m[39]), .Z(n5299) );
  NANDN U7832 ( .A(n5468), .B(creg[39]), .Z(n5298) );
  NAND U7833 ( .A(n5299), .B(n5298), .Z(y[39]) );
  NANDN U7834 ( .A(n5300), .B(n5986), .Z(n5302) );
  NAND U7835 ( .A(n5468), .B(m[3]), .Z(n5301) );
  NAND U7836 ( .A(n5302), .B(n5301), .Z(y[3]) );
  NAND U7837 ( .A(n5468), .B(m[40]), .Z(n5304) );
  NANDN U7838 ( .A(n5468), .B(creg[40]), .Z(n5303) );
  NAND U7839 ( .A(n5304), .B(n5303), .Z(y[40]) );
  NANDN U7840 ( .A(n5305), .B(n5986), .Z(n5307) );
  NAND U7841 ( .A(n5468), .B(m[41]), .Z(n5306) );
  NAND U7842 ( .A(n5307), .B(n5306), .Z(y[41]) );
  NANDN U7843 ( .A(n5308), .B(n5986), .Z(n5310) );
  NAND U7844 ( .A(n5468), .B(m[42]), .Z(n5309) );
  NAND U7845 ( .A(n5310), .B(n5309), .Z(y[42]) );
  NAND U7846 ( .A(n5468), .B(m[43]), .Z(n5312) );
  NANDN U7847 ( .A(n5468), .B(creg[43]), .Z(n5311) );
  NAND U7848 ( .A(n5312), .B(n5311), .Z(y[43]) );
  NAND U7849 ( .A(n5468), .B(m[44]), .Z(n5314) );
  NANDN U7850 ( .A(n5468), .B(creg[44]), .Z(n5313) );
  NAND U7851 ( .A(n5314), .B(n5313), .Z(y[44]) );
  NANDN U7852 ( .A(n5315), .B(n5986), .Z(n5317) );
  NAND U7853 ( .A(n5468), .B(m[45]), .Z(n5316) );
  NAND U7854 ( .A(n5317), .B(n5316), .Z(y[45]) );
  NAND U7855 ( .A(n5468), .B(m[46]), .Z(n5319) );
  NANDN U7856 ( .A(n5468), .B(creg[46]), .Z(n5318) );
  NAND U7857 ( .A(n5319), .B(n5318), .Z(y[46]) );
  NANDN U7858 ( .A(n5320), .B(n5986), .Z(n5322) );
  NAND U7859 ( .A(n5468), .B(m[47]), .Z(n5321) );
  NAND U7860 ( .A(n5322), .B(n5321), .Z(y[47]) );
  NAND U7861 ( .A(n5468), .B(m[48]), .Z(n5324) );
  NANDN U7862 ( .A(n5468), .B(creg[48]), .Z(n5323) );
  NAND U7863 ( .A(n5324), .B(n5323), .Z(y[48]) );
  NANDN U7864 ( .A(n5325), .B(n5986), .Z(n5327) );
  NAND U7865 ( .A(n5468), .B(m[49]), .Z(n5326) );
  NAND U7866 ( .A(n5327), .B(n5326), .Z(y[49]) );
  NANDN U7867 ( .A(n5328), .B(n5986), .Z(n5330) );
  NAND U7868 ( .A(n5468), .B(m[4]), .Z(n5329) );
  NAND U7869 ( .A(n5330), .B(n5329), .Z(y[4]) );
  NAND U7870 ( .A(n5468), .B(m[50]), .Z(n5332) );
  NANDN U7871 ( .A(n5468), .B(creg[50]), .Z(n5331) );
  NAND U7872 ( .A(n5332), .B(n5331), .Z(y[50]) );
  NANDN U7873 ( .A(n5333), .B(n5986), .Z(n5335) );
  NAND U7874 ( .A(n5468), .B(m[51]), .Z(n5334) );
  NAND U7875 ( .A(n5335), .B(n5334), .Z(y[51]) );
  NAND U7876 ( .A(n5468), .B(m[52]), .Z(n5337) );
  NANDN U7877 ( .A(n5468), .B(creg[52]), .Z(n5336) );
  NAND U7878 ( .A(n5337), .B(n5336), .Z(y[52]) );
  NAND U7879 ( .A(n5468), .B(m[53]), .Z(n5339) );
  NANDN U7880 ( .A(n5468), .B(creg[53]), .Z(n5338) );
  NAND U7881 ( .A(n5339), .B(n5338), .Z(y[53]) );
  NANDN U7882 ( .A(n5340), .B(n5986), .Z(n5342) );
  NAND U7883 ( .A(n5468), .B(m[54]), .Z(n5341) );
  NAND U7884 ( .A(n5342), .B(n5341), .Z(y[54]) );
  NANDN U7885 ( .A(n5343), .B(n5986), .Z(n5345) );
  NAND U7886 ( .A(n5468), .B(m[55]), .Z(n5344) );
  NAND U7887 ( .A(n5345), .B(n5344), .Z(y[55]) );
  NANDN U7888 ( .A(n5346), .B(n5986), .Z(n5348) );
  NAND U7889 ( .A(n5468), .B(m[56]), .Z(n5347) );
  NAND U7890 ( .A(n5348), .B(n5347), .Z(y[56]) );
  NAND U7891 ( .A(n5468), .B(m[57]), .Z(n5350) );
  NANDN U7892 ( .A(n5468), .B(creg[57]), .Z(n5349) );
  NAND U7893 ( .A(n5350), .B(n5349), .Z(y[57]) );
  NANDN U7894 ( .A(n5351), .B(n5986), .Z(n5353) );
  NAND U7895 ( .A(n5468), .B(m[58]), .Z(n5352) );
  NAND U7896 ( .A(n5353), .B(n5352), .Z(y[58]) );
  NAND U7897 ( .A(n5468), .B(m[59]), .Z(n5355) );
  NANDN U7898 ( .A(n5468), .B(creg[59]), .Z(n5354) );
  NAND U7899 ( .A(n5355), .B(n5354), .Z(y[59]) );
  NAND U7900 ( .A(n5468), .B(m[5]), .Z(n5357) );
  NANDN U7901 ( .A(n5468), .B(creg[5]), .Z(n5356) );
  NAND U7902 ( .A(n5357), .B(n5356), .Z(y[5]) );
  NANDN U7903 ( .A(n5358), .B(n5986), .Z(n5360) );
  NAND U7904 ( .A(n5468), .B(m[60]), .Z(n5359) );
  NAND U7905 ( .A(n5360), .B(n5359), .Z(y[60]) );
  NAND U7906 ( .A(n5468), .B(m[61]), .Z(n5362) );
  NANDN U7907 ( .A(n5468), .B(creg[61]), .Z(n5361) );
  NAND U7908 ( .A(n5362), .B(n5361), .Z(y[61]) );
  NANDN U7909 ( .A(n5363), .B(n5986), .Z(n5365) );
  NAND U7910 ( .A(n5468), .B(m[62]), .Z(n5364) );
  NAND U7911 ( .A(n5365), .B(n5364), .Z(y[62]) );
  NAND U7912 ( .A(n5468), .B(m[63]), .Z(n5367) );
  NANDN U7913 ( .A(n5468), .B(creg[63]), .Z(n5366) );
  NAND U7914 ( .A(n5367), .B(n5366), .Z(y[63]) );
  NAND U7915 ( .A(n5468), .B(m[64]), .Z(n5369) );
  NANDN U7916 ( .A(n5468), .B(creg[64]), .Z(n5368) );
  NAND U7917 ( .A(n5369), .B(n5368), .Z(y[64]) );
  NAND U7918 ( .A(n5468), .B(m[65]), .Z(n5371) );
  NANDN U7919 ( .A(n5468), .B(creg[65]), .Z(n5370) );
  NAND U7920 ( .A(n5371), .B(n5370), .Z(y[65]) );
  NANDN U7921 ( .A(n5372), .B(n5986), .Z(n5374) );
  NAND U7922 ( .A(n5468), .B(m[66]), .Z(n5373) );
  NAND U7923 ( .A(n5374), .B(n5373), .Z(y[66]) );
  NAND U7924 ( .A(n5468), .B(m[67]), .Z(n5376) );
  NANDN U7925 ( .A(n5468), .B(creg[67]), .Z(n5375) );
  NAND U7926 ( .A(n5376), .B(n5375), .Z(y[67]) );
  NANDN U7927 ( .A(n5377), .B(n5986), .Z(n5379) );
  NAND U7928 ( .A(n5468), .B(m[68]), .Z(n5378) );
  NAND U7929 ( .A(n5379), .B(n5378), .Z(y[68]) );
  NAND U7930 ( .A(n5468), .B(m[69]), .Z(n5381) );
  NANDN U7931 ( .A(n5468), .B(creg[69]), .Z(n5380) );
  NAND U7932 ( .A(n5381), .B(n5380), .Z(y[69]) );
  NAND U7933 ( .A(n5468), .B(m[6]), .Z(n5383) );
  NANDN U7934 ( .A(n5468), .B(creg[6]), .Z(n5382) );
  NAND U7935 ( .A(n5383), .B(n5382), .Z(y[6]) );
  NANDN U7936 ( .A(n5384), .B(n5986), .Z(n5386) );
  NAND U7937 ( .A(n5468), .B(m[70]), .Z(n5385) );
  NAND U7938 ( .A(n5386), .B(n5385), .Z(y[70]) );
  NAND U7939 ( .A(n5468), .B(m[71]), .Z(n5388) );
  NANDN U7940 ( .A(n5468), .B(creg[71]), .Z(n5387) );
  NAND U7941 ( .A(n5388), .B(n5387), .Z(y[71]) );
  NANDN U7942 ( .A(n5389), .B(n5986), .Z(n5391) );
  NAND U7943 ( .A(n5468), .B(m[72]), .Z(n5390) );
  NAND U7944 ( .A(n5391), .B(n5390), .Z(y[72]) );
  NAND U7945 ( .A(n5468), .B(m[73]), .Z(n5393) );
  NANDN U7946 ( .A(n5468), .B(creg[73]), .Z(n5392) );
  NAND U7947 ( .A(n5393), .B(n5392), .Z(y[73]) );
  NANDN U7948 ( .A(n5394), .B(n5986), .Z(n5396) );
  NAND U7949 ( .A(n5468), .B(m[74]), .Z(n5395) );
  NAND U7950 ( .A(n5396), .B(n5395), .Z(y[74]) );
  NANDN U7951 ( .A(n5397), .B(n5986), .Z(n5399) );
  NAND U7952 ( .A(n5468), .B(m[75]), .Z(n5398) );
  NAND U7953 ( .A(n5399), .B(n5398), .Z(y[75]) );
  NANDN U7954 ( .A(n5400), .B(n5986), .Z(n5402) );
  NAND U7955 ( .A(n5468), .B(m[76]), .Z(n5401) );
  NAND U7956 ( .A(n5402), .B(n5401), .Z(y[76]) );
  NANDN U7957 ( .A(n5403), .B(n5986), .Z(n5405) );
  NAND U7958 ( .A(n5468), .B(m[77]), .Z(n5404) );
  NAND U7959 ( .A(n5405), .B(n5404), .Z(y[77]) );
  NAND U7960 ( .A(n5468), .B(m[78]), .Z(n5407) );
  NANDN U7961 ( .A(n5468), .B(creg[78]), .Z(n5406) );
  NAND U7962 ( .A(n5407), .B(n5406), .Z(y[78]) );
  NAND U7963 ( .A(n5468), .B(m[79]), .Z(n5409) );
  NANDN U7964 ( .A(n5468), .B(creg[79]), .Z(n5408) );
  NAND U7965 ( .A(n5409), .B(n5408), .Z(y[79]) );
  NAND U7966 ( .A(n5468), .B(m[7]), .Z(n5411) );
  NANDN U7967 ( .A(n5468), .B(creg[7]), .Z(n5410) );
  NAND U7968 ( .A(n5411), .B(n5410), .Z(y[7]) );
  NANDN U7969 ( .A(n5412), .B(n5986), .Z(n5414) );
  NAND U7970 ( .A(n5468), .B(m[80]), .Z(n5413) );
  NAND U7971 ( .A(n5414), .B(n5413), .Z(y[80]) );
  NANDN U7972 ( .A(n5415), .B(n5986), .Z(n5417) );
  NAND U7973 ( .A(n5468), .B(m[81]), .Z(n5416) );
  NAND U7974 ( .A(n5417), .B(n5416), .Z(y[81]) );
  NANDN U7975 ( .A(n5418), .B(n5986), .Z(n5420) );
  NAND U7976 ( .A(n5468), .B(m[82]), .Z(n5419) );
  NAND U7977 ( .A(n5420), .B(n5419), .Z(y[82]) );
  NANDN U7978 ( .A(n5421), .B(n5986), .Z(n5423) );
  NAND U7979 ( .A(n5468), .B(m[83]), .Z(n5422) );
  NAND U7980 ( .A(n5423), .B(n5422), .Z(y[83]) );
  NAND U7981 ( .A(n5468), .B(m[84]), .Z(n5425) );
  NANDN U7982 ( .A(n5468), .B(creg[84]), .Z(n5424) );
  NAND U7983 ( .A(n5425), .B(n5424), .Z(y[84]) );
  NANDN U7984 ( .A(n5426), .B(n5986), .Z(n5428) );
  NAND U7985 ( .A(n5468), .B(m[85]), .Z(n5427) );
  NAND U7986 ( .A(n5428), .B(n5427), .Z(y[85]) );
  NANDN U7987 ( .A(n5429), .B(n5986), .Z(n5431) );
  NAND U7988 ( .A(n5468), .B(m[86]), .Z(n5430) );
  NAND U7989 ( .A(n5431), .B(n5430), .Z(y[86]) );
  NAND U7990 ( .A(n5468), .B(m[87]), .Z(n5433) );
  NANDN U7991 ( .A(n5468), .B(creg[87]), .Z(n5432) );
  NAND U7992 ( .A(n5433), .B(n5432), .Z(y[87]) );
  NAND U7993 ( .A(n5468), .B(m[88]), .Z(n5435) );
  NANDN U7994 ( .A(n5468), .B(creg[88]), .Z(n5434) );
  NAND U7995 ( .A(n5435), .B(n5434), .Z(y[88]) );
  NAND U7996 ( .A(n5468), .B(m[89]), .Z(n5437) );
  NANDN U7997 ( .A(n5468), .B(creg[89]), .Z(n5436) );
  NAND U7998 ( .A(n5437), .B(n5436), .Z(y[89]) );
  NAND U7999 ( .A(n5468), .B(m[8]), .Z(n5439) );
  NANDN U8000 ( .A(n5468), .B(creg[8]), .Z(n5438) );
  NAND U8001 ( .A(n5439), .B(n5438), .Z(y[8]) );
  NANDN U8002 ( .A(n5440), .B(n5986), .Z(n5442) );
  NAND U8003 ( .A(n5468), .B(m[90]), .Z(n5441) );
  NAND U8004 ( .A(n5442), .B(n5441), .Z(y[90]) );
  NANDN U8005 ( .A(n5443), .B(n5986), .Z(n5445) );
  NAND U8006 ( .A(n5468), .B(m[91]), .Z(n5444) );
  NAND U8007 ( .A(n5445), .B(n5444), .Z(y[91]) );
  NANDN U8008 ( .A(n5446), .B(n5986), .Z(n5448) );
  NAND U8009 ( .A(n5468), .B(m[92]), .Z(n5447) );
  NAND U8010 ( .A(n5448), .B(n5447), .Z(y[92]) );
  NAND U8011 ( .A(n5468), .B(m[93]), .Z(n5450) );
  NANDN U8012 ( .A(n5468), .B(creg[93]), .Z(n5449) );
  NAND U8013 ( .A(n5450), .B(n5449), .Z(y[93]) );
  NANDN U8014 ( .A(n5451), .B(n5986), .Z(n5453) );
  NAND U8015 ( .A(n5468), .B(m[94]), .Z(n5452) );
  NAND U8016 ( .A(n5453), .B(n5452), .Z(y[94]) );
  NANDN U8017 ( .A(n5454), .B(n5986), .Z(n5456) );
  NAND U8018 ( .A(n5468), .B(m[95]), .Z(n5455) );
  NAND U8019 ( .A(n5456), .B(n5455), .Z(y[95]) );
  NANDN U8020 ( .A(n5457), .B(n5986), .Z(n5459) );
  NAND U8021 ( .A(n5468), .B(m[96]), .Z(n5458) );
  NAND U8022 ( .A(n5459), .B(n5458), .Z(y[96]) );
  NANDN U8023 ( .A(n5460), .B(n5986), .Z(n5462) );
  NAND U8024 ( .A(n5468), .B(m[97]), .Z(n5461) );
  NAND U8025 ( .A(n5462), .B(n5461), .Z(y[97]) );
  NANDN U8026 ( .A(n5463), .B(n5986), .Z(n5465) );
  NAND U8027 ( .A(n5468), .B(m[98]), .Z(n5464) );
  NAND U8028 ( .A(n5465), .B(n5464), .Z(y[98]) );
  NAND U8029 ( .A(n5468), .B(m[99]), .Z(n5467) );
  NANDN U8030 ( .A(n5468), .B(creg[99]), .Z(n5466) );
  NAND U8031 ( .A(n5467), .B(n5466), .Z(y[99]) );
  NAND U8032 ( .A(n5468), .B(m[9]), .Z(n5470) );
  NANDN U8033 ( .A(n5468), .B(creg[9]), .Z(n5469) );
  NAND U8034 ( .A(n5470), .B(n5469), .Z(y[9]) );
  ANDN U8035 ( .B(start_reg[511]), .A(n3895), .Z(start_in[511]) );
  AND U8036 ( .A(first_one), .B(start_in[511]), .Z(n5472) );
  NANDN U8037 ( .A(ereg[255]), .B(mul_pow), .Z(n5471) );
  NAND U8038 ( .A(n5472), .B(n5471), .Z(n5983) );
  NAND U8039 ( .A(n3857), .B(o[255]), .Z(n5474) );
  NAND U8040 ( .A(n5983), .B(x[255]), .Z(n5473) );
  NAND U8041 ( .A(n5474), .B(n5473), .Z(n1802) );
  NAND U8042 ( .A(n3857), .B(o[254]), .Z(n5476) );
  NAND U8043 ( .A(n5983), .B(x[254]), .Z(n5475) );
  NAND U8044 ( .A(n5476), .B(n5475), .Z(n1803) );
  NAND U8045 ( .A(n3857), .B(o[253]), .Z(n5478) );
  NAND U8046 ( .A(n5983), .B(x[253]), .Z(n5477) );
  NAND U8047 ( .A(n5478), .B(n5477), .Z(n1804) );
  NAND U8048 ( .A(n3857), .B(o[252]), .Z(n5480) );
  NAND U8049 ( .A(n5983), .B(x[252]), .Z(n5479) );
  NAND U8050 ( .A(n5480), .B(n5479), .Z(n1805) );
  NAND U8051 ( .A(n3857), .B(o[251]), .Z(n5482) );
  NAND U8052 ( .A(n5983), .B(x[251]), .Z(n5481) );
  NAND U8053 ( .A(n5482), .B(n5481), .Z(n1806) );
  NAND U8054 ( .A(n3857), .B(o[250]), .Z(n5484) );
  NAND U8055 ( .A(n5983), .B(x[250]), .Z(n5483) );
  NAND U8056 ( .A(n5484), .B(n5483), .Z(n1807) );
  NAND U8057 ( .A(n3857), .B(o[249]), .Z(n5486) );
  NAND U8058 ( .A(n5983), .B(x[249]), .Z(n5485) );
  NAND U8059 ( .A(n5486), .B(n5485), .Z(n1808) );
  NAND U8060 ( .A(n3857), .B(o[248]), .Z(n5488) );
  NAND U8061 ( .A(n5983), .B(x[248]), .Z(n5487) );
  NAND U8062 ( .A(n5488), .B(n5487), .Z(n1809) );
  NAND U8063 ( .A(n3857), .B(o[247]), .Z(n5490) );
  NAND U8064 ( .A(n5983), .B(x[247]), .Z(n5489) );
  NAND U8065 ( .A(n5490), .B(n5489), .Z(n1810) );
  NAND U8066 ( .A(n3857), .B(o[246]), .Z(n5492) );
  NAND U8067 ( .A(n5983), .B(x[246]), .Z(n5491) );
  NAND U8068 ( .A(n5492), .B(n5491), .Z(n1811) );
  NAND U8069 ( .A(n3857), .B(o[245]), .Z(n5494) );
  NAND U8070 ( .A(n5983), .B(x[245]), .Z(n5493) );
  NAND U8071 ( .A(n5494), .B(n5493), .Z(n1812) );
  NAND U8072 ( .A(n3857), .B(o[244]), .Z(n5496) );
  NAND U8073 ( .A(n5983), .B(x[244]), .Z(n5495) );
  NAND U8074 ( .A(n5496), .B(n5495), .Z(n1813) );
  NAND U8075 ( .A(n3857), .B(o[243]), .Z(n5498) );
  NAND U8076 ( .A(n5983), .B(x[243]), .Z(n5497) );
  NAND U8077 ( .A(n5498), .B(n5497), .Z(n1814) );
  NAND U8078 ( .A(n3857), .B(o[242]), .Z(n5500) );
  NAND U8079 ( .A(n5983), .B(x[242]), .Z(n5499) );
  NAND U8080 ( .A(n5500), .B(n5499), .Z(n1815) );
  NAND U8081 ( .A(n3857), .B(o[241]), .Z(n5502) );
  NAND U8082 ( .A(n5983), .B(x[241]), .Z(n5501) );
  NAND U8083 ( .A(n5502), .B(n5501), .Z(n1816) );
  NAND U8084 ( .A(n3857), .B(o[240]), .Z(n5504) );
  NAND U8085 ( .A(n5983), .B(x[240]), .Z(n5503) );
  NAND U8086 ( .A(n5504), .B(n5503), .Z(n1817) );
  NAND U8087 ( .A(n3857), .B(o[239]), .Z(n5506) );
  NAND U8088 ( .A(n5983), .B(x[239]), .Z(n5505) );
  NAND U8089 ( .A(n5506), .B(n5505), .Z(n1818) );
  NAND U8090 ( .A(n3857), .B(o[238]), .Z(n5508) );
  NAND U8091 ( .A(n5983), .B(x[238]), .Z(n5507) );
  NAND U8092 ( .A(n5508), .B(n5507), .Z(n1819) );
  NAND U8093 ( .A(n3857), .B(o[237]), .Z(n5510) );
  NAND U8094 ( .A(n5983), .B(x[237]), .Z(n5509) );
  NAND U8095 ( .A(n5510), .B(n5509), .Z(n1820) );
  NAND U8096 ( .A(n3857), .B(o[236]), .Z(n5512) );
  NAND U8097 ( .A(n5983), .B(x[236]), .Z(n5511) );
  NAND U8098 ( .A(n5512), .B(n5511), .Z(n1821) );
  NAND U8099 ( .A(n3857), .B(o[235]), .Z(n5514) );
  NAND U8100 ( .A(n5983), .B(x[235]), .Z(n5513) );
  NAND U8101 ( .A(n5514), .B(n5513), .Z(n1822) );
  NAND U8102 ( .A(n3857), .B(o[234]), .Z(n5516) );
  NAND U8103 ( .A(n5983), .B(x[234]), .Z(n5515) );
  NAND U8104 ( .A(n5516), .B(n5515), .Z(n1823) );
  NAND U8105 ( .A(n3857), .B(o[233]), .Z(n5518) );
  NAND U8106 ( .A(n5983), .B(x[233]), .Z(n5517) );
  NAND U8107 ( .A(n5518), .B(n5517), .Z(n1824) );
  NAND U8108 ( .A(n3857), .B(o[232]), .Z(n5520) );
  NAND U8109 ( .A(n5983), .B(x[232]), .Z(n5519) );
  NAND U8110 ( .A(n5520), .B(n5519), .Z(n1825) );
  NAND U8111 ( .A(n3857), .B(o[231]), .Z(n5522) );
  NAND U8112 ( .A(n5983), .B(x[231]), .Z(n5521) );
  NAND U8113 ( .A(n5522), .B(n5521), .Z(n1826) );
  NAND U8114 ( .A(n3857), .B(o[230]), .Z(n5524) );
  NAND U8115 ( .A(n5983), .B(x[230]), .Z(n5523) );
  NAND U8116 ( .A(n5524), .B(n5523), .Z(n1827) );
  NAND U8117 ( .A(n3857), .B(o[229]), .Z(n5526) );
  NAND U8118 ( .A(n5983), .B(x[229]), .Z(n5525) );
  NAND U8119 ( .A(n5526), .B(n5525), .Z(n1828) );
  NAND U8120 ( .A(n3857), .B(o[228]), .Z(n5528) );
  NAND U8121 ( .A(n5983), .B(x[228]), .Z(n5527) );
  NAND U8122 ( .A(n5528), .B(n5527), .Z(n1829) );
  NAND U8123 ( .A(n3857), .B(o[227]), .Z(n5530) );
  NAND U8124 ( .A(n5983), .B(x[227]), .Z(n5529) );
  NAND U8125 ( .A(n5530), .B(n5529), .Z(n1830) );
  NAND U8126 ( .A(n3857), .B(o[226]), .Z(n5532) );
  NAND U8127 ( .A(n5983), .B(x[226]), .Z(n5531) );
  NAND U8128 ( .A(n5532), .B(n5531), .Z(n1831) );
  NAND U8129 ( .A(n3857), .B(o[225]), .Z(n5534) );
  NAND U8130 ( .A(n5983), .B(x[225]), .Z(n5533) );
  NAND U8131 ( .A(n5534), .B(n5533), .Z(n1832) );
  NAND U8132 ( .A(n3857), .B(o[224]), .Z(n5536) );
  NAND U8133 ( .A(n5983), .B(x[224]), .Z(n5535) );
  NAND U8134 ( .A(n5536), .B(n5535), .Z(n1833) );
  NAND U8135 ( .A(n3857), .B(o[223]), .Z(n5538) );
  NAND U8136 ( .A(n5983), .B(x[223]), .Z(n5537) );
  NAND U8137 ( .A(n5538), .B(n5537), .Z(n1834) );
  NAND U8138 ( .A(n3857), .B(o[222]), .Z(n5540) );
  NAND U8139 ( .A(n5983), .B(x[222]), .Z(n5539) );
  NAND U8140 ( .A(n5540), .B(n5539), .Z(n1835) );
  NAND U8141 ( .A(n3857), .B(o[221]), .Z(n5542) );
  NAND U8142 ( .A(n5983), .B(x[221]), .Z(n5541) );
  NAND U8143 ( .A(n5542), .B(n5541), .Z(n1836) );
  NAND U8144 ( .A(n3857), .B(o[220]), .Z(n5544) );
  NAND U8145 ( .A(n5983), .B(x[220]), .Z(n5543) );
  NAND U8146 ( .A(n5544), .B(n5543), .Z(n1837) );
  NAND U8147 ( .A(n3857), .B(o[219]), .Z(n5546) );
  NAND U8148 ( .A(n5983), .B(x[219]), .Z(n5545) );
  NAND U8149 ( .A(n5546), .B(n5545), .Z(n1838) );
  NAND U8150 ( .A(n3857), .B(o[218]), .Z(n5548) );
  NAND U8151 ( .A(n5983), .B(x[218]), .Z(n5547) );
  NAND U8152 ( .A(n5548), .B(n5547), .Z(n1839) );
  NAND U8153 ( .A(n3857), .B(o[217]), .Z(n5550) );
  NAND U8154 ( .A(n5983), .B(x[217]), .Z(n5549) );
  NAND U8155 ( .A(n5550), .B(n5549), .Z(n1840) );
  NAND U8156 ( .A(n3857), .B(o[216]), .Z(n5552) );
  NAND U8157 ( .A(n5983), .B(x[216]), .Z(n5551) );
  NAND U8158 ( .A(n5552), .B(n5551), .Z(n1841) );
  NAND U8159 ( .A(n3857), .B(o[215]), .Z(n5554) );
  NAND U8160 ( .A(n5983), .B(x[215]), .Z(n5553) );
  NAND U8161 ( .A(n5554), .B(n5553), .Z(n1842) );
  NAND U8162 ( .A(n3857), .B(o[214]), .Z(n5556) );
  NAND U8163 ( .A(n5983), .B(x[214]), .Z(n5555) );
  NAND U8164 ( .A(n5556), .B(n5555), .Z(n1843) );
  NAND U8165 ( .A(n3857), .B(o[213]), .Z(n5558) );
  NAND U8166 ( .A(n5983), .B(x[213]), .Z(n5557) );
  NAND U8167 ( .A(n5558), .B(n5557), .Z(n1844) );
  NAND U8168 ( .A(n3857), .B(o[212]), .Z(n5560) );
  NAND U8169 ( .A(n5983), .B(x[212]), .Z(n5559) );
  NAND U8170 ( .A(n5560), .B(n5559), .Z(n1845) );
  NAND U8171 ( .A(n3857), .B(o[211]), .Z(n5562) );
  NAND U8172 ( .A(n5983), .B(x[211]), .Z(n5561) );
  NAND U8173 ( .A(n5562), .B(n5561), .Z(n1846) );
  NAND U8174 ( .A(n3857), .B(o[210]), .Z(n5564) );
  NAND U8175 ( .A(n5983), .B(x[210]), .Z(n5563) );
  NAND U8176 ( .A(n5564), .B(n5563), .Z(n1847) );
  NAND U8177 ( .A(n3857), .B(o[209]), .Z(n5566) );
  NAND U8178 ( .A(n5983), .B(x[209]), .Z(n5565) );
  NAND U8179 ( .A(n5566), .B(n5565), .Z(n1848) );
  NAND U8180 ( .A(n3857), .B(o[208]), .Z(n5568) );
  NAND U8181 ( .A(n5983), .B(x[208]), .Z(n5567) );
  NAND U8182 ( .A(n5568), .B(n5567), .Z(n1849) );
  NAND U8183 ( .A(n3857), .B(o[207]), .Z(n5570) );
  NAND U8184 ( .A(n5983), .B(x[207]), .Z(n5569) );
  NAND U8185 ( .A(n5570), .B(n5569), .Z(n1850) );
  NAND U8186 ( .A(n3857), .B(o[206]), .Z(n5572) );
  NAND U8187 ( .A(n5983), .B(x[206]), .Z(n5571) );
  NAND U8188 ( .A(n5572), .B(n5571), .Z(n1851) );
  NAND U8189 ( .A(n3857), .B(o[205]), .Z(n5574) );
  NAND U8190 ( .A(n5983), .B(x[205]), .Z(n5573) );
  NAND U8191 ( .A(n5574), .B(n5573), .Z(n1852) );
  NAND U8192 ( .A(n3857), .B(o[204]), .Z(n5576) );
  NAND U8193 ( .A(n5983), .B(x[204]), .Z(n5575) );
  NAND U8194 ( .A(n5576), .B(n5575), .Z(n1853) );
  NAND U8195 ( .A(n3857), .B(o[203]), .Z(n5578) );
  NAND U8196 ( .A(n5983), .B(x[203]), .Z(n5577) );
  NAND U8197 ( .A(n5578), .B(n5577), .Z(n1854) );
  NAND U8198 ( .A(n3857), .B(o[202]), .Z(n5580) );
  NAND U8199 ( .A(n5983), .B(x[202]), .Z(n5579) );
  NAND U8200 ( .A(n5580), .B(n5579), .Z(n1855) );
  NAND U8201 ( .A(n3857), .B(o[201]), .Z(n5582) );
  NAND U8202 ( .A(n5983), .B(x[201]), .Z(n5581) );
  NAND U8203 ( .A(n5582), .B(n5581), .Z(n1856) );
  NAND U8204 ( .A(n3857), .B(o[200]), .Z(n5584) );
  NAND U8205 ( .A(n5983), .B(x[200]), .Z(n5583) );
  NAND U8206 ( .A(n5584), .B(n5583), .Z(n1857) );
  NAND U8207 ( .A(n3857), .B(o[199]), .Z(n5586) );
  NAND U8208 ( .A(n5983), .B(x[199]), .Z(n5585) );
  NAND U8209 ( .A(n5586), .B(n5585), .Z(n1858) );
  NAND U8210 ( .A(n3857), .B(o[198]), .Z(n5588) );
  NAND U8211 ( .A(n5983), .B(x[198]), .Z(n5587) );
  NAND U8212 ( .A(n5588), .B(n5587), .Z(n1859) );
  NAND U8213 ( .A(n3857), .B(o[197]), .Z(n5590) );
  NAND U8214 ( .A(n5983), .B(x[197]), .Z(n5589) );
  NAND U8215 ( .A(n5590), .B(n5589), .Z(n1860) );
  NAND U8216 ( .A(n3857), .B(o[196]), .Z(n5592) );
  NAND U8217 ( .A(n5983), .B(x[196]), .Z(n5591) );
  NAND U8218 ( .A(n5592), .B(n5591), .Z(n1861) );
  NAND U8219 ( .A(n3857), .B(o[195]), .Z(n5594) );
  NAND U8220 ( .A(n5983), .B(x[195]), .Z(n5593) );
  NAND U8221 ( .A(n5594), .B(n5593), .Z(n1862) );
  NAND U8222 ( .A(n3857), .B(o[194]), .Z(n5596) );
  NAND U8223 ( .A(n5983), .B(x[194]), .Z(n5595) );
  NAND U8224 ( .A(n5596), .B(n5595), .Z(n1863) );
  NAND U8225 ( .A(n3857), .B(o[193]), .Z(n5598) );
  NAND U8226 ( .A(n5983), .B(x[193]), .Z(n5597) );
  NAND U8227 ( .A(n5598), .B(n5597), .Z(n1864) );
  NAND U8228 ( .A(n3857), .B(o[192]), .Z(n5600) );
  NAND U8229 ( .A(n5983), .B(x[192]), .Z(n5599) );
  NAND U8230 ( .A(n5600), .B(n5599), .Z(n1865) );
  NAND U8231 ( .A(n3857), .B(o[191]), .Z(n5602) );
  NAND U8232 ( .A(n5983), .B(x[191]), .Z(n5601) );
  NAND U8233 ( .A(n5602), .B(n5601), .Z(n1866) );
  NAND U8234 ( .A(n3857), .B(o[190]), .Z(n5604) );
  NAND U8235 ( .A(n5983), .B(x[190]), .Z(n5603) );
  NAND U8236 ( .A(n5604), .B(n5603), .Z(n1867) );
  NAND U8237 ( .A(n3857), .B(o[189]), .Z(n5606) );
  NAND U8238 ( .A(n5983), .B(x[189]), .Z(n5605) );
  NAND U8239 ( .A(n5606), .B(n5605), .Z(n1868) );
  NAND U8240 ( .A(n3857), .B(o[188]), .Z(n5608) );
  NAND U8241 ( .A(n5983), .B(x[188]), .Z(n5607) );
  NAND U8242 ( .A(n5608), .B(n5607), .Z(n1869) );
  NAND U8243 ( .A(n3857), .B(o[187]), .Z(n5610) );
  NAND U8244 ( .A(n5983), .B(x[187]), .Z(n5609) );
  NAND U8245 ( .A(n5610), .B(n5609), .Z(n1870) );
  NAND U8246 ( .A(n3857), .B(o[186]), .Z(n5612) );
  NAND U8247 ( .A(n5983), .B(x[186]), .Z(n5611) );
  NAND U8248 ( .A(n5612), .B(n5611), .Z(n1871) );
  NAND U8249 ( .A(n3857), .B(o[185]), .Z(n5614) );
  NAND U8250 ( .A(n5983), .B(x[185]), .Z(n5613) );
  NAND U8251 ( .A(n5614), .B(n5613), .Z(n1872) );
  NAND U8252 ( .A(n3857), .B(o[184]), .Z(n5616) );
  NAND U8253 ( .A(n5983), .B(x[184]), .Z(n5615) );
  NAND U8254 ( .A(n5616), .B(n5615), .Z(n1873) );
  NAND U8255 ( .A(n3857), .B(o[183]), .Z(n5618) );
  NAND U8256 ( .A(n5983), .B(x[183]), .Z(n5617) );
  NAND U8257 ( .A(n5618), .B(n5617), .Z(n1874) );
  NAND U8258 ( .A(n3857), .B(o[182]), .Z(n5620) );
  NAND U8259 ( .A(n5983), .B(x[182]), .Z(n5619) );
  NAND U8260 ( .A(n5620), .B(n5619), .Z(n1875) );
  NAND U8261 ( .A(n3857), .B(o[181]), .Z(n5622) );
  NAND U8262 ( .A(n5983), .B(x[181]), .Z(n5621) );
  NAND U8263 ( .A(n5622), .B(n5621), .Z(n1876) );
  NAND U8264 ( .A(n3857), .B(o[180]), .Z(n5624) );
  NAND U8265 ( .A(n5983), .B(x[180]), .Z(n5623) );
  NAND U8266 ( .A(n5624), .B(n5623), .Z(n1877) );
  NAND U8267 ( .A(n3857), .B(o[179]), .Z(n5626) );
  NAND U8268 ( .A(n5983), .B(x[179]), .Z(n5625) );
  NAND U8269 ( .A(n5626), .B(n5625), .Z(n1878) );
  NAND U8270 ( .A(n3857), .B(o[178]), .Z(n5628) );
  NAND U8271 ( .A(n5983), .B(x[178]), .Z(n5627) );
  NAND U8272 ( .A(n5628), .B(n5627), .Z(n1879) );
  NAND U8273 ( .A(n3857), .B(o[177]), .Z(n5630) );
  NAND U8274 ( .A(n5983), .B(x[177]), .Z(n5629) );
  NAND U8275 ( .A(n5630), .B(n5629), .Z(n1880) );
  NAND U8276 ( .A(n3857), .B(o[176]), .Z(n5632) );
  NAND U8277 ( .A(n5983), .B(x[176]), .Z(n5631) );
  NAND U8278 ( .A(n5632), .B(n5631), .Z(n1881) );
  NAND U8279 ( .A(n3857), .B(o[175]), .Z(n5634) );
  NAND U8280 ( .A(n5983), .B(x[175]), .Z(n5633) );
  NAND U8281 ( .A(n5634), .B(n5633), .Z(n1882) );
  NAND U8282 ( .A(n3857), .B(o[174]), .Z(n5636) );
  NAND U8283 ( .A(n5983), .B(x[174]), .Z(n5635) );
  NAND U8284 ( .A(n5636), .B(n5635), .Z(n1883) );
  NAND U8285 ( .A(n3857), .B(o[173]), .Z(n5638) );
  NAND U8286 ( .A(n5983), .B(x[173]), .Z(n5637) );
  NAND U8287 ( .A(n5638), .B(n5637), .Z(n1884) );
  NAND U8288 ( .A(n3857), .B(o[172]), .Z(n5640) );
  NAND U8289 ( .A(n5983), .B(x[172]), .Z(n5639) );
  NAND U8290 ( .A(n5640), .B(n5639), .Z(n1885) );
  NAND U8291 ( .A(n3857), .B(o[171]), .Z(n5642) );
  NAND U8292 ( .A(n5983), .B(x[171]), .Z(n5641) );
  NAND U8293 ( .A(n5642), .B(n5641), .Z(n1886) );
  NAND U8294 ( .A(n3857), .B(o[170]), .Z(n5644) );
  NAND U8295 ( .A(n5983), .B(x[170]), .Z(n5643) );
  NAND U8296 ( .A(n5644), .B(n5643), .Z(n1887) );
  NAND U8297 ( .A(n3857), .B(o[169]), .Z(n5646) );
  NAND U8298 ( .A(n5983), .B(x[169]), .Z(n5645) );
  NAND U8299 ( .A(n5646), .B(n5645), .Z(n1888) );
  NAND U8300 ( .A(n3857), .B(o[168]), .Z(n5648) );
  NAND U8301 ( .A(n5983), .B(x[168]), .Z(n5647) );
  NAND U8302 ( .A(n5648), .B(n5647), .Z(n1889) );
  NAND U8303 ( .A(n3857), .B(o[167]), .Z(n5650) );
  NAND U8304 ( .A(n5983), .B(x[167]), .Z(n5649) );
  NAND U8305 ( .A(n5650), .B(n5649), .Z(n1890) );
  NAND U8306 ( .A(n3857), .B(o[166]), .Z(n5652) );
  NAND U8307 ( .A(n5983), .B(x[166]), .Z(n5651) );
  NAND U8308 ( .A(n5652), .B(n5651), .Z(n1891) );
  NAND U8309 ( .A(n3857), .B(o[165]), .Z(n5654) );
  NAND U8310 ( .A(n5983), .B(x[165]), .Z(n5653) );
  NAND U8311 ( .A(n5654), .B(n5653), .Z(n1892) );
  NAND U8312 ( .A(n3857), .B(o[164]), .Z(n5656) );
  NAND U8313 ( .A(n5983), .B(x[164]), .Z(n5655) );
  NAND U8314 ( .A(n5656), .B(n5655), .Z(n1893) );
  NAND U8315 ( .A(n3857), .B(o[163]), .Z(n5658) );
  NAND U8316 ( .A(n5983), .B(x[163]), .Z(n5657) );
  NAND U8317 ( .A(n5658), .B(n5657), .Z(n1894) );
  NAND U8318 ( .A(n3857), .B(o[162]), .Z(n5660) );
  NAND U8319 ( .A(n5983), .B(x[162]), .Z(n5659) );
  NAND U8320 ( .A(n5660), .B(n5659), .Z(n1895) );
  NAND U8321 ( .A(n3857), .B(o[161]), .Z(n5662) );
  NAND U8322 ( .A(n5983), .B(x[161]), .Z(n5661) );
  NAND U8323 ( .A(n5662), .B(n5661), .Z(n1896) );
  NAND U8324 ( .A(n3857), .B(o[160]), .Z(n5664) );
  NAND U8325 ( .A(n5983), .B(x[160]), .Z(n5663) );
  NAND U8326 ( .A(n5664), .B(n5663), .Z(n1897) );
  NAND U8327 ( .A(n3857), .B(o[159]), .Z(n5666) );
  NAND U8328 ( .A(n5983), .B(x[159]), .Z(n5665) );
  NAND U8329 ( .A(n5666), .B(n5665), .Z(n1898) );
  NAND U8330 ( .A(n3857), .B(o[158]), .Z(n5668) );
  NAND U8331 ( .A(n5983), .B(x[158]), .Z(n5667) );
  NAND U8332 ( .A(n5668), .B(n5667), .Z(n1899) );
  NAND U8333 ( .A(n3857), .B(o[157]), .Z(n5670) );
  NAND U8334 ( .A(n5983), .B(x[157]), .Z(n5669) );
  NAND U8335 ( .A(n5670), .B(n5669), .Z(n1900) );
  NAND U8336 ( .A(n3857), .B(o[156]), .Z(n5672) );
  NAND U8337 ( .A(n5983), .B(x[156]), .Z(n5671) );
  NAND U8338 ( .A(n5672), .B(n5671), .Z(n1901) );
  NAND U8339 ( .A(n3857), .B(o[155]), .Z(n5674) );
  NAND U8340 ( .A(n5983), .B(x[155]), .Z(n5673) );
  NAND U8341 ( .A(n5674), .B(n5673), .Z(n1902) );
  NAND U8342 ( .A(n3857), .B(o[154]), .Z(n5676) );
  NAND U8343 ( .A(n5983), .B(x[154]), .Z(n5675) );
  NAND U8344 ( .A(n5676), .B(n5675), .Z(n1903) );
  NAND U8345 ( .A(n3857), .B(o[153]), .Z(n5678) );
  NAND U8346 ( .A(n5983), .B(x[153]), .Z(n5677) );
  NAND U8347 ( .A(n5678), .B(n5677), .Z(n1904) );
  NAND U8348 ( .A(n3857), .B(o[152]), .Z(n5680) );
  NAND U8349 ( .A(n5983), .B(x[152]), .Z(n5679) );
  NAND U8350 ( .A(n5680), .B(n5679), .Z(n1905) );
  NAND U8351 ( .A(n3857), .B(o[151]), .Z(n5682) );
  NAND U8352 ( .A(n5983), .B(x[151]), .Z(n5681) );
  NAND U8353 ( .A(n5682), .B(n5681), .Z(n1906) );
  NAND U8354 ( .A(n3857), .B(o[150]), .Z(n5684) );
  NAND U8355 ( .A(n5983), .B(x[150]), .Z(n5683) );
  NAND U8356 ( .A(n5684), .B(n5683), .Z(n1907) );
  NAND U8357 ( .A(n3857), .B(o[149]), .Z(n5686) );
  NAND U8358 ( .A(n5983), .B(x[149]), .Z(n5685) );
  NAND U8359 ( .A(n5686), .B(n5685), .Z(n1908) );
  NAND U8360 ( .A(n3857), .B(o[148]), .Z(n5688) );
  NAND U8361 ( .A(n5983), .B(x[148]), .Z(n5687) );
  NAND U8362 ( .A(n5688), .B(n5687), .Z(n1909) );
  NAND U8363 ( .A(n3857), .B(o[147]), .Z(n5690) );
  NAND U8364 ( .A(n5983), .B(x[147]), .Z(n5689) );
  NAND U8365 ( .A(n5690), .B(n5689), .Z(n1910) );
  NAND U8366 ( .A(n3857), .B(o[146]), .Z(n5692) );
  NAND U8367 ( .A(n5983), .B(x[146]), .Z(n5691) );
  NAND U8368 ( .A(n5692), .B(n5691), .Z(n1911) );
  NAND U8369 ( .A(n3857), .B(o[145]), .Z(n5694) );
  NAND U8370 ( .A(n5983), .B(x[145]), .Z(n5693) );
  NAND U8371 ( .A(n5694), .B(n5693), .Z(n1912) );
  NAND U8372 ( .A(n3857), .B(o[144]), .Z(n5696) );
  NAND U8373 ( .A(n5983), .B(x[144]), .Z(n5695) );
  NAND U8374 ( .A(n5696), .B(n5695), .Z(n1913) );
  NAND U8375 ( .A(n3857), .B(o[143]), .Z(n5698) );
  NAND U8376 ( .A(n5983), .B(x[143]), .Z(n5697) );
  NAND U8377 ( .A(n5698), .B(n5697), .Z(n1914) );
  NAND U8378 ( .A(n3857), .B(o[142]), .Z(n5700) );
  NAND U8379 ( .A(n5983), .B(x[142]), .Z(n5699) );
  NAND U8380 ( .A(n5700), .B(n5699), .Z(n1915) );
  NAND U8381 ( .A(n3857), .B(o[141]), .Z(n5702) );
  NAND U8382 ( .A(n5983), .B(x[141]), .Z(n5701) );
  NAND U8383 ( .A(n5702), .B(n5701), .Z(n1916) );
  NAND U8384 ( .A(n3857), .B(o[140]), .Z(n5704) );
  NAND U8385 ( .A(n5983), .B(x[140]), .Z(n5703) );
  NAND U8386 ( .A(n5704), .B(n5703), .Z(n1917) );
  NAND U8387 ( .A(n3857), .B(o[139]), .Z(n5706) );
  NAND U8388 ( .A(n5983), .B(x[139]), .Z(n5705) );
  NAND U8389 ( .A(n5706), .B(n5705), .Z(n1918) );
  NAND U8390 ( .A(n3857), .B(o[138]), .Z(n5708) );
  NAND U8391 ( .A(n5983), .B(x[138]), .Z(n5707) );
  NAND U8392 ( .A(n5708), .B(n5707), .Z(n1919) );
  NAND U8393 ( .A(n3857), .B(o[137]), .Z(n5710) );
  NAND U8394 ( .A(n5983), .B(x[137]), .Z(n5709) );
  NAND U8395 ( .A(n5710), .B(n5709), .Z(n1920) );
  NAND U8396 ( .A(n3857), .B(o[136]), .Z(n5712) );
  NAND U8397 ( .A(n5983), .B(x[136]), .Z(n5711) );
  NAND U8398 ( .A(n5712), .B(n5711), .Z(n1921) );
  NAND U8399 ( .A(n3857), .B(o[135]), .Z(n5714) );
  NAND U8400 ( .A(n5983), .B(x[135]), .Z(n5713) );
  NAND U8401 ( .A(n5714), .B(n5713), .Z(n1922) );
  NAND U8402 ( .A(n3857), .B(o[134]), .Z(n5716) );
  NAND U8403 ( .A(n5983), .B(x[134]), .Z(n5715) );
  NAND U8404 ( .A(n5716), .B(n5715), .Z(n1923) );
  NAND U8405 ( .A(n3857), .B(o[133]), .Z(n5718) );
  NAND U8406 ( .A(n5983), .B(x[133]), .Z(n5717) );
  NAND U8407 ( .A(n5718), .B(n5717), .Z(n1924) );
  NAND U8408 ( .A(n3857), .B(o[132]), .Z(n5720) );
  NAND U8409 ( .A(n5983), .B(x[132]), .Z(n5719) );
  NAND U8410 ( .A(n5720), .B(n5719), .Z(n1925) );
  NAND U8411 ( .A(n3857), .B(o[131]), .Z(n5722) );
  NAND U8412 ( .A(n5983), .B(x[131]), .Z(n5721) );
  NAND U8413 ( .A(n5722), .B(n5721), .Z(n1926) );
  NAND U8414 ( .A(n3857), .B(o[130]), .Z(n5724) );
  NAND U8415 ( .A(n5983), .B(x[130]), .Z(n5723) );
  NAND U8416 ( .A(n5724), .B(n5723), .Z(n1927) );
  NAND U8417 ( .A(n3857), .B(o[129]), .Z(n5726) );
  NAND U8418 ( .A(n5983), .B(x[129]), .Z(n5725) );
  NAND U8419 ( .A(n5726), .B(n5725), .Z(n1928) );
  NAND U8420 ( .A(n3857), .B(o[128]), .Z(n5728) );
  NAND U8421 ( .A(n5983), .B(x[128]), .Z(n5727) );
  NAND U8422 ( .A(n5728), .B(n5727), .Z(n1929) );
  NAND U8423 ( .A(n3857), .B(o[127]), .Z(n5730) );
  NAND U8424 ( .A(n5983), .B(x[127]), .Z(n5729) );
  NAND U8425 ( .A(n5730), .B(n5729), .Z(n1930) );
  NAND U8426 ( .A(n3857), .B(o[126]), .Z(n5732) );
  NAND U8427 ( .A(n5983), .B(x[126]), .Z(n5731) );
  NAND U8428 ( .A(n5732), .B(n5731), .Z(n1931) );
  NAND U8429 ( .A(n3857), .B(o[125]), .Z(n5734) );
  NAND U8430 ( .A(n5983), .B(x[125]), .Z(n5733) );
  NAND U8431 ( .A(n5734), .B(n5733), .Z(n1932) );
  NAND U8432 ( .A(n3857), .B(o[124]), .Z(n5736) );
  NAND U8433 ( .A(n5983), .B(x[124]), .Z(n5735) );
  NAND U8434 ( .A(n5736), .B(n5735), .Z(n1933) );
  NAND U8435 ( .A(n3857), .B(o[123]), .Z(n5738) );
  NAND U8436 ( .A(n5983), .B(x[123]), .Z(n5737) );
  NAND U8437 ( .A(n5738), .B(n5737), .Z(n1934) );
  NAND U8438 ( .A(n3857), .B(o[122]), .Z(n5740) );
  NAND U8439 ( .A(n5983), .B(x[122]), .Z(n5739) );
  NAND U8440 ( .A(n5740), .B(n5739), .Z(n1935) );
  NAND U8441 ( .A(n3857), .B(o[121]), .Z(n5742) );
  NAND U8442 ( .A(n5983), .B(x[121]), .Z(n5741) );
  NAND U8443 ( .A(n5742), .B(n5741), .Z(n1936) );
  NAND U8444 ( .A(n3857), .B(o[120]), .Z(n5744) );
  NAND U8445 ( .A(n5983), .B(x[120]), .Z(n5743) );
  NAND U8446 ( .A(n5744), .B(n5743), .Z(n1937) );
  NAND U8447 ( .A(n3857), .B(o[119]), .Z(n5746) );
  NAND U8448 ( .A(n5983), .B(x[119]), .Z(n5745) );
  NAND U8449 ( .A(n5746), .B(n5745), .Z(n1938) );
  NAND U8450 ( .A(n3857), .B(o[118]), .Z(n5748) );
  NAND U8451 ( .A(n5983), .B(x[118]), .Z(n5747) );
  NAND U8452 ( .A(n5748), .B(n5747), .Z(n1939) );
  NAND U8453 ( .A(n3857), .B(o[117]), .Z(n5750) );
  NAND U8454 ( .A(n5983), .B(x[117]), .Z(n5749) );
  NAND U8455 ( .A(n5750), .B(n5749), .Z(n1940) );
  NAND U8456 ( .A(n3857), .B(o[116]), .Z(n5752) );
  NAND U8457 ( .A(n5983), .B(x[116]), .Z(n5751) );
  NAND U8458 ( .A(n5752), .B(n5751), .Z(n1941) );
  NAND U8459 ( .A(n3857), .B(o[115]), .Z(n5754) );
  NAND U8460 ( .A(n5983), .B(x[115]), .Z(n5753) );
  NAND U8461 ( .A(n5754), .B(n5753), .Z(n1942) );
  NAND U8462 ( .A(n3857), .B(o[114]), .Z(n5756) );
  NAND U8463 ( .A(n5983), .B(x[114]), .Z(n5755) );
  NAND U8464 ( .A(n5756), .B(n5755), .Z(n1943) );
  NAND U8465 ( .A(n3857), .B(o[113]), .Z(n5758) );
  NAND U8466 ( .A(n5983), .B(x[113]), .Z(n5757) );
  NAND U8467 ( .A(n5758), .B(n5757), .Z(n1944) );
  NAND U8468 ( .A(n3857), .B(o[112]), .Z(n5760) );
  NAND U8469 ( .A(n5983), .B(x[112]), .Z(n5759) );
  NAND U8470 ( .A(n5760), .B(n5759), .Z(n1945) );
  NAND U8471 ( .A(n3857), .B(o[111]), .Z(n5762) );
  NAND U8472 ( .A(n5983), .B(x[111]), .Z(n5761) );
  NAND U8473 ( .A(n5762), .B(n5761), .Z(n1946) );
  NAND U8474 ( .A(n3857), .B(o[110]), .Z(n5764) );
  NAND U8475 ( .A(n5983), .B(x[110]), .Z(n5763) );
  NAND U8476 ( .A(n5764), .B(n5763), .Z(n1947) );
  NAND U8477 ( .A(n3857), .B(o[109]), .Z(n5766) );
  NAND U8478 ( .A(n5983), .B(x[109]), .Z(n5765) );
  NAND U8479 ( .A(n5766), .B(n5765), .Z(n1948) );
  NAND U8480 ( .A(n3857), .B(o[108]), .Z(n5768) );
  NAND U8481 ( .A(n5983), .B(x[108]), .Z(n5767) );
  NAND U8482 ( .A(n5768), .B(n5767), .Z(n1949) );
  NAND U8483 ( .A(n3857), .B(o[107]), .Z(n5770) );
  NAND U8484 ( .A(n5983), .B(x[107]), .Z(n5769) );
  NAND U8485 ( .A(n5770), .B(n5769), .Z(n1950) );
  NAND U8486 ( .A(n3857), .B(o[106]), .Z(n5772) );
  NAND U8487 ( .A(n5983), .B(x[106]), .Z(n5771) );
  NAND U8488 ( .A(n5772), .B(n5771), .Z(n1951) );
  NAND U8489 ( .A(n3857), .B(o[105]), .Z(n5774) );
  NAND U8490 ( .A(n5983), .B(x[105]), .Z(n5773) );
  NAND U8491 ( .A(n5774), .B(n5773), .Z(n1952) );
  NAND U8492 ( .A(n3857), .B(o[104]), .Z(n5776) );
  NAND U8493 ( .A(n5983), .B(x[104]), .Z(n5775) );
  NAND U8494 ( .A(n5776), .B(n5775), .Z(n1953) );
  NAND U8495 ( .A(n3857), .B(o[103]), .Z(n5778) );
  NAND U8496 ( .A(n5983), .B(x[103]), .Z(n5777) );
  NAND U8497 ( .A(n5778), .B(n5777), .Z(n1954) );
  NAND U8498 ( .A(n3857), .B(o[102]), .Z(n5780) );
  NAND U8499 ( .A(n5983), .B(x[102]), .Z(n5779) );
  NAND U8500 ( .A(n5780), .B(n5779), .Z(n1955) );
  NAND U8501 ( .A(n3857), .B(o[101]), .Z(n5782) );
  NAND U8502 ( .A(n5983), .B(x[101]), .Z(n5781) );
  NAND U8503 ( .A(n5782), .B(n5781), .Z(n1956) );
  NAND U8504 ( .A(n3857), .B(o[100]), .Z(n5784) );
  NAND U8505 ( .A(n5983), .B(x[100]), .Z(n5783) );
  NAND U8506 ( .A(n5784), .B(n5783), .Z(n1957) );
  NAND U8507 ( .A(n3857), .B(o[99]), .Z(n5786) );
  NAND U8508 ( .A(n5983), .B(x[99]), .Z(n5785) );
  NAND U8509 ( .A(n5786), .B(n5785), .Z(n1958) );
  NAND U8510 ( .A(n3857), .B(o[98]), .Z(n5788) );
  NAND U8511 ( .A(n5983), .B(x[98]), .Z(n5787) );
  NAND U8512 ( .A(n5788), .B(n5787), .Z(n1959) );
  NAND U8513 ( .A(n3857), .B(o[97]), .Z(n5790) );
  NAND U8514 ( .A(n5983), .B(x[97]), .Z(n5789) );
  NAND U8515 ( .A(n5790), .B(n5789), .Z(n1960) );
  NAND U8516 ( .A(n3857), .B(o[96]), .Z(n5792) );
  NAND U8517 ( .A(n5983), .B(x[96]), .Z(n5791) );
  NAND U8518 ( .A(n5792), .B(n5791), .Z(n1961) );
  NAND U8519 ( .A(n3857), .B(o[95]), .Z(n5794) );
  NAND U8520 ( .A(n5983), .B(x[95]), .Z(n5793) );
  NAND U8521 ( .A(n5794), .B(n5793), .Z(n1962) );
  NAND U8522 ( .A(n3857), .B(o[94]), .Z(n5796) );
  NAND U8523 ( .A(n5983), .B(x[94]), .Z(n5795) );
  NAND U8524 ( .A(n5796), .B(n5795), .Z(n1963) );
  NAND U8525 ( .A(n3857), .B(o[93]), .Z(n5798) );
  NAND U8526 ( .A(n5983), .B(x[93]), .Z(n5797) );
  NAND U8527 ( .A(n5798), .B(n5797), .Z(n1964) );
  NAND U8528 ( .A(n3857), .B(o[92]), .Z(n5800) );
  NAND U8529 ( .A(n5983), .B(x[92]), .Z(n5799) );
  NAND U8530 ( .A(n5800), .B(n5799), .Z(n1965) );
  NAND U8531 ( .A(n3857), .B(o[91]), .Z(n5802) );
  NAND U8532 ( .A(n5983), .B(x[91]), .Z(n5801) );
  NAND U8533 ( .A(n5802), .B(n5801), .Z(n1966) );
  NAND U8534 ( .A(n3857), .B(o[90]), .Z(n5804) );
  NAND U8535 ( .A(n5983), .B(x[90]), .Z(n5803) );
  NAND U8536 ( .A(n5804), .B(n5803), .Z(n1967) );
  NAND U8537 ( .A(n3857), .B(o[89]), .Z(n5806) );
  NAND U8538 ( .A(n5983), .B(x[89]), .Z(n5805) );
  NAND U8539 ( .A(n5806), .B(n5805), .Z(n1968) );
  NAND U8540 ( .A(n3857), .B(o[88]), .Z(n5808) );
  NAND U8541 ( .A(n5983), .B(x[88]), .Z(n5807) );
  NAND U8542 ( .A(n5808), .B(n5807), .Z(n1969) );
  NAND U8543 ( .A(n3857), .B(o[87]), .Z(n5810) );
  NAND U8544 ( .A(n5983), .B(x[87]), .Z(n5809) );
  NAND U8545 ( .A(n5810), .B(n5809), .Z(n1970) );
  NAND U8546 ( .A(n3857), .B(o[86]), .Z(n5812) );
  NAND U8547 ( .A(n5983), .B(x[86]), .Z(n5811) );
  NAND U8548 ( .A(n5812), .B(n5811), .Z(n1971) );
  NAND U8549 ( .A(n3857), .B(o[85]), .Z(n5814) );
  NAND U8550 ( .A(n5983), .B(x[85]), .Z(n5813) );
  NAND U8551 ( .A(n5814), .B(n5813), .Z(n1972) );
  NAND U8552 ( .A(n3857), .B(o[84]), .Z(n5816) );
  NAND U8553 ( .A(n5983), .B(x[84]), .Z(n5815) );
  NAND U8554 ( .A(n5816), .B(n5815), .Z(n1973) );
  NAND U8555 ( .A(n3857), .B(o[83]), .Z(n5818) );
  NAND U8556 ( .A(n5983), .B(x[83]), .Z(n5817) );
  NAND U8557 ( .A(n5818), .B(n5817), .Z(n1974) );
  NAND U8558 ( .A(n3857), .B(o[82]), .Z(n5820) );
  NAND U8559 ( .A(n5983), .B(x[82]), .Z(n5819) );
  NAND U8560 ( .A(n5820), .B(n5819), .Z(n1975) );
  NAND U8561 ( .A(n3857), .B(o[81]), .Z(n5822) );
  NAND U8562 ( .A(n5983), .B(x[81]), .Z(n5821) );
  NAND U8563 ( .A(n5822), .B(n5821), .Z(n1976) );
  NAND U8564 ( .A(n3857), .B(o[80]), .Z(n5824) );
  NAND U8565 ( .A(n5983), .B(x[80]), .Z(n5823) );
  NAND U8566 ( .A(n5824), .B(n5823), .Z(n1977) );
  NAND U8567 ( .A(n3857), .B(o[79]), .Z(n5826) );
  NAND U8568 ( .A(n5983), .B(x[79]), .Z(n5825) );
  NAND U8569 ( .A(n5826), .B(n5825), .Z(n1978) );
  NAND U8570 ( .A(n3857), .B(o[78]), .Z(n5828) );
  NAND U8571 ( .A(n5983), .B(x[78]), .Z(n5827) );
  NAND U8572 ( .A(n5828), .B(n5827), .Z(n1979) );
  NAND U8573 ( .A(n3857), .B(o[77]), .Z(n5830) );
  NAND U8574 ( .A(n5983), .B(x[77]), .Z(n5829) );
  NAND U8575 ( .A(n5830), .B(n5829), .Z(n1980) );
  NAND U8576 ( .A(n3857), .B(o[76]), .Z(n5832) );
  NAND U8577 ( .A(n5983), .B(x[76]), .Z(n5831) );
  NAND U8578 ( .A(n5832), .B(n5831), .Z(n1981) );
  NAND U8579 ( .A(n3857), .B(o[75]), .Z(n5834) );
  NAND U8580 ( .A(n5983), .B(x[75]), .Z(n5833) );
  NAND U8581 ( .A(n5834), .B(n5833), .Z(n1982) );
  NAND U8582 ( .A(n3857), .B(o[74]), .Z(n5836) );
  NAND U8583 ( .A(n5983), .B(x[74]), .Z(n5835) );
  NAND U8584 ( .A(n5836), .B(n5835), .Z(n1983) );
  NAND U8585 ( .A(n3857), .B(o[73]), .Z(n5838) );
  NAND U8586 ( .A(n5983), .B(x[73]), .Z(n5837) );
  NAND U8587 ( .A(n5838), .B(n5837), .Z(n1984) );
  NAND U8588 ( .A(n3857), .B(o[72]), .Z(n5840) );
  NAND U8589 ( .A(n5983), .B(x[72]), .Z(n5839) );
  NAND U8590 ( .A(n5840), .B(n5839), .Z(n1985) );
  NAND U8591 ( .A(n3857), .B(o[71]), .Z(n5842) );
  NAND U8592 ( .A(n5983), .B(x[71]), .Z(n5841) );
  NAND U8593 ( .A(n5842), .B(n5841), .Z(n1986) );
  NAND U8594 ( .A(n3857), .B(o[70]), .Z(n5844) );
  NAND U8595 ( .A(n5983), .B(x[70]), .Z(n5843) );
  NAND U8596 ( .A(n5844), .B(n5843), .Z(n1987) );
  NAND U8597 ( .A(n3857), .B(o[69]), .Z(n5846) );
  NAND U8598 ( .A(n5983), .B(x[69]), .Z(n5845) );
  NAND U8599 ( .A(n5846), .B(n5845), .Z(n1988) );
  NAND U8600 ( .A(n3857), .B(o[68]), .Z(n5848) );
  NAND U8601 ( .A(n5983), .B(x[68]), .Z(n5847) );
  NAND U8602 ( .A(n5848), .B(n5847), .Z(n1989) );
  NAND U8603 ( .A(n3857), .B(o[67]), .Z(n5850) );
  NAND U8604 ( .A(n5983), .B(x[67]), .Z(n5849) );
  NAND U8605 ( .A(n5850), .B(n5849), .Z(n1990) );
  NAND U8606 ( .A(n3857), .B(o[66]), .Z(n5852) );
  NAND U8607 ( .A(n5983), .B(x[66]), .Z(n5851) );
  NAND U8608 ( .A(n5852), .B(n5851), .Z(n1991) );
  NAND U8609 ( .A(n3857), .B(o[65]), .Z(n5854) );
  NAND U8610 ( .A(n5983), .B(x[65]), .Z(n5853) );
  NAND U8611 ( .A(n5854), .B(n5853), .Z(n1992) );
  NAND U8612 ( .A(n3857), .B(o[64]), .Z(n5856) );
  NAND U8613 ( .A(n5983), .B(x[64]), .Z(n5855) );
  NAND U8614 ( .A(n5856), .B(n5855), .Z(n1993) );
  NAND U8615 ( .A(n3857), .B(o[63]), .Z(n5858) );
  NAND U8616 ( .A(n5983), .B(x[63]), .Z(n5857) );
  NAND U8617 ( .A(n5858), .B(n5857), .Z(n1994) );
  NAND U8618 ( .A(n3857), .B(o[62]), .Z(n5860) );
  NAND U8619 ( .A(n5983), .B(x[62]), .Z(n5859) );
  NAND U8620 ( .A(n5860), .B(n5859), .Z(n1995) );
  NAND U8621 ( .A(n3857), .B(o[61]), .Z(n5862) );
  NAND U8622 ( .A(n5983), .B(x[61]), .Z(n5861) );
  NAND U8623 ( .A(n5862), .B(n5861), .Z(n1996) );
  NAND U8624 ( .A(n3857), .B(o[60]), .Z(n5864) );
  NAND U8625 ( .A(n5983), .B(x[60]), .Z(n5863) );
  NAND U8626 ( .A(n5864), .B(n5863), .Z(n1997) );
  NAND U8627 ( .A(n3857), .B(o[59]), .Z(n5866) );
  NAND U8628 ( .A(n5983), .B(x[59]), .Z(n5865) );
  NAND U8629 ( .A(n5866), .B(n5865), .Z(n1998) );
  NAND U8630 ( .A(n3857), .B(o[58]), .Z(n5868) );
  NAND U8631 ( .A(n5983), .B(x[58]), .Z(n5867) );
  NAND U8632 ( .A(n5868), .B(n5867), .Z(n1999) );
  NAND U8633 ( .A(n3857), .B(o[57]), .Z(n5870) );
  NAND U8634 ( .A(n5983), .B(x[57]), .Z(n5869) );
  NAND U8635 ( .A(n5870), .B(n5869), .Z(n2000) );
  NAND U8636 ( .A(n3857), .B(o[56]), .Z(n5872) );
  NAND U8637 ( .A(n5983), .B(x[56]), .Z(n5871) );
  NAND U8638 ( .A(n5872), .B(n5871), .Z(n2001) );
  NAND U8639 ( .A(n3857), .B(o[55]), .Z(n5874) );
  NAND U8640 ( .A(n5983), .B(x[55]), .Z(n5873) );
  NAND U8641 ( .A(n5874), .B(n5873), .Z(n2002) );
  NAND U8642 ( .A(n3857), .B(o[54]), .Z(n5876) );
  NAND U8643 ( .A(n5983), .B(x[54]), .Z(n5875) );
  NAND U8644 ( .A(n5876), .B(n5875), .Z(n2003) );
  NAND U8645 ( .A(n3857), .B(o[53]), .Z(n5878) );
  NAND U8646 ( .A(n5983), .B(x[53]), .Z(n5877) );
  NAND U8647 ( .A(n5878), .B(n5877), .Z(n2004) );
  NAND U8648 ( .A(n3857), .B(o[52]), .Z(n5880) );
  NAND U8649 ( .A(n5983), .B(x[52]), .Z(n5879) );
  NAND U8650 ( .A(n5880), .B(n5879), .Z(n2005) );
  NAND U8651 ( .A(n3857), .B(o[51]), .Z(n5882) );
  NAND U8652 ( .A(n5983), .B(x[51]), .Z(n5881) );
  NAND U8653 ( .A(n5882), .B(n5881), .Z(n2006) );
  NAND U8654 ( .A(n3857), .B(o[50]), .Z(n5884) );
  NAND U8655 ( .A(n5983), .B(x[50]), .Z(n5883) );
  NAND U8656 ( .A(n5884), .B(n5883), .Z(n2007) );
  NAND U8657 ( .A(n3857), .B(o[49]), .Z(n5886) );
  NAND U8658 ( .A(n5983), .B(x[49]), .Z(n5885) );
  NAND U8659 ( .A(n5886), .B(n5885), .Z(n2008) );
  NAND U8660 ( .A(n3857), .B(o[48]), .Z(n5888) );
  NAND U8661 ( .A(n5983), .B(x[48]), .Z(n5887) );
  NAND U8662 ( .A(n5888), .B(n5887), .Z(n2009) );
  NAND U8663 ( .A(n3857), .B(o[47]), .Z(n5890) );
  NAND U8664 ( .A(n5983), .B(x[47]), .Z(n5889) );
  NAND U8665 ( .A(n5890), .B(n5889), .Z(n2010) );
  NAND U8666 ( .A(n3857), .B(o[46]), .Z(n5892) );
  NAND U8667 ( .A(n5983), .B(x[46]), .Z(n5891) );
  NAND U8668 ( .A(n5892), .B(n5891), .Z(n2011) );
  NAND U8669 ( .A(n3857), .B(o[45]), .Z(n5894) );
  NAND U8670 ( .A(n5983), .B(x[45]), .Z(n5893) );
  NAND U8671 ( .A(n5894), .B(n5893), .Z(n2012) );
  NAND U8672 ( .A(n3857), .B(o[44]), .Z(n5896) );
  NAND U8673 ( .A(n5983), .B(x[44]), .Z(n5895) );
  NAND U8674 ( .A(n5896), .B(n5895), .Z(n2013) );
  NAND U8675 ( .A(n3857), .B(o[43]), .Z(n5898) );
  NAND U8676 ( .A(n5983), .B(x[43]), .Z(n5897) );
  NAND U8677 ( .A(n5898), .B(n5897), .Z(n2014) );
  NAND U8678 ( .A(n3857), .B(o[42]), .Z(n5900) );
  NAND U8679 ( .A(n5983), .B(x[42]), .Z(n5899) );
  NAND U8680 ( .A(n5900), .B(n5899), .Z(n2015) );
  NAND U8681 ( .A(n3857), .B(o[41]), .Z(n5902) );
  NAND U8682 ( .A(n5983), .B(x[41]), .Z(n5901) );
  NAND U8683 ( .A(n5902), .B(n5901), .Z(n2016) );
  NAND U8684 ( .A(n3857), .B(o[40]), .Z(n5904) );
  NAND U8685 ( .A(n5983), .B(x[40]), .Z(n5903) );
  NAND U8686 ( .A(n5904), .B(n5903), .Z(n2017) );
  NAND U8687 ( .A(n3857), .B(o[39]), .Z(n5906) );
  NAND U8688 ( .A(n5983), .B(x[39]), .Z(n5905) );
  NAND U8689 ( .A(n5906), .B(n5905), .Z(n2018) );
  NAND U8690 ( .A(n3857), .B(o[38]), .Z(n5908) );
  NAND U8691 ( .A(n5983), .B(x[38]), .Z(n5907) );
  NAND U8692 ( .A(n5908), .B(n5907), .Z(n2019) );
  NAND U8693 ( .A(n3857), .B(o[37]), .Z(n5910) );
  NAND U8694 ( .A(n5983), .B(x[37]), .Z(n5909) );
  NAND U8695 ( .A(n5910), .B(n5909), .Z(n2020) );
  NAND U8696 ( .A(n3857), .B(o[36]), .Z(n5912) );
  NAND U8697 ( .A(n5983), .B(x[36]), .Z(n5911) );
  NAND U8698 ( .A(n5912), .B(n5911), .Z(n2021) );
  NAND U8699 ( .A(n3857), .B(o[35]), .Z(n5914) );
  NAND U8700 ( .A(n5983), .B(x[35]), .Z(n5913) );
  NAND U8701 ( .A(n5914), .B(n5913), .Z(n2022) );
  NAND U8702 ( .A(n3857), .B(o[34]), .Z(n5916) );
  NAND U8703 ( .A(n5983), .B(x[34]), .Z(n5915) );
  NAND U8704 ( .A(n5916), .B(n5915), .Z(n2023) );
  NAND U8705 ( .A(n3857), .B(o[33]), .Z(n5918) );
  NAND U8706 ( .A(n5983), .B(x[33]), .Z(n5917) );
  NAND U8707 ( .A(n5918), .B(n5917), .Z(n2024) );
  NAND U8708 ( .A(n3857), .B(o[32]), .Z(n5920) );
  NAND U8709 ( .A(n5983), .B(x[32]), .Z(n5919) );
  NAND U8710 ( .A(n5920), .B(n5919), .Z(n2025) );
  NAND U8711 ( .A(n3857), .B(o[31]), .Z(n5922) );
  NAND U8712 ( .A(n5983), .B(x[31]), .Z(n5921) );
  NAND U8713 ( .A(n5922), .B(n5921), .Z(n2026) );
  NAND U8714 ( .A(n3857), .B(o[30]), .Z(n5924) );
  NAND U8715 ( .A(n5983), .B(x[30]), .Z(n5923) );
  NAND U8716 ( .A(n5924), .B(n5923), .Z(n2027) );
  NAND U8717 ( .A(n3857), .B(o[29]), .Z(n5926) );
  NAND U8718 ( .A(n5983), .B(x[29]), .Z(n5925) );
  NAND U8719 ( .A(n5926), .B(n5925), .Z(n2028) );
  NAND U8720 ( .A(n3857), .B(o[28]), .Z(n5928) );
  NAND U8721 ( .A(n5983), .B(x[28]), .Z(n5927) );
  NAND U8722 ( .A(n5928), .B(n5927), .Z(n2029) );
  NAND U8723 ( .A(n3857), .B(o[27]), .Z(n5930) );
  NAND U8724 ( .A(n5983), .B(x[27]), .Z(n5929) );
  NAND U8725 ( .A(n5930), .B(n5929), .Z(n2030) );
  NAND U8726 ( .A(n3857), .B(o[26]), .Z(n5932) );
  NAND U8727 ( .A(n5983), .B(x[26]), .Z(n5931) );
  NAND U8728 ( .A(n5932), .B(n5931), .Z(n2031) );
  NAND U8729 ( .A(n3857), .B(o[25]), .Z(n5934) );
  NAND U8730 ( .A(n5983), .B(x[25]), .Z(n5933) );
  NAND U8731 ( .A(n5934), .B(n5933), .Z(n2032) );
  NAND U8732 ( .A(n3857), .B(o[24]), .Z(n5936) );
  NAND U8733 ( .A(n5983), .B(x[24]), .Z(n5935) );
  NAND U8734 ( .A(n5936), .B(n5935), .Z(n2033) );
  NAND U8735 ( .A(n3857), .B(o[23]), .Z(n5938) );
  NAND U8736 ( .A(n5983), .B(x[23]), .Z(n5937) );
  NAND U8737 ( .A(n5938), .B(n5937), .Z(n2034) );
  NAND U8738 ( .A(n3857), .B(o[22]), .Z(n5940) );
  NAND U8739 ( .A(n5983), .B(x[22]), .Z(n5939) );
  NAND U8740 ( .A(n5940), .B(n5939), .Z(n2035) );
  NAND U8741 ( .A(n3857), .B(o[21]), .Z(n5942) );
  NAND U8742 ( .A(n5983), .B(x[21]), .Z(n5941) );
  NAND U8743 ( .A(n5942), .B(n5941), .Z(n2036) );
  NAND U8744 ( .A(n3857), .B(o[20]), .Z(n5944) );
  NAND U8745 ( .A(n5983), .B(x[20]), .Z(n5943) );
  NAND U8746 ( .A(n5944), .B(n5943), .Z(n2037) );
  NAND U8747 ( .A(n3857), .B(o[19]), .Z(n5946) );
  NAND U8748 ( .A(n5983), .B(x[19]), .Z(n5945) );
  NAND U8749 ( .A(n5946), .B(n5945), .Z(n2038) );
  NAND U8750 ( .A(n3857), .B(o[18]), .Z(n5948) );
  NAND U8751 ( .A(n5983), .B(x[18]), .Z(n5947) );
  NAND U8752 ( .A(n5948), .B(n5947), .Z(n2039) );
  NAND U8753 ( .A(n3857), .B(o[17]), .Z(n5950) );
  NAND U8754 ( .A(n5983), .B(x[17]), .Z(n5949) );
  NAND U8755 ( .A(n5950), .B(n5949), .Z(n2040) );
  NAND U8756 ( .A(n3857), .B(o[16]), .Z(n5952) );
  NAND U8757 ( .A(n5983), .B(x[16]), .Z(n5951) );
  NAND U8758 ( .A(n5952), .B(n5951), .Z(n2041) );
  NAND U8759 ( .A(n3857), .B(o[15]), .Z(n5954) );
  NAND U8760 ( .A(n5983), .B(x[15]), .Z(n5953) );
  NAND U8761 ( .A(n5954), .B(n5953), .Z(n2042) );
  NAND U8762 ( .A(n3857), .B(o[14]), .Z(n5956) );
  NAND U8763 ( .A(n5983), .B(x[14]), .Z(n5955) );
  NAND U8764 ( .A(n5956), .B(n5955), .Z(n2043) );
  NAND U8765 ( .A(n3857), .B(o[13]), .Z(n5958) );
  NAND U8766 ( .A(n5983), .B(x[13]), .Z(n5957) );
  NAND U8767 ( .A(n5958), .B(n5957), .Z(n2044) );
  NAND U8768 ( .A(n3857), .B(o[12]), .Z(n5960) );
  NAND U8769 ( .A(n5983), .B(x[12]), .Z(n5959) );
  NAND U8770 ( .A(n5960), .B(n5959), .Z(n2045) );
  NAND U8771 ( .A(n3857), .B(o[11]), .Z(n5962) );
  NAND U8772 ( .A(n5983), .B(x[11]), .Z(n5961) );
  NAND U8773 ( .A(n5962), .B(n5961), .Z(n2046) );
  NAND U8774 ( .A(n3857), .B(o[10]), .Z(n5964) );
  NAND U8775 ( .A(n5983), .B(x[10]), .Z(n5963) );
  NAND U8776 ( .A(n5964), .B(n5963), .Z(n2047) );
  NAND U8777 ( .A(n3857), .B(o[9]), .Z(n5966) );
  NAND U8778 ( .A(n5983), .B(x[9]), .Z(n5965) );
  NAND U8779 ( .A(n5966), .B(n5965), .Z(n2048) );
  NAND U8780 ( .A(n3857), .B(o[8]), .Z(n5968) );
  NAND U8781 ( .A(n5983), .B(x[8]), .Z(n5967) );
  NAND U8782 ( .A(n5968), .B(n5967), .Z(n2049) );
  NAND U8783 ( .A(n3857), .B(o[7]), .Z(n5970) );
  NAND U8784 ( .A(n5983), .B(x[7]), .Z(n5969) );
  NAND U8785 ( .A(n5970), .B(n5969), .Z(n2050) );
  NAND U8786 ( .A(n3857), .B(o[6]), .Z(n5972) );
  NAND U8787 ( .A(n5983), .B(x[6]), .Z(n5971) );
  NAND U8788 ( .A(n5972), .B(n5971), .Z(n2051) );
  NAND U8789 ( .A(n3857), .B(o[5]), .Z(n5974) );
  NAND U8790 ( .A(n5983), .B(x[5]), .Z(n5973) );
  NAND U8791 ( .A(n5974), .B(n5973), .Z(n2052) );
  NAND U8792 ( .A(n3857), .B(o[4]), .Z(n5976) );
  NAND U8793 ( .A(n5983), .B(x[4]), .Z(n5975) );
  NAND U8794 ( .A(n5976), .B(n5975), .Z(n2053) );
  NAND U8795 ( .A(n3857), .B(o[3]), .Z(n5978) );
  NAND U8796 ( .A(n5983), .B(x[3]), .Z(n5977) );
  NAND U8797 ( .A(n5978), .B(n5977), .Z(n2054) );
  NAND U8798 ( .A(n3857), .B(o[2]), .Z(n5980) );
  NAND U8799 ( .A(n5983), .B(x[2]), .Z(n5979) );
  NAND U8800 ( .A(n5980), .B(n5979), .Z(n2055) );
  NAND U8801 ( .A(n3857), .B(o[1]), .Z(n5982) );
  NAND U8802 ( .A(n5983), .B(x[1]), .Z(n5981) );
  NAND U8803 ( .A(n5982), .B(n5981), .Z(n2056) );
  NAND U8804 ( .A(n3857), .B(o[0]), .Z(n5985) );
  NAND U8805 ( .A(n5983), .B(x[0]), .Z(n5984) );
  NAND U8806 ( .A(n5985), .B(n5984), .Z(n2057) );
  ANDN U8807 ( .B(start_in[511]), .A(n5986), .Z(n7005) );
  NAND U8808 ( .A(n5987), .B(n7005), .Z(n5988) );
  NANDN U8809 ( .A(first_one), .B(n5988), .Z(n2058) );
  NAND U8810 ( .A(n7005), .B(ereg[254]), .Z(n5990) );
  OR U8811 ( .A(n7005), .B(n3896), .Z(n7010) );
  NANDN U8812 ( .A(n7010), .B(ereg[255]), .Z(n5989) );
  AND U8813 ( .A(n5990), .B(n5989), .Z(n5991) );
  NANDN U8814 ( .A(n5992), .B(n5991), .Z(n2059) );
  NAND U8815 ( .A(n7005), .B(ereg[253]), .Z(n5994) );
  NAND U8816 ( .A(n3896), .B(e[254]), .Z(n5993) );
  AND U8817 ( .A(n5994), .B(n5993), .Z(n5996) );
  NANDN U8818 ( .A(n7010), .B(ereg[254]), .Z(n5995) );
  NAND U8819 ( .A(n5996), .B(n5995), .Z(n2060) );
  NAND U8820 ( .A(n7005), .B(ereg[252]), .Z(n5998) );
  NAND U8821 ( .A(n3896), .B(e[253]), .Z(n5997) );
  AND U8822 ( .A(n5998), .B(n5997), .Z(n6000) );
  NANDN U8823 ( .A(n7010), .B(ereg[253]), .Z(n5999) );
  NAND U8824 ( .A(n6000), .B(n5999), .Z(n2061) );
  NAND U8825 ( .A(n7005), .B(ereg[251]), .Z(n6002) );
  NAND U8826 ( .A(n3896), .B(e[252]), .Z(n6001) );
  AND U8827 ( .A(n6002), .B(n6001), .Z(n6004) );
  NANDN U8828 ( .A(n7010), .B(ereg[252]), .Z(n6003) );
  NAND U8829 ( .A(n6004), .B(n6003), .Z(n2062) );
  NAND U8830 ( .A(n7005), .B(ereg[250]), .Z(n6006) );
  NAND U8831 ( .A(n3896), .B(e[251]), .Z(n6005) );
  AND U8832 ( .A(n6006), .B(n6005), .Z(n6008) );
  NANDN U8833 ( .A(n7010), .B(ereg[251]), .Z(n6007) );
  NAND U8834 ( .A(n6008), .B(n6007), .Z(n2063) );
  NAND U8835 ( .A(n7005), .B(ereg[249]), .Z(n6010) );
  NAND U8836 ( .A(n3896), .B(e[250]), .Z(n6009) );
  AND U8837 ( .A(n6010), .B(n6009), .Z(n6012) );
  NANDN U8838 ( .A(n7010), .B(ereg[250]), .Z(n6011) );
  NAND U8839 ( .A(n6012), .B(n6011), .Z(n2064) );
  NAND U8840 ( .A(n7005), .B(ereg[248]), .Z(n6014) );
  NAND U8841 ( .A(n3896), .B(e[249]), .Z(n6013) );
  AND U8842 ( .A(n6014), .B(n6013), .Z(n6016) );
  NANDN U8843 ( .A(n7010), .B(ereg[249]), .Z(n6015) );
  NAND U8844 ( .A(n6016), .B(n6015), .Z(n2065) );
  NAND U8845 ( .A(n7005), .B(ereg[247]), .Z(n6018) );
  NAND U8846 ( .A(n3897), .B(e[248]), .Z(n6017) );
  AND U8847 ( .A(n6018), .B(n6017), .Z(n6020) );
  NANDN U8848 ( .A(n7010), .B(ereg[248]), .Z(n6019) );
  NAND U8849 ( .A(n6020), .B(n6019), .Z(n2066) );
  NAND U8850 ( .A(n7005), .B(ereg[246]), .Z(n6022) );
  NAND U8851 ( .A(n3897), .B(e[247]), .Z(n6021) );
  AND U8852 ( .A(n6022), .B(n6021), .Z(n6024) );
  NANDN U8853 ( .A(n7010), .B(ereg[247]), .Z(n6023) );
  NAND U8854 ( .A(n6024), .B(n6023), .Z(n2067) );
  NAND U8855 ( .A(n7005), .B(ereg[245]), .Z(n6026) );
  NAND U8856 ( .A(n3897), .B(e[246]), .Z(n6025) );
  AND U8857 ( .A(n6026), .B(n6025), .Z(n6028) );
  NANDN U8858 ( .A(n7010), .B(ereg[246]), .Z(n6027) );
  NAND U8859 ( .A(n6028), .B(n6027), .Z(n2068) );
  NAND U8860 ( .A(n7005), .B(ereg[244]), .Z(n6030) );
  NAND U8861 ( .A(n3897), .B(e[245]), .Z(n6029) );
  AND U8862 ( .A(n6030), .B(n6029), .Z(n6032) );
  NANDN U8863 ( .A(n7010), .B(ereg[245]), .Z(n6031) );
  NAND U8864 ( .A(n6032), .B(n6031), .Z(n2069) );
  NAND U8865 ( .A(n7005), .B(ereg[243]), .Z(n6034) );
  NAND U8866 ( .A(n3897), .B(e[244]), .Z(n6033) );
  AND U8867 ( .A(n6034), .B(n6033), .Z(n6036) );
  NANDN U8868 ( .A(n7010), .B(ereg[244]), .Z(n6035) );
  NAND U8869 ( .A(n6036), .B(n6035), .Z(n2070) );
  NAND U8870 ( .A(n7005), .B(ereg[242]), .Z(n6038) );
  NAND U8871 ( .A(n3897), .B(e[243]), .Z(n6037) );
  AND U8872 ( .A(n6038), .B(n6037), .Z(n6040) );
  NANDN U8873 ( .A(n7010), .B(ereg[243]), .Z(n6039) );
  NAND U8874 ( .A(n6040), .B(n6039), .Z(n2071) );
  NAND U8875 ( .A(n7005), .B(ereg[241]), .Z(n6042) );
  NAND U8876 ( .A(n3897), .B(e[242]), .Z(n6041) );
  AND U8877 ( .A(n6042), .B(n6041), .Z(n6044) );
  NANDN U8878 ( .A(n7010), .B(ereg[242]), .Z(n6043) );
  NAND U8879 ( .A(n6044), .B(n6043), .Z(n2072) );
  NAND U8880 ( .A(n7005), .B(ereg[240]), .Z(n6046) );
  NAND U8881 ( .A(n3898), .B(e[241]), .Z(n6045) );
  AND U8882 ( .A(n6046), .B(n6045), .Z(n6048) );
  NANDN U8883 ( .A(n7010), .B(ereg[241]), .Z(n6047) );
  NAND U8884 ( .A(n6048), .B(n6047), .Z(n2073) );
  NAND U8885 ( .A(n7005), .B(ereg[239]), .Z(n6050) );
  NAND U8886 ( .A(n3898), .B(e[240]), .Z(n6049) );
  AND U8887 ( .A(n6050), .B(n6049), .Z(n6052) );
  NANDN U8888 ( .A(n7010), .B(ereg[240]), .Z(n6051) );
  NAND U8889 ( .A(n6052), .B(n6051), .Z(n2074) );
  NAND U8890 ( .A(n7005), .B(ereg[238]), .Z(n6054) );
  NAND U8891 ( .A(n3898), .B(e[239]), .Z(n6053) );
  AND U8892 ( .A(n6054), .B(n6053), .Z(n6056) );
  NANDN U8893 ( .A(n7010), .B(ereg[239]), .Z(n6055) );
  NAND U8894 ( .A(n6056), .B(n6055), .Z(n2075) );
  NAND U8895 ( .A(n7005), .B(ereg[237]), .Z(n6058) );
  NAND U8896 ( .A(n3898), .B(e[238]), .Z(n6057) );
  AND U8897 ( .A(n6058), .B(n6057), .Z(n6060) );
  NANDN U8898 ( .A(n7010), .B(ereg[238]), .Z(n6059) );
  NAND U8899 ( .A(n6060), .B(n6059), .Z(n2076) );
  NAND U8900 ( .A(n7005), .B(ereg[236]), .Z(n6062) );
  NAND U8901 ( .A(n3898), .B(e[237]), .Z(n6061) );
  AND U8902 ( .A(n6062), .B(n6061), .Z(n6064) );
  NANDN U8903 ( .A(n7010), .B(ereg[237]), .Z(n6063) );
  NAND U8904 ( .A(n6064), .B(n6063), .Z(n2077) );
  NAND U8905 ( .A(n7005), .B(ereg[235]), .Z(n6066) );
  NAND U8906 ( .A(n3898), .B(e[236]), .Z(n6065) );
  AND U8907 ( .A(n6066), .B(n6065), .Z(n6068) );
  NANDN U8908 ( .A(n7010), .B(ereg[236]), .Z(n6067) );
  NAND U8909 ( .A(n6068), .B(n6067), .Z(n2078) );
  NAND U8910 ( .A(n7005), .B(ereg[234]), .Z(n6070) );
  NAND U8911 ( .A(n3898), .B(e[235]), .Z(n6069) );
  AND U8912 ( .A(n6070), .B(n6069), .Z(n6072) );
  NANDN U8913 ( .A(n7010), .B(ereg[235]), .Z(n6071) );
  NAND U8914 ( .A(n6072), .B(n6071), .Z(n2079) );
  NAND U8915 ( .A(n7005), .B(ereg[233]), .Z(n6074) );
  NAND U8916 ( .A(n3899), .B(e[234]), .Z(n6073) );
  AND U8917 ( .A(n6074), .B(n6073), .Z(n6076) );
  NANDN U8918 ( .A(n7010), .B(ereg[234]), .Z(n6075) );
  NAND U8919 ( .A(n6076), .B(n6075), .Z(n2080) );
  NAND U8920 ( .A(n7005), .B(ereg[232]), .Z(n6078) );
  NAND U8921 ( .A(n3899), .B(e[233]), .Z(n6077) );
  AND U8922 ( .A(n6078), .B(n6077), .Z(n6080) );
  NANDN U8923 ( .A(n7010), .B(ereg[233]), .Z(n6079) );
  NAND U8924 ( .A(n6080), .B(n6079), .Z(n2081) );
  NAND U8925 ( .A(n7005), .B(ereg[231]), .Z(n6082) );
  NAND U8926 ( .A(n3899), .B(e[232]), .Z(n6081) );
  AND U8927 ( .A(n6082), .B(n6081), .Z(n6084) );
  NANDN U8928 ( .A(n7010), .B(ereg[232]), .Z(n6083) );
  NAND U8929 ( .A(n6084), .B(n6083), .Z(n2082) );
  NAND U8930 ( .A(n7005), .B(ereg[230]), .Z(n6086) );
  NAND U8931 ( .A(n3899), .B(e[231]), .Z(n6085) );
  AND U8932 ( .A(n6086), .B(n6085), .Z(n6088) );
  NANDN U8933 ( .A(n7010), .B(ereg[231]), .Z(n6087) );
  NAND U8934 ( .A(n6088), .B(n6087), .Z(n2083) );
  NAND U8935 ( .A(n7005), .B(ereg[229]), .Z(n6090) );
  NAND U8936 ( .A(n3899), .B(e[230]), .Z(n6089) );
  AND U8937 ( .A(n6090), .B(n6089), .Z(n6092) );
  NANDN U8938 ( .A(n7010), .B(ereg[230]), .Z(n6091) );
  NAND U8939 ( .A(n6092), .B(n6091), .Z(n2084) );
  NAND U8940 ( .A(n7005), .B(ereg[228]), .Z(n6094) );
  NAND U8941 ( .A(n3899), .B(e[229]), .Z(n6093) );
  AND U8942 ( .A(n6094), .B(n6093), .Z(n6096) );
  NANDN U8943 ( .A(n7010), .B(ereg[229]), .Z(n6095) );
  NAND U8944 ( .A(n6096), .B(n6095), .Z(n2085) );
  NAND U8945 ( .A(n7005), .B(ereg[227]), .Z(n6098) );
  NAND U8946 ( .A(n3899), .B(e[228]), .Z(n6097) );
  AND U8947 ( .A(n6098), .B(n6097), .Z(n6100) );
  NANDN U8948 ( .A(n7010), .B(ereg[228]), .Z(n6099) );
  NAND U8949 ( .A(n6100), .B(n6099), .Z(n2086) );
  NAND U8950 ( .A(n7005), .B(ereg[226]), .Z(n6102) );
  NAND U8951 ( .A(n3900), .B(e[227]), .Z(n6101) );
  AND U8952 ( .A(n6102), .B(n6101), .Z(n6104) );
  NANDN U8953 ( .A(n7010), .B(ereg[227]), .Z(n6103) );
  NAND U8954 ( .A(n6104), .B(n6103), .Z(n2087) );
  NAND U8955 ( .A(n7005), .B(ereg[225]), .Z(n6106) );
  NAND U8956 ( .A(n3900), .B(e[226]), .Z(n6105) );
  AND U8957 ( .A(n6106), .B(n6105), .Z(n6108) );
  NANDN U8958 ( .A(n7010), .B(ereg[226]), .Z(n6107) );
  NAND U8959 ( .A(n6108), .B(n6107), .Z(n2088) );
  NAND U8960 ( .A(n7005), .B(ereg[224]), .Z(n6110) );
  NAND U8961 ( .A(n3900), .B(e[225]), .Z(n6109) );
  AND U8962 ( .A(n6110), .B(n6109), .Z(n6112) );
  NANDN U8963 ( .A(n7010), .B(ereg[225]), .Z(n6111) );
  NAND U8964 ( .A(n6112), .B(n6111), .Z(n2089) );
  NAND U8965 ( .A(n7005), .B(ereg[223]), .Z(n6114) );
  NAND U8966 ( .A(n3900), .B(e[224]), .Z(n6113) );
  AND U8967 ( .A(n6114), .B(n6113), .Z(n6116) );
  NANDN U8968 ( .A(n7010), .B(ereg[224]), .Z(n6115) );
  NAND U8969 ( .A(n6116), .B(n6115), .Z(n2090) );
  NAND U8970 ( .A(n7005), .B(ereg[222]), .Z(n6118) );
  NAND U8971 ( .A(n3900), .B(e[223]), .Z(n6117) );
  AND U8972 ( .A(n6118), .B(n6117), .Z(n6120) );
  NANDN U8973 ( .A(n7010), .B(ereg[223]), .Z(n6119) );
  NAND U8974 ( .A(n6120), .B(n6119), .Z(n2091) );
  NAND U8975 ( .A(n7005), .B(ereg[221]), .Z(n6122) );
  NAND U8976 ( .A(n3900), .B(e[222]), .Z(n6121) );
  AND U8977 ( .A(n6122), .B(n6121), .Z(n6124) );
  NANDN U8978 ( .A(n7010), .B(ereg[222]), .Z(n6123) );
  NAND U8979 ( .A(n6124), .B(n6123), .Z(n2092) );
  NAND U8980 ( .A(n7005), .B(ereg[220]), .Z(n6126) );
  NAND U8981 ( .A(n3900), .B(e[221]), .Z(n6125) );
  AND U8982 ( .A(n6126), .B(n6125), .Z(n6128) );
  NANDN U8983 ( .A(n7010), .B(ereg[221]), .Z(n6127) );
  NAND U8984 ( .A(n6128), .B(n6127), .Z(n2093) );
  NAND U8985 ( .A(n7005), .B(ereg[219]), .Z(n6130) );
  NAND U8986 ( .A(n3901), .B(e[220]), .Z(n6129) );
  AND U8987 ( .A(n6130), .B(n6129), .Z(n6132) );
  NANDN U8988 ( .A(n7010), .B(ereg[220]), .Z(n6131) );
  NAND U8989 ( .A(n6132), .B(n6131), .Z(n2094) );
  NAND U8990 ( .A(n7005), .B(ereg[218]), .Z(n6134) );
  NAND U8991 ( .A(n3901), .B(e[219]), .Z(n6133) );
  AND U8992 ( .A(n6134), .B(n6133), .Z(n6136) );
  NANDN U8993 ( .A(n7010), .B(ereg[219]), .Z(n6135) );
  NAND U8994 ( .A(n6136), .B(n6135), .Z(n2095) );
  NAND U8995 ( .A(n7005), .B(ereg[217]), .Z(n6138) );
  NAND U8996 ( .A(n3901), .B(e[218]), .Z(n6137) );
  AND U8997 ( .A(n6138), .B(n6137), .Z(n6140) );
  NANDN U8998 ( .A(n7010), .B(ereg[218]), .Z(n6139) );
  NAND U8999 ( .A(n6140), .B(n6139), .Z(n2096) );
  NAND U9000 ( .A(n7005), .B(ereg[216]), .Z(n6142) );
  NAND U9001 ( .A(n3901), .B(e[217]), .Z(n6141) );
  AND U9002 ( .A(n6142), .B(n6141), .Z(n6144) );
  NANDN U9003 ( .A(n7010), .B(ereg[217]), .Z(n6143) );
  NAND U9004 ( .A(n6144), .B(n6143), .Z(n2097) );
  NAND U9005 ( .A(n7005), .B(ereg[215]), .Z(n6146) );
  NAND U9006 ( .A(n3901), .B(e[216]), .Z(n6145) );
  AND U9007 ( .A(n6146), .B(n6145), .Z(n6148) );
  NANDN U9008 ( .A(n7010), .B(ereg[216]), .Z(n6147) );
  NAND U9009 ( .A(n6148), .B(n6147), .Z(n2098) );
  NAND U9010 ( .A(n7005), .B(ereg[214]), .Z(n6150) );
  NAND U9011 ( .A(n3901), .B(e[215]), .Z(n6149) );
  AND U9012 ( .A(n6150), .B(n6149), .Z(n6152) );
  NANDN U9013 ( .A(n7010), .B(ereg[215]), .Z(n6151) );
  NAND U9014 ( .A(n6152), .B(n6151), .Z(n2099) );
  NAND U9015 ( .A(n7005), .B(ereg[213]), .Z(n6154) );
  NAND U9016 ( .A(n3901), .B(e[214]), .Z(n6153) );
  AND U9017 ( .A(n6154), .B(n6153), .Z(n6156) );
  NANDN U9018 ( .A(n7010), .B(ereg[214]), .Z(n6155) );
  NAND U9019 ( .A(n6156), .B(n6155), .Z(n2100) );
  NAND U9020 ( .A(n7005), .B(ereg[212]), .Z(n6158) );
  NAND U9021 ( .A(n3902), .B(e[213]), .Z(n6157) );
  AND U9022 ( .A(n6158), .B(n6157), .Z(n6160) );
  NANDN U9023 ( .A(n7010), .B(ereg[213]), .Z(n6159) );
  NAND U9024 ( .A(n6160), .B(n6159), .Z(n2101) );
  NAND U9025 ( .A(n7005), .B(ereg[211]), .Z(n6162) );
  NAND U9026 ( .A(n3902), .B(e[212]), .Z(n6161) );
  AND U9027 ( .A(n6162), .B(n6161), .Z(n6164) );
  NANDN U9028 ( .A(n7010), .B(ereg[212]), .Z(n6163) );
  NAND U9029 ( .A(n6164), .B(n6163), .Z(n2102) );
  NAND U9030 ( .A(n7005), .B(ereg[210]), .Z(n6166) );
  NAND U9031 ( .A(n3902), .B(e[211]), .Z(n6165) );
  AND U9032 ( .A(n6166), .B(n6165), .Z(n6168) );
  NANDN U9033 ( .A(n7010), .B(ereg[211]), .Z(n6167) );
  NAND U9034 ( .A(n6168), .B(n6167), .Z(n2103) );
  NAND U9035 ( .A(n7005), .B(ereg[209]), .Z(n6170) );
  NAND U9036 ( .A(n3902), .B(e[210]), .Z(n6169) );
  AND U9037 ( .A(n6170), .B(n6169), .Z(n6172) );
  NANDN U9038 ( .A(n7010), .B(ereg[210]), .Z(n6171) );
  NAND U9039 ( .A(n6172), .B(n6171), .Z(n2104) );
  NAND U9040 ( .A(n7005), .B(ereg[208]), .Z(n6174) );
  NAND U9041 ( .A(n3902), .B(e[209]), .Z(n6173) );
  AND U9042 ( .A(n6174), .B(n6173), .Z(n6176) );
  NANDN U9043 ( .A(n7010), .B(ereg[209]), .Z(n6175) );
  NAND U9044 ( .A(n6176), .B(n6175), .Z(n2105) );
  NAND U9045 ( .A(n7005), .B(ereg[207]), .Z(n6178) );
  NAND U9046 ( .A(n3902), .B(e[208]), .Z(n6177) );
  AND U9047 ( .A(n6178), .B(n6177), .Z(n6180) );
  NANDN U9048 ( .A(n7010), .B(ereg[208]), .Z(n6179) );
  NAND U9049 ( .A(n6180), .B(n6179), .Z(n2106) );
  NAND U9050 ( .A(n7005), .B(ereg[206]), .Z(n6182) );
  NAND U9051 ( .A(n3902), .B(e[207]), .Z(n6181) );
  AND U9052 ( .A(n6182), .B(n6181), .Z(n6184) );
  NANDN U9053 ( .A(n7010), .B(ereg[207]), .Z(n6183) );
  NAND U9054 ( .A(n6184), .B(n6183), .Z(n2107) );
  NAND U9055 ( .A(n7005), .B(ereg[205]), .Z(n6186) );
  NAND U9056 ( .A(n3903), .B(e[206]), .Z(n6185) );
  AND U9057 ( .A(n6186), .B(n6185), .Z(n6188) );
  NANDN U9058 ( .A(n7010), .B(ereg[206]), .Z(n6187) );
  NAND U9059 ( .A(n6188), .B(n6187), .Z(n2108) );
  NAND U9060 ( .A(n7005), .B(ereg[204]), .Z(n6190) );
  NAND U9061 ( .A(n3903), .B(e[205]), .Z(n6189) );
  AND U9062 ( .A(n6190), .B(n6189), .Z(n6192) );
  NANDN U9063 ( .A(n7010), .B(ereg[205]), .Z(n6191) );
  NAND U9064 ( .A(n6192), .B(n6191), .Z(n2109) );
  NAND U9065 ( .A(n7005), .B(ereg[203]), .Z(n6194) );
  NAND U9066 ( .A(n3903), .B(e[204]), .Z(n6193) );
  AND U9067 ( .A(n6194), .B(n6193), .Z(n6196) );
  NANDN U9068 ( .A(n7010), .B(ereg[204]), .Z(n6195) );
  NAND U9069 ( .A(n6196), .B(n6195), .Z(n2110) );
  NAND U9070 ( .A(n7005), .B(ereg[202]), .Z(n6198) );
  NAND U9071 ( .A(n3903), .B(e[203]), .Z(n6197) );
  AND U9072 ( .A(n6198), .B(n6197), .Z(n6200) );
  NANDN U9073 ( .A(n7010), .B(ereg[203]), .Z(n6199) );
  NAND U9074 ( .A(n6200), .B(n6199), .Z(n2111) );
  NAND U9075 ( .A(n7005), .B(ereg[201]), .Z(n6202) );
  NAND U9076 ( .A(n3903), .B(e[202]), .Z(n6201) );
  AND U9077 ( .A(n6202), .B(n6201), .Z(n6204) );
  NANDN U9078 ( .A(n7010), .B(ereg[202]), .Z(n6203) );
  NAND U9079 ( .A(n6204), .B(n6203), .Z(n2112) );
  NAND U9080 ( .A(n7005), .B(ereg[200]), .Z(n6206) );
  NAND U9081 ( .A(n3903), .B(e[201]), .Z(n6205) );
  AND U9082 ( .A(n6206), .B(n6205), .Z(n6208) );
  NANDN U9083 ( .A(n7010), .B(ereg[201]), .Z(n6207) );
  NAND U9084 ( .A(n6208), .B(n6207), .Z(n2113) );
  NAND U9085 ( .A(n7005), .B(ereg[199]), .Z(n6210) );
  NAND U9086 ( .A(n3903), .B(e[200]), .Z(n6209) );
  AND U9087 ( .A(n6210), .B(n6209), .Z(n6212) );
  NANDN U9088 ( .A(n7010), .B(ereg[200]), .Z(n6211) );
  NAND U9089 ( .A(n6212), .B(n6211), .Z(n2114) );
  NAND U9090 ( .A(n7005), .B(ereg[198]), .Z(n6214) );
  NAND U9091 ( .A(n3904), .B(e[199]), .Z(n6213) );
  AND U9092 ( .A(n6214), .B(n6213), .Z(n6216) );
  NANDN U9093 ( .A(n7010), .B(ereg[199]), .Z(n6215) );
  NAND U9094 ( .A(n6216), .B(n6215), .Z(n2115) );
  NAND U9095 ( .A(n7005), .B(ereg[197]), .Z(n6218) );
  NAND U9096 ( .A(n3904), .B(e[198]), .Z(n6217) );
  AND U9097 ( .A(n6218), .B(n6217), .Z(n6220) );
  NANDN U9098 ( .A(n7010), .B(ereg[198]), .Z(n6219) );
  NAND U9099 ( .A(n6220), .B(n6219), .Z(n2116) );
  NAND U9100 ( .A(n7005), .B(ereg[196]), .Z(n6222) );
  NAND U9101 ( .A(n3904), .B(e[197]), .Z(n6221) );
  AND U9102 ( .A(n6222), .B(n6221), .Z(n6224) );
  NANDN U9103 ( .A(n7010), .B(ereg[197]), .Z(n6223) );
  NAND U9104 ( .A(n6224), .B(n6223), .Z(n2117) );
  NAND U9105 ( .A(n7005), .B(ereg[195]), .Z(n6226) );
  NAND U9106 ( .A(n3904), .B(e[196]), .Z(n6225) );
  AND U9107 ( .A(n6226), .B(n6225), .Z(n6228) );
  NANDN U9108 ( .A(n7010), .B(ereg[196]), .Z(n6227) );
  NAND U9109 ( .A(n6228), .B(n6227), .Z(n2118) );
  NAND U9110 ( .A(n7005), .B(ereg[194]), .Z(n6230) );
  NAND U9111 ( .A(n3904), .B(e[195]), .Z(n6229) );
  AND U9112 ( .A(n6230), .B(n6229), .Z(n6232) );
  NANDN U9113 ( .A(n7010), .B(ereg[195]), .Z(n6231) );
  NAND U9114 ( .A(n6232), .B(n6231), .Z(n2119) );
  NAND U9115 ( .A(n7005), .B(ereg[193]), .Z(n6234) );
  NAND U9116 ( .A(n3904), .B(e[194]), .Z(n6233) );
  AND U9117 ( .A(n6234), .B(n6233), .Z(n6236) );
  NANDN U9118 ( .A(n7010), .B(ereg[194]), .Z(n6235) );
  NAND U9119 ( .A(n6236), .B(n6235), .Z(n2120) );
  NAND U9120 ( .A(n7005), .B(ereg[192]), .Z(n6238) );
  NAND U9121 ( .A(n3904), .B(e[193]), .Z(n6237) );
  AND U9122 ( .A(n6238), .B(n6237), .Z(n6240) );
  NANDN U9123 ( .A(n7010), .B(ereg[193]), .Z(n6239) );
  NAND U9124 ( .A(n6240), .B(n6239), .Z(n2121) );
  NAND U9125 ( .A(n7005), .B(ereg[191]), .Z(n6242) );
  NAND U9126 ( .A(n3905), .B(e[192]), .Z(n6241) );
  AND U9127 ( .A(n6242), .B(n6241), .Z(n6244) );
  NANDN U9128 ( .A(n7010), .B(ereg[192]), .Z(n6243) );
  NAND U9129 ( .A(n6244), .B(n6243), .Z(n2122) );
  NAND U9130 ( .A(n7005), .B(ereg[190]), .Z(n6246) );
  NAND U9131 ( .A(n3905), .B(e[191]), .Z(n6245) );
  AND U9132 ( .A(n6246), .B(n6245), .Z(n6248) );
  NANDN U9133 ( .A(n7010), .B(ereg[191]), .Z(n6247) );
  NAND U9134 ( .A(n6248), .B(n6247), .Z(n2123) );
  NAND U9135 ( .A(n7005), .B(ereg[189]), .Z(n6250) );
  NAND U9136 ( .A(n3905), .B(e[190]), .Z(n6249) );
  AND U9137 ( .A(n6250), .B(n6249), .Z(n6252) );
  NANDN U9138 ( .A(n7010), .B(ereg[190]), .Z(n6251) );
  NAND U9139 ( .A(n6252), .B(n6251), .Z(n2124) );
  NAND U9140 ( .A(n7005), .B(ereg[188]), .Z(n6254) );
  NAND U9141 ( .A(n3905), .B(e[189]), .Z(n6253) );
  AND U9142 ( .A(n6254), .B(n6253), .Z(n6256) );
  NANDN U9143 ( .A(n7010), .B(ereg[189]), .Z(n6255) );
  NAND U9144 ( .A(n6256), .B(n6255), .Z(n2125) );
  NAND U9145 ( .A(n7005), .B(ereg[187]), .Z(n6258) );
  NAND U9146 ( .A(n3905), .B(e[188]), .Z(n6257) );
  AND U9147 ( .A(n6258), .B(n6257), .Z(n6260) );
  NANDN U9148 ( .A(n7010), .B(ereg[188]), .Z(n6259) );
  NAND U9149 ( .A(n6260), .B(n6259), .Z(n2126) );
  NAND U9150 ( .A(n7005), .B(ereg[186]), .Z(n6262) );
  NAND U9151 ( .A(n3905), .B(e[187]), .Z(n6261) );
  AND U9152 ( .A(n6262), .B(n6261), .Z(n6264) );
  NANDN U9153 ( .A(n7010), .B(ereg[187]), .Z(n6263) );
  NAND U9154 ( .A(n6264), .B(n6263), .Z(n2127) );
  NAND U9155 ( .A(n7005), .B(ereg[185]), .Z(n6266) );
  NAND U9156 ( .A(n3905), .B(e[186]), .Z(n6265) );
  AND U9157 ( .A(n6266), .B(n6265), .Z(n6268) );
  NANDN U9158 ( .A(n7010), .B(ereg[186]), .Z(n6267) );
  NAND U9159 ( .A(n6268), .B(n6267), .Z(n2128) );
  NAND U9160 ( .A(n7005), .B(ereg[184]), .Z(n6270) );
  NAND U9161 ( .A(n3906), .B(e[185]), .Z(n6269) );
  AND U9162 ( .A(n6270), .B(n6269), .Z(n6272) );
  NANDN U9163 ( .A(n7010), .B(ereg[185]), .Z(n6271) );
  NAND U9164 ( .A(n6272), .B(n6271), .Z(n2129) );
  NAND U9165 ( .A(n7005), .B(ereg[183]), .Z(n6274) );
  NAND U9166 ( .A(n3906), .B(e[184]), .Z(n6273) );
  AND U9167 ( .A(n6274), .B(n6273), .Z(n6276) );
  NANDN U9168 ( .A(n7010), .B(ereg[184]), .Z(n6275) );
  NAND U9169 ( .A(n6276), .B(n6275), .Z(n2130) );
  NAND U9170 ( .A(n7005), .B(ereg[182]), .Z(n6278) );
  NAND U9171 ( .A(n3906), .B(e[183]), .Z(n6277) );
  AND U9172 ( .A(n6278), .B(n6277), .Z(n6280) );
  NANDN U9173 ( .A(n7010), .B(ereg[183]), .Z(n6279) );
  NAND U9174 ( .A(n6280), .B(n6279), .Z(n2131) );
  NAND U9175 ( .A(n7005), .B(ereg[181]), .Z(n6282) );
  NAND U9176 ( .A(n3906), .B(e[182]), .Z(n6281) );
  AND U9177 ( .A(n6282), .B(n6281), .Z(n6284) );
  NANDN U9178 ( .A(n7010), .B(ereg[182]), .Z(n6283) );
  NAND U9179 ( .A(n6284), .B(n6283), .Z(n2132) );
  NAND U9180 ( .A(n7005), .B(ereg[180]), .Z(n6286) );
  NAND U9181 ( .A(n3906), .B(e[181]), .Z(n6285) );
  AND U9182 ( .A(n6286), .B(n6285), .Z(n6288) );
  NANDN U9183 ( .A(n7010), .B(ereg[181]), .Z(n6287) );
  NAND U9184 ( .A(n6288), .B(n6287), .Z(n2133) );
  NAND U9185 ( .A(n7005), .B(ereg[179]), .Z(n6290) );
  NAND U9186 ( .A(n3906), .B(e[180]), .Z(n6289) );
  AND U9187 ( .A(n6290), .B(n6289), .Z(n6292) );
  NANDN U9188 ( .A(n7010), .B(ereg[180]), .Z(n6291) );
  NAND U9189 ( .A(n6292), .B(n6291), .Z(n2134) );
  NAND U9190 ( .A(n7005), .B(ereg[178]), .Z(n6294) );
  NAND U9191 ( .A(n3906), .B(e[179]), .Z(n6293) );
  AND U9192 ( .A(n6294), .B(n6293), .Z(n6296) );
  NANDN U9193 ( .A(n7010), .B(ereg[179]), .Z(n6295) );
  NAND U9194 ( .A(n6296), .B(n6295), .Z(n2135) );
  NAND U9195 ( .A(n7005), .B(ereg[177]), .Z(n6298) );
  NAND U9196 ( .A(n3907), .B(e[178]), .Z(n6297) );
  AND U9197 ( .A(n6298), .B(n6297), .Z(n6300) );
  NANDN U9198 ( .A(n7010), .B(ereg[178]), .Z(n6299) );
  NAND U9199 ( .A(n6300), .B(n6299), .Z(n2136) );
  NAND U9200 ( .A(n7005), .B(ereg[176]), .Z(n6302) );
  NAND U9201 ( .A(n3907), .B(e[177]), .Z(n6301) );
  AND U9202 ( .A(n6302), .B(n6301), .Z(n6304) );
  NANDN U9203 ( .A(n7010), .B(ereg[177]), .Z(n6303) );
  NAND U9204 ( .A(n6304), .B(n6303), .Z(n2137) );
  NAND U9205 ( .A(n7005), .B(ereg[175]), .Z(n6306) );
  NAND U9206 ( .A(n3907), .B(e[176]), .Z(n6305) );
  AND U9207 ( .A(n6306), .B(n6305), .Z(n6308) );
  NANDN U9208 ( .A(n7010), .B(ereg[176]), .Z(n6307) );
  NAND U9209 ( .A(n6308), .B(n6307), .Z(n2138) );
  NAND U9210 ( .A(n7005), .B(ereg[174]), .Z(n6310) );
  NAND U9211 ( .A(n3907), .B(e[175]), .Z(n6309) );
  AND U9212 ( .A(n6310), .B(n6309), .Z(n6312) );
  NANDN U9213 ( .A(n7010), .B(ereg[175]), .Z(n6311) );
  NAND U9214 ( .A(n6312), .B(n6311), .Z(n2139) );
  NAND U9215 ( .A(n7005), .B(ereg[173]), .Z(n6314) );
  NAND U9216 ( .A(n3907), .B(e[174]), .Z(n6313) );
  AND U9217 ( .A(n6314), .B(n6313), .Z(n6316) );
  NANDN U9218 ( .A(n7010), .B(ereg[174]), .Z(n6315) );
  NAND U9219 ( .A(n6316), .B(n6315), .Z(n2140) );
  NAND U9220 ( .A(n7005), .B(ereg[172]), .Z(n6318) );
  NAND U9221 ( .A(n3907), .B(e[173]), .Z(n6317) );
  AND U9222 ( .A(n6318), .B(n6317), .Z(n6320) );
  NANDN U9223 ( .A(n7010), .B(ereg[173]), .Z(n6319) );
  NAND U9224 ( .A(n6320), .B(n6319), .Z(n2141) );
  NAND U9225 ( .A(n7005), .B(ereg[171]), .Z(n6322) );
  NAND U9226 ( .A(n3907), .B(e[172]), .Z(n6321) );
  AND U9227 ( .A(n6322), .B(n6321), .Z(n6324) );
  NANDN U9228 ( .A(n7010), .B(ereg[172]), .Z(n6323) );
  NAND U9229 ( .A(n6324), .B(n6323), .Z(n2142) );
  NAND U9230 ( .A(n7005), .B(ereg[170]), .Z(n6326) );
  NAND U9231 ( .A(n3908), .B(e[171]), .Z(n6325) );
  AND U9232 ( .A(n6326), .B(n6325), .Z(n6328) );
  NANDN U9233 ( .A(n7010), .B(ereg[171]), .Z(n6327) );
  NAND U9234 ( .A(n6328), .B(n6327), .Z(n2143) );
  NAND U9235 ( .A(n7005), .B(ereg[169]), .Z(n6330) );
  NAND U9236 ( .A(n3908), .B(e[170]), .Z(n6329) );
  AND U9237 ( .A(n6330), .B(n6329), .Z(n6332) );
  NANDN U9238 ( .A(n7010), .B(ereg[170]), .Z(n6331) );
  NAND U9239 ( .A(n6332), .B(n6331), .Z(n2144) );
  NAND U9240 ( .A(n7005), .B(ereg[168]), .Z(n6334) );
  NAND U9241 ( .A(n3908), .B(e[169]), .Z(n6333) );
  AND U9242 ( .A(n6334), .B(n6333), .Z(n6336) );
  NANDN U9243 ( .A(n7010), .B(ereg[169]), .Z(n6335) );
  NAND U9244 ( .A(n6336), .B(n6335), .Z(n2145) );
  NAND U9245 ( .A(n7005), .B(ereg[167]), .Z(n6338) );
  NAND U9246 ( .A(n3908), .B(e[168]), .Z(n6337) );
  AND U9247 ( .A(n6338), .B(n6337), .Z(n6340) );
  NANDN U9248 ( .A(n7010), .B(ereg[168]), .Z(n6339) );
  NAND U9249 ( .A(n6340), .B(n6339), .Z(n2146) );
  NAND U9250 ( .A(n7005), .B(ereg[166]), .Z(n6342) );
  NAND U9251 ( .A(n3908), .B(e[167]), .Z(n6341) );
  AND U9252 ( .A(n6342), .B(n6341), .Z(n6344) );
  NANDN U9253 ( .A(n7010), .B(ereg[167]), .Z(n6343) );
  NAND U9254 ( .A(n6344), .B(n6343), .Z(n2147) );
  NAND U9255 ( .A(n7005), .B(ereg[165]), .Z(n6346) );
  NAND U9256 ( .A(n3908), .B(e[166]), .Z(n6345) );
  AND U9257 ( .A(n6346), .B(n6345), .Z(n6348) );
  NANDN U9258 ( .A(n7010), .B(ereg[166]), .Z(n6347) );
  NAND U9259 ( .A(n6348), .B(n6347), .Z(n2148) );
  NAND U9260 ( .A(n7005), .B(ereg[164]), .Z(n6350) );
  NAND U9261 ( .A(n3908), .B(e[165]), .Z(n6349) );
  AND U9262 ( .A(n6350), .B(n6349), .Z(n6352) );
  NANDN U9263 ( .A(n7010), .B(ereg[165]), .Z(n6351) );
  NAND U9264 ( .A(n6352), .B(n6351), .Z(n2149) );
  NAND U9265 ( .A(n7005), .B(ereg[163]), .Z(n6354) );
  NAND U9266 ( .A(n3909), .B(e[164]), .Z(n6353) );
  AND U9267 ( .A(n6354), .B(n6353), .Z(n6356) );
  NANDN U9268 ( .A(n7010), .B(ereg[164]), .Z(n6355) );
  NAND U9269 ( .A(n6356), .B(n6355), .Z(n2150) );
  NAND U9270 ( .A(n7005), .B(ereg[162]), .Z(n6358) );
  NAND U9271 ( .A(n3909), .B(e[163]), .Z(n6357) );
  AND U9272 ( .A(n6358), .B(n6357), .Z(n6360) );
  NANDN U9273 ( .A(n7010), .B(ereg[163]), .Z(n6359) );
  NAND U9274 ( .A(n6360), .B(n6359), .Z(n2151) );
  NAND U9275 ( .A(n7005), .B(ereg[161]), .Z(n6362) );
  NAND U9276 ( .A(n3909), .B(e[162]), .Z(n6361) );
  AND U9277 ( .A(n6362), .B(n6361), .Z(n6364) );
  NANDN U9278 ( .A(n7010), .B(ereg[162]), .Z(n6363) );
  NAND U9279 ( .A(n6364), .B(n6363), .Z(n2152) );
  NAND U9280 ( .A(n7005), .B(ereg[160]), .Z(n6366) );
  NAND U9281 ( .A(n3909), .B(e[161]), .Z(n6365) );
  AND U9282 ( .A(n6366), .B(n6365), .Z(n6368) );
  NANDN U9283 ( .A(n7010), .B(ereg[161]), .Z(n6367) );
  NAND U9284 ( .A(n6368), .B(n6367), .Z(n2153) );
  NAND U9285 ( .A(n7005), .B(ereg[159]), .Z(n6370) );
  NAND U9286 ( .A(n3909), .B(e[160]), .Z(n6369) );
  AND U9287 ( .A(n6370), .B(n6369), .Z(n6372) );
  NANDN U9288 ( .A(n7010), .B(ereg[160]), .Z(n6371) );
  NAND U9289 ( .A(n6372), .B(n6371), .Z(n2154) );
  NAND U9290 ( .A(n7005), .B(ereg[158]), .Z(n6374) );
  NAND U9291 ( .A(n3909), .B(e[159]), .Z(n6373) );
  AND U9292 ( .A(n6374), .B(n6373), .Z(n6376) );
  NANDN U9293 ( .A(n7010), .B(ereg[159]), .Z(n6375) );
  NAND U9294 ( .A(n6376), .B(n6375), .Z(n2155) );
  NAND U9295 ( .A(n7005), .B(ereg[157]), .Z(n6378) );
  NAND U9296 ( .A(n3909), .B(e[158]), .Z(n6377) );
  AND U9297 ( .A(n6378), .B(n6377), .Z(n6380) );
  NANDN U9298 ( .A(n7010), .B(ereg[158]), .Z(n6379) );
  NAND U9299 ( .A(n6380), .B(n6379), .Z(n2156) );
  NAND U9300 ( .A(n7005), .B(ereg[156]), .Z(n6382) );
  NAND U9301 ( .A(n3910), .B(e[157]), .Z(n6381) );
  AND U9302 ( .A(n6382), .B(n6381), .Z(n6384) );
  NANDN U9303 ( .A(n7010), .B(ereg[157]), .Z(n6383) );
  NAND U9304 ( .A(n6384), .B(n6383), .Z(n2157) );
  NAND U9305 ( .A(n7005), .B(ereg[155]), .Z(n6386) );
  NAND U9306 ( .A(n3910), .B(e[156]), .Z(n6385) );
  AND U9307 ( .A(n6386), .B(n6385), .Z(n6388) );
  NANDN U9308 ( .A(n7010), .B(ereg[156]), .Z(n6387) );
  NAND U9309 ( .A(n6388), .B(n6387), .Z(n2158) );
  NAND U9310 ( .A(n7005), .B(ereg[154]), .Z(n6390) );
  NAND U9311 ( .A(n3910), .B(e[155]), .Z(n6389) );
  AND U9312 ( .A(n6390), .B(n6389), .Z(n6392) );
  NANDN U9313 ( .A(n7010), .B(ereg[155]), .Z(n6391) );
  NAND U9314 ( .A(n6392), .B(n6391), .Z(n2159) );
  NAND U9315 ( .A(n7005), .B(ereg[153]), .Z(n6394) );
  NAND U9316 ( .A(n3910), .B(e[154]), .Z(n6393) );
  AND U9317 ( .A(n6394), .B(n6393), .Z(n6396) );
  NANDN U9318 ( .A(n7010), .B(ereg[154]), .Z(n6395) );
  NAND U9319 ( .A(n6396), .B(n6395), .Z(n2160) );
  NAND U9320 ( .A(n7005), .B(ereg[152]), .Z(n6398) );
  NAND U9321 ( .A(n3910), .B(e[153]), .Z(n6397) );
  AND U9322 ( .A(n6398), .B(n6397), .Z(n6400) );
  NANDN U9323 ( .A(n7010), .B(ereg[153]), .Z(n6399) );
  NAND U9324 ( .A(n6400), .B(n6399), .Z(n2161) );
  NAND U9325 ( .A(n7005), .B(ereg[151]), .Z(n6402) );
  NAND U9326 ( .A(n3910), .B(e[152]), .Z(n6401) );
  AND U9327 ( .A(n6402), .B(n6401), .Z(n6404) );
  NANDN U9328 ( .A(n7010), .B(ereg[152]), .Z(n6403) );
  NAND U9329 ( .A(n6404), .B(n6403), .Z(n2162) );
  NAND U9330 ( .A(n7005), .B(ereg[150]), .Z(n6406) );
  NAND U9331 ( .A(n3910), .B(e[151]), .Z(n6405) );
  AND U9332 ( .A(n6406), .B(n6405), .Z(n6408) );
  NANDN U9333 ( .A(n7010), .B(ereg[151]), .Z(n6407) );
  NAND U9334 ( .A(n6408), .B(n6407), .Z(n2163) );
  NAND U9335 ( .A(n7005), .B(ereg[149]), .Z(n6410) );
  NAND U9336 ( .A(n3911), .B(e[150]), .Z(n6409) );
  AND U9337 ( .A(n6410), .B(n6409), .Z(n6412) );
  NANDN U9338 ( .A(n7010), .B(ereg[150]), .Z(n6411) );
  NAND U9339 ( .A(n6412), .B(n6411), .Z(n2164) );
  NAND U9340 ( .A(n7005), .B(ereg[148]), .Z(n6414) );
  NAND U9341 ( .A(n3911), .B(e[149]), .Z(n6413) );
  AND U9342 ( .A(n6414), .B(n6413), .Z(n6416) );
  NANDN U9343 ( .A(n7010), .B(ereg[149]), .Z(n6415) );
  NAND U9344 ( .A(n6416), .B(n6415), .Z(n2165) );
  NAND U9345 ( .A(n7005), .B(ereg[147]), .Z(n6418) );
  NAND U9346 ( .A(n3911), .B(e[148]), .Z(n6417) );
  AND U9347 ( .A(n6418), .B(n6417), .Z(n6420) );
  NANDN U9348 ( .A(n7010), .B(ereg[148]), .Z(n6419) );
  NAND U9349 ( .A(n6420), .B(n6419), .Z(n2166) );
  NAND U9350 ( .A(n7005), .B(ereg[146]), .Z(n6422) );
  NAND U9351 ( .A(n3911), .B(e[147]), .Z(n6421) );
  AND U9352 ( .A(n6422), .B(n6421), .Z(n6424) );
  NANDN U9353 ( .A(n7010), .B(ereg[147]), .Z(n6423) );
  NAND U9354 ( .A(n6424), .B(n6423), .Z(n2167) );
  NAND U9355 ( .A(n7005), .B(ereg[145]), .Z(n6426) );
  NAND U9356 ( .A(n3911), .B(e[146]), .Z(n6425) );
  AND U9357 ( .A(n6426), .B(n6425), .Z(n6428) );
  NANDN U9358 ( .A(n7010), .B(ereg[146]), .Z(n6427) );
  NAND U9359 ( .A(n6428), .B(n6427), .Z(n2168) );
  NAND U9360 ( .A(n7005), .B(ereg[144]), .Z(n6430) );
  NAND U9361 ( .A(n3911), .B(e[145]), .Z(n6429) );
  AND U9362 ( .A(n6430), .B(n6429), .Z(n6432) );
  NANDN U9363 ( .A(n7010), .B(ereg[145]), .Z(n6431) );
  NAND U9364 ( .A(n6432), .B(n6431), .Z(n2169) );
  NAND U9365 ( .A(n7005), .B(ereg[143]), .Z(n6434) );
  NAND U9366 ( .A(n3911), .B(e[144]), .Z(n6433) );
  AND U9367 ( .A(n6434), .B(n6433), .Z(n6436) );
  NANDN U9368 ( .A(n7010), .B(ereg[144]), .Z(n6435) );
  NAND U9369 ( .A(n6436), .B(n6435), .Z(n2170) );
  NAND U9370 ( .A(n7005), .B(ereg[142]), .Z(n6438) );
  NAND U9371 ( .A(n3912), .B(e[143]), .Z(n6437) );
  AND U9372 ( .A(n6438), .B(n6437), .Z(n6440) );
  NANDN U9373 ( .A(n7010), .B(ereg[143]), .Z(n6439) );
  NAND U9374 ( .A(n6440), .B(n6439), .Z(n2171) );
  NAND U9375 ( .A(n7005), .B(ereg[141]), .Z(n6442) );
  NAND U9376 ( .A(n3912), .B(e[142]), .Z(n6441) );
  AND U9377 ( .A(n6442), .B(n6441), .Z(n6444) );
  NANDN U9378 ( .A(n7010), .B(ereg[142]), .Z(n6443) );
  NAND U9379 ( .A(n6444), .B(n6443), .Z(n2172) );
  NAND U9380 ( .A(n7005), .B(ereg[140]), .Z(n6446) );
  NAND U9381 ( .A(n3912), .B(e[141]), .Z(n6445) );
  AND U9382 ( .A(n6446), .B(n6445), .Z(n6448) );
  NANDN U9383 ( .A(n7010), .B(ereg[141]), .Z(n6447) );
  NAND U9384 ( .A(n6448), .B(n6447), .Z(n2173) );
  NAND U9385 ( .A(n7005), .B(ereg[139]), .Z(n6450) );
  NAND U9386 ( .A(n3912), .B(e[140]), .Z(n6449) );
  AND U9387 ( .A(n6450), .B(n6449), .Z(n6452) );
  NANDN U9388 ( .A(n7010), .B(ereg[140]), .Z(n6451) );
  NAND U9389 ( .A(n6452), .B(n6451), .Z(n2174) );
  NAND U9390 ( .A(n7005), .B(ereg[138]), .Z(n6454) );
  NAND U9391 ( .A(n3912), .B(e[139]), .Z(n6453) );
  AND U9392 ( .A(n6454), .B(n6453), .Z(n6456) );
  NANDN U9393 ( .A(n7010), .B(ereg[139]), .Z(n6455) );
  NAND U9394 ( .A(n6456), .B(n6455), .Z(n2175) );
  NAND U9395 ( .A(n7005), .B(ereg[137]), .Z(n6458) );
  NAND U9396 ( .A(n3912), .B(e[138]), .Z(n6457) );
  AND U9397 ( .A(n6458), .B(n6457), .Z(n6460) );
  NANDN U9398 ( .A(n7010), .B(ereg[138]), .Z(n6459) );
  NAND U9399 ( .A(n6460), .B(n6459), .Z(n2176) );
  NAND U9400 ( .A(n7005), .B(ereg[136]), .Z(n6462) );
  NAND U9401 ( .A(n3912), .B(e[137]), .Z(n6461) );
  AND U9402 ( .A(n6462), .B(n6461), .Z(n6464) );
  NANDN U9403 ( .A(n7010), .B(ereg[137]), .Z(n6463) );
  NAND U9404 ( .A(n6464), .B(n6463), .Z(n2177) );
  NAND U9405 ( .A(n7005), .B(ereg[135]), .Z(n6466) );
  NAND U9406 ( .A(n3913), .B(e[136]), .Z(n6465) );
  AND U9407 ( .A(n6466), .B(n6465), .Z(n6468) );
  NANDN U9408 ( .A(n7010), .B(ereg[136]), .Z(n6467) );
  NAND U9409 ( .A(n6468), .B(n6467), .Z(n2178) );
  NAND U9410 ( .A(n7005), .B(ereg[134]), .Z(n6470) );
  NAND U9411 ( .A(n3913), .B(e[135]), .Z(n6469) );
  AND U9412 ( .A(n6470), .B(n6469), .Z(n6472) );
  NANDN U9413 ( .A(n7010), .B(ereg[135]), .Z(n6471) );
  NAND U9414 ( .A(n6472), .B(n6471), .Z(n2179) );
  NAND U9415 ( .A(n7005), .B(ereg[133]), .Z(n6474) );
  NAND U9416 ( .A(n3913), .B(e[134]), .Z(n6473) );
  AND U9417 ( .A(n6474), .B(n6473), .Z(n6476) );
  NANDN U9418 ( .A(n7010), .B(ereg[134]), .Z(n6475) );
  NAND U9419 ( .A(n6476), .B(n6475), .Z(n2180) );
  NAND U9420 ( .A(n7005), .B(ereg[132]), .Z(n6478) );
  NAND U9421 ( .A(n3913), .B(e[133]), .Z(n6477) );
  AND U9422 ( .A(n6478), .B(n6477), .Z(n6480) );
  NANDN U9423 ( .A(n7010), .B(ereg[133]), .Z(n6479) );
  NAND U9424 ( .A(n6480), .B(n6479), .Z(n2181) );
  NAND U9425 ( .A(n7005), .B(ereg[131]), .Z(n6482) );
  NAND U9426 ( .A(n3913), .B(e[132]), .Z(n6481) );
  AND U9427 ( .A(n6482), .B(n6481), .Z(n6484) );
  NANDN U9428 ( .A(n7010), .B(ereg[132]), .Z(n6483) );
  NAND U9429 ( .A(n6484), .B(n6483), .Z(n2182) );
  NAND U9430 ( .A(n7005), .B(ereg[130]), .Z(n6486) );
  NAND U9431 ( .A(n3913), .B(e[131]), .Z(n6485) );
  AND U9432 ( .A(n6486), .B(n6485), .Z(n6488) );
  NANDN U9433 ( .A(n7010), .B(ereg[131]), .Z(n6487) );
  NAND U9434 ( .A(n6488), .B(n6487), .Z(n2183) );
  NAND U9435 ( .A(n7005), .B(ereg[129]), .Z(n6490) );
  NAND U9436 ( .A(n3913), .B(e[130]), .Z(n6489) );
  AND U9437 ( .A(n6490), .B(n6489), .Z(n6492) );
  NANDN U9438 ( .A(n7010), .B(ereg[130]), .Z(n6491) );
  NAND U9439 ( .A(n6492), .B(n6491), .Z(n2184) );
  NAND U9440 ( .A(n7005), .B(ereg[128]), .Z(n6494) );
  NAND U9441 ( .A(n3914), .B(e[129]), .Z(n6493) );
  AND U9442 ( .A(n6494), .B(n6493), .Z(n6496) );
  NANDN U9443 ( .A(n7010), .B(ereg[129]), .Z(n6495) );
  NAND U9444 ( .A(n6496), .B(n6495), .Z(n2185) );
  NAND U9445 ( .A(n7005), .B(ereg[127]), .Z(n6498) );
  NAND U9446 ( .A(n3914), .B(e[128]), .Z(n6497) );
  AND U9447 ( .A(n6498), .B(n6497), .Z(n6500) );
  NANDN U9448 ( .A(n7010), .B(ereg[128]), .Z(n6499) );
  NAND U9449 ( .A(n6500), .B(n6499), .Z(n2186) );
  NAND U9450 ( .A(n7005), .B(ereg[126]), .Z(n6502) );
  NAND U9451 ( .A(n3914), .B(e[127]), .Z(n6501) );
  AND U9452 ( .A(n6502), .B(n6501), .Z(n6504) );
  NANDN U9453 ( .A(n7010), .B(ereg[127]), .Z(n6503) );
  NAND U9454 ( .A(n6504), .B(n6503), .Z(n2187) );
  NAND U9455 ( .A(n7005), .B(ereg[125]), .Z(n6506) );
  NAND U9456 ( .A(n3914), .B(e[126]), .Z(n6505) );
  AND U9457 ( .A(n6506), .B(n6505), .Z(n6508) );
  NANDN U9458 ( .A(n7010), .B(ereg[126]), .Z(n6507) );
  NAND U9459 ( .A(n6508), .B(n6507), .Z(n2188) );
  NAND U9460 ( .A(n7005), .B(ereg[124]), .Z(n6510) );
  NAND U9461 ( .A(n3914), .B(e[125]), .Z(n6509) );
  AND U9462 ( .A(n6510), .B(n6509), .Z(n6512) );
  NANDN U9463 ( .A(n7010), .B(ereg[125]), .Z(n6511) );
  NAND U9464 ( .A(n6512), .B(n6511), .Z(n2189) );
  NAND U9465 ( .A(n7005), .B(ereg[123]), .Z(n6514) );
  NAND U9466 ( .A(n3914), .B(e[124]), .Z(n6513) );
  AND U9467 ( .A(n6514), .B(n6513), .Z(n6516) );
  NANDN U9468 ( .A(n7010), .B(ereg[124]), .Z(n6515) );
  NAND U9469 ( .A(n6516), .B(n6515), .Z(n2190) );
  NAND U9470 ( .A(n7005), .B(ereg[122]), .Z(n6518) );
  NAND U9471 ( .A(n3914), .B(e[123]), .Z(n6517) );
  AND U9472 ( .A(n6518), .B(n6517), .Z(n6520) );
  NANDN U9473 ( .A(n7010), .B(ereg[123]), .Z(n6519) );
  NAND U9474 ( .A(n6520), .B(n6519), .Z(n2191) );
  NAND U9475 ( .A(n7005), .B(ereg[121]), .Z(n6522) );
  NAND U9476 ( .A(n3915), .B(e[122]), .Z(n6521) );
  AND U9477 ( .A(n6522), .B(n6521), .Z(n6524) );
  NANDN U9478 ( .A(n7010), .B(ereg[122]), .Z(n6523) );
  NAND U9479 ( .A(n6524), .B(n6523), .Z(n2192) );
  NAND U9480 ( .A(n7005), .B(ereg[120]), .Z(n6526) );
  NAND U9481 ( .A(n3915), .B(e[121]), .Z(n6525) );
  AND U9482 ( .A(n6526), .B(n6525), .Z(n6528) );
  NANDN U9483 ( .A(n7010), .B(ereg[121]), .Z(n6527) );
  NAND U9484 ( .A(n6528), .B(n6527), .Z(n2193) );
  NAND U9485 ( .A(n7005), .B(ereg[119]), .Z(n6530) );
  NAND U9486 ( .A(n3915), .B(e[120]), .Z(n6529) );
  AND U9487 ( .A(n6530), .B(n6529), .Z(n6532) );
  NANDN U9488 ( .A(n7010), .B(ereg[120]), .Z(n6531) );
  NAND U9489 ( .A(n6532), .B(n6531), .Z(n2194) );
  NAND U9490 ( .A(n7005), .B(ereg[118]), .Z(n6534) );
  NAND U9491 ( .A(n3915), .B(e[119]), .Z(n6533) );
  AND U9492 ( .A(n6534), .B(n6533), .Z(n6536) );
  NANDN U9493 ( .A(n7010), .B(ereg[119]), .Z(n6535) );
  NAND U9494 ( .A(n6536), .B(n6535), .Z(n2195) );
  NAND U9495 ( .A(n7005), .B(ereg[117]), .Z(n6538) );
  NAND U9496 ( .A(n3915), .B(e[118]), .Z(n6537) );
  AND U9497 ( .A(n6538), .B(n6537), .Z(n6540) );
  NANDN U9498 ( .A(n7010), .B(ereg[118]), .Z(n6539) );
  NAND U9499 ( .A(n6540), .B(n6539), .Z(n2196) );
  NAND U9500 ( .A(n7005), .B(ereg[116]), .Z(n6542) );
  NAND U9501 ( .A(n3915), .B(e[117]), .Z(n6541) );
  AND U9502 ( .A(n6542), .B(n6541), .Z(n6544) );
  NANDN U9503 ( .A(n7010), .B(ereg[117]), .Z(n6543) );
  NAND U9504 ( .A(n6544), .B(n6543), .Z(n2197) );
  NAND U9505 ( .A(n7005), .B(ereg[115]), .Z(n6546) );
  NAND U9506 ( .A(n3915), .B(e[116]), .Z(n6545) );
  AND U9507 ( .A(n6546), .B(n6545), .Z(n6548) );
  NANDN U9508 ( .A(n7010), .B(ereg[116]), .Z(n6547) );
  NAND U9509 ( .A(n6548), .B(n6547), .Z(n2198) );
  NAND U9510 ( .A(n7005), .B(ereg[114]), .Z(n6550) );
  NAND U9511 ( .A(n3916), .B(e[115]), .Z(n6549) );
  AND U9512 ( .A(n6550), .B(n6549), .Z(n6552) );
  NANDN U9513 ( .A(n7010), .B(ereg[115]), .Z(n6551) );
  NAND U9514 ( .A(n6552), .B(n6551), .Z(n2199) );
  NAND U9515 ( .A(n7005), .B(ereg[113]), .Z(n6554) );
  NAND U9516 ( .A(n3916), .B(e[114]), .Z(n6553) );
  AND U9517 ( .A(n6554), .B(n6553), .Z(n6556) );
  NANDN U9518 ( .A(n7010), .B(ereg[114]), .Z(n6555) );
  NAND U9519 ( .A(n6556), .B(n6555), .Z(n2200) );
  NAND U9520 ( .A(n7005), .B(ereg[112]), .Z(n6558) );
  NAND U9521 ( .A(n3916), .B(e[113]), .Z(n6557) );
  AND U9522 ( .A(n6558), .B(n6557), .Z(n6560) );
  NANDN U9523 ( .A(n7010), .B(ereg[113]), .Z(n6559) );
  NAND U9524 ( .A(n6560), .B(n6559), .Z(n2201) );
  NAND U9525 ( .A(n7005), .B(ereg[111]), .Z(n6562) );
  NAND U9526 ( .A(n3916), .B(e[112]), .Z(n6561) );
  AND U9527 ( .A(n6562), .B(n6561), .Z(n6564) );
  NANDN U9528 ( .A(n7010), .B(ereg[112]), .Z(n6563) );
  NAND U9529 ( .A(n6564), .B(n6563), .Z(n2202) );
  NAND U9530 ( .A(n7005), .B(ereg[110]), .Z(n6566) );
  NAND U9531 ( .A(n3916), .B(e[111]), .Z(n6565) );
  AND U9532 ( .A(n6566), .B(n6565), .Z(n6568) );
  NANDN U9533 ( .A(n7010), .B(ereg[111]), .Z(n6567) );
  NAND U9534 ( .A(n6568), .B(n6567), .Z(n2203) );
  NAND U9535 ( .A(n7005), .B(ereg[109]), .Z(n6570) );
  NAND U9536 ( .A(n3916), .B(e[110]), .Z(n6569) );
  AND U9537 ( .A(n6570), .B(n6569), .Z(n6572) );
  NANDN U9538 ( .A(n7010), .B(ereg[110]), .Z(n6571) );
  NAND U9539 ( .A(n6572), .B(n6571), .Z(n2204) );
  NAND U9540 ( .A(n7005), .B(ereg[108]), .Z(n6574) );
  NAND U9541 ( .A(n3916), .B(e[109]), .Z(n6573) );
  AND U9542 ( .A(n6574), .B(n6573), .Z(n6576) );
  NANDN U9543 ( .A(n7010), .B(ereg[109]), .Z(n6575) );
  NAND U9544 ( .A(n6576), .B(n6575), .Z(n2205) );
  NAND U9545 ( .A(n7005), .B(ereg[107]), .Z(n6578) );
  NAND U9546 ( .A(n3917), .B(e[108]), .Z(n6577) );
  AND U9547 ( .A(n6578), .B(n6577), .Z(n6580) );
  NANDN U9548 ( .A(n7010), .B(ereg[108]), .Z(n6579) );
  NAND U9549 ( .A(n6580), .B(n6579), .Z(n2206) );
  NAND U9550 ( .A(n7005), .B(ereg[106]), .Z(n6582) );
  NAND U9551 ( .A(n3917), .B(e[107]), .Z(n6581) );
  AND U9552 ( .A(n6582), .B(n6581), .Z(n6584) );
  NANDN U9553 ( .A(n7010), .B(ereg[107]), .Z(n6583) );
  NAND U9554 ( .A(n6584), .B(n6583), .Z(n2207) );
  NAND U9555 ( .A(n7005), .B(ereg[105]), .Z(n6586) );
  NAND U9556 ( .A(n3917), .B(e[106]), .Z(n6585) );
  AND U9557 ( .A(n6586), .B(n6585), .Z(n6588) );
  NANDN U9558 ( .A(n7010), .B(ereg[106]), .Z(n6587) );
  NAND U9559 ( .A(n6588), .B(n6587), .Z(n2208) );
  NAND U9560 ( .A(n7005), .B(ereg[104]), .Z(n6590) );
  NAND U9561 ( .A(n3917), .B(e[105]), .Z(n6589) );
  AND U9562 ( .A(n6590), .B(n6589), .Z(n6592) );
  NANDN U9563 ( .A(n7010), .B(ereg[105]), .Z(n6591) );
  NAND U9564 ( .A(n6592), .B(n6591), .Z(n2209) );
  NAND U9565 ( .A(n7005), .B(ereg[103]), .Z(n6594) );
  NAND U9566 ( .A(n3917), .B(e[104]), .Z(n6593) );
  AND U9567 ( .A(n6594), .B(n6593), .Z(n6596) );
  NANDN U9568 ( .A(n7010), .B(ereg[104]), .Z(n6595) );
  NAND U9569 ( .A(n6596), .B(n6595), .Z(n2210) );
  NAND U9570 ( .A(n7005), .B(ereg[102]), .Z(n6598) );
  NAND U9571 ( .A(n3917), .B(e[103]), .Z(n6597) );
  AND U9572 ( .A(n6598), .B(n6597), .Z(n6600) );
  NANDN U9573 ( .A(n7010), .B(ereg[103]), .Z(n6599) );
  NAND U9574 ( .A(n6600), .B(n6599), .Z(n2211) );
  NAND U9575 ( .A(n7005), .B(ereg[101]), .Z(n6602) );
  NAND U9576 ( .A(n3917), .B(e[102]), .Z(n6601) );
  AND U9577 ( .A(n6602), .B(n6601), .Z(n6604) );
  NANDN U9578 ( .A(n7010), .B(ereg[102]), .Z(n6603) );
  NAND U9579 ( .A(n6604), .B(n6603), .Z(n2212) );
  NAND U9580 ( .A(n7005), .B(ereg[100]), .Z(n6606) );
  NAND U9581 ( .A(n3918), .B(e[101]), .Z(n6605) );
  AND U9582 ( .A(n6606), .B(n6605), .Z(n6608) );
  NANDN U9583 ( .A(n7010), .B(ereg[101]), .Z(n6607) );
  NAND U9584 ( .A(n6608), .B(n6607), .Z(n2213) );
  NAND U9585 ( .A(n7005), .B(ereg[99]), .Z(n6610) );
  NAND U9586 ( .A(n3918), .B(e[100]), .Z(n6609) );
  AND U9587 ( .A(n6610), .B(n6609), .Z(n6612) );
  NANDN U9588 ( .A(n7010), .B(ereg[100]), .Z(n6611) );
  NAND U9589 ( .A(n6612), .B(n6611), .Z(n2214) );
  NAND U9590 ( .A(n7005), .B(ereg[98]), .Z(n6614) );
  NAND U9591 ( .A(n3918), .B(e[99]), .Z(n6613) );
  AND U9592 ( .A(n6614), .B(n6613), .Z(n6616) );
  NANDN U9593 ( .A(n7010), .B(ereg[99]), .Z(n6615) );
  NAND U9594 ( .A(n6616), .B(n6615), .Z(n2215) );
  NAND U9595 ( .A(n7005), .B(ereg[97]), .Z(n6618) );
  NAND U9596 ( .A(n3918), .B(e[98]), .Z(n6617) );
  AND U9597 ( .A(n6618), .B(n6617), .Z(n6620) );
  NANDN U9598 ( .A(n7010), .B(ereg[98]), .Z(n6619) );
  NAND U9599 ( .A(n6620), .B(n6619), .Z(n2216) );
  NAND U9600 ( .A(n7005), .B(ereg[96]), .Z(n6622) );
  NAND U9601 ( .A(n3918), .B(e[97]), .Z(n6621) );
  AND U9602 ( .A(n6622), .B(n6621), .Z(n6624) );
  NANDN U9603 ( .A(n7010), .B(ereg[97]), .Z(n6623) );
  NAND U9604 ( .A(n6624), .B(n6623), .Z(n2217) );
  NAND U9605 ( .A(n7005), .B(ereg[95]), .Z(n6626) );
  NAND U9606 ( .A(n3918), .B(e[96]), .Z(n6625) );
  AND U9607 ( .A(n6626), .B(n6625), .Z(n6628) );
  NANDN U9608 ( .A(n7010), .B(ereg[96]), .Z(n6627) );
  NAND U9609 ( .A(n6628), .B(n6627), .Z(n2218) );
  NAND U9610 ( .A(n7005), .B(ereg[94]), .Z(n6630) );
  NAND U9611 ( .A(n3918), .B(e[95]), .Z(n6629) );
  AND U9612 ( .A(n6630), .B(n6629), .Z(n6632) );
  NANDN U9613 ( .A(n7010), .B(ereg[95]), .Z(n6631) );
  NAND U9614 ( .A(n6632), .B(n6631), .Z(n2219) );
  NAND U9615 ( .A(n7005), .B(ereg[93]), .Z(n6634) );
  NAND U9616 ( .A(n3919), .B(e[94]), .Z(n6633) );
  AND U9617 ( .A(n6634), .B(n6633), .Z(n6636) );
  NANDN U9618 ( .A(n7010), .B(ereg[94]), .Z(n6635) );
  NAND U9619 ( .A(n6636), .B(n6635), .Z(n2220) );
  NAND U9620 ( .A(n7005), .B(ereg[92]), .Z(n6638) );
  NAND U9621 ( .A(n3919), .B(e[93]), .Z(n6637) );
  AND U9622 ( .A(n6638), .B(n6637), .Z(n6640) );
  NANDN U9623 ( .A(n7010), .B(ereg[93]), .Z(n6639) );
  NAND U9624 ( .A(n6640), .B(n6639), .Z(n2221) );
  NAND U9625 ( .A(n7005), .B(ereg[91]), .Z(n6642) );
  NAND U9626 ( .A(n3919), .B(e[92]), .Z(n6641) );
  AND U9627 ( .A(n6642), .B(n6641), .Z(n6644) );
  NANDN U9628 ( .A(n7010), .B(ereg[92]), .Z(n6643) );
  NAND U9629 ( .A(n6644), .B(n6643), .Z(n2222) );
  NAND U9630 ( .A(n7005), .B(ereg[90]), .Z(n6646) );
  NAND U9631 ( .A(n3919), .B(e[91]), .Z(n6645) );
  AND U9632 ( .A(n6646), .B(n6645), .Z(n6648) );
  NANDN U9633 ( .A(n7010), .B(ereg[91]), .Z(n6647) );
  NAND U9634 ( .A(n6648), .B(n6647), .Z(n2223) );
  NAND U9635 ( .A(n7005), .B(ereg[89]), .Z(n6650) );
  NAND U9636 ( .A(n3919), .B(e[90]), .Z(n6649) );
  AND U9637 ( .A(n6650), .B(n6649), .Z(n6652) );
  NANDN U9638 ( .A(n7010), .B(ereg[90]), .Z(n6651) );
  NAND U9639 ( .A(n6652), .B(n6651), .Z(n2224) );
  NAND U9640 ( .A(n7005), .B(ereg[88]), .Z(n6654) );
  NAND U9641 ( .A(n3919), .B(e[89]), .Z(n6653) );
  AND U9642 ( .A(n6654), .B(n6653), .Z(n6656) );
  NANDN U9643 ( .A(n7010), .B(ereg[89]), .Z(n6655) );
  NAND U9644 ( .A(n6656), .B(n6655), .Z(n2225) );
  NAND U9645 ( .A(n7005), .B(ereg[87]), .Z(n6658) );
  NAND U9646 ( .A(n3919), .B(e[88]), .Z(n6657) );
  AND U9647 ( .A(n6658), .B(n6657), .Z(n6660) );
  NANDN U9648 ( .A(n7010), .B(ereg[88]), .Z(n6659) );
  NAND U9649 ( .A(n6660), .B(n6659), .Z(n2226) );
  NAND U9650 ( .A(n7005), .B(ereg[86]), .Z(n6662) );
  NAND U9651 ( .A(n3920), .B(e[87]), .Z(n6661) );
  AND U9652 ( .A(n6662), .B(n6661), .Z(n6664) );
  NANDN U9653 ( .A(n7010), .B(ereg[87]), .Z(n6663) );
  NAND U9654 ( .A(n6664), .B(n6663), .Z(n2227) );
  NAND U9655 ( .A(n7005), .B(ereg[85]), .Z(n6666) );
  NAND U9656 ( .A(n3920), .B(e[86]), .Z(n6665) );
  AND U9657 ( .A(n6666), .B(n6665), .Z(n6668) );
  NANDN U9658 ( .A(n7010), .B(ereg[86]), .Z(n6667) );
  NAND U9659 ( .A(n6668), .B(n6667), .Z(n2228) );
  NAND U9660 ( .A(n7005), .B(ereg[84]), .Z(n6670) );
  NAND U9661 ( .A(n3920), .B(e[85]), .Z(n6669) );
  AND U9662 ( .A(n6670), .B(n6669), .Z(n6672) );
  NANDN U9663 ( .A(n7010), .B(ereg[85]), .Z(n6671) );
  NAND U9664 ( .A(n6672), .B(n6671), .Z(n2229) );
  NAND U9665 ( .A(n7005), .B(ereg[83]), .Z(n6674) );
  NAND U9666 ( .A(n3920), .B(e[84]), .Z(n6673) );
  AND U9667 ( .A(n6674), .B(n6673), .Z(n6676) );
  NANDN U9668 ( .A(n7010), .B(ereg[84]), .Z(n6675) );
  NAND U9669 ( .A(n6676), .B(n6675), .Z(n2230) );
  NAND U9670 ( .A(n7005), .B(ereg[82]), .Z(n6678) );
  NAND U9671 ( .A(n3920), .B(e[83]), .Z(n6677) );
  AND U9672 ( .A(n6678), .B(n6677), .Z(n6680) );
  NANDN U9673 ( .A(n7010), .B(ereg[83]), .Z(n6679) );
  NAND U9674 ( .A(n6680), .B(n6679), .Z(n2231) );
  NAND U9675 ( .A(n7005), .B(ereg[81]), .Z(n6682) );
  NAND U9676 ( .A(n3920), .B(e[82]), .Z(n6681) );
  AND U9677 ( .A(n6682), .B(n6681), .Z(n6684) );
  NANDN U9678 ( .A(n7010), .B(ereg[82]), .Z(n6683) );
  NAND U9679 ( .A(n6684), .B(n6683), .Z(n2232) );
  NAND U9680 ( .A(n7005), .B(ereg[80]), .Z(n6686) );
  NAND U9681 ( .A(n3920), .B(e[81]), .Z(n6685) );
  AND U9682 ( .A(n6686), .B(n6685), .Z(n6688) );
  NANDN U9683 ( .A(n7010), .B(ereg[81]), .Z(n6687) );
  NAND U9684 ( .A(n6688), .B(n6687), .Z(n2233) );
  NAND U9685 ( .A(n7005), .B(ereg[79]), .Z(n6690) );
  NAND U9686 ( .A(n3921), .B(e[80]), .Z(n6689) );
  AND U9687 ( .A(n6690), .B(n6689), .Z(n6692) );
  NANDN U9688 ( .A(n7010), .B(ereg[80]), .Z(n6691) );
  NAND U9689 ( .A(n6692), .B(n6691), .Z(n2234) );
  NAND U9690 ( .A(n7005), .B(ereg[78]), .Z(n6694) );
  NAND U9691 ( .A(n3921), .B(e[79]), .Z(n6693) );
  AND U9692 ( .A(n6694), .B(n6693), .Z(n6696) );
  NANDN U9693 ( .A(n7010), .B(ereg[79]), .Z(n6695) );
  NAND U9694 ( .A(n6696), .B(n6695), .Z(n2235) );
  NAND U9695 ( .A(n7005), .B(ereg[77]), .Z(n6698) );
  NAND U9696 ( .A(n3921), .B(e[78]), .Z(n6697) );
  AND U9697 ( .A(n6698), .B(n6697), .Z(n6700) );
  NANDN U9698 ( .A(n7010), .B(ereg[78]), .Z(n6699) );
  NAND U9699 ( .A(n6700), .B(n6699), .Z(n2236) );
  NAND U9700 ( .A(n7005), .B(ereg[76]), .Z(n6702) );
  NAND U9701 ( .A(n3921), .B(e[77]), .Z(n6701) );
  AND U9702 ( .A(n6702), .B(n6701), .Z(n6704) );
  NANDN U9703 ( .A(n7010), .B(ereg[77]), .Z(n6703) );
  NAND U9704 ( .A(n6704), .B(n6703), .Z(n2237) );
  NAND U9705 ( .A(n7005), .B(ereg[75]), .Z(n6706) );
  NAND U9706 ( .A(n3921), .B(e[76]), .Z(n6705) );
  AND U9707 ( .A(n6706), .B(n6705), .Z(n6708) );
  NANDN U9708 ( .A(n7010), .B(ereg[76]), .Z(n6707) );
  NAND U9709 ( .A(n6708), .B(n6707), .Z(n2238) );
  NAND U9710 ( .A(n7005), .B(ereg[74]), .Z(n6710) );
  NAND U9711 ( .A(n3921), .B(e[75]), .Z(n6709) );
  AND U9712 ( .A(n6710), .B(n6709), .Z(n6712) );
  NANDN U9713 ( .A(n7010), .B(ereg[75]), .Z(n6711) );
  NAND U9714 ( .A(n6712), .B(n6711), .Z(n2239) );
  NAND U9715 ( .A(n7005), .B(ereg[73]), .Z(n6714) );
  NAND U9716 ( .A(n3921), .B(e[74]), .Z(n6713) );
  AND U9717 ( .A(n6714), .B(n6713), .Z(n6716) );
  NANDN U9718 ( .A(n7010), .B(ereg[74]), .Z(n6715) );
  NAND U9719 ( .A(n6716), .B(n6715), .Z(n2240) );
  NAND U9720 ( .A(n7005), .B(ereg[72]), .Z(n6718) );
  NAND U9721 ( .A(n3922), .B(e[73]), .Z(n6717) );
  AND U9722 ( .A(n6718), .B(n6717), .Z(n6720) );
  NANDN U9723 ( .A(n7010), .B(ereg[73]), .Z(n6719) );
  NAND U9724 ( .A(n6720), .B(n6719), .Z(n2241) );
  NAND U9725 ( .A(n7005), .B(ereg[71]), .Z(n6722) );
  NAND U9726 ( .A(n3922), .B(e[72]), .Z(n6721) );
  AND U9727 ( .A(n6722), .B(n6721), .Z(n6724) );
  NANDN U9728 ( .A(n7010), .B(ereg[72]), .Z(n6723) );
  NAND U9729 ( .A(n6724), .B(n6723), .Z(n2242) );
  NAND U9730 ( .A(n7005), .B(ereg[70]), .Z(n6726) );
  NAND U9731 ( .A(n3922), .B(e[71]), .Z(n6725) );
  AND U9732 ( .A(n6726), .B(n6725), .Z(n6728) );
  NANDN U9733 ( .A(n7010), .B(ereg[71]), .Z(n6727) );
  NAND U9734 ( .A(n6728), .B(n6727), .Z(n2243) );
  NAND U9735 ( .A(n7005), .B(ereg[69]), .Z(n6730) );
  NAND U9736 ( .A(n3922), .B(e[70]), .Z(n6729) );
  AND U9737 ( .A(n6730), .B(n6729), .Z(n6732) );
  NANDN U9738 ( .A(n7010), .B(ereg[70]), .Z(n6731) );
  NAND U9739 ( .A(n6732), .B(n6731), .Z(n2244) );
  NAND U9740 ( .A(n7005), .B(ereg[68]), .Z(n6734) );
  NAND U9741 ( .A(n3922), .B(e[69]), .Z(n6733) );
  AND U9742 ( .A(n6734), .B(n6733), .Z(n6736) );
  NANDN U9743 ( .A(n7010), .B(ereg[69]), .Z(n6735) );
  NAND U9744 ( .A(n6736), .B(n6735), .Z(n2245) );
  NAND U9745 ( .A(n7005), .B(ereg[67]), .Z(n6738) );
  NAND U9746 ( .A(n3922), .B(e[68]), .Z(n6737) );
  AND U9747 ( .A(n6738), .B(n6737), .Z(n6740) );
  NANDN U9748 ( .A(n7010), .B(ereg[68]), .Z(n6739) );
  NAND U9749 ( .A(n6740), .B(n6739), .Z(n2246) );
  NAND U9750 ( .A(n7005), .B(ereg[66]), .Z(n6742) );
  NAND U9751 ( .A(n3922), .B(e[67]), .Z(n6741) );
  AND U9752 ( .A(n6742), .B(n6741), .Z(n6744) );
  NANDN U9753 ( .A(n7010), .B(ereg[67]), .Z(n6743) );
  NAND U9754 ( .A(n6744), .B(n6743), .Z(n2247) );
  NAND U9755 ( .A(n7005), .B(ereg[65]), .Z(n6746) );
  NAND U9756 ( .A(n3923), .B(e[66]), .Z(n6745) );
  AND U9757 ( .A(n6746), .B(n6745), .Z(n6748) );
  NANDN U9758 ( .A(n7010), .B(ereg[66]), .Z(n6747) );
  NAND U9759 ( .A(n6748), .B(n6747), .Z(n2248) );
  NAND U9760 ( .A(n7005), .B(ereg[64]), .Z(n6750) );
  NAND U9761 ( .A(n3923), .B(e[65]), .Z(n6749) );
  AND U9762 ( .A(n6750), .B(n6749), .Z(n6752) );
  NANDN U9763 ( .A(n7010), .B(ereg[65]), .Z(n6751) );
  NAND U9764 ( .A(n6752), .B(n6751), .Z(n2249) );
  NAND U9765 ( .A(n7005), .B(ereg[63]), .Z(n6754) );
  NAND U9766 ( .A(n3923), .B(e[64]), .Z(n6753) );
  AND U9767 ( .A(n6754), .B(n6753), .Z(n6756) );
  NANDN U9768 ( .A(n7010), .B(ereg[64]), .Z(n6755) );
  NAND U9769 ( .A(n6756), .B(n6755), .Z(n2250) );
  NAND U9770 ( .A(n7005), .B(ereg[62]), .Z(n6758) );
  NAND U9771 ( .A(n3923), .B(e[63]), .Z(n6757) );
  AND U9772 ( .A(n6758), .B(n6757), .Z(n6760) );
  NANDN U9773 ( .A(n7010), .B(ereg[63]), .Z(n6759) );
  NAND U9774 ( .A(n6760), .B(n6759), .Z(n2251) );
  NAND U9775 ( .A(n7005), .B(ereg[61]), .Z(n6762) );
  NAND U9776 ( .A(n3923), .B(e[62]), .Z(n6761) );
  AND U9777 ( .A(n6762), .B(n6761), .Z(n6764) );
  NANDN U9778 ( .A(n7010), .B(ereg[62]), .Z(n6763) );
  NAND U9779 ( .A(n6764), .B(n6763), .Z(n2252) );
  NAND U9780 ( .A(n7005), .B(ereg[60]), .Z(n6766) );
  NAND U9781 ( .A(n3923), .B(e[61]), .Z(n6765) );
  AND U9782 ( .A(n6766), .B(n6765), .Z(n6768) );
  NANDN U9783 ( .A(n7010), .B(ereg[61]), .Z(n6767) );
  NAND U9784 ( .A(n6768), .B(n6767), .Z(n2253) );
  NAND U9785 ( .A(n7005), .B(ereg[59]), .Z(n6770) );
  NAND U9786 ( .A(n3923), .B(e[60]), .Z(n6769) );
  AND U9787 ( .A(n6770), .B(n6769), .Z(n6772) );
  NANDN U9788 ( .A(n7010), .B(ereg[60]), .Z(n6771) );
  NAND U9789 ( .A(n6772), .B(n6771), .Z(n2254) );
  NAND U9790 ( .A(n7005), .B(ereg[58]), .Z(n6774) );
  NAND U9791 ( .A(n3924), .B(e[59]), .Z(n6773) );
  AND U9792 ( .A(n6774), .B(n6773), .Z(n6776) );
  NANDN U9793 ( .A(n7010), .B(ereg[59]), .Z(n6775) );
  NAND U9794 ( .A(n6776), .B(n6775), .Z(n2255) );
  NAND U9795 ( .A(n7005), .B(ereg[57]), .Z(n6778) );
  NAND U9796 ( .A(n3924), .B(e[58]), .Z(n6777) );
  AND U9797 ( .A(n6778), .B(n6777), .Z(n6780) );
  NANDN U9798 ( .A(n7010), .B(ereg[58]), .Z(n6779) );
  NAND U9799 ( .A(n6780), .B(n6779), .Z(n2256) );
  NAND U9800 ( .A(n7005), .B(ereg[56]), .Z(n6782) );
  NAND U9801 ( .A(n3924), .B(e[57]), .Z(n6781) );
  AND U9802 ( .A(n6782), .B(n6781), .Z(n6784) );
  NANDN U9803 ( .A(n7010), .B(ereg[57]), .Z(n6783) );
  NAND U9804 ( .A(n6784), .B(n6783), .Z(n2257) );
  NAND U9805 ( .A(n7005), .B(ereg[55]), .Z(n6786) );
  NAND U9806 ( .A(n3924), .B(e[56]), .Z(n6785) );
  AND U9807 ( .A(n6786), .B(n6785), .Z(n6788) );
  NANDN U9808 ( .A(n7010), .B(ereg[56]), .Z(n6787) );
  NAND U9809 ( .A(n6788), .B(n6787), .Z(n2258) );
  NAND U9810 ( .A(n7005), .B(ereg[54]), .Z(n6790) );
  NAND U9811 ( .A(n3924), .B(e[55]), .Z(n6789) );
  AND U9812 ( .A(n6790), .B(n6789), .Z(n6792) );
  NANDN U9813 ( .A(n7010), .B(ereg[55]), .Z(n6791) );
  NAND U9814 ( .A(n6792), .B(n6791), .Z(n2259) );
  NAND U9815 ( .A(n7005), .B(ereg[53]), .Z(n6794) );
  NAND U9816 ( .A(n3924), .B(e[54]), .Z(n6793) );
  AND U9817 ( .A(n6794), .B(n6793), .Z(n6796) );
  NANDN U9818 ( .A(n7010), .B(ereg[54]), .Z(n6795) );
  NAND U9819 ( .A(n6796), .B(n6795), .Z(n2260) );
  NAND U9820 ( .A(n7005), .B(ereg[52]), .Z(n6798) );
  NAND U9821 ( .A(n3924), .B(e[53]), .Z(n6797) );
  AND U9822 ( .A(n6798), .B(n6797), .Z(n6800) );
  NANDN U9823 ( .A(n7010), .B(ereg[53]), .Z(n6799) );
  NAND U9824 ( .A(n6800), .B(n6799), .Z(n2261) );
  NAND U9825 ( .A(n7005), .B(ereg[51]), .Z(n6802) );
  NAND U9826 ( .A(n3925), .B(e[52]), .Z(n6801) );
  AND U9827 ( .A(n6802), .B(n6801), .Z(n6804) );
  NANDN U9828 ( .A(n7010), .B(ereg[52]), .Z(n6803) );
  NAND U9829 ( .A(n6804), .B(n6803), .Z(n2262) );
  NAND U9830 ( .A(n7005), .B(ereg[50]), .Z(n6806) );
  NAND U9831 ( .A(n3925), .B(e[51]), .Z(n6805) );
  AND U9832 ( .A(n6806), .B(n6805), .Z(n6808) );
  NANDN U9833 ( .A(n7010), .B(ereg[51]), .Z(n6807) );
  NAND U9834 ( .A(n6808), .B(n6807), .Z(n2263) );
  NAND U9835 ( .A(n7005), .B(ereg[49]), .Z(n6810) );
  NAND U9836 ( .A(n3925), .B(e[50]), .Z(n6809) );
  AND U9837 ( .A(n6810), .B(n6809), .Z(n6812) );
  NANDN U9838 ( .A(n7010), .B(ereg[50]), .Z(n6811) );
  NAND U9839 ( .A(n6812), .B(n6811), .Z(n2264) );
  NAND U9840 ( .A(n7005), .B(ereg[48]), .Z(n6814) );
  NAND U9841 ( .A(n3925), .B(e[49]), .Z(n6813) );
  AND U9842 ( .A(n6814), .B(n6813), .Z(n6816) );
  NANDN U9843 ( .A(n7010), .B(ereg[49]), .Z(n6815) );
  NAND U9844 ( .A(n6816), .B(n6815), .Z(n2265) );
  NAND U9845 ( .A(n7005), .B(ereg[47]), .Z(n6818) );
  NAND U9846 ( .A(n3925), .B(e[48]), .Z(n6817) );
  AND U9847 ( .A(n6818), .B(n6817), .Z(n6820) );
  NANDN U9848 ( .A(n7010), .B(ereg[48]), .Z(n6819) );
  NAND U9849 ( .A(n6820), .B(n6819), .Z(n2266) );
  NAND U9850 ( .A(n7005), .B(ereg[46]), .Z(n6822) );
  NAND U9851 ( .A(n3925), .B(e[47]), .Z(n6821) );
  AND U9852 ( .A(n6822), .B(n6821), .Z(n6824) );
  NANDN U9853 ( .A(n7010), .B(ereg[47]), .Z(n6823) );
  NAND U9854 ( .A(n6824), .B(n6823), .Z(n2267) );
  NAND U9855 ( .A(n7005), .B(ereg[45]), .Z(n6826) );
  NAND U9856 ( .A(n3925), .B(e[46]), .Z(n6825) );
  AND U9857 ( .A(n6826), .B(n6825), .Z(n6828) );
  NANDN U9858 ( .A(n7010), .B(ereg[46]), .Z(n6827) );
  NAND U9859 ( .A(n6828), .B(n6827), .Z(n2268) );
  NAND U9860 ( .A(n7005), .B(ereg[44]), .Z(n6830) );
  NAND U9861 ( .A(n3926), .B(e[45]), .Z(n6829) );
  AND U9862 ( .A(n6830), .B(n6829), .Z(n6832) );
  NANDN U9863 ( .A(n7010), .B(ereg[45]), .Z(n6831) );
  NAND U9864 ( .A(n6832), .B(n6831), .Z(n2269) );
  NAND U9865 ( .A(n7005), .B(ereg[43]), .Z(n6834) );
  NAND U9866 ( .A(n3926), .B(e[44]), .Z(n6833) );
  AND U9867 ( .A(n6834), .B(n6833), .Z(n6836) );
  NANDN U9868 ( .A(n7010), .B(ereg[44]), .Z(n6835) );
  NAND U9869 ( .A(n6836), .B(n6835), .Z(n2270) );
  NAND U9870 ( .A(n7005), .B(ereg[42]), .Z(n6838) );
  NAND U9871 ( .A(n3926), .B(e[43]), .Z(n6837) );
  AND U9872 ( .A(n6838), .B(n6837), .Z(n6840) );
  NANDN U9873 ( .A(n7010), .B(ereg[43]), .Z(n6839) );
  NAND U9874 ( .A(n6840), .B(n6839), .Z(n2271) );
  NAND U9875 ( .A(n7005), .B(ereg[41]), .Z(n6842) );
  NAND U9876 ( .A(n3926), .B(e[42]), .Z(n6841) );
  AND U9877 ( .A(n6842), .B(n6841), .Z(n6844) );
  NANDN U9878 ( .A(n7010), .B(ereg[42]), .Z(n6843) );
  NAND U9879 ( .A(n6844), .B(n6843), .Z(n2272) );
  NAND U9880 ( .A(n7005), .B(ereg[40]), .Z(n6846) );
  NAND U9881 ( .A(n3926), .B(e[41]), .Z(n6845) );
  AND U9882 ( .A(n6846), .B(n6845), .Z(n6848) );
  NANDN U9883 ( .A(n7010), .B(ereg[41]), .Z(n6847) );
  NAND U9884 ( .A(n6848), .B(n6847), .Z(n2273) );
  NAND U9885 ( .A(n7005), .B(ereg[39]), .Z(n6850) );
  NAND U9886 ( .A(n3926), .B(e[40]), .Z(n6849) );
  AND U9887 ( .A(n6850), .B(n6849), .Z(n6852) );
  NANDN U9888 ( .A(n7010), .B(ereg[40]), .Z(n6851) );
  NAND U9889 ( .A(n6852), .B(n6851), .Z(n2274) );
  NAND U9890 ( .A(n7005), .B(ereg[38]), .Z(n6854) );
  NAND U9891 ( .A(n3926), .B(e[39]), .Z(n6853) );
  AND U9892 ( .A(n6854), .B(n6853), .Z(n6856) );
  NANDN U9893 ( .A(n7010), .B(ereg[39]), .Z(n6855) );
  NAND U9894 ( .A(n6856), .B(n6855), .Z(n2275) );
  NAND U9895 ( .A(n7005), .B(ereg[37]), .Z(n6858) );
  NAND U9896 ( .A(n3927), .B(e[38]), .Z(n6857) );
  AND U9897 ( .A(n6858), .B(n6857), .Z(n6860) );
  NANDN U9898 ( .A(n7010), .B(ereg[38]), .Z(n6859) );
  NAND U9899 ( .A(n6860), .B(n6859), .Z(n2276) );
  NAND U9900 ( .A(n7005), .B(ereg[36]), .Z(n6862) );
  NAND U9901 ( .A(n3927), .B(e[37]), .Z(n6861) );
  AND U9902 ( .A(n6862), .B(n6861), .Z(n6864) );
  NANDN U9903 ( .A(n7010), .B(ereg[37]), .Z(n6863) );
  NAND U9904 ( .A(n6864), .B(n6863), .Z(n2277) );
  NAND U9905 ( .A(n7005), .B(ereg[35]), .Z(n6866) );
  NAND U9906 ( .A(n3927), .B(e[36]), .Z(n6865) );
  AND U9907 ( .A(n6866), .B(n6865), .Z(n6868) );
  NANDN U9908 ( .A(n7010), .B(ereg[36]), .Z(n6867) );
  NAND U9909 ( .A(n6868), .B(n6867), .Z(n2278) );
  NAND U9910 ( .A(n7005), .B(ereg[34]), .Z(n6870) );
  NAND U9911 ( .A(n3927), .B(e[35]), .Z(n6869) );
  AND U9912 ( .A(n6870), .B(n6869), .Z(n6872) );
  NANDN U9913 ( .A(n7010), .B(ereg[35]), .Z(n6871) );
  NAND U9914 ( .A(n6872), .B(n6871), .Z(n2279) );
  NAND U9915 ( .A(n7005), .B(ereg[33]), .Z(n6874) );
  NAND U9916 ( .A(n3927), .B(e[34]), .Z(n6873) );
  AND U9917 ( .A(n6874), .B(n6873), .Z(n6876) );
  NANDN U9918 ( .A(n7010), .B(ereg[34]), .Z(n6875) );
  NAND U9919 ( .A(n6876), .B(n6875), .Z(n2280) );
  NAND U9920 ( .A(n7005), .B(ereg[32]), .Z(n6878) );
  NAND U9921 ( .A(n3927), .B(e[33]), .Z(n6877) );
  AND U9922 ( .A(n6878), .B(n6877), .Z(n6880) );
  NANDN U9923 ( .A(n7010), .B(ereg[33]), .Z(n6879) );
  NAND U9924 ( .A(n6880), .B(n6879), .Z(n2281) );
  NAND U9925 ( .A(n7005), .B(ereg[31]), .Z(n6882) );
  NAND U9926 ( .A(n3927), .B(e[32]), .Z(n6881) );
  AND U9927 ( .A(n6882), .B(n6881), .Z(n6884) );
  NANDN U9928 ( .A(n7010), .B(ereg[32]), .Z(n6883) );
  NAND U9929 ( .A(n6884), .B(n6883), .Z(n2282) );
  NAND U9930 ( .A(n7005), .B(ereg[30]), .Z(n6886) );
  NAND U9931 ( .A(n3928), .B(e[31]), .Z(n6885) );
  AND U9932 ( .A(n6886), .B(n6885), .Z(n6888) );
  NANDN U9933 ( .A(n7010), .B(ereg[31]), .Z(n6887) );
  NAND U9934 ( .A(n6888), .B(n6887), .Z(n2283) );
  NAND U9935 ( .A(n7005), .B(ereg[29]), .Z(n6890) );
  NAND U9936 ( .A(n3928), .B(e[30]), .Z(n6889) );
  AND U9937 ( .A(n6890), .B(n6889), .Z(n6892) );
  NANDN U9938 ( .A(n7010), .B(ereg[30]), .Z(n6891) );
  NAND U9939 ( .A(n6892), .B(n6891), .Z(n2284) );
  NAND U9940 ( .A(n7005), .B(ereg[28]), .Z(n6894) );
  NAND U9941 ( .A(n3928), .B(e[29]), .Z(n6893) );
  AND U9942 ( .A(n6894), .B(n6893), .Z(n6896) );
  NANDN U9943 ( .A(n7010), .B(ereg[29]), .Z(n6895) );
  NAND U9944 ( .A(n6896), .B(n6895), .Z(n2285) );
  NAND U9945 ( .A(n7005), .B(ereg[27]), .Z(n6898) );
  NAND U9946 ( .A(n3928), .B(e[28]), .Z(n6897) );
  AND U9947 ( .A(n6898), .B(n6897), .Z(n6900) );
  NANDN U9948 ( .A(n7010), .B(ereg[28]), .Z(n6899) );
  NAND U9949 ( .A(n6900), .B(n6899), .Z(n2286) );
  NAND U9950 ( .A(n7005), .B(ereg[26]), .Z(n6902) );
  NAND U9951 ( .A(n3928), .B(e[27]), .Z(n6901) );
  AND U9952 ( .A(n6902), .B(n6901), .Z(n6904) );
  NANDN U9953 ( .A(n7010), .B(ereg[27]), .Z(n6903) );
  NAND U9954 ( .A(n6904), .B(n6903), .Z(n2287) );
  NAND U9955 ( .A(n7005), .B(ereg[25]), .Z(n6906) );
  NAND U9956 ( .A(n3928), .B(e[26]), .Z(n6905) );
  AND U9957 ( .A(n6906), .B(n6905), .Z(n6908) );
  NANDN U9958 ( .A(n7010), .B(ereg[26]), .Z(n6907) );
  NAND U9959 ( .A(n6908), .B(n6907), .Z(n2288) );
  NAND U9960 ( .A(n7005), .B(ereg[24]), .Z(n6910) );
  NAND U9961 ( .A(n3928), .B(e[25]), .Z(n6909) );
  AND U9962 ( .A(n6910), .B(n6909), .Z(n6912) );
  NANDN U9963 ( .A(n7010), .B(ereg[25]), .Z(n6911) );
  NAND U9964 ( .A(n6912), .B(n6911), .Z(n2289) );
  NAND U9965 ( .A(n7005), .B(ereg[23]), .Z(n6914) );
  NAND U9966 ( .A(n3929), .B(e[24]), .Z(n6913) );
  AND U9967 ( .A(n6914), .B(n6913), .Z(n6916) );
  NANDN U9968 ( .A(n7010), .B(ereg[24]), .Z(n6915) );
  NAND U9969 ( .A(n6916), .B(n6915), .Z(n2290) );
  NAND U9970 ( .A(n7005), .B(ereg[22]), .Z(n6918) );
  NAND U9971 ( .A(n3929), .B(e[23]), .Z(n6917) );
  AND U9972 ( .A(n6918), .B(n6917), .Z(n6920) );
  NANDN U9973 ( .A(n7010), .B(ereg[23]), .Z(n6919) );
  NAND U9974 ( .A(n6920), .B(n6919), .Z(n2291) );
  NAND U9975 ( .A(n7005), .B(ereg[21]), .Z(n6922) );
  NAND U9976 ( .A(n3929), .B(e[22]), .Z(n6921) );
  AND U9977 ( .A(n6922), .B(n6921), .Z(n6924) );
  NANDN U9978 ( .A(n7010), .B(ereg[22]), .Z(n6923) );
  NAND U9979 ( .A(n6924), .B(n6923), .Z(n2292) );
  NAND U9980 ( .A(n7005), .B(ereg[20]), .Z(n6926) );
  NAND U9981 ( .A(n3929), .B(e[21]), .Z(n6925) );
  AND U9982 ( .A(n6926), .B(n6925), .Z(n6928) );
  NANDN U9983 ( .A(n7010), .B(ereg[21]), .Z(n6927) );
  NAND U9984 ( .A(n6928), .B(n6927), .Z(n2293) );
  NAND U9985 ( .A(n7005), .B(ereg[19]), .Z(n6930) );
  NAND U9986 ( .A(n3929), .B(e[20]), .Z(n6929) );
  AND U9987 ( .A(n6930), .B(n6929), .Z(n6932) );
  NANDN U9988 ( .A(n7010), .B(ereg[20]), .Z(n6931) );
  NAND U9989 ( .A(n6932), .B(n6931), .Z(n2294) );
  NAND U9990 ( .A(n7005), .B(ereg[18]), .Z(n6934) );
  NAND U9991 ( .A(n3929), .B(e[19]), .Z(n6933) );
  AND U9992 ( .A(n6934), .B(n6933), .Z(n6936) );
  NANDN U9993 ( .A(n7010), .B(ereg[19]), .Z(n6935) );
  NAND U9994 ( .A(n6936), .B(n6935), .Z(n2295) );
  NAND U9995 ( .A(n7005), .B(ereg[17]), .Z(n6938) );
  NAND U9996 ( .A(n3929), .B(e[18]), .Z(n6937) );
  AND U9997 ( .A(n6938), .B(n6937), .Z(n6940) );
  NANDN U9998 ( .A(n7010), .B(ereg[18]), .Z(n6939) );
  NAND U9999 ( .A(n6940), .B(n6939), .Z(n2296) );
  NAND U10000 ( .A(n7005), .B(ereg[16]), .Z(n6942) );
  NAND U10001 ( .A(n3930), .B(e[17]), .Z(n6941) );
  AND U10002 ( .A(n6942), .B(n6941), .Z(n6944) );
  NANDN U10003 ( .A(n7010), .B(ereg[17]), .Z(n6943) );
  NAND U10004 ( .A(n6944), .B(n6943), .Z(n2297) );
  NAND U10005 ( .A(n7005), .B(ereg[15]), .Z(n6946) );
  NAND U10006 ( .A(n3930), .B(e[16]), .Z(n6945) );
  AND U10007 ( .A(n6946), .B(n6945), .Z(n6948) );
  NANDN U10008 ( .A(n7010), .B(ereg[16]), .Z(n6947) );
  NAND U10009 ( .A(n6948), .B(n6947), .Z(n2298) );
  NAND U10010 ( .A(n7005), .B(ereg[14]), .Z(n6950) );
  NAND U10011 ( .A(n3930), .B(e[15]), .Z(n6949) );
  AND U10012 ( .A(n6950), .B(n6949), .Z(n6952) );
  NANDN U10013 ( .A(n7010), .B(ereg[15]), .Z(n6951) );
  NAND U10014 ( .A(n6952), .B(n6951), .Z(n2299) );
  NAND U10015 ( .A(n7005), .B(ereg[13]), .Z(n6954) );
  NAND U10016 ( .A(n3930), .B(e[14]), .Z(n6953) );
  AND U10017 ( .A(n6954), .B(n6953), .Z(n6956) );
  NANDN U10018 ( .A(n7010), .B(ereg[14]), .Z(n6955) );
  NAND U10019 ( .A(n6956), .B(n6955), .Z(n2300) );
  NAND U10020 ( .A(n7005), .B(ereg[12]), .Z(n6958) );
  NAND U10021 ( .A(n3930), .B(e[13]), .Z(n6957) );
  AND U10022 ( .A(n6958), .B(n6957), .Z(n6960) );
  NANDN U10023 ( .A(n7010), .B(ereg[13]), .Z(n6959) );
  NAND U10024 ( .A(n6960), .B(n6959), .Z(n2301) );
  NAND U10025 ( .A(n7005), .B(ereg[11]), .Z(n6962) );
  NAND U10026 ( .A(n3930), .B(e[12]), .Z(n6961) );
  AND U10027 ( .A(n6962), .B(n6961), .Z(n6964) );
  NANDN U10028 ( .A(n7010), .B(ereg[12]), .Z(n6963) );
  NAND U10029 ( .A(n6964), .B(n6963), .Z(n2302) );
  NAND U10030 ( .A(n7005), .B(ereg[10]), .Z(n6966) );
  NAND U10031 ( .A(n3930), .B(e[11]), .Z(n6965) );
  AND U10032 ( .A(n6966), .B(n6965), .Z(n6968) );
  NANDN U10033 ( .A(n7010), .B(ereg[11]), .Z(n6967) );
  NAND U10034 ( .A(n6968), .B(n6967), .Z(n2303) );
  NAND U10035 ( .A(n7005), .B(ereg[9]), .Z(n6970) );
  NAND U10036 ( .A(n3931), .B(e[10]), .Z(n6969) );
  AND U10037 ( .A(n6970), .B(n6969), .Z(n6972) );
  NANDN U10038 ( .A(n7010), .B(ereg[10]), .Z(n6971) );
  NAND U10039 ( .A(n6972), .B(n6971), .Z(n2304) );
  NAND U10040 ( .A(n7005), .B(ereg[8]), .Z(n6974) );
  NAND U10041 ( .A(n3931), .B(e[9]), .Z(n6973) );
  AND U10042 ( .A(n6974), .B(n6973), .Z(n6976) );
  NANDN U10043 ( .A(n7010), .B(ereg[9]), .Z(n6975) );
  NAND U10044 ( .A(n6976), .B(n6975), .Z(n2305) );
  NAND U10045 ( .A(n7005), .B(ereg[7]), .Z(n6978) );
  NAND U10046 ( .A(n3931), .B(e[8]), .Z(n6977) );
  AND U10047 ( .A(n6978), .B(n6977), .Z(n6980) );
  NANDN U10048 ( .A(n7010), .B(ereg[8]), .Z(n6979) );
  NAND U10049 ( .A(n6980), .B(n6979), .Z(n2306) );
  NAND U10050 ( .A(n7005), .B(ereg[6]), .Z(n6982) );
  NAND U10051 ( .A(n3931), .B(e[7]), .Z(n6981) );
  AND U10052 ( .A(n6982), .B(n6981), .Z(n6984) );
  NANDN U10053 ( .A(n7010), .B(ereg[7]), .Z(n6983) );
  NAND U10054 ( .A(n6984), .B(n6983), .Z(n2307) );
  NAND U10055 ( .A(n7005), .B(ereg[5]), .Z(n6986) );
  NAND U10056 ( .A(n3931), .B(e[6]), .Z(n6985) );
  AND U10057 ( .A(n6986), .B(n6985), .Z(n6988) );
  NANDN U10058 ( .A(n7010), .B(ereg[6]), .Z(n6987) );
  NAND U10059 ( .A(n6988), .B(n6987), .Z(n2308) );
  NAND U10060 ( .A(n7005), .B(ereg[4]), .Z(n6990) );
  NAND U10061 ( .A(n3931), .B(e[5]), .Z(n6989) );
  AND U10062 ( .A(n6990), .B(n6989), .Z(n6992) );
  NANDN U10063 ( .A(n7010), .B(ereg[5]), .Z(n6991) );
  NAND U10064 ( .A(n6992), .B(n6991), .Z(n2309) );
  NAND U10065 ( .A(n7005), .B(ereg[3]), .Z(n6994) );
  NAND U10066 ( .A(n3931), .B(e[4]), .Z(n6993) );
  AND U10067 ( .A(n6994), .B(n6993), .Z(n6996) );
  NANDN U10068 ( .A(n7010), .B(ereg[4]), .Z(n6995) );
  NAND U10069 ( .A(n6996), .B(n6995), .Z(n2310) );
  NAND U10070 ( .A(n7005), .B(ereg[2]), .Z(n6998) );
  NAND U10071 ( .A(n3932), .B(e[3]), .Z(n6997) );
  AND U10072 ( .A(n6998), .B(n6997), .Z(n7000) );
  NANDN U10073 ( .A(n7010), .B(ereg[3]), .Z(n6999) );
  NAND U10074 ( .A(n7000), .B(n6999), .Z(n2311) );
  NAND U10075 ( .A(n7005), .B(ereg[1]), .Z(n7002) );
  NAND U10076 ( .A(n3932), .B(e[2]), .Z(n7001) );
  AND U10077 ( .A(n7002), .B(n7001), .Z(n7004) );
  NANDN U10078 ( .A(n7010), .B(ereg[2]), .Z(n7003) );
  NAND U10079 ( .A(n7004), .B(n7003), .Z(n2312) );
  NAND U10080 ( .A(n7005), .B(ereg[0]), .Z(n7007) );
  NAND U10081 ( .A(n3932), .B(e[1]), .Z(n7006) );
  AND U10082 ( .A(n7007), .B(n7006), .Z(n7009) );
  NANDN U10083 ( .A(n7010), .B(ereg[1]), .Z(n7008) );
  NAND U10084 ( .A(n7009), .B(n7008), .Z(n2313) );
  NAND U10085 ( .A(n3932), .B(e[0]), .Z(n7012) );
  NANDN U10086 ( .A(n7010), .B(ereg[0]), .Z(n7011) );
  NAND U10087 ( .A(n7012), .B(n7011), .Z(n2314) );
  XOR U10088 ( .A(start_in[511]), .B(mul_pow), .Z(n2315) );
endmodule

