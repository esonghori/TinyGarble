
module sum_N1024_CC2 ( clk, rst, a, b, c );
  input [511:0] a;
  input [511:0] b;
  output [511:0] c;
  input clk, rst;
  wire   N1026, N1027, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607;
  wire   [1:0] carry_on;

  DFF \carry_on_reg[1]  ( .D(N1027), .CLK(clk), .RST(rst), .Q(carry_on[1]) );
  DFF \carry_on_reg[0]  ( .D(N1026), .CLK(clk), .RST(rst), .Q(carry_on[0]) );
  DFF \rc_reg[511]  ( .D(n2048), .CLK(clk), .RST(1'b0), .Q(c[511]) );
  DFF \rc_reg[510]  ( .D(n2047), .CLK(clk), .RST(1'b0), .Q(c[510]) );
  DFF \rc_reg[509]  ( .D(n2046), .CLK(clk), .RST(1'b0), .Q(c[509]) );
  DFF \rc_reg[508]  ( .D(n2045), .CLK(clk), .RST(1'b0), .Q(c[508]) );
  DFF \rc_reg[507]  ( .D(n2044), .CLK(clk), .RST(1'b0), .Q(c[507]) );
  DFF \rc_reg[506]  ( .D(n2043), .CLK(clk), .RST(1'b0), .Q(c[506]) );
  DFF \rc_reg[505]  ( .D(n2042), .CLK(clk), .RST(1'b0), .Q(c[505]) );
  DFF \rc_reg[504]  ( .D(n2041), .CLK(clk), .RST(1'b0), .Q(c[504]) );
  DFF \rc_reg[503]  ( .D(n2040), .CLK(clk), .RST(1'b0), .Q(c[503]) );
  DFF \rc_reg[502]  ( .D(n2039), .CLK(clk), .RST(1'b0), .Q(c[502]) );
  DFF \rc_reg[501]  ( .D(n2038), .CLK(clk), .RST(1'b0), .Q(c[501]) );
  DFF \rc_reg[500]  ( .D(n2037), .CLK(clk), .RST(1'b0), .Q(c[500]) );
  DFF \rc_reg[499]  ( .D(n2036), .CLK(clk), .RST(1'b0), .Q(c[499]) );
  DFF \rc_reg[498]  ( .D(n2035), .CLK(clk), .RST(1'b0), .Q(c[498]) );
  DFF \rc_reg[497]  ( .D(n2034), .CLK(clk), .RST(1'b0), .Q(c[497]) );
  DFF \rc_reg[496]  ( .D(n2033), .CLK(clk), .RST(1'b0), .Q(c[496]) );
  DFF \rc_reg[495]  ( .D(n2032), .CLK(clk), .RST(1'b0), .Q(c[495]) );
  DFF \rc_reg[494]  ( .D(n2031), .CLK(clk), .RST(1'b0), .Q(c[494]) );
  DFF \rc_reg[493]  ( .D(n2030), .CLK(clk), .RST(1'b0), .Q(c[493]) );
  DFF \rc_reg[492]  ( .D(n2029), .CLK(clk), .RST(1'b0), .Q(c[492]) );
  DFF \rc_reg[491]  ( .D(n2028), .CLK(clk), .RST(1'b0), .Q(c[491]) );
  DFF \rc_reg[490]  ( .D(n2027), .CLK(clk), .RST(1'b0), .Q(c[490]) );
  DFF \rc_reg[489]  ( .D(n2026), .CLK(clk), .RST(1'b0), .Q(c[489]) );
  DFF \rc_reg[488]  ( .D(n2025), .CLK(clk), .RST(1'b0), .Q(c[488]) );
  DFF \rc_reg[487]  ( .D(n2024), .CLK(clk), .RST(1'b0), .Q(c[487]) );
  DFF \rc_reg[486]  ( .D(n2023), .CLK(clk), .RST(1'b0), .Q(c[486]) );
  DFF \rc_reg[485]  ( .D(n2022), .CLK(clk), .RST(1'b0), .Q(c[485]) );
  DFF \rc_reg[484]  ( .D(n2021), .CLK(clk), .RST(1'b0), .Q(c[484]) );
  DFF \rc_reg[483]  ( .D(n2020), .CLK(clk), .RST(1'b0), .Q(c[483]) );
  DFF \rc_reg[482]  ( .D(n2019), .CLK(clk), .RST(1'b0), .Q(c[482]) );
  DFF \rc_reg[481]  ( .D(n2018), .CLK(clk), .RST(1'b0), .Q(c[481]) );
  DFF \rc_reg[480]  ( .D(n2017), .CLK(clk), .RST(1'b0), .Q(c[480]) );
  DFF \rc_reg[479]  ( .D(n2016), .CLK(clk), .RST(1'b0), .Q(c[479]) );
  DFF \rc_reg[478]  ( .D(n2015), .CLK(clk), .RST(1'b0), .Q(c[478]) );
  DFF \rc_reg[477]  ( .D(n2014), .CLK(clk), .RST(1'b0), .Q(c[477]) );
  DFF \rc_reg[476]  ( .D(n2013), .CLK(clk), .RST(1'b0), .Q(c[476]) );
  DFF \rc_reg[475]  ( .D(n2012), .CLK(clk), .RST(1'b0), .Q(c[475]) );
  DFF \rc_reg[474]  ( .D(n2011), .CLK(clk), .RST(1'b0), .Q(c[474]) );
  DFF \rc_reg[473]  ( .D(n2010), .CLK(clk), .RST(1'b0), .Q(c[473]) );
  DFF \rc_reg[472]  ( .D(n2009), .CLK(clk), .RST(1'b0), .Q(c[472]) );
  DFF \rc_reg[471]  ( .D(n2008), .CLK(clk), .RST(1'b0), .Q(c[471]) );
  DFF \rc_reg[470]  ( .D(n2007), .CLK(clk), .RST(1'b0), .Q(c[470]) );
  DFF \rc_reg[469]  ( .D(n2006), .CLK(clk), .RST(1'b0), .Q(c[469]) );
  DFF \rc_reg[468]  ( .D(n2005), .CLK(clk), .RST(1'b0), .Q(c[468]) );
  DFF \rc_reg[467]  ( .D(n2004), .CLK(clk), .RST(1'b0), .Q(c[467]) );
  DFF \rc_reg[466]  ( .D(n2003), .CLK(clk), .RST(1'b0), .Q(c[466]) );
  DFF \rc_reg[465]  ( .D(n2002), .CLK(clk), .RST(1'b0), .Q(c[465]) );
  DFF \rc_reg[464]  ( .D(n2001), .CLK(clk), .RST(1'b0), .Q(c[464]) );
  DFF \rc_reg[463]  ( .D(n2000), .CLK(clk), .RST(1'b0), .Q(c[463]) );
  DFF \rc_reg[462]  ( .D(n1999), .CLK(clk), .RST(1'b0), .Q(c[462]) );
  DFF \rc_reg[461]  ( .D(n1998), .CLK(clk), .RST(1'b0), .Q(c[461]) );
  DFF \rc_reg[460]  ( .D(n1997), .CLK(clk), .RST(1'b0), .Q(c[460]) );
  DFF \rc_reg[459]  ( .D(n1996), .CLK(clk), .RST(1'b0), .Q(c[459]) );
  DFF \rc_reg[458]  ( .D(n1995), .CLK(clk), .RST(1'b0), .Q(c[458]) );
  DFF \rc_reg[457]  ( .D(n1994), .CLK(clk), .RST(1'b0), .Q(c[457]) );
  DFF \rc_reg[456]  ( .D(n1993), .CLK(clk), .RST(1'b0), .Q(c[456]) );
  DFF \rc_reg[455]  ( .D(n1992), .CLK(clk), .RST(1'b0), .Q(c[455]) );
  DFF \rc_reg[454]  ( .D(n1991), .CLK(clk), .RST(1'b0), .Q(c[454]) );
  DFF \rc_reg[453]  ( .D(n1990), .CLK(clk), .RST(1'b0), .Q(c[453]) );
  DFF \rc_reg[452]  ( .D(n1989), .CLK(clk), .RST(1'b0), .Q(c[452]) );
  DFF \rc_reg[451]  ( .D(n1988), .CLK(clk), .RST(1'b0), .Q(c[451]) );
  DFF \rc_reg[450]  ( .D(n1987), .CLK(clk), .RST(1'b0), .Q(c[450]) );
  DFF \rc_reg[449]  ( .D(n1986), .CLK(clk), .RST(1'b0), .Q(c[449]) );
  DFF \rc_reg[448]  ( .D(n1985), .CLK(clk), .RST(1'b0), .Q(c[448]) );
  DFF \rc_reg[447]  ( .D(n1984), .CLK(clk), .RST(1'b0), .Q(c[447]) );
  DFF \rc_reg[446]  ( .D(n1983), .CLK(clk), .RST(1'b0), .Q(c[446]) );
  DFF \rc_reg[445]  ( .D(n1982), .CLK(clk), .RST(1'b0), .Q(c[445]) );
  DFF \rc_reg[444]  ( .D(n1981), .CLK(clk), .RST(1'b0), .Q(c[444]) );
  DFF \rc_reg[443]  ( .D(n1980), .CLK(clk), .RST(1'b0), .Q(c[443]) );
  DFF \rc_reg[442]  ( .D(n1979), .CLK(clk), .RST(1'b0), .Q(c[442]) );
  DFF \rc_reg[441]  ( .D(n1978), .CLK(clk), .RST(1'b0), .Q(c[441]) );
  DFF \rc_reg[440]  ( .D(n1977), .CLK(clk), .RST(1'b0), .Q(c[440]) );
  DFF \rc_reg[439]  ( .D(n1976), .CLK(clk), .RST(1'b0), .Q(c[439]) );
  DFF \rc_reg[438]  ( .D(n1975), .CLK(clk), .RST(1'b0), .Q(c[438]) );
  DFF \rc_reg[437]  ( .D(n1974), .CLK(clk), .RST(1'b0), .Q(c[437]) );
  DFF \rc_reg[436]  ( .D(n1973), .CLK(clk), .RST(1'b0), .Q(c[436]) );
  DFF \rc_reg[435]  ( .D(n1972), .CLK(clk), .RST(1'b0), .Q(c[435]) );
  DFF \rc_reg[434]  ( .D(n1971), .CLK(clk), .RST(1'b0), .Q(c[434]) );
  DFF \rc_reg[433]  ( .D(n1970), .CLK(clk), .RST(1'b0), .Q(c[433]) );
  DFF \rc_reg[432]  ( .D(n1969), .CLK(clk), .RST(1'b0), .Q(c[432]) );
  DFF \rc_reg[431]  ( .D(n1968), .CLK(clk), .RST(1'b0), .Q(c[431]) );
  DFF \rc_reg[430]  ( .D(n1967), .CLK(clk), .RST(1'b0), .Q(c[430]) );
  DFF \rc_reg[429]  ( .D(n1966), .CLK(clk), .RST(1'b0), .Q(c[429]) );
  DFF \rc_reg[428]  ( .D(n1965), .CLK(clk), .RST(1'b0), .Q(c[428]) );
  DFF \rc_reg[427]  ( .D(n1964), .CLK(clk), .RST(1'b0), .Q(c[427]) );
  DFF \rc_reg[426]  ( .D(n1963), .CLK(clk), .RST(1'b0), .Q(c[426]) );
  DFF \rc_reg[425]  ( .D(n1962), .CLK(clk), .RST(1'b0), .Q(c[425]) );
  DFF \rc_reg[424]  ( .D(n1961), .CLK(clk), .RST(1'b0), .Q(c[424]) );
  DFF \rc_reg[423]  ( .D(n1960), .CLK(clk), .RST(1'b0), .Q(c[423]) );
  DFF \rc_reg[422]  ( .D(n1959), .CLK(clk), .RST(1'b0), .Q(c[422]) );
  DFF \rc_reg[421]  ( .D(n1958), .CLK(clk), .RST(1'b0), .Q(c[421]) );
  DFF \rc_reg[420]  ( .D(n1957), .CLK(clk), .RST(1'b0), .Q(c[420]) );
  DFF \rc_reg[419]  ( .D(n1956), .CLK(clk), .RST(1'b0), .Q(c[419]) );
  DFF \rc_reg[418]  ( .D(n1955), .CLK(clk), .RST(1'b0), .Q(c[418]) );
  DFF \rc_reg[417]  ( .D(n1954), .CLK(clk), .RST(1'b0), .Q(c[417]) );
  DFF \rc_reg[416]  ( .D(n1953), .CLK(clk), .RST(1'b0), .Q(c[416]) );
  DFF \rc_reg[415]  ( .D(n1952), .CLK(clk), .RST(1'b0), .Q(c[415]) );
  DFF \rc_reg[414]  ( .D(n1951), .CLK(clk), .RST(1'b0), .Q(c[414]) );
  DFF \rc_reg[413]  ( .D(n1950), .CLK(clk), .RST(1'b0), .Q(c[413]) );
  DFF \rc_reg[412]  ( .D(n1949), .CLK(clk), .RST(1'b0), .Q(c[412]) );
  DFF \rc_reg[411]  ( .D(n1948), .CLK(clk), .RST(1'b0), .Q(c[411]) );
  DFF \rc_reg[410]  ( .D(n1947), .CLK(clk), .RST(1'b0), .Q(c[410]) );
  DFF \rc_reg[409]  ( .D(n1946), .CLK(clk), .RST(1'b0), .Q(c[409]) );
  DFF \rc_reg[408]  ( .D(n1945), .CLK(clk), .RST(1'b0), .Q(c[408]) );
  DFF \rc_reg[407]  ( .D(n1944), .CLK(clk), .RST(1'b0), .Q(c[407]) );
  DFF \rc_reg[406]  ( .D(n1943), .CLK(clk), .RST(1'b0), .Q(c[406]) );
  DFF \rc_reg[405]  ( .D(n1942), .CLK(clk), .RST(1'b0), .Q(c[405]) );
  DFF \rc_reg[404]  ( .D(n1941), .CLK(clk), .RST(1'b0), .Q(c[404]) );
  DFF \rc_reg[403]  ( .D(n1940), .CLK(clk), .RST(1'b0), .Q(c[403]) );
  DFF \rc_reg[402]  ( .D(n1939), .CLK(clk), .RST(1'b0), .Q(c[402]) );
  DFF \rc_reg[401]  ( .D(n1938), .CLK(clk), .RST(1'b0), .Q(c[401]) );
  DFF \rc_reg[400]  ( .D(n1937), .CLK(clk), .RST(1'b0), .Q(c[400]) );
  DFF \rc_reg[399]  ( .D(n1936), .CLK(clk), .RST(1'b0), .Q(c[399]) );
  DFF \rc_reg[398]  ( .D(n1935), .CLK(clk), .RST(1'b0), .Q(c[398]) );
  DFF \rc_reg[397]  ( .D(n1934), .CLK(clk), .RST(1'b0), .Q(c[397]) );
  DFF \rc_reg[396]  ( .D(n1933), .CLK(clk), .RST(1'b0), .Q(c[396]) );
  DFF \rc_reg[395]  ( .D(n1932), .CLK(clk), .RST(1'b0), .Q(c[395]) );
  DFF \rc_reg[394]  ( .D(n1931), .CLK(clk), .RST(1'b0), .Q(c[394]) );
  DFF \rc_reg[393]  ( .D(n1930), .CLK(clk), .RST(1'b0), .Q(c[393]) );
  DFF \rc_reg[392]  ( .D(n1929), .CLK(clk), .RST(1'b0), .Q(c[392]) );
  DFF \rc_reg[391]  ( .D(n1928), .CLK(clk), .RST(1'b0), .Q(c[391]) );
  DFF \rc_reg[390]  ( .D(n1927), .CLK(clk), .RST(1'b0), .Q(c[390]) );
  DFF \rc_reg[389]  ( .D(n1926), .CLK(clk), .RST(1'b0), .Q(c[389]) );
  DFF \rc_reg[388]  ( .D(n1925), .CLK(clk), .RST(1'b0), .Q(c[388]) );
  DFF \rc_reg[387]  ( .D(n1924), .CLK(clk), .RST(1'b0), .Q(c[387]) );
  DFF \rc_reg[386]  ( .D(n1923), .CLK(clk), .RST(1'b0), .Q(c[386]) );
  DFF \rc_reg[385]  ( .D(n1922), .CLK(clk), .RST(1'b0), .Q(c[385]) );
  DFF \rc_reg[384]  ( .D(n1921), .CLK(clk), .RST(1'b0), .Q(c[384]) );
  DFF \rc_reg[383]  ( .D(n1920), .CLK(clk), .RST(1'b0), .Q(c[383]) );
  DFF \rc_reg[382]  ( .D(n1919), .CLK(clk), .RST(1'b0), .Q(c[382]) );
  DFF \rc_reg[381]  ( .D(n1918), .CLK(clk), .RST(1'b0), .Q(c[381]) );
  DFF \rc_reg[380]  ( .D(n1917), .CLK(clk), .RST(1'b0), .Q(c[380]) );
  DFF \rc_reg[379]  ( .D(n1916), .CLK(clk), .RST(1'b0), .Q(c[379]) );
  DFF \rc_reg[378]  ( .D(n1915), .CLK(clk), .RST(1'b0), .Q(c[378]) );
  DFF \rc_reg[377]  ( .D(n1914), .CLK(clk), .RST(1'b0), .Q(c[377]) );
  DFF \rc_reg[376]  ( .D(n1913), .CLK(clk), .RST(1'b0), .Q(c[376]) );
  DFF \rc_reg[375]  ( .D(n1912), .CLK(clk), .RST(1'b0), .Q(c[375]) );
  DFF \rc_reg[374]  ( .D(n1911), .CLK(clk), .RST(1'b0), .Q(c[374]) );
  DFF \rc_reg[373]  ( .D(n1910), .CLK(clk), .RST(1'b0), .Q(c[373]) );
  DFF \rc_reg[372]  ( .D(n1909), .CLK(clk), .RST(1'b0), .Q(c[372]) );
  DFF \rc_reg[371]  ( .D(n1908), .CLK(clk), .RST(1'b0), .Q(c[371]) );
  DFF \rc_reg[370]  ( .D(n1907), .CLK(clk), .RST(1'b0), .Q(c[370]) );
  DFF \rc_reg[369]  ( .D(n1906), .CLK(clk), .RST(1'b0), .Q(c[369]) );
  DFF \rc_reg[368]  ( .D(n1905), .CLK(clk), .RST(1'b0), .Q(c[368]) );
  DFF \rc_reg[367]  ( .D(n1904), .CLK(clk), .RST(1'b0), .Q(c[367]) );
  DFF \rc_reg[366]  ( .D(n1903), .CLK(clk), .RST(1'b0), .Q(c[366]) );
  DFF \rc_reg[365]  ( .D(n1902), .CLK(clk), .RST(1'b0), .Q(c[365]) );
  DFF \rc_reg[364]  ( .D(n1901), .CLK(clk), .RST(1'b0), .Q(c[364]) );
  DFF \rc_reg[363]  ( .D(n1900), .CLK(clk), .RST(1'b0), .Q(c[363]) );
  DFF \rc_reg[362]  ( .D(n1899), .CLK(clk), .RST(1'b0), .Q(c[362]) );
  DFF \rc_reg[361]  ( .D(n1898), .CLK(clk), .RST(1'b0), .Q(c[361]) );
  DFF \rc_reg[360]  ( .D(n1897), .CLK(clk), .RST(1'b0), .Q(c[360]) );
  DFF \rc_reg[359]  ( .D(n1896), .CLK(clk), .RST(1'b0), .Q(c[359]) );
  DFF \rc_reg[358]  ( .D(n1895), .CLK(clk), .RST(1'b0), .Q(c[358]) );
  DFF \rc_reg[357]  ( .D(n1894), .CLK(clk), .RST(1'b0), .Q(c[357]) );
  DFF \rc_reg[356]  ( .D(n1893), .CLK(clk), .RST(1'b0), .Q(c[356]) );
  DFF \rc_reg[355]  ( .D(n1892), .CLK(clk), .RST(1'b0), .Q(c[355]) );
  DFF \rc_reg[354]  ( .D(n1891), .CLK(clk), .RST(1'b0), .Q(c[354]) );
  DFF \rc_reg[353]  ( .D(n1890), .CLK(clk), .RST(1'b0), .Q(c[353]) );
  DFF \rc_reg[352]  ( .D(n1889), .CLK(clk), .RST(1'b0), .Q(c[352]) );
  DFF \rc_reg[351]  ( .D(n1888), .CLK(clk), .RST(1'b0), .Q(c[351]) );
  DFF \rc_reg[350]  ( .D(n1887), .CLK(clk), .RST(1'b0), .Q(c[350]) );
  DFF \rc_reg[349]  ( .D(n1886), .CLK(clk), .RST(1'b0), .Q(c[349]) );
  DFF \rc_reg[348]  ( .D(n1885), .CLK(clk), .RST(1'b0), .Q(c[348]) );
  DFF \rc_reg[347]  ( .D(n1884), .CLK(clk), .RST(1'b0), .Q(c[347]) );
  DFF \rc_reg[346]  ( .D(n1883), .CLK(clk), .RST(1'b0), .Q(c[346]) );
  DFF \rc_reg[345]  ( .D(n1882), .CLK(clk), .RST(1'b0), .Q(c[345]) );
  DFF \rc_reg[344]  ( .D(n1881), .CLK(clk), .RST(1'b0), .Q(c[344]) );
  DFF \rc_reg[343]  ( .D(n1880), .CLK(clk), .RST(1'b0), .Q(c[343]) );
  DFF \rc_reg[342]  ( .D(n1879), .CLK(clk), .RST(1'b0), .Q(c[342]) );
  DFF \rc_reg[341]  ( .D(n1878), .CLK(clk), .RST(1'b0), .Q(c[341]) );
  DFF \rc_reg[340]  ( .D(n1877), .CLK(clk), .RST(1'b0), .Q(c[340]) );
  DFF \rc_reg[339]  ( .D(n1876), .CLK(clk), .RST(1'b0), .Q(c[339]) );
  DFF \rc_reg[338]  ( .D(n1875), .CLK(clk), .RST(1'b0), .Q(c[338]) );
  DFF \rc_reg[337]  ( .D(n1874), .CLK(clk), .RST(1'b0), .Q(c[337]) );
  DFF \rc_reg[336]  ( .D(n1873), .CLK(clk), .RST(1'b0), .Q(c[336]) );
  DFF \rc_reg[335]  ( .D(n1872), .CLK(clk), .RST(1'b0), .Q(c[335]) );
  DFF \rc_reg[334]  ( .D(n1871), .CLK(clk), .RST(1'b0), .Q(c[334]) );
  DFF \rc_reg[333]  ( .D(n1870), .CLK(clk), .RST(1'b0), .Q(c[333]) );
  DFF \rc_reg[332]  ( .D(n1869), .CLK(clk), .RST(1'b0), .Q(c[332]) );
  DFF \rc_reg[331]  ( .D(n1868), .CLK(clk), .RST(1'b0), .Q(c[331]) );
  DFF \rc_reg[330]  ( .D(n1867), .CLK(clk), .RST(1'b0), .Q(c[330]) );
  DFF \rc_reg[329]  ( .D(n1866), .CLK(clk), .RST(1'b0), .Q(c[329]) );
  DFF \rc_reg[328]  ( .D(n1865), .CLK(clk), .RST(1'b0), .Q(c[328]) );
  DFF \rc_reg[327]  ( .D(n1864), .CLK(clk), .RST(1'b0), .Q(c[327]) );
  DFF \rc_reg[326]  ( .D(n1863), .CLK(clk), .RST(1'b0), .Q(c[326]) );
  DFF \rc_reg[325]  ( .D(n1862), .CLK(clk), .RST(1'b0), .Q(c[325]) );
  DFF \rc_reg[324]  ( .D(n1861), .CLK(clk), .RST(1'b0), .Q(c[324]) );
  DFF \rc_reg[323]  ( .D(n1860), .CLK(clk), .RST(1'b0), .Q(c[323]) );
  DFF \rc_reg[322]  ( .D(n1859), .CLK(clk), .RST(1'b0), .Q(c[322]) );
  DFF \rc_reg[321]  ( .D(n1858), .CLK(clk), .RST(1'b0), .Q(c[321]) );
  DFF \rc_reg[320]  ( .D(n1857), .CLK(clk), .RST(1'b0), .Q(c[320]) );
  DFF \rc_reg[319]  ( .D(n1856), .CLK(clk), .RST(1'b0), .Q(c[319]) );
  DFF \rc_reg[318]  ( .D(n1855), .CLK(clk), .RST(1'b0), .Q(c[318]) );
  DFF \rc_reg[317]  ( .D(n1854), .CLK(clk), .RST(1'b0), .Q(c[317]) );
  DFF \rc_reg[316]  ( .D(n1853), .CLK(clk), .RST(1'b0), .Q(c[316]) );
  DFF \rc_reg[315]  ( .D(n1852), .CLK(clk), .RST(1'b0), .Q(c[315]) );
  DFF \rc_reg[314]  ( .D(n1851), .CLK(clk), .RST(1'b0), .Q(c[314]) );
  DFF \rc_reg[313]  ( .D(n1850), .CLK(clk), .RST(1'b0), .Q(c[313]) );
  DFF \rc_reg[312]  ( .D(n1849), .CLK(clk), .RST(1'b0), .Q(c[312]) );
  DFF \rc_reg[311]  ( .D(n1848), .CLK(clk), .RST(1'b0), .Q(c[311]) );
  DFF \rc_reg[310]  ( .D(n1847), .CLK(clk), .RST(1'b0), .Q(c[310]) );
  DFF \rc_reg[309]  ( .D(n1846), .CLK(clk), .RST(1'b0), .Q(c[309]) );
  DFF \rc_reg[308]  ( .D(n1845), .CLK(clk), .RST(1'b0), .Q(c[308]) );
  DFF \rc_reg[307]  ( .D(n1844), .CLK(clk), .RST(1'b0), .Q(c[307]) );
  DFF \rc_reg[306]  ( .D(n1843), .CLK(clk), .RST(1'b0), .Q(c[306]) );
  DFF \rc_reg[305]  ( .D(n1842), .CLK(clk), .RST(1'b0), .Q(c[305]) );
  DFF \rc_reg[304]  ( .D(n1841), .CLK(clk), .RST(1'b0), .Q(c[304]) );
  DFF \rc_reg[303]  ( .D(n1840), .CLK(clk), .RST(1'b0), .Q(c[303]) );
  DFF \rc_reg[302]  ( .D(n1839), .CLK(clk), .RST(1'b0), .Q(c[302]) );
  DFF \rc_reg[301]  ( .D(n1838), .CLK(clk), .RST(1'b0), .Q(c[301]) );
  DFF \rc_reg[300]  ( .D(n1837), .CLK(clk), .RST(1'b0), .Q(c[300]) );
  DFF \rc_reg[299]  ( .D(n1836), .CLK(clk), .RST(1'b0), .Q(c[299]) );
  DFF \rc_reg[298]  ( .D(n1835), .CLK(clk), .RST(1'b0), .Q(c[298]) );
  DFF \rc_reg[297]  ( .D(n1834), .CLK(clk), .RST(1'b0), .Q(c[297]) );
  DFF \rc_reg[296]  ( .D(n1833), .CLK(clk), .RST(1'b0), .Q(c[296]) );
  DFF \rc_reg[295]  ( .D(n1832), .CLK(clk), .RST(1'b0), .Q(c[295]) );
  DFF \rc_reg[294]  ( .D(n1831), .CLK(clk), .RST(1'b0), .Q(c[294]) );
  DFF \rc_reg[293]  ( .D(n1830), .CLK(clk), .RST(1'b0), .Q(c[293]) );
  DFF \rc_reg[292]  ( .D(n1829), .CLK(clk), .RST(1'b0), .Q(c[292]) );
  DFF \rc_reg[291]  ( .D(n1828), .CLK(clk), .RST(1'b0), .Q(c[291]) );
  DFF \rc_reg[290]  ( .D(n1827), .CLK(clk), .RST(1'b0), .Q(c[290]) );
  DFF \rc_reg[289]  ( .D(n1826), .CLK(clk), .RST(1'b0), .Q(c[289]) );
  DFF \rc_reg[288]  ( .D(n1825), .CLK(clk), .RST(1'b0), .Q(c[288]) );
  DFF \rc_reg[287]  ( .D(n1824), .CLK(clk), .RST(1'b0), .Q(c[287]) );
  DFF \rc_reg[286]  ( .D(n1823), .CLK(clk), .RST(1'b0), .Q(c[286]) );
  DFF \rc_reg[285]  ( .D(n1822), .CLK(clk), .RST(1'b0), .Q(c[285]) );
  DFF \rc_reg[284]  ( .D(n1821), .CLK(clk), .RST(1'b0), .Q(c[284]) );
  DFF \rc_reg[283]  ( .D(n1820), .CLK(clk), .RST(1'b0), .Q(c[283]) );
  DFF \rc_reg[282]  ( .D(n1819), .CLK(clk), .RST(1'b0), .Q(c[282]) );
  DFF \rc_reg[281]  ( .D(n1818), .CLK(clk), .RST(1'b0), .Q(c[281]) );
  DFF \rc_reg[280]  ( .D(n1817), .CLK(clk), .RST(1'b0), .Q(c[280]) );
  DFF \rc_reg[279]  ( .D(n1816), .CLK(clk), .RST(1'b0), .Q(c[279]) );
  DFF \rc_reg[278]  ( .D(n1815), .CLK(clk), .RST(1'b0), .Q(c[278]) );
  DFF \rc_reg[277]  ( .D(n1814), .CLK(clk), .RST(1'b0), .Q(c[277]) );
  DFF \rc_reg[276]  ( .D(n1813), .CLK(clk), .RST(1'b0), .Q(c[276]) );
  DFF \rc_reg[275]  ( .D(n1812), .CLK(clk), .RST(1'b0), .Q(c[275]) );
  DFF \rc_reg[274]  ( .D(n1811), .CLK(clk), .RST(1'b0), .Q(c[274]) );
  DFF \rc_reg[273]  ( .D(n1810), .CLK(clk), .RST(1'b0), .Q(c[273]) );
  DFF \rc_reg[272]  ( .D(n1809), .CLK(clk), .RST(1'b0), .Q(c[272]) );
  DFF \rc_reg[271]  ( .D(n1808), .CLK(clk), .RST(1'b0), .Q(c[271]) );
  DFF \rc_reg[270]  ( .D(n1807), .CLK(clk), .RST(1'b0), .Q(c[270]) );
  DFF \rc_reg[269]  ( .D(n1806), .CLK(clk), .RST(1'b0), .Q(c[269]) );
  DFF \rc_reg[268]  ( .D(n1805), .CLK(clk), .RST(1'b0), .Q(c[268]) );
  DFF \rc_reg[267]  ( .D(n1804), .CLK(clk), .RST(1'b0), .Q(c[267]) );
  DFF \rc_reg[266]  ( .D(n1803), .CLK(clk), .RST(1'b0), .Q(c[266]) );
  DFF \rc_reg[265]  ( .D(n1802), .CLK(clk), .RST(1'b0), .Q(c[265]) );
  DFF \rc_reg[264]  ( .D(n1801), .CLK(clk), .RST(1'b0), .Q(c[264]) );
  DFF \rc_reg[263]  ( .D(n1800), .CLK(clk), .RST(1'b0), .Q(c[263]) );
  DFF \rc_reg[262]  ( .D(n1799), .CLK(clk), .RST(1'b0), .Q(c[262]) );
  DFF \rc_reg[261]  ( .D(n1798), .CLK(clk), .RST(1'b0), .Q(c[261]) );
  DFF \rc_reg[260]  ( .D(n1797), .CLK(clk), .RST(1'b0), .Q(c[260]) );
  DFF \rc_reg[259]  ( .D(n1796), .CLK(clk), .RST(1'b0), .Q(c[259]) );
  DFF \rc_reg[258]  ( .D(n1795), .CLK(clk), .RST(1'b0), .Q(c[258]) );
  DFF \rc_reg[257]  ( .D(n1794), .CLK(clk), .RST(1'b0), .Q(c[257]) );
  DFF \rc_reg[256]  ( .D(n1793), .CLK(clk), .RST(1'b0), .Q(c[256]) );
  DFF \rc_reg[255]  ( .D(n1792), .CLK(clk), .RST(1'b0), .Q(c[255]) );
  DFF \rc_reg[254]  ( .D(n1791), .CLK(clk), .RST(1'b0), .Q(c[254]) );
  DFF \rc_reg[253]  ( .D(n1790), .CLK(clk), .RST(1'b0), .Q(c[253]) );
  DFF \rc_reg[252]  ( .D(n1789), .CLK(clk), .RST(1'b0), .Q(c[252]) );
  DFF \rc_reg[251]  ( .D(n1788), .CLK(clk), .RST(1'b0), .Q(c[251]) );
  DFF \rc_reg[250]  ( .D(n1787), .CLK(clk), .RST(1'b0), .Q(c[250]) );
  DFF \rc_reg[249]  ( .D(n1786), .CLK(clk), .RST(1'b0), .Q(c[249]) );
  DFF \rc_reg[248]  ( .D(n1785), .CLK(clk), .RST(1'b0), .Q(c[248]) );
  DFF \rc_reg[247]  ( .D(n1784), .CLK(clk), .RST(1'b0), .Q(c[247]) );
  DFF \rc_reg[246]  ( .D(n1783), .CLK(clk), .RST(1'b0), .Q(c[246]) );
  DFF \rc_reg[245]  ( .D(n1782), .CLK(clk), .RST(1'b0), .Q(c[245]) );
  DFF \rc_reg[244]  ( .D(n1781), .CLK(clk), .RST(1'b0), .Q(c[244]) );
  DFF \rc_reg[243]  ( .D(n1780), .CLK(clk), .RST(1'b0), .Q(c[243]) );
  DFF \rc_reg[242]  ( .D(n1779), .CLK(clk), .RST(1'b0), .Q(c[242]) );
  DFF \rc_reg[241]  ( .D(n1778), .CLK(clk), .RST(1'b0), .Q(c[241]) );
  DFF \rc_reg[240]  ( .D(n1777), .CLK(clk), .RST(1'b0), .Q(c[240]) );
  DFF \rc_reg[239]  ( .D(n1776), .CLK(clk), .RST(1'b0), .Q(c[239]) );
  DFF \rc_reg[238]  ( .D(n1775), .CLK(clk), .RST(1'b0), .Q(c[238]) );
  DFF \rc_reg[237]  ( .D(n1774), .CLK(clk), .RST(1'b0), .Q(c[237]) );
  DFF \rc_reg[236]  ( .D(n1773), .CLK(clk), .RST(1'b0), .Q(c[236]) );
  DFF \rc_reg[235]  ( .D(n1772), .CLK(clk), .RST(1'b0), .Q(c[235]) );
  DFF \rc_reg[234]  ( .D(n1771), .CLK(clk), .RST(1'b0), .Q(c[234]) );
  DFF \rc_reg[233]  ( .D(n1770), .CLK(clk), .RST(1'b0), .Q(c[233]) );
  DFF \rc_reg[232]  ( .D(n1769), .CLK(clk), .RST(1'b0), .Q(c[232]) );
  DFF \rc_reg[231]  ( .D(n1768), .CLK(clk), .RST(1'b0), .Q(c[231]) );
  DFF \rc_reg[230]  ( .D(n1767), .CLK(clk), .RST(1'b0), .Q(c[230]) );
  DFF \rc_reg[229]  ( .D(n1766), .CLK(clk), .RST(1'b0), .Q(c[229]) );
  DFF \rc_reg[228]  ( .D(n1765), .CLK(clk), .RST(1'b0), .Q(c[228]) );
  DFF \rc_reg[227]  ( .D(n1764), .CLK(clk), .RST(1'b0), .Q(c[227]) );
  DFF \rc_reg[226]  ( .D(n1763), .CLK(clk), .RST(1'b0), .Q(c[226]) );
  DFF \rc_reg[225]  ( .D(n1762), .CLK(clk), .RST(1'b0), .Q(c[225]) );
  DFF \rc_reg[224]  ( .D(n1761), .CLK(clk), .RST(1'b0), .Q(c[224]) );
  DFF \rc_reg[223]  ( .D(n1760), .CLK(clk), .RST(1'b0), .Q(c[223]) );
  DFF \rc_reg[222]  ( .D(n1759), .CLK(clk), .RST(1'b0), .Q(c[222]) );
  DFF \rc_reg[221]  ( .D(n1758), .CLK(clk), .RST(1'b0), .Q(c[221]) );
  DFF \rc_reg[220]  ( .D(n1757), .CLK(clk), .RST(1'b0), .Q(c[220]) );
  DFF \rc_reg[219]  ( .D(n1756), .CLK(clk), .RST(1'b0), .Q(c[219]) );
  DFF \rc_reg[218]  ( .D(n1755), .CLK(clk), .RST(1'b0), .Q(c[218]) );
  DFF \rc_reg[217]  ( .D(n1754), .CLK(clk), .RST(1'b0), .Q(c[217]) );
  DFF \rc_reg[216]  ( .D(n1753), .CLK(clk), .RST(1'b0), .Q(c[216]) );
  DFF \rc_reg[215]  ( .D(n1752), .CLK(clk), .RST(1'b0), .Q(c[215]) );
  DFF \rc_reg[214]  ( .D(n1751), .CLK(clk), .RST(1'b0), .Q(c[214]) );
  DFF \rc_reg[213]  ( .D(n1750), .CLK(clk), .RST(1'b0), .Q(c[213]) );
  DFF \rc_reg[212]  ( .D(n1749), .CLK(clk), .RST(1'b0), .Q(c[212]) );
  DFF \rc_reg[211]  ( .D(n1748), .CLK(clk), .RST(1'b0), .Q(c[211]) );
  DFF \rc_reg[210]  ( .D(n1747), .CLK(clk), .RST(1'b0), .Q(c[210]) );
  DFF \rc_reg[209]  ( .D(n1746), .CLK(clk), .RST(1'b0), .Q(c[209]) );
  DFF \rc_reg[208]  ( .D(n1745), .CLK(clk), .RST(1'b0), .Q(c[208]) );
  DFF \rc_reg[207]  ( .D(n1744), .CLK(clk), .RST(1'b0), .Q(c[207]) );
  DFF \rc_reg[206]  ( .D(n1743), .CLK(clk), .RST(1'b0), .Q(c[206]) );
  DFF \rc_reg[205]  ( .D(n1742), .CLK(clk), .RST(1'b0), .Q(c[205]) );
  DFF \rc_reg[204]  ( .D(n1741), .CLK(clk), .RST(1'b0), .Q(c[204]) );
  DFF \rc_reg[203]  ( .D(n1740), .CLK(clk), .RST(1'b0), .Q(c[203]) );
  DFF \rc_reg[202]  ( .D(n1739), .CLK(clk), .RST(1'b0), .Q(c[202]) );
  DFF \rc_reg[201]  ( .D(n1738), .CLK(clk), .RST(1'b0), .Q(c[201]) );
  DFF \rc_reg[200]  ( .D(n1737), .CLK(clk), .RST(1'b0), .Q(c[200]) );
  DFF \rc_reg[199]  ( .D(n1736), .CLK(clk), .RST(1'b0), .Q(c[199]) );
  DFF \rc_reg[198]  ( .D(n1735), .CLK(clk), .RST(1'b0), .Q(c[198]) );
  DFF \rc_reg[197]  ( .D(n1734), .CLK(clk), .RST(1'b0), .Q(c[197]) );
  DFF \rc_reg[196]  ( .D(n1733), .CLK(clk), .RST(1'b0), .Q(c[196]) );
  DFF \rc_reg[195]  ( .D(n1732), .CLK(clk), .RST(1'b0), .Q(c[195]) );
  DFF \rc_reg[194]  ( .D(n1731), .CLK(clk), .RST(1'b0), .Q(c[194]) );
  DFF \rc_reg[193]  ( .D(n1730), .CLK(clk), .RST(1'b0), .Q(c[193]) );
  DFF \rc_reg[192]  ( .D(n1729), .CLK(clk), .RST(1'b0), .Q(c[192]) );
  DFF \rc_reg[191]  ( .D(n1728), .CLK(clk), .RST(1'b0), .Q(c[191]) );
  DFF \rc_reg[190]  ( .D(n1727), .CLK(clk), .RST(1'b0), .Q(c[190]) );
  DFF \rc_reg[189]  ( .D(n1726), .CLK(clk), .RST(1'b0), .Q(c[189]) );
  DFF \rc_reg[188]  ( .D(n1725), .CLK(clk), .RST(1'b0), .Q(c[188]) );
  DFF \rc_reg[187]  ( .D(n1724), .CLK(clk), .RST(1'b0), .Q(c[187]) );
  DFF \rc_reg[186]  ( .D(n1723), .CLK(clk), .RST(1'b0), .Q(c[186]) );
  DFF \rc_reg[185]  ( .D(n1722), .CLK(clk), .RST(1'b0), .Q(c[185]) );
  DFF \rc_reg[184]  ( .D(n1721), .CLK(clk), .RST(1'b0), .Q(c[184]) );
  DFF \rc_reg[183]  ( .D(n1720), .CLK(clk), .RST(1'b0), .Q(c[183]) );
  DFF \rc_reg[182]  ( .D(n1719), .CLK(clk), .RST(1'b0), .Q(c[182]) );
  DFF \rc_reg[181]  ( .D(n1718), .CLK(clk), .RST(1'b0), .Q(c[181]) );
  DFF \rc_reg[180]  ( .D(n1717), .CLK(clk), .RST(1'b0), .Q(c[180]) );
  DFF \rc_reg[179]  ( .D(n1716), .CLK(clk), .RST(1'b0), .Q(c[179]) );
  DFF \rc_reg[178]  ( .D(n1715), .CLK(clk), .RST(1'b0), .Q(c[178]) );
  DFF \rc_reg[177]  ( .D(n1714), .CLK(clk), .RST(1'b0), .Q(c[177]) );
  DFF \rc_reg[176]  ( .D(n1713), .CLK(clk), .RST(1'b0), .Q(c[176]) );
  DFF \rc_reg[175]  ( .D(n1712), .CLK(clk), .RST(1'b0), .Q(c[175]) );
  DFF \rc_reg[174]  ( .D(n1711), .CLK(clk), .RST(1'b0), .Q(c[174]) );
  DFF \rc_reg[173]  ( .D(n1710), .CLK(clk), .RST(1'b0), .Q(c[173]) );
  DFF \rc_reg[172]  ( .D(n1709), .CLK(clk), .RST(1'b0), .Q(c[172]) );
  DFF \rc_reg[171]  ( .D(n1708), .CLK(clk), .RST(1'b0), .Q(c[171]) );
  DFF \rc_reg[170]  ( .D(n1707), .CLK(clk), .RST(1'b0), .Q(c[170]) );
  DFF \rc_reg[169]  ( .D(n1706), .CLK(clk), .RST(1'b0), .Q(c[169]) );
  DFF \rc_reg[168]  ( .D(n1705), .CLK(clk), .RST(1'b0), .Q(c[168]) );
  DFF \rc_reg[167]  ( .D(n1704), .CLK(clk), .RST(1'b0), .Q(c[167]) );
  DFF \rc_reg[166]  ( .D(n1703), .CLK(clk), .RST(1'b0), .Q(c[166]) );
  DFF \rc_reg[165]  ( .D(n1702), .CLK(clk), .RST(1'b0), .Q(c[165]) );
  DFF \rc_reg[164]  ( .D(n1701), .CLK(clk), .RST(1'b0), .Q(c[164]) );
  DFF \rc_reg[163]  ( .D(n1700), .CLK(clk), .RST(1'b0), .Q(c[163]) );
  DFF \rc_reg[162]  ( .D(n1699), .CLK(clk), .RST(1'b0), .Q(c[162]) );
  DFF \rc_reg[161]  ( .D(n1698), .CLK(clk), .RST(1'b0), .Q(c[161]) );
  DFF \rc_reg[160]  ( .D(n1697), .CLK(clk), .RST(1'b0), .Q(c[160]) );
  DFF \rc_reg[159]  ( .D(n1696), .CLK(clk), .RST(1'b0), .Q(c[159]) );
  DFF \rc_reg[158]  ( .D(n1695), .CLK(clk), .RST(1'b0), .Q(c[158]) );
  DFF \rc_reg[157]  ( .D(n1694), .CLK(clk), .RST(1'b0), .Q(c[157]) );
  DFF \rc_reg[156]  ( .D(n1693), .CLK(clk), .RST(1'b0), .Q(c[156]) );
  DFF \rc_reg[155]  ( .D(n1692), .CLK(clk), .RST(1'b0), .Q(c[155]) );
  DFF \rc_reg[154]  ( .D(n1691), .CLK(clk), .RST(1'b0), .Q(c[154]) );
  DFF \rc_reg[153]  ( .D(n1690), .CLK(clk), .RST(1'b0), .Q(c[153]) );
  DFF \rc_reg[152]  ( .D(n1689), .CLK(clk), .RST(1'b0), .Q(c[152]) );
  DFF \rc_reg[151]  ( .D(n1688), .CLK(clk), .RST(1'b0), .Q(c[151]) );
  DFF \rc_reg[150]  ( .D(n1687), .CLK(clk), .RST(1'b0), .Q(c[150]) );
  DFF \rc_reg[149]  ( .D(n1686), .CLK(clk), .RST(1'b0), .Q(c[149]) );
  DFF \rc_reg[148]  ( .D(n1685), .CLK(clk), .RST(1'b0), .Q(c[148]) );
  DFF \rc_reg[147]  ( .D(n1684), .CLK(clk), .RST(1'b0), .Q(c[147]) );
  DFF \rc_reg[146]  ( .D(n1683), .CLK(clk), .RST(1'b0), .Q(c[146]) );
  DFF \rc_reg[145]  ( .D(n1682), .CLK(clk), .RST(1'b0), .Q(c[145]) );
  DFF \rc_reg[144]  ( .D(n1681), .CLK(clk), .RST(1'b0), .Q(c[144]) );
  DFF \rc_reg[143]  ( .D(n1680), .CLK(clk), .RST(1'b0), .Q(c[143]) );
  DFF \rc_reg[142]  ( .D(n1679), .CLK(clk), .RST(1'b0), .Q(c[142]) );
  DFF \rc_reg[141]  ( .D(n1678), .CLK(clk), .RST(1'b0), .Q(c[141]) );
  DFF \rc_reg[140]  ( .D(n1677), .CLK(clk), .RST(1'b0), .Q(c[140]) );
  DFF \rc_reg[139]  ( .D(n1676), .CLK(clk), .RST(1'b0), .Q(c[139]) );
  DFF \rc_reg[138]  ( .D(n1675), .CLK(clk), .RST(1'b0), .Q(c[138]) );
  DFF \rc_reg[137]  ( .D(n1674), .CLK(clk), .RST(1'b0), .Q(c[137]) );
  DFF \rc_reg[136]  ( .D(n1673), .CLK(clk), .RST(1'b0), .Q(c[136]) );
  DFF \rc_reg[135]  ( .D(n1672), .CLK(clk), .RST(1'b0), .Q(c[135]) );
  DFF \rc_reg[134]  ( .D(n1671), .CLK(clk), .RST(1'b0), .Q(c[134]) );
  DFF \rc_reg[133]  ( .D(n1670), .CLK(clk), .RST(1'b0), .Q(c[133]) );
  DFF \rc_reg[132]  ( .D(n1669), .CLK(clk), .RST(1'b0), .Q(c[132]) );
  DFF \rc_reg[131]  ( .D(n1668), .CLK(clk), .RST(1'b0), .Q(c[131]) );
  DFF \rc_reg[130]  ( .D(n1667), .CLK(clk), .RST(1'b0), .Q(c[130]) );
  DFF \rc_reg[129]  ( .D(n1666), .CLK(clk), .RST(1'b0), .Q(c[129]) );
  DFF \rc_reg[128]  ( .D(n1665), .CLK(clk), .RST(1'b0), .Q(c[128]) );
  DFF \rc_reg[127]  ( .D(n1664), .CLK(clk), .RST(1'b0), .Q(c[127]) );
  DFF \rc_reg[126]  ( .D(n1663), .CLK(clk), .RST(1'b0), .Q(c[126]) );
  DFF \rc_reg[125]  ( .D(n1662), .CLK(clk), .RST(1'b0), .Q(c[125]) );
  DFF \rc_reg[124]  ( .D(n1661), .CLK(clk), .RST(1'b0), .Q(c[124]) );
  DFF \rc_reg[123]  ( .D(n1660), .CLK(clk), .RST(1'b0), .Q(c[123]) );
  DFF \rc_reg[122]  ( .D(n1659), .CLK(clk), .RST(1'b0), .Q(c[122]) );
  DFF \rc_reg[121]  ( .D(n1658), .CLK(clk), .RST(1'b0), .Q(c[121]) );
  DFF \rc_reg[120]  ( .D(n1657), .CLK(clk), .RST(1'b0), .Q(c[120]) );
  DFF \rc_reg[119]  ( .D(n1656), .CLK(clk), .RST(1'b0), .Q(c[119]) );
  DFF \rc_reg[118]  ( .D(n1655), .CLK(clk), .RST(1'b0), .Q(c[118]) );
  DFF \rc_reg[117]  ( .D(n1654), .CLK(clk), .RST(1'b0), .Q(c[117]) );
  DFF \rc_reg[116]  ( .D(n1653), .CLK(clk), .RST(1'b0), .Q(c[116]) );
  DFF \rc_reg[115]  ( .D(n1652), .CLK(clk), .RST(1'b0), .Q(c[115]) );
  DFF \rc_reg[114]  ( .D(n1651), .CLK(clk), .RST(1'b0), .Q(c[114]) );
  DFF \rc_reg[113]  ( .D(n1650), .CLK(clk), .RST(1'b0), .Q(c[113]) );
  DFF \rc_reg[112]  ( .D(n1649), .CLK(clk), .RST(1'b0), .Q(c[112]) );
  DFF \rc_reg[111]  ( .D(n1648), .CLK(clk), .RST(1'b0), .Q(c[111]) );
  DFF \rc_reg[110]  ( .D(n1647), .CLK(clk), .RST(1'b0), .Q(c[110]) );
  DFF \rc_reg[109]  ( .D(n1646), .CLK(clk), .RST(1'b0), .Q(c[109]) );
  DFF \rc_reg[108]  ( .D(n1645), .CLK(clk), .RST(1'b0), .Q(c[108]) );
  DFF \rc_reg[107]  ( .D(n1644), .CLK(clk), .RST(1'b0), .Q(c[107]) );
  DFF \rc_reg[106]  ( .D(n1643), .CLK(clk), .RST(1'b0), .Q(c[106]) );
  DFF \rc_reg[105]  ( .D(n1642), .CLK(clk), .RST(1'b0), .Q(c[105]) );
  DFF \rc_reg[104]  ( .D(n1641), .CLK(clk), .RST(1'b0), .Q(c[104]) );
  DFF \rc_reg[103]  ( .D(n1640), .CLK(clk), .RST(1'b0), .Q(c[103]) );
  DFF \rc_reg[102]  ( .D(n1639), .CLK(clk), .RST(1'b0), .Q(c[102]) );
  DFF \rc_reg[101]  ( .D(n1638), .CLK(clk), .RST(1'b0), .Q(c[101]) );
  DFF \rc_reg[100]  ( .D(n1637), .CLK(clk), .RST(1'b0), .Q(c[100]) );
  DFF \rc_reg[99]  ( .D(n1636), .CLK(clk), .RST(1'b0), .Q(c[99]) );
  DFF \rc_reg[98]  ( .D(n1635), .CLK(clk), .RST(1'b0), .Q(c[98]) );
  DFF \rc_reg[97]  ( .D(n1634), .CLK(clk), .RST(1'b0), .Q(c[97]) );
  DFF \rc_reg[96]  ( .D(n1633), .CLK(clk), .RST(1'b0), .Q(c[96]) );
  DFF \rc_reg[95]  ( .D(n1632), .CLK(clk), .RST(1'b0), .Q(c[95]) );
  DFF \rc_reg[94]  ( .D(n1631), .CLK(clk), .RST(1'b0), .Q(c[94]) );
  DFF \rc_reg[93]  ( .D(n1630), .CLK(clk), .RST(1'b0), .Q(c[93]) );
  DFF \rc_reg[92]  ( .D(n1629), .CLK(clk), .RST(1'b0), .Q(c[92]) );
  DFF \rc_reg[91]  ( .D(n1628), .CLK(clk), .RST(1'b0), .Q(c[91]) );
  DFF \rc_reg[90]  ( .D(n1627), .CLK(clk), .RST(1'b0), .Q(c[90]) );
  DFF \rc_reg[89]  ( .D(n1626), .CLK(clk), .RST(1'b0), .Q(c[89]) );
  DFF \rc_reg[88]  ( .D(n1625), .CLK(clk), .RST(1'b0), .Q(c[88]) );
  DFF \rc_reg[87]  ( .D(n1624), .CLK(clk), .RST(1'b0), .Q(c[87]) );
  DFF \rc_reg[86]  ( .D(n1623), .CLK(clk), .RST(1'b0), .Q(c[86]) );
  DFF \rc_reg[85]  ( .D(n1622), .CLK(clk), .RST(1'b0), .Q(c[85]) );
  DFF \rc_reg[84]  ( .D(n1621), .CLK(clk), .RST(1'b0), .Q(c[84]) );
  DFF \rc_reg[83]  ( .D(n1620), .CLK(clk), .RST(1'b0), .Q(c[83]) );
  DFF \rc_reg[82]  ( .D(n1619), .CLK(clk), .RST(1'b0), .Q(c[82]) );
  DFF \rc_reg[81]  ( .D(n1618), .CLK(clk), .RST(1'b0), .Q(c[81]) );
  DFF \rc_reg[80]  ( .D(n1617), .CLK(clk), .RST(1'b0), .Q(c[80]) );
  DFF \rc_reg[79]  ( .D(n1616), .CLK(clk), .RST(1'b0), .Q(c[79]) );
  DFF \rc_reg[78]  ( .D(n1615), .CLK(clk), .RST(1'b0), .Q(c[78]) );
  DFF \rc_reg[77]  ( .D(n1614), .CLK(clk), .RST(1'b0), .Q(c[77]) );
  DFF \rc_reg[76]  ( .D(n1613), .CLK(clk), .RST(1'b0), .Q(c[76]) );
  DFF \rc_reg[75]  ( .D(n1612), .CLK(clk), .RST(1'b0), .Q(c[75]) );
  DFF \rc_reg[74]  ( .D(n1611), .CLK(clk), .RST(1'b0), .Q(c[74]) );
  DFF \rc_reg[73]  ( .D(n1610), .CLK(clk), .RST(1'b0), .Q(c[73]) );
  DFF \rc_reg[72]  ( .D(n1609), .CLK(clk), .RST(1'b0), .Q(c[72]) );
  DFF \rc_reg[71]  ( .D(n1608), .CLK(clk), .RST(1'b0), .Q(c[71]) );
  DFF \rc_reg[70]  ( .D(n1607), .CLK(clk), .RST(1'b0), .Q(c[70]) );
  DFF \rc_reg[69]  ( .D(n1606), .CLK(clk), .RST(1'b0), .Q(c[69]) );
  DFF \rc_reg[68]  ( .D(n1605), .CLK(clk), .RST(1'b0), .Q(c[68]) );
  DFF \rc_reg[67]  ( .D(n1604), .CLK(clk), .RST(1'b0), .Q(c[67]) );
  DFF \rc_reg[66]  ( .D(n1603), .CLK(clk), .RST(1'b0), .Q(c[66]) );
  DFF \rc_reg[65]  ( .D(n1602), .CLK(clk), .RST(1'b0), .Q(c[65]) );
  DFF \rc_reg[64]  ( .D(n1601), .CLK(clk), .RST(1'b0), .Q(c[64]) );
  DFF \rc_reg[63]  ( .D(n1600), .CLK(clk), .RST(1'b0), .Q(c[63]) );
  DFF \rc_reg[62]  ( .D(n1599), .CLK(clk), .RST(1'b0), .Q(c[62]) );
  DFF \rc_reg[61]  ( .D(n1598), .CLK(clk), .RST(1'b0), .Q(c[61]) );
  DFF \rc_reg[60]  ( .D(n1597), .CLK(clk), .RST(1'b0), .Q(c[60]) );
  DFF \rc_reg[59]  ( .D(n1596), .CLK(clk), .RST(1'b0), .Q(c[59]) );
  DFF \rc_reg[58]  ( .D(n1595), .CLK(clk), .RST(1'b0), .Q(c[58]) );
  DFF \rc_reg[57]  ( .D(n1594), .CLK(clk), .RST(1'b0), .Q(c[57]) );
  DFF \rc_reg[56]  ( .D(n1593), .CLK(clk), .RST(1'b0), .Q(c[56]) );
  DFF \rc_reg[55]  ( .D(n1592), .CLK(clk), .RST(1'b0), .Q(c[55]) );
  DFF \rc_reg[54]  ( .D(n1591), .CLK(clk), .RST(1'b0), .Q(c[54]) );
  DFF \rc_reg[53]  ( .D(n1590), .CLK(clk), .RST(1'b0), .Q(c[53]) );
  DFF \rc_reg[52]  ( .D(n1589), .CLK(clk), .RST(1'b0), .Q(c[52]) );
  DFF \rc_reg[51]  ( .D(n1588), .CLK(clk), .RST(1'b0), .Q(c[51]) );
  DFF \rc_reg[50]  ( .D(n1587), .CLK(clk), .RST(1'b0), .Q(c[50]) );
  DFF \rc_reg[49]  ( .D(n1586), .CLK(clk), .RST(1'b0), .Q(c[49]) );
  DFF \rc_reg[48]  ( .D(n1585), .CLK(clk), .RST(1'b0), .Q(c[48]) );
  DFF \rc_reg[47]  ( .D(n1584), .CLK(clk), .RST(1'b0), .Q(c[47]) );
  DFF \rc_reg[46]  ( .D(n1583), .CLK(clk), .RST(1'b0), .Q(c[46]) );
  DFF \rc_reg[45]  ( .D(n1582), .CLK(clk), .RST(1'b0), .Q(c[45]) );
  DFF \rc_reg[44]  ( .D(n1581), .CLK(clk), .RST(1'b0), .Q(c[44]) );
  DFF \rc_reg[43]  ( .D(n1580), .CLK(clk), .RST(1'b0), .Q(c[43]) );
  DFF \rc_reg[42]  ( .D(n1579), .CLK(clk), .RST(1'b0), .Q(c[42]) );
  DFF \rc_reg[41]  ( .D(n1578), .CLK(clk), .RST(1'b0), .Q(c[41]) );
  DFF \rc_reg[40]  ( .D(n1577), .CLK(clk), .RST(1'b0), .Q(c[40]) );
  DFF \rc_reg[39]  ( .D(n1576), .CLK(clk), .RST(1'b0), .Q(c[39]) );
  DFF \rc_reg[38]  ( .D(n1575), .CLK(clk), .RST(1'b0), .Q(c[38]) );
  DFF \rc_reg[37]  ( .D(n1574), .CLK(clk), .RST(1'b0), .Q(c[37]) );
  DFF \rc_reg[36]  ( .D(n1573), .CLK(clk), .RST(1'b0), .Q(c[36]) );
  DFF \rc_reg[35]  ( .D(n1572), .CLK(clk), .RST(1'b0), .Q(c[35]) );
  DFF \rc_reg[34]  ( .D(n1571), .CLK(clk), .RST(1'b0), .Q(c[34]) );
  DFF \rc_reg[33]  ( .D(n1570), .CLK(clk), .RST(1'b0), .Q(c[33]) );
  DFF \rc_reg[32]  ( .D(n1569), .CLK(clk), .RST(1'b0), .Q(c[32]) );
  DFF \rc_reg[31]  ( .D(n1568), .CLK(clk), .RST(1'b0), .Q(c[31]) );
  DFF \rc_reg[30]  ( .D(n1567), .CLK(clk), .RST(1'b0), .Q(c[30]) );
  DFF \rc_reg[29]  ( .D(n1566), .CLK(clk), .RST(1'b0), .Q(c[29]) );
  DFF \rc_reg[28]  ( .D(n1565), .CLK(clk), .RST(1'b0), .Q(c[28]) );
  DFF \rc_reg[27]  ( .D(n1564), .CLK(clk), .RST(1'b0), .Q(c[27]) );
  DFF \rc_reg[26]  ( .D(n1563), .CLK(clk), .RST(1'b0), .Q(c[26]) );
  DFF \rc_reg[25]  ( .D(n1562), .CLK(clk), .RST(1'b0), .Q(c[25]) );
  DFF \rc_reg[24]  ( .D(n1561), .CLK(clk), .RST(1'b0), .Q(c[24]) );
  DFF \rc_reg[23]  ( .D(n1560), .CLK(clk), .RST(1'b0), .Q(c[23]) );
  DFF \rc_reg[22]  ( .D(n1559), .CLK(clk), .RST(1'b0), .Q(c[22]) );
  DFF \rc_reg[21]  ( .D(n1558), .CLK(clk), .RST(1'b0), .Q(c[21]) );
  DFF \rc_reg[20]  ( .D(n1557), .CLK(clk), .RST(1'b0), .Q(c[20]) );
  DFF \rc_reg[19]  ( .D(n1556), .CLK(clk), .RST(1'b0), .Q(c[19]) );
  DFF \rc_reg[18]  ( .D(n1555), .CLK(clk), .RST(1'b0), .Q(c[18]) );
  DFF \rc_reg[17]  ( .D(n1554), .CLK(clk), .RST(1'b0), .Q(c[17]) );
  DFF \rc_reg[16]  ( .D(n1553), .CLK(clk), .RST(1'b0), .Q(c[16]) );
  DFF \rc_reg[15]  ( .D(n1552), .CLK(clk), .RST(1'b0), .Q(c[15]) );
  DFF \rc_reg[14]  ( .D(n1551), .CLK(clk), .RST(1'b0), .Q(c[14]) );
  DFF \rc_reg[13]  ( .D(n1550), .CLK(clk), .RST(1'b0), .Q(c[13]) );
  DFF \rc_reg[12]  ( .D(n1549), .CLK(clk), .RST(1'b0), .Q(c[12]) );
  DFF \rc_reg[11]  ( .D(n1548), .CLK(clk), .RST(1'b0), .Q(c[11]) );
  DFF \rc_reg[10]  ( .D(n1547), .CLK(clk), .RST(1'b0), .Q(c[10]) );
  DFF \rc_reg[9]  ( .D(n1546), .CLK(clk), .RST(1'b0), .Q(c[9]) );
  DFF \rc_reg[8]  ( .D(n1545), .CLK(clk), .RST(1'b0), .Q(c[8]) );
  DFF \rc_reg[7]  ( .D(n1544), .CLK(clk), .RST(1'b0), .Q(c[7]) );
  DFF \rc_reg[6]  ( .D(n1543), .CLK(clk), .RST(1'b0), .Q(c[6]) );
  DFF \rc_reg[5]  ( .D(n1542), .CLK(clk), .RST(1'b0), .Q(c[5]) );
  DFF \rc_reg[4]  ( .D(n1541), .CLK(clk), .RST(1'b0), .Q(c[4]) );
  DFF \rc_reg[3]  ( .D(n1540), .CLK(clk), .RST(1'b0), .Q(c[3]) );
  DFF \rc_reg[2]  ( .D(n1539), .CLK(clk), .RST(1'b0), .Q(c[2]) );
  DFF \rc_reg[1]  ( .D(n1538), .CLK(clk), .RST(1'b0), .Q(c[1]) );
  DFF \rc_reg[0]  ( .D(n1537), .CLK(clk), .RST(1'b0), .Q(c[0]) );
  NAND U2051 ( .A(n5874), .B(n5873), .Z(n2049) );
  NANDN U2052 ( .A(n3036), .B(n3037), .Z(n2050) );
  NANDN U2053 ( .A(n5869), .B(n5868), .Z(n2051) );
  AND U2054 ( .A(n2050), .B(n2051), .Z(n2052) );
  NANDN U2055 ( .A(n2052), .B(n3038), .Z(n2053) );
  AND U2056 ( .A(n2049), .B(n2053), .Z(n3039) );
  NAND U2057 ( .A(n6514), .B(n6513), .Z(n2054) );
  NANDN U2058 ( .A(n3778), .B(n3779), .Z(n2055) );
  NANDN U2059 ( .A(n6509), .B(n6508), .Z(n2056) );
  AND U2060 ( .A(n2055), .B(n2056), .Z(n2057) );
  NANDN U2061 ( .A(n2057), .B(n3780), .Z(n2058) );
  AND U2062 ( .A(n2054), .B(n2058), .Z(n3781) );
  NANDN U2063 ( .A(n4520), .B(n4521), .Z(n2059) );
  NANDN U2064 ( .A(n7149), .B(n7148), .Z(n2060) );
  AND U2065 ( .A(n2059), .B(n2060), .Z(n2061) );
  NAND U2066 ( .A(n7154), .B(n7153), .Z(n2062) );
  NANDN U2067 ( .A(n2061), .B(n4522), .Z(n2063) );
  AND U2068 ( .A(n2062), .B(n2063), .Z(n4523) );
  XOR U2069 ( .A(n2131), .B(n2130), .Z(n5098) );
  XOR U2070 ( .A(n2155), .B(n2154), .Z(n5118) );
  XOR U2071 ( .A(n2179), .B(n2178), .Z(n5138) );
  XOR U2072 ( .A(n2219), .B(n2218), .Z(n5173) );
  XOR U2073 ( .A(n2259), .B(n2258), .Z(n5208) );
  XOR U2074 ( .A(n2283), .B(n2282), .Z(n5228) );
  XOR U2075 ( .A(n2307), .B(n2306), .Z(n5248) );
  XOR U2076 ( .A(n2331), .B(n2330), .Z(n5268) );
  XOR U2077 ( .A(n2355), .B(n2354), .Z(n5288) );
  XOR U2078 ( .A(n2379), .B(n2378), .Z(n5308) );
  XOR U2079 ( .A(n2403), .B(n2402), .Z(n5328) );
  XOR U2080 ( .A(n2427), .B(n2426), .Z(n5348) );
  XOR U2081 ( .A(n2451), .B(n2450), .Z(n5368) );
  XOR U2082 ( .A(n2475), .B(n2474), .Z(n5388) );
  XOR U2083 ( .A(n2499), .B(n2498), .Z(n5408) );
  XOR U2084 ( .A(n2523), .B(n2522), .Z(n5428) );
  XOR U2085 ( .A(n2547), .B(n2546), .Z(n5448) );
  XOR U2086 ( .A(n2643), .B(n2642), .Z(n5533) );
  XOR U2087 ( .A(n2667), .B(n2666), .Z(n5553) );
  XOR U2088 ( .A(n2691), .B(n2690), .Z(n5573) );
  XOR U2089 ( .A(n2715), .B(n2714), .Z(n5593) );
  XOR U2090 ( .A(n2739), .B(n2738), .Z(n5613) );
  XOR U2091 ( .A(n2763), .B(n2762), .Z(n5633) );
  XOR U2092 ( .A(n2787), .B(n2786), .Z(n5653) );
  XOR U2093 ( .A(n2827), .B(n2826), .Z(n5688) );
  XOR U2094 ( .A(n2851), .B(n2850), .Z(n5708) );
  XOR U2095 ( .A(n2875), .B(n2874), .Z(n5728) );
  XOR U2096 ( .A(n2899), .B(n2898), .Z(n5748) );
  XOR U2097 ( .A(n2923), .B(n2922), .Z(n5768) );
  XOR U2098 ( .A(n2947), .B(n2946), .Z(n5788) );
  XOR U2099 ( .A(n3015), .B(n3014), .Z(n5848) );
  XOR U2100 ( .A(n3058), .B(n3057), .Z(n5893) );
  XOR U2101 ( .A(n3082), .B(n3081), .Z(n5913) );
  XOR U2102 ( .A(n3106), .B(n3105), .Z(n5933) );
  XOR U2103 ( .A(n3130), .B(n3129), .Z(n5953) );
  OR U2104 ( .A(n3159), .B(n3160), .Z(n2064) );
  ANDN U2105 ( .B(n2064), .A(n3162), .Z(n5984) );
  XOR U2106 ( .A(n3197), .B(n3196), .Z(n6013) );
  XOR U2107 ( .A(n3221), .B(n3220), .Z(n6033) );
  XOR U2108 ( .A(n3273), .B(n3272), .Z(n6078) );
  XOR U2109 ( .A(n3297), .B(n3296), .Z(n6098) );
  XOR U2110 ( .A(n3321), .B(n3320), .Z(n6118) );
  XOR U2111 ( .A(n3361), .B(n3360), .Z(n6153) );
  XOR U2112 ( .A(n3385), .B(n3384), .Z(n6173) );
  XOR U2113 ( .A(n3409), .B(n3408), .Z(n6193) );
  XOR U2114 ( .A(n3433), .B(n3432), .Z(n6213) );
  XOR U2115 ( .A(n3473), .B(n3472), .Z(n6248) );
  XOR U2116 ( .A(n3497), .B(n3496), .Z(n6268) );
  XOR U2117 ( .A(n3521), .B(n3520), .Z(n6288) );
  XOR U2118 ( .A(n3545), .B(n3544), .Z(n6308) );
  XOR U2119 ( .A(n3569), .B(n3568), .Z(n6328) );
  XOR U2120 ( .A(n3593), .B(n3592), .Z(n6348) );
  XOR U2121 ( .A(n3617), .B(n3616), .Z(n6368) );
  XOR U2122 ( .A(n3641), .B(n3640), .Z(n6388) );
  XOR U2123 ( .A(n3665), .B(n3664), .Z(n6408) );
  XOR U2124 ( .A(n3689), .B(n3688), .Z(n6428) );
  XOR U2125 ( .A(n3757), .B(n3756), .Z(n6488) );
  XOR U2126 ( .A(n3800), .B(n3799), .Z(n6533) );
  XOR U2127 ( .A(n3824), .B(n3823), .Z(n6553) );
  XOR U2128 ( .A(n3848), .B(n3847), .Z(n6573) );
  XOR U2129 ( .A(n3872), .B(n3871), .Z(n6593) );
  OR U2130 ( .A(n3901), .B(n3902), .Z(n2065) );
  ANDN U2131 ( .B(n2065), .A(n3904), .Z(n6624) );
  XOR U2132 ( .A(n3939), .B(n3938), .Z(n6653) );
  XOR U2133 ( .A(n3963), .B(n3962), .Z(n6673) );
  XOR U2134 ( .A(n4015), .B(n4014), .Z(n6718) );
  XOR U2135 ( .A(n4039), .B(n4038), .Z(n6738) );
  XOR U2136 ( .A(n4063), .B(n4062), .Z(n6758) );
  XOR U2137 ( .A(n4103), .B(n4102), .Z(n6793) );
  XOR U2138 ( .A(n4127), .B(n4126), .Z(n6813) );
  XOR U2139 ( .A(n4151), .B(n4150), .Z(n6833) );
  XOR U2140 ( .A(n4175), .B(n4174), .Z(n6853) );
  XOR U2141 ( .A(n4215), .B(n4214), .Z(n6888) );
  XOR U2142 ( .A(n4239), .B(n4238), .Z(n6908) );
  XOR U2143 ( .A(n4263), .B(n4262), .Z(n6928) );
  XOR U2144 ( .A(n4287), .B(n4286), .Z(n6948) );
  XOR U2145 ( .A(n4311), .B(n4310), .Z(n6968) );
  XOR U2146 ( .A(n4335), .B(n4334), .Z(n6988) );
  XOR U2147 ( .A(n4359), .B(n4358), .Z(n7008) );
  XOR U2148 ( .A(n4383), .B(n4382), .Z(n7028) );
  XOR U2149 ( .A(n4407), .B(n4406), .Z(n7048) );
  XOR U2150 ( .A(n4431), .B(n4430), .Z(n7068) );
  XOR U2151 ( .A(n4499), .B(n4498), .Z(n7128) );
  XOR U2152 ( .A(n4542), .B(n4541), .Z(n7173) );
  XOR U2153 ( .A(n4566), .B(n4565), .Z(n7193) );
  XOR U2154 ( .A(n4590), .B(n4589), .Z(n7213) );
  XOR U2155 ( .A(n4614), .B(n4613), .Z(n7233) );
  OR U2156 ( .A(n4643), .B(n4644), .Z(n2066) );
  ANDN U2157 ( .B(n2066), .A(n4646), .Z(n7264) );
  XOR U2158 ( .A(n4681), .B(n4680), .Z(n7293) );
  XOR U2159 ( .A(n4705), .B(n4704), .Z(n7313) );
  XOR U2160 ( .A(n4757), .B(n4756), .Z(n7358) );
  XOR U2161 ( .A(n4781), .B(n4780), .Z(n7378) );
  XOR U2162 ( .A(n4805), .B(n4804), .Z(n7398) );
  XOR U2163 ( .A(n4845), .B(n4844), .Z(n7433) );
  XOR U2164 ( .A(n4869), .B(n4868), .Z(n7453) );
  XOR U2165 ( .A(n4893), .B(n4892), .Z(n7473) );
  XOR U2166 ( .A(n4917), .B(n4916), .Z(n7493) );
  XOR U2167 ( .A(n4957), .B(n4956), .Z(n7528) );
  XOR U2168 ( .A(n4981), .B(n4980), .Z(n7548) );
  XOR U2169 ( .A(n5005), .B(n5004), .Z(n7568) );
  XOR U2170 ( .A(n5029), .B(n5028), .Z(n7588) );
  NAND U2171 ( .A(n5879), .B(n5878), .Z(n2067) );
  NAND U2172 ( .A(n3041), .B(n3040), .Z(n2068) );
  NAND U2173 ( .A(n2067), .B(n2068), .Z(n2069) );
  ANDN U2174 ( .B(n2069), .A(n3043), .Z(n3045) );
  NAND U2175 ( .A(n6519), .B(n6518), .Z(n2070) );
  NAND U2176 ( .A(n3783), .B(n3782), .Z(n2071) );
  NAND U2177 ( .A(n2070), .B(n2071), .Z(n2072) );
  ANDN U2178 ( .B(n2072), .A(n3785), .Z(n3787) );
  NAND U2179 ( .A(n7159), .B(n7158), .Z(n2073) );
  NAND U2180 ( .A(n4525), .B(n4524), .Z(n2074) );
  NAND U2181 ( .A(n2073), .B(n2074), .Z(n2075) );
  ANDN U2182 ( .B(n2075), .A(n4527), .Z(n4529) );
  XOR U2183 ( .A(n2101), .B(n2102), .Z(n5074) );
  XOR U2184 ( .A(n2119), .B(n2118), .Z(n5088) );
  XOR U2185 ( .A(n2143), .B(n2142), .Z(n5108) );
  XOR U2186 ( .A(n2167), .B(n2166), .Z(n5128) );
  XOR U2187 ( .A(n2191), .B(n2190), .Z(n5148) );
  XOR U2188 ( .A(n2231), .B(n2230), .Z(n5183) );
  XOR U2189 ( .A(n2271), .B(n2270), .Z(n5218) );
  XOR U2190 ( .A(n2295), .B(n2294), .Z(n5238) );
  XOR U2191 ( .A(n2319), .B(n2318), .Z(n5258) );
  XOR U2192 ( .A(n2343), .B(n2342), .Z(n5278) );
  XOR U2193 ( .A(n2367), .B(n2366), .Z(n5298) );
  XOR U2194 ( .A(n2391), .B(n2390), .Z(n5318) );
  XOR U2195 ( .A(n2415), .B(n2414), .Z(n5338) );
  XOR U2196 ( .A(n2439), .B(n2438), .Z(n5358) );
  XOR U2197 ( .A(n2463), .B(n2462), .Z(n5378) );
  XOR U2198 ( .A(n2487), .B(n2486), .Z(n5398) );
  XOR U2199 ( .A(n2511), .B(n2510), .Z(n5418) );
  XOR U2200 ( .A(n2535), .B(n2534), .Z(n5438) );
  XOR U2201 ( .A(n2559), .B(n2558), .Z(n5458) );
  XOR U2202 ( .A(n2587), .B(n2586), .Z(n5483) );
  XOR U2203 ( .A(n2615), .B(n2614), .Z(n5508) );
  XOR U2204 ( .A(n2655), .B(n2654), .Z(n5543) );
  XOR U2205 ( .A(n2679), .B(n2678), .Z(n5563) );
  XOR U2206 ( .A(n2703), .B(n2702), .Z(n5583) );
  XOR U2207 ( .A(n2727), .B(n2726), .Z(n5603) );
  XOR U2208 ( .A(n2751), .B(n2750), .Z(n5623) );
  XOR U2209 ( .A(n2775), .B(n2774), .Z(n5643) );
  XOR U2210 ( .A(n2799), .B(n2798), .Z(n5663) );
  XOR U2211 ( .A(n2839), .B(n2838), .Z(n5698) );
  XOR U2212 ( .A(n2863), .B(n2862), .Z(n5718) );
  XOR U2213 ( .A(n2887), .B(n2886), .Z(n5738) );
  XOR U2214 ( .A(n2911), .B(n2910), .Z(n5758) );
  XOR U2215 ( .A(n2935), .B(n2934), .Z(n5778) );
  XOR U2216 ( .A(n2959), .B(n2958), .Z(n5798) );
  XOR U2217 ( .A(n2987), .B(n2986), .Z(n5823) );
  XOR U2218 ( .A(n3027), .B(n3026), .Z(n5858) );
  XOR U2219 ( .A(n3070), .B(n3069), .Z(n5903) );
  XOR U2220 ( .A(n3094), .B(n3093), .Z(n5923) );
  XOR U2221 ( .A(n3118), .B(n3117), .Z(n5943) );
  XOR U2222 ( .A(n3142), .B(n3141), .Z(n5963) );
  XOR U2223 ( .A(n3169), .B(n3168), .Z(n5988) );
  XOR U2224 ( .A(n3209), .B(n3208), .Z(n6023) );
  XOR U2225 ( .A(n3233), .B(n3232), .Z(n6043) );
  XOR U2226 ( .A(n3261), .B(n3260), .Z(n6068) );
  XOR U2227 ( .A(n3285), .B(n3284), .Z(n6088) );
  XOR U2228 ( .A(n3309), .B(n3308), .Z(n6108) );
  XOR U2229 ( .A(n3333), .B(n3332), .Z(n6128) );
  XOR U2230 ( .A(n3373), .B(n3372), .Z(n6163) );
  XOR U2231 ( .A(n3397), .B(n3396), .Z(n6183) );
  XOR U2232 ( .A(n3421), .B(n3420), .Z(n6203) );
  XOR U2233 ( .A(n3445), .B(n3444), .Z(n6223) );
  XOR U2234 ( .A(n3485), .B(n3484), .Z(n6258) );
  XOR U2235 ( .A(n3509), .B(n3508), .Z(n6278) );
  XOR U2236 ( .A(n3533), .B(n3532), .Z(n6298) );
  XOR U2237 ( .A(n3557), .B(n3556), .Z(n6318) );
  XOR U2238 ( .A(n3581), .B(n3580), .Z(n6338) );
  XOR U2239 ( .A(n3605), .B(n3604), .Z(n6358) );
  XOR U2240 ( .A(n3629), .B(n3628), .Z(n6378) );
  XOR U2241 ( .A(n3653), .B(n3652), .Z(n6398) );
  XOR U2242 ( .A(n3677), .B(n3676), .Z(n6418) );
  XOR U2243 ( .A(n3701), .B(n3700), .Z(n6438) );
  XOR U2244 ( .A(n3729), .B(n3728), .Z(n6463) );
  XOR U2245 ( .A(n3769), .B(n3768), .Z(n6498) );
  XOR U2246 ( .A(n3812), .B(n3811), .Z(n6543) );
  XOR U2247 ( .A(n3836), .B(n3835), .Z(n6563) );
  XOR U2248 ( .A(n3860), .B(n3859), .Z(n6583) );
  XOR U2249 ( .A(n3884), .B(n3883), .Z(n6603) );
  XOR U2250 ( .A(n3911), .B(n3910), .Z(n6628) );
  XOR U2251 ( .A(n3951), .B(n3950), .Z(n6663) );
  XOR U2252 ( .A(n3975), .B(n3974), .Z(n6683) );
  XOR U2253 ( .A(n4003), .B(n4002), .Z(n6708) );
  XOR U2254 ( .A(n4027), .B(n4026), .Z(n6728) );
  XOR U2255 ( .A(n4051), .B(n4050), .Z(n6748) );
  XOR U2256 ( .A(n4075), .B(n4074), .Z(n6768) );
  XOR U2257 ( .A(n4115), .B(n4114), .Z(n6803) );
  XOR U2258 ( .A(n4139), .B(n4138), .Z(n6823) );
  XOR U2259 ( .A(n4163), .B(n4162), .Z(n6843) );
  XOR U2260 ( .A(n4187), .B(n4186), .Z(n6863) );
  XOR U2261 ( .A(n4227), .B(n4226), .Z(n6898) );
  XOR U2262 ( .A(n4251), .B(n4250), .Z(n6918) );
  XOR U2263 ( .A(n4275), .B(n4274), .Z(n6938) );
  XOR U2264 ( .A(n4299), .B(n4298), .Z(n6958) );
  XOR U2265 ( .A(n4323), .B(n4322), .Z(n6978) );
  XOR U2266 ( .A(n4347), .B(n4346), .Z(n6998) );
  XOR U2267 ( .A(n4371), .B(n4370), .Z(n7018) );
  XOR U2268 ( .A(n4395), .B(n4394), .Z(n7038) );
  XOR U2269 ( .A(n4419), .B(n4418), .Z(n7058) );
  XOR U2270 ( .A(n4443), .B(n4442), .Z(n7078) );
  XOR U2271 ( .A(n4471), .B(n4470), .Z(n7103) );
  XOR U2272 ( .A(n4511), .B(n4510), .Z(n7138) );
  XOR U2273 ( .A(n4554), .B(n4553), .Z(n7183) );
  XOR U2274 ( .A(n4578), .B(n4577), .Z(n7203) );
  XOR U2275 ( .A(n4602), .B(n4601), .Z(n7223) );
  XOR U2276 ( .A(n4626), .B(n4625), .Z(n7243) );
  XOR U2277 ( .A(n4653), .B(n4652), .Z(n7268) );
  XOR U2278 ( .A(n4693), .B(n4692), .Z(n7303) );
  XOR U2279 ( .A(n4717), .B(n4716), .Z(n7323) );
  XOR U2280 ( .A(n4745), .B(n4744), .Z(n7348) );
  XOR U2281 ( .A(n4769), .B(n4768), .Z(n7368) );
  XOR U2282 ( .A(n4793), .B(n4792), .Z(n7388) );
  XOR U2283 ( .A(n4817), .B(n4816), .Z(n7408) );
  XOR U2284 ( .A(n4857), .B(n4856), .Z(n7443) );
  XOR U2285 ( .A(n4881), .B(n4880), .Z(n7463) );
  XOR U2286 ( .A(n4905), .B(n4904), .Z(n7483) );
  XOR U2287 ( .A(n4929), .B(n4928), .Z(n7503) );
  XOR U2288 ( .A(n4969), .B(n4968), .Z(n7538) );
  XOR U2289 ( .A(n4993), .B(n4992), .Z(n7558) );
  XOR U2290 ( .A(n5017), .B(n5016), .Z(n7578) );
  XOR U2291 ( .A(n5039), .B(n5040), .Z(n7598) );
  AND U2292 ( .A(a[511]), .B(b[511]), .Z(n5048) );
  NAND U2293 ( .A(a[510]), .B(b[510]), .Z(n5044) );
  NAND U2294 ( .A(a[509]), .B(b[509]), .Z(n5039) );
  NAND U2295 ( .A(a[442]), .B(b[442]), .Z(n4643) );
  NAND U2296 ( .A(a[423]), .B(b[423]), .Z(n4531) );
  NAND U2297 ( .A(a[421]), .B(b[421]), .Z(n4524) );
  NAND U2298 ( .A(a[420]), .B(b[420]), .Z(n4522) );
  AND U2299 ( .A(a[419]), .B(b[419]), .Z(n4520) );
  NAND U2300 ( .A(a[409]), .B(b[409]), .Z(n4460) );
  NAND U2301 ( .A(a[314]), .B(b[314]), .Z(n3901) );
  NAND U2302 ( .A(a[295]), .B(b[295]), .Z(n3789) );
  NAND U2303 ( .A(a[293]), .B(b[293]), .Z(n3782) );
  NAND U2304 ( .A(a[292]), .B(b[292]), .Z(n3780) );
  AND U2305 ( .A(a[291]), .B(b[291]), .Z(n3778) );
  NAND U2306 ( .A(a[281]), .B(b[281]), .Z(n3718) );
  NAND U2307 ( .A(a[186]), .B(b[186]), .Z(n3159) );
  NAND U2308 ( .A(a[167]), .B(b[167]), .Z(n3047) );
  NAND U2309 ( .A(a[165]), .B(b[165]), .Z(n3040) );
  NAND U2310 ( .A(a[164]), .B(b[164]), .Z(n3038) );
  AND U2311 ( .A(a[163]), .B(b[163]), .Z(n3036) );
  NAND U2312 ( .A(a[153]), .B(b[153]), .Z(n2976) );
  NAND U2313 ( .A(a[126]), .B(b[126]), .Z(n2816) );
  NAND U2314 ( .A(a[85]), .B(b[85]), .Z(n2576) );
  NAND U2315 ( .A(a[23]), .B(b[23]), .Z(n2208) );
  AND U2316 ( .A(a[4]), .B(b[4]), .Z(n2101) );
  AND U2317 ( .A(a[3]), .B(b[3]), .Z(n2094) );
  AND U2318 ( .A(a[2]), .B(b[2]), .Z(n2090) );
  XNOR U2319 ( .A(a[1]), .B(b[1]), .Z(n2078) );
  XNOR U2320 ( .A(carry_on[1]), .B(n2078), .Z(n5054) );
  NAND U2321 ( .A(a[0]), .B(b[0]), .Z(n2077) );
  XOR U2322 ( .A(a[0]), .B(b[0]), .Z(n5049) );
  NAND U2323 ( .A(n5049), .B(carry_on[0]), .Z(n2076) );
  NAND U2324 ( .A(n2077), .B(n2076), .Z(n5053) );
  NAND U2325 ( .A(n5054), .B(n5053), .Z(n2080) );
  ANDN U2326 ( .B(carry_on[1]), .A(n2078), .Z(n2081) );
  ANDN U2327 ( .B(n2080), .A(n2081), .Z(n2079) );
  NAND U2328 ( .A(a[1]), .B(b[1]), .Z(n2082) );
  NAND U2329 ( .A(n2079), .B(n2082), .Z(n2086) );
  XNOR U2330 ( .A(n2082), .B(n2080), .Z(n2084) );
  NAND U2331 ( .A(n2082), .B(n2081), .Z(n2083) );
  NAND U2332 ( .A(n2084), .B(n2083), .Z(n5059) );
  XNOR U2333 ( .A(a[2]), .B(b[2]), .Z(n5058) );
  NAND U2334 ( .A(n5059), .B(n5058), .Z(n2085) );
  NAND U2335 ( .A(n2086), .B(n2085), .Z(n2091) );
  ANDN U2336 ( .B(n2090), .A(n2091), .Z(n2087) );
  XNOR U2337 ( .A(n2094), .B(n2087), .Z(n2089) );
  XNOR U2338 ( .A(n2090), .B(n2091), .Z(n5063) );
  XOR U2339 ( .A(a[3]), .B(b[3]), .Z(n5064) );
  NAND U2340 ( .A(n5063), .B(n5064), .Z(n2088) );
  NAND U2341 ( .A(n2089), .B(n2088), .Z(n5069) );
  XNOR U2342 ( .A(a[4]), .B(b[4]), .Z(n5068) );
  NAND U2343 ( .A(n5069), .B(n5068), .Z(n2097) );
  ANDN U2344 ( .B(n2091), .A(n2090), .Z(n2093) );
  ANDN U2345 ( .B(n5063), .A(n5064), .Z(n2092) );
  OR U2346 ( .A(n2093), .B(n2092), .Z(n2095) );
  ANDN U2347 ( .B(n2095), .A(n2094), .Z(n2096) );
  ANDN U2348 ( .B(n2097), .A(n2096), .Z(n2102) );
  NOR U2349 ( .A(n2101), .B(n2102), .Z(n2099) );
  XNOR U2350 ( .A(a[5]), .B(b[5]), .Z(n5073) );
  NAND U2351 ( .A(n5074), .B(n5073), .Z(n2098) );
  NANDN U2352 ( .A(n2099), .B(n2098), .Z(n2100) );
  AND U2353 ( .A(a[5]), .B(b[5]), .Z(n2104) );
  ANDN U2354 ( .B(n2100), .A(n2104), .Z(n2106) );
  AND U2355 ( .A(n2102), .B(n2101), .Z(n2103) );
  NAND U2356 ( .A(n2104), .B(n2103), .Z(n2109) );
  ANDN U2357 ( .B(n2109), .A(n2106), .Z(n5079) );
  XNOR U2358 ( .A(a[6]), .B(b[6]), .Z(n5078) );
  AND U2359 ( .A(n5079), .B(n5078), .Z(n2105) );
  OR U2360 ( .A(n2106), .B(n2105), .Z(n2107) );
  NAND U2361 ( .A(a[6]), .B(b[6]), .Z(n2108) );
  AND U2362 ( .A(n2107), .B(n2108), .Z(n2112) );
  OR U2363 ( .A(n2109), .B(n2108), .Z(n2110) );
  ANDN U2364 ( .B(n2110), .A(n2112), .Z(n5084) );
  XNOR U2365 ( .A(a[7]), .B(b[7]), .Z(n5083) );
  NAND U2366 ( .A(n5084), .B(n5083), .Z(n2111) );
  NANDN U2367 ( .A(n2112), .B(n2111), .Z(n2118) );
  NAND U2368 ( .A(a[7]), .B(b[7]), .Z(n2119) );
  AND U2369 ( .A(n2118), .B(n2119), .Z(n2114) );
  XOR U2370 ( .A(a[8]), .B(b[8]), .Z(n5089) );
  ANDN U2371 ( .B(n5088), .A(n5089), .Z(n2113) );
  OR U2372 ( .A(n2114), .B(n2113), .Z(n2115) );
  AND U2373 ( .A(a[8]), .B(b[8]), .Z(n2117) );
  ANDN U2374 ( .B(n2115), .A(n2117), .Z(n2124) );
  NOR U2375 ( .A(n2119), .B(n2118), .Z(n2116) );
  XNOR U2376 ( .A(n2117), .B(n2116), .Z(n2122) );
  XOR U2377 ( .A(n2119), .B(n2118), .Z(n2120) );
  NAND U2378 ( .A(n2120), .B(n5089), .Z(n2121) );
  NAND U2379 ( .A(n2122), .B(n2121), .Z(n5094) );
  XNOR U2380 ( .A(a[9]), .B(b[9]), .Z(n5093) );
  NAND U2381 ( .A(n5094), .B(n5093), .Z(n2123) );
  NANDN U2382 ( .A(n2124), .B(n2123), .Z(n2130) );
  NAND U2383 ( .A(a[9]), .B(b[9]), .Z(n2131) );
  AND U2384 ( .A(n2130), .B(n2131), .Z(n2126) );
  XOR U2385 ( .A(a[10]), .B(b[10]), .Z(n5099) );
  ANDN U2386 ( .B(n5098), .A(n5099), .Z(n2125) );
  OR U2387 ( .A(n2126), .B(n2125), .Z(n2127) );
  AND U2388 ( .A(a[10]), .B(b[10]), .Z(n2129) );
  ANDN U2389 ( .B(n2127), .A(n2129), .Z(n2136) );
  NOR U2390 ( .A(n2131), .B(n2130), .Z(n2128) );
  XNOR U2391 ( .A(n2129), .B(n2128), .Z(n2134) );
  XOR U2392 ( .A(n2131), .B(n2130), .Z(n2132) );
  NAND U2393 ( .A(n2132), .B(n5099), .Z(n2133) );
  NAND U2394 ( .A(n2134), .B(n2133), .Z(n5104) );
  XNOR U2395 ( .A(a[11]), .B(b[11]), .Z(n5103) );
  NAND U2396 ( .A(n5104), .B(n5103), .Z(n2135) );
  NANDN U2397 ( .A(n2136), .B(n2135), .Z(n2142) );
  NAND U2398 ( .A(a[11]), .B(b[11]), .Z(n2143) );
  AND U2399 ( .A(n2142), .B(n2143), .Z(n2138) );
  XOR U2400 ( .A(a[12]), .B(b[12]), .Z(n5109) );
  ANDN U2401 ( .B(n5108), .A(n5109), .Z(n2137) );
  OR U2402 ( .A(n2138), .B(n2137), .Z(n2139) );
  AND U2403 ( .A(a[12]), .B(b[12]), .Z(n2141) );
  ANDN U2404 ( .B(n2139), .A(n2141), .Z(n2148) );
  NOR U2405 ( .A(n2143), .B(n2142), .Z(n2140) );
  XNOR U2406 ( .A(n2141), .B(n2140), .Z(n2146) );
  XOR U2407 ( .A(n2143), .B(n2142), .Z(n2144) );
  NAND U2408 ( .A(n2144), .B(n5109), .Z(n2145) );
  NAND U2409 ( .A(n2146), .B(n2145), .Z(n5114) );
  XNOR U2410 ( .A(a[13]), .B(b[13]), .Z(n5113) );
  NAND U2411 ( .A(n5114), .B(n5113), .Z(n2147) );
  NANDN U2412 ( .A(n2148), .B(n2147), .Z(n2154) );
  NAND U2413 ( .A(a[13]), .B(b[13]), .Z(n2155) );
  AND U2414 ( .A(n2154), .B(n2155), .Z(n2150) );
  XOR U2415 ( .A(a[14]), .B(b[14]), .Z(n5119) );
  ANDN U2416 ( .B(n5118), .A(n5119), .Z(n2149) );
  OR U2417 ( .A(n2150), .B(n2149), .Z(n2151) );
  AND U2418 ( .A(a[14]), .B(b[14]), .Z(n2153) );
  ANDN U2419 ( .B(n2151), .A(n2153), .Z(n2160) );
  NOR U2420 ( .A(n2155), .B(n2154), .Z(n2152) );
  XNOR U2421 ( .A(n2153), .B(n2152), .Z(n2158) );
  XOR U2422 ( .A(n2155), .B(n2154), .Z(n2156) );
  NAND U2423 ( .A(n2156), .B(n5119), .Z(n2157) );
  NAND U2424 ( .A(n2158), .B(n2157), .Z(n5124) );
  XNOR U2425 ( .A(a[15]), .B(b[15]), .Z(n5123) );
  NAND U2426 ( .A(n5124), .B(n5123), .Z(n2159) );
  NANDN U2427 ( .A(n2160), .B(n2159), .Z(n2166) );
  NAND U2428 ( .A(a[15]), .B(b[15]), .Z(n2167) );
  AND U2429 ( .A(n2166), .B(n2167), .Z(n2162) );
  XOR U2430 ( .A(a[16]), .B(b[16]), .Z(n5129) );
  ANDN U2431 ( .B(n5128), .A(n5129), .Z(n2161) );
  OR U2432 ( .A(n2162), .B(n2161), .Z(n2163) );
  AND U2433 ( .A(a[16]), .B(b[16]), .Z(n2165) );
  ANDN U2434 ( .B(n2163), .A(n2165), .Z(n2172) );
  NOR U2435 ( .A(n2167), .B(n2166), .Z(n2164) );
  XNOR U2436 ( .A(n2165), .B(n2164), .Z(n2170) );
  XOR U2437 ( .A(n2167), .B(n2166), .Z(n2168) );
  NAND U2438 ( .A(n2168), .B(n5129), .Z(n2169) );
  NAND U2439 ( .A(n2170), .B(n2169), .Z(n5134) );
  XNOR U2440 ( .A(a[17]), .B(b[17]), .Z(n5133) );
  NAND U2441 ( .A(n5134), .B(n5133), .Z(n2171) );
  NANDN U2442 ( .A(n2172), .B(n2171), .Z(n2178) );
  NAND U2443 ( .A(a[17]), .B(b[17]), .Z(n2179) );
  AND U2444 ( .A(n2178), .B(n2179), .Z(n2174) );
  XOR U2445 ( .A(a[18]), .B(b[18]), .Z(n5139) );
  ANDN U2446 ( .B(n5138), .A(n5139), .Z(n2173) );
  OR U2447 ( .A(n2174), .B(n2173), .Z(n2175) );
  AND U2448 ( .A(a[18]), .B(b[18]), .Z(n2177) );
  ANDN U2449 ( .B(n2175), .A(n2177), .Z(n2184) );
  NOR U2450 ( .A(n2179), .B(n2178), .Z(n2176) );
  XNOR U2451 ( .A(n2177), .B(n2176), .Z(n2182) );
  XOR U2452 ( .A(n2179), .B(n2178), .Z(n2180) );
  NAND U2453 ( .A(n2180), .B(n5139), .Z(n2181) );
  NAND U2454 ( .A(n2182), .B(n2181), .Z(n5144) );
  XNOR U2455 ( .A(a[19]), .B(b[19]), .Z(n5143) );
  NAND U2456 ( .A(n5144), .B(n5143), .Z(n2183) );
  NANDN U2457 ( .A(n2184), .B(n2183), .Z(n2190) );
  NAND U2458 ( .A(a[19]), .B(b[19]), .Z(n2191) );
  AND U2459 ( .A(n2190), .B(n2191), .Z(n2186) );
  XOR U2460 ( .A(a[20]), .B(b[20]), .Z(n5149) );
  ANDN U2461 ( .B(n5148), .A(n5149), .Z(n2185) );
  OR U2462 ( .A(n2186), .B(n2185), .Z(n2187) );
  AND U2463 ( .A(a[20]), .B(b[20]), .Z(n2189) );
  ANDN U2464 ( .B(n2187), .A(n2189), .Z(n2196) );
  NOR U2465 ( .A(n2191), .B(n2190), .Z(n2188) );
  XNOR U2466 ( .A(n2189), .B(n2188), .Z(n2194) );
  XOR U2467 ( .A(n2191), .B(n2190), .Z(n2192) );
  NAND U2468 ( .A(n2192), .B(n5149), .Z(n2193) );
  NAND U2469 ( .A(n2194), .B(n2193), .Z(n5154) );
  XNOR U2470 ( .A(a[21]), .B(b[21]), .Z(n5153) );
  NAND U2471 ( .A(n5154), .B(n5153), .Z(n2195) );
  NANDN U2472 ( .A(n2196), .B(n2195), .Z(n2197) );
  IV U2473 ( .A(n2197), .Z(n2201) );
  AND U2474 ( .A(a[21]), .B(b[21]), .Z(n2202) );
  NOR U2475 ( .A(n2201), .B(n2202), .Z(n2199) );
  XNOR U2476 ( .A(n2202), .B(n2197), .Z(n5159) );
  XNOR U2477 ( .A(a[22]), .B(b[22]), .Z(n5158) );
  AND U2478 ( .A(n5159), .B(n5158), .Z(n2198) );
  OR U2479 ( .A(n2199), .B(n2198), .Z(n2200) );
  AND U2480 ( .A(a[22]), .B(b[22]), .Z(n2204) );
  ANDN U2481 ( .B(n2200), .A(n2204), .Z(n2206) );
  AND U2482 ( .A(n2202), .B(n2201), .Z(n2203) );
  NAND U2483 ( .A(n2204), .B(n2203), .Z(n2209) );
  ANDN U2484 ( .B(n2209), .A(n2206), .Z(n5164) );
  XNOR U2485 ( .A(a[23]), .B(b[23]), .Z(n5163) );
  AND U2486 ( .A(n5164), .B(n5163), .Z(n2205) );
  OR U2487 ( .A(n2206), .B(n2205), .Z(n2207) );
  AND U2488 ( .A(n2208), .B(n2207), .Z(n2212) );
  OR U2489 ( .A(n2209), .B(n2208), .Z(n2210) );
  ANDN U2490 ( .B(n2210), .A(n2212), .Z(n5169) );
  XNOR U2491 ( .A(a[24]), .B(b[24]), .Z(n5168) );
  NAND U2492 ( .A(n5169), .B(n5168), .Z(n2211) );
  NANDN U2493 ( .A(n2212), .B(n2211), .Z(n2218) );
  NAND U2494 ( .A(a[24]), .B(b[24]), .Z(n2219) );
  AND U2495 ( .A(n2218), .B(n2219), .Z(n2214) );
  XOR U2496 ( .A(a[25]), .B(b[25]), .Z(n5174) );
  ANDN U2497 ( .B(n5173), .A(n5174), .Z(n2213) );
  OR U2498 ( .A(n2214), .B(n2213), .Z(n2215) );
  AND U2499 ( .A(a[25]), .B(b[25]), .Z(n2217) );
  ANDN U2500 ( .B(n2215), .A(n2217), .Z(n2224) );
  NOR U2501 ( .A(n2219), .B(n2218), .Z(n2216) );
  XNOR U2502 ( .A(n2217), .B(n2216), .Z(n2222) );
  XOR U2503 ( .A(n2219), .B(n2218), .Z(n2220) );
  NAND U2504 ( .A(n2220), .B(n5174), .Z(n2221) );
  NAND U2505 ( .A(n2222), .B(n2221), .Z(n5179) );
  XNOR U2506 ( .A(a[26]), .B(b[26]), .Z(n5178) );
  NAND U2507 ( .A(n5179), .B(n5178), .Z(n2223) );
  NANDN U2508 ( .A(n2224), .B(n2223), .Z(n2230) );
  NAND U2509 ( .A(a[26]), .B(b[26]), .Z(n2231) );
  AND U2510 ( .A(n2230), .B(n2231), .Z(n2226) );
  XOR U2511 ( .A(a[27]), .B(b[27]), .Z(n5184) );
  ANDN U2512 ( .B(n5183), .A(n5184), .Z(n2225) );
  OR U2513 ( .A(n2226), .B(n2225), .Z(n2227) );
  AND U2514 ( .A(a[27]), .B(b[27]), .Z(n2229) );
  ANDN U2515 ( .B(n2227), .A(n2229), .Z(n2236) );
  NOR U2516 ( .A(n2231), .B(n2230), .Z(n2228) );
  XNOR U2517 ( .A(n2229), .B(n2228), .Z(n2234) );
  XOR U2518 ( .A(n2231), .B(n2230), .Z(n2232) );
  NAND U2519 ( .A(n2232), .B(n5184), .Z(n2233) );
  NAND U2520 ( .A(n2234), .B(n2233), .Z(n5189) );
  XNOR U2521 ( .A(a[28]), .B(b[28]), .Z(n5188) );
  NAND U2522 ( .A(n5189), .B(n5188), .Z(n2235) );
  NANDN U2523 ( .A(n2236), .B(n2235), .Z(n2237) );
  IV U2524 ( .A(n2237), .Z(n2241) );
  AND U2525 ( .A(a[28]), .B(b[28]), .Z(n2242) );
  NOR U2526 ( .A(n2241), .B(n2242), .Z(n2239) );
  XNOR U2527 ( .A(n2242), .B(n2237), .Z(n5194) );
  XNOR U2528 ( .A(a[29]), .B(b[29]), .Z(n5193) );
  AND U2529 ( .A(n5194), .B(n5193), .Z(n2238) );
  OR U2530 ( .A(n2239), .B(n2238), .Z(n2240) );
  AND U2531 ( .A(a[29]), .B(b[29]), .Z(n2244) );
  ANDN U2532 ( .B(n2240), .A(n2244), .Z(n2246) );
  AND U2533 ( .A(n2242), .B(n2241), .Z(n2243) );
  NAND U2534 ( .A(n2244), .B(n2243), .Z(n2249) );
  ANDN U2535 ( .B(n2249), .A(n2246), .Z(n5199) );
  XNOR U2536 ( .A(a[30]), .B(b[30]), .Z(n5198) );
  AND U2537 ( .A(n5199), .B(n5198), .Z(n2245) );
  OR U2538 ( .A(n2246), .B(n2245), .Z(n2247) );
  AND U2539 ( .A(a[30]), .B(b[30]), .Z(n2248) );
  ANDN U2540 ( .B(n2247), .A(n2248), .Z(n2252) );
  NANDN U2541 ( .A(n2249), .B(n2248), .Z(n2250) );
  ANDN U2542 ( .B(n2250), .A(n2252), .Z(n5204) );
  XNOR U2543 ( .A(a[31]), .B(b[31]), .Z(n5203) );
  NAND U2544 ( .A(n5204), .B(n5203), .Z(n2251) );
  NANDN U2545 ( .A(n2252), .B(n2251), .Z(n2258) );
  NAND U2546 ( .A(a[31]), .B(b[31]), .Z(n2259) );
  AND U2547 ( .A(n2258), .B(n2259), .Z(n2254) );
  XOR U2548 ( .A(a[32]), .B(b[32]), .Z(n5209) );
  ANDN U2549 ( .B(n5208), .A(n5209), .Z(n2253) );
  OR U2550 ( .A(n2254), .B(n2253), .Z(n2255) );
  AND U2551 ( .A(a[32]), .B(b[32]), .Z(n2257) );
  ANDN U2552 ( .B(n2255), .A(n2257), .Z(n2264) );
  NOR U2553 ( .A(n2259), .B(n2258), .Z(n2256) );
  XNOR U2554 ( .A(n2257), .B(n2256), .Z(n2262) );
  XOR U2555 ( .A(n2259), .B(n2258), .Z(n2260) );
  NAND U2556 ( .A(n2260), .B(n5209), .Z(n2261) );
  NAND U2557 ( .A(n2262), .B(n2261), .Z(n5214) );
  XNOR U2558 ( .A(a[33]), .B(b[33]), .Z(n5213) );
  NAND U2559 ( .A(n5214), .B(n5213), .Z(n2263) );
  NANDN U2560 ( .A(n2264), .B(n2263), .Z(n2270) );
  NAND U2561 ( .A(a[33]), .B(b[33]), .Z(n2271) );
  AND U2562 ( .A(n2270), .B(n2271), .Z(n2266) );
  XOR U2563 ( .A(a[34]), .B(b[34]), .Z(n5219) );
  ANDN U2564 ( .B(n5218), .A(n5219), .Z(n2265) );
  OR U2565 ( .A(n2266), .B(n2265), .Z(n2267) );
  AND U2566 ( .A(a[34]), .B(b[34]), .Z(n2269) );
  ANDN U2567 ( .B(n2267), .A(n2269), .Z(n2276) );
  NOR U2568 ( .A(n2271), .B(n2270), .Z(n2268) );
  XNOR U2569 ( .A(n2269), .B(n2268), .Z(n2274) );
  XOR U2570 ( .A(n2271), .B(n2270), .Z(n2272) );
  NAND U2571 ( .A(n2272), .B(n5219), .Z(n2273) );
  NAND U2572 ( .A(n2274), .B(n2273), .Z(n5224) );
  XNOR U2573 ( .A(a[35]), .B(b[35]), .Z(n5223) );
  NAND U2574 ( .A(n5224), .B(n5223), .Z(n2275) );
  NANDN U2575 ( .A(n2276), .B(n2275), .Z(n2282) );
  NAND U2576 ( .A(a[35]), .B(b[35]), .Z(n2283) );
  AND U2577 ( .A(n2282), .B(n2283), .Z(n2278) );
  XOR U2578 ( .A(a[36]), .B(b[36]), .Z(n5229) );
  ANDN U2579 ( .B(n5228), .A(n5229), .Z(n2277) );
  OR U2580 ( .A(n2278), .B(n2277), .Z(n2279) );
  AND U2581 ( .A(a[36]), .B(b[36]), .Z(n2281) );
  ANDN U2582 ( .B(n2279), .A(n2281), .Z(n2288) );
  NOR U2583 ( .A(n2283), .B(n2282), .Z(n2280) );
  XNOR U2584 ( .A(n2281), .B(n2280), .Z(n2286) );
  XOR U2585 ( .A(n2283), .B(n2282), .Z(n2284) );
  NAND U2586 ( .A(n2284), .B(n5229), .Z(n2285) );
  NAND U2587 ( .A(n2286), .B(n2285), .Z(n5234) );
  XNOR U2588 ( .A(a[37]), .B(b[37]), .Z(n5233) );
  NAND U2589 ( .A(n5234), .B(n5233), .Z(n2287) );
  NANDN U2590 ( .A(n2288), .B(n2287), .Z(n2294) );
  NAND U2591 ( .A(a[37]), .B(b[37]), .Z(n2295) );
  AND U2592 ( .A(n2294), .B(n2295), .Z(n2290) );
  XOR U2593 ( .A(a[38]), .B(b[38]), .Z(n5239) );
  ANDN U2594 ( .B(n5238), .A(n5239), .Z(n2289) );
  OR U2595 ( .A(n2290), .B(n2289), .Z(n2291) );
  AND U2596 ( .A(a[38]), .B(b[38]), .Z(n2293) );
  ANDN U2597 ( .B(n2291), .A(n2293), .Z(n2300) );
  NOR U2598 ( .A(n2295), .B(n2294), .Z(n2292) );
  XNOR U2599 ( .A(n2293), .B(n2292), .Z(n2298) );
  XOR U2600 ( .A(n2295), .B(n2294), .Z(n2296) );
  NAND U2601 ( .A(n2296), .B(n5239), .Z(n2297) );
  NAND U2602 ( .A(n2298), .B(n2297), .Z(n5244) );
  XNOR U2603 ( .A(a[39]), .B(b[39]), .Z(n5243) );
  NAND U2604 ( .A(n5244), .B(n5243), .Z(n2299) );
  NANDN U2605 ( .A(n2300), .B(n2299), .Z(n2306) );
  NAND U2606 ( .A(a[39]), .B(b[39]), .Z(n2307) );
  AND U2607 ( .A(n2306), .B(n2307), .Z(n2302) );
  XOR U2608 ( .A(a[40]), .B(b[40]), .Z(n5249) );
  ANDN U2609 ( .B(n5248), .A(n5249), .Z(n2301) );
  OR U2610 ( .A(n2302), .B(n2301), .Z(n2303) );
  AND U2611 ( .A(a[40]), .B(b[40]), .Z(n2305) );
  ANDN U2612 ( .B(n2303), .A(n2305), .Z(n2312) );
  NOR U2613 ( .A(n2307), .B(n2306), .Z(n2304) );
  XNOR U2614 ( .A(n2305), .B(n2304), .Z(n2310) );
  XOR U2615 ( .A(n2307), .B(n2306), .Z(n2308) );
  NAND U2616 ( .A(n2308), .B(n5249), .Z(n2309) );
  NAND U2617 ( .A(n2310), .B(n2309), .Z(n5254) );
  XNOR U2618 ( .A(a[41]), .B(b[41]), .Z(n5253) );
  NAND U2619 ( .A(n5254), .B(n5253), .Z(n2311) );
  NANDN U2620 ( .A(n2312), .B(n2311), .Z(n2318) );
  NAND U2621 ( .A(a[41]), .B(b[41]), .Z(n2319) );
  AND U2622 ( .A(n2318), .B(n2319), .Z(n2314) );
  XOR U2623 ( .A(a[42]), .B(b[42]), .Z(n5259) );
  ANDN U2624 ( .B(n5258), .A(n5259), .Z(n2313) );
  OR U2625 ( .A(n2314), .B(n2313), .Z(n2315) );
  AND U2626 ( .A(a[42]), .B(b[42]), .Z(n2317) );
  ANDN U2627 ( .B(n2315), .A(n2317), .Z(n2324) );
  NOR U2628 ( .A(n2319), .B(n2318), .Z(n2316) );
  XNOR U2629 ( .A(n2317), .B(n2316), .Z(n2322) );
  XOR U2630 ( .A(n2319), .B(n2318), .Z(n2320) );
  NAND U2631 ( .A(n2320), .B(n5259), .Z(n2321) );
  NAND U2632 ( .A(n2322), .B(n2321), .Z(n5264) );
  XNOR U2633 ( .A(a[43]), .B(b[43]), .Z(n5263) );
  NAND U2634 ( .A(n5264), .B(n5263), .Z(n2323) );
  NANDN U2635 ( .A(n2324), .B(n2323), .Z(n2330) );
  NAND U2636 ( .A(a[43]), .B(b[43]), .Z(n2331) );
  AND U2637 ( .A(n2330), .B(n2331), .Z(n2326) );
  XOR U2638 ( .A(a[44]), .B(b[44]), .Z(n5269) );
  ANDN U2639 ( .B(n5268), .A(n5269), .Z(n2325) );
  OR U2640 ( .A(n2326), .B(n2325), .Z(n2327) );
  AND U2641 ( .A(a[44]), .B(b[44]), .Z(n2329) );
  ANDN U2642 ( .B(n2327), .A(n2329), .Z(n2336) );
  NOR U2643 ( .A(n2331), .B(n2330), .Z(n2328) );
  XNOR U2644 ( .A(n2329), .B(n2328), .Z(n2334) );
  XOR U2645 ( .A(n2331), .B(n2330), .Z(n2332) );
  NAND U2646 ( .A(n2332), .B(n5269), .Z(n2333) );
  NAND U2647 ( .A(n2334), .B(n2333), .Z(n5274) );
  XNOR U2648 ( .A(a[45]), .B(b[45]), .Z(n5273) );
  NAND U2649 ( .A(n5274), .B(n5273), .Z(n2335) );
  NANDN U2650 ( .A(n2336), .B(n2335), .Z(n2342) );
  NAND U2651 ( .A(a[45]), .B(b[45]), .Z(n2343) );
  AND U2652 ( .A(n2342), .B(n2343), .Z(n2338) );
  XOR U2653 ( .A(a[46]), .B(b[46]), .Z(n5279) );
  ANDN U2654 ( .B(n5278), .A(n5279), .Z(n2337) );
  OR U2655 ( .A(n2338), .B(n2337), .Z(n2339) );
  AND U2656 ( .A(a[46]), .B(b[46]), .Z(n2341) );
  ANDN U2657 ( .B(n2339), .A(n2341), .Z(n2348) );
  NOR U2658 ( .A(n2343), .B(n2342), .Z(n2340) );
  XNOR U2659 ( .A(n2341), .B(n2340), .Z(n2346) );
  XOR U2660 ( .A(n2343), .B(n2342), .Z(n2344) );
  NAND U2661 ( .A(n2344), .B(n5279), .Z(n2345) );
  NAND U2662 ( .A(n2346), .B(n2345), .Z(n5284) );
  XNOR U2663 ( .A(a[47]), .B(b[47]), .Z(n5283) );
  NAND U2664 ( .A(n5284), .B(n5283), .Z(n2347) );
  NANDN U2665 ( .A(n2348), .B(n2347), .Z(n2354) );
  NAND U2666 ( .A(a[47]), .B(b[47]), .Z(n2355) );
  AND U2667 ( .A(n2354), .B(n2355), .Z(n2350) );
  XOR U2668 ( .A(a[48]), .B(b[48]), .Z(n5289) );
  ANDN U2669 ( .B(n5288), .A(n5289), .Z(n2349) );
  OR U2670 ( .A(n2350), .B(n2349), .Z(n2351) );
  AND U2671 ( .A(a[48]), .B(b[48]), .Z(n2353) );
  ANDN U2672 ( .B(n2351), .A(n2353), .Z(n2360) );
  NOR U2673 ( .A(n2355), .B(n2354), .Z(n2352) );
  XNOR U2674 ( .A(n2353), .B(n2352), .Z(n2358) );
  XOR U2675 ( .A(n2355), .B(n2354), .Z(n2356) );
  NAND U2676 ( .A(n2356), .B(n5289), .Z(n2357) );
  NAND U2677 ( .A(n2358), .B(n2357), .Z(n5294) );
  XNOR U2678 ( .A(a[49]), .B(b[49]), .Z(n5293) );
  NAND U2679 ( .A(n5294), .B(n5293), .Z(n2359) );
  NANDN U2680 ( .A(n2360), .B(n2359), .Z(n2366) );
  NAND U2681 ( .A(a[49]), .B(b[49]), .Z(n2367) );
  AND U2682 ( .A(n2366), .B(n2367), .Z(n2362) );
  XOR U2683 ( .A(a[50]), .B(b[50]), .Z(n5299) );
  ANDN U2684 ( .B(n5298), .A(n5299), .Z(n2361) );
  OR U2685 ( .A(n2362), .B(n2361), .Z(n2363) );
  AND U2686 ( .A(a[50]), .B(b[50]), .Z(n2365) );
  ANDN U2687 ( .B(n2363), .A(n2365), .Z(n2372) );
  NOR U2688 ( .A(n2367), .B(n2366), .Z(n2364) );
  XNOR U2689 ( .A(n2365), .B(n2364), .Z(n2370) );
  XOR U2690 ( .A(n2367), .B(n2366), .Z(n2368) );
  NAND U2691 ( .A(n2368), .B(n5299), .Z(n2369) );
  NAND U2692 ( .A(n2370), .B(n2369), .Z(n5304) );
  XNOR U2693 ( .A(a[51]), .B(b[51]), .Z(n5303) );
  NAND U2694 ( .A(n5304), .B(n5303), .Z(n2371) );
  NANDN U2695 ( .A(n2372), .B(n2371), .Z(n2378) );
  NAND U2696 ( .A(a[51]), .B(b[51]), .Z(n2379) );
  AND U2697 ( .A(n2378), .B(n2379), .Z(n2374) );
  XOR U2698 ( .A(a[52]), .B(b[52]), .Z(n5309) );
  ANDN U2699 ( .B(n5308), .A(n5309), .Z(n2373) );
  OR U2700 ( .A(n2374), .B(n2373), .Z(n2375) );
  AND U2701 ( .A(a[52]), .B(b[52]), .Z(n2377) );
  ANDN U2702 ( .B(n2375), .A(n2377), .Z(n2384) );
  NOR U2703 ( .A(n2379), .B(n2378), .Z(n2376) );
  XNOR U2704 ( .A(n2377), .B(n2376), .Z(n2382) );
  XOR U2705 ( .A(n2379), .B(n2378), .Z(n2380) );
  NAND U2706 ( .A(n2380), .B(n5309), .Z(n2381) );
  NAND U2707 ( .A(n2382), .B(n2381), .Z(n5314) );
  XNOR U2708 ( .A(a[53]), .B(b[53]), .Z(n5313) );
  NAND U2709 ( .A(n5314), .B(n5313), .Z(n2383) );
  NANDN U2710 ( .A(n2384), .B(n2383), .Z(n2390) );
  NAND U2711 ( .A(a[53]), .B(b[53]), .Z(n2391) );
  AND U2712 ( .A(n2390), .B(n2391), .Z(n2386) );
  XOR U2713 ( .A(a[54]), .B(b[54]), .Z(n5319) );
  ANDN U2714 ( .B(n5318), .A(n5319), .Z(n2385) );
  OR U2715 ( .A(n2386), .B(n2385), .Z(n2387) );
  AND U2716 ( .A(a[54]), .B(b[54]), .Z(n2389) );
  ANDN U2717 ( .B(n2387), .A(n2389), .Z(n2396) );
  NOR U2718 ( .A(n2391), .B(n2390), .Z(n2388) );
  XNOR U2719 ( .A(n2389), .B(n2388), .Z(n2394) );
  XOR U2720 ( .A(n2391), .B(n2390), .Z(n2392) );
  NAND U2721 ( .A(n2392), .B(n5319), .Z(n2393) );
  NAND U2722 ( .A(n2394), .B(n2393), .Z(n5324) );
  XNOR U2723 ( .A(a[55]), .B(b[55]), .Z(n5323) );
  NAND U2724 ( .A(n5324), .B(n5323), .Z(n2395) );
  NANDN U2725 ( .A(n2396), .B(n2395), .Z(n2402) );
  NAND U2726 ( .A(a[55]), .B(b[55]), .Z(n2403) );
  AND U2727 ( .A(n2402), .B(n2403), .Z(n2398) );
  XOR U2728 ( .A(a[56]), .B(b[56]), .Z(n5329) );
  ANDN U2729 ( .B(n5328), .A(n5329), .Z(n2397) );
  OR U2730 ( .A(n2398), .B(n2397), .Z(n2399) );
  AND U2731 ( .A(a[56]), .B(b[56]), .Z(n2401) );
  ANDN U2732 ( .B(n2399), .A(n2401), .Z(n2408) );
  NOR U2733 ( .A(n2403), .B(n2402), .Z(n2400) );
  XNOR U2734 ( .A(n2401), .B(n2400), .Z(n2406) );
  XOR U2735 ( .A(n2403), .B(n2402), .Z(n2404) );
  NAND U2736 ( .A(n2404), .B(n5329), .Z(n2405) );
  NAND U2737 ( .A(n2406), .B(n2405), .Z(n5334) );
  XNOR U2738 ( .A(a[57]), .B(b[57]), .Z(n5333) );
  NAND U2739 ( .A(n5334), .B(n5333), .Z(n2407) );
  NANDN U2740 ( .A(n2408), .B(n2407), .Z(n2414) );
  NAND U2741 ( .A(a[57]), .B(b[57]), .Z(n2415) );
  AND U2742 ( .A(n2414), .B(n2415), .Z(n2410) );
  XOR U2743 ( .A(a[58]), .B(b[58]), .Z(n5339) );
  ANDN U2744 ( .B(n5338), .A(n5339), .Z(n2409) );
  OR U2745 ( .A(n2410), .B(n2409), .Z(n2411) );
  AND U2746 ( .A(a[58]), .B(b[58]), .Z(n2413) );
  ANDN U2747 ( .B(n2411), .A(n2413), .Z(n2420) );
  NOR U2748 ( .A(n2415), .B(n2414), .Z(n2412) );
  XNOR U2749 ( .A(n2413), .B(n2412), .Z(n2418) );
  XOR U2750 ( .A(n2415), .B(n2414), .Z(n2416) );
  NAND U2751 ( .A(n2416), .B(n5339), .Z(n2417) );
  NAND U2752 ( .A(n2418), .B(n2417), .Z(n5344) );
  XNOR U2753 ( .A(a[59]), .B(b[59]), .Z(n5343) );
  NAND U2754 ( .A(n5344), .B(n5343), .Z(n2419) );
  NANDN U2755 ( .A(n2420), .B(n2419), .Z(n2426) );
  NAND U2756 ( .A(a[59]), .B(b[59]), .Z(n2427) );
  AND U2757 ( .A(n2426), .B(n2427), .Z(n2422) );
  XOR U2758 ( .A(a[60]), .B(b[60]), .Z(n5349) );
  ANDN U2759 ( .B(n5348), .A(n5349), .Z(n2421) );
  OR U2760 ( .A(n2422), .B(n2421), .Z(n2423) );
  AND U2761 ( .A(a[60]), .B(b[60]), .Z(n2425) );
  ANDN U2762 ( .B(n2423), .A(n2425), .Z(n2432) );
  NOR U2763 ( .A(n2427), .B(n2426), .Z(n2424) );
  XNOR U2764 ( .A(n2425), .B(n2424), .Z(n2430) );
  XOR U2765 ( .A(n2427), .B(n2426), .Z(n2428) );
  NAND U2766 ( .A(n2428), .B(n5349), .Z(n2429) );
  NAND U2767 ( .A(n2430), .B(n2429), .Z(n5354) );
  XNOR U2768 ( .A(a[61]), .B(b[61]), .Z(n5353) );
  NAND U2769 ( .A(n5354), .B(n5353), .Z(n2431) );
  NANDN U2770 ( .A(n2432), .B(n2431), .Z(n2438) );
  NAND U2771 ( .A(a[61]), .B(b[61]), .Z(n2439) );
  AND U2772 ( .A(n2438), .B(n2439), .Z(n2434) );
  XOR U2773 ( .A(a[62]), .B(b[62]), .Z(n5359) );
  ANDN U2774 ( .B(n5358), .A(n5359), .Z(n2433) );
  OR U2775 ( .A(n2434), .B(n2433), .Z(n2435) );
  AND U2776 ( .A(a[62]), .B(b[62]), .Z(n2437) );
  ANDN U2777 ( .B(n2435), .A(n2437), .Z(n2444) );
  NOR U2778 ( .A(n2439), .B(n2438), .Z(n2436) );
  XNOR U2779 ( .A(n2437), .B(n2436), .Z(n2442) );
  XOR U2780 ( .A(n2439), .B(n2438), .Z(n2440) );
  NAND U2781 ( .A(n2440), .B(n5359), .Z(n2441) );
  NAND U2782 ( .A(n2442), .B(n2441), .Z(n5364) );
  XNOR U2783 ( .A(a[63]), .B(b[63]), .Z(n5363) );
  NAND U2784 ( .A(n5364), .B(n5363), .Z(n2443) );
  NANDN U2785 ( .A(n2444), .B(n2443), .Z(n2450) );
  NAND U2786 ( .A(a[63]), .B(b[63]), .Z(n2451) );
  AND U2787 ( .A(n2450), .B(n2451), .Z(n2446) );
  XOR U2788 ( .A(a[64]), .B(b[64]), .Z(n5369) );
  ANDN U2789 ( .B(n5368), .A(n5369), .Z(n2445) );
  OR U2790 ( .A(n2446), .B(n2445), .Z(n2447) );
  AND U2791 ( .A(a[64]), .B(b[64]), .Z(n2449) );
  ANDN U2792 ( .B(n2447), .A(n2449), .Z(n2456) );
  NOR U2793 ( .A(n2451), .B(n2450), .Z(n2448) );
  XNOR U2794 ( .A(n2449), .B(n2448), .Z(n2454) );
  XOR U2795 ( .A(n2451), .B(n2450), .Z(n2452) );
  NAND U2796 ( .A(n2452), .B(n5369), .Z(n2453) );
  NAND U2797 ( .A(n2454), .B(n2453), .Z(n5374) );
  XNOR U2798 ( .A(a[65]), .B(b[65]), .Z(n5373) );
  NAND U2799 ( .A(n5374), .B(n5373), .Z(n2455) );
  NANDN U2800 ( .A(n2456), .B(n2455), .Z(n2462) );
  NAND U2801 ( .A(a[65]), .B(b[65]), .Z(n2463) );
  AND U2802 ( .A(n2462), .B(n2463), .Z(n2458) );
  XOR U2803 ( .A(a[66]), .B(b[66]), .Z(n5379) );
  ANDN U2804 ( .B(n5378), .A(n5379), .Z(n2457) );
  OR U2805 ( .A(n2458), .B(n2457), .Z(n2459) );
  AND U2806 ( .A(a[66]), .B(b[66]), .Z(n2461) );
  ANDN U2807 ( .B(n2459), .A(n2461), .Z(n2468) );
  NOR U2808 ( .A(n2463), .B(n2462), .Z(n2460) );
  XNOR U2809 ( .A(n2461), .B(n2460), .Z(n2466) );
  XOR U2810 ( .A(n2463), .B(n2462), .Z(n2464) );
  NAND U2811 ( .A(n2464), .B(n5379), .Z(n2465) );
  NAND U2812 ( .A(n2466), .B(n2465), .Z(n5384) );
  XNOR U2813 ( .A(a[67]), .B(b[67]), .Z(n5383) );
  NAND U2814 ( .A(n5384), .B(n5383), .Z(n2467) );
  NANDN U2815 ( .A(n2468), .B(n2467), .Z(n2474) );
  NAND U2816 ( .A(a[67]), .B(b[67]), .Z(n2475) );
  AND U2817 ( .A(n2474), .B(n2475), .Z(n2470) );
  XOR U2818 ( .A(a[68]), .B(b[68]), .Z(n5389) );
  ANDN U2819 ( .B(n5388), .A(n5389), .Z(n2469) );
  OR U2820 ( .A(n2470), .B(n2469), .Z(n2471) );
  AND U2821 ( .A(a[68]), .B(b[68]), .Z(n2473) );
  ANDN U2822 ( .B(n2471), .A(n2473), .Z(n2480) );
  NOR U2823 ( .A(n2475), .B(n2474), .Z(n2472) );
  XNOR U2824 ( .A(n2473), .B(n2472), .Z(n2478) );
  XOR U2825 ( .A(n2475), .B(n2474), .Z(n2476) );
  NAND U2826 ( .A(n2476), .B(n5389), .Z(n2477) );
  NAND U2827 ( .A(n2478), .B(n2477), .Z(n5394) );
  XNOR U2828 ( .A(a[69]), .B(b[69]), .Z(n5393) );
  NAND U2829 ( .A(n5394), .B(n5393), .Z(n2479) );
  NANDN U2830 ( .A(n2480), .B(n2479), .Z(n2486) );
  NAND U2831 ( .A(a[69]), .B(b[69]), .Z(n2487) );
  AND U2832 ( .A(n2486), .B(n2487), .Z(n2482) );
  XOR U2833 ( .A(a[70]), .B(b[70]), .Z(n5399) );
  ANDN U2834 ( .B(n5398), .A(n5399), .Z(n2481) );
  OR U2835 ( .A(n2482), .B(n2481), .Z(n2483) );
  AND U2836 ( .A(a[70]), .B(b[70]), .Z(n2485) );
  ANDN U2837 ( .B(n2483), .A(n2485), .Z(n2492) );
  NOR U2838 ( .A(n2487), .B(n2486), .Z(n2484) );
  XNOR U2839 ( .A(n2485), .B(n2484), .Z(n2490) );
  XOR U2840 ( .A(n2487), .B(n2486), .Z(n2488) );
  NAND U2841 ( .A(n2488), .B(n5399), .Z(n2489) );
  NAND U2842 ( .A(n2490), .B(n2489), .Z(n5404) );
  XNOR U2843 ( .A(a[71]), .B(b[71]), .Z(n5403) );
  NAND U2844 ( .A(n5404), .B(n5403), .Z(n2491) );
  NANDN U2845 ( .A(n2492), .B(n2491), .Z(n2498) );
  NAND U2846 ( .A(a[71]), .B(b[71]), .Z(n2499) );
  AND U2847 ( .A(n2498), .B(n2499), .Z(n2494) );
  XOR U2848 ( .A(a[72]), .B(b[72]), .Z(n5409) );
  ANDN U2849 ( .B(n5408), .A(n5409), .Z(n2493) );
  OR U2850 ( .A(n2494), .B(n2493), .Z(n2495) );
  AND U2851 ( .A(a[72]), .B(b[72]), .Z(n2497) );
  ANDN U2852 ( .B(n2495), .A(n2497), .Z(n2504) );
  NOR U2853 ( .A(n2499), .B(n2498), .Z(n2496) );
  XNOR U2854 ( .A(n2497), .B(n2496), .Z(n2502) );
  XOR U2855 ( .A(n2499), .B(n2498), .Z(n2500) );
  NAND U2856 ( .A(n2500), .B(n5409), .Z(n2501) );
  NAND U2857 ( .A(n2502), .B(n2501), .Z(n5414) );
  XNOR U2858 ( .A(a[73]), .B(b[73]), .Z(n5413) );
  NAND U2859 ( .A(n5414), .B(n5413), .Z(n2503) );
  NANDN U2860 ( .A(n2504), .B(n2503), .Z(n2510) );
  NAND U2861 ( .A(a[73]), .B(b[73]), .Z(n2511) );
  AND U2862 ( .A(n2510), .B(n2511), .Z(n2506) );
  XOR U2863 ( .A(a[74]), .B(b[74]), .Z(n5419) );
  ANDN U2864 ( .B(n5418), .A(n5419), .Z(n2505) );
  OR U2865 ( .A(n2506), .B(n2505), .Z(n2507) );
  AND U2866 ( .A(a[74]), .B(b[74]), .Z(n2509) );
  ANDN U2867 ( .B(n2507), .A(n2509), .Z(n2516) );
  NOR U2868 ( .A(n2511), .B(n2510), .Z(n2508) );
  XNOR U2869 ( .A(n2509), .B(n2508), .Z(n2514) );
  XOR U2870 ( .A(n2511), .B(n2510), .Z(n2512) );
  NAND U2871 ( .A(n2512), .B(n5419), .Z(n2513) );
  NAND U2872 ( .A(n2514), .B(n2513), .Z(n5424) );
  XNOR U2873 ( .A(a[75]), .B(b[75]), .Z(n5423) );
  NAND U2874 ( .A(n5424), .B(n5423), .Z(n2515) );
  NANDN U2875 ( .A(n2516), .B(n2515), .Z(n2522) );
  NAND U2876 ( .A(a[75]), .B(b[75]), .Z(n2523) );
  AND U2877 ( .A(n2522), .B(n2523), .Z(n2518) );
  XOR U2878 ( .A(a[76]), .B(b[76]), .Z(n5429) );
  ANDN U2879 ( .B(n5428), .A(n5429), .Z(n2517) );
  OR U2880 ( .A(n2518), .B(n2517), .Z(n2519) );
  AND U2881 ( .A(a[76]), .B(b[76]), .Z(n2521) );
  ANDN U2882 ( .B(n2519), .A(n2521), .Z(n2528) );
  NOR U2883 ( .A(n2523), .B(n2522), .Z(n2520) );
  XNOR U2884 ( .A(n2521), .B(n2520), .Z(n2526) );
  XOR U2885 ( .A(n2523), .B(n2522), .Z(n2524) );
  NAND U2886 ( .A(n2524), .B(n5429), .Z(n2525) );
  NAND U2887 ( .A(n2526), .B(n2525), .Z(n5434) );
  XNOR U2888 ( .A(a[77]), .B(b[77]), .Z(n5433) );
  NAND U2889 ( .A(n5434), .B(n5433), .Z(n2527) );
  NANDN U2890 ( .A(n2528), .B(n2527), .Z(n2534) );
  NAND U2891 ( .A(a[77]), .B(b[77]), .Z(n2535) );
  AND U2892 ( .A(n2534), .B(n2535), .Z(n2530) );
  XOR U2893 ( .A(a[78]), .B(b[78]), .Z(n5439) );
  ANDN U2894 ( .B(n5438), .A(n5439), .Z(n2529) );
  OR U2895 ( .A(n2530), .B(n2529), .Z(n2531) );
  AND U2896 ( .A(a[78]), .B(b[78]), .Z(n2533) );
  ANDN U2897 ( .B(n2531), .A(n2533), .Z(n2540) );
  NOR U2898 ( .A(n2535), .B(n2534), .Z(n2532) );
  XNOR U2899 ( .A(n2533), .B(n2532), .Z(n2538) );
  XOR U2900 ( .A(n2535), .B(n2534), .Z(n2536) );
  NAND U2901 ( .A(n2536), .B(n5439), .Z(n2537) );
  NAND U2902 ( .A(n2538), .B(n2537), .Z(n5444) );
  XNOR U2903 ( .A(a[79]), .B(b[79]), .Z(n5443) );
  NAND U2904 ( .A(n5444), .B(n5443), .Z(n2539) );
  NANDN U2905 ( .A(n2540), .B(n2539), .Z(n2546) );
  NAND U2906 ( .A(a[79]), .B(b[79]), .Z(n2547) );
  AND U2907 ( .A(n2546), .B(n2547), .Z(n2542) );
  XOR U2908 ( .A(a[80]), .B(b[80]), .Z(n5449) );
  ANDN U2909 ( .B(n5448), .A(n5449), .Z(n2541) );
  OR U2910 ( .A(n2542), .B(n2541), .Z(n2543) );
  AND U2911 ( .A(a[80]), .B(b[80]), .Z(n2545) );
  ANDN U2912 ( .B(n2543), .A(n2545), .Z(n2552) );
  NOR U2913 ( .A(n2547), .B(n2546), .Z(n2544) );
  XNOR U2914 ( .A(n2545), .B(n2544), .Z(n2550) );
  XOR U2915 ( .A(n2547), .B(n2546), .Z(n2548) );
  NAND U2916 ( .A(n2548), .B(n5449), .Z(n2549) );
  NAND U2917 ( .A(n2550), .B(n2549), .Z(n5454) );
  XNOR U2918 ( .A(a[81]), .B(b[81]), .Z(n5453) );
  NAND U2919 ( .A(n5454), .B(n5453), .Z(n2551) );
  NANDN U2920 ( .A(n2552), .B(n2551), .Z(n2558) );
  NAND U2921 ( .A(a[81]), .B(b[81]), .Z(n2559) );
  AND U2922 ( .A(n2558), .B(n2559), .Z(n2554) );
  XOR U2923 ( .A(a[82]), .B(b[82]), .Z(n5459) );
  ANDN U2924 ( .B(n5458), .A(n5459), .Z(n2553) );
  OR U2925 ( .A(n2554), .B(n2553), .Z(n2555) );
  AND U2926 ( .A(a[82]), .B(b[82]), .Z(n2557) );
  ANDN U2927 ( .B(n2555), .A(n2557), .Z(n2564) );
  NOR U2928 ( .A(n2559), .B(n2558), .Z(n2556) );
  XNOR U2929 ( .A(n2557), .B(n2556), .Z(n2562) );
  XOR U2930 ( .A(n2559), .B(n2558), .Z(n2560) );
  NAND U2931 ( .A(n2560), .B(n5459), .Z(n2561) );
  NAND U2932 ( .A(n2562), .B(n2561), .Z(n5464) );
  XNOR U2933 ( .A(a[83]), .B(b[83]), .Z(n5463) );
  NAND U2934 ( .A(n5464), .B(n5463), .Z(n2563) );
  NANDN U2935 ( .A(n2564), .B(n2563), .Z(n2565) );
  IV U2936 ( .A(n2565), .Z(n2569) );
  AND U2937 ( .A(a[83]), .B(b[83]), .Z(n2570) );
  NOR U2938 ( .A(n2569), .B(n2570), .Z(n2567) );
  XNOR U2939 ( .A(n2570), .B(n2565), .Z(n5469) );
  XNOR U2940 ( .A(a[84]), .B(b[84]), .Z(n5468) );
  AND U2941 ( .A(n5469), .B(n5468), .Z(n2566) );
  OR U2942 ( .A(n2567), .B(n2566), .Z(n2568) );
  AND U2943 ( .A(a[84]), .B(b[84]), .Z(n2572) );
  ANDN U2944 ( .B(n2568), .A(n2572), .Z(n2574) );
  AND U2945 ( .A(n2570), .B(n2569), .Z(n2571) );
  NAND U2946 ( .A(n2572), .B(n2571), .Z(n2577) );
  ANDN U2947 ( .B(n2577), .A(n2574), .Z(n5474) );
  XNOR U2948 ( .A(a[85]), .B(b[85]), .Z(n5473) );
  AND U2949 ( .A(n5474), .B(n5473), .Z(n2573) );
  OR U2950 ( .A(n2574), .B(n2573), .Z(n2575) );
  AND U2951 ( .A(n2576), .B(n2575), .Z(n2580) );
  OR U2952 ( .A(n2577), .B(n2576), .Z(n2578) );
  ANDN U2953 ( .B(n2578), .A(n2580), .Z(n5479) );
  XNOR U2954 ( .A(a[86]), .B(b[86]), .Z(n5478) );
  NAND U2955 ( .A(n5479), .B(n5478), .Z(n2579) );
  NANDN U2956 ( .A(n2580), .B(n2579), .Z(n2586) );
  NAND U2957 ( .A(a[86]), .B(b[86]), .Z(n2587) );
  AND U2958 ( .A(n2586), .B(n2587), .Z(n2582) );
  XOR U2959 ( .A(a[87]), .B(b[87]), .Z(n5484) );
  ANDN U2960 ( .B(n5483), .A(n5484), .Z(n2581) );
  OR U2961 ( .A(n2582), .B(n2581), .Z(n2583) );
  AND U2962 ( .A(a[87]), .B(b[87]), .Z(n2585) );
  ANDN U2963 ( .B(n2583), .A(n2585), .Z(n2592) );
  NOR U2964 ( .A(n2587), .B(n2586), .Z(n2584) );
  XNOR U2965 ( .A(n2585), .B(n2584), .Z(n2590) );
  XOR U2966 ( .A(n2587), .B(n2586), .Z(n2588) );
  NAND U2967 ( .A(n2588), .B(n5484), .Z(n2589) );
  NAND U2968 ( .A(n2590), .B(n2589), .Z(n5489) );
  XNOR U2969 ( .A(a[88]), .B(b[88]), .Z(n5488) );
  NAND U2970 ( .A(n5489), .B(n5488), .Z(n2591) );
  NANDN U2971 ( .A(n2592), .B(n2591), .Z(n2593) );
  IV U2972 ( .A(n2593), .Z(n2597) );
  AND U2973 ( .A(a[88]), .B(b[88]), .Z(n2598) );
  NOR U2974 ( .A(n2597), .B(n2598), .Z(n2595) );
  XNOR U2975 ( .A(n2598), .B(n2593), .Z(n5494) );
  XNOR U2976 ( .A(a[89]), .B(b[89]), .Z(n5493) );
  AND U2977 ( .A(n5494), .B(n5493), .Z(n2594) );
  OR U2978 ( .A(n2595), .B(n2594), .Z(n2596) );
  AND U2979 ( .A(a[89]), .B(b[89]), .Z(n2600) );
  ANDN U2980 ( .B(n2596), .A(n2600), .Z(n2602) );
  AND U2981 ( .A(n2598), .B(n2597), .Z(n2599) );
  NAND U2982 ( .A(n2600), .B(n2599), .Z(n2605) );
  ANDN U2983 ( .B(n2605), .A(n2602), .Z(n5499) );
  XNOR U2984 ( .A(a[90]), .B(b[90]), .Z(n5498) );
  AND U2985 ( .A(n5499), .B(n5498), .Z(n2601) );
  OR U2986 ( .A(n2602), .B(n2601), .Z(n2603) );
  AND U2987 ( .A(a[90]), .B(b[90]), .Z(n2604) );
  ANDN U2988 ( .B(n2603), .A(n2604), .Z(n2608) );
  NANDN U2989 ( .A(n2605), .B(n2604), .Z(n2606) );
  ANDN U2990 ( .B(n2606), .A(n2608), .Z(n5504) );
  XNOR U2991 ( .A(a[91]), .B(b[91]), .Z(n5503) );
  NAND U2992 ( .A(n5504), .B(n5503), .Z(n2607) );
  NANDN U2993 ( .A(n2608), .B(n2607), .Z(n2614) );
  NAND U2994 ( .A(a[91]), .B(b[91]), .Z(n2615) );
  AND U2995 ( .A(n2614), .B(n2615), .Z(n2610) );
  XOR U2996 ( .A(a[92]), .B(b[92]), .Z(n5509) );
  ANDN U2997 ( .B(n5508), .A(n5509), .Z(n2609) );
  OR U2998 ( .A(n2610), .B(n2609), .Z(n2611) );
  AND U2999 ( .A(a[92]), .B(b[92]), .Z(n2613) );
  ANDN U3000 ( .B(n2611), .A(n2613), .Z(n2620) );
  NOR U3001 ( .A(n2615), .B(n2614), .Z(n2612) );
  XNOR U3002 ( .A(n2613), .B(n2612), .Z(n2618) );
  XOR U3003 ( .A(n2615), .B(n2614), .Z(n2616) );
  NAND U3004 ( .A(n2616), .B(n5509), .Z(n2617) );
  NAND U3005 ( .A(n2618), .B(n2617), .Z(n5514) );
  XNOR U3006 ( .A(a[93]), .B(b[93]), .Z(n5513) );
  NAND U3007 ( .A(n5514), .B(n5513), .Z(n2619) );
  NANDN U3008 ( .A(n2620), .B(n2619), .Z(n2621) );
  IV U3009 ( .A(n2621), .Z(n2625) );
  AND U3010 ( .A(a[93]), .B(b[93]), .Z(n2626) );
  NOR U3011 ( .A(n2625), .B(n2626), .Z(n2623) );
  XNOR U3012 ( .A(n2626), .B(n2621), .Z(n5519) );
  XNOR U3013 ( .A(a[94]), .B(b[94]), .Z(n5518) );
  AND U3014 ( .A(n5519), .B(n5518), .Z(n2622) );
  OR U3015 ( .A(n2623), .B(n2622), .Z(n2624) );
  AND U3016 ( .A(a[94]), .B(b[94]), .Z(n2628) );
  ANDN U3017 ( .B(n2624), .A(n2628), .Z(n2630) );
  AND U3018 ( .A(n2626), .B(n2625), .Z(n2627) );
  NAND U3019 ( .A(n2628), .B(n2627), .Z(n2633) );
  ANDN U3020 ( .B(n2633), .A(n2630), .Z(n5524) );
  XNOR U3021 ( .A(a[95]), .B(b[95]), .Z(n5523) );
  AND U3022 ( .A(n5524), .B(n5523), .Z(n2629) );
  OR U3023 ( .A(n2630), .B(n2629), .Z(n2631) );
  AND U3024 ( .A(a[95]), .B(b[95]), .Z(n2632) );
  ANDN U3025 ( .B(n2631), .A(n2632), .Z(n2636) );
  NANDN U3026 ( .A(n2633), .B(n2632), .Z(n2634) );
  ANDN U3027 ( .B(n2634), .A(n2636), .Z(n5529) );
  XNOR U3028 ( .A(a[96]), .B(b[96]), .Z(n5528) );
  NAND U3029 ( .A(n5529), .B(n5528), .Z(n2635) );
  NANDN U3030 ( .A(n2636), .B(n2635), .Z(n2642) );
  NAND U3031 ( .A(a[96]), .B(b[96]), .Z(n2643) );
  AND U3032 ( .A(n2642), .B(n2643), .Z(n2638) );
  XOR U3033 ( .A(a[97]), .B(b[97]), .Z(n5534) );
  ANDN U3034 ( .B(n5533), .A(n5534), .Z(n2637) );
  OR U3035 ( .A(n2638), .B(n2637), .Z(n2639) );
  AND U3036 ( .A(a[97]), .B(b[97]), .Z(n2641) );
  ANDN U3037 ( .B(n2639), .A(n2641), .Z(n2648) );
  NOR U3038 ( .A(n2643), .B(n2642), .Z(n2640) );
  XNOR U3039 ( .A(n2641), .B(n2640), .Z(n2646) );
  XOR U3040 ( .A(n2643), .B(n2642), .Z(n2644) );
  NAND U3041 ( .A(n2644), .B(n5534), .Z(n2645) );
  NAND U3042 ( .A(n2646), .B(n2645), .Z(n5539) );
  XNOR U3043 ( .A(a[98]), .B(b[98]), .Z(n5538) );
  NAND U3044 ( .A(n5539), .B(n5538), .Z(n2647) );
  NANDN U3045 ( .A(n2648), .B(n2647), .Z(n2654) );
  NAND U3046 ( .A(a[98]), .B(b[98]), .Z(n2655) );
  AND U3047 ( .A(n2654), .B(n2655), .Z(n2650) );
  XOR U3048 ( .A(a[99]), .B(b[99]), .Z(n5544) );
  ANDN U3049 ( .B(n5543), .A(n5544), .Z(n2649) );
  OR U3050 ( .A(n2650), .B(n2649), .Z(n2651) );
  AND U3051 ( .A(a[99]), .B(b[99]), .Z(n2653) );
  ANDN U3052 ( .B(n2651), .A(n2653), .Z(n2660) );
  NOR U3053 ( .A(n2655), .B(n2654), .Z(n2652) );
  XNOR U3054 ( .A(n2653), .B(n2652), .Z(n2658) );
  XOR U3055 ( .A(n2655), .B(n2654), .Z(n2656) );
  NAND U3056 ( .A(n2656), .B(n5544), .Z(n2657) );
  NAND U3057 ( .A(n2658), .B(n2657), .Z(n5549) );
  XNOR U3058 ( .A(a[100]), .B(b[100]), .Z(n5548) );
  NAND U3059 ( .A(n5549), .B(n5548), .Z(n2659) );
  NANDN U3060 ( .A(n2660), .B(n2659), .Z(n2666) );
  NAND U3061 ( .A(a[100]), .B(b[100]), .Z(n2667) );
  AND U3062 ( .A(n2666), .B(n2667), .Z(n2662) );
  XOR U3063 ( .A(a[101]), .B(b[101]), .Z(n5554) );
  ANDN U3064 ( .B(n5553), .A(n5554), .Z(n2661) );
  OR U3065 ( .A(n2662), .B(n2661), .Z(n2663) );
  AND U3066 ( .A(a[101]), .B(b[101]), .Z(n2665) );
  ANDN U3067 ( .B(n2663), .A(n2665), .Z(n2672) );
  NOR U3068 ( .A(n2667), .B(n2666), .Z(n2664) );
  XNOR U3069 ( .A(n2665), .B(n2664), .Z(n2670) );
  XOR U3070 ( .A(n2667), .B(n2666), .Z(n2668) );
  NAND U3071 ( .A(n2668), .B(n5554), .Z(n2669) );
  NAND U3072 ( .A(n2670), .B(n2669), .Z(n5559) );
  XNOR U3073 ( .A(a[102]), .B(b[102]), .Z(n5558) );
  NAND U3074 ( .A(n5559), .B(n5558), .Z(n2671) );
  NANDN U3075 ( .A(n2672), .B(n2671), .Z(n2678) );
  NAND U3076 ( .A(a[102]), .B(b[102]), .Z(n2679) );
  AND U3077 ( .A(n2678), .B(n2679), .Z(n2674) );
  XOR U3078 ( .A(a[103]), .B(b[103]), .Z(n5564) );
  ANDN U3079 ( .B(n5563), .A(n5564), .Z(n2673) );
  OR U3080 ( .A(n2674), .B(n2673), .Z(n2675) );
  AND U3081 ( .A(a[103]), .B(b[103]), .Z(n2677) );
  ANDN U3082 ( .B(n2675), .A(n2677), .Z(n2684) );
  NOR U3083 ( .A(n2679), .B(n2678), .Z(n2676) );
  XNOR U3084 ( .A(n2677), .B(n2676), .Z(n2682) );
  XOR U3085 ( .A(n2679), .B(n2678), .Z(n2680) );
  NAND U3086 ( .A(n2680), .B(n5564), .Z(n2681) );
  NAND U3087 ( .A(n2682), .B(n2681), .Z(n5569) );
  XNOR U3088 ( .A(a[104]), .B(b[104]), .Z(n5568) );
  NAND U3089 ( .A(n5569), .B(n5568), .Z(n2683) );
  NANDN U3090 ( .A(n2684), .B(n2683), .Z(n2690) );
  NAND U3091 ( .A(a[104]), .B(b[104]), .Z(n2691) );
  AND U3092 ( .A(n2690), .B(n2691), .Z(n2686) );
  XOR U3093 ( .A(a[105]), .B(b[105]), .Z(n5574) );
  ANDN U3094 ( .B(n5573), .A(n5574), .Z(n2685) );
  OR U3095 ( .A(n2686), .B(n2685), .Z(n2687) );
  AND U3096 ( .A(a[105]), .B(b[105]), .Z(n2689) );
  ANDN U3097 ( .B(n2687), .A(n2689), .Z(n2696) );
  NOR U3098 ( .A(n2691), .B(n2690), .Z(n2688) );
  XNOR U3099 ( .A(n2689), .B(n2688), .Z(n2694) );
  XOR U3100 ( .A(n2691), .B(n2690), .Z(n2692) );
  NAND U3101 ( .A(n2692), .B(n5574), .Z(n2693) );
  NAND U3102 ( .A(n2694), .B(n2693), .Z(n5579) );
  XNOR U3103 ( .A(a[106]), .B(b[106]), .Z(n5578) );
  NAND U3104 ( .A(n5579), .B(n5578), .Z(n2695) );
  NANDN U3105 ( .A(n2696), .B(n2695), .Z(n2702) );
  NAND U3106 ( .A(a[106]), .B(b[106]), .Z(n2703) );
  AND U3107 ( .A(n2702), .B(n2703), .Z(n2698) );
  XOR U3108 ( .A(a[107]), .B(b[107]), .Z(n5584) );
  ANDN U3109 ( .B(n5583), .A(n5584), .Z(n2697) );
  OR U3110 ( .A(n2698), .B(n2697), .Z(n2699) );
  AND U3111 ( .A(a[107]), .B(b[107]), .Z(n2701) );
  ANDN U3112 ( .B(n2699), .A(n2701), .Z(n2708) );
  NOR U3113 ( .A(n2703), .B(n2702), .Z(n2700) );
  XNOR U3114 ( .A(n2701), .B(n2700), .Z(n2706) );
  XOR U3115 ( .A(n2703), .B(n2702), .Z(n2704) );
  NAND U3116 ( .A(n2704), .B(n5584), .Z(n2705) );
  NAND U3117 ( .A(n2706), .B(n2705), .Z(n5589) );
  XNOR U3118 ( .A(a[108]), .B(b[108]), .Z(n5588) );
  NAND U3119 ( .A(n5589), .B(n5588), .Z(n2707) );
  NANDN U3120 ( .A(n2708), .B(n2707), .Z(n2714) );
  NAND U3121 ( .A(a[108]), .B(b[108]), .Z(n2715) );
  AND U3122 ( .A(n2714), .B(n2715), .Z(n2710) );
  XOR U3123 ( .A(a[109]), .B(b[109]), .Z(n5594) );
  ANDN U3124 ( .B(n5593), .A(n5594), .Z(n2709) );
  OR U3125 ( .A(n2710), .B(n2709), .Z(n2711) );
  AND U3126 ( .A(a[109]), .B(b[109]), .Z(n2713) );
  ANDN U3127 ( .B(n2711), .A(n2713), .Z(n2720) );
  NOR U3128 ( .A(n2715), .B(n2714), .Z(n2712) );
  XNOR U3129 ( .A(n2713), .B(n2712), .Z(n2718) );
  XOR U3130 ( .A(n2715), .B(n2714), .Z(n2716) );
  NAND U3131 ( .A(n2716), .B(n5594), .Z(n2717) );
  NAND U3132 ( .A(n2718), .B(n2717), .Z(n5599) );
  XNOR U3133 ( .A(a[110]), .B(b[110]), .Z(n5598) );
  NAND U3134 ( .A(n5599), .B(n5598), .Z(n2719) );
  NANDN U3135 ( .A(n2720), .B(n2719), .Z(n2726) );
  NAND U3136 ( .A(a[110]), .B(b[110]), .Z(n2727) );
  AND U3137 ( .A(n2726), .B(n2727), .Z(n2722) );
  XOR U3138 ( .A(a[111]), .B(b[111]), .Z(n5604) );
  ANDN U3139 ( .B(n5603), .A(n5604), .Z(n2721) );
  OR U3140 ( .A(n2722), .B(n2721), .Z(n2723) );
  AND U3141 ( .A(a[111]), .B(b[111]), .Z(n2725) );
  ANDN U3142 ( .B(n2723), .A(n2725), .Z(n2732) );
  NOR U3143 ( .A(n2727), .B(n2726), .Z(n2724) );
  XNOR U3144 ( .A(n2725), .B(n2724), .Z(n2730) );
  XOR U3145 ( .A(n2727), .B(n2726), .Z(n2728) );
  NAND U3146 ( .A(n2728), .B(n5604), .Z(n2729) );
  NAND U3147 ( .A(n2730), .B(n2729), .Z(n5609) );
  XNOR U3148 ( .A(a[112]), .B(b[112]), .Z(n5608) );
  NAND U3149 ( .A(n5609), .B(n5608), .Z(n2731) );
  NANDN U3150 ( .A(n2732), .B(n2731), .Z(n2738) );
  NAND U3151 ( .A(a[112]), .B(b[112]), .Z(n2739) );
  AND U3152 ( .A(n2738), .B(n2739), .Z(n2734) );
  XOR U3153 ( .A(a[113]), .B(b[113]), .Z(n5614) );
  ANDN U3154 ( .B(n5613), .A(n5614), .Z(n2733) );
  OR U3155 ( .A(n2734), .B(n2733), .Z(n2735) );
  AND U3156 ( .A(a[113]), .B(b[113]), .Z(n2737) );
  ANDN U3157 ( .B(n2735), .A(n2737), .Z(n2744) );
  NOR U3158 ( .A(n2739), .B(n2738), .Z(n2736) );
  XNOR U3159 ( .A(n2737), .B(n2736), .Z(n2742) );
  XOR U3160 ( .A(n2739), .B(n2738), .Z(n2740) );
  NAND U3161 ( .A(n2740), .B(n5614), .Z(n2741) );
  NAND U3162 ( .A(n2742), .B(n2741), .Z(n5619) );
  XNOR U3163 ( .A(a[114]), .B(b[114]), .Z(n5618) );
  NAND U3164 ( .A(n5619), .B(n5618), .Z(n2743) );
  NANDN U3165 ( .A(n2744), .B(n2743), .Z(n2750) );
  NAND U3166 ( .A(a[114]), .B(b[114]), .Z(n2751) );
  AND U3167 ( .A(n2750), .B(n2751), .Z(n2746) );
  XOR U3168 ( .A(a[115]), .B(b[115]), .Z(n5624) );
  ANDN U3169 ( .B(n5623), .A(n5624), .Z(n2745) );
  OR U3170 ( .A(n2746), .B(n2745), .Z(n2747) );
  AND U3171 ( .A(a[115]), .B(b[115]), .Z(n2749) );
  ANDN U3172 ( .B(n2747), .A(n2749), .Z(n2756) );
  NOR U3173 ( .A(n2751), .B(n2750), .Z(n2748) );
  XNOR U3174 ( .A(n2749), .B(n2748), .Z(n2754) );
  XOR U3175 ( .A(n2751), .B(n2750), .Z(n2752) );
  NAND U3176 ( .A(n2752), .B(n5624), .Z(n2753) );
  NAND U3177 ( .A(n2754), .B(n2753), .Z(n5629) );
  XNOR U3178 ( .A(a[116]), .B(b[116]), .Z(n5628) );
  NAND U3179 ( .A(n5629), .B(n5628), .Z(n2755) );
  NANDN U3180 ( .A(n2756), .B(n2755), .Z(n2762) );
  NAND U3181 ( .A(a[116]), .B(b[116]), .Z(n2763) );
  AND U3182 ( .A(n2762), .B(n2763), .Z(n2758) );
  XOR U3183 ( .A(a[117]), .B(b[117]), .Z(n5634) );
  ANDN U3184 ( .B(n5633), .A(n5634), .Z(n2757) );
  OR U3185 ( .A(n2758), .B(n2757), .Z(n2759) );
  AND U3186 ( .A(a[117]), .B(b[117]), .Z(n2761) );
  ANDN U3187 ( .B(n2759), .A(n2761), .Z(n2768) );
  NOR U3188 ( .A(n2763), .B(n2762), .Z(n2760) );
  XNOR U3189 ( .A(n2761), .B(n2760), .Z(n2766) );
  XOR U3190 ( .A(n2763), .B(n2762), .Z(n2764) );
  NAND U3191 ( .A(n2764), .B(n5634), .Z(n2765) );
  NAND U3192 ( .A(n2766), .B(n2765), .Z(n5639) );
  XNOR U3193 ( .A(a[118]), .B(b[118]), .Z(n5638) );
  NAND U3194 ( .A(n5639), .B(n5638), .Z(n2767) );
  NANDN U3195 ( .A(n2768), .B(n2767), .Z(n2774) );
  NAND U3196 ( .A(a[118]), .B(b[118]), .Z(n2775) );
  AND U3197 ( .A(n2774), .B(n2775), .Z(n2770) );
  XOR U3198 ( .A(a[119]), .B(b[119]), .Z(n5644) );
  ANDN U3199 ( .B(n5643), .A(n5644), .Z(n2769) );
  OR U3200 ( .A(n2770), .B(n2769), .Z(n2771) );
  AND U3201 ( .A(a[119]), .B(b[119]), .Z(n2773) );
  ANDN U3202 ( .B(n2771), .A(n2773), .Z(n2780) );
  NOR U3203 ( .A(n2775), .B(n2774), .Z(n2772) );
  XNOR U3204 ( .A(n2773), .B(n2772), .Z(n2778) );
  XOR U3205 ( .A(n2775), .B(n2774), .Z(n2776) );
  NAND U3206 ( .A(n2776), .B(n5644), .Z(n2777) );
  NAND U3207 ( .A(n2778), .B(n2777), .Z(n5649) );
  XNOR U3208 ( .A(a[120]), .B(b[120]), .Z(n5648) );
  NAND U3209 ( .A(n5649), .B(n5648), .Z(n2779) );
  NANDN U3210 ( .A(n2780), .B(n2779), .Z(n2786) );
  NAND U3211 ( .A(a[120]), .B(b[120]), .Z(n2787) );
  AND U3212 ( .A(n2786), .B(n2787), .Z(n2782) );
  XOR U3213 ( .A(a[121]), .B(b[121]), .Z(n5654) );
  ANDN U3214 ( .B(n5653), .A(n5654), .Z(n2781) );
  OR U3215 ( .A(n2782), .B(n2781), .Z(n2783) );
  AND U3216 ( .A(a[121]), .B(b[121]), .Z(n2785) );
  ANDN U3217 ( .B(n2783), .A(n2785), .Z(n2792) );
  NOR U3218 ( .A(n2787), .B(n2786), .Z(n2784) );
  XNOR U3219 ( .A(n2785), .B(n2784), .Z(n2790) );
  XOR U3220 ( .A(n2787), .B(n2786), .Z(n2788) );
  NAND U3221 ( .A(n2788), .B(n5654), .Z(n2789) );
  NAND U3222 ( .A(n2790), .B(n2789), .Z(n5659) );
  XNOR U3223 ( .A(a[122]), .B(b[122]), .Z(n5658) );
  NAND U3224 ( .A(n5659), .B(n5658), .Z(n2791) );
  NANDN U3225 ( .A(n2792), .B(n2791), .Z(n2798) );
  NAND U3226 ( .A(a[122]), .B(b[122]), .Z(n2799) );
  AND U3227 ( .A(n2798), .B(n2799), .Z(n2794) );
  XOR U3228 ( .A(a[123]), .B(b[123]), .Z(n5664) );
  ANDN U3229 ( .B(n5663), .A(n5664), .Z(n2793) );
  OR U3230 ( .A(n2794), .B(n2793), .Z(n2795) );
  AND U3231 ( .A(a[123]), .B(b[123]), .Z(n2797) );
  ANDN U3232 ( .B(n2795), .A(n2797), .Z(n2804) );
  NOR U3233 ( .A(n2799), .B(n2798), .Z(n2796) );
  XNOR U3234 ( .A(n2797), .B(n2796), .Z(n2802) );
  XOR U3235 ( .A(n2799), .B(n2798), .Z(n2800) );
  NAND U3236 ( .A(n2800), .B(n5664), .Z(n2801) );
  NAND U3237 ( .A(n2802), .B(n2801), .Z(n5669) );
  XNOR U3238 ( .A(a[124]), .B(b[124]), .Z(n5668) );
  NAND U3239 ( .A(n5669), .B(n5668), .Z(n2803) );
  NANDN U3240 ( .A(n2804), .B(n2803), .Z(n2805) );
  IV U3241 ( .A(n2805), .Z(n2809) );
  AND U3242 ( .A(a[124]), .B(b[124]), .Z(n2810) );
  NOR U3243 ( .A(n2809), .B(n2810), .Z(n2807) );
  XNOR U3244 ( .A(n2810), .B(n2805), .Z(n5674) );
  XNOR U3245 ( .A(a[125]), .B(b[125]), .Z(n5673) );
  AND U3246 ( .A(n5674), .B(n5673), .Z(n2806) );
  OR U3247 ( .A(n2807), .B(n2806), .Z(n2808) );
  AND U3248 ( .A(a[125]), .B(b[125]), .Z(n2812) );
  ANDN U3249 ( .B(n2808), .A(n2812), .Z(n2814) );
  AND U3250 ( .A(n2810), .B(n2809), .Z(n2811) );
  NAND U3251 ( .A(n2812), .B(n2811), .Z(n2817) );
  ANDN U3252 ( .B(n2817), .A(n2814), .Z(n5679) );
  XNOR U3253 ( .A(a[126]), .B(b[126]), .Z(n5678) );
  AND U3254 ( .A(n5679), .B(n5678), .Z(n2813) );
  OR U3255 ( .A(n2814), .B(n2813), .Z(n2815) );
  AND U3256 ( .A(n2816), .B(n2815), .Z(n2820) );
  OR U3257 ( .A(n2817), .B(n2816), .Z(n2818) );
  ANDN U3258 ( .B(n2818), .A(n2820), .Z(n5684) );
  XNOR U3259 ( .A(a[127]), .B(b[127]), .Z(n5683) );
  NAND U3260 ( .A(n5684), .B(n5683), .Z(n2819) );
  NANDN U3261 ( .A(n2820), .B(n2819), .Z(n2826) );
  NAND U3262 ( .A(a[127]), .B(b[127]), .Z(n2827) );
  AND U3263 ( .A(n2826), .B(n2827), .Z(n2822) );
  XOR U3264 ( .A(a[128]), .B(b[128]), .Z(n5689) );
  ANDN U3265 ( .B(n5688), .A(n5689), .Z(n2821) );
  OR U3266 ( .A(n2822), .B(n2821), .Z(n2823) );
  AND U3267 ( .A(a[128]), .B(b[128]), .Z(n2825) );
  ANDN U3268 ( .B(n2823), .A(n2825), .Z(n2832) );
  NOR U3269 ( .A(n2827), .B(n2826), .Z(n2824) );
  XNOR U3270 ( .A(n2825), .B(n2824), .Z(n2830) );
  XOR U3271 ( .A(n2827), .B(n2826), .Z(n2828) );
  NAND U3272 ( .A(n2828), .B(n5689), .Z(n2829) );
  NAND U3273 ( .A(n2830), .B(n2829), .Z(n5694) );
  XNOR U3274 ( .A(a[129]), .B(b[129]), .Z(n5693) );
  NAND U3275 ( .A(n5694), .B(n5693), .Z(n2831) );
  NANDN U3276 ( .A(n2832), .B(n2831), .Z(n2838) );
  NAND U3277 ( .A(a[129]), .B(b[129]), .Z(n2839) );
  AND U3278 ( .A(n2838), .B(n2839), .Z(n2834) );
  XOR U3279 ( .A(a[130]), .B(b[130]), .Z(n5699) );
  ANDN U3280 ( .B(n5698), .A(n5699), .Z(n2833) );
  OR U3281 ( .A(n2834), .B(n2833), .Z(n2835) );
  AND U3282 ( .A(a[130]), .B(b[130]), .Z(n2837) );
  ANDN U3283 ( .B(n2835), .A(n2837), .Z(n2844) );
  NOR U3284 ( .A(n2839), .B(n2838), .Z(n2836) );
  XNOR U3285 ( .A(n2837), .B(n2836), .Z(n2842) );
  XOR U3286 ( .A(n2839), .B(n2838), .Z(n2840) );
  NAND U3287 ( .A(n2840), .B(n5699), .Z(n2841) );
  NAND U3288 ( .A(n2842), .B(n2841), .Z(n5704) );
  XNOR U3289 ( .A(a[131]), .B(b[131]), .Z(n5703) );
  NAND U3290 ( .A(n5704), .B(n5703), .Z(n2843) );
  NANDN U3291 ( .A(n2844), .B(n2843), .Z(n2850) );
  NAND U3292 ( .A(a[131]), .B(b[131]), .Z(n2851) );
  AND U3293 ( .A(n2850), .B(n2851), .Z(n2846) );
  XOR U3294 ( .A(a[132]), .B(b[132]), .Z(n5709) );
  ANDN U3295 ( .B(n5708), .A(n5709), .Z(n2845) );
  OR U3296 ( .A(n2846), .B(n2845), .Z(n2847) );
  AND U3297 ( .A(a[132]), .B(b[132]), .Z(n2849) );
  ANDN U3298 ( .B(n2847), .A(n2849), .Z(n2856) );
  NOR U3299 ( .A(n2851), .B(n2850), .Z(n2848) );
  XNOR U3300 ( .A(n2849), .B(n2848), .Z(n2854) );
  XOR U3301 ( .A(n2851), .B(n2850), .Z(n2852) );
  NAND U3302 ( .A(n2852), .B(n5709), .Z(n2853) );
  NAND U3303 ( .A(n2854), .B(n2853), .Z(n5714) );
  XNOR U3304 ( .A(a[133]), .B(b[133]), .Z(n5713) );
  NAND U3305 ( .A(n5714), .B(n5713), .Z(n2855) );
  NANDN U3306 ( .A(n2856), .B(n2855), .Z(n2862) );
  NAND U3307 ( .A(a[133]), .B(b[133]), .Z(n2863) );
  AND U3308 ( .A(n2862), .B(n2863), .Z(n2858) );
  XOR U3309 ( .A(a[134]), .B(b[134]), .Z(n5719) );
  ANDN U3310 ( .B(n5718), .A(n5719), .Z(n2857) );
  OR U3311 ( .A(n2858), .B(n2857), .Z(n2859) );
  AND U3312 ( .A(a[134]), .B(b[134]), .Z(n2861) );
  ANDN U3313 ( .B(n2859), .A(n2861), .Z(n2868) );
  NOR U3314 ( .A(n2863), .B(n2862), .Z(n2860) );
  XNOR U3315 ( .A(n2861), .B(n2860), .Z(n2866) );
  XOR U3316 ( .A(n2863), .B(n2862), .Z(n2864) );
  NAND U3317 ( .A(n2864), .B(n5719), .Z(n2865) );
  NAND U3318 ( .A(n2866), .B(n2865), .Z(n5724) );
  XNOR U3319 ( .A(a[135]), .B(b[135]), .Z(n5723) );
  NAND U3320 ( .A(n5724), .B(n5723), .Z(n2867) );
  NANDN U3321 ( .A(n2868), .B(n2867), .Z(n2874) );
  NAND U3322 ( .A(a[135]), .B(b[135]), .Z(n2875) );
  AND U3323 ( .A(n2874), .B(n2875), .Z(n2870) );
  XOR U3324 ( .A(a[136]), .B(b[136]), .Z(n5729) );
  ANDN U3325 ( .B(n5728), .A(n5729), .Z(n2869) );
  OR U3326 ( .A(n2870), .B(n2869), .Z(n2871) );
  AND U3327 ( .A(a[136]), .B(b[136]), .Z(n2873) );
  ANDN U3328 ( .B(n2871), .A(n2873), .Z(n2880) );
  NOR U3329 ( .A(n2875), .B(n2874), .Z(n2872) );
  XNOR U3330 ( .A(n2873), .B(n2872), .Z(n2878) );
  XOR U3331 ( .A(n2875), .B(n2874), .Z(n2876) );
  NAND U3332 ( .A(n2876), .B(n5729), .Z(n2877) );
  NAND U3333 ( .A(n2878), .B(n2877), .Z(n5734) );
  XNOR U3334 ( .A(a[137]), .B(b[137]), .Z(n5733) );
  NAND U3335 ( .A(n5734), .B(n5733), .Z(n2879) );
  NANDN U3336 ( .A(n2880), .B(n2879), .Z(n2886) );
  NAND U3337 ( .A(a[137]), .B(b[137]), .Z(n2887) );
  AND U3338 ( .A(n2886), .B(n2887), .Z(n2882) );
  XOR U3339 ( .A(a[138]), .B(b[138]), .Z(n5739) );
  ANDN U3340 ( .B(n5738), .A(n5739), .Z(n2881) );
  OR U3341 ( .A(n2882), .B(n2881), .Z(n2883) );
  AND U3342 ( .A(a[138]), .B(b[138]), .Z(n2885) );
  ANDN U3343 ( .B(n2883), .A(n2885), .Z(n2892) );
  NOR U3344 ( .A(n2887), .B(n2886), .Z(n2884) );
  XNOR U3345 ( .A(n2885), .B(n2884), .Z(n2890) );
  XOR U3346 ( .A(n2887), .B(n2886), .Z(n2888) );
  NAND U3347 ( .A(n2888), .B(n5739), .Z(n2889) );
  NAND U3348 ( .A(n2890), .B(n2889), .Z(n5744) );
  XNOR U3349 ( .A(a[139]), .B(b[139]), .Z(n5743) );
  NAND U3350 ( .A(n5744), .B(n5743), .Z(n2891) );
  NANDN U3351 ( .A(n2892), .B(n2891), .Z(n2898) );
  NAND U3352 ( .A(a[139]), .B(b[139]), .Z(n2899) );
  AND U3353 ( .A(n2898), .B(n2899), .Z(n2894) );
  XOR U3354 ( .A(a[140]), .B(b[140]), .Z(n5749) );
  ANDN U3355 ( .B(n5748), .A(n5749), .Z(n2893) );
  OR U3356 ( .A(n2894), .B(n2893), .Z(n2895) );
  AND U3357 ( .A(a[140]), .B(b[140]), .Z(n2897) );
  ANDN U3358 ( .B(n2895), .A(n2897), .Z(n2904) );
  NOR U3359 ( .A(n2899), .B(n2898), .Z(n2896) );
  XNOR U3360 ( .A(n2897), .B(n2896), .Z(n2902) );
  XOR U3361 ( .A(n2899), .B(n2898), .Z(n2900) );
  NAND U3362 ( .A(n2900), .B(n5749), .Z(n2901) );
  NAND U3363 ( .A(n2902), .B(n2901), .Z(n5754) );
  XNOR U3364 ( .A(a[141]), .B(b[141]), .Z(n5753) );
  NAND U3365 ( .A(n5754), .B(n5753), .Z(n2903) );
  NANDN U3366 ( .A(n2904), .B(n2903), .Z(n2910) );
  NAND U3367 ( .A(a[141]), .B(b[141]), .Z(n2911) );
  AND U3368 ( .A(n2910), .B(n2911), .Z(n2906) );
  XOR U3369 ( .A(a[142]), .B(b[142]), .Z(n5759) );
  ANDN U3370 ( .B(n5758), .A(n5759), .Z(n2905) );
  OR U3371 ( .A(n2906), .B(n2905), .Z(n2907) );
  AND U3372 ( .A(a[142]), .B(b[142]), .Z(n2909) );
  ANDN U3373 ( .B(n2907), .A(n2909), .Z(n2916) );
  NOR U3374 ( .A(n2911), .B(n2910), .Z(n2908) );
  XNOR U3375 ( .A(n2909), .B(n2908), .Z(n2914) );
  XOR U3376 ( .A(n2911), .B(n2910), .Z(n2912) );
  NAND U3377 ( .A(n2912), .B(n5759), .Z(n2913) );
  NAND U3378 ( .A(n2914), .B(n2913), .Z(n5764) );
  XNOR U3379 ( .A(a[143]), .B(b[143]), .Z(n5763) );
  NAND U3380 ( .A(n5764), .B(n5763), .Z(n2915) );
  NANDN U3381 ( .A(n2916), .B(n2915), .Z(n2922) );
  NAND U3382 ( .A(a[143]), .B(b[143]), .Z(n2923) );
  AND U3383 ( .A(n2922), .B(n2923), .Z(n2918) );
  XOR U3384 ( .A(a[144]), .B(b[144]), .Z(n5769) );
  ANDN U3385 ( .B(n5768), .A(n5769), .Z(n2917) );
  OR U3386 ( .A(n2918), .B(n2917), .Z(n2919) );
  AND U3387 ( .A(a[144]), .B(b[144]), .Z(n2921) );
  ANDN U3388 ( .B(n2919), .A(n2921), .Z(n2928) );
  NOR U3389 ( .A(n2923), .B(n2922), .Z(n2920) );
  XNOR U3390 ( .A(n2921), .B(n2920), .Z(n2926) );
  XOR U3391 ( .A(n2923), .B(n2922), .Z(n2924) );
  NAND U3392 ( .A(n2924), .B(n5769), .Z(n2925) );
  NAND U3393 ( .A(n2926), .B(n2925), .Z(n5774) );
  XNOR U3394 ( .A(a[145]), .B(b[145]), .Z(n5773) );
  NAND U3395 ( .A(n5774), .B(n5773), .Z(n2927) );
  NANDN U3396 ( .A(n2928), .B(n2927), .Z(n2934) );
  NAND U3397 ( .A(a[145]), .B(b[145]), .Z(n2935) );
  AND U3398 ( .A(n2934), .B(n2935), .Z(n2930) );
  XOR U3399 ( .A(a[146]), .B(b[146]), .Z(n5779) );
  ANDN U3400 ( .B(n5778), .A(n5779), .Z(n2929) );
  OR U3401 ( .A(n2930), .B(n2929), .Z(n2931) );
  AND U3402 ( .A(a[146]), .B(b[146]), .Z(n2933) );
  ANDN U3403 ( .B(n2931), .A(n2933), .Z(n2940) );
  NOR U3404 ( .A(n2935), .B(n2934), .Z(n2932) );
  XNOR U3405 ( .A(n2933), .B(n2932), .Z(n2938) );
  XOR U3406 ( .A(n2935), .B(n2934), .Z(n2936) );
  NAND U3407 ( .A(n2936), .B(n5779), .Z(n2937) );
  NAND U3408 ( .A(n2938), .B(n2937), .Z(n5784) );
  XNOR U3409 ( .A(a[147]), .B(b[147]), .Z(n5783) );
  NAND U3410 ( .A(n5784), .B(n5783), .Z(n2939) );
  NANDN U3411 ( .A(n2940), .B(n2939), .Z(n2946) );
  NAND U3412 ( .A(a[147]), .B(b[147]), .Z(n2947) );
  AND U3413 ( .A(n2946), .B(n2947), .Z(n2942) );
  XOR U3414 ( .A(a[148]), .B(b[148]), .Z(n5789) );
  ANDN U3415 ( .B(n5788), .A(n5789), .Z(n2941) );
  OR U3416 ( .A(n2942), .B(n2941), .Z(n2943) );
  AND U3417 ( .A(a[148]), .B(b[148]), .Z(n2945) );
  ANDN U3418 ( .B(n2943), .A(n2945), .Z(n2952) );
  NOR U3419 ( .A(n2947), .B(n2946), .Z(n2944) );
  XNOR U3420 ( .A(n2945), .B(n2944), .Z(n2950) );
  XOR U3421 ( .A(n2947), .B(n2946), .Z(n2948) );
  NAND U3422 ( .A(n2948), .B(n5789), .Z(n2949) );
  NAND U3423 ( .A(n2950), .B(n2949), .Z(n5794) );
  XNOR U3424 ( .A(a[149]), .B(b[149]), .Z(n5793) );
  NAND U3425 ( .A(n5794), .B(n5793), .Z(n2951) );
  NANDN U3426 ( .A(n2952), .B(n2951), .Z(n2958) );
  NAND U3427 ( .A(a[149]), .B(b[149]), .Z(n2959) );
  AND U3428 ( .A(n2958), .B(n2959), .Z(n2954) );
  XOR U3429 ( .A(a[150]), .B(b[150]), .Z(n5799) );
  ANDN U3430 ( .B(n5798), .A(n5799), .Z(n2953) );
  OR U3431 ( .A(n2954), .B(n2953), .Z(n2955) );
  AND U3432 ( .A(a[150]), .B(b[150]), .Z(n2957) );
  ANDN U3433 ( .B(n2955), .A(n2957), .Z(n2964) );
  NOR U3434 ( .A(n2959), .B(n2958), .Z(n2956) );
  XNOR U3435 ( .A(n2957), .B(n2956), .Z(n2962) );
  XOR U3436 ( .A(n2959), .B(n2958), .Z(n2960) );
  NAND U3437 ( .A(n2960), .B(n5799), .Z(n2961) );
  NAND U3438 ( .A(n2962), .B(n2961), .Z(n5804) );
  XNOR U3439 ( .A(a[151]), .B(b[151]), .Z(n5803) );
  NAND U3440 ( .A(n5804), .B(n5803), .Z(n2963) );
  NANDN U3441 ( .A(n2964), .B(n2963), .Z(n2965) );
  IV U3442 ( .A(n2965), .Z(n2969) );
  AND U3443 ( .A(a[151]), .B(b[151]), .Z(n2970) );
  NOR U3444 ( .A(n2969), .B(n2970), .Z(n2967) );
  XNOR U3445 ( .A(n2970), .B(n2965), .Z(n5809) );
  XNOR U3446 ( .A(a[152]), .B(b[152]), .Z(n5808) );
  AND U3447 ( .A(n5809), .B(n5808), .Z(n2966) );
  OR U3448 ( .A(n2967), .B(n2966), .Z(n2968) );
  AND U3449 ( .A(a[152]), .B(b[152]), .Z(n2972) );
  ANDN U3450 ( .B(n2968), .A(n2972), .Z(n2974) );
  AND U3451 ( .A(n2970), .B(n2969), .Z(n2971) );
  NAND U3452 ( .A(n2972), .B(n2971), .Z(n2977) );
  ANDN U3453 ( .B(n2977), .A(n2974), .Z(n5814) );
  XNOR U3454 ( .A(a[153]), .B(b[153]), .Z(n5813) );
  AND U3455 ( .A(n5814), .B(n5813), .Z(n2973) );
  OR U3456 ( .A(n2974), .B(n2973), .Z(n2975) );
  AND U3457 ( .A(n2976), .B(n2975), .Z(n2980) );
  OR U3458 ( .A(n2977), .B(n2976), .Z(n2978) );
  ANDN U3459 ( .B(n2978), .A(n2980), .Z(n5819) );
  XNOR U3460 ( .A(a[154]), .B(b[154]), .Z(n5818) );
  NAND U3461 ( .A(n5819), .B(n5818), .Z(n2979) );
  NANDN U3462 ( .A(n2980), .B(n2979), .Z(n2986) );
  NAND U3463 ( .A(a[154]), .B(b[154]), .Z(n2987) );
  AND U3464 ( .A(n2986), .B(n2987), .Z(n2982) );
  XOR U3465 ( .A(a[155]), .B(b[155]), .Z(n5824) );
  ANDN U3466 ( .B(n5823), .A(n5824), .Z(n2981) );
  OR U3467 ( .A(n2982), .B(n2981), .Z(n2983) );
  AND U3468 ( .A(a[155]), .B(b[155]), .Z(n2985) );
  ANDN U3469 ( .B(n2983), .A(n2985), .Z(n2992) );
  NOR U3470 ( .A(n2987), .B(n2986), .Z(n2984) );
  XNOR U3471 ( .A(n2985), .B(n2984), .Z(n2990) );
  XOR U3472 ( .A(n2987), .B(n2986), .Z(n2988) );
  NAND U3473 ( .A(n2988), .B(n5824), .Z(n2989) );
  NAND U3474 ( .A(n2990), .B(n2989), .Z(n5829) );
  XNOR U3475 ( .A(a[156]), .B(b[156]), .Z(n5828) );
  NAND U3476 ( .A(n5829), .B(n5828), .Z(n2991) );
  NANDN U3477 ( .A(n2992), .B(n2991), .Z(n2993) );
  IV U3478 ( .A(n2993), .Z(n2997) );
  AND U3479 ( .A(a[156]), .B(b[156]), .Z(n2998) );
  NOR U3480 ( .A(n2997), .B(n2998), .Z(n2995) );
  XNOR U3481 ( .A(n2998), .B(n2993), .Z(n5834) );
  XNOR U3482 ( .A(a[157]), .B(b[157]), .Z(n5833) );
  AND U3483 ( .A(n5834), .B(n5833), .Z(n2994) );
  OR U3484 ( .A(n2995), .B(n2994), .Z(n2996) );
  AND U3485 ( .A(a[157]), .B(b[157]), .Z(n3000) );
  ANDN U3486 ( .B(n2996), .A(n3000), .Z(n3002) );
  AND U3487 ( .A(n2998), .B(n2997), .Z(n2999) );
  NAND U3488 ( .A(n3000), .B(n2999), .Z(n3005) );
  ANDN U3489 ( .B(n3005), .A(n3002), .Z(n5839) );
  XNOR U3490 ( .A(a[158]), .B(b[158]), .Z(n5838) );
  AND U3491 ( .A(n5839), .B(n5838), .Z(n3001) );
  OR U3492 ( .A(n3002), .B(n3001), .Z(n3003) );
  AND U3493 ( .A(a[158]), .B(b[158]), .Z(n3004) );
  ANDN U3494 ( .B(n3003), .A(n3004), .Z(n3008) );
  NANDN U3495 ( .A(n3005), .B(n3004), .Z(n3006) );
  ANDN U3496 ( .B(n3006), .A(n3008), .Z(n5844) );
  XNOR U3497 ( .A(a[159]), .B(b[159]), .Z(n5843) );
  NAND U3498 ( .A(n5844), .B(n5843), .Z(n3007) );
  NANDN U3499 ( .A(n3008), .B(n3007), .Z(n3014) );
  NAND U3500 ( .A(a[159]), .B(b[159]), .Z(n3015) );
  AND U3501 ( .A(n3014), .B(n3015), .Z(n3010) );
  XOR U3502 ( .A(a[160]), .B(b[160]), .Z(n5849) );
  ANDN U3503 ( .B(n5848), .A(n5849), .Z(n3009) );
  OR U3504 ( .A(n3010), .B(n3009), .Z(n3011) );
  AND U3505 ( .A(a[160]), .B(b[160]), .Z(n3013) );
  ANDN U3506 ( .B(n3011), .A(n3013), .Z(n3020) );
  NOR U3507 ( .A(n3015), .B(n3014), .Z(n3012) );
  XNOR U3508 ( .A(n3013), .B(n3012), .Z(n3018) );
  XOR U3509 ( .A(n3015), .B(n3014), .Z(n3016) );
  NAND U3510 ( .A(n3016), .B(n5849), .Z(n3017) );
  NAND U3511 ( .A(n3018), .B(n3017), .Z(n5854) );
  XNOR U3512 ( .A(a[161]), .B(b[161]), .Z(n5853) );
  NAND U3513 ( .A(n5854), .B(n5853), .Z(n3019) );
  NANDN U3514 ( .A(n3020), .B(n3019), .Z(n3026) );
  NAND U3515 ( .A(a[161]), .B(b[161]), .Z(n3027) );
  AND U3516 ( .A(n3026), .B(n3027), .Z(n3022) );
  XOR U3517 ( .A(a[162]), .B(b[162]), .Z(n5859) );
  ANDN U3518 ( .B(n5858), .A(n5859), .Z(n3021) );
  OR U3519 ( .A(n3022), .B(n3021), .Z(n3023) );
  AND U3520 ( .A(a[162]), .B(b[162]), .Z(n3025) );
  ANDN U3521 ( .B(n3023), .A(n3025), .Z(n3032) );
  NOR U3522 ( .A(n3027), .B(n3026), .Z(n3024) );
  XNOR U3523 ( .A(n3025), .B(n3024), .Z(n3030) );
  XOR U3524 ( .A(n3027), .B(n3026), .Z(n3028) );
  NAND U3525 ( .A(n3028), .B(n5859), .Z(n3029) );
  NAND U3526 ( .A(n3030), .B(n3029), .Z(n5864) );
  XNOR U3527 ( .A(a[163]), .B(b[163]), .Z(n5863) );
  NAND U3528 ( .A(n5864), .B(n5863), .Z(n3031) );
  NANDN U3529 ( .A(n3032), .B(n3031), .Z(n3037) );
  ANDN U3530 ( .B(n3036), .A(n3037), .Z(n3033) );
  XOR U3531 ( .A(n3038), .B(n3033), .Z(n3035) );
  XOR U3532 ( .A(a[164]), .B(b[164]), .Z(n5869) );
  XNOR U3533 ( .A(n3036), .B(n3037), .Z(n5868) );
  NAND U3534 ( .A(n5869), .B(n5868), .Z(n3034) );
  NAND U3535 ( .A(n3035), .B(n3034), .Z(n5874) );
  XNOR U3536 ( .A(a[165]), .B(b[165]), .Z(n5873) );
  IV U3537 ( .A(n3039), .Z(n3041) );
  XNOR U3538 ( .A(n3040), .B(n3039), .Z(n5879) );
  XNOR U3539 ( .A(a[166]), .B(b[166]), .Z(n5878) );
  AND U3540 ( .A(a[166]), .B(b[166]), .Z(n3043) );
  NOR U3541 ( .A(n3041), .B(n3040), .Z(n3042) );
  NAND U3542 ( .A(n3043), .B(n3042), .Z(n3048) );
  ANDN U3543 ( .B(n3048), .A(n3045), .Z(n5884) );
  XNOR U3544 ( .A(a[167]), .B(b[167]), .Z(n5883) );
  NAND U3545 ( .A(n5884), .B(n5883), .Z(n3044) );
  NANDN U3546 ( .A(n3045), .B(n3044), .Z(n3046) );
  AND U3547 ( .A(n3047), .B(n3046), .Z(n3051) );
  OR U3548 ( .A(n3048), .B(n3047), .Z(n3049) );
  ANDN U3549 ( .B(n3049), .A(n3051), .Z(n5889) );
  XNOR U3550 ( .A(a[168]), .B(b[168]), .Z(n5888) );
  NAND U3551 ( .A(n5889), .B(n5888), .Z(n3050) );
  NANDN U3552 ( .A(n3051), .B(n3050), .Z(n3057) );
  NAND U3553 ( .A(a[168]), .B(b[168]), .Z(n3058) );
  AND U3554 ( .A(n3057), .B(n3058), .Z(n3053) );
  XOR U3555 ( .A(a[169]), .B(b[169]), .Z(n5894) );
  ANDN U3556 ( .B(n5893), .A(n5894), .Z(n3052) );
  OR U3557 ( .A(n3053), .B(n3052), .Z(n3054) );
  AND U3558 ( .A(a[169]), .B(b[169]), .Z(n3056) );
  ANDN U3559 ( .B(n3054), .A(n3056), .Z(n3063) );
  NOR U3560 ( .A(n3058), .B(n3057), .Z(n3055) );
  XNOR U3561 ( .A(n3056), .B(n3055), .Z(n3061) );
  XOR U3562 ( .A(n3058), .B(n3057), .Z(n3059) );
  NAND U3563 ( .A(n3059), .B(n5894), .Z(n3060) );
  NAND U3564 ( .A(n3061), .B(n3060), .Z(n5899) );
  XNOR U3565 ( .A(a[170]), .B(b[170]), .Z(n5898) );
  NAND U3566 ( .A(n5899), .B(n5898), .Z(n3062) );
  NANDN U3567 ( .A(n3063), .B(n3062), .Z(n3069) );
  NAND U3568 ( .A(a[170]), .B(b[170]), .Z(n3070) );
  AND U3569 ( .A(n3069), .B(n3070), .Z(n3065) );
  XOR U3570 ( .A(a[171]), .B(b[171]), .Z(n5904) );
  ANDN U3571 ( .B(n5903), .A(n5904), .Z(n3064) );
  OR U3572 ( .A(n3065), .B(n3064), .Z(n3066) );
  AND U3573 ( .A(a[171]), .B(b[171]), .Z(n3068) );
  ANDN U3574 ( .B(n3066), .A(n3068), .Z(n3075) );
  NOR U3575 ( .A(n3070), .B(n3069), .Z(n3067) );
  XNOR U3576 ( .A(n3068), .B(n3067), .Z(n3073) );
  XOR U3577 ( .A(n3070), .B(n3069), .Z(n3071) );
  NAND U3578 ( .A(n3071), .B(n5904), .Z(n3072) );
  NAND U3579 ( .A(n3073), .B(n3072), .Z(n5909) );
  XNOR U3580 ( .A(a[172]), .B(b[172]), .Z(n5908) );
  NAND U3581 ( .A(n5909), .B(n5908), .Z(n3074) );
  NANDN U3582 ( .A(n3075), .B(n3074), .Z(n3081) );
  NAND U3583 ( .A(a[172]), .B(b[172]), .Z(n3082) );
  AND U3584 ( .A(n3081), .B(n3082), .Z(n3077) );
  XOR U3585 ( .A(a[173]), .B(b[173]), .Z(n5914) );
  ANDN U3586 ( .B(n5913), .A(n5914), .Z(n3076) );
  OR U3587 ( .A(n3077), .B(n3076), .Z(n3078) );
  AND U3588 ( .A(a[173]), .B(b[173]), .Z(n3080) );
  ANDN U3589 ( .B(n3078), .A(n3080), .Z(n3087) );
  NOR U3590 ( .A(n3082), .B(n3081), .Z(n3079) );
  XNOR U3591 ( .A(n3080), .B(n3079), .Z(n3085) );
  XOR U3592 ( .A(n3082), .B(n3081), .Z(n3083) );
  NAND U3593 ( .A(n3083), .B(n5914), .Z(n3084) );
  NAND U3594 ( .A(n3085), .B(n3084), .Z(n5919) );
  XNOR U3595 ( .A(a[174]), .B(b[174]), .Z(n5918) );
  NAND U3596 ( .A(n5919), .B(n5918), .Z(n3086) );
  NANDN U3597 ( .A(n3087), .B(n3086), .Z(n3093) );
  NAND U3598 ( .A(a[174]), .B(b[174]), .Z(n3094) );
  AND U3599 ( .A(n3093), .B(n3094), .Z(n3089) );
  XOR U3600 ( .A(a[175]), .B(b[175]), .Z(n5924) );
  ANDN U3601 ( .B(n5923), .A(n5924), .Z(n3088) );
  OR U3602 ( .A(n3089), .B(n3088), .Z(n3090) );
  AND U3603 ( .A(a[175]), .B(b[175]), .Z(n3092) );
  ANDN U3604 ( .B(n3090), .A(n3092), .Z(n3099) );
  NOR U3605 ( .A(n3094), .B(n3093), .Z(n3091) );
  XNOR U3606 ( .A(n3092), .B(n3091), .Z(n3097) );
  XOR U3607 ( .A(n3094), .B(n3093), .Z(n3095) );
  NAND U3608 ( .A(n3095), .B(n5924), .Z(n3096) );
  NAND U3609 ( .A(n3097), .B(n3096), .Z(n5929) );
  XNOR U3610 ( .A(a[176]), .B(b[176]), .Z(n5928) );
  NAND U3611 ( .A(n5929), .B(n5928), .Z(n3098) );
  NANDN U3612 ( .A(n3099), .B(n3098), .Z(n3105) );
  NAND U3613 ( .A(a[176]), .B(b[176]), .Z(n3106) );
  AND U3614 ( .A(n3105), .B(n3106), .Z(n3101) );
  XOR U3615 ( .A(a[177]), .B(b[177]), .Z(n5934) );
  ANDN U3616 ( .B(n5933), .A(n5934), .Z(n3100) );
  OR U3617 ( .A(n3101), .B(n3100), .Z(n3102) );
  AND U3618 ( .A(a[177]), .B(b[177]), .Z(n3104) );
  ANDN U3619 ( .B(n3102), .A(n3104), .Z(n3111) );
  NOR U3620 ( .A(n3106), .B(n3105), .Z(n3103) );
  XNOR U3621 ( .A(n3104), .B(n3103), .Z(n3109) );
  XOR U3622 ( .A(n3106), .B(n3105), .Z(n3107) );
  NAND U3623 ( .A(n3107), .B(n5934), .Z(n3108) );
  NAND U3624 ( .A(n3109), .B(n3108), .Z(n5939) );
  XNOR U3625 ( .A(a[178]), .B(b[178]), .Z(n5938) );
  NAND U3626 ( .A(n5939), .B(n5938), .Z(n3110) );
  NANDN U3627 ( .A(n3111), .B(n3110), .Z(n3117) );
  NAND U3628 ( .A(a[178]), .B(b[178]), .Z(n3118) );
  AND U3629 ( .A(n3117), .B(n3118), .Z(n3113) );
  XOR U3630 ( .A(a[179]), .B(b[179]), .Z(n5944) );
  ANDN U3631 ( .B(n5943), .A(n5944), .Z(n3112) );
  OR U3632 ( .A(n3113), .B(n3112), .Z(n3114) );
  AND U3633 ( .A(a[179]), .B(b[179]), .Z(n3116) );
  ANDN U3634 ( .B(n3114), .A(n3116), .Z(n3123) );
  NOR U3635 ( .A(n3118), .B(n3117), .Z(n3115) );
  XNOR U3636 ( .A(n3116), .B(n3115), .Z(n3121) );
  XOR U3637 ( .A(n3118), .B(n3117), .Z(n3119) );
  NAND U3638 ( .A(n3119), .B(n5944), .Z(n3120) );
  NAND U3639 ( .A(n3121), .B(n3120), .Z(n5949) );
  XNOR U3640 ( .A(a[180]), .B(b[180]), .Z(n5948) );
  NAND U3641 ( .A(n5949), .B(n5948), .Z(n3122) );
  NANDN U3642 ( .A(n3123), .B(n3122), .Z(n3129) );
  NAND U3643 ( .A(a[180]), .B(b[180]), .Z(n3130) );
  AND U3644 ( .A(n3129), .B(n3130), .Z(n3125) );
  XOR U3645 ( .A(a[181]), .B(b[181]), .Z(n5954) );
  ANDN U3646 ( .B(n5953), .A(n5954), .Z(n3124) );
  OR U3647 ( .A(n3125), .B(n3124), .Z(n3126) );
  AND U3648 ( .A(a[181]), .B(b[181]), .Z(n3128) );
  ANDN U3649 ( .B(n3126), .A(n3128), .Z(n3135) );
  NOR U3650 ( .A(n3130), .B(n3129), .Z(n3127) );
  XNOR U3651 ( .A(n3128), .B(n3127), .Z(n3133) );
  XOR U3652 ( .A(n3130), .B(n3129), .Z(n3131) );
  NAND U3653 ( .A(n3131), .B(n5954), .Z(n3132) );
  NAND U3654 ( .A(n3133), .B(n3132), .Z(n5959) );
  XNOR U3655 ( .A(a[182]), .B(b[182]), .Z(n5958) );
  NAND U3656 ( .A(n5959), .B(n5958), .Z(n3134) );
  NANDN U3657 ( .A(n3135), .B(n3134), .Z(n3141) );
  NAND U3658 ( .A(a[182]), .B(b[182]), .Z(n3142) );
  AND U3659 ( .A(n3141), .B(n3142), .Z(n3137) );
  XOR U3660 ( .A(a[183]), .B(b[183]), .Z(n5964) );
  ANDN U3661 ( .B(n5963), .A(n5964), .Z(n3136) );
  OR U3662 ( .A(n3137), .B(n3136), .Z(n3138) );
  AND U3663 ( .A(a[183]), .B(b[183]), .Z(n3140) );
  ANDN U3664 ( .B(n3138), .A(n3140), .Z(n3147) );
  NOR U3665 ( .A(n3142), .B(n3141), .Z(n3139) );
  XNOR U3666 ( .A(n3140), .B(n3139), .Z(n3145) );
  XOR U3667 ( .A(n3142), .B(n3141), .Z(n3143) );
  NAND U3668 ( .A(n3143), .B(n5964), .Z(n3144) );
  NAND U3669 ( .A(n3145), .B(n3144), .Z(n5969) );
  XNOR U3670 ( .A(a[184]), .B(b[184]), .Z(n5968) );
  NAND U3671 ( .A(n5969), .B(n5968), .Z(n3146) );
  NANDN U3672 ( .A(n3147), .B(n3146), .Z(n3148) );
  IV U3673 ( .A(n3148), .Z(n3152) );
  AND U3674 ( .A(a[184]), .B(b[184]), .Z(n3153) );
  NOR U3675 ( .A(n3152), .B(n3153), .Z(n3150) );
  XNOR U3676 ( .A(n3153), .B(n3148), .Z(n5974) );
  XNOR U3677 ( .A(a[185]), .B(b[185]), .Z(n5973) );
  AND U3678 ( .A(n5974), .B(n5973), .Z(n3149) );
  OR U3679 ( .A(n3150), .B(n3149), .Z(n3151) );
  AND U3680 ( .A(a[185]), .B(b[185]), .Z(n3155) );
  ANDN U3681 ( .B(n3151), .A(n3155), .Z(n3157) );
  AND U3682 ( .A(n3153), .B(n3152), .Z(n3154) );
  NAND U3683 ( .A(n3155), .B(n3154), .Z(n3160) );
  ANDN U3684 ( .B(n3160), .A(n3157), .Z(n5979) );
  XNOR U3685 ( .A(a[186]), .B(b[186]), .Z(n5978) );
  AND U3686 ( .A(n5979), .B(n5978), .Z(n3156) );
  OR U3687 ( .A(n3157), .B(n3156), .Z(n3158) );
  AND U3688 ( .A(n3159), .B(n3158), .Z(n3162) );
  XNOR U3689 ( .A(a[187]), .B(b[187]), .Z(n5983) );
  NAND U3690 ( .A(n5984), .B(n5983), .Z(n3161) );
  NANDN U3691 ( .A(n3162), .B(n3161), .Z(n3168) );
  NAND U3692 ( .A(a[187]), .B(b[187]), .Z(n3169) );
  AND U3693 ( .A(n3168), .B(n3169), .Z(n3164) );
  XOR U3694 ( .A(a[188]), .B(b[188]), .Z(n5989) );
  ANDN U3695 ( .B(n5988), .A(n5989), .Z(n3163) );
  OR U3696 ( .A(n3164), .B(n3163), .Z(n3165) );
  AND U3697 ( .A(a[188]), .B(b[188]), .Z(n3167) );
  ANDN U3698 ( .B(n3165), .A(n3167), .Z(n3174) );
  NOR U3699 ( .A(n3169), .B(n3168), .Z(n3166) );
  XNOR U3700 ( .A(n3167), .B(n3166), .Z(n3172) );
  XOR U3701 ( .A(n3169), .B(n3168), .Z(n3170) );
  NAND U3702 ( .A(n3170), .B(n5989), .Z(n3171) );
  NAND U3703 ( .A(n3172), .B(n3171), .Z(n5994) );
  XNOR U3704 ( .A(a[189]), .B(b[189]), .Z(n5993) );
  NAND U3705 ( .A(n5994), .B(n5993), .Z(n3173) );
  NANDN U3706 ( .A(n3174), .B(n3173), .Z(n3175) );
  IV U3707 ( .A(n3175), .Z(n3179) );
  AND U3708 ( .A(a[189]), .B(b[189]), .Z(n3180) );
  NOR U3709 ( .A(n3179), .B(n3180), .Z(n3177) );
  XNOR U3710 ( .A(n3180), .B(n3175), .Z(n5999) );
  XNOR U3711 ( .A(a[190]), .B(b[190]), .Z(n5998) );
  AND U3712 ( .A(n5999), .B(n5998), .Z(n3176) );
  OR U3713 ( .A(n3177), .B(n3176), .Z(n3178) );
  AND U3714 ( .A(a[190]), .B(b[190]), .Z(n3182) );
  ANDN U3715 ( .B(n3178), .A(n3182), .Z(n3184) );
  AND U3716 ( .A(n3180), .B(n3179), .Z(n3181) );
  NAND U3717 ( .A(n3182), .B(n3181), .Z(n3187) );
  ANDN U3718 ( .B(n3187), .A(n3184), .Z(n6004) );
  XNOR U3719 ( .A(a[191]), .B(b[191]), .Z(n6003) );
  AND U3720 ( .A(n6004), .B(n6003), .Z(n3183) );
  OR U3721 ( .A(n3184), .B(n3183), .Z(n3185) );
  AND U3722 ( .A(a[191]), .B(b[191]), .Z(n3186) );
  ANDN U3723 ( .B(n3185), .A(n3186), .Z(n3190) );
  NANDN U3724 ( .A(n3187), .B(n3186), .Z(n3188) );
  ANDN U3725 ( .B(n3188), .A(n3190), .Z(n6009) );
  XNOR U3726 ( .A(a[192]), .B(b[192]), .Z(n6008) );
  NAND U3727 ( .A(n6009), .B(n6008), .Z(n3189) );
  NANDN U3728 ( .A(n3190), .B(n3189), .Z(n3196) );
  NAND U3729 ( .A(a[192]), .B(b[192]), .Z(n3197) );
  AND U3730 ( .A(n3196), .B(n3197), .Z(n3192) );
  XOR U3731 ( .A(a[193]), .B(b[193]), .Z(n6014) );
  ANDN U3732 ( .B(n6013), .A(n6014), .Z(n3191) );
  OR U3733 ( .A(n3192), .B(n3191), .Z(n3193) );
  AND U3734 ( .A(a[193]), .B(b[193]), .Z(n3195) );
  ANDN U3735 ( .B(n3193), .A(n3195), .Z(n3202) );
  NOR U3736 ( .A(n3197), .B(n3196), .Z(n3194) );
  XNOR U3737 ( .A(n3195), .B(n3194), .Z(n3200) );
  XOR U3738 ( .A(n3197), .B(n3196), .Z(n3198) );
  NAND U3739 ( .A(n3198), .B(n6014), .Z(n3199) );
  NAND U3740 ( .A(n3200), .B(n3199), .Z(n6019) );
  XNOR U3741 ( .A(a[194]), .B(b[194]), .Z(n6018) );
  NAND U3742 ( .A(n6019), .B(n6018), .Z(n3201) );
  NANDN U3743 ( .A(n3202), .B(n3201), .Z(n3208) );
  NAND U3744 ( .A(a[194]), .B(b[194]), .Z(n3209) );
  AND U3745 ( .A(n3208), .B(n3209), .Z(n3204) );
  XOR U3746 ( .A(a[195]), .B(b[195]), .Z(n6024) );
  ANDN U3747 ( .B(n6023), .A(n6024), .Z(n3203) );
  OR U3748 ( .A(n3204), .B(n3203), .Z(n3205) );
  AND U3749 ( .A(a[195]), .B(b[195]), .Z(n3207) );
  ANDN U3750 ( .B(n3205), .A(n3207), .Z(n3214) );
  NOR U3751 ( .A(n3209), .B(n3208), .Z(n3206) );
  XNOR U3752 ( .A(n3207), .B(n3206), .Z(n3212) );
  XOR U3753 ( .A(n3209), .B(n3208), .Z(n3210) );
  NAND U3754 ( .A(n3210), .B(n6024), .Z(n3211) );
  NAND U3755 ( .A(n3212), .B(n3211), .Z(n6029) );
  XNOR U3756 ( .A(a[196]), .B(b[196]), .Z(n6028) );
  NAND U3757 ( .A(n6029), .B(n6028), .Z(n3213) );
  NANDN U3758 ( .A(n3214), .B(n3213), .Z(n3220) );
  NAND U3759 ( .A(a[196]), .B(b[196]), .Z(n3221) );
  AND U3760 ( .A(n3220), .B(n3221), .Z(n3216) );
  XOR U3761 ( .A(a[197]), .B(b[197]), .Z(n6034) );
  ANDN U3762 ( .B(n6033), .A(n6034), .Z(n3215) );
  OR U3763 ( .A(n3216), .B(n3215), .Z(n3217) );
  AND U3764 ( .A(a[197]), .B(b[197]), .Z(n3219) );
  ANDN U3765 ( .B(n3217), .A(n3219), .Z(n3226) );
  NOR U3766 ( .A(n3221), .B(n3220), .Z(n3218) );
  XNOR U3767 ( .A(n3219), .B(n3218), .Z(n3224) );
  XOR U3768 ( .A(n3221), .B(n3220), .Z(n3222) );
  NAND U3769 ( .A(n3222), .B(n6034), .Z(n3223) );
  NAND U3770 ( .A(n3224), .B(n3223), .Z(n6039) );
  XNOR U3771 ( .A(a[198]), .B(b[198]), .Z(n6038) );
  NAND U3772 ( .A(n6039), .B(n6038), .Z(n3225) );
  NANDN U3773 ( .A(n3226), .B(n3225), .Z(n3232) );
  NAND U3774 ( .A(a[198]), .B(b[198]), .Z(n3233) );
  AND U3775 ( .A(n3232), .B(n3233), .Z(n3228) );
  XOR U3776 ( .A(a[199]), .B(b[199]), .Z(n6044) );
  ANDN U3777 ( .B(n6043), .A(n6044), .Z(n3227) );
  OR U3778 ( .A(n3228), .B(n3227), .Z(n3229) );
  AND U3779 ( .A(a[199]), .B(b[199]), .Z(n3231) );
  ANDN U3780 ( .B(n3229), .A(n3231), .Z(n3238) );
  NOR U3781 ( .A(n3233), .B(n3232), .Z(n3230) );
  XNOR U3782 ( .A(n3231), .B(n3230), .Z(n3236) );
  XOR U3783 ( .A(n3233), .B(n3232), .Z(n3234) );
  NAND U3784 ( .A(n3234), .B(n6044), .Z(n3235) );
  NAND U3785 ( .A(n3236), .B(n3235), .Z(n6049) );
  XNOR U3786 ( .A(a[200]), .B(b[200]), .Z(n6048) );
  NAND U3787 ( .A(n6049), .B(n6048), .Z(n3237) );
  NANDN U3788 ( .A(n3238), .B(n3237), .Z(n3239) );
  IV U3789 ( .A(n3239), .Z(n3243) );
  AND U3790 ( .A(a[200]), .B(b[200]), .Z(n3244) );
  NOR U3791 ( .A(n3243), .B(n3244), .Z(n3241) );
  XNOR U3792 ( .A(n3244), .B(n3239), .Z(n6054) );
  XNOR U3793 ( .A(a[201]), .B(b[201]), .Z(n6053) );
  AND U3794 ( .A(n6054), .B(n6053), .Z(n3240) );
  OR U3795 ( .A(n3241), .B(n3240), .Z(n3242) );
  AND U3796 ( .A(a[201]), .B(b[201]), .Z(n3246) );
  ANDN U3797 ( .B(n3242), .A(n3246), .Z(n3248) );
  AND U3798 ( .A(n3244), .B(n3243), .Z(n3245) );
  NAND U3799 ( .A(n3246), .B(n3245), .Z(n3251) );
  ANDN U3800 ( .B(n3251), .A(n3248), .Z(n6059) );
  XNOR U3801 ( .A(a[202]), .B(b[202]), .Z(n6058) );
  AND U3802 ( .A(n6059), .B(n6058), .Z(n3247) );
  OR U3803 ( .A(n3248), .B(n3247), .Z(n3249) );
  AND U3804 ( .A(a[202]), .B(b[202]), .Z(n3250) );
  ANDN U3805 ( .B(n3249), .A(n3250), .Z(n3254) );
  NANDN U3806 ( .A(n3251), .B(n3250), .Z(n3252) );
  ANDN U3807 ( .B(n3252), .A(n3254), .Z(n6064) );
  XNOR U3808 ( .A(a[203]), .B(b[203]), .Z(n6063) );
  NAND U3809 ( .A(n6064), .B(n6063), .Z(n3253) );
  NANDN U3810 ( .A(n3254), .B(n3253), .Z(n3260) );
  NAND U3811 ( .A(a[203]), .B(b[203]), .Z(n3261) );
  AND U3812 ( .A(n3260), .B(n3261), .Z(n3256) );
  XOR U3813 ( .A(a[204]), .B(b[204]), .Z(n6069) );
  ANDN U3814 ( .B(n6068), .A(n6069), .Z(n3255) );
  OR U3815 ( .A(n3256), .B(n3255), .Z(n3257) );
  AND U3816 ( .A(a[204]), .B(b[204]), .Z(n3259) );
  ANDN U3817 ( .B(n3257), .A(n3259), .Z(n3266) );
  NOR U3818 ( .A(n3261), .B(n3260), .Z(n3258) );
  XNOR U3819 ( .A(n3259), .B(n3258), .Z(n3264) );
  XOR U3820 ( .A(n3261), .B(n3260), .Z(n3262) );
  NAND U3821 ( .A(n3262), .B(n6069), .Z(n3263) );
  NAND U3822 ( .A(n3264), .B(n3263), .Z(n6074) );
  XNOR U3823 ( .A(a[205]), .B(b[205]), .Z(n6073) );
  NAND U3824 ( .A(n6074), .B(n6073), .Z(n3265) );
  NANDN U3825 ( .A(n3266), .B(n3265), .Z(n3272) );
  NAND U3826 ( .A(a[205]), .B(b[205]), .Z(n3273) );
  AND U3827 ( .A(n3272), .B(n3273), .Z(n3268) );
  XOR U3828 ( .A(a[206]), .B(b[206]), .Z(n6079) );
  ANDN U3829 ( .B(n6078), .A(n6079), .Z(n3267) );
  OR U3830 ( .A(n3268), .B(n3267), .Z(n3269) );
  AND U3831 ( .A(a[206]), .B(b[206]), .Z(n3271) );
  ANDN U3832 ( .B(n3269), .A(n3271), .Z(n3278) );
  NOR U3833 ( .A(n3273), .B(n3272), .Z(n3270) );
  XNOR U3834 ( .A(n3271), .B(n3270), .Z(n3276) );
  XOR U3835 ( .A(n3273), .B(n3272), .Z(n3274) );
  NAND U3836 ( .A(n3274), .B(n6079), .Z(n3275) );
  NAND U3837 ( .A(n3276), .B(n3275), .Z(n6084) );
  XNOR U3838 ( .A(a[207]), .B(b[207]), .Z(n6083) );
  NAND U3839 ( .A(n6084), .B(n6083), .Z(n3277) );
  NANDN U3840 ( .A(n3278), .B(n3277), .Z(n3284) );
  NAND U3841 ( .A(a[207]), .B(b[207]), .Z(n3285) );
  AND U3842 ( .A(n3284), .B(n3285), .Z(n3280) );
  XOR U3843 ( .A(a[208]), .B(b[208]), .Z(n6089) );
  ANDN U3844 ( .B(n6088), .A(n6089), .Z(n3279) );
  OR U3845 ( .A(n3280), .B(n3279), .Z(n3281) );
  AND U3846 ( .A(a[208]), .B(b[208]), .Z(n3283) );
  ANDN U3847 ( .B(n3281), .A(n3283), .Z(n3290) );
  NOR U3848 ( .A(n3285), .B(n3284), .Z(n3282) );
  XNOR U3849 ( .A(n3283), .B(n3282), .Z(n3288) );
  XOR U3850 ( .A(n3285), .B(n3284), .Z(n3286) );
  NAND U3851 ( .A(n3286), .B(n6089), .Z(n3287) );
  NAND U3852 ( .A(n3288), .B(n3287), .Z(n6094) );
  XNOR U3853 ( .A(a[209]), .B(b[209]), .Z(n6093) );
  NAND U3854 ( .A(n6094), .B(n6093), .Z(n3289) );
  NANDN U3855 ( .A(n3290), .B(n3289), .Z(n3296) );
  NAND U3856 ( .A(a[209]), .B(b[209]), .Z(n3297) );
  AND U3857 ( .A(n3296), .B(n3297), .Z(n3292) );
  XOR U3858 ( .A(a[210]), .B(b[210]), .Z(n6099) );
  ANDN U3859 ( .B(n6098), .A(n6099), .Z(n3291) );
  OR U3860 ( .A(n3292), .B(n3291), .Z(n3293) );
  AND U3861 ( .A(a[210]), .B(b[210]), .Z(n3295) );
  ANDN U3862 ( .B(n3293), .A(n3295), .Z(n3302) );
  NOR U3863 ( .A(n3297), .B(n3296), .Z(n3294) );
  XNOR U3864 ( .A(n3295), .B(n3294), .Z(n3300) );
  XOR U3865 ( .A(n3297), .B(n3296), .Z(n3298) );
  NAND U3866 ( .A(n3298), .B(n6099), .Z(n3299) );
  NAND U3867 ( .A(n3300), .B(n3299), .Z(n6104) );
  XNOR U3868 ( .A(a[211]), .B(b[211]), .Z(n6103) );
  NAND U3869 ( .A(n6104), .B(n6103), .Z(n3301) );
  NANDN U3870 ( .A(n3302), .B(n3301), .Z(n3308) );
  NAND U3871 ( .A(a[211]), .B(b[211]), .Z(n3309) );
  AND U3872 ( .A(n3308), .B(n3309), .Z(n3304) );
  XOR U3873 ( .A(a[212]), .B(b[212]), .Z(n6109) );
  ANDN U3874 ( .B(n6108), .A(n6109), .Z(n3303) );
  OR U3875 ( .A(n3304), .B(n3303), .Z(n3305) );
  AND U3876 ( .A(a[212]), .B(b[212]), .Z(n3307) );
  ANDN U3877 ( .B(n3305), .A(n3307), .Z(n3314) );
  NOR U3878 ( .A(n3309), .B(n3308), .Z(n3306) );
  XNOR U3879 ( .A(n3307), .B(n3306), .Z(n3312) );
  XOR U3880 ( .A(n3309), .B(n3308), .Z(n3310) );
  NAND U3881 ( .A(n3310), .B(n6109), .Z(n3311) );
  NAND U3882 ( .A(n3312), .B(n3311), .Z(n6114) );
  XNOR U3883 ( .A(a[213]), .B(b[213]), .Z(n6113) );
  NAND U3884 ( .A(n6114), .B(n6113), .Z(n3313) );
  NANDN U3885 ( .A(n3314), .B(n3313), .Z(n3320) );
  NAND U3886 ( .A(a[213]), .B(b[213]), .Z(n3321) );
  AND U3887 ( .A(n3320), .B(n3321), .Z(n3316) );
  XOR U3888 ( .A(a[214]), .B(b[214]), .Z(n6119) );
  ANDN U3889 ( .B(n6118), .A(n6119), .Z(n3315) );
  OR U3890 ( .A(n3316), .B(n3315), .Z(n3317) );
  AND U3891 ( .A(a[214]), .B(b[214]), .Z(n3319) );
  ANDN U3892 ( .B(n3317), .A(n3319), .Z(n3326) );
  NOR U3893 ( .A(n3321), .B(n3320), .Z(n3318) );
  XNOR U3894 ( .A(n3319), .B(n3318), .Z(n3324) );
  XOR U3895 ( .A(n3321), .B(n3320), .Z(n3322) );
  NAND U3896 ( .A(n3322), .B(n6119), .Z(n3323) );
  NAND U3897 ( .A(n3324), .B(n3323), .Z(n6124) );
  XNOR U3898 ( .A(a[215]), .B(b[215]), .Z(n6123) );
  NAND U3899 ( .A(n6124), .B(n6123), .Z(n3325) );
  NANDN U3900 ( .A(n3326), .B(n3325), .Z(n3332) );
  NAND U3901 ( .A(a[215]), .B(b[215]), .Z(n3333) );
  AND U3902 ( .A(n3332), .B(n3333), .Z(n3328) );
  XOR U3903 ( .A(a[216]), .B(b[216]), .Z(n6129) );
  ANDN U3904 ( .B(n6128), .A(n6129), .Z(n3327) );
  OR U3905 ( .A(n3328), .B(n3327), .Z(n3329) );
  AND U3906 ( .A(a[216]), .B(b[216]), .Z(n3331) );
  ANDN U3907 ( .B(n3329), .A(n3331), .Z(n3338) );
  NOR U3908 ( .A(n3333), .B(n3332), .Z(n3330) );
  XNOR U3909 ( .A(n3331), .B(n3330), .Z(n3336) );
  XOR U3910 ( .A(n3333), .B(n3332), .Z(n3334) );
  NAND U3911 ( .A(n3334), .B(n6129), .Z(n3335) );
  NAND U3912 ( .A(n3336), .B(n3335), .Z(n6134) );
  XNOR U3913 ( .A(a[217]), .B(b[217]), .Z(n6133) );
  NAND U3914 ( .A(n6134), .B(n6133), .Z(n3337) );
  NANDN U3915 ( .A(n3338), .B(n3337), .Z(n3339) );
  IV U3916 ( .A(n3339), .Z(n3343) );
  AND U3917 ( .A(a[217]), .B(b[217]), .Z(n3344) );
  NOR U3918 ( .A(n3343), .B(n3344), .Z(n3341) );
  XNOR U3919 ( .A(n3344), .B(n3339), .Z(n6139) );
  XNOR U3920 ( .A(a[218]), .B(b[218]), .Z(n6138) );
  AND U3921 ( .A(n6139), .B(n6138), .Z(n3340) );
  OR U3922 ( .A(n3341), .B(n3340), .Z(n3342) );
  AND U3923 ( .A(a[218]), .B(b[218]), .Z(n3346) );
  ANDN U3924 ( .B(n3342), .A(n3346), .Z(n3348) );
  AND U3925 ( .A(n3344), .B(n3343), .Z(n3345) );
  NAND U3926 ( .A(n3346), .B(n3345), .Z(n3351) );
  ANDN U3927 ( .B(n3351), .A(n3348), .Z(n6144) );
  XNOR U3928 ( .A(a[219]), .B(b[219]), .Z(n6143) );
  AND U3929 ( .A(n6144), .B(n6143), .Z(n3347) );
  OR U3930 ( .A(n3348), .B(n3347), .Z(n3349) );
  AND U3931 ( .A(a[219]), .B(b[219]), .Z(n3350) );
  ANDN U3932 ( .B(n3349), .A(n3350), .Z(n3354) );
  NANDN U3933 ( .A(n3351), .B(n3350), .Z(n3352) );
  ANDN U3934 ( .B(n3352), .A(n3354), .Z(n6149) );
  XNOR U3935 ( .A(a[220]), .B(b[220]), .Z(n6148) );
  NAND U3936 ( .A(n6149), .B(n6148), .Z(n3353) );
  NANDN U3937 ( .A(n3354), .B(n3353), .Z(n3360) );
  NAND U3938 ( .A(a[220]), .B(b[220]), .Z(n3361) );
  AND U3939 ( .A(n3360), .B(n3361), .Z(n3356) );
  XOR U3940 ( .A(a[221]), .B(b[221]), .Z(n6154) );
  ANDN U3941 ( .B(n6153), .A(n6154), .Z(n3355) );
  OR U3942 ( .A(n3356), .B(n3355), .Z(n3357) );
  AND U3943 ( .A(a[221]), .B(b[221]), .Z(n3359) );
  ANDN U3944 ( .B(n3357), .A(n3359), .Z(n3366) );
  NOR U3945 ( .A(n3361), .B(n3360), .Z(n3358) );
  XNOR U3946 ( .A(n3359), .B(n3358), .Z(n3364) );
  XOR U3947 ( .A(n3361), .B(n3360), .Z(n3362) );
  NAND U3948 ( .A(n3362), .B(n6154), .Z(n3363) );
  NAND U3949 ( .A(n3364), .B(n3363), .Z(n6159) );
  XNOR U3950 ( .A(a[222]), .B(b[222]), .Z(n6158) );
  NAND U3951 ( .A(n6159), .B(n6158), .Z(n3365) );
  NANDN U3952 ( .A(n3366), .B(n3365), .Z(n3372) );
  NAND U3953 ( .A(a[222]), .B(b[222]), .Z(n3373) );
  AND U3954 ( .A(n3372), .B(n3373), .Z(n3368) );
  XOR U3955 ( .A(a[223]), .B(b[223]), .Z(n6164) );
  ANDN U3956 ( .B(n6163), .A(n6164), .Z(n3367) );
  OR U3957 ( .A(n3368), .B(n3367), .Z(n3369) );
  AND U3958 ( .A(a[223]), .B(b[223]), .Z(n3371) );
  ANDN U3959 ( .B(n3369), .A(n3371), .Z(n3378) );
  NOR U3960 ( .A(n3373), .B(n3372), .Z(n3370) );
  XNOR U3961 ( .A(n3371), .B(n3370), .Z(n3376) );
  XOR U3962 ( .A(n3373), .B(n3372), .Z(n3374) );
  NAND U3963 ( .A(n3374), .B(n6164), .Z(n3375) );
  NAND U3964 ( .A(n3376), .B(n3375), .Z(n6169) );
  XNOR U3965 ( .A(a[224]), .B(b[224]), .Z(n6168) );
  NAND U3966 ( .A(n6169), .B(n6168), .Z(n3377) );
  NANDN U3967 ( .A(n3378), .B(n3377), .Z(n3384) );
  NAND U3968 ( .A(a[224]), .B(b[224]), .Z(n3385) );
  AND U3969 ( .A(n3384), .B(n3385), .Z(n3380) );
  XOR U3970 ( .A(a[225]), .B(b[225]), .Z(n6174) );
  ANDN U3971 ( .B(n6173), .A(n6174), .Z(n3379) );
  OR U3972 ( .A(n3380), .B(n3379), .Z(n3381) );
  AND U3973 ( .A(a[225]), .B(b[225]), .Z(n3383) );
  ANDN U3974 ( .B(n3381), .A(n3383), .Z(n3390) );
  NOR U3975 ( .A(n3385), .B(n3384), .Z(n3382) );
  XNOR U3976 ( .A(n3383), .B(n3382), .Z(n3388) );
  XOR U3977 ( .A(n3385), .B(n3384), .Z(n3386) );
  NAND U3978 ( .A(n3386), .B(n6174), .Z(n3387) );
  NAND U3979 ( .A(n3388), .B(n3387), .Z(n6179) );
  XNOR U3980 ( .A(a[226]), .B(b[226]), .Z(n6178) );
  NAND U3981 ( .A(n6179), .B(n6178), .Z(n3389) );
  NANDN U3982 ( .A(n3390), .B(n3389), .Z(n3396) );
  NAND U3983 ( .A(a[226]), .B(b[226]), .Z(n3397) );
  AND U3984 ( .A(n3396), .B(n3397), .Z(n3392) );
  XOR U3985 ( .A(a[227]), .B(b[227]), .Z(n6184) );
  ANDN U3986 ( .B(n6183), .A(n6184), .Z(n3391) );
  OR U3987 ( .A(n3392), .B(n3391), .Z(n3393) );
  AND U3988 ( .A(a[227]), .B(b[227]), .Z(n3395) );
  ANDN U3989 ( .B(n3393), .A(n3395), .Z(n3402) );
  NOR U3990 ( .A(n3397), .B(n3396), .Z(n3394) );
  XNOR U3991 ( .A(n3395), .B(n3394), .Z(n3400) );
  XOR U3992 ( .A(n3397), .B(n3396), .Z(n3398) );
  NAND U3993 ( .A(n3398), .B(n6184), .Z(n3399) );
  NAND U3994 ( .A(n3400), .B(n3399), .Z(n6189) );
  XNOR U3995 ( .A(a[228]), .B(b[228]), .Z(n6188) );
  NAND U3996 ( .A(n6189), .B(n6188), .Z(n3401) );
  NANDN U3997 ( .A(n3402), .B(n3401), .Z(n3408) );
  NAND U3998 ( .A(a[228]), .B(b[228]), .Z(n3409) );
  AND U3999 ( .A(n3408), .B(n3409), .Z(n3404) );
  XOR U4000 ( .A(a[229]), .B(b[229]), .Z(n6194) );
  ANDN U4001 ( .B(n6193), .A(n6194), .Z(n3403) );
  OR U4002 ( .A(n3404), .B(n3403), .Z(n3405) );
  AND U4003 ( .A(a[229]), .B(b[229]), .Z(n3407) );
  ANDN U4004 ( .B(n3405), .A(n3407), .Z(n3414) );
  NOR U4005 ( .A(n3409), .B(n3408), .Z(n3406) );
  XNOR U4006 ( .A(n3407), .B(n3406), .Z(n3412) );
  XOR U4007 ( .A(n3409), .B(n3408), .Z(n3410) );
  NAND U4008 ( .A(n3410), .B(n6194), .Z(n3411) );
  NAND U4009 ( .A(n3412), .B(n3411), .Z(n6199) );
  XNOR U4010 ( .A(a[230]), .B(b[230]), .Z(n6198) );
  NAND U4011 ( .A(n6199), .B(n6198), .Z(n3413) );
  NANDN U4012 ( .A(n3414), .B(n3413), .Z(n3420) );
  NAND U4013 ( .A(a[230]), .B(b[230]), .Z(n3421) );
  AND U4014 ( .A(n3420), .B(n3421), .Z(n3416) );
  XOR U4015 ( .A(a[231]), .B(b[231]), .Z(n6204) );
  ANDN U4016 ( .B(n6203), .A(n6204), .Z(n3415) );
  OR U4017 ( .A(n3416), .B(n3415), .Z(n3417) );
  AND U4018 ( .A(a[231]), .B(b[231]), .Z(n3419) );
  ANDN U4019 ( .B(n3417), .A(n3419), .Z(n3426) );
  NOR U4020 ( .A(n3421), .B(n3420), .Z(n3418) );
  XNOR U4021 ( .A(n3419), .B(n3418), .Z(n3424) );
  XOR U4022 ( .A(n3421), .B(n3420), .Z(n3422) );
  NAND U4023 ( .A(n3422), .B(n6204), .Z(n3423) );
  NAND U4024 ( .A(n3424), .B(n3423), .Z(n6209) );
  XNOR U4025 ( .A(a[232]), .B(b[232]), .Z(n6208) );
  NAND U4026 ( .A(n6209), .B(n6208), .Z(n3425) );
  NANDN U4027 ( .A(n3426), .B(n3425), .Z(n3432) );
  NAND U4028 ( .A(a[232]), .B(b[232]), .Z(n3433) );
  AND U4029 ( .A(n3432), .B(n3433), .Z(n3428) );
  XOR U4030 ( .A(a[233]), .B(b[233]), .Z(n6214) );
  ANDN U4031 ( .B(n6213), .A(n6214), .Z(n3427) );
  OR U4032 ( .A(n3428), .B(n3427), .Z(n3429) );
  AND U4033 ( .A(a[233]), .B(b[233]), .Z(n3431) );
  ANDN U4034 ( .B(n3429), .A(n3431), .Z(n3438) );
  NOR U4035 ( .A(n3433), .B(n3432), .Z(n3430) );
  XNOR U4036 ( .A(n3431), .B(n3430), .Z(n3436) );
  XOR U4037 ( .A(n3433), .B(n3432), .Z(n3434) );
  NAND U4038 ( .A(n3434), .B(n6214), .Z(n3435) );
  NAND U4039 ( .A(n3436), .B(n3435), .Z(n6219) );
  XNOR U4040 ( .A(a[234]), .B(b[234]), .Z(n6218) );
  NAND U4041 ( .A(n6219), .B(n6218), .Z(n3437) );
  NANDN U4042 ( .A(n3438), .B(n3437), .Z(n3444) );
  NAND U4043 ( .A(a[234]), .B(b[234]), .Z(n3445) );
  AND U4044 ( .A(n3444), .B(n3445), .Z(n3440) );
  XOR U4045 ( .A(a[235]), .B(b[235]), .Z(n6224) );
  ANDN U4046 ( .B(n6223), .A(n6224), .Z(n3439) );
  OR U4047 ( .A(n3440), .B(n3439), .Z(n3441) );
  AND U4048 ( .A(a[235]), .B(b[235]), .Z(n3443) );
  ANDN U4049 ( .B(n3441), .A(n3443), .Z(n3450) );
  NOR U4050 ( .A(n3445), .B(n3444), .Z(n3442) );
  XNOR U4051 ( .A(n3443), .B(n3442), .Z(n3448) );
  XOR U4052 ( .A(n3445), .B(n3444), .Z(n3446) );
  NAND U4053 ( .A(n3446), .B(n6224), .Z(n3447) );
  NAND U4054 ( .A(n3448), .B(n3447), .Z(n6229) );
  XNOR U4055 ( .A(a[236]), .B(b[236]), .Z(n6228) );
  NAND U4056 ( .A(n6229), .B(n6228), .Z(n3449) );
  NANDN U4057 ( .A(n3450), .B(n3449), .Z(n3451) );
  IV U4058 ( .A(n3451), .Z(n3455) );
  AND U4059 ( .A(a[236]), .B(b[236]), .Z(n3456) );
  NOR U4060 ( .A(n3455), .B(n3456), .Z(n3453) );
  XNOR U4061 ( .A(n3456), .B(n3451), .Z(n6234) );
  XNOR U4062 ( .A(a[237]), .B(b[237]), .Z(n6233) );
  AND U4063 ( .A(n6234), .B(n6233), .Z(n3452) );
  OR U4064 ( .A(n3453), .B(n3452), .Z(n3454) );
  AND U4065 ( .A(a[237]), .B(b[237]), .Z(n3458) );
  ANDN U4066 ( .B(n3454), .A(n3458), .Z(n3460) );
  AND U4067 ( .A(n3456), .B(n3455), .Z(n3457) );
  NAND U4068 ( .A(n3458), .B(n3457), .Z(n3463) );
  ANDN U4069 ( .B(n3463), .A(n3460), .Z(n6239) );
  XNOR U4070 ( .A(a[238]), .B(b[238]), .Z(n6238) );
  AND U4071 ( .A(n6239), .B(n6238), .Z(n3459) );
  OR U4072 ( .A(n3460), .B(n3459), .Z(n3461) );
  AND U4073 ( .A(a[238]), .B(b[238]), .Z(n3462) );
  ANDN U4074 ( .B(n3461), .A(n3462), .Z(n3466) );
  NANDN U4075 ( .A(n3463), .B(n3462), .Z(n3464) );
  ANDN U4076 ( .B(n3464), .A(n3466), .Z(n6244) );
  XNOR U4077 ( .A(a[239]), .B(b[239]), .Z(n6243) );
  NAND U4078 ( .A(n6244), .B(n6243), .Z(n3465) );
  NANDN U4079 ( .A(n3466), .B(n3465), .Z(n3472) );
  NAND U4080 ( .A(a[239]), .B(b[239]), .Z(n3473) );
  AND U4081 ( .A(n3472), .B(n3473), .Z(n3468) );
  XOR U4082 ( .A(a[240]), .B(b[240]), .Z(n6249) );
  ANDN U4083 ( .B(n6248), .A(n6249), .Z(n3467) );
  OR U4084 ( .A(n3468), .B(n3467), .Z(n3469) );
  AND U4085 ( .A(a[240]), .B(b[240]), .Z(n3471) );
  ANDN U4086 ( .B(n3469), .A(n3471), .Z(n3478) );
  NOR U4087 ( .A(n3473), .B(n3472), .Z(n3470) );
  XNOR U4088 ( .A(n3471), .B(n3470), .Z(n3476) );
  XOR U4089 ( .A(n3473), .B(n3472), .Z(n3474) );
  NAND U4090 ( .A(n3474), .B(n6249), .Z(n3475) );
  NAND U4091 ( .A(n3476), .B(n3475), .Z(n6254) );
  XNOR U4092 ( .A(a[241]), .B(b[241]), .Z(n6253) );
  NAND U4093 ( .A(n6254), .B(n6253), .Z(n3477) );
  NANDN U4094 ( .A(n3478), .B(n3477), .Z(n3484) );
  NAND U4095 ( .A(a[241]), .B(b[241]), .Z(n3485) );
  AND U4096 ( .A(n3484), .B(n3485), .Z(n3480) );
  XOR U4097 ( .A(a[242]), .B(b[242]), .Z(n6259) );
  ANDN U4098 ( .B(n6258), .A(n6259), .Z(n3479) );
  OR U4099 ( .A(n3480), .B(n3479), .Z(n3481) );
  AND U4100 ( .A(a[242]), .B(b[242]), .Z(n3483) );
  ANDN U4101 ( .B(n3481), .A(n3483), .Z(n3490) );
  NOR U4102 ( .A(n3485), .B(n3484), .Z(n3482) );
  XNOR U4103 ( .A(n3483), .B(n3482), .Z(n3488) );
  XOR U4104 ( .A(n3485), .B(n3484), .Z(n3486) );
  NAND U4105 ( .A(n3486), .B(n6259), .Z(n3487) );
  NAND U4106 ( .A(n3488), .B(n3487), .Z(n6264) );
  XNOR U4107 ( .A(a[243]), .B(b[243]), .Z(n6263) );
  NAND U4108 ( .A(n6264), .B(n6263), .Z(n3489) );
  NANDN U4109 ( .A(n3490), .B(n3489), .Z(n3496) );
  NAND U4110 ( .A(a[243]), .B(b[243]), .Z(n3497) );
  AND U4111 ( .A(n3496), .B(n3497), .Z(n3492) );
  XOR U4112 ( .A(a[244]), .B(b[244]), .Z(n6269) );
  ANDN U4113 ( .B(n6268), .A(n6269), .Z(n3491) );
  OR U4114 ( .A(n3492), .B(n3491), .Z(n3493) );
  AND U4115 ( .A(a[244]), .B(b[244]), .Z(n3495) );
  ANDN U4116 ( .B(n3493), .A(n3495), .Z(n3502) );
  NOR U4117 ( .A(n3497), .B(n3496), .Z(n3494) );
  XNOR U4118 ( .A(n3495), .B(n3494), .Z(n3500) );
  XOR U4119 ( .A(n3497), .B(n3496), .Z(n3498) );
  NAND U4120 ( .A(n3498), .B(n6269), .Z(n3499) );
  NAND U4121 ( .A(n3500), .B(n3499), .Z(n6274) );
  XNOR U4122 ( .A(a[245]), .B(b[245]), .Z(n6273) );
  NAND U4123 ( .A(n6274), .B(n6273), .Z(n3501) );
  NANDN U4124 ( .A(n3502), .B(n3501), .Z(n3508) );
  NAND U4125 ( .A(a[245]), .B(b[245]), .Z(n3509) );
  AND U4126 ( .A(n3508), .B(n3509), .Z(n3504) );
  XOR U4127 ( .A(a[246]), .B(b[246]), .Z(n6279) );
  ANDN U4128 ( .B(n6278), .A(n6279), .Z(n3503) );
  OR U4129 ( .A(n3504), .B(n3503), .Z(n3505) );
  AND U4130 ( .A(a[246]), .B(b[246]), .Z(n3507) );
  ANDN U4131 ( .B(n3505), .A(n3507), .Z(n3514) );
  NOR U4132 ( .A(n3509), .B(n3508), .Z(n3506) );
  XNOR U4133 ( .A(n3507), .B(n3506), .Z(n3512) );
  XOR U4134 ( .A(n3509), .B(n3508), .Z(n3510) );
  NAND U4135 ( .A(n3510), .B(n6279), .Z(n3511) );
  NAND U4136 ( .A(n3512), .B(n3511), .Z(n6284) );
  XNOR U4137 ( .A(a[247]), .B(b[247]), .Z(n6283) );
  NAND U4138 ( .A(n6284), .B(n6283), .Z(n3513) );
  NANDN U4139 ( .A(n3514), .B(n3513), .Z(n3520) );
  NAND U4140 ( .A(a[247]), .B(b[247]), .Z(n3521) );
  AND U4141 ( .A(n3520), .B(n3521), .Z(n3516) );
  XOR U4142 ( .A(a[248]), .B(b[248]), .Z(n6289) );
  ANDN U4143 ( .B(n6288), .A(n6289), .Z(n3515) );
  OR U4144 ( .A(n3516), .B(n3515), .Z(n3517) );
  AND U4145 ( .A(a[248]), .B(b[248]), .Z(n3519) );
  ANDN U4146 ( .B(n3517), .A(n3519), .Z(n3526) );
  NOR U4147 ( .A(n3521), .B(n3520), .Z(n3518) );
  XNOR U4148 ( .A(n3519), .B(n3518), .Z(n3524) );
  XOR U4149 ( .A(n3521), .B(n3520), .Z(n3522) );
  NAND U4150 ( .A(n3522), .B(n6289), .Z(n3523) );
  NAND U4151 ( .A(n3524), .B(n3523), .Z(n6294) );
  XNOR U4152 ( .A(a[249]), .B(b[249]), .Z(n6293) );
  NAND U4153 ( .A(n6294), .B(n6293), .Z(n3525) );
  NANDN U4154 ( .A(n3526), .B(n3525), .Z(n3532) );
  NAND U4155 ( .A(a[249]), .B(b[249]), .Z(n3533) );
  AND U4156 ( .A(n3532), .B(n3533), .Z(n3528) );
  XOR U4157 ( .A(a[250]), .B(b[250]), .Z(n6299) );
  ANDN U4158 ( .B(n6298), .A(n6299), .Z(n3527) );
  OR U4159 ( .A(n3528), .B(n3527), .Z(n3529) );
  AND U4160 ( .A(a[250]), .B(b[250]), .Z(n3531) );
  ANDN U4161 ( .B(n3529), .A(n3531), .Z(n3538) );
  NOR U4162 ( .A(n3533), .B(n3532), .Z(n3530) );
  XNOR U4163 ( .A(n3531), .B(n3530), .Z(n3536) );
  XOR U4164 ( .A(n3533), .B(n3532), .Z(n3534) );
  NAND U4165 ( .A(n3534), .B(n6299), .Z(n3535) );
  NAND U4166 ( .A(n3536), .B(n3535), .Z(n6304) );
  XNOR U4167 ( .A(a[251]), .B(b[251]), .Z(n6303) );
  NAND U4168 ( .A(n6304), .B(n6303), .Z(n3537) );
  NANDN U4169 ( .A(n3538), .B(n3537), .Z(n3544) );
  NAND U4170 ( .A(a[251]), .B(b[251]), .Z(n3545) );
  AND U4171 ( .A(n3544), .B(n3545), .Z(n3540) );
  XOR U4172 ( .A(a[252]), .B(b[252]), .Z(n6309) );
  ANDN U4173 ( .B(n6308), .A(n6309), .Z(n3539) );
  OR U4174 ( .A(n3540), .B(n3539), .Z(n3541) );
  AND U4175 ( .A(a[252]), .B(b[252]), .Z(n3543) );
  ANDN U4176 ( .B(n3541), .A(n3543), .Z(n3550) );
  NOR U4177 ( .A(n3545), .B(n3544), .Z(n3542) );
  XNOR U4178 ( .A(n3543), .B(n3542), .Z(n3548) );
  XOR U4179 ( .A(n3545), .B(n3544), .Z(n3546) );
  NAND U4180 ( .A(n3546), .B(n6309), .Z(n3547) );
  NAND U4181 ( .A(n3548), .B(n3547), .Z(n6314) );
  XNOR U4182 ( .A(a[253]), .B(b[253]), .Z(n6313) );
  NAND U4183 ( .A(n6314), .B(n6313), .Z(n3549) );
  NANDN U4184 ( .A(n3550), .B(n3549), .Z(n3556) );
  NAND U4185 ( .A(a[253]), .B(b[253]), .Z(n3557) );
  AND U4186 ( .A(n3556), .B(n3557), .Z(n3552) );
  XOR U4187 ( .A(a[254]), .B(b[254]), .Z(n6319) );
  ANDN U4188 ( .B(n6318), .A(n6319), .Z(n3551) );
  OR U4189 ( .A(n3552), .B(n3551), .Z(n3553) );
  AND U4190 ( .A(a[254]), .B(b[254]), .Z(n3555) );
  ANDN U4191 ( .B(n3553), .A(n3555), .Z(n3562) );
  NOR U4192 ( .A(n3557), .B(n3556), .Z(n3554) );
  XNOR U4193 ( .A(n3555), .B(n3554), .Z(n3560) );
  XOR U4194 ( .A(n3557), .B(n3556), .Z(n3558) );
  NAND U4195 ( .A(n3558), .B(n6319), .Z(n3559) );
  NAND U4196 ( .A(n3560), .B(n3559), .Z(n6324) );
  XNOR U4197 ( .A(a[255]), .B(b[255]), .Z(n6323) );
  NAND U4198 ( .A(n6324), .B(n6323), .Z(n3561) );
  NANDN U4199 ( .A(n3562), .B(n3561), .Z(n3568) );
  NAND U4200 ( .A(a[255]), .B(b[255]), .Z(n3569) );
  AND U4201 ( .A(n3568), .B(n3569), .Z(n3564) );
  XOR U4202 ( .A(a[256]), .B(b[256]), .Z(n6329) );
  ANDN U4203 ( .B(n6328), .A(n6329), .Z(n3563) );
  OR U4204 ( .A(n3564), .B(n3563), .Z(n3565) );
  AND U4205 ( .A(a[256]), .B(b[256]), .Z(n3567) );
  ANDN U4206 ( .B(n3565), .A(n3567), .Z(n3574) );
  NOR U4207 ( .A(n3569), .B(n3568), .Z(n3566) );
  XNOR U4208 ( .A(n3567), .B(n3566), .Z(n3572) );
  XOR U4209 ( .A(n3569), .B(n3568), .Z(n3570) );
  NAND U4210 ( .A(n3570), .B(n6329), .Z(n3571) );
  NAND U4211 ( .A(n3572), .B(n3571), .Z(n6334) );
  XNOR U4212 ( .A(a[257]), .B(b[257]), .Z(n6333) );
  NAND U4213 ( .A(n6334), .B(n6333), .Z(n3573) );
  NANDN U4214 ( .A(n3574), .B(n3573), .Z(n3580) );
  NAND U4215 ( .A(a[257]), .B(b[257]), .Z(n3581) );
  AND U4216 ( .A(n3580), .B(n3581), .Z(n3576) );
  XOR U4217 ( .A(a[258]), .B(b[258]), .Z(n6339) );
  ANDN U4218 ( .B(n6338), .A(n6339), .Z(n3575) );
  OR U4219 ( .A(n3576), .B(n3575), .Z(n3577) );
  AND U4220 ( .A(a[258]), .B(b[258]), .Z(n3579) );
  ANDN U4221 ( .B(n3577), .A(n3579), .Z(n3586) );
  NOR U4222 ( .A(n3581), .B(n3580), .Z(n3578) );
  XNOR U4223 ( .A(n3579), .B(n3578), .Z(n3584) );
  XOR U4224 ( .A(n3581), .B(n3580), .Z(n3582) );
  NAND U4225 ( .A(n3582), .B(n6339), .Z(n3583) );
  NAND U4226 ( .A(n3584), .B(n3583), .Z(n6344) );
  XNOR U4227 ( .A(a[259]), .B(b[259]), .Z(n6343) );
  NAND U4228 ( .A(n6344), .B(n6343), .Z(n3585) );
  NANDN U4229 ( .A(n3586), .B(n3585), .Z(n3592) );
  NAND U4230 ( .A(a[259]), .B(b[259]), .Z(n3593) );
  AND U4231 ( .A(n3592), .B(n3593), .Z(n3588) );
  XOR U4232 ( .A(a[260]), .B(b[260]), .Z(n6349) );
  ANDN U4233 ( .B(n6348), .A(n6349), .Z(n3587) );
  OR U4234 ( .A(n3588), .B(n3587), .Z(n3589) );
  AND U4235 ( .A(a[260]), .B(b[260]), .Z(n3591) );
  ANDN U4236 ( .B(n3589), .A(n3591), .Z(n3598) );
  NOR U4237 ( .A(n3593), .B(n3592), .Z(n3590) );
  XNOR U4238 ( .A(n3591), .B(n3590), .Z(n3596) );
  XOR U4239 ( .A(n3593), .B(n3592), .Z(n3594) );
  NAND U4240 ( .A(n3594), .B(n6349), .Z(n3595) );
  NAND U4241 ( .A(n3596), .B(n3595), .Z(n6354) );
  XNOR U4242 ( .A(a[261]), .B(b[261]), .Z(n6353) );
  NAND U4243 ( .A(n6354), .B(n6353), .Z(n3597) );
  NANDN U4244 ( .A(n3598), .B(n3597), .Z(n3604) );
  NAND U4245 ( .A(a[261]), .B(b[261]), .Z(n3605) );
  AND U4246 ( .A(n3604), .B(n3605), .Z(n3600) );
  XOR U4247 ( .A(a[262]), .B(b[262]), .Z(n6359) );
  ANDN U4248 ( .B(n6358), .A(n6359), .Z(n3599) );
  OR U4249 ( .A(n3600), .B(n3599), .Z(n3601) );
  AND U4250 ( .A(a[262]), .B(b[262]), .Z(n3603) );
  ANDN U4251 ( .B(n3601), .A(n3603), .Z(n3610) );
  NOR U4252 ( .A(n3605), .B(n3604), .Z(n3602) );
  XNOR U4253 ( .A(n3603), .B(n3602), .Z(n3608) );
  XOR U4254 ( .A(n3605), .B(n3604), .Z(n3606) );
  NAND U4255 ( .A(n3606), .B(n6359), .Z(n3607) );
  NAND U4256 ( .A(n3608), .B(n3607), .Z(n6364) );
  XNOR U4257 ( .A(a[263]), .B(b[263]), .Z(n6363) );
  NAND U4258 ( .A(n6364), .B(n6363), .Z(n3609) );
  NANDN U4259 ( .A(n3610), .B(n3609), .Z(n3616) );
  NAND U4260 ( .A(a[263]), .B(b[263]), .Z(n3617) );
  AND U4261 ( .A(n3616), .B(n3617), .Z(n3612) );
  XOR U4262 ( .A(a[264]), .B(b[264]), .Z(n6369) );
  ANDN U4263 ( .B(n6368), .A(n6369), .Z(n3611) );
  OR U4264 ( .A(n3612), .B(n3611), .Z(n3613) );
  AND U4265 ( .A(a[264]), .B(b[264]), .Z(n3615) );
  ANDN U4266 ( .B(n3613), .A(n3615), .Z(n3622) );
  NOR U4267 ( .A(n3617), .B(n3616), .Z(n3614) );
  XNOR U4268 ( .A(n3615), .B(n3614), .Z(n3620) );
  XOR U4269 ( .A(n3617), .B(n3616), .Z(n3618) );
  NAND U4270 ( .A(n3618), .B(n6369), .Z(n3619) );
  NAND U4271 ( .A(n3620), .B(n3619), .Z(n6374) );
  XNOR U4272 ( .A(a[265]), .B(b[265]), .Z(n6373) );
  NAND U4273 ( .A(n6374), .B(n6373), .Z(n3621) );
  NANDN U4274 ( .A(n3622), .B(n3621), .Z(n3628) );
  NAND U4275 ( .A(a[265]), .B(b[265]), .Z(n3629) );
  AND U4276 ( .A(n3628), .B(n3629), .Z(n3624) );
  XOR U4277 ( .A(a[266]), .B(b[266]), .Z(n6379) );
  ANDN U4278 ( .B(n6378), .A(n6379), .Z(n3623) );
  OR U4279 ( .A(n3624), .B(n3623), .Z(n3625) );
  AND U4280 ( .A(a[266]), .B(b[266]), .Z(n3627) );
  ANDN U4281 ( .B(n3625), .A(n3627), .Z(n3634) );
  NOR U4282 ( .A(n3629), .B(n3628), .Z(n3626) );
  XNOR U4283 ( .A(n3627), .B(n3626), .Z(n3632) );
  XOR U4284 ( .A(n3629), .B(n3628), .Z(n3630) );
  NAND U4285 ( .A(n3630), .B(n6379), .Z(n3631) );
  NAND U4286 ( .A(n3632), .B(n3631), .Z(n6384) );
  XNOR U4287 ( .A(a[267]), .B(b[267]), .Z(n6383) );
  NAND U4288 ( .A(n6384), .B(n6383), .Z(n3633) );
  NANDN U4289 ( .A(n3634), .B(n3633), .Z(n3640) );
  NAND U4290 ( .A(a[267]), .B(b[267]), .Z(n3641) );
  AND U4291 ( .A(n3640), .B(n3641), .Z(n3636) );
  XOR U4292 ( .A(a[268]), .B(b[268]), .Z(n6389) );
  ANDN U4293 ( .B(n6388), .A(n6389), .Z(n3635) );
  OR U4294 ( .A(n3636), .B(n3635), .Z(n3637) );
  AND U4295 ( .A(a[268]), .B(b[268]), .Z(n3639) );
  ANDN U4296 ( .B(n3637), .A(n3639), .Z(n3646) );
  NOR U4297 ( .A(n3641), .B(n3640), .Z(n3638) );
  XNOR U4298 ( .A(n3639), .B(n3638), .Z(n3644) );
  XOR U4299 ( .A(n3641), .B(n3640), .Z(n3642) );
  NAND U4300 ( .A(n3642), .B(n6389), .Z(n3643) );
  NAND U4301 ( .A(n3644), .B(n3643), .Z(n6394) );
  XNOR U4302 ( .A(a[269]), .B(b[269]), .Z(n6393) );
  NAND U4303 ( .A(n6394), .B(n6393), .Z(n3645) );
  NANDN U4304 ( .A(n3646), .B(n3645), .Z(n3652) );
  NAND U4305 ( .A(a[269]), .B(b[269]), .Z(n3653) );
  AND U4306 ( .A(n3652), .B(n3653), .Z(n3648) );
  XOR U4307 ( .A(a[270]), .B(b[270]), .Z(n6399) );
  ANDN U4308 ( .B(n6398), .A(n6399), .Z(n3647) );
  OR U4309 ( .A(n3648), .B(n3647), .Z(n3649) );
  AND U4310 ( .A(a[270]), .B(b[270]), .Z(n3651) );
  ANDN U4311 ( .B(n3649), .A(n3651), .Z(n3658) );
  NOR U4312 ( .A(n3653), .B(n3652), .Z(n3650) );
  XNOR U4313 ( .A(n3651), .B(n3650), .Z(n3656) );
  XOR U4314 ( .A(n3653), .B(n3652), .Z(n3654) );
  NAND U4315 ( .A(n3654), .B(n6399), .Z(n3655) );
  NAND U4316 ( .A(n3656), .B(n3655), .Z(n6404) );
  XNOR U4317 ( .A(a[271]), .B(b[271]), .Z(n6403) );
  NAND U4318 ( .A(n6404), .B(n6403), .Z(n3657) );
  NANDN U4319 ( .A(n3658), .B(n3657), .Z(n3664) );
  NAND U4320 ( .A(a[271]), .B(b[271]), .Z(n3665) );
  AND U4321 ( .A(n3664), .B(n3665), .Z(n3660) );
  XOR U4322 ( .A(a[272]), .B(b[272]), .Z(n6409) );
  ANDN U4323 ( .B(n6408), .A(n6409), .Z(n3659) );
  OR U4324 ( .A(n3660), .B(n3659), .Z(n3661) );
  AND U4325 ( .A(a[272]), .B(b[272]), .Z(n3663) );
  ANDN U4326 ( .B(n3661), .A(n3663), .Z(n3670) );
  NOR U4327 ( .A(n3665), .B(n3664), .Z(n3662) );
  XNOR U4328 ( .A(n3663), .B(n3662), .Z(n3668) );
  XOR U4329 ( .A(n3665), .B(n3664), .Z(n3666) );
  NAND U4330 ( .A(n3666), .B(n6409), .Z(n3667) );
  NAND U4331 ( .A(n3668), .B(n3667), .Z(n6414) );
  XNOR U4332 ( .A(a[273]), .B(b[273]), .Z(n6413) );
  NAND U4333 ( .A(n6414), .B(n6413), .Z(n3669) );
  NANDN U4334 ( .A(n3670), .B(n3669), .Z(n3676) );
  NAND U4335 ( .A(a[273]), .B(b[273]), .Z(n3677) );
  AND U4336 ( .A(n3676), .B(n3677), .Z(n3672) );
  XOR U4337 ( .A(a[274]), .B(b[274]), .Z(n6419) );
  ANDN U4338 ( .B(n6418), .A(n6419), .Z(n3671) );
  OR U4339 ( .A(n3672), .B(n3671), .Z(n3673) );
  AND U4340 ( .A(a[274]), .B(b[274]), .Z(n3675) );
  ANDN U4341 ( .B(n3673), .A(n3675), .Z(n3682) );
  NOR U4342 ( .A(n3677), .B(n3676), .Z(n3674) );
  XNOR U4343 ( .A(n3675), .B(n3674), .Z(n3680) );
  XOR U4344 ( .A(n3677), .B(n3676), .Z(n3678) );
  NAND U4345 ( .A(n3678), .B(n6419), .Z(n3679) );
  NAND U4346 ( .A(n3680), .B(n3679), .Z(n6424) );
  XNOR U4347 ( .A(a[275]), .B(b[275]), .Z(n6423) );
  NAND U4348 ( .A(n6424), .B(n6423), .Z(n3681) );
  NANDN U4349 ( .A(n3682), .B(n3681), .Z(n3688) );
  NAND U4350 ( .A(a[275]), .B(b[275]), .Z(n3689) );
  AND U4351 ( .A(n3688), .B(n3689), .Z(n3684) );
  XOR U4352 ( .A(a[276]), .B(b[276]), .Z(n6429) );
  ANDN U4353 ( .B(n6428), .A(n6429), .Z(n3683) );
  OR U4354 ( .A(n3684), .B(n3683), .Z(n3685) );
  AND U4355 ( .A(a[276]), .B(b[276]), .Z(n3687) );
  ANDN U4356 ( .B(n3685), .A(n3687), .Z(n3694) );
  NOR U4357 ( .A(n3689), .B(n3688), .Z(n3686) );
  XNOR U4358 ( .A(n3687), .B(n3686), .Z(n3692) );
  XOR U4359 ( .A(n3689), .B(n3688), .Z(n3690) );
  NAND U4360 ( .A(n3690), .B(n6429), .Z(n3691) );
  NAND U4361 ( .A(n3692), .B(n3691), .Z(n6434) );
  XNOR U4362 ( .A(a[277]), .B(b[277]), .Z(n6433) );
  NAND U4363 ( .A(n6434), .B(n6433), .Z(n3693) );
  NANDN U4364 ( .A(n3694), .B(n3693), .Z(n3700) );
  NAND U4365 ( .A(a[277]), .B(b[277]), .Z(n3701) );
  AND U4366 ( .A(n3700), .B(n3701), .Z(n3696) );
  XOR U4367 ( .A(a[278]), .B(b[278]), .Z(n6439) );
  ANDN U4368 ( .B(n6438), .A(n6439), .Z(n3695) );
  OR U4369 ( .A(n3696), .B(n3695), .Z(n3697) );
  AND U4370 ( .A(a[278]), .B(b[278]), .Z(n3699) );
  ANDN U4371 ( .B(n3697), .A(n3699), .Z(n3706) );
  NOR U4372 ( .A(n3701), .B(n3700), .Z(n3698) );
  XNOR U4373 ( .A(n3699), .B(n3698), .Z(n3704) );
  XOR U4374 ( .A(n3701), .B(n3700), .Z(n3702) );
  NAND U4375 ( .A(n3702), .B(n6439), .Z(n3703) );
  NAND U4376 ( .A(n3704), .B(n3703), .Z(n6444) );
  XNOR U4377 ( .A(a[279]), .B(b[279]), .Z(n6443) );
  NAND U4378 ( .A(n6444), .B(n6443), .Z(n3705) );
  NANDN U4379 ( .A(n3706), .B(n3705), .Z(n3707) );
  IV U4380 ( .A(n3707), .Z(n3711) );
  AND U4381 ( .A(a[279]), .B(b[279]), .Z(n3712) );
  NOR U4382 ( .A(n3711), .B(n3712), .Z(n3709) );
  XNOR U4383 ( .A(n3712), .B(n3707), .Z(n6449) );
  XNOR U4384 ( .A(a[280]), .B(b[280]), .Z(n6448) );
  AND U4385 ( .A(n6449), .B(n6448), .Z(n3708) );
  OR U4386 ( .A(n3709), .B(n3708), .Z(n3710) );
  AND U4387 ( .A(a[280]), .B(b[280]), .Z(n3714) );
  ANDN U4388 ( .B(n3710), .A(n3714), .Z(n3716) );
  AND U4389 ( .A(n3712), .B(n3711), .Z(n3713) );
  NAND U4390 ( .A(n3714), .B(n3713), .Z(n3719) );
  ANDN U4391 ( .B(n3719), .A(n3716), .Z(n6454) );
  XNOR U4392 ( .A(a[281]), .B(b[281]), .Z(n6453) );
  AND U4393 ( .A(n6454), .B(n6453), .Z(n3715) );
  OR U4394 ( .A(n3716), .B(n3715), .Z(n3717) );
  AND U4395 ( .A(n3718), .B(n3717), .Z(n3722) );
  OR U4396 ( .A(n3719), .B(n3718), .Z(n3720) );
  ANDN U4397 ( .B(n3720), .A(n3722), .Z(n6459) );
  XNOR U4398 ( .A(a[282]), .B(b[282]), .Z(n6458) );
  NAND U4399 ( .A(n6459), .B(n6458), .Z(n3721) );
  NANDN U4400 ( .A(n3722), .B(n3721), .Z(n3728) );
  NAND U4401 ( .A(a[282]), .B(b[282]), .Z(n3729) );
  AND U4402 ( .A(n3728), .B(n3729), .Z(n3724) );
  XOR U4403 ( .A(a[283]), .B(b[283]), .Z(n6464) );
  ANDN U4404 ( .B(n6463), .A(n6464), .Z(n3723) );
  OR U4405 ( .A(n3724), .B(n3723), .Z(n3725) );
  AND U4406 ( .A(a[283]), .B(b[283]), .Z(n3727) );
  ANDN U4407 ( .B(n3725), .A(n3727), .Z(n3734) );
  NOR U4408 ( .A(n3729), .B(n3728), .Z(n3726) );
  XNOR U4409 ( .A(n3727), .B(n3726), .Z(n3732) );
  XOR U4410 ( .A(n3729), .B(n3728), .Z(n3730) );
  NAND U4411 ( .A(n3730), .B(n6464), .Z(n3731) );
  NAND U4412 ( .A(n3732), .B(n3731), .Z(n6469) );
  XNOR U4413 ( .A(a[284]), .B(b[284]), .Z(n6468) );
  NAND U4414 ( .A(n6469), .B(n6468), .Z(n3733) );
  NANDN U4415 ( .A(n3734), .B(n3733), .Z(n3735) );
  IV U4416 ( .A(n3735), .Z(n3739) );
  AND U4417 ( .A(a[284]), .B(b[284]), .Z(n3740) );
  NOR U4418 ( .A(n3739), .B(n3740), .Z(n3737) );
  XNOR U4419 ( .A(n3740), .B(n3735), .Z(n6474) );
  XNOR U4420 ( .A(a[285]), .B(b[285]), .Z(n6473) );
  AND U4421 ( .A(n6474), .B(n6473), .Z(n3736) );
  OR U4422 ( .A(n3737), .B(n3736), .Z(n3738) );
  AND U4423 ( .A(a[285]), .B(b[285]), .Z(n3742) );
  ANDN U4424 ( .B(n3738), .A(n3742), .Z(n3744) );
  AND U4425 ( .A(n3740), .B(n3739), .Z(n3741) );
  NAND U4426 ( .A(n3742), .B(n3741), .Z(n3747) );
  ANDN U4427 ( .B(n3747), .A(n3744), .Z(n6479) );
  XNOR U4428 ( .A(a[286]), .B(b[286]), .Z(n6478) );
  AND U4429 ( .A(n6479), .B(n6478), .Z(n3743) );
  OR U4430 ( .A(n3744), .B(n3743), .Z(n3745) );
  AND U4431 ( .A(a[286]), .B(b[286]), .Z(n3746) );
  ANDN U4432 ( .B(n3745), .A(n3746), .Z(n3750) );
  NANDN U4433 ( .A(n3747), .B(n3746), .Z(n3748) );
  ANDN U4434 ( .B(n3748), .A(n3750), .Z(n6484) );
  XNOR U4435 ( .A(a[287]), .B(b[287]), .Z(n6483) );
  NAND U4436 ( .A(n6484), .B(n6483), .Z(n3749) );
  NANDN U4437 ( .A(n3750), .B(n3749), .Z(n3756) );
  NAND U4438 ( .A(a[287]), .B(b[287]), .Z(n3757) );
  AND U4439 ( .A(n3756), .B(n3757), .Z(n3752) );
  XOR U4440 ( .A(a[288]), .B(b[288]), .Z(n6489) );
  ANDN U4441 ( .B(n6488), .A(n6489), .Z(n3751) );
  OR U4442 ( .A(n3752), .B(n3751), .Z(n3753) );
  AND U4443 ( .A(a[288]), .B(b[288]), .Z(n3755) );
  ANDN U4444 ( .B(n3753), .A(n3755), .Z(n3762) );
  NOR U4445 ( .A(n3757), .B(n3756), .Z(n3754) );
  XNOR U4446 ( .A(n3755), .B(n3754), .Z(n3760) );
  XOR U4447 ( .A(n3757), .B(n3756), .Z(n3758) );
  NAND U4448 ( .A(n3758), .B(n6489), .Z(n3759) );
  NAND U4449 ( .A(n3760), .B(n3759), .Z(n6494) );
  XNOR U4450 ( .A(a[289]), .B(b[289]), .Z(n6493) );
  NAND U4451 ( .A(n6494), .B(n6493), .Z(n3761) );
  NANDN U4452 ( .A(n3762), .B(n3761), .Z(n3768) );
  NAND U4453 ( .A(a[289]), .B(b[289]), .Z(n3769) );
  AND U4454 ( .A(n3768), .B(n3769), .Z(n3764) );
  XOR U4455 ( .A(a[290]), .B(b[290]), .Z(n6499) );
  ANDN U4456 ( .B(n6498), .A(n6499), .Z(n3763) );
  OR U4457 ( .A(n3764), .B(n3763), .Z(n3765) );
  AND U4458 ( .A(a[290]), .B(b[290]), .Z(n3767) );
  ANDN U4459 ( .B(n3765), .A(n3767), .Z(n3774) );
  NOR U4460 ( .A(n3769), .B(n3768), .Z(n3766) );
  XNOR U4461 ( .A(n3767), .B(n3766), .Z(n3772) );
  XOR U4462 ( .A(n3769), .B(n3768), .Z(n3770) );
  NAND U4463 ( .A(n3770), .B(n6499), .Z(n3771) );
  NAND U4464 ( .A(n3772), .B(n3771), .Z(n6504) );
  XNOR U4465 ( .A(a[291]), .B(b[291]), .Z(n6503) );
  NAND U4466 ( .A(n6504), .B(n6503), .Z(n3773) );
  NANDN U4467 ( .A(n3774), .B(n3773), .Z(n3779) );
  ANDN U4468 ( .B(n3778), .A(n3779), .Z(n3775) );
  XOR U4469 ( .A(n3780), .B(n3775), .Z(n3777) );
  XOR U4470 ( .A(a[292]), .B(b[292]), .Z(n6509) );
  XNOR U4471 ( .A(n3778), .B(n3779), .Z(n6508) );
  NAND U4472 ( .A(n6509), .B(n6508), .Z(n3776) );
  NAND U4473 ( .A(n3777), .B(n3776), .Z(n6514) );
  XNOR U4474 ( .A(a[293]), .B(b[293]), .Z(n6513) );
  IV U4475 ( .A(n3781), .Z(n3783) );
  XNOR U4476 ( .A(n3782), .B(n3781), .Z(n6519) );
  XNOR U4477 ( .A(a[294]), .B(b[294]), .Z(n6518) );
  AND U4478 ( .A(a[294]), .B(b[294]), .Z(n3785) );
  NOR U4479 ( .A(n3783), .B(n3782), .Z(n3784) );
  NAND U4480 ( .A(n3785), .B(n3784), .Z(n3790) );
  ANDN U4481 ( .B(n3790), .A(n3787), .Z(n6524) );
  XNOR U4482 ( .A(a[295]), .B(b[295]), .Z(n6523) );
  NAND U4483 ( .A(n6524), .B(n6523), .Z(n3786) );
  NANDN U4484 ( .A(n3787), .B(n3786), .Z(n3788) );
  AND U4485 ( .A(n3789), .B(n3788), .Z(n3793) );
  OR U4486 ( .A(n3790), .B(n3789), .Z(n3791) );
  ANDN U4487 ( .B(n3791), .A(n3793), .Z(n6529) );
  XNOR U4488 ( .A(a[296]), .B(b[296]), .Z(n6528) );
  NAND U4489 ( .A(n6529), .B(n6528), .Z(n3792) );
  NANDN U4490 ( .A(n3793), .B(n3792), .Z(n3799) );
  NAND U4491 ( .A(a[296]), .B(b[296]), .Z(n3800) );
  AND U4492 ( .A(n3799), .B(n3800), .Z(n3795) );
  XOR U4493 ( .A(a[297]), .B(b[297]), .Z(n6534) );
  ANDN U4494 ( .B(n6533), .A(n6534), .Z(n3794) );
  OR U4495 ( .A(n3795), .B(n3794), .Z(n3796) );
  AND U4496 ( .A(a[297]), .B(b[297]), .Z(n3798) );
  ANDN U4497 ( .B(n3796), .A(n3798), .Z(n3805) );
  NOR U4498 ( .A(n3800), .B(n3799), .Z(n3797) );
  XNOR U4499 ( .A(n3798), .B(n3797), .Z(n3803) );
  XOR U4500 ( .A(n3800), .B(n3799), .Z(n3801) );
  NAND U4501 ( .A(n3801), .B(n6534), .Z(n3802) );
  NAND U4502 ( .A(n3803), .B(n3802), .Z(n6539) );
  XNOR U4503 ( .A(a[298]), .B(b[298]), .Z(n6538) );
  NAND U4504 ( .A(n6539), .B(n6538), .Z(n3804) );
  NANDN U4505 ( .A(n3805), .B(n3804), .Z(n3811) );
  NAND U4506 ( .A(a[298]), .B(b[298]), .Z(n3812) );
  AND U4507 ( .A(n3811), .B(n3812), .Z(n3807) );
  XOR U4508 ( .A(a[299]), .B(b[299]), .Z(n6544) );
  ANDN U4509 ( .B(n6543), .A(n6544), .Z(n3806) );
  OR U4510 ( .A(n3807), .B(n3806), .Z(n3808) );
  AND U4511 ( .A(a[299]), .B(b[299]), .Z(n3810) );
  ANDN U4512 ( .B(n3808), .A(n3810), .Z(n3817) );
  NOR U4513 ( .A(n3812), .B(n3811), .Z(n3809) );
  XNOR U4514 ( .A(n3810), .B(n3809), .Z(n3815) );
  XOR U4515 ( .A(n3812), .B(n3811), .Z(n3813) );
  NAND U4516 ( .A(n3813), .B(n6544), .Z(n3814) );
  NAND U4517 ( .A(n3815), .B(n3814), .Z(n6549) );
  XNOR U4518 ( .A(a[300]), .B(b[300]), .Z(n6548) );
  NAND U4519 ( .A(n6549), .B(n6548), .Z(n3816) );
  NANDN U4520 ( .A(n3817), .B(n3816), .Z(n3823) );
  NAND U4521 ( .A(a[300]), .B(b[300]), .Z(n3824) );
  AND U4522 ( .A(n3823), .B(n3824), .Z(n3819) );
  XOR U4523 ( .A(a[301]), .B(b[301]), .Z(n6554) );
  ANDN U4524 ( .B(n6553), .A(n6554), .Z(n3818) );
  OR U4525 ( .A(n3819), .B(n3818), .Z(n3820) );
  AND U4526 ( .A(a[301]), .B(b[301]), .Z(n3822) );
  ANDN U4527 ( .B(n3820), .A(n3822), .Z(n3829) );
  NOR U4528 ( .A(n3824), .B(n3823), .Z(n3821) );
  XNOR U4529 ( .A(n3822), .B(n3821), .Z(n3827) );
  XOR U4530 ( .A(n3824), .B(n3823), .Z(n3825) );
  NAND U4531 ( .A(n3825), .B(n6554), .Z(n3826) );
  NAND U4532 ( .A(n3827), .B(n3826), .Z(n6559) );
  XNOR U4533 ( .A(a[302]), .B(b[302]), .Z(n6558) );
  NAND U4534 ( .A(n6559), .B(n6558), .Z(n3828) );
  NANDN U4535 ( .A(n3829), .B(n3828), .Z(n3835) );
  NAND U4536 ( .A(a[302]), .B(b[302]), .Z(n3836) );
  AND U4537 ( .A(n3835), .B(n3836), .Z(n3831) );
  XOR U4538 ( .A(a[303]), .B(b[303]), .Z(n6564) );
  ANDN U4539 ( .B(n6563), .A(n6564), .Z(n3830) );
  OR U4540 ( .A(n3831), .B(n3830), .Z(n3832) );
  AND U4541 ( .A(a[303]), .B(b[303]), .Z(n3834) );
  ANDN U4542 ( .B(n3832), .A(n3834), .Z(n3841) );
  NOR U4543 ( .A(n3836), .B(n3835), .Z(n3833) );
  XNOR U4544 ( .A(n3834), .B(n3833), .Z(n3839) );
  XOR U4545 ( .A(n3836), .B(n3835), .Z(n3837) );
  NAND U4546 ( .A(n3837), .B(n6564), .Z(n3838) );
  NAND U4547 ( .A(n3839), .B(n3838), .Z(n6569) );
  XNOR U4548 ( .A(a[304]), .B(b[304]), .Z(n6568) );
  NAND U4549 ( .A(n6569), .B(n6568), .Z(n3840) );
  NANDN U4550 ( .A(n3841), .B(n3840), .Z(n3847) );
  NAND U4551 ( .A(a[304]), .B(b[304]), .Z(n3848) );
  AND U4552 ( .A(n3847), .B(n3848), .Z(n3843) );
  XOR U4553 ( .A(a[305]), .B(b[305]), .Z(n6574) );
  ANDN U4554 ( .B(n6573), .A(n6574), .Z(n3842) );
  OR U4555 ( .A(n3843), .B(n3842), .Z(n3844) );
  AND U4556 ( .A(a[305]), .B(b[305]), .Z(n3846) );
  ANDN U4557 ( .B(n3844), .A(n3846), .Z(n3853) );
  NOR U4558 ( .A(n3848), .B(n3847), .Z(n3845) );
  XNOR U4559 ( .A(n3846), .B(n3845), .Z(n3851) );
  XOR U4560 ( .A(n3848), .B(n3847), .Z(n3849) );
  NAND U4561 ( .A(n3849), .B(n6574), .Z(n3850) );
  NAND U4562 ( .A(n3851), .B(n3850), .Z(n6579) );
  XNOR U4563 ( .A(a[306]), .B(b[306]), .Z(n6578) );
  NAND U4564 ( .A(n6579), .B(n6578), .Z(n3852) );
  NANDN U4565 ( .A(n3853), .B(n3852), .Z(n3859) );
  NAND U4566 ( .A(a[306]), .B(b[306]), .Z(n3860) );
  AND U4567 ( .A(n3859), .B(n3860), .Z(n3855) );
  XOR U4568 ( .A(a[307]), .B(b[307]), .Z(n6584) );
  ANDN U4569 ( .B(n6583), .A(n6584), .Z(n3854) );
  OR U4570 ( .A(n3855), .B(n3854), .Z(n3856) );
  AND U4571 ( .A(a[307]), .B(b[307]), .Z(n3858) );
  ANDN U4572 ( .B(n3856), .A(n3858), .Z(n3865) );
  NOR U4573 ( .A(n3860), .B(n3859), .Z(n3857) );
  XNOR U4574 ( .A(n3858), .B(n3857), .Z(n3863) );
  XOR U4575 ( .A(n3860), .B(n3859), .Z(n3861) );
  NAND U4576 ( .A(n3861), .B(n6584), .Z(n3862) );
  NAND U4577 ( .A(n3863), .B(n3862), .Z(n6589) );
  XNOR U4578 ( .A(a[308]), .B(b[308]), .Z(n6588) );
  NAND U4579 ( .A(n6589), .B(n6588), .Z(n3864) );
  NANDN U4580 ( .A(n3865), .B(n3864), .Z(n3871) );
  NAND U4581 ( .A(a[308]), .B(b[308]), .Z(n3872) );
  AND U4582 ( .A(n3871), .B(n3872), .Z(n3867) );
  XOR U4583 ( .A(a[309]), .B(b[309]), .Z(n6594) );
  ANDN U4584 ( .B(n6593), .A(n6594), .Z(n3866) );
  OR U4585 ( .A(n3867), .B(n3866), .Z(n3868) );
  AND U4586 ( .A(a[309]), .B(b[309]), .Z(n3870) );
  ANDN U4587 ( .B(n3868), .A(n3870), .Z(n3877) );
  NOR U4588 ( .A(n3872), .B(n3871), .Z(n3869) );
  XNOR U4589 ( .A(n3870), .B(n3869), .Z(n3875) );
  XOR U4590 ( .A(n3872), .B(n3871), .Z(n3873) );
  NAND U4591 ( .A(n3873), .B(n6594), .Z(n3874) );
  NAND U4592 ( .A(n3875), .B(n3874), .Z(n6599) );
  XNOR U4593 ( .A(a[310]), .B(b[310]), .Z(n6598) );
  NAND U4594 ( .A(n6599), .B(n6598), .Z(n3876) );
  NANDN U4595 ( .A(n3877), .B(n3876), .Z(n3883) );
  NAND U4596 ( .A(a[310]), .B(b[310]), .Z(n3884) );
  AND U4597 ( .A(n3883), .B(n3884), .Z(n3879) );
  XOR U4598 ( .A(a[311]), .B(b[311]), .Z(n6604) );
  ANDN U4599 ( .B(n6603), .A(n6604), .Z(n3878) );
  OR U4600 ( .A(n3879), .B(n3878), .Z(n3880) );
  AND U4601 ( .A(a[311]), .B(b[311]), .Z(n3882) );
  ANDN U4602 ( .B(n3880), .A(n3882), .Z(n3889) );
  NOR U4603 ( .A(n3884), .B(n3883), .Z(n3881) );
  XNOR U4604 ( .A(n3882), .B(n3881), .Z(n3887) );
  XOR U4605 ( .A(n3884), .B(n3883), .Z(n3885) );
  NAND U4606 ( .A(n3885), .B(n6604), .Z(n3886) );
  NAND U4607 ( .A(n3887), .B(n3886), .Z(n6609) );
  XNOR U4608 ( .A(a[312]), .B(b[312]), .Z(n6608) );
  NAND U4609 ( .A(n6609), .B(n6608), .Z(n3888) );
  NANDN U4610 ( .A(n3889), .B(n3888), .Z(n3890) );
  IV U4611 ( .A(n3890), .Z(n3894) );
  AND U4612 ( .A(a[312]), .B(b[312]), .Z(n3895) );
  NOR U4613 ( .A(n3894), .B(n3895), .Z(n3892) );
  XNOR U4614 ( .A(n3895), .B(n3890), .Z(n6614) );
  XNOR U4615 ( .A(a[313]), .B(b[313]), .Z(n6613) );
  AND U4616 ( .A(n6614), .B(n6613), .Z(n3891) );
  OR U4617 ( .A(n3892), .B(n3891), .Z(n3893) );
  AND U4618 ( .A(a[313]), .B(b[313]), .Z(n3897) );
  ANDN U4619 ( .B(n3893), .A(n3897), .Z(n3899) );
  AND U4620 ( .A(n3895), .B(n3894), .Z(n3896) );
  NAND U4621 ( .A(n3897), .B(n3896), .Z(n3902) );
  ANDN U4622 ( .B(n3902), .A(n3899), .Z(n6619) );
  XNOR U4623 ( .A(a[314]), .B(b[314]), .Z(n6618) );
  AND U4624 ( .A(n6619), .B(n6618), .Z(n3898) );
  OR U4625 ( .A(n3899), .B(n3898), .Z(n3900) );
  AND U4626 ( .A(n3901), .B(n3900), .Z(n3904) );
  XNOR U4627 ( .A(a[315]), .B(b[315]), .Z(n6623) );
  NAND U4628 ( .A(n6624), .B(n6623), .Z(n3903) );
  NANDN U4629 ( .A(n3904), .B(n3903), .Z(n3910) );
  NAND U4630 ( .A(a[315]), .B(b[315]), .Z(n3911) );
  AND U4631 ( .A(n3910), .B(n3911), .Z(n3906) );
  XOR U4632 ( .A(a[316]), .B(b[316]), .Z(n6629) );
  ANDN U4633 ( .B(n6628), .A(n6629), .Z(n3905) );
  OR U4634 ( .A(n3906), .B(n3905), .Z(n3907) );
  AND U4635 ( .A(a[316]), .B(b[316]), .Z(n3909) );
  ANDN U4636 ( .B(n3907), .A(n3909), .Z(n3916) );
  NOR U4637 ( .A(n3911), .B(n3910), .Z(n3908) );
  XNOR U4638 ( .A(n3909), .B(n3908), .Z(n3914) );
  XOR U4639 ( .A(n3911), .B(n3910), .Z(n3912) );
  NAND U4640 ( .A(n3912), .B(n6629), .Z(n3913) );
  NAND U4641 ( .A(n3914), .B(n3913), .Z(n6634) );
  XNOR U4642 ( .A(a[317]), .B(b[317]), .Z(n6633) );
  NAND U4643 ( .A(n6634), .B(n6633), .Z(n3915) );
  NANDN U4644 ( .A(n3916), .B(n3915), .Z(n3917) );
  IV U4645 ( .A(n3917), .Z(n3921) );
  AND U4646 ( .A(a[317]), .B(b[317]), .Z(n3922) );
  NOR U4647 ( .A(n3921), .B(n3922), .Z(n3919) );
  XNOR U4648 ( .A(n3922), .B(n3917), .Z(n6639) );
  XNOR U4649 ( .A(a[318]), .B(b[318]), .Z(n6638) );
  AND U4650 ( .A(n6639), .B(n6638), .Z(n3918) );
  OR U4651 ( .A(n3919), .B(n3918), .Z(n3920) );
  AND U4652 ( .A(a[318]), .B(b[318]), .Z(n3924) );
  ANDN U4653 ( .B(n3920), .A(n3924), .Z(n3926) );
  AND U4654 ( .A(n3922), .B(n3921), .Z(n3923) );
  NAND U4655 ( .A(n3924), .B(n3923), .Z(n3929) );
  ANDN U4656 ( .B(n3929), .A(n3926), .Z(n6644) );
  XNOR U4657 ( .A(a[319]), .B(b[319]), .Z(n6643) );
  AND U4658 ( .A(n6644), .B(n6643), .Z(n3925) );
  OR U4659 ( .A(n3926), .B(n3925), .Z(n3927) );
  AND U4660 ( .A(a[319]), .B(b[319]), .Z(n3928) );
  ANDN U4661 ( .B(n3927), .A(n3928), .Z(n3932) );
  NANDN U4662 ( .A(n3929), .B(n3928), .Z(n3930) );
  ANDN U4663 ( .B(n3930), .A(n3932), .Z(n6649) );
  XNOR U4664 ( .A(a[320]), .B(b[320]), .Z(n6648) );
  NAND U4665 ( .A(n6649), .B(n6648), .Z(n3931) );
  NANDN U4666 ( .A(n3932), .B(n3931), .Z(n3938) );
  NAND U4667 ( .A(a[320]), .B(b[320]), .Z(n3939) );
  AND U4668 ( .A(n3938), .B(n3939), .Z(n3934) );
  XOR U4669 ( .A(a[321]), .B(b[321]), .Z(n6654) );
  ANDN U4670 ( .B(n6653), .A(n6654), .Z(n3933) );
  OR U4671 ( .A(n3934), .B(n3933), .Z(n3935) );
  AND U4672 ( .A(a[321]), .B(b[321]), .Z(n3937) );
  ANDN U4673 ( .B(n3935), .A(n3937), .Z(n3944) );
  NOR U4674 ( .A(n3939), .B(n3938), .Z(n3936) );
  XNOR U4675 ( .A(n3937), .B(n3936), .Z(n3942) );
  XOR U4676 ( .A(n3939), .B(n3938), .Z(n3940) );
  NAND U4677 ( .A(n3940), .B(n6654), .Z(n3941) );
  NAND U4678 ( .A(n3942), .B(n3941), .Z(n6659) );
  XNOR U4679 ( .A(a[322]), .B(b[322]), .Z(n6658) );
  NAND U4680 ( .A(n6659), .B(n6658), .Z(n3943) );
  NANDN U4681 ( .A(n3944), .B(n3943), .Z(n3950) );
  NAND U4682 ( .A(a[322]), .B(b[322]), .Z(n3951) );
  AND U4683 ( .A(n3950), .B(n3951), .Z(n3946) );
  XOR U4684 ( .A(a[323]), .B(b[323]), .Z(n6664) );
  ANDN U4685 ( .B(n6663), .A(n6664), .Z(n3945) );
  OR U4686 ( .A(n3946), .B(n3945), .Z(n3947) );
  AND U4687 ( .A(a[323]), .B(b[323]), .Z(n3949) );
  ANDN U4688 ( .B(n3947), .A(n3949), .Z(n3956) );
  NOR U4689 ( .A(n3951), .B(n3950), .Z(n3948) );
  XNOR U4690 ( .A(n3949), .B(n3948), .Z(n3954) );
  XOR U4691 ( .A(n3951), .B(n3950), .Z(n3952) );
  NAND U4692 ( .A(n3952), .B(n6664), .Z(n3953) );
  NAND U4693 ( .A(n3954), .B(n3953), .Z(n6669) );
  XNOR U4694 ( .A(a[324]), .B(b[324]), .Z(n6668) );
  NAND U4695 ( .A(n6669), .B(n6668), .Z(n3955) );
  NANDN U4696 ( .A(n3956), .B(n3955), .Z(n3962) );
  NAND U4697 ( .A(a[324]), .B(b[324]), .Z(n3963) );
  AND U4698 ( .A(n3962), .B(n3963), .Z(n3958) );
  XOR U4699 ( .A(a[325]), .B(b[325]), .Z(n6674) );
  ANDN U4700 ( .B(n6673), .A(n6674), .Z(n3957) );
  OR U4701 ( .A(n3958), .B(n3957), .Z(n3959) );
  AND U4702 ( .A(a[325]), .B(b[325]), .Z(n3961) );
  ANDN U4703 ( .B(n3959), .A(n3961), .Z(n3968) );
  NOR U4704 ( .A(n3963), .B(n3962), .Z(n3960) );
  XNOR U4705 ( .A(n3961), .B(n3960), .Z(n3966) );
  XOR U4706 ( .A(n3963), .B(n3962), .Z(n3964) );
  NAND U4707 ( .A(n3964), .B(n6674), .Z(n3965) );
  NAND U4708 ( .A(n3966), .B(n3965), .Z(n6679) );
  XNOR U4709 ( .A(a[326]), .B(b[326]), .Z(n6678) );
  NAND U4710 ( .A(n6679), .B(n6678), .Z(n3967) );
  NANDN U4711 ( .A(n3968), .B(n3967), .Z(n3974) );
  NAND U4712 ( .A(a[326]), .B(b[326]), .Z(n3975) );
  AND U4713 ( .A(n3974), .B(n3975), .Z(n3970) );
  XOR U4714 ( .A(a[327]), .B(b[327]), .Z(n6684) );
  ANDN U4715 ( .B(n6683), .A(n6684), .Z(n3969) );
  OR U4716 ( .A(n3970), .B(n3969), .Z(n3971) );
  AND U4717 ( .A(a[327]), .B(b[327]), .Z(n3973) );
  ANDN U4718 ( .B(n3971), .A(n3973), .Z(n3980) );
  NOR U4719 ( .A(n3975), .B(n3974), .Z(n3972) );
  XNOR U4720 ( .A(n3973), .B(n3972), .Z(n3978) );
  XOR U4721 ( .A(n3975), .B(n3974), .Z(n3976) );
  NAND U4722 ( .A(n3976), .B(n6684), .Z(n3977) );
  NAND U4723 ( .A(n3978), .B(n3977), .Z(n6689) );
  XNOR U4724 ( .A(a[328]), .B(b[328]), .Z(n6688) );
  NAND U4725 ( .A(n6689), .B(n6688), .Z(n3979) );
  NANDN U4726 ( .A(n3980), .B(n3979), .Z(n3981) );
  IV U4727 ( .A(n3981), .Z(n3985) );
  AND U4728 ( .A(a[328]), .B(b[328]), .Z(n3986) );
  NOR U4729 ( .A(n3985), .B(n3986), .Z(n3983) );
  XNOR U4730 ( .A(n3986), .B(n3981), .Z(n6694) );
  XNOR U4731 ( .A(a[329]), .B(b[329]), .Z(n6693) );
  AND U4732 ( .A(n6694), .B(n6693), .Z(n3982) );
  OR U4733 ( .A(n3983), .B(n3982), .Z(n3984) );
  AND U4734 ( .A(a[329]), .B(b[329]), .Z(n3988) );
  ANDN U4735 ( .B(n3984), .A(n3988), .Z(n3990) );
  AND U4736 ( .A(n3986), .B(n3985), .Z(n3987) );
  NAND U4737 ( .A(n3988), .B(n3987), .Z(n3993) );
  ANDN U4738 ( .B(n3993), .A(n3990), .Z(n6699) );
  XNOR U4739 ( .A(a[330]), .B(b[330]), .Z(n6698) );
  AND U4740 ( .A(n6699), .B(n6698), .Z(n3989) );
  OR U4741 ( .A(n3990), .B(n3989), .Z(n3991) );
  AND U4742 ( .A(a[330]), .B(b[330]), .Z(n3992) );
  ANDN U4743 ( .B(n3991), .A(n3992), .Z(n3996) );
  NANDN U4744 ( .A(n3993), .B(n3992), .Z(n3994) );
  ANDN U4745 ( .B(n3994), .A(n3996), .Z(n6704) );
  XNOR U4746 ( .A(a[331]), .B(b[331]), .Z(n6703) );
  NAND U4747 ( .A(n6704), .B(n6703), .Z(n3995) );
  NANDN U4748 ( .A(n3996), .B(n3995), .Z(n4002) );
  NAND U4749 ( .A(a[331]), .B(b[331]), .Z(n4003) );
  AND U4750 ( .A(n4002), .B(n4003), .Z(n3998) );
  XOR U4751 ( .A(a[332]), .B(b[332]), .Z(n6709) );
  ANDN U4752 ( .B(n6708), .A(n6709), .Z(n3997) );
  OR U4753 ( .A(n3998), .B(n3997), .Z(n3999) );
  AND U4754 ( .A(a[332]), .B(b[332]), .Z(n4001) );
  ANDN U4755 ( .B(n3999), .A(n4001), .Z(n4008) );
  NOR U4756 ( .A(n4003), .B(n4002), .Z(n4000) );
  XNOR U4757 ( .A(n4001), .B(n4000), .Z(n4006) );
  XOR U4758 ( .A(n4003), .B(n4002), .Z(n4004) );
  NAND U4759 ( .A(n4004), .B(n6709), .Z(n4005) );
  NAND U4760 ( .A(n4006), .B(n4005), .Z(n6714) );
  XNOR U4761 ( .A(a[333]), .B(b[333]), .Z(n6713) );
  NAND U4762 ( .A(n6714), .B(n6713), .Z(n4007) );
  NANDN U4763 ( .A(n4008), .B(n4007), .Z(n4014) );
  NAND U4764 ( .A(a[333]), .B(b[333]), .Z(n4015) );
  AND U4765 ( .A(n4014), .B(n4015), .Z(n4010) );
  XOR U4766 ( .A(a[334]), .B(b[334]), .Z(n6719) );
  ANDN U4767 ( .B(n6718), .A(n6719), .Z(n4009) );
  OR U4768 ( .A(n4010), .B(n4009), .Z(n4011) );
  AND U4769 ( .A(a[334]), .B(b[334]), .Z(n4013) );
  ANDN U4770 ( .B(n4011), .A(n4013), .Z(n4020) );
  NOR U4771 ( .A(n4015), .B(n4014), .Z(n4012) );
  XNOR U4772 ( .A(n4013), .B(n4012), .Z(n4018) );
  XOR U4773 ( .A(n4015), .B(n4014), .Z(n4016) );
  NAND U4774 ( .A(n4016), .B(n6719), .Z(n4017) );
  NAND U4775 ( .A(n4018), .B(n4017), .Z(n6724) );
  XNOR U4776 ( .A(a[335]), .B(b[335]), .Z(n6723) );
  NAND U4777 ( .A(n6724), .B(n6723), .Z(n4019) );
  NANDN U4778 ( .A(n4020), .B(n4019), .Z(n4026) );
  NAND U4779 ( .A(a[335]), .B(b[335]), .Z(n4027) );
  AND U4780 ( .A(n4026), .B(n4027), .Z(n4022) );
  XOR U4781 ( .A(a[336]), .B(b[336]), .Z(n6729) );
  ANDN U4782 ( .B(n6728), .A(n6729), .Z(n4021) );
  OR U4783 ( .A(n4022), .B(n4021), .Z(n4023) );
  AND U4784 ( .A(a[336]), .B(b[336]), .Z(n4025) );
  ANDN U4785 ( .B(n4023), .A(n4025), .Z(n4032) );
  NOR U4786 ( .A(n4027), .B(n4026), .Z(n4024) );
  XNOR U4787 ( .A(n4025), .B(n4024), .Z(n4030) );
  XOR U4788 ( .A(n4027), .B(n4026), .Z(n4028) );
  NAND U4789 ( .A(n4028), .B(n6729), .Z(n4029) );
  NAND U4790 ( .A(n4030), .B(n4029), .Z(n6734) );
  XNOR U4791 ( .A(a[337]), .B(b[337]), .Z(n6733) );
  NAND U4792 ( .A(n6734), .B(n6733), .Z(n4031) );
  NANDN U4793 ( .A(n4032), .B(n4031), .Z(n4038) );
  NAND U4794 ( .A(a[337]), .B(b[337]), .Z(n4039) );
  AND U4795 ( .A(n4038), .B(n4039), .Z(n4034) );
  XOR U4796 ( .A(a[338]), .B(b[338]), .Z(n6739) );
  ANDN U4797 ( .B(n6738), .A(n6739), .Z(n4033) );
  OR U4798 ( .A(n4034), .B(n4033), .Z(n4035) );
  AND U4799 ( .A(a[338]), .B(b[338]), .Z(n4037) );
  ANDN U4800 ( .B(n4035), .A(n4037), .Z(n4044) );
  NOR U4801 ( .A(n4039), .B(n4038), .Z(n4036) );
  XNOR U4802 ( .A(n4037), .B(n4036), .Z(n4042) );
  XOR U4803 ( .A(n4039), .B(n4038), .Z(n4040) );
  NAND U4804 ( .A(n4040), .B(n6739), .Z(n4041) );
  NAND U4805 ( .A(n4042), .B(n4041), .Z(n6744) );
  XNOR U4806 ( .A(a[339]), .B(b[339]), .Z(n6743) );
  NAND U4807 ( .A(n6744), .B(n6743), .Z(n4043) );
  NANDN U4808 ( .A(n4044), .B(n4043), .Z(n4050) );
  NAND U4809 ( .A(a[339]), .B(b[339]), .Z(n4051) );
  AND U4810 ( .A(n4050), .B(n4051), .Z(n4046) );
  XOR U4811 ( .A(a[340]), .B(b[340]), .Z(n6749) );
  ANDN U4812 ( .B(n6748), .A(n6749), .Z(n4045) );
  OR U4813 ( .A(n4046), .B(n4045), .Z(n4047) );
  AND U4814 ( .A(a[340]), .B(b[340]), .Z(n4049) );
  ANDN U4815 ( .B(n4047), .A(n4049), .Z(n4056) );
  NOR U4816 ( .A(n4051), .B(n4050), .Z(n4048) );
  XNOR U4817 ( .A(n4049), .B(n4048), .Z(n4054) );
  XOR U4818 ( .A(n4051), .B(n4050), .Z(n4052) );
  NAND U4819 ( .A(n4052), .B(n6749), .Z(n4053) );
  NAND U4820 ( .A(n4054), .B(n4053), .Z(n6754) );
  XNOR U4821 ( .A(a[341]), .B(b[341]), .Z(n6753) );
  NAND U4822 ( .A(n6754), .B(n6753), .Z(n4055) );
  NANDN U4823 ( .A(n4056), .B(n4055), .Z(n4062) );
  NAND U4824 ( .A(a[341]), .B(b[341]), .Z(n4063) );
  AND U4825 ( .A(n4062), .B(n4063), .Z(n4058) );
  XOR U4826 ( .A(a[342]), .B(b[342]), .Z(n6759) );
  ANDN U4827 ( .B(n6758), .A(n6759), .Z(n4057) );
  OR U4828 ( .A(n4058), .B(n4057), .Z(n4059) );
  AND U4829 ( .A(a[342]), .B(b[342]), .Z(n4061) );
  ANDN U4830 ( .B(n4059), .A(n4061), .Z(n4068) );
  NOR U4831 ( .A(n4063), .B(n4062), .Z(n4060) );
  XNOR U4832 ( .A(n4061), .B(n4060), .Z(n4066) );
  XOR U4833 ( .A(n4063), .B(n4062), .Z(n4064) );
  NAND U4834 ( .A(n4064), .B(n6759), .Z(n4065) );
  NAND U4835 ( .A(n4066), .B(n4065), .Z(n6764) );
  XNOR U4836 ( .A(a[343]), .B(b[343]), .Z(n6763) );
  NAND U4837 ( .A(n6764), .B(n6763), .Z(n4067) );
  NANDN U4838 ( .A(n4068), .B(n4067), .Z(n4074) );
  NAND U4839 ( .A(a[343]), .B(b[343]), .Z(n4075) );
  AND U4840 ( .A(n4074), .B(n4075), .Z(n4070) );
  XOR U4841 ( .A(a[344]), .B(b[344]), .Z(n6769) );
  ANDN U4842 ( .B(n6768), .A(n6769), .Z(n4069) );
  OR U4843 ( .A(n4070), .B(n4069), .Z(n4071) );
  AND U4844 ( .A(a[344]), .B(b[344]), .Z(n4073) );
  ANDN U4845 ( .B(n4071), .A(n4073), .Z(n4080) );
  NOR U4846 ( .A(n4075), .B(n4074), .Z(n4072) );
  XNOR U4847 ( .A(n4073), .B(n4072), .Z(n4078) );
  XOR U4848 ( .A(n4075), .B(n4074), .Z(n4076) );
  NAND U4849 ( .A(n4076), .B(n6769), .Z(n4077) );
  NAND U4850 ( .A(n4078), .B(n4077), .Z(n6774) );
  XNOR U4851 ( .A(a[345]), .B(b[345]), .Z(n6773) );
  NAND U4852 ( .A(n6774), .B(n6773), .Z(n4079) );
  NANDN U4853 ( .A(n4080), .B(n4079), .Z(n4081) );
  IV U4854 ( .A(n4081), .Z(n4085) );
  AND U4855 ( .A(a[345]), .B(b[345]), .Z(n4086) );
  NOR U4856 ( .A(n4085), .B(n4086), .Z(n4083) );
  XNOR U4857 ( .A(n4086), .B(n4081), .Z(n6779) );
  XNOR U4858 ( .A(a[346]), .B(b[346]), .Z(n6778) );
  AND U4859 ( .A(n6779), .B(n6778), .Z(n4082) );
  OR U4860 ( .A(n4083), .B(n4082), .Z(n4084) );
  AND U4861 ( .A(a[346]), .B(b[346]), .Z(n4088) );
  ANDN U4862 ( .B(n4084), .A(n4088), .Z(n4090) );
  AND U4863 ( .A(n4086), .B(n4085), .Z(n4087) );
  NAND U4864 ( .A(n4088), .B(n4087), .Z(n4093) );
  ANDN U4865 ( .B(n4093), .A(n4090), .Z(n6784) );
  XNOR U4866 ( .A(a[347]), .B(b[347]), .Z(n6783) );
  AND U4867 ( .A(n6784), .B(n6783), .Z(n4089) );
  OR U4868 ( .A(n4090), .B(n4089), .Z(n4091) );
  AND U4869 ( .A(a[347]), .B(b[347]), .Z(n4092) );
  ANDN U4870 ( .B(n4091), .A(n4092), .Z(n4096) );
  NANDN U4871 ( .A(n4093), .B(n4092), .Z(n4094) );
  ANDN U4872 ( .B(n4094), .A(n4096), .Z(n6789) );
  XNOR U4873 ( .A(a[348]), .B(b[348]), .Z(n6788) );
  NAND U4874 ( .A(n6789), .B(n6788), .Z(n4095) );
  NANDN U4875 ( .A(n4096), .B(n4095), .Z(n4102) );
  NAND U4876 ( .A(a[348]), .B(b[348]), .Z(n4103) );
  AND U4877 ( .A(n4102), .B(n4103), .Z(n4098) );
  XOR U4878 ( .A(a[349]), .B(b[349]), .Z(n6794) );
  ANDN U4879 ( .B(n6793), .A(n6794), .Z(n4097) );
  OR U4880 ( .A(n4098), .B(n4097), .Z(n4099) );
  AND U4881 ( .A(a[349]), .B(b[349]), .Z(n4101) );
  ANDN U4882 ( .B(n4099), .A(n4101), .Z(n4108) );
  NOR U4883 ( .A(n4103), .B(n4102), .Z(n4100) );
  XNOR U4884 ( .A(n4101), .B(n4100), .Z(n4106) );
  XOR U4885 ( .A(n4103), .B(n4102), .Z(n4104) );
  NAND U4886 ( .A(n4104), .B(n6794), .Z(n4105) );
  NAND U4887 ( .A(n4106), .B(n4105), .Z(n6799) );
  XNOR U4888 ( .A(a[350]), .B(b[350]), .Z(n6798) );
  NAND U4889 ( .A(n6799), .B(n6798), .Z(n4107) );
  NANDN U4890 ( .A(n4108), .B(n4107), .Z(n4114) );
  NAND U4891 ( .A(a[350]), .B(b[350]), .Z(n4115) );
  AND U4892 ( .A(n4114), .B(n4115), .Z(n4110) );
  XOR U4893 ( .A(a[351]), .B(b[351]), .Z(n6804) );
  ANDN U4894 ( .B(n6803), .A(n6804), .Z(n4109) );
  OR U4895 ( .A(n4110), .B(n4109), .Z(n4111) );
  AND U4896 ( .A(a[351]), .B(b[351]), .Z(n4113) );
  ANDN U4897 ( .B(n4111), .A(n4113), .Z(n4120) );
  NOR U4898 ( .A(n4115), .B(n4114), .Z(n4112) );
  XNOR U4899 ( .A(n4113), .B(n4112), .Z(n4118) );
  XOR U4900 ( .A(n4115), .B(n4114), .Z(n4116) );
  NAND U4901 ( .A(n4116), .B(n6804), .Z(n4117) );
  NAND U4902 ( .A(n4118), .B(n4117), .Z(n6809) );
  XNOR U4903 ( .A(a[352]), .B(b[352]), .Z(n6808) );
  NAND U4904 ( .A(n6809), .B(n6808), .Z(n4119) );
  NANDN U4905 ( .A(n4120), .B(n4119), .Z(n4126) );
  NAND U4906 ( .A(a[352]), .B(b[352]), .Z(n4127) );
  AND U4907 ( .A(n4126), .B(n4127), .Z(n4122) );
  XOR U4908 ( .A(a[353]), .B(b[353]), .Z(n6814) );
  ANDN U4909 ( .B(n6813), .A(n6814), .Z(n4121) );
  OR U4910 ( .A(n4122), .B(n4121), .Z(n4123) );
  AND U4911 ( .A(a[353]), .B(b[353]), .Z(n4125) );
  ANDN U4912 ( .B(n4123), .A(n4125), .Z(n4132) );
  NOR U4913 ( .A(n4127), .B(n4126), .Z(n4124) );
  XNOR U4914 ( .A(n4125), .B(n4124), .Z(n4130) );
  XOR U4915 ( .A(n4127), .B(n4126), .Z(n4128) );
  NAND U4916 ( .A(n4128), .B(n6814), .Z(n4129) );
  NAND U4917 ( .A(n4130), .B(n4129), .Z(n6819) );
  XNOR U4918 ( .A(a[354]), .B(b[354]), .Z(n6818) );
  NAND U4919 ( .A(n6819), .B(n6818), .Z(n4131) );
  NANDN U4920 ( .A(n4132), .B(n4131), .Z(n4138) );
  NAND U4921 ( .A(a[354]), .B(b[354]), .Z(n4139) );
  AND U4922 ( .A(n4138), .B(n4139), .Z(n4134) );
  XOR U4923 ( .A(a[355]), .B(b[355]), .Z(n6824) );
  ANDN U4924 ( .B(n6823), .A(n6824), .Z(n4133) );
  OR U4925 ( .A(n4134), .B(n4133), .Z(n4135) );
  AND U4926 ( .A(a[355]), .B(b[355]), .Z(n4137) );
  ANDN U4927 ( .B(n4135), .A(n4137), .Z(n4144) );
  NOR U4928 ( .A(n4139), .B(n4138), .Z(n4136) );
  XNOR U4929 ( .A(n4137), .B(n4136), .Z(n4142) );
  XOR U4930 ( .A(n4139), .B(n4138), .Z(n4140) );
  NAND U4931 ( .A(n4140), .B(n6824), .Z(n4141) );
  NAND U4932 ( .A(n4142), .B(n4141), .Z(n6829) );
  XNOR U4933 ( .A(a[356]), .B(b[356]), .Z(n6828) );
  NAND U4934 ( .A(n6829), .B(n6828), .Z(n4143) );
  NANDN U4935 ( .A(n4144), .B(n4143), .Z(n4150) );
  NAND U4936 ( .A(a[356]), .B(b[356]), .Z(n4151) );
  AND U4937 ( .A(n4150), .B(n4151), .Z(n4146) );
  XOR U4938 ( .A(a[357]), .B(b[357]), .Z(n6834) );
  ANDN U4939 ( .B(n6833), .A(n6834), .Z(n4145) );
  OR U4940 ( .A(n4146), .B(n4145), .Z(n4147) );
  AND U4941 ( .A(a[357]), .B(b[357]), .Z(n4149) );
  ANDN U4942 ( .B(n4147), .A(n4149), .Z(n4156) );
  NOR U4943 ( .A(n4151), .B(n4150), .Z(n4148) );
  XNOR U4944 ( .A(n4149), .B(n4148), .Z(n4154) );
  XOR U4945 ( .A(n4151), .B(n4150), .Z(n4152) );
  NAND U4946 ( .A(n4152), .B(n6834), .Z(n4153) );
  NAND U4947 ( .A(n4154), .B(n4153), .Z(n6839) );
  XNOR U4948 ( .A(a[358]), .B(b[358]), .Z(n6838) );
  NAND U4949 ( .A(n6839), .B(n6838), .Z(n4155) );
  NANDN U4950 ( .A(n4156), .B(n4155), .Z(n4162) );
  NAND U4951 ( .A(a[358]), .B(b[358]), .Z(n4163) );
  AND U4952 ( .A(n4162), .B(n4163), .Z(n4158) );
  XOR U4953 ( .A(a[359]), .B(b[359]), .Z(n6844) );
  ANDN U4954 ( .B(n6843), .A(n6844), .Z(n4157) );
  OR U4955 ( .A(n4158), .B(n4157), .Z(n4159) );
  AND U4956 ( .A(a[359]), .B(b[359]), .Z(n4161) );
  ANDN U4957 ( .B(n4159), .A(n4161), .Z(n4168) );
  NOR U4958 ( .A(n4163), .B(n4162), .Z(n4160) );
  XNOR U4959 ( .A(n4161), .B(n4160), .Z(n4166) );
  XOR U4960 ( .A(n4163), .B(n4162), .Z(n4164) );
  NAND U4961 ( .A(n4164), .B(n6844), .Z(n4165) );
  NAND U4962 ( .A(n4166), .B(n4165), .Z(n6849) );
  XNOR U4963 ( .A(a[360]), .B(b[360]), .Z(n6848) );
  NAND U4964 ( .A(n6849), .B(n6848), .Z(n4167) );
  NANDN U4965 ( .A(n4168), .B(n4167), .Z(n4174) );
  NAND U4966 ( .A(a[360]), .B(b[360]), .Z(n4175) );
  AND U4967 ( .A(n4174), .B(n4175), .Z(n4170) );
  XOR U4968 ( .A(a[361]), .B(b[361]), .Z(n6854) );
  ANDN U4969 ( .B(n6853), .A(n6854), .Z(n4169) );
  OR U4970 ( .A(n4170), .B(n4169), .Z(n4171) );
  AND U4971 ( .A(a[361]), .B(b[361]), .Z(n4173) );
  ANDN U4972 ( .B(n4171), .A(n4173), .Z(n4180) );
  NOR U4973 ( .A(n4175), .B(n4174), .Z(n4172) );
  XNOR U4974 ( .A(n4173), .B(n4172), .Z(n4178) );
  XOR U4975 ( .A(n4175), .B(n4174), .Z(n4176) );
  NAND U4976 ( .A(n4176), .B(n6854), .Z(n4177) );
  NAND U4977 ( .A(n4178), .B(n4177), .Z(n6859) );
  XNOR U4978 ( .A(a[362]), .B(b[362]), .Z(n6858) );
  NAND U4979 ( .A(n6859), .B(n6858), .Z(n4179) );
  NANDN U4980 ( .A(n4180), .B(n4179), .Z(n4186) );
  NAND U4981 ( .A(a[362]), .B(b[362]), .Z(n4187) );
  AND U4982 ( .A(n4186), .B(n4187), .Z(n4182) );
  XOR U4983 ( .A(a[363]), .B(b[363]), .Z(n6864) );
  ANDN U4984 ( .B(n6863), .A(n6864), .Z(n4181) );
  OR U4985 ( .A(n4182), .B(n4181), .Z(n4183) );
  AND U4986 ( .A(a[363]), .B(b[363]), .Z(n4185) );
  ANDN U4987 ( .B(n4183), .A(n4185), .Z(n4192) );
  NOR U4988 ( .A(n4187), .B(n4186), .Z(n4184) );
  XNOR U4989 ( .A(n4185), .B(n4184), .Z(n4190) );
  XOR U4990 ( .A(n4187), .B(n4186), .Z(n4188) );
  NAND U4991 ( .A(n4188), .B(n6864), .Z(n4189) );
  NAND U4992 ( .A(n4190), .B(n4189), .Z(n6869) );
  XNOR U4993 ( .A(a[364]), .B(b[364]), .Z(n6868) );
  NAND U4994 ( .A(n6869), .B(n6868), .Z(n4191) );
  NANDN U4995 ( .A(n4192), .B(n4191), .Z(n4193) );
  IV U4996 ( .A(n4193), .Z(n4197) );
  AND U4997 ( .A(a[364]), .B(b[364]), .Z(n4198) );
  NOR U4998 ( .A(n4197), .B(n4198), .Z(n4195) );
  XNOR U4999 ( .A(n4198), .B(n4193), .Z(n6874) );
  XNOR U5000 ( .A(a[365]), .B(b[365]), .Z(n6873) );
  AND U5001 ( .A(n6874), .B(n6873), .Z(n4194) );
  OR U5002 ( .A(n4195), .B(n4194), .Z(n4196) );
  AND U5003 ( .A(a[365]), .B(b[365]), .Z(n4200) );
  ANDN U5004 ( .B(n4196), .A(n4200), .Z(n4202) );
  AND U5005 ( .A(n4198), .B(n4197), .Z(n4199) );
  NAND U5006 ( .A(n4200), .B(n4199), .Z(n4205) );
  ANDN U5007 ( .B(n4205), .A(n4202), .Z(n6879) );
  XNOR U5008 ( .A(a[366]), .B(b[366]), .Z(n6878) );
  AND U5009 ( .A(n6879), .B(n6878), .Z(n4201) );
  OR U5010 ( .A(n4202), .B(n4201), .Z(n4203) );
  AND U5011 ( .A(a[366]), .B(b[366]), .Z(n4204) );
  ANDN U5012 ( .B(n4203), .A(n4204), .Z(n4208) );
  NANDN U5013 ( .A(n4205), .B(n4204), .Z(n4206) );
  ANDN U5014 ( .B(n4206), .A(n4208), .Z(n6884) );
  XNOR U5015 ( .A(a[367]), .B(b[367]), .Z(n6883) );
  NAND U5016 ( .A(n6884), .B(n6883), .Z(n4207) );
  NANDN U5017 ( .A(n4208), .B(n4207), .Z(n4214) );
  NAND U5018 ( .A(a[367]), .B(b[367]), .Z(n4215) );
  AND U5019 ( .A(n4214), .B(n4215), .Z(n4210) );
  XOR U5020 ( .A(a[368]), .B(b[368]), .Z(n6889) );
  ANDN U5021 ( .B(n6888), .A(n6889), .Z(n4209) );
  OR U5022 ( .A(n4210), .B(n4209), .Z(n4211) );
  AND U5023 ( .A(a[368]), .B(b[368]), .Z(n4213) );
  ANDN U5024 ( .B(n4211), .A(n4213), .Z(n4220) );
  NOR U5025 ( .A(n4215), .B(n4214), .Z(n4212) );
  XNOR U5026 ( .A(n4213), .B(n4212), .Z(n4218) );
  XOR U5027 ( .A(n4215), .B(n4214), .Z(n4216) );
  NAND U5028 ( .A(n4216), .B(n6889), .Z(n4217) );
  NAND U5029 ( .A(n4218), .B(n4217), .Z(n6894) );
  XNOR U5030 ( .A(a[369]), .B(b[369]), .Z(n6893) );
  NAND U5031 ( .A(n6894), .B(n6893), .Z(n4219) );
  NANDN U5032 ( .A(n4220), .B(n4219), .Z(n4226) );
  NAND U5033 ( .A(a[369]), .B(b[369]), .Z(n4227) );
  AND U5034 ( .A(n4226), .B(n4227), .Z(n4222) );
  XOR U5035 ( .A(a[370]), .B(b[370]), .Z(n6899) );
  ANDN U5036 ( .B(n6898), .A(n6899), .Z(n4221) );
  OR U5037 ( .A(n4222), .B(n4221), .Z(n4223) );
  AND U5038 ( .A(a[370]), .B(b[370]), .Z(n4225) );
  ANDN U5039 ( .B(n4223), .A(n4225), .Z(n4232) );
  NOR U5040 ( .A(n4227), .B(n4226), .Z(n4224) );
  XNOR U5041 ( .A(n4225), .B(n4224), .Z(n4230) );
  XOR U5042 ( .A(n4227), .B(n4226), .Z(n4228) );
  NAND U5043 ( .A(n4228), .B(n6899), .Z(n4229) );
  NAND U5044 ( .A(n4230), .B(n4229), .Z(n6904) );
  XNOR U5045 ( .A(a[371]), .B(b[371]), .Z(n6903) );
  NAND U5046 ( .A(n6904), .B(n6903), .Z(n4231) );
  NANDN U5047 ( .A(n4232), .B(n4231), .Z(n4238) );
  NAND U5048 ( .A(a[371]), .B(b[371]), .Z(n4239) );
  AND U5049 ( .A(n4238), .B(n4239), .Z(n4234) );
  XOR U5050 ( .A(a[372]), .B(b[372]), .Z(n6909) );
  ANDN U5051 ( .B(n6908), .A(n6909), .Z(n4233) );
  OR U5052 ( .A(n4234), .B(n4233), .Z(n4235) );
  AND U5053 ( .A(a[372]), .B(b[372]), .Z(n4237) );
  ANDN U5054 ( .B(n4235), .A(n4237), .Z(n4244) );
  NOR U5055 ( .A(n4239), .B(n4238), .Z(n4236) );
  XNOR U5056 ( .A(n4237), .B(n4236), .Z(n4242) );
  XOR U5057 ( .A(n4239), .B(n4238), .Z(n4240) );
  NAND U5058 ( .A(n4240), .B(n6909), .Z(n4241) );
  NAND U5059 ( .A(n4242), .B(n4241), .Z(n6914) );
  XNOR U5060 ( .A(a[373]), .B(b[373]), .Z(n6913) );
  NAND U5061 ( .A(n6914), .B(n6913), .Z(n4243) );
  NANDN U5062 ( .A(n4244), .B(n4243), .Z(n4250) );
  NAND U5063 ( .A(a[373]), .B(b[373]), .Z(n4251) );
  AND U5064 ( .A(n4250), .B(n4251), .Z(n4246) );
  XOR U5065 ( .A(a[374]), .B(b[374]), .Z(n6919) );
  ANDN U5066 ( .B(n6918), .A(n6919), .Z(n4245) );
  OR U5067 ( .A(n4246), .B(n4245), .Z(n4247) );
  AND U5068 ( .A(a[374]), .B(b[374]), .Z(n4249) );
  ANDN U5069 ( .B(n4247), .A(n4249), .Z(n4256) );
  NOR U5070 ( .A(n4251), .B(n4250), .Z(n4248) );
  XNOR U5071 ( .A(n4249), .B(n4248), .Z(n4254) );
  XOR U5072 ( .A(n4251), .B(n4250), .Z(n4252) );
  NAND U5073 ( .A(n4252), .B(n6919), .Z(n4253) );
  NAND U5074 ( .A(n4254), .B(n4253), .Z(n6924) );
  XNOR U5075 ( .A(a[375]), .B(b[375]), .Z(n6923) );
  NAND U5076 ( .A(n6924), .B(n6923), .Z(n4255) );
  NANDN U5077 ( .A(n4256), .B(n4255), .Z(n4262) );
  NAND U5078 ( .A(a[375]), .B(b[375]), .Z(n4263) );
  AND U5079 ( .A(n4262), .B(n4263), .Z(n4258) );
  XOR U5080 ( .A(a[376]), .B(b[376]), .Z(n6929) );
  ANDN U5081 ( .B(n6928), .A(n6929), .Z(n4257) );
  OR U5082 ( .A(n4258), .B(n4257), .Z(n4259) );
  AND U5083 ( .A(a[376]), .B(b[376]), .Z(n4261) );
  ANDN U5084 ( .B(n4259), .A(n4261), .Z(n4268) );
  NOR U5085 ( .A(n4263), .B(n4262), .Z(n4260) );
  XNOR U5086 ( .A(n4261), .B(n4260), .Z(n4266) );
  XOR U5087 ( .A(n4263), .B(n4262), .Z(n4264) );
  NAND U5088 ( .A(n4264), .B(n6929), .Z(n4265) );
  NAND U5089 ( .A(n4266), .B(n4265), .Z(n6934) );
  XNOR U5090 ( .A(a[377]), .B(b[377]), .Z(n6933) );
  NAND U5091 ( .A(n6934), .B(n6933), .Z(n4267) );
  NANDN U5092 ( .A(n4268), .B(n4267), .Z(n4274) );
  NAND U5093 ( .A(a[377]), .B(b[377]), .Z(n4275) );
  AND U5094 ( .A(n4274), .B(n4275), .Z(n4270) );
  XOR U5095 ( .A(a[378]), .B(b[378]), .Z(n6939) );
  ANDN U5096 ( .B(n6938), .A(n6939), .Z(n4269) );
  OR U5097 ( .A(n4270), .B(n4269), .Z(n4271) );
  AND U5098 ( .A(a[378]), .B(b[378]), .Z(n4273) );
  ANDN U5099 ( .B(n4271), .A(n4273), .Z(n4280) );
  NOR U5100 ( .A(n4275), .B(n4274), .Z(n4272) );
  XNOR U5101 ( .A(n4273), .B(n4272), .Z(n4278) );
  XOR U5102 ( .A(n4275), .B(n4274), .Z(n4276) );
  NAND U5103 ( .A(n4276), .B(n6939), .Z(n4277) );
  NAND U5104 ( .A(n4278), .B(n4277), .Z(n6944) );
  XNOR U5105 ( .A(a[379]), .B(b[379]), .Z(n6943) );
  NAND U5106 ( .A(n6944), .B(n6943), .Z(n4279) );
  NANDN U5107 ( .A(n4280), .B(n4279), .Z(n4286) );
  NAND U5108 ( .A(a[379]), .B(b[379]), .Z(n4287) );
  AND U5109 ( .A(n4286), .B(n4287), .Z(n4282) );
  XOR U5110 ( .A(a[380]), .B(b[380]), .Z(n6949) );
  ANDN U5111 ( .B(n6948), .A(n6949), .Z(n4281) );
  OR U5112 ( .A(n4282), .B(n4281), .Z(n4283) );
  AND U5113 ( .A(a[380]), .B(b[380]), .Z(n4285) );
  ANDN U5114 ( .B(n4283), .A(n4285), .Z(n4292) );
  NOR U5115 ( .A(n4287), .B(n4286), .Z(n4284) );
  XNOR U5116 ( .A(n4285), .B(n4284), .Z(n4290) );
  XOR U5117 ( .A(n4287), .B(n4286), .Z(n4288) );
  NAND U5118 ( .A(n4288), .B(n6949), .Z(n4289) );
  NAND U5119 ( .A(n4290), .B(n4289), .Z(n6954) );
  XNOR U5120 ( .A(a[381]), .B(b[381]), .Z(n6953) );
  NAND U5121 ( .A(n6954), .B(n6953), .Z(n4291) );
  NANDN U5122 ( .A(n4292), .B(n4291), .Z(n4298) );
  NAND U5123 ( .A(a[381]), .B(b[381]), .Z(n4299) );
  AND U5124 ( .A(n4298), .B(n4299), .Z(n4294) );
  XOR U5125 ( .A(a[382]), .B(b[382]), .Z(n6959) );
  ANDN U5126 ( .B(n6958), .A(n6959), .Z(n4293) );
  OR U5127 ( .A(n4294), .B(n4293), .Z(n4295) );
  AND U5128 ( .A(a[382]), .B(b[382]), .Z(n4297) );
  ANDN U5129 ( .B(n4295), .A(n4297), .Z(n4304) );
  NOR U5130 ( .A(n4299), .B(n4298), .Z(n4296) );
  XNOR U5131 ( .A(n4297), .B(n4296), .Z(n4302) );
  XOR U5132 ( .A(n4299), .B(n4298), .Z(n4300) );
  NAND U5133 ( .A(n4300), .B(n6959), .Z(n4301) );
  NAND U5134 ( .A(n4302), .B(n4301), .Z(n6964) );
  XNOR U5135 ( .A(a[383]), .B(b[383]), .Z(n6963) );
  NAND U5136 ( .A(n6964), .B(n6963), .Z(n4303) );
  NANDN U5137 ( .A(n4304), .B(n4303), .Z(n4310) );
  NAND U5138 ( .A(a[383]), .B(b[383]), .Z(n4311) );
  AND U5139 ( .A(n4310), .B(n4311), .Z(n4306) );
  XOR U5140 ( .A(a[384]), .B(b[384]), .Z(n6969) );
  ANDN U5141 ( .B(n6968), .A(n6969), .Z(n4305) );
  OR U5142 ( .A(n4306), .B(n4305), .Z(n4307) );
  AND U5143 ( .A(a[384]), .B(b[384]), .Z(n4309) );
  ANDN U5144 ( .B(n4307), .A(n4309), .Z(n4316) );
  NOR U5145 ( .A(n4311), .B(n4310), .Z(n4308) );
  XNOR U5146 ( .A(n4309), .B(n4308), .Z(n4314) );
  XOR U5147 ( .A(n4311), .B(n4310), .Z(n4312) );
  NAND U5148 ( .A(n4312), .B(n6969), .Z(n4313) );
  NAND U5149 ( .A(n4314), .B(n4313), .Z(n6974) );
  XNOR U5150 ( .A(a[385]), .B(b[385]), .Z(n6973) );
  NAND U5151 ( .A(n6974), .B(n6973), .Z(n4315) );
  NANDN U5152 ( .A(n4316), .B(n4315), .Z(n4322) );
  NAND U5153 ( .A(a[385]), .B(b[385]), .Z(n4323) );
  AND U5154 ( .A(n4322), .B(n4323), .Z(n4318) );
  XOR U5155 ( .A(a[386]), .B(b[386]), .Z(n6979) );
  ANDN U5156 ( .B(n6978), .A(n6979), .Z(n4317) );
  OR U5157 ( .A(n4318), .B(n4317), .Z(n4319) );
  AND U5158 ( .A(a[386]), .B(b[386]), .Z(n4321) );
  ANDN U5159 ( .B(n4319), .A(n4321), .Z(n4328) );
  NOR U5160 ( .A(n4323), .B(n4322), .Z(n4320) );
  XNOR U5161 ( .A(n4321), .B(n4320), .Z(n4326) );
  XOR U5162 ( .A(n4323), .B(n4322), .Z(n4324) );
  NAND U5163 ( .A(n4324), .B(n6979), .Z(n4325) );
  NAND U5164 ( .A(n4326), .B(n4325), .Z(n6984) );
  XNOR U5165 ( .A(a[387]), .B(b[387]), .Z(n6983) );
  NAND U5166 ( .A(n6984), .B(n6983), .Z(n4327) );
  NANDN U5167 ( .A(n4328), .B(n4327), .Z(n4334) );
  NAND U5168 ( .A(a[387]), .B(b[387]), .Z(n4335) );
  AND U5169 ( .A(n4334), .B(n4335), .Z(n4330) );
  XOR U5170 ( .A(a[388]), .B(b[388]), .Z(n6989) );
  ANDN U5171 ( .B(n6988), .A(n6989), .Z(n4329) );
  OR U5172 ( .A(n4330), .B(n4329), .Z(n4331) );
  AND U5173 ( .A(a[388]), .B(b[388]), .Z(n4333) );
  ANDN U5174 ( .B(n4331), .A(n4333), .Z(n4340) );
  NOR U5175 ( .A(n4335), .B(n4334), .Z(n4332) );
  XNOR U5176 ( .A(n4333), .B(n4332), .Z(n4338) );
  XOR U5177 ( .A(n4335), .B(n4334), .Z(n4336) );
  NAND U5178 ( .A(n4336), .B(n6989), .Z(n4337) );
  NAND U5179 ( .A(n4338), .B(n4337), .Z(n6994) );
  XNOR U5180 ( .A(a[389]), .B(b[389]), .Z(n6993) );
  NAND U5181 ( .A(n6994), .B(n6993), .Z(n4339) );
  NANDN U5182 ( .A(n4340), .B(n4339), .Z(n4346) );
  NAND U5183 ( .A(a[389]), .B(b[389]), .Z(n4347) );
  AND U5184 ( .A(n4346), .B(n4347), .Z(n4342) );
  XOR U5185 ( .A(a[390]), .B(b[390]), .Z(n6999) );
  ANDN U5186 ( .B(n6998), .A(n6999), .Z(n4341) );
  OR U5187 ( .A(n4342), .B(n4341), .Z(n4343) );
  AND U5188 ( .A(a[390]), .B(b[390]), .Z(n4345) );
  ANDN U5189 ( .B(n4343), .A(n4345), .Z(n4352) );
  NOR U5190 ( .A(n4347), .B(n4346), .Z(n4344) );
  XNOR U5191 ( .A(n4345), .B(n4344), .Z(n4350) );
  XOR U5192 ( .A(n4347), .B(n4346), .Z(n4348) );
  NAND U5193 ( .A(n4348), .B(n6999), .Z(n4349) );
  NAND U5194 ( .A(n4350), .B(n4349), .Z(n7004) );
  XNOR U5195 ( .A(a[391]), .B(b[391]), .Z(n7003) );
  NAND U5196 ( .A(n7004), .B(n7003), .Z(n4351) );
  NANDN U5197 ( .A(n4352), .B(n4351), .Z(n4358) );
  NAND U5198 ( .A(a[391]), .B(b[391]), .Z(n4359) );
  AND U5199 ( .A(n4358), .B(n4359), .Z(n4354) );
  XOR U5200 ( .A(a[392]), .B(b[392]), .Z(n7009) );
  ANDN U5201 ( .B(n7008), .A(n7009), .Z(n4353) );
  OR U5202 ( .A(n4354), .B(n4353), .Z(n4355) );
  AND U5203 ( .A(a[392]), .B(b[392]), .Z(n4357) );
  ANDN U5204 ( .B(n4355), .A(n4357), .Z(n4364) );
  NOR U5205 ( .A(n4359), .B(n4358), .Z(n4356) );
  XNOR U5206 ( .A(n4357), .B(n4356), .Z(n4362) );
  XOR U5207 ( .A(n4359), .B(n4358), .Z(n4360) );
  NAND U5208 ( .A(n4360), .B(n7009), .Z(n4361) );
  NAND U5209 ( .A(n4362), .B(n4361), .Z(n7014) );
  XNOR U5210 ( .A(a[393]), .B(b[393]), .Z(n7013) );
  NAND U5211 ( .A(n7014), .B(n7013), .Z(n4363) );
  NANDN U5212 ( .A(n4364), .B(n4363), .Z(n4370) );
  NAND U5213 ( .A(a[393]), .B(b[393]), .Z(n4371) );
  AND U5214 ( .A(n4370), .B(n4371), .Z(n4366) );
  XOR U5215 ( .A(a[394]), .B(b[394]), .Z(n7019) );
  ANDN U5216 ( .B(n7018), .A(n7019), .Z(n4365) );
  OR U5217 ( .A(n4366), .B(n4365), .Z(n4367) );
  AND U5218 ( .A(a[394]), .B(b[394]), .Z(n4369) );
  ANDN U5219 ( .B(n4367), .A(n4369), .Z(n4376) );
  NOR U5220 ( .A(n4371), .B(n4370), .Z(n4368) );
  XNOR U5221 ( .A(n4369), .B(n4368), .Z(n4374) );
  XOR U5222 ( .A(n4371), .B(n4370), .Z(n4372) );
  NAND U5223 ( .A(n4372), .B(n7019), .Z(n4373) );
  NAND U5224 ( .A(n4374), .B(n4373), .Z(n7024) );
  XNOR U5225 ( .A(a[395]), .B(b[395]), .Z(n7023) );
  NAND U5226 ( .A(n7024), .B(n7023), .Z(n4375) );
  NANDN U5227 ( .A(n4376), .B(n4375), .Z(n4382) );
  NAND U5228 ( .A(a[395]), .B(b[395]), .Z(n4383) );
  AND U5229 ( .A(n4382), .B(n4383), .Z(n4378) );
  XOR U5230 ( .A(a[396]), .B(b[396]), .Z(n7029) );
  ANDN U5231 ( .B(n7028), .A(n7029), .Z(n4377) );
  OR U5232 ( .A(n4378), .B(n4377), .Z(n4379) );
  AND U5233 ( .A(a[396]), .B(b[396]), .Z(n4381) );
  ANDN U5234 ( .B(n4379), .A(n4381), .Z(n4388) );
  NOR U5235 ( .A(n4383), .B(n4382), .Z(n4380) );
  XNOR U5236 ( .A(n4381), .B(n4380), .Z(n4386) );
  XOR U5237 ( .A(n4383), .B(n4382), .Z(n4384) );
  NAND U5238 ( .A(n4384), .B(n7029), .Z(n4385) );
  NAND U5239 ( .A(n4386), .B(n4385), .Z(n7034) );
  XNOR U5240 ( .A(a[397]), .B(b[397]), .Z(n7033) );
  NAND U5241 ( .A(n7034), .B(n7033), .Z(n4387) );
  NANDN U5242 ( .A(n4388), .B(n4387), .Z(n4394) );
  NAND U5243 ( .A(a[397]), .B(b[397]), .Z(n4395) );
  AND U5244 ( .A(n4394), .B(n4395), .Z(n4390) );
  XOR U5245 ( .A(a[398]), .B(b[398]), .Z(n7039) );
  ANDN U5246 ( .B(n7038), .A(n7039), .Z(n4389) );
  OR U5247 ( .A(n4390), .B(n4389), .Z(n4391) );
  AND U5248 ( .A(a[398]), .B(b[398]), .Z(n4393) );
  ANDN U5249 ( .B(n4391), .A(n4393), .Z(n4400) );
  NOR U5250 ( .A(n4395), .B(n4394), .Z(n4392) );
  XNOR U5251 ( .A(n4393), .B(n4392), .Z(n4398) );
  XOR U5252 ( .A(n4395), .B(n4394), .Z(n4396) );
  NAND U5253 ( .A(n4396), .B(n7039), .Z(n4397) );
  NAND U5254 ( .A(n4398), .B(n4397), .Z(n7044) );
  XNOR U5255 ( .A(a[399]), .B(b[399]), .Z(n7043) );
  NAND U5256 ( .A(n7044), .B(n7043), .Z(n4399) );
  NANDN U5257 ( .A(n4400), .B(n4399), .Z(n4406) );
  NAND U5258 ( .A(a[399]), .B(b[399]), .Z(n4407) );
  AND U5259 ( .A(n4406), .B(n4407), .Z(n4402) );
  XOR U5260 ( .A(a[400]), .B(b[400]), .Z(n7049) );
  ANDN U5261 ( .B(n7048), .A(n7049), .Z(n4401) );
  OR U5262 ( .A(n4402), .B(n4401), .Z(n4403) );
  AND U5263 ( .A(a[400]), .B(b[400]), .Z(n4405) );
  ANDN U5264 ( .B(n4403), .A(n4405), .Z(n4412) );
  NOR U5265 ( .A(n4407), .B(n4406), .Z(n4404) );
  XNOR U5266 ( .A(n4405), .B(n4404), .Z(n4410) );
  XOR U5267 ( .A(n4407), .B(n4406), .Z(n4408) );
  NAND U5268 ( .A(n4408), .B(n7049), .Z(n4409) );
  NAND U5269 ( .A(n4410), .B(n4409), .Z(n7054) );
  XNOR U5270 ( .A(a[401]), .B(b[401]), .Z(n7053) );
  NAND U5271 ( .A(n7054), .B(n7053), .Z(n4411) );
  NANDN U5272 ( .A(n4412), .B(n4411), .Z(n4418) );
  NAND U5273 ( .A(a[401]), .B(b[401]), .Z(n4419) );
  AND U5274 ( .A(n4418), .B(n4419), .Z(n4414) );
  XOR U5275 ( .A(a[402]), .B(b[402]), .Z(n7059) );
  ANDN U5276 ( .B(n7058), .A(n7059), .Z(n4413) );
  OR U5277 ( .A(n4414), .B(n4413), .Z(n4415) );
  AND U5278 ( .A(a[402]), .B(b[402]), .Z(n4417) );
  ANDN U5279 ( .B(n4415), .A(n4417), .Z(n4424) );
  NOR U5280 ( .A(n4419), .B(n4418), .Z(n4416) );
  XNOR U5281 ( .A(n4417), .B(n4416), .Z(n4422) );
  XOR U5282 ( .A(n4419), .B(n4418), .Z(n4420) );
  NAND U5283 ( .A(n4420), .B(n7059), .Z(n4421) );
  NAND U5284 ( .A(n4422), .B(n4421), .Z(n7064) );
  XNOR U5285 ( .A(a[403]), .B(b[403]), .Z(n7063) );
  NAND U5286 ( .A(n7064), .B(n7063), .Z(n4423) );
  NANDN U5287 ( .A(n4424), .B(n4423), .Z(n4430) );
  NAND U5288 ( .A(a[403]), .B(b[403]), .Z(n4431) );
  AND U5289 ( .A(n4430), .B(n4431), .Z(n4426) );
  XOR U5290 ( .A(a[404]), .B(b[404]), .Z(n7069) );
  ANDN U5291 ( .B(n7068), .A(n7069), .Z(n4425) );
  OR U5292 ( .A(n4426), .B(n4425), .Z(n4427) );
  AND U5293 ( .A(a[404]), .B(b[404]), .Z(n4429) );
  ANDN U5294 ( .B(n4427), .A(n4429), .Z(n4436) );
  NOR U5295 ( .A(n4431), .B(n4430), .Z(n4428) );
  XNOR U5296 ( .A(n4429), .B(n4428), .Z(n4434) );
  XOR U5297 ( .A(n4431), .B(n4430), .Z(n4432) );
  NAND U5298 ( .A(n4432), .B(n7069), .Z(n4433) );
  NAND U5299 ( .A(n4434), .B(n4433), .Z(n7074) );
  XNOR U5300 ( .A(a[405]), .B(b[405]), .Z(n7073) );
  NAND U5301 ( .A(n7074), .B(n7073), .Z(n4435) );
  NANDN U5302 ( .A(n4436), .B(n4435), .Z(n4442) );
  NAND U5303 ( .A(a[405]), .B(b[405]), .Z(n4443) );
  AND U5304 ( .A(n4442), .B(n4443), .Z(n4438) );
  XOR U5305 ( .A(a[406]), .B(b[406]), .Z(n7079) );
  ANDN U5306 ( .B(n7078), .A(n7079), .Z(n4437) );
  OR U5307 ( .A(n4438), .B(n4437), .Z(n4439) );
  AND U5308 ( .A(a[406]), .B(b[406]), .Z(n4441) );
  ANDN U5309 ( .B(n4439), .A(n4441), .Z(n4448) );
  NOR U5310 ( .A(n4443), .B(n4442), .Z(n4440) );
  XNOR U5311 ( .A(n4441), .B(n4440), .Z(n4446) );
  XOR U5312 ( .A(n4443), .B(n4442), .Z(n4444) );
  NAND U5313 ( .A(n4444), .B(n7079), .Z(n4445) );
  NAND U5314 ( .A(n4446), .B(n4445), .Z(n7084) );
  XNOR U5315 ( .A(a[407]), .B(b[407]), .Z(n7083) );
  NAND U5316 ( .A(n7084), .B(n7083), .Z(n4447) );
  NANDN U5317 ( .A(n4448), .B(n4447), .Z(n4449) );
  IV U5318 ( .A(n4449), .Z(n4453) );
  AND U5319 ( .A(a[407]), .B(b[407]), .Z(n4454) );
  NOR U5320 ( .A(n4453), .B(n4454), .Z(n4451) );
  XNOR U5321 ( .A(n4454), .B(n4449), .Z(n7089) );
  XNOR U5322 ( .A(a[408]), .B(b[408]), .Z(n7088) );
  AND U5323 ( .A(n7089), .B(n7088), .Z(n4450) );
  OR U5324 ( .A(n4451), .B(n4450), .Z(n4452) );
  AND U5325 ( .A(a[408]), .B(b[408]), .Z(n4456) );
  ANDN U5326 ( .B(n4452), .A(n4456), .Z(n4458) );
  AND U5327 ( .A(n4454), .B(n4453), .Z(n4455) );
  NAND U5328 ( .A(n4456), .B(n4455), .Z(n4461) );
  ANDN U5329 ( .B(n4461), .A(n4458), .Z(n7094) );
  XNOR U5330 ( .A(a[409]), .B(b[409]), .Z(n7093) );
  AND U5331 ( .A(n7094), .B(n7093), .Z(n4457) );
  OR U5332 ( .A(n4458), .B(n4457), .Z(n4459) );
  AND U5333 ( .A(n4460), .B(n4459), .Z(n4464) );
  OR U5334 ( .A(n4461), .B(n4460), .Z(n4462) );
  ANDN U5335 ( .B(n4462), .A(n4464), .Z(n7099) );
  XNOR U5336 ( .A(a[410]), .B(b[410]), .Z(n7098) );
  NAND U5337 ( .A(n7099), .B(n7098), .Z(n4463) );
  NANDN U5338 ( .A(n4464), .B(n4463), .Z(n4470) );
  NAND U5339 ( .A(a[410]), .B(b[410]), .Z(n4471) );
  AND U5340 ( .A(n4470), .B(n4471), .Z(n4466) );
  XOR U5341 ( .A(a[411]), .B(b[411]), .Z(n7104) );
  ANDN U5342 ( .B(n7103), .A(n7104), .Z(n4465) );
  OR U5343 ( .A(n4466), .B(n4465), .Z(n4467) );
  AND U5344 ( .A(a[411]), .B(b[411]), .Z(n4469) );
  ANDN U5345 ( .B(n4467), .A(n4469), .Z(n4476) );
  NOR U5346 ( .A(n4471), .B(n4470), .Z(n4468) );
  XNOR U5347 ( .A(n4469), .B(n4468), .Z(n4474) );
  XOR U5348 ( .A(n4471), .B(n4470), .Z(n4472) );
  NAND U5349 ( .A(n4472), .B(n7104), .Z(n4473) );
  NAND U5350 ( .A(n4474), .B(n4473), .Z(n7109) );
  XNOR U5351 ( .A(a[412]), .B(b[412]), .Z(n7108) );
  NAND U5352 ( .A(n7109), .B(n7108), .Z(n4475) );
  NANDN U5353 ( .A(n4476), .B(n4475), .Z(n4477) );
  IV U5354 ( .A(n4477), .Z(n4481) );
  AND U5355 ( .A(a[412]), .B(b[412]), .Z(n4482) );
  NOR U5356 ( .A(n4481), .B(n4482), .Z(n4479) );
  XNOR U5357 ( .A(n4482), .B(n4477), .Z(n7114) );
  XNOR U5358 ( .A(a[413]), .B(b[413]), .Z(n7113) );
  AND U5359 ( .A(n7114), .B(n7113), .Z(n4478) );
  OR U5360 ( .A(n4479), .B(n4478), .Z(n4480) );
  AND U5361 ( .A(a[413]), .B(b[413]), .Z(n4484) );
  ANDN U5362 ( .B(n4480), .A(n4484), .Z(n4486) );
  AND U5363 ( .A(n4482), .B(n4481), .Z(n4483) );
  NAND U5364 ( .A(n4484), .B(n4483), .Z(n4489) );
  ANDN U5365 ( .B(n4489), .A(n4486), .Z(n7119) );
  XNOR U5366 ( .A(a[414]), .B(b[414]), .Z(n7118) );
  AND U5367 ( .A(n7119), .B(n7118), .Z(n4485) );
  OR U5368 ( .A(n4486), .B(n4485), .Z(n4487) );
  AND U5369 ( .A(a[414]), .B(b[414]), .Z(n4488) );
  ANDN U5370 ( .B(n4487), .A(n4488), .Z(n4492) );
  NANDN U5371 ( .A(n4489), .B(n4488), .Z(n4490) );
  ANDN U5372 ( .B(n4490), .A(n4492), .Z(n7124) );
  XNOR U5373 ( .A(a[415]), .B(b[415]), .Z(n7123) );
  NAND U5374 ( .A(n7124), .B(n7123), .Z(n4491) );
  NANDN U5375 ( .A(n4492), .B(n4491), .Z(n4498) );
  NAND U5376 ( .A(a[415]), .B(b[415]), .Z(n4499) );
  AND U5377 ( .A(n4498), .B(n4499), .Z(n4494) );
  XOR U5378 ( .A(a[416]), .B(b[416]), .Z(n7129) );
  ANDN U5379 ( .B(n7128), .A(n7129), .Z(n4493) );
  OR U5380 ( .A(n4494), .B(n4493), .Z(n4495) );
  AND U5381 ( .A(a[416]), .B(b[416]), .Z(n4497) );
  ANDN U5382 ( .B(n4495), .A(n4497), .Z(n4504) );
  NOR U5383 ( .A(n4499), .B(n4498), .Z(n4496) );
  XNOR U5384 ( .A(n4497), .B(n4496), .Z(n4502) );
  XOR U5385 ( .A(n4499), .B(n4498), .Z(n4500) );
  NAND U5386 ( .A(n4500), .B(n7129), .Z(n4501) );
  NAND U5387 ( .A(n4502), .B(n4501), .Z(n7134) );
  XNOR U5388 ( .A(a[417]), .B(b[417]), .Z(n7133) );
  NAND U5389 ( .A(n7134), .B(n7133), .Z(n4503) );
  NANDN U5390 ( .A(n4504), .B(n4503), .Z(n4510) );
  NAND U5391 ( .A(a[417]), .B(b[417]), .Z(n4511) );
  AND U5392 ( .A(n4510), .B(n4511), .Z(n4506) );
  XOR U5393 ( .A(a[418]), .B(b[418]), .Z(n7139) );
  ANDN U5394 ( .B(n7138), .A(n7139), .Z(n4505) );
  OR U5395 ( .A(n4506), .B(n4505), .Z(n4507) );
  AND U5396 ( .A(a[418]), .B(b[418]), .Z(n4509) );
  ANDN U5397 ( .B(n4507), .A(n4509), .Z(n4516) );
  NOR U5398 ( .A(n4511), .B(n4510), .Z(n4508) );
  XNOR U5399 ( .A(n4509), .B(n4508), .Z(n4514) );
  XOR U5400 ( .A(n4511), .B(n4510), .Z(n4512) );
  NAND U5401 ( .A(n4512), .B(n7139), .Z(n4513) );
  NAND U5402 ( .A(n4514), .B(n4513), .Z(n7144) );
  XNOR U5403 ( .A(a[419]), .B(b[419]), .Z(n7143) );
  NAND U5404 ( .A(n7144), .B(n7143), .Z(n4515) );
  NANDN U5405 ( .A(n4516), .B(n4515), .Z(n4521) );
  ANDN U5406 ( .B(n4520), .A(n4521), .Z(n4517) );
  XOR U5407 ( .A(n4522), .B(n4517), .Z(n4519) );
  XOR U5408 ( .A(a[420]), .B(b[420]), .Z(n7149) );
  XNOR U5409 ( .A(n4520), .B(n4521), .Z(n7148) );
  NAND U5410 ( .A(n7149), .B(n7148), .Z(n4518) );
  NAND U5411 ( .A(n4519), .B(n4518), .Z(n7154) );
  XNOR U5412 ( .A(a[421]), .B(b[421]), .Z(n7153) );
  IV U5413 ( .A(n4523), .Z(n4525) );
  XNOR U5414 ( .A(n4524), .B(n4523), .Z(n7159) );
  XNOR U5415 ( .A(a[422]), .B(b[422]), .Z(n7158) );
  AND U5416 ( .A(a[422]), .B(b[422]), .Z(n4527) );
  NOR U5417 ( .A(n4525), .B(n4524), .Z(n4526) );
  NAND U5418 ( .A(n4527), .B(n4526), .Z(n4532) );
  ANDN U5419 ( .B(n4532), .A(n4529), .Z(n7164) );
  XNOR U5420 ( .A(a[423]), .B(b[423]), .Z(n7163) );
  NAND U5421 ( .A(n7164), .B(n7163), .Z(n4528) );
  NANDN U5422 ( .A(n4529), .B(n4528), .Z(n4530) );
  AND U5423 ( .A(n4531), .B(n4530), .Z(n4535) );
  OR U5424 ( .A(n4532), .B(n4531), .Z(n4533) );
  ANDN U5425 ( .B(n4533), .A(n4535), .Z(n7169) );
  XNOR U5426 ( .A(a[424]), .B(b[424]), .Z(n7168) );
  NAND U5427 ( .A(n7169), .B(n7168), .Z(n4534) );
  NANDN U5428 ( .A(n4535), .B(n4534), .Z(n4541) );
  NAND U5429 ( .A(a[424]), .B(b[424]), .Z(n4542) );
  AND U5430 ( .A(n4541), .B(n4542), .Z(n4537) );
  XOR U5431 ( .A(a[425]), .B(b[425]), .Z(n7174) );
  ANDN U5432 ( .B(n7173), .A(n7174), .Z(n4536) );
  OR U5433 ( .A(n4537), .B(n4536), .Z(n4538) );
  AND U5434 ( .A(a[425]), .B(b[425]), .Z(n4540) );
  ANDN U5435 ( .B(n4538), .A(n4540), .Z(n4547) );
  NOR U5436 ( .A(n4542), .B(n4541), .Z(n4539) );
  XNOR U5437 ( .A(n4540), .B(n4539), .Z(n4545) );
  XOR U5438 ( .A(n4542), .B(n4541), .Z(n4543) );
  NAND U5439 ( .A(n4543), .B(n7174), .Z(n4544) );
  NAND U5440 ( .A(n4545), .B(n4544), .Z(n7179) );
  XNOR U5441 ( .A(a[426]), .B(b[426]), .Z(n7178) );
  NAND U5442 ( .A(n7179), .B(n7178), .Z(n4546) );
  NANDN U5443 ( .A(n4547), .B(n4546), .Z(n4553) );
  NAND U5444 ( .A(a[426]), .B(b[426]), .Z(n4554) );
  AND U5445 ( .A(n4553), .B(n4554), .Z(n4549) );
  XOR U5446 ( .A(a[427]), .B(b[427]), .Z(n7184) );
  ANDN U5447 ( .B(n7183), .A(n7184), .Z(n4548) );
  OR U5448 ( .A(n4549), .B(n4548), .Z(n4550) );
  AND U5449 ( .A(a[427]), .B(b[427]), .Z(n4552) );
  ANDN U5450 ( .B(n4550), .A(n4552), .Z(n4559) );
  NOR U5451 ( .A(n4554), .B(n4553), .Z(n4551) );
  XNOR U5452 ( .A(n4552), .B(n4551), .Z(n4557) );
  XOR U5453 ( .A(n4554), .B(n4553), .Z(n4555) );
  NAND U5454 ( .A(n4555), .B(n7184), .Z(n4556) );
  NAND U5455 ( .A(n4557), .B(n4556), .Z(n7189) );
  XNOR U5456 ( .A(a[428]), .B(b[428]), .Z(n7188) );
  NAND U5457 ( .A(n7189), .B(n7188), .Z(n4558) );
  NANDN U5458 ( .A(n4559), .B(n4558), .Z(n4565) );
  NAND U5459 ( .A(a[428]), .B(b[428]), .Z(n4566) );
  AND U5460 ( .A(n4565), .B(n4566), .Z(n4561) );
  XOR U5461 ( .A(a[429]), .B(b[429]), .Z(n7194) );
  ANDN U5462 ( .B(n7193), .A(n7194), .Z(n4560) );
  OR U5463 ( .A(n4561), .B(n4560), .Z(n4562) );
  AND U5464 ( .A(a[429]), .B(b[429]), .Z(n4564) );
  ANDN U5465 ( .B(n4562), .A(n4564), .Z(n4571) );
  NOR U5466 ( .A(n4566), .B(n4565), .Z(n4563) );
  XNOR U5467 ( .A(n4564), .B(n4563), .Z(n4569) );
  XOR U5468 ( .A(n4566), .B(n4565), .Z(n4567) );
  NAND U5469 ( .A(n4567), .B(n7194), .Z(n4568) );
  NAND U5470 ( .A(n4569), .B(n4568), .Z(n7199) );
  XNOR U5471 ( .A(a[430]), .B(b[430]), .Z(n7198) );
  NAND U5472 ( .A(n7199), .B(n7198), .Z(n4570) );
  NANDN U5473 ( .A(n4571), .B(n4570), .Z(n4577) );
  NAND U5474 ( .A(a[430]), .B(b[430]), .Z(n4578) );
  AND U5475 ( .A(n4577), .B(n4578), .Z(n4573) );
  XOR U5476 ( .A(a[431]), .B(b[431]), .Z(n7204) );
  ANDN U5477 ( .B(n7203), .A(n7204), .Z(n4572) );
  OR U5478 ( .A(n4573), .B(n4572), .Z(n4574) );
  AND U5479 ( .A(a[431]), .B(b[431]), .Z(n4576) );
  ANDN U5480 ( .B(n4574), .A(n4576), .Z(n4583) );
  NOR U5481 ( .A(n4578), .B(n4577), .Z(n4575) );
  XNOR U5482 ( .A(n4576), .B(n4575), .Z(n4581) );
  XOR U5483 ( .A(n4578), .B(n4577), .Z(n4579) );
  NAND U5484 ( .A(n4579), .B(n7204), .Z(n4580) );
  NAND U5485 ( .A(n4581), .B(n4580), .Z(n7209) );
  XNOR U5486 ( .A(a[432]), .B(b[432]), .Z(n7208) );
  NAND U5487 ( .A(n7209), .B(n7208), .Z(n4582) );
  NANDN U5488 ( .A(n4583), .B(n4582), .Z(n4589) );
  NAND U5489 ( .A(a[432]), .B(b[432]), .Z(n4590) );
  AND U5490 ( .A(n4589), .B(n4590), .Z(n4585) );
  XOR U5491 ( .A(a[433]), .B(b[433]), .Z(n7214) );
  ANDN U5492 ( .B(n7213), .A(n7214), .Z(n4584) );
  OR U5493 ( .A(n4585), .B(n4584), .Z(n4586) );
  AND U5494 ( .A(a[433]), .B(b[433]), .Z(n4588) );
  ANDN U5495 ( .B(n4586), .A(n4588), .Z(n4595) );
  NOR U5496 ( .A(n4590), .B(n4589), .Z(n4587) );
  XNOR U5497 ( .A(n4588), .B(n4587), .Z(n4593) );
  XOR U5498 ( .A(n4590), .B(n4589), .Z(n4591) );
  NAND U5499 ( .A(n4591), .B(n7214), .Z(n4592) );
  NAND U5500 ( .A(n4593), .B(n4592), .Z(n7219) );
  XNOR U5501 ( .A(a[434]), .B(b[434]), .Z(n7218) );
  NAND U5502 ( .A(n7219), .B(n7218), .Z(n4594) );
  NANDN U5503 ( .A(n4595), .B(n4594), .Z(n4601) );
  NAND U5504 ( .A(a[434]), .B(b[434]), .Z(n4602) );
  AND U5505 ( .A(n4601), .B(n4602), .Z(n4597) );
  XOR U5506 ( .A(a[435]), .B(b[435]), .Z(n7224) );
  ANDN U5507 ( .B(n7223), .A(n7224), .Z(n4596) );
  OR U5508 ( .A(n4597), .B(n4596), .Z(n4598) );
  AND U5509 ( .A(a[435]), .B(b[435]), .Z(n4600) );
  ANDN U5510 ( .B(n4598), .A(n4600), .Z(n4607) );
  NOR U5511 ( .A(n4602), .B(n4601), .Z(n4599) );
  XNOR U5512 ( .A(n4600), .B(n4599), .Z(n4605) );
  XOR U5513 ( .A(n4602), .B(n4601), .Z(n4603) );
  NAND U5514 ( .A(n4603), .B(n7224), .Z(n4604) );
  NAND U5515 ( .A(n4605), .B(n4604), .Z(n7229) );
  XNOR U5516 ( .A(a[436]), .B(b[436]), .Z(n7228) );
  NAND U5517 ( .A(n7229), .B(n7228), .Z(n4606) );
  NANDN U5518 ( .A(n4607), .B(n4606), .Z(n4613) );
  NAND U5519 ( .A(a[436]), .B(b[436]), .Z(n4614) );
  AND U5520 ( .A(n4613), .B(n4614), .Z(n4609) );
  XOR U5521 ( .A(a[437]), .B(b[437]), .Z(n7234) );
  ANDN U5522 ( .B(n7233), .A(n7234), .Z(n4608) );
  OR U5523 ( .A(n4609), .B(n4608), .Z(n4610) );
  AND U5524 ( .A(a[437]), .B(b[437]), .Z(n4612) );
  ANDN U5525 ( .B(n4610), .A(n4612), .Z(n4619) );
  NOR U5526 ( .A(n4614), .B(n4613), .Z(n4611) );
  XNOR U5527 ( .A(n4612), .B(n4611), .Z(n4617) );
  XOR U5528 ( .A(n4614), .B(n4613), .Z(n4615) );
  NAND U5529 ( .A(n4615), .B(n7234), .Z(n4616) );
  NAND U5530 ( .A(n4617), .B(n4616), .Z(n7239) );
  XNOR U5531 ( .A(a[438]), .B(b[438]), .Z(n7238) );
  NAND U5532 ( .A(n7239), .B(n7238), .Z(n4618) );
  NANDN U5533 ( .A(n4619), .B(n4618), .Z(n4625) );
  NAND U5534 ( .A(a[438]), .B(b[438]), .Z(n4626) );
  AND U5535 ( .A(n4625), .B(n4626), .Z(n4621) );
  XOR U5536 ( .A(a[439]), .B(b[439]), .Z(n7244) );
  ANDN U5537 ( .B(n7243), .A(n7244), .Z(n4620) );
  OR U5538 ( .A(n4621), .B(n4620), .Z(n4622) );
  AND U5539 ( .A(a[439]), .B(b[439]), .Z(n4624) );
  ANDN U5540 ( .B(n4622), .A(n4624), .Z(n4631) );
  NOR U5541 ( .A(n4626), .B(n4625), .Z(n4623) );
  XNOR U5542 ( .A(n4624), .B(n4623), .Z(n4629) );
  XOR U5543 ( .A(n4626), .B(n4625), .Z(n4627) );
  NAND U5544 ( .A(n4627), .B(n7244), .Z(n4628) );
  NAND U5545 ( .A(n4629), .B(n4628), .Z(n7249) );
  XNOR U5546 ( .A(a[440]), .B(b[440]), .Z(n7248) );
  NAND U5547 ( .A(n7249), .B(n7248), .Z(n4630) );
  NANDN U5548 ( .A(n4631), .B(n4630), .Z(n4632) );
  IV U5549 ( .A(n4632), .Z(n4636) );
  AND U5550 ( .A(a[440]), .B(b[440]), .Z(n4637) );
  NOR U5551 ( .A(n4636), .B(n4637), .Z(n4634) );
  XNOR U5552 ( .A(n4637), .B(n4632), .Z(n7254) );
  XNOR U5553 ( .A(a[441]), .B(b[441]), .Z(n7253) );
  AND U5554 ( .A(n7254), .B(n7253), .Z(n4633) );
  OR U5555 ( .A(n4634), .B(n4633), .Z(n4635) );
  AND U5556 ( .A(a[441]), .B(b[441]), .Z(n4639) );
  ANDN U5557 ( .B(n4635), .A(n4639), .Z(n4641) );
  AND U5558 ( .A(n4637), .B(n4636), .Z(n4638) );
  NAND U5559 ( .A(n4639), .B(n4638), .Z(n4644) );
  ANDN U5560 ( .B(n4644), .A(n4641), .Z(n7259) );
  XNOR U5561 ( .A(a[442]), .B(b[442]), .Z(n7258) );
  AND U5562 ( .A(n7259), .B(n7258), .Z(n4640) );
  OR U5563 ( .A(n4641), .B(n4640), .Z(n4642) );
  AND U5564 ( .A(n4643), .B(n4642), .Z(n4646) );
  XNOR U5565 ( .A(a[443]), .B(b[443]), .Z(n7263) );
  NAND U5566 ( .A(n7264), .B(n7263), .Z(n4645) );
  NANDN U5567 ( .A(n4646), .B(n4645), .Z(n4652) );
  NAND U5568 ( .A(a[443]), .B(b[443]), .Z(n4653) );
  AND U5569 ( .A(n4652), .B(n4653), .Z(n4648) );
  XOR U5570 ( .A(a[444]), .B(b[444]), .Z(n7269) );
  ANDN U5571 ( .B(n7268), .A(n7269), .Z(n4647) );
  OR U5572 ( .A(n4648), .B(n4647), .Z(n4649) );
  AND U5573 ( .A(a[444]), .B(b[444]), .Z(n4651) );
  ANDN U5574 ( .B(n4649), .A(n4651), .Z(n4658) );
  NOR U5575 ( .A(n4653), .B(n4652), .Z(n4650) );
  XNOR U5576 ( .A(n4651), .B(n4650), .Z(n4656) );
  XOR U5577 ( .A(n4653), .B(n4652), .Z(n4654) );
  NAND U5578 ( .A(n4654), .B(n7269), .Z(n4655) );
  NAND U5579 ( .A(n4656), .B(n4655), .Z(n7274) );
  XNOR U5580 ( .A(a[445]), .B(b[445]), .Z(n7273) );
  NAND U5581 ( .A(n7274), .B(n7273), .Z(n4657) );
  NANDN U5582 ( .A(n4658), .B(n4657), .Z(n4659) );
  IV U5583 ( .A(n4659), .Z(n4663) );
  AND U5584 ( .A(a[445]), .B(b[445]), .Z(n4664) );
  NOR U5585 ( .A(n4663), .B(n4664), .Z(n4661) );
  XNOR U5586 ( .A(n4664), .B(n4659), .Z(n7279) );
  XNOR U5587 ( .A(a[446]), .B(b[446]), .Z(n7278) );
  AND U5588 ( .A(n7279), .B(n7278), .Z(n4660) );
  OR U5589 ( .A(n4661), .B(n4660), .Z(n4662) );
  AND U5590 ( .A(a[446]), .B(b[446]), .Z(n4666) );
  ANDN U5591 ( .B(n4662), .A(n4666), .Z(n4668) );
  AND U5592 ( .A(n4664), .B(n4663), .Z(n4665) );
  NAND U5593 ( .A(n4666), .B(n4665), .Z(n4671) );
  ANDN U5594 ( .B(n4671), .A(n4668), .Z(n7284) );
  XNOR U5595 ( .A(a[447]), .B(b[447]), .Z(n7283) );
  AND U5596 ( .A(n7284), .B(n7283), .Z(n4667) );
  OR U5597 ( .A(n4668), .B(n4667), .Z(n4669) );
  AND U5598 ( .A(a[447]), .B(b[447]), .Z(n4670) );
  ANDN U5599 ( .B(n4669), .A(n4670), .Z(n4674) );
  NANDN U5600 ( .A(n4671), .B(n4670), .Z(n4672) );
  ANDN U5601 ( .B(n4672), .A(n4674), .Z(n7289) );
  XNOR U5602 ( .A(a[448]), .B(b[448]), .Z(n7288) );
  NAND U5603 ( .A(n7289), .B(n7288), .Z(n4673) );
  NANDN U5604 ( .A(n4674), .B(n4673), .Z(n4680) );
  NAND U5605 ( .A(a[448]), .B(b[448]), .Z(n4681) );
  AND U5606 ( .A(n4680), .B(n4681), .Z(n4676) );
  XOR U5607 ( .A(a[449]), .B(b[449]), .Z(n7294) );
  ANDN U5608 ( .B(n7293), .A(n7294), .Z(n4675) );
  OR U5609 ( .A(n4676), .B(n4675), .Z(n4677) );
  AND U5610 ( .A(a[449]), .B(b[449]), .Z(n4679) );
  ANDN U5611 ( .B(n4677), .A(n4679), .Z(n4686) );
  NOR U5612 ( .A(n4681), .B(n4680), .Z(n4678) );
  XNOR U5613 ( .A(n4679), .B(n4678), .Z(n4684) );
  XOR U5614 ( .A(n4681), .B(n4680), .Z(n4682) );
  NAND U5615 ( .A(n4682), .B(n7294), .Z(n4683) );
  NAND U5616 ( .A(n4684), .B(n4683), .Z(n7299) );
  XNOR U5617 ( .A(a[450]), .B(b[450]), .Z(n7298) );
  NAND U5618 ( .A(n7299), .B(n7298), .Z(n4685) );
  NANDN U5619 ( .A(n4686), .B(n4685), .Z(n4692) );
  NAND U5620 ( .A(a[450]), .B(b[450]), .Z(n4693) );
  AND U5621 ( .A(n4692), .B(n4693), .Z(n4688) );
  XOR U5622 ( .A(a[451]), .B(b[451]), .Z(n7304) );
  ANDN U5623 ( .B(n7303), .A(n7304), .Z(n4687) );
  OR U5624 ( .A(n4688), .B(n4687), .Z(n4689) );
  AND U5625 ( .A(a[451]), .B(b[451]), .Z(n4691) );
  ANDN U5626 ( .B(n4689), .A(n4691), .Z(n4698) );
  NOR U5627 ( .A(n4693), .B(n4692), .Z(n4690) );
  XNOR U5628 ( .A(n4691), .B(n4690), .Z(n4696) );
  XOR U5629 ( .A(n4693), .B(n4692), .Z(n4694) );
  NAND U5630 ( .A(n4694), .B(n7304), .Z(n4695) );
  NAND U5631 ( .A(n4696), .B(n4695), .Z(n7309) );
  XNOR U5632 ( .A(a[452]), .B(b[452]), .Z(n7308) );
  NAND U5633 ( .A(n7309), .B(n7308), .Z(n4697) );
  NANDN U5634 ( .A(n4698), .B(n4697), .Z(n4704) );
  NAND U5635 ( .A(a[452]), .B(b[452]), .Z(n4705) );
  AND U5636 ( .A(n4704), .B(n4705), .Z(n4700) );
  XOR U5637 ( .A(a[453]), .B(b[453]), .Z(n7314) );
  ANDN U5638 ( .B(n7313), .A(n7314), .Z(n4699) );
  OR U5639 ( .A(n4700), .B(n4699), .Z(n4701) );
  AND U5640 ( .A(a[453]), .B(b[453]), .Z(n4703) );
  ANDN U5641 ( .B(n4701), .A(n4703), .Z(n4710) );
  NOR U5642 ( .A(n4705), .B(n4704), .Z(n4702) );
  XNOR U5643 ( .A(n4703), .B(n4702), .Z(n4708) );
  XOR U5644 ( .A(n4705), .B(n4704), .Z(n4706) );
  NAND U5645 ( .A(n4706), .B(n7314), .Z(n4707) );
  NAND U5646 ( .A(n4708), .B(n4707), .Z(n7319) );
  XNOR U5647 ( .A(a[454]), .B(b[454]), .Z(n7318) );
  NAND U5648 ( .A(n7319), .B(n7318), .Z(n4709) );
  NANDN U5649 ( .A(n4710), .B(n4709), .Z(n4716) );
  NAND U5650 ( .A(a[454]), .B(b[454]), .Z(n4717) );
  AND U5651 ( .A(n4716), .B(n4717), .Z(n4712) );
  XOR U5652 ( .A(a[455]), .B(b[455]), .Z(n7324) );
  ANDN U5653 ( .B(n7323), .A(n7324), .Z(n4711) );
  OR U5654 ( .A(n4712), .B(n4711), .Z(n4713) );
  AND U5655 ( .A(a[455]), .B(b[455]), .Z(n4715) );
  ANDN U5656 ( .B(n4713), .A(n4715), .Z(n4722) );
  NOR U5657 ( .A(n4717), .B(n4716), .Z(n4714) );
  XNOR U5658 ( .A(n4715), .B(n4714), .Z(n4720) );
  XOR U5659 ( .A(n4717), .B(n4716), .Z(n4718) );
  NAND U5660 ( .A(n4718), .B(n7324), .Z(n4719) );
  NAND U5661 ( .A(n4720), .B(n4719), .Z(n7329) );
  XNOR U5662 ( .A(a[456]), .B(b[456]), .Z(n7328) );
  NAND U5663 ( .A(n7329), .B(n7328), .Z(n4721) );
  NANDN U5664 ( .A(n4722), .B(n4721), .Z(n4723) );
  IV U5665 ( .A(n4723), .Z(n4727) );
  AND U5666 ( .A(a[456]), .B(b[456]), .Z(n4728) );
  NOR U5667 ( .A(n4727), .B(n4728), .Z(n4725) );
  XNOR U5668 ( .A(n4728), .B(n4723), .Z(n7334) );
  XNOR U5669 ( .A(a[457]), .B(b[457]), .Z(n7333) );
  AND U5670 ( .A(n7334), .B(n7333), .Z(n4724) );
  OR U5671 ( .A(n4725), .B(n4724), .Z(n4726) );
  AND U5672 ( .A(a[457]), .B(b[457]), .Z(n4730) );
  ANDN U5673 ( .B(n4726), .A(n4730), .Z(n4732) );
  AND U5674 ( .A(n4728), .B(n4727), .Z(n4729) );
  NAND U5675 ( .A(n4730), .B(n4729), .Z(n4735) );
  ANDN U5676 ( .B(n4735), .A(n4732), .Z(n7339) );
  XNOR U5677 ( .A(a[458]), .B(b[458]), .Z(n7338) );
  AND U5678 ( .A(n7339), .B(n7338), .Z(n4731) );
  OR U5679 ( .A(n4732), .B(n4731), .Z(n4733) );
  AND U5680 ( .A(a[458]), .B(b[458]), .Z(n4734) );
  ANDN U5681 ( .B(n4733), .A(n4734), .Z(n4738) );
  NANDN U5682 ( .A(n4735), .B(n4734), .Z(n4736) );
  ANDN U5683 ( .B(n4736), .A(n4738), .Z(n7344) );
  XNOR U5684 ( .A(a[459]), .B(b[459]), .Z(n7343) );
  NAND U5685 ( .A(n7344), .B(n7343), .Z(n4737) );
  NANDN U5686 ( .A(n4738), .B(n4737), .Z(n4744) );
  NAND U5687 ( .A(a[459]), .B(b[459]), .Z(n4745) );
  AND U5688 ( .A(n4744), .B(n4745), .Z(n4740) );
  XOR U5689 ( .A(a[460]), .B(b[460]), .Z(n7349) );
  ANDN U5690 ( .B(n7348), .A(n7349), .Z(n4739) );
  OR U5691 ( .A(n4740), .B(n4739), .Z(n4741) );
  AND U5692 ( .A(a[460]), .B(b[460]), .Z(n4743) );
  ANDN U5693 ( .B(n4741), .A(n4743), .Z(n4750) );
  NOR U5694 ( .A(n4745), .B(n4744), .Z(n4742) );
  XNOR U5695 ( .A(n4743), .B(n4742), .Z(n4748) );
  XOR U5696 ( .A(n4745), .B(n4744), .Z(n4746) );
  NAND U5697 ( .A(n4746), .B(n7349), .Z(n4747) );
  NAND U5698 ( .A(n4748), .B(n4747), .Z(n7354) );
  XNOR U5699 ( .A(a[461]), .B(b[461]), .Z(n7353) );
  NAND U5700 ( .A(n7354), .B(n7353), .Z(n4749) );
  NANDN U5701 ( .A(n4750), .B(n4749), .Z(n4756) );
  NAND U5702 ( .A(a[461]), .B(b[461]), .Z(n4757) );
  AND U5703 ( .A(n4756), .B(n4757), .Z(n4752) );
  XOR U5704 ( .A(a[462]), .B(b[462]), .Z(n7359) );
  ANDN U5705 ( .B(n7358), .A(n7359), .Z(n4751) );
  OR U5706 ( .A(n4752), .B(n4751), .Z(n4753) );
  AND U5707 ( .A(a[462]), .B(b[462]), .Z(n4755) );
  ANDN U5708 ( .B(n4753), .A(n4755), .Z(n4762) );
  NOR U5709 ( .A(n4757), .B(n4756), .Z(n4754) );
  XNOR U5710 ( .A(n4755), .B(n4754), .Z(n4760) );
  XOR U5711 ( .A(n4757), .B(n4756), .Z(n4758) );
  NAND U5712 ( .A(n4758), .B(n7359), .Z(n4759) );
  NAND U5713 ( .A(n4760), .B(n4759), .Z(n7364) );
  XNOR U5714 ( .A(a[463]), .B(b[463]), .Z(n7363) );
  NAND U5715 ( .A(n7364), .B(n7363), .Z(n4761) );
  NANDN U5716 ( .A(n4762), .B(n4761), .Z(n4768) );
  NAND U5717 ( .A(a[463]), .B(b[463]), .Z(n4769) );
  AND U5718 ( .A(n4768), .B(n4769), .Z(n4764) );
  XOR U5719 ( .A(a[464]), .B(b[464]), .Z(n7369) );
  ANDN U5720 ( .B(n7368), .A(n7369), .Z(n4763) );
  OR U5721 ( .A(n4764), .B(n4763), .Z(n4765) );
  AND U5722 ( .A(a[464]), .B(b[464]), .Z(n4767) );
  ANDN U5723 ( .B(n4765), .A(n4767), .Z(n4774) );
  NOR U5724 ( .A(n4769), .B(n4768), .Z(n4766) );
  XNOR U5725 ( .A(n4767), .B(n4766), .Z(n4772) );
  XOR U5726 ( .A(n4769), .B(n4768), .Z(n4770) );
  NAND U5727 ( .A(n4770), .B(n7369), .Z(n4771) );
  NAND U5728 ( .A(n4772), .B(n4771), .Z(n7374) );
  XNOR U5729 ( .A(a[465]), .B(b[465]), .Z(n7373) );
  NAND U5730 ( .A(n7374), .B(n7373), .Z(n4773) );
  NANDN U5731 ( .A(n4774), .B(n4773), .Z(n4780) );
  NAND U5732 ( .A(a[465]), .B(b[465]), .Z(n4781) );
  AND U5733 ( .A(n4780), .B(n4781), .Z(n4776) );
  XOR U5734 ( .A(a[466]), .B(b[466]), .Z(n7379) );
  ANDN U5735 ( .B(n7378), .A(n7379), .Z(n4775) );
  OR U5736 ( .A(n4776), .B(n4775), .Z(n4777) );
  AND U5737 ( .A(a[466]), .B(b[466]), .Z(n4779) );
  ANDN U5738 ( .B(n4777), .A(n4779), .Z(n4786) );
  NOR U5739 ( .A(n4781), .B(n4780), .Z(n4778) );
  XNOR U5740 ( .A(n4779), .B(n4778), .Z(n4784) );
  XOR U5741 ( .A(n4781), .B(n4780), .Z(n4782) );
  NAND U5742 ( .A(n4782), .B(n7379), .Z(n4783) );
  NAND U5743 ( .A(n4784), .B(n4783), .Z(n7384) );
  XNOR U5744 ( .A(a[467]), .B(b[467]), .Z(n7383) );
  NAND U5745 ( .A(n7384), .B(n7383), .Z(n4785) );
  NANDN U5746 ( .A(n4786), .B(n4785), .Z(n4792) );
  NAND U5747 ( .A(a[467]), .B(b[467]), .Z(n4793) );
  AND U5748 ( .A(n4792), .B(n4793), .Z(n4788) );
  XOR U5749 ( .A(a[468]), .B(b[468]), .Z(n7389) );
  ANDN U5750 ( .B(n7388), .A(n7389), .Z(n4787) );
  OR U5751 ( .A(n4788), .B(n4787), .Z(n4789) );
  AND U5752 ( .A(a[468]), .B(b[468]), .Z(n4791) );
  ANDN U5753 ( .B(n4789), .A(n4791), .Z(n4798) );
  NOR U5754 ( .A(n4793), .B(n4792), .Z(n4790) );
  XNOR U5755 ( .A(n4791), .B(n4790), .Z(n4796) );
  XOR U5756 ( .A(n4793), .B(n4792), .Z(n4794) );
  NAND U5757 ( .A(n4794), .B(n7389), .Z(n4795) );
  NAND U5758 ( .A(n4796), .B(n4795), .Z(n7394) );
  XNOR U5759 ( .A(a[469]), .B(b[469]), .Z(n7393) );
  NAND U5760 ( .A(n7394), .B(n7393), .Z(n4797) );
  NANDN U5761 ( .A(n4798), .B(n4797), .Z(n4804) );
  NAND U5762 ( .A(a[469]), .B(b[469]), .Z(n4805) );
  AND U5763 ( .A(n4804), .B(n4805), .Z(n4800) );
  XOR U5764 ( .A(a[470]), .B(b[470]), .Z(n7399) );
  ANDN U5765 ( .B(n7398), .A(n7399), .Z(n4799) );
  OR U5766 ( .A(n4800), .B(n4799), .Z(n4801) );
  AND U5767 ( .A(a[470]), .B(b[470]), .Z(n4803) );
  ANDN U5768 ( .B(n4801), .A(n4803), .Z(n4810) );
  NOR U5769 ( .A(n4805), .B(n4804), .Z(n4802) );
  XNOR U5770 ( .A(n4803), .B(n4802), .Z(n4808) );
  XOR U5771 ( .A(n4805), .B(n4804), .Z(n4806) );
  NAND U5772 ( .A(n4806), .B(n7399), .Z(n4807) );
  NAND U5773 ( .A(n4808), .B(n4807), .Z(n7404) );
  XNOR U5774 ( .A(a[471]), .B(b[471]), .Z(n7403) );
  NAND U5775 ( .A(n7404), .B(n7403), .Z(n4809) );
  NANDN U5776 ( .A(n4810), .B(n4809), .Z(n4816) );
  NAND U5777 ( .A(a[471]), .B(b[471]), .Z(n4817) );
  AND U5778 ( .A(n4816), .B(n4817), .Z(n4812) );
  XOR U5779 ( .A(a[472]), .B(b[472]), .Z(n7409) );
  ANDN U5780 ( .B(n7408), .A(n7409), .Z(n4811) );
  OR U5781 ( .A(n4812), .B(n4811), .Z(n4813) );
  AND U5782 ( .A(a[472]), .B(b[472]), .Z(n4815) );
  ANDN U5783 ( .B(n4813), .A(n4815), .Z(n4822) );
  NOR U5784 ( .A(n4817), .B(n4816), .Z(n4814) );
  XNOR U5785 ( .A(n4815), .B(n4814), .Z(n4820) );
  XOR U5786 ( .A(n4817), .B(n4816), .Z(n4818) );
  NAND U5787 ( .A(n4818), .B(n7409), .Z(n4819) );
  NAND U5788 ( .A(n4820), .B(n4819), .Z(n7414) );
  XNOR U5789 ( .A(a[473]), .B(b[473]), .Z(n7413) );
  NAND U5790 ( .A(n7414), .B(n7413), .Z(n4821) );
  NANDN U5791 ( .A(n4822), .B(n4821), .Z(n4823) );
  IV U5792 ( .A(n4823), .Z(n4827) );
  AND U5793 ( .A(a[473]), .B(b[473]), .Z(n4828) );
  NOR U5794 ( .A(n4827), .B(n4828), .Z(n4825) );
  XNOR U5795 ( .A(n4828), .B(n4823), .Z(n7419) );
  XNOR U5796 ( .A(a[474]), .B(b[474]), .Z(n7418) );
  AND U5797 ( .A(n7419), .B(n7418), .Z(n4824) );
  OR U5798 ( .A(n4825), .B(n4824), .Z(n4826) );
  AND U5799 ( .A(a[474]), .B(b[474]), .Z(n4830) );
  ANDN U5800 ( .B(n4826), .A(n4830), .Z(n4832) );
  AND U5801 ( .A(n4828), .B(n4827), .Z(n4829) );
  NAND U5802 ( .A(n4830), .B(n4829), .Z(n4835) );
  ANDN U5803 ( .B(n4835), .A(n4832), .Z(n7424) );
  XNOR U5804 ( .A(a[475]), .B(b[475]), .Z(n7423) );
  AND U5805 ( .A(n7424), .B(n7423), .Z(n4831) );
  OR U5806 ( .A(n4832), .B(n4831), .Z(n4833) );
  AND U5807 ( .A(a[475]), .B(b[475]), .Z(n4834) );
  ANDN U5808 ( .B(n4833), .A(n4834), .Z(n4838) );
  NANDN U5809 ( .A(n4835), .B(n4834), .Z(n4836) );
  ANDN U5810 ( .B(n4836), .A(n4838), .Z(n7429) );
  XNOR U5811 ( .A(a[476]), .B(b[476]), .Z(n7428) );
  NAND U5812 ( .A(n7429), .B(n7428), .Z(n4837) );
  NANDN U5813 ( .A(n4838), .B(n4837), .Z(n4844) );
  NAND U5814 ( .A(a[476]), .B(b[476]), .Z(n4845) );
  AND U5815 ( .A(n4844), .B(n4845), .Z(n4840) );
  XOR U5816 ( .A(a[477]), .B(b[477]), .Z(n7434) );
  ANDN U5817 ( .B(n7433), .A(n7434), .Z(n4839) );
  OR U5818 ( .A(n4840), .B(n4839), .Z(n4841) );
  AND U5819 ( .A(a[477]), .B(b[477]), .Z(n4843) );
  ANDN U5820 ( .B(n4841), .A(n4843), .Z(n4850) );
  NOR U5821 ( .A(n4845), .B(n4844), .Z(n4842) );
  XNOR U5822 ( .A(n4843), .B(n4842), .Z(n4848) );
  XOR U5823 ( .A(n4845), .B(n4844), .Z(n4846) );
  NAND U5824 ( .A(n4846), .B(n7434), .Z(n4847) );
  NAND U5825 ( .A(n4848), .B(n4847), .Z(n7439) );
  XNOR U5826 ( .A(a[478]), .B(b[478]), .Z(n7438) );
  NAND U5827 ( .A(n7439), .B(n7438), .Z(n4849) );
  NANDN U5828 ( .A(n4850), .B(n4849), .Z(n4856) );
  NAND U5829 ( .A(a[478]), .B(b[478]), .Z(n4857) );
  AND U5830 ( .A(n4856), .B(n4857), .Z(n4852) );
  XOR U5831 ( .A(a[479]), .B(b[479]), .Z(n7444) );
  ANDN U5832 ( .B(n7443), .A(n7444), .Z(n4851) );
  OR U5833 ( .A(n4852), .B(n4851), .Z(n4853) );
  AND U5834 ( .A(a[479]), .B(b[479]), .Z(n4855) );
  ANDN U5835 ( .B(n4853), .A(n4855), .Z(n4862) );
  NOR U5836 ( .A(n4857), .B(n4856), .Z(n4854) );
  XNOR U5837 ( .A(n4855), .B(n4854), .Z(n4860) );
  XOR U5838 ( .A(n4857), .B(n4856), .Z(n4858) );
  NAND U5839 ( .A(n4858), .B(n7444), .Z(n4859) );
  NAND U5840 ( .A(n4860), .B(n4859), .Z(n7449) );
  XNOR U5841 ( .A(a[480]), .B(b[480]), .Z(n7448) );
  NAND U5842 ( .A(n7449), .B(n7448), .Z(n4861) );
  NANDN U5843 ( .A(n4862), .B(n4861), .Z(n4868) );
  NAND U5844 ( .A(a[480]), .B(b[480]), .Z(n4869) );
  AND U5845 ( .A(n4868), .B(n4869), .Z(n4864) );
  XOR U5846 ( .A(a[481]), .B(b[481]), .Z(n7454) );
  ANDN U5847 ( .B(n7453), .A(n7454), .Z(n4863) );
  OR U5848 ( .A(n4864), .B(n4863), .Z(n4865) );
  AND U5849 ( .A(a[481]), .B(b[481]), .Z(n4867) );
  ANDN U5850 ( .B(n4865), .A(n4867), .Z(n4874) );
  NOR U5851 ( .A(n4869), .B(n4868), .Z(n4866) );
  XNOR U5852 ( .A(n4867), .B(n4866), .Z(n4872) );
  XOR U5853 ( .A(n4869), .B(n4868), .Z(n4870) );
  NAND U5854 ( .A(n4870), .B(n7454), .Z(n4871) );
  NAND U5855 ( .A(n4872), .B(n4871), .Z(n7459) );
  XNOR U5856 ( .A(a[482]), .B(b[482]), .Z(n7458) );
  NAND U5857 ( .A(n7459), .B(n7458), .Z(n4873) );
  NANDN U5858 ( .A(n4874), .B(n4873), .Z(n4880) );
  NAND U5859 ( .A(a[482]), .B(b[482]), .Z(n4881) );
  AND U5860 ( .A(n4880), .B(n4881), .Z(n4876) );
  XOR U5861 ( .A(a[483]), .B(b[483]), .Z(n7464) );
  ANDN U5862 ( .B(n7463), .A(n7464), .Z(n4875) );
  OR U5863 ( .A(n4876), .B(n4875), .Z(n4877) );
  AND U5864 ( .A(a[483]), .B(b[483]), .Z(n4879) );
  ANDN U5865 ( .B(n4877), .A(n4879), .Z(n4886) );
  NOR U5866 ( .A(n4881), .B(n4880), .Z(n4878) );
  XNOR U5867 ( .A(n4879), .B(n4878), .Z(n4884) );
  XOR U5868 ( .A(n4881), .B(n4880), .Z(n4882) );
  NAND U5869 ( .A(n4882), .B(n7464), .Z(n4883) );
  NAND U5870 ( .A(n4884), .B(n4883), .Z(n7469) );
  XNOR U5871 ( .A(a[484]), .B(b[484]), .Z(n7468) );
  NAND U5872 ( .A(n7469), .B(n7468), .Z(n4885) );
  NANDN U5873 ( .A(n4886), .B(n4885), .Z(n4892) );
  NAND U5874 ( .A(a[484]), .B(b[484]), .Z(n4893) );
  AND U5875 ( .A(n4892), .B(n4893), .Z(n4888) );
  XOR U5876 ( .A(a[485]), .B(b[485]), .Z(n7474) );
  ANDN U5877 ( .B(n7473), .A(n7474), .Z(n4887) );
  OR U5878 ( .A(n4888), .B(n4887), .Z(n4889) );
  AND U5879 ( .A(a[485]), .B(b[485]), .Z(n4891) );
  ANDN U5880 ( .B(n4889), .A(n4891), .Z(n4898) );
  NOR U5881 ( .A(n4893), .B(n4892), .Z(n4890) );
  XNOR U5882 ( .A(n4891), .B(n4890), .Z(n4896) );
  XOR U5883 ( .A(n4893), .B(n4892), .Z(n4894) );
  NAND U5884 ( .A(n4894), .B(n7474), .Z(n4895) );
  NAND U5885 ( .A(n4896), .B(n4895), .Z(n7479) );
  XNOR U5886 ( .A(a[486]), .B(b[486]), .Z(n7478) );
  NAND U5887 ( .A(n7479), .B(n7478), .Z(n4897) );
  NANDN U5888 ( .A(n4898), .B(n4897), .Z(n4904) );
  NAND U5889 ( .A(a[486]), .B(b[486]), .Z(n4905) );
  AND U5890 ( .A(n4904), .B(n4905), .Z(n4900) );
  XOR U5891 ( .A(a[487]), .B(b[487]), .Z(n7484) );
  ANDN U5892 ( .B(n7483), .A(n7484), .Z(n4899) );
  OR U5893 ( .A(n4900), .B(n4899), .Z(n4901) );
  AND U5894 ( .A(a[487]), .B(b[487]), .Z(n4903) );
  ANDN U5895 ( .B(n4901), .A(n4903), .Z(n4910) );
  NOR U5896 ( .A(n4905), .B(n4904), .Z(n4902) );
  XNOR U5897 ( .A(n4903), .B(n4902), .Z(n4908) );
  XOR U5898 ( .A(n4905), .B(n4904), .Z(n4906) );
  NAND U5899 ( .A(n4906), .B(n7484), .Z(n4907) );
  NAND U5900 ( .A(n4908), .B(n4907), .Z(n7489) );
  XNOR U5901 ( .A(a[488]), .B(b[488]), .Z(n7488) );
  NAND U5902 ( .A(n7489), .B(n7488), .Z(n4909) );
  NANDN U5903 ( .A(n4910), .B(n4909), .Z(n4916) );
  NAND U5904 ( .A(a[488]), .B(b[488]), .Z(n4917) );
  AND U5905 ( .A(n4916), .B(n4917), .Z(n4912) );
  XOR U5906 ( .A(a[489]), .B(b[489]), .Z(n7494) );
  ANDN U5907 ( .B(n7493), .A(n7494), .Z(n4911) );
  OR U5908 ( .A(n4912), .B(n4911), .Z(n4913) );
  AND U5909 ( .A(a[489]), .B(b[489]), .Z(n4915) );
  ANDN U5910 ( .B(n4913), .A(n4915), .Z(n4922) );
  NOR U5911 ( .A(n4917), .B(n4916), .Z(n4914) );
  XNOR U5912 ( .A(n4915), .B(n4914), .Z(n4920) );
  XOR U5913 ( .A(n4917), .B(n4916), .Z(n4918) );
  NAND U5914 ( .A(n4918), .B(n7494), .Z(n4919) );
  NAND U5915 ( .A(n4920), .B(n4919), .Z(n7499) );
  XNOR U5916 ( .A(a[490]), .B(b[490]), .Z(n7498) );
  NAND U5917 ( .A(n7499), .B(n7498), .Z(n4921) );
  NANDN U5918 ( .A(n4922), .B(n4921), .Z(n4928) );
  NAND U5919 ( .A(a[490]), .B(b[490]), .Z(n4929) );
  AND U5920 ( .A(n4928), .B(n4929), .Z(n4924) );
  XOR U5921 ( .A(a[491]), .B(b[491]), .Z(n7504) );
  ANDN U5922 ( .B(n7503), .A(n7504), .Z(n4923) );
  OR U5923 ( .A(n4924), .B(n4923), .Z(n4925) );
  AND U5924 ( .A(a[491]), .B(b[491]), .Z(n4927) );
  ANDN U5925 ( .B(n4925), .A(n4927), .Z(n4934) );
  NOR U5926 ( .A(n4929), .B(n4928), .Z(n4926) );
  XNOR U5927 ( .A(n4927), .B(n4926), .Z(n4932) );
  XOR U5928 ( .A(n4929), .B(n4928), .Z(n4930) );
  NAND U5929 ( .A(n4930), .B(n7504), .Z(n4931) );
  NAND U5930 ( .A(n4932), .B(n4931), .Z(n7509) );
  XNOR U5931 ( .A(a[492]), .B(b[492]), .Z(n7508) );
  NAND U5932 ( .A(n7509), .B(n7508), .Z(n4933) );
  NANDN U5933 ( .A(n4934), .B(n4933), .Z(n4935) );
  IV U5934 ( .A(n4935), .Z(n4939) );
  AND U5935 ( .A(a[492]), .B(b[492]), .Z(n4940) );
  NOR U5936 ( .A(n4939), .B(n4940), .Z(n4937) );
  XNOR U5937 ( .A(n4940), .B(n4935), .Z(n7514) );
  XNOR U5938 ( .A(a[493]), .B(b[493]), .Z(n7513) );
  AND U5939 ( .A(n7514), .B(n7513), .Z(n4936) );
  OR U5940 ( .A(n4937), .B(n4936), .Z(n4938) );
  AND U5941 ( .A(a[493]), .B(b[493]), .Z(n4942) );
  ANDN U5942 ( .B(n4938), .A(n4942), .Z(n4944) );
  AND U5943 ( .A(n4940), .B(n4939), .Z(n4941) );
  NAND U5944 ( .A(n4942), .B(n4941), .Z(n4947) );
  ANDN U5945 ( .B(n4947), .A(n4944), .Z(n7519) );
  XNOR U5946 ( .A(a[494]), .B(b[494]), .Z(n7518) );
  AND U5947 ( .A(n7519), .B(n7518), .Z(n4943) );
  OR U5948 ( .A(n4944), .B(n4943), .Z(n4945) );
  AND U5949 ( .A(a[494]), .B(b[494]), .Z(n4946) );
  ANDN U5950 ( .B(n4945), .A(n4946), .Z(n4950) );
  NANDN U5951 ( .A(n4947), .B(n4946), .Z(n4948) );
  ANDN U5952 ( .B(n4948), .A(n4950), .Z(n7524) );
  XNOR U5953 ( .A(a[495]), .B(b[495]), .Z(n7523) );
  NAND U5954 ( .A(n7524), .B(n7523), .Z(n4949) );
  NANDN U5955 ( .A(n4950), .B(n4949), .Z(n4956) );
  NAND U5956 ( .A(a[495]), .B(b[495]), .Z(n4957) );
  AND U5957 ( .A(n4956), .B(n4957), .Z(n4952) );
  XOR U5958 ( .A(a[496]), .B(b[496]), .Z(n7529) );
  ANDN U5959 ( .B(n7528), .A(n7529), .Z(n4951) );
  OR U5960 ( .A(n4952), .B(n4951), .Z(n4953) );
  AND U5961 ( .A(a[496]), .B(b[496]), .Z(n4955) );
  ANDN U5962 ( .B(n4953), .A(n4955), .Z(n4962) );
  NOR U5963 ( .A(n4957), .B(n4956), .Z(n4954) );
  XNOR U5964 ( .A(n4955), .B(n4954), .Z(n4960) );
  XOR U5965 ( .A(n4957), .B(n4956), .Z(n4958) );
  NAND U5966 ( .A(n4958), .B(n7529), .Z(n4959) );
  NAND U5967 ( .A(n4960), .B(n4959), .Z(n7534) );
  XNOR U5968 ( .A(a[497]), .B(b[497]), .Z(n7533) );
  NAND U5969 ( .A(n7534), .B(n7533), .Z(n4961) );
  NANDN U5970 ( .A(n4962), .B(n4961), .Z(n4968) );
  NAND U5971 ( .A(a[497]), .B(b[497]), .Z(n4969) );
  AND U5972 ( .A(n4968), .B(n4969), .Z(n4964) );
  XOR U5973 ( .A(a[498]), .B(b[498]), .Z(n7539) );
  ANDN U5974 ( .B(n7538), .A(n7539), .Z(n4963) );
  OR U5975 ( .A(n4964), .B(n4963), .Z(n4965) );
  AND U5976 ( .A(a[498]), .B(b[498]), .Z(n4967) );
  ANDN U5977 ( .B(n4965), .A(n4967), .Z(n4974) );
  NOR U5978 ( .A(n4969), .B(n4968), .Z(n4966) );
  XNOR U5979 ( .A(n4967), .B(n4966), .Z(n4972) );
  XOR U5980 ( .A(n4969), .B(n4968), .Z(n4970) );
  NAND U5981 ( .A(n4970), .B(n7539), .Z(n4971) );
  NAND U5982 ( .A(n4972), .B(n4971), .Z(n7544) );
  XNOR U5983 ( .A(a[499]), .B(b[499]), .Z(n7543) );
  NAND U5984 ( .A(n7544), .B(n7543), .Z(n4973) );
  NANDN U5985 ( .A(n4974), .B(n4973), .Z(n4980) );
  NAND U5986 ( .A(a[499]), .B(b[499]), .Z(n4981) );
  AND U5987 ( .A(n4980), .B(n4981), .Z(n4976) );
  XOR U5988 ( .A(a[500]), .B(b[500]), .Z(n7549) );
  ANDN U5989 ( .B(n7548), .A(n7549), .Z(n4975) );
  OR U5990 ( .A(n4976), .B(n4975), .Z(n4977) );
  AND U5991 ( .A(a[500]), .B(b[500]), .Z(n4979) );
  ANDN U5992 ( .B(n4977), .A(n4979), .Z(n4986) );
  NOR U5993 ( .A(n4981), .B(n4980), .Z(n4978) );
  XNOR U5994 ( .A(n4979), .B(n4978), .Z(n4984) );
  XOR U5995 ( .A(n4981), .B(n4980), .Z(n4982) );
  NAND U5996 ( .A(n4982), .B(n7549), .Z(n4983) );
  NAND U5997 ( .A(n4984), .B(n4983), .Z(n7554) );
  XNOR U5998 ( .A(a[501]), .B(b[501]), .Z(n7553) );
  NAND U5999 ( .A(n7554), .B(n7553), .Z(n4985) );
  NANDN U6000 ( .A(n4986), .B(n4985), .Z(n4992) );
  NAND U6001 ( .A(a[501]), .B(b[501]), .Z(n4993) );
  AND U6002 ( .A(n4992), .B(n4993), .Z(n4988) );
  XOR U6003 ( .A(a[502]), .B(b[502]), .Z(n7559) );
  ANDN U6004 ( .B(n7558), .A(n7559), .Z(n4987) );
  OR U6005 ( .A(n4988), .B(n4987), .Z(n4989) );
  AND U6006 ( .A(a[502]), .B(b[502]), .Z(n4991) );
  ANDN U6007 ( .B(n4989), .A(n4991), .Z(n4998) );
  NOR U6008 ( .A(n4993), .B(n4992), .Z(n4990) );
  XNOR U6009 ( .A(n4991), .B(n4990), .Z(n4996) );
  XOR U6010 ( .A(n4993), .B(n4992), .Z(n4994) );
  NAND U6011 ( .A(n4994), .B(n7559), .Z(n4995) );
  NAND U6012 ( .A(n4996), .B(n4995), .Z(n7564) );
  XNOR U6013 ( .A(a[503]), .B(b[503]), .Z(n7563) );
  NAND U6014 ( .A(n7564), .B(n7563), .Z(n4997) );
  NANDN U6015 ( .A(n4998), .B(n4997), .Z(n5004) );
  NAND U6016 ( .A(a[503]), .B(b[503]), .Z(n5005) );
  AND U6017 ( .A(n5004), .B(n5005), .Z(n5000) );
  XOR U6018 ( .A(a[504]), .B(b[504]), .Z(n7569) );
  ANDN U6019 ( .B(n7568), .A(n7569), .Z(n4999) );
  OR U6020 ( .A(n5000), .B(n4999), .Z(n5001) );
  AND U6021 ( .A(a[504]), .B(b[504]), .Z(n5003) );
  ANDN U6022 ( .B(n5001), .A(n5003), .Z(n5010) );
  NOR U6023 ( .A(n5005), .B(n5004), .Z(n5002) );
  XNOR U6024 ( .A(n5003), .B(n5002), .Z(n5008) );
  XOR U6025 ( .A(n5005), .B(n5004), .Z(n5006) );
  NAND U6026 ( .A(n5006), .B(n7569), .Z(n5007) );
  NAND U6027 ( .A(n5008), .B(n5007), .Z(n7574) );
  XNOR U6028 ( .A(a[505]), .B(b[505]), .Z(n7573) );
  NAND U6029 ( .A(n7574), .B(n7573), .Z(n5009) );
  NANDN U6030 ( .A(n5010), .B(n5009), .Z(n5016) );
  NAND U6031 ( .A(a[505]), .B(b[505]), .Z(n5017) );
  AND U6032 ( .A(n5016), .B(n5017), .Z(n5012) );
  XOR U6033 ( .A(a[506]), .B(b[506]), .Z(n7579) );
  ANDN U6034 ( .B(n7578), .A(n7579), .Z(n5011) );
  OR U6035 ( .A(n5012), .B(n5011), .Z(n5013) );
  AND U6036 ( .A(a[506]), .B(b[506]), .Z(n5015) );
  ANDN U6037 ( .B(n5013), .A(n5015), .Z(n5022) );
  NOR U6038 ( .A(n5017), .B(n5016), .Z(n5014) );
  XNOR U6039 ( .A(n5015), .B(n5014), .Z(n5020) );
  XOR U6040 ( .A(n5017), .B(n5016), .Z(n5018) );
  NAND U6041 ( .A(n5018), .B(n7579), .Z(n5019) );
  NAND U6042 ( .A(n5020), .B(n5019), .Z(n7584) );
  XNOR U6043 ( .A(a[507]), .B(b[507]), .Z(n7583) );
  NAND U6044 ( .A(n7584), .B(n7583), .Z(n5021) );
  NANDN U6045 ( .A(n5022), .B(n5021), .Z(n5028) );
  NAND U6046 ( .A(a[507]), .B(b[507]), .Z(n5029) );
  AND U6047 ( .A(n5028), .B(n5029), .Z(n5024) );
  XOR U6048 ( .A(a[508]), .B(b[508]), .Z(n7589) );
  ANDN U6049 ( .B(n7588), .A(n7589), .Z(n5023) );
  OR U6050 ( .A(n5024), .B(n5023), .Z(n5025) );
  AND U6051 ( .A(a[508]), .B(b[508]), .Z(n5027) );
  ANDN U6052 ( .B(n5025), .A(n5027), .Z(n5034) );
  NOR U6053 ( .A(n5029), .B(n5028), .Z(n5026) );
  XNOR U6054 ( .A(n5027), .B(n5026), .Z(n5032) );
  XOR U6055 ( .A(n5029), .B(n5028), .Z(n5030) );
  NAND U6056 ( .A(n5030), .B(n7589), .Z(n5031) );
  NAND U6057 ( .A(n5032), .B(n5031), .Z(n7594) );
  XNOR U6058 ( .A(a[509]), .B(b[509]), .Z(n7593) );
  NAND U6059 ( .A(n7594), .B(n7593), .Z(n5033) );
  NANDN U6060 ( .A(n5034), .B(n5033), .Z(n5040) );
  NOR U6061 ( .A(n5039), .B(n5040), .Z(n5035) );
  XOR U6062 ( .A(n5044), .B(n5035), .Z(n5038) );
  XNOR U6063 ( .A(a[510]), .B(b[510]), .Z(n7599) );
  XOR U6064 ( .A(n5039), .B(n5040), .Z(n5036) );
  NANDN U6065 ( .A(n7599), .B(n5036), .Z(n5037) );
  NAND U6066 ( .A(n5038), .B(n5037), .Z(n7604) );
  XNOR U6067 ( .A(a[511]), .B(b[511]), .Z(n7603) );
  NAND U6068 ( .A(n7604), .B(n7603), .Z(n5046) );
  AND U6069 ( .A(n5040), .B(n5039), .Z(n5042) );
  AND U6070 ( .A(n7598), .B(n7599), .Z(n5041) );
  OR U6071 ( .A(n5042), .B(n5041), .Z(n5043) );
  AND U6072 ( .A(n5044), .B(n5043), .Z(n5045) );
  ANDN U6073 ( .B(n5046), .A(n5045), .Z(n5047) );
  XOR U6074 ( .A(n5048), .B(n5047), .Z(N1026) );
  AND U6075 ( .A(n5048), .B(n5047), .Z(N1027) );
  NAND U6077 ( .A(c[0]), .B(rst), .Z(n5052) );
  XOR U6078 ( .A(n5049), .B(carry_on[0]), .Z(n5050) );
  NANDN U6079 ( .A(rst), .B(n5050), .Z(n5051) );
  NAND U6080 ( .A(n5052), .B(n5051), .Z(n1537) );
  NAND U6081 ( .A(c[1]), .B(rst), .Z(n5057) );
  XOR U6082 ( .A(n5054), .B(n5053), .Z(n5055) );
  NANDN U6083 ( .A(rst), .B(n5055), .Z(n5056) );
  NAND U6084 ( .A(n5057), .B(n5056), .Z(n1538) );
  NAND U6085 ( .A(c[2]), .B(rst), .Z(n5062) );
  XNOR U6086 ( .A(n5059), .B(n5058), .Z(n5060) );
  NANDN U6087 ( .A(rst), .B(n5060), .Z(n5061) );
  NAND U6088 ( .A(n5062), .B(n5061), .Z(n1539) );
  NAND U6089 ( .A(c[3]), .B(rst), .Z(n5067) );
  XOR U6090 ( .A(n5064), .B(n5063), .Z(n5065) );
  NANDN U6091 ( .A(rst), .B(n5065), .Z(n5066) );
  NAND U6092 ( .A(n5067), .B(n5066), .Z(n1540) );
  NAND U6093 ( .A(c[4]), .B(rst), .Z(n5072) );
  XNOR U6094 ( .A(n5069), .B(n5068), .Z(n5070) );
  NANDN U6095 ( .A(rst), .B(n5070), .Z(n5071) );
  NAND U6096 ( .A(n5072), .B(n5071), .Z(n1541) );
  NAND U6097 ( .A(c[5]), .B(rst), .Z(n5077) );
  XNOR U6098 ( .A(n5074), .B(n5073), .Z(n5075) );
  NANDN U6099 ( .A(rst), .B(n5075), .Z(n5076) );
  NAND U6100 ( .A(n5077), .B(n5076), .Z(n1542) );
  NAND U6101 ( .A(c[6]), .B(rst), .Z(n5082) );
  XNOR U6102 ( .A(n5079), .B(n5078), .Z(n5080) );
  NANDN U6103 ( .A(rst), .B(n5080), .Z(n5081) );
  NAND U6104 ( .A(n5082), .B(n5081), .Z(n1543) );
  NAND U6105 ( .A(c[7]), .B(rst), .Z(n5087) );
  XNOR U6106 ( .A(n5084), .B(n5083), .Z(n5085) );
  NANDN U6107 ( .A(rst), .B(n5085), .Z(n5086) );
  NAND U6108 ( .A(n5087), .B(n5086), .Z(n1544) );
  NAND U6109 ( .A(c[8]), .B(rst), .Z(n5092) );
  XOR U6110 ( .A(n5089), .B(n5088), .Z(n5090) );
  NANDN U6111 ( .A(rst), .B(n5090), .Z(n5091) );
  NAND U6112 ( .A(n5092), .B(n5091), .Z(n1545) );
  NAND U6113 ( .A(c[9]), .B(rst), .Z(n5097) );
  XNOR U6114 ( .A(n5094), .B(n5093), .Z(n5095) );
  NANDN U6115 ( .A(rst), .B(n5095), .Z(n5096) );
  NAND U6116 ( .A(n5097), .B(n5096), .Z(n1546) );
  NAND U6117 ( .A(c[10]), .B(rst), .Z(n5102) );
  XOR U6118 ( .A(n5099), .B(n5098), .Z(n5100) );
  NANDN U6119 ( .A(rst), .B(n5100), .Z(n5101) );
  NAND U6120 ( .A(n5102), .B(n5101), .Z(n1547) );
  NAND U6121 ( .A(c[11]), .B(rst), .Z(n5107) );
  XNOR U6122 ( .A(n5104), .B(n5103), .Z(n5105) );
  NANDN U6123 ( .A(rst), .B(n5105), .Z(n5106) );
  NAND U6124 ( .A(n5107), .B(n5106), .Z(n1548) );
  NAND U6125 ( .A(c[12]), .B(rst), .Z(n5112) );
  XOR U6126 ( .A(n5109), .B(n5108), .Z(n5110) );
  NANDN U6127 ( .A(rst), .B(n5110), .Z(n5111) );
  NAND U6128 ( .A(n5112), .B(n5111), .Z(n1549) );
  NAND U6129 ( .A(c[13]), .B(rst), .Z(n5117) );
  XNOR U6130 ( .A(n5114), .B(n5113), .Z(n5115) );
  NANDN U6131 ( .A(rst), .B(n5115), .Z(n5116) );
  NAND U6132 ( .A(n5117), .B(n5116), .Z(n1550) );
  NAND U6133 ( .A(c[14]), .B(rst), .Z(n5122) );
  XOR U6134 ( .A(n5119), .B(n5118), .Z(n5120) );
  NANDN U6135 ( .A(rst), .B(n5120), .Z(n5121) );
  NAND U6136 ( .A(n5122), .B(n5121), .Z(n1551) );
  NAND U6137 ( .A(c[15]), .B(rst), .Z(n5127) );
  XNOR U6138 ( .A(n5124), .B(n5123), .Z(n5125) );
  NANDN U6139 ( .A(rst), .B(n5125), .Z(n5126) );
  NAND U6140 ( .A(n5127), .B(n5126), .Z(n1552) );
  NAND U6141 ( .A(c[16]), .B(rst), .Z(n5132) );
  XOR U6142 ( .A(n5129), .B(n5128), .Z(n5130) );
  NANDN U6143 ( .A(rst), .B(n5130), .Z(n5131) );
  NAND U6144 ( .A(n5132), .B(n5131), .Z(n1553) );
  NAND U6145 ( .A(c[17]), .B(rst), .Z(n5137) );
  XNOR U6146 ( .A(n5134), .B(n5133), .Z(n5135) );
  NANDN U6147 ( .A(rst), .B(n5135), .Z(n5136) );
  NAND U6148 ( .A(n5137), .B(n5136), .Z(n1554) );
  NAND U6149 ( .A(c[18]), .B(rst), .Z(n5142) );
  XOR U6150 ( .A(n5139), .B(n5138), .Z(n5140) );
  NANDN U6151 ( .A(rst), .B(n5140), .Z(n5141) );
  NAND U6152 ( .A(n5142), .B(n5141), .Z(n1555) );
  NAND U6153 ( .A(c[19]), .B(rst), .Z(n5147) );
  XNOR U6154 ( .A(n5144), .B(n5143), .Z(n5145) );
  NANDN U6155 ( .A(rst), .B(n5145), .Z(n5146) );
  NAND U6156 ( .A(n5147), .B(n5146), .Z(n1556) );
  NAND U6157 ( .A(c[20]), .B(rst), .Z(n5152) );
  XOR U6158 ( .A(n5149), .B(n5148), .Z(n5150) );
  NANDN U6159 ( .A(rst), .B(n5150), .Z(n5151) );
  NAND U6160 ( .A(n5152), .B(n5151), .Z(n1557) );
  NAND U6161 ( .A(c[21]), .B(rst), .Z(n5157) );
  XNOR U6162 ( .A(n5154), .B(n5153), .Z(n5155) );
  NANDN U6163 ( .A(rst), .B(n5155), .Z(n5156) );
  NAND U6164 ( .A(n5157), .B(n5156), .Z(n1558) );
  NAND U6165 ( .A(c[22]), .B(rst), .Z(n5162) );
  XNOR U6166 ( .A(n5159), .B(n5158), .Z(n5160) );
  NANDN U6167 ( .A(rst), .B(n5160), .Z(n5161) );
  NAND U6168 ( .A(n5162), .B(n5161), .Z(n1559) );
  NAND U6169 ( .A(c[23]), .B(rst), .Z(n5167) );
  XNOR U6170 ( .A(n5164), .B(n5163), .Z(n5165) );
  NANDN U6171 ( .A(rst), .B(n5165), .Z(n5166) );
  NAND U6172 ( .A(n5167), .B(n5166), .Z(n1560) );
  NAND U6173 ( .A(c[24]), .B(rst), .Z(n5172) );
  XNOR U6174 ( .A(n5169), .B(n5168), .Z(n5170) );
  NANDN U6175 ( .A(rst), .B(n5170), .Z(n5171) );
  NAND U6176 ( .A(n5172), .B(n5171), .Z(n1561) );
  NAND U6177 ( .A(c[25]), .B(rst), .Z(n5177) );
  XOR U6178 ( .A(n5174), .B(n5173), .Z(n5175) );
  NANDN U6179 ( .A(rst), .B(n5175), .Z(n5176) );
  NAND U6180 ( .A(n5177), .B(n5176), .Z(n1562) );
  NAND U6181 ( .A(c[26]), .B(rst), .Z(n5182) );
  XNOR U6182 ( .A(n5179), .B(n5178), .Z(n5180) );
  NANDN U6183 ( .A(rst), .B(n5180), .Z(n5181) );
  NAND U6184 ( .A(n5182), .B(n5181), .Z(n1563) );
  NAND U6185 ( .A(c[27]), .B(rst), .Z(n5187) );
  XOR U6186 ( .A(n5184), .B(n5183), .Z(n5185) );
  NANDN U6187 ( .A(rst), .B(n5185), .Z(n5186) );
  NAND U6188 ( .A(n5187), .B(n5186), .Z(n1564) );
  NAND U6189 ( .A(c[28]), .B(rst), .Z(n5192) );
  XNOR U6190 ( .A(n5189), .B(n5188), .Z(n5190) );
  NANDN U6191 ( .A(rst), .B(n5190), .Z(n5191) );
  NAND U6192 ( .A(n5192), .B(n5191), .Z(n1565) );
  NAND U6193 ( .A(c[29]), .B(rst), .Z(n5197) );
  XNOR U6194 ( .A(n5194), .B(n5193), .Z(n5195) );
  NANDN U6195 ( .A(rst), .B(n5195), .Z(n5196) );
  NAND U6196 ( .A(n5197), .B(n5196), .Z(n1566) );
  NAND U6197 ( .A(c[30]), .B(rst), .Z(n5202) );
  XNOR U6198 ( .A(n5199), .B(n5198), .Z(n5200) );
  NANDN U6199 ( .A(rst), .B(n5200), .Z(n5201) );
  NAND U6200 ( .A(n5202), .B(n5201), .Z(n1567) );
  NAND U6201 ( .A(c[31]), .B(rst), .Z(n5207) );
  XNOR U6202 ( .A(n5204), .B(n5203), .Z(n5205) );
  NANDN U6203 ( .A(rst), .B(n5205), .Z(n5206) );
  NAND U6204 ( .A(n5207), .B(n5206), .Z(n1568) );
  NAND U6205 ( .A(c[32]), .B(rst), .Z(n5212) );
  XOR U6206 ( .A(n5209), .B(n5208), .Z(n5210) );
  NANDN U6207 ( .A(rst), .B(n5210), .Z(n5211) );
  NAND U6208 ( .A(n5212), .B(n5211), .Z(n1569) );
  NAND U6209 ( .A(c[33]), .B(rst), .Z(n5217) );
  XNOR U6210 ( .A(n5214), .B(n5213), .Z(n5215) );
  NANDN U6211 ( .A(rst), .B(n5215), .Z(n5216) );
  NAND U6212 ( .A(n5217), .B(n5216), .Z(n1570) );
  NAND U6213 ( .A(c[34]), .B(rst), .Z(n5222) );
  XOR U6214 ( .A(n5219), .B(n5218), .Z(n5220) );
  NANDN U6215 ( .A(rst), .B(n5220), .Z(n5221) );
  NAND U6216 ( .A(n5222), .B(n5221), .Z(n1571) );
  NAND U6217 ( .A(c[35]), .B(rst), .Z(n5227) );
  XNOR U6218 ( .A(n5224), .B(n5223), .Z(n5225) );
  NANDN U6219 ( .A(rst), .B(n5225), .Z(n5226) );
  NAND U6220 ( .A(n5227), .B(n5226), .Z(n1572) );
  NAND U6221 ( .A(c[36]), .B(rst), .Z(n5232) );
  XOR U6222 ( .A(n5229), .B(n5228), .Z(n5230) );
  NANDN U6223 ( .A(rst), .B(n5230), .Z(n5231) );
  NAND U6224 ( .A(n5232), .B(n5231), .Z(n1573) );
  NAND U6225 ( .A(c[37]), .B(rst), .Z(n5237) );
  XNOR U6226 ( .A(n5234), .B(n5233), .Z(n5235) );
  NANDN U6227 ( .A(rst), .B(n5235), .Z(n5236) );
  NAND U6228 ( .A(n5237), .B(n5236), .Z(n1574) );
  NAND U6229 ( .A(c[38]), .B(rst), .Z(n5242) );
  XOR U6230 ( .A(n5239), .B(n5238), .Z(n5240) );
  NANDN U6231 ( .A(rst), .B(n5240), .Z(n5241) );
  NAND U6232 ( .A(n5242), .B(n5241), .Z(n1575) );
  NAND U6233 ( .A(c[39]), .B(rst), .Z(n5247) );
  XNOR U6234 ( .A(n5244), .B(n5243), .Z(n5245) );
  NANDN U6235 ( .A(rst), .B(n5245), .Z(n5246) );
  NAND U6236 ( .A(n5247), .B(n5246), .Z(n1576) );
  NAND U6237 ( .A(c[40]), .B(rst), .Z(n5252) );
  XOR U6238 ( .A(n5249), .B(n5248), .Z(n5250) );
  NANDN U6239 ( .A(rst), .B(n5250), .Z(n5251) );
  NAND U6240 ( .A(n5252), .B(n5251), .Z(n1577) );
  NAND U6241 ( .A(c[41]), .B(rst), .Z(n5257) );
  XNOR U6242 ( .A(n5254), .B(n5253), .Z(n5255) );
  NANDN U6243 ( .A(rst), .B(n5255), .Z(n5256) );
  NAND U6244 ( .A(n5257), .B(n5256), .Z(n1578) );
  NAND U6245 ( .A(c[42]), .B(rst), .Z(n5262) );
  XOR U6246 ( .A(n5259), .B(n5258), .Z(n5260) );
  NANDN U6247 ( .A(rst), .B(n5260), .Z(n5261) );
  NAND U6248 ( .A(n5262), .B(n5261), .Z(n1579) );
  NAND U6249 ( .A(c[43]), .B(rst), .Z(n5267) );
  XNOR U6250 ( .A(n5264), .B(n5263), .Z(n5265) );
  NANDN U6251 ( .A(rst), .B(n5265), .Z(n5266) );
  NAND U6252 ( .A(n5267), .B(n5266), .Z(n1580) );
  NAND U6253 ( .A(c[44]), .B(rst), .Z(n5272) );
  XOR U6254 ( .A(n5269), .B(n5268), .Z(n5270) );
  NANDN U6255 ( .A(rst), .B(n5270), .Z(n5271) );
  NAND U6256 ( .A(n5272), .B(n5271), .Z(n1581) );
  NAND U6257 ( .A(c[45]), .B(rst), .Z(n5277) );
  XNOR U6258 ( .A(n5274), .B(n5273), .Z(n5275) );
  NANDN U6259 ( .A(rst), .B(n5275), .Z(n5276) );
  NAND U6260 ( .A(n5277), .B(n5276), .Z(n1582) );
  NAND U6261 ( .A(c[46]), .B(rst), .Z(n5282) );
  XOR U6262 ( .A(n5279), .B(n5278), .Z(n5280) );
  NANDN U6263 ( .A(rst), .B(n5280), .Z(n5281) );
  NAND U6264 ( .A(n5282), .B(n5281), .Z(n1583) );
  NAND U6265 ( .A(c[47]), .B(rst), .Z(n5287) );
  XNOR U6266 ( .A(n5284), .B(n5283), .Z(n5285) );
  NANDN U6267 ( .A(rst), .B(n5285), .Z(n5286) );
  NAND U6268 ( .A(n5287), .B(n5286), .Z(n1584) );
  NAND U6269 ( .A(c[48]), .B(rst), .Z(n5292) );
  XOR U6270 ( .A(n5289), .B(n5288), .Z(n5290) );
  NANDN U6271 ( .A(rst), .B(n5290), .Z(n5291) );
  NAND U6272 ( .A(n5292), .B(n5291), .Z(n1585) );
  NAND U6273 ( .A(c[49]), .B(rst), .Z(n5297) );
  XNOR U6274 ( .A(n5294), .B(n5293), .Z(n5295) );
  NANDN U6275 ( .A(rst), .B(n5295), .Z(n5296) );
  NAND U6276 ( .A(n5297), .B(n5296), .Z(n1586) );
  NAND U6277 ( .A(c[50]), .B(rst), .Z(n5302) );
  XOR U6278 ( .A(n5299), .B(n5298), .Z(n5300) );
  NANDN U6279 ( .A(rst), .B(n5300), .Z(n5301) );
  NAND U6280 ( .A(n5302), .B(n5301), .Z(n1587) );
  NAND U6281 ( .A(c[51]), .B(rst), .Z(n5307) );
  XNOR U6282 ( .A(n5304), .B(n5303), .Z(n5305) );
  NANDN U6283 ( .A(rst), .B(n5305), .Z(n5306) );
  NAND U6284 ( .A(n5307), .B(n5306), .Z(n1588) );
  NAND U6285 ( .A(c[52]), .B(rst), .Z(n5312) );
  XOR U6286 ( .A(n5309), .B(n5308), .Z(n5310) );
  NANDN U6287 ( .A(rst), .B(n5310), .Z(n5311) );
  NAND U6288 ( .A(n5312), .B(n5311), .Z(n1589) );
  NAND U6289 ( .A(c[53]), .B(rst), .Z(n5317) );
  XNOR U6290 ( .A(n5314), .B(n5313), .Z(n5315) );
  NANDN U6291 ( .A(rst), .B(n5315), .Z(n5316) );
  NAND U6292 ( .A(n5317), .B(n5316), .Z(n1590) );
  NAND U6293 ( .A(c[54]), .B(rst), .Z(n5322) );
  XOR U6294 ( .A(n5319), .B(n5318), .Z(n5320) );
  NANDN U6295 ( .A(rst), .B(n5320), .Z(n5321) );
  NAND U6296 ( .A(n5322), .B(n5321), .Z(n1591) );
  NAND U6297 ( .A(c[55]), .B(rst), .Z(n5327) );
  XNOR U6298 ( .A(n5324), .B(n5323), .Z(n5325) );
  NANDN U6299 ( .A(rst), .B(n5325), .Z(n5326) );
  NAND U6300 ( .A(n5327), .B(n5326), .Z(n1592) );
  NAND U6301 ( .A(c[56]), .B(rst), .Z(n5332) );
  XOR U6302 ( .A(n5329), .B(n5328), .Z(n5330) );
  NANDN U6303 ( .A(rst), .B(n5330), .Z(n5331) );
  NAND U6304 ( .A(n5332), .B(n5331), .Z(n1593) );
  NAND U6305 ( .A(c[57]), .B(rst), .Z(n5337) );
  XNOR U6306 ( .A(n5334), .B(n5333), .Z(n5335) );
  NANDN U6307 ( .A(rst), .B(n5335), .Z(n5336) );
  NAND U6308 ( .A(n5337), .B(n5336), .Z(n1594) );
  NAND U6309 ( .A(c[58]), .B(rst), .Z(n5342) );
  XOR U6310 ( .A(n5339), .B(n5338), .Z(n5340) );
  NANDN U6311 ( .A(rst), .B(n5340), .Z(n5341) );
  NAND U6312 ( .A(n5342), .B(n5341), .Z(n1595) );
  NAND U6313 ( .A(c[59]), .B(rst), .Z(n5347) );
  XNOR U6314 ( .A(n5344), .B(n5343), .Z(n5345) );
  NANDN U6315 ( .A(rst), .B(n5345), .Z(n5346) );
  NAND U6316 ( .A(n5347), .B(n5346), .Z(n1596) );
  NAND U6317 ( .A(c[60]), .B(rst), .Z(n5352) );
  XOR U6318 ( .A(n5349), .B(n5348), .Z(n5350) );
  NANDN U6319 ( .A(rst), .B(n5350), .Z(n5351) );
  NAND U6320 ( .A(n5352), .B(n5351), .Z(n1597) );
  NAND U6321 ( .A(c[61]), .B(rst), .Z(n5357) );
  XNOR U6322 ( .A(n5354), .B(n5353), .Z(n5355) );
  NANDN U6323 ( .A(rst), .B(n5355), .Z(n5356) );
  NAND U6324 ( .A(n5357), .B(n5356), .Z(n1598) );
  NAND U6325 ( .A(c[62]), .B(rst), .Z(n5362) );
  XOR U6326 ( .A(n5359), .B(n5358), .Z(n5360) );
  NANDN U6327 ( .A(rst), .B(n5360), .Z(n5361) );
  NAND U6328 ( .A(n5362), .B(n5361), .Z(n1599) );
  NAND U6329 ( .A(c[63]), .B(rst), .Z(n5367) );
  XNOR U6330 ( .A(n5364), .B(n5363), .Z(n5365) );
  NANDN U6331 ( .A(rst), .B(n5365), .Z(n5366) );
  NAND U6332 ( .A(n5367), .B(n5366), .Z(n1600) );
  NAND U6333 ( .A(c[64]), .B(rst), .Z(n5372) );
  XOR U6334 ( .A(n5369), .B(n5368), .Z(n5370) );
  NANDN U6335 ( .A(rst), .B(n5370), .Z(n5371) );
  NAND U6336 ( .A(n5372), .B(n5371), .Z(n1601) );
  NAND U6337 ( .A(c[65]), .B(rst), .Z(n5377) );
  XNOR U6338 ( .A(n5374), .B(n5373), .Z(n5375) );
  NANDN U6339 ( .A(rst), .B(n5375), .Z(n5376) );
  NAND U6340 ( .A(n5377), .B(n5376), .Z(n1602) );
  NAND U6341 ( .A(c[66]), .B(rst), .Z(n5382) );
  XOR U6342 ( .A(n5379), .B(n5378), .Z(n5380) );
  NANDN U6343 ( .A(rst), .B(n5380), .Z(n5381) );
  NAND U6344 ( .A(n5382), .B(n5381), .Z(n1603) );
  NAND U6345 ( .A(c[67]), .B(rst), .Z(n5387) );
  XNOR U6346 ( .A(n5384), .B(n5383), .Z(n5385) );
  NANDN U6347 ( .A(rst), .B(n5385), .Z(n5386) );
  NAND U6348 ( .A(n5387), .B(n5386), .Z(n1604) );
  NAND U6349 ( .A(c[68]), .B(rst), .Z(n5392) );
  XOR U6350 ( .A(n5389), .B(n5388), .Z(n5390) );
  NANDN U6351 ( .A(rst), .B(n5390), .Z(n5391) );
  NAND U6352 ( .A(n5392), .B(n5391), .Z(n1605) );
  NAND U6353 ( .A(c[69]), .B(rst), .Z(n5397) );
  XNOR U6354 ( .A(n5394), .B(n5393), .Z(n5395) );
  NANDN U6355 ( .A(rst), .B(n5395), .Z(n5396) );
  NAND U6356 ( .A(n5397), .B(n5396), .Z(n1606) );
  NAND U6357 ( .A(c[70]), .B(rst), .Z(n5402) );
  XOR U6358 ( .A(n5399), .B(n5398), .Z(n5400) );
  NANDN U6359 ( .A(rst), .B(n5400), .Z(n5401) );
  NAND U6360 ( .A(n5402), .B(n5401), .Z(n1607) );
  NAND U6361 ( .A(c[71]), .B(rst), .Z(n5407) );
  XNOR U6362 ( .A(n5404), .B(n5403), .Z(n5405) );
  NANDN U6363 ( .A(rst), .B(n5405), .Z(n5406) );
  NAND U6364 ( .A(n5407), .B(n5406), .Z(n1608) );
  NAND U6365 ( .A(c[72]), .B(rst), .Z(n5412) );
  XOR U6366 ( .A(n5409), .B(n5408), .Z(n5410) );
  NANDN U6367 ( .A(rst), .B(n5410), .Z(n5411) );
  NAND U6368 ( .A(n5412), .B(n5411), .Z(n1609) );
  NAND U6369 ( .A(c[73]), .B(rst), .Z(n5417) );
  XNOR U6370 ( .A(n5414), .B(n5413), .Z(n5415) );
  NANDN U6371 ( .A(rst), .B(n5415), .Z(n5416) );
  NAND U6372 ( .A(n5417), .B(n5416), .Z(n1610) );
  NAND U6373 ( .A(c[74]), .B(rst), .Z(n5422) );
  XOR U6374 ( .A(n5419), .B(n5418), .Z(n5420) );
  NANDN U6375 ( .A(rst), .B(n5420), .Z(n5421) );
  NAND U6376 ( .A(n5422), .B(n5421), .Z(n1611) );
  NAND U6377 ( .A(c[75]), .B(rst), .Z(n5427) );
  XNOR U6378 ( .A(n5424), .B(n5423), .Z(n5425) );
  NANDN U6379 ( .A(rst), .B(n5425), .Z(n5426) );
  NAND U6380 ( .A(n5427), .B(n5426), .Z(n1612) );
  NAND U6381 ( .A(c[76]), .B(rst), .Z(n5432) );
  XOR U6382 ( .A(n5429), .B(n5428), .Z(n5430) );
  NANDN U6383 ( .A(rst), .B(n5430), .Z(n5431) );
  NAND U6384 ( .A(n5432), .B(n5431), .Z(n1613) );
  NAND U6385 ( .A(c[77]), .B(rst), .Z(n5437) );
  XNOR U6386 ( .A(n5434), .B(n5433), .Z(n5435) );
  NANDN U6387 ( .A(rst), .B(n5435), .Z(n5436) );
  NAND U6388 ( .A(n5437), .B(n5436), .Z(n1614) );
  NAND U6389 ( .A(c[78]), .B(rst), .Z(n5442) );
  XOR U6390 ( .A(n5439), .B(n5438), .Z(n5440) );
  NANDN U6391 ( .A(rst), .B(n5440), .Z(n5441) );
  NAND U6392 ( .A(n5442), .B(n5441), .Z(n1615) );
  NAND U6393 ( .A(c[79]), .B(rst), .Z(n5447) );
  XNOR U6394 ( .A(n5444), .B(n5443), .Z(n5445) );
  NANDN U6395 ( .A(rst), .B(n5445), .Z(n5446) );
  NAND U6396 ( .A(n5447), .B(n5446), .Z(n1616) );
  NAND U6397 ( .A(c[80]), .B(rst), .Z(n5452) );
  XOR U6398 ( .A(n5449), .B(n5448), .Z(n5450) );
  NANDN U6399 ( .A(rst), .B(n5450), .Z(n5451) );
  NAND U6400 ( .A(n5452), .B(n5451), .Z(n1617) );
  NAND U6401 ( .A(c[81]), .B(rst), .Z(n5457) );
  XNOR U6402 ( .A(n5454), .B(n5453), .Z(n5455) );
  NANDN U6403 ( .A(rst), .B(n5455), .Z(n5456) );
  NAND U6404 ( .A(n5457), .B(n5456), .Z(n1618) );
  NAND U6405 ( .A(c[82]), .B(rst), .Z(n5462) );
  XOR U6406 ( .A(n5459), .B(n5458), .Z(n5460) );
  NANDN U6407 ( .A(rst), .B(n5460), .Z(n5461) );
  NAND U6408 ( .A(n5462), .B(n5461), .Z(n1619) );
  NAND U6409 ( .A(c[83]), .B(rst), .Z(n5467) );
  XNOR U6410 ( .A(n5464), .B(n5463), .Z(n5465) );
  NANDN U6411 ( .A(rst), .B(n5465), .Z(n5466) );
  NAND U6412 ( .A(n5467), .B(n5466), .Z(n1620) );
  NAND U6413 ( .A(c[84]), .B(rst), .Z(n5472) );
  XNOR U6414 ( .A(n5469), .B(n5468), .Z(n5470) );
  NANDN U6415 ( .A(rst), .B(n5470), .Z(n5471) );
  NAND U6416 ( .A(n5472), .B(n5471), .Z(n1621) );
  NAND U6417 ( .A(c[85]), .B(rst), .Z(n5477) );
  XNOR U6418 ( .A(n5474), .B(n5473), .Z(n5475) );
  NANDN U6419 ( .A(rst), .B(n5475), .Z(n5476) );
  NAND U6420 ( .A(n5477), .B(n5476), .Z(n1622) );
  NAND U6421 ( .A(c[86]), .B(rst), .Z(n5482) );
  XNOR U6422 ( .A(n5479), .B(n5478), .Z(n5480) );
  NANDN U6423 ( .A(rst), .B(n5480), .Z(n5481) );
  NAND U6424 ( .A(n5482), .B(n5481), .Z(n1623) );
  NAND U6425 ( .A(c[87]), .B(rst), .Z(n5487) );
  XOR U6426 ( .A(n5484), .B(n5483), .Z(n5485) );
  NANDN U6427 ( .A(rst), .B(n5485), .Z(n5486) );
  NAND U6428 ( .A(n5487), .B(n5486), .Z(n1624) );
  NAND U6429 ( .A(c[88]), .B(rst), .Z(n5492) );
  XNOR U6430 ( .A(n5489), .B(n5488), .Z(n5490) );
  NANDN U6431 ( .A(rst), .B(n5490), .Z(n5491) );
  NAND U6432 ( .A(n5492), .B(n5491), .Z(n1625) );
  NAND U6433 ( .A(c[89]), .B(rst), .Z(n5497) );
  XNOR U6434 ( .A(n5494), .B(n5493), .Z(n5495) );
  NANDN U6435 ( .A(rst), .B(n5495), .Z(n5496) );
  NAND U6436 ( .A(n5497), .B(n5496), .Z(n1626) );
  NAND U6437 ( .A(c[90]), .B(rst), .Z(n5502) );
  XNOR U6438 ( .A(n5499), .B(n5498), .Z(n5500) );
  NANDN U6439 ( .A(rst), .B(n5500), .Z(n5501) );
  NAND U6440 ( .A(n5502), .B(n5501), .Z(n1627) );
  NAND U6441 ( .A(c[91]), .B(rst), .Z(n5507) );
  XNOR U6442 ( .A(n5504), .B(n5503), .Z(n5505) );
  NANDN U6443 ( .A(rst), .B(n5505), .Z(n5506) );
  NAND U6444 ( .A(n5507), .B(n5506), .Z(n1628) );
  NAND U6445 ( .A(c[92]), .B(rst), .Z(n5512) );
  XOR U6446 ( .A(n5509), .B(n5508), .Z(n5510) );
  NANDN U6447 ( .A(rst), .B(n5510), .Z(n5511) );
  NAND U6448 ( .A(n5512), .B(n5511), .Z(n1629) );
  NAND U6449 ( .A(c[93]), .B(rst), .Z(n5517) );
  XNOR U6450 ( .A(n5514), .B(n5513), .Z(n5515) );
  NANDN U6451 ( .A(rst), .B(n5515), .Z(n5516) );
  NAND U6452 ( .A(n5517), .B(n5516), .Z(n1630) );
  NAND U6453 ( .A(c[94]), .B(rst), .Z(n5522) );
  XNOR U6454 ( .A(n5519), .B(n5518), .Z(n5520) );
  NANDN U6455 ( .A(rst), .B(n5520), .Z(n5521) );
  NAND U6456 ( .A(n5522), .B(n5521), .Z(n1631) );
  NAND U6457 ( .A(c[95]), .B(rst), .Z(n5527) );
  XNOR U6458 ( .A(n5524), .B(n5523), .Z(n5525) );
  NANDN U6459 ( .A(rst), .B(n5525), .Z(n5526) );
  NAND U6460 ( .A(n5527), .B(n5526), .Z(n1632) );
  NAND U6461 ( .A(c[96]), .B(rst), .Z(n5532) );
  XNOR U6462 ( .A(n5529), .B(n5528), .Z(n5530) );
  NANDN U6463 ( .A(rst), .B(n5530), .Z(n5531) );
  NAND U6464 ( .A(n5532), .B(n5531), .Z(n1633) );
  NAND U6465 ( .A(c[97]), .B(rst), .Z(n5537) );
  XOR U6466 ( .A(n5534), .B(n5533), .Z(n5535) );
  NANDN U6467 ( .A(rst), .B(n5535), .Z(n5536) );
  NAND U6468 ( .A(n5537), .B(n5536), .Z(n1634) );
  NAND U6469 ( .A(c[98]), .B(rst), .Z(n5542) );
  XNOR U6470 ( .A(n5539), .B(n5538), .Z(n5540) );
  NANDN U6471 ( .A(rst), .B(n5540), .Z(n5541) );
  NAND U6472 ( .A(n5542), .B(n5541), .Z(n1635) );
  NAND U6473 ( .A(c[99]), .B(rst), .Z(n5547) );
  XOR U6474 ( .A(n5544), .B(n5543), .Z(n5545) );
  NANDN U6475 ( .A(rst), .B(n5545), .Z(n5546) );
  NAND U6476 ( .A(n5547), .B(n5546), .Z(n1636) );
  NAND U6477 ( .A(c[100]), .B(rst), .Z(n5552) );
  XNOR U6478 ( .A(n5549), .B(n5548), .Z(n5550) );
  NANDN U6479 ( .A(rst), .B(n5550), .Z(n5551) );
  NAND U6480 ( .A(n5552), .B(n5551), .Z(n1637) );
  NAND U6481 ( .A(c[101]), .B(rst), .Z(n5557) );
  XOR U6482 ( .A(n5554), .B(n5553), .Z(n5555) );
  NANDN U6483 ( .A(rst), .B(n5555), .Z(n5556) );
  NAND U6484 ( .A(n5557), .B(n5556), .Z(n1638) );
  NAND U6485 ( .A(c[102]), .B(rst), .Z(n5562) );
  XNOR U6486 ( .A(n5559), .B(n5558), .Z(n5560) );
  NANDN U6487 ( .A(rst), .B(n5560), .Z(n5561) );
  NAND U6488 ( .A(n5562), .B(n5561), .Z(n1639) );
  NAND U6489 ( .A(c[103]), .B(rst), .Z(n5567) );
  XOR U6490 ( .A(n5564), .B(n5563), .Z(n5565) );
  NANDN U6491 ( .A(rst), .B(n5565), .Z(n5566) );
  NAND U6492 ( .A(n5567), .B(n5566), .Z(n1640) );
  NAND U6493 ( .A(c[104]), .B(rst), .Z(n5572) );
  XNOR U6494 ( .A(n5569), .B(n5568), .Z(n5570) );
  NANDN U6495 ( .A(rst), .B(n5570), .Z(n5571) );
  NAND U6496 ( .A(n5572), .B(n5571), .Z(n1641) );
  NAND U6497 ( .A(c[105]), .B(rst), .Z(n5577) );
  XOR U6498 ( .A(n5574), .B(n5573), .Z(n5575) );
  NANDN U6499 ( .A(rst), .B(n5575), .Z(n5576) );
  NAND U6500 ( .A(n5577), .B(n5576), .Z(n1642) );
  NAND U6501 ( .A(c[106]), .B(rst), .Z(n5582) );
  XNOR U6502 ( .A(n5579), .B(n5578), .Z(n5580) );
  NANDN U6503 ( .A(rst), .B(n5580), .Z(n5581) );
  NAND U6504 ( .A(n5582), .B(n5581), .Z(n1643) );
  NAND U6505 ( .A(c[107]), .B(rst), .Z(n5587) );
  XOR U6506 ( .A(n5584), .B(n5583), .Z(n5585) );
  NANDN U6507 ( .A(rst), .B(n5585), .Z(n5586) );
  NAND U6508 ( .A(n5587), .B(n5586), .Z(n1644) );
  NAND U6509 ( .A(c[108]), .B(rst), .Z(n5592) );
  XNOR U6510 ( .A(n5589), .B(n5588), .Z(n5590) );
  NANDN U6511 ( .A(rst), .B(n5590), .Z(n5591) );
  NAND U6512 ( .A(n5592), .B(n5591), .Z(n1645) );
  NAND U6513 ( .A(c[109]), .B(rst), .Z(n5597) );
  XOR U6514 ( .A(n5594), .B(n5593), .Z(n5595) );
  NANDN U6515 ( .A(rst), .B(n5595), .Z(n5596) );
  NAND U6516 ( .A(n5597), .B(n5596), .Z(n1646) );
  NAND U6517 ( .A(c[110]), .B(rst), .Z(n5602) );
  XNOR U6518 ( .A(n5599), .B(n5598), .Z(n5600) );
  NANDN U6519 ( .A(rst), .B(n5600), .Z(n5601) );
  NAND U6520 ( .A(n5602), .B(n5601), .Z(n1647) );
  NAND U6521 ( .A(c[111]), .B(rst), .Z(n5607) );
  XOR U6522 ( .A(n5604), .B(n5603), .Z(n5605) );
  NANDN U6523 ( .A(rst), .B(n5605), .Z(n5606) );
  NAND U6524 ( .A(n5607), .B(n5606), .Z(n1648) );
  NAND U6525 ( .A(c[112]), .B(rst), .Z(n5612) );
  XNOR U6526 ( .A(n5609), .B(n5608), .Z(n5610) );
  NANDN U6527 ( .A(rst), .B(n5610), .Z(n5611) );
  NAND U6528 ( .A(n5612), .B(n5611), .Z(n1649) );
  NAND U6529 ( .A(c[113]), .B(rst), .Z(n5617) );
  XOR U6530 ( .A(n5614), .B(n5613), .Z(n5615) );
  NANDN U6531 ( .A(rst), .B(n5615), .Z(n5616) );
  NAND U6532 ( .A(n5617), .B(n5616), .Z(n1650) );
  NAND U6533 ( .A(c[114]), .B(rst), .Z(n5622) );
  XNOR U6534 ( .A(n5619), .B(n5618), .Z(n5620) );
  NANDN U6535 ( .A(rst), .B(n5620), .Z(n5621) );
  NAND U6536 ( .A(n5622), .B(n5621), .Z(n1651) );
  NAND U6537 ( .A(c[115]), .B(rst), .Z(n5627) );
  XOR U6538 ( .A(n5624), .B(n5623), .Z(n5625) );
  NANDN U6539 ( .A(rst), .B(n5625), .Z(n5626) );
  NAND U6540 ( .A(n5627), .B(n5626), .Z(n1652) );
  NAND U6541 ( .A(c[116]), .B(rst), .Z(n5632) );
  XNOR U6542 ( .A(n5629), .B(n5628), .Z(n5630) );
  NANDN U6543 ( .A(rst), .B(n5630), .Z(n5631) );
  NAND U6544 ( .A(n5632), .B(n5631), .Z(n1653) );
  NAND U6545 ( .A(c[117]), .B(rst), .Z(n5637) );
  XOR U6546 ( .A(n5634), .B(n5633), .Z(n5635) );
  NANDN U6547 ( .A(rst), .B(n5635), .Z(n5636) );
  NAND U6548 ( .A(n5637), .B(n5636), .Z(n1654) );
  NAND U6549 ( .A(c[118]), .B(rst), .Z(n5642) );
  XNOR U6550 ( .A(n5639), .B(n5638), .Z(n5640) );
  NANDN U6551 ( .A(rst), .B(n5640), .Z(n5641) );
  NAND U6552 ( .A(n5642), .B(n5641), .Z(n1655) );
  NAND U6553 ( .A(c[119]), .B(rst), .Z(n5647) );
  XOR U6554 ( .A(n5644), .B(n5643), .Z(n5645) );
  NANDN U6555 ( .A(rst), .B(n5645), .Z(n5646) );
  NAND U6556 ( .A(n5647), .B(n5646), .Z(n1656) );
  NAND U6557 ( .A(c[120]), .B(rst), .Z(n5652) );
  XNOR U6558 ( .A(n5649), .B(n5648), .Z(n5650) );
  NANDN U6559 ( .A(rst), .B(n5650), .Z(n5651) );
  NAND U6560 ( .A(n5652), .B(n5651), .Z(n1657) );
  NAND U6561 ( .A(c[121]), .B(rst), .Z(n5657) );
  XOR U6562 ( .A(n5654), .B(n5653), .Z(n5655) );
  NANDN U6563 ( .A(rst), .B(n5655), .Z(n5656) );
  NAND U6564 ( .A(n5657), .B(n5656), .Z(n1658) );
  NAND U6565 ( .A(c[122]), .B(rst), .Z(n5662) );
  XNOR U6566 ( .A(n5659), .B(n5658), .Z(n5660) );
  NANDN U6567 ( .A(rst), .B(n5660), .Z(n5661) );
  NAND U6568 ( .A(n5662), .B(n5661), .Z(n1659) );
  NAND U6569 ( .A(c[123]), .B(rst), .Z(n5667) );
  XOR U6570 ( .A(n5664), .B(n5663), .Z(n5665) );
  NANDN U6571 ( .A(rst), .B(n5665), .Z(n5666) );
  NAND U6572 ( .A(n5667), .B(n5666), .Z(n1660) );
  NAND U6573 ( .A(c[124]), .B(rst), .Z(n5672) );
  XNOR U6574 ( .A(n5669), .B(n5668), .Z(n5670) );
  NANDN U6575 ( .A(rst), .B(n5670), .Z(n5671) );
  NAND U6576 ( .A(n5672), .B(n5671), .Z(n1661) );
  NAND U6577 ( .A(c[125]), .B(rst), .Z(n5677) );
  XNOR U6578 ( .A(n5674), .B(n5673), .Z(n5675) );
  NANDN U6579 ( .A(rst), .B(n5675), .Z(n5676) );
  NAND U6580 ( .A(n5677), .B(n5676), .Z(n1662) );
  NAND U6581 ( .A(c[126]), .B(rst), .Z(n5682) );
  XNOR U6582 ( .A(n5679), .B(n5678), .Z(n5680) );
  NANDN U6583 ( .A(rst), .B(n5680), .Z(n5681) );
  NAND U6584 ( .A(n5682), .B(n5681), .Z(n1663) );
  NAND U6585 ( .A(c[127]), .B(rst), .Z(n5687) );
  XNOR U6586 ( .A(n5684), .B(n5683), .Z(n5685) );
  NANDN U6587 ( .A(rst), .B(n5685), .Z(n5686) );
  NAND U6588 ( .A(n5687), .B(n5686), .Z(n1664) );
  NAND U6589 ( .A(c[128]), .B(rst), .Z(n5692) );
  XOR U6590 ( .A(n5689), .B(n5688), .Z(n5690) );
  NANDN U6591 ( .A(rst), .B(n5690), .Z(n5691) );
  NAND U6592 ( .A(n5692), .B(n5691), .Z(n1665) );
  NAND U6593 ( .A(c[129]), .B(rst), .Z(n5697) );
  XNOR U6594 ( .A(n5694), .B(n5693), .Z(n5695) );
  NANDN U6595 ( .A(rst), .B(n5695), .Z(n5696) );
  NAND U6596 ( .A(n5697), .B(n5696), .Z(n1666) );
  NAND U6597 ( .A(c[130]), .B(rst), .Z(n5702) );
  XOR U6598 ( .A(n5699), .B(n5698), .Z(n5700) );
  NANDN U6599 ( .A(rst), .B(n5700), .Z(n5701) );
  NAND U6600 ( .A(n5702), .B(n5701), .Z(n1667) );
  NAND U6601 ( .A(c[131]), .B(rst), .Z(n5707) );
  XNOR U6602 ( .A(n5704), .B(n5703), .Z(n5705) );
  NANDN U6603 ( .A(rst), .B(n5705), .Z(n5706) );
  NAND U6604 ( .A(n5707), .B(n5706), .Z(n1668) );
  NAND U6605 ( .A(c[132]), .B(rst), .Z(n5712) );
  XOR U6606 ( .A(n5709), .B(n5708), .Z(n5710) );
  NANDN U6607 ( .A(rst), .B(n5710), .Z(n5711) );
  NAND U6608 ( .A(n5712), .B(n5711), .Z(n1669) );
  NAND U6609 ( .A(c[133]), .B(rst), .Z(n5717) );
  XNOR U6610 ( .A(n5714), .B(n5713), .Z(n5715) );
  NANDN U6611 ( .A(rst), .B(n5715), .Z(n5716) );
  NAND U6612 ( .A(n5717), .B(n5716), .Z(n1670) );
  NAND U6613 ( .A(c[134]), .B(rst), .Z(n5722) );
  XOR U6614 ( .A(n5719), .B(n5718), .Z(n5720) );
  NANDN U6615 ( .A(rst), .B(n5720), .Z(n5721) );
  NAND U6616 ( .A(n5722), .B(n5721), .Z(n1671) );
  NAND U6617 ( .A(c[135]), .B(rst), .Z(n5727) );
  XNOR U6618 ( .A(n5724), .B(n5723), .Z(n5725) );
  NANDN U6619 ( .A(rst), .B(n5725), .Z(n5726) );
  NAND U6620 ( .A(n5727), .B(n5726), .Z(n1672) );
  NAND U6621 ( .A(c[136]), .B(rst), .Z(n5732) );
  XOR U6622 ( .A(n5729), .B(n5728), .Z(n5730) );
  NANDN U6623 ( .A(rst), .B(n5730), .Z(n5731) );
  NAND U6624 ( .A(n5732), .B(n5731), .Z(n1673) );
  NAND U6625 ( .A(c[137]), .B(rst), .Z(n5737) );
  XNOR U6626 ( .A(n5734), .B(n5733), .Z(n5735) );
  NANDN U6627 ( .A(rst), .B(n5735), .Z(n5736) );
  NAND U6628 ( .A(n5737), .B(n5736), .Z(n1674) );
  NAND U6629 ( .A(c[138]), .B(rst), .Z(n5742) );
  XOR U6630 ( .A(n5739), .B(n5738), .Z(n5740) );
  NANDN U6631 ( .A(rst), .B(n5740), .Z(n5741) );
  NAND U6632 ( .A(n5742), .B(n5741), .Z(n1675) );
  NAND U6633 ( .A(c[139]), .B(rst), .Z(n5747) );
  XNOR U6634 ( .A(n5744), .B(n5743), .Z(n5745) );
  NANDN U6635 ( .A(rst), .B(n5745), .Z(n5746) );
  NAND U6636 ( .A(n5747), .B(n5746), .Z(n1676) );
  NAND U6637 ( .A(c[140]), .B(rst), .Z(n5752) );
  XOR U6638 ( .A(n5749), .B(n5748), .Z(n5750) );
  NANDN U6639 ( .A(rst), .B(n5750), .Z(n5751) );
  NAND U6640 ( .A(n5752), .B(n5751), .Z(n1677) );
  NAND U6641 ( .A(c[141]), .B(rst), .Z(n5757) );
  XNOR U6642 ( .A(n5754), .B(n5753), .Z(n5755) );
  NANDN U6643 ( .A(rst), .B(n5755), .Z(n5756) );
  NAND U6644 ( .A(n5757), .B(n5756), .Z(n1678) );
  NAND U6645 ( .A(c[142]), .B(rst), .Z(n5762) );
  XOR U6646 ( .A(n5759), .B(n5758), .Z(n5760) );
  NANDN U6647 ( .A(rst), .B(n5760), .Z(n5761) );
  NAND U6648 ( .A(n5762), .B(n5761), .Z(n1679) );
  NAND U6649 ( .A(c[143]), .B(rst), .Z(n5767) );
  XNOR U6650 ( .A(n5764), .B(n5763), .Z(n5765) );
  NANDN U6651 ( .A(rst), .B(n5765), .Z(n5766) );
  NAND U6652 ( .A(n5767), .B(n5766), .Z(n1680) );
  NAND U6653 ( .A(c[144]), .B(rst), .Z(n5772) );
  XOR U6654 ( .A(n5769), .B(n5768), .Z(n5770) );
  NANDN U6655 ( .A(rst), .B(n5770), .Z(n5771) );
  NAND U6656 ( .A(n5772), .B(n5771), .Z(n1681) );
  NAND U6657 ( .A(c[145]), .B(rst), .Z(n5777) );
  XNOR U6658 ( .A(n5774), .B(n5773), .Z(n5775) );
  NANDN U6659 ( .A(rst), .B(n5775), .Z(n5776) );
  NAND U6660 ( .A(n5777), .B(n5776), .Z(n1682) );
  NAND U6661 ( .A(c[146]), .B(rst), .Z(n5782) );
  XOR U6662 ( .A(n5779), .B(n5778), .Z(n5780) );
  NANDN U6663 ( .A(rst), .B(n5780), .Z(n5781) );
  NAND U6664 ( .A(n5782), .B(n5781), .Z(n1683) );
  NAND U6665 ( .A(c[147]), .B(rst), .Z(n5787) );
  XNOR U6666 ( .A(n5784), .B(n5783), .Z(n5785) );
  NANDN U6667 ( .A(rst), .B(n5785), .Z(n5786) );
  NAND U6668 ( .A(n5787), .B(n5786), .Z(n1684) );
  NAND U6669 ( .A(c[148]), .B(rst), .Z(n5792) );
  XOR U6670 ( .A(n5789), .B(n5788), .Z(n5790) );
  NANDN U6671 ( .A(rst), .B(n5790), .Z(n5791) );
  NAND U6672 ( .A(n5792), .B(n5791), .Z(n1685) );
  NAND U6673 ( .A(c[149]), .B(rst), .Z(n5797) );
  XNOR U6674 ( .A(n5794), .B(n5793), .Z(n5795) );
  NANDN U6675 ( .A(rst), .B(n5795), .Z(n5796) );
  NAND U6676 ( .A(n5797), .B(n5796), .Z(n1686) );
  NAND U6677 ( .A(c[150]), .B(rst), .Z(n5802) );
  XOR U6678 ( .A(n5799), .B(n5798), .Z(n5800) );
  NANDN U6679 ( .A(rst), .B(n5800), .Z(n5801) );
  NAND U6680 ( .A(n5802), .B(n5801), .Z(n1687) );
  NAND U6681 ( .A(c[151]), .B(rst), .Z(n5807) );
  XNOR U6682 ( .A(n5804), .B(n5803), .Z(n5805) );
  NANDN U6683 ( .A(rst), .B(n5805), .Z(n5806) );
  NAND U6684 ( .A(n5807), .B(n5806), .Z(n1688) );
  NAND U6685 ( .A(c[152]), .B(rst), .Z(n5812) );
  XNOR U6686 ( .A(n5809), .B(n5808), .Z(n5810) );
  NANDN U6687 ( .A(rst), .B(n5810), .Z(n5811) );
  NAND U6688 ( .A(n5812), .B(n5811), .Z(n1689) );
  NAND U6689 ( .A(c[153]), .B(rst), .Z(n5817) );
  XNOR U6690 ( .A(n5814), .B(n5813), .Z(n5815) );
  NANDN U6691 ( .A(rst), .B(n5815), .Z(n5816) );
  NAND U6692 ( .A(n5817), .B(n5816), .Z(n1690) );
  NAND U6693 ( .A(c[154]), .B(rst), .Z(n5822) );
  XNOR U6694 ( .A(n5819), .B(n5818), .Z(n5820) );
  NANDN U6695 ( .A(rst), .B(n5820), .Z(n5821) );
  NAND U6696 ( .A(n5822), .B(n5821), .Z(n1691) );
  NAND U6697 ( .A(c[155]), .B(rst), .Z(n5827) );
  XOR U6698 ( .A(n5824), .B(n5823), .Z(n5825) );
  NANDN U6699 ( .A(rst), .B(n5825), .Z(n5826) );
  NAND U6700 ( .A(n5827), .B(n5826), .Z(n1692) );
  NAND U6701 ( .A(c[156]), .B(rst), .Z(n5832) );
  XNOR U6702 ( .A(n5829), .B(n5828), .Z(n5830) );
  NANDN U6703 ( .A(rst), .B(n5830), .Z(n5831) );
  NAND U6704 ( .A(n5832), .B(n5831), .Z(n1693) );
  NAND U6705 ( .A(c[157]), .B(rst), .Z(n5837) );
  XNOR U6706 ( .A(n5834), .B(n5833), .Z(n5835) );
  NANDN U6707 ( .A(rst), .B(n5835), .Z(n5836) );
  NAND U6708 ( .A(n5837), .B(n5836), .Z(n1694) );
  NAND U6709 ( .A(c[158]), .B(rst), .Z(n5842) );
  XNOR U6710 ( .A(n5839), .B(n5838), .Z(n5840) );
  NANDN U6711 ( .A(rst), .B(n5840), .Z(n5841) );
  NAND U6712 ( .A(n5842), .B(n5841), .Z(n1695) );
  NAND U6713 ( .A(c[159]), .B(rst), .Z(n5847) );
  XNOR U6714 ( .A(n5844), .B(n5843), .Z(n5845) );
  NANDN U6715 ( .A(rst), .B(n5845), .Z(n5846) );
  NAND U6716 ( .A(n5847), .B(n5846), .Z(n1696) );
  NAND U6717 ( .A(c[160]), .B(rst), .Z(n5852) );
  XOR U6718 ( .A(n5849), .B(n5848), .Z(n5850) );
  NANDN U6719 ( .A(rst), .B(n5850), .Z(n5851) );
  NAND U6720 ( .A(n5852), .B(n5851), .Z(n1697) );
  NAND U6721 ( .A(c[161]), .B(rst), .Z(n5857) );
  XNOR U6722 ( .A(n5854), .B(n5853), .Z(n5855) );
  NANDN U6723 ( .A(rst), .B(n5855), .Z(n5856) );
  NAND U6724 ( .A(n5857), .B(n5856), .Z(n1698) );
  NAND U6725 ( .A(c[162]), .B(rst), .Z(n5862) );
  XOR U6726 ( .A(n5859), .B(n5858), .Z(n5860) );
  NANDN U6727 ( .A(rst), .B(n5860), .Z(n5861) );
  NAND U6728 ( .A(n5862), .B(n5861), .Z(n1699) );
  NAND U6729 ( .A(c[163]), .B(rst), .Z(n5867) );
  XNOR U6730 ( .A(n5864), .B(n5863), .Z(n5865) );
  NANDN U6731 ( .A(rst), .B(n5865), .Z(n5866) );
  NAND U6732 ( .A(n5867), .B(n5866), .Z(n1700) );
  NAND U6733 ( .A(c[164]), .B(rst), .Z(n5872) );
  XOR U6734 ( .A(n5869), .B(n5868), .Z(n5870) );
  NANDN U6735 ( .A(rst), .B(n5870), .Z(n5871) );
  NAND U6736 ( .A(n5872), .B(n5871), .Z(n1701) );
  NAND U6737 ( .A(c[165]), .B(rst), .Z(n5877) );
  XNOR U6738 ( .A(n5874), .B(n5873), .Z(n5875) );
  NANDN U6739 ( .A(rst), .B(n5875), .Z(n5876) );
  NAND U6740 ( .A(n5877), .B(n5876), .Z(n1702) );
  NAND U6741 ( .A(c[166]), .B(rst), .Z(n5882) );
  XNOR U6742 ( .A(n5879), .B(n5878), .Z(n5880) );
  NANDN U6743 ( .A(rst), .B(n5880), .Z(n5881) );
  NAND U6744 ( .A(n5882), .B(n5881), .Z(n1703) );
  NAND U6745 ( .A(c[167]), .B(rst), .Z(n5887) );
  XNOR U6746 ( .A(n5884), .B(n5883), .Z(n5885) );
  NANDN U6747 ( .A(rst), .B(n5885), .Z(n5886) );
  NAND U6748 ( .A(n5887), .B(n5886), .Z(n1704) );
  NAND U6749 ( .A(c[168]), .B(rst), .Z(n5892) );
  XNOR U6750 ( .A(n5889), .B(n5888), .Z(n5890) );
  NANDN U6751 ( .A(rst), .B(n5890), .Z(n5891) );
  NAND U6752 ( .A(n5892), .B(n5891), .Z(n1705) );
  NAND U6753 ( .A(c[169]), .B(rst), .Z(n5897) );
  XOR U6754 ( .A(n5894), .B(n5893), .Z(n5895) );
  NANDN U6755 ( .A(rst), .B(n5895), .Z(n5896) );
  NAND U6756 ( .A(n5897), .B(n5896), .Z(n1706) );
  NAND U6757 ( .A(c[170]), .B(rst), .Z(n5902) );
  XNOR U6758 ( .A(n5899), .B(n5898), .Z(n5900) );
  NANDN U6759 ( .A(rst), .B(n5900), .Z(n5901) );
  NAND U6760 ( .A(n5902), .B(n5901), .Z(n1707) );
  NAND U6761 ( .A(c[171]), .B(rst), .Z(n5907) );
  XOR U6762 ( .A(n5904), .B(n5903), .Z(n5905) );
  NANDN U6763 ( .A(rst), .B(n5905), .Z(n5906) );
  NAND U6764 ( .A(n5907), .B(n5906), .Z(n1708) );
  NAND U6765 ( .A(c[172]), .B(rst), .Z(n5912) );
  XNOR U6766 ( .A(n5909), .B(n5908), .Z(n5910) );
  NANDN U6767 ( .A(rst), .B(n5910), .Z(n5911) );
  NAND U6768 ( .A(n5912), .B(n5911), .Z(n1709) );
  NAND U6769 ( .A(c[173]), .B(rst), .Z(n5917) );
  XOR U6770 ( .A(n5914), .B(n5913), .Z(n5915) );
  NANDN U6771 ( .A(rst), .B(n5915), .Z(n5916) );
  NAND U6772 ( .A(n5917), .B(n5916), .Z(n1710) );
  NAND U6773 ( .A(c[174]), .B(rst), .Z(n5922) );
  XNOR U6774 ( .A(n5919), .B(n5918), .Z(n5920) );
  NANDN U6775 ( .A(rst), .B(n5920), .Z(n5921) );
  NAND U6776 ( .A(n5922), .B(n5921), .Z(n1711) );
  NAND U6777 ( .A(c[175]), .B(rst), .Z(n5927) );
  XOR U6778 ( .A(n5924), .B(n5923), .Z(n5925) );
  NANDN U6779 ( .A(rst), .B(n5925), .Z(n5926) );
  NAND U6780 ( .A(n5927), .B(n5926), .Z(n1712) );
  NAND U6781 ( .A(c[176]), .B(rst), .Z(n5932) );
  XNOR U6782 ( .A(n5929), .B(n5928), .Z(n5930) );
  NANDN U6783 ( .A(rst), .B(n5930), .Z(n5931) );
  NAND U6784 ( .A(n5932), .B(n5931), .Z(n1713) );
  NAND U6785 ( .A(c[177]), .B(rst), .Z(n5937) );
  XOR U6786 ( .A(n5934), .B(n5933), .Z(n5935) );
  NANDN U6787 ( .A(rst), .B(n5935), .Z(n5936) );
  NAND U6788 ( .A(n5937), .B(n5936), .Z(n1714) );
  NAND U6789 ( .A(c[178]), .B(rst), .Z(n5942) );
  XNOR U6790 ( .A(n5939), .B(n5938), .Z(n5940) );
  NANDN U6791 ( .A(rst), .B(n5940), .Z(n5941) );
  NAND U6792 ( .A(n5942), .B(n5941), .Z(n1715) );
  NAND U6793 ( .A(c[179]), .B(rst), .Z(n5947) );
  XOR U6794 ( .A(n5944), .B(n5943), .Z(n5945) );
  NANDN U6795 ( .A(rst), .B(n5945), .Z(n5946) );
  NAND U6796 ( .A(n5947), .B(n5946), .Z(n1716) );
  NAND U6797 ( .A(c[180]), .B(rst), .Z(n5952) );
  XNOR U6798 ( .A(n5949), .B(n5948), .Z(n5950) );
  NANDN U6799 ( .A(rst), .B(n5950), .Z(n5951) );
  NAND U6800 ( .A(n5952), .B(n5951), .Z(n1717) );
  NAND U6801 ( .A(c[181]), .B(rst), .Z(n5957) );
  XOR U6802 ( .A(n5954), .B(n5953), .Z(n5955) );
  NANDN U6803 ( .A(rst), .B(n5955), .Z(n5956) );
  NAND U6804 ( .A(n5957), .B(n5956), .Z(n1718) );
  NAND U6805 ( .A(c[182]), .B(rst), .Z(n5962) );
  XNOR U6806 ( .A(n5959), .B(n5958), .Z(n5960) );
  NANDN U6807 ( .A(rst), .B(n5960), .Z(n5961) );
  NAND U6808 ( .A(n5962), .B(n5961), .Z(n1719) );
  NAND U6809 ( .A(c[183]), .B(rst), .Z(n5967) );
  XOR U6810 ( .A(n5964), .B(n5963), .Z(n5965) );
  NANDN U6811 ( .A(rst), .B(n5965), .Z(n5966) );
  NAND U6812 ( .A(n5967), .B(n5966), .Z(n1720) );
  NAND U6813 ( .A(c[184]), .B(rst), .Z(n5972) );
  XNOR U6814 ( .A(n5969), .B(n5968), .Z(n5970) );
  NANDN U6815 ( .A(rst), .B(n5970), .Z(n5971) );
  NAND U6816 ( .A(n5972), .B(n5971), .Z(n1721) );
  NAND U6817 ( .A(c[185]), .B(rst), .Z(n5977) );
  XNOR U6818 ( .A(n5974), .B(n5973), .Z(n5975) );
  NANDN U6819 ( .A(rst), .B(n5975), .Z(n5976) );
  NAND U6820 ( .A(n5977), .B(n5976), .Z(n1722) );
  NAND U6821 ( .A(c[186]), .B(rst), .Z(n5982) );
  XNOR U6822 ( .A(n5979), .B(n5978), .Z(n5980) );
  NANDN U6823 ( .A(rst), .B(n5980), .Z(n5981) );
  NAND U6824 ( .A(n5982), .B(n5981), .Z(n1723) );
  NAND U6825 ( .A(c[187]), .B(rst), .Z(n5987) );
  XNOR U6826 ( .A(n5984), .B(n5983), .Z(n5985) );
  NANDN U6827 ( .A(rst), .B(n5985), .Z(n5986) );
  NAND U6828 ( .A(n5987), .B(n5986), .Z(n1724) );
  NAND U6829 ( .A(c[188]), .B(rst), .Z(n5992) );
  XOR U6830 ( .A(n5989), .B(n5988), .Z(n5990) );
  NANDN U6831 ( .A(rst), .B(n5990), .Z(n5991) );
  NAND U6832 ( .A(n5992), .B(n5991), .Z(n1725) );
  NAND U6833 ( .A(c[189]), .B(rst), .Z(n5997) );
  XNOR U6834 ( .A(n5994), .B(n5993), .Z(n5995) );
  NANDN U6835 ( .A(rst), .B(n5995), .Z(n5996) );
  NAND U6836 ( .A(n5997), .B(n5996), .Z(n1726) );
  NAND U6837 ( .A(c[190]), .B(rst), .Z(n6002) );
  XNOR U6838 ( .A(n5999), .B(n5998), .Z(n6000) );
  NANDN U6839 ( .A(rst), .B(n6000), .Z(n6001) );
  NAND U6840 ( .A(n6002), .B(n6001), .Z(n1727) );
  NAND U6841 ( .A(c[191]), .B(rst), .Z(n6007) );
  XNOR U6842 ( .A(n6004), .B(n6003), .Z(n6005) );
  NANDN U6843 ( .A(rst), .B(n6005), .Z(n6006) );
  NAND U6844 ( .A(n6007), .B(n6006), .Z(n1728) );
  NAND U6845 ( .A(c[192]), .B(rst), .Z(n6012) );
  XNOR U6846 ( .A(n6009), .B(n6008), .Z(n6010) );
  NANDN U6847 ( .A(rst), .B(n6010), .Z(n6011) );
  NAND U6848 ( .A(n6012), .B(n6011), .Z(n1729) );
  NAND U6849 ( .A(c[193]), .B(rst), .Z(n6017) );
  XOR U6850 ( .A(n6014), .B(n6013), .Z(n6015) );
  NANDN U6851 ( .A(rst), .B(n6015), .Z(n6016) );
  NAND U6852 ( .A(n6017), .B(n6016), .Z(n1730) );
  NAND U6853 ( .A(c[194]), .B(rst), .Z(n6022) );
  XNOR U6854 ( .A(n6019), .B(n6018), .Z(n6020) );
  NANDN U6855 ( .A(rst), .B(n6020), .Z(n6021) );
  NAND U6856 ( .A(n6022), .B(n6021), .Z(n1731) );
  NAND U6857 ( .A(c[195]), .B(rst), .Z(n6027) );
  XOR U6858 ( .A(n6024), .B(n6023), .Z(n6025) );
  NANDN U6859 ( .A(rst), .B(n6025), .Z(n6026) );
  NAND U6860 ( .A(n6027), .B(n6026), .Z(n1732) );
  NAND U6861 ( .A(c[196]), .B(rst), .Z(n6032) );
  XNOR U6862 ( .A(n6029), .B(n6028), .Z(n6030) );
  NANDN U6863 ( .A(rst), .B(n6030), .Z(n6031) );
  NAND U6864 ( .A(n6032), .B(n6031), .Z(n1733) );
  NAND U6865 ( .A(c[197]), .B(rst), .Z(n6037) );
  XOR U6866 ( .A(n6034), .B(n6033), .Z(n6035) );
  NANDN U6867 ( .A(rst), .B(n6035), .Z(n6036) );
  NAND U6868 ( .A(n6037), .B(n6036), .Z(n1734) );
  NAND U6869 ( .A(c[198]), .B(rst), .Z(n6042) );
  XNOR U6870 ( .A(n6039), .B(n6038), .Z(n6040) );
  NANDN U6871 ( .A(rst), .B(n6040), .Z(n6041) );
  NAND U6872 ( .A(n6042), .B(n6041), .Z(n1735) );
  NAND U6873 ( .A(c[199]), .B(rst), .Z(n6047) );
  XOR U6874 ( .A(n6044), .B(n6043), .Z(n6045) );
  NANDN U6875 ( .A(rst), .B(n6045), .Z(n6046) );
  NAND U6876 ( .A(n6047), .B(n6046), .Z(n1736) );
  NAND U6877 ( .A(c[200]), .B(rst), .Z(n6052) );
  XNOR U6878 ( .A(n6049), .B(n6048), .Z(n6050) );
  NANDN U6879 ( .A(rst), .B(n6050), .Z(n6051) );
  NAND U6880 ( .A(n6052), .B(n6051), .Z(n1737) );
  NAND U6881 ( .A(c[201]), .B(rst), .Z(n6057) );
  XNOR U6882 ( .A(n6054), .B(n6053), .Z(n6055) );
  NANDN U6883 ( .A(rst), .B(n6055), .Z(n6056) );
  NAND U6884 ( .A(n6057), .B(n6056), .Z(n1738) );
  NAND U6885 ( .A(c[202]), .B(rst), .Z(n6062) );
  XNOR U6886 ( .A(n6059), .B(n6058), .Z(n6060) );
  NANDN U6887 ( .A(rst), .B(n6060), .Z(n6061) );
  NAND U6888 ( .A(n6062), .B(n6061), .Z(n1739) );
  NAND U6889 ( .A(c[203]), .B(rst), .Z(n6067) );
  XNOR U6890 ( .A(n6064), .B(n6063), .Z(n6065) );
  NANDN U6891 ( .A(rst), .B(n6065), .Z(n6066) );
  NAND U6892 ( .A(n6067), .B(n6066), .Z(n1740) );
  NAND U6893 ( .A(c[204]), .B(rst), .Z(n6072) );
  XOR U6894 ( .A(n6069), .B(n6068), .Z(n6070) );
  NANDN U6895 ( .A(rst), .B(n6070), .Z(n6071) );
  NAND U6896 ( .A(n6072), .B(n6071), .Z(n1741) );
  NAND U6897 ( .A(c[205]), .B(rst), .Z(n6077) );
  XNOR U6898 ( .A(n6074), .B(n6073), .Z(n6075) );
  NANDN U6899 ( .A(rst), .B(n6075), .Z(n6076) );
  NAND U6900 ( .A(n6077), .B(n6076), .Z(n1742) );
  NAND U6901 ( .A(c[206]), .B(rst), .Z(n6082) );
  XOR U6902 ( .A(n6079), .B(n6078), .Z(n6080) );
  NANDN U6903 ( .A(rst), .B(n6080), .Z(n6081) );
  NAND U6904 ( .A(n6082), .B(n6081), .Z(n1743) );
  NAND U6905 ( .A(c[207]), .B(rst), .Z(n6087) );
  XNOR U6906 ( .A(n6084), .B(n6083), .Z(n6085) );
  NANDN U6907 ( .A(rst), .B(n6085), .Z(n6086) );
  NAND U6908 ( .A(n6087), .B(n6086), .Z(n1744) );
  NAND U6909 ( .A(c[208]), .B(rst), .Z(n6092) );
  XOR U6910 ( .A(n6089), .B(n6088), .Z(n6090) );
  NANDN U6911 ( .A(rst), .B(n6090), .Z(n6091) );
  NAND U6912 ( .A(n6092), .B(n6091), .Z(n1745) );
  NAND U6913 ( .A(c[209]), .B(rst), .Z(n6097) );
  XNOR U6914 ( .A(n6094), .B(n6093), .Z(n6095) );
  NANDN U6915 ( .A(rst), .B(n6095), .Z(n6096) );
  NAND U6916 ( .A(n6097), .B(n6096), .Z(n1746) );
  NAND U6917 ( .A(c[210]), .B(rst), .Z(n6102) );
  XOR U6918 ( .A(n6099), .B(n6098), .Z(n6100) );
  NANDN U6919 ( .A(rst), .B(n6100), .Z(n6101) );
  NAND U6920 ( .A(n6102), .B(n6101), .Z(n1747) );
  NAND U6921 ( .A(c[211]), .B(rst), .Z(n6107) );
  XNOR U6922 ( .A(n6104), .B(n6103), .Z(n6105) );
  NANDN U6923 ( .A(rst), .B(n6105), .Z(n6106) );
  NAND U6924 ( .A(n6107), .B(n6106), .Z(n1748) );
  NAND U6925 ( .A(c[212]), .B(rst), .Z(n6112) );
  XOR U6926 ( .A(n6109), .B(n6108), .Z(n6110) );
  NANDN U6927 ( .A(rst), .B(n6110), .Z(n6111) );
  NAND U6928 ( .A(n6112), .B(n6111), .Z(n1749) );
  NAND U6929 ( .A(c[213]), .B(rst), .Z(n6117) );
  XNOR U6930 ( .A(n6114), .B(n6113), .Z(n6115) );
  NANDN U6931 ( .A(rst), .B(n6115), .Z(n6116) );
  NAND U6932 ( .A(n6117), .B(n6116), .Z(n1750) );
  NAND U6933 ( .A(c[214]), .B(rst), .Z(n6122) );
  XOR U6934 ( .A(n6119), .B(n6118), .Z(n6120) );
  NANDN U6935 ( .A(rst), .B(n6120), .Z(n6121) );
  NAND U6936 ( .A(n6122), .B(n6121), .Z(n1751) );
  NAND U6937 ( .A(c[215]), .B(rst), .Z(n6127) );
  XNOR U6938 ( .A(n6124), .B(n6123), .Z(n6125) );
  NANDN U6939 ( .A(rst), .B(n6125), .Z(n6126) );
  NAND U6940 ( .A(n6127), .B(n6126), .Z(n1752) );
  NAND U6941 ( .A(c[216]), .B(rst), .Z(n6132) );
  XOR U6942 ( .A(n6129), .B(n6128), .Z(n6130) );
  NANDN U6943 ( .A(rst), .B(n6130), .Z(n6131) );
  NAND U6944 ( .A(n6132), .B(n6131), .Z(n1753) );
  NAND U6945 ( .A(c[217]), .B(rst), .Z(n6137) );
  XNOR U6946 ( .A(n6134), .B(n6133), .Z(n6135) );
  NANDN U6947 ( .A(rst), .B(n6135), .Z(n6136) );
  NAND U6948 ( .A(n6137), .B(n6136), .Z(n1754) );
  NAND U6949 ( .A(c[218]), .B(rst), .Z(n6142) );
  XNOR U6950 ( .A(n6139), .B(n6138), .Z(n6140) );
  NANDN U6951 ( .A(rst), .B(n6140), .Z(n6141) );
  NAND U6952 ( .A(n6142), .B(n6141), .Z(n1755) );
  NAND U6953 ( .A(c[219]), .B(rst), .Z(n6147) );
  XNOR U6954 ( .A(n6144), .B(n6143), .Z(n6145) );
  NANDN U6955 ( .A(rst), .B(n6145), .Z(n6146) );
  NAND U6956 ( .A(n6147), .B(n6146), .Z(n1756) );
  NAND U6957 ( .A(c[220]), .B(rst), .Z(n6152) );
  XNOR U6958 ( .A(n6149), .B(n6148), .Z(n6150) );
  NANDN U6959 ( .A(rst), .B(n6150), .Z(n6151) );
  NAND U6960 ( .A(n6152), .B(n6151), .Z(n1757) );
  NAND U6961 ( .A(c[221]), .B(rst), .Z(n6157) );
  XOR U6962 ( .A(n6154), .B(n6153), .Z(n6155) );
  NANDN U6963 ( .A(rst), .B(n6155), .Z(n6156) );
  NAND U6964 ( .A(n6157), .B(n6156), .Z(n1758) );
  NAND U6965 ( .A(c[222]), .B(rst), .Z(n6162) );
  XNOR U6966 ( .A(n6159), .B(n6158), .Z(n6160) );
  NANDN U6967 ( .A(rst), .B(n6160), .Z(n6161) );
  NAND U6968 ( .A(n6162), .B(n6161), .Z(n1759) );
  NAND U6969 ( .A(c[223]), .B(rst), .Z(n6167) );
  XOR U6970 ( .A(n6164), .B(n6163), .Z(n6165) );
  NANDN U6971 ( .A(rst), .B(n6165), .Z(n6166) );
  NAND U6972 ( .A(n6167), .B(n6166), .Z(n1760) );
  NAND U6973 ( .A(c[224]), .B(rst), .Z(n6172) );
  XNOR U6974 ( .A(n6169), .B(n6168), .Z(n6170) );
  NANDN U6975 ( .A(rst), .B(n6170), .Z(n6171) );
  NAND U6976 ( .A(n6172), .B(n6171), .Z(n1761) );
  NAND U6977 ( .A(c[225]), .B(rst), .Z(n6177) );
  XOR U6978 ( .A(n6174), .B(n6173), .Z(n6175) );
  NANDN U6979 ( .A(rst), .B(n6175), .Z(n6176) );
  NAND U6980 ( .A(n6177), .B(n6176), .Z(n1762) );
  NAND U6981 ( .A(c[226]), .B(rst), .Z(n6182) );
  XNOR U6982 ( .A(n6179), .B(n6178), .Z(n6180) );
  NANDN U6983 ( .A(rst), .B(n6180), .Z(n6181) );
  NAND U6984 ( .A(n6182), .B(n6181), .Z(n1763) );
  NAND U6985 ( .A(c[227]), .B(rst), .Z(n6187) );
  XOR U6986 ( .A(n6184), .B(n6183), .Z(n6185) );
  NANDN U6987 ( .A(rst), .B(n6185), .Z(n6186) );
  NAND U6988 ( .A(n6187), .B(n6186), .Z(n1764) );
  NAND U6989 ( .A(c[228]), .B(rst), .Z(n6192) );
  XNOR U6990 ( .A(n6189), .B(n6188), .Z(n6190) );
  NANDN U6991 ( .A(rst), .B(n6190), .Z(n6191) );
  NAND U6992 ( .A(n6192), .B(n6191), .Z(n1765) );
  NAND U6993 ( .A(c[229]), .B(rst), .Z(n6197) );
  XOR U6994 ( .A(n6194), .B(n6193), .Z(n6195) );
  NANDN U6995 ( .A(rst), .B(n6195), .Z(n6196) );
  NAND U6996 ( .A(n6197), .B(n6196), .Z(n1766) );
  NAND U6997 ( .A(c[230]), .B(rst), .Z(n6202) );
  XNOR U6998 ( .A(n6199), .B(n6198), .Z(n6200) );
  NANDN U6999 ( .A(rst), .B(n6200), .Z(n6201) );
  NAND U7000 ( .A(n6202), .B(n6201), .Z(n1767) );
  NAND U7001 ( .A(c[231]), .B(rst), .Z(n6207) );
  XOR U7002 ( .A(n6204), .B(n6203), .Z(n6205) );
  NANDN U7003 ( .A(rst), .B(n6205), .Z(n6206) );
  NAND U7004 ( .A(n6207), .B(n6206), .Z(n1768) );
  NAND U7005 ( .A(c[232]), .B(rst), .Z(n6212) );
  XNOR U7006 ( .A(n6209), .B(n6208), .Z(n6210) );
  NANDN U7007 ( .A(rst), .B(n6210), .Z(n6211) );
  NAND U7008 ( .A(n6212), .B(n6211), .Z(n1769) );
  NAND U7009 ( .A(c[233]), .B(rst), .Z(n6217) );
  XOR U7010 ( .A(n6214), .B(n6213), .Z(n6215) );
  NANDN U7011 ( .A(rst), .B(n6215), .Z(n6216) );
  NAND U7012 ( .A(n6217), .B(n6216), .Z(n1770) );
  NAND U7013 ( .A(c[234]), .B(rst), .Z(n6222) );
  XNOR U7014 ( .A(n6219), .B(n6218), .Z(n6220) );
  NANDN U7015 ( .A(rst), .B(n6220), .Z(n6221) );
  NAND U7016 ( .A(n6222), .B(n6221), .Z(n1771) );
  NAND U7017 ( .A(c[235]), .B(rst), .Z(n6227) );
  XOR U7018 ( .A(n6224), .B(n6223), .Z(n6225) );
  NANDN U7019 ( .A(rst), .B(n6225), .Z(n6226) );
  NAND U7020 ( .A(n6227), .B(n6226), .Z(n1772) );
  NAND U7021 ( .A(c[236]), .B(rst), .Z(n6232) );
  XNOR U7022 ( .A(n6229), .B(n6228), .Z(n6230) );
  NANDN U7023 ( .A(rst), .B(n6230), .Z(n6231) );
  NAND U7024 ( .A(n6232), .B(n6231), .Z(n1773) );
  NAND U7025 ( .A(c[237]), .B(rst), .Z(n6237) );
  XNOR U7026 ( .A(n6234), .B(n6233), .Z(n6235) );
  NANDN U7027 ( .A(rst), .B(n6235), .Z(n6236) );
  NAND U7028 ( .A(n6237), .B(n6236), .Z(n1774) );
  NAND U7029 ( .A(c[238]), .B(rst), .Z(n6242) );
  XNOR U7030 ( .A(n6239), .B(n6238), .Z(n6240) );
  NANDN U7031 ( .A(rst), .B(n6240), .Z(n6241) );
  NAND U7032 ( .A(n6242), .B(n6241), .Z(n1775) );
  NAND U7033 ( .A(c[239]), .B(rst), .Z(n6247) );
  XNOR U7034 ( .A(n6244), .B(n6243), .Z(n6245) );
  NANDN U7035 ( .A(rst), .B(n6245), .Z(n6246) );
  NAND U7036 ( .A(n6247), .B(n6246), .Z(n1776) );
  NAND U7037 ( .A(c[240]), .B(rst), .Z(n6252) );
  XOR U7038 ( .A(n6249), .B(n6248), .Z(n6250) );
  NANDN U7039 ( .A(rst), .B(n6250), .Z(n6251) );
  NAND U7040 ( .A(n6252), .B(n6251), .Z(n1777) );
  NAND U7041 ( .A(c[241]), .B(rst), .Z(n6257) );
  XNOR U7042 ( .A(n6254), .B(n6253), .Z(n6255) );
  NANDN U7043 ( .A(rst), .B(n6255), .Z(n6256) );
  NAND U7044 ( .A(n6257), .B(n6256), .Z(n1778) );
  NAND U7045 ( .A(c[242]), .B(rst), .Z(n6262) );
  XOR U7046 ( .A(n6259), .B(n6258), .Z(n6260) );
  NANDN U7047 ( .A(rst), .B(n6260), .Z(n6261) );
  NAND U7048 ( .A(n6262), .B(n6261), .Z(n1779) );
  NAND U7049 ( .A(c[243]), .B(rst), .Z(n6267) );
  XNOR U7050 ( .A(n6264), .B(n6263), .Z(n6265) );
  NANDN U7051 ( .A(rst), .B(n6265), .Z(n6266) );
  NAND U7052 ( .A(n6267), .B(n6266), .Z(n1780) );
  NAND U7053 ( .A(c[244]), .B(rst), .Z(n6272) );
  XOR U7054 ( .A(n6269), .B(n6268), .Z(n6270) );
  NANDN U7055 ( .A(rst), .B(n6270), .Z(n6271) );
  NAND U7056 ( .A(n6272), .B(n6271), .Z(n1781) );
  NAND U7057 ( .A(c[245]), .B(rst), .Z(n6277) );
  XNOR U7058 ( .A(n6274), .B(n6273), .Z(n6275) );
  NANDN U7059 ( .A(rst), .B(n6275), .Z(n6276) );
  NAND U7060 ( .A(n6277), .B(n6276), .Z(n1782) );
  NAND U7061 ( .A(c[246]), .B(rst), .Z(n6282) );
  XOR U7062 ( .A(n6279), .B(n6278), .Z(n6280) );
  NANDN U7063 ( .A(rst), .B(n6280), .Z(n6281) );
  NAND U7064 ( .A(n6282), .B(n6281), .Z(n1783) );
  NAND U7065 ( .A(c[247]), .B(rst), .Z(n6287) );
  XNOR U7066 ( .A(n6284), .B(n6283), .Z(n6285) );
  NANDN U7067 ( .A(rst), .B(n6285), .Z(n6286) );
  NAND U7068 ( .A(n6287), .B(n6286), .Z(n1784) );
  NAND U7069 ( .A(c[248]), .B(rst), .Z(n6292) );
  XOR U7070 ( .A(n6289), .B(n6288), .Z(n6290) );
  NANDN U7071 ( .A(rst), .B(n6290), .Z(n6291) );
  NAND U7072 ( .A(n6292), .B(n6291), .Z(n1785) );
  NAND U7073 ( .A(c[249]), .B(rst), .Z(n6297) );
  XNOR U7074 ( .A(n6294), .B(n6293), .Z(n6295) );
  NANDN U7075 ( .A(rst), .B(n6295), .Z(n6296) );
  NAND U7076 ( .A(n6297), .B(n6296), .Z(n1786) );
  NAND U7077 ( .A(c[250]), .B(rst), .Z(n6302) );
  XOR U7078 ( .A(n6299), .B(n6298), .Z(n6300) );
  NANDN U7079 ( .A(rst), .B(n6300), .Z(n6301) );
  NAND U7080 ( .A(n6302), .B(n6301), .Z(n1787) );
  NAND U7081 ( .A(c[251]), .B(rst), .Z(n6307) );
  XNOR U7082 ( .A(n6304), .B(n6303), .Z(n6305) );
  NANDN U7083 ( .A(rst), .B(n6305), .Z(n6306) );
  NAND U7084 ( .A(n6307), .B(n6306), .Z(n1788) );
  NAND U7085 ( .A(c[252]), .B(rst), .Z(n6312) );
  XOR U7086 ( .A(n6309), .B(n6308), .Z(n6310) );
  NANDN U7087 ( .A(rst), .B(n6310), .Z(n6311) );
  NAND U7088 ( .A(n6312), .B(n6311), .Z(n1789) );
  NAND U7089 ( .A(c[253]), .B(rst), .Z(n6317) );
  XNOR U7090 ( .A(n6314), .B(n6313), .Z(n6315) );
  NANDN U7091 ( .A(rst), .B(n6315), .Z(n6316) );
  NAND U7092 ( .A(n6317), .B(n6316), .Z(n1790) );
  NAND U7093 ( .A(c[254]), .B(rst), .Z(n6322) );
  XOR U7094 ( .A(n6319), .B(n6318), .Z(n6320) );
  NANDN U7095 ( .A(rst), .B(n6320), .Z(n6321) );
  NAND U7096 ( .A(n6322), .B(n6321), .Z(n1791) );
  NAND U7097 ( .A(c[255]), .B(rst), .Z(n6327) );
  XNOR U7098 ( .A(n6324), .B(n6323), .Z(n6325) );
  NANDN U7099 ( .A(rst), .B(n6325), .Z(n6326) );
  NAND U7100 ( .A(n6327), .B(n6326), .Z(n1792) );
  NAND U7101 ( .A(c[256]), .B(rst), .Z(n6332) );
  XOR U7102 ( .A(n6329), .B(n6328), .Z(n6330) );
  NANDN U7103 ( .A(rst), .B(n6330), .Z(n6331) );
  NAND U7104 ( .A(n6332), .B(n6331), .Z(n1793) );
  NAND U7105 ( .A(c[257]), .B(rst), .Z(n6337) );
  XNOR U7106 ( .A(n6334), .B(n6333), .Z(n6335) );
  NANDN U7107 ( .A(rst), .B(n6335), .Z(n6336) );
  NAND U7108 ( .A(n6337), .B(n6336), .Z(n1794) );
  NAND U7109 ( .A(c[258]), .B(rst), .Z(n6342) );
  XOR U7110 ( .A(n6339), .B(n6338), .Z(n6340) );
  NANDN U7111 ( .A(rst), .B(n6340), .Z(n6341) );
  NAND U7112 ( .A(n6342), .B(n6341), .Z(n1795) );
  NAND U7113 ( .A(c[259]), .B(rst), .Z(n6347) );
  XNOR U7114 ( .A(n6344), .B(n6343), .Z(n6345) );
  NANDN U7115 ( .A(rst), .B(n6345), .Z(n6346) );
  NAND U7116 ( .A(n6347), .B(n6346), .Z(n1796) );
  NAND U7117 ( .A(c[260]), .B(rst), .Z(n6352) );
  XOR U7118 ( .A(n6349), .B(n6348), .Z(n6350) );
  NANDN U7119 ( .A(rst), .B(n6350), .Z(n6351) );
  NAND U7120 ( .A(n6352), .B(n6351), .Z(n1797) );
  NAND U7121 ( .A(c[261]), .B(rst), .Z(n6357) );
  XNOR U7122 ( .A(n6354), .B(n6353), .Z(n6355) );
  NANDN U7123 ( .A(rst), .B(n6355), .Z(n6356) );
  NAND U7124 ( .A(n6357), .B(n6356), .Z(n1798) );
  NAND U7125 ( .A(c[262]), .B(rst), .Z(n6362) );
  XOR U7126 ( .A(n6359), .B(n6358), .Z(n6360) );
  NANDN U7127 ( .A(rst), .B(n6360), .Z(n6361) );
  NAND U7128 ( .A(n6362), .B(n6361), .Z(n1799) );
  NAND U7129 ( .A(c[263]), .B(rst), .Z(n6367) );
  XNOR U7130 ( .A(n6364), .B(n6363), .Z(n6365) );
  NANDN U7131 ( .A(rst), .B(n6365), .Z(n6366) );
  NAND U7132 ( .A(n6367), .B(n6366), .Z(n1800) );
  NAND U7133 ( .A(c[264]), .B(rst), .Z(n6372) );
  XOR U7134 ( .A(n6369), .B(n6368), .Z(n6370) );
  NANDN U7135 ( .A(rst), .B(n6370), .Z(n6371) );
  NAND U7136 ( .A(n6372), .B(n6371), .Z(n1801) );
  NAND U7137 ( .A(c[265]), .B(rst), .Z(n6377) );
  XNOR U7138 ( .A(n6374), .B(n6373), .Z(n6375) );
  NANDN U7139 ( .A(rst), .B(n6375), .Z(n6376) );
  NAND U7140 ( .A(n6377), .B(n6376), .Z(n1802) );
  NAND U7141 ( .A(c[266]), .B(rst), .Z(n6382) );
  XOR U7142 ( .A(n6379), .B(n6378), .Z(n6380) );
  NANDN U7143 ( .A(rst), .B(n6380), .Z(n6381) );
  NAND U7144 ( .A(n6382), .B(n6381), .Z(n1803) );
  NAND U7145 ( .A(c[267]), .B(rst), .Z(n6387) );
  XNOR U7146 ( .A(n6384), .B(n6383), .Z(n6385) );
  NANDN U7147 ( .A(rst), .B(n6385), .Z(n6386) );
  NAND U7148 ( .A(n6387), .B(n6386), .Z(n1804) );
  NAND U7149 ( .A(c[268]), .B(rst), .Z(n6392) );
  XOR U7150 ( .A(n6389), .B(n6388), .Z(n6390) );
  NANDN U7151 ( .A(rst), .B(n6390), .Z(n6391) );
  NAND U7152 ( .A(n6392), .B(n6391), .Z(n1805) );
  NAND U7153 ( .A(c[269]), .B(rst), .Z(n6397) );
  XNOR U7154 ( .A(n6394), .B(n6393), .Z(n6395) );
  NANDN U7155 ( .A(rst), .B(n6395), .Z(n6396) );
  NAND U7156 ( .A(n6397), .B(n6396), .Z(n1806) );
  NAND U7157 ( .A(c[270]), .B(rst), .Z(n6402) );
  XOR U7158 ( .A(n6399), .B(n6398), .Z(n6400) );
  NANDN U7159 ( .A(rst), .B(n6400), .Z(n6401) );
  NAND U7160 ( .A(n6402), .B(n6401), .Z(n1807) );
  NAND U7161 ( .A(c[271]), .B(rst), .Z(n6407) );
  XNOR U7162 ( .A(n6404), .B(n6403), .Z(n6405) );
  NANDN U7163 ( .A(rst), .B(n6405), .Z(n6406) );
  NAND U7164 ( .A(n6407), .B(n6406), .Z(n1808) );
  NAND U7165 ( .A(c[272]), .B(rst), .Z(n6412) );
  XOR U7166 ( .A(n6409), .B(n6408), .Z(n6410) );
  NANDN U7167 ( .A(rst), .B(n6410), .Z(n6411) );
  NAND U7168 ( .A(n6412), .B(n6411), .Z(n1809) );
  NAND U7169 ( .A(c[273]), .B(rst), .Z(n6417) );
  XNOR U7170 ( .A(n6414), .B(n6413), .Z(n6415) );
  NANDN U7171 ( .A(rst), .B(n6415), .Z(n6416) );
  NAND U7172 ( .A(n6417), .B(n6416), .Z(n1810) );
  NAND U7173 ( .A(c[274]), .B(rst), .Z(n6422) );
  XOR U7174 ( .A(n6419), .B(n6418), .Z(n6420) );
  NANDN U7175 ( .A(rst), .B(n6420), .Z(n6421) );
  NAND U7176 ( .A(n6422), .B(n6421), .Z(n1811) );
  NAND U7177 ( .A(c[275]), .B(rst), .Z(n6427) );
  XNOR U7178 ( .A(n6424), .B(n6423), .Z(n6425) );
  NANDN U7179 ( .A(rst), .B(n6425), .Z(n6426) );
  NAND U7180 ( .A(n6427), .B(n6426), .Z(n1812) );
  NAND U7181 ( .A(c[276]), .B(rst), .Z(n6432) );
  XOR U7182 ( .A(n6429), .B(n6428), .Z(n6430) );
  NANDN U7183 ( .A(rst), .B(n6430), .Z(n6431) );
  NAND U7184 ( .A(n6432), .B(n6431), .Z(n1813) );
  NAND U7185 ( .A(c[277]), .B(rst), .Z(n6437) );
  XNOR U7186 ( .A(n6434), .B(n6433), .Z(n6435) );
  NANDN U7187 ( .A(rst), .B(n6435), .Z(n6436) );
  NAND U7188 ( .A(n6437), .B(n6436), .Z(n1814) );
  NAND U7189 ( .A(c[278]), .B(rst), .Z(n6442) );
  XOR U7190 ( .A(n6439), .B(n6438), .Z(n6440) );
  NANDN U7191 ( .A(rst), .B(n6440), .Z(n6441) );
  NAND U7192 ( .A(n6442), .B(n6441), .Z(n1815) );
  NAND U7193 ( .A(c[279]), .B(rst), .Z(n6447) );
  XNOR U7194 ( .A(n6444), .B(n6443), .Z(n6445) );
  NANDN U7195 ( .A(rst), .B(n6445), .Z(n6446) );
  NAND U7196 ( .A(n6447), .B(n6446), .Z(n1816) );
  NAND U7197 ( .A(c[280]), .B(rst), .Z(n6452) );
  XNOR U7198 ( .A(n6449), .B(n6448), .Z(n6450) );
  NANDN U7199 ( .A(rst), .B(n6450), .Z(n6451) );
  NAND U7200 ( .A(n6452), .B(n6451), .Z(n1817) );
  NAND U7201 ( .A(c[281]), .B(rst), .Z(n6457) );
  XNOR U7202 ( .A(n6454), .B(n6453), .Z(n6455) );
  NANDN U7203 ( .A(rst), .B(n6455), .Z(n6456) );
  NAND U7204 ( .A(n6457), .B(n6456), .Z(n1818) );
  NAND U7205 ( .A(c[282]), .B(rst), .Z(n6462) );
  XNOR U7206 ( .A(n6459), .B(n6458), .Z(n6460) );
  NANDN U7207 ( .A(rst), .B(n6460), .Z(n6461) );
  NAND U7208 ( .A(n6462), .B(n6461), .Z(n1819) );
  NAND U7209 ( .A(c[283]), .B(rst), .Z(n6467) );
  XOR U7210 ( .A(n6464), .B(n6463), .Z(n6465) );
  NANDN U7211 ( .A(rst), .B(n6465), .Z(n6466) );
  NAND U7212 ( .A(n6467), .B(n6466), .Z(n1820) );
  NAND U7213 ( .A(c[284]), .B(rst), .Z(n6472) );
  XNOR U7214 ( .A(n6469), .B(n6468), .Z(n6470) );
  NANDN U7215 ( .A(rst), .B(n6470), .Z(n6471) );
  NAND U7216 ( .A(n6472), .B(n6471), .Z(n1821) );
  NAND U7217 ( .A(c[285]), .B(rst), .Z(n6477) );
  XNOR U7218 ( .A(n6474), .B(n6473), .Z(n6475) );
  NANDN U7219 ( .A(rst), .B(n6475), .Z(n6476) );
  NAND U7220 ( .A(n6477), .B(n6476), .Z(n1822) );
  NAND U7221 ( .A(c[286]), .B(rst), .Z(n6482) );
  XNOR U7222 ( .A(n6479), .B(n6478), .Z(n6480) );
  NANDN U7223 ( .A(rst), .B(n6480), .Z(n6481) );
  NAND U7224 ( .A(n6482), .B(n6481), .Z(n1823) );
  NAND U7225 ( .A(c[287]), .B(rst), .Z(n6487) );
  XNOR U7226 ( .A(n6484), .B(n6483), .Z(n6485) );
  NANDN U7227 ( .A(rst), .B(n6485), .Z(n6486) );
  NAND U7228 ( .A(n6487), .B(n6486), .Z(n1824) );
  NAND U7229 ( .A(c[288]), .B(rst), .Z(n6492) );
  XOR U7230 ( .A(n6489), .B(n6488), .Z(n6490) );
  NANDN U7231 ( .A(rst), .B(n6490), .Z(n6491) );
  NAND U7232 ( .A(n6492), .B(n6491), .Z(n1825) );
  NAND U7233 ( .A(c[289]), .B(rst), .Z(n6497) );
  XNOR U7234 ( .A(n6494), .B(n6493), .Z(n6495) );
  NANDN U7235 ( .A(rst), .B(n6495), .Z(n6496) );
  NAND U7236 ( .A(n6497), .B(n6496), .Z(n1826) );
  NAND U7237 ( .A(c[290]), .B(rst), .Z(n6502) );
  XOR U7238 ( .A(n6499), .B(n6498), .Z(n6500) );
  NANDN U7239 ( .A(rst), .B(n6500), .Z(n6501) );
  NAND U7240 ( .A(n6502), .B(n6501), .Z(n1827) );
  NAND U7241 ( .A(c[291]), .B(rst), .Z(n6507) );
  XNOR U7242 ( .A(n6504), .B(n6503), .Z(n6505) );
  NANDN U7243 ( .A(rst), .B(n6505), .Z(n6506) );
  NAND U7244 ( .A(n6507), .B(n6506), .Z(n1828) );
  NAND U7245 ( .A(c[292]), .B(rst), .Z(n6512) );
  XOR U7246 ( .A(n6509), .B(n6508), .Z(n6510) );
  NANDN U7247 ( .A(rst), .B(n6510), .Z(n6511) );
  NAND U7248 ( .A(n6512), .B(n6511), .Z(n1829) );
  NAND U7249 ( .A(c[293]), .B(rst), .Z(n6517) );
  XNOR U7250 ( .A(n6514), .B(n6513), .Z(n6515) );
  NANDN U7251 ( .A(rst), .B(n6515), .Z(n6516) );
  NAND U7252 ( .A(n6517), .B(n6516), .Z(n1830) );
  NAND U7253 ( .A(c[294]), .B(rst), .Z(n6522) );
  XNOR U7254 ( .A(n6519), .B(n6518), .Z(n6520) );
  NANDN U7255 ( .A(rst), .B(n6520), .Z(n6521) );
  NAND U7256 ( .A(n6522), .B(n6521), .Z(n1831) );
  NAND U7257 ( .A(c[295]), .B(rst), .Z(n6527) );
  XNOR U7258 ( .A(n6524), .B(n6523), .Z(n6525) );
  NANDN U7259 ( .A(rst), .B(n6525), .Z(n6526) );
  NAND U7260 ( .A(n6527), .B(n6526), .Z(n1832) );
  NAND U7261 ( .A(c[296]), .B(rst), .Z(n6532) );
  XNOR U7262 ( .A(n6529), .B(n6528), .Z(n6530) );
  NANDN U7263 ( .A(rst), .B(n6530), .Z(n6531) );
  NAND U7264 ( .A(n6532), .B(n6531), .Z(n1833) );
  NAND U7265 ( .A(c[297]), .B(rst), .Z(n6537) );
  XOR U7266 ( .A(n6534), .B(n6533), .Z(n6535) );
  NANDN U7267 ( .A(rst), .B(n6535), .Z(n6536) );
  NAND U7268 ( .A(n6537), .B(n6536), .Z(n1834) );
  NAND U7269 ( .A(c[298]), .B(rst), .Z(n6542) );
  XNOR U7270 ( .A(n6539), .B(n6538), .Z(n6540) );
  NANDN U7271 ( .A(rst), .B(n6540), .Z(n6541) );
  NAND U7272 ( .A(n6542), .B(n6541), .Z(n1835) );
  NAND U7273 ( .A(c[299]), .B(rst), .Z(n6547) );
  XOR U7274 ( .A(n6544), .B(n6543), .Z(n6545) );
  NANDN U7275 ( .A(rst), .B(n6545), .Z(n6546) );
  NAND U7276 ( .A(n6547), .B(n6546), .Z(n1836) );
  NAND U7277 ( .A(c[300]), .B(rst), .Z(n6552) );
  XNOR U7278 ( .A(n6549), .B(n6548), .Z(n6550) );
  NANDN U7279 ( .A(rst), .B(n6550), .Z(n6551) );
  NAND U7280 ( .A(n6552), .B(n6551), .Z(n1837) );
  NAND U7281 ( .A(c[301]), .B(rst), .Z(n6557) );
  XOR U7282 ( .A(n6554), .B(n6553), .Z(n6555) );
  NANDN U7283 ( .A(rst), .B(n6555), .Z(n6556) );
  NAND U7284 ( .A(n6557), .B(n6556), .Z(n1838) );
  NAND U7285 ( .A(c[302]), .B(rst), .Z(n6562) );
  XNOR U7286 ( .A(n6559), .B(n6558), .Z(n6560) );
  NANDN U7287 ( .A(rst), .B(n6560), .Z(n6561) );
  NAND U7288 ( .A(n6562), .B(n6561), .Z(n1839) );
  NAND U7289 ( .A(c[303]), .B(rst), .Z(n6567) );
  XOR U7290 ( .A(n6564), .B(n6563), .Z(n6565) );
  NANDN U7291 ( .A(rst), .B(n6565), .Z(n6566) );
  NAND U7292 ( .A(n6567), .B(n6566), .Z(n1840) );
  NAND U7293 ( .A(c[304]), .B(rst), .Z(n6572) );
  XNOR U7294 ( .A(n6569), .B(n6568), .Z(n6570) );
  NANDN U7295 ( .A(rst), .B(n6570), .Z(n6571) );
  NAND U7296 ( .A(n6572), .B(n6571), .Z(n1841) );
  NAND U7297 ( .A(c[305]), .B(rst), .Z(n6577) );
  XOR U7298 ( .A(n6574), .B(n6573), .Z(n6575) );
  NANDN U7299 ( .A(rst), .B(n6575), .Z(n6576) );
  NAND U7300 ( .A(n6577), .B(n6576), .Z(n1842) );
  NAND U7301 ( .A(c[306]), .B(rst), .Z(n6582) );
  XNOR U7302 ( .A(n6579), .B(n6578), .Z(n6580) );
  NANDN U7303 ( .A(rst), .B(n6580), .Z(n6581) );
  NAND U7304 ( .A(n6582), .B(n6581), .Z(n1843) );
  NAND U7305 ( .A(c[307]), .B(rst), .Z(n6587) );
  XOR U7306 ( .A(n6584), .B(n6583), .Z(n6585) );
  NANDN U7307 ( .A(rst), .B(n6585), .Z(n6586) );
  NAND U7308 ( .A(n6587), .B(n6586), .Z(n1844) );
  NAND U7309 ( .A(c[308]), .B(rst), .Z(n6592) );
  XNOR U7310 ( .A(n6589), .B(n6588), .Z(n6590) );
  NANDN U7311 ( .A(rst), .B(n6590), .Z(n6591) );
  NAND U7312 ( .A(n6592), .B(n6591), .Z(n1845) );
  NAND U7313 ( .A(c[309]), .B(rst), .Z(n6597) );
  XOR U7314 ( .A(n6594), .B(n6593), .Z(n6595) );
  NANDN U7315 ( .A(rst), .B(n6595), .Z(n6596) );
  NAND U7316 ( .A(n6597), .B(n6596), .Z(n1846) );
  NAND U7317 ( .A(c[310]), .B(rst), .Z(n6602) );
  XNOR U7318 ( .A(n6599), .B(n6598), .Z(n6600) );
  NANDN U7319 ( .A(rst), .B(n6600), .Z(n6601) );
  NAND U7320 ( .A(n6602), .B(n6601), .Z(n1847) );
  NAND U7321 ( .A(c[311]), .B(rst), .Z(n6607) );
  XOR U7322 ( .A(n6604), .B(n6603), .Z(n6605) );
  NANDN U7323 ( .A(rst), .B(n6605), .Z(n6606) );
  NAND U7324 ( .A(n6607), .B(n6606), .Z(n1848) );
  NAND U7325 ( .A(c[312]), .B(rst), .Z(n6612) );
  XNOR U7326 ( .A(n6609), .B(n6608), .Z(n6610) );
  NANDN U7327 ( .A(rst), .B(n6610), .Z(n6611) );
  NAND U7328 ( .A(n6612), .B(n6611), .Z(n1849) );
  NAND U7329 ( .A(c[313]), .B(rst), .Z(n6617) );
  XNOR U7330 ( .A(n6614), .B(n6613), .Z(n6615) );
  NANDN U7331 ( .A(rst), .B(n6615), .Z(n6616) );
  NAND U7332 ( .A(n6617), .B(n6616), .Z(n1850) );
  NAND U7333 ( .A(c[314]), .B(rst), .Z(n6622) );
  XNOR U7334 ( .A(n6619), .B(n6618), .Z(n6620) );
  NANDN U7335 ( .A(rst), .B(n6620), .Z(n6621) );
  NAND U7336 ( .A(n6622), .B(n6621), .Z(n1851) );
  NAND U7337 ( .A(c[315]), .B(rst), .Z(n6627) );
  XNOR U7338 ( .A(n6624), .B(n6623), .Z(n6625) );
  NANDN U7339 ( .A(rst), .B(n6625), .Z(n6626) );
  NAND U7340 ( .A(n6627), .B(n6626), .Z(n1852) );
  NAND U7341 ( .A(c[316]), .B(rst), .Z(n6632) );
  XOR U7342 ( .A(n6629), .B(n6628), .Z(n6630) );
  NANDN U7343 ( .A(rst), .B(n6630), .Z(n6631) );
  NAND U7344 ( .A(n6632), .B(n6631), .Z(n1853) );
  NAND U7345 ( .A(c[317]), .B(rst), .Z(n6637) );
  XNOR U7346 ( .A(n6634), .B(n6633), .Z(n6635) );
  NANDN U7347 ( .A(rst), .B(n6635), .Z(n6636) );
  NAND U7348 ( .A(n6637), .B(n6636), .Z(n1854) );
  NAND U7349 ( .A(c[318]), .B(rst), .Z(n6642) );
  XNOR U7350 ( .A(n6639), .B(n6638), .Z(n6640) );
  NANDN U7351 ( .A(rst), .B(n6640), .Z(n6641) );
  NAND U7352 ( .A(n6642), .B(n6641), .Z(n1855) );
  NAND U7353 ( .A(c[319]), .B(rst), .Z(n6647) );
  XNOR U7354 ( .A(n6644), .B(n6643), .Z(n6645) );
  NANDN U7355 ( .A(rst), .B(n6645), .Z(n6646) );
  NAND U7356 ( .A(n6647), .B(n6646), .Z(n1856) );
  NAND U7357 ( .A(c[320]), .B(rst), .Z(n6652) );
  XNOR U7358 ( .A(n6649), .B(n6648), .Z(n6650) );
  NANDN U7359 ( .A(rst), .B(n6650), .Z(n6651) );
  NAND U7360 ( .A(n6652), .B(n6651), .Z(n1857) );
  NAND U7361 ( .A(c[321]), .B(rst), .Z(n6657) );
  XOR U7362 ( .A(n6654), .B(n6653), .Z(n6655) );
  NANDN U7363 ( .A(rst), .B(n6655), .Z(n6656) );
  NAND U7364 ( .A(n6657), .B(n6656), .Z(n1858) );
  NAND U7365 ( .A(c[322]), .B(rst), .Z(n6662) );
  XNOR U7366 ( .A(n6659), .B(n6658), .Z(n6660) );
  NANDN U7367 ( .A(rst), .B(n6660), .Z(n6661) );
  NAND U7368 ( .A(n6662), .B(n6661), .Z(n1859) );
  NAND U7369 ( .A(c[323]), .B(rst), .Z(n6667) );
  XOR U7370 ( .A(n6664), .B(n6663), .Z(n6665) );
  NANDN U7371 ( .A(rst), .B(n6665), .Z(n6666) );
  NAND U7372 ( .A(n6667), .B(n6666), .Z(n1860) );
  NAND U7373 ( .A(c[324]), .B(rst), .Z(n6672) );
  XNOR U7374 ( .A(n6669), .B(n6668), .Z(n6670) );
  NANDN U7375 ( .A(rst), .B(n6670), .Z(n6671) );
  NAND U7376 ( .A(n6672), .B(n6671), .Z(n1861) );
  NAND U7377 ( .A(c[325]), .B(rst), .Z(n6677) );
  XOR U7378 ( .A(n6674), .B(n6673), .Z(n6675) );
  NANDN U7379 ( .A(rst), .B(n6675), .Z(n6676) );
  NAND U7380 ( .A(n6677), .B(n6676), .Z(n1862) );
  NAND U7381 ( .A(c[326]), .B(rst), .Z(n6682) );
  XNOR U7382 ( .A(n6679), .B(n6678), .Z(n6680) );
  NANDN U7383 ( .A(rst), .B(n6680), .Z(n6681) );
  NAND U7384 ( .A(n6682), .B(n6681), .Z(n1863) );
  NAND U7385 ( .A(c[327]), .B(rst), .Z(n6687) );
  XOR U7386 ( .A(n6684), .B(n6683), .Z(n6685) );
  NANDN U7387 ( .A(rst), .B(n6685), .Z(n6686) );
  NAND U7388 ( .A(n6687), .B(n6686), .Z(n1864) );
  NAND U7389 ( .A(c[328]), .B(rst), .Z(n6692) );
  XNOR U7390 ( .A(n6689), .B(n6688), .Z(n6690) );
  NANDN U7391 ( .A(rst), .B(n6690), .Z(n6691) );
  NAND U7392 ( .A(n6692), .B(n6691), .Z(n1865) );
  NAND U7393 ( .A(c[329]), .B(rst), .Z(n6697) );
  XNOR U7394 ( .A(n6694), .B(n6693), .Z(n6695) );
  NANDN U7395 ( .A(rst), .B(n6695), .Z(n6696) );
  NAND U7396 ( .A(n6697), .B(n6696), .Z(n1866) );
  NAND U7397 ( .A(c[330]), .B(rst), .Z(n6702) );
  XNOR U7398 ( .A(n6699), .B(n6698), .Z(n6700) );
  NANDN U7399 ( .A(rst), .B(n6700), .Z(n6701) );
  NAND U7400 ( .A(n6702), .B(n6701), .Z(n1867) );
  NAND U7401 ( .A(c[331]), .B(rst), .Z(n6707) );
  XNOR U7402 ( .A(n6704), .B(n6703), .Z(n6705) );
  NANDN U7403 ( .A(rst), .B(n6705), .Z(n6706) );
  NAND U7404 ( .A(n6707), .B(n6706), .Z(n1868) );
  NAND U7405 ( .A(c[332]), .B(rst), .Z(n6712) );
  XOR U7406 ( .A(n6709), .B(n6708), .Z(n6710) );
  NANDN U7407 ( .A(rst), .B(n6710), .Z(n6711) );
  NAND U7408 ( .A(n6712), .B(n6711), .Z(n1869) );
  NAND U7409 ( .A(c[333]), .B(rst), .Z(n6717) );
  XNOR U7410 ( .A(n6714), .B(n6713), .Z(n6715) );
  NANDN U7411 ( .A(rst), .B(n6715), .Z(n6716) );
  NAND U7412 ( .A(n6717), .B(n6716), .Z(n1870) );
  NAND U7413 ( .A(c[334]), .B(rst), .Z(n6722) );
  XOR U7414 ( .A(n6719), .B(n6718), .Z(n6720) );
  NANDN U7415 ( .A(rst), .B(n6720), .Z(n6721) );
  NAND U7416 ( .A(n6722), .B(n6721), .Z(n1871) );
  NAND U7417 ( .A(c[335]), .B(rst), .Z(n6727) );
  XNOR U7418 ( .A(n6724), .B(n6723), .Z(n6725) );
  NANDN U7419 ( .A(rst), .B(n6725), .Z(n6726) );
  NAND U7420 ( .A(n6727), .B(n6726), .Z(n1872) );
  NAND U7421 ( .A(c[336]), .B(rst), .Z(n6732) );
  XOR U7422 ( .A(n6729), .B(n6728), .Z(n6730) );
  NANDN U7423 ( .A(rst), .B(n6730), .Z(n6731) );
  NAND U7424 ( .A(n6732), .B(n6731), .Z(n1873) );
  NAND U7425 ( .A(c[337]), .B(rst), .Z(n6737) );
  XNOR U7426 ( .A(n6734), .B(n6733), .Z(n6735) );
  NANDN U7427 ( .A(rst), .B(n6735), .Z(n6736) );
  NAND U7428 ( .A(n6737), .B(n6736), .Z(n1874) );
  NAND U7429 ( .A(c[338]), .B(rst), .Z(n6742) );
  XOR U7430 ( .A(n6739), .B(n6738), .Z(n6740) );
  NANDN U7431 ( .A(rst), .B(n6740), .Z(n6741) );
  NAND U7432 ( .A(n6742), .B(n6741), .Z(n1875) );
  NAND U7433 ( .A(c[339]), .B(rst), .Z(n6747) );
  XNOR U7434 ( .A(n6744), .B(n6743), .Z(n6745) );
  NANDN U7435 ( .A(rst), .B(n6745), .Z(n6746) );
  NAND U7436 ( .A(n6747), .B(n6746), .Z(n1876) );
  NAND U7437 ( .A(c[340]), .B(rst), .Z(n6752) );
  XOR U7438 ( .A(n6749), .B(n6748), .Z(n6750) );
  NANDN U7439 ( .A(rst), .B(n6750), .Z(n6751) );
  NAND U7440 ( .A(n6752), .B(n6751), .Z(n1877) );
  NAND U7441 ( .A(c[341]), .B(rst), .Z(n6757) );
  XNOR U7442 ( .A(n6754), .B(n6753), .Z(n6755) );
  NANDN U7443 ( .A(rst), .B(n6755), .Z(n6756) );
  NAND U7444 ( .A(n6757), .B(n6756), .Z(n1878) );
  NAND U7445 ( .A(c[342]), .B(rst), .Z(n6762) );
  XOR U7446 ( .A(n6759), .B(n6758), .Z(n6760) );
  NANDN U7447 ( .A(rst), .B(n6760), .Z(n6761) );
  NAND U7448 ( .A(n6762), .B(n6761), .Z(n1879) );
  NAND U7449 ( .A(c[343]), .B(rst), .Z(n6767) );
  XNOR U7450 ( .A(n6764), .B(n6763), .Z(n6765) );
  NANDN U7451 ( .A(rst), .B(n6765), .Z(n6766) );
  NAND U7452 ( .A(n6767), .B(n6766), .Z(n1880) );
  NAND U7453 ( .A(c[344]), .B(rst), .Z(n6772) );
  XOR U7454 ( .A(n6769), .B(n6768), .Z(n6770) );
  NANDN U7455 ( .A(rst), .B(n6770), .Z(n6771) );
  NAND U7456 ( .A(n6772), .B(n6771), .Z(n1881) );
  NAND U7457 ( .A(c[345]), .B(rst), .Z(n6777) );
  XNOR U7458 ( .A(n6774), .B(n6773), .Z(n6775) );
  NANDN U7459 ( .A(rst), .B(n6775), .Z(n6776) );
  NAND U7460 ( .A(n6777), .B(n6776), .Z(n1882) );
  NAND U7461 ( .A(c[346]), .B(rst), .Z(n6782) );
  XNOR U7462 ( .A(n6779), .B(n6778), .Z(n6780) );
  NANDN U7463 ( .A(rst), .B(n6780), .Z(n6781) );
  NAND U7464 ( .A(n6782), .B(n6781), .Z(n1883) );
  NAND U7465 ( .A(c[347]), .B(rst), .Z(n6787) );
  XNOR U7466 ( .A(n6784), .B(n6783), .Z(n6785) );
  NANDN U7467 ( .A(rst), .B(n6785), .Z(n6786) );
  NAND U7468 ( .A(n6787), .B(n6786), .Z(n1884) );
  NAND U7469 ( .A(c[348]), .B(rst), .Z(n6792) );
  XNOR U7470 ( .A(n6789), .B(n6788), .Z(n6790) );
  NANDN U7471 ( .A(rst), .B(n6790), .Z(n6791) );
  NAND U7472 ( .A(n6792), .B(n6791), .Z(n1885) );
  NAND U7473 ( .A(c[349]), .B(rst), .Z(n6797) );
  XOR U7474 ( .A(n6794), .B(n6793), .Z(n6795) );
  NANDN U7475 ( .A(rst), .B(n6795), .Z(n6796) );
  NAND U7476 ( .A(n6797), .B(n6796), .Z(n1886) );
  NAND U7477 ( .A(c[350]), .B(rst), .Z(n6802) );
  XNOR U7478 ( .A(n6799), .B(n6798), .Z(n6800) );
  NANDN U7479 ( .A(rst), .B(n6800), .Z(n6801) );
  NAND U7480 ( .A(n6802), .B(n6801), .Z(n1887) );
  NAND U7481 ( .A(c[351]), .B(rst), .Z(n6807) );
  XOR U7482 ( .A(n6804), .B(n6803), .Z(n6805) );
  NANDN U7483 ( .A(rst), .B(n6805), .Z(n6806) );
  NAND U7484 ( .A(n6807), .B(n6806), .Z(n1888) );
  NAND U7485 ( .A(c[352]), .B(rst), .Z(n6812) );
  XNOR U7486 ( .A(n6809), .B(n6808), .Z(n6810) );
  NANDN U7487 ( .A(rst), .B(n6810), .Z(n6811) );
  NAND U7488 ( .A(n6812), .B(n6811), .Z(n1889) );
  NAND U7489 ( .A(c[353]), .B(rst), .Z(n6817) );
  XOR U7490 ( .A(n6814), .B(n6813), .Z(n6815) );
  NANDN U7491 ( .A(rst), .B(n6815), .Z(n6816) );
  NAND U7492 ( .A(n6817), .B(n6816), .Z(n1890) );
  NAND U7493 ( .A(c[354]), .B(rst), .Z(n6822) );
  XNOR U7494 ( .A(n6819), .B(n6818), .Z(n6820) );
  NANDN U7495 ( .A(rst), .B(n6820), .Z(n6821) );
  NAND U7496 ( .A(n6822), .B(n6821), .Z(n1891) );
  NAND U7497 ( .A(c[355]), .B(rst), .Z(n6827) );
  XOR U7498 ( .A(n6824), .B(n6823), .Z(n6825) );
  NANDN U7499 ( .A(rst), .B(n6825), .Z(n6826) );
  NAND U7500 ( .A(n6827), .B(n6826), .Z(n1892) );
  NAND U7501 ( .A(c[356]), .B(rst), .Z(n6832) );
  XNOR U7502 ( .A(n6829), .B(n6828), .Z(n6830) );
  NANDN U7503 ( .A(rst), .B(n6830), .Z(n6831) );
  NAND U7504 ( .A(n6832), .B(n6831), .Z(n1893) );
  NAND U7505 ( .A(c[357]), .B(rst), .Z(n6837) );
  XOR U7506 ( .A(n6834), .B(n6833), .Z(n6835) );
  NANDN U7507 ( .A(rst), .B(n6835), .Z(n6836) );
  NAND U7508 ( .A(n6837), .B(n6836), .Z(n1894) );
  NAND U7509 ( .A(c[358]), .B(rst), .Z(n6842) );
  XNOR U7510 ( .A(n6839), .B(n6838), .Z(n6840) );
  NANDN U7511 ( .A(rst), .B(n6840), .Z(n6841) );
  NAND U7512 ( .A(n6842), .B(n6841), .Z(n1895) );
  NAND U7513 ( .A(c[359]), .B(rst), .Z(n6847) );
  XOR U7514 ( .A(n6844), .B(n6843), .Z(n6845) );
  NANDN U7515 ( .A(rst), .B(n6845), .Z(n6846) );
  NAND U7516 ( .A(n6847), .B(n6846), .Z(n1896) );
  NAND U7517 ( .A(c[360]), .B(rst), .Z(n6852) );
  XNOR U7518 ( .A(n6849), .B(n6848), .Z(n6850) );
  NANDN U7519 ( .A(rst), .B(n6850), .Z(n6851) );
  NAND U7520 ( .A(n6852), .B(n6851), .Z(n1897) );
  NAND U7521 ( .A(c[361]), .B(rst), .Z(n6857) );
  XOR U7522 ( .A(n6854), .B(n6853), .Z(n6855) );
  NANDN U7523 ( .A(rst), .B(n6855), .Z(n6856) );
  NAND U7524 ( .A(n6857), .B(n6856), .Z(n1898) );
  NAND U7525 ( .A(c[362]), .B(rst), .Z(n6862) );
  XNOR U7526 ( .A(n6859), .B(n6858), .Z(n6860) );
  NANDN U7527 ( .A(rst), .B(n6860), .Z(n6861) );
  NAND U7528 ( .A(n6862), .B(n6861), .Z(n1899) );
  NAND U7529 ( .A(c[363]), .B(rst), .Z(n6867) );
  XOR U7530 ( .A(n6864), .B(n6863), .Z(n6865) );
  NANDN U7531 ( .A(rst), .B(n6865), .Z(n6866) );
  NAND U7532 ( .A(n6867), .B(n6866), .Z(n1900) );
  NAND U7533 ( .A(c[364]), .B(rst), .Z(n6872) );
  XNOR U7534 ( .A(n6869), .B(n6868), .Z(n6870) );
  NANDN U7535 ( .A(rst), .B(n6870), .Z(n6871) );
  NAND U7536 ( .A(n6872), .B(n6871), .Z(n1901) );
  NAND U7537 ( .A(c[365]), .B(rst), .Z(n6877) );
  XNOR U7538 ( .A(n6874), .B(n6873), .Z(n6875) );
  NANDN U7539 ( .A(rst), .B(n6875), .Z(n6876) );
  NAND U7540 ( .A(n6877), .B(n6876), .Z(n1902) );
  NAND U7541 ( .A(c[366]), .B(rst), .Z(n6882) );
  XNOR U7542 ( .A(n6879), .B(n6878), .Z(n6880) );
  NANDN U7543 ( .A(rst), .B(n6880), .Z(n6881) );
  NAND U7544 ( .A(n6882), .B(n6881), .Z(n1903) );
  NAND U7545 ( .A(c[367]), .B(rst), .Z(n6887) );
  XNOR U7546 ( .A(n6884), .B(n6883), .Z(n6885) );
  NANDN U7547 ( .A(rst), .B(n6885), .Z(n6886) );
  NAND U7548 ( .A(n6887), .B(n6886), .Z(n1904) );
  NAND U7549 ( .A(c[368]), .B(rst), .Z(n6892) );
  XOR U7550 ( .A(n6889), .B(n6888), .Z(n6890) );
  NANDN U7551 ( .A(rst), .B(n6890), .Z(n6891) );
  NAND U7552 ( .A(n6892), .B(n6891), .Z(n1905) );
  NAND U7553 ( .A(c[369]), .B(rst), .Z(n6897) );
  XNOR U7554 ( .A(n6894), .B(n6893), .Z(n6895) );
  NANDN U7555 ( .A(rst), .B(n6895), .Z(n6896) );
  NAND U7556 ( .A(n6897), .B(n6896), .Z(n1906) );
  NAND U7557 ( .A(c[370]), .B(rst), .Z(n6902) );
  XOR U7558 ( .A(n6899), .B(n6898), .Z(n6900) );
  NANDN U7559 ( .A(rst), .B(n6900), .Z(n6901) );
  NAND U7560 ( .A(n6902), .B(n6901), .Z(n1907) );
  NAND U7561 ( .A(c[371]), .B(rst), .Z(n6907) );
  XNOR U7562 ( .A(n6904), .B(n6903), .Z(n6905) );
  NANDN U7563 ( .A(rst), .B(n6905), .Z(n6906) );
  NAND U7564 ( .A(n6907), .B(n6906), .Z(n1908) );
  NAND U7565 ( .A(c[372]), .B(rst), .Z(n6912) );
  XOR U7566 ( .A(n6909), .B(n6908), .Z(n6910) );
  NANDN U7567 ( .A(rst), .B(n6910), .Z(n6911) );
  NAND U7568 ( .A(n6912), .B(n6911), .Z(n1909) );
  NAND U7569 ( .A(c[373]), .B(rst), .Z(n6917) );
  XNOR U7570 ( .A(n6914), .B(n6913), .Z(n6915) );
  NANDN U7571 ( .A(rst), .B(n6915), .Z(n6916) );
  NAND U7572 ( .A(n6917), .B(n6916), .Z(n1910) );
  NAND U7573 ( .A(c[374]), .B(rst), .Z(n6922) );
  XOR U7574 ( .A(n6919), .B(n6918), .Z(n6920) );
  NANDN U7575 ( .A(rst), .B(n6920), .Z(n6921) );
  NAND U7576 ( .A(n6922), .B(n6921), .Z(n1911) );
  NAND U7577 ( .A(c[375]), .B(rst), .Z(n6927) );
  XNOR U7578 ( .A(n6924), .B(n6923), .Z(n6925) );
  NANDN U7579 ( .A(rst), .B(n6925), .Z(n6926) );
  NAND U7580 ( .A(n6927), .B(n6926), .Z(n1912) );
  NAND U7581 ( .A(c[376]), .B(rst), .Z(n6932) );
  XOR U7582 ( .A(n6929), .B(n6928), .Z(n6930) );
  NANDN U7583 ( .A(rst), .B(n6930), .Z(n6931) );
  NAND U7584 ( .A(n6932), .B(n6931), .Z(n1913) );
  NAND U7585 ( .A(c[377]), .B(rst), .Z(n6937) );
  XNOR U7586 ( .A(n6934), .B(n6933), .Z(n6935) );
  NANDN U7587 ( .A(rst), .B(n6935), .Z(n6936) );
  NAND U7588 ( .A(n6937), .B(n6936), .Z(n1914) );
  NAND U7589 ( .A(c[378]), .B(rst), .Z(n6942) );
  XOR U7590 ( .A(n6939), .B(n6938), .Z(n6940) );
  NANDN U7591 ( .A(rst), .B(n6940), .Z(n6941) );
  NAND U7592 ( .A(n6942), .B(n6941), .Z(n1915) );
  NAND U7593 ( .A(c[379]), .B(rst), .Z(n6947) );
  XNOR U7594 ( .A(n6944), .B(n6943), .Z(n6945) );
  NANDN U7595 ( .A(rst), .B(n6945), .Z(n6946) );
  NAND U7596 ( .A(n6947), .B(n6946), .Z(n1916) );
  NAND U7597 ( .A(c[380]), .B(rst), .Z(n6952) );
  XOR U7598 ( .A(n6949), .B(n6948), .Z(n6950) );
  NANDN U7599 ( .A(rst), .B(n6950), .Z(n6951) );
  NAND U7600 ( .A(n6952), .B(n6951), .Z(n1917) );
  NAND U7601 ( .A(c[381]), .B(rst), .Z(n6957) );
  XNOR U7602 ( .A(n6954), .B(n6953), .Z(n6955) );
  NANDN U7603 ( .A(rst), .B(n6955), .Z(n6956) );
  NAND U7604 ( .A(n6957), .B(n6956), .Z(n1918) );
  NAND U7605 ( .A(c[382]), .B(rst), .Z(n6962) );
  XOR U7606 ( .A(n6959), .B(n6958), .Z(n6960) );
  NANDN U7607 ( .A(rst), .B(n6960), .Z(n6961) );
  NAND U7608 ( .A(n6962), .B(n6961), .Z(n1919) );
  NAND U7609 ( .A(c[383]), .B(rst), .Z(n6967) );
  XNOR U7610 ( .A(n6964), .B(n6963), .Z(n6965) );
  NANDN U7611 ( .A(rst), .B(n6965), .Z(n6966) );
  NAND U7612 ( .A(n6967), .B(n6966), .Z(n1920) );
  NAND U7613 ( .A(c[384]), .B(rst), .Z(n6972) );
  XOR U7614 ( .A(n6969), .B(n6968), .Z(n6970) );
  NANDN U7615 ( .A(rst), .B(n6970), .Z(n6971) );
  NAND U7616 ( .A(n6972), .B(n6971), .Z(n1921) );
  NAND U7617 ( .A(c[385]), .B(rst), .Z(n6977) );
  XNOR U7618 ( .A(n6974), .B(n6973), .Z(n6975) );
  NANDN U7619 ( .A(rst), .B(n6975), .Z(n6976) );
  NAND U7620 ( .A(n6977), .B(n6976), .Z(n1922) );
  NAND U7621 ( .A(c[386]), .B(rst), .Z(n6982) );
  XOR U7622 ( .A(n6979), .B(n6978), .Z(n6980) );
  NANDN U7623 ( .A(rst), .B(n6980), .Z(n6981) );
  NAND U7624 ( .A(n6982), .B(n6981), .Z(n1923) );
  NAND U7625 ( .A(c[387]), .B(rst), .Z(n6987) );
  XNOR U7626 ( .A(n6984), .B(n6983), .Z(n6985) );
  NANDN U7627 ( .A(rst), .B(n6985), .Z(n6986) );
  NAND U7628 ( .A(n6987), .B(n6986), .Z(n1924) );
  NAND U7629 ( .A(c[388]), .B(rst), .Z(n6992) );
  XOR U7630 ( .A(n6989), .B(n6988), .Z(n6990) );
  NANDN U7631 ( .A(rst), .B(n6990), .Z(n6991) );
  NAND U7632 ( .A(n6992), .B(n6991), .Z(n1925) );
  NAND U7633 ( .A(c[389]), .B(rst), .Z(n6997) );
  XNOR U7634 ( .A(n6994), .B(n6993), .Z(n6995) );
  NANDN U7635 ( .A(rst), .B(n6995), .Z(n6996) );
  NAND U7636 ( .A(n6997), .B(n6996), .Z(n1926) );
  NAND U7637 ( .A(c[390]), .B(rst), .Z(n7002) );
  XOR U7638 ( .A(n6999), .B(n6998), .Z(n7000) );
  NANDN U7639 ( .A(rst), .B(n7000), .Z(n7001) );
  NAND U7640 ( .A(n7002), .B(n7001), .Z(n1927) );
  NAND U7641 ( .A(c[391]), .B(rst), .Z(n7007) );
  XNOR U7642 ( .A(n7004), .B(n7003), .Z(n7005) );
  NANDN U7643 ( .A(rst), .B(n7005), .Z(n7006) );
  NAND U7644 ( .A(n7007), .B(n7006), .Z(n1928) );
  NAND U7645 ( .A(c[392]), .B(rst), .Z(n7012) );
  XOR U7646 ( .A(n7009), .B(n7008), .Z(n7010) );
  NANDN U7647 ( .A(rst), .B(n7010), .Z(n7011) );
  NAND U7648 ( .A(n7012), .B(n7011), .Z(n1929) );
  NAND U7649 ( .A(c[393]), .B(rst), .Z(n7017) );
  XNOR U7650 ( .A(n7014), .B(n7013), .Z(n7015) );
  NANDN U7651 ( .A(rst), .B(n7015), .Z(n7016) );
  NAND U7652 ( .A(n7017), .B(n7016), .Z(n1930) );
  NAND U7653 ( .A(c[394]), .B(rst), .Z(n7022) );
  XOR U7654 ( .A(n7019), .B(n7018), .Z(n7020) );
  NANDN U7655 ( .A(rst), .B(n7020), .Z(n7021) );
  NAND U7656 ( .A(n7022), .B(n7021), .Z(n1931) );
  NAND U7657 ( .A(c[395]), .B(rst), .Z(n7027) );
  XNOR U7658 ( .A(n7024), .B(n7023), .Z(n7025) );
  NANDN U7659 ( .A(rst), .B(n7025), .Z(n7026) );
  NAND U7660 ( .A(n7027), .B(n7026), .Z(n1932) );
  NAND U7661 ( .A(c[396]), .B(rst), .Z(n7032) );
  XOR U7662 ( .A(n7029), .B(n7028), .Z(n7030) );
  NANDN U7663 ( .A(rst), .B(n7030), .Z(n7031) );
  NAND U7664 ( .A(n7032), .B(n7031), .Z(n1933) );
  NAND U7665 ( .A(c[397]), .B(rst), .Z(n7037) );
  XNOR U7666 ( .A(n7034), .B(n7033), .Z(n7035) );
  NANDN U7667 ( .A(rst), .B(n7035), .Z(n7036) );
  NAND U7668 ( .A(n7037), .B(n7036), .Z(n1934) );
  NAND U7669 ( .A(c[398]), .B(rst), .Z(n7042) );
  XOR U7670 ( .A(n7039), .B(n7038), .Z(n7040) );
  NANDN U7671 ( .A(rst), .B(n7040), .Z(n7041) );
  NAND U7672 ( .A(n7042), .B(n7041), .Z(n1935) );
  NAND U7673 ( .A(c[399]), .B(rst), .Z(n7047) );
  XNOR U7674 ( .A(n7044), .B(n7043), .Z(n7045) );
  NANDN U7675 ( .A(rst), .B(n7045), .Z(n7046) );
  NAND U7676 ( .A(n7047), .B(n7046), .Z(n1936) );
  NAND U7677 ( .A(c[400]), .B(rst), .Z(n7052) );
  XOR U7678 ( .A(n7049), .B(n7048), .Z(n7050) );
  NANDN U7679 ( .A(rst), .B(n7050), .Z(n7051) );
  NAND U7680 ( .A(n7052), .B(n7051), .Z(n1937) );
  NAND U7681 ( .A(c[401]), .B(rst), .Z(n7057) );
  XNOR U7682 ( .A(n7054), .B(n7053), .Z(n7055) );
  NANDN U7683 ( .A(rst), .B(n7055), .Z(n7056) );
  NAND U7684 ( .A(n7057), .B(n7056), .Z(n1938) );
  NAND U7685 ( .A(c[402]), .B(rst), .Z(n7062) );
  XOR U7686 ( .A(n7059), .B(n7058), .Z(n7060) );
  NANDN U7687 ( .A(rst), .B(n7060), .Z(n7061) );
  NAND U7688 ( .A(n7062), .B(n7061), .Z(n1939) );
  NAND U7689 ( .A(c[403]), .B(rst), .Z(n7067) );
  XNOR U7690 ( .A(n7064), .B(n7063), .Z(n7065) );
  NANDN U7691 ( .A(rst), .B(n7065), .Z(n7066) );
  NAND U7692 ( .A(n7067), .B(n7066), .Z(n1940) );
  NAND U7693 ( .A(c[404]), .B(rst), .Z(n7072) );
  XOR U7694 ( .A(n7069), .B(n7068), .Z(n7070) );
  NANDN U7695 ( .A(rst), .B(n7070), .Z(n7071) );
  NAND U7696 ( .A(n7072), .B(n7071), .Z(n1941) );
  NAND U7697 ( .A(c[405]), .B(rst), .Z(n7077) );
  XNOR U7698 ( .A(n7074), .B(n7073), .Z(n7075) );
  NANDN U7699 ( .A(rst), .B(n7075), .Z(n7076) );
  NAND U7700 ( .A(n7077), .B(n7076), .Z(n1942) );
  NAND U7701 ( .A(c[406]), .B(rst), .Z(n7082) );
  XOR U7702 ( .A(n7079), .B(n7078), .Z(n7080) );
  NANDN U7703 ( .A(rst), .B(n7080), .Z(n7081) );
  NAND U7704 ( .A(n7082), .B(n7081), .Z(n1943) );
  NAND U7705 ( .A(c[407]), .B(rst), .Z(n7087) );
  XNOR U7706 ( .A(n7084), .B(n7083), .Z(n7085) );
  NANDN U7707 ( .A(rst), .B(n7085), .Z(n7086) );
  NAND U7708 ( .A(n7087), .B(n7086), .Z(n1944) );
  NAND U7709 ( .A(c[408]), .B(rst), .Z(n7092) );
  XNOR U7710 ( .A(n7089), .B(n7088), .Z(n7090) );
  NANDN U7711 ( .A(rst), .B(n7090), .Z(n7091) );
  NAND U7712 ( .A(n7092), .B(n7091), .Z(n1945) );
  NAND U7713 ( .A(c[409]), .B(rst), .Z(n7097) );
  XNOR U7714 ( .A(n7094), .B(n7093), .Z(n7095) );
  NANDN U7715 ( .A(rst), .B(n7095), .Z(n7096) );
  NAND U7716 ( .A(n7097), .B(n7096), .Z(n1946) );
  NAND U7717 ( .A(c[410]), .B(rst), .Z(n7102) );
  XNOR U7718 ( .A(n7099), .B(n7098), .Z(n7100) );
  NANDN U7719 ( .A(rst), .B(n7100), .Z(n7101) );
  NAND U7720 ( .A(n7102), .B(n7101), .Z(n1947) );
  NAND U7721 ( .A(c[411]), .B(rst), .Z(n7107) );
  XOR U7722 ( .A(n7104), .B(n7103), .Z(n7105) );
  NANDN U7723 ( .A(rst), .B(n7105), .Z(n7106) );
  NAND U7724 ( .A(n7107), .B(n7106), .Z(n1948) );
  NAND U7725 ( .A(c[412]), .B(rst), .Z(n7112) );
  XNOR U7726 ( .A(n7109), .B(n7108), .Z(n7110) );
  NANDN U7727 ( .A(rst), .B(n7110), .Z(n7111) );
  NAND U7728 ( .A(n7112), .B(n7111), .Z(n1949) );
  NAND U7729 ( .A(c[413]), .B(rst), .Z(n7117) );
  XNOR U7730 ( .A(n7114), .B(n7113), .Z(n7115) );
  NANDN U7731 ( .A(rst), .B(n7115), .Z(n7116) );
  NAND U7732 ( .A(n7117), .B(n7116), .Z(n1950) );
  NAND U7733 ( .A(c[414]), .B(rst), .Z(n7122) );
  XNOR U7734 ( .A(n7119), .B(n7118), .Z(n7120) );
  NANDN U7735 ( .A(rst), .B(n7120), .Z(n7121) );
  NAND U7736 ( .A(n7122), .B(n7121), .Z(n1951) );
  NAND U7737 ( .A(c[415]), .B(rst), .Z(n7127) );
  XNOR U7738 ( .A(n7124), .B(n7123), .Z(n7125) );
  NANDN U7739 ( .A(rst), .B(n7125), .Z(n7126) );
  NAND U7740 ( .A(n7127), .B(n7126), .Z(n1952) );
  NAND U7741 ( .A(c[416]), .B(rst), .Z(n7132) );
  XOR U7742 ( .A(n7129), .B(n7128), .Z(n7130) );
  NANDN U7743 ( .A(rst), .B(n7130), .Z(n7131) );
  NAND U7744 ( .A(n7132), .B(n7131), .Z(n1953) );
  NAND U7745 ( .A(c[417]), .B(rst), .Z(n7137) );
  XNOR U7746 ( .A(n7134), .B(n7133), .Z(n7135) );
  NANDN U7747 ( .A(rst), .B(n7135), .Z(n7136) );
  NAND U7748 ( .A(n7137), .B(n7136), .Z(n1954) );
  NAND U7749 ( .A(c[418]), .B(rst), .Z(n7142) );
  XOR U7750 ( .A(n7139), .B(n7138), .Z(n7140) );
  NANDN U7751 ( .A(rst), .B(n7140), .Z(n7141) );
  NAND U7752 ( .A(n7142), .B(n7141), .Z(n1955) );
  NAND U7753 ( .A(c[419]), .B(rst), .Z(n7147) );
  XNOR U7754 ( .A(n7144), .B(n7143), .Z(n7145) );
  NANDN U7755 ( .A(rst), .B(n7145), .Z(n7146) );
  NAND U7756 ( .A(n7147), .B(n7146), .Z(n1956) );
  NAND U7757 ( .A(c[420]), .B(rst), .Z(n7152) );
  XOR U7758 ( .A(n7149), .B(n7148), .Z(n7150) );
  NANDN U7759 ( .A(rst), .B(n7150), .Z(n7151) );
  NAND U7760 ( .A(n7152), .B(n7151), .Z(n1957) );
  NAND U7761 ( .A(c[421]), .B(rst), .Z(n7157) );
  XNOR U7762 ( .A(n7154), .B(n7153), .Z(n7155) );
  NANDN U7763 ( .A(rst), .B(n7155), .Z(n7156) );
  NAND U7764 ( .A(n7157), .B(n7156), .Z(n1958) );
  NAND U7765 ( .A(c[422]), .B(rst), .Z(n7162) );
  XNOR U7766 ( .A(n7159), .B(n7158), .Z(n7160) );
  NANDN U7767 ( .A(rst), .B(n7160), .Z(n7161) );
  NAND U7768 ( .A(n7162), .B(n7161), .Z(n1959) );
  NAND U7769 ( .A(c[423]), .B(rst), .Z(n7167) );
  XNOR U7770 ( .A(n7164), .B(n7163), .Z(n7165) );
  NANDN U7771 ( .A(rst), .B(n7165), .Z(n7166) );
  NAND U7772 ( .A(n7167), .B(n7166), .Z(n1960) );
  NAND U7773 ( .A(c[424]), .B(rst), .Z(n7172) );
  XNOR U7774 ( .A(n7169), .B(n7168), .Z(n7170) );
  NANDN U7775 ( .A(rst), .B(n7170), .Z(n7171) );
  NAND U7776 ( .A(n7172), .B(n7171), .Z(n1961) );
  NAND U7777 ( .A(c[425]), .B(rst), .Z(n7177) );
  XOR U7778 ( .A(n7174), .B(n7173), .Z(n7175) );
  NANDN U7779 ( .A(rst), .B(n7175), .Z(n7176) );
  NAND U7780 ( .A(n7177), .B(n7176), .Z(n1962) );
  NAND U7781 ( .A(c[426]), .B(rst), .Z(n7182) );
  XNOR U7782 ( .A(n7179), .B(n7178), .Z(n7180) );
  NANDN U7783 ( .A(rst), .B(n7180), .Z(n7181) );
  NAND U7784 ( .A(n7182), .B(n7181), .Z(n1963) );
  NAND U7785 ( .A(c[427]), .B(rst), .Z(n7187) );
  XOR U7786 ( .A(n7184), .B(n7183), .Z(n7185) );
  NANDN U7787 ( .A(rst), .B(n7185), .Z(n7186) );
  NAND U7788 ( .A(n7187), .B(n7186), .Z(n1964) );
  NAND U7789 ( .A(c[428]), .B(rst), .Z(n7192) );
  XNOR U7790 ( .A(n7189), .B(n7188), .Z(n7190) );
  NANDN U7791 ( .A(rst), .B(n7190), .Z(n7191) );
  NAND U7792 ( .A(n7192), .B(n7191), .Z(n1965) );
  NAND U7793 ( .A(c[429]), .B(rst), .Z(n7197) );
  XOR U7794 ( .A(n7194), .B(n7193), .Z(n7195) );
  NANDN U7795 ( .A(rst), .B(n7195), .Z(n7196) );
  NAND U7796 ( .A(n7197), .B(n7196), .Z(n1966) );
  NAND U7797 ( .A(c[430]), .B(rst), .Z(n7202) );
  XNOR U7798 ( .A(n7199), .B(n7198), .Z(n7200) );
  NANDN U7799 ( .A(rst), .B(n7200), .Z(n7201) );
  NAND U7800 ( .A(n7202), .B(n7201), .Z(n1967) );
  NAND U7801 ( .A(c[431]), .B(rst), .Z(n7207) );
  XOR U7802 ( .A(n7204), .B(n7203), .Z(n7205) );
  NANDN U7803 ( .A(rst), .B(n7205), .Z(n7206) );
  NAND U7804 ( .A(n7207), .B(n7206), .Z(n1968) );
  NAND U7805 ( .A(c[432]), .B(rst), .Z(n7212) );
  XNOR U7806 ( .A(n7209), .B(n7208), .Z(n7210) );
  NANDN U7807 ( .A(rst), .B(n7210), .Z(n7211) );
  NAND U7808 ( .A(n7212), .B(n7211), .Z(n1969) );
  NAND U7809 ( .A(c[433]), .B(rst), .Z(n7217) );
  XOR U7810 ( .A(n7214), .B(n7213), .Z(n7215) );
  NANDN U7811 ( .A(rst), .B(n7215), .Z(n7216) );
  NAND U7812 ( .A(n7217), .B(n7216), .Z(n1970) );
  NAND U7813 ( .A(c[434]), .B(rst), .Z(n7222) );
  XNOR U7814 ( .A(n7219), .B(n7218), .Z(n7220) );
  NANDN U7815 ( .A(rst), .B(n7220), .Z(n7221) );
  NAND U7816 ( .A(n7222), .B(n7221), .Z(n1971) );
  NAND U7817 ( .A(c[435]), .B(rst), .Z(n7227) );
  XOR U7818 ( .A(n7224), .B(n7223), .Z(n7225) );
  NANDN U7819 ( .A(rst), .B(n7225), .Z(n7226) );
  NAND U7820 ( .A(n7227), .B(n7226), .Z(n1972) );
  NAND U7821 ( .A(c[436]), .B(rst), .Z(n7232) );
  XNOR U7822 ( .A(n7229), .B(n7228), .Z(n7230) );
  NANDN U7823 ( .A(rst), .B(n7230), .Z(n7231) );
  NAND U7824 ( .A(n7232), .B(n7231), .Z(n1973) );
  NAND U7825 ( .A(c[437]), .B(rst), .Z(n7237) );
  XOR U7826 ( .A(n7234), .B(n7233), .Z(n7235) );
  NANDN U7827 ( .A(rst), .B(n7235), .Z(n7236) );
  NAND U7828 ( .A(n7237), .B(n7236), .Z(n1974) );
  NAND U7829 ( .A(c[438]), .B(rst), .Z(n7242) );
  XNOR U7830 ( .A(n7239), .B(n7238), .Z(n7240) );
  NANDN U7831 ( .A(rst), .B(n7240), .Z(n7241) );
  NAND U7832 ( .A(n7242), .B(n7241), .Z(n1975) );
  NAND U7833 ( .A(c[439]), .B(rst), .Z(n7247) );
  XOR U7834 ( .A(n7244), .B(n7243), .Z(n7245) );
  NANDN U7835 ( .A(rst), .B(n7245), .Z(n7246) );
  NAND U7836 ( .A(n7247), .B(n7246), .Z(n1976) );
  NAND U7837 ( .A(c[440]), .B(rst), .Z(n7252) );
  XNOR U7838 ( .A(n7249), .B(n7248), .Z(n7250) );
  NANDN U7839 ( .A(rst), .B(n7250), .Z(n7251) );
  NAND U7840 ( .A(n7252), .B(n7251), .Z(n1977) );
  NAND U7841 ( .A(c[441]), .B(rst), .Z(n7257) );
  XNOR U7842 ( .A(n7254), .B(n7253), .Z(n7255) );
  NANDN U7843 ( .A(rst), .B(n7255), .Z(n7256) );
  NAND U7844 ( .A(n7257), .B(n7256), .Z(n1978) );
  NAND U7845 ( .A(c[442]), .B(rst), .Z(n7262) );
  XNOR U7846 ( .A(n7259), .B(n7258), .Z(n7260) );
  NANDN U7847 ( .A(rst), .B(n7260), .Z(n7261) );
  NAND U7848 ( .A(n7262), .B(n7261), .Z(n1979) );
  NAND U7849 ( .A(c[443]), .B(rst), .Z(n7267) );
  XNOR U7850 ( .A(n7264), .B(n7263), .Z(n7265) );
  NANDN U7851 ( .A(rst), .B(n7265), .Z(n7266) );
  NAND U7852 ( .A(n7267), .B(n7266), .Z(n1980) );
  NAND U7853 ( .A(c[444]), .B(rst), .Z(n7272) );
  XOR U7854 ( .A(n7269), .B(n7268), .Z(n7270) );
  NANDN U7855 ( .A(rst), .B(n7270), .Z(n7271) );
  NAND U7856 ( .A(n7272), .B(n7271), .Z(n1981) );
  NAND U7857 ( .A(c[445]), .B(rst), .Z(n7277) );
  XNOR U7858 ( .A(n7274), .B(n7273), .Z(n7275) );
  NANDN U7859 ( .A(rst), .B(n7275), .Z(n7276) );
  NAND U7860 ( .A(n7277), .B(n7276), .Z(n1982) );
  NAND U7861 ( .A(c[446]), .B(rst), .Z(n7282) );
  XNOR U7862 ( .A(n7279), .B(n7278), .Z(n7280) );
  NANDN U7863 ( .A(rst), .B(n7280), .Z(n7281) );
  NAND U7864 ( .A(n7282), .B(n7281), .Z(n1983) );
  NAND U7865 ( .A(c[447]), .B(rst), .Z(n7287) );
  XNOR U7866 ( .A(n7284), .B(n7283), .Z(n7285) );
  NANDN U7867 ( .A(rst), .B(n7285), .Z(n7286) );
  NAND U7868 ( .A(n7287), .B(n7286), .Z(n1984) );
  NAND U7869 ( .A(c[448]), .B(rst), .Z(n7292) );
  XNOR U7870 ( .A(n7289), .B(n7288), .Z(n7290) );
  NANDN U7871 ( .A(rst), .B(n7290), .Z(n7291) );
  NAND U7872 ( .A(n7292), .B(n7291), .Z(n1985) );
  NAND U7873 ( .A(c[449]), .B(rst), .Z(n7297) );
  XOR U7874 ( .A(n7294), .B(n7293), .Z(n7295) );
  NANDN U7875 ( .A(rst), .B(n7295), .Z(n7296) );
  NAND U7876 ( .A(n7297), .B(n7296), .Z(n1986) );
  NAND U7877 ( .A(c[450]), .B(rst), .Z(n7302) );
  XNOR U7878 ( .A(n7299), .B(n7298), .Z(n7300) );
  NANDN U7879 ( .A(rst), .B(n7300), .Z(n7301) );
  NAND U7880 ( .A(n7302), .B(n7301), .Z(n1987) );
  NAND U7881 ( .A(c[451]), .B(rst), .Z(n7307) );
  XOR U7882 ( .A(n7304), .B(n7303), .Z(n7305) );
  NANDN U7883 ( .A(rst), .B(n7305), .Z(n7306) );
  NAND U7884 ( .A(n7307), .B(n7306), .Z(n1988) );
  NAND U7885 ( .A(c[452]), .B(rst), .Z(n7312) );
  XNOR U7886 ( .A(n7309), .B(n7308), .Z(n7310) );
  NANDN U7887 ( .A(rst), .B(n7310), .Z(n7311) );
  NAND U7888 ( .A(n7312), .B(n7311), .Z(n1989) );
  NAND U7889 ( .A(c[453]), .B(rst), .Z(n7317) );
  XOR U7890 ( .A(n7314), .B(n7313), .Z(n7315) );
  NANDN U7891 ( .A(rst), .B(n7315), .Z(n7316) );
  NAND U7892 ( .A(n7317), .B(n7316), .Z(n1990) );
  NAND U7893 ( .A(c[454]), .B(rst), .Z(n7322) );
  XNOR U7894 ( .A(n7319), .B(n7318), .Z(n7320) );
  NANDN U7895 ( .A(rst), .B(n7320), .Z(n7321) );
  NAND U7896 ( .A(n7322), .B(n7321), .Z(n1991) );
  NAND U7897 ( .A(c[455]), .B(rst), .Z(n7327) );
  XOR U7898 ( .A(n7324), .B(n7323), .Z(n7325) );
  NANDN U7899 ( .A(rst), .B(n7325), .Z(n7326) );
  NAND U7900 ( .A(n7327), .B(n7326), .Z(n1992) );
  NAND U7901 ( .A(c[456]), .B(rst), .Z(n7332) );
  XNOR U7902 ( .A(n7329), .B(n7328), .Z(n7330) );
  NANDN U7903 ( .A(rst), .B(n7330), .Z(n7331) );
  NAND U7904 ( .A(n7332), .B(n7331), .Z(n1993) );
  NAND U7905 ( .A(c[457]), .B(rst), .Z(n7337) );
  XNOR U7906 ( .A(n7334), .B(n7333), .Z(n7335) );
  NANDN U7907 ( .A(rst), .B(n7335), .Z(n7336) );
  NAND U7908 ( .A(n7337), .B(n7336), .Z(n1994) );
  NAND U7909 ( .A(c[458]), .B(rst), .Z(n7342) );
  XNOR U7910 ( .A(n7339), .B(n7338), .Z(n7340) );
  NANDN U7911 ( .A(rst), .B(n7340), .Z(n7341) );
  NAND U7912 ( .A(n7342), .B(n7341), .Z(n1995) );
  NAND U7913 ( .A(c[459]), .B(rst), .Z(n7347) );
  XNOR U7914 ( .A(n7344), .B(n7343), .Z(n7345) );
  NANDN U7915 ( .A(rst), .B(n7345), .Z(n7346) );
  NAND U7916 ( .A(n7347), .B(n7346), .Z(n1996) );
  NAND U7917 ( .A(c[460]), .B(rst), .Z(n7352) );
  XOR U7918 ( .A(n7349), .B(n7348), .Z(n7350) );
  NANDN U7919 ( .A(rst), .B(n7350), .Z(n7351) );
  NAND U7920 ( .A(n7352), .B(n7351), .Z(n1997) );
  NAND U7921 ( .A(c[461]), .B(rst), .Z(n7357) );
  XNOR U7922 ( .A(n7354), .B(n7353), .Z(n7355) );
  NANDN U7923 ( .A(rst), .B(n7355), .Z(n7356) );
  NAND U7924 ( .A(n7357), .B(n7356), .Z(n1998) );
  NAND U7925 ( .A(c[462]), .B(rst), .Z(n7362) );
  XOR U7926 ( .A(n7359), .B(n7358), .Z(n7360) );
  NANDN U7927 ( .A(rst), .B(n7360), .Z(n7361) );
  NAND U7928 ( .A(n7362), .B(n7361), .Z(n1999) );
  NAND U7929 ( .A(c[463]), .B(rst), .Z(n7367) );
  XNOR U7930 ( .A(n7364), .B(n7363), .Z(n7365) );
  NANDN U7931 ( .A(rst), .B(n7365), .Z(n7366) );
  NAND U7932 ( .A(n7367), .B(n7366), .Z(n2000) );
  NAND U7933 ( .A(c[464]), .B(rst), .Z(n7372) );
  XOR U7934 ( .A(n7369), .B(n7368), .Z(n7370) );
  NANDN U7935 ( .A(rst), .B(n7370), .Z(n7371) );
  NAND U7936 ( .A(n7372), .B(n7371), .Z(n2001) );
  NAND U7937 ( .A(c[465]), .B(rst), .Z(n7377) );
  XNOR U7938 ( .A(n7374), .B(n7373), .Z(n7375) );
  NANDN U7939 ( .A(rst), .B(n7375), .Z(n7376) );
  NAND U7940 ( .A(n7377), .B(n7376), .Z(n2002) );
  NAND U7941 ( .A(c[466]), .B(rst), .Z(n7382) );
  XOR U7942 ( .A(n7379), .B(n7378), .Z(n7380) );
  NANDN U7943 ( .A(rst), .B(n7380), .Z(n7381) );
  NAND U7944 ( .A(n7382), .B(n7381), .Z(n2003) );
  NAND U7945 ( .A(c[467]), .B(rst), .Z(n7387) );
  XNOR U7946 ( .A(n7384), .B(n7383), .Z(n7385) );
  NANDN U7947 ( .A(rst), .B(n7385), .Z(n7386) );
  NAND U7948 ( .A(n7387), .B(n7386), .Z(n2004) );
  NAND U7949 ( .A(c[468]), .B(rst), .Z(n7392) );
  XOR U7950 ( .A(n7389), .B(n7388), .Z(n7390) );
  NANDN U7951 ( .A(rst), .B(n7390), .Z(n7391) );
  NAND U7952 ( .A(n7392), .B(n7391), .Z(n2005) );
  NAND U7953 ( .A(c[469]), .B(rst), .Z(n7397) );
  XNOR U7954 ( .A(n7394), .B(n7393), .Z(n7395) );
  NANDN U7955 ( .A(rst), .B(n7395), .Z(n7396) );
  NAND U7956 ( .A(n7397), .B(n7396), .Z(n2006) );
  NAND U7957 ( .A(c[470]), .B(rst), .Z(n7402) );
  XOR U7958 ( .A(n7399), .B(n7398), .Z(n7400) );
  NANDN U7959 ( .A(rst), .B(n7400), .Z(n7401) );
  NAND U7960 ( .A(n7402), .B(n7401), .Z(n2007) );
  NAND U7961 ( .A(c[471]), .B(rst), .Z(n7407) );
  XNOR U7962 ( .A(n7404), .B(n7403), .Z(n7405) );
  NANDN U7963 ( .A(rst), .B(n7405), .Z(n7406) );
  NAND U7964 ( .A(n7407), .B(n7406), .Z(n2008) );
  NAND U7965 ( .A(c[472]), .B(rst), .Z(n7412) );
  XOR U7966 ( .A(n7409), .B(n7408), .Z(n7410) );
  NANDN U7967 ( .A(rst), .B(n7410), .Z(n7411) );
  NAND U7968 ( .A(n7412), .B(n7411), .Z(n2009) );
  NAND U7969 ( .A(c[473]), .B(rst), .Z(n7417) );
  XNOR U7970 ( .A(n7414), .B(n7413), .Z(n7415) );
  NANDN U7971 ( .A(rst), .B(n7415), .Z(n7416) );
  NAND U7972 ( .A(n7417), .B(n7416), .Z(n2010) );
  NAND U7973 ( .A(c[474]), .B(rst), .Z(n7422) );
  XNOR U7974 ( .A(n7419), .B(n7418), .Z(n7420) );
  NANDN U7975 ( .A(rst), .B(n7420), .Z(n7421) );
  NAND U7976 ( .A(n7422), .B(n7421), .Z(n2011) );
  NAND U7977 ( .A(c[475]), .B(rst), .Z(n7427) );
  XNOR U7978 ( .A(n7424), .B(n7423), .Z(n7425) );
  NANDN U7979 ( .A(rst), .B(n7425), .Z(n7426) );
  NAND U7980 ( .A(n7427), .B(n7426), .Z(n2012) );
  NAND U7981 ( .A(c[476]), .B(rst), .Z(n7432) );
  XNOR U7982 ( .A(n7429), .B(n7428), .Z(n7430) );
  NANDN U7983 ( .A(rst), .B(n7430), .Z(n7431) );
  NAND U7984 ( .A(n7432), .B(n7431), .Z(n2013) );
  NAND U7985 ( .A(c[477]), .B(rst), .Z(n7437) );
  XOR U7986 ( .A(n7434), .B(n7433), .Z(n7435) );
  NANDN U7987 ( .A(rst), .B(n7435), .Z(n7436) );
  NAND U7988 ( .A(n7437), .B(n7436), .Z(n2014) );
  NAND U7989 ( .A(c[478]), .B(rst), .Z(n7442) );
  XNOR U7990 ( .A(n7439), .B(n7438), .Z(n7440) );
  NANDN U7991 ( .A(rst), .B(n7440), .Z(n7441) );
  NAND U7992 ( .A(n7442), .B(n7441), .Z(n2015) );
  NAND U7993 ( .A(c[479]), .B(rst), .Z(n7447) );
  XOR U7994 ( .A(n7444), .B(n7443), .Z(n7445) );
  NANDN U7995 ( .A(rst), .B(n7445), .Z(n7446) );
  NAND U7996 ( .A(n7447), .B(n7446), .Z(n2016) );
  NAND U7997 ( .A(c[480]), .B(rst), .Z(n7452) );
  XNOR U7998 ( .A(n7449), .B(n7448), .Z(n7450) );
  NANDN U7999 ( .A(rst), .B(n7450), .Z(n7451) );
  NAND U8000 ( .A(n7452), .B(n7451), .Z(n2017) );
  NAND U8001 ( .A(c[481]), .B(rst), .Z(n7457) );
  XOR U8002 ( .A(n7454), .B(n7453), .Z(n7455) );
  NANDN U8003 ( .A(rst), .B(n7455), .Z(n7456) );
  NAND U8004 ( .A(n7457), .B(n7456), .Z(n2018) );
  NAND U8005 ( .A(c[482]), .B(rst), .Z(n7462) );
  XNOR U8006 ( .A(n7459), .B(n7458), .Z(n7460) );
  NANDN U8007 ( .A(rst), .B(n7460), .Z(n7461) );
  NAND U8008 ( .A(n7462), .B(n7461), .Z(n2019) );
  NAND U8009 ( .A(c[483]), .B(rst), .Z(n7467) );
  XOR U8010 ( .A(n7464), .B(n7463), .Z(n7465) );
  NANDN U8011 ( .A(rst), .B(n7465), .Z(n7466) );
  NAND U8012 ( .A(n7467), .B(n7466), .Z(n2020) );
  NAND U8013 ( .A(c[484]), .B(rst), .Z(n7472) );
  XNOR U8014 ( .A(n7469), .B(n7468), .Z(n7470) );
  NANDN U8015 ( .A(rst), .B(n7470), .Z(n7471) );
  NAND U8016 ( .A(n7472), .B(n7471), .Z(n2021) );
  NAND U8017 ( .A(c[485]), .B(rst), .Z(n7477) );
  XOR U8018 ( .A(n7474), .B(n7473), .Z(n7475) );
  NANDN U8019 ( .A(rst), .B(n7475), .Z(n7476) );
  NAND U8020 ( .A(n7477), .B(n7476), .Z(n2022) );
  NAND U8021 ( .A(c[486]), .B(rst), .Z(n7482) );
  XNOR U8022 ( .A(n7479), .B(n7478), .Z(n7480) );
  NANDN U8023 ( .A(rst), .B(n7480), .Z(n7481) );
  NAND U8024 ( .A(n7482), .B(n7481), .Z(n2023) );
  NAND U8025 ( .A(c[487]), .B(rst), .Z(n7487) );
  XOR U8026 ( .A(n7484), .B(n7483), .Z(n7485) );
  NANDN U8027 ( .A(rst), .B(n7485), .Z(n7486) );
  NAND U8028 ( .A(n7487), .B(n7486), .Z(n2024) );
  NAND U8029 ( .A(c[488]), .B(rst), .Z(n7492) );
  XNOR U8030 ( .A(n7489), .B(n7488), .Z(n7490) );
  NANDN U8031 ( .A(rst), .B(n7490), .Z(n7491) );
  NAND U8032 ( .A(n7492), .B(n7491), .Z(n2025) );
  NAND U8033 ( .A(c[489]), .B(rst), .Z(n7497) );
  XOR U8034 ( .A(n7494), .B(n7493), .Z(n7495) );
  NANDN U8035 ( .A(rst), .B(n7495), .Z(n7496) );
  NAND U8036 ( .A(n7497), .B(n7496), .Z(n2026) );
  NAND U8037 ( .A(c[490]), .B(rst), .Z(n7502) );
  XNOR U8038 ( .A(n7499), .B(n7498), .Z(n7500) );
  NANDN U8039 ( .A(rst), .B(n7500), .Z(n7501) );
  NAND U8040 ( .A(n7502), .B(n7501), .Z(n2027) );
  NAND U8041 ( .A(c[491]), .B(rst), .Z(n7507) );
  XOR U8042 ( .A(n7504), .B(n7503), .Z(n7505) );
  NANDN U8043 ( .A(rst), .B(n7505), .Z(n7506) );
  NAND U8044 ( .A(n7507), .B(n7506), .Z(n2028) );
  NAND U8045 ( .A(c[492]), .B(rst), .Z(n7512) );
  XNOR U8046 ( .A(n7509), .B(n7508), .Z(n7510) );
  NANDN U8047 ( .A(rst), .B(n7510), .Z(n7511) );
  NAND U8048 ( .A(n7512), .B(n7511), .Z(n2029) );
  NAND U8049 ( .A(c[493]), .B(rst), .Z(n7517) );
  XNOR U8050 ( .A(n7514), .B(n7513), .Z(n7515) );
  NANDN U8051 ( .A(rst), .B(n7515), .Z(n7516) );
  NAND U8052 ( .A(n7517), .B(n7516), .Z(n2030) );
  NAND U8053 ( .A(c[494]), .B(rst), .Z(n7522) );
  XNOR U8054 ( .A(n7519), .B(n7518), .Z(n7520) );
  NANDN U8055 ( .A(rst), .B(n7520), .Z(n7521) );
  NAND U8056 ( .A(n7522), .B(n7521), .Z(n2031) );
  NAND U8057 ( .A(c[495]), .B(rst), .Z(n7527) );
  XNOR U8058 ( .A(n7524), .B(n7523), .Z(n7525) );
  NANDN U8059 ( .A(rst), .B(n7525), .Z(n7526) );
  NAND U8060 ( .A(n7527), .B(n7526), .Z(n2032) );
  NAND U8061 ( .A(c[496]), .B(rst), .Z(n7532) );
  XOR U8062 ( .A(n7529), .B(n7528), .Z(n7530) );
  NANDN U8063 ( .A(rst), .B(n7530), .Z(n7531) );
  NAND U8064 ( .A(n7532), .B(n7531), .Z(n2033) );
  NAND U8065 ( .A(c[497]), .B(rst), .Z(n7537) );
  XNOR U8066 ( .A(n7534), .B(n7533), .Z(n7535) );
  NANDN U8067 ( .A(rst), .B(n7535), .Z(n7536) );
  NAND U8068 ( .A(n7537), .B(n7536), .Z(n2034) );
  NAND U8069 ( .A(c[498]), .B(rst), .Z(n7542) );
  XOR U8070 ( .A(n7539), .B(n7538), .Z(n7540) );
  NANDN U8071 ( .A(rst), .B(n7540), .Z(n7541) );
  NAND U8072 ( .A(n7542), .B(n7541), .Z(n2035) );
  NAND U8073 ( .A(c[499]), .B(rst), .Z(n7547) );
  XNOR U8074 ( .A(n7544), .B(n7543), .Z(n7545) );
  NANDN U8075 ( .A(rst), .B(n7545), .Z(n7546) );
  NAND U8076 ( .A(n7547), .B(n7546), .Z(n2036) );
  NAND U8077 ( .A(c[500]), .B(rst), .Z(n7552) );
  XOR U8078 ( .A(n7549), .B(n7548), .Z(n7550) );
  NANDN U8079 ( .A(rst), .B(n7550), .Z(n7551) );
  NAND U8080 ( .A(n7552), .B(n7551), .Z(n2037) );
  NAND U8081 ( .A(c[501]), .B(rst), .Z(n7557) );
  XNOR U8082 ( .A(n7554), .B(n7553), .Z(n7555) );
  NANDN U8083 ( .A(rst), .B(n7555), .Z(n7556) );
  NAND U8084 ( .A(n7557), .B(n7556), .Z(n2038) );
  NAND U8085 ( .A(c[502]), .B(rst), .Z(n7562) );
  XOR U8086 ( .A(n7559), .B(n7558), .Z(n7560) );
  NANDN U8087 ( .A(rst), .B(n7560), .Z(n7561) );
  NAND U8088 ( .A(n7562), .B(n7561), .Z(n2039) );
  NAND U8089 ( .A(c[503]), .B(rst), .Z(n7567) );
  XNOR U8090 ( .A(n7564), .B(n7563), .Z(n7565) );
  NANDN U8091 ( .A(rst), .B(n7565), .Z(n7566) );
  NAND U8092 ( .A(n7567), .B(n7566), .Z(n2040) );
  NAND U8093 ( .A(c[504]), .B(rst), .Z(n7572) );
  XOR U8094 ( .A(n7569), .B(n7568), .Z(n7570) );
  NANDN U8095 ( .A(rst), .B(n7570), .Z(n7571) );
  NAND U8096 ( .A(n7572), .B(n7571), .Z(n2041) );
  NAND U8097 ( .A(c[505]), .B(rst), .Z(n7577) );
  XNOR U8098 ( .A(n7574), .B(n7573), .Z(n7575) );
  NANDN U8099 ( .A(rst), .B(n7575), .Z(n7576) );
  NAND U8100 ( .A(n7577), .B(n7576), .Z(n2042) );
  NAND U8101 ( .A(c[506]), .B(rst), .Z(n7582) );
  XOR U8102 ( .A(n7579), .B(n7578), .Z(n7580) );
  NANDN U8103 ( .A(rst), .B(n7580), .Z(n7581) );
  NAND U8104 ( .A(n7582), .B(n7581), .Z(n2043) );
  NAND U8105 ( .A(c[507]), .B(rst), .Z(n7587) );
  XNOR U8106 ( .A(n7584), .B(n7583), .Z(n7585) );
  NANDN U8107 ( .A(rst), .B(n7585), .Z(n7586) );
  NAND U8108 ( .A(n7587), .B(n7586), .Z(n2044) );
  NAND U8109 ( .A(c[508]), .B(rst), .Z(n7592) );
  XOR U8110 ( .A(n7589), .B(n7588), .Z(n7590) );
  NANDN U8111 ( .A(rst), .B(n7590), .Z(n7591) );
  NAND U8112 ( .A(n7592), .B(n7591), .Z(n2045) );
  NAND U8113 ( .A(c[509]), .B(rst), .Z(n7597) );
  XNOR U8114 ( .A(n7594), .B(n7593), .Z(n7595) );
  NANDN U8115 ( .A(rst), .B(n7595), .Z(n7596) );
  NAND U8116 ( .A(n7597), .B(n7596), .Z(n2046) );
  NAND U8117 ( .A(c[510]), .B(rst), .Z(n7602) );
  XNOR U8118 ( .A(n7599), .B(n7598), .Z(n7600) );
  NANDN U8119 ( .A(rst), .B(n7600), .Z(n7601) );
  NAND U8120 ( .A(n7602), .B(n7601), .Z(n2047) );
  NAND U8121 ( .A(c[511]), .B(rst), .Z(n7607) );
  XNOR U8122 ( .A(n7604), .B(n7603), .Z(n7605) );
  NANDN U8123 ( .A(rst), .B(n7605), .Z(n7606) );
  NAND U8124 ( .A(n7607), .B(n7606), .Z(n2048) );
endmodule

