
module matrixMult_N_M_0_N3_M8 ( clk, rst, x, y, o );
  input [71:0] x;
  input [71:0] y;
  output [71:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067;

  XNOR U1 ( .A(n792), .B(n791), .Z(n773) );
  XOR U2 ( .A(n932), .B(n931), .Z(n929) );
  NAND U3 ( .A(n3020), .B(n3085), .Z(n1) );
  NANDN U4 ( .A(n3021), .B(n3022), .Z(n2) );
  AND U5 ( .A(n1), .B(n2), .Z(n3065) );
  XOR U6 ( .A(n3921), .B(n3920), .Z(n3918) );
  XOR U7 ( .A(n516), .B(n515), .Z(n503) );
  NAND U8 ( .A(n950), .B(n857), .Z(n3) );
  NANDN U9 ( .A(n858), .B(n859), .Z(n4) );
  AND U10 ( .A(n3), .B(n4), .Z(n918) );
  NANDN U11 ( .A(n1726), .B(n1725), .Z(n5) );
  NANDN U12 ( .A(n1723), .B(n1724), .Z(n6) );
  AND U13 ( .A(n5), .B(n6), .Z(n1770) );
  NAND U14 ( .A(n3838), .B(n3939), .Z(n7) );
  NANDN U15 ( .A(n3839), .B(n3840), .Z(n8) );
  AND U16 ( .A(n7), .B(n8), .Z(n3907) );
  XOR U17 ( .A(n3769), .B(n3768), .Z(n3806) );
  NAND U18 ( .A(n776), .B(n775), .Z(n9) );
  NANDN U19 ( .A(n773), .B(n774), .Z(n10) );
  AND U20 ( .A(n9), .B(n10), .Z(n841) );
  XOR U21 ( .A(n1649), .B(n1648), .Z(n1650) );
  XOR U22 ( .A(n2097), .B(n2098), .Z(n2107) );
  XOR U23 ( .A(n2082), .B(n2081), .Z(n2113) );
  XOR U24 ( .A(n2905), .B(n2904), .Z(n2943) );
  XNOR U25 ( .A(n2940), .B(n2939), .Z(n2949) );
  XOR U26 ( .A(n524), .B(n523), .Z(n521) );
  NAND U27 ( .A(n877), .B(n876), .Z(n11) );
  NANDN U28 ( .A(n878), .B(n879), .Z(n12) );
  NAND U29 ( .A(n11), .B(n12), .Z(n1041) );
  XOR U30 ( .A(n938), .B(n937), .Z(n935) );
  NAND U31 ( .A(n898), .B(n897), .Z(n13) );
  NANDN U32 ( .A(n895), .B(n896), .Z(n14) );
  AND U33 ( .A(n13), .B(n14), .Z(n925) );
  XOR U34 ( .A(n1351), .B(n1350), .Z(n1348) );
  XOR U35 ( .A(n2236), .B(n2235), .Z(n2233) );
  NANDN U36 ( .A(n2517), .B(n2518), .Z(n15) );
  NANDN U37 ( .A(n2520), .B(n2519), .Z(n16) );
  NAND U38 ( .A(n15), .B(n16), .Z(n2608) );
  AND U39 ( .A(y[66]), .B(x[45]), .Z(n17) );
  NAND U40 ( .A(n2744), .B(n2745), .Z(n18) );
  NAND U41 ( .A(n2746), .B(n2747), .Z(n19) );
  AND U42 ( .A(n18), .B(n19), .Z(n20) );
  AND U43 ( .A(y[22]), .B(x[25]), .Z(n21) );
  NAND U44 ( .A(x[46]), .B(y[65]), .Z(n22) );
  XNOR U45 ( .A(n21), .B(n22), .Z(n23) );
  AND U46 ( .A(x[47]), .B(y[64]), .Z(n24) );
  NAND U47 ( .A(y[67]), .B(x[44]), .Z(n25) );
  XNOR U48 ( .A(n24), .B(n25), .Z(n26) );
  XOR U49 ( .A(n23), .B(n26), .Z(n27) );
  XNOR U50 ( .A(n2748), .B(n20), .Z(n28) );
  XNOR U51 ( .A(n27), .B(n28), .Z(n29) );
  NANDN U52 ( .A(n2743), .B(n17), .Z(n30) );
  XNOR U53 ( .A(n29), .B(n30), .Z(n2749) );
  XOR U54 ( .A(n3075), .B(n3074), .Z(n3072) );
  XNOR U55 ( .A(n3514), .B(n3513), .Z(n3512) );
  NAND U56 ( .A(n3848), .B(n3847), .Z(n31) );
  NANDN U57 ( .A(n3849), .B(n3850), .Z(n32) );
  NAND U58 ( .A(n31), .B(n32), .Z(n4047) );
  NAND U59 ( .A(n3867), .B(n3989), .Z(n33) );
  NANDN U60 ( .A(n3868), .B(n3869), .Z(n34) );
  AND U61 ( .A(n33), .B(n34), .Z(n3919) );
  XOR U62 ( .A(n500), .B(n499), .Z(n497) );
  XOR U63 ( .A(n1062), .B(n1061), .Z(n1060) );
  NANDN U64 ( .A(n1255), .B(n1254), .Z(n35) );
  NANDN U65 ( .A(n1252), .B(n1253), .Z(n36) );
  AND U66 ( .A(n35), .B(n36), .Z(n1327) );
  XOR U67 ( .A(n1794), .B(n1793), .Z(n1767) );
  NAND U68 ( .A(n3161), .B(n2997), .Z(n37) );
  NANDN U69 ( .A(n2998), .B(n2999), .Z(n38) );
  AND U70 ( .A(n37), .B(n38), .Z(n3049) );
  XOR U71 ( .A(n4067), .B(n4066), .Z(n4064) );
  XNOR U72 ( .A(n1210), .B(n1209), .Z(n1180) );
  XOR U73 ( .A(n1194), .B(n1193), .Z(n1173) );
  XOR U74 ( .A(n3763), .B(n3762), .Z(n3807) );
  XNOR U75 ( .A(n1272), .B(n1271), .Z(n1308) );
  XNOR U76 ( .A(n1645), .B(n1644), .Z(n1654) );
  XOR U77 ( .A(n2080), .B(n2079), .Z(n2081) );
  XOR U78 ( .A(n2093), .B(n2092), .Z(n2114) );
  XNOR U79 ( .A(n2110), .B(n2109), .Z(n2068) );
  XOR U80 ( .A(n2938), .B(n2937), .Z(n2939) );
  XOR U81 ( .A(n2944), .B(n2943), .Z(n2945) );
  XOR U82 ( .A(n518), .B(n517), .Z(n515) );
  NAND U83 ( .A(n866), .B(n865), .Z(n39) );
  NANDN U84 ( .A(n867), .B(n1019), .Z(n40) );
  AND U85 ( .A(n39), .B(n40), .Z(n936) );
  XOR U86 ( .A(n926), .B(n925), .Z(n923) );
  NANDN U87 ( .A(n842), .B(n841), .Z(n41) );
  NANDN U88 ( .A(n843), .B(n844), .Z(n42) );
  NAND U89 ( .A(n41), .B(n42), .Z(n1050) );
  XOR U90 ( .A(n1683), .B(n1682), .Z(n1684) );
  XOR U91 ( .A(n1788), .B(n1787), .Z(n1785) );
  XNOR U92 ( .A(n2128), .B(n2127), .Z(n2196) );
  XNOR U93 ( .A(n2228), .B(n2227), .Z(n2226) );
  NANDN U94 ( .A(n2516), .B(n2515), .Z(n43) );
  NANDN U95 ( .A(n2513), .B(n2514), .Z(n44) );
  AND U96 ( .A(n43), .B(n44), .Z(n2609) );
  XOR U97 ( .A(n2665), .B(n2664), .Z(n2662) );
  NAND U98 ( .A(n3109), .B(n3037), .Z(n45) );
  NANDN U99 ( .A(n3038), .B(n3039), .Z(n46) );
  AND U100 ( .A(n45), .B(n46), .Z(n3054) );
  NAND U101 ( .A(n2988), .B(n2987), .Z(n47) );
  NANDN U102 ( .A(n2989), .B(n2990), .Z(n48) );
  AND U103 ( .A(n47), .B(n48), .Z(n3189) );
  XNOR U104 ( .A(n3061), .B(n3060), .Z(n3059) );
  XNOR U105 ( .A(n3472), .B(n3471), .Z(n3465) );
  XOR U106 ( .A(n3500), .B(n3499), .Z(n3497) );
  XOR U107 ( .A(n3893), .B(n3892), .Z(n3895) );
  XNOR U108 ( .A(n3927), .B(n3926), .Z(n3925) );
  NAND U109 ( .A(n3881), .B(n3974), .Z(n49) );
  NANDN U110 ( .A(n3882), .B(n3883), .Z(n50) );
  AND U111 ( .A(n49), .B(n50), .Z(n3914) );
  NANDN U112 ( .A(n477), .B(n478), .Z(n51) );
  NANDN U113 ( .A(n480), .B(n479), .Z(n52) );
  NAND U114 ( .A(n51), .B(n52), .Z(n654) );
  XOR U115 ( .A(n922), .B(n921), .Z(n919) );
  XOR U116 ( .A(n1349), .B(n1348), .Z(n1325) );
  XOR U117 ( .A(n1764), .B(n1763), .Z(n1761) );
  NANDN U118 ( .A(n2972), .B(n2971), .Z(n53) );
  NANDN U119 ( .A(n2973), .B(n2974), .Z(n54) );
  NAND U120 ( .A(n53), .B(n54), .Z(n3205) );
  XNOR U121 ( .A(n3624), .B(n3623), .Z(n3636) );
  NAND U122 ( .A(n3981), .B(n3842), .Z(n55) );
  NANDN U123 ( .A(n3843), .B(n3844), .Z(n56) );
  AND U124 ( .A(n55), .B(n56), .Z(n3908) );
  XOR U125 ( .A(n325), .B(n324), .Z(n326) );
  XOR U126 ( .A(n786), .B(n785), .Z(n774) );
  XOR U127 ( .A(n1134), .B(n1133), .Z(n1167) );
  XOR U128 ( .A(n1152), .B(n1151), .Z(n1161) );
  XOR U129 ( .A(n1180), .B(n1179), .Z(n1182) );
  XOR U130 ( .A(n1188), .B(n1187), .Z(n1174) );
  XOR U131 ( .A(n2073), .B(n2072), .Z(n2074) );
  AND U132 ( .A(x[67]), .B(y[64]), .Z(n57) );
  NAND U133 ( .A(y[67]), .B(x[64]), .Z(n58) );
  XNOR U134 ( .A(n57), .B(n58), .Z(n59) );
  XNOR U135 ( .A(n59), .B(n3733), .Z(n3744) );
  XOR U136 ( .A(n3727), .B(n3726), .Z(n3738) );
  XOR U137 ( .A(n1307), .B(n1306), .Z(n1309) );
  XOR U138 ( .A(n1313), .B(n1312), .Z(n1315) );
  XOR U139 ( .A(n2903), .B(n2902), .Z(n2904) );
  NANDN U140 ( .A(n377), .B(n378), .Z(n60) );
  NANDN U141 ( .A(n376), .B(n375), .Z(n61) );
  AND U142 ( .A(n60), .B(n61), .Z(n440) );
  AND U143 ( .A(y[50]), .B(x[21]), .Z(n62) );
  NAND U144 ( .A(n610), .B(n611), .Z(n63) );
  NAND U145 ( .A(n612), .B(n613), .Z(n64) );
  AND U146 ( .A(n63), .B(n64), .Z(n65) );
  AND U147 ( .A(x[12]), .B(y[27]), .Z(n66) );
  NAND U148 ( .A(x[7]), .B(y[0]), .Z(n67) );
  XNOR U149 ( .A(n66), .B(n67), .Z(n68) );
  AND U150 ( .A(y[53]), .B(x[18]), .Z(n69) );
  NAND U151 ( .A(x[15]), .B(y[24]), .Z(n70) );
  XNOR U152 ( .A(n69), .B(n70), .Z(n71) );
  XOR U153 ( .A(n68), .B(n71), .Z(n72) );
  XNOR U154 ( .A(n614), .B(n65), .Z(n73) );
  XNOR U155 ( .A(n72), .B(n73), .Z(n74) );
  NANDN U156 ( .A(n615), .B(n62), .Z(n75) );
  XNOR U157 ( .A(n74), .B(n75), .Z(n616) );
  XOR U158 ( .A(n852), .B(n851), .Z(n854) );
  NANDN U159 ( .A(n888), .B(n889), .Z(n76) );
  NANDN U160 ( .A(n886), .B(n887), .Z(n77) );
  AND U161 ( .A(n76), .B(n77), .Z(n1036) );
  AND U162 ( .A(y[58]), .B(x[21]), .Z(n78) );
  NAND U163 ( .A(n1016), .B(n1017), .Z(n79) );
  NAND U164 ( .A(n1018), .B(n1019), .Z(n80) );
  AND U165 ( .A(n79), .B(n80), .Z(n81) );
  AND U166 ( .A(y[61]), .B(x[18]), .Z(n82) );
  NAND U167 ( .A(x[22]), .B(y[57]), .Z(n83) );
  XNOR U168 ( .A(n82), .B(n83), .Z(n84) );
  AND U169 ( .A(x[5]), .B(y[10]), .Z(n85) );
  NAND U170 ( .A(x[15]), .B(y[32]), .Z(n86) );
  XNOR U171 ( .A(n85), .B(n86), .Z(n87) );
  XOR U172 ( .A(n84), .B(n87), .Z(n88) );
  XNOR U173 ( .A(n1020), .B(n81), .Z(n89) );
  XNOR U174 ( .A(n88), .B(n89), .Z(n90) );
  NAND U175 ( .A(y[57]), .B(x[20]), .Z(n91) );
  NAND U176 ( .A(n78), .B(n91), .Z(n92) );
  XNOR U177 ( .A(n90), .B(n92), .Z(n1021) );
  NAND U178 ( .A(n890), .B(n1001), .Z(n93) );
  NANDN U179 ( .A(n891), .B(n892), .Z(n94) );
  AND U180 ( .A(n93), .B(n94), .Z(n924) );
  NAND U181 ( .A(n1237), .B(n1235), .Z(n95) );
  XOR U182 ( .A(n1237), .B(n1235), .Z(n96) );
  NANDN U183 ( .A(n1236), .B(n96), .Z(n97) );
  NAND U184 ( .A(n95), .B(n97), .Z(n1238) );
  NANDN U185 ( .A(n1656), .B(n1657), .Z(n98) );
  NANDN U186 ( .A(n1654), .B(n1655), .Z(n99) );
  AND U187 ( .A(n98), .B(n99), .Z(n1676) );
  XOR U188 ( .A(n1796), .B(n1795), .Z(n1793) );
  XOR U189 ( .A(n2184), .B(n2183), .Z(n2185) );
  NANDN U190 ( .A(n2068), .B(n2069), .Z(n100) );
  NANDN U191 ( .A(n2071), .B(n2070), .Z(n101) );
  NAND U192 ( .A(n100), .B(n101), .Z(n2119) );
  XNOR U193 ( .A(n2222), .B(n2221), .Z(n2220) );
  NANDN U194 ( .A(n2522), .B(n2521), .Z(n102) );
  NANDN U195 ( .A(n2523), .B(n2524), .Z(n103) );
  AND U196 ( .A(n102), .B(n103), .Z(n2620) );
  XOR U197 ( .A(n2657), .B(n2656), .Z(n2654) );
  NANDN U198 ( .A(n2951), .B(n2952), .Z(n104) );
  NANDN U199 ( .A(n2949), .B(n2950), .Z(n105) );
  AND U200 ( .A(n104), .B(n105), .Z(n2971) );
  XOR U201 ( .A(n3055), .B(n3054), .Z(n3052) );
  NAND U202 ( .A(n3000), .B(n3080), .Z(n106) );
  NANDN U203 ( .A(n3001), .B(n3002), .Z(n107) );
  AND U204 ( .A(n106), .B(n107), .Z(n3073) );
  NAND U205 ( .A(n3259), .B(n3258), .Z(n108) );
  NANDN U206 ( .A(n3256), .B(n3257), .Z(n109) );
  AND U207 ( .A(n108), .B(n109), .Z(n3291) );
  XOR U208 ( .A(n3494), .B(n3493), .Z(n3491) );
  XNOR U209 ( .A(n3506), .B(n3505), .Z(n3504) );
  XOR U210 ( .A(n3899), .B(n3898), .Z(n3900) );
  NAND U211 ( .A(n3825), .B(n3824), .Z(n110) );
  XOR U212 ( .A(n3825), .B(n3824), .Z(n111) );
  NANDN U213 ( .A(n3826), .B(n111), .Z(n112) );
  NAND U214 ( .A(n110), .B(n112), .Z(n3827) );
  NANDN U215 ( .A(n3865), .B(n3866), .Z(n113) );
  NANDN U216 ( .A(n3863), .B(n3864), .Z(n114) );
  AND U217 ( .A(n113), .B(n114), .Z(n4041) );
  NAND U218 ( .A(n3834), .B(n3833), .Z(n115) );
  NANDN U219 ( .A(n3835), .B(n3995), .Z(n116) );
  AND U220 ( .A(n115), .B(n116), .Z(n3924) );
  XOR U221 ( .A(n3915), .B(n3914), .Z(n3912) );
  XNOR U222 ( .A(n4065), .B(n4064), .Z(n4054) );
  NANDN U223 ( .A(n482), .B(n481), .Z(n117) );
  NANDN U224 ( .A(n483), .B(n484), .Z(n118) );
  AND U225 ( .A(n117), .B(n118), .Z(n655) );
  XOR U226 ( .A(n1050), .B(n1049), .Z(n1048) );
  NAND U227 ( .A(n1007), .B(n861), .Z(n119) );
  NANDN U228 ( .A(n862), .B(n863), .Z(n120) );
  AND U229 ( .A(n119), .B(n120), .Z(n920) );
  XOR U230 ( .A(n1501), .B(n1500), .Z(n1498) );
  XOR U231 ( .A(n1934), .B(n1933), .Z(n1931) );
  XOR U232 ( .A(n2358), .B(n2357), .Z(n2209) );
  XOR U233 ( .A(n2633), .B(n2632), .Z(n2630) );
  NAND U234 ( .A(n3189), .B(n3188), .Z(n121) );
  NANDN U235 ( .A(n3186), .B(n3187), .Z(n122) );
  AND U236 ( .A(n121), .B(n122), .Z(n3197) );
  NANDN U237 ( .A(n3476), .B(n3475), .Z(n123) );
  NANDN U238 ( .A(n3477), .B(n3478), .Z(n124) );
  NAND U239 ( .A(n123), .B(n124), .Z(n3487) );
  XNOR U240 ( .A(n3911), .B(n3910), .Z(n3909) );
  XOR U241 ( .A(n751), .B(n750), .Z(n752) );
  XOR U242 ( .A(n1150), .B(n1149), .Z(n1151) );
  XOR U243 ( .A(n3725), .B(n3724), .Z(n3726) );
  XOR U244 ( .A(n809), .B(n808), .Z(n778) );
  XOR U245 ( .A(n1192), .B(n1191), .Z(n1193) );
  XOR U246 ( .A(n1199), .B(n1198), .Z(n1185) );
  XOR U247 ( .A(n1589), .B(n1588), .Z(n1590) );
  XOR U248 ( .A(n2028), .B(n2027), .Z(n2029) );
  XOR U249 ( .A(n2457), .B(n2456), .Z(n2458) );
  XOR U250 ( .A(n2880), .B(n2879), .Z(n2881) );
  XOR U251 ( .A(n3313), .B(n3312), .Z(n3314) );
  XOR U252 ( .A(n537), .B(n451), .Z(n452) );
  XOR U253 ( .A(n556), .B(n419), .Z(n420) );
  XOR U254 ( .A(n790), .B(n789), .Z(n791) );
  XOR U255 ( .A(n797), .B(n796), .Z(n783) );
  XOR U256 ( .A(n1287), .B(n1400), .Z(n1288) );
  XOR U257 ( .A(n1643), .B(n1642), .Z(n1644) );
  XOR U258 ( .A(n1651), .B(n1650), .Z(n1655) );
  XOR U259 ( .A(n1807), .B(n1727), .Z(n1728) );
  XOR U260 ( .A(n2116), .B(n2115), .Z(n2069) );
  XNOR U261 ( .A(n2086), .B(n2085), .Z(n2063) );
  XOR U262 ( .A(n2582), .B(n2504), .Z(n2505) );
  XOR U263 ( .A(n2946), .B(n2945), .Z(n2950) );
  XOR U264 ( .A(n2917), .B(n2916), .Z(n2954) );
  XOR U265 ( .A(n3000), .B(n3080), .Z(n3002) );
  XOR U266 ( .A(n3524), .B(n3413), .Z(n3414) );
  XOR U267 ( .A(n3767), .B(n3766), .Z(n3768) );
  XOR U268 ( .A(n3774), .B(n3773), .Z(n3760) );
  NAND U269 ( .A(n250), .B(n248), .Z(n125) );
  XOR U270 ( .A(n250), .B(n248), .Z(n126) );
  NANDN U271 ( .A(n249), .B(n126), .Z(n127) );
  NAND U272 ( .A(n125), .B(n127), .Z(n269) );
  NANDN U273 ( .A(n302), .B(n301), .Z(n128) );
  NANDN U274 ( .A(n299), .B(n300), .Z(n129) );
  AND U275 ( .A(n128), .B(n129), .Z(n354) );
  XOR U276 ( .A(n512), .B(n511), .Z(n509) );
  NANDN U277 ( .A(n362), .B(n361), .Z(n130) );
  NANDN U278 ( .A(n359), .B(n360), .Z(n131) );
  AND U279 ( .A(n130), .B(n131), .Z(n486) );
  XOR U280 ( .A(n532), .B(n531), .Z(n529) );
  NAND U281 ( .A(n671), .B(n672), .Z(n132) );
  XOR U282 ( .A(n671), .B(n672), .Z(n133) );
  NANDN U283 ( .A(n670), .B(n133), .Z(n134) );
  NAND U284 ( .A(n132), .B(n134), .Z(n692) );
  XOR U285 ( .A(n1319), .B(n1318), .Z(n1321) );
  XOR U286 ( .A(n1270), .B(n1269), .Z(n1271) );
  XNOR U287 ( .A(n1345), .B(n1344), .Z(n1343) );
  XNOR U288 ( .A(n1339), .B(n1338), .Z(n1337) );
  XOR U289 ( .A(n1256), .B(n1433), .Z(n1257) );
  XNOR U290 ( .A(n1489), .B(n1488), .Z(n1487) );
  XOR U291 ( .A(n1514), .B(n1513), .Z(n135) );
  NANDN U292 ( .A(n1512), .B(n135), .Z(n136) );
  NAND U293 ( .A(n1514), .B(n1513), .Z(n137) );
  AND U294 ( .A(n136), .B(n137), .Z(n1534) );
  NANDN U295 ( .A(n1566), .B(n1565), .Z(n138) );
  NANDN U296 ( .A(n1563), .B(n1564), .Z(n139) );
  AND U297 ( .A(n138), .B(n139), .Z(n1671) );
  NANDN U298 ( .A(n1641), .B(n1640), .Z(n140) );
  NANDN U299 ( .A(n1638), .B(n1639), .Z(n141) );
  NAND U300 ( .A(n140), .B(n141), .Z(n1750) );
  XNOR U301 ( .A(n1776), .B(n1775), .Z(n1774) );
  XNOR U302 ( .A(n1685), .B(n1684), .Z(n1679) );
  NANDN U303 ( .A(n1697), .B(n1696), .Z(n142) );
  NANDN U304 ( .A(n1694), .B(n1695), .Z(n143) );
  AND U305 ( .A(n142), .B(n143), .Z(n1916) );
  XNOR U306 ( .A(n1782), .B(n1781), .Z(n1780) );
  XOR U307 ( .A(n1951), .B(n1950), .Z(n144) );
  NANDN U308 ( .A(n1949), .B(n144), .Z(n145) );
  NAND U309 ( .A(n1951), .B(n1950), .Z(n146) );
  AND U310 ( .A(n145), .B(n146), .Z(n1972) );
  NANDN U311 ( .A(n2005), .B(n2004), .Z(n147) );
  NANDN U312 ( .A(n2002), .B(n2003), .Z(n148) );
  AND U313 ( .A(n147), .B(n148), .Z(n2057) );
  XOR U314 ( .A(n2158), .B(n2157), .Z(n2186) );
  XNOR U315 ( .A(n2196), .B(n2195), .Z(n2198) );
  XOR U316 ( .A(n2190), .B(n2189), .Z(n2192) );
  XOR U317 ( .A(n2216), .B(n2215), .Z(n2213) );
  AND U318 ( .A(x[37]), .B(y[34]), .Z(n149) );
  NAND U319 ( .A(y[15]), .B(x[24]), .Z(n150) );
  XNOR U320 ( .A(n149), .B(n150), .Z(n151) );
  AND U321 ( .A(x[29]), .B(y[10]), .Z(n152) );
  NAND U322 ( .A(x[31]), .B(y[8]), .Z(n153) );
  XNOR U323 ( .A(n152), .B(n153), .Z(n154) );
  AND U324 ( .A(y[58]), .B(x[45]), .Z(n155) );
  AND U325 ( .A(y[57]), .B(x[46]), .Z(n156) );
  NANDN U326 ( .A(n2280), .B(n155), .Z(n157) );
  XNOR U327 ( .A(n156), .B(n157), .Z(n158) );
  AND U328 ( .A(x[36]), .B(y[35]), .Z(n159) );
  NAND U329 ( .A(y[60]), .B(x[43]), .Z(n160) );
  XNOR U330 ( .A(n159), .B(n160), .Z(n161) );
  XOR U331 ( .A(n158), .B(n161), .Z(n162) );
  XNOR U332 ( .A(n151), .B(n154), .Z(n163) );
  XNOR U333 ( .A(n162), .B(n163), .Z(n2320) );
  XOR U334 ( .A(n2381), .B(n2380), .Z(n164) );
  NANDN U335 ( .A(n2379), .B(n164), .Z(n165) );
  NAND U336 ( .A(n2381), .B(n2380), .Z(n166) );
  AND U337 ( .A(n165), .B(n166), .Z(n2401) );
  NANDN U338 ( .A(n2434), .B(n2433), .Z(n167) );
  NANDN U339 ( .A(n2431), .B(n2432), .Z(n168) );
  AND U340 ( .A(n167), .B(n168), .Z(n2538) );
  XNOR U341 ( .A(n2645), .B(n2644), .Z(n2643) );
  XOR U342 ( .A(n2655), .B(n2654), .Z(n2762) );
  XOR U343 ( .A(n2651), .B(n2650), .Z(n2648) );
  XOR U344 ( .A(n2805), .B(n2804), .Z(n169) );
  NANDN U345 ( .A(n2803), .B(n169), .Z(n170) );
  NAND U346 ( .A(n2805), .B(n2804), .Z(n171) );
  AND U347 ( .A(n170), .B(n171), .Z(n2825) );
  NANDN U348 ( .A(n2857), .B(n2856), .Z(n172) );
  NANDN U349 ( .A(n2854), .B(n2855), .Z(n173) );
  AND U350 ( .A(n172), .B(n173), .Z(n2966) );
  XOR U351 ( .A(n2982), .B(n2981), .Z(n2984) );
  XOR U352 ( .A(n3161), .B(n3160), .Z(n3053) );
  NANDN U353 ( .A(n3018), .B(n3019), .Z(n174) );
  NANDN U354 ( .A(n3016), .B(n3017), .Z(n175) );
  AND U355 ( .A(n174), .B(n175), .Z(n3193) );
  NAND U356 ( .A(n3006), .B(n3005), .Z(n176) );
  NANDN U357 ( .A(n3007), .B(n3098), .Z(n177) );
  AND U358 ( .A(n176), .B(n177), .Z(n3058) );
  NANDN U359 ( .A(n3353), .B(n3352), .Z(n178) );
  NANDN U360 ( .A(n3350), .B(n3351), .Z(n179) );
  NAND U361 ( .A(n178), .B(n179), .Z(n3430) );
  NANDN U362 ( .A(n3425), .B(n3426), .Z(n180) );
  NANDN U363 ( .A(n3428), .B(n3427), .Z(n181) );
  NAND U364 ( .A(n180), .B(n181), .Z(n3625) );
  XOR U365 ( .A(n3492), .B(n3491), .Z(n3617) );
  AND U366 ( .A(y[58]), .B(x[69]), .Z(n182) );
  NAND U367 ( .A(n3592), .B(n3593), .Z(n183) );
  NAND U368 ( .A(n3594), .B(n3595), .Z(n184) );
  AND U369 ( .A(n183), .B(n184), .Z(n185) );
  AND U370 ( .A(x[68]), .B(y[59]), .Z(n186) );
  NAND U371 ( .A(x[70]), .B(y[57]), .Z(n187) );
  XNOR U372 ( .A(n186), .B(n187), .Z(n188) );
  AND U373 ( .A(y[39]), .B(x[56]), .Z(n189) );
  NAND U374 ( .A(x[49]), .B(y[14]), .Z(n190) );
  XNOR U375 ( .A(n189), .B(n190), .Z(n191) );
  XOR U376 ( .A(n191), .B(n3596), .Z(n192) );
  XNOR U377 ( .A(n185), .B(n188), .Z(n193) );
  XNOR U378 ( .A(n192), .B(n193), .Z(n194) );
  NAND U379 ( .A(x[68]), .B(y[57]), .Z(n195) );
  NAND U380 ( .A(n182), .B(n195), .Z(n196) );
  XNOR U381 ( .A(n194), .B(n196), .Z(n3597) );
  NAND U382 ( .A(n3398), .B(n3400), .Z(n197) );
  XOR U383 ( .A(n3398), .B(n3400), .Z(n198) );
  NANDN U384 ( .A(n3399), .B(n198), .Z(n199) );
  NAND U385 ( .A(n197), .B(n199), .Z(n3479) );
  XNOR U386 ( .A(n655), .B(n654), .Z(n653) );
  NANDN U387 ( .A(n1131), .B(n1130), .Z(n200) );
  NANDN U388 ( .A(n1128), .B(n1129), .Z(n201) );
  AND U389 ( .A(n200), .B(n201), .Z(n1235) );
  XOR U390 ( .A(n1333), .B(n1332), .Z(n1330) );
  XOR U391 ( .A(n1932), .B(n1931), .Z(n1927) );
  XOR U392 ( .A(n2210), .B(n2209), .Z(n2208) );
  NANDN U393 ( .A(n2621), .B(n2620), .Z(n202) );
  NANDN U394 ( .A(n2622), .B(n2623), .Z(n203) );
  NAND U395 ( .A(n202), .B(n203), .Z(n2781) );
  XOR U396 ( .A(n3205), .B(n3204), .Z(n3203) );
  XNOR U397 ( .A(n3642), .B(n3641), .Z(n3488) );
  NANDN U398 ( .A(n3752), .B(n3751), .Z(n204) );
  NANDN U399 ( .A(n3749), .B(n3750), .Z(n205) );
  AND U400 ( .A(n204), .B(n205), .Z(n3825) );
  NAND U401 ( .A(n918), .B(n917), .Z(n206) );
  NANDN U402 ( .A(n915), .B(n916), .Z(n207) );
  AND U403 ( .A(n206), .B(n207), .Z(n208) );
  NAND U404 ( .A(n920), .B(n919), .Z(n209) );
  NAND U405 ( .A(n922), .B(n921), .Z(n210) );
  AND U406 ( .A(n209), .B(n210), .Z(n211) );
  XOR U407 ( .A(n1046), .B(n1045), .Z(n212) );
  XNOR U408 ( .A(n1032), .B(n1031), .Z(n213) );
  XNOR U409 ( .A(n212), .B(n213), .Z(n214) );
  AND U410 ( .A(n1058), .B(n1057), .Z(n215) );
  NAND U411 ( .A(n1052), .B(n1051), .Z(n216) );
  XNOR U412 ( .A(n215), .B(n216), .Z(n217) );
  XOR U413 ( .A(n214), .B(n217), .Z(n218) );
  XNOR U414 ( .A(n208), .B(n211), .Z(n219) );
  XNOR U415 ( .A(n218), .B(n219), .Z(n220) );
  NAND U416 ( .A(n1059), .B(n1060), .Z(n221) );
  NAND U417 ( .A(n1062), .B(n1061), .Z(n222) );
  NAND U418 ( .A(n221), .B(n222), .Z(n223) );
  XNOR U419 ( .A(n220), .B(n223), .Z(o[15]) );
  NAND U420 ( .A(n3907), .B(n3906), .Z(n224) );
  NANDN U421 ( .A(n3904), .B(n3905), .Z(n225) );
  AND U422 ( .A(n224), .B(n225), .Z(n226) );
  NAND U423 ( .A(n3911), .B(n3910), .Z(n227) );
  NANDN U424 ( .A(n3909), .B(n3908), .Z(n228) );
  AND U425 ( .A(n227), .B(n228), .Z(n229) );
  XOR U426 ( .A(n4051), .B(n4050), .Z(n230) );
  XNOR U427 ( .A(n4037), .B(n4036), .Z(n231) );
  XNOR U428 ( .A(n230), .B(n231), .Z(n232) );
  AND U429 ( .A(n4063), .B(n4062), .Z(n233) );
  NAND U430 ( .A(n4057), .B(n4056), .Z(n234) );
  XNOR U431 ( .A(n233), .B(n234), .Z(n235) );
  XOR U432 ( .A(n232), .B(n235), .Z(n236) );
  XNOR U433 ( .A(n226), .B(n229), .Z(n237) );
  XNOR U434 ( .A(n236), .B(n237), .Z(n238) );
  NAND U435 ( .A(n4064), .B(n4065), .Z(n239) );
  NAND U436 ( .A(n4067), .B(n4066), .Z(n240) );
  NAND U437 ( .A(n239), .B(n240), .Z(n241) );
  XNOR U438 ( .A(n238), .B(n241), .Z(o[71]) );
  AND U439 ( .A(y[24]), .B(x[8]), .Z(n243) );
  NAND U440 ( .A(y[0]), .B(x[0]), .Z(n242) );
  XNOR U441 ( .A(n243), .B(n242), .Z(n244) );
  NAND U442 ( .A(y[48]), .B(x[16]), .Z(n330) );
  XNOR U443 ( .A(n244), .B(n330), .Z(o[0]) );
  AND U444 ( .A(y[24]), .B(x[9]), .Z(n317) );
  AND U445 ( .A(y[25]), .B(x[8]), .Z(n254) );
  AND U446 ( .A(y[48]), .B(x[17]), .Z(n253) );
  XOR U447 ( .A(n254), .B(n253), .Z(n255) );
  XNOR U448 ( .A(n317), .B(n255), .Z(n250) );
  AND U449 ( .A(y[1]), .B(x[0]), .Z(n281) );
  AND U450 ( .A(y[49]), .B(x[16]), .Z(n288) );
  AND U451 ( .A(x[1]), .B(y[0]), .Z(n258) );
  XOR U452 ( .A(n288), .B(n258), .Z(n259) );
  XNOR U453 ( .A(n281), .B(n259), .Z(n248) );
  NANDN U454 ( .A(n243), .B(n242), .Z(n246) );
  NAND U455 ( .A(n244), .B(n330), .Z(n245) );
  AND U456 ( .A(n246), .B(n245), .Z(n249) );
  XNOR U457 ( .A(n248), .B(n249), .Z(n247) );
  XNOR U458 ( .A(n250), .B(n247), .Z(o[1]) );
  AND U459 ( .A(x[0]), .B(y[2]), .Z(n252) );
  NAND U460 ( .A(y[1]), .B(x[1]), .Z(n251) );
  XNOR U461 ( .A(n252), .B(n251), .Z(n283) );
  AND U462 ( .A(y[24]), .B(x[10]), .Z(n282) );
  XOR U463 ( .A(n283), .B(n282), .Z(n296) );
  AND U464 ( .A(y[26]), .B(x[8]), .Z(n294) );
  NAND U465 ( .A(y[25]), .B(x[9]), .Z(n293) );
  XNOR U466 ( .A(n294), .B(n293), .Z(n295) );
  XOR U467 ( .A(n296), .B(n295), .Z(n270) );
  XNOR U468 ( .A(n269), .B(n270), .Z(n272) );
  NAND U469 ( .A(n254), .B(n253), .Z(n257) );
  NAND U470 ( .A(n317), .B(n255), .Z(n256) );
  NAND U471 ( .A(n257), .B(n256), .Z(n265) );
  NAND U472 ( .A(n288), .B(n258), .Z(n261) );
  NAND U473 ( .A(n281), .B(n259), .Z(n260) );
  NAND U474 ( .A(n261), .B(n260), .Z(n263) );
  AND U475 ( .A(y[0]), .B(x[2]), .Z(n309) );
  NAND U476 ( .A(x[18]), .B(y[48]), .Z(n275) );
  XNOR U477 ( .A(n309), .B(n275), .Z(n277) );
  AND U478 ( .A(x[17]), .B(y[49]), .Z(n323) );
  NAND U479 ( .A(x[16]), .B(y[50]), .Z(n262) );
  XNOR U480 ( .A(n323), .B(n262), .Z(n276) );
  XOR U481 ( .A(n277), .B(n276), .Z(n264) );
  XNOR U482 ( .A(n263), .B(n264), .Z(n266) );
  XOR U483 ( .A(n265), .B(n266), .Z(n271) );
  XNOR U484 ( .A(n272), .B(n271), .Z(o[2]) );
  NAND U485 ( .A(n264), .B(n263), .Z(n268) );
  NANDN U486 ( .A(n266), .B(n265), .Z(n267) );
  AND U487 ( .A(n268), .B(n267), .Z(n304) );
  NANDN U488 ( .A(n270), .B(n269), .Z(n274) );
  NAND U489 ( .A(n272), .B(n271), .Z(n273) );
  AND U490 ( .A(n274), .B(n273), .Z(n303) );
  XNOR U491 ( .A(n304), .B(n303), .Z(n306) );
  NANDN U492 ( .A(n275), .B(n309), .Z(n279) );
  NAND U493 ( .A(n277), .B(n276), .Z(n278) );
  NAND U494 ( .A(n279), .B(n278), .Z(n337) );
  AND U495 ( .A(y[27]), .B(x[8]), .Z(n324) );
  AND U496 ( .A(x[1]), .B(y[2]), .Z(n325) );
  NAND U497 ( .A(y[3]), .B(x[0]), .Z(n327) );
  XNOR U498 ( .A(n326), .B(n327), .Z(n336) );
  AND U499 ( .A(x[9]), .B(y[26]), .Z(n386) );
  NAND U500 ( .A(x[11]), .B(y[24]), .Z(n280) );
  XNOR U501 ( .A(n386), .B(n280), .Z(n319) );
  AND U502 ( .A(y[25]), .B(x[10]), .Z(n318) );
  XOR U503 ( .A(n319), .B(n318), .Z(n335) );
  XOR U504 ( .A(n336), .B(n335), .Z(n338) );
  XOR U505 ( .A(n337), .B(n338), .Z(n300) );
  NAND U506 ( .A(n325), .B(n281), .Z(n285) );
  NAND U507 ( .A(n283), .B(n282), .Z(n284) );
  NAND U508 ( .A(n285), .B(n284), .Z(n343) );
  AND U509 ( .A(y[1]), .B(x[2]), .Z(n287) );
  NAND U510 ( .A(x[3]), .B(y[0]), .Z(n286) );
  XNOR U511 ( .A(n287), .B(n286), .Z(n310) );
  AND U512 ( .A(x[17]), .B(y[50]), .Z(n292) );
  NAND U513 ( .A(n288), .B(n292), .Z(n311) );
  XNOR U514 ( .A(n310), .B(n311), .Z(n342) );
  AND U515 ( .A(x[19]), .B(y[48]), .Z(n290) );
  NAND U516 ( .A(x[16]), .B(y[51]), .Z(n289) );
  XNOR U517 ( .A(n290), .B(n289), .Z(n332) );
  NAND U518 ( .A(y[49]), .B(x[18]), .Z(n291) );
  XNOR U519 ( .A(n292), .B(n291), .Z(n331) );
  XOR U520 ( .A(n332), .B(n331), .Z(n341) );
  XOR U521 ( .A(n342), .B(n341), .Z(n344) );
  XNOR U522 ( .A(n343), .B(n344), .Z(n299) );
  XNOR U523 ( .A(n300), .B(n299), .Z(n301) );
  NANDN U524 ( .A(n294), .B(n293), .Z(n298) );
  NANDN U525 ( .A(n296), .B(n295), .Z(n297) );
  NAND U526 ( .A(n298), .B(n297), .Z(n302) );
  XNOR U527 ( .A(n301), .B(n302), .Z(n305) );
  XOR U528 ( .A(n306), .B(n305), .Z(o[3]) );
  NANDN U529 ( .A(n304), .B(n303), .Z(n308) );
  NAND U530 ( .A(n306), .B(n305), .Z(n307) );
  NAND U531 ( .A(n308), .B(n307), .Z(n353) );
  XNOR U532 ( .A(n354), .B(n353), .Z(n356) );
  AND U533 ( .A(x[3]), .B(y[1]), .Z(n377) );
  NAND U534 ( .A(n377), .B(n309), .Z(n313) );
  NANDN U535 ( .A(n311), .B(n310), .Z(n312) );
  AND U536 ( .A(n313), .B(n312), .Z(n409) );
  AND U537 ( .A(x[19]), .B(y[49]), .Z(n432) );
  NAND U538 ( .A(y[50]), .B(x[18]), .Z(n314) );
  XNOR U539 ( .A(n432), .B(n314), .Z(n369) );
  NAND U540 ( .A(y[48]), .B(x[20]), .Z(n370) );
  XNOR U541 ( .A(n369), .B(n370), .Z(n371) );
  NAND U542 ( .A(y[51]), .B(x[17]), .Z(n372) );
  XNOR U543 ( .A(n371), .B(n372), .Z(n406) );
  AND U544 ( .A(y[27]), .B(x[9]), .Z(n316) );
  NAND U545 ( .A(x[10]), .B(y[26]), .Z(n315) );
  XNOR U546 ( .A(n316), .B(n315), .Z(n387) );
  NAND U547 ( .A(y[25]), .B(x[11]), .Z(n388) );
  XOR U548 ( .A(n387), .B(n388), .Z(n407) );
  XNOR U549 ( .A(n406), .B(n407), .Z(n408) );
  XNOR U550 ( .A(n409), .B(n408), .Z(n363) );
  AND U551 ( .A(y[26]), .B(x[11]), .Z(n419) );
  NAND U552 ( .A(n419), .B(n317), .Z(n321) );
  NAND U553 ( .A(n319), .B(n318), .Z(n320) );
  AND U554 ( .A(n321), .B(n320), .Z(n403) );
  AND U555 ( .A(y[52]), .B(x[16]), .Z(n446) );
  AND U556 ( .A(x[18]), .B(y[50]), .Z(n322) );
  AND U557 ( .A(n323), .B(n322), .Z(n379) );
  NAND U558 ( .A(y[0]), .B(x[4]), .Z(n380) );
  XOR U559 ( .A(n379), .B(n380), .Z(n381) );
  XNOR U560 ( .A(n446), .B(n381), .Z(n400) );
  AND U561 ( .A(y[24]), .B(x[12]), .Z(n435) );
  AND U562 ( .A(y[28]), .B(x[8]), .Z(n391) );
  XOR U563 ( .A(n435), .B(n391), .Z(n393) );
  NAND U564 ( .A(x[1]), .B(y[3]), .Z(n392) );
  XOR U565 ( .A(n393), .B(n392), .Z(n401) );
  XNOR U566 ( .A(n400), .B(n401), .Z(n402) );
  XOR U567 ( .A(n403), .B(n402), .Z(n364) );
  XNOR U568 ( .A(n363), .B(n364), .Z(n365) );
  NAND U569 ( .A(n325), .B(n324), .Z(n329) );
  NANDN U570 ( .A(n327), .B(n326), .Z(n328) );
  AND U571 ( .A(n329), .B(n328), .Z(n362) );
  AND U572 ( .A(y[2]), .B(x[2]), .Z(n376) );
  NAND U573 ( .A(y[4]), .B(x[0]), .Z(n378) );
  XNOR U574 ( .A(n377), .B(n378), .Z(n375) );
  XNOR U575 ( .A(n376), .B(n375), .Z(n359) );
  AND U576 ( .A(y[51]), .B(x[19]), .Z(n602) );
  NANDN U577 ( .A(n330), .B(n602), .Z(n334) );
  NAND U578 ( .A(n332), .B(n331), .Z(n333) );
  NAND U579 ( .A(n334), .B(n333), .Z(n360) );
  XNOR U580 ( .A(n359), .B(n360), .Z(n361) );
  XOR U581 ( .A(n362), .B(n361), .Z(n366) );
  XOR U582 ( .A(n365), .B(n366), .Z(n349) );
  NAND U583 ( .A(n336), .B(n335), .Z(n340) );
  NAND U584 ( .A(n338), .B(n337), .Z(n339) );
  AND U585 ( .A(n340), .B(n339), .Z(n348) );
  NAND U586 ( .A(n342), .B(n341), .Z(n346) );
  NAND U587 ( .A(n344), .B(n343), .Z(n345) );
  AND U588 ( .A(n346), .B(n345), .Z(n347) );
  XOR U589 ( .A(n348), .B(n347), .Z(n350) );
  XNOR U590 ( .A(n349), .B(n350), .Z(n355) );
  XOR U591 ( .A(n356), .B(n355), .Z(o[4]) );
  NAND U592 ( .A(n348), .B(n347), .Z(n352) );
  NAND U593 ( .A(n350), .B(n349), .Z(n351) );
  AND U594 ( .A(n352), .B(n351), .Z(n492) );
  NANDN U595 ( .A(n354), .B(n353), .Z(n358) );
  NAND U596 ( .A(n356), .B(n355), .Z(n357) );
  AND U597 ( .A(n358), .B(n357), .Z(n491) );
  XNOR U598 ( .A(n492), .B(n491), .Z(n494) );
  NANDN U599 ( .A(n364), .B(n363), .Z(n368) );
  NANDN U600 ( .A(n366), .B(n365), .Z(n367) );
  NAND U601 ( .A(n368), .B(n367), .Z(n485) );
  XNOR U602 ( .A(n486), .B(n485), .Z(n488) );
  NANDN U603 ( .A(n370), .B(n369), .Z(n374) );
  NANDN U604 ( .A(n372), .B(n371), .Z(n373) );
  AND U605 ( .A(n374), .B(n373), .Z(n441) );
  XNOR U606 ( .A(n441), .B(n440), .Z(n442) );
  NANDN U607 ( .A(n380), .B(n379), .Z(n383) );
  NANDN U608 ( .A(n381), .B(n446), .Z(n382) );
  AND U609 ( .A(n383), .B(n382), .Z(n416) );
  AND U610 ( .A(y[24]), .B(x[13]), .Z(n385) );
  NAND U611 ( .A(x[12]), .B(y[25]), .Z(n384) );
  XNOR U612 ( .A(n385), .B(n384), .Z(n437) );
  AND U613 ( .A(y[4]), .B(x[1]), .Z(n436) );
  XOR U614 ( .A(n437), .B(n436), .Z(n413) );
  AND U615 ( .A(y[51]), .B(x[18]), .Z(n427) );
  AND U616 ( .A(y[48]), .B(x[21]), .Z(n426) );
  XOR U617 ( .A(n427), .B(n426), .Z(n429) );
  AND U618 ( .A(x[20]), .B(y[49]), .Z(n615) );
  AND U619 ( .A(x[19]), .B(y[50]), .Z(n397) );
  XOR U620 ( .A(n615), .B(n397), .Z(n428) );
  XNOR U621 ( .A(n429), .B(n428), .Z(n412) );
  XNOR U622 ( .A(n413), .B(n412), .Z(n415) );
  XOR U623 ( .A(n416), .B(n415), .Z(n443) );
  XOR U624 ( .A(n442), .B(n443), .Z(n479) );
  AND U625 ( .A(x[10]), .B(y[27]), .Z(n451) );
  NAND U626 ( .A(n451), .B(n386), .Z(n390) );
  NANDN U627 ( .A(n388), .B(n387), .Z(n389) );
  AND U628 ( .A(n390), .B(n389), .Z(n474) );
  AND U629 ( .A(y[0]), .B(x[5]), .Z(n537) );
  NAND U630 ( .A(x[4]), .B(y[1]), .Z(n453) );
  XNOR U631 ( .A(n452), .B(n453), .Z(n471) );
  AND U632 ( .A(y[28]), .B(x[9]), .Z(n613) );
  AND U633 ( .A(x[0]), .B(y[5]), .Z(n458) );
  NAND U634 ( .A(y[29]), .B(x[8]), .Z(n459) );
  XOR U635 ( .A(n458), .B(n459), .Z(n460) );
  XOR U636 ( .A(n613), .B(n460), .Z(n472) );
  XNOR U637 ( .A(n471), .B(n472), .Z(n473) );
  XNOR U638 ( .A(n474), .B(n473), .Z(n477) );
  NAND U639 ( .A(n435), .B(n391), .Z(n395) );
  ANDN U640 ( .B(n393), .A(n392), .Z(n394) );
  ANDN U641 ( .B(n395), .A(n394), .Z(n468) );
  AND U642 ( .A(x[18]), .B(y[49]), .Z(n396) );
  AND U643 ( .A(n397), .B(n396), .Z(n447) );
  AND U644 ( .A(y[53]), .B(x[16]), .Z(n399) );
  NAND U645 ( .A(y[52]), .B(x[17]), .Z(n398) );
  XOR U646 ( .A(n399), .B(n398), .Z(n448) );
  XNOR U647 ( .A(n447), .B(n448), .Z(n465) );
  AND U648 ( .A(y[2]), .B(x[3]), .Z(n556) );
  NAND U649 ( .A(y[3]), .B(x[2]), .Z(n421) );
  XOR U650 ( .A(n420), .B(n421), .Z(n466) );
  XNOR U651 ( .A(n465), .B(n466), .Z(n467) );
  XOR U652 ( .A(n468), .B(n467), .Z(n478) );
  XOR U653 ( .A(n477), .B(n478), .Z(n480) );
  XNOR U654 ( .A(n479), .B(n480), .Z(n483) );
  NANDN U655 ( .A(n401), .B(n400), .Z(n405) );
  NANDN U656 ( .A(n403), .B(n402), .Z(n404) );
  AND U657 ( .A(n405), .B(n404), .Z(n482) );
  NANDN U658 ( .A(n407), .B(n406), .Z(n411) );
  NANDN U659 ( .A(n409), .B(n408), .Z(n410) );
  NAND U660 ( .A(n411), .B(n410), .Z(n481) );
  XNOR U661 ( .A(n482), .B(n481), .Z(n484) );
  XNOR U662 ( .A(n483), .B(n484), .Z(n487) );
  XNOR U663 ( .A(n488), .B(n487), .Z(n493) );
  XNOR U664 ( .A(n494), .B(n493), .Z(o[5]) );
  IV U665 ( .A(n412), .Z(n414) );
  NAND U666 ( .A(n414), .B(n413), .Z(n418) );
  NANDN U667 ( .A(n416), .B(n415), .Z(n417) );
  AND U668 ( .A(n418), .B(n417), .Z(n506) );
  NAND U669 ( .A(n556), .B(n419), .Z(n423) );
  NANDN U670 ( .A(n421), .B(n420), .Z(n422) );
  AND U671 ( .A(n423), .B(n422), .Z(n522) );
  AND U672 ( .A(y[29]), .B(x[9]), .Z(n425) );
  NAND U673 ( .A(x[10]), .B(y[28]), .Z(n424) );
  XNOR U674 ( .A(n425), .B(n424), .Z(n611) );
  AND U675 ( .A(y[4]), .B(x[2]), .Z(n610) );
  XNOR U676 ( .A(n611), .B(n610), .Z(n524) );
  NAND U677 ( .A(n427), .B(n426), .Z(n431) );
  NAND U678 ( .A(n429), .B(n428), .Z(n430) );
  AND U679 ( .A(n431), .B(n430), .Z(n523) );
  XOR U680 ( .A(n522), .B(n521), .Z(n505) );
  XOR U681 ( .A(n506), .B(n505), .Z(n504) );
  AND U682 ( .A(x[17]), .B(y[53]), .Z(n585) );
  AND U683 ( .A(y[50]), .B(x[20]), .Z(n457) );
  AND U684 ( .A(n457), .B(n432), .Z(n587) );
  AND U685 ( .A(x[18]), .B(y[52]), .Z(n586) );
  XOR U686 ( .A(n587), .B(n586), .Z(n584) );
  XNOR U687 ( .A(n585), .B(n584), .Z(n516) );
  AND U688 ( .A(y[3]), .B(x[3]), .Z(n434) );
  NAND U689 ( .A(y[2]), .B(x[4]), .Z(n433) );
  XNOR U690 ( .A(n434), .B(n433), .Z(n555) );
  AND U691 ( .A(x[12]), .B(y[26]), .Z(n554) );
  XNOR U692 ( .A(n555), .B(n554), .Z(n518) );
  AND U693 ( .A(y[25]), .B(x[13]), .Z(n541) );
  NAND U694 ( .A(n541), .B(n435), .Z(n439) );
  NAND U695 ( .A(n437), .B(n436), .Z(n438) );
  AND U696 ( .A(n439), .B(n438), .Z(n517) );
  XNOR U697 ( .A(n504), .B(n503), .Z(n500) );
  NANDN U698 ( .A(n441), .B(n440), .Z(n445) );
  NANDN U699 ( .A(n443), .B(n442), .Z(n444) );
  NAND U700 ( .A(n445), .B(n444), .Z(n499) );
  NAND U701 ( .A(n446), .B(n585), .Z(n450) );
  NANDN U702 ( .A(n448), .B(n447), .Z(n449) );
  AND U703 ( .A(n450), .B(n449), .Z(n637) );
  NAND U704 ( .A(n537), .B(n451), .Z(n455) );
  NANDN U705 ( .A(n453), .B(n452), .Z(n454) );
  AND U706 ( .A(n455), .B(n454), .Z(n510) );
  AND U707 ( .A(y[24]), .B(x[14]), .Z(n543) );
  AND U708 ( .A(x[0]), .B(y[6]), .Z(n542) );
  XOR U709 ( .A(n543), .B(n542), .Z(n540) );
  XNOR U710 ( .A(n541), .B(n540), .Z(n512) );
  NAND U711 ( .A(y[49]), .B(x[21]), .Z(n456) );
  XNOR U712 ( .A(n457), .B(n456), .Z(n605) );
  AND U713 ( .A(y[48]), .B(x[22]), .Z(n604) );
  XOR U714 ( .A(n605), .B(n604), .Z(n603) );
  XNOR U715 ( .A(n603), .B(n602), .Z(n511) );
  XOR U716 ( .A(n510), .B(n509), .Z(n636) );
  XOR U717 ( .A(n637), .B(n636), .Z(n635) );
  NANDN U718 ( .A(n459), .B(n458), .Z(n462) );
  NANDN U719 ( .A(n460), .B(n613), .Z(n461) );
  AND U720 ( .A(n462), .B(n461), .Z(n530) );
  AND U721 ( .A(x[5]), .B(y[1]), .Z(n464) );
  NAND U722 ( .A(x[6]), .B(y[0]), .Z(n463) );
  XNOR U723 ( .A(n464), .B(n463), .Z(n536) );
  AND U724 ( .A(x[11]), .B(y[27]), .Z(n535) );
  XNOR U725 ( .A(n536), .B(n535), .Z(n532) );
  AND U726 ( .A(x[1]), .B(y[5]), .Z(n549) );
  AND U727 ( .A(x[16]), .B(y[54]), .Z(n551) );
  AND U728 ( .A(x[8]), .B(y[30]), .Z(n550) );
  XOR U729 ( .A(n551), .B(n550), .Z(n548) );
  XNOR U730 ( .A(n549), .B(n548), .Z(n531) );
  XOR U731 ( .A(n530), .B(n529), .Z(n634) );
  XOR U732 ( .A(n635), .B(n634), .Z(n629) );
  NANDN U733 ( .A(n466), .B(n465), .Z(n470) );
  NANDN U734 ( .A(n468), .B(n467), .Z(n469) );
  NAND U735 ( .A(n470), .B(n469), .Z(n631) );
  NANDN U736 ( .A(n472), .B(n471), .Z(n476) );
  NANDN U737 ( .A(n474), .B(n473), .Z(n475) );
  NAND U738 ( .A(n476), .B(n475), .Z(n630) );
  XOR U739 ( .A(n631), .B(n630), .Z(n628) );
  XNOR U740 ( .A(n629), .B(n628), .Z(n498) );
  XNOR U741 ( .A(n497), .B(n498), .Z(n652) );
  XOR U742 ( .A(n652), .B(n653), .Z(n649) );
  NANDN U743 ( .A(n486), .B(n485), .Z(n490) );
  NAND U744 ( .A(n488), .B(n487), .Z(n489) );
  NAND U745 ( .A(n490), .B(n489), .Z(n648) );
  XOR U746 ( .A(n649), .B(n648), .Z(n647) );
  NANDN U747 ( .A(n492), .B(n491), .Z(n496) );
  NAND U748 ( .A(n494), .B(n493), .Z(n495) );
  AND U749 ( .A(n496), .B(n495), .Z(n646) );
  XOR U750 ( .A(n647), .B(n646), .Z(o[6]) );
  NAND U751 ( .A(n498), .B(n497), .Z(n502) );
  NAND U752 ( .A(n500), .B(n499), .Z(n501) );
  AND U753 ( .A(n502), .B(n501), .Z(n663) );
  NAND U754 ( .A(n504), .B(n503), .Z(n508) );
  NAND U755 ( .A(n506), .B(n505), .Z(n507) );
  AND U756 ( .A(n508), .B(n507), .Z(n645) );
  NAND U757 ( .A(n510), .B(n509), .Z(n514) );
  NAND U758 ( .A(n512), .B(n511), .Z(n513) );
  AND U759 ( .A(n514), .B(n513), .Z(n627) );
  NAND U760 ( .A(n516), .B(n515), .Z(n520) );
  NAND U761 ( .A(n518), .B(n517), .Z(n519) );
  AND U762 ( .A(n520), .B(n519), .Z(n528) );
  NAND U763 ( .A(n522), .B(n521), .Z(n526) );
  NAND U764 ( .A(n524), .B(n523), .Z(n525) );
  NAND U765 ( .A(n526), .B(n525), .Z(n527) );
  XNOR U766 ( .A(n528), .B(n527), .Z(n625) );
  NAND U767 ( .A(n530), .B(n529), .Z(n534) );
  NAND U768 ( .A(n532), .B(n531), .Z(n533) );
  AND U769 ( .A(n534), .B(n533), .Z(n623) );
  NAND U770 ( .A(n536), .B(n535), .Z(n539) );
  AND U771 ( .A(y[1]), .B(x[6]), .Z(n614) );
  NAND U772 ( .A(n537), .B(n614), .Z(n538) );
  AND U773 ( .A(n539), .B(n538), .Z(n547) );
  NAND U774 ( .A(n541), .B(n540), .Z(n545) );
  NAND U775 ( .A(n543), .B(n542), .Z(n544) );
  NAND U776 ( .A(n545), .B(n544), .Z(n546) );
  XNOR U777 ( .A(n547), .B(n546), .Z(n562) );
  NAND U778 ( .A(n549), .B(n548), .Z(n553) );
  NAND U779 ( .A(n551), .B(n550), .Z(n552) );
  AND U780 ( .A(n553), .B(n552), .Z(n560) );
  NAND U781 ( .A(n555), .B(n554), .Z(n558) );
  AND U782 ( .A(x[4]), .B(y[3]), .Z(n571) );
  NAND U783 ( .A(n556), .B(n571), .Z(n557) );
  NAND U784 ( .A(n558), .B(n557), .Z(n559) );
  XNOR U785 ( .A(n560), .B(n559), .Z(n561) );
  XOR U786 ( .A(n562), .B(n561), .Z(n601) );
  AND U787 ( .A(x[23]), .B(y[48]), .Z(n564) );
  NAND U788 ( .A(x[20]), .B(y[51]), .Z(n563) );
  XNOR U789 ( .A(n564), .B(n563), .Z(n575) );
  AND U790 ( .A(y[31]), .B(x[8]), .Z(n566) );
  NAND U791 ( .A(y[55]), .B(x[16]), .Z(n565) );
  XNOR U792 ( .A(n566), .B(n565), .Z(n570) );
  AND U793 ( .A(y[6]), .B(x[1]), .Z(n568) );
  NAND U794 ( .A(x[3]), .B(y[4]), .Z(n567) );
  XNOR U795 ( .A(n568), .B(n567), .Z(n569) );
  XOR U796 ( .A(n570), .B(n569), .Z(n573) );
  AND U797 ( .A(y[29]), .B(x[10]), .Z(n612) );
  XNOR U798 ( .A(n612), .B(n571), .Z(n572) );
  XNOR U799 ( .A(n573), .B(n572), .Z(n574) );
  XOR U800 ( .A(n575), .B(n574), .Z(n583) );
  AND U801 ( .A(y[7]), .B(x[0]), .Z(n577) );
  NAND U802 ( .A(y[52]), .B(x[19]), .Z(n576) );
  XNOR U803 ( .A(n577), .B(n576), .Z(n581) );
  AND U804 ( .A(y[26]), .B(x[13]), .Z(n579) );
  NAND U805 ( .A(x[14]), .B(y[25]), .Z(n578) );
  XNOR U806 ( .A(n579), .B(n578), .Z(n580) );
  XNOR U807 ( .A(n581), .B(n580), .Z(n582) );
  XNOR U808 ( .A(n583), .B(n582), .Z(n599) );
  NAND U809 ( .A(n585), .B(n584), .Z(n589) );
  NAND U810 ( .A(n587), .B(n586), .Z(n588) );
  AND U811 ( .A(n589), .B(n588), .Z(n597) );
  AND U812 ( .A(y[5]), .B(x[2]), .Z(n591) );
  NAND U813 ( .A(y[54]), .B(x[17]), .Z(n590) );
  XNOR U814 ( .A(n591), .B(n590), .Z(n595) );
  AND U815 ( .A(y[30]), .B(x[9]), .Z(n593) );
  NAND U816 ( .A(x[22]), .B(y[49]), .Z(n592) );
  XNOR U817 ( .A(n593), .B(n592), .Z(n594) );
  XNOR U818 ( .A(n595), .B(n594), .Z(n596) );
  XNOR U819 ( .A(n597), .B(n596), .Z(n598) );
  XNOR U820 ( .A(n599), .B(n598), .Z(n600) );
  XNOR U821 ( .A(n601), .B(n600), .Z(n621) );
  NAND U822 ( .A(n603), .B(n602), .Z(n607) );
  NAND U823 ( .A(n605), .B(n604), .Z(n606) );
  AND U824 ( .A(n607), .B(n606), .Z(n619) );
  AND U825 ( .A(x[5]), .B(y[2]), .Z(n609) );
  NAND U826 ( .A(y[28]), .B(x[11]), .Z(n608) );
  XNOR U827 ( .A(n609), .B(n608), .Z(n617) );
  XNOR U828 ( .A(n617), .B(n616), .Z(n618) );
  XNOR U829 ( .A(n619), .B(n618), .Z(n620) );
  XNOR U830 ( .A(n621), .B(n620), .Z(n622) );
  XNOR U831 ( .A(n623), .B(n622), .Z(n624) );
  XNOR U832 ( .A(n625), .B(n624), .Z(n626) );
  XNOR U833 ( .A(n627), .B(n626), .Z(n643) );
  NANDN U834 ( .A(n629), .B(n628), .Z(n633) );
  NAND U835 ( .A(n631), .B(n630), .Z(n632) );
  AND U836 ( .A(n633), .B(n632), .Z(n641) );
  NAND U837 ( .A(n635), .B(n634), .Z(n639) );
  NAND U838 ( .A(n637), .B(n636), .Z(n638) );
  NAND U839 ( .A(n639), .B(n638), .Z(n640) );
  XNOR U840 ( .A(n641), .B(n640), .Z(n642) );
  XNOR U841 ( .A(n643), .B(n642), .Z(n644) );
  XNOR U842 ( .A(n645), .B(n644), .Z(n661) );
  NAND U843 ( .A(n647), .B(n646), .Z(n651) );
  NAND U844 ( .A(n649), .B(n648), .Z(n650) );
  AND U845 ( .A(n651), .B(n650), .Z(n659) );
  NANDN U846 ( .A(n653), .B(n652), .Z(n657) );
  NAND U847 ( .A(n655), .B(n654), .Z(n656) );
  NAND U848 ( .A(n657), .B(n656), .Z(n658) );
  XNOR U849 ( .A(n659), .B(n658), .Z(n660) );
  XNOR U850 ( .A(n661), .B(n660), .Z(n662) );
  XNOR U851 ( .A(n663), .B(n662), .Z(o[7]) );
  AND U852 ( .A(x[8]), .B(y[32]), .Z(n665) );
  NAND U853 ( .A(x[0]), .B(y[8]), .Z(n664) );
  XNOR U854 ( .A(n665), .B(n664), .Z(n666) );
  NAND U855 ( .A(x[16]), .B(y[56]), .Z(n756) );
  XNOR U856 ( .A(n666), .B(n756), .Z(o[8]) );
  AND U857 ( .A(x[9]), .B(y[32]), .Z(n743) );
  AND U858 ( .A(x[17]), .B(y[56]), .Z(n795) );
  AND U859 ( .A(x[8]), .B(y[33]), .Z(n675) );
  XOR U860 ( .A(n795), .B(n675), .Z(n676) );
  XOR U861 ( .A(n743), .B(n676), .Z(n672) );
  NANDN U862 ( .A(n665), .B(n664), .Z(n668) );
  NAND U863 ( .A(n666), .B(n756), .Z(n667) );
  NAND U864 ( .A(n668), .B(n667), .Z(n670) );
  AND U865 ( .A(x[0]), .B(y[9]), .Z(n703) );
  AND U866 ( .A(x[16]), .B(y[57]), .Z(n710) );
  AND U867 ( .A(x[1]), .B(y[8]), .Z(n679) );
  XOR U868 ( .A(n710), .B(n679), .Z(n680) );
  XOR U869 ( .A(n703), .B(n680), .Z(n671) );
  XOR U870 ( .A(n670), .B(n671), .Z(n669) );
  XNOR U871 ( .A(n672), .B(n669), .Z(o[9]) );
  AND U872 ( .A(y[10]), .B(x[0]), .Z(n674) );
  NAND U873 ( .A(y[9]), .B(x[1]), .Z(n673) );
  XNOR U874 ( .A(n674), .B(n673), .Z(n704) );
  NAND U875 ( .A(x[10]), .B(y[32]), .Z(n705) );
  XOR U876 ( .A(n704), .B(n705), .Z(n717) );
  NAND U877 ( .A(x[8]), .B(y[34]), .Z(n716) );
  NAND U878 ( .A(x[9]), .B(y[33]), .Z(n715) );
  XOR U879 ( .A(n716), .B(n715), .Z(n718) );
  XOR U880 ( .A(n717), .B(n718), .Z(n691) );
  XNOR U881 ( .A(n692), .B(n691), .Z(n694) );
  NAND U882 ( .A(n795), .B(n675), .Z(n678) );
  NAND U883 ( .A(n743), .B(n676), .Z(n677) );
  NAND U884 ( .A(n678), .B(n677), .Z(n687) );
  NAND U885 ( .A(n710), .B(n679), .Z(n682) );
  NAND U886 ( .A(n703), .B(n680), .Z(n681) );
  NAND U887 ( .A(n682), .B(n681), .Z(n685) );
  AND U888 ( .A(x[2]), .B(y[8]), .Z(n733) );
  NAND U889 ( .A(x[18]), .B(y[56]), .Z(n697) );
  XNOR U890 ( .A(n733), .B(n697), .Z(n699) );
  AND U891 ( .A(y[58]), .B(x[16]), .Z(n684) );
  NAND U892 ( .A(y[57]), .B(x[17]), .Z(n683) );
  XNOR U893 ( .A(n684), .B(n683), .Z(n698) );
  XOR U894 ( .A(n699), .B(n698), .Z(n686) );
  XNOR U895 ( .A(n685), .B(n686), .Z(n688) );
  XOR U896 ( .A(n687), .B(n688), .Z(n693) );
  XNOR U897 ( .A(n694), .B(n693), .Z(o[10]) );
  NAND U898 ( .A(n686), .B(n685), .Z(n690) );
  NANDN U899 ( .A(n688), .B(n687), .Z(n689) );
  AND U900 ( .A(n690), .B(n689), .Z(n722) );
  NANDN U901 ( .A(n692), .B(n691), .Z(n696) );
  NAND U902 ( .A(n694), .B(n693), .Z(n695) );
  AND U903 ( .A(n696), .B(n695), .Z(n721) );
  XNOR U904 ( .A(n722), .B(n721), .Z(n724) );
  NANDN U905 ( .A(n697), .B(n733), .Z(n701) );
  NAND U906 ( .A(n699), .B(n698), .Z(n700) );
  AND U907 ( .A(n701), .B(n700), .Z(n764) );
  AND U908 ( .A(x[8]), .B(y[35]), .Z(n750) );
  AND U909 ( .A(x[1]), .B(y[10]), .Z(n751) );
  NAND U910 ( .A(x[0]), .B(y[11]), .Z(n753) );
  XNOR U911 ( .A(n752), .B(n753), .Z(n761) );
  AND U912 ( .A(y[34]), .B(x[9]), .Z(n814) );
  NAND U913 ( .A(y[32]), .B(x[11]), .Z(n702) );
  XNOR U914 ( .A(n814), .B(n702), .Z(n744) );
  NAND U915 ( .A(x[10]), .B(y[33]), .Z(n745) );
  XOR U916 ( .A(n744), .B(n745), .Z(n762) );
  XNOR U917 ( .A(n761), .B(n762), .Z(n763) );
  XNOR U918 ( .A(n764), .B(n763), .Z(n728) );
  NAND U919 ( .A(n751), .B(n703), .Z(n707) );
  NANDN U920 ( .A(n705), .B(n704), .Z(n706) );
  AND U921 ( .A(n707), .B(n706), .Z(n769) );
  AND U922 ( .A(y[9]), .B(x[2]), .Z(n709) );
  NAND U923 ( .A(y[8]), .B(x[3]), .Z(n708) );
  XNOR U924 ( .A(n709), .B(n708), .Z(n734) );
  AND U925 ( .A(x[17]), .B(y[58]), .Z(n714) );
  NAND U926 ( .A(n710), .B(n714), .Z(n735) );
  XNOR U927 ( .A(n734), .B(n735), .Z(n767) );
  AND U928 ( .A(y[59]), .B(x[16]), .Z(n712) );
  NAND U929 ( .A(y[56]), .B(x[19]), .Z(n711) );
  XNOR U930 ( .A(n712), .B(n711), .Z(n757) );
  NAND U931 ( .A(y[57]), .B(x[18]), .Z(n713) );
  XOR U932 ( .A(n714), .B(n713), .Z(n758) );
  XOR U933 ( .A(n757), .B(n758), .Z(n768) );
  XOR U934 ( .A(n767), .B(n768), .Z(n770) );
  XOR U935 ( .A(n769), .B(n770), .Z(n727) );
  XOR U936 ( .A(n728), .B(n727), .Z(n730) );
  NAND U937 ( .A(n716), .B(n715), .Z(n720) );
  NAND U938 ( .A(n718), .B(n717), .Z(n719) );
  AND U939 ( .A(n720), .B(n719), .Z(n729) );
  XOR U940 ( .A(n730), .B(n729), .Z(n723) );
  XOR U941 ( .A(n724), .B(n723), .Z(o[11]) );
  NANDN U942 ( .A(n722), .B(n721), .Z(n726) );
  NAND U943 ( .A(n724), .B(n723), .Z(n725) );
  AND U944 ( .A(n726), .B(n725), .Z(n835) );
  NAND U945 ( .A(n728), .B(n727), .Z(n732) );
  NAND U946 ( .A(n730), .B(n729), .Z(n731) );
  NAND U947 ( .A(n732), .B(n731), .Z(n836) );
  XNOR U948 ( .A(n835), .B(n836), .Z(n838) );
  NAND U949 ( .A(x[3]), .B(y[9]), .Z(n811) );
  NANDN U950 ( .A(n811), .B(n733), .Z(n737) );
  NANDN U951 ( .A(n735), .B(n734), .Z(n736) );
  NAND U952 ( .A(n737), .B(n736), .Z(n786) );
  AND U953 ( .A(y[34]), .B(x[10]), .Z(n739) );
  NAND U954 ( .A(y[35]), .B(x[9]), .Z(n738) );
  XNOR U955 ( .A(n739), .B(n738), .Z(n815) );
  NAND U956 ( .A(x[11]), .B(y[33]), .Z(n816) );
  XNOR U957 ( .A(n815), .B(n816), .Z(n784) );
  AND U958 ( .A(y[59]), .B(x[17]), .Z(n741) );
  NAND U959 ( .A(y[56]), .B(x[20]), .Z(n740) );
  XNOR U960 ( .A(n741), .B(n740), .Z(n796) );
  AND U961 ( .A(y[57]), .B(x[19]), .Z(n900) );
  NAND U962 ( .A(y[58]), .B(x[18]), .Z(n742) );
  XNOR U963 ( .A(n900), .B(n742), .Z(n797) );
  XOR U964 ( .A(n784), .B(n783), .Z(n785) );
  NAND U965 ( .A(x[11]), .B(y[34]), .Z(n828) );
  IV U966 ( .A(n828), .Z(n890) );
  NAND U967 ( .A(n890), .B(n743), .Z(n747) );
  NANDN U968 ( .A(n745), .B(n744), .Z(n746) );
  NAND U969 ( .A(n747), .B(n746), .Z(n792) );
  AND U970 ( .A(x[16]), .B(y[60]), .Z(n857) );
  AND U971 ( .A(x[18]), .B(y[58]), .Z(n749) );
  AND U972 ( .A(x[17]), .B(y[57]), .Z(n748) );
  AND U973 ( .A(n749), .B(n748), .Z(n800) );
  NAND U974 ( .A(x[4]), .B(y[8]), .Z(n801) );
  XOR U975 ( .A(n800), .B(n801), .Z(n802) );
  XNOR U976 ( .A(n857), .B(n802), .Z(n789) );
  AND U977 ( .A(x[12]), .B(y[32]), .Z(n903) );
  AND U978 ( .A(x[8]), .B(y[36]), .Z(n819) );
  XOR U979 ( .A(n903), .B(n819), .Z(n820) );
  NAND U980 ( .A(x[1]), .B(y[11]), .Z(n821) );
  XNOR U981 ( .A(n820), .B(n821), .Z(n790) );
  XNOR U982 ( .A(n774), .B(n773), .Z(n776) );
  NAND U983 ( .A(n751), .B(n750), .Z(n755) );
  NANDN U984 ( .A(n753), .B(n752), .Z(n754) );
  NAND U985 ( .A(n755), .B(n754), .Z(n779) );
  NAND U986 ( .A(x[2]), .B(y[10]), .Z(n809) );
  NAND U987 ( .A(x[0]), .B(y[12]), .Z(n810) );
  XOR U988 ( .A(n811), .B(n810), .Z(n808) );
  AND U989 ( .A(x[19]), .B(y[59]), .Z(n943) );
  NANDN U990 ( .A(n756), .B(n943), .Z(n760) );
  NANDN U991 ( .A(n758), .B(n757), .Z(n759) );
  NAND U992 ( .A(n760), .B(n759), .Z(n777) );
  XNOR U993 ( .A(n778), .B(n777), .Z(n780) );
  XOR U994 ( .A(n779), .B(n780), .Z(n775) );
  XOR U995 ( .A(n776), .B(n775), .Z(n832) );
  NANDN U996 ( .A(n762), .B(n761), .Z(n766) );
  NANDN U997 ( .A(n764), .B(n763), .Z(n765) );
  AND U998 ( .A(n766), .B(n765), .Z(n829) );
  NANDN U999 ( .A(n768), .B(n767), .Z(n772) );
  OR U1000 ( .A(n770), .B(n769), .Z(n771) );
  NAND U1001 ( .A(n772), .B(n771), .Z(n830) );
  XNOR U1002 ( .A(n829), .B(n830), .Z(n831) );
  XNOR U1003 ( .A(n832), .B(n831), .Z(n837) );
  XNOR U1004 ( .A(n838), .B(n837), .Z(o[12]) );
  NANDN U1005 ( .A(n778), .B(n777), .Z(n782) );
  NAND U1006 ( .A(n780), .B(n779), .Z(n781) );
  NAND U1007 ( .A(n782), .B(n781), .Z(n842) );
  XNOR U1008 ( .A(n841), .B(n842), .Z(n844) );
  NAND U1009 ( .A(n784), .B(n783), .Z(n788) );
  NAND U1010 ( .A(n786), .B(n785), .Z(n787) );
  AND U1011 ( .A(n788), .B(n787), .Z(n851) );
  NAND U1012 ( .A(n790), .B(n789), .Z(n794) );
  NAND U1013 ( .A(n792), .B(n791), .Z(n793) );
  AND U1014 ( .A(n794), .B(n793), .Z(n852) );
  AND U1015 ( .A(x[20]), .B(y[59]), .Z(n1020) );
  NAND U1016 ( .A(n1020), .B(n795), .Z(n799) );
  NAND U1017 ( .A(n797), .B(n796), .Z(n798) );
  NAND U1018 ( .A(n799), .B(n798), .Z(n882) );
  NANDN U1019 ( .A(n801), .B(n800), .Z(n804) );
  NANDN U1020 ( .A(n802), .B(n857), .Z(n803) );
  AND U1021 ( .A(n804), .B(n803), .Z(n888) );
  AND U1022 ( .A(y[33]), .B(x[12]), .Z(n806) );
  NAND U1023 ( .A(y[32]), .B(x[13]), .Z(n805) );
  XNOR U1024 ( .A(n806), .B(n805), .Z(n905) );
  NAND U1025 ( .A(x[1]), .B(y[12]), .Z(n904) );
  XNOR U1026 ( .A(n905), .B(n904), .Z(n887) );
  AND U1027 ( .A(x[18]), .B(y[59]), .Z(n896) );
  NAND U1028 ( .A(x[21]), .B(y[56]), .Z(n895) );
  XNOR U1029 ( .A(n896), .B(n895), .Z(n898) );
  AND U1030 ( .A(y[58]), .B(x[19]), .Z(n826) );
  NAND U1031 ( .A(y[57]), .B(x[20]), .Z(n807) );
  XNOR U1032 ( .A(n826), .B(n807), .Z(n897) );
  XNOR U1033 ( .A(n898), .B(n897), .Z(n886) );
  XNOR U1034 ( .A(n887), .B(n886), .Z(n889) );
  XNOR U1035 ( .A(n888), .B(n889), .Z(n881) );
  NAND U1036 ( .A(n809), .B(n808), .Z(n813) );
  AND U1037 ( .A(n811), .B(n810), .Z(n812) );
  ANDN U1038 ( .B(n813), .A(n812), .Z(n880) );
  XOR U1039 ( .A(n881), .B(n880), .Z(n883) );
  XNOR U1040 ( .A(n882), .B(n883), .Z(n847) );
  AND U1041 ( .A(x[10]), .B(y[35]), .Z(n861) );
  NAND U1042 ( .A(n861), .B(n814), .Z(n818) );
  NANDN U1043 ( .A(n816), .B(n815), .Z(n817) );
  NAND U1044 ( .A(n818), .B(n817), .Z(n879) );
  NAND U1045 ( .A(x[5]), .B(y[8]), .Z(n860) );
  XNOR U1046 ( .A(n861), .B(n860), .Z(n863) );
  NAND U1047 ( .A(x[4]), .B(y[9]), .Z(n862) );
  XNOR U1048 ( .A(n863), .B(n862), .Z(n877) );
  AND U1049 ( .A(x[9]), .B(y[36]), .Z(n1019) );
  AND U1050 ( .A(x[0]), .B(y[13]), .Z(n866) );
  AND U1051 ( .A(x[8]), .B(y[37]), .Z(n865) );
  XNOR U1052 ( .A(n866), .B(n865), .Z(n867) );
  XNOR U1053 ( .A(n1019), .B(n867), .Z(n876) );
  XNOR U1054 ( .A(n877), .B(n876), .Z(n878) );
  XOR U1055 ( .A(n879), .B(n878), .Z(n846) );
  AND U1056 ( .A(n903), .B(n819), .Z(n823) );
  NANDN U1057 ( .A(n821), .B(n820), .Z(n822) );
  NANDN U1058 ( .A(n823), .B(n822), .Z(n872) );
  AND U1059 ( .A(y[61]), .B(x[16]), .Z(n825) );
  NAND U1060 ( .A(y[60]), .B(x[17]), .Z(n824) );
  XNOR U1061 ( .A(n825), .B(n824), .Z(n859) );
  AND U1062 ( .A(x[18]), .B(y[57]), .Z(n827) );
  NAND U1063 ( .A(n827), .B(n826), .Z(n858) );
  XNOR U1064 ( .A(n859), .B(n858), .Z(n871) );
  AND U1065 ( .A(x[3]), .B(y[10]), .Z(n1001) );
  XNOR U1066 ( .A(n1001), .B(n828), .Z(n892) );
  NAND U1067 ( .A(x[2]), .B(y[11]), .Z(n891) );
  XNOR U1068 ( .A(n892), .B(n891), .Z(n870) );
  XNOR U1069 ( .A(n871), .B(n870), .Z(n873) );
  XOR U1070 ( .A(n872), .B(n873), .Z(n845) );
  XOR U1071 ( .A(n846), .B(n845), .Z(n848) );
  XOR U1072 ( .A(n847), .B(n848), .Z(n853) );
  XNOR U1073 ( .A(n854), .B(n853), .Z(n843) );
  XNOR U1074 ( .A(n844), .B(n843), .Z(n912) );
  NANDN U1075 ( .A(n830), .B(n829), .Z(n834) );
  NANDN U1076 ( .A(n832), .B(n831), .Z(n833) );
  AND U1077 ( .A(n834), .B(n833), .Z(n910) );
  NANDN U1078 ( .A(n836), .B(n835), .Z(n840) );
  NAND U1079 ( .A(n838), .B(n837), .Z(n839) );
  NAND U1080 ( .A(n840), .B(n839), .Z(n909) );
  XNOR U1081 ( .A(n910), .B(n909), .Z(n911) );
  XNOR U1082 ( .A(n912), .B(n911), .Z(o[13]) );
  NAND U1083 ( .A(n846), .B(n845), .Z(n850) );
  NAND U1084 ( .A(n848), .B(n847), .Z(n849) );
  NAND U1085 ( .A(n850), .B(n849), .Z(n1062) );
  NAND U1086 ( .A(n852), .B(n851), .Z(n856) );
  NAND U1087 ( .A(n854), .B(n853), .Z(n855) );
  NAND U1088 ( .A(n856), .B(n855), .Z(n1061) );
  AND U1089 ( .A(x[17]), .B(y[61]), .Z(n950) );
  IV U1090 ( .A(n860), .Z(n1007) );
  AND U1091 ( .A(x[13]), .B(y[33]), .Z(n991) );
  AND U1092 ( .A(x[14]), .B(y[32]), .Z(n993) );
  AND U1093 ( .A(x[0]), .B(y[14]), .Z(n992) );
  XOR U1094 ( .A(n993), .B(n992), .Z(n990) );
  XNOR U1095 ( .A(n991), .B(n990), .Z(n922) );
  AND U1096 ( .A(x[20]), .B(y[58]), .Z(n899) );
  NAND U1097 ( .A(y[57]), .B(x[21]), .Z(n864) );
  XNOR U1098 ( .A(n899), .B(n864), .Z(n946) );
  AND U1099 ( .A(x[22]), .B(y[56]), .Z(n945) );
  XOR U1100 ( .A(n946), .B(n945), .Z(n944) );
  XNOR U1101 ( .A(n944), .B(n943), .Z(n921) );
  XOR U1102 ( .A(n920), .B(n919), .Z(n917) );
  XOR U1103 ( .A(n918), .B(n917), .Z(n916) );
  AND U1104 ( .A(y[8]), .B(x[6]), .Z(n869) );
  NAND U1105 ( .A(y[9]), .B(x[5]), .Z(n868) );
  XNOR U1106 ( .A(n869), .B(n868), .Z(n1005) );
  AND U1107 ( .A(x[11]), .B(y[35]), .Z(n1004) );
  XNOR U1108 ( .A(n1005), .B(n1004), .Z(n938) );
  AND U1109 ( .A(x[1]), .B(y[13]), .Z(n985) );
  AND U1110 ( .A(x[16]), .B(y[62]), .Z(n987) );
  AND U1111 ( .A(x[8]), .B(y[38]), .Z(n986) );
  XOR U1112 ( .A(n987), .B(n986), .Z(n984) );
  XNOR U1113 ( .A(n985), .B(n984), .Z(n937) );
  XNOR U1114 ( .A(n936), .B(n935), .Z(n915) );
  XNOR U1115 ( .A(n916), .B(n915), .Z(n1040) );
  NAND U1116 ( .A(n871), .B(n870), .Z(n875) );
  NANDN U1117 ( .A(n873), .B(n872), .Z(n874) );
  NAND U1118 ( .A(n875), .B(n874), .Z(n1042) );
  XOR U1119 ( .A(n1042), .B(n1041), .Z(n1039) );
  XOR U1120 ( .A(n1040), .B(n1039), .Z(n1053) );
  NAND U1121 ( .A(n881), .B(n880), .Z(n885) );
  NAND U1122 ( .A(n883), .B(n882), .Z(n884) );
  AND U1123 ( .A(n885), .B(n884), .Z(n1056) );
  AND U1124 ( .A(y[36]), .B(x[10]), .Z(n894) );
  NAND U1125 ( .A(y[37]), .B(x[9]), .Z(n893) );
  XNOR U1126 ( .A(n894), .B(n893), .Z(n1017) );
  AND U1127 ( .A(x[2]), .B(y[12]), .Z(n1016) );
  XNOR U1128 ( .A(n1017), .B(n1016), .Z(n926) );
  XOR U1129 ( .A(n924), .B(n923), .Z(n1035) );
  XOR U1130 ( .A(n1036), .B(n1035), .Z(n1034) );
  AND U1131 ( .A(n900), .B(n899), .Z(n952) );
  AND U1132 ( .A(x[18]), .B(y[60]), .Z(n951) );
  XOR U1133 ( .A(n952), .B(n951), .Z(n949) );
  XOR U1134 ( .A(n950), .B(n949), .Z(n930) );
  AND U1135 ( .A(y[11]), .B(x[3]), .Z(n902) );
  NAND U1136 ( .A(y[10]), .B(x[4]), .Z(n901) );
  XNOR U1137 ( .A(n902), .B(n901), .Z(n999) );
  AND U1138 ( .A(x[12]), .B(y[34]), .Z(n998) );
  XNOR U1139 ( .A(n999), .B(n998), .Z(n932) );
  NAND U1140 ( .A(n903), .B(n991), .Z(n908) );
  IV U1141 ( .A(n904), .Z(n906) );
  NAND U1142 ( .A(n906), .B(n905), .Z(n907) );
  AND U1143 ( .A(n908), .B(n907), .Z(n931) );
  XNOR U1144 ( .A(n930), .B(n929), .Z(n1033) );
  XOR U1145 ( .A(n1034), .B(n1033), .Z(n1055) );
  XOR U1146 ( .A(n1056), .B(n1055), .Z(n1054) );
  XOR U1147 ( .A(n1053), .B(n1054), .Z(n1059) );
  XOR U1148 ( .A(n1060), .B(n1059), .Z(n1049) );
  NANDN U1149 ( .A(n910), .B(n909), .Z(n914) );
  NAND U1150 ( .A(n912), .B(n911), .Z(n913) );
  NAND U1151 ( .A(n914), .B(n913), .Z(n1047) );
  XNOR U1152 ( .A(n1048), .B(n1047), .Z(o[14]) );
  NAND U1153 ( .A(n924), .B(n923), .Z(n928) );
  NAND U1154 ( .A(n926), .B(n925), .Z(n927) );
  AND U1155 ( .A(n928), .B(n927), .Z(n1032) );
  NANDN U1156 ( .A(n930), .B(n929), .Z(n934) );
  NAND U1157 ( .A(n932), .B(n931), .Z(n933) );
  AND U1158 ( .A(n934), .B(n933), .Z(n942) );
  NAND U1159 ( .A(n936), .B(n935), .Z(n940) );
  NAND U1160 ( .A(n938), .B(n937), .Z(n939) );
  NAND U1161 ( .A(n940), .B(n939), .Z(n941) );
  XNOR U1162 ( .A(n942), .B(n941), .Z(n1030) );
  NAND U1163 ( .A(n944), .B(n943), .Z(n948) );
  NAND U1164 ( .A(n946), .B(n945), .Z(n947) );
  AND U1165 ( .A(n948), .B(n947), .Z(n1028) );
  NAND U1166 ( .A(n950), .B(n949), .Z(n954) );
  NAND U1167 ( .A(n952), .B(n951), .Z(n953) );
  AND U1168 ( .A(n954), .B(n953), .Z(n983) );
  AND U1169 ( .A(y[39]), .B(x[8]), .Z(n956) );
  NAND U1170 ( .A(y[14]), .B(x[1]), .Z(n955) );
  XNOR U1171 ( .A(n956), .B(n955), .Z(n963) );
  AND U1172 ( .A(y[60]), .B(x[19]), .Z(n961) );
  AND U1173 ( .A(x[4]), .B(y[11]), .Z(n1000) );
  AND U1174 ( .A(y[12]), .B(x[3]), .Z(n958) );
  NAND U1175 ( .A(y[63]), .B(x[16]), .Z(n957) );
  XNOR U1176 ( .A(n958), .B(n957), .Z(n959) );
  XNOR U1177 ( .A(n1000), .B(n959), .Z(n960) );
  XNOR U1178 ( .A(n961), .B(n960), .Z(n962) );
  XOR U1179 ( .A(n963), .B(n962), .Z(n965) );
  AND U1180 ( .A(x[6]), .B(y[9]), .Z(n1006) );
  AND U1181 ( .A(x[10]), .B(y[37]), .Z(n1018) );
  XNOR U1182 ( .A(n1006), .B(n1018), .Z(n964) );
  XNOR U1183 ( .A(n965), .B(n964), .Z(n981) );
  AND U1184 ( .A(y[56]), .B(x[23]), .Z(n967) );
  NAND U1185 ( .A(y[38]), .B(x[9]), .Z(n966) );
  XNOR U1186 ( .A(n967), .B(n966), .Z(n971) );
  AND U1187 ( .A(y[36]), .B(x[11]), .Z(n969) );
  NAND U1188 ( .A(y[35]), .B(x[12]), .Z(n968) );
  XNOR U1189 ( .A(n969), .B(n968), .Z(n970) );
  XOR U1190 ( .A(n971), .B(n970), .Z(n979) );
  AND U1191 ( .A(y[33]), .B(x[14]), .Z(n973) );
  NAND U1192 ( .A(y[62]), .B(x[17]), .Z(n972) );
  XNOR U1193 ( .A(n973), .B(n972), .Z(n977) );
  AND U1194 ( .A(y[13]), .B(x[2]), .Z(n975) );
  NAND U1195 ( .A(y[34]), .B(x[13]), .Z(n974) );
  XNOR U1196 ( .A(n975), .B(n974), .Z(n976) );
  XNOR U1197 ( .A(n977), .B(n976), .Z(n978) );
  XNOR U1198 ( .A(n979), .B(n978), .Z(n980) );
  XNOR U1199 ( .A(n981), .B(n980), .Z(n982) );
  XNOR U1200 ( .A(n983), .B(n982), .Z(n1026) );
  NAND U1201 ( .A(n985), .B(n984), .Z(n989) );
  NAND U1202 ( .A(n987), .B(n986), .Z(n988) );
  AND U1203 ( .A(n989), .B(n988), .Z(n997) );
  NAND U1204 ( .A(n991), .B(n990), .Z(n995) );
  NAND U1205 ( .A(n993), .B(n992), .Z(n994) );
  NAND U1206 ( .A(n995), .B(n994), .Z(n996) );
  XNOR U1207 ( .A(n997), .B(n996), .Z(n1013) );
  NAND U1208 ( .A(n999), .B(n998), .Z(n1003) );
  NAND U1209 ( .A(n1001), .B(n1000), .Z(n1002) );
  AND U1210 ( .A(n1003), .B(n1002), .Z(n1011) );
  NAND U1211 ( .A(n1005), .B(n1004), .Z(n1009) );
  NAND U1212 ( .A(n1007), .B(n1006), .Z(n1008) );
  NAND U1213 ( .A(n1009), .B(n1008), .Z(n1010) );
  XNOR U1214 ( .A(n1011), .B(n1010), .Z(n1012) );
  XOR U1215 ( .A(n1013), .B(n1012), .Z(n1024) );
  AND U1216 ( .A(y[8]), .B(x[7]), .Z(n1015) );
  NAND U1217 ( .A(y[15]), .B(x[0]), .Z(n1014) );
  XNOR U1218 ( .A(n1015), .B(n1014), .Z(n1022) );
  XNOR U1219 ( .A(n1022), .B(n1021), .Z(n1023) );
  XNOR U1220 ( .A(n1024), .B(n1023), .Z(n1025) );
  XNOR U1221 ( .A(n1026), .B(n1025), .Z(n1027) );
  XNOR U1222 ( .A(n1028), .B(n1027), .Z(n1029) );
  XNOR U1223 ( .A(n1030), .B(n1029), .Z(n1031) );
  NAND U1224 ( .A(n1034), .B(n1033), .Z(n1038) );
  NAND U1225 ( .A(n1036), .B(n1035), .Z(n1037) );
  AND U1226 ( .A(n1038), .B(n1037), .Z(n1046) );
  NANDN U1227 ( .A(n1040), .B(n1039), .Z(n1044) );
  NAND U1228 ( .A(n1042), .B(n1041), .Z(n1043) );
  NAND U1229 ( .A(n1044), .B(n1043), .Z(n1045) );
  NAND U1230 ( .A(n1048), .B(n1047), .Z(n1052) );
  NAND U1231 ( .A(n1050), .B(n1049), .Z(n1051) );
  NAND U1232 ( .A(n1054), .B(n1053), .Z(n1058) );
  NAND U1233 ( .A(n1056), .B(n1055), .Z(n1057) );
  AND U1234 ( .A(x[8]), .B(y[40]), .Z(n1064) );
  NAND U1235 ( .A(x[0]), .B(y[16]), .Z(n1063) );
  XNOR U1236 ( .A(n1064), .B(n1063), .Z(n1065) );
  NAND U1237 ( .A(x[16]), .B(y[64]), .Z(n1155) );
  XNOR U1238 ( .A(n1065), .B(n1155), .Z(o[16]) );
  AND U1239 ( .A(x[0]), .B(y[17]), .Z(n1104) );
  AND U1240 ( .A(x[16]), .B(y[65]), .Z(n1111) );
  AND U1241 ( .A(x[1]), .B(y[16]), .Z(n1080) );
  XOR U1242 ( .A(n1111), .B(n1080), .Z(n1081) );
  XOR U1243 ( .A(n1104), .B(n1081), .Z(n1068) );
  NANDN U1244 ( .A(n1064), .B(n1063), .Z(n1067) );
  NAND U1245 ( .A(n1155), .B(n1065), .Z(n1066) );
  NAND U1246 ( .A(n1067), .B(n1066), .Z(n1069) );
  XNOR U1247 ( .A(n1068), .B(n1069), .Z(n1071) );
  AND U1248 ( .A(x[9]), .B(y[40]), .Z(n1142) );
  AND U1249 ( .A(x[17]), .B(y[64]), .Z(n1197) );
  AND U1250 ( .A(x[8]), .B(y[41]), .Z(n1076) );
  XOR U1251 ( .A(n1197), .B(n1076), .Z(n1077) );
  XOR U1252 ( .A(n1142), .B(n1077), .Z(n1070) );
  XOR U1253 ( .A(n1071), .B(n1070), .Z(o[17]) );
  NANDN U1254 ( .A(n1069), .B(n1068), .Z(n1073) );
  NAND U1255 ( .A(n1071), .B(n1070), .Z(n1072) );
  AND U1256 ( .A(n1073), .B(n1072), .Z(n1092) );
  AND U1257 ( .A(y[18]), .B(x[0]), .Z(n1075) );
  NAND U1258 ( .A(y[17]), .B(x[1]), .Z(n1074) );
  XNOR U1259 ( .A(n1075), .B(n1074), .Z(n1106) );
  AND U1260 ( .A(x[10]), .B(y[40]), .Z(n1105) );
  XOR U1261 ( .A(n1106), .B(n1105), .Z(n1119) );
  AND U1262 ( .A(x[8]), .B(y[42]), .Z(n1117) );
  NAND U1263 ( .A(x[9]), .B(y[41]), .Z(n1116) );
  XNOR U1264 ( .A(n1117), .B(n1116), .Z(n1118) );
  XOR U1265 ( .A(n1119), .B(n1118), .Z(n1093) );
  XNOR U1266 ( .A(n1092), .B(n1093), .Z(n1095) );
  NAND U1267 ( .A(n1197), .B(n1076), .Z(n1079) );
  NAND U1268 ( .A(n1142), .B(n1077), .Z(n1078) );
  NAND U1269 ( .A(n1079), .B(n1078), .Z(n1088) );
  NAND U1270 ( .A(n1111), .B(n1080), .Z(n1083) );
  NAND U1271 ( .A(n1104), .B(n1081), .Z(n1082) );
  NAND U1272 ( .A(n1083), .B(n1082), .Z(n1086) );
  AND U1273 ( .A(x[2]), .B(y[16]), .Z(n1132) );
  NAND U1274 ( .A(x[18]), .B(y[64]), .Z(n1098) );
  XNOR U1275 ( .A(n1132), .B(n1098), .Z(n1100) );
  AND U1276 ( .A(y[66]), .B(x[16]), .Z(n1085) );
  NAND U1277 ( .A(y[65]), .B(x[17]), .Z(n1084) );
  XNOR U1278 ( .A(n1085), .B(n1084), .Z(n1099) );
  XOR U1279 ( .A(n1100), .B(n1099), .Z(n1087) );
  XNOR U1280 ( .A(n1086), .B(n1087), .Z(n1089) );
  XOR U1281 ( .A(n1088), .B(n1089), .Z(n1094) );
  XNOR U1282 ( .A(n1095), .B(n1094), .Z(o[18]) );
  NAND U1283 ( .A(n1087), .B(n1086), .Z(n1091) );
  NANDN U1284 ( .A(n1089), .B(n1088), .Z(n1090) );
  AND U1285 ( .A(n1091), .B(n1090), .Z(n1123) );
  NANDN U1286 ( .A(n1093), .B(n1092), .Z(n1097) );
  NAND U1287 ( .A(n1095), .B(n1094), .Z(n1096) );
  AND U1288 ( .A(n1097), .B(n1096), .Z(n1122) );
  XNOR U1289 ( .A(n1123), .B(n1122), .Z(n1125) );
  NANDN U1290 ( .A(n1098), .B(n1132), .Z(n1102) );
  NAND U1291 ( .A(n1100), .B(n1099), .Z(n1101) );
  NAND U1292 ( .A(n1102), .B(n1101), .Z(n1162) );
  AND U1293 ( .A(x[8]), .B(y[43]), .Z(n1149) );
  AND U1294 ( .A(x[1]), .B(y[18]), .Z(n1150) );
  AND U1295 ( .A(x[0]), .B(y[19]), .Z(n1152) );
  AND U1296 ( .A(y[42]), .B(x[9]), .Z(n1215) );
  NAND U1297 ( .A(y[40]), .B(x[11]), .Z(n1103) );
  XNOR U1298 ( .A(n1215), .B(n1103), .Z(n1144) );
  AND U1299 ( .A(x[10]), .B(y[41]), .Z(n1143) );
  XOR U1300 ( .A(n1144), .B(n1143), .Z(n1160) );
  XOR U1301 ( .A(n1161), .B(n1160), .Z(n1163) );
  XOR U1302 ( .A(n1162), .B(n1163), .Z(n1129) );
  NAND U1303 ( .A(n1150), .B(n1104), .Z(n1108) );
  NAND U1304 ( .A(n1106), .B(n1105), .Z(n1107) );
  NAND U1305 ( .A(n1108), .B(n1107), .Z(n1168) );
  AND U1306 ( .A(y[17]), .B(x[2]), .Z(n1110) );
  NAND U1307 ( .A(y[16]), .B(x[3]), .Z(n1109) );
  XNOR U1308 ( .A(n1110), .B(n1109), .Z(n1133) );
  AND U1309 ( .A(y[66]), .B(x[17]), .Z(n1115) );
  AND U1310 ( .A(n1111), .B(n1115), .Z(n1134) );
  AND U1311 ( .A(y[67]), .B(x[16]), .Z(n1113) );
  NAND U1312 ( .A(y[64]), .B(x[19]), .Z(n1112) );
  XNOR U1313 ( .A(n1113), .B(n1112), .Z(n1157) );
  NAND U1314 ( .A(y[65]), .B(x[18]), .Z(n1114) );
  XNOR U1315 ( .A(n1115), .B(n1114), .Z(n1156) );
  XOR U1316 ( .A(n1157), .B(n1156), .Z(n1166) );
  XOR U1317 ( .A(n1167), .B(n1166), .Z(n1169) );
  XNOR U1318 ( .A(n1168), .B(n1169), .Z(n1128) );
  XNOR U1319 ( .A(n1129), .B(n1128), .Z(n1130) );
  NANDN U1320 ( .A(n1117), .B(n1116), .Z(n1121) );
  NANDN U1321 ( .A(n1119), .B(n1118), .Z(n1120) );
  NAND U1322 ( .A(n1121), .B(n1120), .Z(n1131) );
  XNOR U1323 ( .A(n1130), .B(n1131), .Z(n1124) );
  XOR U1324 ( .A(n1125), .B(n1124), .Z(o[19]) );
  NANDN U1325 ( .A(n1123), .B(n1122), .Z(n1127) );
  NAND U1326 ( .A(n1125), .B(n1124), .Z(n1126) );
  NAND U1327 ( .A(n1127), .B(n1126), .Z(n1236) );
  NAND U1328 ( .A(x[3]), .B(y[17]), .Z(n1212) );
  NANDN U1329 ( .A(n1212), .B(n1132), .Z(n1136) );
  NAND U1330 ( .A(n1134), .B(n1133), .Z(n1135) );
  NAND U1331 ( .A(n1136), .B(n1135), .Z(n1188) );
  AND U1332 ( .A(y[42]), .B(x[10]), .Z(n1138) );
  NAND U1333 ( .A(y[43]), .B(x[9]), .Z(n1137) );
  XNOR U1334 ( .A(n1138), .B(n1137), .Z(n1216) );
  NAND U1335 ( .A(x[11]), .B(y[41]), .Z(n1217) );
  XNOR U1336 ( .A(n1216), .B(n1217), .Z(n1186) );
  AND U1337 ( .A(y[67]), .B(x[17]), .Z(n1140) );
  NAND U1338 ( .A(y[64]), .B(x[20]), .Z(n1139) );
  XNOR U1339 ( .A(n1140), .B(n1139), .Z(n1198) );
  AND U1340 ( .A(y[65]), .B(x[19]), .Z(n1251) );
  NAND U1341 ( .A(y[66]), .B(x[18]), .Z(n1141) );
  XNOR U1342 ( .A(n1251), .B(n1141), .Z(n1199) );
  XOR U1343 ( .A(n1186), .B(n1185), .Z(n1187) );
  AND U1344 ( .A(x[11]), .B(y[42]), .Z(n1256) );
  NAND U1345 ( .A(n1256), .B(n1142), .Z(n1146) );
  NAND U1346 ( .A(n1144), .B(n1143), .Z(n1145) );
  NAND U1347 ( .A(n1146), .B(n1145), .Z(n1194) );
  AND U1348 ( .A(x[4]), .B(y[16]), .Z(n1202) );
  AND U1349 ( .A(x[17]), .B(y[65]), .Z(n1148) );
  AND U1350 ( .A(x[18]), .B(y[66]), .Z(n1147) );
  NAND U1351 ( .A(n1148), .B(n1147), .Z(n1203) );
  XNOR U1352 ( .A(n1202), .B(n1203), .Z(n1204) );
  NAND U1353 ( .A(x[16]), .B(y[68]), .Z(n1282) );
  XNOR U1354 ( .A(n1204), .B(n1282), .Z(n1191) );
  AND U1355 ( .A(x[12]), .B(y[40]), .Z(n1246) );
  AND U1356 ( .A(x[8]), .B(y[44]), .Z(n1220) );
  XOR U1357 ( .A(n1246), .B(n1220), .Z(n1222) );
  NAND U1358 ( .A(x[1]), .B(y[19]), .Z(n1221) );
  XNOR U1359 ( .A(n1222), .B(n1221), .Z(n1192) );
  XOR U1360 ( .A(n1174), .B(n1173), .Z(n1176) );
  NAND U1361 ( .A(n1150), .B(n1149), .Z(n1154) );
  NAND U1362 ( .A(n1152), .B(n1151), .Z(n1153) );
  NAND U1363 ( .A(n1154), .B(n1153), .Z(n1181) );
  NAND U1364 ( .A(x[2]), .B(y[18]), .Z(n1210) );
  NAND U1365 ( .A(x[0]), .B(y[20]), .Z(n1211) );
  XOR U1366 ( .A(n1212), .B(n1211), .Z(n1209) );
  AND U1367 ( .A(x[19]), .B(y[67]), .Z(n1357) );
  NANDN U1368 ( .A(n1155), .B(n1357), .Z(n1159) );
  NAND U1369 ( .A(n1157), .B(n1156), .Z(n1158) );
  NAND U1370 ( .A(n1159), .B(n1158), .Z(n1179) );
  XOR U1371 ( .A(n1181), .B(n1182), .Z(n1175) );
  XOR U1372 ( .A(n1176), .B(n1175), .Z(n1232) );
  NAND U1373 ( .A(n1161), .B(n1160), .Z(n1165) );
  NAND U1374 ( .A(n1163), .B(n1162), .Z(n1164) );
  AND U1375 ( .A(n1165), .B(n1164), .Z(n1230) );
  NAND U1376 ( .A(n1167), .B(n1166), .Z(n1171) );
  NAND U1377 ( .A(n1169), .B(n1168), .Z(n1170) );
  AND U1378 ( .A(n1171), .B(n1170), .Z(n1229) );
  XOR U1379 ( .A(n1230), .B(n1229), .Z(n1231) );
  XNOR U1380 ( .A(n1232), .B(n1231), .Z(n1237) );
  XNOR U1381 ( .A(n1235), .B(n1237), .Z(n1172) );
  XNOR U1382 ( .A(n1236), .B(n1172), .Z(o[20]) );
  NAND U1383 ( .A(n1174), .B(n1173), .Z(n1178) );
  NAND U1384 ( .A(n1176), .B(n1175), .Z(n1177) );
  AND U1385 ( .A(n1178), .B(n1177), .Z(n1318) );
  NAND U1386 ( .A(n1180), .B(n1179), .Z(n1184) );
  NAND U1387 ( .A(n1182), .B(n1181), .Z(n1183) );
  AND U1388 ( .A(n1184), .B(n1183), .Z(n1319) );
  NAND U1389 ( .A(n1186), .B(n1185), .Z(n1190) );
  NAND U1390 ( .A(n1188), .B(n1187), .Z(n1189) );
  AND U1391 ( .A(n1190), .B(n1189), .Z(n1312) );
  NAND U1392 ( .A(n1192), .B(n1191), .Z(n1196) );
  NAND U1393 ( .A(n1194), .B(n1193), .Z(n1195) );
  AND U1394 ( .A(n1196), .B(n1195), .Z(n1313) );
  AND U1395 ( .A(x[20]), .B(y[67]), .Z(n1377) );
  NAND U1396 ( .A(n1377), .B(n1197), .Z(n1201) );
  NAND U1397 ( .A(n1199), .B(n1198), .Z(n1200) );
  NAND U1398 ( .A(n1201), .B(n1200), .Z(n1272) );
  NANDN U1399 ( .A(n1203), .B(n1202), .Z(n1206) );
  NANDN U1400 ( .A(n1282), .B(n1204), .Z(n1205) );
  AND U1401 ( .A(n1206), .B(n1205), .Z(n1255) );
  AND U1402 ( .A(y[41]), .B(x[12]), .Z(n1208) );
  NAND U1403 ( .A(y[40]), .B(x[13]), .Z(n1207) );
  XNOR U1404 ( .A(n1208), .B(n1207), .Z(n1247) );
  NAND U1405 ( .A(x[1]), .B(y[20]), .Z(n1248) );
  XNOR U1406 ( .A(n1247), .B(n1248), .Z(n1253) );
  AND U1407 ( .A(x[18]), .B(y[67]), .Z(n1264) );
  AND U1408 ( .A(x[21]), .B(y[64]), .Z(n1263) );
  XOR U1409 ( .A(n1264), .B(n1263), .Z(n1266) );
  AND U1410 ( .A(x[19]), .B(y[66]), .Z(n1226) );
  AND U1411 ( .A(x[20]), .B(y[65]), .Z(n1430) );
  XOR U1412 ( .A(n1226), .B(n1430), .Z(n1265) );
  XNOR U1413 ( .A(n1266), .B(n1265), .Z(n1252) );
  XNOR U1414 ( .A(n1253), .B(n1252), .Z(n1254) );
  XNOR U1415 ( .A(n1255), .B(n1254), .Z(n1269) );
  NAND U1416 ( .A(n1210), .B(n1209), .Z(n1214) );
  AND U1417 ( .A(n1212), .B(n1211), .Z(n1213) );
  ANDN U1418 ( .B(n1214), .A(n1213), .Z(n1270) );
  AND U1419 ( .A(x[10]), .B(y[43]), .Z(n1287) );
  NAND U1420 ( .A(n1287), .B(n1215), .Z(n1219) );
  NANDN U1421 ( .A(n1217), .B(n1216), .Z(n1218) );
  AND U1422 ( .A(n1219), .B(n1218), .Z(n1296) );
  AND U1423 ( .A(x[9]), .B(y[44]), .Z(n1406) );
  AND U1424 ( .A(x[0]), .B(y[21]), .Z(n1275) );
  NAND U1425 ( .A(x[8]), .B(y[45]), .Z(n1276) );
  XOR U1426 ( .A(n1275), .B(n1276), .Z(n1277) );
  XNOR U1427 ( .A(n1406), .B(n1277), .Z(n1294) );
  AND U1428 ( .A(x[5]), .B(y[16]), .Z(n1400) );
  NAND U1429 ( .A(x[4]), .B(y[17]), .Z(n1289) );
  XOR U1430 ( .A(n1288), .B(n1289), .Z(n1295) );
  XOR U1431 ( .A(n1294), .B(n1295), .Z(n1297) );
  XNOR U1432 ( .A(n1296), .B(n1297), .Z(n1307) );
  NAND U1433 ( .A(n1246), .B(n1220), .Z(n1224) );
  ANDN U1434 ( .B(n1222), .A(n1221), .Z(n1223) );
  ANDN U1435 ( .B(n1224), .A(n1223), .Z(n1302) );
  AND U1436 ( .A(x[18]), .B(y[65]), .Z(n1225) );
  AND U1437 ( .A(n1226), .B(n1225), .Z(n1283) );
  AND U1438 ( .A(y[69]), .B(x[16]), .Z(n1228) );
  NAND U1439 ( .A(y[68]), .B(x[17]), .Z(n1227) );
  XOR U1440 ( .A(n1228), .B(n1227), .Z(n1284) );
  XNOR U1441 ( .A(n1283), .B(n1284), .Z(n1300) );
  AND U1442 ( .A(x[3]), .B(y[18]), .Z(n1433) );
  NAND U1443 ( .A(x[2]), .B(y[19]), .Z(n1258) );
  XOR U1444 ( .A(n1257), .B(n1258), .Z(n1301) );
  XOR U1445 ( .A(n1300), .B(n1301), .Z(n1303) );
  XNOR U1446 ( .A(n1302), .B(n1303), .Z(n1306) );
  XOR U1447 ( .A(n1308), .B(n1309), .Z(n1314) );
  XOR U1448 ( .A(n1315), .B(n1314), .Z(n1320) );
  XOR U1449 ( .A(n1321), .B(n1320), .Z(n1241) );
  NAND U1450 ( .A(n1230), .B(n1229), .Z(n1234) );
  NANDN U1451 ( .A(n1232), .B(n1231), .Z(n1233) );
  AND U1452 ( .A(n1234), .B(n1233), .Z(n1239) );
  XNOR U1453 ( .A(n1239), .B(n1238), .Z(n1240) );
  XNOR U1454 ( .A(n1241), .B(n1240), .Z(o[21]) );
  NANDN U1455 ( .A(n1239), .B(n1238), .Z(n1243) );
  NAND U1456 ( .A(n1241), .B(n1240), .Z(n1242) );
  AND U1457 ( .A(n1243), .B(n1242), .Z(n1481) );
  AND U1458 ( .A(y[19]), .B(x[3]), .Z(n1245) );
  NAND U1459 ( .A(y[18]), .B(x[4]), .Z(n1244) );
  XNOR U1460 ( .A(n1245), .B(n1244), .Z(n1432) );
  AND U1461 ( .A(x[12]), .B(y[42]), .Z(n1431) );
  XNOR U1462 ( .A(n1432), .B(n1431), .Z(n1351) );
  AND U1463 ( .A(x[13]), .B(y[41]), .Z(n1412) );
  NAND U1464 ( .A(n1246), .B(n1412), .Z(n1250) );
  NANDN U1465 ( .A(n1248), .B(n1247), .Z(n1249) );
  AND U1466 ( .A(n1250), .B(n1249), .Z(n1350) );
  AND U1467 ( .A(x[17]), .B(y[69]), .Z(n1363) );
  AND U1468 ( .A(x[18]), .B(y[68]), .Z(n1365) );
  AND U1469 ( .A(y[66]), .B(x[20]), .Z(n1293) );
  AND U1470 ( .A(n1293), .B(n1251), .Z(n1364) );
  XOR U1471 ( .A(n1365), .B(n1364), .Z(n1362) );
  XNOR U1472 ( .A(n1363), .B(n1362), .Z(n1349) );
  NAND U1473 ( .A(n1256), .B(n1433), .Z(n1260) );
  NANDN U1474 ( .A(n1258), .B(n1257), .Z(n1259) );
  AND U1475 ( .A(n1260), .B(n1259), .Z(n1331) );
  AND U1476 ( .A(y[44]), .B(x[10]), .Z(n1262) );
  NAND U1477 ( .A(y[45]), .B(x[9]), .Z(n1261) );
  XNOR U1478 ( .A(n1262), .B(n1261), .Z(n1405) );
  AND U1479 ( .A(x[2]), .B(y[20]), .Z(n1404) );
  XNOR U1480 ( .A(n1405), .B(n1404), .Z(n1333) );
  NAND U1481 ( .A(n1264), .B(n1263), .Z(n1268) );
  NAND U1482 ( .A(n1266), .B(n1265), .Z(n1267) );
  AND U1483 ( .A(n1268), .B(n1267), .Z(n1332) );
  XOR U1484 ( .A(n1331), .B(n1330), .Z(n1326) );
  XOR U1485 ( .A(n1327), .B(n1326), .Z(n1324) );
  XNOR U1486 ( .A(n1325), .B(n1324), .Z(n1501) );
  NAND U1487 ( .A(n1270), .B(n1269), .Z(n1274) );
  NAND U1488 ( .A(n1272), .B(n1271), .Z(n1273) );
  NAND U1489 ( .A(n1274), .B(n1273), .Z(n1500) );
  NANDN U1490 ( .A(n1276), .B(n1275), .Z(n1279) );
  NANDN U1491 ( .A(n1277), .B(n1406), .Z(n1278) );
  AND U1492 ( .A(n1279), .B(n1278), .Z(n1342) );
  AND U1493 ( .A(y[16]), .B(x[6]), .Z(n1281) );
  NAND U1494 ( .A(y[17]), .B(x[5]), .Z(n1280) );
  XNOR U1495 ( .A(n1281), .B(n1280), .Z(n1399) );
  AND U1496 ( .A(x[11]), .B(y[43]), .Z(n1398) );
  XNOR U1497 ( .A(n1399), .B(n1398), .Z(n1345) );
  AND U1498 ( .A(x[1]), .B(y[21]), .Z(n1418) );
  AND U1499 ( .A(x[16]), .B(y[70]), .Z(n1420) );
  AND U1500 ( .A(x[8]), .B(y[46]), .Z(n1419) );
  XOR U1501 ( .A(n1420), .B(n1419), .Z(n1417) );
  XNOR U1502 ( .A(n1418), .B(n1417), .Z(n1344) );
  XNOR U1503 ( .A(n1342), .B(n1343), .Z(n1469) );
  NANDN U1504 ( .A(n1282), .B(n1363), .Z(n1286) );
  NANDN U1505 ( .A(n1284), .B(n1283), .Z(n1285) );
  AND U1506 ( .A(n1286), .B(n1285), .Z(n1471) );
  NAND U1507 ( .A(n1287), .B(n1400), .Z(n1291) );
  NANDN U1508 ( .A(n1289), .B(n1288), .Z(n1290) );
  AND U1509 ( .A(n1291), .B(n1290), .Z(n1336) );
  AND U1510 ( .A(x[14]), .B(y[40]), .Z(n1414) );
  AND U1511 ( .A(x[0]), .B(y[22]), .Z(n1413) );
  XOR U1512 ( .A(n1414), .B(n1413), .Z(n1411) );
  XNOR U1513 ( .A(n1412), .B(n1411), .Z(n1339) );
  NAND U1514 ( .A(y[65]), .B(x[21]), .Z(n1292) );
  XNOR U1515 ( .A(n1293), .B(n1292), .Z(n1359) );
  AND U1516 ( .A(x[22]), .B(y[64]), .Z(n1358) );
  XOR U1517 ( .A(n1359), .B(n1358), .Z(n1356) );
  XNOR U1518 ( .A(n1357), .B(n1356), .Z(n1338) );
  XNOR U1519 ( .A(n1336), .B(n1337), .Z(n1470) );
  XOR U1520 ( .A(n1471), .B(n1470), .Z(n1468) );
  XOR U1521 ( .A(n1469), .B(n1468), .Z(n1463) );
  NANDN U1522 ( .A(n1295), .B(n1294), .Z(n1299) );
  OR U1523 ( .A(n1297), .B(n1296), .Z(n1298) );
  NAND U1524 ( .A(n1299), .B(n1298), .Z(n1465) );
  NANDN U1525 ( .A(n1301), .B(n1300), .Z(n1305) );
  OR U1526 ( .A(n1303), .B(n1302), .Z(n1304) );
  NAND U1527 ( .A(n1305), .B(n1304), .Z(n1464) );
  XOR U1528 ( .A(n1465), .B(n1464), .Z(n1462) );
  XNOR U1529 ( .A(n1463), .B(n1462), .Z(n1499) );
  XNOR U1530 ( .A(n1498), .B(n1499), .Z(n1486) );
  NAND U1531 ( .A(n1307), .B(n1306), .Z(n1311) );
  NAND U1532 ( .A(n1309), .B(n1308), .Z(n1310) );
  NAND U1533 ( .A(n1311), .B(n1310), .Z(n1489) );
  NAND U1534 ( .A(n1313), .B(n1312), .Z(n1317) );
  NAND U1535 ( .A(n1315), .B(n1314), .Z(n1316) );
  NAND U1536 ( .A(n1317), .B(n1316), .Z(n1488) );
  XOR U1537 ( .A(n1486), .B(n1487), .Z(n1482) );
  NAND U1538 ( .A(n1319), .B(n1318), .Z(n1323) );
  NAND U1539 ( .A(n1321), .B(n1320), .Z(n1322) );
  AND U1540 ( .A(n1323), .B(n1322), .Z(n1483) );
  XOR U1541 ( .A(n1482), .B(n1483), .Z(n1480) );
  XOR U1542 ( .A(n1481), .B(n1480), .Z(o[22]) );
  NAND U1543 ( .A(n1325), .B(n1324), .Z(n1329) );
  NAND U1544 ( .A(n1327), .B(n1326), .Z(n1328) );
  AND U1545 ( .A(n1329), .B(n1328), .Z(n1497) );
  NAND U1546 ( .A(n1331), .B(n1330), .Z(n1335) );
  NAND U1547 ( .A(n1333), .B(n1332), .Z(n1334) );
  AND U1548 ( .A(n1335), .B(n1334), .Z(n1479) );
  NANDN U1549 ( .A(n1337), .B(n1336), .Z(n1341) );
  NAND U1550 ( .A(n1339), .B(n1338), .Z(n1340) );
  AND U1551 ( .A(n1341), .B(n1340), .Z(n1461) );
  NANDN U1552 ( .A(n1343), .B(n1342), .Z(n1347) );
  NAND U1553 ( .A(n1345), .B(n1344), .Z(n1346) );
  AND U1554 ( .A(n1347), .B(n1346), .Z(n1355) );
  NAND U1555 ( .A(n1349), .B(n1348), .Z(n1353) );
  NAND U1556 ( .A(n1351), .B(n1350), .Z(n1352) );
  NAND U1557 ( .A(n1353), .B(n1352), .Z(n1354) );
  XNOR U1558 ( .A(n1355), .B(n1354), .Z(n1459) );
  NAND U1559 ( .A(n1357), .B(n1356), .Z(n1361) );
  NAND U1560 ( .A(n1359), .B(n1358), .Z(n1360) );
  AND U1561 ( .A(n1361), .B(n1360), .Z(n1457) );
  NAND U1562 ( .A(n1363), .B(n1362), .Z(n1367) );
  NAND U1563 ( .A(n1365), .B(n1364), .Z(n1366) );
  AND U1564 ( .A(n1367), .B(n1366), .Z(n1397) );
  AND U1565 ( .A(y[18]), .B(x[5]), .Z(n1369) );
  NAND U1566 ( .A(y[46]), .B(x[9]), .Z(n1368) );
  XNOR U1567 ( .A(n1369), .B(n1368), .Z(n1376) );
  AND U1568 ( .A(y[42]), .B(x[13]), .Z(n1374) );
  AND U1569 ( .A(x[21]), .B(y[66]), .Z(n1429) );
  AND U1570 ( .A(y[23]), .B(x[0]), .Z(n1371) );
  NAND U1571 ( .A(y[21]), .B(x[2]), .Z(n1370) );
  XNOR U1572 ( .A(n1371), .B(n1370), .Z(n1372) );
  XNOR U1573 ( .A(n1429), .B(n1372), .Z(n1373) );
  XNOR U1574 ( .A(n1374), .B(n1373), .Z(n1375) );
  XOR U1575 ( .A(n1376), .B(n1375), .Z(n1379) );
  AND U1576 ( .A(x[6]), .B(y[17]), .Z(n1401) );
  XNOR U1577 ( .A(n1377), .B(n1401), .Z(n1378) );
  XNOR U1578 ( .A(n1379), .B(n1378), .Z(n1395) );
  AND U1579 ( .A(y[65]), .B(x[22]), .Z(n1381) );
  NAND U1580 ( .A(y[44]), .B(x[11]), .Z(n1380) );
  XNOR U1581 ( .A(n1381), .B(n1380), .Z(n1385) );
  AND U1582 ( .A(y[69]), .B(x[18]), .Z(n1383) );
  NAND U1583 ( .A(y[43]), .B(x[12]), .Z(n1382) );
  XNOR U1584 ( .A(n1383), .B(n1382), .Z(n1384) );
  XOR U1585 ( .A(n1385), .B(n1384), .Z(n1393) );
  AND U1586 ( .A(y[70]), .B(x[17]), .Z(n1387) );
  NAND U1587 ( .A(y[68]), .B(x[19]), .Z(n1386) );
  XNOR U1588 ( .A(n1387), .B(n1386), .Z(n1391) );
  AND U1589 ( .A(y[40]), .B(x[15]), .Z(n1389) );
  NAND U1590 ( .A(y[16]), .B(x[7]), .Z(n1388) );
  XNOR U1591 ( .A(n1389), .B(n1388), .Z(n1390) );
  XNOR U1592 ( .A(n1391), .B(n1390), .Z(n1392) );
  XNOR U1593 ( .A(n1393), .B(n1392), .Z(n1394) );
  XNOR U1594 ( .A(n1395), .B(n1394), .Z(n1396) );
  XNOR U1595 ( .A(n1397), .B(n1396), .Z(n1455) );
  NAND U1596 ( .A(n1399), .B(n1398), .Z(n1403) );
  NAND U1597 ( .A(n1401), .B(n1400), .Z(n1402) );
  AND U1598 ( .A(n1403), .B(n1402), .Z(n1410) );
  NAND U1599 ( .A(n1405), .B(n1404), .Z(n1408) );
  AND U1600 ( .A(x[10]), .B(y[45]), .Z(n1446) );
  NAND U1601 ( .A(n1446), .B(n1406), .Z(n1407) );
  NAND U1602 ( .A(n1408), .B(n1407), .Z(n1409) );
  XNOR U1603 ( .A(n1410), .B(n1409), .Z(n1426) );
  NAND U1604 ( .A(n1412), .B(n1411), .Z(n1416) );
  NAND U1605 ( .A(n1414), .B(n1413), .Z(n1415) );
  AND U1606 ( .A(n1416), .B(n1415), .Z(n1424) );
  NAND U1607 ( .A(n1418), .B(n1417), .Z(n1422) );
  NAND U1608 ( .A(n1420), .B(n1419), .Z(n1421) );
  NAND U1609 ( .A(n1422), .B(n1421), .Z(n1423) );
  XNOR U1610 ( .A(n1424), .B(n1423), .Z(n1425) );
  XOR U1611 ( .A(n1426), .B(n1425), .Z(n1453) );
  AND U1612 ( .A(y[20]), .B(x[3]), .Z(n1428) );
  NAND U1613 ( .A(y[22]), .B(x[1]), .Z(n1427) );
  XNOR U1614 ( .A(n1428), .B(n1427), .Z(n1451) );
  AND U1615 ( .A(n1430), .B(n1429), .Z(n1445) );
  NAND U1616 ( .A(n1432), .B(n1431), .Z(n1435) );
  AND U1617 ( .A(x[4]), .B(y[19]), .Z(n1447) );
  NAND U1618 ( .A(n1447), .B(n1433), .Z(n1434) );
  AND U1619 ( .A(n1435), .B(n1434), .Z(n1443) );
  AND U1620 ( .A(y[47]), .B(x[8]), .Z(n1437) );
  NAND U1621 ( .A(y[71]), .B(x[16]), .Z(n1436) );
  XNOR U1622 ( .A(n1437), .B(n1436), .Z(n1441) );
  AND U1623 ( .A(y[64]), .B(x[23]), .Z(n1439) );
  NAND U1624 ( .A(y[41]), .B(x[14]), .Z(n1438) );
  XNOR U1625 ( .A(n1439), .B(n1438), .Z(n1440) );
  XNOR U1626 ( .A(n1441), .B(n1440), .Z(n1442) );
  XNOR U1627 ( .A(n1443), .B(n1442), .Z(n1444) );
  XOR U1628 ( .A(n1445), .B(n1444), .Z(n1449) );
  XNOR U1629 ( .A(n1447), .B(n1446), .Z(n1448) );
  XNOR U1630 ( .A(n1449), .B(n1448), .Z(n1450) );
  XNOR U1631 ( .A(n1451), .B(n1450), .Z(n1452) );
  XNOR U1632 ( .A(n1453), .B(n1452), .Z(n1454) );
  XNOR U1633 ( .A(n1455), .B(n1454), .Z(n1456) );
  XNOR U1634 ( .A(n1457), .B(n1456), .Z(n1458) );
  XNOR U1635 ( .A(n1459), .B(n1458), .Z(n1460) );
  XNOR U1636 ( .A(n1461), .B(n1460), .Z(n1477) );
  NANDN U1637 ( .A(n1463), .B(n1462), .Z(n1467) );
  NAND U1638 ( .A(n1465), .B(n1464), .Z(n1466) );
  AND U1639 ( .A(n1467), .B(n1466), .Z(n1475) );
  NAND U1640 ( .A(n1469), .B(n1468), .Z(n1473) );
  NAND U1641 ( .A(n1471), .B(n1470), .Z(n1472) );
  NAND U1642 ( .A(n1473), .B(n1472), .Z(n1474) );
  XNOR U1643 ( .A(n1475), .B(n1474), .Z(n1476) );
  XNOR U1644 ( .A(n1477), .B(n1476), .Z(n1478) );
  XNOR U1645 ( .A(n1479), .B(n1478), .Z(n1495) );
  NAND U1646 ( .A(n1481), .B(n1480), .Z(n1485) );
  NAND U1647 ( .A(n1483), .B(n1482), .Z(n1484) );
  AND U1648 ( .A(n1485), .B(n1484), .Z(n1493) );
  NANDN U1649 ( .A(n1487), .B(n1486), .Z(n1491) );
  NAND U1650 ( .A(n1489), .B(n1488), .Z(n1490) );
  NAND U1651 ( .A(n1491), .B(n1490), .Z(n1492) );
  XNOR U1652 ( .A(n1493), .B(n1492), .Z(n1494) );
  XNOR U1653 ( .A(n1495), .B(n1494), .Z(n1496) );
  XNOR U1654 ( .A(n1497), .B(n1496), .Z(n1505) );
  NAND U1655 ( .A(n1499), .B(n1498), .Z(n1503) );
  NAND U1656 ( .A(n1501), .B(n1500), .Z(n1502) );
  NAND U1657 ( .A(n1503), .B(n1502), .Z(n1504) );
  XNOR U1658 ( .A(n1505), .B(n1504), .Z(o[23]) );
  AND U1659 ( .A(y[24]), .B(x[32]), .Z(n1507) );
  NAND U1660 ( .A(y[0]), .B(x[24]), .Z(n1506) );
  XNOR U1661 ( .A(n1507), .B(n1506), .Z(n1508) );
  NAND U1662 ( .A(y[48]), .B(x[40]), .Z(n1594) );
  XNOR U1663 ( .A(n1508), .B(n1594), .Z(o[24]) );
  AND U1664 ( .A(y[24]), .B(x[33]), .Z(n1581) );
  AND U1665 ( .A(y[25]), .B(x[32]), .Z(n1518) );
  AND U1666 ( .A(y[48]), .B(x[41]), .Z(n1517) );
  XOR U1667 ( .A(n1518), .B(n1517), .Z(n1519) );
  XNOR U1668 ( .A(n1581), .B(n1519), .Z(n1514) );
  NANDN U1669 ( .A(n1507), .B(n1506), .Z(n1510) );
  NAND U1670 ( .A(n1508), .B(n1594), .Z(n1509) );
  AND U1671 ( .A(n1510), .B(n1509), .Z(n1512) );
  AND U1672 ( .A(y[1]), .B(x[24]), .Z(n1545) );
  AND U1673 ( .A(y[49]), .B(x[40]), .Z(n1553) );
  AND U1674 ( .A(y[0]), .B(x[25]), .Z(n1522) );
  XOR U1675 ( .A(n1553), .B(n1522), .Z(n1523) );
  XNOR U1676 ( .A(n1545), .B(n1523), .Z(n1513) );
  XNOR U1677 ( .A(n1512), .B(n1513), .Z(n1511) );
  XNOR U1678 ( .A(n1514), .B(n1511), .Z(o[25]) );
  AND U1679 ( .A(x[25]), .B(y[1]), .Z(n1516) );
  NAND U1680 ( .A(x[24]), .B(y[2]), .Z(n1515) );
  XNOR U1681 ( .A(n1516), .B(n1515), .Z(n1547) );
  AND U1682 ( .A(y[24]), .B(x[34]), .Z(n1546) );
  XOR U1683 ( .A(n1547), .B(n1546), .Z(n1560) );
  AND U1684 ( .A(y[26]), .B(x[32]), .Z(n1558) );
  NAND U1685 ( .A(y[25]), .B(x[33]), .Z(n1557) );
  XNOR U1686 ( .A(n1558), .B(n1557), .Z(n1559) );
  XNOR U1687 ( .A(n1560), .B(n1559), .Z(n1533) );
  XNOR U1688 ( .A(n1534), .B(n1533), .Z(n1536) );
  NAND U1689 ( .A(n1518), .B(n1517), .Z(n1521) );
  NAND U1690 ( .A(n1581), .B(n1519), .Z(n1520) );
  NAND U1691 ( .A(n1521), .B(n1520), .Z(n1529) );
  NAND U1692 ( .A(n1553), .B(n1522), .Z(n1525) );
  NAND U1693 ( .A(n1545), .B(n1523), .Z(n1524) );
  NAND U1694 ( .A(n1525), .B(n1524), .Z(n1527) );
  AND U1695 ( .A(y[0]), .B(x[26]), .Z(n1573) );
  NAND U1696 ( .A(y[48]), .B(x[42]), .Z(n1539) );
  XNOR U1697 ( .A(n1573), .B(n1539), .Z(n1541) );
  AND U1698 ( .A(x[41]), .B(y[49]), .Z(n1587) );
  NAND U1699 ( .A(x[40]), .B(y[50]), .Z(n1526) );
  XNOR U1700 ( .A(n1587), .B(n1526), .Z(n1540) );
  XOR U1701 ( .A(n1541), .B(n1540), .Z(n1528) );
  XNOR U1702 ( .A(n1527), .B(n1528), .Z(n1530) );
  XOR U1703 ( .A(n1529), .B(n1530), .Z(n1535) );
  XNOR U1704 ( .A(n1536), .B(n1535), .Z(o[26]) );
  NAND U1705 ( .A(n1528), .B(n1527), .Z(n1532) );
  NANDN U1706 ( .A(n1530), .B(n1529), .Z(n1531) );
  AND U1707 ( .A(n1532), .B(n1531), .Z(n1568) );
  NANDN U1708 ( .A(n1534), .B(n1533), .Z(n1538) );
  NAND U1709 ( .A(n1536), .B(n1535), .Z(n1537) );
  AND U1710 ( .A(n1538), .B(n1537), .Z(n1567) );
  XNOR U1711 ( .A(n1568), .B(n1567), .Z(n1570) );
  NANDN U1712 ( .A(n1539), .B(n1573), .Z(n1543) );
  NAND U1713 ( .A(n1541), .B(n1540), .Z(n1542) );
  NAND U1714 ( .A(n1543), .B(n1542), .Z(n1601) );
  AND U1715 ( .A(y[27]), .B(x[32]), .Z(n1588) );
  AND U1716 ( .A(y[2]), .B(x[25]), .Z(n1589) );
  NAND U1717 ( .A(y[3]), .B(x[24]), .Z(n1591) );
  XNOR U1718 ( .A(n1590), .B(n1591), .Z(n1600) );
  AND U1719 ( .A(x[33]), .B(y[26]), .Z(n1611) );
  NAND U1720 ( .A(x[35]), .B(y[24]), .Z(n1544) );
  XNOR U1721 ( .A(n1611), .B(n1544), .Z(n1583) );
  AND U1722 ( .A(y[25]), .B(x[34]), .Z(n1582) );
  XOR U1723 ( .A(n1583), .B(n1582), .Z(n1599) );
  XOR U1724 ( .A(n1600), .B(n1599), .Z(n1602) );
  XOR U1725 ( .A(n1601), .B(n1602), .Z(n1564) );
  NAND U1726 ( .A(n1589), .B(n1545), .Z(n1549) );
  NAND U1727 ( .A(n1547), .B(n1546), .Z(n1548) );
  NAND U1728 ( .A(n1549), .B(n1548), .Z(n1607) );
  AND U1729 ( .A(x[26]), .B(y[1]), .Z(n1551) );
  NAND U1730 ( .A(x[27]), .B(y[0]), .Z(n1550) );
  XNOR U1731 ( .A(n1551), .B(n1550), .Z(n1574) );
  AND U1732 ( .A(y[50]), .B(x[41]), .Z(n1552) );
  NAND U1733 ( .A(n1553), .B(n1552), .Z(n1575) );
  XNOR U1734 ( .A(n1574), .B(n1575), .Z(n1606) );
  AND U1735 ( .A(x[43]), .B(y[48]), .Z(n1555) );
  NAND U1736 ( .A(x[40]), .B(y[51]), .Z(n1554) );
  XNOR U1737 ( .A(n1555), .B(n1554), .Z(n1596) );
  AND U1738 ( .A(x[42]), .B(y[49]), .Z(n1621) );
  NAND U1739 ( .A(x[41]), .B(y[50]), .Z(n1556) );
  XNOR U1740 ( .A(n1621), .B(n1556), .Z(n1595) );
  XOR U1741 ( .A(n1596), .B(n1595), .Z(n1605) );
  XOR U1742 ( .A(n1606), .B(n1605), .Z(n1608) );
  XNOR U1743 ( .A(n1607), .B(n1608), .Z(n1563) );
  XNOR U1744 ( .A(n1564), .B(n1563), .Z(n1565) );
  NANDN U1745 ( .A(n1558), .B(n1557), .Z(n1562) );
  NANDN U1746 ( .A(n1560), .B(n1559), .Z(n1561) );
  NAND U1747 ( .A(n1562), .B(n1561), .Z(n1566) );
  XNOR U1748 ( .A(n1565), .B(n1566), .Z(n1569) );
  XOR U1749 ( .A(n1570), .B(n1569), .Z(o[27]) );
  NANDN U1750 ( .A(n1568), .B(n1567), .Z(n1572) );
  NAND U1751 ( .A(n1570), .B(n1569), .Z(n1571) );
  NAND U1752 ( .A(n1572), .B(n1571), .Z(n1670) );
  XNOR U1753 ( .A(n1671), .B(n1670), .Z(n1673) );
  AND U1754 ( .A(y[1]), .B(x[27]), .Z(n1638) );
  NAND U1755 ( .A(n1638), .B(n1573), .Z(n1577) );
  NANDN U1756 ( .A(n1575), .B(n1574), .Z(n1576) );
  NAND U1757 ( .A(n1577), .B(n1576), .Z(n1651) );
  AND U1758 ( .A(x[43]), .B(y[49]), .Z(n1748) );
  NAND U1759 ( .A(x[42]), .B(y[50]), .Z(n1578) );
  XNOR U1760 ( .A(n1748), .B(n1578), .Z(n1624) );
  NAND U1761 ( .A(y[51]), .B(x[41]), .Z(n1625) );
  XNOR U1762 ( .A(n1624), .B(n1625), .Z(n1626) );
  NAND U1763 ( .A(y[48]), .B(x[44]), .Z(n1627) );
  XNOR U1764 ( .A(n1626), .B(n1627), .Z(n1648) );
  AND U1765 ( .A(x[33]), .B(y[27]), .Z(n1580) );
  NAND U1766 ( .A(x[34]), .B(y[26]), .Z(n1579) );
  XNOR U1767 ( .A(n1580), .B(n1579), .Z(n1612) );
  NAND U1768 ( .A(y[25]), .B(x[35]), .Z(n1613) );
  XNOR U1769 ( .A(n1612), .B(n1613), .Z(n1649) );
  AND U1770 ( .A(y[26]), .B(x[35]), .Z(n1727) );
  NAND U1771 ( .A(n1727), .B(n1581), .Z(n1585) );
  NAND U1772 ( .A(n1583), .B(n1582), .Z(n1584) );
  NAND U1773 ( .A(n1585), .B(n1584), .Z(n1645) );
  AND U1774 ( .A(y[52]), .B(x[40]), .Z(n1711) );
  AND U1775 ( .A(y[0]), .B(x[28]), .Z(n1630) );
  AND U1776 ( .A(y[50]), .B(x[42]), .Z(n1586) );
  NAND U1777 ( .A(n1587), .B(n1586), .Z(n1631) );
  XOR U1778 ( .A(n1630), .B(n1631), .Z(n1632) );
  XNOR U1779 ( .A(n1711), .B(n1632), .Z(n1642) );
  AND U1780 ( .A(y[24]), .B(x[36]), .Z(n1742) );
  AND U1781 ( .A(y[28]), .B(x[32]), .Z(n1616) );
  XOR U1782 ( .A(n1742), .B(n1616), .Z(n1618) );
  NAND U1783 ( .A(y[3]), .B(x[25]), .Z(n1617) );
  XNOR U1784 ( .A(n1618), .B(n1617), .Z(n1643) );
  XNOR U1785 ( .A(n1655), .B(n1654), .Z(n1657) );
  NAND U1786 ( .A(n1589), .B(n1588), .Z(n1593) );
  NANDN U1787 ( .A(n1591), .B(n1590), .Z(n1592) );
  NAND U1788 ( .A(n1593), .B(n1592), .Z(n1660) );
  AND U1789 ( .A(y[2]), .B(x[26]), .Z(n1641) );
  NAND U1790 ( .A(y[4]), .B(x[24]), .Z(n1639) );
  XNOR U1791 ( .A(n1638), .B(n1639), .Z(n1640) );
  XOR U1792 ( .A(n1641), .B(n1640), .Z(n1659) );
  AND U1793 ( .A(y[51]), .B(x[43]), .Z(n1866) );
  NANDN U1794 ( .A(n1594), .B(n1866), .Z(n1598) );
  NAND U1795 ( .A(n1596), .B(n1595), .Z(n1597) );
  NAND U1796 ( .A(n1598), .B(n1597), .Z(n1658) );
  XOR U1797 ( .A(n1659), .B(n1658), .Z(n1661) );
  XNOR U1798 ( .A(n1660), .B(n1661), .Z(n1656) );
  XNOR U1799 ( .A(n1657), .B(n1656), .Z(n1667) );
  NAND U1800 ( .A(n1600), .B(n1599), .Z(n1604) );
  NAND U1801 ( .A(n1602), .B(n1601), .Z(n1603) );
  AND U1802 ( .A(n1604), .B(n1603), .Z(n1665) );
  NAND U1803 ( .A(n1606), .B(n1605), .Z(n1610) );
  NAND U1804 ( .A(n1608), .B(n1607), .Z(n1609) );
  AND U1805 ( .A(n1610), .B(n1609), .Z(n1664) );
  XOR U1806 ( .A(n1665), .B(n1664), .Z(n1666) );
  XOR U1807 ( .A(n1667), .B(n1666), .Z(n1672) );
  XOR U1808 ( .A(n1673), .B(n1672), .Z(o[28]) );
  AND U1809 ( .A(y[27]), .B(x[34]), .Z(n1716) );
  NAND U1810 ( .A(n1716), .B(n1611), .Z(n1615) );
  NANDN U1811 ( .A(n1613), .B(n1612), .Z(n1614) );
  AND U1812 ( .A(n1615), .B(n1614), .Z(n1697) );
  AND U1813 ( .A(y[0]), .B(x[29]), .Z(n1820) );
  XOR U1814 ( .A(n1820), .B(n1716), .Z(n1718) );
  AND U1815 ( .A(y[1]), .B(x[28]), .Z(n1717) );
  XOR U1816 ( .A(n1718), .B(n1717), .Z(n1695) );
  AND U1817 ( .A(y[28]), .B(x[33]), .Z(n1878) );
  AND U1818 ( .A(y[5]), .B(x[24]), .Z(n1705) );
  AND U1819 ( .A(y[29]), .B(x[32]), .Z(n1704) );
  XOR U1820 ( .A(n1705), .B(n1704), .Z(n1706) );
  XNOR U1821 ( .A(n1878), .B(n1706), .Z(n1694) );
  XNOR U1822 ( .A(n1695), .B(n1694), .Z(n1696) );
  XOR U1823 ( .A(n1697), .B(n1696), .Z(n1689) );
  NAND U1824 ( .A(n1742), .B(n1616), .Z(n1620) );
  ANDN U1825 ( .B(n1618), .A(n1617), .Z(n1619) );
  ANDN U1826 ( .B(n1620), .A(n1619), .Z(n1700) );
  AND U1827 ( .A(x[43]), .B(y[50]), .Z(n1637) );
  AND U1828 ( .A(n1637), .B(n1621), .Z(n1713) );
  AND U1829 ( .A(x[40]), .B(y[53]), .Z(n1623) );
  AND U1830 ( .A(x[41]), .B(y[52]), .Z(n1622) );
  XOR U1831 ( .A(n1623), .B(n1622), .Z(n1712) );
  XOR U1832 ( .A(n1713), .B(n1712), .Z(n1698) );
  AND U1833 ( .A(y[2]), .B(x[27]), .Z(n1807) );
  NAND U1834 ( .A(y[3]), .B(x[26]), .Z(n1729) );
  XOR U1835 ( .A(n1728), .B(n1729), .Z(n1699) );
  XOR U1836 ( .A(n1698), .B(n1699), .Z(n1701) );
  XNOR U1837 ( .A(n1700), .B(n1701), .Z(n1688) );
  XOR U1838 ( .A(n1689), .B(n1688), .Z(n1691) );
  NANDN U1839 ( .A(n1625), .B(n1624), .Z(n1629) );
  NANDN U1840 ( .A(n1627), .B(n1626), .Z(n1628) );
  AND U1841 ( .A(n1629), .B(n1628), .Z(n1751) );
  NANDN U1842 ( .A(n1631), .B(n1630), .Z(n1634) );
  NANDN U1843 ( .A(n1632), .B(n1711), .Z(n1633) );
  AND U1844 ( .A(n1634), .B(n1633), .Z(n1726) );
  AND U1845 ( .A(x[37]), .B(y[24]), .Z(n1636) );
  NAND U1846 ( .A(x[36]), .B(y[25]), .Z(n1635) );
  XNOR U1847 ( .A(n1636), .B(n1635), .Z(n1744) );
  AND U1848 ( .A(y[4]), .B(x[25]), .Z(n1743) );
  XOR U1849 ( .A(n1744), .B(n1743), .Z(n1724) );
  AND U1850 ( .A(y[51]), .B(x[42]), .Z(n1735) );
  AND U1851 ( .A(y[48]), .B(x[45]), .Z(n1734) );
  XOR U1852 ( .A(n1735), .B(n1734), .Z(n1737) );
  AND U1853 ( .A(y[49]), .B(x[44]), .Z(n1875) );
  XOR U1854 ( .A(n1875), .B(n1637), .Z(n1736) );
  XNOR U1855 ( .A(n1737), .B(n1736), .Z(n1723) );
  XNOR U1856 ( .A(n1724), .B(n1723), .Z(n1725) );
  XNOR U1857 ( .A(n1726), .B(n1725), .Z(n1749) );
  XOR U1858 ( .A(n1749), .B(n1750), .Z(n1752) );
  XNOR U1859 ( .A(n1751), .B(n1752), .Z(n1690) );
  XNOR U1860 ( .A(n1691), .B(n1690), .Z(n1685) );
  NAND U1861 ( .A(n1643), .B(n1642), .Z(n1647) );
  NAND U1862 ( .A(n1645), .B(n1644), .Z(n1646) );
  NAND U1863 ( .A(n1647), .B(n1646), .Z(n1683) );
  NAND U1864 ( .A(n1649), .B(n1648), .Z(n1653) );
  NAND U1865 ( .A(n1651), .B(n1650), .Z(n1652) );
  NAND U1866 ( .A(n1653), .B(n1652), .Z(n1682) );
  NAND U1867 ( .A(n1659), .B(n1658), .Z(n1663) );
  NAND U1868 ( .A(n1661), .B(n1660), .Z(n1662) );
  NAND U1869 ( .A(n1663), .B(n1662), .Z(n1677) );
  XNOR U1870 ( .A(n1676), .B(n1677), .Z(n1678) );
  XOR U1871 ( .A(n1679), .B(n1678), .Z(n1758) );
  NAND U1872 ( .A(n1665), .B(n1664), .Z(n1669) );
  NANDN U1873 ( .A(n1667), .B(n1666), .Z(n1668) );
  AND U1874 ( .A(n1669), .B(n1668), .Z(n1756) );
  NANDN U1875 ( .A(n1671), .B(n1670), .Z(n1675) );
  NAND U1876 ( .A(n1673), .B(n1672), .Z(n1674) );
  AND U1877 ( .A(n1675), .B(n1674), .Z(n1755) );
  XNOR U1878 ( .A(n1756), .B(n1755), .Z(n1757) );
  XNOR U1879 ( .A(n1758), .B(n1757), .Z(o[29]) );
  NANDN U1880 ( .A(n1677), .B(n1676), .Z(n1681) );
  NAND U1881 ( .A(n1679), .B(n1678), .Z(n1680) );
  AND U1882 ( .A(n1681), .B(n1680), .Z(n1928) );
  NAND U1883 ( .A(n1683), .B(n1682), .Z(n1687) );
  NAND U1884 ( .A(n1685), .B(n1684), .Z(n1686) );
  NAND U1885 ( .A(n1687), .B(n1686), .Z(n1934) );
  NAND U1886 ( .A(n1689), .B(n1688), .Z(n1693) );
  NAND U1887 ( .A(n1691), .B(n1690), .Z(n1692) );
  AND U1888 ( .A(n1693), .B(n1692), .Z(n1933) );
  NANDN U1889 ( .A(n1699), .B(n1698), .Z(n1703) );
  OR U1890 ( .A(n1701), .B(n1700), .Z(n1702) );
  AND U1891 ( .A(n1703), .B(n1702), .Z(n1915) );
  XOR U1892 ( .A(n1916), .B(n1915), .Z(n1914) );
  NAND U1893 ( .A(n1705), .B(n1704), .Z(n1708) );
  NAND U1894 ( .A(n1878), .B(n1706), .Z(n1707) );
  AND U1895 ( .A(n1708), .B(n1707), .Z(n1779) );
  AND U1896 ( .A(x[29]), .B(y[1]), .Z(n1710) );
  NAND U1897 ( .A(x[30]), .B(y[0]), .Z(n1709) );
  XNOR U1898 ( .A(n1710), .B(n1709), .Z(n1819) );
  AND U1899 ( .A(y[27]), .B(x[35]), .Z(n1818) );
  XNOR U1900 ( .A(n1819), .B(n1818), .Z(n1782) );
  AND U1901 ( .A(y[5]), .B(x[25]), .Z(n1800) );
  AND U1902 ( .A(y[54]), .B(x[40]), .Z(n1802) );
  AND U1903 ( .A(y[30]), .B(x[32]), .Z(n1801) );
  XOR U1904 ( .A(n1802), .B(n1801), .Z(n1799) );
  XNOR U1905 ( .A(n1800), .B(n1799), .Z(n1781) );
  XNOR U1906 ( .A(n1779), .B(n1780), .Z(n1908) );
  AND U1907 ( .A(y[53]), .B(x[41]), .Z(n1849) );
  NAND U1908 ( .A(n1711), .B(n1849), .Z(n1715) );
  NAND U1909 ( .A(n1713), .B(n1712), .Z(n1714) );
  AND U1910 ( .A(n1715), .B(n1714), .Z(n1910) );
  NAND U1911 ( .A(n1820), .B(n1716), .Z(n1720) );
  NAND U1912 ( .A(n1718), .B(n1717), .Z(n1719) );
  AND U1913 ( .A(n1720), .B(n1719), .Z(n1773) );
  AND U1914 ( .A(y[25]), .B(x[37]), .Z(n1813) );
  AND U1915 ( .A(y[24]), .B(x[38]), .Z(n1815) );
  AND U1916 ( .A(y[6]), .B(x[24]), .Z(n1814) );
  XOR U1917 ( .A(n1815), .B(n1814), .Z(n1812) );
  XNOR U1918 ( .A(n1813), .B(n1812), .Z(n1776) );
  AND U1919 ( .A(x[45]), .B(y[49]), .Z(n1722) );
  NAND U1920 ( .A(x[44]), .B(y[50]), .Z(n1721) );
  XNOR U1921 ( .A(n1722), .B(n1721), .Z(n1869) );
  AND U1922 ( .A(y[48]), .B(x[46]), .Z(n1868) );
  XOR U1923 ( .A(n1869), .B(n1868), .Z(n1867) );
  XNOR U1924 ( .A(n1867), .B(n1866), .Z(n1775) );
  XNOR U1925 ( .A(n1773), .B(n1774), .Z(n1909) );
  XOR U1926 ( .A(n1910), .B(n1909), .Z(n1907) );
  XOR U1927 ( .A(n1908), .B(n1907), .Z(n1913) );
  XOR U1928 ( .A(n1914), .B(n1913), .Z(n1762) );
  NAND U1929 ( .A(n1807), .B(n1727), .Z(n1731) );
  NANDN U1930 ( .A(n1729), .B(n1728), .Z(n1730) );
  AND U1931 ( .A(n1731), .B(n1730), .Z(n1786) );
  AND U1932 ( .A(x[33]), .B(y[29]), .Z(n1733) );
  NAND U1933 ( .A(x[34]), .B(y[28]), .Z(n1732) );
  XNOR U1934 ( .A(n1733), .B(n1732), .Z(n1877) );
  AND U1935 ( .A(y[4]), .B(x[26]), .Z(n1876) );
  XNOR U1936 ( .A(n1877), .B(n1876), .Z(n1788) );
  NAND U1937 ( .A(n1735), .B(n1734), .Z(n1739) );
  NAND U1938 ( .A(n1737), .B(n1736), .Z(n1738) );
  AND U1939 ( .A(n1739), .B(n1738), .Z(n1787) );
  XOR U1940 ( .A(n1786), .B(n1785), .Z(n1769) );
  XOR U1941 ( .A(n1770), .B(n1769), .Z(n1768) );
  AND U1942 ( .A(x[27]), .B(y[3]), .Z(n1741) );
  NAND U1943 ( .A(x[28]), .B(y[2]), .Z(n1740) );
  XNOR U1944 ( .A(n1741), .B(n1740), .Z(n1806) );
  AND U1945 ( .A(y[26]), .B(x[36]), .Z(n1805) );
  XNOR U1946 ( .A(n1806), .B(n1805), .Z(n1796) );
  NAND U1947 ( .A(n1813), .B(n1742), .Z(n1746) );
  NAND U1948 ( .A(n1744), .B(n1743), .Z(n1745) );
  AND U1949 ( .A(n1746), .B(n1745), .Z(n1795) );
  AND U1950 ( .A(y[50]), .B(x[44]), .Z(n1747) );
  AND U1951 ( .A(n1748), .B(n1747), .Z(n1851) );
  AND U1952 ( .A(y[52]), .B(x[42]), .Z(n1850) );
  XOR U1953 ( .A(n1851), .B(n1850), .Z(n1848) );
  XNOR U1954 ( .A(n1849), .B(n1848), .Z(n1794) );
  XNOR U1955 ( .A(n1768), .B(n1767), .Z(n1764) );
  NANDN U1956 ( .A(n1750), .B(n1749), .Z(n1754) );
  OR U1957 ( .A(n1752), .B(n1751), .Z(n1753) );
  NAND U1958 ( .A(n1754), .B(n1753), .Z(n1763) );
  XNOR U1959 ( .A(n1762), .B(n1761), .Z(n1932) );
  XOR U1960 ( .A(n1928), .B(n1927), .Z(n1926) );
  NANDN U1961 ( .A(n1756), .B(n1755), .Z(n1760) );
  NAND U1962 ( .A(n1758), .B(n1757), .Z(n1759) );
  AND U1963 ( .A(n1760), .B(n1759), .Z(n1925) );
  XOR U1964 ( .A(n1926), .B(n1925), .Z(o[30]) );
  NANDN U1965 ( .A(n1762), .B(n1761), .Z(n1766) );
  NAND U1966 ( .A(n1764), .B(n1763), .Z(n1765) );
  AND U1967 ( .A(n1766), .B(n1765), .Z(n1942) );
  NAND U1968 ( .A(n1768), .B(n1767), .Z(n1772) );
  NAND U1969 ( .A(n1770), .B(n1769), .Z(n1771) );
  AND U1970 ( .A(n1772), .B(n1771), .Z(n1924) );
  NANDN U1971 ( .A(n1774), .B(n1773), .Z(n1778) );
  NAND U1972 ( .A(n1776), .B(n1775), .Z(n1777) );
  AND U1973 ( .A(n1778), .B(n1777), .Z(n1906) );
  NANDN U1974 ( .A(n1780), .B(n1779), .Z(n1784) );
  NAND U1975 ( .A(n1782), .B(n1781), .Z(n1783) );
  AND U1976 ( .A(n1784), .B(n1783), .Z(n1792) );
  NAND U1977 ( .A(n1786), .B(n1785), .Z(n1790) );
  NAND U1978 ( .A(n1788), .B(n1787), .Z(n1789) );
  NAND U1979 ( .A(n1790), .B(n1789), .Z(n1791) );
  XNOR U1980 ( .A(n1792), .B(n1791), .Z(n1904) );
  NAND U1981 ( .A(n1794), .B(n1793), .Z(n1798) );
  NAND U1982 ( .A(n1796), .B(n1795), .Z(n1797) );
  AND U1983 ( .A(n1798), .B(n1797), .Z(n1902) );
  NAND U1984 ( .A(n1800), .B(n1799), .Z(n1804) );
  NAND U1985 ( .A(n1802), .B(n1801), .Z(n1803) );
  AND U1986 ( .A(n1804), .B(n1803), .Z(n1811) );
  NAND U1987 ( .A(n1806), .B(n1805), .Z(n1809) );
  AND U1988 ( .A(y[3]), .B(x[28]), .Z(n1891) );
  NAND U1989 ( .A(n1807), .B(n1891), .Z(n1808) );
  NAND U1990 ( .A(n1809), .B(n1808), .Z(n1810) );
  XNOR U1991 ( .A(n1811), .B(n1810), .Z(n1826) );
  NAND U1992 ( .A(n1813), .B(n1812), .Z(n1817) );
  NAND U1993 ( .A(n1815), .B(n1814), .Z(n1816) );
  AND U1994 ( .A(n1817), .B(n1816), .Z(n1824) );
  NAND U1995 ( .A(n1819), .B(n1818), .Z(n1822) );
  AND U1996 ( .A(y[1]), .B(x[30]), .Z(n1835) );
  NAND U1997 ( .A(n1820), .B(n1835), .Z(n1821) );
  NAND U1998 ( .A(n1822), .B(n1821), .Z(n1823) );
  XNOR U1999 ( .A(n1824), .B(n1823), .Z(n1825) );
  XOR U2000 ( .A(n1826), .B(n1825), .Z(n1865) );
  AND U2001 ( .A(x[26]), .B(y[5]), .Z(n1828) );
  NAND U2002 ( .A(x[37]), .B(y[26]), .Z(n1827) );
  XNOR U2003 ( .A(n1828), .B(n1827), .Z(n1839) );
  AND U2004 ( .A(x[41]), .B(y[54]), .Z(n1830) );
  NAND U2005 ( .A(x[38]), .B(y[25]), .Z(n1829) );
  XNOR U2006 ( .A(n1830), .B(n1829), .Z(n1834) );
  AND U2007 ( .A(x[24]), .B(y[7]), .Z(n1832) );
  NAND U2008 ( .A(x[31]), .B(y[0]), .Z(n1831) );
  XNOR U2009 ( .A(n1832), .B(n1831), .Z(n1833) );
  XOR U2010 ( .A(n1834), .B(n1833), .Z(n1837) );
  AND U2011 ( .A(y[50]), .B(x[45]), .Z(n1874) );
  XNOR U2012 ( .A(n1835), .B(n1874), .Z(n1836) );
  XNOR U2013 ( .A(n1837), .B(n1836), .Z(n1838) );
  XOR U2014 ( .A(n1839), .B(n1838), .Z(n1847) );
  AND U2015 ( .A(x[33]), .B(y[30]), .Z(n1841) );
  NAND U2016 ( .A(x[47]), .B(y[48]), .Z(n1840) );
  XNOR U2017 ( .A(n1841), .B(n1840), .Z(n1845) );
  AND U2018 ( .A(x[46]), .B(y[49]), .Z(n1843) );
  NAND U2019 ( .A(x[44]), .B(y[51]), .Z(n1842) );
  XNOR U2020 ( .A(n1843), .B(n1842), .Z(n1844) );
  XNOR U2021 ( .A(n1845), .B(n1844), .Z(n1846) );
  XNOR U2022 ( .A(n1847), .B(n1846), .Z(n1863) );
  NAND U2023 ( .A(n1849), .B(n1848), .Z(n1853) );
  NAND U2024 ( .A(n1851), .B(n1850), .Z(n1852) );
  AND U2025 ( .A(n1853), .B(n1852), .Z(n1861) );
  AND U2026 ( .A(x[32]), .B(y[31]), .Z(n1855) );
  NAND U2027 ( .A(x[25]), .B(y[6]), .Z(n1854) );
  XNOR U2028 ( .A(n1855), .B(n1854), .Z(n1859) );
  AND U2029 ( .A(x[40]), .B(y[55]), .Z(n1857) );
  NAND U2030 ( .A(x[27]), .B(y[4]), .Z(n1856) );
  XNOR U2031 ( .A(n1857), .B(n1856), .Z(n1858) );
  XNOR U2032 ( .A(n1859), .B(n1858), .Z(n1860) );
  XNOR U2033 ( .A(n1861), .B(n1860), .Z(n1862) );
  XNOR U2034 ( .A(n1863), .B(n1862), .Z(n1864) );
  XNOR U2035 ( .A(n1865), .B(n1864), .Z(n1900) );
  NAND U2036 ( .A(n1867), .B(n1866), .Z(n1871) );
  NAND U2037 ( .A(n1869), .B(n1868), .Z(n1870) );
  AND U2038 ( .A(n1871), .B(n1870), .Z(n1898) );
  AND U2039 ( .A(x[42]), .B(y[53]), .Z(n1873) );
  NAND U2040 ( .A(x[43]), .B(y[52]), .Z(n1872) );
  XNOR U2041 ( .A(n1873), .B(n1872), .Z(n1896) );
  AND U2042 ( .A(n1875), .B(n1874), .Z(n1890) );
  NAND U2043 ( .A(n1877), .B(n1876), .Z(n1880) );
  AND U2044 ( .A(y[29]), .B(x[34]), .Z(n1892) );
  NAND U2045 ( .A(n1892), .B(n1878), .Z(n1879) );
  AND U2046 ( .A(n1880), .B(n1879), .Z(n1888) );
  AND U2047 ( .A(x[36]), .B(y[27]), .Z(n1882) );
  NAND U2048 ( .A(x[29]), .B(y[2]), .Z(n1881) );
  XNOR U2049 ( .A(n1882), .B(n1881), .Z(n1886) );
  AND U2050 ( .A(x[35]), .B(y[28]), .Z(n1884) );
  NAND U2051 ( .A(x[39]), .B(y[24]), .Z(n1883) );
  XNOR U2052 ( .A(n1884), .B(n1883), .Z(n1885) );
  XNOR U2053 ( .A(n1886), .B(n1885), .Z(n1887) );
  XNOR U2054 ( .A(n1888), .B(n1887), .Z(n1889) );
  XOR U2055 ( .A(n1890), .B(n1889), .Z(n1894) );
  XNOR U2056 ( .A(n1892), .B(n1891), .Z(n1893) );
  XNOR U2057 ( .A(n1894), .B(n1893), .Z(n1895) );
  XNOR U2058 ( .A(n1896), .B(n1895), .Z(n1897) );
  XNOR U2059 ( .A(n1898), .B(n1897), .Z(n1899) );
  XNOR U2060 ( .A(n1900), .B(n1899), .Z(n1901) );
  XNOR U2061 ( .A(n1902), .B(n1901), .Z(n1903) );
  XNOR U2062 ( .A(n1904), .B(n1903), .Z(n1905) );
  XNOR U2063 ( .A(n1906), .B(n1905), .Z(n1922) );
  NAND U2064 ( .A(n1908), .B(n1907), .Z(n1912) );
  NAND U2065 ( .A(n1910), .B(n1909), .Z(n1911) );
  AND U2066 ( .A(n1912), .B(n1911), .Z(n1920) );
  NAND U2067 ( .A(n1914), .B(n1913), .Z(n1918) );
  NAND U2068 ( .A(n1916), .B(n1915), .Z(n1917) );
  NAND U2069 ( .A(n1918), .B(n1917), .Z(n1919) );
  XNOR U2070 ( .A(n1920), .B(n1919), .Z(n1921) );
  XNOR U2071 ( .A(n1922), .B(n1921), .Z(n1923) );
  XNOR U2072 ( .A(n1924), .B(n1923), .Z(n1940) );
  NAND U2073 ( .A(n1926), .B(n1925), .Z(n1930) );
  NAND U2074 ( .A(n1928), .B(n1927), .Z(n1929) );
  AND U2075 ( .A(n1930), .B(n1929), .Z(n1938) );
  NAND U2076 ( .A(n1932), .B(n1931), .Z(n1936) );
  NAND U2077 ( .A(n1934), .B(n1933), .Z(n1935) );
  NAND U2078 ( .A(n1936), .B(n1935), .Z(n1937) );
  XNOR U2079 ( .A(n1938), .B(n1937), .Z(n1939) );
  XNOR U2080 ( .A(n1940), .B(n1939), .Z(n1941) );
  XNOR U2081 ( .A(n1942), .B(n1941), .Z(o[31]) );
  AND U2082 ( .A(y[32]), .B(x[32]), .Z(n1944) );
  NAND U2083 ( .A(y[8]), .B(x[24]), .Z(n1943) );
  XNOR U2084 ( .A(n1944), .B(n1943), .Z(n1945) );
  NAND U2085 ( .A(y[56]), .B(x[40]), .Z(n2033) );
  XNOR U2086 ( .A(n1945), .B(n2033), .Z(o[32]) );
  AND U2087 ( .A(y[32]), .B(x[33]), .Z(n2020) );
  AND U2088 ( .A(y[33]), .B(x[32]), .Z(n1955) );
  AND U2089 ( .A(y[56]), .B(x[41]), .Z(n1954) );
  XOR U2090 ( .A(n1955), .B(n1954), .Z(n1956) );
  XNOR U2091 ( .A(n2020), .B(n1956), .Z(n1951) );
  NANDN U2092 ( .A(n1944), .B(n1943), .Z(n1947) );
  NAND U2093 ( .A(n1945), .B(n2033), .Z(n1946) );
  AND U2094 ( .A(n1947), .B(n1946), .Z(n1949) );
  AND U2095 ( .A(y[9]), .B(x[24]), .Z(n1984) );
  AND U2096 ( .A(y[57]), .B(x[40]), .Z(n1991) );
  AND U2097 ( .A(y[8]), .B(x[25]), .Z(n1959) );
  XOR U2098 ( .A(n1991), .B(n1959), .Z(n1960) );
  XNOR U2099 ( .A(n1984), .B(n1960), .Z(n1950) );
  XNOR U2100 ( .A(n1949), .B(n1950), .Z(n1948) );
  XNOR U2101 ( .A(n1951), .B(n1948), .Z(o[33]) );
  AND U2102 ( .A(x[24]), .B(y[10]), .Z(n1953) );
  NAND U2103 ( .A(x[25]), .B(y[9]), .Z(n1952) );
  XNOR U2104 ( .A(n1953), .B(n1952), .Z(n1986) );
  AND U2105 ( .A(y[32]), .B(x[34]), .Z(n1985) );
  XOR U2106 ( .A(n1986), .B(n1985), .Z(n1999) );
  AND U2107 ( .A(y[34]), .B(x[32]), .Z(n1997) );
  NAND U2108 ( .A(y[33]), .B(x[33]), .Z(n1996) );
  XNOR U2109 ( .A(n1997), .B(n1996), .Z(n1998) );
  XNOR U2110 ( .A(n1999), .B(n1998), .Z(n1971) );
  XNOR U2111 ( .A(n1972), .B(n1971), .Z(n1974) );
  NAND U2112 ( .A(n1955), .B(n1954), .Z(n1958) );
  NAND U2113 ( .A(n2020), .B(n1956), .Z(n1957) );
  NAND U2114 ( .A(n1958), .B(n1957), .Z(n1967) );
  NAND U2115 ( .A(n1991), .B(n1959), .Z(n1962) );
  NAND U2116 ( .A(n1984), .B(n1960), .Z(n1961) );
  NAND U2117 ( .A(n1962), .B(n1961), .Z(n1965) );
  AND U2118 ( .A(y[8]), .B(x[26]), .Z(n2012) );
  NAND U2119 ( .A(y[56]), .B(x[42]), .Z(n1977) );
  XNOR U2120 ( .A(n2012), .B(n1977), .Z(n1979) );
  AND U2121 ( .A(x[40]), .B(y[58]), .Z(n1964) );
  NAND U2122 ( .A(x[41]), .B(y[57]), .Z(n1963) );
  XNOR U2123 ( .A(n1964), .B(n1963), .Z(n1978) );
  XOR U2124 ( .A(n1979), .B(n1978), .Z(n1966) );
  XNOR U2125 ( .A(n1965), .B(n1966), .Z(n1968) );
  XOR U2126 ( .A(n1967), .B(n1968), .Z(n1973) );
  XNOR U2127 ( .A(n1974), .B(n1973), .Z(o[34]) );
  NAND U2128 ( .A(n1966), .B(n1965), .Z(n1970) );
  NANDN U2129 ( .A(n1968), .B(n1967), .Z(n1969) );
  AND U2130 ( .A(n1970), .B(n1969), .Z(n2007) );
  NANDN U2131 ( .A(n1972), .B(n1971), .Z(n1976) );
  NAND U2132 ( .A(n1974), .B(n1973), .Z(n1975) );
  AND U2133 ( .A(n1976), .B(n1975), .Z(n2006) );
  XNOR U2134 ( .A(n2007), .B(n2006), .Z(n2009) );
  NANDN U2135 ( .A(n1977), .B(n2012), .Z(n1981) );
  NAND U2136 ( .A(n1979), .B(n1978), .Z(n1980) );
  NAND U2137 ( .A(n1981), .B(n1980), .Z(n2040) );
  AND U2138 ( .A(y[35]), .B(x[32]), .Z(n2027) );
  AND U2139 ( .A(y[10]), .B(x[25]), .Z(n2028) );
  NAND U2140 ( .A(y[11]), .B(x[24]), .Z(n2030) );
  XNOR U2141 ( .A(n2029), .B(n2030), .Z(n2039) );
  AND U2142 ( .A(x[35]), .B(y[32]), .Z(n1983) );
  NAND U2143 ( .A(x[33]), .B(y[34]), .Z(n1982) );
  XNOR U2144 ( .A(n1983), .B(n1982), .Z(n2022) );
  AND U2145 ( .A(y[33]), .B(x[34]), .Z(n2021) );
  XOR U2146 ( .A(n2022), .B(n2021), .Z(n2038) );
  XOR U2147 ( .A(n2039), .B(n2038), .Z(n2041) );
  XOR U2148 ( .A(n2040), .B(n2041), .Z(n2003) );
  NAND U2149 ( .A(n2028), .B(n1984), .Z(n1988) );
  NAND U2150 ( .A(n1986), .B(n1985), .Z(n1987) );
  NAND U2151 ( .A(n1988), .B(n1987), .Z(n2046) );
  AND U2152 ( .A(x[26]), .B(y[9]), .Z(n1990) );
  NAND U2153 ( .A(x[27]), .B(y[8]), .Z(n1989) );
  XNOR U2154 ( .A(n1990), .B(n1989), .Z(n2013) );
  AND U2155 ( .A(y[58]), .B(x[41]), .Z(n1995) );
  NAND U2156 ( .A(n1991), .B(n1995), .Z(n2014) );
  XNOR U2157 ( .A(n2013), .B(n2014), .Z(n2045) );
  AND U2158 ( .A(x[43]), .B(y[56]), .Z(n1993) );
  NAND U2159 ( .A(x[40]), .B(y[59]), .Z(n1992) );
  XNOR U2160 ( .A(n1993), .B(n1992), .Z(n2035) );
  NAND U2161 ( .A(x[42]), .B(y[57]), .Z(n1994) );
  XNOR U2162 ( .A(n1995), .B(n1994), .Z(n2034) );
  XOR U2163 ( .A(n2035), .B(n2034), .Z(n2044) );
  XOR U2164 ( .A(n2045), .B(n2044), .Z(n2047) );
  XNOR U2165 ( .A(n2046), .B(n2047), .Z(n2002) );
  XNOR U2166 ( .A(n2003), .B(n2002), .Z(n2004) );
  NANDN U2167 ( .A(n1997), .B(n1996), .Z(n2001) );
  NANDN U2168 ( .A(n1999), .B(n1998), .Z(n2000) );
  NAND U2169 ( .A(n2001), .B(n2000), .Z(n2005) );
  XNOR U2170 ( .A(n2004), .B(n2005), .Z(n2008) );
  XOR U2171 ( .A(n2009), .B(n2008), .Z(o[35]) );
  NANDN U2172 ( .A(n2007), .B(n2006), .Z(n2011) );
  NAND U2173 ( .A(n2009), .B(n2008), .Z(n2010) );
  NAND U2174 ( .A(n2011), .B(n2010), .Z(n2056) );
  XNOR U2175 ( .A(n2057), .B(n2056), .Z(n2059) );
  NAND U2176 ( .A(y[9]), .B(x[27]), .Z(n2088) );
  NANDN U2177 ( .A(n2088), .B(n2012), .Z(n2016) );
  NANDN U2178 ( .A(n2014), .B(n2013), .Z(n2015) );
  NAND U2179 ( .A(n2016), .B(n2015), .Z(n2116) );
  AND U2180 ( .A(x[34]), .B(y[34]), .Z(n2018) );
  NAND U2181 ( .A(x[33]), .B(y[35]), .Z(n2017) );
  XNOR U2182 ( .A(n2018), .B(n2017), .Z(n2092) );
  AND U2183 ( .A(y[33]), .B(x[35]), .Z(n2093) );
  AND U2184 ( .A(x[42]), .B(y[58]), .Z(n2025) );
  NAND U2185 ( .A(x[43]), .B(y[57]), .Z(n2019) );
  XNOR U2186 ( .A(n2025), .B(n2019), .Z(n2079) );
  AND U2187 ( .A(y[56]), .B(x[44]), .Z(n2080) );
  AND U2188 ( .A(y[59]), .B(x[41]), .Z(n2082) );
  XOR U2189 ( .A(n2114), .B(n2113), .Z(n2115) );
  NAND U2190 ( .A(y[34]), .B(x[35]), .Z(n2106) );
  IV U2191 ( .A(n2106), .Z(n2161) );
  NAND U2192 ( .A(n2161), .B(n2020), .Z(n2024) );
  NAND U2193 ( .A(n2022), .B(n2021), .Z(n2023) );
  NAND U2194 ( .A(n2024), .B(n2023), .Z(n2110) );
  AND U2195 ( .A(y[60]), .B(x[40]), .Z(n2137) );
  AND U2196 ( .A(y[57]), .B(x[41]), .Z(n2026) );
  AND U2197 ( .A(n2026), .B(n2025), .Z(n2072) );
  AND U2198 ( .A(y[8]), .B(x[28]), .Z(n2073) );
  XOR U2199 ( .A(n2137), .B(n2074), .Z(n2108) );
  AND U2200 ( .A(y[32]), .B(x[36]), .Z(n2178) );
  AND U2201 ( .A(y[36]), .B(x[32]), .Z(n2099) );
  XOR U2202 ( .A(n2178), .B(n2099), .Z(n2098) );
  AND U2203 ( .A(y[11]), .B(x[25]), .Z(n2097) );
  XOR U2204 ( .A(n2108), .B(n2107), .Z(n2109) );
  XNOR U2205 ( .A(n2069), .B(n2068), .Z(n2070) );
  NAND U2206 ( .A(n2028), .B(n2027), .Z(n2032) );
  NANDN U2207 ( .A(n2030), .B(n2029), .Z(n2031) );
  AND U2208 ( .A(n2032), .B(n2031), .Z(n2065) );
  NAND U2209 ( .A(y[10]), .B(x[26]), .Z(n2086) );
  NAND U2210 ( .A(y[12]), .B(x[24]), .Z(n2087) );
  XOR U2211 ( .A(n2088), .B(n2087), .Z(n2085) );
  AND U2212 ( .A(y[59]), .B(x[43]), .Z(n2281) );
  NANDN U2213 ( .A(n2033), .B(n2281), .Z(n2037) );
  NAND U2214 ( .A(n2035), .B(n2034), .Z(n2036) );
  NAND U2215 ( .A(n2037), .B(n2036), .Z(n2062) );
  XOR U2216 ( .A(n2063), .B(n2062), .Z(n2064) );
  XOR U2217 ( .A(n2065), .B(n2064), .Z(n2071) );
  XOR U2218 ( .A(n2070), .B(n2071), .Z(n2052) );
  NAND U2219 ( .A(n2039), .B(n2038), .Z(n2043) );
  NAND U2220 ( .A(n2041), .B(n2040), .Z(n2042) );
  AND U2221 ( .A(n2043), .B(n2042), .Z(n2051) );
  NAND U2222 ( .A(n2045), .B(n2044), .Z(n2049) );
  NAND U2223 ( .A(n2047), .B(n2046), .Z(n2048) );
  AND U2224 ( .A(n2049), .B(n2048), .Z(n2050) );
  XOR U2225 ( .A(n2051), .B(n2050), .Z(n2053) );
  XNOR U2226 ( .A(n2052), .B(n2053), .Z(n2058) );
  XOR U2227 ( .A(n2059), .B(n2058), .Z(o[36]) );
  NAND U2228 ( .A(n2051), .B(n2050), .Z(n2055) );
  NAND U2229 ( .A(n2053), .B(n2052), .Z(n2054) );
  AND U2230 ( .A(n2055), .B(n2054), .Z(n2202) );
  NANDN U2231 ( .A(n2057), .B(n2056), .Z(n2061) );
  NAND U2232 ( .A(n2059), .B(n2058), .Z(n2060) );
  AND U2233 ( .A(n2061), .B(n2060), .Z(n2201) );
  XNOR U2234 ( .A(n2202), .B(n2201), .Z(n2204) );
  NAND U2235 ( .A(n2063), .B(n2062), .Z(n2067) );
  NANDN U2236 ( .A(n2065), .B(n2064), .Z(n2066) );
  AND U2237 ( .A(n2067), .B(n2066), .Z(n2120) );
  XNOR U2238 ( .A(n2120), .B(n2119), .Z(n2122) );
  NAND U2239 ( .A(n2073), .B(n2072), .Z(n2076) );
  NAND U2240 ( .A(n2137), .B(n2074), .Z(n2075) );
  NAND U2241 ( .A(n2076), .B(n2075), .Z(n2158) );
  AND U2242 ( .A(x[37]), .B(y[32]), .Z(n2078) );
  NAND U2243 ( .A(x[36]), .B(y[33]), .Z(n2077) );
  XNOR U2244 ( .A(n2078), .B(n2077), .Z(n2180) );
  AND U2245 ( .A(y[12]), .B(x[25]), .Z(n2179) );
  XOR U2246 ( .A(n2180), .B(n2179), .Z(n2156) );
  AND U2247 ( .A(y[59]), .B(x[42]), .Z(n2169) );
  AND U2248 ( .A(y[56]), .B(x[45]), .Z(n2168) );
  XOR U2249 ( .A(n2169), .B(n2168), .Z(n2171) );
  AND U2250 ( .A(y[58]), .B(x[43]), .Z(n2103) );
  AND U2251 ( .A(y[57]), .B(x[44]), .Z(n2280) );
  XOR U2252 ( .A(n2103), .B(n2280), .Z(n2170) );
  XOR U2253 ( .A(n2171), .B(n2170), .Z(n2155) );
  XOR U2254 ( .A(n2156), .B(n2155), .Z(n2157) );
  NAND U2255 ( .A(n2080), .B(n2079), .Z(n2084) );
  NAND U2256 ( .A(n2082), .B(n2081), .Z(n2083) );
  NAND U2257 ( .A(n2084), .B(n2083), .Z(n2184) );
  NAND U2258 ( .A(n2086), .B(n2085), .Z(n2090) );
  AND U2259 ( .A(n2088), .B(n2087), .Z(n2089) );
  ANDN U2260 ( .B(n2090), .A(n2089), .Z(n2183) );
  XNOR U2261 ( .A(n2186), .B(n2185), .Z(n2197) );
  NAND U2262 ( .A(y[35]), .B(x[34]), .Z(n2096) );
  IV U2263 ( .A(n2096), .Z(n2142) );
  AND U2264 ( .A(y[34]), .B(x[33]), .Z(n2091) );
  NAND U2265 ( .A(n2142), .B(n2091), .Z(n2095) );
  NAND U2266 ( .A(n2093), .B(n2092), .Z(n2094) );
  NAND U2267 ( .A(n2095), .B(n2094), .Z(n2128) );
  AND U2268 ( .A(y[8]), .B(x[29]), .Z(n2277) );
  XNOR U2269 ( .A(n2277), .B(n2096), .Z(n2144) );
  AND U2270 ( .A(y[9]), .B(x[28]), .Z(n2143) );
  XOR U2271 ( .A(n2144), .B(n2143), .Z(n2126) );
  AND U2272 ( .A(y[36]), .B(x[33]), .Z(n2310) );
  AND U2273 ( .A(y[13]), .B(x[24]), .Z(n2149) );
  AND U2274 ( .A(y[37]), .B(x[32]), .Z(n2148) );
  XOR U2275 ( .A(n2149), .B(n2148), .Z(n2150) );
  XOR U2276 ( .A(n2310), .B(n2150), .Z(n2125) );
  XOR U2277 ( .A(n2126), .B(n2125), .Z(n2127) );
  AND U2278 ( .A(n2098), .B(n2097), .Z(n2101) );
  NAND U2279 ( .A(n2178), .B(n2099), .Z(n2100) );
  NANDN U2280 ( .A(n2101), .B(n2100), .Z(n2134) );
  AND U2281 ( .A(y[57]), .B(x[42]), .Z(n2102) );
  AND U2282 ( .A(n2103), .B(n2102), .Z(n2139) );
  AND U2283 ( .A(y[60]), .B(x[41]), .Z(n2105) );
  AND U2284 ( .A(x[40]), .B(y[61]), .Z(n2104) );
  XOR U2285 ( .A(n2105), .B(n2104), .Z(n2138) );
  XOR U2286 ( .A(n2139), .B(n2138), .Z(n2132) );
  AND U2287 ( .A(y[10]), .B(x[27]), .Z(n2304) );
  XNOR U2288 ( .A(n2304), .B(n2106), .Z(n2163) );
  AND U2289 ( .A(y[11]), .B(x[26]), .Z(n2162) );
  XOR U2290 ( .A(n2163), .B(n2162), .Z(n2131) );
  XOR U2291 ( .A(n2132), .B(n2131), .Z(n2133) );
  XNOR U2292 ( .A(n2134), .B(n2133), .Z(n2195) );
  XOR U2293 ( .A(n2197), .B(n2198), .Z(n2191) );
  NAND U2294 ( .A(n2108), .B(n2107), .Z(n2112) );
  NAND U2295 ( .A(n2110), .B(n2109), .Z(n2111) );
  NAND U2296 ( .A(n2112), .B(n2111), .Z(n2190) );
  NAND U2297 ( .A(n2114), .B(n2113), .Z(n2118) );
  NAND U2298 ( .A(n2116), .B(n2115), .Z(n2117) );
  NAND U2299 ( .A(n2118), .B(n2117), .Z(n2189) );
  XOR U2300 ( .A(n2191), .B(n2192), .Z(n2121) );
  XNOR U2301 ( .A(n2122), .B(n2121), .Z(n2203) );
  XNOR U2302 ( .A(n2204), .B(n2203), .Z(o[37]) );
  NANDN U2303 ( .A(n2120), .B(n2119), .Z(n2124) );
  NAND U2304 ( .A(n2122), .B(n2121), .Z(n2123) );
  NAND U2305 ( .A(n2124), .B(n2123), .Z(n2210) );
  NAND U2306 ( .A(n2126), .B(n2125), .Z(n2130) );
  NAND U2307 ( .A(n2128), .B(n2127), .Z(n2129) );
  AND U2308 ( .A(n2130), .B(n2129), .Z(n2342) );
  NAND U2309 ( .A(n2132), .B(n2131), .Z(n2136) );
  NAND U2310 ( .A(n2134), .B(n2133), .Z(n2135) );
  AND U2311 ( .A(n2136), .B(n2135), .Z(n2341) );
  XOR U2312 ( .A(n2342), .B(n2341), .Z(n2340) );
  AND U2313 ( .A(y[61]), .B(x[41]), .Z(n2240) );
  NAND U2314 ( .A(n2240), .B(n2137), .Z(n2141) );
  NAND U2315 ( .A(n2139), .B(n2138), .Z(n2140) );
  AND U2316 ( .A(n2141), .B(n2140), .Z(n2334) );
  NAND U2317 ( .A(n2142), .B(n2277), .Z(n2146) );
  NAND U2318 ( .A(n2144), .B(n2143), .Z(n2145) );
  AND U2319 ( .A(n2146), .B(n2145), .Z(n2234) );
  AND U2320 ( .A(y[33]), .B(x[37]), .Z(n2294) );
  AND U2321 ( .A(y[32]), .B(x[38]), .Z(n2296) );
  AND U2322 ( .A(y[14]), .B(x[24]), .Z(n2295) );
  XOR U2323 ( .A(n2296), .B(n2295), .Z(n2293) );
  XNOR U2324 ( .A(n2294), .B(n2293), .Z(n2236) );
  AND U2325 ( .A(y[58]), .B(x[44]), .Z(n2175) );
  NAND U2326 ( .A(x[45]), .B(y[57]), .Z(n2147) );
  XNOR U2327 ( .A(n2175), .B(n2147), .Z(n2284) );
  AND U2328 ( .A(y[56]), .B(x[46]), .Z(n2283) );
  XOR U2329 ( .A(n2284), .B(n2283), .Z(n2282) );
  XNOR U2330 ( .A(n2282), .B(n2281), .Z(n2235) );
  XOR U2331 ( .A(n2234), .B(n2233), .Z(n2333) );
  XOR U2332 ( .A(n2334), .B(n2333), .Z(n2332) );
  NAND U2333 ( .A(n2149), .B(n2148), .Z(n2152) );
  NAND U2334 ( .A(n2310), .B(n2150), .Z(n2151) );
  AND U2335 ( .A(n2152), .B(n2151), .Z(n2219) );
  AND U2336 ( .A(x[29]), .B(y[9]), .Z(n2154) );
  NAND U2337 ( .A(x[30]), .B(y[8]), .Z(n2153) );
  XNOR U2338 ( .A(n2154), .B(n2153), .Z(n2275) );
  AND U2339 ( .A(y[35]), .B(x[35]), .Z(n2274) );
  XNOR U2340 ( .A(n2275), .B(n2274), .Z(n2222) );
  AND U2341 ( .A(y[62]), .B(x[40]), .Z(n2290) );
  AND U2342 ( .A(y[38]), .B(x[32]), .Z(n2289) );
  XOR U2343 ( .A(n2290), .B(n2289), .Z(n2288) );
  AND U2344 ( .A(y[13]), .B(x[25]), .Z(n2287) );
  XNOR U2345 ( .A(n2288), .B(n2287), .Z(n2221) );
  XNOR U2346 ( .A(n2219), .B(n2220), .Z(n2331) );
  XOR U2347 ( .A(n2332), .B(n2331), .Z(n2339) );
  XOR U2348 ( .A(n2340), .B(n2339), .Z(n2364) );
  NAND U2349 ( .A(n2156), .B(n2155), .Z(n2160) );
  NAND U2350 ( .A(n2158), .B(n2157), .Z(n2159) );
  AND U2351 ( .A(n2160), .B(n2159), .Z(n2348) );
  NAND U2352 ( .A(n2161), .B(n2304), .Z(n2165) );
  NAND U2353 ( .A(n2163), .B(n2162), .Z(n2164) );
  AND U2354 ( .A(n2165), .B(n2164), .Z(n2214) );
  AND U2355 ( .A(x[33]), .B(y[37]), .Z(n2167) );
  NAND U2356 ( .A(x[34]), .B(y[36]), .Z(n2166) );
  XNOR U2357 ( .A(n2167), .B(n2166), .Z(n2308) );
  AND U2358 ( .A(y[12]), .B(x[26]), .Z(n2307) );
  XNOR U2359 ( .A(n2308), .B(n2307), .Z(n2216) );
  NAND U2360 ( .A(n2169), .B(n2168), .Z(n2173) );
  NAND U2361 ( .A(n2171), .B(n2170), .Z(n2172) );
  AND U2362 ( .A(n2173), .B(n2172), .Z(n2215) );
  XOR U2363 ( .A(n2214), .B(n2213), .Z(n2347) );
  XOR U2364 ( .A(n2348), .B(n2347), .Z(n2345) );
  AND U2365 ( .A(y[57]), .B(x[43]), .Z(n2174) );
  AND U2366 ( .A(n2175), .B(n2174), .Z(n2242) );
  AND U2367 ( .A(y[60]), .B(x[42]), .Z(n2241) );
  XOR U2368 ( .A(n2242), .B(n2241), .Z(n2239) );
  XNOR U2369 ( .A(n2239), .B(n2240), .Z(n2225) );
  AND U2370 ( .A(x[28]), .B(y[10]), .Z(n2177) );
  NAND U2371 ( .A(x[27]), .B(y[11]), .Z(n2176) );
  XNOR U2372 ( .A(n2177), .B(n2176), .Z(n2302) );
  AND U2373 ( .A(y[34]), .B(x[36]), .Z(n2301) );
  XNOR U2374 ( .A(n2302), .B(n2301), .Z(n2228) );
  NAND U2375 ( .A(n2178), .B(n2294), .Z(n2182) );
  NAND U2376 ( .A(n2180), .B(n2179), .Z(n2181) );
  AND U2377 ( .A(n2182), .B(n2181), .Z(n2227) );
  XOR U2378 ( .A(n2225), .B(n2226), .Z(n2346) );
  XNOR U2379 ( .A(n2345), .B(n2346), .Z(n2366) );
  NAND U2380 ( .A(n2184), .B(n2183), .Z(n2188) );
  NAND U2381 ( .A(n2186), .B(n2185), .Z(n2187) );
  AND U2382 ( .A(n2188), .B(n2187), .Z(n2365) );
  XOR U2383 ( .A(n2366), .B(n2365), .Z(n2363) );
  XNOR U2384 ( .A(n2364), .B(n2363), .Z(n2358) );
  NAND U2385 ( .A(n2190), .B(n2189), .Z(n2194) );
  NAND U2386 ( .A(n2192), .B(n2191), .Z(n2193) );
  NAND U2387 ( .A(n2194), .B(n2193), .Z(n2359) );
  NAND U2388 ( .A(n2196), .B(n2195), .Z(n2200) );
  NANDN U2389 ( .A(n2198), .B(n2197), .Z(n2199) );
  AND U2390 ( .A(n2200), .B(n2199), .Z(n2360) );
  XOR U2391 ( .A(n2359), .B(n2360), .Z(n2357) );
  NANDN U2392 ( .A(n2202), .B(n2201), .Z(n2206) );
  NAND U2393 ( .A(n2204), .B(n2203), .Z(n2205) );
  AND U2394 ( .A(n2206), .B(n2205), .Z(n2207) );
  XOR U2395 ( .A(n2208), .B(n2207), .Z(o[38]) );
  NAND U2396 ( .A(n2208), .B(n2207), .Z(n2212) );
  NAND U2397 ( .A(n2210), .B(n2209), .Z(n2211) );
  AND U2398 ( .A(n2212), .B(n2211), .Z(n2356) );
  NAND U2399 ( .A(n2214), .B(n2213), .Z(n2218) );
  NAND U2400 ( .A(n2216), .B(n2215), .Z(n2217) );
  AND U2401 ( .A(n2218), .B(n2217), .Z(n2330) );
  NANDN U2402 ( .A(n2220), .B(n2219), .Z(n2224) );
  NAND U2403 ( .A(n2222), .B(n2221), .Z(n2223) );
  AND U2404 ( .A(n2224), .B(n2223), .Z(n2232) );
  NANDN U2405 ( .A(n2226), .B(n2225), .Z(n2230) );
  NAND U2406 ( .A(n2228), .B(n2227), .Z(n2229) );
  NAND U2407 ( .A(n2230), .B(n2229), .Z(n2231) );
  XNOR U2408 ( .A(n2232), .B(n2231), .Z(n2328) );
  NAND U2409 ( .A(n2234), .B(n2233), .Z(n2238) );
  NAND U2410 ( .A(n2236), .B(n2235), .Z(n2237) );
  AND U2411 ( .A(n2238), .B(n2237), .Z(n2326) );
  NAND U2412 ( .A(n2240), .B(n2239), .Z(n2244) );
  NAND U2413 ( .A(n2242), .B(n2241), .Z(n2243) );
  AND U2414 ( .A(n2244), .B(n2243), .Z(n2273) );
  AND U2415 ( .A(x[38]), .B(y[33]), .Z(n2249) );
  AND U2416 ( .A(y[37]), .B(x[34]), .Z(n2309) );
  AND U2417 ( .A(x[33]), .B(y[38]), .Z(n2246) );
  NAND U2418 ( .A(x[39]), .B(y[32]), .Z(n2245) );
  XNOR U2419 ( .A(n2246), .B(n2245), .Z(n2247) );
  XNOR U2420 ( .A(n2309), .B(n2247), .Z(n2248) );
  XNOR U2421 ( .A(n2249), .B(n2248), .Z(n2271) );
  AND U2422 ( .A(x[47]), .B(y[56]), .Z(n2251) );
  NAND U2423 ( .A(x[44]), .B(y[59]), .Z(n2250) );
  XNOR U2424 ( .A(n2251), .B(n2250), .Z(n2261) );
  AND U2425 ( .A(x[32]), .B(y[39]), .Z(n2253) );
  NAND U2426 ( .A(x[25]), .B(y[14]), .Z(n2252) );
  XNOR U2427 ( .A(n2253), .B(n2252), .Z(n2257) );
  AND U2428 ( .A(x[40]), .B(y[63]), .Z(n2255) );
  NAND U2429 ( .A(x[27]), .B(y[12]), .Z(n2254) );
  XNOR U2430 ( .A(n2255), .B(n2254), .Z(n2256) );
  XOR U2431 ( .A(n2257), .B(n2256), .Z(n2259) );
  AND U2432 ( .A(y[11]), .B(x[28]), .Z(n2303) );
  AND U2433 ( .A(y[9]), .B(x[30]), .Z(n2276) );
  XNOR U2434 ( .A(n2303), .B(n2276), .Z(n2258) );
  XNOR U2435 ( .A(n2259), .B(n2258), .Z(n2260) );
  XOR U2436 ( .A(n2261), .B(n2260), .Z(n2269) );
  AND U2437 ( .A(x[41]), .B(y[62]), .Z(n2263) );
  NAND U2438 ( .A(x[26]), .B(y[13]), .Z(n2262) );
  XNOR U2439 ( .A(n2263), .B(n2262), .Z(n2267) );
  AND U2440 ( .A(x[42]), .B(y[61]), .Z(n2265) );
  NAND U2441 ( .A(x[35]), .B(y[36]), .Z(n2264) );
  XNOR U2442 ( .A(n2265), .B(n2264), .Z(n2266) );
  XNOR U2443 ( .A(n2267), .B(n2266), .Z(n2268) );
  XNOR U2444 ( .A(n2269), .B(n2268), .Z(n2270) );
  XNOR U2445 ( .A(n2271), .B(n2270), .Z(n2272) );
  XNOR U2446 ( .A(n2273), .B(n2272), .Z(n2324) );
  NAND U2447 ( .A(n2275), .B(n2274), .Z(n2279) );
  NAND U2448 ( .A(n2277), .B(n2276), .Z(n2278) );
  AND U2449 ( .A(n2279), .B(n2278), .Z(n2322) );
  NAND U2450 ( .A(n2282), .B(n2281), .Z(n2286) );
  NAND U2451 ( .A(n2284), .B(n2283), .Z(n2285) );
  AND U2452 ( .A(n2286), .B(n2285), .Z(n2318) );
  NAND U2453 ( .A(n2288), .B(n2287), .Z(n2292) );
  NAND U2454 ( .A(n2290), .B(n2289), .Z(n2291) );
  AND U2455 ( .A(n2292), .B(n2291), .Z(n2300) );
  NAND U2456 ( .A(n2294), .B(n2293), .Z(n2298) );
  NAND U2457 ( .A(n2296), .B(n2295), .Z(n2297) );
  NAND U2458 ( .A(n2298), .B(n2297), .Z(n2299) );
  XNOR U2459 ( .A(n2300), .B(n2299), .Z(n2316) );
  NAND U2460 ( .A(n2302), .B(n2301), .Z(n2306) );
  NAND U2461 ( .A(n2304), .B(n2303), .Z(n2305) );
  AND U2462 ( .A(n2306), .B(n2305), .Z(n2314) );
  NAND U2463 ( .A(n2308), .B(n2307), .Z(n2312) );
  NAND U2464 ( .A(n2310), .B(n2309), .Z(n2311) );
  NAND U2465 ( .A(n2312), .B(n2311), .Z(n2313) );
  XNOR U2466 ( .A(n2314), .B(n2313), .Z(n2315) );
  XNOR U2467 ( .A(n2316), .B(n2315), .Z(n2317) );
  XNOR U2468 ( .A(n2318), .B(n2317), .Z(n2319) );
  XNOR U2469 ( .A(n2320), .B(n2319), .Z(n2321) );
  XNOR U2470 ( .A(n2322), .B(n2321), .Z(n2323) );
  XNOR U2471 ( .A(n2324), .B(n2323), .Z(n2325) );
  XNOR U2472 ( .A(n2326), .B(n2325), .Z(n2327) );
  XNOR U2473 ( .A(n2328), .B(n2327), .Z(n2329) );
  XNOR U2474 ( .A(n2330), .B(n2329), .Z(n2338) );
  NAND U2475 ( .A(n2332), .B(n2331), .Z(n2336) );
  NAND U2476 ( .A(n2334), .B(n2333), .Z(n2335) );
  NAND U2477 ( .A(n2336), .B(n2335), .Z(n2337) );
  XNOR U2478 ( .A(n2338), .B(n2337), .Z(n2354) );
  NAND U2479 ( .A(n2340), .B(n2339), .Z(n2344) );
  NAND U2480 ( .A(n2342), .B(n2341), .Z(n2343) );
  AND U2481 ( .A(n2344), .B(n2343), .Z(n2352) );
  NANDN U2482 ( .A(n2346), .B(n2345), .Z(n2350) );
  NAND U2483 ( .A(n2348), .B(n2347), .Z(n2349) );
  NAND U2484 ( .A(n2350), .B(n2349), .Z(n2351) );
  XNOR U2485 ( .A(n2352), .B(n2351), .Z(n2353) );
  XNOR U2486 ( .A(n2354), .B(n2353), .Z(n2355) );
  XNOR U2487 ( .A(n2356), .B(n2355), .Z(n2372) );
  NAND U2488 ( .A(n2358), .B(n2357), .Z(n2362) );
  NAND U2489 ( .A(n2360), .B(n2359), .Z(n2361) );
  AND U2490 ( .A(n2362), .B(n2361), .Z(n2370) );
  NAND U2491 ( .A(n2364), .B(n2363), .Z(n2368) );
  NAND U2492 ( .A(n2366), .B(n2365), .Z(n2367) );
  NAND U2493 ( .A(n2368), .B(n2367), .Z(n2369) );
  XNOR U2494 ( .A(n2370), .B(n2369), .Z(n2371) );
  XNOR U2495 ( .A(n2372), .B(n2371), .Z(o[39]) );
  AND U2496 ( .A(y[40]), .B(x[32]), .Z(n2374) );
  NAND U2497 ( .A(y[16]), .B(x[24]), .Z(n2373) );
  XNOR U2498 ( .A(n2374), .B(n2373), .Z(n2375) );
  NAND U2499 ( .A(y[64]), .B(x[40]), .Z(n2462) );
  XNOR U2500 ( .A(n2375), .B(n2462), .Z(o[40]) );
  AND U2501 ( .A(y[40]), .B(x[33]), .Z(n2449) );
  AND U2502 ( .A(y[41]), .B(x[32]), .Z(n2385) );
  AND U2503 ( .A(y[64]), .B(x[41]), .Z(n2384) );
  XOR U2504 ( .A(n2385), .B(n2384), .Z(n2386) );
  XNOR U2505 ( .A(n2449), .B(n2386), .Z(n2381) );
  NANDN U2506 ( .A(n2374), .B(n2373), .Z(n2377) );
  NAND U2507 ( .A(n2375), .B(n2462), .Z(n2376) );
  AND U2508 ( .A(n2377), .B(n2376), .Z(n2379) );
  AND U2509 ( .A(y[17]), .B(x[24]), .Z(n2413) );
  AND U2510 ( .A(y[65]), .B(x[40]), .Z(n2421) );
  AND U2511 ( .A(y[16]), .B(x[25]), .Z(n2389) );
  XOR U2512 ( .A(n2421), .B(n2389), .Z(n2390) );
  XNOR U2513 ( .A(n2413), .B(n2390), .Z(n2380) );
  XNOR U2514 ( .A(n2379), .B(n2380), .Z(n2378) );
  XNOR U2515 ( .A(n2381), .B(n2378), .Z(o[41]) );
  AND U2516 ( .A(x[25]), .B(y[17]), .Z(n2383) );
  NAND U2517 ( .A(x[24]), .B(y[18]), .Z(n2382) );
  XNOR U2518 ( .A(n2383), .B(n2382), .Z(n2415) );
  AND U2519 ( .A(y[40]), .B(x[34]), .Z(n2414) );
  XOR U2520 ( .A(n2415), .B(n2414), .Z(n2428) );
  AND U2521 ( .A(y[42]), .B(x[32]), .Z(n2426) );
  NAND U2522 ( .A(y[41]), .B(x[33]), .Z(n2425) );
  XNOR U2523 ( .A(n2426), .B(n2425), .Z(n2427) );
  XNOR U2524 ( .A(n2428), .B(n2427), .Z(n2400) );
  XNOR U2525 ( .A(n2401), .B(n2400), .Z(n2403) );
  NAND U2526 ( .A(n2385), .B(n2384), .Z(n2388) );
  NAND U2527 ( .A(n2449), .B(n2386), .Z(n2387) );
  NAND U2528 ( .A(n2388), .B(n2387), .Z(n2396) );
  NAND U2529 ( .A(n2421), .B(n2389), .Z(n2392) );
  NAND U2530 ( .A(n2413), .B(n2390), .Z(n2391) );
  NAND U2531 ( .A(n2392), .B(n2391), .Z(n2394) );
  AND U2532 ( .A(y[16]), .B(x[26]), .Z(n2441) );
  NAND U2533 ( .A(y[64]), .B(x[42]), .Z(n2406) );
  XNOR U2534 ( .A(n2441), .B(n2406), .Z(n2408) );
  AND U2535 ( .A(x[41]), .B(y[65]), .Z(n2455) );
  NAND U2536 ( .A(x[40]), .B(y[66]), .Z(n2393) );
  XNOR U2537 ( .A(n2455), .B(n2393), .Z(n2407) );
  XOR U2538 ( .A(n2408), .B(n2407), .Z(n2395) );
  XNOR U2539 ( .A(n2394), .B(n2395), .Z(n2397) );
  XOR U2540 ( .A(n2396), .B(n2397), .Z(n2402) );
  XNOR U2541 ( .A(n2403), .B(n2402), .Z(o[42]) );
  NAND U2542 ( .A(n2395), .B(n2394), .Z(n2399) );
  NANDN U2543 ( .A(n2397), .B(n2396), .Z(n2398) );
  AND U2544 ( .A(n2399), .B(n2398), .Z(n2436) );
  NANDN U2545 ( .A(n2401), .B(n2400), .Z(n2405) );
  NAND U2546 ( .A(n2403), .B(n2402), .Z(n2404) );
  AND U2547 ( .A(n2405), .B(n2404), .Z(n2435) );
  XNOR U2548 ( .A(n2436), .B(n2435), .Z(n2438) );
  NANDN U2549 ( .A(n2406), .B(n2441), .Z(n2410) );
  NAND U2550 ( .A(n2408), .B(n2407), .Z(n2409) );
  NAND U2551 ( .A(n2410), .B(n2409), .Z(n2469) );
  AND U2552 ( .A(y[43]), .B(x[32]), .Z(n2456) );
  AND U2553 ( .A(y[18]), .B(x[25]), .Z(n2457) );
  NAND U2554 ( .A(y[19]), .B(x[24]), .Z(n2459) );
  XNOR U2555 ( .A(n2458), .B(n2459), .Z(n2468) );
  AND U2556 ( .A(x[35]), .B(y[40]), .Z(n2412) );
  NAND U2557 ( .A(x[33]), .B(y[42]), .Z(n2411) );
  XNOR U2558 ( .A(n2412), .B(n2411), .Z(n2451) );
  AND U2559 ( .A(y[41]), .B(x[34]), .Z(n2450) );
  XOR U2560 ( .A(n2451), .B(n2450), .Z(n2467) );
  XOR U2561 ( .A(n2468), .B(n2467), .Z(n2470) );
  XOR U2562 ( .A(n2469), .B(n2470), .Z(n2432) );
  NAND U2563 ( .A(n2457), .B(n2413), .Z(n2417) );
  NAND U2564 ( .A(n2415), .B(n2414), .Z(n2416) );
  NAND U2565 ( .A(n2417), .B(n2416), .Z(n2475) );
  AND U2566 ( .A(x[26]), .B(y[17]), .Z(n2419) );
  NAND U2567 ( .A(x[27]), .B(y[16]), .Z(n2418) );
  XNOR U2568 ( .A(n2419), .B(n2418), .Z(n2442) );
  AND U2569 ( .A(y[66]), .B(x[41]), .Z(n2420) );
  NAND U2570 ( .A(n2421), .B(n2420), .Z(n2443) );
  XNOR U2571 ( .A(n2442), .B(n2443), .Z(n2474) );
  AND U2572 ( .A(x[43]), .B(y[64]), .Z(n2423) );
  NAND U2573 ( .A(x[40]), .B(y[67]), .Z(n2422) );
  XNOR U2574 ( .A(n2423), .B(n2422), .Z(n2464) );
  AND U2575 ( .A(x[42]), .B(y[65]), .Z(n2510) );
  NAND U2576 ( .A(x[41]), .B(y[66]), .Z(n2424) );
  XNOR U2577 ( .A(n2510), .B(n2424), .Z(n2463) );
  XOR U2578 ( .A(n2464), .B(n2463), .Z(n2473) );
  XOR U2579 ( .A(n2474), .B(n2473), .Z(n2476) );
  XNOR U2580 ( .A(n2475), .B(n2476), .Z(n2431) );
  XNOR U2581 ( .A(n2432), .B(n2431), .Z(n2433) );
  NANDN U2582 ( .A(n2426), .B(n2425), .Z(n2430) );
  NANDN U2583 ( .A(n2428), .B(n2427), .Z(n2429) );
  NAND U2584 ( .A(n2430), .B(n2429), .Z(n2434) );
  XNOR U2585 ( .A(n2433), .B(n2434), .Z(n2437) );
  XOR U2586 ( .A(n2438), .B(n2437), .Z(o[43]) );
  NANDN U2587 ( .A(n2436), .B(n2435), .Z(n2440) );
  NAND U2588 ( .A(n2438), .B(n2437), .Z(n2439) );
  NAND U2589 ( .A(n2440), .B(n2439), .Z(n2537) );
  XNOR U2590 ( .A(n2538), .B(n2537), .Z(n2540) );
  NAND U2591 ( .A(y[17]), .B(x[27]), .Z(n2496) );
  NANDN U2592 ( .A(n2496), .B(n2441), .Z(n2445) );
  NANDN U2593 ( .A(n2443), .B(n2442), .Z(n2444) );
  AND U2594 ( .A(n2445), .B(n2444), .Z(n2520) );
  AND U2595 ( .A(y[65]), .B(x[43]), .Z(n2588) );
  NAND U2596 ( .A(x[42]), .B(y[66]), .Z(n2446) );
  XNOR U2597 ( .A(n2588), .B(n2446), .Z(n2479) );
  NAND U2598 ( .A(y[67]), .B(x[41]), .Z(n2480) );
  XNOR U2599 ( .A(n2479), .B(n2480), .Z(n2481) );
  NAND U2600 ( .A(y[64]), .B(x[44]), .Z(n2482) );
  XNOR U2601 ( .A(n2481), .B(n2482), .Z(n2518) );
  AND U2602 ( .A(x[33]), .B(y[43]), .Z(n2448) );
  NAND U2603 ( .A(x[34]), .B(y[42]), .Z(n2447) );
  XNOR U2604 ( .A(n2448), .B(n2447), .Z(n2500) );
  NAND U2605 ( .A(y[41]), .B(x[35]), .Z(n2501) );
  XOR U2606 ( .A(n2500), .B(n2501), .Z(n2517) );
  XNOR U2607 ( .A(n2518), .B(n2517), .Z(n2519) );
  XNOR U2608 ( .A(n2520), .B(n2519), .Z(n2521) );
  AND U2609 ( .A(y[42]), .B(x[35]), .Z(n2595) );
  NAND U2610 ( .A(n2595), .B(n2449), .Z(n2453) );
  NAND U2611 ( .A(n2451), .B(n2450), .Z(n2452) );
  AND U2612 ( .A(n2453), .B(n2452), .Z(n2516) );
  AND U2613 ( .A(y[68]), .B(x[40]), .Z(n2562) );
  AND U2614 ( .A(y[66]), .B(x[42]), .Z(n2454) );
  AND U2615 ( .A(n2455), .B(n2454), .Z(n2485) );
  NAND U2616 ( .A(y[16]), .B(x[28]), .Z(n2486) );
  XNOR U2617 ( .A(n2485), .B(n2486), .Z(n2487) );
  XOR U2618 ( .A(n2562), .B(n2487), .Z(n2514) );
  AND U2619 ( .A(y[44]), .B(x[32]), .Z(n2504) );
  AND U2620 ( .A(y[40]), .B(x[36]), .Z(n2582) );
  NAND U2621 ( .A(y[19]), .B(x[25]), .Z(n2506) );
  XOR U2622 ( .A(n2505), .B(n2506), .Z(n2513) );
  XNOR U2623 ( .A(n2514), .B(n2513), .Z(n2515) );
  XOR U2624 ( .A(n2516), .B(n2515), .Z(n2522) );
  XNOR U2625 ( .A(n2521), .B(n2522), .Z(n2524) );
  NAND U2626 ( .A(n2457), .B(n2456), .Z(n2461) );
  NANDN U2627 ( .A(n2459), .B(n2458), .Z(n2460) );
  NAND U2628 ( .A(n2461), .B(n2460), .Z(n2527) );
  AND U2629 ( .A(y[18]), .B(x[26]), .Z(n2494) );
  NAND U2630 ( .A(y[20]), .B(x[24]), .Z(n2495) );
  XOR U2631 ( .A(n2496), .B(n2495), .Z(n2493) );
  XOR U2632 ( .A(n2494), .B(n2493), .Z(n2526) );
  AND U2633 ( .A(y[67]), .B(x[43]), .Z(n2735) );
  NANDN U2634 ( .A(n2462), .B(n2735), .Z(n2466) );
  NAND U2635 ( .A(n2464), .B(n2463), .Z(n2465) );
  NAND U2636 ( .A(n2466), .B(n2465), .Z(n2525) );
  XOR U2637 ( .A(n2526), .B(n2525), .Z(n2528) );
  XNOR U2638 ( .A(n2527), .B(n2528), .Z(n2523) );
  XNOR U2639 ( .A(n2524), .B(n2523), .Z(n2534) );
  NAND U2640 ( .A(n2468), .B(n2467), .Z(n2472) );
  NAND U2641 ( .A(n2470), .B(n2469), .Z(n2471) );
  AND U2642 ( .A(n2472), .B(n2471), .Z(n2532) );
  NAND U2643 ( .A(n2474), .B(n2473), .Z(n2478) );
  NAND U2644 ( .A(n2476), .B(n2475), .Z(n2477) );
  AND U2645 ( .A(n2478), .B(n2477), .Z(n2531) );
  XOR U2646 ( .A(n2532), .B(n2531), .Z(n2533) );
  XOR U2647 ( .A(n2534), .B(n2533), .Z(n2539) );
  XOR U2648 ( .A(n2540), .B(n2539), .Z(o[44]) );
  NANDN U2649 ( .A(n2480), .B(n2479), .Z(n2484) );
  NANDN U2650 ( .A(n2482), .B(n2481), .Z(n2483) );
  NAND U2651 ( .A(n2484), .B(n2483), .Z(n2576) );
  NANDN U2652 ( .A(n2486), .B(n2485), .Z(n2489) );
  NAND U2653 ( .A(n2562), .B(n2487), .Z(n2488) );
  NAND U2654 ( .A(n2489), .B(n2488), .Z(n2591) );
  AND U2655 ( .A(x[36]), .B(y[41]), .Z(n2491) );
  NAND U2656 ( .A(x[37]), .B(y[40]), .Z(n2490) );
  XNOR U2657 ( .A(n2491), .B(n2490), .Z(n2584) );
  AND U2658 ( .A(y[20]), .B(x[25]), .Z(n2583) );
  XOR U2659 ( .A(n2584), .B(n2583), .Z(n2590) );
  AND U2660 ( .A(y[67]), .B(x[42]), .Z(n2603) );
  AND U2661 ( .A(y[64]), .B(x[45]), .Z(n2602) );
  XOR U2662 ( .A(n2603), .B(n2602), .Z(n2605) );
  AND U2663 ( .A(y[65]), .B(x[44]), .Z(n2743) );
  NAND U2664 ( .A(x[43]), .B(y[66]), .Z(n2492) );
  XNOR U2665 ( .A(n2743), .B(n2492), .Z(n2604) );
  XOR U2666 ( .A(n2605), .B(n2604), .Z(n2589) );
  XOR U2667 ( .A(n2590), .B(n2589), .Z(n2592) );
  XOR U2668 ( .A(n2591), .B(n2592), .Z(n2575) );
  NANDN U2669 ( .A(n2494), .B(n2493), .Z(n2498) );
  AND U2670 ( .A(n2496), .B(n2495), .Z(n2497) );
  ANDN U2671 ( .B(n2498), .A(n2497), .Z(n2574) );
  XOR U2672 ( .A(n2575), .B(n2574), .Z(n2577) );
  XNOR U2673 ( .A(n2576), .B(n2577), .Z(n2616) );
  AND U2674 ( .A(y[42]), .B(x[33]), .Z(n2499) );
  AND U2675 ( .A(y[43]), .B(x[34]), .Z(n2567) );
  NAND U2676 ( .A(n2499), .B(n2567), .Z(n2503) );
  NANDN U2677 ( .A(n2501), .B(n2500), .Z(n2502) );
  NAND U2678 ( .A(n2503), .B(n2502), .Z(n2545) );
  AND U2679 ( .A(y[16]), .B(x[29]), .Z(n2676) );
  XOR U2680 ( .A(n2567), .B(n2676), .Z(n2569) );
  AND U2681 ( .A(y[17]), .B(x[28]), .Z(n2568) );
  XOR U2682 ( .A(n2569), .B(n2568), .Z(n2544) );
  AND U2683 ( .A(y[21]), .B(x[24]), .Z(n2556) );
  AND U2684 ( .A(y[45]), .B(x[32]), .Z(n2555) );
  XOR U2685 ( .A(n2556), .B(n2555), .Z(n2557) );
  AND U2686 ( .A(y[44]), .B(x[33]), .Z(n2683) );
  XOR U2687 ( .A(n2557), .B(n2683), .Z(n2543) );
  XOR U2688 ( .A(n2544), .B(n2543), .Z(n2546) );
  XNOR U2689 ( .A(n2545), .B(n2546), .Z(n2615) );
  NAND U2690 ( .A(n2582), .B(n2504), .Z(n2508) );
  NANDN U2691 ( .A(n2506), .B(n2505), .Z(n2507) );
  NAND U2692 ( .A(n2508), .B(n2507), .Z(n2551) );
  AND U2693 ( .A(y[66]), .B(x[43]), .Z(n2509) );
  AND U2694 ( .A(n2510), .B(n2509), .Z(n2564) );
  AND U2695 ( .A(y[68]), .B(x[41]), .Z(n2512) );
  AND U2696 ( .A(x[40]), .B(y[69]), .Z(n2511) );
  XOR U2697 ( .A(n2512), .B(n2511), .Z(n2563) );
  XOR U2698 ( .A(n2564), .B(n2563), .Z(n2550) );
  AND U2699 ( .A(y[18]), .B(x[27]), .Z(n2747) );
  XOR U2700 ( .A(n2595), .B(n2747), .Z(n2597) );
  AND U2701 ( .A(y[19]), .B(x[26]), .Z(n2596) );
  XOR U2702 ( .A(n2597), .B(n2596), .Z(n2549) );
  XOR U2703 ( .A(n2550), .B(n2549), .Z(n2552) );
  XNOR U2704 ( .A(n2551), .B(n2552), .Z(n2614) );
  XOR U2705 ( .A(n2615), .B(n2614), .Z(n2617) );
  XNOR U2706 ( .A(n2616), .B(n2617), .Z(n2610) );
  XOR U2707 ( .A(n2609), .B(n2608), .Z(n2611) );
  XNOR U2708 ( .A(n2610), .B(n2611), .Z(n2622) );
  NAND U2709 ( .A(n2526), .B(n2525), .Z(n2530) );
  NAND U2710 ( .A(n2528), .B(n2527), .Z(n2529) );
  NAND U2711 ( .A(n2530), .B(n2529), .Z(n2621) );
  XNOR U2712 ( .A(n2620), .B(n2621), .Z(n2623) );
  XNOR U2713 ( .A(n2622), .B(n2623), .Z(n2627) );
  NAND U2714 ( .A(n2532), .B(n2531), .Z(n2536) );
  NANDN U2715 ( .A(n2534), .B(n2533), .Z(n2535) );
  AND U2716 ( .A(n2536), .B(n2535), .Z(n2625) );
  NANDN U2717 ( .A(n2538), .B(n2537), .Z(n2542) );
  NAND U2718 ( .A(n2540), .B(n2539), .Z(n2541) );
  AND U2719 ( .A(n2542), .B(n2541), .Z(n2624) );
  XNOR U2720 ( .A(n2625), .B(n2624), .Z(n2626) );
  XNOR U2721 ( .A(n2627), .B(n2626), .Z(o[45]) );
  NAND U2722 ( .A(n2544), .B(n2543), .Z(n2548) );
  NAND U2723 ( .A(n2546), .B(n2545), .Z(n2547) );
  AND U2724 ( .A(n2548), .B(n2547), .Z(n2639) );
  NAND U2725 ( .A(n2550), .B(n2549), .Z(n2554) );
  NAND U2726 ( .A(n2552), .B(n2551), .Z(n2553) );
  AND U2727 ( .A(n2554), .B(n2553), .Z(n2638) );
  XOR U2728 ( .A(n2639), .B(n2638), .Z(n2637) );
  NAND U2729 ( .A(n2556), .B(n2555), .Z(n2559) );
  NAND U2730 ( .A(n2557), .B(n2683), .Z(n2558) );
  AND U2731 ( .A(n2559), .B(n2558), .Z(n2642) );
  AND U2732 ( .A(x[29]), .B(y[17]), .Z(n2561) );
  NAND U2733 ( .A(x[30]), .B(y[16]), .Z(n2560) );
  XNOR U2734 ( .A(n2561), .B(n2560), .Z(n2675) );
  AND U2735 ( .A(y[43]), .B(x[35]), .Z(n2674) );
  XNOR U2736 ( .A(n2675), .B(n2674), .Z(n2645) );
  AND U2737 ( .A(y[21]), .B(x[25]), .Z(n2669) );
  AND U2738 ( .A(y[70]), .B(x[40]), .Z(n2671) );
  AND U2739 ( .A(y[46]), .B(x[32]), .Z(n2670) );
  XOR U2740 ( .A(n2671), .B(n2670), .Z(n2668) );
  XNOR U2741 ( .A(n2669), .B(n2668), .Z(n2644) );
  XNOR U2742 ( .A(n2642), .B(n2643), .Z(n2768) );
  AND U2743 ( .A(y[69]), .B(x[41]), .Z(n2718) );
  NAND U2744 ( .A(n2562), .B(n2718), .Z(n2566) );
  NAND U2745 ( .A(n2564), .B(n2563), .Z(n2565) );
  AND U2746 ( .A(n2566), .B(n2565), .Z(n2770) );
  NAND U2747 ( .A(n2567), .B(n2676), .Z(n2571) );
  NAND U2748 ( .A(n2569), .B(n2568), .Z(n2570) );
  AND U2749 ( .A(n2571), .B(n2570), .Z(n2663) );
  AND U2750 ( .A(y[41]), .B(x[37]), .Z(n2687) );
  AND U2751 ( .A(y[40]), .B(x[38]), .Z(n2689) );
  AND U2752 ( .A(y[22]), .B(x[24]), .Z(n2688) );
  XOR U2753 ( .A(n2689), .B(n2688), .Z(n2686) );
  XNOR U2754 ( .A(n2687), .B(n2686), .Z(n2665) );
  AND U2755 ( .A(x[45]), .B(y[65]), .Z(n2573) );
  NAND U2756 ( .A(x[44]), .B(y[66]), .Z(n2572) );
  XNOR U2757 ( .A(n2573), .B(n2572), .Z(n2738) );
  AND U2758 ( .A(y[64]), .B(x[46]), .Z(n2737) );
  XOR U2759 ( .A(n2738), .B(n2737), .Z(n2736) );
  XNOR U2760 ( .A(n2736), .B(n2735), .Z(n2664) );
  XOR U2761 ( .A(n2663), .B(n2662), .Z(n2769) );
  XOR U2762 ( .A(n2770), .B(n2769), .Z(n2767) );
  XOR U2763 ( .A(n2768), .B(n2767), .Z(n2636) );
  XOR U2764 ( .A(n2637), .B(n2636), .Z(n2786) );
  NAND U2765 ( .A(n2575), .B(n2574), .Z(n2579) );
  NAND U2766 ( .A(n2577), .B(n2576), .Z(n2578) );
  AND U2767 ( .A(n2579), .B(n2578), .Z(n2788) );
  AND U2768 ( .A(x[28]), .B(y[18]), .Z(n2581) );
  NAND U2769 ( .A(x[27]), .B(y[19]), .Z(n2580) );
  XNOR U2770 ( .A(n2581), .B(n2580), .Z(n2745) );
  AND U2771 ( .A(y[42]), .B(x[36]), .Z(n2744) );
  XNOR U2772 ( .A(n2745), .B(n2744), .Z(n2657) );
  NAND U2773 ( .A(n2582), .B(n2687), .Z(n2586) );
  NAND U2774 ( .A(n2584), .B(n2583), .Z(n2585) );
  AND U2775 ( .A(n2586), .B(n2585), .Z(n2656) );
  AND U2776 ( .A(y[66]), .B(x[44]), .Z(n2587) );
  AND U2777 ( .A(n2588), .B(n2587), .Z(n2720) );
  AND U2778 ( .A(y[68]), .B(x[42]), .Z(n2719) );
  XOR U2779 ( .A(n2720), .B(n2719), .Z(n2717) );
  XNOR U2780 ( .A(n2718), .B(n2717), .Z(n2655) );
  NAND U2781 ( .A(n2590), .B(n2589), .Z(n2594) );
  NAND U2782 ( .A(n2592), .B(n2591), .Z(n2593) );
  AND U2783 ( .A(n2594), .B(n2593), .Z(n2764) );
  NAND U2784 ( .A(n2595), .B(n2747), .Z(n2599) );
  NAND U2785 ( .A(n2597), .B(n2596), .Z(n2598) );
  AND U2786 ( .A(n2599), .B(n2598), .Z(n2649) );
  AND U2787 ( .A(x[34]), .B(y[44]), .Z(n2601) );
  NAND U2788 ( .A(x[33]), .B(y[45]), .Z(n2600) );
  XNOR U2789 ( .A(n2601), .B(n2600), .Z(n2682) );
  AND U2790 ( .A(y[20]), .B(x[26]), .Z(n2681) );
  XNOR U2791 ( .A(n2682), .B(n2681), .Z(n2651) );
  NAND U2792 ( .A(n2603), .B(n2602), .Z(n2607) );
  NAND U2793 ( .A(n2605), .B(n2604), .Z(n2606) );
  AND U2794 ( .A(n2607), .B(n2606), .Z(n2650) );
  XOR U2795 ( .A(n2649), .B(n2648), .Z(n2763) );
  XOR U2796 ( .A(n2764), .B(n2763), .Z(n2761) );
  XOR U2797 ( .A(n2762), .B(n2761), .Z(n2787) );
  XOR U2798 ( .A(n2788), .B(n2787), .Z(n2785) );
  XOR U2799 ( .A(n2786), .B(n2785), .Z(n2631) );
  NANDN U2800 ( .A(n2609), .B(n2608), .Z(n2613) );
  NANDN U2801 ( .A(n2611), .B(n2610), .Z(n2612) );
  NAND U2802 ( .A(n2613), .B(n2612), .Z(n2633) );
  NAND U2803 ( .A(n2615), .B(n2614), .Z(n2619) );
  NAND U2804 ( .A(n2617), .B(n2616), .Z(n2618) );
  AND U2805 ( .A(n2619), .B(n2618), .Z(n2632) );
  XOR U2806 ( .A(n2631), .B(n2630), .Z(n2782) );
  XOR U2807 ( .A(n2782), .B(n2781), .Z(n2780) );
  NANDN U2808 ( .A(n2625), .B(n2624), .Z(n2629) );
  NAND U2809 ( .A(n2627), .B(n2626), .Z(n2628) );
  NAND U2810 ( .A(n2629), .B(n2628), .Z(n2779) );
  XNOR U2811 ( .A(n2780), .B(n2779), .Z(o[46]) );
  NANDN U2812 ( .A(n2631), .B(n2630), .Z(n2635) );
  NAND U2813 ( .A(n2633), .B(n2632), .Z(n2634) );
  AND U2814 ( .A(n2635), .B(n2634), .Z(n2796) );
  NAND U2815 ( .A(n2637), .B(n2636), .Z(n2641) );
  NAND U2816 ( .A(n2639), .B(n2638), .Z(n2640) );
  AND U2817 ( .A(n2641), .B(n2640), .Z(n2778) );
  NANDN U2818 ( .A(n2643), .B(n2642), .Z(n2647) );
  NAND U2819 ( .A(n2645), .B(n2644), .Z(n2646) );
  AND U2820 ( .A(n2647), .B(n2646), .Z(n2760) );
  NAND U2821 ( .A(n2649), .B(n2648), .Z(n2653) );
  NAND U2822 ( .A(n2651), .B(n2650), .Z(n2652) );
  AND U2823 ( .A(n2653), .B(n2652), .Z(n2661) );
  NAND U2824 ( .A(n2655), .B(n2654), .Z(n2659) );
  NAND U2825 ( .A(n2657), .B(n2656), .Z(n2658) );
  NAND U2826 ( .A(n2659), .B(n2658), .Z(n2660) );
  XNOR U2827 ( .A(n2661), .B(n2660), .Z(n2758) );
  NAND U2828 ( .A(n2663), .B(n2662), .Z(n2667) );
  NAND U2829 ( .A(n2665), .B(n2664), .Z(n2666) );
  AND U2830 ( .A(n2667), .B(n2666), .Z(n2756) );
  NAND U2831 ( .A(n2669), .B(n2668), .Z(n2673) );
  NAND U2832 ( .A(n2671), .B(n2670), .Z(n2672) );
  AND U2833 ( .A(n2673), .B(n2672), .Z(n2680) );
  NAND U2834 ( .A(n2675), .B(n2674), .Z(n2678) );
  AND U2835 ( .A(y[17]), .B(x[30]), .Z(n2748) );
  NAND U2836 ( .A(n2676), .B(n2748), .Z(n2677) );
  NAND U2837 ( .A(n2678), .B(n2677), .Z(n2679) );
  XNOR U2838 ( .A(n2680), .B(n2679), .Z(n2695) );
  NAND U2839 ( .A(n2682), .B(n2681), .Z(n2685) );
  AND U2840 ( .A(y[45]), .B(x[34]), .Z(n2704) );
  NAND U2841 ( .A(n2683), .B(n2704), .Z(n2684) );
  AND U2842 ( .A(n2685), .B(n2684), .Z(n2693) );
  NAND U2843 ( .A(n2687), .B(n2686), .Z(n2691) );
  NAND U2844 ( .A(n2689), .B(n2688), .Z(n2690) );
  NAND U2845 ( .A(n2691), .B(n2690), .Z(n2692) );
  XNOR U2846 ( .A(n2693), .B(n2692), .Z(n2694) );
  XOR U2847 ( .A(n2695), .B(n2694), .Z(n2734) );
  AND U2848 ( .A(x[33]), .B(y[46]), .Z(n2697) );
  NAND U2849 ( .A(x[39]), .B(y[40]), .Z(n2696) );
  XNOR U2850 ( .A(n2697), .B(n2696), .Z(n2708) );
  AND U2851 ( .A(x[31]), .B(y[16]), .Z(n2699) );
  NAND U2852 ( .A(x[43]), .B(y[68]), .Z(n2698) );
  XNOR U2853 ( .A(n2699), .B(n2698), .Z(n2703) );
  AND U2854 ( .A(x[24]), .B(y[23]), .Z(n2701) );
  NAND U2855 ( .A(x[29]), .B(y[18]), .Z(n2700) );
  XNOR U2856 ( .A(n2701), .B(n2700), .Z(n2702) );
  XOR U2857 ( .A(n2703), .B(n2702), .Z(n2706) );
  AND U2858 ( .A(y[19]), .B(x[28]), .Z(n2746) );
  XNOR U2859 ( .A(n2746), .B(n2704), .Z(n2705) );
  XNOR U2860 ( .A(n2706), .B(n2705), .Z(n2707) );
  XOR U2861 ( .A(n2708), .B(n2707), .Z(n2716) );
  AND U2862 ( .A(x[32]), .B(y[47]), .Z(n2710) );
  NAND U2863 ( .A(x[36]), .B(y[43]), .Z(n2709) );
  XNOR U2864 ( .A(n2710), .B(n2709), .Z(n2714) );
  AND U2865 ( .A(x[40]), .B(y[71]), .Z(n2712) );
  NAND U2866 ( .A(x[27]), .B(y[20]), .Z(n2711) );
  XNOR U2867 ( .A(n2712), .B(n2711), .Z(n2713) );
  XNOR U2868 ( .A(n2714), .B(n2713), .Z(n2715) );
  XNOR U2869 ( .A(n2716), .B(n2715), .Z(n2732) );
  NAND U2870 ( .A(n2718), .B(n2717), .Z(n2722) );
  NAND U2871 ( .A(n2720), .B(n2719), .Z(n2721) );
  AND U2872 ( .A(n2722), .B(n2721), .Z(n2730) );
  AND U2873 ( .A(x[26]), .B(y[21]), .Z(n2724) );
  NAND U2874 ( .A(x[35]), .B(y[44]), .Z(n2723) );
  XNOR U2875 ( .A(n2724), .B(n2723), .Z(n2728) );
  AND U2876 ( .A(x[41]), .B(y[70]), .Z(n2726) );
  NAND U2877 ( .A(x[42]), .B(y[69]), .Z(n2725) );
  XNOR U2878 ( .A(n2726), .B(n2725), .Z(n2727) );
  XNOR U2879 ( .A(n2728), .B(n2727), .Z(n2729) );
  XNOR U2880 ( .A(n2730), .B(n2729), .Z(n2731) );
  XNOR U2881 ( .A(n2732), .B(n2731), .Z(n2733) );
  XNOR U2882 ( .A(n2734), .B(n2733), .Z(n2754) );
  NAND U2883 ( .A(n2736), .B(n2735), .Z(n2740) );
  NAND U2884 ( .A(n2738), .B(n2737), .Z(n2739) );
  AND U2885 ( .A(n2740), .B(n2739), .Z(n2752) );
  AND U2886 ( .A(x[38]), .B(y[41]), .Z(n2742) );
  NAND U2887 ( .A(x[37]), .B(y[42]), .Z(n2741) );
  XNOR U2888 ( .A(n2742), .B(n2741), .Z(n2750) );
  XNOR U2889 ( .A(n2750), .B(n2749), .Z(n2751) );
  XNOR U2890 ( .A(n2752), .B(n2751), .Z(n2753) );
  XNOR U2891 ( .A(n2754), .B(n2753), .Z(n2755) );
  XNOR U2892 ( .A(n2756), .B(n2755), .Z(n2757) );
  XNOR U2893 ( .A(n2758), .B(n2757), .Z(n2759) );
  XNOR U2894 ( .A(n2760), .B(n2759), .Z(n2776) );
  NAND U2895 ( .A(n2762), .B(n2761), .Z(n2766) );
  NAND U2896 ( .A(n2764), .B(n2763), .Z(n2765) );
  AND U2897 ( .A(n2766), .B(n2765), .Z(n2774) );
  NAND U2898 ( .A(n2768), .B(n2767), .Z(n2772) );
  NAND U2899 ( .A(n2770), .B(n2769), .Z(n2771) );
  NAND U2900 ( .A(n2772), .B(n2771), .Z(n2773) );
  XNOR U2901 ( .A(n2774), .B(n2773), .Z(n2775) );
  XNOR U2902 ( .A(n2776), .B(n2775), .Z(n2777) );
  XNOR U2903 ( .A(n2778), .B(n2777), .Z(n2794) );
  NAND U2904 ( .A(n2780), .B(n2779), .Z(n2784) );
  NAND U2905 ( .A(n2782), .B(n2781), .Z(n2783) );
  AND U2906 ( .A(n2784), .B(n2783), .Z(n2792) );
  NAND U2907 ( .A(n2786), .B(n2785), .Z(n2790) );
  NAND U2908 ( .A(n2788), .B(n2787), .Z(n2789) );
  NAND U2909 ( .A(n2790), .B(n2789), .Z(n2791) );
  XNOR U2910 ( .A(n2792), .B(n2791), .Z(n2793) );
  XNOR U2911 ( .A(n2794), .B(n2793), .Z(n2795) );
  XNOR U2912 ( .A(n2796), .B(n2795), .Z(o[47]) );
  AND U2913 ( .A(y[24]), .B(x[56]), .Z(n2798) );
  NAND U2914 ( .A(y[0]), .B(x[48]), .Z(n2797) );
  XNOR U2915 ( .A(n2798), .B(n2797), .Z(n2799) );
  NAND U2916 ( .A(y[48]), .B(x[64]), .Z(n2885) );
  XNOR U2917 ( .A(n2799), .B(n2885), .Z(o[48]) );
  AND U2918 ( .A(y[24]), .B(x[57]), .Z(n2872) );
  AND U2919 ( .A(y[25]), .B(x[56]), .Z(n2809) );
  AND U2920 ( .A(y[48]), .B(x[65]), .Z(n2808) );
  XOR U2921 ( .A(n2809), .B(n2808), .Z(n2810) );
  XNOR U2922 ( .A(n2872), .B(n2810), .Z(n2805) );
  NANDN U2923 ( .A(n2798), .B(n2797), .Z(n2801) );
  NAND U2924 ( .A(n2799), .B(n2885), .Z(n2800) );
  AND U2925 ( .A(n2801), .B(n2800), .Z(n2803) );
  AND U2926 ( .A(y[1]), .B(x[48]), .Z(n2836) );
  AND U2927 ( .A(y[49]), .B(x[64]), .Z(n2844) );
  AND U2928 ( .A(y[0]), .B(x[49]), .Z(n2813) );
  XOR U2929 ( .A(n2844), .B(n2813), .Z(n2814) );
  XNOR U2930 ( .A(n2836), .B(n2814), .Z(n2804) );
  XNOR U2931 ( .A(n2803), .B(n2804), .Z(n2802) );
  XNOR U2932 ( .A(n2805), .B(n2802), .Z(o[49]) );
  AND U2933 ( .A(x[49]), .B(y[1]), .Z(n2807) );
  NAND U2934 ( .A(x[48]), .B(y[2]), .Z(n2806) );
  XNOR U2935 ( .A(n2807), .B(n2806), .Z(n2838) );
  AND U2936 ( .A(y[24]), .B(x[58]), .Z(n2837) );
  XOR U2937 ( .A(n2838), .B(n2837), .Z(n2851) );
  AND U2938 ( .A(y[26]), .B(x[56]), .Z(n2849) );
  NAND U2939 ( .A(y[25]), .B(x[57]), .Z(n2848) );
  XNOR U2940 ( .A(n2849), .B(n2848), .Z(n2850) );
  XNOR U2941 ( .A(n2851), .B(n2850), .Z(n2824) );
  XNOR U2942 ( .A(n2825), .B(n2824), .Z(n2827) );
  NAND U2943 ( .A(n2809), .B(n2808), .Z(n2812) );
  NAND U2944 ( .A(n2872), .B(n2810), .Z(n2811) );
  NAND U2945 ( .A(n2812), .B(n2811), .Z(n2820) );
  NAND U2946 ( .A(n2844), .B(n2813), .Z(n2816) );
  NAND U2947 ( .A(n2836), .B(n2814), .Z(n2815) );
  NAND U2948 ( .A(n2816), .B(n2815), .Z(n2818) );
  AND U2949 ( .A(y[0]), .B(x[50]), .Z(n2864) );
  NAND U2950 ( .A(y[48]), .B(x[66]), .Z(n2830) );
  XNOR U2951 ( .A(n2864), .B(n2830), .Z(n2832) );
  AND U2952 ( .A(x[65]), .B(y[49]), .Z(n2878) );
  NAND U2953 ( .A(x[64]), .B(y[50]), .Z(n2817) );
  XNOR U2954 ( .A(n2878), .B(n2817), .Z(n2831) );
  XOR U2955 ( .A(n2832), .B(n2831), .Z(n2819) );
  XNOR U2956 ( .A(n2818), .B(n2819), .Z(n2821) );
  XOR U2957 ( .A(n2820), .B(n2821), .Z(n2826) );
  XNOR U2958 ( .A(n2827), .B(n2826), .Z(o[50]) );
  NAND U2959 ( .A(n2819), .B(n2818), .Z(n2823) );
  NANDN U2960 ( .A(n2821), .B(n2820), .Z(n2822) );
  AND U2961 ( .A(n2823), .B(n2822), .Z(n2859) );
  NANDN U2962 ( .A(n2825), .B(n2824), .Z(n2829) );
  NAND U2963 ( .A(n2827), .B(n2826), .Z(n2828) );
  AND U2964 ( .A(n2829), .B(n2828), .Z(n2858) );
  XNOR U2965 ( .A(n2859), .B(n2858), .Z(n2861) );
  NANDN U2966 ( .A(n2830), .B(n2864), .Z(n2834) );
  NAND U2967 ( .A(n2832), .B(n2831), .Z(n2833) );
  NAND U2968 ( .A(n2834), .B(n2833), .Z(n2892) );
  AND U2969 ( .A(y[27]), .B(x[56]), .Z(n2879) );
  AND U2970 ( .A(y[2]), .B(x[49]), .Z(n2880) );
  NAND U2971 ( .A(y[3]), .B(x[48]), .Z(n2882) );
  XNOR U2972 ( .A(n2881), .B(n2882), .Z(n2891) );
  AND U2973 ( .A(x[57]), .B(y[26]), .Z(n2922) );
  NAND U2974 ( .A(x[59]), .B(y[24]), .Z(n2835) );
  XNOR U2975 ( .A(n2922), .B(n2835), .Z(n2874) );
  AND U2976 ( .A(y[25]), .B(x[58]), .Z(n2873) );
  XOR U2977 ( .A(n2874), .B(n2873), .Z(n2890) );
  XOR U2978 ( .A(n2891), .B(n2890), .Z(n2893) );
  XOR U2979 ( .A(n2892), .B(n2893), .Z(n2855) );
  NAND U2980 ( .A(n2880), .B(n2836), .Z(n2840) );
  NAND U2981 ( .A(n2838), .B(n2837), .Z(n2839) );
  NAND U2982 ( .A(n2840), .B(n2839), .Z(n2898) );
  AND U2983 ( .A(x[50]), .B(y[1]), .Z(n2842) );
  NAND U2984 ( .A(x[51]), .B(y[0]), .Z(n2841) );
  XNOR U2985 ( .A(n2842), .B(n2841), .Z(n2865) );
  AND U2986 ( .A(y[50]), .B(x[65]), .Z(n2843) );
  NAND U2987 ( .A(n2844), .B(n2843), .Z(n2866) );
  XNOR U2988 ( .A(n2865), .B(n2866), .Z(n2897) );
  AND U2989 ( .A(x[67]), .B(y[48]), .Z(n2846) );
  NAND U2990 ( .A(x[64]), .B(y[51]), .Z(n2845) );
  XNOR U2991 ( .A(n2846), .B(n2845), .Z(n2887) );
  AND U2992 ( .A(x[66]), .B(y[49]), .Z(n2932) );
  NAND U2993 ( .A(x[65]), .B(y[50]), .Z(n2847) );
  XNOR U2994 ( .A(n2932), .B(n2847), .Z(n2886) );
  XOR U2995 ( .A(n2887), .B(n2886), .Z(n2896) );
  XOR U2996 ( .A(n2897), .B(n2896), .Z(n2899) );
  XNOR U2997 ( .A(n2898), .B(n2899), .Z(n2854) );
  XNOR U2998 ( .A(n2855), .B(n2854), .Z(n2856) );
  NANDN U2999 ( .A(n2849), .B(n2848), .Z(n2853) );
  NANDN U3000 ( .A(n2851), .B(n2850), .Z(n2852) );
  NAND U3001 ( .A(n2853), .B(n2852), .Z(n2857) );
  XNOR U3002 ( .A(n2856), .B(n2857), .Z(n2860) );
  XOR U3003 ( .A(n2861), .B(n2860), .Z(o[51]) );
  NANDN U3004 ( .A(n2859), .B(n2858), .Z(n2863) );
  NAND U3005 ( .A(n2861), .B(n2860), .Z(n2862) );
  NAND U3006 ( .A(n2863), .B(n2862), .Z(n2965) );
  XNOR U3007 ( .A(n2966), .B(n2965), .Z(n2968) );
  NAND U3008 ( .A(y[1]), .B(x[51]), .Z(n2919) );
  NANDN U3009 ( .A(n2919), .B(n2864), .Z(n2868) );
  NANDN U3010 ( .A(n2866), .B(n2865), .Z(n2867) );
  NAND U3011 ( .A(n2868), .B(n2867), .Z(n2946) );
  AND U3012 ( .A(x[67]), .B(y[49]), .Z(n3033) );
  NAND U3013 ( .A(x[66]), .B(y[50]), .Z(n2869) );
  XNOR U3014 ( .A(n3033), .B(n2869), .Z(n2902) );
  AND U3015 ( .A(y[51]), .B(x[65]), .Z(n2903) );
  AND U3016 ( .A(y[48]), .B(x[68]), .Z(n2905) );
  AND U3017 ( .A(x[57]), .B(y[27]), .Z(n2871) );
  NAND U3018 ( .A(x[58]), .B(y[26]), .Z(n2870) );
  XNOR U3019 ( .A(n2871), .B(n2870), .Z(n2923) );
  NAND U3020 ( .A(y[25]), .B(x[59]), .Z(n2924) );
  XNOR U3021 ( .A(n2923), .B(n2924), .Z(n2944) );
  NAND U3022 ( .A(y[26]), .B(x[59]), .Z(n2936) );
  IV U3023 ( .A(n2936), .Z(n3020) );
  NAND U3024 ( .A(n3020), .B(n2872), .Z(n2876) );
  NAND U3025 ( .A(n2874), .B(n2873), .Z(n2875) );
  NAND U3026 ( .A(n2876), .B(n2875), .Z(n2940) );
  AND U3027 ( .A(y[52]), .B(x[64]), .Z(n2997) );
  AND U3028 ( .A(y[0]), .B(x[52]), .Z(n2908) );
  AND U3029 ( .A(y[50]), .B(x[66]), .Z(n2877) );
  NAND U3030 ( .A(n2878), .B(n2877), .Z(n2909) );
  XOR U3031 ( .A(n2908), .B(n2909), .Z(n2910) );
  XNOR U3032 ( .A(n2997), .B(n2910), .Z(n2937) );
  AND U3033 ( .A(y[24]), .B(x[60]), .Z(n3037) );
  AND U3034 ( .A(y[28]), .B(x[56]), .Z(n2927) );
  XOR U3035 ( .A(n3037), .B(n2927), .Z(n2928) );
  NAND U3036 ( .A(y[3]), .B(x[49]), .Z(n2929) );
  XNOR U3037 ( .A(n2928), .B(n2929), .Z(n2938) );
  XNOR U3038 ( .A(n2950), .B(n2949), .Z(n2952) );
  NAND U3039 ( .A(n2880), .B(n2879), .Z(n2884) );
  NANDN U3040 ( .A(n2882), .B(n2881), .Z(n2883) );
  NAND U3041 ( .A(n2884), .B(n2883), .Z(n2955) );
  NAND U3042 ( .A(y[2]), .B(x[50]), .Z(n2917) );
  NAND U3043 ( .A(y[4]), .B(x[48]), .Z(n2918) );
  XOR U3044 ( .A(n2919), .B(n2918), .Z(n2916) );
  AND U3045 ( .A(y[51]), .B(x[67]), .Z(n3132) );
  NANDN U3046 ( .A(n2885), .B(n3132), .Z(n2889) );
  NAND U3047 ( .A(n2887), .B(n2886), .Z(n2888) );
  NAND U3048 ( .A(n2889), .B(n2888), .Z(n2953) );
  XNOR U3049 ( .A(n2954), .B(n2953), .Z(n2956) );
  XNOR U3050 ( .A(n2955), .B(n2956), .Z(n2951) );
  XNOR U3051 ( .A(n2952), .B(n2951), .Z(n2962) );
  NAND U3052 ( .A(n2891), .B(n2890), .Z(n2895) );
  NAND U3053 ( .A(n2893), .B(n2892), .Z(n2894) );
  AND U3054 ( .A(n2895), .B(n2894), .Z(n2960) );
  NAND U3055 ( .A(n2897), .B(n2896), .Z(n2901) );
  NAND U3056 ( .A(n2899), .B(n2898), .Z(n2900) );
  AND U3057 ( .A(n2901), .B(n2900), .Z(n2959) );
  XOR U3058 ( .A(n2960), .B(n2959), .Z(n2961) );
  XOR U3059 ( .A(n2962), .B(n2961), .Z(n2967) );
  XOR U3060 ( .A(n2968), .B(n2967), .Z(o[52]) );
  NAND U3061 ( .A(n2903), .B(n2902), .Z(n2907) );
  NAND U3062 ( .A(n2905), .B(n2904), .Z(n2906) );
  NAND U3063 ( .A(n2907), .B(n2906), .Z(n3012) );
  NANDN U3064 ( .A(n2909), .B(n2908), .Z(n2912) );
  NANDN U3065 ( .A(n2910), .B(n2997), .Z(n2911) );
  AND U3066 ( .A(n2912), .B(n2911), .Z(n3018) );
  AND U3067 ( .A(x[61]), .B(y[24]), .Z(n2914) );
  NAND U3068 ( .A(x[60]), .B(y[25]), .Z(n2913) );
  XNOR U3069 ( .A(n2914), .B(n2913), .Z(n3039) );
  NAND U3070 ( .A(y[4]), .B(x[49]), .Z(n3038) );
  XNOR U3071 ( .A(n3039), .B(n3038), .Z(n3017) );
  AND U3072 ( .A(y[51]), .B(x[66]), .Z(n3026) );
  NAND U3073 ( .A(y[48]), .B(x[69]), .Z(n3025) );
  XNOR U3074 ( .A(n3026), .B(n3025), .Z(n3029) );
  AND U3075 ( .A(y[49]), .B(x[68]), .Z(n3107) );
  NAND U3076 ( .A(x[67]), .B(y[50]), .Z(n2915) );
  XNOR U3077 ( .A(n3107), .B(n2915), .Z(n3028) );
  XNOR U3078 ( .A(n3029), .B(n3028), .Z(n3016) );
  XNOR U3079 ( .A(n3017), .B(n3016), .Z(n3019) );
  XNOR U3080 ( .A(n3018), .B(n3019), .Z(n3011) );
  NAND U3081 ( .A(n2917), .B(n2916), .Z(n2921) );
  AND U3082 ( .A(n2919), .B(n2918), .Z(n2920) );
  ANDN U3083 ( .B(n2921), .A(n2920), .Z(n3010) );
  XOR U3084 ( .A(n3011), .B(n3010), .Z(n3013) );
  XNOR U3085 ( .A(n3012), .B(n3013), .Z(n2977) );
  AND U3086 ( .A(y[27]), .B(x[58]), .Z(n3000) );
  NAND U3087 ( .A(n3000), .B(n2922), .Z(n2926) );
  NANDN U3088 ( .A(n2924), .B(n2923), .Z(n2925) );
  NAND U3089 ( .A(n2926), .B(n2925), .Z(n2990) );
  AND U3090 ( .A(y[0]), .B(x[53]), .Z(n3080) );
  NAND U3091 ( .A(y[1]), .B(x[52]), .Z(n3001) );
  XNOR U3092 ( .A(n3002), .B(n3001), .Z(n2988) );
  AND U3093 ( .A(y[28]), .B(x[57]), .Z(n3098) );
  AND U3094 ( .A(y[5]), .B(x[48]), .Z(n3006) );
  AND U3095 ( .A(y[29]), .B(x[56]), .Z(n3005) );
  XNOR U3096 ( .A(n3006), .B(n3005), .Z(n3007) );
  XNOR U3097 ( .A(n3098), .B(n3007), .Z(n2987) );
  XNOR U3098 ( .A(n2988), .B(n2987), .Z(n2989) );
  XOR U3099 ( .A(n2990), .B(n2989), .Z(n2976) );
  AND U3100 ( .A(n3037), .B(n2927), .Z(n2931) );
  NANDN U3101 ( .A(n2929), .B(n2928), .Z(n2930) );
  NANDN U3102 ( .A(n2931), .B(n2930), .Z(n2993) );
  AND U3103 ( .A(y[50]), .B(x[67]), .Z(n2933) );
  AND U3104 ( .A(n2933), .B(n2932), .Z(n2999) );
  AND U3105 ( .A(x[64]), .B(y[53]), .Z(n2935) );
  AND U3106 ( .A(x[65]), .B(y[52]), .Z(n2934) );
  XNOR U3107 ( .A(n2935), .B(n2934), .Z(n2998) );
  XNOR U3108 ( .A(n2999), .B(n2998), .Z(n2992) );
  AND U3109 ( .A(y[2]), .B(x[51]), .Z(n3085) );
  XNOR U3110 ( .A(n3085), .B(n2936), .Z(n3022) );
  NAND U3111 ( .A(y[3]), .B(x[50]), .Z(n3021) );
  XNOR U3112 ( .A(n3022), .B(n3021), .Z(n2991) );
  XNOR U3113 ( .A(n2992), .B(n2991), .Z(n2994) );
  XOR U3114 ( .A(n2993), .B(n2994), .Z(n2975) );
  XOR U3115 ( .A(n2976), .B(n2975), .Z(n2978) );
  XNOR U3116 ( .A(n2977), .B(n2978), .Z(n2983) );
  NAND U3117 ( .A(n2938), .B(n2937), .Z(n2942) );
  NAND U3118 ( .A(n2940), .B(n2939), .Z(n2941) );
  NAND U3119 ( .A(n2942), .B(n2941), .Z(n2982) );
  NAND U3120 ( .A(n2944), .B(n2943), .Z(n2948) );
  NAND U3121 ( .A(n2946), .B(n2945), .Z(n2947) );
  NAND U3122 ( .A(n2948), .B(n2947), .Z(n2981) );
  XOR U3123 ( .A(n2983), .B(n2984), .Z(n2973) );
  NANDN U3124 ( .A(n2954), .B(n2953), .Z(n2958) );
  NAND U3125 ( .A(n2956), .B(n2955), .Z(n2957) );
  NAND U3126 ( .A(n2958), .B(n2957), .Z(n2972) );
  XNOR U3127 ( .A(n2971), .B(n2972), .Z(n2974) );
  XNOR U3128 ( .A(n2973), .B(n2974), .Z(n3043) );
  NAND U3129 ( .A(n2960), .B(n2959), .Z(n2964) );
  NANDN U3130 ( .A(n2962), .B(n2961), .Z(n2963) );
  AND U3131 ( .A(n2964), .B(n2963), .Z(n3041) );
  NANDN U3132 ( .A(n2966), .B(n2965), .Z(n2970) );
  NAND U3133 ( .A(n2968), .B(n2967), .Z(n2969) );
  AND U3134 ( .A(n2970), .B(n2969), .Z(n3040) );
  XNOR U3135 ( .A(n3041), .B(n3040), .Z(n3042) );
  XNOR U3136 ( .A(n3043), .B(n3042), .Z(o[53]) );
  NAND U3137 ( .A(n2976), .B(n2975), .Z(n2980) );
  NAND U3138 ( .A(n2978), .B(n2977), .Z(n2979) );
  NAND U3139 ( .A(n2980), .B(n2979), .Z(n3212) );
  NAND U3140 ( .A(n2982), .B(n2981), .Z(n2986) );
  NAND U3141 ( .A(n2984), .B(n2983), .Z(n2985) );
  AND U3142 ( .A(n2986), .B(n2985), .Z(n3213) );
  XOR U3143 ( .A(n3212), .B(n3213), .Z(n3211) );
  NAND U3144 ( .A(n2992), .B(n2991), .Z(n2996) );
  NANDN U3145 ( .A(n2994), .B(n2993), .Z(n2995) );
  AND U3146 ( .A(n2996), .B(n2995), .Z(n3188) );
  XOR U3147 ( .A(n3189), .B(n3188), .Z(n3187) );
  AND U3148 ( .A(y[53]), .B(x[65]), .Z(n3161) );
  AND U3149 ( .A(y[25]), .B(x[61]), .Z(n3109) );
  AND U3150 ( .A(y[24]), .B(x[62]), .Z(n3111) );
  AND U3151 ( .A(y[6]), .B(x[48]), .Z(n3110) );
  XOR U3152 ( .A(n3111), .B(n3110), .Z(n3108) );
  XNOR U3153 ( .A(n3109), .B(n3108), .Z(n3075) );
  AND U3154 ( .A(x[69]), .B(y[49]), .Z(n3004) );
  NAND U3155 ( .A(x[68]), .B(y[50]), .Z(n3003) );
  XNOR U3156 ( .A(n3004), .B(n3003), .Z(n3135) );
  AND U3157 ( .A(y[48]), .B(x[70]), .Z(n3134) );
  XOR U3158 ( .A(n3135), .B(n3134), .Z(n3133) );
  XNOR U3159 ( .A(n3133), .B(n3132), .Z(n3074) );
  XOR U3160 ( .A(n3073), .B(n3072), .Z(n3048) );
  XOR U3161 ( .A(n3049), .B(n3048), .Z(n3047) );
  AND U3162 ( .A(x[53]), .B(y[1]), .Z(n3009) );
  NAND U3163 ( .A(x[54]), .B(y[0]), .Z(n3008) );
  XNOR U3164 ( .A(n3009), .B(n3008), .Z(n3079) );
  AND U3165 ( .A(y[27]), .B(x[59]), .Z(n3078) );
  XNOR U3166 ( .A(n3079), .B(n3078), .Z(n3061) );
  AND U3167 ( .A(y[54]), .B(x[64]), .Z(n3093) );
  AND U3168 ( .A(y[30]), .B(x[56]), .Z(n3092) );
  XOR U3169 ( .A(n3093), .B(n3092), .Z(n3091) );
  AND U3170 ( .A(y[5]), .B(x[49]), .Z(n3090) );
  XNOR U3171 ( .A(n3091), .B(n3090), .Z(n3060) );
  XNOR U3172 ( .A(n3058), .B(n3059), .Z(n3046) );
  XNOR U3173 ( .A(n3047), .B(n3046), .Z(n3186) );
  XNOR U3174 ( .A(n3187), .B(n3186), .Z(n3217) );
  NAND U3175 ( .A(n3011), .B(n3010), .Z(n3015) );
  NAND U3176 ( .A(n3013), .B(n3012), .Z(n3014) );
  AND U3177 ( .A(n3015), .B(n3014), .Z(n3219) );
  AND U3178 ( .A(x[57]), .B(y[29]), .Z(n3024) );
  NAND U3179 ( .A(x[58]), .B(y[28]), .Z(n3023) );
  XNOR U3180 ( .A(n3024), .B(n3023), .Z(n3097) );
  AND U3181 ( .A(y[4]), .B(x[50]), .Z(n3096) );
  XNOR U3182 ( .A(n3097), .B(n3096), .Z(n3067) );
  IV U3183 ( .A(n3067), .Z(n3032) );
  IV U3184 ( .A(n3025), .Z(n3027) );
  NAND U3185 ( .A(n3027), .B(n3026), .Z(n3031) );
  NAND U3186 ( .A(n3029), .B(n3028), .Z(n3030) );
  AND U3187 ( .A(n3031), .B(n3030), .Z(n3066) );
  XNOR U3188 ( .A(n3032), .B(n3066), .Z(n3064) );
  XOR U3189 ( .A(n3065), .B(n3064), .Z(n3192) );
  XOR U3190 ( .A(n3193), .B(n3192), .Z(n3191) );
  AND U3191 ( .A(y[50]), .B(x[68]), .Z(n3034) );
  AND U3192 ( .A(n3034), .B(n3033), .Z(n3163) );
  AND U3193 ( .A(y[52]), .B(x[66]), .Z(n3162) );
  XOR U3194 ( .A(n3163), .B(n3162), .Z(n3160) );
  AND U3195 ( .A(x[51]), .B(y[3]), .Z(n3036) );
  NAND U3196 ( .A(x[52]), .B(y[2]), .Z(n3035) );
  XNOR U3197 ( .A(n3036), .B(n3035), .Z(n3084) );
  AND U3198 ( .A(y[26]), .B(x[60]), .Z(n3083) );
  XNOR U3199 ( .A(n3084), .B(n3083), .Z(n3055) );
  XNOR U3200 ( .A(n3053), .B(n3052), .Z(n3190) );
  XOR U3201 ( .A(n3191), .B(n3190), .Z(n3218) );
  XOR U3202 ( .A(n3219), .B(n3218), .Z(n3216) );
  XOR U3203 ( .A(n3217), .B(n3216), .Z(n3210) );
  XOR U3204 ( .A(n3211), .B(n3210), .Z(n3204) );
  NANDN U3205 ( .A(n3041), .B(n3040), .Z(n3045) );
  NAND U3206 ( .A(n3043), .B(n3042), .Z(n3044) );
  NAND U3207 ( .A(n3045), .B(n3044), .Z(n3202) );
  XNOR U3208 ( .A(n3203), .B(n3202), .Z(o[54]) );
  NAND U3209 ( .A(n3047), .B(n3046), .Z(n3051) );
  NAND U3210 ( .A(n3049), .B(n3048), .Z(n3050) );
  AND U3211 ( .A(n3051), .B(n3050), .Z(n3201) );
  NANDN U3212 ( .A(n3053), .B(n3052), .Z(n3057) );
  NAND U3213 ( .A(n3055), .B(n3054), .Z(n3056) );
  AND U3214 ( .A(n3057), .B(n3056), .Z(n3185) );
  NANDN U3215 ( .A(n3059), .B(n3058), .Z(n3063) );
  NAND U3216 ( .A(n3061), .B(n3060), .Z(n3062) );
  AND U3217 ( .A(n3063), .B(n3062), .Z(n3071) );
  NAND U3218 ( .A(n3065), .B(n3064), .Z(n3069) );
  NAND U3219 ( .A(n3067), .B(n3066), .Z(n3068) );
  NAND U3220 ( .A(n3069), .B(n3068), .Z(n3070) );
  XNOR U3221 ( .A(n3071), .B(n3070), .Z(n3183) );
  NAND U3222 ( .A(n3073), .B(n3072), .Z(n3077) );
  NAND U3223 ( .A(n3075), .B(n3074), .Z(n3076) );
  AND U3224 ( .A(n3077), .B(n3076), .Z(n3181) );
  NAND U3225 ( .A(n3079), .B(n3078), .Z(n3082) );
  AND U3226 ( .A(y[1]), .B(x[54]), .Z(n3143) );
  NAND U3227 ( .A(n3080), .B(n3143), .Z(n3081) );
  AND U3228 ( .A(n3082), .B(n3081), .Z(n3089) );
  NAND U3229 ( .A(n3084), .B(n3083), .Z(n3087) );
  AND U3230 ( .A(y[3]), .B(x[52]), .Z(n3124) );
  NAND U3231 ( .A(n3085), .B(n3124), .Z(n3086) );
  NAND U3232 ( .A(n3087), .B(n3086), .Z(n3088) );
  XNOR U3233 ( .A(n3089), .B(n3088), .Z(n3104) );
  NAND U3234 ( .A(n3091), .B(n3090), .Z(n3095) );
  NAND U3235 ( .A(n3093), .B(n3092), .Z(n3094) );
  AND U3236 ( .A(n3095), .B(n3094), .Z(n3102) );
  NAND U3237 ( .A(n3097), .B(n3096), .Z(n3100) );
  AND U3238 ( .A(y[29]), .B(x[58]), .Z(n3125) );
  NAND U3239 ( .A(n3125), .B(n3098), .Z(n3099) );
  NAND U3240 ( .A(n3100), .B(n3099), .Z(n3101) );
  XNOR U3241 ( .A(n3102), .B(n3101), .Z(n3103) );
  XOR U3242 ( .A(n3104), .B(n3103), .Z(n3131) );
  AND U3243 ( .A(x[71]), .B(y[48]), .Z(n3106) );
  NAND U3244 ( .A(x[68]), .B(y[51]), .Z(n3105) );
  XNOR U3245 ( .A(n3106), .B(n3105), .Z(n3129) );
  AND U3246 ( .A(y[50]), .B(x[69]), .Z(n3147) );
  AND U3247 ( .A(n3107), .B(n3147), .Z(n3123) );
  NAND U3248 ( .A(n3109), .B(n3108), .Z(n3113) );
  NAND U3249 ( .A(n3111), .B(n3110), .Z(n3112) );
  AND U3250 ( .A(n3113), .B(n3112), .Z(n3121) );
  AND U3251 ( .A(x[64]), .B(y[55]), .Z(n3115) );
  NAND U3252 ( .A(x[70]), .B(y[49]), .Z(n3114) );
  XNOR U3253 ( .A(n3115), .B(n3114), .Z(n3119) );
  AND U3254 ( .A(x[49]), .B(y[6]), .Z(n3117) );
  NAND U3255 ( .A(x[51]), .B(y[4]), .Z(n3116) );
  XNOR U3256 ( .A(n3117), .B(n3116), .Z(n3118) );
  XNOR U3257 ( .A(n3119), .B(n3118), .Z(n3120) );
  XNOR U3258 ( .A(n3121), .B(n3120), .Z(n3122) );
  XOR U3259 ( .A(n3123), .B(n3122), .Z(n3127) );
  XNOR U3260 ( .A(n3125), .B(n3124), .Z(n3126) );
  XNOR U3261 ( .A(n3127), .B(n3126), .Z(n3128) );
  XNOR U3262 ( .A(n3129), .B(n3128), .Z(n3130) );
  XNOR U3263 ( .A(n3131), .B(n3130), .Z(n3179) );
  NAND U3264 ( .A(n3133), .B(n3132), .Z(n3137) );
  AND U3265 ( .A(n3135), .B(n3134), .Z(n3136) );
  ANDN U3266 ( .B(n3137), .A(n3136), .Z(n3177) );
  AND U3267 ( .A(x[48]), .B(y[7]), .Z(n3139) );
  NAND U3268 ( .A(x[53]), .B(y[2]), .Z(n3138) );
  XNOR U3269 ( .A(n3139), .B(n3138), .Z(n3151) );
  AND U3270 ( .A(x[59]), .B(y[28]), .Z(n3149) );
  AND U3271 ( .A(x[60]), .B(y[27]), .Z(n3145) );
  AND U3272 ( .A(x[67]), .B(y[52]), .Z(n3141) );
  NAND U3273 ( .A(x[55]), .B(y[0]), .Z(n3140) );
  XNOR U3274 ( .A(n3141), .B(n3140), .Z(n3142) );
  XNOR U3275 ( .A(n3143), .B(n3142), .Z(n3144) );
  XNOR U3276 ( .A(n3145), .B(n3144), .Z(n3146) );
  XNOR U3277 ( .A(n3147), .B(n3146), .Z(n3148) );
  XNOR U3278 ( .A(n3149), .B(n3148), .Z(n3150) );
  XOR U3279 ( .A(n3151), .B(n3150), .Z(n3159) );
  AND U3280 ( .A(x[56]), .B(y[31]), .Z(n3153) );
  NAND U3281 ( .A(x[57]), .B(y[30]), .Z(n3152) );
  XNOR U3282 ( .A(n3153), .B(n3152), .Z(n3157) );
  AND U3283 ( .A(x[66]), .B(y[53]), .Z(n3155) );
  NAND U3284 ( .A(x[63]), .B(y[24]), .Z(n3154) );
  XNOR U3285 ( .A(n3155), .B(n3154), .Z(n3156) );
  XNOR U3286 ( .A(n3157), .B(n3156), .Z(n3158) );
  XNOR U3287 ( .A(n3159), .B(n3158), .Z(n3175) );
  NAND U3288 ( .A(n3161), .B(n3160), .Z(n3165) );
  NAND U3289 ( .A(n3163), .B(n3162), .Z(n3164) );
  AND U3290 ( .A(n3165), .B(n3164), .Z(n3173) );
  AND U3291 ( .A(x[61]), .B(y[26]), .Z(n3167) );
  NAND U3292 ( .A(x[62]), .B(y[25]), .Z(n3166) );
  XNOR U3293 ( .A(n3167), .B(n3166), .Z(n3171) );
  AND U3294 ( .A(x[65]), .B(y[54]), .Z(n3169) );
  NAND U3295 ( .A(x[50]), .B(y[5]), .Z(n3168) );
  XNOR U3296 ( .A(n3169), .B(n3168), .Z(n3170) );
  XNOR U3297 ( .A(n3171), .B(n3170), .Z(n3172) );
  XNOR U3298 ( .A(n3173), .B(n3172), .Z(n3174) );
  XNOR U3299 ( .A(n3175), .B(n3174), .Z(n3176) );
  XNOR U3300 ( .A(n3177), .B(n3176), .Z(n3178) );
  XNOR U3301 ( .A(n3179), .B(n3178), .Z(n3180) );
  XNOR U3302 ( .A(n3181), .B(n3180), .Z(n3182) );
  XNOR U3303 ( .A(n3183), .B(n3182), .Z(n3184) );
  XNOR U3304 ( .A(n3185), .B(n3184), .Z(n3199) );
  NAND U3305 ( .A(n3191), .B(n3190), .Z(n3195) );
  NAND U3306 ( .A(n3193), .B(n3192), .Z(n3194) );
  NAND U3307 ( .A(n3195), .B(n3194), .Z(n3196) );
  XNOR U3308 ( .A(n3197), .B(n3196), .Z(n3198) );
  XNOR U3309 ( .A(n3199), .B(n3198), .Z(n3200) );
  XNOR U3310 ( .A(n3201), .B(n3200), .Z(n3209) );
  NAND U3311 ( .A(n3203), .B(n3202), .Z(n3207) );
  NAND U3312 ( .A(n3205), .B(n3204), .Z(n3206) );
  NAND U3313 ( .A(n3207), .B(n3206), .Z(n3208) );
  XNOR U3314 ( .A(n3209), .B(n3208), .Z(n3225) );
  NAND U3315 ( .A(n3211), .B(n3210), .Z(n3215) );
  NAND U3316 ( .A(n3213), .B(n3212), .Z(n3214) );
  AND U3317 ( .A(n3215), .B(n3214), .Z(n3223) );
  NAND U3318 ( .A(n3217), .B(n3216), .Z(n3221) );
  NAND U3319 ( .A(n3219), .B(n3218), .Z(n3220) );
  NAND U3320 ( .A(n3221), .B(n3220), .Z(n3222) );
  XNOR U3321 ( .A(n3223), .B(n3222), .Z(n3224) );
  XNOR U3322 ( .A(n3225), .B(n3224), .Z(o[55]) );
  AND U3323 ( .A(y[32]), .B(x[56]), .Z(n3227) );
  NAND U3324 ( .A(y[8]), .B(x[48]), .Z(n3226) );
  XNOR U3325 ( .A(n3227), .B(n3226), .Z(n3228) );
  NAND U3326 ( .A(y[56]), .B(x[64]), .Z(n3318) );
  XNOR U3327 ( .A(n3228), .B(n3318), .Z(o[56]) );
  AND U3328 ( .A(y[9]), .B(x[48]), .Z(n3267) );
  AND U3329 ( .A(y[57]), .B(x[64]), .Z(n3274) );
  AND U3330 ( .A(y[8]), .B(x[49]), .Z(n3244) );
  XOR U3331 ( .A(n3274), .B(n3244), .Z(n3245) );
  XOR U3332 ( .A(n3267), .B(n3245), .Z(n3231) );
  NANDN U3333 ( .A(n3227), .B(n3226), .Z(n3230) );
  NAND U3334 ( .A(n3228), .B(n3318), .Z(n3229) );
  NAND U3335 ( .A(n3230), .B(n3229), .Z(n3232) );
  XNOR U3336 ( .A(n3231), .B(n3232), .Z(n3234) );
  AND U3337 ( .A(y[32]), .B(x[57]), .Z(n3305) );
  AND U3338 ( .A(y[33]), .B(x[56]), .Z(n3240) );
  AND U3339 ( .A(y[56]), .B(x[65]), .Z(n3239) );
  XOR U3340 ( .A(n3240), .B(n3239), .Z(n3241) );
  XOR U3341 ( .A(n3305), .B(n3241), .Z(n3233) );
  XOR U3342 ( .A(n3234), .B(n3233), .Z(o[57]) );
  NANDN U3343 ( .A(n3232), .B(n3231), .Z(n3236) );
  NAND U3344 ( .A(n3234), .B(n3233), .Z(n3235) );
  AND U3345 ( .A(n3236), .B(n3235), .Z(n3257) );
  AND U3346 ( .A(x[48]), .B(y[10]), .Z(n3238) );
  NAND U3347 ( .A(x[49]), .B(y[9]), .Z(n3237) );
  XNOR U3348 ( .A(n3238), .B(n3237), .Z(n3268) );
  NAND U3349 ( .A(y[32]), .B(x[58]), .Z(n3269) );
  XOR U3350 ( .A(n3268), .B(n3269), .Z(n3281) );
  NAND U3351 ( .A(y[34]), .B(x[56]), .Z(n3280) );
  NAND U3352 ( .A(y[33]), .B(x[57]), .Z(n3279) );
  XOR U3353 ( .A(n3280), .B(n3279), .Z(n3282) );
  XNOR U3354 ( .A(n3281), .B(n3282), .Z(n3256) );
  XNOR U3355 ( .A(n3257), .B(n3256), .Z(n3259) );
  NAND U3356 ( .A(n3240), .B(n3239), .Z(n3243) );
  NAND U3357 ( .A(n3305), .B(n3241), .Z(n3242) );
  NAND U3358 ( .A(n3243), .B(n3242), .Z(n3252) );
  NAND U3359 ( .A(n3274), .B(n3244), .Z(n3247) );
  NAND U3360 ( .A(n3267), .B(n3245), .Z(n3246) );
  NAND U3361 ( .A(n3247), .B(n3246), .Z(n3250) );
  AND U3362 ( .A(y[8]), .B(x[50]), .Z(n3297) );
  NAND U3363 ( .A(y[56]), .B(x[66]), .Z(n3260) );
  XNOR U3364 ( .A(n3297), .B(n3260), .Z(n3262) );
  AND U3365 ( .A(x[64]), .B(y[58]), .Z(n3249) );
  NAND U3366 ( .A(x[65]), .B(y[57]), .Z(n3248) );
  XNOR U3367 ( .A(n3249), .B(n3248), .Z(n3261) );
  XOR U3368 ( .A(n3262), .B(n3261), .Z(n3251) );
  XNOR U3369 ( .A(n3250), .B(n3251), .Z(n3253) );
  XOR U3370 ( .A(n3252), .B(n3253), .Z(n3258) );
  XNOR U3371 ( .A(n3259), .B(n3258), .Z(o[58]) );
  NAND U3372 ( .A(n3251), .B(n3250), .Z(n3255) );
  NANDN U3373 ( .A(n3253), .B(n3252), .Z(n3254) );
  AND U3374 ( .A(n3255), .B(n3254), .Z(n3292) );
  XNOR U3375 ( .A(n3292), .B(n3291), .Z(n3294) );
  NANDN U3376 ( .A(n3260), .B(n3297), .Z(n3264) );
  NAND U3377 ( .A(n3262), .B(n3261), .Z(n3263) );
  AND U3378 ( .A(n3264), .B(n3263), .Z(n3326) );
  AND U3379 ( .A(y[35]), .B(x[56]), .Z(n3312) );
  AND U3380 ( .A(y[10]), .B(x[49]), .Z(n3313) );
  NAND U3381 ( .A(y[11]), .B(x[48]), .Z(n3315) );
  XNOR U3382 ( .A(n3314), .B(n3315), .Z(n3323) );
  AND U3383 ( .A(x[59]), .B(y[32]), .Z(n3266) );
  NAND U3384 ( .A(x[57]), .B(y[34]), .Z(n3265) );
  XNOR U3385 ( .A(n3266), .B(n3265), .Z(n3306) );
  NAND U3386 ( .A(y[33]), .B(x[58]), .Z(n3307) );
  XOR U3387 ( .A(n3306), .B(n3307), .Z(n3324) );
  XNOR U3388 ( .A(n3323), .B(n3324), .Z(n3325) );
  XNOR U3389 ( .A(n3326), .B(n3325), .Z(n3286) );
  NAND U3390 ( .A(n3313), .B(n3267), .Z(n3271) );
  NANDN U3391 ( .A(n3269), .B(n3268), .Z(n3270) );
  AND U3392 ( .A(n3271), .B(n3270), .Z(n3331) );
  AND U3393 ( .A(x[50]), .B(y[9]), .Z(n3273) );
  NAND U3394 ( .A(x[51]), .B(y[8]), .Z(n3272) );
  XNOR U3395 ( .A(n3273), .B(n3272), .Z(n3298) );
  AND U3396 ( .A(x[65]), .B(y[58]), .Z(n3278) );
  NAND U3397 ( .A(n3274), .B(n3278), .Z(n3299) );
  XNOR U3398 ( .A(n3298), .B(n3299), .Z(n3329) );
  AND U3399 ( .A(x[67]), .B(y[56]), .Z(n3276) );
  NAND U3400 ( .A(x[64]), .B(y[59]), .Z(n3275) );
  XNOR U3401 ( .A(n3276), .B(n3275), .Z(n3319) );
  NAND U3402 ( .A(x[66]), .B(y[57]), .Z(n3277) );
  XOR U3403 ( .A(n3278), .B(n3277), .Z(n3320) );
  XOR U3404 ( .A(n3319), .B(n3320), .Z(n3330) );
  XOR U3405 ( .A(n3329), .B(n3330), .Z(n3332) );
  XOR U3406 ( .A(n3331), .B(n3332), .Z(n3285) );
  XOR U3407 ( .A(n3286), .B(n3285), .Z(n3288) );
  NAND U3408 ( .A(n3280), .B(n3279), .Z(n3284) );
  NAND U3409 ( .A(n3282), .B(n3281), .Z(n3283) );
  AND U3410 ( .A(n3284), .B(n3283), .Z(n3287) );
  XOR U3411 ( .A(n3288), .B(n3287), .Z(n3293) );
  XOR U3412 ( .A(n3294), .B(n3293), .Z(o[59]) );
  NAND U3413 ( .A(n3286), .B(n3285), .Z(n3290) );
  NAND U3414 ( .A(n3288), .B(n3287), .Z(n3289) );
  NAND U3415 ( .A(n3290), .B(n3289), .Z(n3399) );
  NANDN U3416 ( .A(n3292), .B(n3291), .Z(n3296) );
  NAND U3417 ( .A(n3294), .B(n3293), .Z(n3295) );
  AND U3418 ( .A(n3296), .B(n3295), .Z(n3398) );
  AND U3419 ( .A(y[9]), .B(x[51]), .Z(n3350) );
  NAND U3420 ( .A(n3350), .B(n3297), .Z(n3301) );
  NANDN U3421 ( .A(n3299), .B(n3298), .Z(n3300) );
  AND U3422 ( .A(n3301), .B(n3300), .Z(n3377) );
  AND U3423 ( .A(x[66]), .B(y[58]), .Z(n3310) );
  NAND U3424 ( .A(x[67]), .B(y[57]), .Z(n3302) );
  XNOR U3425 ( .A(n3310), .B(n3302), .Z(n3336) );
  NAND U3426 ( .A(y[59]), .B(x[65]), .Z(n3337) );
  XNOR U3427 ( .A(n3336), .B(n3337), .Z(n3338) );
  NAND U3428 ( .A(y[56]), .B(x[68]), .Z(n3339) );
  XNOR U3429 ( .A(n3338), .B(n3339), .Z(n3374) );
  AND U3430 ( .A(x[58]), .B(y[34]), .Z(n3304) );
  NAND U3431 ( .A(x[57]), .B(y[35]), .Z(n3303) );
  XNOR U3432 ( .A(n3304), .B(n3303), .Z(n3355) );
  NAND U3433 ( .A(y[33]), .B(x[59]), .Z(n3356) );
  XOR U3434 ( .A(n3355), .B(n3356), .Z(n3375) );
  XNOR U3435 ( .A(n3374), .B(n3375), .Z(n3376) );
  XNOR U3436 ( .A(n3377), .B(n3376), .Z(n3380) );
  AND U3437 ( .A(y[34]), .B(x[59]), .Z(n3441) );
  NAND U3438 ( .A(n3441), .B(n3305), .Z(n3309) );
  NANDN U3439 ( .A(n3307), .B(n3306), .Z(n3308) );
  AND U3440 ( .A(n3309), .B(n3308), .Z(n3371) );
  AND U3441 ( .A(y[57]), .B(x[65]), .Z(n3311) );
  AND U3442 ( .A(n3311), .B(n3310), .Z(n3342) );
  NAND U3443 ( .A(y[8]), .B(x[52]), .Z(n3343) );
  XNOR U3444 ( .A(n3342), .B(n3343), .Z(n3344) );
  NAND U3445 ( .A(y[60]), .B(x[64]), .Z(n3408) );
  XNOR U3446 ( .A(n3344), .B(n3408), .Z(n3368) );
  AND U3447 ( .A(y[32]), .B(x[60]), .Z(n3456) );
  AND U3448 ( .A(y[36]), .B(x[56]), .Z(n3359) );
  XOR U3449 ( .A(n3456), .B(n3359), .Z(n3361) );
  NAND U3450 ( .A(y[11]), .B(x[49]), .Z(n3360) );
  XOR U3451 ( .A(n3361), .B(n3360), .Z(n3369) );
  XNOR U3452 ( .A(n3368), .B(n3369), .Z(n3370) );
  XOR U3453 ( .A(n3371), .B(n3370), .Z(n3381) );
  XNOR U3454 ( .A(n3380), .B(n3381), .Z(n3383) );
  NAND U3455 ( .A(n3313), .B(n3312), .Z(n3317) );
  NANDN U3456 ( .A(n3315), .B(n3314), .Z(n3316) );
  NAND U3457 ( .A(n3317), .B(n3316), .Z(n3388) );
  AND U3458 ( .A(y[10]), .B(x[50]), .Z(n3353) );
  NAND U3459 ( .A(y[12]), .B(x[48]), .Z(n3351) );
  XNOR U3460 ( .A(n3350), .B(n3351), .Z(n3352) );
  XOR U3461 ( .A(n3353), .B(n3352), .Z(n3387) );
  AND U3462 ( .A(y[59]), .B(x[67]), .Z(n3584) );
  NANDN U3463 ( .A(n3318), .B(n3584), .Z(n3322) );
  NANDN U3464 ( .A(n3320), .B(n3319), .Z(n3321) );
  NAND U3465 ( .A(n3322), .B(n3321), .Z(n3386) );
  XOR U3466 ( .A(n3387), .B(n3386), .Z(n3389) );
  XOR U3467 ( .A(n3388), .B(n3389), .Z(n3382) );
  XOR U3468 ( .A(n3383), .B(n3382), .Z(n3395) );
  NANDN U3469 ( .A(n3324), .B(n3323), .Z(n3328) );
  NANDN U3470 ( .A(n3326), .B(n3325), .Z(n3327) );
  AND U3471 ( .A(n3328), .B(n3327), .Z(n3392) );
  NANDN U3472 ( .A(n3330), .B(n3329), .Z(n3334) );
  OR U3473 ( .A(n3332), .B(n3331), .Z(n3333) );
  NAND U3474 ( .A(n3334), .B(n3333), .Z(n3393) );
  XNOR U3475 ( .A(n3392), .B(n3393), .Z(n3394) );
  XNOR U3476 ( .A(n3395), .B(n3394), .Z(n3400) );
  XNOR U3477 ( .A(n3398), .B(n3400), .Z(n3335) );
  XNOR U3478 ( .A(n3399), .B(n3335), .Z(o[60]) );
  NANDN U3479 ( .A(n3337), .B(n3336), .Z(n3341) );
  NANDN U3480 ( .A(n3339), .B(n3338), .Z(n3340) );
  AND U3481 ( .A(n3341), .B(n3340), .Z(n3432) );
  NANDN U3482 ( .A(n3343), .B(n3342), .Z(n3346) );
  NANDN U3483 ( .A(n3408), .B(n3344), .Z(n3345) );
  NAND U3484 ( .A(n3346), .B(n3345), .Z(n3437) );
  AND U3485 ( .A(x[61]), .B(y[32]), .Z(n3348) );
  NAND U3486 ( .A(x[60]), .B(y[33]), .Z(n3347) );
  XNOR U3487 ( .A(n3348), .B(n3347), .Z(n3458) );
  AND U3488 ( .A(y[12]), .B(x[49]), .Z(n3457) );
  XOR U3489 ( .A(n3458), .B(n3457), .Z(n3436) );
  AND U3490 ( .A(y[59]), .B(x[66]), .Z(n3449) );
  AND U3491 ( .A(y[56]), .B(x[69]), .Z(n3448) );
  XOR U3492 ( .A(n3449), .B(n3448), .Z(n3451) );
  AND U3493 ( .A(x[67]), .B(y[58]), .Z(n3364) );
  NAND U3494 ( .A(x[68]), .B(y[57]), .Z(n3349) );
  XNOR U3495 ( .A(n3364), .B(n3349), .Z(n3450) );
  XOR U3496 ( .A(n3451), .B(n3450), .Z(n3435) );
  XOR U3497 ( .A(n3436), .B(n3435), .Z(n3438) );
  XOR U3498 ( .A(n3437), .B(n3438), .Z(n3429) );
  XNOR U3499 ( .A(n3429), .B(n3430), .Z(n3431) );
  XOR U3500 ( .A(n3432), .B(n3431), .Z(n3471) );
  AND U3501 ( .A(y[34]), .B(x[57]), .Z(n3354) );
  AND U3502 ( .A(y[35]), .B(x[58]), .Z(n3413) );
  NAND U3503 ( .A(n3354), .B(n3413), .Z(n3358) );
  NANDN U3504 ( .A(n3356), .B(n3355), .Z(n3357) );
  AND U3505 ( .A(n3358), .B(n3357), .Z(n3422) );
  AND U3506 ( .A(y[8]), .B(x[53]), .Z(n3524) );
  NAND U3507 ( .A(y[9]), .B(x[52]), .Z(n3415) );
  XNOR U3508 ( .A(n3414), .B(n3415), .Z(n3419) );
  AND U3509 ( .A(y[36]), .B(x[57]), .Z(n3519) );
  AND U3510 ( .A(y[13]), .B(x[48]), .Z(n3401) );
  NAND U3511 ( .A(y[37]), .B(x[56]), .Z(n3402) );
  XOR U3512 ( .A(n3401), .B(n3402), .Z(n3403) );
  XOR U3513 ( .A(n3519), .B(n3403), .Z(n3420) );
  XNOR U3514 ( .A(n3419), .B(n3420), .Z(n3421) );
  XOR U3515 ( .A(n3422), .B(n3421), .Z(n3470) );
  NAND U3516 ( .A(n3456), .B(n3359), .Z(n3363) );
  ANDN U3517 ( .B(n3361), .A(n3360), .Z(n3362) );
  ANDN U3518 ( .B(n3363), .A(n3362), .Z(n3428) );
  AND U3519 ( .A(y[57]), .B(x[66]), .Z(n3365) );
  AND U3520 ( .A(n3365), .B(n3364), .Z(n3409) );
  AND U3521 ( .A(x[65]), .B(y[60]), .Z(n3367) );
  NAND U3522 ( .A(x[64]), .B(y[61]), .Z(n3366) );
  XOR U3523 ( .A(n3367), .B(n3366), .Z(n3410) );
  XNOR U3524 ( .A(n3409), .B(n3410), .Z(n3426) );
  AND U3525 ( .A(y[10]), .B(x[51]), .Z(n3531) );
  XOR U3526 ( .A(n3441), .B(n3531), .Z(n3443) );
  AND U3527 ( .A(y[11]), .B(x[50]), .Z(n3442) );
  XNOR U3528 ( .A(n3443), .B(n3442), .Z(n3425) );
  XNOR U3529 ( .A(n3426), .B(n3425), .Z(n3427) );
  XOR U3530 ( .A(n3428), .B(n3427), .Z(n3469) );
  XOR U3531 ( .A(n3470), .B(n3469), .Z(n3472) );
  NANDN U3532 ( .A(n3369), .B(n3368), .Z(n3373) );
  NANDN U3533 ( .A(n3371), .B(n3370), .Z(n3372) );
  AND U3534 ( .A(n3373), .B(n3372), .Z(n3464) );
  NANDN U3535 ( .A(n3375), .B(n3374), .Z(n3379) );
  NANDN U3536 ( .A(n3377), .B(n3376), .Z(n3378) );
  NAND U3537 ( .A(n3379), .B(n3378), .Z(n3463) );
  XOR U3538 ( .A(n3464), .B(n3463), .Z(n3466) );
  XNOR U3539 ( .A(n3465), .B(n3466), .Z(n3477) );
  NANDN U3540 ( .A(n3381), .B(n3380), .Z(n3385) );
  NAND U3541 ( .A(n3383), .B(n3382), .Z(n3384) );
  AND U3542 ( .A(n3385), .B(n3384), .Z(n3475) );
  NAND U3543 ( .A(n3387), .B(n3386), .Z(n3391) );
  NAND U3544 ( .A(n3389), .B(n3388), .Z(n3390) );
  NAND U3545 ( .A(n3391), .B(n3390), .Z(n3476) );
  XNOR U3546 ( .A(n3475), .B(n3476), .Z(n3478) );
  XNOR U3547 ( .A(n3477), .B(n3478), .Z(n3482) );
  NANDN U3548 ( .A(n3393), .B(n3392), .Z(n3397) );
  NANDN U3549 ( .A(n3395), .B(n3394), .Z(n3396) );
  AND U3550 ( .A(n3397), .B(n3396), .Z(n3480) );
  XNOR U3551 ( .A(n3480), .B(n3479), .Z(n3481) );
  XNOR U3552 ( .A(n3482), .B(n3481), .Z(o[61]) );
  NANDN U3553 ( .A(n3402), .B(n3401), .Z(n3405) );
  NANDN U3554 ( .A(n3403), .B(n3519), .Z(n3404) );
  AND U3555 ( .A(n3405), .B(n3404), .Z(n3503) );
  AND U3556 ( .A(x[53]), .B(y[9]), .Z(n3407) );
  NAND U3557 ( .A(x[54]), .B(y[8]), .Z(n3406) );
  XNOR U3558 ( .A(n3407), .B(n3406), .Z(n3523) );
  AND U3559 ( .A(y[35]), .B(x[59]), .Z(n3522) );
  XNOR U3560 ( .A(n3523), .B(n3522), .Z(n3506) );
  AND U3561 ( .A(y[13]), .B(x[49]), .Z(n3535) );
  AND U3562 ( .A(y[62]), .B(x[64]), .Z(n3537) );
  AND U3563 ( .A(y[38]), .B(x[56]), .Z(n3536) );
  XOR U3564 ( .A(n3537), .B(n3536), .Z(n3534) );
  XNOR U3565 ( .A(n3535), .B(n3534), .Z(n3505) );
  XNOR U3566 ( .A(n3503), .B(n3504), .Z(n3610) );
  AND U3567 ( .A(y[61]), .B(x[65]), .Z(n3567) );
  NANDN U3568 ( .A(n3408), .B(n3567), .Z(n3412) );
  NANDN U3569 ( .A(n3410), .B(n3409), .Z(n3411) );
  AND U3570 ( .A(n3412), .B(n3411), .Z(n3612) );
  NAND U3571 ( .A(n3524), .B(n3413), .Z(n3417) );
  NANDN U3572 ( .A(n3415), .B(n3414), .Z(n3416) );
  AND U3573 ( .A(n3417), .B(n3416), .Z(n3511) );
  AND U3574 ( .A(y[33]), .B(x[61]), .Z(n3593) );
  AND U3575 ( .A(y[32]), .B(x[62]), .Z(n3595) );
  AND U3576 ( .A(y[14]), .B(x[48]), .Z(n3594) );
  XOR U3577 ( .A(n3595), .B(n3594), .Z(n3592) );
  XNOR U3578 ( .A(n3593), .B(n3592), .Z(n3514) );
  AND U3579 ( .A(y[58]), .B(x[68]), .Z(n3461) );
  NAND U3580 ( .A(x[69]), .B(y[57]), .Z(n3418) );
  XNOR U3581 ( .A(n3461), .B(n3418), .Z(n3587) );
  AND U3582 ( .A(y[56]), .B(x[70]), .Z(n3586) );
  XOR U3583 ( .A(n3587), .B(n3586), .Z(n3585) );
  XNOR U3584 ( .A(n3585), .B(n3584), .Z(n3513) );
  XNOR U3585 ( .A(n3511), .B(n3512), .Z(n3611) );
  XOR U3586 ( .A(n3612), .B(n3611), .Z(n3609) );
  XNOR U3587 ( .A(n3610), .B(n3609), .Z(n3624) );
  NANDN U3588 ( .A(n3420), .B(n3419), .Z(n3424) );
  NANDN U3589 ( .A(n3422), .B(n3421), .Z(n3423) );
  NAND U3590 ( .A(n3424), .B(n3423), .Z(n3626) );
  XOR U3591 ( .A(n3626), .B(n3625), .Z(n3623) );
  NANDN U3592 ( .A(n3430), .B(n3429), .Z(n3434) );
  NANDN U3593 ( .A(n3432), .B(n3431), .Z(n3433) );
  AND U3594 ( .A(n3434), .B(n3433), .Z(n3638) );
  NAND U3595 ( .A(n3436), .B(n3435), .Z(n3440) );
  NAND U3596 ( .A(n3438), .B(n3437), .Z(n3439) );
  AND U3597 ( .A(n3440), .B(n3439), .Z(n3620) );
  NAND U3598 ( .A(n3441), .B(n3531), .Z(n3445) );
  NAND U3599 ( .A(n3443), .B(n3442), .Z(n3444) );
  AND U3600 ( .A(n3445), .B(n3444), .Z(n3498) );
  AND U3601 ( .A(x[57]), .B(y[37]), .Z(n3447) );
  NAND U3602 ( .A(x[58]), .B(y[36]), .Z(n3446) );
  XNOR U3603 ( .A(n3447), .B(n3446), .Z(n3518) );
  AND U3604 ( .A(y[12]), .B(x[50]), .Z(n3517) );
  XNOR U3605 ( .A(n3518), .B(n3517), .Z(n3500) );
  NAND U3606 ( .A(n3449), .B(n3448), .Z(n3453) );
  NAND U3607 ( .A(n3451), .B(n3450), .Z(n3452) );
  AND U3608 ( .A(n3453), .B(n3452), .Z(n3499) );
  XOR U3609 ( .A(n3498), .B(n3497), .Z(n3619) );
  XOR U3610 ( .A(n3620), .B(n3619), .Z(n3618) );
  AND U3611 ( .A(x[52]), .B(y[10]), .Z(n3455) );
  NAND U3612 ( .A(x[51]), .B(y[11]), .Z(n3454) );
  XNOR U3613 ( .A(n3455), .B(n3454), .Z(n3530) );
  AND U3614 ( .A(y[34]), .B(x[60]), .Z(n3529) );
  XNOR U3615 ( .A(n3530), .B(n3529), .Z(n3494) );
  NAND U3616 ( .A(n3456), .B(n3593), .Z(n3460) );
  NAND U3617 ( .A(n3458), .B(n3457), .Z(n3459) );
  AND U3618 ( .A(n3460), .B(n3459), .Z(n3493) );
  AND U3619 ( .A(y[57]), .B(x[67]), .Z(n3462) );
  AND U3620 ( .A(n3462), .B(n3461), .Z(n3569) );
  AND U3621 ( .A(y[60]), .B(x[66]), .Z(n3568) );
  XOR U3622 ( .A(n3569), .B(n3568), .Z(n3566) );
  XNOR U3623 ( .A(n3567), .B(n3566), .Z(n3492) );
  XOR U3624 ( .A(n3618), .B(n3617), .Z(n3637) );
  XOR U3625 ( .A(n3638), .B(n3637), .Z(n3635) );
  XNOR U3626 ( .A(n3636), .B(n3635), .Z(n3641) );
  NANDN U3627 ( .A(n3464), .B(n3463), .Z(n3468) );
  NANDN U3628 ( .A(n3466), .B(n3465), .Z(n3467) );
  NAND U3629 ( .A(n3468), .B(n3467), .Z(n3643) );
  NAND U3630 ( .A(n3470), .B(n3469), .Z(n3474) );
  NAND U3631 ( .A(n3472), .B(n3471), .Z(n3473) );
  AND U3632 ( .A(n3474), .B(n3473), .Z(n3644) );
  XOR U3633 ( .A(n3643), .B(n3644), .Z(n3642) );
  XOR U3634 ( .A(n3488), .B(n3487), .Z(n3486) );
  NANDN U3635 ( .A(n3480), .B(n3479), .Z(n3484) );
  NAND U3636 ( .A(n3482), .B(n3481), .Z(n3483) );
  NAND U3637 ( .A(n3484), .B(n3483), .Z(n3485) );
  XNOR U3638 ( .A(n3486), .B(n3485), .Z(o[62]) );
  NAND U3639 ( .A(n3486), .B(n3485), .Z(n3490) );
  NAND U3640 ( .A(n3488), .B(n3487), .Z(n3489) );
  AND U3641 ( .A(n3490), .B(n3489), .Z(n3634) );
  NAND U3642 ( .A(n3492), .B(n3491), .Z(n3496) );
  NAND U3643 ( .A(n3494), .B(n3493), .Z(n3495) );
  AND U3644 ( .A(n3496), .B(n3495), .Z(n3608) );
  NAND U3645 ( .A(n3498), .B(n3497), .Z(n3502) );
  NAND U3646 ( .A(n3500), .B(n3499), .Z(n3501) );
  AND U3647 ( .A(n3502), .B(n3501), .Z(n3510) );
  NANDN U3648 ( .A(n3504), .B(n3503), .Z(n3508) );
  NAND U3649 ( .A(n3506), .B(n3505), .Z(n3507) );
  NAND U3650 ( .A(n3508), .B(n3507), .Z(n3509) );
  XNOR U3651 ( .A(n3510), .B(n3509), .Z(n3606) );
  NANDN U3652 ( .A(n3512), .B(n3511), .Z(n3516) );
  NAND U3653 ( .A(n3514), .B(n3513), .Z(n3515) );
  AND U3654 ( .A(n3516), .B(n3515), .Z(n3604) );
  NAND U3655 ( .A(n3518), .B(n3517), .Z(n3521) );
  AND U3656 ( .A(y[37]), .B(x[58]), .Z(n3553) );
  NAND U3657 ( .A(n3519), .B(n3553), .Z(n3520) );
  AND U3658 ( .A(n3521), .B(n3520), .Z(n3528) );
  NAND U3659 ( .A(n3523), .B(n3522), .Z(n3526) );
  AND U3660 ( .A(y[9]), .B(x[54]), .Z(n3596) );
  NAND U3661 ( .A(n3524), .B(n3596), .Z(n3525) );
  NAND U3662 ( .A(n3526), .B(n3525), .Z(n3527) );
  XNOR U3663 ( .A(n3528), .B(n3527), .Z(n3543) );
  NAND U3664 ( .A(n3530), .B(n3529), .Z(n3533) );
  AND U3665 ( .A(y[11]), .B(x[52]), .Z(n3552) );
  NAND U3666 ( .A(n3531), .B(n3552), .Z(n3532) );
  AND U3667 ( .A(n3533), .B(n3532), .Z(n3541) );
  NAND U3668 ( .A(n3535), .B(n3534), .Z(n3539) );
  NAND U3669 ( .A(n3537), .B(n3536), .Z(n3538) );
  NAND U3670 ( .A(n3539), .B(n3538), .Z(n3540) );
  XNOR U3671 ( .A(n3541), .B(n3540), .Z(n3542) );
  XOR U3672 ( .A(n3543), .B(n3542), .Z(n3583) );
  AND U3673 ( .A(x[63]), .B(y[32]), .Z(n3545) );
  NAND U3674 ( .A(x[55]), .B(y[8]), .Z(n3544) );
  XNOR U3675 ( .A(n3545), .B(n3544), .Z(n3557) );
  AND U3676 ( .A(x[48]), .B(y[15]), .Z(n3547) );
  NAND U3677 ( .A(x[67]), .B(y[60]), .Z(n3546) );
  XNOR U3678 ( .A(n3547), .B(n3546), .Z(n3551) );
  AND U3679 ( .A(x[53]), .B(y[10]), .Z(n3549) );
  NAND U3680 ( .A(x[66]), .B(y[61]), .Z(n3548) );
  XNOR U3681 ( .A(n3549), .B(n3548), .Z(n3550) );
  XOR U3682 ( .A(n3551), .B(n3550), .Z(n3555) );
  XNOR U3683 ( .A(n3553), .B(n3552), .Z(n3554) );
  XNOR U3684 ( .A(n3555), .B(n3554), .Z(n3556) );
  XOR U3685 ( .A(n3557), .B(n3556), .Z(n3565) );
  AND U3686 ( .A(x[71]), .B(y[56]), .Z(n3559) );
  NAND U3687 ( .A(x[60]), .B(y[35]), .Z(n3558) );
  XNOR U3688 ( .A(n3559), .B(n3558), .Z(n3563) );
  AND U3689 ( .A(x[59]), .B(y[36]), .Z(n3561) );
  NAND U3690 ( .A(x[61]), .B(y[34]), .Z(n3560) );
  XNOR U3691 ( .A(n3561), .B(n3560), .Z(n3562) );
  XNOR U3692 ( .A(n3563), .B(n3562), .Z(n3564) );
  XNOR U3693 ( .A(n3565), .B(n3564), .Z(n3581) );
  NAND U3694 ( .A(n3567), .B(n3566), .Z(n3571) );
  NAND U3695 ( .A(n3569), .B(n3568), .Z(n3570) );
  AND U3696 ( .A(n3571), .B(n3570), .Z(n3579) );
  AND U3697 ( .A(x[65]), .B(y[62]), .Z(n3573) );
  NAND U3698 ( .A(x[62]), .B(y[33]), .Z(n3572) );
  XNOR U3699 ( .A(n3573), .B(n3572), .Z(n3577) );
  AND U3700 ( .A(x[57]), .B(y[38]), .Z(n3575) );
  NAND U3701 ( .A(x[50]), .B(y[13]), .Z(n3574) );
  XNOR U3702 ( .A(n3575), .B(n3574), .Z(n3576) );
  XNOR U3703 ( .A(n3577), .B(n3576), .Z(n3578) );
  XNOR U3704 ( .A(n3579), .B(n3578), .Z(n3580) );
  XNOR U3705 ( .A(n3581), .B(n3580), .Z(n3582) );
  XNOR U3706 ( .A(n3583), .B(n3582), .Z(n3602) );
  NAND U3707 ( .A(n3585), .B(n3584), .Z(n3589) );
  NAND U3708 ( .A(n3587), .B(n3586), .Z(n3588) );
  AND U3709 ( .A(n3589), .B(n3588), .Z(n3600) );
  AND U3710 ( .A(x[64]), .B(y[63]), .Z(n3591) );
  NAND U3711 ( .A(x[51]), .B(y[12]), .Z(n3590) );
  XNOR U3712 ( .A(n3591), .B(n3590), .Z(n3598) );
  XNOR U3713 ( .A(n3598), .B(n3597), .Z(n3599) );
  XNOR U3714 ( .A(n3600), .B(n3599), .Z(n3601) );
  XNOR U3715 ( .A(n3602), .B(n3601), .Z(n3603) );
  XNOR U3716 ( .A(n3604), .B(n3603), .Z(n3605) );
  XNOR U3717 ( .A(n3606), .B(n3605), .Z(n3607) );
  XNOR U3718 ( .A(n3608), .B(n3607), .Z(n3616) );
  NAND U3719 ( .A(n3610), .B(n3609), .Z(n3614) );
  NAND U3720 ( .A(n3612), .B(n3611), .Z(n3613) );
  NAND U3721 ( .A(n3614), .B(n3613), .Z(n3615) );
  XNOR U3722 ( .A(n3616), .B(n3615), .Z(n3632) );
  NAND U3723 ( .A(n3618), .B(n3617), .Z(n3622) );
  NAND U3724 ( .A(n3620), .B(n3619), .Z(n3621) );
  AND U3725 ( .A(n3622), .B(n3621), .Z(n3630) );
  NAND U3726 ( .A(n3624), .B(n3623), .Z(n3628) );
  NAND U3727 ( .A(n3626), .B(n3625), .Z(n3627) );
  NAND U3728 ( .A(n3628), .B(n3627), .Z(n3629) );
  XNOR U3729 ( .A(n3630), .B(n3629), .Z(n3631) );
  XNOR U3730 ( .A(n3632), .B(n3631), .Z(n3633) );
  XNOR U3731 ( .A(n3634), .B(n3633), .Z(n3650) );
  NAND U3732 ( .A(n3636), .B(n3635), .Z(n3640) );
  NAND U3733 ( .A(n3638), .B(n3637), .Z(n3639) );
  AND U3734 ( .A(n3640), .B(n3639), .Z(n3648) );
  NAND U3735 ( .A(n3642), .B(n3641), .Z(n3646) );
  NAND U3736 ( .A(n3644), .B(n3643), .Z(n3645) );
  NAND U3737 ( .A(n3646), .B(n3645), .Z(n3647) );
  XNOR U3738 ( .A(n3648), .B(n3647), .Z(n3649) );
  XNOR U3739 ( .A(n3650), .B(n3649), .Z(o[63]) );
  AND U3740 ( .A(y[40]), .B(x[56]), .Z(n3652) );
  NAND U3741 ( .A(y[16]), .B(x[48]), .Z(n3651) );
  XNOR U3742 ( .A(n3652), .B(n3651), .Z(n3653) );
  NAND U3743 ( .A(y[64]), .B(x[64]), .Z(n3730) );
  XNOR U3744 ( .A(n3653), .B(n3730), .Z(o[64]) );
  AND U3745 ( .A(y[17]), .B(x[48]), .Z(n3692) );
  AND U3746 ( .A(y[65]), .B(x[64]), .Z(n3700) );
  AND U3747 ( .A(y[16]), .B(x[49]), .Z(n3668) );
  XOR U3748 ( .A(n3700), .B(n3668), .Z(n3669) );
  XOR U3749 ( .A(n3692), .B(n3669), .Z(n3656) );
  NANDN U3750 ( .A(n3652), .B(n3651), .Z(n3655) );
  NAND U3751 ( .A(n3730), .B(n3653), .Z(n3654) );
  NAND U3752 ( .A(n3655), .B(n3654), .Z(n3657) );
  XNOR U3753 ( .A(n3656), .B(n3657), .Z(n3659) );
  AND U3754 ( .A(y[40]), .B(x[57]), .Z(n3717) );
  AND U3755 ( .A(y[64]), .B(x[65]), .Z(n3772) );
  AND U3756 ( .A(y[41]), .B(x[56]), .Z(n3664) );
  XOR U3757 ( .A(n3772), .B(n3664), .Z(n3665) );
  XOR U3758 ( .A(n3717), .B(n3665), .Z(n3658) );
  XOR U3759 ( .A(n3659), .B(n3658), .Z(o[65]) );
  NANDN U3760 ( .A(n3657), .B(n3656), .Z(n3661) );
  NAND U3761 ( .A(n3659), .B(n3658), .Z(n3660) );
  AND U3762 ( .A(n3661), .B(n3660), .Z(n3679) );
  AND U3763 ( .A(x[49]), .B(y[17]), .Z(n3663) );
  NAND U3764 ( .A(x[48]), .B(y[18]), .Z(n3662) );
  XNOR U3765 ( .A(n3663), .B(n3662), .Z(n3694) );
  AND U3766 ( .A(y[40]), .B(x[58]), .Z(n3693) );
  XOR U3767 ( .A(n3694), .B(n3693), .Z(n3704) );
  AND U3768 ( .A(y[42]), .B(x[56]), .Z(n3702) );
  NAND U3769 ( .A(y[41]), .B(x[57]), .Z(n3701) );
  XNOR U3770 ( .A(n3702), .B(n3701), .Z(n3703) );
  XOR U3771 ( .A(n3704), .B(n3703), .Z(n3680) );
  XNOR U3772 ( .A(n3679), .B(n3680), .Z(n3682) );
  NAND U3773 ( .A(n3772), .B(n3664), .Z(n3667) );
  NAND U3774 ( .A(n3717), .B(n3665), .Z(n3666) );
  NAND U3775 ( .A(n3667), .B(n3666), .Z(n3675) );
  NAND U3776 ( .A(n3700), .B(n3668), .Z(n3671) );
  NAND U3777 ( .A(n3692), .B(n3669), .Z(n3670) );
  NAND U3778 ( .A(n3671), .B(n3670), .Z(n3673) );
  AND U3779 ( .A(y[16]), .B(x[50]), .Z(n3707) );
  NAND U3780 ( .A(y[64]), .B(x[66]), .Z(n3685) );
  XNOR U3781 ( .A(n3707), .B(n3685), .Z(n3687) );
  AND U3782 ( .A(x[65]), .B(y[65]), .Z(n3722) );
  NAND U3783 ( .A(x[64]), .B(y[66]), .Z(n3672) );
  XNOR U3784 ( .A(n3722), .B(n3672), .Z(n3686) );
  XOR U3785 ( .A(n3687), .B(n3686), .Z(n3674) );
  XNOR U3786 ( .A(n3673), .B(n3674), .Z(n3676) );
  XOR U3787 ( .A(n3675), .B(n3676), .Z(n3681) );
  XNOR U3788 ( .A(n3682), .B(n3681), .Z(o[66]) );
  NAND U3789 ( .A(n3674), .B(n3673), .Z(n3678) );
  NANDN U3790 ( .A(n3676), .B(n3675), .Z(n3677) );
  AND U3791 ( .A(n3678), .B(n3677), .Z(n3754) );
  NANDN U3792 ( .A(n3680), .B(n3679), .Z(n3684) );
  NAND U3793 ( .A(n3682), .B(n3681), .Z(n3683) );
  AND U3794 ( .A(n3684), .B(n3683), .Z(n3753) );
  XNOR U3795 ( .A(n3754), .B(n3753), .Z(n3756) );
  NANDN U3796 ( .A(n3685), .B(n3707), .Z(n3689) );
  NAND U3797 ( .A(n3687), .B(n3686), .Z(n3688) );
  NAND U3798 ( .A(n3689), .B(n3688), .Z(n3739) );
  AND U3799 ( .A(y[43]), .B(x[56]), .Z(n3724) );
  AND U3800 ( .A(y[18]), .B(x[49]), .Z(n3725) );
  AND U3801 ( .A(y[19]), .B(x[48]), .Z(n3727) );
  AND U3802 ( .A(x[59]), .B(y[40]), .Z(n3691) );
  NAND U3803 ( .A(x[57]), .B(y[42]), .Z(n3690) );
  XNOR U3804 ( .A(n3691), .B(n3690), .Z(n3719) );
  AND U3805 ( .A(y[41]), .B(x[58]), .Z(n3718) );
  XOR U3806 ( .A(n3719), .B(n3718), .Z(n3737) );
  XOR U3807 ( .A(n3738), .B(n3737), .Z(n3740) );
  XOR U3808 ( .A(n3739), .B(n3740), .Z(n3750) );
  NAND U3809 ( .A(n3725), .B(n3692), .Z(n3696) );
  NAND U3810 ( .A(n3694), .B(n3693), .Z(n3695) );
  NAND U3811 ( .A(n3696), .B(n3695), .Z(n3745) );
  AND U3812 ( .A(x[66]), .B(y[65]), .Z(n3804) );
  AND U3813 ( .A(y[66]), .B(x[65]), .Z(n3699) );
  XNOR U3814 ( .A(n3804), .B(n3699), .Z(n3733) );
  AND U3815 ( .A(x[50]), .B(y[17]), .Z(n3698) );
  NAND U3816 ( .A(x[51]), .B(y[16]), .Z(n3697) );
  XNOR U3817 ( .A(n3698), .B(n3697), .Z(n3709) );
  AND U3818 ( .A(n3700), .B(n3699), .Z(n3708) );
  XOR U3819 ( .A(n3709), .B(n3708), .Z(n3743) );
  XOR U3820 ( .A(n3744), .B(n3743), .Z(n3746) );
  XNOR U3821 ( .A(n3745), .B(n3746), .Z(n3749) );
  XNOR U3822 ( .A(n3750), .B(n3749), .Z(n3751) );
  NANDN U3823 ( .A(n3702), .B(n3701), .Z(n3706) );
  NANDN U3824 ( .A(n3704), .B(n3703), .Z(n3705) );
  NAND U3825 ( .A(n3706), .B(n3705), .Z(n3752) );
  XNOR U3826 ( .A(n3751), .B(n3752), .Z(n3755) );
  XOR U3827 ( .A(n3756), .B(n3755), .Z(o[67]) );
  NAND U3828 ( .A(y[17]), .B(x[51]), .Z(n3788) );
  NANDN U3829 ( .A(n3788), .B(n3707), .Z(n3711) );
  NAND U3830 ( .A(n3709), .B(n3708), .Z(n3710) );
  NAND U3831 ( .A(n3711), .B(n3710), .Z(n3763) );
  AND U3832 ( .A(x[57]), .B(y[43]), .Z(n3713) );
  NAND U3833 ( .A(x[58]), .B(y[42]), .Z(n3712) );
  XNOR U3834 ( .A(n3713), .B(n3712), .Z(n3792) );
  NAND U3835 ( .A(y[41]), .B(x[59]), .Z(n3793) );
  XNOR U3836 ( .A(n3792), .B(n3793), .Z(n3761) );
  AND U3837 ( .A(x[68]), .B(y[64]), .Z(n3715) );
  NAND U3838 ( .A(x[65]), .B(y[67]), .Z(n3714) );
  XNOR U3839 ( .A(n3715), .B(n3714), .Z(n3773) );
  AND U3840 ( .A(x[67]), .B(y[65]), .Z(n3885) );
  NAND U3841 ( .A(x[66]), .B(y[66]), .Z(n3716) );
  XNOR U3842 ( .A(n3885), .B(n3716), .Z(n3774) );
  XOR U3843 ( .A(n3761), .B(n3760), .Z(n3762) );
  NAND U3844 ( .A(y[42]), .B(x[59]), .Z(n3805) );
  IV U3845 ( .A(n3805), .Z(n3867) );
  NAND U3846 ( .A(n3867), .B(n3717), .Z(n3721) );
  NAND U3847 ( .A(n3719), .B(n3718), .Z(n3720) );
  NAND U3848 ( .A(n3721), .B(n3720), .Z(n3769) );
  AND U3849 ( .A(y[68]), .B(x[64]), .Z(n3838) );
  AND U3850 ( .A(y[66]), .B(x[66]), .Z(n3723) );
  AND U3851 ( .A(n3723), .B(n3722), .Z(n3777) );
  NAND U3852 ( .A(y[16]), .B(x[52]), .Z(n3778) );
  XOR U3853 ( .A(n3777), .B(n3778), .Z(n3779) );
  XNOR U3854 ( .A(n3838), .B(n3779), .Z(n3766) );
  AND U3855 ( .A(y[40]), .B(x[60]), .Z(n3881) );
  AND U3856 ( .A(y[44]), .B(x[56]), .Z(n3796) );
  XOR U3857 ( .A(n3881), .B(n3796), .Z(n3797) );
  NAND U3858 ( .A(y[19]), .B(x[49]), .Z(n3798) );
  XNOR U3859 ( .A(n3797), .B(n3798), .Z(n3767) );
  XOR U3860 ( .A(n3807), .B(n3806), .Z(n3809) );
  NAND U3861 ( .A(n3725), .B(n3724), .Z(n3729) );
  NAND U3862 ( .A(n3727), .B(n3726), .Z(n3728) );
  NAND U3863 ( .A(n3729), .B(n3728), .Z(n3814) );
  AND U3864 ( .A(y[67]), .B(x[67]), .Z(n3933) );
  NANDN U3865 ( .A(n3730), .B(n3933), .Z(n3736) );
  NAND U3866 ( .A(x[67]), .B(y[64]), .Z(n3732) );
  NAND U3867 ( .A(x[64]), .B(y[67]), .Z(n3731) );
  AND U3868 ( .A(n3732), .B(n3731), .Z(n3734) );
  OR U3869 ( .A(n3734), .B(n3733), .Z(n3735) );
  AND U3870 ( .A(n3736), .B(n3735), .Z(n3813) );
  AND U3871 ( .A(y[18]), .B(x[50]), .Z(n3786) );
  NAND U3872 ( .A(y[20]), .B(x[48]), .Z(n3787) );
  XOR U3873 ( .A(n3788), .B(n3787), .Z(n3785) );
  XOR U3874 ( .A(n3786), .B(n3785), .Z(n3812) );
  XNOR U3875 ( .A(n3813), .B(n3812), .Z(n3815) );
  XOR U3876 ( .A(n3814), .B(n3815), .Z(n3808) );
  XOR U3877 ( .A(n3809), .B(n3808), .Z(n3821) );
  NAND U3878 ( .A(n3738), .B(n3737), .Z(n3742) );
  NAND U3879 ( .A(n3740), .B(n3739), .Z(n3741) );
  AND U3880 ( .A(n3742), .B(n3741), .Z(n3819) );
  NAND U3881 ( .A(n3744), .B(n3743), .Z(n3748) );
  NAND U3882 ( .A(n3746), .B(n3745), .Z(n3747) );
  AND U3883 ( .A(n3748), .B(n3747), .Z(n3818) );
  XOR U3884 ( .A(n3819), .B(n3818), .Z(n3820) );
  XOR U3885 ( .A(n3821), .B(n3820), .Z(n3826) );
  NANDN U3886 ( .A(n3754), .B(n3753), .Z(n3758) );
  NAND U3887 ( .A(n3756), .B(n3755), .Z(n3757) );
  AND U3888 ( .A(n3758), .B(n3757), .Z(n3824) );
  XNOR U3889 ( .A(n3825), .B(n3824), .Z(n3759) );
  XNOR U3890 ( .A(n3826), .B(n3759), .Z(o[68]) );
  NAND U3891 ( .A(n3761), .B(n3760), .Z(n3765) );
  NAND U3892 ( .A(n3763), .B(n3762), .Z(n3764) );
  AND U3893 ( .A(n3765), .B(n3764), .Z(n3892) );
  NAND U3894 ( .A(n3767), .B(n3766), .Z(n3771) );
  NAND U3895 ( .A(n3769), .B(n3768), .Z(n3770) );
  AND U3896 ( .A(n3771), .B(n3770), .Z(n3893) );
  AND U3897 ( .A(y[67]), .B(x[68]), .Z(n4023) );
  NAND U3898 ( .A(n4023), .B(n3772), .Z(n3776) );
  NAND U3899 ( .A(n3774), .B(n3773), .Z(n3775) );
  NAND U3900 ( .A(n3776), .B(n3775), .Z(n3859) );
  NANDN U3901 ( .A(n3778), .B(n3777), .Z(n3781) );
  NANDN U3902 ( .A(n3779), .B(n3838), .Z(n3780) );
  AND U3903 ( .A(n3781), .B(n3780), .Z(n3865) );
  AND U3904 ( .A(x[60]), .B(y[41]), .Z(n3783) );
  NAND U3905 ( .A(x[61]), .B(y[40]), .Z(n3782) );
  XNOR U3906 ( .A(n3783), .B(n3782), .Z(n3883) );
  NAND U3907 ( .A(y[20]), .B(x[49]), .Z(n3882) );
  XNOR U3908 ( .A(n3883), .B(n3882), .Z(n3864) );
  AND U3909 ( .A(y[67]), .B(x[66]), .Z(n3873) );
  NAND U3910 ( .A(y[64]), .B(x[69]), .Z(n3872) );
  XNOR U3911 ( .A(n3873), .B(n3872), .Z(n3876) );
  AND U3912 ( .A(y[65]), .B(x[68]), .Z(n4005) );
  NAND U3913 ( .A(x[67]), .B(y[66]), .Z(n3784) );
  XNOR U3914 ( .A(n4005), .B(n3784), .Z(n3875) );
  XNOR U3915 ( .A(n3876), .B(n3875), .Z(n3863) );
  XNOR U3916 ( .A(n3864), .B(n3863), .Z(n3866) );
  XNOR U3917 ( .A(n3865), .B(n3866), .Z(n3858) );
  NANDN U3918 ( .A(n3786), .B(n3785), .Z(n3790) );
  AND U3919 ( .A(n3788), .B(n3787), .Z(n3789) );
  ANDN U3920 ( .B(n3790), .A(n3789), .Z(n3857) );
  XOR U3921 ( .A(n3858), .B(n3857), .Z(n3860) );
  XNOR U3922 ( .A(n3859), .B(n3860), .Z(n3888) );
  AND U3923 ( .A(y[43]), .B(x[58]), .Z(n3842) );
  AND U3924 ( .A(y[42]), .B(x[57]), .Z(n3791) );
  NAND U3925 ( .A(n3842), .B(n3791), .Z(n3795) );
  NANDN U3926 ( .A(n3793), .B(n3792), .Z(n3794) );
  NAND U3927 ( .A(n3795), .B(n3794), .Z(n3850) );
  NAND U3928 ( .A(y[16]), .B(x[53]), .Z(n3841) );
  XNOR U3929 ( .A(n3842), .B(n3841), .Z(n3844) );
  NAND U3930 ( .A(y[17]), .B(x[52]), .Z(n3843) );
  XNOR U3931 ( .A(n3844), .B(n3843), .Z(n3848) );
  AND U3932 ( .A(y[44]), .B(x[57]), .Z(n3995) );
  AND U3933 ( .A(y[21]), .B(x[48]), .Z(n3834) );
  AND U3934 ( .A(y[45]), .B(x[56]), .Z(n3833) );
  XNOR U3935 ( .A(n3834), .B(n3833), .Z(n3835) );
  XNOR U3936 ( .A(n3995), .B(n3835), .Z(n3847) );
  XNOR U3937 ( .A(n3848), .B(n3847), .Z(n3849) );
  XOR U3938 ( .A(n3850), .B(n3849), .Z(n3887) );
  AND U3939 ( .A(n3881), .B(n3796), .Z(n3800) );
  NANDN U3940 ( .A(n3798), .B(n3797), .Z(n3799) );
  NANDN U3941 ( .A(n3800), .B(n3799), .Z(n3853) );
  AND U3942 ( .A(x[65]), .B(y[68]), .Z(n3802) );
  NAND U3943 ( .A(x[64]), .B(y[69]), .Z(n3801) );
  XNOR U3944 ( .A(n3802), .B(n3801), .Z(n3840) );
  AND U3945 ( .A(y[66]), .B(x[67]), .Z(n3803) );
  NAND U3946 ( .A(n3804), .B(n3803), .Z(n3839) );
  XNOR U3947 ( .A(n3840), .B(n3839), .Z(n3852) );
  AND U3948 ( .A(y[18]), .B(x[51]), .Z(n3989) );
  XNOR U3949 ( .A(n3989), .B(n3805), .Z(n3869) );
  NAND U3950 ( .A(y[19]), .B(x[50]), .Z(n3868) );
  XNOR U3951 ( .A(n3869), .B(n3868), .Z(n3851) );
  XNOR U3952 ( .A(n3852), .B(n3851), .Z(n3854) );
  XOR U3953 ( .A(n3853), .B(n3854), .Z(n3886) );
  XOR U3954 ( .A(n3887), .B(n3886), .Z(n3889) );
  XOR U3955 ( .A(n3888), .B(n3889), .Z(n3894) );
  XOR U3956 ( .A(n3895), .B(n3894), .Z(n3901) );
  NAND U3957 ( .A(n3807), .B(n3806), .Z(n3811) );
  NAND U3958 ( .A(n3809), .B(n3808), .Z(n3810) );
  AND U3959 ( .A(n3811), .B(n3810), .Z(n3898) );
  NANDN U3960 ( .A(n3813), .B(n3812), .Z(n3817) );
  NAND U3961 ( .A(n3815), .B(n3814), .Z(n3816) );
  AND U3962 ( .A(n3817), .B(n3816), .Z(n3899) );
  XOR U3963 ( .A(n3901), .B(n3900), .Z(n3830) );
  NAND U3964 ( .A(n3819), .B(n3818), .Z(n3823) );
  NANDN U3965 ( .A(n3821), .B(n3820), .Z(n3822) );
  AND U3966 ( .A(n3823), .B(n3822), .Z(n3828) );
  XNOR U3967 ( .A(n3828), .B(n3827), .Z(n3829) );
  XNOR U3968 ( .A(n3830), .B(n3829), .Z(o[69]) );
  NANDN U3969 ( .A(n3828), .B(n3827), .Z(n3832) );
  NAND U3970 ( .A(n3830), .B(n3829), .Z(n3831) );
  AND U3971 ( .A(n3832), .B(n3831), .Z(n4053) );
  AND U3972 ( .A(x[53]), .B(y[17]), .Z(n3837) );
  NAND U3973 ( .A(x[54]), .B(y[16]), .Z(n3836) );
  XNOR U3974 ( .A(n3837), .B(n3836), .Z(n3980) );
  AND U3975 ( .A(y[43]), .B(x[59]), .Z(n3979) );
  XNOR U3976 ( .A(n3980), .B(n3979), .Z(n3927) );
  AND U3977 ( .A(y[21]), .B(x[49]), .Z(n4007) );
  AND U3978 ( .A(y[70]), .B(x[64]), .Z(n4009) );
  AND U3979 ( .A(y[46]), .B(x[56]), .Z(n4008) );
  XOR U3980 ( .A(n4009), .B(n4008), .Z(n4006) );
  XNOR U3981 ( .A(n4007), .B(n4006), .Z(n3926) );
  XNOR U3982 ( .A(n3924), .B(n3925), .Z(n3905) );
  AND U3983 ( .A(y[69]), .B(x[65]), .Z(n3939) );
  IV U3984 ( .A(n3841), .Z(n3981) );
  AND U3985 ( .A(y[41]), .B(x[61]), .Z(n3974) );
  AND U3986 ( .A(y[40]), .B(x[62]), .Z(n3976) );
  AND U3987 ( .A(y[22]), .B(x[48]), .Z(n3975) );
  XOR U3988 ( .A(n3976), .B(n3975), .Z(n3973) );
  XNOR U3989 ( .A(n3974), .B(n3973), .Z(n3911) );
  AND U3990 ( .A(x[69]), .B(y[65]), .Z(n3846) );
  NAND U3991 ( .A(x[68]), .B(y[66]), .Z(n3845) );
  XNOR U3992 ( .A(n3846), .B(n3845), .Z(n3935) );
  AND U3993 ( .A(y[64]), .B(x[70]), .Z(n3934) );
  XOR U3994 ( .A(n3935), .B(n3934), .Z(n3932) );
  XNOR U3995 ( .A(n3933), .B(n3932), .Z(n3910) );
  XNOR U3996 ( .A(n3908), .B(n3909), .Z(n3906) );
  XNOR U3997 ( .A(n3907), .B(n3906), .Z(n3904) );
  XNOR U3998 ( .A(n3905), .B(n3904), .Z(n4045) );
  NAND U3999 ( .A(n3852), .B(n3851), .Z(n3856) );
  NANDN U4000 ( .A(n3854), .B(n3853), .Z(n3855) );
  NAND U4001 ( .A(n3856), .B(n3855), .Z(n4046) );
  XOR U4002 ( .A(n4047), .B(n4046), .Z(n4044) );
  XNOR U4003 ( .A(n4045), .B(n4044), .Z(n4059) );
  NAND U4004 ( .A(n3858), .B(n3857), .Z(n3862) );
  NAND U4005 ( .A(n3860), .B(n3859), .Z(n3861) );
  NAND U4006 ( .A(n3862), .B(n3861), .Z(n4061) );
  AND U4007 ( .A(x[58]), .B(y[44]), .Z(n3871) );
  NAND U4008 ( .A(x[57]), .B(y[45]), .Z(n3870) );
  XNOR U4009 ( .A(n3871), .B(n3870), .Z(n3993) );
  AND U4010 ( .A(y[20]), .B(x[50]), .Z(n3992) );
  XNOR U4011 ( .A(n3993), .B(n3992), .Z(n3921) );
  IV U4012 ( .A(n3872), .Z(n3874) );
  NAND U4013 ( .A(n3874), .B(n3873), .Z(n3878) );
  NAND U4014 ( .A(n3876), .B(n3875), .Z(n3877) );
  AND U4015 ( .A(n3878), .B(n3877), .Z(n3920) );
  XOR U4016 ( .A(n3919), .B(n3918), .Z(n4040) );
  XOR U4017 ( .A(n4041), .B(n4040), .Z(n4039) );
  AND U4018 ( .A(x[52]), .B(y[18]), .Z(n3880) );
  NAND U4019 ( .A(x[51]), .B(y[19]), .Z(n3879) );
  XNOR U4020 ( .A(n3880), .B(n3879), .Z(n3987) );
  AND U4021 ( .A(y[42]), .B(x[60]), .Z(n3986) );
  XNOR U4022 ( .A(n3987), .B(n3986), .Z(n3915) );
  AND U4023 ( .A(y[66]), .B(x[68]), .Z(n3884) );
  AND U4024 ( .A(n3885), .B(n3884), .Z(n3941) );
  AND U4025 ( .A(y[68]), .B(x[66]), .Z(n3940) );
  XOR U4026 ( .A(n3941), .B(n3940), .Z(n3938) );
  XOR U4027 ( .A(n3939), .B(n3938), .Z(n3913) );
  XNOR U4028 ( .A(n3912), .B(n3913), .Z(n4038) );
  XNOR U4029 ( .A(n4039), .B(n4038), .Z(n4060) );
  XOR U4030 ( .A(n4061), .B(n4060), .Z(n4058) );
  XNOR U4031 ( .A(n4059), .B(n4058), .Z(n4065) );
  NAND U4032 ( .A(n3887), .B(n3886), .Z(n3891) );
  NAND U4033 ( .A(n3889), .B(n3888), .Z(n3890) );
  NAND U4034 ( .A(n3891), .B(n3890), .Z(n4067) );
  NAND U4035 ( .A(n3893), .B(n3892), .Z(n3897) );
  NAND U4036 ( .A(n3895), .B(n3894), .Z(n3896) );
  NAND U4037 ( .A(n3897), .B(n3896), .Z(n4066) );
  NAND U4038 ( .A(n3899), .B(n3898), .Z(n3903) );
  NAND U4039 ( .A(n3901), .B(n3900), .Z(n3902) );
  AND U4040 ( .A(n3903), .B(n3902), .Z(n4055) );
  XOR U4041 ( .A(n4054), .B(n4055), .Z(n4052) );
  XOR U4042 ( .A(n4053), .B(n4052), .Z(o[70]) );
  NANDN U4043 ( .A(n3913), .B(n3912), .Z(n3917) );
  NAND U4044 ( .A(n3915), .B(n3914), .Z(n3916) );
  AND U4045 ( .A(n3917), .B(n3916), .Z(n4037) );
  NAND U4046 ( .A(n3919), .B(n3918), .Z(n3923) );
  NAND U4047 ( .A(n3921), .B(n3920), .Z(n3922) );
  AND U4048 ( .A(n3923), .B(n3922), .Z(n3931) );
  NANDN U4049 ( .A(n3925), .B(n3924), .Z(n3929) );
  NAND U4050 ( .A(n3927), .B(n3926), .Z(n3928) );
  NAND U4051 ( .A(n3929), .B(n3928), .Z(n3930) );
  XNOR U4052 ( .A(n3931), .B(n3930), .Z(n4035) );
  NAND U4053 ( .A(n3933), .B(n3932), .Z(n3937) );
  NAND U4054 ( .A(n3935), .B(n3934), .Z(n3936) );
  AND U4055 ( .A(n3937), .B(n3936), .Z(n4033) );
  NAND U4056 ( .A(n3939), .B(n3938), .Z(n3943) );
  NAND U4057 ( .A(n3941), .B(n3940), .Z(n3942) );
  AND U4058 ( .A(n3943), .B(n3942), .Z(n3972) );
  AND U4059 ( .A(x[64]), .B(y[71]), .Z(n3945) );
  NAND U4060 ( .A(x[59]), .B(y[44]), .Z(n3944) );
  XNOR U4061 ( .A(n3945), .B(n3944), .Z(n3952) );
  AND U4062 ( .A(x[51]), .B(y[20]), .Z(n3950) );
  AND U4063 ( .A(y[19]), .B(x[52]), .Z(n3988) );
  AND U4064 ( .A(x[49]), .B(y[22]), .Z(n3947) );
  NAND U4065 ( .A(x[60]), .B(y[43]), .Z(n3946) );
  XNOR U4066 ( .A(n3947), .B(n3946), .Z(n3948) );
  XNOR U4067 ( .A(n3988), .B(n3948), .Z(n3949) );
  XNOR U4068 ( .A(n3950), .B(n3949), .Z(n3951) );
  XOR U4069 ( .A(n3952), .B(n3951), .Z(n3954) );
  AND U4070 ( .A(y[66]), .B(x[69]), .Z(n4004) );
  AND U4071 ( .A(y[45]), .B(x[58]), .Z(n3994) );
  XNOR U4072 ( .A(n4004), .B(n3994), .Z(n3953) );
  XNOR U4073 ( .A(n3954), .B(n3953), .Z(n3970) );
  AND U4074 ( .A(x[67]), .B(y[68]), .Z(n3956) );
  NAND U4075 ( .A(x[53]), .B(y[18]), .Z(n3955) );
  XNOR U4076 ( .A(n3956), .B(n3955), .Z(n3960) );
  AND U4077 ( .A(x[55]), .B(y[16]), .Z(n3958) );
  NAND U4078 ( .A(x[66]), .B(y[69]), .Z(n3957) );
  XNOR U4079 ( .A(n3958), .B(n3957), .Z(n3959) );
  XOR U4080 ( .A(n3960), .B(n3959), .Z(n3968) );
  AND U4081 ( .A(x[71]), .B(y[64]), .Z(n3962) );
  NAND U4082 ( .A(x[61]), .B(y[42]), .Z(n3961) );
  XNOR U4083 ( .A(n3962), .B(n3961), .Z(n3966) );
  AND U4084 ( .A(x[56]), .B(y[47]), .Z(n3964) );
  NAND U4085 ( .A(x[70]), .B(y[65]), .Z(n3963) );
  XNOR U4086 ( .A(n3964), .B(n3963), .Z(n3965) );
  XNOR U4087 ( .A(n3966), .B(n3965), .Z(n3967) );
  XNOR U4088 ( .A(n3968), .B(n3967), .Z(n3969) );
  XNOR U4089 ( .A(n3970), .B(n3969), .Z(n3971) );
  XNOR U4090 ( .A(n3972), .B(n3971), .Z(n4031) );
  NAND U4091 ( .A(n3974), .B(n3973), .Z(n3978) );
  NAND U4092 ( .A(n3976), .B(n3975), .Z(n3977) );
  AND U4093 ( .A(n3978), .B(n3977), .Z(n3985) );
  NAND U4094 ( .A(n3980), .B(n3979), .Z(n3983) );
  AND U4095 ( .A(y[17]), .B(x[54]), .Z(n4022) );
  NAND U4096 ( .A(n3981), .B(n4022), .Z(n3982) );
  NAND U4097 ( .A(n3983), .B(n3982), .Z(n3984) );
  XNOR U4098 ( .A(n3985), .B(n3984), .Z(n4001) );
  NAND U4099 ( .A(n3987), .B(n3986), .Z(n3991) );
  NAND U4100 ( .A(n3989), .B(n3988), .Z(n3990) );
  AND U4101 ( .A(n3991), .B(n3990), .Z(n3999) );
  NAND U4102 ( .A(n3993), .B(n3992), .Z(n3997) );
  NAND U4103 ( .A(n3995), .B(n3994), .Z(n3996) );
  NAND U4104 ( .A(n3997), .B(n3996), .Z(n3998) );
  XNOR U4105 ( .A(n3999), .B(n3998), .Z(n4000) );
  XOR U4106 ( .A(n4001), .B(n4000), .Z(n4029) );
  AND U4107 ( .A(x[65]), .B(y[70]), .Z(n4003) );
  NAND U4108 ( .A(x[62]), .B(y[41]), .Z(n4002) );
  XNOR U4109 ( .A(n4003), .B(n4002), .Z(n4027) );
  AND U4110 ( .A(n4005), .B(n4004), .Z(n4021) );
  NAND U4111 ( .A(n4007), .B(n4006), .Z(n4011) );
  NAND U4112 ( .A(n4009), .B(n4008), .Z(n4010) );
  AND U4113 ( .A(n4011), .B(n4010), .Z(n4019) );
  AND U4114 ( .A(x[48]), .B(y[23]), .Z(n4013) );
  NAND U4115 ( .A(x[57]), .B(y[46]), .Z(n4012) );
  XNOR U4116 ( .A(n4013), .B(n4012), .Z(n4017) );
  AND U4117 ( .A(x[50]), .B(y[21]), .Z(n4015) );
  NAND U4118 ( .A(x[63]), .B(y[40]), .Z(n4014) );
  XNOR U4119 ( .A(n4015), .B(n4014), .Z(n4016) );
  XNOR U4120 ( .A(n4017), .B(n4016), .Z(n4018) );
  XNOR U4121 ( .A(n4019), .B(n4018), .Z(n4020) );
  XOR U4122 ( .A(n4021), .B(n4020), .Z(n4025) );
  XNOR U4123 ( .A(n4023), .B(n4022), .Z(n4024) );
  XNOR U4124 ( .A(n4025), .B(n4024), .Z(n4026) );
  XNOR U4125 ( .A(n4027), .B(n4026), .Z(n4028) );
  XNOR U4126 ( .A(n4029), .B(n4028), .Z(n4030) );
  XNOR U4127 ( .A(n4031), .B(n4030), .Z(n4032) );
  XNOR U4128 ( .A(n4033), .B(n4032), .Z(n4034) );
  XNOR U4129 ( .A(n4035), .B(n4034), .Z(n4036) );
  NAND U4130 ( .A(n4039), .B(n4038), .Z(n4043) );
  NAND U4131 ( .A(n4041), .B(n4040), .Z(n4042) );
  AND U4132 ( .A(n4043), .B(n4042), .Z(n4051) );
  NANDN U4133 ( .A(n4045), .B(n4044), .Z(n4049) );
  NAND U4134 ( .A(n4047), .B(n4046), .Z(n4048) );
  NAND U4135 ( .A(n4049), .B(n4048), .Z(n4050) );
  NAND U4136 ( .A(n4053), .B(n4052), .Z(n4057) );
  NAND U4137 ( .A(n4055), .B(n4054), .Z(n4056) );
  NAND U4138 ( .A(n4059), .B(n4058), .Z(n4063) );
  NAND U4139 ( .A(n4061), .B(n4060), .Z(n4062) );
endmodule

