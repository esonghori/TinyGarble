
module matrixMult_N_M_1_N5_M32 ( clk, rst, x, y, o );
  input [159:0] x;
  input [799:0] y;
  output [159:0] o;
  input clk, rst;
  wire   N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N161, N162, N163, N164, N165, N166, N167, N168, N169, N170,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N225, N226, N227, N228, N229, N230, N231, N232, N233, N234, N235,
         N236, N237, N238, N239, N240, N241, N242, N243, N244, N245, N246,
         N247, N248, N249, N250, N251, N252, N253, N254, N255, N256, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201,
         n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212,
         n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223,
         n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278,
         n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085;

  DFF \oi_reg[0][31]  ( .D(N64), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \oi_reg[0][30]  ( .D(N63), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \oi_reg[0][29]  ( .D(N62), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \oi_reg[0][28]  ( .D(N61), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \oi_reg[0][27]  ( .D(N60), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \oi_reg[0][26]  ( .D(N59), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \oi_reg[0][25]  ( .D(N58), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \oi_reg[0][24]  ( .D(N57), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \oi_reg[0][23]  ( .D(N56), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \oi_reg[0][22]  ( .D(N55), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \oi_reg[0][21]  ( .D(N54), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \oi_reg[0][20]  ( .D(N53), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \oi_reg[0][19]  ( .D(N52), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \oi_reg[0][18]  ( .D(N51), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \oi_reg[0][17]  ( .D(N50), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \oi_reg[0][16]  ( .D(N49), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \oi_reg[0][15]  ( .D(N48), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \oi_reg[0][14]  ( .D(N47), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \oi_reg[0][13]  ( .D(N46), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \oi_reg[0][12]  ( .D(N45), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \oi_reg[0][11]  ( .D(N44), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \oi_reg[0][10]  ( .D(N43), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \oi_reg[0][9]  ( .D(N42), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \oi_reg[0][8]  ( .D(N41), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \oi_reg[0][7]  ( .D(N40), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \oi_reg[0][6]  ( .D(N39), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \oi_reg[0][5]  ( .D(N38), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \oi_reg[0][4]  ( .D(N37), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \oi_reg[0][3]  ( .D(N36), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \oi_reg[0][2]  ( .D(N35), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \oi_reg[0][1]  ( .D(N34), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \oi_reg[0][0]  ( .D(N33), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \oi_reg[1][31]  ( .D(N128), .CLK(clk), .RST(rst), .Q(o[63]) );
  DFF \oi_reg[1][30]  ( .D(N127), .CLK(clk), .RST(rst), .Q(o[62]) );
  DFF \oi_reg[1][29]  ( .D(N126), .CLK(clk), .RST(rst), .Q(o[61]) );
  DFF \oi_reg[1][28]  ( .D(N125), .CLK(clk), .RST(rst), .Q(o[60]) );
  DFF \oi_reg[1][27]  ( .D(N124), .CLK(clk), .RST(rst), .Q(o[59]) );
  DFF \oi_reg[1][26]  ( .D(N123), .CLK(clk), .RST(rst), .Q(o[58]) );
  DFF \oi_reg[1][25]  ( .D(N122), .CLK(clk), .RST(rst), .Q(o[57]) );
  DFF \oi_reg[1][24]  ( .D(N121), .CLK(clk), .RST(rst), .Q(o[56]) );
  DFF \oi_reg[1][23]  ( .D(N120), .CLK(clk), .RST(rst), .Q(o[55]) );
  DFF \oi_reg[1][22]  ( .D(N119), .CLK(clk), .RST(rst), .Q(o[54]) );
  DFF \oi_reg[1][21]  ( .D(N118), .CLK(clk), .RST(rst), .Q(o[53]) );
  DFF \oi_reg[1][20]  ( .D(N117), .CLK(clk), .RST(rst), .Q(o[52]) );
  DFF \oi_reg[1][19]  ( .D(N116), .CLK(clk), .RST(rst), .Q(o[51]) );
  DFF \oi_reg[1][18]  ( .D(N115), .CLK(clk), .RST(rst), .Q(o[50]) );
  DFF \oi_reg[1][17]  ( .D(N114), .CLK(clk), .RST(rst), .Q(o[49]) );
  DFF \oi_reg[1][16]  ( .D(N113), .CLK(clk), .RST(rst), .Q(o[48]) );
  DFF \oi_reg[1][15]  ( .D(N112), .CLK(clk), .RST(rst), .Q(o[47]) );
  DFF \oi_reg[1][14]  ( .D(N111), .CLK(clk), .RST(rst), .Q(o[46]) );
  DFF \oi_reg[1][13]  ( .D(N110), .CLK(clk), .RST(rst), .Q(o[45]) );
  DFF \oi_reg[1][12]  ( .D(N109), .CLK(clk), .RST(rst), .Q(o[44]) );
  DFF \oi_reg[1][11]  ( .D(N108), .CLK(clk), .RST(rst), .Q(o[43]) );
  DFF \oi_reg[1][10]  ( .D(N107), .CLK(clk), .RST(rst), .Q(o[42]) );
  DFF \oi_reg[1][9]  ( .D(N106), .CLK(clk), .RST(rst), .Q(o[41]) );
  DFF \oi_reg[1][8]  ( .D(N105), .CLK(clk), .RST(rst), .Q(o[40]) );
  DFF \oi_reg[1][7]  ( .D(N104), .CLK(clk), .RST(rst), .Q(o[39]) );
  DFF \oi_reg[1][6]  ( .D(N103), .CLK(clk), .RST(rst), .Q(o[38]) );
  DFF \oi_reg[1][5]  ( .D(N102), .CLK(clk), .RST(rst), .Q(o[37]) );
  DFF \oi_reg[1][4]  ( .D(N101), .CLK(clk), .RST(rst), .Q(o[36]) );
  DFF \oi_reg[1][3]  ( .D(N100), .CLK(clk), .RST(rst), .Q(o[35]) );
  DFF \oi_reg[1][2]  ( .D(N99), .CLK(clk), .RST(rst), .Q(o[34]) );
  DFF \oi_reg[1][1]  ( .D(N98), .CLK(clk), .RST(rst), .Q(o[33]) );
  DFF \oi_reg[1][0]  ( .D(N97), .CLK(clk), .RST(rst), .Q(o[32]) );
  DFF \oi_reg[2][31]  ( .D(N192), .CLK(clk), .RST(rst), .Q(o[95]) );
  DFF \oi_reg[2][30]  ( .D(N191), .CLK(clk), .RST(rst), .Q(o[94]) );
  DFF \oi_reg[2][29]  ( .D(N190), .CLK(clk), .RST(rst), .Q(o[93]) );
  DFF \oi_reg[2][28]  ( .D(N189), .CLK(clk), .RST(rst), .Q(o[92]) );
  DFF \oi_reg[2][27]  ( .D(N188), .CLK(clk), .RST(rst), .Q(o[91]) );
  DFF \oi_reg[2][26]  ( .D(N187), .CLK(clk), .RST(rst), .Q(o[90]) );
  DFF \oi_reg[2][25]  ( .D(N186), .CLK(clk), .RST(rst), .Q(o[89]) );
  DFF \oi_reg[2][24]  ( .D(N185), .CLK(clk), .RST(rst), .Q(o[88]) );
  DFF \oi_reg[2][23]  ( .D(N184), .CLK(clk), .RST(rst), .Q(o[87]) );
  DFF \oi_reg[2][22]  ( .D(N183), .CLK(clk), .RST(rst), .Q(o[86]) );
  DFF \oi_reg[2][21]  ( .D(N182), .CLK(clk), .RST(rst), .Q(o[85]) );
  DFF \oi_reg[2][20]  ( .D(N181), .CLK(clk), .RST(rst), .Q(o[84]) );
  DFF \oi_reg[2][19]  ( .D(N180), .CLK(clk), .RST(rst), .Q(o[83]) );
  DFF \oi_reg[2][18]  ( .D(N179), .CLK(clk), .RST(rst), .Q(o[82]) );
  DFF \oi_reg[2][17]  ( .D(N178), .CLK(clk), .RST(rst), .Q(o[81]) );
  DFF \oi_reg[2][16]  ( .D(N177), .CLK(clk), .RST(rst), .Q(o[80]) );
  DFF \oi_reg[2][15]  ( .D(N176), .CLK(clk), .RST(rst), .Q(o[79]) );
  DFF \oi_reg[2][14]  ( .D(N175), .CLK(clk), .RST(rst), .Q(o[78]) );
  DFF \oi_reg[2][13]  ( .D(N174), .CLK(clk), .RST(rst), .Q(o[77]) );
  DFF \oi_reg[2][12]  ( .D(N173), .CLK(clk), .RST(rst), .Q(o[76]) );
  DFF \oi_reg[2][11]  ( .D(N172), .CLK(clk), .RST(rst), .Q(o[75]) );
  DFF \oi_reg[2][10]  ( .D(N171), .CLK(clk), .RST(rst), .Q(o[74]) );
  DFF \oi_reg[2][9]  ( .D(N170), .CLK(clk), .RST(rst), .Q(o[73]) );
  DFF \oi_reg[2][8]  ( .D(N169), .CLK(clk), .RST(rst), .Q(o[72]) );
  DFF \oi_reg[2][7]  ( .D(N168), .CLK(clk), .RST(rst), .Q(o[71]) );
  DFF \oi_reg[2][6]  ( .D(N167), .CLK(clk), .RST(rst), .Q(o[70]) );
  DFF \oi_reg[2][5]  ( .D(N166), .CLK(clk), .RST(rst), .Q(o[69]) );
  DFF \oi_reg[2][4]  ( .D(N165), .CLK(clk), .RST(rst), .Q(o[68]) );
  DFF \oi_reg[2][3]  ( .D(N164), .CLK(clk), .RST(rst), .Q(o[67]) );
  DFF \oi_reg[2][2]  ( .D(N163), .CLK(clk), .RST(rst), .Q(o[66]) );
  DFF \oi_reg[2][1]  ( .D(N162), .CLK(clk), .RST(rst), .Q(o[65]) );
  DFF \oi_reg[2][0]  ( .D(N161), .CLK(clk), .RST(rst), .Q(o[64]) );
  DFF \oi_reg[3][31]  ( .D(N256), .CLK(clk), .RST(rst), .Q(o[127]) );
  DFF \oi_reg[3][30]  ( .D(N255), .CLK(clk), .RST(rst), .Q(o[126]) );
  DFF \oi_reg[3][29]  ( .D(N254), .CLK(clk), .RST(rst), .Q(o[125]) );
  DFF \oi_reg[3][28]  ( .D(N253), .CLK(clk), .RST(rst), .Q(o[124]) );
  DFF \oi_reg[3][27]  ( .D(N252), .CLK(clk), .RST(rst), .Q(o[123]) );
  DFF \oi_reg[3][26]  ( .D(N251), .CLK(clk), .RST(rst), .Q(o[122]) );
  DFF \oi_reg[3][25]  ( .D(N250), .CLK(clk), .RST(rst), .Q(o[121]) );
  DFF \oi_reg[3][24]  ( .D(N249), .CLK(clk), .RST(rst), .Q(o[120]) );
  DFF \oi_reg[3][23]  ( .D(N248), .CLK(clk), .RST(rst), .Q(o[119]) );
  DFF \oi_reg[3][22]  ( .D(N247), .CLK(clk), .RST(rst), .Q(o[118]) );
  DFF \oi_reg[3][21]  ( .D(N246), .CLK(clk), .RST(rst), .Q(o[117]) );
  DFF \oi_reg[3][20]  ( .D(N245), .CLK(clk), .RST(rst), .Q(o[116]) );
  DFF \oi_reg[3][19]  ( .D(N244), .CLK(clk), .RST(rst), .Q(o[115]) );
  DFF \oi_reg[3][18]  ( .D(N243), .CLK(clk), .RST(rst), .Q(o[114]) );
  DFF \oi_reg[3][17]  ( .D(N242), .CLK(clk), .RST(rst), .Q(o[113]) );
  DFF \oi_reg[3][16]  ( .D(N241), .CLK(clk), .RST(rst), .Q(o[112]) );
  DFF \oi_reg[3][15]  ( .D(N240), .CLK(clk), .RST(rst), .Q(o[111]) );
  DFF \oi_reg[3][14]  ( .D(N239), .CLK(clk), .RST(rst), .Q(o[110]) );
  DFF \oi_reg[3][13]  ( .D(N238), .CLK(clk), .RST(rst), .Q(o[109]) );
  DFF \oi_reg[3][12]  ( .D(N237), .CLK(clk), .RST(rst), .Q(o[108]) );
  DFF \oi_reg[3][11]  ( .D(N236), .CLK(clk), .RST(rst), .Q(o[107]) );
  DFF \oi_reg[3][10]  ( .D(N235), .CLK(clk), .RST(rst), .Q(o[106]) );
  DFF \oi_reg[3][9]  ( .D(N234), .CLK(clk), .RST(rst), .Q(o[105]) );
  DFF \oi_reg[3][8]  ( .D(N233), .CLK(clk), .RST(rst), .Q(o[104]) );
  DFF \oi_reg[3][7]  ( .D(N232), .CLK(clk), .RST(rst), .Q(o[103]) );
  DFF \oi_reg[3][6]  ( .D(N231), .CLK(clk), .RST(rst), .Q(o[102]) );
  DFF \oi_reg[3][5]  ( .D(N230), .CLK(clk), .RST(rst), .Q(o[101]) );
  DFF \oi_reg[3][4]  ( .D(N229), .CLK(clk), .RST(rst), .Q(o[100]) );
  DFF \oi_reg[3][3]  ( .D(N228), .CLK(clk), .RST(rst), .Q(o[99]) );
  DFF \oi_reg[3][2]  ( .D(N227), .CLK(clk), .RST(rst), .Q(o[98]) );
  DFF \oi_reg[3][1]  ( .D(N226), .CLK(clk), .RST(rst), .Q(o[97]) );
  DFF \oi_reg[3][0]  ( .D(N225), .CLK(clk), .RST(rst), .Q(o[96]) );
  DFF \oi_reg[4][31]  ( .D(N320), .CLK(clk), .RST(rst), .Q(o[159]) );
  DFF \oi_reg[4][30]  ( .D(N319), .CLK(clk), .RST(rst), .Q(o[158]) );
  DFF \oi_reg[4][29]  ( .D(N318), .CLK(clk), .RST(rst), .Q(o[157]) );
  DFF \oi_reg[4][28]  ( .D(N317), .CLK(clk), .RST(rst), .Q(o[156]) );
  DFF \oi_reg[4][27]  ( .D(N316), .CLK(clk), .RST(rst), .Q(o[155]) );
  DFF \oi_reg[4][26]  ( .D(N315), .CLK(clk), .RST(rst), .Q(o[154]) );
  DFF \oi_reg[4][25]  ( .D(N314), .CLK(clk), .RST(rst), .Q(o[153]) );
  DFF \oi_reg[4][24]  ( .D(N313), .CLK(clk), .RST(rst), .Q(o[152]) );
  DFF \oi_reg[4][23]  ( .D(N312), .CLK(clk), .RST(rst), .Q(o[151]) );
  DFF \oi_reg[4][22]  ( .D(N311), .CLK(clk), .RST(rst), .Q(o[150]) );
  DFF \oi_reg[4][21]  ( .D(N310), .CLK(clk), .RST(rst), .Q(o[149]) );
  DFF \oi_reg[4][20]  ( .D(N309), .CLK(clk), .RST(rst), .Q(o[148]) );
  DFF \oi_reg[4][19]  ( .D(N308), .CLK(clk), .RST(rst), .Q(o[147]) );
  DFF \oi_reg[4][18]  ( .D(N307), .CLK(clk), .RST(rst), .Q(o[146]) );
  DFF \oi_reg[4][17]  ( .D(N306), .CLK(clk), .RST(rst), .Q(o[145]) );
  DFF \oi_reg[4][16]  ( .D(N305), .CLK(clk), .RST(rst), .Q(o[144]) );
  DFF \oi_reg[4][15]  ( .D(N304), .CLK(clk), .RST(rst), .Q(o[143]) );
  DFF \oi_reg[4][14]  ( .D(N303), .CLK(clk), .RST(rst), .Q(o[142]) );
  DFF \oi_reg[4][13]  ( .D(N302), .CLK(clk), .RST(rst), .Q(o[141]) );
  DFF \oi_reg[4][12]  ( .D(N301), .CLK(clk), .RST(rst), .Q(o[140]) );
  DFF \oi_reg[4][11]  ( .D(N300), .CLK(clk), .RST(rst), .Q(o[139]) );
  DFF \oi_reg[4][10]  ( .D(N299), .CLK(clk), .RST(rst), .Q(o[138]) );
  DFF \oi_reg[4][9]  ( .D(N298), .CLK(clk), .RST(rst), .Q(o[137]) );
  DFF \oi_reg[4][8]  ( .D(N297), .CLK(clk), .RST(rst), .Q(o[136]) );
  DFF \oi_reg[4][7]  ( .D(N296), .CLK(clk), .RST(rst), .Q(o[135]) );
  DFF \oi_reg[4][6]  ( .D(N295), .CLK(clk), .RST(rst), .Q(o[134]) );
  DFF \oi_reg[4][5]  ( .D(N294), .CLK(clk), .RST(rst), .Q(o[133]) );
  DFF \oi_reg[4][4]  ( .D(N293), .CLK(clk), .RST(rst), .Q(o[132]) );
  DFF \oi_reg[4][3]  ( .D(N292), .CLK(clk), .RST(rst), .Q(o[131]) );
  DFF \oi_reg[4][2]  ( .D(N291), .CLK(clk), .RST(rst), .Q(o[130]) );
  DFF \oi_reg[4][1]  ( .D(N290), .CLK(clk), .RST(rst), .Q(o[129]) );
  DFF \oi_reg[4][0]  ( .D(N289), .CLK(clk), .RST(rst), .Q(o[128]) );
  NAND U3 ( .A(n13912), .B(n13911), .Z(n1) );
  NAND U4 ( .A(n13909), .B(n13910), .Z(n2) );
  NAND U5 ( .A(n1), .B(n2), .Z(n14046) );
  AND U6 ( .A(n10258), .B(n10257), .Z(n3) );
  AND U7 ( .A(n10660), .B(y[743]), .Z(n4) );
  NAND U8 ( .A(x[144]), .B(n4), .Z(n5) );
  NANDN U9 ( .A(n3), .B(n5), .Z(n10419) );
  NAND U10 ( .A(n4323), .B(n4322), .Z(n6) );
  NAND U11 ( .A(n4521), .B(n5090), .Z(n7) );
  NAND U12 ( .A(n6), .B(n7), .Z(n4427) );
  XNOR U13 ( .A(n12957), .B(n12956), .Z(n12958) );
  NAND U14 ( .A(n13491), .B(n13490), .Z(n8) );
  NAND U15 ( .A(n13488), .B(n13489), .Z(n9) );
  NAND U16 ( .A(n8), .B(n9), .Z(n13634) );
  NAND U17 ( .A(n13888), .B(n13887), .Z(n10) );
  NAND U18 ( .A(n13885), .B(n13886), .Z(n11) );
  NAND U19 ( .A(n10), .B(n11), .Z(n14010) );
  XOR U20 ( .A(n9013), .B(n9012), .Z(n9015) );
  NAND U21 ( .A(n4425), .B(n4424), .Z(n12) );
  NAND U22 ( .A(n4422), .B(n4423), .Z(n13) );
  AND U23 ( .A(n12), .B(n13), .Z(n4563) );
  NAND U24 ( .A(n5724), .B(n5723), .Z(n14) );
  NAND U25 ( .A(n5721), .B(n5722), .Z(n15) );
  NAND U26 ( .A(n14), .B(n15), .Z(n5837) );
  XNOR U27 ( .A(n2322), .B(n2321), .Z(n2323) );
  XNOR U28 ( .A(n14737), .B(n14736), .Z(n14738) );
  XNOR U29 ( .A(n11903), .B(n11902), .Z(n11794) );
  NAND U30 ( .A(n8967), .B(n8966), .Z(n16) );
  NAND U31 ( .A(n8965), .B(n9085), .Z(n17) );
  NAND U32 ( .A(n16), .B(n17), .Z(n9079) );
  NAND U33 ( .A(n5889), .B(n5888), .Z(n18) );
  NAND U34 ( .A(n5886), .B(n5887), .Z(n19) );
  NAND U35 ( .A(n18), .B(n19), .Z(n6006) );
  NAND U36 ( .A(n5757), .B(n5756), .Z(n20) );
  NAND U37 ( .A(n5754), .B(n5755), .Z(n21) );
  NAND U38 ( .A(n20), .B(n21), .Z(n5923) );
  NAND U39 ( .A(n6038), .B(n6037), .Z(n22) );
  NAND U40 ( .A(n6035), .B(n6036), .Z(n23) );
  NAND U41 ( .A(n22), .B(n23), .Z(n6126) );
  NAND U42 ( .A(n13648), .B(n13647), .Z(n24) );
  NAND U43 ( .A(n13645), .B(n13646), .Z(n25) );
  NAND U44 ( .A(n24), .B(n25), .Z(n13868) );
  NAND U45 ( .A(n5933), .B(n5932), .Z(n26) );
  NAND U46 ( .A(n5930), .B(n5931), .Z(n27) );
  NAND U47 ( .A(n26), .B(n27), .Z(n6051) );
  NAND U48 ( .A(n6302), .B(n6301), .Z(n28) );
  NAND U49 ( .A(n6299), .B(n6300), .Z(n29) );
  NAND U50 ( .A(n28), .B(n29), .Z(n6303) );
  XNOR U51 ( .A(n1093), .B(n1092), .Z(n1100) );
  XNOR U52 ( .A(n6097), .B(n6096), .Z(n6094) );
  NAND U53 ( .A(n3122), .B(n3121), .Z(n30) );
  NANDN U54 ( .A(n3120), .B(n3119), .Z(n31) );
  AND U55 ( .A(n30), .B(n31), .Z(n3274) );
  XNOR U56 ( .A(n8328), .B(o[89]), .Z(n8298) );
  NAND U57 ( .A(n13938), .B(n13939), .Z(n32) );
  NAND U58 ( .A(n13940), .B(n13941), .Z(n33) );
  NAND U59 ( .A(n32), .B(n33), .Z(n14032) );
  XNOR U60 ( .A(n8460), .B(n8461), .Z(n8485) );
  XNOR U61 ( .A(n1609), .B(n1608), .Z(n1652) );
  XNOR U62 ( .A(n1994), .B(n1993), .Z(n1970) );
  NAND U63 ( .A(n13469), .B(n13331), .Z(n34) );
  NANDN U64 ( .A(n13431), .B(n13330), .Z(n35) );
  NAND U65 ( .A(n34), .B(n35), .Z(n13437) );
  AND U66 ( .A(n13348), .B(n13347), .Z(n36) );
  AND U67 ( .A(n14214), .B(y[770]), .Z(n37) );
  NAND U68 ( .A(x[138]), .B(n37), .Z(n38) );
  NANDN U69 ( .A(n36), .B(n38), .Z(n13481) );
  NAND U70 ( .A(n13816), .B(n13815), .Z(n39) );
  NAND U71 ( .A(n13813), .B(n13814), .Z(n40) );
  NAND U72 ( .A(n39), .B(n40), .Z(n13886) );
  NAND U73 ( .A(n13804), .B(n13803), .Z(n41) );
  NAND U74 ( .A(n13801), .B(n13802), .Z(n42) );
  NAND U75 ( .A(n41), .B(n42), .Z(n13973) );
  NAND U76 ( .A(n13898), .B(n13897), .Z(n43) );
  NAND U77 ( .A(n13895), .B(n13896), .Z(n44) );
  AND U78 ( .A(n43), .B(n44), .Z(n14041) );
  XNOR U79 ( .A(n14229), .B(n14228), .Z(n14264) );
  NAND U80 ( .A(n14103), .B(n14102), .Z(n45) );
  NAND U81 ( .A(n14100), .B(n14101), .Z(n46) );
  NAND U82 ( .A(n45), .B(n46), .Z(n14186) );
  NAND U83 ( .A(n10302), .B(n10301), .Z(n47) );
  NAND U84 ( .A(n10299), .B(n10300), .Z(n48) );
  NAND U85 ( .A(n47), .B(n48), .Z(n10410) );
  OR U86 ( .A(n4319), .B(n4447), .Z(n49) );
  NAND U87 ( .A(n4320), .B(n4321), .Z(n50) );
  NAND U88 ( .A(n49), .B(n50), .Z(n4426) );
  XNOR U89 ( .A(n12959), .B(n12958), .Z(n12950) );
  XNOR U90 ( .A(n12987), .B(n12986), .Z(n13028) );
  XNOR U91 ( .A(n12965), .B(n12964), .Z(n12945) );
  XNOR U92 ( .A(n14123), .B(n14122), .Z(n14117) );
  XNOR U93 ( .A(n14530), .B(n14722), .Z(n14531) );
  NAND U94 ( .A(n10107), .B(n10106), .Z(n51) );
  NAND U95 ( .A(n10104), .B(n10105), .Z(n52) );
  NAND U96 ( .A(n51), .B(n52), .Z(n10218) );
  NAND U97 ( .A(n10200), .B(n10199), .Z(n53) );
  NANDN U98 ( .A(n11139), .B(n10267), .Z(n54) );
  NAND U99 ( .A(n53), .B(n54), .Z(n10315) );
  NAND U100 ( .A(n10422), .B(n10421), .Z(n55) );
  NAND U101 ( .A(n10419), .B(n10420), .Z(n56) );
  AND U102 ( .A(n55), .B(n56), .Z(n10556) );
  XNOR U103 ( .A(n11500), .B(n11499), .Z(n11565) );
  XNOR U104 ( .A(n6856), .B(n6855), .Z(n6859) );
  XNOR U105 ( .A(n7085), .B(n7084), .Z(n7086) );
  XNOR U106 ( .A(n7264), .B(n7263), .Z(n7314) );
  XNOR U107 ( .A(n8838), .B(n8837), .Z(n8734) );
  XNOR U108 ( .A(n8830), .B(n8829), .Z(n8831) );
  XNOR U109 ( .A(n4107), .B(n4106), .Z(n4056) );
  NAND U110 ( .A(n4421), .B(n4420), .Z(n57) );
  NAND U111 ( .A(n4418), .B(n4419), .Z(n58) );
  AND U112 ( .A(n57), .B(n58), .Z(n4564) );
  NAND U113 ( .A(n5874), .B(n5873), .Z(n59) );
  NAND U114 ( .A(n5872), .B(n6020), .Z(n60) );
  AND U115 ( .A(n59), .B(n60), .Z(n6075) );
  NAND U116 ( .A(n5843), .B(n5842), .Z(n61) );
  NAND U117 ( .A(n5840), .B(n5841), .Z(n62) );
  NAND U118 ( .A(n61), .B(n62), .Z(n6089) );
  NAND U119 ( .A(n5720), .B(n5719), .Z(n63) );
  NAND U120 ( .A(n5717), .B(n5718), .Z(n64) );
  NAND U121 ( .A(n63), .B(n64), .Z(n5836) );
  XOR U122 ( .A(n1769), .B(n1768), .Z(n1773) );
  XOR U123 ( .A(n1898), .B(n1897), .Z(n1902) );
  XNOR U124 ( .A(n2174), .B(n2173), .Z(n2178) );
  XNOR U125 ( .A(n2306), .B(n2305), .Z(n2324) );
  XNOR U126 ( .A(n14538), .B(n14537), .Z(n14599) );
  XNOR U127 ( .A(n14515), .B(n14514), .Z(n14605) );
  XNOR U128 ( .A(n9870), .B(n9869), .Z(n9871) );
  NAND U129 ( .A(n10225), .B(n10224), .Z(n65) );
  NAND U130 ( .A(n10222), .B(n10223), .Z(n66) );
  NAND U131 ( .A(n65), .B(n66), .Z(n10241) );
  NAND U132 ( .A(n10247), .B(n10246), .Z(n67) );
  NANDN U133 ( .A(n10245), .B(n10244), .Z(n68) );
  AND U134 ( .A(n67), .B(n68), .Z(n10443) );
  XOR U135 ( .A(n8725), .B(n8724), .Z(n8711) );
  XNOR U136 ( .A(n9242), .B(n9241), .Z(n9239) );
  XOR U137 ( .A(n5821), .B(n5820), .Z(n5807) );
  NAND U138 ( .A(n5753), .B(n5752), .Z(n69) );
  NAND U139 ( .A(n5750), .B(n5751), .Z(n70) );
  NAND U140 ( .A(n69), .B(n70), .Z(n5922) );
  NAND U141 ( .A(n6069), .B(n6068), .Z(n71) );
  NANDN U142 ( .A(n6071), .B(n6070), .Z(n72) );
  AND U143 ( .A(n71), .B(n72), .Z(n6301) );
  NAND U144 ( .A(n5859), .B(n5858), .Z(n73) );
  NAND U145 ( .A(n5856), .B(n5857), .Z(n74) );
  AND U146 ( .A(n73), .B(n74), .Z(n6058) );
  XNOR U147 ( .A(n1033), .B(n1032), .Z(n1034) );
  XNOR U148 ( .A(n2318), .B(n2317), .Z(n2198) );
  OR U149 ( .A(n13643), .B(n13644), .Z(n75) );
  NAND U150 ( .A(n13642), .B(n13641), .Z(n76) );
  AND U151 ( .A(n75), .B(n76), .Z(n13871) );
  NAND U152 ( .A(n14272), .B(n14271), .Z(n77) );
  NAND U153 ( .A(n14269), .B(n14270), .Z(n78) );
  NAND U154 ( .A(n77), .B(n78), .Z(n14283) );
  XOR U155 ( .A(n12208), .B(n12207), .Z(n79) );
  XNOR U156 ( .A(n12209), .B(n79), .Z(n12193) );
  XNOR U157 ( .A(n9268), .B(n9267), .Z(n9265) );
  XNOR U158 ( .A(n4806), .B(n4805), .Z(n4821) );
  NAND U159 ( .A(n5929), .B(n5928), .Z(n80) );
  NAND U160 ( .A(n5926), .B(n5927), .Z(n81) );
  NAND U161 ( .A(n80), .B(n81), .Z(n6050) );
  NAND U162 ( .A(n5982), .B(n5981), .Z(n82) );
  NANDN U163 ( .A(n5984), .B(n5983), .Z(n83) );
  AND U164 ( .A(n82), .B(n83), .Z(n6333) );
  NAND U165 ( .A(n6118), .B(n6119), .Z(n84) );
  NAND U166 ( .A(n6120), .B(n6121), .Z(n85) );
  AND U167 ( .A(n84), .B(n85), .Z(n86) );
  NANDN U168 ( .A(n6125), .B(n6124), .Z(n87) );
  NANDN U169 ( .A(n6123), .B(n6122), .Z(n88) );
  AND U170 ( .A(n87), .B(n88), .Z(n89) );
  NAND U171 ( .A(n6127), .B(n6126), .Z(n90) );
  NAND U172 ( .A(n6128), .B(n6129), .Z(n91) );
  AND U173 ( .A(n90), .B(n91), .Z(n92) );
  XOR U174 ( .A(n6259), .B(n6258), .Z(n93) );
  XNOR U175 ( .A(n6205), .B(n6204), .Z(n94) );
  XNOR U176 ( .A(n93), .B(n94), .Z(n95) );
  AND U177 ( .A(n6134), .B(n6133), .Z(n96) );
  XNOR U178 ( .A(n6290), .B(n95), .Z(n97) );
  XNOR U179 ( .A(n96), .B(n97), .Z(n98) );
  XOR U180 ( .A(n92), .B(n98), .Z(n99) );
  XNOR U181 ( .A(n86), .B(n89), .Z(n100) );
  XNOR U182 ( .A(n99), .B(n100), .Z(n6291) );
  XOR U183 ( .A(n1100), .B(n1099), .Z(n1102) );
  XNOR U184 ( .A(n3133), .B(n3132), .Z(n3123) );
  XNOR U185 ( .A(n15043), .B(n15042), .Z(n14786) );
  XNOR U186 ( .A(n11942), .B(n11941), .Z(n11939) );
  XNOR U187 ( .A(n6443), .B(n6442), .Z(n6448) );
  XNOR U188 ( .A(n9042), .B(n9041), .Z(n9039) );
  XNOR U189 ( .A(n3621), .B(n3620), .Z(n3626) );
  XOR U190 ( .A(n6365), .B(n6364), .Z(n6363) );
  XOR U191 ( .A(n3548), .B(n3549), .Z(n3550) );
  XNOR U192 ( .A(n13087), .B(n13086), .Z(n13101) );
  XNOR U193 ( .A(n11147), .B(n11146), .Z(n11152) );
  XNOR U194 ( .A(n8301), .B(n8300), .Z(n8311) );
  XNOR U195 ( .A(n8507), .B(n8506), .Z(n8508) );
  XNOR U196 ( .A(n1631), .B(n1630), .Z(n1646) );
  XNOR U197 ( .A(n1618), .B(n1617), .Z(n1653) );
  XNOR U198 ( .A(n1702), .B(n1701), .Z(n1683) );
  XNOR U199 ( .A(n1743), .B(n1742), .Z(n1744) );
  XNOR U200 ( .A(n1960), .B(n1959), .Z(n1971) );
  XNOR U201 ( .A(n1979), .B(n1978), .Z(n2016) );
  XNOR U202 ( .A(n2006), .B(n2005), .Z(n2026) );
  XNOR U203 ( .A(n2518), .B(n2517), .Z(n2523) );
  XNOR U204 ( .A(n12850), .B(n12849), .Z(n12822) );
  XNOR U205 ( .A(n13096), .B(n13095), .Z(n13145) );
  NAND U206 ( .A(n13424), .B(n13423), .Z(n101) );
  NAND U207 ( .A(n13422), .B(n14835), .Z(n102) );
  NAND U208 ( .A(n101), .B(n102), .Z(n13616) );
  NAND U209 ( .A(n13335), .B(n13334), .Z(n103) );
  NAND U210 ( .A(n13332), .B(n13333), .Z(n104) );
  NAND U211 ( .A(n103), .B(n104), .Z(n13435) );
  NAND U212 ( .A(n13313), .B(n13312), .Z(n105) );
  NAND U213 ( .A(n13311), .B(n14208), .Z(n106) );
  NAND U214 ( .A(n105), .B(n106), .Z(n13445) );
  NAND U215 ( .A(n13776), .B(n13775), .Z(n107) );
  NAND U216 ( .A(n13773), .B(n13774), .Z(n108) );
  NAND U217 ( .A(n107), .B(n108), .Z(n13889) );
  XNOR U218 ( .A(n14217), .B(n14216), .Z(n14198) );
  XNOR U219 ( .A(n14264), .B(n14263), .Z(n14265) );
  XNOR U220 ( .A(n10535), .B(n10534), .Z(n10489) );
  XNOR U221 ( .A(n11414), .B(n11413), .Z(n11415) );
  XNOR U222 ( .A(n7270), .B(n7269), .Z(n7275) );
  XNOR U223 ( .A(n8435), .B(n8434), .Z(n8471) );
  XNOR U224 ( .A(n8586), .B(n8585), .Z(n8587) );
  XNOR U225 ( .A(n4349), .B(n4348), .Z(n4350) );
  NAND U226 ( .A(n4327), .B(n4326), .Z(n109) );
  NAND U227 ( .A(n4324), .B(n4325), .Z(n110) );
  NAND U228 ( .A(n109), .B(n110), .Z(n4425) );
  XNOR U229 ( .A(n4667), .B(n4666), .Z(n4668) );
  NAND U230 ( .A(n4861), .B(n4860), .Z(n111) );
  NANDN U231 ( .A(n4863), .B(n4862), .Z(n112) );
  NAND U232 ( .A(n111), .B(n112), .Z(n4963) );
  XNOR U233 ( .A(n1710), .B(n1709), .Z(n1748) );
  XNOR U234 ( .A(n12675), .B(n12674), .Z(n12668) );
  XNOR U235 ( .A(n13060), .B(n13059), .Z(n13030) );
  XOR U236 ( .A(n13370), .B(n13369), .Z(n13364) );
  NAND U237 ( .A(n13432), .B(n13431), .Z(n113) );
  NANDN U238 ( .A(n13434), .B(n13433), .Z(n114) );
  NAND U239 ( .A(n113), .B(n114), .Z(n13612) );
  XOR U240 ( .A(n13637), .B(n13636), .Z(n13631) );
  XNOR U241 ( .A(n14121), .B(n14120), .Z(n14122) );
  NAND U242 ( .A(n13973), .B(n13972), .Z(n115) );
  NANDN U243 ( .A(n13975), .B(n13974), .Z(n116) );
  AND U244 ( .A(n115), .B(n116), .Z(n14118) );
  NAND U245 ( .A(n14045), .B(n14044), .Z(n117) );
  NAND U246 ( .A(n14042), .B(n14043), .Z(n118) );
  AND U247 ( .A(n117), .B(n118), .Z(n14144) );
  OR U248 ( .A(n14048), .B(n14049), .Z(n119) );
  NAND U249 ( .A(n14046), .B(n14047), .Z(n120) );
  NAND U250 ( .A(n119), .B(n120), .Z(n14190) );
  XNOR U251 ( .A(n14543), .B(n14542), .Z(n14544) );
  XNOR U252 ( .A(n9696), .B(n9695), .Z(n9699) );
  NAND U253 ( .A(n10103), .B(n10102), .Z(n121) );
  NAND U254 ( .A(n10100), .B(n10101), .Z(n122) );
  NAND U255 ( .A(n121), .B(n122), .Z(n10220) );
  NAND U256 ( .A(n10179), .B(n10178), .Z(n123) );
  NANDN U257 ( .A(n10181), .B(n10180), .Z(n124) );
  AND U258 ( .A(n123), .B(n124), .Z(n10303) );
  XNOR U259 ( .A(n10316), .B(n10315), .Z(n10318) );
  XNOR U260 ( .A(n10322), .B(n10321), .Z(n10324) );
  NAND U261 ( .A(n10412), .B(n10411), .Z(n125) );
  NAND U262 ( .A(n10409), .B(n10410), .Z(n126) );
  AND U263 ( .A(n125), .B(n126), .Z(n10559) );
  XNOR U264 ( .A(n11685), .B(n11684), .Z(n11687) );
  XNOR U265 ( .A(n11566), .B(n11565), .Z(n11568) );
  XNOR U266 ( .A(n6854), .B(n6853), .Z(n6855) );
  XNOR U267 ( .A(n7087), .B(n7086), .Z(n7078) );
  XNOR U268 ( .A(n7091), .B(n7090), .Z(n7092) );
  XNOR U269 ( .A(n8771), .B(n8770), .Z(n8819) );
  XNOR U270 ( .A(n8970), .B(n8969), .Z(n9000) );
  NAND U271 ( .A(n8615), .B(n8614), .Z(n127) );
  NANDN U272 ( .A(n8613), .B(n8612), .Z(n128) );
  NAND U273 ( .A(n127), .B(n128), .Z(n8740) );
  XOR U274 ( .A(n3930), .B(n3929), .Z(n3932) );
  XNOR U275 ( .A(n4004), .B(n4609), .Z(n3982) );
  XNOR U276 ( .A(n3972), .B(n3971), .Z(n3965) );
  XNOR U277 ( .A(n4065), .B(n4064), .Z(n4057) );
  XNOR U278 ( .A(n4510), .B(n4509), .Z(n4575) );
  NAND U279 ( .A(n4794), .B(n4793), .Z(n129) );
  NANDN U280 ( .A(n4796), .B(n4795), .Z(n130) );
  NAND U281 ( .A(n129), .B(n130), .Z(n4924) );
  NAND U282 ( .A(n4838), .B(n4837), .Z(n131) );
  NANDN U283 ( .A(n4836), .B(n4835), .Z(n132) );
  AND U284 ( .A(n131), .B(n132), .Z(n4960) );
  NAND U285 ( .A(n5711), .B(n5710), .Z(n133) );
  NAND U286 ( .A(n5708), .B(n5709), .Z(n134) );
  NAND U287 ( .A(n133), .B(n134), .Z(n5896) );
  XNOR U288 ( .A(n6000), .B(n5999), .Z(n6001) );
  XNOR U289 ( .A(n935), .B(n934), .Z(n961) );
  XNOR U290 ( .A(n985), .B(n984), .Z(n986) );
  XNOR U291 ( .A(n975), .B(n974), .Z(n978) );
  XNOR U292 ( .A(n1908), .B(n1907), .Z(n1909) );
  XNOR U293 ( .A(n2178), .B(n2177), .Z(n2180) );
  XOR U294 ( .A(n3025), .B(n3024), .Z(n3027) );
  XNOR U295 ( .A(n3439), .B(n3438), .Z(n3436) );
  NAND U296 ( .A(n12430), .B(n13232), .Z(n135) );
  NANDN U297 ( .A(n12432), .B(n12431), .Z(n136) );
  AND U298 ( .A(n135), .B(n136), .Z(n12461) );
  XNOR U299 ( .A(n13388), .B(n13387), .Z(n13391) );
  XNOR U300 ( .A(n14565), .B(n14564), .Z(n14586) );
  XNOR U301 ( .A(n14551), .B(n14550), .Z(n14598) );
  XNOR U302 ( .A(n14518), .B(n14519), .Z(n14604) );
  XNOR U303 ( .A(n14647), .B(n14646), .Z(n14653) );
  XNOR U304 ( .A(n14781), .B(n14780), .Z(n14743) );
  XOR U305 ( .A(n14766), .B(n14767), .Z(n137) );
  NANDN U306 ( .A(n14873), .B(n137), .Z(n138) );
  NAND U307 ( .A(n14766), .B(n14767), .Z(n139) );
  AND U308 ( .A(n138), .B(n139), .Z(n15008) );
  XNOR U309 ( .A(n11699), .B(n11698), .Z(n11732) );
  XNOR U310 ( .A(n6868), .B(n6867), .Z(n6861) );
  XNOR U311 ( .A(n7321), .B(n7320), .Z(n7322) );
  XNOR U312 ( .A(n8693), .B(n8692), .Z(n8550) );
  XNOR U313 ( .A(n8826), .B(n8825), .Z(n8729) );
  XOR U314 ( .A(n9080), .B(n9079), .Z(n9078) );
  XNOR U315 ( .A(n8888), .B(n8887), .Z(n8890) );
  XNOR U316 ( .A(n8882), .B(n8881), .Z(n8884) );
  XNOR U317 ( .A(n4112), .B(n4111), .Z(n4113) );
  XNOR U318 ( .A(n4491), .B(n4490), .Z(n4493) );
  NAND U319 ( .A(n5893), .B(n5892), .Z(n140) );
  NANDN U320 ( .A(n5891), .B(n5890), .Z(n141) );
  NAND U321 ( .A(n140), .B(n141), .Z(n5982) );
  NAND U322 ( .A(n6090), .B(n6089), .Z(n142) );
  NANDN U323 ( .A(n6092), .B(n6091), .Z(n143) );
  AND U324 ( .A(n142), .B(n143), .Z(n6294) );
  NAND U325 ( .A(n6041), .B(n6040), .Z(n144) );
  NAND U326 ( .A(n6039), .B(n6231), .Z(n145) );
  NAND U327 ( .A(n144), .B(n145), .Z(n6129) );
  NAND U328 ( .A(n5839), .B(n5838), .Z(n146) );
  NAND U329 ( .A(n5836), .B(n5837), .Z(n147) );
  AND U330 ( .A(n146), .B(n147), .Z(n6060) );
  XNOR U331 ( .A(n2312), .B(n2311), .Z(n2200) );
  XOR U332 ( .A(n2946), .B(n2945), .Z(n2932) );
  NAND U333 ( .A(n2867), .B(n2866), .Z(n148) );
  NANDN U334 ( .A(n2869), .B(n2868), .Z(n149) );
  NAND U335 ( .A(n148), .B(n149), .Z(n3044) );
  XNOR U336 ( .A(n3269), .B(n3268), .Z(n3184) );
  XNOR U337 ( .A(n3309), .B(n3308), .Z(n3306) );
  XNOR U338 ( .A(n3493), .B(n3492), .Z(n3490) );
  XNOR U339 ( .A(n12288), .B(n12287), .Z(n12292) );
  XOR U340 ( .A(n12947), .B(n12946), .Z(n12968) );
  XNOR U341 ( .A(n12981), .B(n12980), .Z(n13068) );
  XNOR U342 ( .A(n9358), .B(n9357), .Z(n9362) );
  XNOR U343 ( .A(n9523), .B(n9522), .Z(n9524) );
  XNOR U344 ( .A(n9872), .B(n9871), .Z(n9946) );
  XNOR U345 ( .A(n10563), .B(n10562), .Z(n10564) );
  XNOR U346 ( .A(n11885), .B(n11884), .Z(n11780) );
  XNOR U347 ( .A(n11946), .B(n11945), .Z(n12178) );
  NAND U348 ( .A(n6454), .B(n6453), .Z(n150) );
  XOR U349 ( .A(n6454), .B(n6453), .Z(n151) );
  NANDN U350 ( .A(n6514), .B(n151), .Z(n152) );
  NAND U351 ( .A(n150), .B(n152), .Z(n6490) );
  XOR U352 ( .A(n6596), .B(n6595), .Z(n6637) );
  XNOR U353 ( .A(n6932), .B(n6931), .Z(n7009) );
  XNOR U354 ( .A(n8985), .B(n8984), .Z(n8902) );
  XNOR U355 ( .A(n9048), .B(n9047), .Z(n9272) );
  NAND U356 ( .A(n3632), .B(n3631), .Z(n153) );
  XOR U357 ( .A(n3632), .B(n3631), .Z(n154) );
  NANDN U358 ( .A(n3692), .B(n154), .Z(n155) );
  NAND U359 ( .A(n153), .B(n155), .Z(n3668) );
  XOR U360 ( .A(n3836), .B(n3835), .Z(n3883) );
  XOR U361 ( .A(n4261), .B(n4260), .Z(n4282) );
  XNOR U362 ( .A(n5341), .B(n5340), .Z(n5342) );
  NAND U363 ( .A(n5925), .B(n5924), .Z(n156) );
  NAND U364 ( .A(n5922), .B(n5923), .Z(n157) );
  NAND U365 ( .A(n156), .B(n157), .Z(n6052) );
  NAND U366 ( .A(n5980), .B(n5979), .Z(n158) );
  NANDN U367 ( .A(n5978), .B(n5977), .Z(n159) );
  AND U368 ( .A(n158), .B(n159), .Z(n6346) );
  XOR U369 ( .A(n6336), .B(n6335), .Z(n6334) );
  NAND U370 ( .A(n5992), .B(n5991), .Z(n160) );
  NAND U371 ( .A(n5989), .B(n5990), .Z(n161) );
  NAND U372 ( .A(n160), .B(n161), .Z(n6106) );
  XNOR U373 ( .A(n1787), .B(n1786), .Z(n1790) );
  XNOR U374 ( .A(n3521), .B(n3520), .Z(n3518) );
  XNOR U375 ( .A(n3293), .B(n3292), .Z(n3290) );
  XNOR U376 ( .A(n3499), .B(n3498), .Z(n3497) );
  XNOR U377 ( .A(n3178), .B(n3177), .Z(n3137) );
  XNOR U378 ( .A(n12800), .B(n12799), .Z(n12806) );
  NAND U379 ( .A(n13746), .B(n13747), .Z(n162) );
  XOR U380 ( .A(n13746), .B(n13747), .Z(n163) );
  NANDN U381 ( .A(n13745), .B(n163), .Z(n164) );
  NAND U382 ( .A(n162), .B(n164), .Z(n13866) );
  NAND U383 ( .A(n13871), .B(n13870), .Z(n165) );
  NAND U384 ( .A(n13868), .B(n13869), .Z(n166) );
  AND U385 ( .A(n165), .B(n166), .Z(n13989) );
  NAND U386 ( .A(n14290), .B(n14291), .Z(n167) );
  XOR U387 ( .A(n14290), .B(n14291), .Z(n168) );
  NANDN U388 ( .A(n14289), .B(n168), .Z(n169) );
  NAND U389 ( .A(n167), .B(n169), .Z(n14450) );
  XNOR U390 ( .A(n14787), .B(n14786), .Z(n14784) );
  NAND U391 ( .A(n9866), .B(n9867), .Z(n170) );
  XOR U392 ( .A(n9866), .B(n9867), .Z(n171) );
  NANDN U393 ( .A(n9865), .B(n171), .Z(n172) );
  NAND U394 ( .A(n170), .B(n172), .Z(n9951) );
  NAND U395 ( .A(n10440), .B(n10441), .Z(n173) );
  XOR U396 ( .A(n10440), .B(n10441), .Z(n174) );
  NANDN U397 ( .A(n10439), .B(n174), .Z(n175) );
  NAND U398 ( .A(n173), .B(n175), .Z(n10569) );
  XNOR U399 ( .A(n12194), .B(n12193), .Z(n12221) );
  NAND U400 ( .A(n6448), .B(n6447), .Z(n176) );
  XOR U401 ( .A(n6448), .B(n6447), .Z(n177) );
  NANDN U402 ( .A(n6446), .B(n177), .Z(n178) );
  NAND U403 ( .A(n176), .B(n178), .Z(n6497) );
  XOR U404 ( .A(n9301), .B(n9302), .Z(n9303) );
  NAND U405 ( .A(n3626), .B(n3625), .Z(n179) );
  XOR U406 ( .A(n3626), .B(n3625), .Z(n180) );
  NANDN U407 ( .A(n3624), .B(n180), .Z(n181) );
  NAND U408 ( .A(n179), .B(n181), .Z(n3675) );
  XOR U409 ( .A(n4703), .B(n4702), .Z(n182) );
  NANDN U410 ( .A(n4704), .B(n182), .Z(n183) );
  NAND U411 ( .A(n4703), .B(n4702), .Z(n184) );
  AND U412 ( .A(n183), .B(n184), .Z(n4815) );
  NAND U413 ( .A(n4821), .B(n4820), .Z(n185) );
  NAND U414 ( .A(n4818), .B(n4819), .Z(n186) );
  AND U415 ( .A(n185), .B(n186), .Z(n4931) );
  XOR U416 ( .A(n5208), .B(n5207), .Z(n187) );
  NANDN U417 ( .A(n5206), .B(n187), .Z(n188) );
  NAND U418 ( .A(n5208), .B(n5207), .Z(n189) );
  AND U419 ( .A(n188), .B(n189), .Z(n5346) );
  NAND U420 ( .A(n5944), .B(n5945), .Z(n190) );
  XOR U421 ( .A(n5944), .B(n5945), .Z(n191) );
  NANDN U422 ( .A(n5946), .B(n191), .Z(n192) );
  NAND U423 ( .A(n190), .B(n192), .Z(n6356) );
  NAND U424 ( .A(n1107), .B(n1106), .Z(n193) );
  XOR U425 ( .A(n1107), .B(n1106), .Z(n194) );
  NANDN U426 ( .A(n1108), .B(n194), .Z(n195) );
  NAND U427 ( .A(n193), .B(n195), .Z(n1265) );
  XNOR U428 ( .A(n1919), .B(n1918), .Z(n1915) );
  NAND U429 ( .A(n2620), .B(n2621), .Z(n196) );
  XOR U430 ( .A(n2620), .B(n2621), .Z(n197) );
  NANDN U431 ( .A(n2619), .B(n197), .Z(n198) );
  NAND U432 ( .A(n196), .B(n198), .Z(n2777) );
  XNOR U433 ( .A(n3533), .B(n3532), .Z(n3531) );
  XNOR U434 ( .A(n11011), .B(n11010), .Z(n11074) );
  XNOR U435 ( .A(n1622), .B(n1621), .Z(n1624) );
  XNOR U436 ( .A(n2404), .B(n2403), .Z(n2405) );
  XNOR U437 ( .A(n13722), .B(n13721), .Z(n13688) );
  NAND U438 ( .A(n13683), .B(n13684), .Z(n199) );
  NAND U439 ( .A(n13685), .B(n13686), .Z(n200) );
  NAND U440 ( .A(n199), .B(n200), .Z(n13797) );
  NAND U441 ( .A(n13762), .B(n13761), .Z(n201) );
  NAND U442 ( .A(n13899), .B(n14165), .Z(n202) );
  AND U443 ( .A(n201), .B(n202), .Z(n13917) );
  NAND U444 ( .A(n13937), .B(n13936), .Z(n203) );
  NAND U445 ( .A(n13934), .B(n13935), .Z(n204) );
  NAND U446 ( .A(n203), .B(n204), .Z(n14033) );
  NAND U447 ( .A(n10269), .B(n10268), .Z(n205) );
  NANDN U448 ( .A(n11349), .B(n10267), .Z(n206) );
  AND U449 ( .A(n205), .B(n206), .Z(n10380) );
  XNOR U450 ( .A(n10356), .B(n10355), .Z(n10337) );
  XNOR U451 ( .A(n10674), .B(n10673), .Z(n10618) );
  XNOR U452 ( .A(n8465), .B(n8464), .Z(n8467) );
  XNOR U453 ( .A(n8495), .B(n8494), .Z(n8496) );
  XNOR U454 ( .A(n8415), .B(n8414), .Z(n8417) );
  XNOR U455 ( .A(n8502), .B(n8501), .Z(n8482) );
  XOR U456 ( .A(n8439), .B(n8438), .Z(n8441) );
  XNOR U457 ( .A(n1999), .B(n1998), .Z(n2001) );
  XOR U458 ( .A(n1956), .B(n1955), .Z(n1972) );
  XNOR U459 ( .A(n2015), .B(n2014), .Z(n2017) );
  XNOR U460 ( .A(n2522), .B(n2521), .Z(n2524) );
  XNOR U461 ( .A(n12859), .B(n13085), .Z(n12868) );
  XOR U462 ( .A(n12906), .B(n12905), .Z(n12940) );
  XNOR U463 ( .A(n12919), .B(n12918), .Z(n12921) );
  XNOR U464 ( .A(n12985), .B(n12984), .Z(n12986) );
  XNOR U465 ( .A(n13196), .B(n13195), .Z(n13197) );
  XNOR U466 ( .A(n13456), .B(n13455), .Z(n13434) );
  XNOR U467 ( .A(n13704), .B(n13703), .Z(n13665) );
  NAND U468 ( .A(n13928), .B(n13927), .Z(n207) );
  NANDN U469 ( .A(n14020), .B(n13926), .Z(n208) );
  NAND U470 ( .A(n207), .B(n208), .Z(n14042) );
  XOR U471 ( .A(n14233), .B(n14232), .Z(n14235) );
  XNOR U472 ( .A(n14878), .B(n14697), .Z(n14698) );
  XNOR U473 ( .A(n9553), .B(o[105]), .Z(n9543) );
  XNOR U474 ( .A(n9623), .B(n9622), .Z(n9597) );
  NAND U475 ( .A(n10209), .B(n10208), .Z(n209) );
  NANDN U476 ( .A(n10211), .B(n10210), .Z(n210) );
  AND U477 ( .A(n209), .B(n210), .Z(n10248) );
  AND U478 ( .A(n10256), .B(n10255), .Z(n211) );
  AND U479 ( .A(n10254), .B(y[749]), .Z(n212) );
  NAND U480 ( .A(x[134]), .B(n212), .Z(n213) );
  NANDN U481 ( .A(n211), .B(n213), .Z(n10421) );
  NAND U482 ( .A(n10298), .B(n10297), .Z(n214) );
  NAND U483 ( .A(n10295), .B(n10296), .Z(n215) );
  NAND U484 ( .A(n214), .B(n215), .Z(n10409) );
  XNOR U485 ( .A(n10541), .B(n10540), .Z(n10491) );
  XNOR U486 ( .A(n11404), .B(o[122]), .Z(n11358) );
  XNOR U487 ( .A(n11406), .B(n11405), .Z(n11407) );
  XNOR U488 ( .A(n11396), .B(n11395), .Z(n11344) );
  XNOR U489 ( .A(n11390), .B(n11389), .Z(n11320) );
  XNOR U490 ( .A(n11422), .B(n11421), .Z(n11369) );
  XNOR U491 ( .A(n6794), .B(n6793), .Z(n6787) );
  XNOR U492 ( .A(n6969), .B(n6968), .Z(n6941) );
  XNOR U493 ( .A(n7274), .B(n7273), .Z(n7276) );
  XNOR U494 ( .A(n7465), .B(n7464), .Z(n7446) );
  XNOR U495 ( .A(n8034), .B(n8033), .Z(n8035) );
  XNOR U496 ( .A(n8054), .B(n8053), .Z(n7991) );
  XNOR U497 ( .A(n8184), .B(n8183), .Z(n8186) );
  XNOR U498 ( .A(n8313), .B(n8312), .Z(n8284) );
  XNOR U499 ( .A(n8471), .B(n8470), .Z(n8472) );
  XNOR U500 ( .A(n8515), .B(n8514), .Z(n8517) );
  XNOR U501 ( .A(n8588), .B(n8587), .Z(n8575) );
  XOR U502 ( .A(n8625), .B(n8624), .Z(n8685) );
  XOR U503 ( .A(n8669), .B(n8668), .Z(n8679) );
  XNOR U504 ( .A(n4063), .B(n4062), .Z(n4064) );
  XNOR U505 ( .A(n4679), .B(n4678), .Z(n4681) );
  XNOR U506 ( .A(n6283), .B(n6042), .Z(n6043) );
  XNOR U507 ( .A(n952), .B(n951), .Z(n926) );
  XOR U508 ( .A(n1751), .B(n1750), .Z(n1761) );
  XNOR U509 ( .A(n1767), .B(n1766), .Z(n1768) );
  XNOR U510 ( .A(n1755), .B(n1754), .Z(n1757) );
  XNOR U511 ( .A(n1801), .B(n1800), .Z(n1803) );
  XNOR U512 ( .A(n2098), .B(n2097), .Z(n2085) );
  XNOR U513 ( .A(n2092), .B(n2091), .Z(n2165) );
  XNOR U514 ( .A(n2078), .B(n2077), .Z(n2079) );
  XNOR U515 ( .A(n2280), .B(n2279), .Z(n2281) );
  XNOR U516 ( .A(n2300), .B(n2299), .Z(n2237) );
  XNOR U517 ( .A(n2727), .B(n2726), .Z(n2728) );
  XNOR U518 ( .A(n2765), .B(n2764), .Z(n2766) );
  XOR U519 ( .A(n2903), .B(n2902), .Z(n2913) );
  XNOR U520 ( .A(n12685), .B(n12686), .Z(n12671) );
  XNOR U521 ( .A(n12823), .B(n12822), .Z(n12824) );
  XNOR U522 ( .A(n12951), .B(n12950), .Z(n12952) );
  XNOR U523 ( .A(n13264), .B(n13263), .Z(n13189) );
  XNOR U524 ( .A(n13368), .B(n13367), .Z(n13369) );
  NAND U525 ( .A(n13619), .B(n13618), .Z(n216) );
  NANDN U526 ( .A(n13617), .B(n13616), .Z(n217) );
  AND U527 ( .A(n216), .B(n217), .Z(n13651) );
  NAND U528 ( .A(n13438), .B(n13437), .Z(n218) );
  NAND U529 ( .A(n13435), .B(n13436), .Z(n219) );
  AND U530 ( .A(n218), .B(n219), .Z(n13614) );
  NAND U531 ( .A(n13487), .B(n13486), .Z(n220) );
  NAND U532 ( .A(n13484), .B(n13485), .Z(n221) );
  NAND U533 ( .A(n220), .B(n221), .Z(n13635) );
  NAND U534 ( .A(n13728), .B(n13727), .Z(n222) );
  NANDN U535 ( .A(n13726), .B(n13725), .Z(n223) );
  AND U536 ( .A(n222), .B(n223), .Z(n13856) );
  OR U537 ( .A(n14039), .B(n14038), .Z(n224) );
  NAND U538 ( .A(n14041), .B(n14040), .Z(n225) );
  NAND U539 ( .A(n224), .B(n225), .Z(n14145) );
  NAND U540 ( .A(n14157), .B(n14156), .Z(n226) );
  NAND U541 ( .A(n14154), .B(n14155), .Z(n227) );
  AND U542 ( .A(n226), .B(n227), .Z(n14433) );
  NAND U543 ( .A(n14187), .B(n14186), .Z(n228) );
  NAND U544 ( .A(n14184), .B(n14185), .Z(n229) );
  AND U545 ( .A(n228), .B(n229), .Z(n14306) );
  XNOR U546 ( .A(n14532), .B(n14531), .Z(n14562) );
  XNOR U547 ( .A(n14536), .B(n14535), .Z(n14537) );
  XNOR U548 ( .A(n14507), .B(n14506), .Z(n14508) );
  XNOR U549 ( .A(n9700), .B(n9699), .Z(n9701) );
  XNOR U550 ( .A(n9766), .B(n10349), .Z(n9744) );
  XNOR U551 ( .A(n9734), .B(n9733), .Z(n9727) );
  XNOR U552 ( .A(n10306), .B(n10305), .Z(n10244) );
  XNOR U553 ( .A(n11416), .B(n11415), .Z(n11378) );
  XNOR U554 ( .A(n11245), .B(n11244), .Z(n11249) );
  XNOR U555 ( .A(n11482), .B(n11481), .Z(n11554) );
  XNOR U556 ( .A(n7079), .B(n7078), .Z(n7080) );
  XNOR U557 ( .A(n7093), .B(n7092), .Z(n7073) );
  XNOR U558 ( .A(n9126), .B(n8968), .Z(n8969) );
  NAND U559 ( .A(n8605), .B(n8604), .Z(n230) );
  NAND U560 ( .A(n8603), .B(n8805), .Z(n231) );
  AND U561 ( .A(n230), .B(n231), .Z(n8743) );
  XNOR U562 ( .A(n8735), .B(n8734), .Z(n8737) );
  XNOR U563 ( .A(n8824), .B(n8823), .Z(n8825) );
  XNOR U564 ( .A(n8842), .B(n8841), .Z(n8843) );
  XNOR U565 ( .A(n3982), .B(n3983), .Z(n3968) );
  XNOR U566 ( .A(n4369), .B(n4368), .Z(n4338) );
  NAND U567 ( .A(n4412), .B(n4411), .Z(n232) );
  NAND U568 ( .A(n4409), .B(n4410), .Z(n233) );
  NAND U569 ( .A(n232), .B(n233), .Z(n4576) );
  XNOR U570 ( .A(n4560), .B(n4559), .Z(n4568) );
  XOR U571 ( .A(n4669), .B(n4668), .Z(n4592) );
  XNOR U572 ( .A(n5490), .B(n5489), .Z(n5493) );
  XNOR U573 ( .A(n5728), .B(n5727), .Z(n5785) );
  XOR U574 ( .A(n5769), .B(n5768), .Z(n5779) );
  NAND U575 ( .A(n5864), .B(n5865), .Z(n234) );
  NAND U576 ( .A(n5866), .B(n5867), .Z(n235) );
  NAND U577 ( .A(n234), .B(n235), .Z(n6069) );
  XNOR U578 ( .A(n6247), .B(n6246), .Z(n6244) );
  NAND U579 ( .A(n5761), .B(n5760), .Z(n236) );
  NAND U580 ( .A(n5758), .B(n5759), .Z(n237) );
  NAND U581 ( .A(n236), .B(n237), .Z(n5858) );
  XNOR U582 ( .A(n961), .B(n960), .Z(n962) );
  XNOR U583 ( .A(n979), .B(n978), .Z(n980) );
  XNOR U584 ( .A(n1051), .B(n1050), .Z(n1044) );
  XNOR U585 ( .A(n1441), .B(n1440), .Z(n1443) );
  XNOR U586 ( .A(n1592), .B(n1591), .Z(n1593) );
  XNOR U587 ( .A(n1837), .B(n1836), .Z(n1895) );
  XOR U588 ( .A(n1781), .B(n1780), .Z(n1785) );
  XNOR U589 ( .A(n1930), .B(n1929), .Z(n1931) );
  XNOR U590 ( .A(n2304), .B(n2303), .Z(n2305) );
  NAND U591 ( .A(n2834), .B(n2833), .Z(n238) );
  NAND U592 ( .A(n2831), .B(n2832), .Z(n239) );
  NAND U593 ( .A(n238), .B(n239), .Z(n3026) );
  NAND U594 ( .A(n12307), .B(n12306), .Z(n240) );
  XOR U595 ( .A(n12307), .B(n12306), .Z(n241) );
  NANDN U596 ( .A(n12380), .B(n241), .Z(n242) );
  NAND U597 ( .A(n240), .B(n242), .Z(n12328) );
  XNOR U598 ( .A(n12979), .B(n12978), .Z(n12980) );
  XNOR U599 ( .A(n13386), .B(n13385), .Z(n13387) );
  XNOR U600 ( .A(n13499), .B(n13498), .Z(n13501) );
  NAND U601 ( .A(n13633), .B(n13632), .Z(n243) );
  NANDN U602 ( .A(n13631), .B(n13630), .Z(n244) );
  NAND U603 ( .A(n243), .B(n244), .Z(n13641) );
  NAND U604 ( .A(n14013), .B(n14012), .Z(n245) );
  NAND U605 ( .A(n14010), .B(n14011), .Z(n246) );
  NAND U606 ( .A(n245), .B(n246), .Z(n14271) );
  NAND U607 ( .A(n14119), .B(n14118), .Z(n247) );
  NAND U608 ( .A(n14116), .B(n14117), .Z(n248) );
  AND U609 ( .A(n247), .B(n248), .Z(n14141) );
  XNOR U610 ( .A(n14293), .B(n14292), .Z(n14294) );
  XOR U611 ( .A(n14545), .B(n14544), .Z(n14587) );
  XOR U612 ( .A(n14761), .B(n14760), .Z(n14762) );
  XNOR U613 ( .A(n14743), .B(n14742), .Z(n14745) );
  XNOR U614 ( .A(n15009), .B(n15008), .Z(n15007) );
  XOR U615 ( .A(n9654), .B(n9653), .Z(n9683) );
  XNOR U616 ( .A(n9716), .B(n9715), .Z(n9717) );
  XNOR U617 ( .A(n9808), .B(n9807), .Z(n9795) );
  NAND U618 ( .A(n10221), .B(n10220), .Z(n249) );
  NAND U619 ( .A(n10218), .B(n10219), .Z(n250) );
  NAND U620 ( .A(n249), .B(n250), .Z(n10240) );
  XNOR U621 ( .A(n10430), .B(n10429), .Z(n10433) );
  XNOR U622 ( .A(n10704), .B(n10703), .Z(n10706) );
  XNOR U623 ( .A(n10698), .B(n10697), .Z(n10699) );
  XOR U624 ( .A(n11631), .B(n11630), .Z(n11729) );
  XNOR U625 ( .A(n11798), .B(n11797), .Z(n11799) );
  XNOR U626 ( .A(n11733), .B(n11732), .Z(n11734) );
  XOR U627 ( .A(n11596), .B(n11595), .Z(n11590) );
  XNOR U628 ( .A(n6529), .B(n6528), .Z(n6536) );
  XNOR U629 ( .A(n6930), .B(n6929), .Z(n6931) );
  XNOR U630 ( .A(n7111), .B(n7110), .Z(n7112) );
  XNOR U631 ( .A(n7550), .B(n7549), .Z(n7437) );
  XNOR U632 ( .A(n8558), .B(n8557), .Z(n8540) );
  XNOR U633 ( .A(n8832), .B(n8831), .Z(n8728) );
  XNOR U634 ( .A(n3828), .B(n3827), .Z(n3829) );
  XOR U635 ( .A(n4461), .B(n4460), .Z(n4383) );
  NAND U636 ( .A(n4574), .B(n4573), .Z(n251) );
  NAND U637 ( .A(n4571), .B(n4572), .Z(n252) );
  NAND U638 ( .A(n251), .B(n252), .Z(n4685) );
  NAND U639 ( .A(n4566), .B(n4565), .Z(n253) );
  NAND U640 ( .A(n4563), .B(n4564), .Z(n254) );
  AND U641 ( .A(n253), .B(n254), .Z(n4690) );
  XNOR U642 ( .A(n5071), .B(n5070), .Z(n5073) );
  XNOR U643 ( .A(n5793), .B(n5792), .Z(n5669) );
  XNOR U644 ( .A(n5917), .B(n5916), .Z(n5919) );
  NAND U645 ( .A(n5885), .B(n5884), .Z(n255) );
  NAND U646 ( .A(n5882), .B(n5883), .Z(n256) );
  NAND U647 ( .A(n255), .B(n256), .Z(n6005) );
  XNOR U648 ( .A(n5907), .B(n5906), .Z(n5824) );
  XNOR U649 ( .A(n6002), .B(n6001), .Z(n6028) );
  NAND U650 ( .A(n6084), .B(n6083), .Z(n257) );
  NAND U651 ( .A(n6081), .B(n6082), .Z(n258) );
  NAND U652 ( .A(n257), .B(n258), .Z(n6118) );
  NAND U653 ( .A(n5871), .B(n5870), .Z(n259) );
  NAND U654 ( .A(n5868), .B(n5869), .Z(n260) );
  NAND U655 ( .A(n259), .B(n260), .Z(n5988) );
  XNOR U656 ( .A(n987), .B(n986), .Z(n1017) );
  XNOR U657 ( .A(n2198), .B(n2197), .Z(n2199) );
  XNOR U658 ( .A(n2454), .B(n2453), .Z(n2455) );
  NAND U659 ( .A(n2863), .B(n2862), .Z(n261) );
  NANDN U660 ( .A(n2865), .B(n2864), .Z(n262) );
  AND U661 ( .A(n261), .B(n262), .Z(n3045) );
  XNOR U662 ( .A(n3151), .B(n3150), .Z(n3269) );
  XNOR U663 ( .A(n12322), .B(n12321), .Z(n12323) );
  XNOR U664 ( .A(n13067), .B(n13066), .Z(n13069) );
  XOR U665 ( .A(n14873), .B(n14766), .Z(n263) );
  XNOR U666 ( .A(n14767), .B(n263), .Z(n14682) );
  XNOR U667 ( .A(n14732), .B(n14731), .Z(n14626) );
  XNOR U668 ( .A(n14757), .B(n14756), .Z(n14647) );
  XNOR U669 ( .A(n14797), .B(n14796), .Z(n15033) );
  XNOR U670 ( .A(n9392), .B(n9391), .Z(n9393) );
  XOR U671 ( .A(n9776), .B(n9775), .Z(n9780) );
  XNOR U672 ( .A(n10040), .B(n10039), .Z(n10041) );
  NAND U673 ( .A(n10690), .B(n10689), .Z(n264) );
  NANDN U674 ( .A(n10692), .B(n10691), .Z(n265) );
  AND U675 ( .A(n264), .B(n265), .Z(n10819) );
  XNOR U676 ( .A(n11930), .B(n11929), .Z(n11889) );
  XOR U677 ( .A(n12202), .B(n12201), .Z(n12200) );
  XNOR U678 ( .A(n11954), .B(n11953), .Z(n11951) );
  NAND U679 ( .A(n6380), .B(n6379), .Z(n266) );
  NAND U680 ( .A(n6387), .B(n6378), .Z(n267) );
  AND U681 ( .A(n266), .B(n267), .Z(n6393) );
  XNOR U682 ( .A(n6701), .B(n6700), .Z(n6703) );
  XNOR U683 ( .A(n7008), .B(n7007), .Z(n7010) );
  XNOR U684 ( .A(n7323), .B(n7322), .Z(n7423) );
  XOR U685 ( .A(n9282), .B(n9281), .Z(n9275) );
  XNOR U686 ( .A(n9298), .B(n9297), .Z(n9296) );
  NAND U687 ( .A(n8867), .B(n8868), .Z(n268) );
  XOR U688 ( .A(n8867), .B(n8868), .Z(n269) );
  NANDN U689 ( .A(n8866), .B(n269), .Z(n270) );
  NAND U690 ( .A(n268), .B(n270), .Z(n9292) );
  NAND U691 ( .A(n3558), .B(n3557), .Z(n271) );
  NAND U692 ( .A(n3565), .B(n3556), .Z(n272) );
  AND U693 ( .A(n271), .B(n272), .Z(n3571) );
  XNOR U694 ( .A(n3890), .B(n3889), .Z(n3891) );
  XOR U695 ( .A(n4114), .B(n4113), .Z(n4196) );
  XNOR U696 ( .A(n4391), .B(n4390), .Z(n4478) );
  XNOR U697 ( .A(n4487), .B(n4486), .Z(n4581) );
  XNOR U698 ( .A(n4934), .B(n4933), .Z(n4936) );
  NAND U699 ( .A(n4956), .B(n4955), .Z(n273) );
  NANDN U700 ( .A(n4954), .B(n4953), .Z(n274) );
  AND U701 ( .A(n273), .B(n274), .Z(n5202) );
  NAND U702 ( .A(n6057), .B(n6056), .Z(n275) );
  NAND U703 ( .A(n6054), .B(n6055), .Z(n276) );
  NAND U704 ( .A(n275), .B(n276), .Z(n6329) );
  XOR U705 ( .A(n6312), .B(n6311), .Z(n6310) );
  XNOR U706 ( .A(n641), .B(n640), .Z(n652) );
  XNOR U707 ( .A(n1110), .B(n1109), .Z(n1111) );
  XNOR U708 ( .A(n1904), .B(n1903), .Z(n1919) );
  NAND U709 ( .A(n2958), .B(n2957), .Z(n277) );
  NANDN U710 ( .A(n2956), .B(n2955), .Z(n278) );
  AND U711 ( .A(n277), .B(n278), .Z(n3124) );
  XNOR U712 ( .A(n3539), .B(n3538), .Z(n3537) );
  XOR U713 ( .A(n3098), .B(n3099), .Z(n279) );
  NANDN U714 ( .A(n3100), .B(n279), .Z(n280) );
  NAND U715 ( .A(n3098), .B(n3099), .Z(n281) );
  AND U716 ( .A(n280), .B(n281), .Z(n3532) );
  NANDN U717 ( .A(n12297), .B(n12299), .Z(n282) );
  OR U718 ( .A(n12299), .B(n12300), .Z(n283) );
  NAND U719 ( .A(n12298), .B(n283), .Z(n284) );
  NAND U720 ( .A(n282), .B(n284), .Z(n12318) );
  XNOR U721 ( .A(n12513), .B(n12512), .Z(n12506) );
  XOR U722 ( .A(n12633), .B(n12634), .Z(n285) );
  NANDN U723 ( .A(n12635), .B(n285), .Z(n286) );
  NAND U724 ( .A(n12633), .B(n12634), .Z(n287) );
  AND U725 ( .A(n286), .B(n287), .Z(n12650) );
  NAND U726 ( .A(n12975), .B(n12976), .Z(n288) );
  XOR U727 ( .A(n12975), .B(n12976), .Z(n289) );
  NANDN U728 ( .A(n12974), .B(n289), .Z(n290) );
  NAND U729 ( .A(n288), .B(n290), .Z(n13063) );
  NAND U730 ( .A(n13531), .B(n13532), .Z(n291) );
  XOR U731 ( .A(n13531), .B(n13532), .Z(n292) );
  NANDN U732 ( .A(n13530), .B(n292), .Z(n293) );
  NAND U733 ( .A(n291), .B(n293), .Z(n13746) );
  XOR U734 ( .A(n13989), .B(n13988), .Z(n294) );
  NANDN U735 ( .A(n13990), .B(n294), .Z(n295) );
  NAND U736 ( .A(n13989), .B(n13988), .Z(n296) );
  AND U737 ( .A(n295), .B(n296), .Z(n14127) );
  XOR U738 ( .A(n14451), .B(n14450), .Z(n297) );
  NANDN U739 ( .A(n14452), .B(n297), .Z(n298) );
  NAND U740 ( .A(n14451), .B(n14450), .Z(n299) );
  AND U741 ( .A(n298), .B(n299), .Z(n14612) );
  XNOR U742 ( .A(n14793), .B(n14792), .Z(n14791) );
  NANDN U743 ( .A(n9367), .B(n9369), .Z(n300) );
  OR U744 ( .A(n9369), .B(n9370), .Z(n301) );
  NAND U745 ( .A(n9368), .B(n301), .Z(n302) );
  NAND U746 ( .A(n300), .B(n302), .Z(n9388) );
  XNOR U747 ( .A(n9525), .B(n9524), .Z(n9521) );
  NAND U748 ( .A(n9951), .B(n9952), .Z(n303) );
  XOR U749 ( .A(n9951), .B(n9952), .Z(n304) );
  NANDN U750 ( .A(n9950), .B(n304), .Z(n305) );
  NAND U751 ( .A(n303), .B(n305), .Z(n10036) );
  NAND U752 ( .A(n10571), .B(n10568), .Z(n306) );
  NANDN U753 ( .A(n10571), .B(n10570), .Z(n307) );
  NANDN U754 ( .A(n10569), .B(n307), .Z(n308) );
  NAND U755 ( .A(n306), .B(n308), .Z(n10694) );
  NAND U756 ( .A(n11111), .B(n11112), .Z(n309) );
  XOR U757 ( .A(n11111), .B(n11112), .Z(n310) );
  NANDN U758 ( .A(n11110), .B(n310), .Z(n311) );
  NAND U759 ( .A(n309), .B(n311), .Z(n11254) );
  XOR U760 ( .A(n11579), .B(n11578), .Z(n312) );
  NANDN U761 ( .A(n11577), .B(n312), .Z(n313) );
  NAND U762 ( .A(n11579), .B(n11578), .Z(n314) );
  AND U763 ( .A(n313), .B(n314), .Z(n11744) );
  NANDN U764 ( .A(n12208), .B(n12207), .Z(n12212) );
  NAND U765 ( .A(n6497), .B(n6498), .Z(n315) );
  XOR U766 ( .A(n6497), .B(n6498), .Z(n316) );
  NANDN U767 ( .A(n6496), .B(n316), .Z(n317) );
  NAND U768 ( .A(n315), .B(n317), .Z(n6532) );
  NAND U769 ( .A(n6642), .B(n6643), .Z(n318) );
  XOR U770 ( .A(n6642), .B(n6643), .Z(n319) );
  NANDN U771 ( .A(n6641), .B(n319), .Z(n320) );
  NAND U772 ( .A(n318), .B(n320), .Z(n6697) );
  NAND U773 ( .A(n6920), .B(n6921), .Z(n321) );
  XOR U774 ( .A(n6920), .B(n6921), .Z(n322) );
  NANDN U775 ( .A(n6919), .B(n322), .Z(n323) );
  NAND U776 ( .A(n321), .B(n323), .Z(n7004) );
  XNOR U777 ( .A(n7677), .B(n7676), .Z(n7670) );
  XOR U778 ( .A(n8233), .B(n8234), .Z(n324) );
  NANDN U779 ( .A(n8235), .B(n324), .Z(n325) );
  NAND U780 ( .A(n8233), .B(n8234), .Z(n326) );
  AND U781 ( .A(n325), .B(n326), .Z(n8533) );
  NAND U782 ( .A(n9054), .B(n9053), .Z(n327) );
  NANDN U783 ( .A(n9056), .B(n9055), .Z(n328) );
  AND U784 ( .A(n327), .B(n328), .Z(n329) );
  AND U785 ( .A(n9264), .B(n9263), .Z(n330) );
  NAND U786 ( .A(n9258), .B(n9257), .Z(n331) );
  XNOR U787 ( .A(n330), .B(n331), .Z(n332) );
  AND U788 ( .A(n9062), .B(n9061), .Z(n333) );
  XNOR U789 ( .A(n9252), .B(n9251), .Z(n334) );
  XNOR U790 ( .A(n333), .B(n334), .Z(n335) );
  NAND U791 ( .A(n9266), .B(n9265), .Z(n336) );
  NANDN U792 ( .A(n9268), .B(n9267), .Z(n337) );
  AND U793 ( .A(n336), .B(n337), .Z(n338) );
  NAND U794 ( .A(n9272), .B(n9271), .Z(n339) );
  NANDN U795 ( .A(n9270), .B(n9269), .Z(n340) );
  AND U796 ( .A(n339), .B(n340), .Z(n341) );
  XOR U797 ( .A(n338), .B(n341), .Z(n342) );
  XNOR U798 ( .A(n332), .B(n335), .Z(n343) );
  XNOR U799 ( .A(n342), .B(n343), .Z(n344) );
  XNOR U800 ( .A(n329), .B(n344), .Z(n9273) );
  NAND U801 ( .A(n3675), .B(n3676), .Z(n345) );
  XOR U802 ( .A(n3675), .B(n3676), .Z(n346) );
  NANDN U803 ( .A(n3674), .B(n346), .Z(n347) );
  NAND U804 ( .A(n345), .B(n347), .Z(n3710) );
  NAND U805 ( .A(n3880), .B(n3881), .Z(n348) );
  XOR U806 ( .A(n3880), .B(n3881), .Z(n349) );
  NANDN U807 ( .A(n3879), .B(n349), .Z(n350) );
  NAND U808 ( .A(n348), .B(n350), .Z(n3895) );
  XOR U809 ( .A(n4373), .B(n4372), .Z(n351) );
  NANDN U810 ( .A(n4374), .B(n351), .Z(n352) );
  NAND U811 ( .A(n4373), .B(n4372), .Z(n353) );
  AND U812 ( .A(n352), .B(n353), .Z(n4472) );
  XOR U813 ( .A(n4815), .B(n4816), .Z(n354) );
  NANDN U814 ( .A(n4817), .B(n354), .Z(n355) );
  NAND U815 ( .A(n4815), .B(n4816), .Z(n356) );
  AND U816 ( .A(n355), .B(n356), .Z(n4930) );
  XOR U817 ( .A(n5357), .B(n5356), .Z(n357) );
  NANDN U818 ( .A(n5358), .B(n357), .Z(n358) );
  NAND U819 ( .A(n5357), .B(n5356), .Z(n359) );
  AND U820 ( .A(n358), .B(n359), .Z(n5649) );
  XOR U821 ( .A(n5940), .B(n5941), .Z(n360) );
  NANDN U822 ( .A(n5942), .B(n360), .Z(n361) );
  NAND U823 ( .A(n5940), .B(n5941), .Z(n362) );
  AND U824 ( .A(n361), .B(n362), .Z(n5944) );
  NAND U825 ( .A(n6051), .B(n6050), .Z(n363) );
  NANDN U826 ( .A(n6053), .B(n6052), .Z(n364) );
  AND U827 ( .A(n363), .B(n364), .Z(n6347) );
  XOR U828 ( .A(n1096), .B(n1097), .Z(n365) );
  NANDN U829 ( .A(n1098), .B(n365), .Z(n366) );
  NAND U830 ( .A(n1096), .B(n1097), .Z(n367) );
  AND U831 ( .A(n366), .B(n367), .Z(n1107) );
  XOR U832 ( .A(n1350), .B(n1351), .Z(n368) );
  NANDN U833 ( .A(n1352), .B(n368), .Z(n369) );
  NAND U834 ( .A(n1350), .B(n1351), .Z(n370) );
  AND U835 ( .A(n369), .B(n370), .Z(n1453) );
  NAND U836 ( .A(n1797), .B(n1798), .Z(n371) );
  XOR U837 ( .A(n1797), .B(n1798), .Z(n372) );
  NANDN U838 ( .A(n1796), .B(n372), .Z(n373) );
  NAND U839 ( .A(n371), .B(n373), .Z(n1913) );
  NAND U840 ( .A(n2777), .B(n2778), .Z(n374) );
  XOR U841 ( .A(n2777), .B(n2778), .Z(n375) );
  NANDN U842 ( .A(n2776), .B(n375), .Z(n376) );
  NAND U843 ( .A(n374), .B(n376), .Z(n2786) );
  NANDN U844 ( .A(n3291), .B(n3290), .Z(n377) );
  NANDN U845 ( .A(n3293), .B(n3292), .Z(n378) );
  AND U846 ( .A(n377), .B(n378), .Z(n379) );
  AND U847 ( .A(n3501), .B(n3500), .Z(n380) );
  NAND U848 ( .A(n3495), .B(n3494), .Z(n381) );
  XNOR U849 ( .A(n380), .B(n381), .Z(n382) );
  AND U850 ( .A(n3299), .B(n3298), .Z(n383) );
  XNOR U851 ( .A(n3489), .B(n3488), .Z(n384) );
  XNOR U852 ( .A(n383), .B(n384), .Z(n385) );
  NAND U853 ( .A(n3503), .B(n3502), .Z(n386) );
  NANDN U854 ( .A(n3505), .B(n3504), .Z(n387) );
  AND U855 ( .A(n386), .B(n387), .Z(n388) );
  NAND U856 ( .A(n3507), .B(n3506), .Z(n389) );
  NAND U857 ( .A(n3508), .B(n3509), .Z(n390) );
  AND U858 ( .A(n389), .B(n390), .Z(n391) );
  XOR U859 ( .A(n388), .B(n391), .Z(n392) );
  XNOR U860 ( .A(n382), .B(n385), .Z(n393) );
  XNOR U861 ( .A(n392), .B(n393), .Z(n394) );
  XNOR U862 ( .A(n379), .B(n394), .Z(n3510) );
  XNOR U863 ( .A(n11009), .B(n11008), .Z(n11010) );
  XNOR U864 ( .A(n8299), .B(n8298), .Z(n8300) );
  AND U865 ( .A(n13246), .B(o[146]), .Z(n13335) );
  AND U866 ( .A(n13719), .B(o[150]), .Z(n13776) );
  NAND U867 ( .A(n13808), .B(n13807), .Z(n395) );
  NAND U868 ( .A(n13805), .B(n13806), .Z(n396) );
  NAND U869 ( .A(n395), .B(n396), .Z(n13897) );
  NAND U870 ( .A(n13767), .B(n13766), .Z(n397) );
  NAND U871 ( .A(n13764), .B(n13765), .Z(n398) );
  NAND U872 ( .A(n397), .B(n398), .Z(n13911) );
  NAND U873 ( .A(n13945), .B(n13944), .Z(n399) );
  NAND U874 ( .A(n13942), .B(n13943), .Z(n400) );
  NAND U875 ( .A(n399), .B(n400), .Z(n14028) );
  NAND U876 ( .A(n13901), .B(n13900), .Z(n401) );
  NANDN U877 ( .A(n14878), .B(n13899), .Z(n402) );
  NAND U878 ( .A(n401), .B(n402), .Z(n14106) );
  XNOR U879 ( .A(n10196), .B(n10195), .Z(n10208) );
  XNOR U880 ( .A(n10351), .B(n10350), .Z(n10377) );
  XNOR U881 ( .A(n10401), .B(n10400), .Z(n10338) );
  XNOR U882 ( .A(n10618), .B(n10617), .Z(n10600) );
  XNOR U883 ( .A(n10998), .B(n10999), .Z(n11081) );
  XNOR U884 ( .A(n11151), .B(n11150), .Z(n11153) );
  XNOR U885 ( .A(n7183), .B(n7182), .Z(n7185) );
  XNOR U886 ( .A(n8149), .B(n8148), .Z(n8143) );
  XOR U887 ( .A(n8332), .B(n8331), .Z(n8310) );
  XOR U888 ( .A(n8360), .B(n8359), .Z(n8362) );
  XNOR U889 ( .A(n8354), .B(n8353), .Z(n8356) );
  XNOR U890 ( .A(n8421), .B(n8420), .Z(n8423) );
  XNOR U891 ( .A(n8490), .B(n8491), .Z(n8427) );
  NAND U892 ( .A(n4780), .B(n4779), .Z(n403) );
  NANDN U893 ( .A(n4778), .B(n4777), .Z(n404) );
  NAND U894 ( .A(n403), .B(n404), .Z(n4902) );
  XNOR U895 ( .A(n5060), .B(n5059), .Z(n5024) );
  XNOR U896 ( .A(n5042), .B(n5041), .Z(n4999) );
  XNOR U897 ( .A(n1527), .B(n1526), .Z(n1504) );
  XNOR U898 ( .A(n1827), .B(o[20]), .Z(n1818) );
  XNOR U899 ( .A(n1640), .B(n1639), .Z(n1599) );
  XNOR U900 ( .A(n1954), .B(n1953), .Z(n1955) );
  XNOR U901 ( .A(n2156), .B(n2155), .Z(n2120) );
  XNOR U902 ( .A(n2218), .B(n2217), .Z(n2255) );
  XNOR U903 ( .A(n2406), .B(n2405), .Z(n2346) );
  XNOR U904 ( .A(n2393), .B(n2394), .Z(n2370) );
  XNOR U905 ( .A(n2733), .B(n2732), .Z(n2734) );
  XNOR U906 ( .A(n12874), .B(n12873), .Z(n12876) );
  XNOR U907 ( .A(n12910), .B(n12909), .Z(n12939) );
  XNOR U908 ( .A(n12925), .B(n12924), .Z(n12926) );
  NAND U909 ( .A(n13627), .B(n13626), .Z(n405) );
  NANDN U910 ( .A(n13629), .B(n13628), .Z(n406) );
  NAND U911 ( .A(n405), .B(n406), .Z(n13649) );
  NAND U912 ( .A(n13689), .B(n13688), .Z(n407) );
  NANDN U913 ( .A(n13691), .B(n13690), .Z(n408) );
  AND U914 ( .A(n407), .B(n408), .Z(n13792) );
  NAND U915 ( .A(n13772), .B(n13771), .Z(n409) );
  NAND U916 ( .A(n13770), .B(n14021), .Z(n410) );
  AND U917 ( .A(n409), .B(n410), .Z(n13890) );
  NAND U918 ( .A(n13812), .B(n13811), .Z(n411) );
  NAND U919 ( .A(n13809), .B(n13810), .Z(n412) );
  NAND U920 ( .A(n411), .B(n412), .Z(n13885) );
  NAND U921 ( .A(n13780), .B(n13779), .Z(n413) );
  NAND U922 ( .A(n13777), .B(n13778), .Z(n414) );
  AND U923 ( .A(n413), .B(n414), .Z(n13961) );
  NAND U924 ( .A(n13800), .B(n13799), .Z(n415) );
  NANDN U925 ( .A(n13798), .B(n13797), .Z(n416) );
  NAND U926 ( .A(n415), .B(n416), .Z(n13974) );
  NAND U927 ( .A(n10079), .B(n10078), .Z(n417) );
  NANDN U928 ( .A(n10911), .B(n10267), .Z(n418) );
  NAND U929 ( .A(n417), .B(n418), .Z(n10188) );
  XNOR U930 ( .A(n10365), .B(n10364), .Z(n10371) );
  XNOR U931 ( .A(n10490), .B(n10489), .Z(n10492) );
  XNOR U932 ( .A(n10527), .B(n10526), .Z(n10529) );
  XNOR U933 ( .A(n10869), .B(n10868), .Z(n10937) );
  XNOR U934 ( .A(n11054), .B(n11053), .Z(n11040) );
  XNOR U935 ( .A(n11394), .B(n11393), .Z(n11395) );
  XNOR U936 ( .A(n11408), .B(n11407), .Z(n11296) );
  XNOR U937 ( .A(n11420), .B(n11419), .Z(n11421) );
  XOR U938 ( .A(n6805), .B(n6804), .Z(n6789) );
  XNOR U939 ( .A(n7123), .B(n7122), .Z(n7125) );
  XNOR U940 ( .A(n7497), .B(n7496), .Z(n7447) );
  XNOR U941 ( .A(n7473), .B(n7472), .Z(n7511) );
  XNOR U942 ( .A(n8048), .B(n8047), .Z(n8036) );
  XNOR U943 ( .A(n8042), .B(n8041), .Z(n7993) );
  XNOR U944 ( .A(n8509), .B(n8508), .Z(n8403) );
  XNOR U945 ( .A(n8497), .B(n8496), .Z(n8451) );
  XNOR U946 ( .A(n8410), .B(n8411), .Z(n8445) );
  XNOR U947 ( .A(n8568), .B(n8567), .Z(n8569) );
  XNOR U948 ( .A(n8623), .B(n8622), .Z(n8624) );
  XNOR U949 ( .A(n8629), .B(n8628), .Z(n8631) );
  XNOR U950 ( .A(n8617), .B(n8616), .Z(n8619) );
  XNOR U951 ( .A(n8574), .B(n8573), .Z(n8576) );
  XNOR U952 ( .A(n3928), .B(o[43]), .Z(n3909) );
  XNOR U953 ( .A(n4307), .B(n4306), .Z(n4344) );
  XNOR U954 ( .A(n4616), .B(n4615), .Z(n4597) );
  XNOR U955 ( .A(n4624), .B(n4623), .Z(n4660) );
  NAND U956 ( .A(n4637), .B(n4636), .Z(n419) );
  NANDN U957 ( .A(n4635), .B(n4634), .Z(n420) );
  AND U958 ( .A(n419), .B(n420), .Z(n4735) );
  NAND U959 ( .A(n4859), .B(n4858), .Z(n421) );
  NAND U960 ( .A(n4856), .B(n4857), .Z(n422) );
  AND U961 ( .A(n421), .B(n422), .Z(n4964) );
  XNOR U962 ( .A(n5293), .B(n5292), .Z(n5295) );
  XNOR U963 ( .A(n5402), .B(n5401), .Z(n5403) );
  XNOR U964 ( .A(n5604), .B(n5605), .Z(n5607) );
  AND U965 ( .A(n5621), .B(o[58]), .Z(n5724) );
  XNOR U966 ( .A(n1323), .B(n1322), .Z(n1302) );
  XNOR U967 ( .A(n1605), .B(n1604), .Z(n1677) );
  XNOR U968 ( .A(n1649), .B(n1648), .Z(n1672) );
  XNOR U969 ( .A(n1655), .B(n1654), .Z(n1665) );
  XOR U970 ( .A(n1745), .B(n1744), .Z(n1762) );
  XNOR U971 ( .A(n1686), .B(n1685), .Z(n1766) );
  XNOR U972 ( .A(n2127), .B(n2126), .Z(n2095) );
  XNOR U973 ( .A(n2084), .B(n2083), .Z(n2086) );
  XNOR U974 ( .A(n2160), .B(n2159), .Z(n2162) );
  XNOR U975 ( .A(n2294), .B(n2293), .Z(n2282) );
  XNOR U976 ( .A(n2288), .B(n2287), .Z(n2239) );
  XOR U977 ( .A(n12671), .B(n12670), .Z(n12665) );
  XNOR U978 ( .A(n12963), .B(n12962), .Z(n12964) );
  XNOR U979 ( .A(n13029), .B(n13028), .Z(n13031) );
  XOR U980 ( .A(n12953), .B(n12952), .Z(n12944) );
  XNOR U981 ( .A(n13262), .B(n13261), .Z(n13263) );
  XNOR U982 ( .A(n13274), .B(n13273), .Z(n13276) );
  XNOR U983 ( .A(n13280), .B(n13279), .Z(n13282) );
  XNOR U984 ( .A(n13268), .B(n13267), .Z(n13270) );
  XNOR U985 ( .A(n13198), .B(n13197), .Z(n13192) );
  XOR U986 ( .A(n13380), .B(n13379), .Z(n13382) );
  NAND U987 ( .A(n13481), .B(n13480), .Z(n423) );
  NANDN U988 ( .A(n13483), .B(n13482), .Z(n424) );
  NAND U989 ( .A(n423), .B(n424), .Z(n13636) );
  NAND U990 ( .A(n13448), .B(n13447), .Z(n425) );
  NAND U991 ( .A(n13445), .B(n13446), .Z(n426) );
  NAND U992 ( .A(n425), .B(n426), .Z(n13632) );
  NAND U993 ( .A(n13658), .B(n13657), .Z(n427) );
  NANDN U994 ( .A(n13656), .B(n13655), .Z(n428) );
  AND U995 ( .A(n427), .B(n428), .Z(n13844) );
  NAND U996 ( .A(n14199), .B(n14198), .Z(n429) );
  NANDN U997 ( .A(n14201), .B(n14200), .Z(n430) );
  AND U998 ( .A(n429), .B(n430), .Z(n14420) );
  XNOR U999 ( .A(n14434), .B(n14433), .Z(n14305) );
  XNOR U1000 ( .A(n14513), .B(n14512), .Z(n14514) );
  XNOR U1001 ( .A(n14699), .B(n14698), .Z(n14748) );
  XNOR U1002 ( .A(n14993), .B(n14992), .Z(n14990) );
  XNOR U1003 ( .A(n9632), .B(n9631), .Z(n9633) );
  XNOR U1004 ( .A(n9600), .B(n9599), .Z(n9591) );
  XNOR U1005 ( .A(n9652), .B(n9651), .Z(n9653) );
  XOR U1006 ( .A(n9744), .B(n9745), .Z(n9729) );
  XNOR U1007 ( .A(n9856), .B(n9855), .Z(n9805) );
  XNOR U1008 ( .A(n10304), .B(n10303), .Z(n10305) );
  XNOR U1009 ( .A(n10310), .B(n10309), .Z(n10312) );
  XNOR U1010 ( .A(n10586), .B(n10585), .Z(n10588) );
  XNOR U1011 ( .A(n10957), .B(n10956), .Z(n10943) );
  XNOR U1012 ( .A(n11243), .B(n11242), .Z(n11244) );
  XOR U1013 ( .A(n11458), .B(n11457), .Z(n11512) );
  XOR U1014 ( .A(n11550), .B(n11549), .Z(n11560) );
  XNOR U1015 ( .A(n11439), .B(n11438), .Z(n11441) );
  XNOR U1016 ( .A(n11574), .B(n11573), .Z(n11427) );
  XNOR U1017 ( .A(n6692), .B(n6691), .Z(n6693) );
  XNOR U1018 ( .A(n6916), .B(n6915), .Z(n6865) );
  XOR U1019 ( .A(n7081), .B(n7080), .Z(n7072) );
  XNOR U1020 ( .A(n7327), .B(n7326), .Z(n7329) );
  XOR U1021 ( .A(n7544), .B(n7543), .Z(n7548) );
  XNOR U1022 ( .A(n7662), .B(n7661), .Z(n7663) );
  XNOR U1023 ( .A(n8368), .B(n8367), .Z(n8371) );
  XNOR U1024 ( .A(n8391), .B(n8390), .Z(n8393) );
  XNOR U1025 ( .A(n8562), .B(n8561), .Z(n8564) );
  XNOR U1026 ( .A(n9003), .B(n9002), .Z(n9035) );
  XNOR U1027 ( .A(n8844), .B(n8843), .Z(n8736) );
  XNOR U1028 ( .A(n8836), .B(n8835), .Z(n8837) );
  XNOR U1029 ( .A(n3874), .B(n3873), .Z(n3875) );
  XNOR U1030 ( .A(n3804), .B(n3803), .Z(n3805) );
  XOR U1031 ( .A(n3810), .B(n3809), .Z(n3798) );
  XOR U1032 ( .A(n3968), .B(n3967), .Z(n3962) );
  XNOR U1033 ( .A(n4118), .B(n4117), .Z(n4119) );
  XNOR U1034 ( .A(n4331), .B(n4330), .Z(n4332) );
  XOR U1035 ( .A(n4351), .B(n4350), .Z(n4366) );
  XNOR U1036 ( .A(n4459), .B(n4458), .Z(n4460) );
  XNOR U1037 ( .A(n4554), .B(n4553), .Z(n4573) );
  NAND U1038 ( .A(n4427), .B(n4426), .Z(n431) );
  NANDN U1039 ( .A(n4429), .B(n4428), .Z(n432) );
  AND U1040 ( .A(n431), .B(n432), .Z(n4565) );
  XNOR U1041 ( .A(n4812), .B(n4811), .Z(n4803) );
  XNOR U1042 ( .A(n5740), .B(n5739), .Z(n5683) );
  XNOR U1043 ( .A(n5689), .B(n5688), .Z(n5773) );
  NAND U1044 ( .A(n5707), .B(n5706), .Z(n433) );
  NANDN U1045 ( .A(n5705), .B(n5704), .Z(n434) );
  NAND U1046 ( .A(n433), .B(n434), .Z(n5892) );
  NAND U1047 ( .A(n5863), .B(n5862), .Z(n435) );
  NAND U1048 ( .A(n5860), .B(n5861), .Z(n436) );
  NAND U1049 ( .A(n435), .B(n436), .Z(n6068) );
  XNOR U1050 ( .A(n6044), .B(n6043), .Z(n6062) );
  XNOR U1051 ( .A(n884), .B(o[9]), .Z(n874) );
  XOR U1052 ( .A(n1061), .B(n1062), .Z(n1046) );
  XNOR U1053 ( .A(n1896), .B(n1895), .Z(n1897) );
  XNOR U1054 ( .A(n2080), .B(n2079), .Z(n2071) );
  XNOR U1055 ( .A(n2316), .B(n2315), .Z(n2317) );
  XNOR U1056 ( .A(n2729), .B(n2728), .Z(n2723) );
  XNOR U1057 ( .A(n2767), .B(n2766), .Z(n2635) );
  NAND U1058 ( .A(n2890), .B(n2889), .Z(n437) );
  NANDN U1059 ( .A(n2888), .B(n2887), .Z(n438) );
  NAND U1060 ( .A(n437), .B(n438), .Z(n3066) );
  XNOR U1061 ( .A(n3328), .B(n3327), .Z(n3325) );
  XNOR U1062 ( .A(n12279), .B(o[132]), .Z(n12283) );
  XOR U1063 ( .A(n12451), .B(n12450), .Z(n12413) );
  XOR U1064 ( .A(n12831), .B(n12830), .Z(n12880) );
  XOR U1065 ( .A(n13082), .B(n13081), .Z(n13177) );
  NAND U1066 ( .A(n13615), .B(n13614), .Z(n439) );
  NANDN U1067 ( .A(n13613), .B(n13612), .Z(n440) );
  NAND U1068 ( .A(n439), .B(n440), .Z(n13645) );
  NAND U1069 ( .A(n13742), .B(n13741), .Z(n441) );
  NANDN U1070 ( .A(n13744), .B(n13743), .Z(n442) );
  AND U1071 ( .A(n441), .B(n442), .Z(n13756) );
  NAND U1072 ( .A(n14145), .B(n14144), .Z(n443) );
  NANDN U1073 ( .A(n14147), .B(n14146), .Z(n444) );
  NAND U1074 ( .A(n443), .B(n444), .Z(n14298) );
  NAND U1075 ( .A(n14191), .B(n14190), .Z(n445) );
  NANDN U1076 ( .A(n14189), .B(n14188), .Z(n446) );
  AND U1077 ( .A(n445), .B(n446), .Z(n14295) );
  XNOR U1078 ( .A(n14549), .B(n14548), .Z(n14550) );
  XNOR U1079 ( .A(n14509), .B(n14508), .Z(n14589) );
  XNOR U1080 ( .A(n14651), .B(n14650), .Z(n14652) );
  XNOR U1081 ( .A(n14987), .B(n14986), .Z(n14984) );
  XOR U1082 ( .A(n14811), .B(n14810), .Z(n14809) );
  XOR U1083 ( .A(n14823), .B(n14822), .Z(n14821) );
  XNOR U1084 ( .A(n9476), .B(n9475), .Z(n9478) );
  XOR U1085 ( .A(n9463), .B(n9376), .Z(n447) );
  NANDN U1086 ( .A(n9377), .B(n447), .Z(n448) );
  NAND U1087 ( .A(n9463), .B(n9376), .Z(n449) );
  AND U1088 ( .A(n448), .B(n449), .Z(n9429) );
  XOR U1089 ( .A(n9702), .B(n9701), .Z(n9684) );
  XNOR U1090 ( .A(n10428), .B(n10427), .Z(n10429) );
  OR U1091 ( .A(n10424), .B(n10423), .Z(n450) );
  NAND U1092 ( .A(n10425), .B(n10426), .Z(n451) );
  AND U1093 ( .A(n450), .B(n451), .Z(n10552) );
  XNOR U1094 ( .A(n10700), .B(n10699), .Z(n10823) );
  XOR U1095 ( .A(n11121), .B(n11120), .Z(n11123) );
  XNOR U1096 ( .A(n11284), .B(n11283), .Z(n11286) );
  XOR U1097 ( .A(n11705), .B(n11704), .Z(n11600) );
  XNOR U1098 ( .A(n11697), .B(n11696), .Z(n11698) );
  XNOR U1099 ( .A(n11727), .B(n11726), .Z(n11728) );
  XNOR U1100 ( .A(n11794), .B(n11793), .Z(n11800) );
  XNOR U1101 ( .A(n11960), .B(n11959), .Z(n11957) );
  XNOR U1102 ( .A(n11870), .B(n11869), .Z(n11894) );
  XOR U1103 ( .A(n11974), .B(n11973), .Z(n11972) );
  XOR U1104 ( .A(n11966), .B(n11965), .Z(n11964) );
  XOR U1105 ( .A(n11741), .B(n11740), .Z(n11588) );
  XNOR U1106 ( .A(n6527), .B(n6526), .Z(n6528) );
  XNOR U1107 ( .A(n6860), .B(n6859), .Z(n6862) );
  XOR U1108 ( .A(n7316), .B(n7315), .Z(n7229) );
  XNOR U1109 ( .A(n8243), .B(n8242), .Z(n8245) );
  XNOR U1110 ( .A(n8550), .B(n8549), .Z(n8552) );
  XNOR U1111 ( .A(n8729), .B(n8728), .Z(n8730) );
  XNOR U1112 ( .A(n8983), .B(n8982), .Z(n8984) );
  NAND U1113 ( .A(n8820), .B(n8819), .Z(n452) );
  NANDN U1114 ( .A(n8822), .B(n8821), .Z(n453) );
  NAND U1115 ( .A(n452), .B(n453), .Z(n8988) );
  XOR U1116 ( .A(n9072), .B(n9071), .Z(n9070) );
  XOR U1117 ( .A(n9060), .B(n9059), .Z(n9058) );
  XNOR U1118 ( .A(n9262), .B(n9261), .Z(n9260) );
  XOR U1119 ( .A(n9236), .B(n9235), .Z(n9234) );
  XNOR U1120 ( .A(n9090), .B(n8935), .Z(n8936) );
  XNOR U1121 ( .A(n8941), .B(n8940), .Z(n8942) );
  XOR U1122 ( .A(n3761), .B(n3760), .Z(n3721) );
  XNOR U1123 ( .A(n3834), .B(n3833), .Z(n3835) );
  XNOR U1124 ( .A(n4084), .B(n4083), .Z(n4051) );
  XNOR U1125 ( .A(n4059), .B(n4058), .Z(n4046) );
  NAND U1126 ( .A(n4570), .B(n4569), .Z(n454) );
  NAND U1127 ( .A(n4567), .B(n4568), .Z(n455) );
  NAND U1128 ( .A(n454), .B(n455), .Z(n4686) );
  XNOR U1129 ( .A(n4594), .B(n4593), .Z(n4693) );
  NAND U1130 ( .A(n4921), .B(n4920), .Z(n456) );
  NANDN U1131 ( .A(n4923), .B(n4922), .Z(n457) );
  AND U1132 ( .A(n456), .B(n457), .Z(n4954) );
  XNOR U1133 ( .A(n5366), .B(n5365), .Z(n5368) );
  XOR U1134 ( .A(n5360), .B(n5359), .Z(n5362) );
  XNOR U1135 ( .A(n5669), .B(n5668), .Z(n5671) );
  XNOR U1136 ( .A(n5663), .B(n5662), .Z(n5664) );
  XOR U1137 ( .A(n5815), .B(n5814), .Z(n5809) );
  XNOR U1138 ( .A(n5825), .B(n5824), .Z(n5826) );
  NAND U1139 ( .A(n5745), .B(n5744), .Z(n458) );
  NAND U1140 ( .A(n5743), .B(n6180), .Z(n459) );
  NAND U1141 ( .A(n458), .B(n459), .Z(n5932) );
  NAND U1142 ( .A(n5749), .B(n5748), .Z(n460) );
  NAND U1143 ( .A(n5746), .B(n5747), .Z(n461) );
  NAND U1144 ( .A(n460), .B(n461), .Z(n5928) );
  NAND U1145 ( .A(n5897), .B(n5896), .Z(n462) );
  NAND U1146 ( .A(n5894), .B(n5895), .Z(n463) );
  NAND U1147 ( .A(n462), .B(n463), .Z(n6055) );
  XNOR U1148 ( .A(n6253), .B(n6252), .Z(n6250) );
  XOR U1149 ( .A(n6115), .B(n6114), .Z(n6113) );
  NAND U1150 ( .A(n5878), .B(n5877), .Z(n464) );
  NAND U1151 ( .A(n5875), .B(n5876), .Z(n465) );
  NAND U1152 ( .A(n464), .B(n465), .Z(n6030) );
  OR U1153 ( .A(n6073), .B(n6072), .Z(n466) );
  NAND U1154 ( .A(n6075), .B(n6074), .Z(n467) );
  NAND U1155 ( .A(n466), .B(n467), .Z(n6299) );
  XNOR U1156 ( .A(n6296), .B(n6295), .Z(n6293) );
  XOR U1157 ( .A(n6125), .B(n6124), .Z(n6123) );
  XNOR U1158 ( .A(n861), .B(n860), .Z(n863) );
  XNOR U1159 ( .A(n929), .B(n928), .Z(n920) );
  XOR U1160 ( .A(n1017), .B(n1016), .Z(n1019) );
  XOR U1161 ( .A(n1467), .B(n1466), .Z(n1469) );
  XOR U1162 ( .A(n1461), .B(n1460), .Z(n1463) );
  XNOR U1163 ( .A(n1775), .B(n1774), .Z(n1787) );
  XNOR U1164 ( .A(n1594), .B(n1593), .Z(n1587) );
  XOR U1165 ( .A(n1932), .B(n1931), .Z(n1925) );
  XNOR U1166 ( .A(n2200), .B(n2199), .Z(n2184) );
  XNOR U1167 ( .A(n2448), .B(n2447), .Z(n2449) );
  XNOR U1168 ( .A(n2480), .B(n2479), .Z(n2482) );
  XNOR U1169 ( .A(n2927), .B(n2926), .Z(n2790) );
  XOR U1170 ( .A(n2940), .B(n2939), .Z(n2934) );
  NAND U1171 ( .A(n2861), .B(n2860), .Z(n468) );
  NANDN U1172 ( .A(n2859), .B(n2858), .Z(n469) );
  AND U1173 ( .A(n468), .B(n469), .Z(n3047) );
  XNOR U1174 ( .A(n3267), .B(n3266), .Z(n3268) );
  XNOR U1175 ( .A(n3303), .B(n3302), .Z(n3300) );
  XOR U1176 ( .A(n3297), .B(n3296), .Z(n3295) );
  XNOR U1177 ( .A(n3317), .B(n3316), .Z(n3314) );
  XNOR U1178 ( .A(n12329), .B(n12328), .Z(n12331) );
  XNOR U1179 ( .A(n13511), .B(n13510), .Z(n13512) );
  NAND U1180 ( .A(n14143), .B(n14142), .Z(n470) );
  NAND U1181 ( .A(n14140), .B(n14141), .Z(n471) );
  NAND U1182 ( .A(n470), .B(n471), .Z(n14285) );
  XNOR U1183 ( .A(n14739), .B(n14738), .Z(n14638) );
  XNOR U1184 ( .A(n14645), .B(n14644), .Z(n14646) );
  XNOR U1185 ( .A(n14730), .B(n14729), .Z(n14731) );
  XOR U1186 ( .A(n15051), .B(n15050), .Z(n15049) );
  XNOR U1187 ( .A(n15027), .B(n15026), .Z(n15024) );
  XNOR U1188 ( .A(n9718), .B(n9717), .Z(n9781) );
  XNOR U1189 ( .A(n9860), .B(n9859), .Z(n9861) );
  OR U1190 ( .A(n10242), .B(n10243), .Z(n472) );
  NAND U1191 ( .A(n10240), .B(n10241), .Z(n473) );
  NAND U1192 ( .A(n472), .B(n473), .Z(n10444) );
  XNOR U1193 ( .A(n10961), .B(n10960), .Z(n10962) );
  XNOR U1194 ( .A(n11889), .B(n11888), .Z(n11891) );
  XNOR U1195 ( .A(n12184), .B(n12183), .Z(n12182) );
  XNOR U1196 ( .A(n12160), .B(n12159), .Z(n12158) );
  XOR U1197 ( .A(n6408), .B(n6407), .Z(n474) );
  NANDN U1198 ( .A(n6409), .B(n474), .Z(n475) );
  NAND U1199 ( .A(n6408), .B(n6407), .Z(n476) );
  AND U1200 ( .A(n475), .B(n476), .Z(n6434) );
  XNOR U1201 ( .A(n7113), .B(n7112), .Z(n7205) );
  XOR U1202 ( .A(n3586), .B(n3585), .Z(n477) );
  NANDN U1203 ( .A(n3587), .B(n477), .Z(n478) );
  NAND U1204 ( .A(n3586), .B(n3585), .Z(n479) );
  AND U1205 ( .A(n478), .B(n479), .Z(n3612) );
  XNOR U1206 ( .A(n4025), .B(n4024), .Z(n4027) );
  XNOR U1207 ( .A(n4376), .B(n4375), .Z(n4378) );
  XOR U1208 ( .A(n5960), .B(n5959), .Z(n5962) );
  NAND U1209 ( .A(n6006), .B(n6005), .Z(n480) );
  NANDN U1210 ( .A(n6008), .B(n6007), .Z(n481) );
  AND U1211 ( .A(n480), .B(n481), .Z(n6093) );
  XOR U1212 ( .A(n6347), .B(n6346), .Z(n482) );
  XNOR U1213 ( .A(n6348), .B(n482), .Z(n6328) );
  NAND U1214 ( .A(n6059), .B(n6058), .Z(n483) );
  NANDN U1215 ( .A(n6061), .B(n6060), .Z(n484) );
  AND U1216 ( .A(n483), .B(n484), .Z(n6309) );
  NAND U1217 ( .A(n5988), .B(n5987), .Z(n485) );
  NAND U1218 ( .A(n5985), .B(n5986), .Z(n486) );
  AND U1219 ( .A(n485), .B(n486), .Z(n6096) );
  XNOR U1220 ( .A(n1035), .B(n1034), .Z(n1101) );
  XNOR U1221 ( .A(n2046), .B(n2045), .Z(n2048) );
  XNOR U1222 ( .A(n2053), .B(n2052), .Z(n2054) );
  XOR U1223 ( .A(n2456), .B(n2455), .Z(n2467) );
  NAND U1224 ( .A(n3065), .B(n3064), .Z(n487) );
  NAND U1225 ( .A(n3062), .B(n3063), .Z(n488) );
  NAND U1226 ( .A(n487), .B(n488), .Z(n3114) );
  XNOR U1227 ( .A(n3515), .B(n3514), .Z(n3513) );
  XNOR U1228 ( .A(n3505), .B(n3504), .Z(n3502) );
  XNOR U1229 ( .A(n3137), .B(n3136), .Z(n3139) );
  XOR U1230 ( .A(n12318), .B(n12319), .Z(n489) );
  NANDN U1231 ( .A(n12320), .B(n489), .Z(n490) );
  NAND U1232 ( .A(n12318), .B(n12319), .Z(n491) );
  AND U1233 ( .A(n490), .B(n491), .Z(n12336) );
  NAND U1234 ( .A(n12570), .B(n12571), .Z(n492) );
  XOR U1235 ( .A(n12570), .B(n12571), .Z(n493) );
  NANDN U1236 ( .A(n12569), .B(n493), .Z(n494) );
  NAND U1237 ( .A(n492), .B(n494), .Z(n12633) );
  XOR U1238 ( .A(n12727), .B(n12728), .Z(n495) );
  NANDN U1239 ( .A(n12729), .B(n495), .Z(n496) );
  NAND U1240 ( .A(n12727), .B(n12728), .Z(n497) );
  AND U1241 ( .A(n496), .B(n497), .Z(n12804) );
  XOR U1242 ( .A(n13063), .B(n13064), .Z(n498) );
  NANDN U1243 ( .A(n13065), .B(n498), .Z(n499) );
  NAND U1244 ( .A(n13063), .B(n13064), .Z(n500) );
  AND U1245 ( .A(n499), .B(n500), .Z(n13171) );
  XNOR U1246 ( .A(n13527), .B(n13526), .Z(n13532) );
  NAND U1247 ( .A(n13866), .B(n13867), .Z(n501) );
  XOR U1248 ( .A(n13866), .B(n13867), .Z(n502) );
  NANDN U1249 ( .A(n13865), .B(n502), .Z(n503) );
  NAND U1250 ( .A(n501), .B(n503), .Z(n13988) );
  XOR U1251 ( .A(n14273), .B(n14274), .Z(n504) );
  NANDN U1252 ( .A(n14275), .B(n504), .Z(n505) );
  NAND U1253 ( .A(n14273), .B(n14274), .Z(n506) );
  AND U1254 ( .A(n505), .B(n506), .Z(n14290) );
  NAND U1255 ( .A(n14612), .B(n14613), .Z(n507) );
  XOR U1256 ( .A(n14612), .B(n14613), .Z(n508) );
  NANDN U1257 ( .A(n14611), .B(n508), .Z(n509) );
  NAND U1258 ( .A(n507), .B(n509), .Z(n15071) );
  XOR U1259 ( .A(n9388), .B(n9389), .Z(n510) );
  NANDN U1260 ( .A(n9390), .B(n510), .Z(n511) );
  NAND U1261 ( .A(n9388), .B(n9389), .Z(n512) );
  AND U1262 ( .A(n511), .B(n512), .Z(n9424) );
  XOR U1263 ( .A(n9519), .B(n9520), .Z(n513) );
  NANDN U1264 ( .A(n9521), .B(n513), .Z(n514) );
  NAND U1265 ( .A(n9519), .B(n9520), .Z(n515) );
  AND U1266 ( .A(n514), .B(n515), .Z(n9573) );
  XOR U1267 ( .A(n9705), .B(n9706), .Z(n516) );
  NANDN U1268 ( .A(n9707), .B(n516), .Z(n517) );
  NAND U1269 ( .A(n9705), .B(n9706), .Z(n518) );
  AND U1270 ( .A(n517), .B(n518), .Z(n9786) );
  XOR U1271 ( .A(n10036), .B(n10037), .Z(n519) );
  NANDN U1272 ( .A(n10038), .B(n519), .Z(n520) );
  NAND U1273 ( .A(n10036), .B(n10037), .Z(n521) );
  AND U1274 ( .A(n520), .B(n521), .Z(n10128) );
  XOR U1275 ( .A(n10327), .B(n10328), .Z(n522) );
  NANDN U1276 ( .A(n10329), .B(n522), .Z(n523) );
  NAND U1277 ( .A(n10327), .B(n10328), .Z(n524) );
  AND U1278 ( .A(n523), .B(n524), .Z(n10440) );
  NAND U1279 ( .A(n10694), .B(n10695), .Z(n525) );
  XOR U1280 ( .A(n10694), .B(n10695), .Z(n526) );
  NANDN U1281 ( .A(n10693), .B(n526), .Z(n527) );
  NAND U1282 ( .A(n525), .B(n527), .Z(n10820) );
  XOR U1283 ( .A(n11254), .B(n11255), .Z(n528) );
  NANDN U1284 ( .A(n11256), .B(n528), .Z(n529) );
  NAND U1285 ( .A(n11254), .B(n11255), .Z(n530) );
  AND U1286 ( .A(n529), .B(n530), .Z(n11272) );
  XOR U1287 ( .A(n11744), .B(n11745), .Z(n531) );
  NANDN U1288 ( .A(n11746), .B(n531), .Z(n532) );
  NAND U1289 ( .A(n11744), .B(n11745), .Z(n533) );
  AND U1290 ( .A(n532), .B(n533), .Z(n11755) );
  XNOR U1291 ( .A(n12222), .B(n12221), .Z(n12219) );
  NAND U1292 ( .A(n6430), .B(n6429), .Z(n534) );
  NANDN U1293 ( .A(n6432), .B(n6431), .Z(n535) );
  NAND U1294 ( .A(n534), .B(n535), .Z(n6447) );
  XOR U1295 ( .A(n6532), .B(n6533), .Z(n536) );
  NANDN U1296 ( .A(n6534), .B(n536), .Z(n537) );
  NAND U1297 ( .A(n6532), .B(n6533), .Z(n538) );
  AND U1298 ( .A(n537), .B(n538), .Z(n6586) );
  XOR U1299 ( .A(n6697), .B(n6698), .Z(n539) );
  NANDN U1300 ( .A(n6699), .B(n539), .Z(n540) );
  NAND U1301 ( .A(n6697), .B(n6698), .Z(n541) );
  AND U1302 ( .A(n540), .B(n541), .Z(n6763) );
  XOR U1303 ( .A(n7004), .B(n7005), .Z(n542) );
  NANDN U1304 ( .A(n7006), .B(n542), .Z(n543) );
  NAND U1305 ( .A(n7004), .B(n7005), .Z(n544) );
  AND U1306 ( .A(n543), .B(n544), .Z(n7098) );
  XNOR U1307 ( .A(n7213), .B(n7212), .Z(n7219) );
  XOR U1308 ( .A(n7443), .B(n7444), .Z(n545) );
  NANDN U1309 ( .A(n7445), .B(n545), .Z(n546) );
  NAND U1310 ( .A(n7443), .B(n7444), .Z(n547) );
  AND U1311 ( .A(n546), .B(n547), .Z(n7669) );
  XOR U1312 ( .A(n7948), .B(n7949), .Z(n548) );
  NANDN U1313 ( .A(n7950), .B(n548), .Z(n549) );
  NAND U1314 ( .A(n7948), .B(n7949), .Z(n550) );
  AND U1315 ( .A(n549), .B(n550), .Z(n8220) );
  XOR U1316 ( .A(n8546), .B(n8547), .Z(n551) );
  NANDN U1317 ( .A(n8548), .B(n551), .Z(n552) );
  NAND U1318 ( .A(n8546), .B(n8547), .Z(n553) );
  AND U1319 ( .A(n552), .B(n553), .Z(n8704) );
  NAND U1320 ( .A(n3608), .B(n3607), .Z(n554) );
  NANDN U1321 ( .A(n3610), .B(n3609), .Z(n555) );
  NAND U1322 ( .A(n554), .B(n555), .Z(n3625) );
  XOR U1323 ( .A(n3710), .B(n3711), .Z(n556) );
  NANDN U1324 ( .A(n3712), .B(n556), .Z(n557) );
  NAND U1325 ( .A(n3710), .B(n3711), .Z(n558) );
  AND U1326 ( .A(n557), .B(n558), .Z(n3728) );
  XNOR U1327 ( .A(n3823), .B(n3822), .Z(n3816) );
  XOR U1328 ( .A(n3895), .B(n3896), .Z(n559) );
  NANDN U1329 ( .A(n3897), .B(n559), .Z(n560) );
  NAND U1330 ( .A(n3895), .B(n3896), .Z(n561) );
  AND U1331 ( .A(n560), .B(n561), .Z(n4019) );
  NAND U1332 ( .A(n4289), .B(n4288), .Z(n562) );
  XOR U1333 ( .A(n4289), .B(n4288), .Z(n563) );
  NANDN U1334 ( .A(n4290), .B(n563), .Z(n564) );
  NAND U1335 ( .A(n562), .B(n564), .Z(n4373) );
  XOR U1336 ( .A(n4589), .B(n4588), .Z(n565) );
  NANDN U1337 ( .A(n4587), .B(n565), .Z(n566) );
  NAND U1338 ( .A(n4589), .B(n4588), .Z(n567) );
  AND U1339 ( .A(n566), .B(n567), .Z(n4703) );
  XOR U1340 ( .A(n4931), .B(n4930), .Z(n568) );
  NANDN U1341 ( .A(n4932), .B(n568), .Z(n569) );
  NAND U1342 ( .A(n4931), .B(n4930), .Z(n570) );
  AND U1343 ( .A(n569), .B(n570), .Z(n4948) );
  NAND U1344 ( .A(n5347), .B(n5346), .Z(n571) );
  XOR U1345 ( .A(n5347), .B(n5346), .Z(n572) );
  NANDN U1346 ( .A(n5348), .B(n572), .Z(n573) );
  NAND U1347 ( .A(n571), .B(n573), .Z(n5357) );
  NAND U1348 ( .A(n5797), .B(n5798), .Z(n574) );
  XOR U1349 ( .A(n5797), .B(n5798), .Z(n575) );
  NANDN U1350 ( .A(n5796), .B(n575), .Z(n576) );
  NAND U1351 ( .A(n574), .B(n576), .Z(n5940) );
  XNOR U1352 ( .A(n6357), .B(n6356), .Z(n6355) );
  XOR U1353 ( .A(n649), .B(n648), .Z(n577) );
  NANDN U1354 ( .A(n650), .B(n577), .Z(n578) );
  NAND U1355 ( .A(n649), .B(n648), .Z(n579) );
  AND U1356 ( .A(n578), .B(n579), .Z(n672) );
  XOR U1357 ( .A(n787), .B(n788), .Z(n580) );
  NANDN U1358 ( .A(n789), .B(n580), .Z(n581) );
  NAND U1359 ( .A(n787), .B(n788), .Z(n582) );
  AND U1360 ( .A(n581), .B(n582), .Z(n805) );
  XOR U1361 ( .A(n1029), .B(n1028), .Z(n583) );
  NANDN U1362 ( .A(n1030), .B(n583), .Z(n584) );
  NAND U1363 ( .A(n1029), .B(n1028), .Z(n585) );
  AND U1364 ( .A(n584), .B(n585), .Z(n1096) );
  XOR U1365 ( .A(n1265), .B(n1264), .Z(n586) );
  NANDN U1366 ( .A(n1266), .B(n586), .Z(n587) );
  NAND U1367 ( .A(n1265), .B(n1264), .Z(n588) );
  AND U1368 ( .A(n587), .B(n588), .Z(n1350) );
  XOR U1369 ( .A(n1556), .B(n1557), .Z(n589) );
  NANDN U1370 ( .A(n1558), .B(n589), .Z(n590) );
  NAND U1371 ( .A(n1556), .B(n1557), .Z(n591) );
  AND U1372 ( .A(n590), .B(n591), .Z(n1573) );
  XOR U1373 ( .A(n1913), .B(n1914), .Z(n592) );
  NANDN U1374 ( .A(n1915), .B(n592), .Z(n593) );
  NAND U1375 ( .A(n1913), .B(n1914), .Z(n594) );
  AND U1376 ( .A(n593), .B(n594), .Z(n2040) );
  XOR U1377 ( .A(n2786), .B(n2787), .Z(n595) );
  NANDN U1378 ( .A(n2788), .B(n595), .Z(n596) );
  NAND U1379 ( .A(n2786), .B(n2787), .Z(n597) );
  AND U1380 ( .A(n596), .B(n597), .Z(n3091) );
  XNOR U1381 ( .A(n3281), .B(n3280), .Z(n3278) );
  NAND U1382 ( .A(n9040), .B(n9039), .Z(n598) );
  NANDN U1383 ( .A(n9042), .B(n9041), .Z(n599) );
  AND U1384 ( .A(n598), .B(n599), .Z(n600) );
  NAND U1385 ( .A(n9043), .B(n9044), .Z(n601) );
  NAND U1386 ( .A(n9045), .B(n9046), .Z(n602) );
  AND U1387 ( .A(n601), .B(n602), .Z(n603) );
  XOR U1388 ( .A(n9288), .B(n9287), .Z(n604) );
  XNOR U1389 ( .A(n9274), .B(n9273), .Z(n605) );
  XNOR U1390 ( .A(n604), .B(n605), .Z(n606) );
  AND U1391 ( .A(n9300), .B(n9299), .Z(n607) );
  NAND U1392 ( .A(n9294), .B(n9293), .Z(n608) );
  XNOR U1393 ( .A(n607), .B(n608), .Z(n609) );
  XOR U1394 ( .A(n606), .B(n609), .Z(n610) );
  XNOR U1395 ( .A(n600), .B(n603), .Z(n611) );
  XNOR U1396 ( .A(n610), .B(n611), .Z(n612) );
  NANDN U1397 ( .A(n9303), .B(n9304), .Z(n613) );
  NANDN U1398 ( .A(n9301), .B(n9302), .Z(n614) );
  AND U1399 ( .A(n613), .B(n614), .Z(n615) );
  XNOR U1400 ( .A(n612), .B(n615), .Z(N192) );
  AND U1401 ( .A(x[128]), .B(y[640]), .Z(n1273) );
  XOR U1402 ( .A(n1273), .B(o[0]), .Z(N33) );
  NAND U1403 ( .A(x[129]), .B(y[640]), .Z(n616) );
  AND U1404 ( .A(y[641]), .B(x[128]), .Z(n624) );
  XNOR U1405 ( .A(n624), .B(o[1]), .Z(n617) );
  XOR U1406 ( .A(n616), .B(n617), .Z(n619) );
  NAND U1407 ( .A(n1273), .B(o[0]), .Z(n618) );
  XNOR U1408 ( .A(n619), .B(n618), .Z(N34) );
  IV U1409 ( .A(n616), .Z(n628) );
  NANDN U1410 ( .A(n628), .B(n617), .Z(n621) );
  NAND U1411 ( .A(n619), .B(n618), .Z(n620) );
  AND U1412 ( .A(n621), .B(n620), .Z(n634) );
  AND U1413 ( .A(y[642]), .B(x[128]), .Z(n627) );
  XNOR U1414 ( .A(n627), .B(o[2]), .Z(n633) );
  XNOR U1415 ( .A(n634), .B(n633), .Z(n636) );
  AND U1416 ( .A(y[640]), .B(x[130]), .Z(n623) );
  NAND U1417 ( .A(x[129]), .B(y[641]), .Z(n622) );
  XNOR U1418 ( .A(n623), .B(n622), .Z(n630) );
  AND U1419 ( .A(n624), .B(o[1]), .Z(n629) );
  XNOR U1420 ( .A(n630), .B(n629), .Z(n635) );
  XNOR U1421 ( .A(n636), .B(n635), .Z(N35) );
  AND U1422 ( .A(y[642]), .B(x[129]), .Z(n760) );
  NAND U1423 ( .A(y[641]), .B(x[130]), .Z(n646) );
  XNOR U1424 ( .A(o[3]), .B(n646), .Z(n651) );
  XOR U1425 ( .A(n760), .B(n651), .Z(n653) );
  AND U1426 ( .A(y[643]), .B(x[128]), .Z(n626) );
  NAND U1427 ( .A(y[640]), .B(x[131]), .Z(n625) );
  XNOR U1428 ( .A(n626), .B(n625), .Z(n640) );
  NAND U1429 ( .A(n627), .B(o[2]), .Z(n641) );
  XNOR U1430 ( .A(n653), .B(n652), .Z(n650) );
  NANDN U1431 ( .A(n646), .B(n628), .Z(n632) );
  NAND U1432 ( .A(n630), .B(n629), .Z(n631) );
  NAND U1433 ( .A(n632), .B(n631), .Z(n648) );
  NANDN U1434 ( .A(n634), .B(n633), .Z(n638) );
  NAND U1435 ( .A(n636), .B(n635), .Z(n637) );
  AND U1436 ( .A(n638), .B(n637), .Z(n649) );
  XOR U1437 ( .A(n648), .B(n649), .Z(n639) );
  XNOR U1438 ( .A(n650), .B(n639), .Z(N36) );
  AND U1439 ( .A(x[131]), .B(y[643]), .Z(n701) );
  NAND U1440 ( .A(n1273), .B(n701), .Z(n643) );
  NANDN U1441 ( .A(n641), .B(n640), .Z(n642) );
  AND U1442 ( .A(n643), .B(n642), .Z(n680) );
  AND U1443 ( .A(y[640]), .B(x[132]), .Z(n645) );
  NAND U1444 ( .A(x[128]), .B(y[644]), .Z(n644) );
  XNOR U1445 ( .A(n645), .B(n644), .Z(n667) );
  ANDN U1446 ( .B(o[3]), .A(n646), .Z(n666) );
  XOR U1447 ( .A(n667), .B(n666), .Z(n678) );
  AND U1448 ( .A(y[643]), .B(x[129]), .Z(n878) );
  NAND U1449 ( .A(x[130]), .B(y[642]), .Z(n647) );
  XNOR U1450 ( .A(n878), .B(n647), .Z(n663) );
  NAND U1451 ( .A(y[641]), .B(x[131]), .Z(n661) );
  XNOR U1452 ( .A(o[4]), .B(n661), .Z(n662) );
  XOR U1453 ( .A(n663), .B(n662), .Z(n677) );
  XOR U1454 ( .A(n678), .B(n677), .Z(n679) );
  XOR U1455 ( .A(n680), .B(n679), .Z(n673) );
  NAND U1456 ( .A(n760), .B(n651), .Z(n655) );
  NAND U1457 ( .A(n653), .B(n652), .Z(n654) );
  NAND U1458 ( .A(n655), .B(n654), .Z(n671) );
  IV U1459 ( .A(n671), .Z(n670) );
  XOR U1460 ( .A(n672), .B(n670), .Z(n656) );
  XNOR U1461 ( .A(n673), .B(n656), .Z(N37) );
  AND U1462 ( .A(x[130]), .B(y[643]), .Z(n769) );
  AND U1463 ( .A(x[129]), .B(y[644]), .Z(n658) );
  NAND U1464 ( .A(x[131]), .B(y[642]), .Z(n657) );
  XNOR U1465 ( .A(n658), .B(n657), .Z(n685) );
  NAND U1466 ( .A(y[641]), .B(x[132]), .Z(n699) );
  XNOR U1467 ( .A(o[5]), .B(n699), .Z(n684) );
  XOR U1468 ( .A(n685), .B(n684), .Z(n688) );
  XOR U1469 ( .A(n769), .B(n688), .Z(n690) );
  AND U1470 ( .A(y[640]), .B(x[133]), .Z(n660) );
  NAND U1471 ( .A(x[128]), .B(y[645]), .Z(n659) );
  XNOR U1472 ( .A(n660), .B(n659), .Z(n694) );
  ANDN U1473 ( .B(o[4]), .A(n661), .Z(n693) );
  XOR U1474 ( .A(n694), .B(n693), .Z(n689) );
  XOR U1475 ( .A(n690), .B(n689), .Z(n713) );
  NAND U1476 ( .A(n769), .B(n760), .Z(n665) );
  NAND U1477 ( .A(n663), .B(n662), .Z(n664) );
  AND U1478 ( .A(n665), .B(n664), .Z(n711) );
  AND U1479 ( .A(y[644]), .B(x[132]), .Z(n1476) );
  NAND U1480 ( .A(n1476), .B(n1273), .Z(n669) );
  NAND U1481 ( .A(n667), .B(n666), .Z(n668) );
  NAND U1482 ( .A(n669), .B(n668), .Z(n710) );
  XNOR U1483 ( .A(n711), .B(n710), .Z(n712) );
  XNOR U1484 ( .A(n713), .B(n712), .Z(n706) );
  OR U1485 ( .A(n672), .B(n670), .Z(n676) );
  ANDN U1486 ( .B(n672), .A(n671), .Z(n674) );
  OR U1487 ( .A(n674), .B(n673), .Z(n675) );
  AND U1488 ( .A(n676), .B(n675), .Z(n705) );
  NAND U1489 ( .A(n678), .B(n677), .Z(n682) );
  NANDN U1490 ( .A(n680), .B(n679), .Z(n681) );
  NAND U1491 ( .A(n682), .B(n681), .Z(n704) );
  IV U1492 ( .A(n704), .Z(n703) );
  XOR U1493 ( .A(n705), .B(n703), .Z(n683) );
  XNOR U1494 ( .A(n706), .B(n683), .Z(N38) );
  AND U1495 ( .A(y[644]), .B(x[131]), .Z(n770) );
  NAND U1496 ( .A(n770), .B(n760), .Z(n687) );
  NAND U1497 ( .A(n685), .B(n684), .Z(n686) );
  AND U1498 ( .A(n687), .B(n686), .Z(n741) );
  NAND U1499 ( .A(n769), .B(n688), .Z(n692) );
  NAND U1500 ( .A(n690), .B(n689), .Z(n691) );
  NAND U1501 ( .A(n692), .B(n691), .Z(n740) );
  XNOR U1502 ( .A(n741), .B(n740), .Z(n743) );
  AND U1503 ( .A(y[645]), .B(x[133]), .Z(n956) );
  NAND U1504 ( .A(n1273), .B(n956), .Z(n696) );
  NAND U1505 ( .A(n694), .B(n693), .Z(n695) );
  NAND U1506 ( .A(n696), .B(n695), .Z(n717) );
  AND U1507 ( .A(y[640]), .B(x[134]), .Z(n698) );
  NAND U1508 ( .A(x[128]), .B(y[646]), .Z(n697) );
  XNOR U1509 ( .A(n698), .B(n697), .Z(n725) );
  ANDN U1510 ( .B(o[5]), .A(n699), .Z(n724) );
  XOR U1511 ( .A(n725), .B(n724), .Z(n718) );
  XOR U1512 ( .A(n717), .B(n718), .Z(n720) );
  NAND U1513 ( .A(x[130]), .B(y[644]), .Z(n700) );
  XNOR U1514 ( .A(n701), .B(n700), .Z(n729) );
  AND U1515 ( .A(x[129]), .B(y[645]), .Z(n994) );
  NAND U1516 ( .A(x[132]), .B(y[642]), .Z(n702) );
  XNOR U1517 ( .A(n994), .B(n702), .Z(n733) );
  AND U1518 ( .A(y[641]), .B(x[133]), .Z(n739) );
  XOR U1519 ( .A(n739), .B(o[6]), .Z(n732) );
  XOR U1520 ( .A(n733), .B(n732), .Z(n728) );
  XOR U1521 ( .A(n729), .B(n728), .Z(n719) );
  XOR U1522 ( .A(n720), .B(n719), .Z(n742) );
  XOR U1523 ( .A(n743), .B(n742), .Z(n749) );
  OR U1524 ( .A(n705), .B(n703), .Z(n709) );
  ANDN U1525 ( .B(n705), .A(n704), .Z(n707) );
  OR U1526 ( .A(n707), .B(n706), .Z(n708) );
  AND U1527 ( .A(n709), .B(n708), .Z(n747) );
  NANDN U1528 ( .A(n711), .B(n710), .Z(n715) );
  NAND U1529 ( .A(n713), .B(n712), .Z(n714) );
  AND U1530 ( .A(n715), .B(n714), .Z(n748) );
  IV U1531 ( .A(n748), .Z(n746) );
  XOR U1532 ( .A(n747), .B(n746), .Z(n716) );
  XNOR U1533 ( .A(n749), .B(n716), .Z(N39) );
  NAND U1534 ( .A(n718), .B(n717), .Z(n722) );
  NAND U1535 ( .A(n720), .B(n719), .Z(n721) );
  AND U1536 ( .A(n722), .B(n721), .Z(n793) );
  AND U1537 ( .A(x[129]), .B(y[646]), .Z(n1132) );
  NAND U1538 ( .A(x[133]), .B(y[642]), .Z(n723) );
  XNOR U1539 ( .A(n1132), .B(n723), .Z(n763) );
  NAND U1540 ( .A(y[641]), .B(x[134]), .Z(n767) );
  XNOR U1541 ( .A(o[7]), .B(n767), .Z(n762) );
  XOR U1542 ( .A(n763), .B(n762), .Z(n782) );
  AND U1543 ( .A(y[646]), .B(x[134]), .Z(n1014) );
  NAND U1544 ( .A(n1273), .B(n1014), .Z(n727) );
  NAND U1545 ( .A(n725), .B(n724), .Z(n726) );
  AND U1546 ( .A(n727), .B(n726), .Z(n781) );
  XNOR U1547 ( .A(n782), .B(n781), .Z(n783) );
  NAND U1548 ( .A(n769), .B(n770), .Z(n731) );
  NAND U1549 ( .A(n729), .B(n728), .Z(n730) );
  NAND U1550 ( .A(n731), .B(n730), .Z(n784) );
  XNOR U1551 ( .A(n783), .B(n784), .Z(n791) );
  AND U1552 ( .A(y[645]), .B(x[132]), .Z(n1278) );
  NAND U1553 ( .A(n1278), .B(n760), .Z(n735) );
  NAND U1554 ( .A(n733), .B(n732), .Z(n734) );
  AND U1555 ( .A(n735), .B(n734), .Z(n757) );
  AND U1556 ( .A(y[643]), .B(x[132]), .Z(n932) );
  NAND U1557 ( .A(x[130]), .B(y[645]), .Z(n736) );
  XNOR U1558 ( .A(n932), .B(n736), .Z(n771) );
  XOR U1559 ( .A(n771), .B(n770), .Z(n755) );
  AND U1560 ( .A(y[647]), .B(x[128]), .Z(n738) );
  NAND U1561 ( .A(y[640]), .B(x[135]), .Z(n737) );
  XNOR U1562 ( .A(n738), .B(n737), .Z(n776) );
  AND U1563 ( .A(n739), .B(o[6]), .Z(n775) );
  XNOR U1564 ( .A(n776), .B(n775), .Z(n754) );
  XNOR U1565 ( .A(n755), .B(n754), .Z(n756) );
  XOR U1566 ( .A(n757), .B(n756), .Z(n790) );
  XOR U1567 ( .A(n791), .B(n790), .Z(n792) );
  XOR U1568 ( .A(n793), .B(n792), .Z(n789) );
  NANDN U1569 ( .A(n741), .B(n740), .Z(n745) );
  NAND U1570 ( .A(n743), .B(n742), .Z(n744) );
  NAND U1571 ( .A(n745), .B(n744), .Z(n788) );
  NANDN U1572 ( .A(n746), .B(n747), .Z(n752) );
  NOR U1573 ( .A(n748), .B(n747), .Z(n750) );
  OR U1574 ( .A(n750), .B(n749), .Z(n751) );
  AND U1575 ( .A(n752), .B(n751), .Z(n787) );
  XOR U1576 ( .A(n788), .B(n787), .Z(n753) );
  XNOR U1577 ( .A(n789), .B(n753), .Z(N40) );
  NANDN U1578 ( .A(n755), .B(n754), .Z(n759) );
  NAND U1579 ( .A(n757), .B(n756), .Z(n758) );
  AND U1580 ( .A(n759), .B(n758), .Z(n843) );
  AND U1581 ( .A(y[646]), .B(x[133]), .Z(n761) );
  NAND U1582 ( .A(n761), .B(n760), .Z(n765) );
  NAND U1583 ( .A(n763), .B(n762), .Z(n764) );
  NAND U1584 ( .A(n765), .B(n764), .Z(n841) );
  AND U1585 ( .A(y[643]), .B(x[133]), .Z(n1378) );
  NAND U1586 ( .A(y[647]), .B(x[129]), .Z(n766) );
  XNOR U1587 ( .A(n1378), .B(n766), .Z(n822) );
  ANDN U1588 ( .B(o[7]), .A(n767), .Z(n821) );
  XOR U1589 ( .A(n822), .B(n821), .Z(n827) );
  NAND U1590 ( .A(y[645]), .B(x[131]), .Z(n1629) );
  AND U1591 ( .A(x[130]), .B(y[646]), .Z(n1700) );
  NAND U1592 ( .A(x[134]), .B(y[642]), .Z(n768) );
  XNOR U1593 ( .A(n1700), .B(n768), .Z(n831) );
  XNOR U1594 ( .A(n1476), .B(n831), .Z(n825) );
  XOR U1595 ( .A(n1629), .B(n825), .Z(n826) );
  XOR U1596 ( .A(n827), .B(n826), .Z(n840) );
  XOR U1597 ( .A(n841), .B(n840), .Z(n842) );
  XOR U1598 ( .A(n843), .B(n842), .Z(n800) );
  NAND U1599 ( .A(n1278), .B(n769), .Z(n773) );
  NAND U1600 ( .A(n771), .B(n770), .Z(n772) );
  NAND U1601 ( .A(n773), .B(n772), .Z(n836) );
  AND U1602 ( .A(x[135]), .B(y[647]), .Z(n774) );
  NAND U1603 ( .A(n1273), .B(n774), .Z(n778) );
  NAND U1604 ( .A(n776), .B(n775), .Z(n777) );
  NAND U1605 ( .A(n778), .B(n777), .Z(n834) );
  AND U1606 ( .A(y[648]), .B(x[128]), .Z(n780) );
  NAND U1607 ( .A(y[640]), .B(x[136]), .Z(n779) );
  XNOR U1608 ( .A(n780), .B(n779), .Z(n812) );
  NAND U1609 ( .A(x[135]), .B(y[641]), .Z(n817) );
  XNOR U1610 ( .A(o[8]), .B(n817), .Z(n811) );
  XOR U1611 ( .A(n812), .B(n811), .Z(n835) );
  XNOR U1612 ( .A(n834), .B(n835), .Z(n837) );
  XOR U1613 ( .A(n836), .B(n837), .Z(n798) );
  NANDN U1614 ( .A(n782), .B(n781), .Z(n786) );
  NANDN U1615 ( .A(n784), .B(n783), .Z(n785) );
  NAND U1616 ( .A(n786), .B(n785), .Z(n797) );
  XOR U1617 ( .A(n798), .B(n797), .Z(n799) );
  XNOR U1618 ( .A(n800), .B(n799), .Z(n806) );
  NAND U1619 ( .A(n791), .B(n790), .Z(n795) );
  NAND U1620 ( .A(n793), .B(n792), .Z(n794) );
  AND U1621 ( .A(n795), .B(n794), .Z(n804) );
  IV U1622 ( .A(n804), .Z(n803) );
  XOR U1623 ( .A(n805), .B(n803), .Z(n796) );
  XNOR U1624 ( .A(n806), .B(n796), .Z(N41) );
  NAND U1625 ( .A(n798), .B(n797), .Z(n802) );
  NANDN U1626 ( .A(n800), .B(n799), .Z(n801) );
  NAND U1627 ( .A(n802), .B(n801), .Z(n855) );
  IV U1628 ( .A(n855), .Z(n853) );
  OR U1629 ( .A(n805), .B(n803), .Z(n809) );
  ANDN U1630 ( .B(n805), .A(n804), .Z(n807) );
  OR U1631 ( .A(n807), .B(n806), .Z(n808) );
  AND U1632 ( .A(n809), .B(n808), .Z(n854) );
  AND U1633 ( .A(x[136]), .B(y[648]), .Z(n810) );
  NAND U1634 ( .A(n810), .B(n1273), .Z(n814) );
  NAND U1635 ( .A(n812), .B(n811), .Z(n813) );
  AND U1636 ( .A(n814), .B(n813), .Z(n895) );
  AND U1637 ( .A(x[133]), .B(y[644]), .Z(n816) );
  NAND U1638 ( .A(y[642]), .B(x[135]), .Z(n815) );
  XNOR U1639 ( .A(n816), .B(n815), .Z(n869) );
  ANDN U1640 ( .B(o[8]), .A(n817), .Z(n868) );
  XOR U1641 ( .A(n869), .B(n868), .Z(n893) );
  AND U1642 ( .A(x[137]), .B(y[640]), .Z(n819) );
  NAND U1643 ( .A(x[128]), .B(y[649]), .Z(n818) );
  XNOR U1644 ( .A(n819), .B(n818), .Z(n875) );
  NAND U1645 ( .A(y[641]), .B(x[136]), .Z(n884) );
  XNOR U1646 ( .A(n875), .B(n874), .Z(n892) );
  XNOR U1647 ( .A(n893), .B(n892), .Z(n894) );
  XOR U1648 ( .A(n895), .B(n894), .Z(n889) );
  AND U1649 ( .A(y[648]), .B(x[129]), .Z(n1616) );
  NAND U1650 ( .A(y[643]), .B(x[134]), .Z(n820) );
  XNOR U1651 ( .A(n1616), .B(n820), .Z(n879) );
  XOR U1652 ( .A(n1278), .B(n879), .Z(n899) );
  NAND U1653 ( .A(x[130]), .B(y[647]), .Z(n1525) );
  NAND U1654 ( .A(y[646]), .B(x[131]), .Z(n1231) );
  XOR U1655 ( .A(n1525), .B(n1231), .Z(n898) );
  XOR U1656 ( .A(n899), .B(n898), .Z(n887) );
  NAND U1657 ( .A(x[133]), .B(y[647]), .Z(n1060) );
  NANDN U1658 ( .A(n1060), .B(n878), .Z(n824) );
  NAND U1659 ( .A(n822), .B(n821), .Z(n823) );
  NAND U1660 ( .A(n824), .B(n823), .Z(n886) );
  XOR U1661 ( .A(n887), .B(n886), .Z(n888) );
  XOR U1662 ( .A(n889), .B(n888), .Z(n862) );
  NAND U1663 ( .A(n1629), .B(n825), .Z(n829) );
  NANDN U1664 ( .A(n827), .B(n826), .Z(n828) );
  AND U1665 ( .A(n829), .B(n828), .Z(n861) );
  AND U1666 ( .A(y[642]), .B(x[130]), .Z(n830) );
  NAND U1667 ( .A(n1014), .B(n830), .Z(n833) );
  NAND U1668 ( .A(n1476), .B(n831), .Z(n832) );
  AND U1669 ( .A(n833), .B(n832), .Z(n860) );
  XOR U1670 ( .A(n862), .B(n863), .Z(n850) );
  NAND U1671 ( .A(n835), .B(n834), .Z(n839) );
  NANDN U1672 ( .A(n837), .B(n836), .Z(n838) );
  NAND U1673 ( .A(n839), .B(n838), .Z(n848) );
  NAND U1674 ( .A(n841), .B(n840), .Z(n845) );
  NAND U1675 ( .A(n843), .B(n842), .Z(n844) );
  NAND U1676 ( .A(n845), .B(n844), .Z(n847) );
  XOR U1677 ( .A(n848), .B(n847), .Z(n849) );
  XNOR U1678 ( .A(n850), .B(n849), .Z(n856) );
  XNOR U1679 ( .A(n854), .B(n856), .Z(n846) );
  XOR U1680 ( .A(n853), .B(n846), .Z(N42) );
  NAND U1681 ( .A(n848), .B(n847), .Z(n852) );
  NANDN U1682 ( .A(n850), .B(n849), .Z(n851) );
  AND U1683 ( .A(n852), .B(n851), .Z(n903) );
  NANDN U1684 ( .A(n853), .B(n854), .Z(n859) );
  NOR U1685 ( .A(n855), .B(n854), .Z(n857) );
  OR U1686 ( .A(n857), .B(n856), .Z(n858) );
  AND U1687 ( .A(n859), .B(n858), .Z(n902) );
  XNOR U1688 ( .A(n903), .B(n902), .Z(n905) );
  NANDN U1689 ( .A(n861), .B(n860), .Z(n865) );
  NAND U1690 ( .A(n863), .B(n862), .Z(n864) );
  AND U1691 ( .A(n865), .B(n864), .Z(n911) );
  AND U1692 ( .A(x[135]), .B(y[644]), .Z(n867) );
  AND U1693 ( .A(y[642]), .B(x[133]), .Z(n866) );
  NAND U1694 ( .A(n867), .B(n866), .Z(n871) );
  NAND U1695 ( .A(n869), .B(n868), .Z(n870) );
  AND U1696 ( .A(n871), .B(n870), .Z(n963) );
  AND U1697 ( .A(x[132]), .B(y[646]), .Z(n873) );
  NAND U1698 ( .A(y[643]), .B(x[135]), .Z(n872) );
  XNOR U1699 ( .A(n873), .B(n872), .Z(n934) );
  NAND U1700 ( .A(y[644]), .B(x[134]), .Z(n935) );
  AND U1701 ( .A(y[642]), .B(x[136]), .Z(n1127) );
  NAND U1702 ( .A(y[641]), .B(x[137]), .Z(n944) );
  XNOR U1703 ( .A(o[10]), .B(n944), .Z(n955) );
  XOR U1704 ( .A(n1127), .B(n955), .Z(n957) );
  XNOR U1705 ( .A(n957), .B(n956), .Z(n960) );
  XOR U1706 ( .A(n963), .B(n962), .Z(n923) );
  AND U1707 ( .A(y[649]), .B(x[137]), .Z(n1485) );
  NAND U1708 ( .A(n1485), .B(n1273), .Z(n877) );
  NAND U1709 ( .A(n875), .B(n874), .Z(n876) );
  AND U1710 ( .A(n877), .B(n876), .Z(n921) );
  AND U1711 ( .A(x[134]), .B(y[648]), .Z(n1163) );
  NAND U1712 ( .A(n1163), .B(n878), .Z(n881) );
  NAND U1713 ( .A(n1278), .B(n879), .Z(n880) );
  AND U1714 ( .A(n881), .B(n880), .Z(n929) );
  AND U1715 ( .A(x[128]), .B(y[650]), .Z(n883) );
  NAND U1716 ( .A(y[640]), .B(x[138]), .Z(n882) );
  XNOR U1717 ( .A(n883), .B(n882), .Z(n939) );
  ANDN U1718 ( .B(o[9]), .A(n884), .Z(n938) );
  XOR U1719 ( .A(n939), .B(n938), .Z(n927) );
  AND U1720 ( .A(y[647]), .B(x[131]), .Z(n1851) );
  NAND U1721 ( .A(x[129]), .B(y[649]), .Z(n885) );
  XNOR U1722 ( .A(n1851), .B(n885), .Z(n951) );
  NAND U1723 ( .A(x[130]), .B(y[648]), .Z(n952) );
  XOR U1724 ( .A(n927), .B(n926), .Z(n928) );
  XNOR U1725 ( .A(n921), .B(n920), .Z(n922) );
  XOR U1726 ( .A(n923), .B(n922), .Z(n909) );
  NAND U1727 ( .A(n887), .B(n886), .Z(n891) );
  NANDN U1728 ( .A(n889), .B(n888), .Z(n890) );
  AND U1729 ( .A(n891), .B(n890), .Z(n917) );
  NANDN U1730 ( .A(n893), .B(n892), .Z(n897) );
  NAND U1731 ( .A(n895), .B(n894), .Z(n896) );
  AND U1732 ( .A(n897), .B(n896), .Z(n914) );
  AND U1733 ( .A(n1525), .B(n1231), .Z(n901) );
  NANDN U1734 ( .A(n899), .B(n898), .Z(n900) );
  NANDN U1735 ( .A(n901), .B(n900), .Z(n915) );
  XNOR U1736 ( .A(n914), .B(n915), .Z(n916) );
  XOR U1737 ( .A(n917), .B(n916), .Z(n908) );
  XOR U1738 ( .A(n909), .B(n908), .Z(n910) );
  XOR U1739 ( .A(n911), .B(n910), .Z(n904) );
  XOR U1740 ( .A(n905), .B(n904), .Z(N43) );
  NANDN U1741 ( .A(n903), .B(n902), .Z(n907) );
  NAND U1742 ( .A(n905), .B(n904), .Z(n906) );
  AND U1743 ( .A(n907), .B(n906), .Z(n1029) );
  NAND U1744 ( .A(n909), .B(n908), .Z(n913) );
  NANDN U1745 ( .A(n911), .B(n910), .Z(n912) );
  NAND U1746 ( .A(n913), .B(n912), .Z(n1028) );
  NANDN U1747 ( .A(n915), .B(n914), .Z(n919) );
  NANDN U1748 ( .A(n917), .B(n916), .Z(n918) );
  AND U1749 ( .A(n919), .B(n918), .Z(n1025) );
  NANDN U1750 ( .A(n921), .B(n920), .Z(n925) );
  NANDN U1751 ( .A(n923), .B(n922), .Z(n924) );
  AND U1752 ( .A(n925), .B(n924), .Z(n1023) );
  NAND U1753 ( .A(n927), .B(n926), .Z(n931) );
  NANDN U1754 ( .A(n929), .B(n928), .Z(n930) );
  NAND U1755 ( .A(n931), .B(n930), .Z(n981) );
  AND U1756 ( .A(x[135]), .B(y[646]), .Z(n933) );
  NAND U1757 ( .A(n933), .B(n932), .Z(n937) );
  NANDN U1758 ( .A(n935), .B(n934), .Z(n936) );
  AND U1759 ( .A(n937), .B(n936), .Z(n979) );
  AND U1760 ( .A(x[138]), .B(y[650]), .Z(n1706) );
  NAND U1761 ( .A(n1706), .B(n1273), .Z(n941) );
  NAND U1762 ( .A(n939), .B(n938), .Z(n940) );
  AND U1763 ( .A(n941), .B(n940), .Z(n975) );
  AND U1764 ( .A(y[640]), .B(x[139]), .Z(n943) );
  NAND U1765 ( .A(x[128]), .B(y[651]), .Z(n942) );
  XNOR U1766 ( .A(n943), .B(n942), .Z(n1006) );
  ANDN U1767 ( .B(o[10]), .A(n944), .Z(n1005) );
  XOR U1768 ( .A(n1006), .B(n1005), .Z(n973) );
  AND U1769 ( .A(x[129]), .B(y[650]), .Z(n946) );
  NAND U1770 ( .A(x[134]), .B(y[645]), .Z(n945) );
  XNOR U1771 ( .A(n946), .B(n945), .Z(n996) );
  NAND U1772 ( .A(x[138]), .B(y[641]), .Z(n1015) );
  XNOR U1773 ( .A(o[11]), .B(n1015), .Z(n995) );
  XOR U1774 ( .A(n996), .B(n995), .Z(n972) );
  XOR U1775 ( .A(n973), .B(n972), .Z(n974) );
  XNOR U1776 ( .A(n981), .B(n980), .Z(n1018) );
  AND U1777 ( .A(x[131]), .B(y[648]), .Z(n1992) );
  AND U1778 ( .A(x[130]), .B(y[649]), .Z(n948) );
  NAND U1779 ( .A(x[133]), .B(y[646]), .Z(n947) );
  XNOR U1780 ( .A(n948), .B(n947), .Z(n991) );
  AND U1781 ( .A(x[132]), .B(y[647]), .Z(n990) );
  XNOR U1782 ( .A(n991), .B(n990), .Z(n967) );
  XNOR U1783 ( .A(n1992), .B(n967), .Z(n969) );
  AND U1784 ( .A(x[137]), .B(y[642]), .Z(n950) );
  NAND U1785 ( .A(y[644]), .B(x[135]), .Z(n949) );
  XNOR U1786 ( .A(n950), .B(n949), .Z(n1010) );
  AND U1787 ( .A(x[136]), .B(y[643]), .Z(n1009) );
  XNOR U1788 ( .A(n1010), .B(n1009), .Z(n968) );
  XOR U1789 ( .A(n969), .B(n968), .Z(n987) );
  NAND U1790 ( .A(y[649]), .B(x[131]), .Z(n1051) );
  AND U1791 ( .A(x[129]), .B(y[647]), .Z(n1268) );
  NANDN U1792 ( .A(n1051), .B(n1268), .Z(n954) );
  NANDN U1793 ( .A(n952), .B(n951), .Z(n953) );
  AND U1794 ( .A(n954), .B(n953), .Z(n985) );
  NAND U1795 ( .A(n1127), .B(n955), .Z(n959) );
  NAND U1796 ( .A(n957), .B(n956), .Z(n958) );
  NAND U1797 ( .A(n959), .B(n958), .Z(n984) );
  NANDN U1798 ( .A(n961), .B(n960), .Z(n965) );
  NAND U1799 ( .A(n963), .B(n962), .Z(n964) );
  NAND U1800 ( .A(n965), .B(n964), .Z(n1016) );
  XOR U1801 ( .A(n1018), .B(n1019), .Z(n1022) );
  XNOR U1802 ( .A(n1023), .B(n1022), .Z(n1024) );
  XNOR U1803 ( .A(n1025), .B(n1024), .Z(n1030) );
  XOR U1804 ( .A(n1028), .B(n1030), .Z(n966) );
  XOR U1805 ( .A(n1029), .B(n966), .Z(N44) );
  NANDN U1806 ( .A(n1992), .B(n967), .Z(n971) );
  NAND U1807 ( .A(n969), .B(n968), .Z(n970) );
  AND U1808 ( .A(n971), .B(n970), .Z(n1033) );
  NAND U1809 ( .A(n973), .B(n972), .Z(n977) );
  NANDN U1810 ( .A(n975), .B(n974), .Z(n976) );
  AND U1811 ( .A(n977), .B(n976), .Z(n1032) );
  NANDN U1812 ( .A(n979), .B(n978), .Z(n983) );
  NAND U1813 ( .A(n981), .B(n980), .Z(n982) );
  NAND U1814 ( .A(n983), .B(n982), .Z(n1035) );
  NANDN U1815 ( .A(n985), .B(n984), .Z(n989) );
  NANDN U1816 ( .A(n987), .B(n986), .Z(n988) );
  AND U1817 ( .A(n989), .B(n988), .Z(n1093) );
  AND U1818 ( .A(y[649]), .B(x[133]), .Z(n1516) );
  NAND U1819 ( .A(n1700), .B(n1516), .Z(n993) );
  NAND U1820 ( .A(n991), .B(n990), .Z(n992) );
  AND U1821 ( .A(n993), .B(n992), .Z(n1039) );
  AND U1822 ( .A(x[134]), .B(y[650]), .Z(n1285) );
  NAND U1823 ( .A(n1285), .B(n994), .Z(n998) );
  NAND U1824 ( .A(n996), .B(n995), .Z(n997) );
  NAND U1825 ( .A(n998), .B(n997), .Z(n1038) );
  XNOR U1826 ( .A(n1039), .B(n1038), .Z(n1041) );
  AND U1827 ( .A(x[137]), .B(y[643]), .Z(n1695) );
  AND U1828 ( .A(y[648]), .B(x[132]), .Z(n1000) );
  NAND U1829 ( .A(y[642]), .B(x[138]), .Z(n999) );
  XOR U1830 ( .A(n1000), .B(n999), .Z(n1083) );
  XNOR U1831 ( .A(n1695), .B(n1083), .Z(n1061) );
  NAND U1832 ( .A(x[135]), .B(y[645]), .Z(n1059) );
  XOR U1833 ( .A(n1060), .B(n1059), .Z(n1062) );
  AND U1834 ( .A(x[128]), .B(y[652]), .Z(n1002) );
  NAND U1835 ( .A(y[640]), .B(x[140]), .Z(n1001) );
  XNOR U1836 ( .A(n1002), .B(n1001), .Z(n1076) );
  NAND U1837 ( .A(x[139]), .B(y[641]), .Z(n1056) );
  XNOR U1838 ( .A(o[12]), .B(n1056), .Z(n1075) );
  XOR U1839 ( .A(n1076), .B(n1075), .Z(n1045) );
  AND U1840 ( .A(x[130]), .B(y[650]), .Z(n1004) );
  NAND U1841 ( .A(y[644]), .B(x[136]), .Z(n1003) );
  XNOR U1842 ( .A(n1004), .B(n1003), .Z(n1050) );
  XOR U1843 ( .A(n1045), .B(n1044), .Z(n1047) );
  XOR U1844 ( .A(n1046), .B(n1047), .Z(n1040) );
  XOR U1845 ( .A(n1041), .B(n1040), .Z(n1091) );
  AND U1846 ( .A(y[651]), .B(x[139]), .Z(n2116) );
  NAND U1847 ( .A(n2116), .B(n1273), .Z(n1008) );
  NAND U1848 ( .A(n1006), .B(n1005), .Z(n1007) );
  AND U1849 ( .A(n1008), .B(n1007), .Z(n1068) );
  AND U1850 ( .A(x[135]), .B(y[642]), .Z(n1207) );
  AND U1851 ( .A(y[644]), .B(x[137]), .Z(n1058) );
  NAND U1852 ( .A(n1207), .B(n1058), .Z(n1012) );
  NAND U1853 ( .A(n1010), .B(n1009), .Z(n1011) );
  AND U1854 ( .A(n1012), .B(n1011), .Z(n1066) );
  NAND U1855 ( .A(x[129]), .B(y[651]), .Z(n1013) );
  XNOR U1856 ( .A(n1014), .B(n1013), .Z(n1072) );
  ANDN U1857 ( .B(o[11]), .A(n1015), .Z(n1071) );
  XOR U1858 ( .A(n1072), .B(n1071), .Z(n1065) );
  XNOR U1859 ( .A(n1066), .B(n1065), .Z(n1067) );
  XNOR U1860 ( .A(n1068), .B(n1067), .Z(n1090) );
  XOR U1861 ( .A(n1091), .B(n1090), .Z(n1092) );
  NANDN U1862 ( .A(n1017), .B(n1016), .Z(n1021) );
  NANDN U1863 ( .A(n1019), .B(n1018), .Z(n1020) );
  NAND U1864 ( .A(n1021), .B(n1020), .Z(n1099) );
  XNOR U1865 ( .A(n1101), .B(n1102), .Z(n1098) );
  NANDN U1866 ( .A(n1023), .B(n1022), .Z(n1027) );
  NANDN U1867 ( .A(n1025), .B(n1024), .Z(n1026) );
  NAND U1868 ( .A(n1027), .B(n1026), .Z(n1097) );
  XOR U1869 ( .A(n1097), .B(n1096), .Z(n1031) );
  XNOR U1870 ( .A(n1098), .B(n1031), .Z(N45) );
  NANDN U1871 ( .A(n1033), .B(n1032), .Z(n1037) );
  NANDN U1872 ( .A(n1035), .B(n1034), .Z(n1036) );
  AND U1873 ( .A(n1037), .B(n1036), .Z(n1112) );
  NANDN U1874 ( .A(n1039), .B(n1038), .Z(n1043) );
  NAND U1875 ( .A(n1041), .B(n1040), .Z(n1042) );
  AND U1876 ( .A(n1043), .B(n1042), .Z(n1171) );
  NAND U1877 ( .A(n1045), .B(n1044), .Z(n1049) );
  NAND U1878 ( .A(n1047), .B(n1046), .Z(n1048) );
  NAND U1879 ( .A(n1049), .B(n1048), .Z(n1178) );
  AND U1880 ( .A(x[136]), .B(y[650]), .Z(n2386) );
  AND U1881 ( .A(y[644]), .B(x[130]), .Z(n1216) );
  NAND U1882 ( .A(n2386), .B(n1216), .Z(n1053) );
  NANDN U1883 ( .A(n1051), .B(n1050), .Z(n1052) );
  AND U1884 ( .A(n1053), .B(n1052), .Z(n1143) );
  AND U1885 ( .A(x[129]), .B(y[652]), .Z(n1055) );
  NAND U1886 ( .A(y[646]), .B(x[135]), .Z(n1054) );
  XNOR U1887 ( .A(n1055), .B(n1054), .Z(n1134) );
  ANDN U1888 ( .B(o[12]), .A(n1056), .Z(n1133) );
  XOR U1889 ( .A(n1134), .B(n1133), .Z(n1141) );
  AND U1890 ( .A(x[134]), .B(y[647]), .Z(n2154) );
  NAND U1891 ( .A(x[130]), .B(y[651]), .Z(n1057) );
  XOR U1892 ( .A(n1058), .B(n1057), .Z(n1147) );
  XNOR U1893 ( .A(n2154), .B(n1147), .Z(n1140) );
  XOR U1894 ( .A(n1141), .B(n1140), .Z(n1142) );
  XNOR U1895 ( .A(n1143), .B(n1142), .Z(n1177) );
  NAND U1896 ( .A(n1060), .B(n1059), .Z(n1064) );
  ANDN U1897 ( .B(n1062), .A(n1061), .Z(n1063) );
  ANDN U1898 ( .B(n1064), .A(n1063), .Z(n1176) );
  XOR U1899 ( .A(n1177), .B(n1176), .Z(n1179) );
  XOR U1900 ( .A(n1178), .B(n1179), .Z(n1170) );
  XNOR U1901 ( .A(n1171), .B(n1170), .Z(n1173) );
  NANDN U1902 ( .A(n1066), .B(n1065), .Z(n1070) );
  NANDN U1903 ( .A(n1068), .B(n1067), .Z(n1069) );
  AND U1904 ( .A(n1070), .B(n1069), .Z(n1118) );
  AND U1905 ( .A(y[651]), .B(x[134]), .Z(n1437) );
  IV U1906 ( .A(n1437), .Z(n1518) );
  NANDN U1907 ( .A(n1518), .B(n1132), .Z(n1074) );
  NAND U1908 ( .A(n1072), .B(n1071), .Z(n1073) );
  AND U1909 ( .A(n1074), .B(n1073), .Z(n1124) );
  AND U1910 ( .A(x[140]), .B(y[652]), .Z(n2392) );
  NAND U1911 ( .A(n2392), .B(n1273), .Z(n1078) );
  NAND U1912 ( .A(n1076), .B(n1075), .Z(n1077) );
  AND U1913 ( .A(n1078), .B(n1077), .Z(n1122) );
  AND U1914 ( .A(x[138]), .B(y[643]), .Z(n2004) );
  AND U1915 ( .A(y[645]), .B(x[136]), .Z(n1080) );
  NAND U1916 ( .A(y[642]), .B(x[139]), .Z(n1079) );
  XOR U1917 ( .A(n1080), .B(n1079), .Z(n1129) );
  XNOR U1918 ( .A(n2004), .B(n1129), .Z(n1121) );
  XNOR U1919 ( .A(n1122), .B(n1121), .Z(n1123) );
  XNOR U1920 ( .A(n1124), .B(n1123), .Z(n1116) );
  AND U1921 ( .A(x[138]), .B(y[648]), .Z(n1082) );
  AND U1922 ( .A(y[642]), .B(x[132]), .Z(n1081) );
  NAND U1923 ( .A(n1082), .B(n1081), .Z(n1085) );
  NANDN U1924 ( .A(n1083), .B(n1695), .Z(n1084) );
  AND U1925 ( .A(n1085), .B(n1084), .Z(n1167) );
  AND U1926 ( .A(y[640]), .B(x[141]), .Z(n1087) );
  NAND U1927 ( .A(x[128]), .B(y[653]), .Z(n1086) );
  XNOR U1928 ( .A(n1087), .B(n1086), .Z(n1159) );
  NAND U1929 ( .A(x[140]), .B(y[641]), .Z(n1152) );
  XNOR U1930 ( .A(o[13]), .B(n1152), .Z(n1158) );
  XOR U1931 ( .A(n1159), .B(n1158), .Z(n1165) );
  AND U1932 ( .A(y[648]), .B(x[133]), .Z(n1089) );
  NAND U1933 ( .A(x[131]), .B(y[650]), .Z(n1088) );
  XNOR U1934 ( .A(n1089), .B(n1088), .Z(n1154) );
  NAND U1935 ( .A(x[132]), .B(y[649]), .Z(n1155) );
  XNOR U1936 ( .A(n1154), .B(n1155), .Z(n1164) );
  XOR U1937 ( .A(n1165), .B(n1164), .Z(n1166) );
  XNOR U1938 ( .A(n1167), .B(n1166), .Z(n1115) );
  XOR U1939 ( .A(n1116), .B(n1115), .Z(n1117) );
  XNOR U1940 ( .A(n1118), .B(n1117), .Z(n1172) );
  XOR U1941 ( .A(n1173), .B(n1172), .Z(n1110) );
  NAND U1942 ( .A(n1091), .B(n1090), .Z(n1095) );
  NANDN U1943 ( .A(n1093), .B(n1092), .Z(n1094) );
  AND U1944 ( .A(n1095), .B(n1094), .Z(n1109) );
  XOR U1945 ( .A(n1112), .B(n1111), .Z(n1108) );
  NANDN U1946 ( .A(n1100), .B(n1099), .Z(n1104) );
  NANDN U1947 ( .A(n1102), .B(n1101), .Z(n1103) );
  NAND U1948 ( .A(n1104), .B(n1103), .Z(n1106) );
  XNOR U1949 ( .A(n1107), .B(n1106), .Z(n1105) );
  XNOR U1950 ( .A(n1108), .B(n1105), .Z(N46) );
  NANDN U1951 ( .A(n1110), .B(n1109), .Z(n1114) );
  NANDN U1952 ( .A(n1112), .B(n1111), .Z(n1113) );
  NAND U1953 ( .A(n1114), .B(n1113), .Z(n1264) );
  NAND U1954 ( .A(n1116), .B(n1115), .Z(n1120) );
  NANDN U1955 ( .A(n1118), .B(n1117), .Z(n1119) );
  AND U1956 ( .A(n1120), .B(n1119), .Z(n1186) );
  NANDN U1957 ( .A(n1122), .B(n1121), .Z(n1126) );
  NANDN U1958 ( .A(n1124), .B(n1123), .Z(n1125) );
  AND U1959 ( .A(n1126), .B(n1125), .Z(n1192) );
  AND U1960 ( .A(x[139]), .B(y[645]), .Z(n1128) );
  NAND U1961 ( .A(n1128), .B(n1127), .Z(n1131) );
  NANDN U1962 ( .A(n1129), .B(n2004), .Z(n1130) );
  AND U1963 ( .A(n1131), .B(n1130), .Z(n1247) );
  NAND U1964 ( .A(x[135]), .B(y[652]), .Z(n1710) );
  NANDN U1965 ( .A(n1710), .B(n1132), .Z(n1136) );
  NAND U1966 ( .A(n1134), .B(n1133), .Z(n1135) );
  NAND U1967 ( .A(n1136), .B(n1135), .Z(n1246) );
  XNOR U1968 ( .A(n1247), .B(n1246), .Z(n1249) );
  AND U1969 ( .A(x[132]), .B(y[650]), .Z(n1638) );
  AND U1970 ( .A(y[646]), .B(x[136]), .Z(n1138) );
  NAND U1971 ( .A(x[131]), .B(y[651]), .Z(n1137) );
  XOR U1972 ( .A(n1138), .B(n1137), .Z(n1232) );
  XNOR U1973 ( .A(n1516), .B(n1232), .Z(n1241) );
  XOR U1974 ( .A(n1638), .B(n1241), .Z(n1243) );
  AND U1975 ( .A(y[645]), .B(x[137]), .Z(n1822) );
  AND U1976 ( .A(x[130]), .B(y[652]), .Z(n1139) );
  AND U1977 ( .A(y[644]), .B(x[138]), .Z(n1846) );
  XOR U1978 ( .A(n1139), .B(n1846), .Z(n1217) );
  XOR U1979 ( .A(n1822), .B(n1217), .Z(n1242) );
  XOR U1980 ( .A(n1243), .B(n1242), .Z(n1248) );
  XOR U1981 ( .A(n1249), .B(n1248), .Z(n1190) );
  NAND U1982 ( .A(n1141), .B(n1140), .Z(n1145) );
  NANDN U1983 ( .A(n1143), .B(n1142), .Z(n1144) );
  AND U1984 ( .A(n1145), .B(n1144), .Z(n1189) );
  XNOR U1985 ( .A(n1190), .B(n1189), .Z(n1191) );
  XOR U1986 ( .A(n1192), .B(n1191), .Z(n1184) );
  AND U1987 ( .A(y[651]), .B(x[137]), .Z(n1146) );
  NAND U1988 ( .A(n1146), .B(n1216), .Z(n1149) );
  NANDN U1989 ( .A(n1147), .B(n2154), .Z(n1148) );
  AND U1990 ( .A(n1149), .B(n1148), .Z(n1204) );
  AND U1991 ( .A(y[640]), .B(x[142]), .Z(n1151) );
  NAND U1992 ( .A(x[128]), .B(y[654]), .Z(n1150) );
  XNOR U1993 ( .A(n1151), .B(n1150), .Z(n1227) );
  ANDN U1994 ( .B(o[13]), .A(n1152), .Z(n1226) );
  XOR U1995 ( .A(n1227), .B(n1226), .Z(n1202) );
  AND U1996 ( .A(y[642]), .B(x[140]), .Z(n1812) );
  NAND U1997 ( .A(y[647]), .B(x[135]), .Z(n1153) );
  XNOR U1998 ( .A(n1812), .B(n1153), .Z(n1209) );
  NAND U1999 ( .A(y[641]), .B(x[141]), .Z(n1215) );
  XNOR U2000 ( .A(o[14]), .B(n1215), .Z(n1208) );
  XOR U2001 ( .A(n1209), .B(n1208), .Z(n1201) );
  XOR U2002 ( .A(n1202), .B(n1201), .Z(n1203) );
  XOR U2003 ( .A(n1204), .B(n1203), .Z(n1253) );
  NAND U2004 ( .A(y[650]), .B(x[133]), .Z(n1286) );
  NANDN U2005 ( .A(n1286), .B(n1992), .Z(n1157) );
  NANDN U2006 ( .A(n1155), .B(n1154), .Z(n1156) );
  AND U2007 ( .A(n1157), .B(n1156), .Z(n1198) );
  AND U2008 ( .A(y[653]), .B(x[141]), .Z(n2739) );
  NAND U2009 ( .A(n2739), .B(n1273), .Z(n1161) );
  NAND U2010 ( .A(n1159), .B(n1158), .Z(n1160) );
  AND U2011 ( .A(n1161), .B(n1160), .Z(n1196) );
  NAND U2012 ( .A(y[643]), .B(x[139]), .Z(n1162) );
  XNOR U2013 ( .A(n1163), .B(n1162), .Z(n1222) );
  NAND U2014 ( .A(y[653]), .B(x[129]), .Z(n1223) );
  XNOR U2015 ( .A(n1222), .B(n1223), .Z(n1195) );
  XNOR U2016 ( .A(n1196), .B(n1195), .Z(n1197) );
  XOR U2017 ( .A(n1198), .B(n1197), .Z(n1252) );
  XOR U2018 ( .A(n1253), .B(n1252), .Z(n1255) );
  NAND U2019 ( .A(n1165), .B(n1164), .Z(n1169) );
  NANDN U2020 ( .A(n1167), .B(n1166), .Z(n1168) );
  AND U2021 ( .A(n1169), .B(n1168), .Z(n1254) );
  XNOR U2022 ( .A(n1255), .B(n1254), .Z(n1183) );
  XNOR U2023 ( .A(n1184), .B(n1183), .Z(n1185) );
  XNOR U2024 ( .A(n1186), .B(n1185), .Z(n1261) );
  NANDN U2025 ( .A(n1171), .B(n1170), .Z(n1175) );
  NAND U2026 ( .A(n1173), .B(n1172), .Z(n1174) );
  AND U2027 ( .A(n1175), .B(n1174), .Z(n1259) );
  NAND U2028 ( .A(n1177), .B(n1176), .Z(n1181) );
  NAND U2029 ( .A(n1179), .B(n1178), .Z(n1180) );
  NAND U2030 ( .A(n1181), .B(n1180), .Z(n1258) );
  XNOR U2031 ( .A(n1259), .B(n1258), .Z(n1260) );
  XOR U2032 ( .A(n1261), .B(n1260), .Z(n1266) );
  XOR U2033 ( .A(n1264), .B(n1266), .Z(n1182) );
  XOR U2034 ( .A(n1265), .B(n1182), .Z(N47) );
  NANDN U2035 ( .A(n1184), .B(n1183), .Z(n1188) );
  NANDN U2036 ( .A(n1186), .B(n1185), .Z(n1187) );
  AND U2037 ( .A(n1188), .B(n1187), .Z(n1356) );
  NANDN U2038 ( .A(n1190), .B(n1189), .Z(n1194) );
  NAND U2039 ( .A(n1192), .B(n1191), .Z(n1193) );
  AND U2040 ( .A(n1194), .B(n1193), .Z(n1329) );
  NANDN U2041 ( .A(n1196), .B(n1195), .Z(n1200) );
  NANDN U2042 ( .A(n1198), .B(n1197), .Z(n1199) );
  AND U2043 ( .A(n1200), .B(n1199), .Z(n1335) );
  NAND U2044 ( .A(n1202), .B(n1201), .Z(n1206) );
  NANDN U2045 ( .A(n1204), .B(n1203), .Z(n1205) );
  AND U2046 ( .A(n1206), .B(n1205), .Z(n1333) );
  NAND U2047 ( .A(x[140]), .B(y[647]), .Z(n1702) );
  NANDN U2048 ( .A(n1702), .B(n1207), .Z(n1211) );
  NAND U2049 ( .A(n1209), .B(n1208), .Z(n1210) );
  AND U2050 ( .A(n1211), .B(n1210), .Z(n1309) );
  AND U2051 ( .A(x[141]), .B(y[642]), .Z(n2142) );
  NAND U2052 ( .A(y[644]), .B(x[139]), .Z(n1212) );
  XNOR U2053 ( .A(n2142), .B(n1212), .Z(n1313) );
  AND U2054 ( .A(x[140]), .B(y[643]), .Z(n1312) );
  XOR U2055 ( .A(n1313), .B(n1312), .Z(n1307) );
  AND U2056 ( .A(x[128]), .B(y[655]), .Z(n1214) );
  NAND U2057 ( .A(y[640]), .B(x[143]), .Z(n1213) );
  XNOR U2058 ( .A(n1214), .B(n1213), .Z(n1275) );
  ANDN U2059 ( .B(o[14]), .A(n1215), .Z(n1274) );
  XNOR U2060 ( .A(n1275), .B(n1274), .Z(n1306) );
  XNOR U2061 ( .A(n1307), .B(n1306), .Z(n1308) );
  XOR U2062 ( .A(n1309), .B(n1308), .Z(n1341) );
  NAND U2063 ( .A(x[138]), .B(y[652]), .Z(n2156) );
  NANDN U2064 ( .A(n2156), .B(n1216), .Z(n1219) );
  NAND U2065 ( .A(n1822), .B(n1217), .Z(n1218) );
  AND U2066 ( .A(n1219), .B(n1218), .Z(n1339) );
  AND U2067 ( .A(x[139]), .B(y[648]), .Z(n1221) );
  AND U2068 ( .A(x[134]), .B(y[643]), .Z(n1220) );
  NAND U2069 ( .A(n1221), .B(n1220), .Z(n1225) );
  NANDN U2070 ( .A(n1223), .B(n1222), .Z(n1224) );
  NAND U2071 ( .A(n1225), .B(n1224), .Z(n1338) );
  XNOR U2072 ( .A(n1339), .B(n1338), .Z(n1340) );
  XNOR U2073 ( .A(n1341), .B(n1340), .Z(n1332) );
  XNOR U2074 ( .A(n1333), .B(n1332), .Z(n1334) );
  XOR U2075 ( .A(n1335), .B(n1334), .Z(n1326) );
  AND U2076 ( .A(y[654]), .B(x[142]), .Z(n3003) );
  NAND U2077 ( .A(n3003), .B(n1273), .Z(n1229) );
  NAND U2078 ( .A(n1227), .B(n1226), .Z(n1228) );
  AND U2079 ( .A(n1229), .B(n1228), .Z(n1301) );
  AND U2080 ( .A(y[651]), .B(x[136]), .Z(n1230) );
  NANDN U2081 ( .A(n1231), .B(n1230), .Z(n1234) );
  NANDN U2082 ( .A(n1232), .B(n1516), .Z(n1233) );
  NAND U2083 ( .A(n1234), .B(n1233), .Z(n1300) );
  XNOR U2084 ( .A(n1301), .B(n1300), .Z(n1303) );
  AND U2085 ( .A(y[645]), .B(x[138]), .Z(n1236) );
  NAND U2086 ( .A(x[132]), .B(y[651]), .Z(n1235) );
  XNOR U2087 ( .A(n1236), .B(n1235), .Z(n1281) );
  AND U2088 ( .A(x[135]), .B(y[648]), .Z(n1280) );
  XOR U2089 ( .A(n1281), .B(n1280), .Z(n1288) );
  AND U2090 ( .A(x[134]), .B(y[649]), .Z(n1387) );
  XNOR U2091 ( .A(n1387), .B(n1286), .Z(n1287) );
  XNOR U2092 ( .A(n1288), .B(n1287), .Z(n1323) );
  AND U2093 ( .A(x[137]), .B(y[646]), .Z(n1238) );
  NAND U2094 ( .A(x[130]), .B(y[653]), .Z(n1237) );
  XNOR U2095 ( .A(n1238), .B(n1237), .Z(n1291) );
  NAND U2096 ( .A(y[652]), .B(x[131]), .Z(n1292) );
  XNOR U2097 ( .A(n1291), .B(n1292), .Z(n1321) );
  AND U2098 ( .A(x[129]), .B(y[654]), .Z(n1240) );
  NAND U2099 ( .A(y[647]), .B(x[136]), .Z(n1239) );
  XNOR U2100 ( .A(n1240), .B(n1239), .Z(n1270) );
  NAND U2101 ( .A(y[641]), .B(x[142]), .Z(n1297) );
  XNOR U2102 ( .A(o[15]), .B(n1297), .Z(n1269) );
  XOR U2103 ( .A(n1270), .B(n1269), .Z(n1320) );
  XOR U2104 ( .A(n1321), .B(n1320), .Z(n1322) );
  XOR U2105 ( .A(n1303), .B(n1302), .Z(n1345) );
  NAND U2106 ( .A(n1638), .B(n1241), .Z(n1245) );
  NAND U2107 ( .A(n1243), .B(n1242), .Z(n1244) );
  AND U2108 ( .A(n1245), .B(n1244), .Z(n1344) );
  XNOR U2109 ( .A(n1345), .B(n1344), .Z(n1346) );
  NANDN U2110 ( .A(n1247), .B(n1246), .Z(n1251) );
  NAND U2111 ( .A(n1249), .B(n1248), .Z(n1250) );
  NAND U2112 ( .A(n1251), .B(n1250), .Z(n1347) );
  XNOR U2113 ( .A(n1346), .B(n1347), .Z(n1327) );
  XOR U2114 ( .A(n1326), .B(n1327), .Z(n1328) );
  XOR U2115 ( .A(n1329), .B(n1328), .Z(n1353) );
  NAND U2116 ( .A(n1253), .B(n1252), .Z(n1257) );
  NAND U2117 ( .A(n1255), .B(n1254), .Z(n1256) );
  AND U2118 ( .A(n1257), .B(n1256), .Z(n1354) );
  XOR U2119 ( .A(n1353), .B(n1354), .Z(n1355) );
  XOR U2120 ( .A(n1356), .B(n1355), .Z(n1352) );
  NANDN U2121 ( .A(n1259), .B(n1258), .Z(n1263) );
  NAND U2122 ( .A(n1261), .B(n1260), .Z(n1262) );
  NAND U2123 ( .A(n1263), .B(n1262), .Z(n1351) );
  XOR U2124 ( .A(n1351), .B(n1350), .Z(n1267) );
  XNOR U2125 ( .A(n1352), .B(n1267), .Z(N48) );
  AND U2126 ( .A(x[136]), .B(y[654]), .Z(n2013) );
  NAND U2127 ( .A(n2013), .B(n1268), .Z(n1272) );
  NAND U2128 ( .A(n1270), .B(n1269), .Z(n1271) );
  AND U2129 ( .A(n1272), .B(n1271), .Z(n1417) );
  AND U2130 ( .A(x[143]), .B(y[655]), .Z(n3399) );
  NAND U2131 ( .A(n3399), .B(n1273), .Z(n1277) );
  NAND U2132 ( .A(n1275), .B(n1274), .Z(n1276) );
  NAND U2133 ( .A(n1277), .B(n1276), .Z(n1416) );
  XNOR U2134 ( .A(n1417), .B(n1416), .Z(n1419) );
  AND U2135 ( .A(y[651]), .B(x[138]), .Z(n1279) );
  NAND U2136 ( .A(n1279), .B(n1278), .Z(n1283) );
  NAND U2137 ( .A(n1281), .B(n1280), .Z(n1282) );
  NAND U2138 ( .A(n1283), .B(n1282), .Z(n1374) );
  AND U2139 ( .A(y[656]), .B(x[128]), .Z(n1396) );
  NAND U2140 ( .A(x[144]), .B(y[640]), .Z(n1397) );
  XNOR U2141 ( .A(n1396), .B(n1397), .Z(n1399) );
  NAND U2142 ( .A(y[641]), .B(x[143]), .Z(n1384) );
  XNOR U2143 ( .A(o[16]), .B(n1384), .Z(n1398) );
  XOR U2144 ( .A(n1399), .B(n1398), .Z(n1373) );
  NAND U2145 ( .A(y[649]), .B(x[135]), .Z(n1284) );
  XNOR U2146 ( .A(n1285), .B(n1284), .Z(n1389) );
  AND U2147 ( .A(x[138]), .B(y[646]), .Z(n1388) );
  XOR U2148 ( .A(n1389), .B(n1388), .Z(n1372) );
  XOR U2149 ( .A(n1373), .B(n1372), .Z(n1375) );
  XOR U2150 ( .A(n1374), .B(n1375), .Z(n1418) );
  XOR U2151 ( .A(n1419), .B(n1418), .Z(n1369) );
  NANDN U2152 ( .A(n1387), .B(n1286), .Z(n1290) );
  NANDN U2153 ( .A(n1288), .B(n1287), .Z(n1289) );
  AND U2154 ( .A(n1290), .B(n1289), .Z(n1367) );
  NAND U2155 ( .A(y[653]), .B(x[137]), .Z(n2127) );
  NANDN U2156 ( .A(n2127), .B(n1700), .Z(n1294) );
  NANDN U2157 ( .A(n1292), .B(n1291), .Z(n1293) );
  NAND U2158 ( .A(n1294), .B(n1293), .Z(n1406) );
  AND U2159 ( .A(x[129]), .B(y[655]), .Z(n1296) );
  NAND U2160 ( .A(y[648]), .B(x[136]), .Z(n1295) );
  XNOR U2161 ( .A(n1296), .B(n1295), .Z(n1393) );
  ANDN U2162 ( .B(o[15]), .A(n1297), .Z(n1392) );
  XOR U2163 ( .A(n1393), .B(n1392), .Z(n1405) );
  AND U2164 ( .A(x[142]), .B(y[642]), .Z(n1299) );
  NAND U2165 ( .A(y[645]), .B(x[139]), .Z(n1298) );
  XNOR U2166 ( .A(n1299), .B(n1298), .Z(n1428) );
  NAND U2167 ( .A(x[132]), .B(y[652]), .Z(n1429) );
  XNOR U2168 ( .A(n1428), .B(n1429), .Z(n1404) );
  XOR U2169 ( .A(n1405), .B(n1404), .Z(n1407) );
  XNOR U2170 ( .A(n1406), .B(n1407), .Z(n1366) );
  XNOR U2171 ( .A(n1367), .B(n1366), .Z(n1368) );
  XNOR U2172 ( .A(n1369), .B(n1368), .Z(n1410) );
  NANDN U2173 ( .A(n1301), .B(n1300), .Z(n1305) );
  NAND U2174 ( .A(n1303), .B(n1302), .Z(n1304) );
  NAND U2175 ( .A(n1305), .B(n1304), .Z(n1411) );
  XNOR U2176 ( .A(n1410), .B(n1411), .Z(n1413) );
  NANDN U2177 ( .A(n1307), .B(n1306), .Z(n1311) );
  NAND U2178 ( .A(n1309), .B(n1308), .Z(n1310) );
  NAND U2179 ( .A(n1311), .B(n1310), .Z(n1442) );
  AND U2180 ( .A(x[139]), .B(y[642]), .Z(n1965) );
  AND U2181 ( .A(y[644]), .B(x[141]), .Z(n1439) );
  NAND U2182 ( .A(n1965), .B(n1439), .Z(n1315) );
  NAND U2183 ( .A(n1313), .B(n1312), .Z(n1314) );
  AND U2184 ( .A(n1315), .B(n1314), .Z(n1425) );
  AND U2185 ( .A(y[647]), .B(x[137]), .Z(n1317) );
  NAND U2186 ( .A(x[130]), .B(y[654]), .Z(n1316) );
  XNOR U2187 ( .A(n1317), .B(n1316), .Z(n1432) );
  NAND U2188 ( .A(y[653]), .B(x[131]), .Z(n1433) );
  XNOR U2189 ( .A(n1432), .B(n1433), .Z(n1423) );
  AND U2190 ( .A(x[140]), .B(y[644]), .Z(n2131) );
  AND U2191 ( .A(y[643]), .B(x[141]), .Z(n1319) );
  NAND U2192 ( .A(x[133]), .B(y[651]), .Z(n1318) );
  XOR U2193 ( .A(n1319), .B(n1318), .Z(n1379) );
  XNOR U2194 ( .A(n2131), .B(n1379), .Z(n1422) );
  XOR U2195 ( .A(n1423), .B(n1422), .Z(n1424) );
  XNOR U2196 ( .A(n1425), .B(n1424), .Z(n1441) );
  NAND U2197 ( .A(n1321), .B(n1320), .Z(n1325) );
  NANDN U2198 ( .A(n1323), .B(n1322), .Z(n1324) );
  AND U2199 ( .A(n1325), .B(n1324), .Z(n1440) );
  XOR U2200 ( .A(n1442), .B(n1443), .Z(n1412) );
  XOR U2201 ( .A(n1413), .B(n1412), .Z(n1447) );
  NAND U2202 ( .A(n1327), .B(n1326), .Z(n1331) );
  NANDN U2203 ( .A(n1329), .B(n1328), .Z(n1330) );
  AND U2204 ( .A(n1331), .B(n1330), .Z(n1446) );
  XNOR U2205 ( .A(n1447), .B(n1446), .Z(n1449) );
  NANDN U2206 ( .A(n1333), .B(n1332), .Z(n1337) );
  NANDN U2207 ( .A(n1335), .B(n1334), .Z(n1336) );
  AND U2208 ( .A(n1337), .B(n1336), .Z(n1363) );
  NANDN U2209 ( .A(n1339), .B(n1338), .Z(n1343) );
  NANDN U2210 ( .A(n1341), .B(n1340), .Z(n1342) );
  AND U2211 ( .A(n1343), .B(n1342), .Z(n1361) );
  NANDN U2212 ( .A(n1345), .B(n1344), .Z(n1349) );
  NANDN U2213 ( .A(n1347), .B(n1346), .Z(n1348) );
  AND U2214 ( .A(n1349), .B(n1348), .Z(n1360) );
  XNOR U2215 ( .A(n1361), .B(n1360), .Z(n1362) );
  XNOR U2216 ( .A(n1363), .B(n1362), .Z(n1448) );
  XOR U2217 ( .A(n1449), .B(n1448), .Z(n1455) );
  NAND U2218 ( .A(n1354), .B(n1353), .Z(n1358) );
  NANDN U2219 ( .A(n1356), .B(n1355), .Z(n1357) );
  AND U2220 ( .A(n1358), .B(n1357), .Z(n1454) );
  IV U2221 ( .A(n1454), .Z(n1452) );
  XOR U2222 ( .A(n1453), .B(n1452), .Z(n1359) );
  XNOR U2223 ( .A(n1455), .B(n1359), .Z(N49) );
  NANDN U2224 ( .A(n1361), .B(n1360), .Z(n1365) );
  NANDN U2225 ( .A(n1363), .B(n1362), .Z(n1364) );
  AND U2226 ( .A(n1365), .B(n1364), .Z(n1562) );
  NANDN U2227 ( .A(n1367), .B(n1366), .Z(n1371) );
  NANDN U2228 ( .A(n1369), .B(n1368), .Z(n1370) );
  NAND U2229 ( .A(n1371), .B(n1370), .Z(n1468) );
  NAND U2230 ( .A(n1373), .B(n1372), .Z(n1377) );
  NAND U2231 ( .A(n1375), .B(n1374), .Z(n1376) );
  AND U2232 ( .A(n1377), .B(n1376), .Z(n1553) );
  AND U2233 ( .A(y[651]), .B(x[141]), .Z(n2400) );
  NAND U2234 ( .A(n2400), .B(n1378), .Z(n1381) );
  NANDN U2235 ( .A(n1379), .B(n2131), .Z(n1380) );
  AND U2236 ( .A(n1381), .B(n1380), .Z(n1501) );
  AND U2237 ( .A(y[648]), .B(x[137]), .Z(n1383) );
  NAND U2238 ( .A(x[129]), .B(y[656]), .Z(n1382) );
  XNOR U2239 ( .A(n1383), .B(n1382), .Z(n1522) );
  ANDN U2240 ( .B(o[16]), .A(n1384), .Z(n1521) );
  XOR U2241 ( .A(n1522), .B(n1521), .Z(n1499) );
  AND U2242 ( .A(x[143]), .B(y[642]), .Z(n1386) );
  NAND U2243 ( .A(y[645]), .B(x[140]), .Z(n1385) );
  XNOR U2244 ( .A(n1386), .B(n1385), .Z(n1473) );
  AND U2245 ( .A(x[142]), .B(y[643]), .Z(n1472) );
  XOR U2246 ( .A(n1473), .B(n1472), .Z(n1498) );
  XOR U2247 ( .A(n1499), .B(n1498), .Z(n1500) );
  XNOR U2248 ( .A(n1501), .B(n1500), .Z(n1551) );
  NAND U2249 ( .A(x[135]), .B(y[650]), .Z(n1533) );
  NANDN U2250 ( .A(n1533), .B(n1387), .Z(n1391) );
  NAND U2251 ( .A(n1389), .B(n1388), .Z(n1390) );
  AND U2252 ( .A(n1391), .B(n1390), .Z(n1511) );
  NAND U2253 ( .A(x[136]), .B(y[655]), .Z(n2218) );
  NANDN U2254 ( .A(n2218), .B(n1616), .Z(n1395) );
  NAND U2255 ( .A(n1393), .B(n1392), .Z(n1394) );
  NAND U2256 ( .A(n1395), .B(n1394), .Z(n1510) );
  XNOR U2257 ( .A(n1511), .B(n1510), .Z(n1513) );
  NANDN U2258 ( .A(n1397), .B(n1396), .Z(n1401) );
  NAND U2259 ( .A(n1399), .B(n1398), .Z(n1400) );
  AND U2260 ( .A(n1401), .B(n1400), .Z(n1507) );
  AND U2261 ( .A(y[657]), .B(x[128]), .Z(n1487) );
  AND U2262 ( .A(x[145]), .B(y[640]), .Z(n1486) );
  XOR U2263 ( .A(n1487), .B(n1486), .Z(n1489) );
  AND U2264 ( .A(x[144]), .B(y[641]), .Z(n1483) );
  XOR U2265 ( .A(n1483), .B(o[17]), .Z(n1488) );
  XOR U2266 ( .A(n1489), .B(n1488), .Z(n1505) );
  AND U2267 ( .A(x[130]), .B(y[655]), .Z(n1403) );
  NAND U2268 ( .A(y[647]), .B(x[138]), .Z(n1402) );
  XNOR U2269 ( .A(n1403), .B(n1402), .Z(n1526) );
  NAND U2270 ( .A(y[654]), .B(x[131]), .Z(n1527) );
  XOR U2271 ( .A(n1505), .B(n1504), .Z(n1506) );
  XNOR U2272 ( .A(n1507), .B(n1506), .Z(n1512) );
  XOR U2273 ( .A(n1513), .B(n1512), .Z(n1550) );
  XOR U2274 ( .A(n1551), .B(n1550), .Z(n1552) );
  XNOR U2275 ( .A(n1553), .B(n1552), .Z(n1467) );
  NAND U2276 ( .A(n1405), .B(n1404), .Z(n1409) );
  NAND U2277 ( .A(n1407), .B(n1406), .Z(n1408) );
  AND U2278 ( .A(n1409), .B(n1408), .Z(n1466) );
  XOR U2279 ( .A(n1468), .B(n1469), .Z(n1560) );
  NANDN U2280 ( .A(n1411), .B(n1410), .Z(n1415) );
  NAND U2281 ( .A(n1413), .B(n1412), .Z(n1414) );
  NAND U2282 ( .A(n1415), .B(n1414), .Z(n1462) );
  NANDN U2283 ( .A(n1417), .B(n1416), .Z(n1421) );
  NAND U2284 ( .A(n1419), .B(n1418), .Z(n1420) );
  AND U2285 ( .A(n1421), .B(n1420), .Z(n1547) );
  NAND U2286 ( .A(n1423), .B(n1422), .Z(n1427) );
  NANDN U2287 ( .A(n1425), .B(n1424), .Z(n1426) );
  AND U2288 ( .A(n1427), .B(n1426), .Z(n1545) );
  NAND U2289 ( .A(y[645]), .B(x[142]), .Z(n1734) );
  NANDN U2290 ( .A(n1734), .B(n1965), .Z(n1431) );
  NANDN U2291 ( .A(n1429), .B(n1428), .Z(n1430) );
  AND U2292 ( .A(n1431), .B(n1430), .Z(n1539) );
  AND U2293 ( .A(x[137]), .B(y[654]), .Z(n2381) );
  NANDN U2294 ( .A(n1525), .B(n2381), .Z(n1435) );
  NANDN U2295 ( .A(n1433), .B(n1432), .Z(n1434) );
  NAND U2296 ( .A(n1435), .B(n1434), .Z(n1538) );
  XNOR U2297 ( .A(n1539), .B(n1538), .Z(n1541) );
  AND U2298 ( .A(y[652]), .B(x[133]), .Z(n1597) );
  NAND U2299 ( .A(y[649]), .B(x[136]), .Z(n1436) );
  XNOR U2300 ( .A(n1597), .B(n1436), .Z(n1517) );
  XOR U2301 ( .A(n1517), .B(n1437), .Z(n1532) );
  XNOR U2302 ( .A(n1532), .B(n1533), .Z(n1535) );
  NAND U2303 ( .A(x[132]), .B(y[653]), .Z(n1438) );
  XNOR U2304 ( .A(n1439), .B(n1438), .Z(n1477) );
  NAND U2305 ( .A(x[139]), .B(y[646]), .Z(n1478) );
  XNOR U2306 ( .A(n1477), .B(n1478), .Z(n1534) );
  XOR U2307 ( .A(n1535), .B(n1534), .Z(n1540) );
  XOR U2308 ( .A(n1541), .B(n1540), .Z(n1544) );
  XNOR U2309 ( .A(n1545), .B(n1544), .Z(n1546) );
  XNOR U2310 ( .A(n1547), .B(n1546), .Z(n1461) );
  NANDN U2311 ( .A(n1441), .B(n1440), .Z(n1445) );
  NAND U2312 ( .A(n1443), .B(n1442), .Z(n1444) );
  NAND U2313 ( .A(n1445), .B(n1444), .Z(n1460) );
  XOR U2314 ( .A(n1462), .B(n1463), .Z(n1559) );
  XOR U2315 ( .A(n1560), .B(n1559), .Z(n1561) );
  XOR U2316 ( .A(n1562), .B(n1561), .Z(n1558) );
  NANDN U2317 ( .A(n1447), .B(n1446), .Z(n1451) );
  NAND U2318 ( .A(n1449), .B(n1448), .Z(n1450) );
  NAND U2319 ( .A(n1451), .B(n1450), .Z(n1557) );
  NANDN U2320 ( .A(n1452), .B(n1453), .Z(n1458) );
  NOR U2321 ( .A(n1454), .B(n1453), .Z(n1456) );
  OR U2322 ( .A(n1456), .B(n1455), .Z(n1457) );
  AND U2323 ( .A(n1458), .B(n1457), .Z(n1556) );
  XOR U2324 ( .A(n1557), .B(n1556), .Z(n1459) );
  XNOR U2325 ( .A(n1558), .B(n1459), .Z(N50) );
  NANDN U2326 ( .A(n1461), .B(n1460), .Z(n1465) );
  NANDN U2327 ( .A(n1463), .B(n1462), .Z(n1464) );
  AND U2328 ( .A(n1465), .B(n1464), .Z(n1569) );
  NANDN U2329 ( .A(n1467), .B(n1466), .Z(n1471) );
  NANDN U2330 ( .A(n1469), .B(n1468), .Z(n1470) );
  AND U2331 ( .A(n1471), .B(n1470), .Z(n1567) );
  AND U2332 ( .A(x[143]), .B(y[645]), .Z(n1708) );
  NAND U2333 ( .A(n1708), .B(n1812), .Z(n1475) );
  NAND U2334 ( .A(n1473), .B(n1472), .Z(n1474) );
  NAND U2335 ( .A(n1475), .B(n1474), .Z(n1664) );
  NAND U2336 ( .A(n2739), .B(n1476), .Z(n1480) );
  NANDN U2337 ( .A(n1478), .B(n1477), .Z(n1479) );
  AND U2338 ( .A(n1480), .B(n1479), .Z(n1655) );
  AND U2339 ( .A(x[129]), .B(y[657]), .Z(n1482) );
  NAND U2340 ( .A(y[648]), .B(x[138]), .Z(n1481) );
  XNOR U2341 ( .A(n1482), .B(n1481), .Z(n1617) );
  NAND U2342 ( .A(n1483), .B(o[17]), .Z(n1618) );
  NAND U2343 ( .A(y[643]), .B(x[143]), .Z(n1484) );
  XNOR U2344 ( .A(n1485), .B(n1484), .Z(n1608) );
  NAND U2345 ( .A(y[644]), .B(x[142]), .Z(n1609) );
  XOR U2346 ( .A(n1653), .B(n1652), .Z(n1654) );
  XOR U2347 ( .A(n1664), .B(n1665), .Z(n1667) );
  NAND U2348 ( .A(n1487), .B(n1486), .Z(n1491) );
  NAND U2349 ( .A(n1489), .B(n1488), .Z(n1490) );
  NAND U2350 ( .A(n1491), .B(n1490), .Z(n1676) );
  AND U2351 ( .A(y[647]), .B(x[139]), .Z(n1493) );
  NAND U2352 ( .A(y[642]), .B(x[144]), .Z(n1492) );
  XNOR U2353 ( .A(n1493), .B(n1492), .Z(n1604) );
  NAND U2354 ( .A(y[656]), .B(x[130]), .Z(n1605) );
  XOR U2355 ( .A(n1676), .B(n1677), .Z(n1679) );
  AND U2356 ( .A(y[652]), .B(x[134]), .Z(n1495) );
  NAND U2357 ( .A(x[133]), .B(y[653]), .Z(n1494) );
  XNOR U2358 ( .A(n1495), .B(n1494), .Z(n1600) );
  AND U2359 ( .A(y[654]), .B(x[132]), .Z(n1497) );
  NAND U2360 ( .A(y[650]), .B(x[136]), .Z(n1496) );
  XNOR U2361 ( .A(n1497), .B(n1496), .Z(n1639) );
  NAND U2362 ( .A(y[651]), .B(x[135]), .Z(n1640) );
  XOR U2363 ( .A(n1600), .B(n1599), .Z(n1678) );
  XOR U2364 ( .A(n1679), .B(n1678), .Z(n1666) );
  XOR U2365 ( .A(n1667), .B(n1666), .Z(n1586) );
  NAND U2366 ( .A(n1499), .B(n1498), .Z(n1503) );
  NANDN U2367 ( .A(n1501), .B(n1500), .Z(n1502) );
  AND U2368 ( .A(n1503), .B(n1502), .Z(n1659) );
  NAND U2369 ( .A(n1505), .B(n1504), .Z(n1509) );
  NANDN U2370 ( .A(n1507), .B(n1506), .Z(n1508) );
  AND U2371 ( .A(n1509), .B(n1508), .Z(n1658) );
  XOR U2372 ( .A(n1659), .B(n1658), .Z(n1661) );
  NANDN U2373 ( .A(n1511), .B(n1510), .Z(n1515) );
  NAND U2374 ( .A(n1513), .B(n1512), .Z(n1514) );
  AND U2375 ( .A(n1515), .B(n1514), .Z(n1660) );
  XOR U2376 ( .A(n1661), .B(n1660), .Z(n1585) );
  XNOR U2377 ( .A(n1586), .B(n1585), .Z(n1588) );
  AND U2378 ( .A(x[136]), .B(y[652]), .Z(n1852) );
  NAND U2379 ( .A(n1852), .B(n1516), .Z(n1520) );
  NANDN U2380 ( .A(n1518), .B(n1517), .Z(n1519) );
  NAND U2381 ( .A(n1520), .B(n1519), .Z(n1671) );
  NAND U2382 ( .A(y[656]), .B(x[137]), .Z(n2509) );
  NANDN U2383 ( .A(n2509), .B(n1616), .Z(n1524) );
  NAND U2384 ( .A(n1522), .B(n1521), .Z(n1523) );
  NAND U2385 ( .A(n1524), .B(n1523), .Z(n1670) );
  XOR U2386 ( .A(n1671), .B(n1670), .Z(n1673) );
  NAND U2387 ( .A(x[138]), .B(y[655]), .Z(n2409) );
  IV U2388 ( .A(n2409), .Z(n2510) );
  NANDN U2389 ( .A(n1525), .B(n2510), .Z(n1529) );
  NANDN U2390 ( .A(n1527), .B(n1526), .Z(n1528) );
  AND U2391 ( .A(n1529), .B(n1528), .Z(n1649) );
  AND U2392 ( .A(x[128]), .B(y[658]), .Z(n1621) );
  NAND U2393 ( .A(x[146]), .B(y[640]), .Z(n1622) );
  NAND U2394 ( .A(y[641]), .B(x[145]), .Z(n1643) );
  XNOR U2395 ( .A(o[18]), .B(n1643), .Z(n1623) );
  XOR U2396 ( .A(n1624), .B(n1623), .Z(n1647) );
  AND U2397 ( .A(x[131]), .B(y[655]), .Z(n1531) );
  NAND U2398 ( .A(x[141]), .B(y[645]), .Z(n1530) );
  XNOR U2399 ( .A(n1531), .B(n1530), .Z(n1630) );
  NAND U2400 ( .A(x[140]), .B(y[646]), .Z(n1631) );
  XOR U2401 ( .A(n1647), .B(n1646), .Z(n1648) );
  XOR U2402 ( .A(n1673), .B(n1672), .Z(n1592) );
  NANDN U2403 ( .A(n1533), .B(n1532), .Z(n1537) );
  NAND U2404 ( .A(n1535), .B(n1534), .Z(n1536) );
  AND U2405 ( .A(n1537), .B(n1536), .Z(n1591) );
  NANDN U2406 ( .A(n1539), .B(n1538), .Z(n1543) );
  NAND U2407 ( .A(n1541), .B(n1540), .Z(n1542) );
  NAND U2408 ( .A(n1543), .B(n1542), .Z(n1594) );
  XOR U2409 ( .A(n1588), .B(n1587), .Z(n1582) );
  NANDN U2410 ( .A(n1545), .B(n1544), .Z(n1549) );
  NANDN U2411 ( .A(n1547), .B(n1546), .Z(n1548) );
  AND U2412 ( .A(n1549), .B(n1548), .Z(n1580) );
  NAND U2413 ( .A(n1551), .B(n1550), .Z(n1555) );
  NANDN U2414 ( .A(n1553), .B(n1552), .Z(n1554) );
  NAND U2415 ( .A(n1555), .B(n1554), .Z(n1579) );
  XNOR U2416 ( .A(n1580), .B(n1579), .Z(n1581) );
  XNOR U2417 ( .A(n1582), .B(n1581), .Z(n1566) );
  XOR U2418 ( .A(n1567), .B(n1566), .Z(n1568) );
  XOR U2419 ( .A(n1569), .B(n1568), .Z(n1575) );
  NAND U2420 ( .A(n1560), .B(n1559), .Z(n1564) );
  NANDN U2421 ( .A(n1562), .B(n1561), .Z(n1563) );
  AND U2422 ( .A(n1564), .B(n1563), .Z(n1574) );
  IV U2423 ( .A(n1574), .Z(n1572) );
  XOR U2424 ( .A(n1573), .B(n1572), .Z(n1565) );
  XNOR U2425 ( .A(n1575), .B(n1565), .Z(N51) );
  NAND U2426 ( .A(n1567), .B(n1566), .Z(n1571) );
  NAND U2427 ( .A(n1569), .B(n1568), .Z(n1570) );
  AND U2428 ( .A(n1571), .B(n1570), .Z(n1796) );
  NANDN U2429 ( .A(n1572), .B(n1573), .Z(n1578) );
  NOR U2430 ( .A(n1574), .B(n1573), .Z(n1576) );
  OR U2431 ( .A(n1576), .B(n1575), .Z(n1577) );
  AND U2432 ( .A(n1578), .B(n1577), .Z(n1797) );
  NANDN U2433 ( .A(n1580), .B(n1579), .Z(n1584) );
  NANDN U2434 ( .A(n1582), .B(n1581), .Z(n1583) );
  AND U2435 ( .A(n1584), .B(n1583), .Z(n1793) );
  NANDN U2436 ( .A(n1586), .B(n1585), .Z(n1590) );
  NAND U2437 ( .A(n1588), .B(n1587), .Z(n1589) );
  AND U2438 ( .A(n1590), .B(n1589), .Z(n1791) );
  NANDN U2439 ( .A(n1592), .B(n1591), .Z(n1596) );
  NANDN U2440 ( .A(n1594), .B(n1593), .Z(n1595) );
  AND U2441 ( .A(n1596), .B(n1595), .Z(n1775) );
  AND U2442 ( .A(y[653]), .B(x[134]), .Z(n1598) );
  NAND U2443 ( .A(n1598), .B(n1597), .Z(n1602) );
  NAND U2444 ( .A(n1600), .B(n1599), .Z(n1601) );
  AND U2445 ( .A(n1602), .B(n1601), .Z(n1769) );
  AND U2446 ( .A(x[144]), .B(y[647]), .Z(n1603) );
  NAND U2447 ( .A(n1603), .B(n1965), .Z(n1607) );
  NANDN U2448 ( .A(n1605), .B(n1604), .Z(n1606) );
  AND U2449 ( .A(n1607), .B(n1606), .Z(n1767) );
  AND U2450 ( .A(x[143]), .B(y[649]), .Z(n2412) );
  NAND U2451 ( .A(n2412), .B(n1695), .Z(n1611) );
  NANDN U2452 ( .A(n1609), .B(n1608), .Z(n1610) );
  AND U2453 ( .A(n1611), .B(n1610), .Z(n1686) );
  AND U2454 ( .A(y[658]), .B(x[129]), .Z(n1613) );
  NAND U2455 ( .A(x[136]), .B(y[651]), .Z(n1612) );
  XNOR U2456 ( .A(n1613), .B(n1612), .Z(n1733) );
  XNOR U2457 ( .A(n1733), .B(n1734), .Z(n1684) );
  AND U2458 ( .A(x[141]), .B(y[646]), .Z(n1615) );
  NAND U2459 ( .A(x[130]), .B(y[657]), .Z(n1614) );
  XNOR U2460 ( .A(n1615), .B(n1614), .Z(n1701) );
  XOR U2461 ( .A(n1684), .B(n1683), .Z(n1685) );
  NAND U2462 ( .A(x[138]), .B(y[657]), .Z(n2831) );
  NANDN U2463 ( .A(n2831), .B(n1616), .Z(n1620) );
  NANDN U2464 ( .A(n1618), .B(n1617), .Z(n1619) );
  AND U2465 ( .A(n1620), .B(n1619), .Z(n1745) );
  NANDN U2466 ( .A(n1622), .B(n1621), .Z(n1626) );
  NAND U2467 ( .A(n1624), .B(n1623), .Z(n1625) );
  AND U2468 ( .A(n1626), .B(n1625), .Z(n1743) );
  AND U2469 ( .A(x[137]), .B(y[650]), .Z(n1628) );
  NAND U2470 ( .A(y[643]), .B(x[144]), .Z(n1627) );
  XNOR U2471 ( .A(n1628), .B(n1627), .Z(n1696) );
  NAND U2472 ( .A(x[143]), .B(y[644]), .Z(n1697) );
  XNOR U2473 ( .A(n1696), .B(n1697), .Z(n1742) );
  AND U2474 ( .A(x[141]), .B(y[655]), .Z(n3031) );
  NANDN U2475 ( .A(n1629), .B(n3031), .Z(n1633) );
  NANDN U2476 ( .A(n1631), .B(n1630), .Z(n1632) );
  AND U2477 ( .A(n1633), .B(n1632), .Z(n1751) );
  AND U2478 ( .A(x[145]), .B(y[642]), .Z(n1635) );
  NAND U2479 ( .A(y[649]), .B(x[138]), .Z(n1634) );
  XNOR U2480 ( .A(n1635), .B(n1634), .Z(n1739) );
  NAND U2481 ( .A(y[641]), .B(x[146]), .Z(n1715) );
  XNOR U2482 ( .A(o[19]), .B(n1715), .Z(n1738) );
  XOR U2483 ( .A(n1739), .B(n1738), .Z(n1749) );
  AND U2484 ( .A(x[131]), .B(y[656]), .Z(n1637) );
  NAND U2485 ( .A(y[648]), .B(x[139]), .Z(n1636) );
  XNOR U2486 ( .A(n1637), .B(n1636), .Z(n1709) );
  XOR U2487 ( .A(n1749), .B(n1748), .Z(n1750) );
  NAND U2488 ( .A(n2013), .B(n1638), .Z(n1642) );
  NANDN U2489 ( .A(n1640), .B(n1639), .Z(n1641) );
  AND U2490 ( .A(n1642), .B(n1641), .Z(n1692) );
  AND U2491 ( .A(y[659]), .B(x[128]), .Z(n1720) );
  NAND U2492 ( .A(x[147]), .B(y[640]), .Z(n1721) );
  XNOR U2493 ( .A(n1720), .B(n1721), .Z(n1723) );
  ANDN U2494 ( .B(o[18]), .A(n1643), .Z(n1722) );
  XOR U2495 ( .A(n1723), .B(n1722), .Z(n1690) );
  AND U2496 ( .A(x[132]), .B(y[655]), .Z(n1866) );
  AND U2497 ( .A(x[133]), .B(y[654]), .Z(n1645) );
  NAND U2498 ( .A(x[134]), .B(y[653]), .Z(n1644) );
  XOR U2499 ( .A(n1645), .B(n1644), .Z(n1717) );
  XNOR U2500 ( .A(n1866), .B(n1717), .Z(n1689) );
  XOR U2501 ( .A(n1690), .B(n1689), .Z(n1691) );
  XOR U2502 ( .A(n1692), .B(n1691), .Z(n1760) );
  XOR U2503 ( .A(n1761), .B(n1760), .Z(n1763) );
  XNOR U2504 ( .A(n1762), .B(n1763), .Z(n1756) );
  NAND U2505 ( .A(n1647), .B(n1646), .Z(n1651) );
  NANDN U2506 ( .A(n1649), .B(n1648), .Z(n1650) );
  AND U2507 ( .A(n1651), .B(n1650), .Z(n1755) );
  NAND U2508 ( .A(n1653), .B(n1652), .Z(n1657) );
  NANDN U2509 ( .A(n1655), .B(n1654), .Z(n1656) );
  NAND U2510 ( .A(n1657), .B(n1656), .Z(n1754) );
  XNOR U2511 ( .A(n1756), .B(n1757), .Z(n1772) );
  XOR U2512 ( .A(n1773), .B(n1772), .Z(n1774) );
  NAND U2513 ( .A(n1659), .B(n1658), .Z(n1663) );
  NAND U2514 ( .A(n1661), .B(n1660), .Z(n1662) );
  AND U2515 ( .A(n1663), .B(n1662), .Z(n1784) );
  NAND U2516 ( .A(n1665), .B(n1664), .Z(n1669) );
  NAND U2517 ( .A(n1667), .B(n1666), .Z(n1668) );
  NAND U2518 ( .A(n1669), .B(n1668), .Z(n1780) );
  NAND U2519 ( .A(n1671), .B(n1670), .Z(n1675) );
  NAND U2520 ( .A(n1673), .B(n1672), .Z(n1674) );
  NAND U2521 ( .A(n1675), .B(n1674), .Z(n1779) );
  NAND U2522 ( .A(n1677), .B(n1676), .Z(n1681) );
  NAND U2523 ( .A(n1679), .B(n1678), .Z(n1680) );
  NAND U2524 ( .A(n1681), .B(n1680), .Z(n1778) );
  XNOR U2525 ( .A(n1779), .B(n1778), .Z(n1781) );
  XNOR U2526 ( .A(n1784), .B(n1785), .Z(n1786) );
  XOR U2527 ( .A(n1791), .B(n1790), .Z(n1792) );
  XNOR U2528 ( .A(n1793), .B(n1792), .Z(n1798) );
  XNOR U2529 ( .A(n1797), .B(n1798), .Z(n1682) );
  XOR U2530 ( .A(n1796), .B(n1682), .Z(N52) );
  NAND U2531 ( .A(n1684), .B(n1683), .Z(n1688) );
  NANDN U2532 ( .A(n1686), .B(n1685), .Z(n1687) );
  AND U2533 ( .A(n1688), .B(n1687), .Z(n1801) );
  NAND U2534 ( .A(n1690), .B(n1689), .Z(n1694) );
  NANDN U2535 ( .A(n1692), .B(n1691), .Z(n1693) );
  NAND U2536 ( .A(n1694), .B(n1693), .Z(n1800) );
  AND U2537 ( .A(x[144]), .B(y[650]), .Z(n2659) );
  NAND U2538 ( .A(n2659), .B(n1695), .Z(n1699) );
  NANDN U2539 ( .A(n1697), .B(n1696), .Z(n1698) );
  AND U2540 ( .A(n1699), .B(n1698), .Z(n1841) );
  AND U2541 ( .A(y[657]), .B(x[141]), .Z(n3171) );
  NAND U2542 ( .A(n3171), .B(n1700), .Z(n1704) );
  NANDN U2543 ( .A(n1702), .B(n1701), .Z(n1703) );
  AND U2544 ( .A(n1704), .B(n1703), .Z(n1886) );
  NAND U2545 ( .A(y[644]), .B(x[144]), .Z(n1705) );
  XNOR U2546 ( .A(n1706), .B(n1705), .Z(n1847) );
  NAND U2547 ( .A(x[130]), .B(y[658]), .Z(n1848) );
  XNOR U2548 ( .A(n1847), .B(n1848), .Z(n1884) );
  NAND U2549 ( .A(x[137]), .B(y[651]), .Z(n1707) );
  XNOR U2550 ( .A(n1708), .B(n1707), .Z(n1823) );
  NAND U2551 ( .A(y[646]), .B(x[142]), .Z(n1824) );
  XNOR U2552 ( .A(n1823), .B(n1824), .Z(n1883) );
  XOR U2553 ( .A(n1884), .B(n1883), .Z(n1885) );
  XNOR U2554 ( .A(n1886), .B(n1885), .Z(n1840) );
  XNOR U2555 ( .A(n1841), .B(n1840), .Z(n1843) );
  NAND U2556 ( .A(x[139]), .B(y[656]), .Z(n2833) );
  NANDN U2557 ( .A(n2833), .B(n1992), .Z(n1712) );
  NANDN U2558 ( .A(n1710), .B(n1709), .Z(n1711) );
  AND U2559 ( .A(n1712), .B(n1711), .Z(n1892) );
  AND U2560 ( .A(x[129]), .B(y[659]), .Z(n1714) );
  NAND U2561 ( .A(y[649]), .B(x[139]), .Z(n1713) );
  XNOR U2562 ( .A(n1714), .B(n1713), .Z(n1819) );
  NAND U2563 ( .A(y[641]), .B(x[147]), .Z(n1827) );
  XOR U2564 ( .A(n1819), .B(n1818), .Z(n1890) );
  AND U2565 ( .A(x[128]), .B(y[660]), .Z(n1871) );
  NAND U2566 ( .A(y[640]), .B(x[148]), .Z(n1872) );
  XNOR U2567 ( .A(n1871), .B(n1872), .Z(n1874) );
  ANDN U2568 ( .B(o[19]), .A(n1715), .Z(n1873) );
  XOR U2569 ( .A(n1874), .B(n1873), .Z(n1889) );
  XOR U2570 ( .A(n1890), .B(n1889), .Z(n1891) );
  XNOR U2571 ( .A(n1892), .B(n1891), .Z(n1842) );
  XOR U2572 ( .A(n1843), .B(n1842), .Z(n1802) );
  XOR U2573 ( .A(n1803), .B(n1802), .Z(n1898) );
  AND U2574 ( .A(x[134]), .B(y[654]), .Z(n1807) );
  AND U2575 ( .A(y[653]), .B(x[133]), .Z(n1716) );
  NAND U2576 ( .A(n1807), .B(n1716), .Z(n1719) );
  NANDN U2577 ( .A(n1717), .B(n1866), .Z(n1718) );
  AND U2578 ( .A(n1719), .B(n1718), .Z(n1831) );
  NANDN U2579 ( .A(n1721), .B(n1720), .Z(n1725) );
  NAND U2580 ( .A(n1723), .B(n1722), .Z(n1724) );
  AND U2581 ( .A(n1725), .B(n1724), .Z(n1829) );
  AND U2582 ( .A(x[146]), .B(y[642]), .Z(n1727) );
  NAND U2583 ( .A(y[648]), .B(x[140]), .Z(n1726) );
  XNOR U2584 ( .A(n1727), .B(n1726), .Z(n1813) );
  NAND U2585 ( .A(x[145]), .B(y[643]), .Z(n1814) );
  XNOR U2586 ( .A(n1813), .B(n1814), .Z(n1828) );
  XNOR U2587 ( .A(n1829), .B(n1828), .Z(n1830) );
  XOR U2588 ( .A(n1831), .B(n1830), .Z(n1835) );
  AND U2589 ( .A(y[647]), .B(x[141]), .Z(n1729) );
  NAND U2590 ( .A(x[131]), .B(y[657]), .Z(n1728) );
  XNOR U2591 ( .A(n1729), .B(n1728), .Z(n1853) );
  XOR U2592 ( .A(n1853), .B(n1852), .Z(n1809) );
  AND U2593 ( .A(x[133]), .B(y[655]), .Z(n1731) );
  NAND U2594 ( .A(x[132]), .B(y[656]), .Z(n1730) );
  XNOR U2595 ( .A(n1731), .B(n1730), .Z(n1868) );
  AND U2596 ( .A(x[135]), .B(y[653]), .Z(n1867) );
  XNOR U2597 ( .A(n1868), .B(n1867), .Z(n1806) );
  XNOR U2598 ( .A(n1807), .B(n1806), .Z(n1808) );
  XOR U2599 ( .A(n1809), .B(n1808), .Z(n1879) );
  AND U2600 ( .A(x[136]), .B(y[658]), .Z(n2977) );
  AND U2601 ( .A(y[651]), .B(x[129]), .Z(n1732) );
  NAND U2602 ( .A(n2977), .B(n1732), .Z(n1736) );
  NANDN U2603 ( .A(n1734), .B(n1733), .Z(n1735) );
  AND U2604 ( .A(n1736), .B(n1735), .Z(n1878) );
  AND U2605 ( .A(x[145]), .B(y[649]), .Z(n2665) );
  AND U2606 ( .A(x[138]), .B(y[642]), .Z(n1737) );
  NAND U2607 ( .A(n2665), .B(n1737), .Z(n1741) );
  NAND U2608 ( .A(n1739), .B(n1738), .Z(n1740) );
  NAND U2609 ( .A(n1741), .B(n1740), .Z(n1877) );
  XNOR U2610 ( .A(n1878), .B(n1877), .Z(n1880) );
  XNOR U2611 ( .A(n1879), .B(n1880), .Z(n1834) );
  XOR U2612 ( .A(n1835), .B(n1834), .Z(n1836) );
  NANDN U2613 ( .A(n1743), .B(n1742), .Z(n1747) );
  NANDN U2614 ( .A(n1745), .B(n1744), .Z(n1746) );
  NAND U2615 ( .A(n1747), .B(n1746), .Z(n1837) );
  NAND U2616 ( .A(n1749), .B(n1748), .Z(n1753) );
  NANDN U2617 ( .A(n1751), .B(n1750), .Z(n1752) );
  NAND U2618 ( .A(n1753), .B(n1752), .Z(n1896) );
  NANDN U2619 ( .A(n1755), .B(n1754), .Z(n1759) );
  NAND U2620 ( .A(n1757), .B(n1756), .Z(n1758) );
  AND U2621 ( .A(n1759), .B(n1758), .Z(n1910) );
  NAND U2622 ( .A(n1761), .B(n1760), .Z(n1765) );
  NAND U2623 ( .A(n1763), .B(n1762), .Z(n1764) );
  AND U2624 ( .A(n1765), .B(n1764), .Z(n1908) );
  NANDN U2625 ( .A(n1767), .B(n1766), .Z(n1771) );
  NANDN U2626 ( .A(n1769), .B(n1768), .Z(n1770) );
  AND U2627 ( .A(n1771), .B(n1770), .Z(n1907) );
  XNOR U2628 ( .A(n1910), .B(n1909), .Z(n1901) );
  XOR U2629 ( .A(n1902), .B(n1901), .Z(n1903) );
  NAND U2630 ( .A(n1773), .B(n1772), .Z(n1777) );
  NANDN U2631 ( .A(n1775), .B(n1774), .Z(n1776) );
  NAND U2632 ( .A(n1777), .B(n1776), .Z(n1904) );
  NAND U2633 ( .A(n1779), .B(n1778), .Z(n1783) );
  NANDN U2634 ( .A(n1781), .B(n1780), .Z(n1782) );
  AND U2635 ( .A(n1783), .B(n1782), .Z(n1917) );
  NANDN U2636 ( .A(n1785), .B(n1784), .Z(n1789) );
  NANDN U2637 ( .A(n1787), .B(n1786), .Z(n1788) );
  AND U2638 ( .A(n1789), .B(n1788), .Z(n1916) );
  XOR U2639 ( .A(n1917), .B(n1916), .Z(n1918) );
  NAND U2640 ( .A(n1791), .B(n1790), .Z(n1795) );
  NANDN U2641 ( .A(n1793), .B(n1792), .Z(n1794) );
  NAND U2642 ( .A(n1795), .B(n1794), .Z(n1914) );
  XOR U2643 ( .A(n1914), .B(n1913), .Z(n1799) );
  XNOR U2644 ( .A(n1915), .B(n1799), .Z(N53) );
  NANDN U2645 ( .A(n1801), .B(n1800), .Z(n1805) );
  NAND U2646 ( .A(n1803), .B(n1802), .Z(n1804) );
  AND U2647 ( .A(n1805), .B(n1804), .Z(n1932) );
  NANDN U2648 ( .A(n1807), .B(n1806), .Z(n1811) );
  NANDN U2649 ( .A(n1809), .B(n1808), .Z(n1810) );
  AND U2650 ( .A(n1811), .B(n1810), .Z(n2033) );
  AND U2651 ( .A(x[146]), .B(y[648]), .Z(n2667) );
  NAND U2652 ( .A(n2667), .B(n1812), .Z(n1816) );
  NANDN U2653 ( .A(n1814), .B(n1813), .Z(n1815) );
  AND U2654 ( .A(n1816), .B(n1815), .Z(n2015) );
  AND U2655 ( .A(x[139]), .B(y[659]), .Z(n3459) );
  AND U2656 ( .A(y[649]), .B(x[129]), .Z(n1817) );
  NAND U2657 ( .A(n3459), .B(n1817), .Z(n1821) );
  NAND U2658 ( .A(n1819), .B(n1818), .Z(n1820) );
  NAND U2659 ( .A(n1821), .B(n1820), .Z(n2014) );
  AND U2660 ( .A(y[651]), .B(x[143]), .Z(n2654) );
  NAND U2661 ( .A(n2654), .B(n1822), .Z(n1826) );
  NANDN U2662 ( .A(n1824), .B(n1823), .Z(n1825) );
  AND U2663 ( .A(n1826), .B(n1825), .Z(n1979) );
  AND U2664 ( .A(y[661]), .B(x[128]), .Z(n1998) );
  NAND U2665 ( .A(y[640]), .B(x[149]), .Z(n1999) );
  ANDN U2666 ( .B(o[20]), .A(n1827), .Z(n2000) );
  XOR U2667 ( .A(n2001), .B(n2000), .Z(n1977) );
  AND U2668 ( .A(y[656]), .B(x[133]), .Z(n1983) );
  AND U2669 ( .A(x[144]), .B(y[645]), .Z(n1982) );
  XOR U2670 ( .A(n1983), .B(n1982), .Z(n1985) );
  NAND U2671 ( .A(x[143]), .B(y[646]), .Z(n1984) );
  XNOR U2672 ( .A(n1985), .B(n1984), .Z(n1976) );
  XOR U2673 ( .A(n1977), .B(n1976), .Z(n1978) );
  XNOR U2674 ( .A(n2017), .B(n2016), .Z(n2032) );
  XNOR U2675 ( .A(n2033), .B(n2032), .Z(n2035) );
  NANDN U2676 ( .A(n1829), .B(n1828), .Z(n1833) );
  NANDN U2677 ( .A(n1831), .B(n1830), .Z(n1832) );
  AND U2678 ( .A(n1833), .B(n1832), .Z(n2034) );
  XOR U2679 ( .A(n2035), .B(n2034), .Z(n1930) );
  NAND U2680 ( .A(n1835), .B(n1834), .Z(n1839) );
  NANDN U2681 ( .A(n1837), .B(n1836), .Z(n1838) );
  AND U2682 ( .A(n1839), .B(n1838), .Z(n1929) );
  NANDN U2683 ( .A(n1841), .B(n1840), .Z(n1845) );
  NAND U2684 ( .A(n1843), .B(n1842), .Z(n1844) );
  AND U2685 ( .A(n1845), .B(n1844), .Z(n1938) );
  NAND U2686 ( .A(n2659), .B(n1846), .Z(n1850) );
  NANDN U2687 ( .A(n1848), .B(n1847), .Z(n1849) );
  AND U2688 ( .A(n1850), .B(n1849), .Z(n1948) );
  NAND U2689 ( .A(n3171), .B(n1851), .Z(n1855) );
  NAND U2690 ( .A(n1853), .B(n1852), .Z(n1854) );
  AND U2691 ( .A(n1855), .B(n1854), .Z(n2029) );
  AND U2692 ( .A(x[147]), .B(y[642]), .Z(n1857) );
  NAND U2693 ( .A(y[650]), .B(x[139]), .Z(n1856) );
  XNOR U2694 ( .A(n1857), .B(n1856), .Z(n1967) );
  NAND U2695 ( .A(y[641]), .B(x[148]), .Z(n1997) );
  XNOR U2696 ( .A(o[21]), .B(n1997), .Z(n1966) );
  XOR U2697 ( .A(n1967), .B(n1966), .Z(n2027) );
  AND U2698 ( .A(y[643]), .B(x[146]), .Z(n1859) );
  NAND U2699 ( .A(x[138]), .B(y[651]), .Z(n1858) );
  XNOR U2700 ( .A(n1859), .B(n1858), .Z(n2005) );
  NAND U2701 ( .A(x[129]), .B(y[660]), .Z(n2006) );
  XOR U2702 ( .A(n2027), .B(n2026), .Z(n2028) );
  XNOR U2703 ( .A(n2029), .B(n2028), .Z(n1947) );
  XNOR U2704 ( .A(n1948), .B(n1947), .Z(n1950) );
  AND U2705 ( .A(x[135]), .B(y[654]), .Z(n2216) );
  AND U2706 ( .A(y[647]), .B(x[142]), .Z(n1861) );
  NAND U2707 ( .A(y[655]), .B(x[134]), .Z(n1860) );
  XNOR U2708 ( .A(n1861), .B(n1860), .Z(n2009) );
  XOR U2709 ( .A(n2216), .B(n2009), .Z(n1956) );
  AND U2710 ( .A(y[652]), .B(x[137]), .Z(n1954) );
  NAND U2711 ( .A(y[653]), .B(x[136]), .Z(n1953) );
  AND U2712 ( .A(x[145]), .B(y[644]), .Z(n1863) );
  NAND U2713 ( .A(y[649]), .B(x[140]), .Z(n1862) );
  XNOR U2714 ( .A(n1863), .B(n1862), .Z(n1959) );
  NAND U2715 ( .A(y[659]), .B(x[130]), .Z(n1960) );
  AND U2716 ( .A(y[658]), .B(x[131]), .Z(n1865) );
  NAND U2717 ( .A(y[648]), .B(x[141]), .Z(n1864) );
  XNOR U2718 ( .A(n1865), .B(n1864), .Z(n1993) );
  NAND U2719 ( .A(y[657]), .B(x[132]), .Z(n1994) );
  XOR U2720 ( .A(n1971), .B(n1970), .Z(n1973) );
  XOR U2721 ( .A(n1972), .B(n1973), .Z(n2023) );
  NAND U2722 ( .A(n1983), .B(n1866), .Z(n1870) );
  NAND U2723 ( .A(n1868), .B(n1867), .Z(n1869) );
  AND U2724 ( .A(n1870), .B(n1869), .Z(n2021) );
  NANDN U2725 ( .A(n1872), .B(n1871), .Z(n1876) );
  NAND U2726 ( .A(n1874), .B(n1873), .Z(n1875) );
  NAND U2727 ( .A(n1876), .B(n1875), .Z(n2020) );
  XNOR U2728 ( .A(n2021), .B(n2020), .Z(n2022) );
  XOR U2729 ( .A(n2023), .B(n2022), .Z(n1949) );
  XOR U2730 ( .A(n1950), .B(n1949), .Z(n1936) );
  NANDN U2731 ( .A(n1878), .B(n1877), .Z(n1882) );
  NAND U2732 ( .A(n1880), .B(n1879), .Z(n1881) );
  NAND U2733 ( .A(n1882), .B(n1881), .Z(n1943) );
  NAND U2734 ( .A(n1884), .B(n1883), .Z(n1888) );
  NANDN U2735 ( .A(n1886), .B(n1885), .Z(n1887) );
  NAND U2736 ( .A(n1888), .B(n1887), .Z(n1942) );
  NAND U2737 ( .A(n1890), .B(n1889), .Z(n1894) );
  NANDN U2738 ( .A(n1892), .B(n1891), .Z(n1893) );
  NAND U2739 ( .A(n1894), .B(n1893), .Z(n1941) );
  XOR U2740 ( .A(n1942), .B(n1941), .Z(n1944) );
  XOR U2741 ( .A(n1943), .B(n1944), .Z(n1935) );
  XOR U2742 ( .A(n1936), .B(n1935), .Z(n1937) );
  XOR U2743 ( .A(n1938), .B(n1937), .Z(n1924) );
  NANDN U2744 ( .A(n1896), .B(n1895), .Z(n1900) );
  NANDN U2745 ( .A(n1898), .B(n1897), .Z(n1899) );
  NAND U2746 ( .A(n1900), .B(n1899), .Z(n1923) );
  XOR U2747 ( .A(n1924), .B(n1923), .Z(n1926) );
  XNOR U2748 ( .A(n1925), .B(n1926), .Z(n2047) );
  NAND U2749 ( .A(n1902), .B(n1901), .Z(n1906) );
  NANDN U2750 ( .A(n1904), .B(n1903), .Z(n1905) );
  AND U2751 ( .A(n1906), .B(n1905), .Z(n2046) );
  NANDN U2752 ( .A(n1908), .B(n1907), .Z(n1912) );
  NAND U2753 ( .A(n1910), .B(n1909), .Z(n1911) );
  AND U2754 ( .A(n1912), .B(n1911), .Z(n2045) );
  XNOR U2755 ( .A(n2047), .B(n2048), .Z(n2041) );
  NAND U2756 ( .A(n1917), .B(n1916), .Z(n1921) );
  NANDN U2757 ( .A(n1919), .B(n1918), .Z(n1920) );
  AND U2758 ( .A(n1921), .B(n1920), .Z(n2039) );
  IV U2759 ( .A(n2039), .Z(n2038) );
  XOR U2760 ( .A(n2040), .B(n2038), .Z(n1922) );
  XNOR U2761 ( .A(n2041), .B(n1922), .Z(N54) );
  NAND U2762 ( .A(n1924), .B(n1923), .Z(n1928) );
  NAND U2763 ( .A(n1926), .B(n1925), .Z(n1927) );
  AND U2764 ( .A(n1928), .B(n1927), .Z(n2055) );
  NANDN U2765 ( .A(n1930), .B(n1929), .Z(n1934) );
  NANDN U2766 ( .A(n1932), .B(n1931), .Z(n1933) );
  AND U2767 ( .A(n1934), .B(n1933), .Z(n2053) );
  NAND U2768 ( .A(n1936), .B(n1935), .Z(n1940) );
  NANDN U2769 ( .A(n1938), .B(n1937), .Z(n1939) );
  AND U2770 ( .A(n1940), .B(n1939), .Z(n2066) );
  NAND U2771 ( .A(n1942), .B(n1941), .Z(n1946) );
  NAND U2772 ( .A(n1944), .B(n1943), .Z(n1945) );
  NAND U2773 ( .A(n1946), .B(n1945), .Z(n2065) );
  XNOR U2774 ( .A(n2066), .B(n2065), .Z(n2068) );
  NANDN U2775 ( .A(n1948), .B(n1947), .Z(n1952) );
  NAND U2776 ( .A(n1950), .B(n1949), .Z(n1951) );
  NAND U2777 ( .A(n1952), .B(n1951), .Z(n2179) );
  NANDN U2778 ( .A(n1954), .B(n1953), .Z(n1958) );
  NANDN U2779 ( .A(n1956), .B(n1955), .Z(n1957) );
  AND U2780 ( .A(n1958), .B(n1957), .Z(n2174) );
  NAND U2781 ( .A(n2665), .B(n2131), .Z(n1962) );
  NANDN U2782 ( .A(n1960), .B(n1959), .Z(n1961) );
  NAND U2783 ( .A(n1962), .B(n1961), .Z(n2103) );
  AND U2784 ( .A(y[657]), .B(x[133]), .Z(n2147) );
  NAND U2785 ( .A(y[645]), .B(x[145]), .Z(n2148) );
  XNOR U2786 ( .A(n2147), .B(n2148), .Z(n2149) );
  NAND U2787 ( .A(x[144]), .B(y[646]), .Z(n2150) );
  XNOR U2788 ( .A(n2149), .B(n2150), .Z(n2102) );
  AND U2789 ( .A(x[146]), .B(y[644]), .Z(n1964) );
  NAND U2790 ( .A(y[650]), .B(x[140]), .Z(n1963) );
  XNOR U2791 ( .A(n1964), .B(n1963), .Z(n2132) );
  NAND U2792 ( .A(x[132]), .B(y[658]), .Z(n2133) );
  XNOR U2793 ( .A(n2132), .B(n2133), .Z(n2101) );
  XOR U2794 ( .A(n2102), .B(n2101), .Z(n2104) );
  XNOR U2795 ( .A(n2103), .B(n2104), .Z(n2171) );
  AND U2796 ( .A(x[147]), .B(y[650]), .Z(n3205) );
  NAND U2797 ( .A(n3205), .B(n1965), .Z(n1969) );
  NAND U2798 ( .A(n1967), .B(n1966), .Z(n1968) );
  AND U2799 ( .A(n1969), .B(n1968), .Z(n2172) );
  XOR U2800 ( .A(n2171), .B(n2172), .Z(n2173) );
  NAND U2801 ( .A(n1971), .B(n1970), .Z(n1975) );
  NAND U2802 ( .A(n1973), .B(n1972), .Z(n1974) );
  AND U2803 ( .A(n1975), .B(n1974), .Z(n2160) );
  NAND U2804 ( .A(n1977), .B(n1976), .Z(n1981) );
  NANDN U2805 ( .A(n1979), .B(n1978), .Z(n1980) );
  NAND U2806 ( .A(n1981), .B(n1980), .Z(n2159) );
  NAND U2807 ( .A(n1983), .B(n1982), .Z(n1987) );
  ANDN U2808 ( .B(n1985), .A(n1984), .Z(n1986) );
  ANDN U2809 ( .B(n1987), .A(n1986), .Z(n2123) );
  AND U2810 ( .A(x[141]), .B(y[649]), .Z(n1989) );
  NAND U2811 ( .A(x[148]), .B(y[642]), .Z(n1988) );
  XNOR U2812 ( .A(n1989), .B(n1988), .Z(n2143) );
  NAND U2813 ( .A(x[130]), .B(y[660]), .Z(n2144) );
  XNOR U2814 ( .A(n2143), .B(n2144), .Z(n2121) );
  AND U2815 ( .A(y[647]), .B(x[143]), .Z(n1991) );
  NAND U2816 ( .A(x[134]), .B(y[656]), .Z(n1990) );
  XNOR U2817 ( .A(n1991), .B(n1990), .Z(n2155) );
  XOR U2818 ( .A(n2121), .B(n2120), .Z(n2122) );
  XNOR U2819 ( .A(n2123), .B(n2122), .Z(n2166) );
  AND U2820 ( .A(x[141]), .B(y[658]), .Z(n3460) );
  NAND U2821 ( .A(n1992), .B(n3460), .Z(n1996) );
  NANDN U2822 ( .A(n1994), .B(n1993), .Z(n1995) );
  AND U2823 ( .A(n1996), .B(n1995), .Z(n2092) );
  AND U2824 ( .A(y[661]), .B(x[129]), .Z(n2115) );
  XOR U2825 ( .A(n2116), .B(n2115), .Z(n2114) );
  ANDN U2826 ( .B(o[21]), .A(n1997), .Z(n2113) );
  XOR U2827 ( .A(n2114), .B(n2113), .Z(n2090) );
  AND U2828 ( .A(x[142]), .B(y[648]), .Z(n2107) );
  NAND U2829 ( .A(y[659]), .B(x[131]), .Z(n2108) );
  XNOR U2830 ( .A(n2107), .B(n2108), .Z(n2109) );
  NAND U2831 ( .A(x[147]), .B(y[643]), .Z(n2110) );
  XNOR U2832 ( .A(n2109), .B(n2110), .Z(n2089) );
  XOR U2833 ( .A(n2090), .B(n2089), .Z(n2091) );
  XOR U2834 ( .A(n2166), .B(n2165), .Z(n2168) );
  NANDN U2835 ( .A(n1999), .B(n1998), .Z(n2003) );
  NAND U2836 ( .A(n2001), .B(n2000), .Z(n2002) );
  AND U2837 ( .A(n2003), .B(n2002), .Z(n2084) );
  AND U2838 ( .A(y[651]), .B(x[146]), .Z(n3208) );
  NAND U2839 ( .A(n3208), .B(n2004), .Z(n2008) );
  NANDN U2840 ( .A(n2006), .B(n2005), .Z(n2007) );
  NAND U2841 ( .A(n2008), .B(n2007), .Z(n2083) );
  AND U2842 ( .A(y[655]), .B(x[142]), .Z(n3218) );
  NAND U2843 ( .A(n3218), .B(n2154), .Z(n2011) );
  NAND U2844 ( .A(n2216), .B(n2009), .Z(n2010) );
  AND U2845 ( .A(n2011), .B(n2010), .Z(n2098) );
  AND U2846 ( .A(y[662]), .B(x[128]), .Z(n2136) );
  NAND U2847 ( .A(x[150]), .B(y[640]), .Z(n2137) );
  XNOR U2848 ( .A(n2136), .B(n2137), .Z(n2139) );
  NAND U2849 ( .A(y[641]), .B(x[149]), .Z(n2153) );
  XNOR U2850 ( .A(o[22]), .B(n2153), .Z(n2138) );
  XOR U2851 ( .A(n2139), .B(n2138), .Z(n2096) );
  NAND U2852 ( .A(y[655]), .B(x[135]), .Z(n2012) );
  XNOR U2853 ( .A(n2013), .B(n2012), .Z(n2126) );
  XOR U2854 ( .A(n2096), .B(n2095), .Z(n2097) );
  XOR U2855 ( .A(n2086), .B(n2085), .Z(n2167) );
  XOR U2856 ( .A(n2168), .B(n2167), .Z(n2161) );
  XOR U2857 ( .A(n2162), .B(n2161), .Z(n2177) );
  XOR U2858 ( .A(n2179), .B(n2180), .Z(n2074) );
  NANDN U2859 ( .A(n2015), .B(n2014), .Z(n2019) );
  NAND U2860 ( .A(n2017), .B(n2016), .Z(n2018) );
  AND U2861 ( .A(n2019), .B(n2018), .Z(n2080) );
  NANDN U2862 ( .A(n2021), .B(n2020), .Z(n2025) );
  NAND U2863 ( .A(n2023), .B(n2022), .Z(n2024) );
  AND U2864 ( .A(n2025), .B(n2024), .Z(n2078) );
  NAND U2865 ( .A(n2027), .B(n2026), .Z(n2031) );
  NANDN U2866 ( .A(n2029), .B(n2028), .Z(n2030) );
  NAND U2867 ( .A(n2031), .B(n2030), .Z(n2077) );
  NANDN U2868 ( .A(n2033), .B(n2032), .Z(n2037) );
  NAND U2869 ( .A(n2035), .B(n2034), .Z(n2036) );
  NAND U2870 ( .A(n2037), .B(n2036), .Z(n2072) );
  XNOR U2871 ( .A(n2071), .B(n2072), .Z(n2073) );
  XOR U2872 ( .A(n2074), .B(n2073), .Z(n2067) );
  XOR U2873 ( .A(n2068), .B(n2067), .Z(n2052) );
  XNOR U2874 ( .A(n2055), .B(n2054), .Z(n2061) );
  OR U2875 ( .A(n2040), .B(n2038), .Z(n2044) );
  ANDN U2876 ( .B(n2040), .A(n2039), .Z(n2042) );
  OR U2877 ( .A(n2042), .B(n2041), .Z(n2043) );
  AND U2878 ( .A(n2044), .B(n2043), .Z(n2060) );
  NANDN U2879 ( .A(n2046), .B(n2045), .Z(n2050) );
  NAND U2880 ( .A(n2048), .B(n2047), .Z(n2049) );
  NAND U2881 ( .A(n2050), .B(n2049), .Z(n2059) );
  IV U2882 ( .A(n2059), .Z(n2058) );
  XOR U2883 ( .A(n2060), .B(n2058), .Z(n2051) );
  XNOR U2884 ( .A(n2061), .B(n2051), .Z(N55) );
  NANDN U2885 ( .A(n2053), .B(n2052), .Z(n2057) );
  NAND U2886 ( .A(n2055), .B(n2054), .Z(n2056) );
  NAND U2887 ( .A(n2057), .B(n2056), .Z(n2191) );
  IV U2888 ( .A(n2191), .Z(n2190) );
  OR U2889 ( .A(n2060), .B(n2058), .Z(n2064) );
  ANDN U2890 ( .B(n2060), .A(n2059), .Z(n2062) );
  OR U2891 ( .A(n2062), .B(n2061), .Z(n2063) );
  AND U2892 ( .A(n2064), .B(n2063), .Z(n2192) );
  NANDN U2893 ( .A(n2066), .B(n2065), .Z(n2070) );
  NAND U2894 ( .A(n2068), .B(n2067), .Z(n2069) );
  AND U2895 ( .A(n2070), .B(n2069), .Z(n2187) );
  NANDN U2896 ( .A(n2072), .B(n2071), .Z(n2076) );
  NAND U2897 ( .A(n2074), .B(n2073), .Z(n2075) );
  AND U2898 ( .A(n2076), .B(n2075), .Z(n2185) );
  NANDN U2899 ( .A(n2078), .B(n2077), .Z(n2082) );
  NANDN U2900 ( .A(n2080), .B(n2079), .Z(n2081) );
  AND U2901 ( .A(n2082), .B(n2081), .Z(n2312) );
  NANDN U2902 ( .A(n2084), .B(n2083), .Z(n2088) );
  NAND U2903 ( .A(n2086), .B(n2085), .Z(n2087) );
  AND U2904 ( .A(n2088), .B(n2087), .Z(n2306) );
  NAND U2905 ( .A(n2090), .B(n2089), .Z(n2094) );
  NANDN U2906 ( .A(n2092), .B(n2091), .Z(n2093) );
  AND U2907 ( .A(n2094), .B(n2093), .Z(n2304) );
  NAND U2908 ( .A(n2096), .B(n2095), .Z(n2100) );
  NANDN U2909 ( .A(n2098), .B(n2097), .Z(n2099) );
  NAND U2910 ( .A(n2100), .B(n2099), .Z(n2303) );
  NAND U2911 ( .A(n2102), .B(n2101), .Z(n2106) );
  NAND U2912 ( .A(n2104), .B(n2103), .Z(n2105) );
  AND U2913 ( .A(n2106), .B(n2105), .Z(n2322) );
  NANDN U2914 ( .A(n2108), .B(n2107), .Z(n2112) );
  NANDN U2915 ( .A(n2110), .B(n2109), .Z(n2111) );
  AND U2916 ( .A(n2112), .B(n2111), .Z(n2250) );
  AND U2917 ( .A(n2114), .B(n2113), .Z(n2118) );
  NAND U2918 ( .A(n2116), .B(n2115), .Z(n2117) );
  NANDN U2919 ( .A(n2118), .B(n2117), .Z(n2249) );
  XNOR U2920 ( .A(n2250), .B(n2249), .Z(n2252) );
  NAND U2921 ( .A(x[135]), .B(y[656]), .Z(n2119) );
  XNOR U2922 ( .A(n2381), .B(n2119), .Z(n2217) );
  NAND U2923 ( .A(x[138]), .B(y[653]), .Z(n2256) );
  XNOR U2924 ( .A(n2255), .B(n2256), .Z(n2258) );
  AND U2925 ( .A(y[657]), .B(x[134]), .Z(n2208) );
  NAND U2926 ( .A(x[143]), .B(y[648]), .Z(n2209) );
  XNOR U2927 ( .A(n2208), .B(n2209), .Z(n2210) );
  NAND U2928 ( .A(x[139]), .B(y[652]), .Z(n2211) );
  XNOR U2929 ( .A(n2210), .B(n2211), .Z(n2257) );
  XOR U2930 ( .A(n2258), .B(n2257), .Z(n2251) );
  XOR U2931 ( .A(n2252), .B(n2251), .Z(n2321) );
  XOR U2932 ( .A(n2324), .B(n2323), .Z(n2310) );
  NAND U2933 ( .A(n2121), .B(n2120), .Z(n2125) );
  NANDN U2934 ( .A(n2123), .B(n2122), .Z(n2124) );
  AND U2935 ( .A(n2125), .B(n2124), .Z(n2244) );
  NANDN U2936 ( .A(n2218), .B(n2216), .Z(n2129) );
  NANDN U2937 ( .A(n2127), .B(n2126), .Z(n2128) );
  AND U2938 ( .A(n2129), .B(n2128), .Z(n2294) );
  AND U2939 ( .A(y[663]), .B(x[128]), .Z(n2227) );
  NAND U2940 ( .A(x[151]), .B(y[640]), .Z(n2228) );
  XNOR U2941 ( .A(n2227), .B(n2228), .Z(n2230) );
  NAND U2942 ( .A(y[641]), .B(x[150]), .Z(n2207) );
  XNOR U2943 ( .A(o[23]), .B(n2207), .Z(n2229) );
  XOR U2944 ( .A(n2230), .B(n2229), .Z(n2292) );
  AND U2945 ( .A(x[148]), .B(y[643]), .Z(n2870) );
  NAND U2946 ( .A(y[647]), .B(x[144]), .Z(n2130) );
  XNOR U2947 ( .A(n2870), .B(n2130), .Z(n2203) );
  NAND U2948 ( .A(y[644]), .B(x[147]), .Z(n2204) );
  XNOR U2949 ( .A(n2203), .B(n2204), .Z(n2291) );
  XOR U2950 ( .A(n2292), .B(n2291), .Z(n2293) );
  AND U2951 ( .A(x[146]), .B(y[650]), .Z(n3013) );
  NAND U2952 ( .A(n3013), .B(n2131), .Z(n2135) );
  NANDN U2953 ( .A(n2133), .B(n2132), .Z(n2134) );
  AND U2954 ( .A(n2135), .B(n2134), .Z(n2280) );
  NANDN U2955 ( .A(n2137), .B(n2136), .Z(n2141) );
  NAND U2956 ( .A(n2139), .B(n2138), .Z(n2140) );
  NAND U2957 ( .A(n2141), .B(n2140), .Z(n2279) );
  XOR U2958 ( .A(n2282), .B(n2281), .Z(n2243) );
  XNOR U2959 ( .A(n2244), .B(n2243), .Z(n2246) );
  AND U2960 ( .A(y[649]), .B(x[148]), .Z(n3229) );
  NAND U2961 ( .A(n3229), .B(n2142), .Z(n2146) );
  NANDN U2962 ( .A(n2144), .B(n2143), .Z(n2145) );
  AND U2963 ( .A(n2146), .B(n2145), .Z(n2238) );
  NANDN U2964 ( .A(n2148), .B(n2147), .Z(n2152) );
  NANDN U2965 ( .A(n2150), .B(n2149), .Z(n2151) );
  AND U2966 ( .A(n2152), .B(n2151), .Z(n2300) );
  AND U2967 ( .A(y[650]), .B(x[141]), .Z(n2273) );
  NAND U2968 ( .A(y[661]), .B(x[130]), .Z(n2274) );
  XNOR U2969 ( .A(n2273), .B(n2274), .Z(n2275) );
  NAND U2970 ( .A(y[642]), .B(x[149]), .Z(n2276) );
  XNOR U2971 ( .A(n2275), .B(n2276), .Z(n2298) );
  AND U2972 ( .A(y[651]), .B(x[140]), .Z(n2221) );
  NAND U2973 ( .A(y[662]), .B(x[129]), .Z(n2222) );
  XNOR U2974 ( .A(n2221), .B(n2222), .Z(n2224) );
  ANDN U2975 ( .B(o[22]), .A(n2153), .Z(n2223) );
  XOR U2976 ( .A(n2224), .B(n2223), .Z(n2297) );
  XOR U2977 ( .A(n2298), .B(n2297), .Z(n2299) );
  XNOR U2978 ( .A(n2238), .B(n2237), .Z(n2240) );
  AND U2979 ( .A(y[656]), .B(x[143]), .Z(n3359) );
  NAND U2980 ( .A(n3359), .B(n2154), .Z(n2158) );
  NANDN U2981 ( .A(n2156), .B(n2155), .Z(n2157) );
  AND U2982 ( .A(n2158), .B(n2157), .Z(n2288) );
  AND U2983 ( .A(y[649]), .B(x[142]), .Z(n2267) );
  NAND U2984 ( .A(x[131]), .B(y[660]), .Z(n2268) );
  XNOR U2985 ( .A(n2267), .B(n2268), .Z(n2269) );
  NAND U2986 ( .A(y[659]), .B(x[132]), .Z(n2270) );
  XNOR U2987 ( .A(n2269), .B(n2270), .Z(n2286) );
  AND U2988 ( .A(x[133]), .B(y[658]), .Z(n2261) );
  NAND U2989 ( .A(y[645]), .B(x[146]), .Z(n2262) );
  XNOR U2990 ( .A(n2261), .B(n2262), .Z(n2263) );
  NAND U2991 ( .A(x[145]), .B(y[646]), .Z(n2264) );
  XNOR U2992 ( .A(n2263), .B(n2264), .Z(n2285) );
  XOR U2993 ( .A(n2286), .B(n2285), .Z(n2287) );
  XOR U2994 ( .A(n2240), .B(n2239), .Z(n2245) );
  XOR U2995 ( .A(n2246), .B(n2245), .Z(n2309) );
  XOR U2996 ( .A(n2310), .B(n2309), .Z(n2311) );
  NANDN U2997 ( .A(n2160), .B(n2159), .Z(n2164) );
  NAND U2998 ( .A(n2162), .B(n2161), .Z(n2163) );
  AND U2999 ( .A(n2164), .B(n2163), .Z(n2318) );
  NAND U3000 ( .A(n2166), .B(n2165), .Z(n2170) );
  NAND U3001 ( .A(n2168), .B(n2167), .Z(n2169) );
  AND U3002 ( .A(n2170), .B(n2169), .Z(n2316) );
  NAND U3003 ( .A(n2172), .B(n2171), .Z(n2176) );
  NANDN U3004 ( .A(n2174), .B(n2173), .Z(n2175) );
  AND U3005 ( .A(n2176), .B(n2175), .Z(n2315) );
  NANDN U3006 ( .A(n2178), .B(n2177), .Z(n2182) );
  NAND U3007 ( .A(n2180), .B(n2179), .Z(n2181) );
  AND U3008 ( .A(n2182), .B(n2181), .Z(n2197) );
  XOR U3009 ( .A(n2185), .B(n2184), .Z(n2186) );
  XOR U3010 ( .A(n2187), .B(n2186), .Z(n2193) );
  XNOR U3011 ( .A(n2192), .B(n2193), .Z(n2183) );
  XOR U3012 ( .A(n2190), .B(n2183), .Z(N56) );
  NAND U3013 ( .A(n2185), .B(n2184), .Z(n2189) );
  NAND U3014 ( .A(n2187), .B(n2186), .Z(n2188) );
  NAND U3015 ( .A(n2189), .B(n2188), .Z(n2461) );
  IV U3016 ( .A(n2461), .Z(n2459) );
  OR U3017 ( .A(n2192), .B(n2190), .Z(n2196) );
  ANDN U3018 ( .B(n2192), .A(n2191), .Z(n2194) );
  OR U3019 ( .A(n2194), .B(n2193), .Z(n2195) );
  AND U3020 ( .A(n2196), .B(n2195), .Z(n2460) );
  NANDN U3021 ( .A(n2198), .B(n2197), .Z(n2202) );
  NANDN U3022 ( .A(n2200), .B(n2199), .Z(n2201) );
  AND U3023 ( .A(n2202), .B(n2201), .Z(n2468) );
  AND U3024 ( .A(y[647]), .B(x[148]), .Z(n2763) );
  AND U3025 ( .A(x[144]), .B(y[643]), .Z(n2352) );
  NAND U3026 ( .A(n2763), .B(n2352), .Z(n2206) );
  NANDN U3027 ( .A(n2204), .B(n2203), .Z(n2205) );
  AND U3028 ( .A(n2206), .B(n2205), .Z(n2372) );
  AND U3029 ( .A(y[642]), .B(x[150]), .Z(n2391) );
  XOR U3030 ( .A(n2392), .B(n2391), .Z(n2394) );
  NAND U3031 ( .A(y[662]), .B(x[130]), .Z(n2393) );
  AND U3032 ( .A(x[129]), .B(y[663]), .Z(n2399) );
  XOR U3033 ( .A(n2400), .B(n2399), .Z(n2398) );
  ANDN U3034 ( .B(o[23]), .A(n2207), .Z(n2397) );
  XOR U3035 ( .A(n2398), .B(n2397), .Z(n2369) );
  XOR U3036 ( .A(n2370), .B(n2369), .Z(n2371) );
  XNOR U3037 ( .A(n2372), .B(n2371), .Z(n2430) );
  NANDN U3038 ( .A(n2209), .B(n2208), .Z(n2213) );
  NANDN U3039 ( .A(n2211), .B(n2210), .Z(n2212) );
  AND U3040 ( .A(n2213), .B(n2212), .Z(n2366) );
  AND U3041 ( .A(y[643]), .B(x[149]), .Z(n2215) );
  NAND U3042 ( .A(y[648]), .B(x[144]), .Z(n2214) );
  XNOR U3043 ( .A(n2215), .B(n2214), .Z(n2353) );
  NAND U3044 ( .A(y[659]), .B(x[133]), .Z(n2354) );
  XNOR U3045 ( .A(n2353), .B(n2354), .Z(n2364) );
  AND U3046 ( .A(x[134]), .B(y[658]), .Z(n2750) );
  NAND U3047 ( .A(y[644]), .B(x[148]), .Z(n2584) );
  XNOR U3048 ( .A(n2750), .B(n2584), .Z(n2359) );
  NAND U3049 ( .A(y[645]), .B(x[147]), .Z(n2360) );
  XNOR U3050 ( .A(n2359), .B(n2360), .Z(n2363) );
  XOR U3051 ( .A(n2364), .B(n2363), .Z(n2365) );
  XNOR U3052 ( .A(n2366), .B(n2365), .Z(n2343) );
  NANDN U3053 ( .A(n2509), .B(n2216), .Z(n2220) );
  NANDN U3054 ( .A(n2218), .B(n2217), .Z(n2219) );
  AND U3055 ( .A(n2220), .B(n2219), .Z(n2341) );
  NANDN U3056 ( .A(n2222), .B(n2221), .Z(n2226) );
  NAND U3057 ( .A(n2224), .B(n2223), .Z(n2225) );
  NAND U3058 ( .A(n2226), .B(n2225), .Z(n2340) );
  XNOR U3059 ( .A(n2341), .B(n2340), .Z(n2342) );
  XOR U3060 ( .A(n2343), .B(n2342), .Z(n2429) );
  XOR U3061 ( .A(n2430), .B(n2429), .Z(n2432) );
  NANDN U3062 ( .A(n2228), .B(n2227), .Z(n2232) );
  NAND U3063 ( .A(n2230), .B(n2229), .Z(n2231) );
  AND U3064 ( .A(n2232), .B(n2231), .Z(n2424) );
  AND U3065 ( .A(y[661]), .B(x[131]), .Z(n2411) );
  XOR U3066 ( .A(n2412), .B(n2411), .Z(n2414) );
  NAND U3067 ( .A(x[132]), .B(y[660]), .Z(n2413) );
  XNOR U3068 ( .A(n2414), .B(n2413), .Z(n2423) );
  XNOR U3069 ( .A(n2424), .B(n2423), .Z(n2426) );
  AND U3070 ( .A(x[137]), .B(y[655]), .Z(n2234) );
  NAND U3071 ( .A(y[654]), .B(x[138]), .Z(n2233) );
  XNOR U3072 ( .A(n2234), .B(n2233), .Z(n2383) );
  AND U3073 ( .A(x[142]), .B(y[650]), .Z(n2236) );
  NAND U3074 ( .A(x[136]), .B(y[656]), .Z(n2235) );
  XNOR U3075 ( .A(n2236), .B(n2235), .Z(n2387) );
  NAND U3076 ( .A(x[139]), .B(y[653]), .Z(n2388) );
  XNOR U3077 ( .A(n2387), .B(n2388), .Z(n2382) );
  XOR U3078 ( .A(n2383), .B(n2382), .Z(n2425) );
  XOR U3079 ( .A(n2426), .B(n2425), .Z(n2431) );
  XOR U3080 ( .A(n2432), .B(n2431), .Z(n2442) );
  NANDN U3081 ( .A(n2238), .B(n2237), .Z(n2242) );
  NAND U3082 ( .A(n2240), .B(n2239), .Z(n2241) );
  AND U3083 ( .A(n2242), .B(n2241), .Z(n2441) );
  XNOR U3084 ( .A(n2442), .B(n2441), .Z(n2443) );
  NANDN U3085 ( .A(n2244), .B(n2243), .Z(n2248) );
  NAND U3086 ( .A(n2246), .B(n2245), .Z(n2247) );
  NAND U3087 ( .A(n2248), .B(n2247), .Z(n2444) );
  XNOR U3088 ( .A(n2443), .B(n2444), .Z(n2450) );
  NANDN U3089 ( .A(n2250), .B(n2249), .Z(n2254) );
  NAND U3090 ( .A(n2252), .B(n2251), .Z(n2253) );
  AND U3091 ( .A(n2254), .B(n2253), .Z(n2438) );
  NANDN U3092 ( .A(n2256), .B(n2255), .Z(n2260) );
  NAND U3093 ( .A(n2258), .B(n2257), .Z(n2259) );
  AND U3094 ( .A(n2260), .B(n2259), .Z(n2436) );
  NANDN U3095 ( .A(n2262), .B(n2261), .Z(n2266) );
  NANDN U3096 ( .A(n2264), .B(n2263), .Z(n2265) );
  AND U3097 ( .A(n2266), .B(n2265), .Z(n2349) );
  AND U3098 ( .A(y[664]), .B(x[128]), .Z(n2417) );
  NAND U3099 ( .A(y[640]), .B(x[152]), .Z(n2418) );
  XNOR U3100 ( .A(n2417), .B(n2418), .Z(n2420) );
  NAND U3101 ( .A(y[641]), .B(x[151]), .Z(n2410) );
  XNOR U3102 ( .A(o[24]), .B(n2410), .Z(n2419) );
  XOR U3103 ( .A(n2420), .B(n2419), .Z(n2347) );
  AND U3104 ( .A(y[657]), .B(x[135]), .Z(n2403) );
  NAND U3105 ( .A(y[646]), .B(x[146]), .Z(n2404) );
  NAND U3106 ( .A(x[145]), .B(y[647]), .Z(n2406) );
  XOR U3107 ( .A(n2347), .B(n2346), .Z(n2348) );
  XNOR U3108 ( .A(n2349), .B(n2348), .Z(n2337) );
  NANDN U3109 ( .A(n2268), .B(n2267), .Z(n2272) );
  NANDN U3110 ( .A(n2270), .B(n2269), .Z(n2271) );
  AND U3111 ( .A(n2272), .B(n2271), .Z(n2335) );
  NANDN U3112 ( .A(n2274), .B(n2273), .Z(n2278) );
  NANDN U3113 ( .A(n2276), .B(n2275), .Z(n2277) );
  NAND U3114 ( .A(n2278), .B(n2277), .Z(n2334) );
  XNOR U3115 ( .A(n2335), .B(n2334), .Z(n2336) );
  XOR U3116 ( .A(n2337), .B(n2336), .Z(n2435) );
  XNOR U3117 ( .A(n2436), .B(n2435), .Z(n2437) );
  XOR U3118 ( .A(n2438), .B(n2437), .Z(n2377) );
  NANDN U3119 ( .A(n2280), .B(n2279), .Z(n2284) );
  NAND U3120 ( .A(n2282), .B(n2281), .Z(n2283) );
  AND U3121 ( .A(n2284), .B(n2283), .Z(n2331) );
  NAND U3122 ( .A(n2286), .B(n2285), .Z(n2290) );
  NANDN U3123 ( .A(n2288), .B(n2287), .Z(n2289) );
  AND U3124 ( .A(n2290), .B(n2289), .Z(n2328) );
  NAND U3125 ( .A(n2292), .B(n2291), .Z(n2296) );
  NANDN U3126 ( .A(n2294), .B(n2293), .Z(n2295) );
  NAND U3127 ( .A(n2296), .B(n2295), .Z(n2329) );
  XNOR U3128 ( .A(n2328), .B(n2329), .Z(n2330) );
  XOR U3129 ( .A(n2331), .B(n2330), .Z(n2375) );
  NAND U3130 ( .A(n2298), .B(n2297), .Z(n2302) );
  NANDN U3131 ( .A(n2300), .B(n2299), .Z(n2301) );
  NAND U3132 ( .A(n2302), .B(n2301), .Z(n2376) );
  XNOR U3133 ( .A(n2375), .B(n2376), .Z(n2378) );
  XOR U3134 ( .A(n2377), .B(n2378), .Z(n2447) );
  NANDN U3135 ( .A(n2304), .B(n2303), .Z(n2308) );
  NANDN U3136 ( .A(n2306), .B(n2305), .Z(n2307) );
  NAND U3137 ( .A(n2308), .B(n2307), .Z(n2448) );
  XNOR U3138 ( .A(n2450), .B(n2449), .Z(n2466) );
  NAND U3139 ( .A(n2310), .B(n2309), .Z(n2314) );
  NANDN U3140 ( .A(n2312), .B(n2311), .Z(n2313) );
  AND U3141 ( .A(n2314), .B(n2313), .Z(n2456) );
  NANDN U3142 ( .A(n2316), .B(n2315), .Z(n2320) );
  NANDN U3143 ( .A(n2318), .B(n2317), .Z(n2319) );
  AND U3144 ( .A(n2320), .B(n2319), .Z(n2454) );
  NANDN U3145 ( .A(n2322), .B(n2321), .Z(n2326) );
  NAND U3146 ( .A(n2324), .B(n2323), .Z(n2325) );
  NAND U3147 ( .A(n2326), .B(n2325), .Z(n2453) );
  XOR U3148 ( .A(n2466), .B(n2467), .Z(n2469) );
  XNOR U3149 ( .A(n2468), .B(n2469), .Z(n2462) );
  XNOR U3150 ( .A(n2460), .B(n2462), .Z(n2327) );
  XOR U3151 ( .A(n2459), .B(n2327), .Z(N57) );
  NANDN U3152 ( .A(n2329), .B(n2328), .Z(n2333) );
  NAND U3153 ( .A(n2331), .B(n2330), .Z(n2332) );
  AND U3154 ( .A(n2333), .B(n2332), .Z(n2480) );
  NANDN U3155 ( .A(n2335), .B(n2334), .Z(n2339) );
  NAND U3156 ( .A(n2337), .B(n2336), .Z(n2338) );
  AND U3157 ( .A(n2339), .B(n2338), .Z(n2498) );
  NANDN U3158 ( .A(n2341), .B(n2340), .Z(n2345) );
  NAND U3159 ( .A(n2343), .B(n2342), .Z(n2344) );
  NAND U3160 ( .A(n2345), .B(n2344), .Z(n2497) );
  XNOR U3161 ( .A(n2498), .B(n2497), .Z(n2500) );
  NAND U3162 ( .A(n2347), .B(n2346), .Z(n2351) );
  NANDN U3163 ( .A(n2349), .B(n2348), .Z(n2350) );
  AND U3164 ( .A(n2351), .B(n2350), .Z(n2530) );
  AND U3165 ( .A(x[149]), .B(y[648]), .Z(n3469) );
  NAND U3166 ( .A(n3469), .B(n2352), .Z(n2356) );
  NANDN U3167 ( .A(n2354), .B(n2353), .Z(n2355) );
  AND U3168 ( .A(n2356), .B(n2355), .Z(n2604) );
  NAND U3169 ( .A(x[150]), .B(y[643]), .Z(n2573) );
  NAND U3170 ( .A(x[133]), .B(y[660]), .Z(n2572) );
  NAND U3171 ( .A(x[145]), .B(y[648]), .Z(n2571) );
  XNOR U3172 ( .A(n2572), .B(n2571), .Z(n2574) );
  XOR U3173 ( .A(n2573), .B(n2574), .Z(n2601) );
  AND U3174 ( .A(x[148]), .B(y[645]), .Z(n2358) );
  NAND U3175 ( .A(x[149]), .B(y[644]), .Z(n2357) );
  XNOR U3176 ( .A(n2358), .B(n2357), .Z(n2586) );
  AND U3177 ( .A(y[646]), .B(x[147]), .Z(n2585) );
  XOR U3178 ( .A(n2586), .B(n2585), .Z(n2602) );
  XOR U3179 ( .A(n2601), .B(n2602), .Z(n2603) );
  XOR U3180 ( .A(n2604), .B(n2603), .Z(n2528) );
  NANDN U3181 ( .A(n2584), .B(n2750), .Z(n2362) );
  NANDN U3182 ( .A(n2360), .B(n2359), .Z(n2361) );
  AND U3183 ( .A(n2362), .B(n2361), .Z(n2610) );
  NAND U3184 ( .A(x[143]), .B(y[650]), .Z(n2591) );
  NAND U3185 ( .A(x[146]), .B(y[647]), .Z(n2590) );
  NAND U3186 ( .A(y[659]), .B(x[134]), .Z(n2589) );
  XNOR U3187 ( .A(n2590), .B(n2589), .Z(n2592) );
  XOR U3188 ( .A(n2591), .B(n2592), .Z(n2608) );
  NAND U3189 ( .A(y[642]), .B(x[151]), .Z(n2567) );
  NAND U3190 ( .A(y[661]), .B(x[132]), .Z(n2566) );
  NAND U3191 ( .A(x[144]), .B(y[649]), .Z(n2565) );
  XNOR U3192 ( .A(n2566), .B(n2565), .Z(n2568) );
  XOR U3193 ( .A(n2567), .B(n2568), .Z(n2607) );
  XOR U3194 ( .A(n2608), .B(n2607), .Z(n2609) );
  XOR U3195 ( .A(n2610), .B(n2609), .Z(n2527) );
  XOR U3196 ( .A(n2528), .B(n2527), .Z(n2529) );
  XOR U3197 ( .A(n2530), .B(n2529), .Z(n2542) );
  NAND U3198 ( .A(n2364), .B(n2363), .Z(n2368) );
  NANDN U3199 ( .A(n2366), .B(n2365), .Z(n2367) );
  AND U3200 ( .A(n2368), .B(n2367), .Z(n2540) );
  NAND U3201 ( .A(n2370), .B(n2369), .Z(n2374) );
  NANDN U3202 ( .A(n2372), .B(n2371), .Z(n2373) );
  NAND U3203 ( .A(n2374), .B(n2373), .Z(n2539) );
  XNOR U3204 ( .A(n2540), .B(n2539), .Z(n2541) );
  XNOR U3205 ( .A(n2542), .B(n2541), .Z(n2499) );
  XNOR U3206 ( .A(n2500), .B(n2499), .Z(n2479) );
  NANDN U3207 ( .A(n2376), .B(n2375), .Z(n2380) );
  NAND U3208 ( .A(n2378), .B(n2377), .Z(n2379) );
  NAND U3209 ( .A(n2380), .B(n2379), .Z(n2481) );
  XOR U3210 ( .A(n2482), .B(n2481), .Z(n2476) );
  NANDN U3211 ( .A(n2409), .B(n2381), .Z(n2385) );
  NAND U3212 ( .A(n2383), .B(n2382), .Z(n2384) );
  AND U3213 ( .A(n2385), .B(n2384), .Z(n2534) );
  AND U3214 ( .A(y[656]), .B(x[142]), .Z(n3407) );
  NAND U3215 ( .A(n3407), .B(n2386), .Z(n2390) );
  NANDN U3216 ( .A(n2388), .B(n2387), .Z(n2389) );
  NAND U3217 ( .A(n2390), .B(n2389), .Z(n2561) );
  NAND U3218 ( .A(x[139]), .B(y[654]), .Z(n2580) );
  NAND U3219 ( .A(x[140]), .B(y[653]), .Z(n2579) );
  NAND U3220 ( .A(x[135]), .B(y[658]), .Z(n2578) );
  XOR U3221 ( .A(n2579), .B(n2578), .Z(n2581) );
  XOR U3222 ( .A(n2580), .B(n2581), .Z(n2560) );
  NAND U3223 ( .A(y[641]), .B(x[152]), .Z(n2577) );
  XNOR U3224 ( .A(o[25]), .B(n2577), .Z(n2548) );
  AND U3225 ( .A(y[664]), .B(x[129]), .Z(n2547) );
  XOR U3226 ( .A(n2548), .B(n2547), .Z(n2550) );
  AND U3227 ( .A(x[141]), .B(y[652]), .Z(n2549) );
  XOR U3228 ( .A(n2550), .B(n2549), .Z(n2559) );
  XNOR U3229 ( .A(n2560), .B(n2559), .Z(n2562) );
  XOR U3230 ( .A(n2561), .B(n2562), .Z(n2533) );
  XNOR U3231 ( .A(n2534), .B(n2533), .Z(n2536) );
  NAND U3232 ( .A(n2392), .B(n2391), .Z(n2396) );
  ANDN U3233 ( .B(n2394), .A(n2393), .Z(n2395) );
  ANDN U3234 ( .B(n2396), .A(n2395), .Z(n2522) );
  AND U3235 ( .A(n2398), .B(n2397), .Z(n2402) );
  NAND U3236 ( .A(n2400), .B(n2399), .Z(n2401) );
  NANDN U3237 ( .A(n2402), .B(n2401), .Z(n2521) );
  NANDN U3238 ( .A(n2404), .B(n2403), .Z(n2408) );
  NANDN U3239 ( .A(n2406), .B(n2405), .Z(n2407) );
  AND U3240 ( .A(n2408), .B(n2407), .Z(n2518) );
  NAND U3241 ( .A(y[657]), .B(x[136]), .Z(n2511) );
  XNOR U3242 ( .A(n2509), .B(n2409), .Z(n2512) );
  XOR U3243 ( .A(n2511), .B(n2512), .Z(n2516) );
  NANDN U3244 ( .A(n2410), .B(o[24]), .Z(n2505) );
  NAND U3245 ( .A(x[153]), .B(y[640]), .Z(n2504) );
  NAND U3246 ( .A(y[665]), .B(x[128]), .Z(n2503) );
  XNOR U3247 ( .A(n2504), .B(n2503), .Z(n2506) );
  XOR U3248 ( .A(n2505), .B(n2506), .Z(n2515) );
  XOR U3249 ( .A(n2516), .B(n2515), .Z(n2517) );
  XOR U3250 ( .A(n2524), .B(n2523), .Z(n2535) );
  XOR U3251 ( .A(n2536), .B(n2535), .Z(n2494) );
  NAND U3252 ( .A(n2412), .B(n2411), .Z(n2416) );
  ANDN U3253 ( .B(n2414), .A(n2413), .Z(n2415) );
  ANDN U3254 ( .B(n2416), .A(n2415), .Z(n2598) );
  NANDN U3255 ( .A(n2418), .B(n2417), .Z(n2422) );
  NAND U3256 ( .A(n2420), .B(n2419), .Z(n2421) );
  AND U3257 ( .A(n2422), .B(n2421), .Z(n2596) );
  AND U3258 ( .A(y[651]), .B(x[142]), .Z(n2554) );
  AND U3259 ( .A(x[130]), .B(y[663]), .Z(n2553) );
  XOR U3260 ( .A(n2554), .B(n2553), .Z(n2556) );
  AND U3261 ( .A(y[662]), .B(x[131]), .Z(n2555) );
  XOR U3262 ( .A(n2556), .B(n2555), .Z(n2595) );
  XNOR U3263 ( .A(n2596), .B(n2595), .Z(n2597) );
  XNOR U3264 ( .A(n2598), .B(n2597), .Z(n2492) );
  NANDN U3265 ( .A(n2424), .B(n2423), .Z(n2428) );
  NAND U3266 ( .A(n2426), .B(n2425), .Z(n2427) );
  AND U3267 ( .A(n2428), .B(n2427), .Z(n2491) );
  XNOR U3268 ( .A(n2492), .B(n2491), .Z(n2493) );
  XNOR U3269 ( .A(n2494), .B(n2493), .Z(n2485) );
  NAND U3270 ( .A(n2430), .B(n2429), .Z(n2434) );
  NAND U3271 ( .A(n2432), .B(n2431), .Z(n2433) );
  NAND U3272 ( .A(n2434), .B(n2433), .Z(n2486) );
  XNOR U3273 ( .A(n2485), .B(n2486), .Z(n2488) );
  NANDN U3274 ( .A(n2436), .B(n2435), .Z(n2440) );
  NANDN U3275 ( .A(n2438), .B(n2437), .Z(n2439) );
  AND U3276 ( .A(n2440), .B(n2439), .Z(n2487) );
  XOR U3277 ( .A(n2488), .B(n2487), .Z(n2474) );
  NANDN U3278 ( .A(n2442), .B(n2441), .Z(n2446) );
  NANDN U3279 ( .A(n2444), .B(n2443), .Z(n2445) );
  AND U3280 ( .A(n2446), .B(n2445), .Z(n2473) );
  XNOR U3281 ( .A(n2474), .B(n2473), .Z(n2475) );
  XOR U3282 ( .A(n2476), .B(n2475), .Z(n2614) );
  NANDN U3283 ( .A(n2448), .B(n2447), .Z(n2452) );
  NAND U3284 ( .A(n2450), .B(n2449), .Z(n2451) );
  NAND U3285 ( .A(n2452), .B(n2451), .Z(n2613) );
  XOR U3286 ( .A(n2614), .B(n2613), .Z(n2616) );
  NANDN U3287 ( .A(n2454), .B(n2453), .Z(n2458) );
  NANDN U3288 ( .A(n2456), .B(n2455), .Z(n2457) );
  AND U3289 ( .A(n2458), .B(n2457), .Z(n2615) );
  XNOR U3290 ( .A(n2616), .B(n2615), .Z(n2621) );
  NANDN U3291 ( .A(n2459), .B(n2460), .Z(n2465) );
  NOR U3292 ( .A(n2461), .B(n2460), .Z(n2463) );
  OR U3293 ( .A(n2463), .B(n2462), .Z(n2464) );
  AND U3294 ( .A(n2465), .B(n2464), .Z(n2620) );
  NANDN U3295 ( .A(n2467), .B(n2466), .Z(n2471) );
  NANDN U3296 ( .A(n2469), .B(n2468), .Z(n2470) );
  AND U3297 ( .A(n2471), .B(n2470), .Z(n2619) );
  XOR U3298 ( .A(n2620), .B(n2619), .Z(n2472) );
  XNOR U3299 ( .A(n2621), .B(n2472), .Z(N58) );
  NANDN U3300 ( .A(n2474), .B(n2473), .Z(n2478) );
  NANDN U3301 ( .A(n2476), .B(n2475), .Z(n2477) );
  AND U3302 ( .A(n2478), .B(n2477), .Z(n2771) );
  NANDN U3303 ( .A(n2480), .B(n2479), .Z(n2484) );
  NAND U3304 ( .A(n2482), .B(n2481), .Z(n2483) );
  AND U3305 ( .A(n2484), .B(n2483), .Z(n2770) );
  XNOR U3306 ( .A(n2771), .B(n2770), .Z(n2773) );
  NANDN U3307 ( .A(n2486), .B(n2485), .Z(n2490) );
  NAND U3308 ( .A(n2488), .B(n2487), .Z(n2489) );
  AND U3309 ( .A(n2490), .B(n2489), .Z(n2623) );
  NANDN U3310 ( .A(n2492), .B(n2491), .Z(n2496) );
  NANDN U3311 ( .A(n2494), .B(n2493), .Z(n2495) );
  NAND U3312 ( .A(n2496), .B(n2495), .Z(n2624) );
  XNOR U3313 ( .A(n2623), .B(n2624), .Z(n2626) );
  NANDN U3314 ( .A(n2498), .B(n2497), .Z(n2502) );
  NAND U3315 ( .A(n2500), .B(n2499), .Z(n2501) );
  AND U3316 ( .A(n2502), .B(n2501), .Z(n2632) );
  AND U3317 ( .A(y[664]), .B(x[130]), .Z(n2653) );
  XOR U3318 ( .A(n2654), .B(n2653), .Z(n2656) );
  NAND U3319 ( .A(y[642]), .B(x[152]), .Z(n2655) );
  XNOR U3320 ( .A(n2656), .B(n2655), .Z(n2690) );
  NAND U3321 ( .A(n2504), .B(n2503), .Z(n2508) );
  NANDN U3322 ( .A(n2506), .B(n2505), .Z(n2507) );
  AND U3323 ( .A(n2508), .B(n2507), .Z(n2689) );
  XOR U3324 ( .A(n2690), .B(n2689), .Z(n2692) );
  NANDN U3325 ( .A(n2510), .B(n2509), .Z(n2514) );
  NANDN U3326 ( .A(n2512), .B(n2511), .Z(n2513) );
  AND U3327 ( .A(n2514), .B(n2513), .Z(n2691) );
  XOR U3328 ( .A(n2692), .B(n2691), .Z(n2727) );
  NAND U3329 ( .A(n2516), .B(n2515), .Z(n2520) );
  NANDN U3330 ( .A(n2518), .B(n2517), .Z(n2519) );
  AND U3331 ( .A(n2520), .B(n2519), .Z(n2726) );
  NANDN U3332 ( .A(n2522), .B(n2521), .Z(n2526) );
  NAND U3333 ( .A(n2524), .B(n2523), .Z(n2525) );
  NAND U3334 ( .A(n2526), .B(n2525), .Z(n2729) );
  NAND U3335 ( .A(n2528), .B(n2527), .Z(n2532) );
  NAND U3336 ( .A(n2530), .B(n2529), .Z(n2531) );
  AND U3337 ( .A(n2532), .B(n2531), .Z(n2721) );
  NANDN U3338 ( .A(n2534), .B(n2533), .Z(n2538) );
  NAND U3339 ( .A(n2536), .B(n2535), .Z(n2537) );
  AND U3340 ( .A(n2538), .B(n2537), .Z(n2720) );
  XNOR U3341 ( .A(n2721), .B(n2720), .Z(n2722) );
  XOR U3342 ( .A(n2723), .B(n2722), .Z(n2630) );
  NANDN U3343 ( .A(n2540), .B(n2539), .Z(n2544) );
  NANDN U3344 ( .A(n2542), .B(n2541), .Z(n2543) );
  AND U3345 ( .A(n2544), .B(n2543), .Z(n2638) );
  AND U3346 ( .A(x[140]), .B(y[654]), .Z(n2841) );
  AND U3347 ( .A(y[661]), .B(x[133]), .Z(n2703) );
  XOR U3348 ( .A(n2841), .B(n2703), .Z(n2705) );
  NAND U3349 ( .A(x[138]), .B(y[656]), .Z(n2704) );
  XNOR U3350 ( .A(n2705), .B(n2704), .Z(n2735) );
  AND U3351 ( .A(x[135]), .B(y[659]), .Z(n2732) );
  AND U3352 ( .A(y[660]), .B(x[134]), .Z(n2546) );
  NAND U3353 ( .A(y[658]), .B(x[136]), .Z(n2545) );
  XNOR U3354 ( .A(n2546), .B(n2545), .Z(n2751) );
  NAND U3355 ( .A(y[657]), .B(x[137]), .Z(n2752) );
  XOR U3356 ( .A(n2751), .B(n2752), .Z(n2733) );
  XOR U3357 ( .A(n2735), .B(n2734), .Z(n2679) );
  NAND U3358 ( .A(n2548), .B(n2547), .Z(n2552) );
  NAND U3359 ( .A(n2550), .B(n2549), .Z(n2551) );
  NAND U3360 ( .A(n2552), .B(n2551), .Z(n2678) );
  NAND U3361 ( .A(n2554), .B(n2553), .Z(n2558) );
  NAND U3362 ( .A(n2556), .B(n2555), .Z(n2557) );
  NAND U3363 ( .A(n2558), .B(n2557), .Z(n2677) );
  XNOR U3364 ( .A(n2678), .B(n2677), .Z(n2680) );
  XNOR U3365 ( .A(n2679), .B(n2680), .Z(n2715) );
  NANDN U3366 ( .A(n2560), .B(n2559), .Z(n2564) );
  NAND U3367 ( .A(n2562), .B(n2561), .Z(n2563) );
  AND U3368 ( .A(n2564), .B(n2563), .Z(n2714) );
  XNOR U3369 ( .A(n2715), .B(n2714), .Z(n2717) );
  NAND U3370 ( .A(n2566), .B(n2565), .Z(n2570) );
  NANDN U3371 ( .A(n2568), .B(n2567), .Z(n2569) );
  AND U3372 ( .A(n2570), .B(n2569), .Z(n2642) );
  NAND U3373 ( .A(n2572), .B(n2571), .Z(n2576) );
  NANDN U3374 ( .A(n2574), .B(n2573), .Z(n2575) );
  AND U3375 ( .A(n2576), .B(n2575), .Z(n2641) );
  XOR U3376 ( .A(n2642), .B(n2641), .Z(n2644) );
  ANDN U3377 ( .B(o[25]), .A(n2577), .Z(n2744) );
  NAND U3378 ( .A(y[652]), .B(x[142]), .Z(n2745) );
  XNOR U3379 ( .A(n2744), .B(n2745), .Z(n2746) );
  NAND U3380 ( .A(y[665]), .B(x[129]), .Z(n2747) );
  XNOR U3381 ( .A(n2746), .B(n2747), .Z(n2696) );
  NAND U3382 ( .A(y[641]), .B(x[153]), .Z(n2755) );
  XNOR U3383 ( .A(o[26]), .B(n2755), .Z(n2708) );
  NAND U3384 ( .A(x[154]), .B(y[640]), .Z(n2709) );
  XNOR U3385 ( .A(n2708), .B(n2709), .Z(n2711) );
  AND U3386 ( .A(y[666]), .B(x[128]), .Z(n2710) );
  XOR U3387 ( .A(n2711), .B(n2710), .Z(n2695) );
  XOR U3388 ( .A(n2696), .B(n2695), .Z(n2698) );
  NAND U3389 ( .A(n2579), .B(n2578), .Z(n2583) );
  NAND U3390 ( .A(n2581), .B(n2580), .Z(n2582) );
  AND U3391 ( .A(n2583), .B(n2582), .Z(n2697) );
  XOR U3392 ( .A(n2698), .B(n2697), .Z(n2643) );
  XOR U3393 ( .A(n2644), .B(n2643), .Z(n2686) );
  AND U3394 ( .A(y[645]), .B(x[149]), .Z(n2738) );
  NANDN U3395 ( .A(n2584), .B(n2738), .Z(n2588) );
  NAND U3396 ( .A(n2586), .B(n2585), .Z(n2587) );
  NAND U3397 ( .A(n2588), .B(n2587), .Z(n2673) );
  XOR U3398 ( .A(n2739), .B(n2738), .Z(n2741) );
  NAND U3399 ( .A(y[646]), .B(x[148]), .Z(n2740) );
  XNOR U3400 ( .A(n2741), .B(n2740), .Z(n2672) );
  NAND U3401 ( .A(x[151]), .B(y[643]), .Z(n2660) );
  XNOR U3402 ( .A(n2659), .B(n2660), .Z(n2662) );
  AND U3403 ( .A(y[644]), .B(x[150]), .Z(n2661) );
  XOR U3404 ( .A(n2662), .B(n2661), .Z(n2671) );
  XOR U3405 ( .A(n2672), .B(n2671), .Z(n2674) );
  XOR U3406 ( .A(n2673), .B(n2674), .Z(n2684) );
  AND U3407 ( .A(x[147]), .B(y[647]), .Z(n2756) );
  NAND U3408 ( .A(x[131]), .B(y[663]), .Z(n2757) );
  XNOR U3409 ( .A(n2756), .B(n2757), .Z(n2758) );
  NAND U3410 ( .A(x[139]), .B(y[655]), .Z(n2759) );
  XNOR U3411 ( .A(n2758), .B(n2759), .Z(n2648) );
  NAND U3412 ( .A(x[132]), .B(y[662]), .Z(n2666) );
  XNOR U3413 ( .A(n2665), .B(n2666), .Z(n2668) );
  XOR U3414 ( .A(n2668), .B(n2667), .Z(n2647) );
  XOR U3415 ( .A(n2648), .B(n2647), .Z(n2650) );
  NAND U3416 ( .A(n2590), .B(n2589), .Z(n2594) );
  NANDN U3417 ( .A(n2592), .B(n2591), .Z(n2593) );
  AND U3418 ( .A(n2594), .B(n2593), .Z(n2649) );
  XNOR U3419 ( .A(n2650), .B(n2649), .Z(n2683) );
  XNOR U3420 ( .A(n2684), .B(n2683), .Z(n2685) );
  XNOR U3421 ( .A(n2686), .B(n2685), .Z(n2716) );
  XOR U3422 ( .A(n2717), .B(n2716), .Z(n2636) );
  NANDN U3423 ( .A(n2596), .B(n2595), .Z(n2600) );
  NANDN U3424 ( .A(n2598), .B(n2597), .Z(n2599) );
  AND U3425 ( .A(n2600), .B(n2599), .Z(n2767) );
  NAND U3426 ( .A(n2602), .B(n2601), .Z(n2606) );
  NANDN U3427 ( .A(n2604), .B(n2603), .Z(n2605) );
  AND U3428 ( .A(n2606), .B(n2605), .Z(n2765) );
  NAND U3429 ( .A(n2608), .B(n2607), .Z(n2612) );
  NANDN U3430 ( .A(n2610), .B(n2609), .Z(n2611) );
  NAND U3431 ( .A(n2612), .B(n2611), .Z(n2764) );
  XNOR U3432 ( .A(n2636), .B(n2635), .Z(n2637) );
  XNOR U3433 ( .A(n2638), .B(n2637), .Z(n2629) );
  XNOR U3434 ( .A(n2630), .B(n2629), .Z(n2631) );
  XNOR U3435 ( .A(n2632), .B(n2631), .Z(n2625) );
  XOR U3436 ( .A(n2626), .B(n2625), .Z(n2772) );
  XOR U3437 ( .A(n2773), .B(n2772), .Z(n2778) );
  NAND U3438 ( .A(n2614), .B(n2613), .Z(n2618) );
  NAND U3439 ( .A(n2616), .B(n2615), .Z(n2617) );
  NAND U3440 ( .A(n2618), .B(n2617), .Z(n2776) );
  XOR U3441 ( .A(n2776), .B(n2777), .Z(n2622) );
  XNOR U3442 ( .A(n2778), .B(n2622), .Z(N59) );
  NANDN U3443 ( .A(n2624), .B(n2623), .Z(n2628) );
  NAND U3444 ( .A(n2626), .B(n2625), .Z(n2627) );
  AND U3445 ( .A(n2628), .B(n2627), .Z(n2783) );
  NANDN U3446 ( .A(n2630), .B(n2629), .Z(n2634) );
  NANDN U3447 ( .A(n2632), .B(n2631), .Z(n2633) );
  AND U3448 ( .A(n2634), .B(n2633), .Z(n2781) );
  NANDN U3449 ( .A(n2636), .B(n2635), .Z(n2640) );
  NANDN U3450 ( .A(n2638), .B(n2637), .Z(n2639) );
  NAND U3451 ( .A(n2640), .B(n2639), .Z(n2791) );
  NAND U3452 ( .A(n2642), .B(n2641), .Z(n2646) );
  NAND U3453 ( .A(n2644), .B(n2643), .Z(n2645) );
  NAND U3454 ( .A(n2646), .B(n2645), .Z(n2908) );
  NAND U3455 ( .A(n2648), .B(n2647), .Z(n2652) );
  NAND U3456 ( .A(n2650), .B(n2649), .Z(n2651) );
  NAND U3457 ( .A(n2652), .B(n2651), .Z(n2906) );
  NAND U3458 ( .A(n2654), .B(n2653), .Z(n2658) );
  ANDN U3459 ( .B(n2656), .A(n2655), .Z(n2657) );
  ANDN U3460 ( .B(n2658), .A(n2657), .Z(n2814) );
  NANDN U3461 ( .A(n2660), .B(n2659), .Z(n2664) );
  NAND U3462 ( .A(n2662), .B(n2661), .Z(n2663) );
  NAND U3463 ( .A(n2664), .B(n2663), .Z(n2813) );
  XNOR U3464 ( .A(n2814), .B(n2813), .Z(n2815) );
  NANDN U3465 ( .A(n2666), .B(n2665), .Z(n2670) );
  NAND U3466 ( .A(n2668), .B(n2667), .Z(n2669) );
  AND U3467 ( .A(n2670), .B(n2669), .Z(n2828) );
  AND U3468 ( .A(x[128]), .B(y[667]), .Z(n2887) );
  NAND U3469 ( .A(x[155]), .B(y[640]), .Z(n2888) );
  XNOR U3470 ( .A(n2887), .B(n2888), .Z(n2890) );
  AND U3471 ( .A(y[641]), .B(x[154]), .Z(n2897) );
  XOR U3472 ( .A(o[27]), .B(n2897), .Z(n2889) );
  XOR U3473 ( .A(n2890), .B(n2889), .Z(n2825) );
  AND U3474 ( .A(x[137]), .B(y[658]), .Z(n2891) );
  NAND U3475 ( .A(y[646]), .B(x[149]), .Z(n2892) );
  XNOR U3476 ( .A(n2891), .B(n2892), .Z(n2893) );
  NAND U3477 ( .A(y[649]), .B(x[146]), .Z(n2894) );
  XOR U3478 ( .A(n2893), .B(n2894), .Z(n2826) );
  XNOR U3479 ( .A(n2825), .B(n2826), .Z(n2827) );
  XOR U3480 ( .A(n2828), .B(n2827), .Z(n2816) );
  XNOR U3481 ( .A(n2815), .B(n2816), .Z(n2907) );
  XOR U3482 ( .A(n2906), .B(n2907), .Z(n2909) );
  XOR U3483 ( .A(n2908), .B(n2909), .Z(n2927) );
  NAND U3484 ( .A(n2672), .B(n2671), .Z(n2676) );
  NAND U3485 ( .A(n2674), .B(n2673), .Z(n2675) );
  AND U3486 ( .A(n2676), .B(n2675), .Z(n2925) );
  NAND U3487 ( .A(n2678), .B(n2677), .Z(n2682) );
  NANDN U3488 ( .A(n2680), .B(n2679), .Z(n2681) );
  AND U3489 ( .A(n2682), .B(n2681), .Z(n2924) );
  XOR U3490 ( .A(n2925), .B(n2924), .Z(n2926) );
  NANDN U3491 ( .A(n2684), .B(n2683), .Z(n2688) );
  NANDN U3492 ( .A(n2686), .B(n2685), .Z(n2687) );
  AND U3493 ( .A(n2688), .B(n2687), .Z(n2912) );
  NAND U3494 ( .A(n2690), .B(n2689), .Z(n2694) );
  NAND U3495 ( .A(n2692), .B(n2691), .Z(n2693) );
  NAND U3496 ( .A(n2694), .B(n2693), .Z(n2902) );
  NAND U3497 ( .A(n2696), .B(n2695), .Z(n2700) );
  NAND U3498 ( .A(n2698), .B(n2697), .Z(n2699) );
  NAND U3499 ( .A(n2700), .B(n2699), .Z(n2900) );
  AND U3500 ( .A(x[147]), .B(y[648]), .Z(n2875) );
  NAND U3501 ( .A(y[642]), .B(x[153]), .Z(n2876) );
  XNOR U3502 ( .A(n2875), .B(n2876), .Z(n2877) );
  NAND U3503 ( .A(y[661]), .B(x[134]), .Z(n2878) );
  XNOR U3504 ( .A(n2877), .B(n2878), .Z(n2867) );
  AND U3505 ( .A(x[143]), .B(y[652]), .Z(n2846) );
  AND U3506 ( .A(x[130]), .B(y[665]), .Z(n2847) );
  XOR U3507 ( .A(n2846), .B(n2847), .Z(n2848) );
  AND U3508 ( .A(y[664]), .B(x[131]), .Z(n2849) );
  XOR U3509 ( .A(n2848), .B(n2849), .Z(n2866) );
  XOR U3510 ( .A(n2867), .B(n2866), .Z(n2868) );
  NAND U3511 ( .A(x[144]), .B(y[651]), .Z(n2832) );
  XOR U3512 ( .A(n2832), .B(n2831), .Z(n2834) );
  XOR U3513 ( .A(n2833), .B(n2834), .Z(n2843) );
  AND U3514 ( .A(y[654]), .B(x[141]), .Z(n2702) );
  NAND U3515 ( .A(y[655]), .B(x[140]), .Z(n2701) );
  XNOR U3516 ( .A(n2702), .B(n2701), .Z(n2842) );
  XOR U3517 ( .A(n2843), .B(n2842), .Z(n2869) );
  XNOR U3518 ( .A(n2868), .B(n2869), .Z(n2810) );
  NAND U3519 ( .A(n2841), .B(n2703), .Z(n2707) );
  ANDN U3520 ( .B(n2705), .A(n2704), .Z(n2706) );
  ANDN U3521 ( .B(n2707), .A(n2706), .Z(n2808) );
  NANDN U3522 ( .A(n2709), .B(n2708), .Z(n2713) );
  NAND U3523 ( .A(n2711), .B(n2710), .Z(n2712) );
  NAND U3524 ( .A(n2713), .B(n2712), .Z(n2807) );
  XNOR U3525 ( .A(n2808), .B(n2807), .Z(n2809) );
  XOR U3526 ( .A(n2810), .B(n2809), .Z(n2901) );
  XNOR U3527 ( .A(n2900), .B(n2901), .Z(n2903) );
  XNOR U3528 ( .A(n2912), .B(n2913), .Z(n2915) );
  NANDN U3529 ( .A(n2715), .B(n2714), .Z(n2719) );
  NAND U3530 ( .A(n2717), .B(n2716), .Z(n2718) );
  AND U3531 ( .A(n2719), .B(n2718), .Z(n2914) );
  XOR U3532 ( .A(n2915), .B(n2914), .Z(n2789) );
  XOR U3533 ( .A(n2790), .B(n2789), .Z(n2792) );
  XOR U3534 ( .A(n2791), .B(n2792), .Z(n2797) );
  NANDN U3535 ( .A(n2721), .B(n2720), .Z(n2725) );
  NAND U3536 ( .A(n2723), .B(n2722), .Z(n2724) );
  AND U3537 ( .A(n2725), .B(n2724), .Z(n2796) );
  NANDN U3538 ( .A(n2727), .B(n2726), .Z(n2731) );
  NANDN U3539 ( .A(n2729), .B(n2728), .Z(n2730) );
  NAND U3540 ( .A(n2731), .B(n2730), .Z(n2802) );
  NANDN U3541 ( .A(n2733), .B(n2732), .Z(n2737) );
  NAND U3542 ( .A(n2735), .B(n2734), .Z(n2736) );
  NAND U3543 ( .A(n2737), .B(n2736), .Z(n2920) );
  NAND U3544 ( .A(n2739), .B(n2738), .Z(n2743) );
  ANDN U3545 ( .B(n2741), .A(n2740), .Z(n2742) );
  ANDN U3546 ( .B(n2743), .A(n2742), .Z(n2859) );
  NANDN U3547 ( .A(n2745), .B(n2744), .Z(n2749) );
  NANDN U3548 ( .A(n2747), .B(n2746), .Z(n2748) );
  NAND U3549 ( .A(n2749), .B(n2748), .Z(n2858) );
  XNOR U3550 ( .A(n2859), .B(n2858), .Z(n2861) );
  AND U3551 ( .A(y[660]), .B(x[136]), .Z(n2899) );
  NAND U3552 ( .A(n2899), .B(n2750), .Z(n2754) );
  NANDN U3553 ( .A(n2752), .B(n2751), .Z(n2753) );
  NAND U3554 ( .A(n2754), .B(n2753), .Z(n2822) );
  AND U3555 ( .A(y[653]), .B(x[142]), .Z(n2852) );
  AND U3556 ( .A(x[129]), .B(y[666]), .Z(n2853) );
  XOR U3557 ( .A(n2852), .B(n2853), .Z(n2854) );
  ANDN U3558 ( .B(o[26]), .A(n2755), .Z(n2855) );
  XOR U3559 ( .A(n2854), .B(n2855), .Z(n2819) );
  AND U3560 ( .A(x[145]), .B(y[650]), .Z(n2881) );
  NAND U3561 ( .A(x[132]), .B(y[663]), .Z(n2882) );
  XNOR U3562 ( .A(n2881), .B(n2882), .Z(n2884) );
  AND U3563 ( .A(y[662]), .B(x[133]), .Z(n2883) );
  XOR U3564 ( .A(n2884), .B(n2883), .Z(n2820) );
  XOR U3565 ( .A(n2819), .B(n2820), .Z(n2821) );
  XOR U3566 ( .A(n2822), .B(n2821), .Z(n2860) );
  XOR U3567 ( .A(n2861), .B(n2860), .Z(n2919) );
  NANDN U3568 ( .A(n2757), .B(n2756), .Z(n2761) );
  NANDN U3569 ( .A(n2759), .B(n2758), .Z(n2760) );
  AND U3570 ( .A(n2761), .B(n2760), .Z(n2865) );
  NAND U3571 ( .A(x[152]), .B(y[643]), .Z(n2762) );
  XNOR U3572 ( .A(n2763), .B(n2762), .Z(n2871) );
  NAND U3573 ( .A(x[135]), .B(y[660]), .Z(n2872) );
  XNOR U3574 ( .A(n2871), .B(n2872), .Z(n2863) );
  AND U3575 ( .A(x[136]), .B(y[659]), .Z(n2835) );
  AND U3576 ( .A(x[151]), .B(y[644]), .Z(n2836) );
  XOR U3577 ( .A(n2835), .B(n2836), .Z(n2837) );
  AND U3578 ( .A(x[150]), .B(y[645]), .Z(n2838) );
  XOR U3579 ( .A(n2837), .B(n2838), .Z(n2862) );
  XOR U3580 ( .A(n2863), .B(n2862), .Z(n2864) );
  XNOR U3581 ( .A(n2865), .B(n2864), .Z(n2918) );
  XOR U3582 ( .A(n2919), .B(n2918), .Z(n2921) );
  XNOR U3583 ( .A(n2920), .B(n2921), .Z(n2801) );
  XOR U3584 ( .A(n2802), .B(n2801), .Z(n2804) );
  NANDN U3585 ( .A(n2765), .B(n2764), .Z(n2769) );
  NANDN U3586 ( .A(n2767), .B(n2766), .Z(n2768) );
  AND U3587 ( .A(n2769), .B(n2768), .Z(n2803) );
  XOR U3588 ( .A(n2804), .B(n2803), .Z(n2795) );
  XNOR U3589 ( .A(n2796), .B(n2795), .Z(n2798) );
  XOR U3590 ( .A(n2797), .B(n2798), .Z(n2780) );
  XOR U3591 ( .A(n2781), .B(n2780), .Z(n2782) );
  XOR U3592 ( .A(n2783), .B(n2782), .Z(n2788) );
  NANDN U3593 ( .A(n2771), .B(n2770), .Z(n2775) );
  NAND U3594 ( .A(n2773), .B(n2772), .Z(n2774) );
  NAND U3595 ( .A(n2775), .B(n2774), .Z(n2787) );
  XOR U3596 ( .A(n2787), .B(n2786), .Z(n2779) );
  XNOR U3597 ( .A(n2788), .B(n2779), .Z(N60) );
  NAND U3598 ( .A(n2781), .B(n2780), .Z(n2785) );
  NAND U3599 ( .A(n2783), .B(n2782), .Z(n2784) );
  NAND U3600 ( .A(n2785), .B(n2784), .Z(n3092) );
  IV U3601 ( .A(n3092), .Z(n3090) );
  NANDN U3602 ( .A(n2790), .B(n2789), .Z(n2794) );
  NANDN U3603 ( .A(n2792), .B(n2791), .Z(n2793) );
  AND U3604 ( .A(n2794), .B(n2793), .Z(n3085) );
  NANDN U3605 ( .A(n2796), .B(n2795), .Z(n2800) );
  NAND U3606 ( .A(n2798), .B(n2797), .Z(n2799) );
  AND U3607 ( .A(n2800), .B(n2799), .Z(n3084) );
  XNOR U3608 ( .A(n3085), .B(n3084), .Z(n3087) );
  NAND U3609 ( .A(n2802), .B(n2801), .Z(n2806) );
  NAND U3610 ( .A(n2804), .B(n2803), .Z(n2805) );
  AND U3611 ( .A(n2806), .B(n2805), .Z(n2931) );
  NANDN U3612 ( .A(n2808), .B(n2807), .Z(n2812) );
  NAND U3613 ( .A(n2810), .B(n2809), .Z(n2811) );
  AND U3614 ( .A(n2812), .B(n2811), .Z(n2956) );
  NANDN U3615 ( .A(n2814), .B(n2813), .Z(n2818) );
  NANDN U3616 ( .A(n2816), .B(n2815), .Z(n2817) );
  AND U3617 ( .A(n2818), .B(n2817), .Z(n3059) );
  NAND U3618 ( .A(n2820), .B(n2819), .Z(n2824) );
  NAND U3619 ( .A(n2822), .B(n2821), .Z(n2823) );
  AND U3620 ( .A(n2824), .B(n2823), .Z(n3057) );
  NANDN U3621 ( .A(n2826), .B(n2825), .Z(n2830) );
  NANDN U3622 ( .A(n2828), .B(n2827), .Z(n2829) );
  NAND U3623 ( .A(n2830), .B(n2829), .Z(n3056) );
  XNOR U3624 ( .A(n3057), .B(n3056), .Z(n3058) );
  XNOR U3625 ( .A(n3059), .B(n3058), .Z(n2955) );
  XNOR U3626 ( .A(n2956), .B(n2955), .Z(n2958) );
  AND U3627 ( .A(x[135]), .B(y[661]), .Z(n3007) );
  AND U3628 ( .A(y[656]), .B(x[140]), .Z(n3006) );
  XOR U3629 ( .A(n3007), .B(n3006), .Z(n3009) );
  AND U3630 ( .A(y[657]), .B(x[139]), .Z(n3008) );
  XOR U3631 ( .A(n3009), .B(n3008), .Z(n3025) );
  AND U3632 ( .A(x[155]), .B(y[641]), .Z(n3023) );
  XOR U3633 ( .A(o[28]), .B(n3023), .Z(n3037) );
  AND U3634 ( .A(x[154]), .B(y[642]), .Z(n3036) );
  XOR U3635 ( .A(n3037), .B(n3036), .Z(n3039) );
  AND U3636 ( .A(x[143]), .B(y[653]), .Z(n3038) );
  XNOR U3637 ( .A(n3039), .B(n3038), .Z(n3024) );
  XOR U3638 ( .A(n3026), .B(n3027), .Z(n3063) );
  NAND U3639 ( .A(n2836), .B(n2835), .Z(n2840) );
  NAND U3640 ( .A(n2838), .B(n2837), .Z(n2839) );
  NAND U3641 ( .A(n2840), .B(n2839), .Z(n2990) );
  AND U3642 ( .A(y[651]), .B(x[145]), .Z(n2966) );
  AND U3643 ( .A(x[150]), .B(y[646]), .Z(n2965) );
  XOR U3644 ( .A(n2966), .B(n2965), .Z(n2968) );
  AND U3645 ( .A(x[132]), .B(y[664]), .Z(n2967) );
  XOR U3646 ( .A(n2968), .B(n2967), .Z(n2989) );
  AND U3647 ( .A(x[134]), .B(y[662]), .Z(n3247) );
  AND U3648 ( .A(x[147]), .B(y[649]), .Z(n3012) );
  XOR U3649 ( .A(n3247), .B(n3012), .Z(n3014) );
  XOR U3650 ( .A(n3014), .B(n3013), .Z(n2988) );
  XOR U3651 ( .A(n2989), .B(n2988), .Z(n2991) );
  XOR U3652 ( .A(n2990), .B(n2991), .Z(n3062) );
  XOR U3653 ( .A(n3063), .B(n3062), .Z(n3065) );
  NAND U3654 ( .A(n3031), .B(n2841), .Z(n2845) );
  NANDN U3655 ( .A(n2843), .B(n2842), .Z(n2844) );
  NAND U3656 ( .A(n2845), .B(n2844), .Z(n2984) );
  NAND U3657 ( .A(n2847), .B(n2846), .Z(n2851) );
  NAND U3658 ( .A(n2849), .B(n2848), .Z(n2850) );
  NAND U3659 ( .A(n2851), .B(n2850), .Z(n2983) );
  NAND U3660 ( .A(n2853), .B(n2852), .Z(n2857) );
  NAND U3661 ( .A(n2855), .B(n2854), .Z(n2856) );
  NAND U3662 ( .A(n2857), .B(n2856), .Z(n2982) );
  XOR U3663 ( .A(n2983), .B(n2982), .Z(n2985) );
  XOR U3664 ( .A(n2984), .B(n2985), .Z(n3064) );
  XOR U3665 ( .A(n3065), .B(n3064), .Z(n2957) );
  XNOR U3666 ( .A(n2958), .B(n2957), .Z(n2952) );
  XNOR U3667 ( .A(n3045), .B(n3044), .Z(n3046) );
  XOR U3668 ( .A(n3047), .B(n3046), .Z(n2949) );
  AND U3669 ( .A(x[152]), .B(y[647]), .Z(n3347) );
  NAND U3670 ( .A(n3347), .B(n2870), .Z(n2874) );
  NANDN U3671 ( .A(n2872), .B(n2871), .Z(n2873) );
  NAND U3672 ( .A(n2874), .B(n2873), .Z(n3074) );
  AND U3673 ( .A(x[153]), .B(y[643]), .Z(n3002) );
  XOR U3674 ( .A(n3003), .B(n3002), .Z(n3001) );
  AND U3675 ( .A(x[129]), .B(y[667]), .Z(n3000) );
  XOR U3676 ( .A(n3001), .B(n3000), .Z(n3073) );
  AND U3677 ( .A(x[144]), .B(y[652]), .Z(n2995) );
  AND U3678 ( .A(y[644]), .B(x[152]), .Z(n2994) );
  XOR U3679 ( .A(n2995), .B(n2994), .Z(n2997) );
  AND U3680 ( .A(x[130]), .B(y[666]), .Z(n2996) );
  XOR U3681 ( .A(n2997), .B(n2996), .Z(n3072) );
  XOR U3682 ( .A(n3073), .B(n3072), .Z(n3075) );
  XNOR U3683 ( .A(n3074), .B(n3075), .Z(n3053) );
  NANDN U3684 ( .A(n2876), .B(n2875), .Z(n2880) );
  NANDN U3685 ( .A(n2878), .B(n2877), .Z(n2879) );
  NAND U3686 ( .A(n2880), .B(n2879), .Z(n3080) );
  AND U3687 ( .A(y[665]), .B(x[131]), .Z(n3030) );
  XOR U3688 ( .A(n3031), .B(n3030), .Z(n3033) );
  AND U3689 ( .A(x[151]), .B(y[645]), .Z(n3032) );
  XOR U3690 ( .A(n3033), .B(n3032), .Z(n3079) );
  AND U3691 ( .A(y[663]), .B(x[133]), .Z(n3018) );
  AND U3692 ( .A(x[149]), .B(y[647]), .Z(n3017) );
  XOR U3693 ( .A(n3018), .B(n3017), .Z(n3020) );
  AND U3694 ( .A(x[148]), .B(y[648]), .Z(n3019) );
  XOR U3695 ( .A(n3020), .B(n3019), .Z(n3078) );
  XOR U3696 ( .A(n3079), .B(n3078), .Z(n3081) );
  XNOR U3697 ( .A(n3080), .B(n3081), .Z(n3051) );
  NANDN U3698 ( .A(n2882), .B(n2881), .Z(n2886) );
  NAND U3699 ( .A(n2884), .B(n2883), .Z(n2885) );
  NAND U3700 ( .A(n2886), .B(n2885), .Z(n3067) );
  XOR U3701 ( .A(n3067), .B(n3066), .Z(n3069) );
  NANDN U3702 ( .A(n2892), .B(n2891), .Z(n2896) );
  NANDN U3703 ( .A(n2894), .B(n2893), .Z(n2895) );
  NAND U3704 ( .A(n2896), .B(n2895), .Z(n2961) );
  AND U3705 ( .A(n2897), .B(o[27]), .Z(n2974) );
  AND U3706 ( .A(x[128]), .B(y[668]), .Z(n2972) );
  AND U3707 ( .A(y[640]), .B(x[156]), .Z(n2971) );
  XOR U3708 ( .A(n2972), .B(n2971), .Z(n2973) );
  XOR U3709 ( .A(n2974), .B(n2973), .Z(n2960) );
  NAND U3710 ( .A(y[658]), .B(x[138]), .Z(n2898) );
  XNOR U3711 ( .A(n2899), .B(n2898), .Z(n2979) );
  AND U3712 ( .A(y[659]), .B(x[137]), .Z(n2978) );
  XOR U3713 ( .A(n2979), .B(n2978), .Z(n2959) );
  XOR U3714 ( .A(n2960), .B(n2959), .Z(n2962) );
  XOR U3715 ( .A(n2961), .B(n2962), .Z(n3068) );
  XNOR U3716 ( .A(n3069), .B(n3068), .Z(n3050) );
  XOR U3717 ( .A(n3051), .B(n3050), .Z(n3052) );
  XOR U3718 ( .A(n3053), .B(n3052), .Z(n2950) );
  XOR U3719 ( .A(n2949), .B(n2950), .Z(n2951) );
  XNOR U3720 ( .A(n2952), .B(n2951), .Z(n2945) );
  NAND U3721 ( .A(n2901), .B(n2900), .Z(n2905) );
  NANDN U3722 ( .A(n2903), .B(n2902), .Z(n2904) );
  NAND U3723 ( .A(n2905), .B(n2904), .Z(n2944) );
  NAND U3724 ( .A(n2907), .B(n2906), .Z(n2911) );
  NAND U3725 ( .A(n2909), .B(n2908), .Z(n2910) );
  NAND U3726 ( .A(n2911), .B(n2910), .Z(n2943) );
  XNOR U3727 ( .A(n2944), .B(n2943), .Z(n2946) );
  XNOR U3728 ( .A(n2931), .B(n2932), .Z(n2933) );
  NANDN U3729 ( .A(n2913), .B(n2912), .Z(n2917) );
  NAND U3730 ( .A(n2915), .B(n2914), .Z(n2916) );
  NAND U3731 ( .A(n2917), .B(n2916), .Z(n2939) );
  NAND U3732 ( .A(n2919), .B(n2918), .Z(n2923) );
  NAND U3733 ( .A(n2921), .B(n2920), .Z(n2922) );
  NAND U3734 ( .A(n2923), .B(n2922), .Z(n2937) );
  NAND U3735 ( .A(n2925), .B(n2924), .Z(n2929) );
  NANDN U3736 ( .A(n2927), .B(n2926), .Z(n2928) );
  AND U3737 ( .A(n2929), .B(n2928), .Z(n2938) );
  XNOR U3738 ( .A(n2937), .B(n2938), .Z(n2940) );
  XNOR U3739 ( .A(n2933), .B(n2934), .Z(n3086) );
  XOR U3740 ( .A(n3087), .B(n3086), .Z(n3093) );
  XNOR U3741 ( .A(n3091), .B(n3093), .Z(n2930) );
  XOR U3742 ( .A(n3090), .B(n2930), .Z(N61) );
  NANDN U3743 ( .A(n2932), .B(n2931), .Z(n2936) );
  NANDN U3744 ( .A(n2934), .B(n2933), .Z(n2935) );
  NAND U3745 ( .A(n2936), .B(n2935), .Z(n3103) );
  NAND U3746 ( .A(n2938), .B(n2937), .Z(n2942) );
  NANDN U3747 ( .A(n2940), .B(n2939), .Z(n2941) );
  NAND U3748 ( .A(n2942), .B(n2941), .Z(n3101) );
  NAND U3749 ( .A(n2944), .B(n2943), .Z(n2948) );
  NANDN U3750 ( .A(n2946), .B(n2945), .Z(n2947) );
  NAND U3751 ( .A(n2948), .B(n2947), .Z(n3107) );
  NAND U3752 ( .A(n2950), .B(n2949), .Z(n2954) );
  NAND U3753 ( .A(n2952), .B(n2951), .Z(n2953) );
  AND U3754 ( .A(n2954), .B(n2953), .Z(n3108) );
  XOR U3755 ( .A(n3107), .B(n3108), .Z(n3110) );
  NAND U3756 ( .A(n2960), .B(n2959), .Z(n2964) );
  NAND U3757 ( .A(n2962), .B(n2961), .Z(n2963) );
  AND U3758 ( .A(n2964), .B(n2963), .Z(n3136) );
  NAND U3759 ( .A(n2966), .B(n2965), .Z(n2970) );
  NAND U3760 ( .A(n2968), .B(n2967), .Z(n2969) );
  NAND U3761 ( .A(n2970), .B(n2969), .Z(n3176) );
  NAND U3762 ( .A(n2972), .B(n2971), .Z(n2976) );
  NAND U3763 ( .A(n2974), .B(n2973), .Z(n2975) );
  NAND U3764 ( .A(n2976), .B(n2975), .Z(n3175) );
  XOR U3765 ( .A(n3176), .B(n3175), .Z(n3177) );
  AND U3766 ( .A(y[660]), .B(x[138]), .Z(n3173) );
  NAND U3767 ( .A(n3173), .B(n2977), .Z(n2981) );
  NAND U3768 ( .A(n2979), .B(n2978), .Z(n2980) );
  NAND U3769 ( .A(n2981), .B(n2980), .Z(n3144) );
  AND U3770 ( .A(x[150]), .B(y[647]), .Z(n3225) );
  AND U3771 ( .A(y[657]), .B(x[140]), .Z(n3461) );
  AND U3772 ( .A(x[129]), .B(y[668]), .Z(n3223) );
  XOR U3773 ( .A(n3461), .B(n3223), .Z(n3224) );
  XOR U3774 ( .A(n3225), .B(n3224), .Z(n3143) );
  AND U3775 ( .A(x[143]), .B(y[654]), .Z(n3228) );
  XOR U3776 ( .A(n3228), .B(n3469), .Z(n3230) );
  XOR U3777 ( .A(n3230), .B(n3229), .Z(n3142) );
  XOR U3778 ( .A(n3143), .B(n3142), .Z(n3145) );
  XNOR U3779 ( .A(n3144), .B(n3145), .Z(n3178) );
  NAND U3780 ( .A(n2983), .B(n2982), .Z(n2987) );
  NAND U3781 ( .A(n2985), .B(n2984), .Z(n2986) );
  AND U3782 ( .A(n2987), .B(n2986), .Z(n3138) );
  XOR U3783 ( .A(n3139), .B(n3138), .Z(n3133) );
  NAND U3784 ( .A(n2989), .B(n2988), .Z(n2993) );
  NAND U3785 ( .A(n2991), .B(n2990), .Z(n2992) );
  NAND U3786 ( .A(n2993), .B(n2992), .Z(n3131) );
  NAND U3787 ( .A(n2995), .B(n2994), .Z(n2999) );
  NAND U3788 ( .A(n2997), .B(n2996), .Z(n2998) );
  NAND U3789 ( .A(n2999), .B(n2998), .Z(n3149) );
  AND U3790 ( .A(n3001), .B(n3000), .Z(n3005) );
  NAND U3791 ( .A(n3003), .B(n3002), .Z(n3004) );
  NANDN U3792 ( .A(n3005), .B(n3004), .Z(n3148) );
  XOR U3793 ( .A(n3149), .B(n3148), .Z(n3150) );
  NAND U3794 ( .A(n3007), .B(n3006), .Z(n3011) );
  NAND U3795 ( .A(n3009), .B(n3008), .Z(n3010) );
  NAND U3796 ( .A(n3011), .B(n3010), .Z(n3189) );
  AND U3797 ( .A(x[139]), .B(y[658]), .Z(n3244) );
  AND U3798 ( .A(x[131]), .B(y[666]), .Z(n3242) );
  AND U3799 ( .A(x[145]), .B(y[652]), .Z(n3241) );
  XOR U3800 ( .A(n3242), .B(n3241), .Z(n3243) );
  XOR U3801 ( .A(n3244), .B(n3243), .Z(n3188) );
  AND U3802 ( .A(x[151]), .B(y[646]), .Z(n3238) );
  AND U3803 ( .A(y[656]), .B(x[141]), .Z(n3236) );
  AND U3804 ( .A(y[645]), .B(x[152]), .Z(n3455) );
  XOR U3805 ( .A(n3236), .B(n3455), .Z(n3237) );
  XOR U3806 ( .A(n3238), .B(n3237), .Z(n3187) );
  XOR U3807 ( .A(n3188), .B(n3187), .Z(n3190) );
  XNOR U3808 ( .A(n3189), .B(n3190), .Z(n3151) );
  NAND U3809 ( .A(n3247), .B(n3012), .Z(n3016) );
  NAND U3810 ( .A(n3014), .B(n3013), .Z(n3015) );
  NAND U3811 ( .A(n3016), .B(n3015), .Z(n3157) );
  AND U3812 ( .A(y[641]), .B(x[156]), .Z(n3235) );
  XOR U3813 ( .A(o[29]), .B(n3235), .Z(n3168) );
  AND U3814 ( .A(x[128]), .B(y[669]), .Z(n3166) );
  AND U3815 ( .A(y[640]), .B(x[157]), .Z(n3165) );
  XOR U3816 ( .A(n3166), .B(n3165), .Z(n3167) );
  XOR U3817 ( .A(n3168), .B(n3167), .Z(n3155) );
  AND U3818 ( .A(y[644]), .B(x[153]), .Z(n3220) );
  AND U3819 ( .A(x[154]), .B(y[643]), .Z(n3217) );
  XOR U3820 ( .A(n3218), .B(n3217), .Z(n3219) );
  XOR U3821 ( .A(n3220), .B(n3219), .Z(n3154) );
  XOR U3822 ( .A(n3155), .B(n3154), .Z(n3156) );
  XOR U3823 ( .A(n3157), .B(n3156), .Z(n3267) );
  NAND U3824 ( .A(n3018), .B(n3017), .Z(n3022) );
  NAND U3825 ( .A(n3020), .B(n3019), .Z(n3021) );
  NAND U3826 ( .A(n3022), .B(n3021), .Z(n3256) );
  AND U3827 ( .A(x[130]), .B(y[667]), .Z(n3206) );
  XOR U3828 ( .A(n3206), .B(n3205), .Z(n3207) );
  XOR U3829 ( .A(n3208), .B(n3207), .Z(n3255) );
  AND U3830 ( .A(n3023), .B(o[28]), .Z(n3196) );
  AND U3831 ( .A(x[144]), .B(y[653]), .Z(n3194) );
  AND U3832 ( .A(x[155]), .B(y[642]), .Z(n3193) );
  XOR U3833 ( .A(n3194), .B(n3193), .Z(n3195) );
  XOR U3834 ( .A(n3196), .B(n3195), .Z(n3254) );
  XOR U3835 ( .A(n3255), .B(n3254), .Z(n3257) );
  XNOR U3836 ( .A(n3256), .B(n3257), .Z(n3266) );
  NANDN U3837 ( .A(n3025), .B(n3024), .Z(n3029) );
  NANDN U3838 ( .A(n3027), .B(n3026), .Z(n3028) );
  NAND U3839 ( .A(n3029), .B(n3028), .Z(n3182) );
  NAND U3840 ( .A(n3031), .B(n3030), .Z(n3035) );
  NAND U3841 ( .A(n3033), .B(n3032), .Z(n3034) );
  NAND U3842 ( .A(n3035), .B(n3034), .Z(n3212) );
  NAND U3843 ( .A(n3037), .B(n3036), .Z(n3041) );
  NAND U3844 ( .A(n3039), .B(n3038), .Z(n3040) );
  NAND U3845 ( .A(n3041), .B(n3040), .Z(n3211) );
  XOR U3846 ( .A(n3212), .B(n3211), .Z(n3214) );
  AND U3847 ( .A(y[661]), .B(x[136]), .Z(n3249) );
  AND U3848 ( .A(y[663]), .B(x[134]), .Z(n3043) );
  AND U3849 ( .A(y[662]), .B(x[135]), .Z(n3042) );
  XOR U3850 ( .A(n3043), .B(n3042), .Z(n3248) );
  XOR U3851 ( .A(n3249), .B(n3248), .Z(n3160) );
  AND U3852 ( .A(x[137]), .B(y[660]), .Z(n3322) );
  XOR U3853 ( .A(n3160), .B(n3322), .Z(n3162) );
  AND U3854 ( .A(y[664]), .B(x[133]), .Z(n3202) );
  AND U3855 ( .A(x[132]), .B(y[665]), .Z(n3200) );
  AND U3856 ( .A(x[138]), .B(y[659]), .Z(n3199) );
  XOR U3857 ( .A(n3200), .B(n3199), .Z(n3201) );
  XOR U3858 ( .A(n3202), .B(n3201), .Z(n3161) );
  XOR U3859 ( .A(n3162), .B(n3161), .Z(n3213) );
  XNOR U3860 ( .A(n3214), .B(n3213), .Z(n3181) );
  XOR U3861 ( .A(n3182), .B(n3181), .Z(n3183) );
  XNOR U3862 ( .A(n3184), .B(n3183), .Z(n3130) );
  XOR U3863 ( .A(n3131), .B(n3130), .Z(n3132) );
  XNOR U3864 ( .A(n3124), .B(n3123), .Z(n3126) );
  NANDN U3865 ( .A(n3045), .B(n3044), .Z(n3049) );
  NANDN U3866 ( .A(n3047), .B(n3046), .Z(n3048) );
  AND U3867 ( .A(n3049), .B(n3048), .Z(n3120) );
  NAND U3868 ( .A(n3051), .B(n3050), .Z(n3055) );
  NAND U3869 ( .A(n3053), .B(n3052), .Z(n3054) );
  AND U3870 ( .A(n3055), .B(n3054), .Z(n3119) );
  XNOR U3871 ( .A(n3120), .B(n3119), .Z(n3122) );
  NANDN U3872 ( .A(n3057), .B(n3056), .Z(n3061) );
  NANDN U3873 ( .A(n3059), .B(n3058), .Z(n3060) );
  NAND U3874 ( .A(n3061), .B(n3060), .Z(n3116) );
  NAND U3875 ( .A(n3067), .B(n3066), .Z(n3071) );
  NAND U3876 ( .A(n3069), .B(n3068), .Z(n3070) );
  NAND U3877 ( .A(n3071), .B(n3070), .Z(n3262) );
  NAND U3878 ( .A(n3073), .B(n3072), .Z(n3077) );
  NAND U3879 ( .A(n3075), .B(n3074), .Z(n3076) );
  NAND U3880 ( .A(n3077), .B(n3076), .Z(n3261) );
  NAND U3881 ( .A(n3079), .B(n3078), .Z(n3083) );
  NAND U3882 ( .A(n3081), .B(n3080), .Z(n3082) );
  NAND U3883 ( .A(n3083), .B(n3082), .Z(n3260) );
  XOR U3884 ( .A(n3261), .B(n3260), .Z(n3263) );
  XOR U3885 ( .A(n3262), .B(n3263), .Z(n3113) );
  XOR U3886 ( .A(n3114), .B(n3113), .Z(n3115) );
  XOR U3887 ( .A(n3116), .B(n3115), .Z(n3121) );
  XOR U3888 ( .A(n3122), .B(n3121), .Z(n3125) );
  XOR U3889 ( .A(n3126), .B(n3125), .Z(n3109) );
  XOR U3890 ( .A(n3110), .B(n3109), .Z(n3102) );
  XNOR U3891 ( .A(n3101), .B(n3102), .Z(n3104) );
  XOR U3892 ( .A(n3103), .B(n3104), .Z(n3100) );
  NANDN U3893 ( .A(n3085), .B(n3084), .Z(n3089) );
  NAND U3894 ( .A(n3087), .B(n3086), .Z(n3088) );
  NAND U3895 ( .A(n3089), .B(n3088), .Z(n3099) );
  NANDN U3896 ( .A(n3090), .B(n3091), .Z(n3096) );
  NOR U3897 ( .A(n3092), .B(n3091), .Z(n3094) );
  OR U3898 ( .A(n3094), .B(n3093), .Z(n3095) );
  AND U3899 ( .A(n3096), .B(n3095), .Z(n3098) );
  XOR U3900 ( .A(n3099), .B(n3098), .Z(n3097) );
  XNOR U3901 ( .A(n3100), .B(n3097), .Z(N62) );
  NAND U3902 ( .A(n3102), .B(n3101), .Z(n3106) );
  NANDN U3903 ( .A(n3104), .B(n3103), .Z(n3105) );
  NAND U3904 ( .A(n3106), .B(n3105), .Z(n3533) );
  NAND U3905 ( .A(n3108), .B(n3107), .Z(n3112) );
  NAND U3906 ( .A(n3110), .B(n3109), .Z(n3111) );
  NAND U3907 ( .A(n3112), .B(n3111), .Z(n3551) );
  NAND U3908 ( .A(n3114), .B(n3113), .Z(n3118) );
  NAND U3909 ( .A(n3116), .B(n3115), .Z(n3117) );
  AND U3910 ( .A(n3118), .B(n3117), .Z(n3272) );
  NANDN U3911 ( .A(n3124), .B(n3123), .Z(n3129) );
  IV U3912 ( .A(n3125), .Z(n3127) );
  NANDN U3913 ( .A(n3127), .B(n3126), .Z(n3128) );
  NAND U3914 ( .A(n3129), .B(n3128), .Z(n3275) );
  XNOR U3915 ( .A(n3274), .B(n3275), .Z(n3273) );
  XNOR U3916 ( .A(n3272), .B(n3273), .Z(n3549) );
  NAND U3917 ( .A(n3131), .B(n3130), .Z(n3135) );
  NANDN U3918 ( .A(n3133), .B(n3132), .Z(n3134) );
  AND U3919 ( .A(n3135), .B(n3134), .Z(n3538) );
  NANDN U3920 ( .A(n3137), .B(n3136), .Z(n3141) );
  NAND U3921 ( .A(n3139), .B(n3138), .Z(n3140) );
  AND U3922 ( .A(n3141), .B(n3140), .Z(n3279) );
  NAND U3923 ( .A(n3143), .B(n3142), .Z(n3147) );
  NAND U3924 ( .A(n3145), .B(n3144), .Z(n3146) );
  AND U3925 ( .A(n3147), .B(n3146), .Z(n3287) );
  NAND U3926 ( .A(n3149), .B(n3148), .Z(n3153) );
  NANDN U3927 ( .A(n3151), .B(n3150), .Z(n3152) );
  AND U3928 ( .A(n3153), .B(n3152), .Z(n3286) );
  XOR U3929 ( .A(n3287), .B(n3286), .Z(n3285) );
  NAND U3930 ( .A(n3155), .B(n3154), .Z(n3159) );
  NAND U3931 ( .A(n3157), .B(n3156), .Z(n3158) );
  AND U3932 ( .A(n3159), .B(n3158), .Z(n3284) );
  XOR U3933 ( .A(n3285), .B(n3284), .Z(n3281) );
  NAND U3934 ( .A(n3160), .B(n3322), .Z(n3164) );
  NAND U3935 ( .A(n3162), .B(n3161), .Z(n3163) );
  AND U3936 ( .A(n3164), .B(n3163), .Z(n3498) );
  NAND U3937 ( .A(n3166), .B(n3165), .Z(n3170) );
  NAND U3938 ( .A(n3168), .B(n3167), .Z(n3169) );
  NAND U3939 ( .A(n3170), .B(n3169), .Z(n3442) );
  AND U3940 ( .A(y[658]), .B(x[140]), .Z(n3172) );
  XOR U3941 ( .A(n3172), .B(n3171), .Z(n3458) );
  XOR U3942 ( .A(n3459), .B(n3458), .Z(n3321) );
  AND U3943 ( .A(y[661]), .B(x[137]), .Z(n3174) );
  XOR U3944 ( .A(n3174), .B(n3173), .Z(n3320) );
  XOR U3945 ( .A(n3321), .B(n3320), .Z(n3445) );
  AND U3946 ( .A(x[155]), .B(y[643]), .Z(n3401) );
  AND U3947 ( .A(x[129]), .B(y[669]), .Z(n3400) );
  XOR U3948 ( .A(n3401), .B(n3400), .Z(n3398) );
  XOR U3949 ( .A(n3399), .B(n3398), .Z(n3444) );
  XOR U3950 ( .A(n3445), .B(n3444), .Z(n3443) );
  XOR U3951 ( .A(n3442), .B(n3443), .Z(n3499) );
  NAND U3952 ( .A(n3176), .B(n3175), .Z(n3180) );
  NANDN U3953 ( .A(n3178), .B(n3177), .Z(n3179) );
  AND U3954 ( .A(n3180), .B(n3179), .Z(n3496) );
  XNOR U3955 ( .A(n3497), .B(n3496), .Z(n3280) );
  XOR U3956 ( .A(n3279), .B(n3278), .Z(n3539) );
  NAND U3957 ( .A(n3182), .B(n3181), .Z(n3186) );
  NAND U3958 ( .A(n3184), .B(n3183), .Z(n3185) );
  AND U3959 ( .A(n3186), .B(n3185), .Z(n3519) );
  NAND U3960 ( .A(n3188), .B(n3187), .Z(n3192) );
  NAND U3961 ( .A(n3190), .B(n3189), .Z(n3191) );
  AND U3962 ( .A(n3192), .B(n3191), .Z(n3509) );
  NAND U3963 ( .A(n3194), .B(n3193), .Z(n3198) );
  NAND U3964 ( .A(n3196), .B(n3195), .Z(n3197) );
  AND U3965 ( .A(n3198), .B(n3197), .Z(n3291) );
  NAND U3966 ( .A(n3200), .B(n3199), .Z(n3204) );
  NAND U3967 ( .A(n3202), .B(n3201), .Z(n3203) );
  AND U3968 ( .A(n3204), .B(n3203), .Z(n3293) );
  AND U3969 ( .A(y[664]), .B(x[134]), .Z(n3411) );
  AND U3970 ( .A(y[665]), .B(x[133]), .Z(n3413) );
  AND U3971 ( .A(y[651]), .B(x[147]), .Z(n3412) );
  XOR U3972 ( .A(n3413), .B(n3412), .Z(n3410) );
  XNOR U3973 ( .A(n3411), .B(n3410), .Z(n3294) );
  AND U3974 ( .A(x[132]), .B(y[666]), .Z(n3473) );
  AND U3975 ( .A(x[131]), .B(y[667]), .Z(n3475) );
  AND U3976 ( .A(x[146]), .B(y[652]), .Z(n3474) );
  XOR U3977 ( .A(n3475), .B(n3474), .Z(n3472) );
  XOR U3978 ( .A(n3473), .B(n3472), .Z(n3297) );
  NAND U3979 ( .A(n3206), .B(n3205), .Z(n3210) );
  NAND U3980 ( .A(n3208), .B(n3207), .Z(n3209) );
  AND U3981 ( .A(n3210), .B(n3209), .Z(n3296) );
  XOR U3982 ( .A(n3294), .B(n3295), .Z(n3292) );
  XOR U3983 ( .A(n3291), .B(n3290), .Z(n3508) );
  XOR U3984 ( .A(n3509), .B(n3508), .Z(n3507) );
  NAND U3985 ( .A(n3212), .B(n3211), .Z(n3216) );
  NAND U3986 ( .A(n3214), .B(n3213), .Z(n3215) );
  AND U3987 ( .A(n3216), .B(n3215), .Z(n3506) );
  XOR U3988 ( .A(n3507), .B(n3506), .Z(n3521) );
  NAND U3989 ( .A(n3218), .B(n3217), .Z(n3222) );
  AND U3990 ( .A(n3220), .B(n3219), .Z(n3221) );
  ANDN U3991 ( .B(n3222), .A(n3221), .Z(n3315) );
  NAND U3992 ( .A(n3461), .B(n3223), .Z(n3227) );
  AND U3993 ( .A(n3225), .B(n3224), .Z(n3226) );
  ANDN U3994 ( .B(n3227), .A(n3226), .Z(n3317) );
  NAND U3995 ( .A(n3228), .B(n3469), .Z(n3232) );
  NAND U3996 ( .A(n3230), .B(n3229), .Z(n3231) );
  AND U3997 ( .A(n3232), .B(n3231), .Z(n3307) );
  AND U3998 ( .A(x[151]), .B(y[647]), .Z(n3453) );
  AND U3999 ( .A(x[152]), .B(y[646]), .Z(n3234) );
  NAND U4000 ( .A(x[153]), .B(y[645]), .Z(n3233) );
  XNOR U4001 ( .A(n3234), .B(n3233), .Z(n3452) );
  XOR U4002 ( .A(n3453), .B(n3452), .Z(n3309) );
  AND U4003 ( .A(n3235), .B(o[29]), .Z(n3332) );
  AND U4004 ( .A(y[642]), .B(x[156]), .Z(n3334) );
  AND U4005 ( .A(x[144]), .B(y[654]), .Z(n3333) );
  XOR U4006 ( .A(n3334), .B(n3333), .Z(n3331) );
  XNOR U4007 ( .A(n3332), .B(n3331), .Z(n3308) );
  XNOR U4008 ( .A(n3307), .B(n3306), .Z(n3316) );
  XNOR U4009 ( .A(n3315), .B(n3314), .Z(n3503) );
  NAND U4010 ( .A(n3236), .B(n3455), .Z(n3240) );
  NAND U4011 ( .A(n3238), .B(n3237), .Z(n3239) );
  AND U4012 ( .A(n3240), .B(n3239), .Z(n3493) );
  NAND U4013 ( .A(n3242), .B(n3241), .Z(n3246) );
  NAND U4014 ( .A(n3244), .B(n3243), .Z(n3245) );
  AND U4015 ( .A(n3246), .B(n3245), .Z(n3301) );
  AND U4016 ( .A(x[128]), .B(y[670]), .Z(n3340) );
  AND U4017 ( .A(y[641]), .B(x[157]), .Z(n3345) );
  XOR U4018 ( .A(o[30]), .B(n3345), .Z(n3342) );
  AND U4019 ( .A(y[640]), .B(x[158]), .Z(n3341) );
  XOR U4020 ( .A(n3342), .B(n3341), .Z(n3339) );
  XOR U4021 ( .A(n3340), .B(n3339), .Z(n3303) );
  AND U4022 ( .A(y[650]), .B(x[148]), .Z(n3406) );
  XOR U4023 ( .A(n3407), .B(n3406), .Z(n3405) );
  AND U4024 ( .A(x[136]), .B(y[662]), .Z(n3404) );
  XNOR U4025 ( .A(n3405), .B(n3404), .Z(n3302) );
  XNOR U4026 ( .A(n3301), .B(n3300), .Z(n3492) );
  AND U4027 ( .A(x[135]), .B(y[663]), .Z(n3467) );
  NAND U4028 ( .A(n3247), .B(n3467), .Z(n3251) );
  NAND U4029 ( .A(n3249), .B(n3248), .Z(n3250) );
  AND U4030 ( .A(n3251), .B(n3250), .Z(n3437) );
  AND U4031 ( .A(x[149]), .B(y[649]), .Z(n3253) );
  NAND U4032 ( .A(y[648]), .B(x[150]), .Z(n3252) );
  XNOR U4033 ( .A(n3253), .B(n3252), .Z(n3466) );
  XOR U4034 ( .A(n3467), .B(n3466), .Z(n3439) );
  AND U4035 ( .A(y[653]), .B(x[145]), .Z(n3326) );
  AND U4036 ( .A(x[130]), .B(y[668]), .Z(n3327) );
  NAND U4037 ( .A(x[154]), .B(y[644]), .Z(n3328) );
  XNOR U4038 ( .A(n3326), .B(n3325), .Z(n3438) );
  XOR U4039 ( .A(n3437), .B(n3436), .Z(n3491) );
  XNOR U4040 ( .A(n3490), .B(n3491), .Z(n3504) );
  NAND U4041 ( .A(n3255), .B(n3254), .Z(n3259) );
  NAND U4042 ( .A(n3257), .B(n3256), .Z(n3258) );
  AND U4043 ( .A(n3259), .B(n3258), .Z(n3505) );
  XOR U4044 ( .A(n3503), .B(n3502), .Z(n3520) );
  XOR U4045 ( .A(n3519), .B(n3518), .Z(n3515) );
  NAND U4046 ( .A(n3261), .B(n3260), .Z(n3265) );
  NAND U4047 ( .A(n3263), .B(n3262), .Z(n3264) );
  AND U4048 ( .A(n3265), .B(n3264), .Z(n3514) );
  NANDN U4049 ( .A(n3267), .B(n3266), .Z(n3271) );
  NANDN U4050 ( .A(n3269), .B(n3268), .Z(n3270) );
  NAND U4051 ( .A(n3271), .B(n3270), .Z(n3512) );
  XOR U4052 ( .A(n3513), .B(n3512), .Z(n3536) );
  XOR U4053 ( .A(n3537), .B(n3536), .Z(n3548) );
  XOR U4054 ( .A(n3551), .B(n3550), .Z(n3530) );
  XNOR U4055 ( .A(n3531), .B(n3530), .Z(N63) );
  NAND U4056 ( .A(n3273), .B(n3272), .Z(n3277) );
  NANDN U4057 ( .A(n3275), .B(n3274), .Z(n3276) );
  AND U4058 ( .A(n3277), .B(n3276), .Z(n3547) );
  NAND U4059 ( .A(n3279), .B(n3278), .Z(n3283) );
  NANDN U4060 ( .A(n3281), .B(n3280), .Z(n3282) );
  AND U4061 ( .A(n3283), .B(n3282), .Z(n3529) );
  NAND U4062 ( .A(n3285), .B(n3284), .Z(n3289) );
  NAND U4063 ( .A(n3287), .B(n3286), .Z(n3288) );
  AND U4064 ( .A(n3289), .B(n3288), .Z(n3511) );
  NANDN U4065 ( .A(n3295), .B(n3294), .Z(n3299) );
  NANDN U4066 ( .A(n3297), .B(n3296), .Z(n3298) );
  NAND U4067 ( .A(n3301), .B(n3300), .Z(n3305) );
  NANDN U4068 ( .A(n3303), .B(n3302), .Z(n3304) );
  AND U4069 ( .A(n3305), .B(n3304), .Z(n3313) );
  NAND U4070 ( .A(n3307), .B(n3306), .Z(n3311) );
  NANDN U4071 ( .A(n3309), .B(n3308), .Z(n3310) );
  NAND U4072 ( .A(n3311), .B(n3310), .Z(n3312) );
  XNOR U4073 ( .A(n3313), .B(n3312), .Z(n3489) );
  NANDN U4074 ( .A(n3315), .B(n3314), .Z(n3319) );
  NANDN U4075 ( .A(n3317), .B(n3316), .Z(n3318) );
  AND U4076 ( .A(n3319), .B(n3318), .Z(n3487) );
  NAND U4077 ( .A(n3321), .B(n3320), .Z(n3324) );
  AND U4078 ( .A(x[138]), .B(y[661]), .Z(n3346) );
  NAND U4079 ( .A(n3322), .B(n3346), .Z(n3323) );
  AND U4080 ( .A(n3324), .B(n3323), .Z(n3397) );
  NAND U4081 ( .A(n3326), .B(n3325), .Z(n3330) );
  NANDN U4082 ( .A(n3328), .B(n3327), .Z(n3329) );
  AND U4083 ( .A(n3330), .B(n3329), .Z(n3338) );
  NAND U4084 ( .A(n3332), .B(n3331), .Z(n3336) );
  NAND U4085 ( .A(n3334), .B(n3333), .Z(n3335) );
  NAND U4086 ( .A(n3336), .B(n3335), .Z(n3337) );
  XNOR U4087 ( .A(n3338), .B(n3337), .Z(n3395) );
  NAND U4088 ( .A(n3340), .B(n3339), .Z(n3344) );
  NAND U4089 ( .A(n3342), .B(n3341), .Z(n3343) );
  AND U4090 ( .A(n3344), .B(n3343), .Z(n3393) );
  AND U4091 ( .A(x[149]), .B(y[650]), .Z(n3353) );
  AND U4092 ( .A(n3345), .B(o[30]), .Z(n3351) );
  XOR U4093 ( .A(n3346), .B(o[31]), .Z(n3349) );
  XNOR U4094 ( .A(n3347), .B(n3460), .Z(n3348) );
  XNOR U4095 ( .A(n3349), .B(n3348), .Z(n3350) );
  XNOR U4096 ( .A(n3351), .B(n3350), .Z(n3352) );
  XNOR U4097 ( .A(n3353), .B(n3352), .Z(n3391) );
  AND U4098 ( .A(y[652]), .B(x[147]), .Z(n3355) );
  NAND U4099 ( .A(y[663]), .B(x[136]), .Z(n3354) );
  XNOR U4100 ( .A(n3355), .B(n3354), .Z(n3363) );
  AND U4101 ( .A(y[659]), .B(x[140]), .Z(n3361) );
  AND U4102 ( .A(x[157]), .B(y[642]), .Z(n3357) );
  NAND U4103 ( .A(y[645]), .B(x[154]), .Z(n3356) );
  XNOR U4104 ( .A(n3357), .B(n3356), .Z(n3358) );
  XNOR U4105 ( .A(n3359), .B(n3358), .Z(n3360) );
  XNOR U4106 ( .A(n3361), .B(n3360), .Z(n3362) );
  XOR U4107 ( .A(n3363), .B(n3362), .Z(n3365) );
  AND U4108 ( .A(y[646]), .B(x[153]), .Z(n3454) );
  AND U4109 ( .A(x[150]), .B(y[649]), .Z(n3468) );
  XNOR U4110 ( .A(n3454), .B(n3468), .Z(n3364) );
  XNOR U4111 ( .A(n3365), .B(n3364), .Z(n3381) );
  AND U4112 ( .A(y[660]), .B(x[139]), .Z(n3367) );
  NAND U4113 ( .A(x[142]), .B(y[657]), .Z(n3366) );
  XNOR U4114 ( .A(n3367), .B(n3366), .Z(n3371) );
  AND U4115 ( .A(y[665]), .B(x[134]), .Z(n3369) );
  NAND U4116 ( .A(y[664]), .B(x[135]), .Z(n3368) );
  XNOR U4117 ( .A(n3369), .B(n3368), .Z(n3370) );
  XOR U4118 ( .A(n3371), .B(n3370), .Z(n3379) );
  AND U4119 ( .A(x[158]), .B(y[641]), .Z(n3373) );
  NAND U4120 ( .A(y[655]), .B(x[144]), .Z(n3372) );
  XNOR U4121 ( .A(n3373), .B(n3372), .Z(n3377) );
  AND U4122 ( .A(x[137]), .B(y[662]), .Z(n3375) );
  NAND U4123 ( .A(x[148]), .B(y[651]), .Z(n3374) );
  XNOR U4124 ( .A(n3375), .B(n3374), .Z(n3376) );
  XNOR U4125 ( .A(n3377), .B(n3376), .Z(n3378) );
  XNOR U4126 ( .A(n3379), .B(n3378), .Z(n3380) );
  XOR U4127 ( .A(n3381), .B(n3380), .Z(n3389) );
  AND U4128 ( .A(y[643]), .B(x[156]), .Z(n3383) );
  NAND U4129 ( .A(y[670]), .B(x[129]), .Z(n3382) );
  XNOR U4130 ( .A(n3383), .B(n3382), .Z(n3387) );
  AND U4131 ( .A(y[671]), .B(x[128]), .Z(n3385) );
  NAND U4132 ( .A(y[654]), .B(x[145]), .Z(n3384) );
  XNOR U4133 ( .A(n3385), .B(n3384), .Z(n3386) );
  XNOR U4134 ( .A(n3387), .B(n3386), .Z(n3388) );
  XNOR U4135 ( .A(n3389), .B(n3388), .Z(n3390) );
  XNOR U4136 ( .A(n3391), .B(n3390), .Z(n3392) );
  XNOR U4137 ( .A(n3393), .B(n3392), .Z(n3394) );
  XNOR U4138 ( .A(n3395), .B(n3394), .Z(n3396) );
  XNOR U4139 ( .A(n3397), .B(n3396), .Z(n3485) );
  NAND U4140 ( .A(n3399), .B(n3398), .Z(n3403) );
  NAND U4141 ( .A(n3401), .B(n3400), .Z(n3402) );
  AND U4142 ( .A(n3403), .B(n3402), .Z(n3435) );
  NAND U4143 ( .A(n3405), .B(n3404), .Z(n3409) );
  NAND U4144 ( .A(n3407), .B(n3406), .Z(n3408) );
  AND U4145 ( .A(n3409), .B(n3408), .Z(n3417) );
  NAND U4146 ( .A(n3411), .B(n3410), .Z(n3415) );
  NAND U4147 ( .A(n3413), .B(n3412), .Z(n3414) );
  NAND U4148 ( .A(n3415), .B(n3414), .Z(n3416) );
  XNOR U4149 ( .A(n3417), .B(n3416), .Z(n3433) );
  AND U4150 ( .A(y[668]), .B(x[131]), .Z(n3419) );
  NAND U4151 ( .A(y[667]), .B(x[132]), .Z(n3418) );
  XNOR U4152 ( .A(n3419), .B(n3418), .Z(n3423) );
  AND U4153 ( .A(x[133]), .B(y[666]), .Z(n3421) );
  NAND U4154 ( .A(x[146]), .B(y[653]), .Z(n3420) );
  XNOR U4155 ( .A(n3421), .B(n3420), .Z(n3422) );
  XOR U4156 ( .A(n3423), .B(n3422), .Z(n3431) );
  AND U4157 ( .A(x[159]), .B(y[640]), .Z(n3425) );
  NAND U4158 ( .A(y[648]), .B(x[151]), .Z(n3424) );
  XNOR U4159 ( .A(n3425), .B(n3424), .Z(n3429) );
  AND U4160 ( .A(y[669]), .B(x[130]), .Z(n3427) );
  NAND U4161 ( .A(y[644]), .B(x[155]), .Z(n3426) );
  XNOR U4162 ( .A(n3427), .B(n3426), .Z(n3428) );
  XNOR U4163 ( .A(n3429), .B(n3428), .Z(n3430) );
  XNOR U4164 ( .A(n3431), .B(n3430), .Z(n3432) );
  XNOR U4165 ( .A(n3433), .B(n3432), .Z(n3434) );
  XNOR U4166 ( .A(n3435), .B(n3434), .Z(n3451) );
  NAND U4167 ( .A(n3437), .B(n3436), .Z(n3441) );
  NANDN U4168 ( .A(n3439), .B(n3438), .Z(n3440) );
  AND U4169 ( .A(n3441), .B(n3440), .Z(n3449) );
  NAND U4170 ( .A(n3443), .B(n3442), .Z(n3447) );
  NAND U4171 ( .A(n3445), .B(n3444), .Z(n3446) );
  NAND U4172 ( .A(n3447), .B(n3446), .Z(n3448) );
  XNOR U4173 ( .A(n3449), .B(n3448), .Z(n3450) );
  XOR U4174 ( .A(n3451), .B(n3450), .Z(n3483) );
  NAND U4175 ( .A(n3453), .B(n3452), .Z(n3457) );
  NAND U4176 ( .A(n3455), .B(n3454), .Z(n3456) );
  AND U4177 ( .A(n3457), .B(n3456), .Z(n3465) );
  NAND U4178 ( .A(n3459), .B(n3458), .Z(n3463) );
  NAND U4179 ( .A(n3461), .B(n3460), .Z(n3462) );
  NAND U4180 ( .A(n3463), .B(n3462), .Z(n3464) );
  XNOR U4181 ( .A(n3465), .B(n3464), .Z(n3481) );
  NAND U4182 ( .A(n3467), .B(n3466), .Z(n3471) );
  NAND U4183 ( .A(n3469), .B(n3468), .Z(n3470) );
  AND U4184 ( .A(n3471), .B(n3470), .Z(n3479) );
  NAND U4185 ( .A(n3473), .B(n3472), .Z(n3477) );
  NAND U4186 ( .A(n3475), .B(n3474), .Z(n3476) );
  NAND U4187 ( .A(n3477), .B(n3476), .Z(n3478) );
  XNOR U4188 ( .A(n3479), .B(n3478), .Z(n3480) );
  XNOR U4189 ( .A(n3481), .B(n3480), .Z(n3482) );
  XNOR U4190 ( .A(n3483), .B(n3482), .Z(n3484) );
  XNOR U4191 ( .A(n3485), .B(n3484), .Z(n3486) );
  XNOR U4192 ( .A(n3487), .B(n3486), .Z(n3488) );
  NANDN U4193 ( .A(n3491), .B(n3490), .Z(n3495) );
  NANDN U4194 ( .A(n3493), .B(n3492), .Z(n3494) );
  NAND U4195 ( .A(n3497), .B(n3496), .Z(n3501) );
  NANDN U4196 ( .A(n3499), .B(n3498), .Z(n3500) );
  XNOR U4197 ( .A(n3511), .B(n3510), .Z(n3527) );
  NAND U4198 ( .A(n3513), .B(n3512), .Z(n3517) );
  NANDN U4199 ( .A(n3515), .B(n3514), .Z(n3516) );
  AND U4200 ( .A(n3517), .B(n3516), .Z(n3525) );
  NAND U4201 ( .A(n3519), .B(n3518), .Z(n3523) );
  NANDN U4202 ( .A(n3521), .B(n3520), .Z(n3522) );
  NAND U4203 ( .A(n3523), .B(n3522), .Z(n3524) );
  XNOR U4204 ( .A(n3525), .B(n3524), .Z(n3526) );
  XNOR U4205 ( .A(n3527), .B(n3526), .Z(n3528) );
  XNOR U4206 ( .A(n3529), .B(n3528), .Z(n3545) );
  NAND U4207 ( .A(n3531), .B(n3530), .Z(n3535) );
  NANDN U4208 ( .A(n3533), .B(n3532), .Z(n3534) );
  AND U4209 ( .A(n3535), .B(n3534), .Z(n3543) );
  NAND U4210 ( .A(n3537), .B(n3536), .Z(n3541) );
  NANDN U4211 ( .A(n3539), .B(n3538), .Z(n3540) );
  NAND U4212 ( .A(n3541), .B(n3540), .Z(n3542) );
  XNOR U4213 ( .A(n3543), .B(n3542), .Z(n3544) );
  XNOR U4214 ( .A(n3545), .B(n3544), .Z(n3546) );
  XNOR U4215 ( .A(n3547), .B(n3546), .Z(n3555) );
  ANDN U4216 ( .B(n3549), .A(n3548), .Z(n3553) );
  ANDN U4217 ( .B(n3551), .A(n3550), .Z(n3552) );
  NOR U4218 ( .A(n3553), .B(n3552), .Z(n3554) );
  XNOR U4219 ( .A(n3555), .B(n3554), .Z(N64) );
  AND U4220 ( .A(x[128]), .B(y[672]), .Z(n4205) );
  XOR U4221 ( .A(n4205), .B(o[32]), .Z(N97) );
  NAND U4222 ( .A(x[129]), .B(y[672]), .Z(n3565) );
  AND U4223 ( .A(x[128]), .B(y[673]), .Z(n3561) );
  XNOR U4224 ( .A(n3561), .B(o[33]), .Z(n3556) );
  XOR U4225 ( .A(n3565), .B(n3556), .Z(n3558) );
  NAND U4226 ( .A(n4205), .B(o[32]), .Z(n3557) );
  XNOR U4227 ( .A(n3558), .B(n3557), .Z(N98) );
  AND U4228 ( .A(x[128]), .B(y[674]), .Z(n3564) );
  XNOR U4229 ( .A(n3564), .B(o[34]), .Z(n3570) );
  XNOR U4230 ( .A(n3571), .B(n3570), .Z(n3573) );
  AND U4231 ( .A(y[673]), .B(x[129]), .Z(n3560) );
  NAND U4232 ( .A(y[672]), .B(x[130]), .Z(n3559) );
  XNOR U4233 ( .A(n3560), .B(n3559), .Z(n3567) );
  AND U4234 ( .A(n3561), .B(o[33]), .Z(n3566) );
  XNOR U4235 ( .A(n3567), .B(n3566), .Z(n3572) );
  XNOR U4236 ( .A(n3573), .B(n3572), .Z(N99) );
  AND U4237 ( .A(x[129]), .B(y[674]), .Z(n3684) );
  AND U4238 ( .A(x[130]), .B(y[673]), .Z(n3583) );
  XOR U4239 ( .A(n3583), .B(o[35]), .Z(n3588) );
  XOR U4240 ( .A(n3684), .B(n3588), .Z(n3590) );
  AND U4241 ( .A(y[675]), .B(x[128]), .Z(n3563) );
  NAND U4242 ( .A(y[672]), .B(x[131]), .Z(n3562) );
  XNOR U4243 ( .A(n3563), .B(n3562), .Z(n3577) );
  NAND U4244 ( .A(n3564), .B(o[34]), .Z(n3578) );
  XNOR U4245 ( .A(n3577), .B(n3578), .Z(n3589) );
  XNOR U4246 ( .A(n3590), .B(n3589), .Z(n3587) );
  NANDN U4247 ( .A(n3565), .B(n3583), .Z(n3569) );
  NAND U4248 ( .A(n3567), .B(n3566), .Z(n3568) );
  NAND U4249 ( .A(n3569), .B(n3568), .Z(n3585) );
  NANDN U4250 ( .A(n3571), .B(n3570), .Z(n3575) );
  NAND U4251 ( .A(n3573), .B(n3572), .Z(n3574) );
  AND U4252 ( .A(n3575), .B(n3574), .Z(n3586) );
  XOR U4253 ( .A(n3585), .B(n3586), .Z(n3576) );
  XNOR U4254 ( .A(n3587), .B(n3576), .Z(N100) );
  AND U4255 ( .A(x[131]), .B(y[675]), .Z(n3641) );
  NAND U4256 ( .A(n4205), .B(n3641), .Z(n3580) );
  NANDN U4257 ( .A(n3578), .B(n3577), .Z(n3579) );
  AND U4258 ( .A(n3580), .B(n3579), .Z(n3610) );
  AND U4259 ( .A(y[676]), .B(x[128]), .Z(n3582) );
  NAND U4260 ( .A(y[672]), .B(x[132]), .Z(n3581) );
  XNOR U4261 ( .A(n3582), .B(n3581), .Z(n3604) );
  AND U4262 ( .A(n3583), .B(o[35]), .Z(n3603) );
  XOR U4263 ( .A(n3604), .B(n3603), .Z(n3608) );
  AND U4264 ( .A(y[675]), .B(x[129]), .Z(n3789) );
  NAND U4265 ( .A(y[674]), .B(x[130]), .Z(n3584) );
  XNOR U4266 ( .A(n3789), .B(n3584), .Z(n3600) );
  AND U4267 ( .A(x[131]), .B(y[673]), .Z(n3595) );
  XOR U4268 ( .A(n3595), .B(o[36]), .Z(n3599) );
  XOR U4269 ( .A(n3600), .B(n3599), .Z(n3607) );
  XOR U4270 ( .A(n3608), .B(n3607), .Z(n3609) );
  XNOR U4271 ( .A(n3610), .B(n3609), .Z(n3614) );
  NAND U4272 ( .A(n3684), .B(n3588), .Z(n3592) );
  NAND U4273 ( .A(n3590), .B(n3589), .Z(n3591) );
  NAND U4274 ( .A(n3592), .B(n3591), .Z(n3611) );
  XNOR U4275 ( .A(n3612), .B(n3611), .Z(n3613) );
  XOR U4276 ( .A(n3614), .B(n3613), .Z(N101) );
  AND U4277 ( .A(y[677]), .B(x[128]), .Z(n3594) );
  NAND U4278 ( .A(y[672]), .B(x[133]), .Z(n3593) );
  XNOR U4279 ( .A(n3594), .B(n3593), .Z(n3634) );
  AND U4280 ( .A(n3595), .B(o[36]), .Z(n3633) );
  XOR U4281 ( .A(n3634), .B(n3633), .Z(n3632) );
  NAND U4282 ( .A(x[130]), .B(y[675]), .Z(n3692) );
  AND U4283 ( .A(y[676]), .B(x[129]), .Z(n3597) );
  NAND U4284 ( .A(y[674]), .B(x[131]), .Z(n3596) );
  XNOR U4285 ( .A(n3597), .B(n3596), .Z(n3628) );
  AND U4286 ( .A(x[132]), .B(y[673]), .Z(n3639) );
  XOR U4287 ( .A(n3639), .B(o[37]), .Z(n3627) );
  XOR U4288 ( .A(n3628), .B(n3627), .Z(n3631) );
  XOR U4289 ( .A(n3692), .B(n3631), .Z(n3598) );
  XNOR U4290 ( .A(n3632), .B(n3598), .Z(n3620) );
  NANDN U4291 ( .A(n3692), .B(n3684), .Z(n3602) );
  NAND U4292 ( .A(n3600), .B(n3599), .Z(n3601) );
  NAND U4293 ( .A(n3602), .B(n3601), .Z(n3619) );
  AND U4294 ( .A(x[132]), .B(y[676]), .Z(n4399) );
  NAND U4295 ( .A(n4399), .B(n4205), .Z(n3606) );
  NAND U4296 ( .A(n3604), .B(n3603), .Z(n3605) );
  NAND U4297 ( .A(n3606), .B(n3605), .Z(n3618) );
  XNOR U4298 ( .A(n3619), .B(n3618), .Z(n3621) );
  NANDN U4299 ( .A(n3612), .B(n3611), .Z(n3616) );
  NAND U4300 ( .A(n3614), .B(n3613), .Z(n3615) );
  AND U4301 ( .A(n3616), .B(n3615), .Z(n3624) );
  XOR U4302 ( .A(n3625), .B(n3624), .Z(n3617) );
  XNOR U4303 ( .A(n3626), .B(n3617), .Z(N102) );
  NAND U4304 ( .A(n3619), .B(n3618), .Z(n3623) );
  NANDN U4305 ( .A(n3621), .B(n3620), .Z(n3622) );
  AND U4306 ( .A(n3623), .B(n3622), .Z(n3674) );
  AND U4307 ( .A(x[131]), .B(y[676]), .Z(n3693) );
  NAND U4308 ( .A(n3693), .B(n3684), .Z(n3630) );
  NAND U4309 ( .A(n3628), .B(n3627), .Z(n3629) );
  AND U4310 ( .A(n3630), .B(n3629), .Z(n3669) );
  XNOR U4311 ( .A(n3669), .B(n3668), .Z(n3671) );
  AND U4312 ( .A(x[133]), .B(y[677]), .Z(n3869) );
  NAND U4313 ( .A(n4205), .B(n3869), .Z(n3636) );
  NAND U4314 ( .A(n3634), .B(n3633), .Z(n3635) );
  NAND U4315 ( .A(n3636), .B(n3635), .Z(n3644) );
  AND U4316 ( .A(y[678]), .B(x[128]), .Z(n3638) );
  NAND U4317 ( .A(y[672]), .B(x[134]), .Z(n3637) );
  XNOR U4318 ( .A(n3638), .B(n3637), .Z(n3651) );
  NAND U4319 ( .A(n3639), .B(o[37]), .Z(n3652) );
  XNOR U4320 ( .A(n3651), .B(n3652), .Z(n3645) );
  XOR U4321 ( .A(n3644), .B(n3645), .Z(n3647) );
  NAND U4322 ( .A(y[676]), .B(x[130]), .Z(n3640) );
  XNOR U4323 ( .A(n3641), .B(n3640), .Z(n3656) );
  AND U4324 ( .A(y[677]), .B(x[129]), .Z(n3908) );
  NAND U4325 ( .A(y[674]), .B(x[132]), .Z(n3642) );
  XNOR U4326 ( .A(n3908), .B(n3642), .Z(n3660) );
  AND U4327 ( .A(x[133]), .B(y[673]), .Z(n3667) );
  XOR U4328 ( .A(n3667), .B(o[38]), .Z(n3659) );
  XOR U4329 ( .A(n3660), .B(n3659), .Z(n3655) );
  XOR U4330 ( .A(n3656), .B(n3655), .Z(n3646) );
  XOR U4331 ( .A(n3647), .B(n3646), .Z(n3670) );
  XOR U4332 ( .A(n3671), .B(n3670), .Z(n3676) );
  XNOR U4333 ( .A(n3675), .B(n3676), .Z(n3643) );
  XOR U4334 ( .A(n3674), .B(n3643), .Z(N103) );
  NAND U4335 ( .A(n3645), .B(n3644), .Z(n3649) );
  NAND U4336 ( .A(n3647), .B(n3646), .Z(n3648) );
  AND U4337 ( .A(n3649), .B(n3648), .Z(n3716) );
  AND U4338 ( .A(y[674]), .B(x[133]), .Z(n3777) );
  NAND U4339 ( .A(y[678]), .B(x[129]), .Z(n3650) );
  XNOR U4340 ( .A(n3777), .B(n3650), .Z(n3686) );
  NAND U4341 ( .A(x[134]), .B(y[673]), .Z(n3690) );
  XNOR U4342 ( .A(o[39]), .B(n3690), .Z(n3685) );
  XOR U4343 ( .A(n3686), .B(n3685), .Z(n3705) );
  AND U4344 ( .A(x[134]), .B(y[678]), .Z(n3754) );
  NAND U4345 ( .A(n4205), .B(n3754), .Z(n3654) );
  NANDN U4346 ( .A(n3652), .B(n3651), .Z(n3653) );
  AND U4347 ( .A(n3654), .B(n3653), .Z(n3704) );
  XNOR U4348 ( .A(n3705), .B(n3704), .Z(n3706) );
  NANDN U4349 ( .A(n3692), .B(n3693), .Z(n3658) );
  NAND U4350 ( .A(n3656), .B(n3655), .Z(n3657) );
  NAND U4351 ( .A(n3658), .B(n3657), .Z(n3707) );
  XNOR U4352 ( .A(n3706), .B(n3707), .Z(n3714) );
  AND U4353 ( .A(x[132]), .B(y[677]), .Z(n4210) );
  NAND U4354 ( .A(n4210), .B(n3684), .Z(n3662) );
  NAND U4355 ( .A(n3660), .B(n3659), .Z(n3661) );
  AND U4356 ( .A(n3662), .B(n3661), .Z(n3681) );
  AND U4357 ( .A(y[677]), .B(x[130]), .Z(n3664) );
  NAND U4358 ( .A(y[675]), .B(x[132]), .Z(n3663) );
  XNOR U4359 ( .A(n3664), .B(n3663), .Z(n3694) );
  XOR U4360 ( .A(n3694), .B(n3693), .Z(n3679) );
  AND U4361 ( .A(y[679]), .B(x[128]), .Z(n3666) );
  NAND U4362 ( .A(y[672]), .B(x[135]), .Z(n3665) );
  XNOR U4363 ( .A(n3666), .B(n3665), .Z(n3699) );
  AND U4364 ( .A(n3667), .B(o[38]), .Z(n3698) );
  XNOR U4365 ( .A(n3699), .B(n3698), .Z(n3678) );
  XNOR U4366 ( .A(n3679), .B(n3678), .Z(n3680) );
  XOR U4367 ( .A(n3681), .B(n3680), .Z(n3713) );
  XOR U4368 ( .A(n3714), .B(n3713), .Z(n3715) );
  XOR U4369 ( .A(n3716), .B(n3715), .Z(n3712) );
  NANDN U4370 ( .A(n3669), .B(n3668), .Z(n3673) );
  NAND U4371 ( .A(n3671), .B(n3670), .Z(n3672) );
  NAND U4372 ( .A(n3673), .B(n3672), .Z(n3711) );
  XOR U4373 ( .A(n3711), .B(n3710), .Z(n3677) );
  XNOR U4374 ( .A(n3712), .B(n3677), .Z(N104) );
  NANDN U4375 ( .A(n3679), .B(n3678), .Z(n3683) );
  NAND U4376 ( .A(n3681), .B(n3680), .Z(n3682) );
  AND U4377 ( .A(n3683), .B(n3682), .Z(n3767) );
  AND U4378 ( .A(x[133]), .B(y[678]), .Z(n3861) );
  NAND U4379 ( .A(n3861), .B(n3684), .Z(n3688) );
  NAND U4380 ( .A(n3686), .B(n3685), .Z(n3687) );
  NAND U4381 ( .A(n3688), .B(n3687), .Z(n3765) );
  AND U4382 ( .A(y[675]), .B(x[133]), .Z(n4310) );
  NAND U4383 ( .A(y[679]), .B(x[129]), .Z(n3689) );
  XNOR U4384 ( .A(n4310), .B(n3689), .Z(n3745) );
  ANDN U4385 ( .B(o[39]), .A(n3690), .Z(n3744) );
  XOR U4386 ( .A(n3745), .B(n3744), .Z(n3750) );
  NAND U4387 ( .A(x[131]), .B(y[677]), .Z(n4534) );
  AND U4388 ( .A(y[678]), .B(x[130]), .Z(n4614) );
  NAND U4389 ( .A(y[674]), .B(x[134]), .Z(n3691) );
  XNOR U4390 ( .A(n4614), .B(n3691), .Z(n3755) );
  XNOR U4391 ( .A(n4399), .B(n3755), .Z(n3748) );
  XOR U4392 ( .A(n4534), .B(n3748), .Z(n3749) );
  XOR U4393 ( .A(n3750), .B(n3749), .Z(n3764) );
  XOR U4394 ( .A(n3765), .B(n3764), .Z(n3766) );
  XOR U4395 ( .A(n3767), .B(n3766), .Z(n3723) );
  NANDN U4396 ( .A(n3692), .B(n4210), .Z(n3696) );
  NAND U4397 ( .A(n3694), .B(n3693), .Z(n3695) );
  NAND U4398 ( .A(n3696), .B(n3695), .Z(n3760) );
  AND U4399 ( .A(x[135]), .B(y[679]), .Z(n3697) );
  NAND U4400 ( .A(n4205), .B(n3697), .Z(n3701) );
  NAND U4401 ( .A(n3699), .B(n3698), .Z(n3700) );
  NAND U4402 ( .A(n3701), .B(n3700), .Z(n3758) );
  AND U4403 ( .A(y[680]), .B(x[128]), .Z(n3703) );
  NAND U4404 ( .A(y[672]), .B(x[136]), .Z(n3702) );
  XNOR U4405 ( .A(n3703), .B(n3702), .Z(n3735) );
  NAND U4406 ( .A(x[135]), .B(y[673]), .Z(n3740) );
  XNOR U4407 ( .A(o[40]), .B(n3740), .Z(n3734) );
  XOR U4408 ( .A(n3735), .B(n3734), .Z(n3759) );
  XNOR U4409 ( .A(n3758), .B(n3759), .Z(n3761) );
  NANDN U4410 ( .A(n3705), .B(n3704), .Z(n3709) );
  NANDN U4411 ( .A(n3707), .B(n3706), .Z(n3708) );
  NAND U4412 ( .A(n3709), .B(n3708), .Z(n3720) );
  XOR U4413 ( .A(n3721), .B(n3720), .Z(n3722) );
  XNOR U4414 ( .A(n3723), .B(n3722), .Z(n3729) );
  NAND U4415 ( .A(n3714), .B(n3713), .Z(n3718) );
  NAND U4416 ( .A(n3716), .B(n3715), .Z(n3717) );
  AND U4417 ( .A(n3718), .B(n3717), .Z(n3727) );
  IV U4418 ( .A(n3727), .Z(n3726) );
  XOR U4419 ( .A(n3728), .B(n3726), .Z(n3719) );
  XNOR U4420 ( .A(n3729), .B(n3719), .Z(N105) );
  NAND U4421 ( .A(n3721), .B(n3720), .Z(n3725) );
  NANDN U4422 ( .A(n3723), .B(n3722), .Z(n3724) );
  NAND U4423 ( .A(n3725), .B(n3724), .Z(n3815) );
  IV U4424 ( .A(n3815), .Z(n3813) );
  OR U4425 ( .A(n3728), .B(n3726), .Z(n3732) );
  ANDN U4426 ( .B(n3728), .A(n3727), .Z(n3730) );
  OR U4427 ( .A(n3730), .B(n3729), .Z(n3731) );
  AND U4428 ( .A(n3732), .B(n3731), .Z(n3814) );
  AND U4429 ( .A(x[136]), .B(y[680]), .Z(n3733) );
  NAND U4430 ( .A(n3733), .B(n4205), .Z(n3737) );
  NAND U4431 ( .A(n3735), .B(n3734), .Z(n3736) );
  AND U4432 ( .A(n3737), .B(n3736), .Z(n3806) );
  AND U4433 ( .A(y[676]), .B(x[133]), .Z(n3739) );
  NAND U4434 ( .A(y[674]), .B(x[135]), .Z(n3738) );
  XNOR U4435 ( .A(n3739), .B(n3738), .Z(n3780) );
  ANDN U4436 ( .B(o[40]), .A(n3740), .Z(n3779) );
  XOR U4437 ( .A(n3780), .B(n3779), .Z(n3804) );
  AND U4438 ( .A(y[672]), .B(x[137]), .Z(n3742) );
  NAND U4439 ( .A(y[681]), .B(x[128]), .Z(n3741) );
  XNOR U4440 ( .A(n3742), .B(n3741), .Z(n3786) );
  NAND U4441 ( .A(x[136]), .B(y[673]), .Z(n3795) );
  XNOR U4442 ( .A(o[41]), .B(n3795), .Z(n3785) );
  XNOR U4443 ( .A(n3786), .B(n3785), .Z(n3803) );
  XOR U4444 ( .A(n3806), .B(n3805), .Z(n3800) );
  AND U4445 ( .A(y[680]), .B(x[129]), .Z(n4521) );
  NAND U4446 ( .A(y[675]), .B(x[134]), .Z(n3743) );
  XNOR U4447 ( .A(n4521), .B(n3743), .Z(n3790) );
  XOR U4448 ( .A(n4210), .B(n3790), .Z(n3810) );
  AND U4449 ( .A(x[130]), .B(y[679]), .Z(n4439) );
  NAND U4450 ( .A(x[131]), .B(y[678]), .Z(n4159) );
  XNOR U4451 ( .A(n4439), .B(n4159), .Z(n3809) );
  NAND U4452 ( .A(x[133]), .B(y[679]), .Z(n3981) );
  NANDN U4453 ( .A(n3981), .B(n3789), .Z(n3747) );
  NAND U4454 ( .A(n3745), .B(n3744), .Z(n3746) );
  NAND U4455 ( .A(n3747), .B(n3746), .Z(n3797) );
  XOR U4456 ( .A(n3798), .B(n3797), .Z(n3799) );
  XOR U4457 ( .A(n3800), .B(n3799), .Z(n3773) );
  NAND U4458 ( .A(n4534), .B(n3748), .Z(n3752) );
  NANDN U4459 ( .A(n3750), .B(n3749), .Z(n3751) );
  AND U4460 ( .A(n3752), .B(n3751), .Z(n3772) );
  AND U4461 ( .A(x[130]), .B(y[674]), .Z(n3753) );
  NAND U4462 ( .A(n3754), .B(n3753), .Z(n3757) );
  NAND U4463 ( .A(n4399), .B(n3755), .Z(n3756) );
  AND U4464 ( .A(n3757), .B(n3756), .Z(n3771) );
  XNOR U4465 ( .A(n3772), .B(n3771), .Z(n3774) );
  XOR U4466 ( .A(n3773), .B(n3774), .Z(n3823) );
  NAND U4467 ( .A(n3759), .B(n3758), .Z(n3763) );
  NANDN U4468 ( .A(n3761), .B(n3760), .Z(n3762) );
  NAND U4469 ( .A(n3763), .B(n3762), .Z(n3821) );
  NAND U4470 ( .A(n3765), .B(n3764), .Z(n3769) );
  NAND U4471 ( .A(n3767), .B(n3766), .Z(n3768) );
  NAND U4472 ( .A(n3769), .B(n3768), .Z(n3820) );
  XOR U4473 ( .A(n3821), .B(n3820), .Z(n3822) );
  XNOR U4474 ( .A(n3814), .B(n3816), .Z(n3770) );
  XOR U4475 ( .A(n3813), .B(n3770), .Z(N106) );
  NANDN U4476 ( .A(n3772), .B(n3771), .Z(n3776) );
  NAND U4477 ( .A(n3774), .B(n3773), .Z(n3775) );
  AND U4478 ( .A(n3776), .B(n3775), .Z(n3885) );
  AND U4479 ( .A(x[135]), .B(y[676]), .Z(n3778) );
  NAND U4480 ( .A(n3778), .B(n3777), .Z(n3782) );
  NAND U4481 ( .A(n3780), .B(n3779), .Z(n3781) );
  AND U4482 ( .A(n3782), .B(n3781), .Z(n3876) );
  AND U4483 ( .A(y[678]), .B(x[132]), .Z(n3784) );
  NAND U4484 ( .A(y[675]), .B(x[135]), .Z(n3783) );
  XNOR U4485 ( .A(n3784), .B(n3783), .Z(n3847) );
  NAND U4486 ( .A(x[134]), .B(y[676]), .Z(n3848) );
  XNOR U4487 ( .A(n3847), .B(n3848), .Z(n3874) );
  AND U4488 ( .A(x[136]), .B(y[674]), .Z(n4068) );
  NAND U4489 ( .A(x[137]), .B(y[673]), .Z(n3857) );
  XNOR U4490 ( .A(o[42]), .B(n3857), .Z(n3868) );
  XOR U4491 ( .A(n4068), .B(n3868), .Z(n3870) );
  XNOR U4492 ( .A(n3870), .B(n3869), .Z(n3873) );
  XOR U4493 ( .A(n3876), .B(n3875), .Z(n3836) );
  AND U4494 ( .A(x[137]), .B(y[681]), .Z(n4408) );
  NAND U4495 ( .A(n4408), .B(n4205), .Z(n3788) );
  NAND U4496 ( .A(n3786), .B(n3785), .Z(n3787) );
  AND U4497 ( .A(n3788), .B(n3787), .Z(n3834) );
  AND U4498 ( .A(x[134]), .B(y[680]), .Z(n4103) );
  NAND U4499 ( .A(n4103), .B(n3789), .Z(n3792) );
  NAND U4500 ( .A(n4210), .B(n3790), .Z(n3791) );
  AND U4501 ( .A(n3792), .B(n3791), .Z(n3842) );
  AND U4502 ( .A(y[682]), .B(x[128]), .Z(n3794) );
  NAND U4503 ( .A(y[672]), .B(x[138]), .Z(n3793) );
  XNOR U4504 ( .A(n3794), .B(n3793), .Z(n3852) );
  ANDN U4505 ( .B(o[41]), .A(n3795), .Z(n3851) );
  XOR U4506 ( .A(n3852), .B(n3851), .Z(n3840) );
  AND U4507 ( .A(y[681]), .B(x[129]), .Z(n4717) );
  NAND U4508 ( .A(y[679]), .B(x[131]), .Z(n3796) );
  XNOR U4509 ( .A(n4717), .B(n3796), .Z(n3864) );
  NAND U4510 ( .A(x[130]), .B(y[680]), .Z(n3865) );
  XNOR U4511 ( .A(n3864), .B(n3865), .Z(n3839) );
  XOR U4512 ( .A(n3840), .B(n3839), .Z(n3841) );
  XNOR U4513 ( .A(n3842), .B(n3841), .Z(n3833) );
  NAND U4514 ( .A(n3798), .B(n3797), .Z(n3802) );
  NANDN U4515 ( .A(n3800), .B(n3799), .Z(n3801) );
  AND U4516 ( .A(n3802), .B(n3801), .Z(n3830) );
  NANDN U4517 ( .A(n3804), .B(n3803), .Z(n3808) );
  NAND U4518 ( .A(n3806), .B(n3805), .Z(n3807) );
  AND U4519 ( .A(n3808), .B(n3807), .Z(n3827) );
  ANDN U4520 ( .B(n4159), .A(n4439), .Z(n3812) );
  NANDN U4521 ( .A(n3810), .B(n3809), .Z(n3811) );
  NANDN U4522 ( .A(n3812), .B(n3811), .Z(n3828) );
  XOR U4523 ( .A(n3830), .B(n3829), .Z(n3882) );
  XOR U4524 ( .A(n3883), .B(n3882), .Z(n3884) );
  XOR U4525 ( .A(n3885), .B(n3884), .Z(n3881) );
  NANDN U4526 ( .A(n3813), .B(n3814), .Z(n3819) );
  NOR U4527 ( .A(n3815), .B(n3814), .Z(n3817) );
  OR U4528 ( .A(n3817), .B(n3816), .Z(n3818) );
  AND U4529 ( .A(n3819), .B(n3818), .Z(n3880) );
  NAND U4530 ( .A(n3821), .B(n3820), .Z(n3825) );
  NANDN U4531 ( .A(n3823), .B(n3822), .Z(n3824) );
  AND U4532 ( .A(n3825), .B(n3824), .Z(n3879) );
  XOR U4533 ( .A(n3880), .B(n3879), .Z(n3826) );
  XNOR U4534 ( .A(n3881), .B(n3826), .Z(N107) );
  NANDN U4535 ( .A(n3828), .B(n3827), .Z(n3832) );
  NANDN U4536 ( .A(n3830), .B(n3829), .Z(n3831) );
  AND U4537 ( .A(n3832), .B(n3831), .Z(n3892) );
  NANDN U4538 ( .A(n3834), .B(n3833), .Z(n3838) );
  NANDN U4539 ( .A(n3836), .B(n3835), .Z(n3837) );
  AND U4540 ( .A(n3838), .B(n3837), .Z(n3890) );
  NAND U4541 ( .A(n3840), .B(n3839), .Z(n3844) );
  NANDN U4542 ( .A(n3842), .B(n3841), .Z(n3843) );
  NAND U4543 ( .A(n3844), .B(n3843), .Z(n3949) );
  AND U4544 ( .A(x[135]), .B(y[678]), .Z(n3846) );
  AND U4545 ( .A(x[132]), .B(y[675]), .Z(n3845) );
  NAND U4546 ( .A(n3846), .B(n3845), .Z(n3850) );
  NANDN U4547 ( .A(n3848), .B(n3847), .Z(n3849) );
  AND U4548 ( .A(n3850), .B(n3849), .Z(n3947) );
  AND U4549 ( .A(x[138]), .B(y[682]), .Z(n4620) );
  NAND U4550 ( .A(n4620), .B(n4205), .Z(n3854) );
  NAND U4551 ( .A(n3852), .B(n3851), .Z(n3853) );
  AND U4552 ( .A(n3854), .B(n3853), .Z(n3943) );
  AND U4553 ( .A(y[683]), .B(x[128]), .Z(n3856) );
  NAND U4554 ( .A(y[672]), .B(x[139]), .Z(n3855) );
  XNOR U4555 ( .A(n3856), .B(n3855), .Z(n3920) );
  ANDN U4556 ( .B(o[42]), .A(n3857), .Z(n3919) );
  XOR U4557 ( .A(n3920), .B(n3919), .Z(n3941) );
  AND U4558 ( .A(y[682]), .B(x[129]), .Z(n3859) );
  NAND U4559 ( .A(y[677]), .B(x[134]), .Z(n3858) );
  XNOR U4560 ( .A(n3859), .B(n3858), .Z(n3910) );
  NAND U4561 ( .A(x[138]), .B(y[673]), .Z(n3928) );
  XOR U4562 ( .A(n3910), .B(n3909), .Z(n3940) );
  XOR U4563 ( .A(n3941), .B(n3940), .Z(n3942) );
  XNOR U4564 ( .A(n3943), .B(n3942), .Z(n3946) );
  XNOR U4565 ( .A(n3947), .B(n3946), .Z(n3948) );
  XNOR U4566 ( .A(n3949), .B(n3948), .Z(n3931) );
  AND U4567 ( .A(x[131]), .B(y[680]), .Z(n4874) );
  NAND U4568 ( .A(y[681]), .B(x[130]), .Z(n3860) );
  XNOR U4569 ( .A(n3861), .B(n3860), .Z(n3905) );
  AND U4570 ( .A(x[132]), .B(y[679]), .Z(n3904) );
  XNOR U4571 ( .A(n3905), .B(n3904), .Z(n3935) );
  XNOR U4572 ( .A(n4874), .B(n3935), .Z(n3937) );
  AND U4573 ( .A(y[674]), .B(x[137]), .Z(n3863) );
  NAND U4574 ( .A(y[676]), .B(x[135]), .Z(n3862) );
  XNOR U4575 ( .A(n3863), .B(n3862), .Z(n3924) );
  AND U4576 ( .A(x[136]), .B(y[675]), .Z(n3923) );
  XNOR U4577 ( .A(n3924), .B(n3923), .Z(n3936) );
  XOR U4578 ( .A(n3937), .B(n3936), .Z(n3901) );
  NAND U4579 ( .A(x[131]), .B(y[681]), .Z(n3972) );
  AND U4580 ( .A(x[129]), .B(y[679]), .Z(n4200) );
  NANDN U4581 ( .A(n3972), .B(n4200), .Z(n3867) );
  NANDN U4582 ( .A(n3865), .B(n3864), .Z(n3866) );
  AND U4583 ( .A(n3867), .B(n3866), .Z(n3899) );
  NAND U4584 ( .A(n4068), .B(n3868), .Z(n3872) );
  NAND U4585 ( .A(n3870), .B(n3869), .Z(n3871) );
  NAND U4586 ( .A(n3872), .B(n3871), .Z(n3898) );
  XNOR U4587 ( .A(n3899), .B(n3898), .Z(n3900) );
  XNOR U4588 ( .A(n3901), .B(n3900), .Z(n3930) );
  NANDN U4589 ( .A(n3874), .B(n3873), .Z(n3878) );
  NAND U4590 ( .A(n3876), .B(n3875), .Z(n3877) );
  NAND U4591 ( .A(n3878), .B(n3877), .Z(n3929) );
  XOR U4592 ( .A(n3931), .B(n3932), .Z(n3889) );
  XOR U4593 ( .A(n3892), .B(n3891), .Z(n3897) );
  NAND U4594 ( .A(n3883), .B(n3882), .Z(n3887) );
  NANDN U4595 ( .A(n3885), .B(n3884), .Z(n3886) );
  AND U4596 ( .A(n3887), .B(n3886), .Z(n3896) );
  XOR U4597 ( .A(n3895), .B(n3896), .Z(n3888) );
  XNOR U4598 ( .A(n3897), .B(n3888), .Z(N108) );
  NANDN U4599 ( .A(n3890), .B(n3889), .Z(n3894) );
  NANDN U4600 ( .A(n3892), .B(n3891), .Z(n3893) );
  NAND U4601 ( .A(n3894), .B(n3893), .Z(n4018) );
  IV U4602 ( .A(n4018), .Z(n4017) );
  NANDN U4603 ( .A(n3899), .B(n3898), .Z(n3903) );
  NANDN U4604 ( .A(n3901), .B(n3900), .Z(n3902) );
  AND U4605 ( .A(n3903), .B(n3902), .Z(n4014) );
  AND U4606 ( .A(x[133]), .B(y[681]), .Z(n4430) );
  NAND U4607 ( .A(n4614), .B(n4430), .Z(n3907) );
  NAND U4608 ( .A(n3905), .B(n3904), .Z(n3906) );
  NAND U4609 ( .A(n3907), .B(n3906), .Z(n3960) );
  AND U4610 ( .A(x[134]), .B(y[682]), .Z(n4217) );
  NAND U4611 ( .A(n4217), .B(n3908), .Z(n3912) );
  NAND U4612 ( .A(n3910), .B(n3909), .Z(n3911) );
  NAND U4613 ( .A(n3912), .B(n3911), .Z(n3959) );
  XOR U4614 ( .A(n3960), .B(n3959), .Z(n3961) );
  AND U4615 ( .A(x[137]), .B(y[675]), .Z(n4609) );
  AND U4616 ( .A(y[680]), .B(x[132]), .Z(n3914) );
  NAND U4617 ( .A(y[674]), .B(x[138]), .Z(n3913) );
  XOR U4618 ( .A(n3914), .B(n3913), .Z(n4004) );
  NAND U4619 ( .A(x[135]), .B(y[677]), .Z(n3980) );
  XOR U4620 ( .A(n3981), .B(n3980), .Z(n3983) );
  AND U4621 ( .A(y[684]), .B(x[128]), .Z(n3916) );
  NAND U4622 ( .A(y[672]), .B(x[140]), .Z(n3915) );
  XNOR U4623 ( .A(n3916), .B(n3915), .Z(n3997) );
  NAND U4624 ( .A(x[139]), .B(y[673]), .Z(n3977) );
  XNOR U4625 ( .A(o[44]), .B(n3977), .Z(n3996) );
  XOR U4626 ( .A(n3997), .B(n3996), .Z(n3966) );
  AND U4627 ( .A(y[682]), .B(x[130]), .Z(n3918) );
  NAND U4628 ( .A(y[676]), .B(x[136]), .Z(n3917) );
  XNOR U4629 ( .A(n3918), .B(n3917), .Z(n3971) );
  XOR U4630 ( .A(n3966), .B(n3965), .Z(n3967) );
  XNOR U4631 ( .A(n3961), .B(n3962), .Z(n4012) );
  AND U4632 ( .A(x[139]), .B(y[683]), .Z(n5020) );
  NAND U4633 ( .A(n5020), .B(n4205), .Z(n3922) );
  NAND U4634 ( .A(n3920), .B(n3919), .Z(n3921) );
  AND U4635 ( .A(n3922), .B(n3921), .Z(n3989) );
  AND U4636 ( .A(x[135]), .B(y[674]), .Z(n4135) );
  AND U4637 ( .A(x[137]), .B(y[676]), .Z(n3979) );
  NAND U4638 ( .A(n4135), .B(n3979), .Z(n3926) );
  NAND U4639 ( .A(n3924), .B(n3923), .Z(n3925) );
  AND U4640 ( .A(n3926), .B(n3925), .Z(n3987) );
  AND U4641 ( .A(y[683]), .B(x[129]), .Z(n4644) );
  NAND U4642 ( .A(y[678]), .B(x[134]), .Z(n3927) );
  XNOR U4643 ( .A(n4644), .B(n3927), .Z(n3993) );
  ANDN U4644 ( .B(o[43]), .A(n3928), .Z(n3992) );
  XOR U4645 ( .A(n3993), .B(n3992), .Z(n3986) );
  XNOR U4646 ( .A(n3987), .B(n3986), .Z(n3988) );
  XNOR U4647 ( .A(n3989), .B(n3988), .Z(n4011) );
  XOR U4648 ( .A(n4012), .B(n4011), .Z(n4013) );
  XNOR U4649 ( .A(n4014), .B(n4013), .Z(n4025) );
  NANDN U4650 ( .A(n3930), .B(n3929), .Z(n3934) );
  NANDN U4651 ( .A(n3932), .B(n3931), .Z(n3933) );
  NAND U4652 ( .A(n3934), .B(n3933), .Z(n4024) );
  NANDN U4653 ( .A(n4874), .B(n3935), .Z(n3939) );
  NAND U4654 ( .A(n3937), .B(n3936), .Z(n3938) );
  AND U4655 ( .A(n3939), .B(n3938), .Z(n3954) );
  NAND U4656 ( .A(n3941), .B(n3940), .Z(n3945) );
  NANDN U4657 ( .A(n3943), .B(n3942), .Z(n3944) );
  AND U4658 ( .A(n3945), .B(n3944), .Z(n3953) );
  XNOR U4659 ( .A(n3954), .B(n3953), .Z(n3956) );
  NANDN U4660 ( .A(n3947), .B(n3946), .Z(n3951) );
  NAND U4661 ( .A(n3949), .B(n3948), .Z(n3950) );
  AND U4662 ( .A(n3951), .B(n3950), .Z(n3955) );
  XOR U4663 ( .A(n3956), .B(n3955), .Z(n4026) );
  XOR U4664 ( .A(n4027), .B(n4026), .Z(n4020) );
  XNOR U4665 ( .A(n4019), .B(n4020), .Z(n3952) );
  XOR U4666 ( .A(n4017), .B(n3952), .Z(N109) );
  NANDN U4667 ( .A(n3954), .B(n3953), .Z(n3958) );
  NAND U4668 ( .A(n3956), .B(n3955), .Z(n3957) );
  AND U4669 ( .A(n3958), .B(n3957), .Z(n4034) );
  NAND U4670 ( .A(n3960), .B(n3959), .Z(n3964) );
  NANDN U4671 ( .A(n3962), .B(n3961), .Z(n3963) );
  NAND U4672 ( .A(n3964), .B(n3963), .Z(n4044) );
  NAND U4673 ( .A(n3966), .B(n3965), .Z(n3970) );
  NANDN U4674 ( .A(n3968), .B(n3967), .Z(n3969) );
  NAND U4675 ( .A(n3970), .B(n3969), .Z(n4052) );
  AND U4676 ( .A(x[136]), .B(y[682]), .Z(n5268) );
  AND U4677 ( .A(x[130]), .B(y[676]), .Z(n4144) );
  NAND U4678 ( .A(n5268), .B(n4144), .Z(n3974) );
  NANDN U4679 ( .A(n3972), .B(n3971), .Z(n3973) );
  AND U4680 ( .A(n3974), .B(n3973), .Z(n4084) );
  AND U4681 ( .A(y[684]), .B(x[129]), .Z(n3976) );
  NAND U4682 ( .A(y[678]), .B(x[135]), .Z(n3975) );
  XNOR U4683 ( .A(n3976), .B(n3975), .Z(n4075) );
  ANDN U4684 ( .B(o[44]), .A(n3977), .Z(n4074) );
  XOR U4685 ( .A(n4075), .B(n4074), .Z(n4082) );
  AND U4686 ( .A(x[134]), .B(y[679]), .Z(n5058) );
  NAND U4687 ( .A(y[683]), .B(x[130]), .Z(n3978) );
  XOR U4688 ( .A(n3979), .B(n3978), .Z(n4087) );
  XNOR U4689 ( .A(n5058), .B(n4087), .Z(n4081) );
  XOR U4690 ( .A(n4082), .B(n4081), .Z(n4083) );
  NAND U4691 ( .A(n3981), .B(n3980), .Z(n3985) );
  ANDN U4692 ( .B(n3983), .A(n3982), .Z(n3984) );
  ANDN U4693 ( .B(n3985), .A(n3984), .Z(n4050) );
  XOR U4694 ( .A(n4051), .B(n4050), .Z(n4053) );
  XOR U4695 ( .A(n4052), .B(n4053), .Z(n4045) );
  XOR U4696 ( .A(n4044), .B(n4045), .Z(n4047) );
  NANDN U4697 ( .A(n3987), .B(n3986), .Z(n3991) );
  NANDN U4698 ( .A(n3989), .B(n3988), .Z(n3990) );
  AND U4699 ( .A(n3991), .B(n3990), .Z(n4059) );
  AND U4700 ( .A(x[134]), .B(y[683]), .Z(n4363) );
  IV U4701 ( .A(n4363), .Z(n4432) );
  AND U4702 ( .A(x[129]), .B(y[678]), .Z(n4073) );
  NANDN U4703 ( .A(n4432), .B(n4073), .Z(n3995) );
  NAND U4704 ( .A(n3993), .B(n3992), .Z(n3994) );
  AND U4705 ( .A(n3995), .B(n3994), .Z(n4065) );
  AND U4706 ( .A(x[140]), .B(y[684]), .Z(n5274) );
  NAND U4707 ( .A(n5274), .B(n4205), .Z(n3999) );
  NAND U4708 ( .A(n3997), .B(n3996), .Z(n3998) );
  AND U4709 ( .A(n3999), .B(n3998), .Z(n4063) );
  AND U4710 ( .A(x[138]), .B(y[675]), .Z(n4886) );
  AND U4711 ( .A(y[677]), .B(x[136]), .Z(n4001) );
  NAND U4712 ( .A(y[674]), .B(x[139]), .Z(n4000) );
  XOR U4713 ( .A(n4001), .B(n4000), .Z(n4070) );
  XNOR U4714 ( .A(n4886), .B(n4070), .Z(n4062) );
  AND U4715 ( .A(x[138]), .B(y[680]), .Z(n4003) );
  AND U4716 ( .A(x[132]), .B(y[674]), .Z(n4002) );
  NAND U4717 ( .A(n4003), .B(n4002), .Z(n4006) );
  NANDN U4718 ( .A(n4004), .B(n4609), .Z(n4005) );
  AND U4719 ( .A(n4006), .B(n4005), .Z(n4107) );
  AND U4720 ( .A(y[685]), .B(x[128]), .Z(n4008) );
  NAND U4721 ( .A(y[672]), .B(x[141]), .Z(n4007) );
  XNOR U4722 ( .A(n4008), .B(n4007), .Z(n4099) );
  NAND U4723 ( .A(x[140]), .B(y[673]), .Z(n4092) );
  XNOR U4724 ( .A(o[45]), .B(n4092), .Z(n4098) );
  XOR U4725 ( .A(n4099), .B(n4098), .Z(n4105) );
  AND U4726 ( .A(y[680]), .B(x[133]), .Z(n4010) );
  NAND U4727 ( .A(y[682]), .B(x[131]), .Z(n4009) );
  XNOR U4728 ( .A(n4010), .B(n4009), .Z(n4094) );
  NAND U4729 ( .A(x[132]), .B(y[681]), .Z(n4095) );
  XNOR U4730 ( .A(n4094), .B(n4095), .Z(n4104) );
  XOR U4731 ( .A(n4105), .B(n4104), .Z(n4106) );
  XOR U4732 ( .A(n4057), .B(n4056), .Z(n4058) );
  XOR U4733 ( .A(n4047), .B(n4046), .Z(n4032) );
  NAND U4734 ( .A(n4012), .B(n4011), .Z(n4016) );
  NANDN U4735 ( .A(n4014), .B(n4013), .Z(n4015) );
  AND U4736 ( .A(n4016), .B(n4015), .Z(n4031) );
  XNOR U4737 ( .A(n4032), .B(n4031), .Z(n4033) );
  XNOR U4738 ( .A(n4034), .B(n4033), .Z(n4040) );
  OR U4739 ( .A(n4019), .B(n4017), .Z(n4023) );
  ANDN U4740 ( .B(n4019), .A(n4018), .Z(n4021) );
  OR U4741 ( .A(n4021), .B(n4020), .Z(n4022) );
  AND U4742 ( .A(n4023), .B(n4022), .Z(n4039) );
  NANDN U4743 ( .A(n4025), .B(n4024), .Z(n4029) );
  NAND U4744 ( .A(n4027), .B(n4026), .Z(n4028) );
  AND U4745 ( .A(n4029), .B(n4028), .Z(n4038) );
  IV U4746 ( .A(n4038), .Z(n4037) );
  XOR U4747 ( .A(n4039), .B(n4037), .Z(n4030) );
  XNOR U4748 ( .A(n4040), .B(n4030), .Z(N110) );
  NANDN U4749 ( .A(n4032), .B(n4031), .Z(n4036) );
  NANDN U4750 ( .A(n4034), .B(n4033), .Z(n4035) );
  NAND U4751 ( .A(n4036), .B(n4035), .Z(n4188) );
  IV U4752 ( .A(n4188), .Z(n4186) );
  OR U4753 ( .A(n4039), .B(n4037), .Z(n4043) );
  ANDN U4754 ( .B(n4039), .A(n4038), .Z(n4041) );
  OR U4755 ( .A(n4041), .B(n4040), .Z(n4042) );
  AND U4756 ( .A(n4043), .B(n4042), .Z(n4187) );
  NAND U4757 ( .A(n4045), .B(n4044), .Z(n4049) );
  NAND U4758 ( .A(n4047), .B(n4046), .Z(n4048) );
  NAND U4759 ( .A(n4049), .B(n4048), .Z(n4194) );
  NAND U4760 ( .A(n4051), .B(n4050), .Z(n4055) );
  NAND U4761 ( .A(n4053), .B(n4052), .Z(n4054) );
  NAND U4762 ( .A(n4055), .B(n4054), .Z(n4193) );
  XOR U4763 ( .A(n4194), .B(n4193), .Z(n4195) );
  NAND U4764 ( .A(n4057), .B(n4056), .Z(n4061) );
  NANDN U4765 ( .A(n4059), .B(n4058), .Z(n4060) );
  AND U4766 ( .A(n4061), .B(n4060), .Z(n4114) );
  NANDN U4767 ( .A(n4063), .B(n4062), .Z(n4067) );
  NANDN U4768 ( .A(n4065), .B(n4064), .Z(n4066) );
  AND U4769 ( .A(n4067), .B(n4066), .Z(n4120) );
  AND U4770 ( .A(x[139]), .B(y[677]), .Z(n4069) );
  NAND U4771 ( .A(n4069), .B(n4068), .Z(n4072) );
  NANDN U4772 ( .A(n4070), .B(n4886), .Z(n4071) );
  AND U4773 ( .A(n4072), .B(n4071), .Z(n4175) );
  NAND U4774 ( .A(x[135]), .B(y[684]), .Z(n4624) );
  NANDN U4775 ( .A(n4624), .B(n4073), .Z(n4077) );
  NAND U4776 ( .A(n4075), .B(n4074), .Z(n4076) );
  NAND U4777 ( .A(n4077), .B(n4076), .Z(n4174) );
  XNOR U4778 ( .A(n4175), .B(n4174), .Z(n4177) );
  AND U4779 ( .A(x[132]), .B(y[682]), .Z(n4543) );
  AND U4780 ( .A(y[683]), .B(x[131]), .Z(n4079) );
  NAND U4781 ( .A(y[678]), .B(x[136]), .Z(n4078) );
  XOR U4782 ( .A(n4079), .B(n4078), .Z(n4160) );
  XNOR U4783 ( .A(n4430), .B(n4160), .Z(n4169) );
  XOR U4784 ( .A(n4543), .B(n4169), .Z(n4171) );
  AND U4785 ( .A(x[137]), .B(y[677]), .Z(n4722) );
  AND U4786 ( .A(y[684]), .B(x[130]), .Z(n4080) );
  AND U4787 ( .A(y[676]), .B(x[138]), .Z(n4752) );
  XOR U4788 ( .A(n4080), .B(n4752), .Z(n4145) );
  XOR U4789 ( .A(n4722), .B(n4145), .Z(n4170) );
  XOR U4790 ( .A(n4171), .B(n4170), .Z(n4176) );
  XOR U4791 ( .A(n4177), .B(n4176), .Z(n4118) );
  NAND U4792 ( .A(n4082), .B(n4081), .Z(n4086) );
  NANDN U4793 ( .A(n4084), .B(n4083), .Z(n4085) );
  AND U4794 ( .A(n4086), .B(n4085), .Z(n4117) );
  XOR U4795 ( .A(n4120), .B(n4119), .Z(n4112) );
  AND U4796 ( .A(x[137]), .B(y[683]), .Z(n4622) );
  NAND U4797 ( .A(n4622), .B(n4144), .Z(n4089) );
  NANDN U4798 ( .A(n4087), .B(n5058), .Z(n4088) );
  AND U4799 ( .A(n4089), .B(n4088), .Z(n4132) );
  AND U4800 ( .A(y[686]), .B(x[128]), .Z(n4091) );
  NAND U4801 ( .A(y[672]), .B(x[142]), .Z(n4090) );
  XNOR U4802 ( .A(n4091), .B(n4090), .Z(n4155) );
  ANDN U4803 ( .B(o[45]), .A(n4092), .Z(n4154) );
  XOR U4804 ( .A(n4155), .B(n4154), .Z(n4130) );
  AND U4805 ( .A(y[674]), .B(x[140]), .Z(n4712) );
  NAND U4806 ( .A(y[679]), .B(x[135]), .Z(n4093) );
  XNOR U4807 ( .A(n4712), .B(n4093), .Z(n4137) );
  NAND U4808 ( .A(x[141]), .B(y[673]), .Z(n4143) );
  XNOR U4809 ( .A(o[46]), .B(n4143), .Z(n4136) );
  XOR U4810 ( .A(n4137), .B(n4136), .Z(n4129) );
  XOR U4811 ( .A(n4130), .B(n4129), .Z(n4131) );
  XOR U4812 ( .A(n4132), .B(n4131), .Z(n4181) );
  AND U4813 ( .A(x[133]), .B(y[682]), .Z(n4218) );
  NAND U4814 ( .A(n4874), .B(n4218), .Z(n4097) );
  NANDN U4815 ( .A(n4095), .B(n4094), .Z(n4096) );
  AND U4816 ( .A(n4097), .B(n4096), .Z(n4126) );
  AND U4817 ( .A(x[141]), .B(y[685]), .Z(n5605) );
  NAND U4818 ( .A(n5605), .B(n4205), .Z(n4101) );
  NAND U4819 ( .A(n4099), .B(n4098), .Z(n4100) );
  AND U4820 ( .A(n4101), .B(n4100), .Z(n4124) );
  NAND U4821 ( .A(y[675]), .B(x[139]), .Z(n4102) );
  XNOR U4822 ( .A(n4103), .B(n4102), .Z(n4151) );
  AND U4823 ( .A(x[129]), .B(y[685]), .Z(n4150) );
  XOR U4824 ( .A(n4151), .B(n4150), .Z(n4123) );
  XNOR U4825 ( .A(n4124), .B(n4123), .Z(n4125) );
  XOR U4826 ( .A(n4126), .B(n4125), .Z(n4180) );
  XOR U4827 ( .A(n4181), .B(n4180), .Z(n4183) );
  NAND U4828 ( .A(n4105), .B(n4104), .Z(n4109) );
  NANDN U4829 ( .A(n4107), .B(n4106), .Z(n4108) );
  AND U4830 ( .A(n4109), .B(n4108), .Z(n4182) );
  XNOR U4831 ( .A(n4183), .B(n4182), .Z(n4111) );
  XNOR U4832 ( .A(n4195), .B(n4196), .Z(n4189) );
  XNOR U4833 ( .A(n4187), .B(n4189), .Z(n4110) );
  XOR U4834 ( .A(n4186), .B(n4110), .Z(N111) );
  NANDN U4835 ( .A(n4112), .B(n4111), .Z(n4116) );
  NANDN U4836 ( .A(n4114), .B(n4113), .Z(n4115) );
  AND U4837 ( .A(n4116), .B(n4115), .Z(n4285) );
  NANDN U4838 ( .A(n4118), .B(n4117), .Z(n4122) );
  NAND U4839 ( .A(n4120), .B(n4119), .Z(n4121) );
  AND U4840 ( .A(n4122), .B(n4121), .Z(n4261) );
  NANDN U4841 ( .A(n4124), .B(n4123), .Z(n4128) );
  NANDN U4842 ( .A(n4126), .B(n4125), .Z(n4127) );
  NAND U4843 ( .A(n4128), .B(n4127), .Z(n4266) );
  NAND U4844 ( .A(n4130), .B(n4129), .Z(n4134) );
  NANDN U4845 ( .A(n4132), .B(n4131), .Z(n4133) );
  NAND U4846 ( .A(n4134), .B(n4133), .Z(n4264) );
  NAND U4847 ( .A(x[140]), .B(y[679]), .Z(n4616) );
  NANDN U4848 ( .A(n4616), .B(n4135), .Z(n4139) );
  NAND U4849 ( .A(n4137), .B(n4136), .Z(n4138) );
  AND U4850 ( .A(n4139), .B(n4138), .Z(n4241) );
  AND U4851 ( .A(y[674]), .B(x[141]), .Z(n5046) );
  NAND U4852 ( .A(y[676]), .B(x[139]), .Z(n4140) );
  XNOR U4853 ( .A(n5046), .B(n4140), .Z(n4245) );
  AND U4854 ( .A(x[140]), .B(y[675]), .Z(n4244) );
  XOR U4855 ( .A(n4245), .B(n4244), .Z(n4239) );
  AND U4856 ( .A(y[687]), .B(x[128]), .Z(n4142) );
  NAND U4857 ( .A(y[672]), .B(x[143]), .Z(n4141) );
  XNOR U4858 ( .A(n4142), .B(n4141), .Z(n4207) );
  ANDN U4859 ( .B(o[46]), .A(n4143), .Z(n4206) );
  XNOR U4860 ( .A(n4207), .B(n4206), .Z(n4238) );
  XNOR U4861 ( .A(n4239), .B(n4238), .Z(n4240) );
  XNOR U4862 ( .A(n4241), .B(n4240), .Z(n4272) );
  NAND U4863 ( .A(x[138]), .B(y[684]), .Z(n5060) );
  NANDN U4864 ( .A(n5060), .B(n4144), .Z(n4147) );
  NAND U4865 ( .A(n4722), .B(n4145), .Z(n4146) );
  NAND U4866 ( .A(n4147), .B(n4146), .Z(n4271) );
  AND U4867 ( .A(x[139]), .B(y[680]), .Z(n4149) );
  AND U4868 ( .A(x[134]), .B(y[675]), .Z(n4148) );
  NAND U4869 ( .A(n4149), .B(n4148), .Z(n4153) );
  NAND U4870 ( .A(n4151), .B(n4150), .Z(n4152) );
  NAND U4871 ( .A(n4153), .B(n4152), .Z(n4270) );
  XNOR U4872 ( .A(n4271), .B(n4270), .Z(n4273) );
  XOR U4873 ( .A(n4272), .B(n4273), .Z(n4265) );
  XOR U4874 ( .A(n4264), .B(n4265), .Z(n4267) );
  XOR U4875 ( .A(n4266), .B(n4267), .Z(n4258) );
  AND U4876 ( .A(x[142]), .B(y[686]), .Z(n5867) );
  NAND U4877 ( .A(n5867), .B(n4205), .Z(n4157) );
  NAND U4878 ( .A(n4155), .B(n4154), .Z(n4156) );
  AND U4879 ( .A(n4157), .B(n4156), .Z(n4233) );
  AND U4880 ( .A(x[136]), .B(y[683]), .Z(n4158) );
  NANDN U4881 ( .A(n4159), .B(n4158), .Z(n4162) );
  NANDN U4882 ( .A(n4160), .B(n4430), .Z(n4161) );
  NAND U4883 ( .A(n4162), .B(n4161), .Z(n4232) );
  XNOR U4884 ( .A(n4233), .B(n4232), .Z(n4235) );
  AND U4885 ( .A(y[683]), .B(x[132]), .Z(n4164) );
  NAND U4886 ( .A(y[677]), .B(x[138]), .Z(n4163) );
  XNOR U4887 ( .A(n4164), .B(n4163), .Z(n4213) );
  AND U4888 ( .A(x[135]), .B(y[680]), .Z(n4212) );
  XOR U4889 ( .A(n4213), .B(n4212), .Z(n4220) );
  NAND U4890 ( .A(x[134]), .B(y[681]), .Z(n4319) );
  XNOR U4891 ( .A(n4319), .B(n4218), .Z(n4219) );
  XOR U4892 ( .A(n4220), .B(n4219), .Z(n4254) );
  AND U4893 ( .A(y[678]), .B(x[137]), .Z(n4166) );
  NAND U4894 ( .A(y[685]), .B(x[130]), .Z(n4165) );
  XNOR U4895 ( .A(n4166), .B(n4165), .Z(n4223) );
  NAND U4896 ( .A(x[131]), .B(y[684]), .Z(n4224) );
  XNOR U4897 ( .A(n4223), .B(n4224), .Z(n4253) );
  AND U4898 ( .A(y[686]), .B(x[129]), .Z(n4168) );
  NAND U4899 ( .A(y[679]), .B(x[136]), .Z(n4167) );
  XNOR U4900 ( .A(n4168), .B(n4167), .Z(n4201) );
  NAND U4901 ( .A(x[142]), .B(y[673]), .Z(n4229) );
  XOR U4902 ( .A(o[47]), .B(n4229), .Z(n4202) );
  XNOR U4903 ( .A(n4201), .B(n4202), .Z(n4252) );
  XOR U4904 ( .A(n4253), .B(n4252), .Z(n4255) );
  XOR U4905 ( .A(n4254), .B(n4255), .Z(n4234) );
  XOR U4906 ( .A(n4235), .B(n4234), .Z(n4277) );
  NAND U4907 ( .A(n4543), .B(n4169), .Z(n4173) );
  NAND U4908 ( .A(n4171), .B(n4170), .Z(n4172) );
  AND U4909 ( .A(n4173), .B(n4172), .Z(n4276) );
  XNOR U4910 ( .A(n4277), .B(n4276), .Z(n4279) );
  NANDN U4911 ( .A(n4175), .B(n4174), .Z(n4179) );
  NAND U4912 ( .A(n4177), .B(n4176), .Z(n4178) );
  AND U4913 ( .A(n4179), .B(n4178), .Z(n4278) );
  XOR U4914 ( .A(n4279), .B(n4278), .Z(n4259) );
  XOR U4915 ( .A(n4258), .B(n4259), .Z(n4260) );
  NAND U4916 ( .A(n4181), .B(n4180), .Z(n4185) );
  NAND U4917 ( .A(n4183), .B(n4182), .Z(n4184) );
  AND U4918 ( .A(n4185), .B(n4184), .Z(n4283) );
  XOR U4919 ( .A(n4282), .B(n4283), .Z(n4284) );
  XOR U4920 ( .A(n4285), .B(n4284), .Z(n4290) );
  NANDN U4921 ( .A(n4186), .B(n4187), .Z(n4192) );
  NOR U4922 ( .A(n4188), .B(n4187), .Z(n4190) );
  OR U4923 ( .A(n4190), .B(n4189), .Z(n4191) );
  AND U4924 ( .A(n4192), .B(n4191), .Z(n4289) );
  NAND U4925 ( .A(n4194), .B(n4193), .Z(n4198) );
  NANDN U4926 ( .A(n4196), .B(n4195), .Z(n4197) );
  NAND U4927 ( .A(n4198), .B(n4197), .Z(n4288) );
  XOR U4928 ( .A(n4289), .B(n4288), .Z(n4199) );
  XNOR U4929 ( .A(n4290), .B(n4199), .Z(N112) );
  AND U4930 ( .A(x[136]), .B(y[686]), .Z(n4895) );
  NAND U4931 ( .A(n4895), .B(n4200), .Z(n4204) );
  NANDN U4932 ( .A(n4202), .B(n4201), .Z(n4203) );
  NAND U4933 ( .A(n4204), .B(n4203), .Z(n4343) );
  AND U4934 ( .A(x[143]), .B(y[687]), .Z(n6261) );
  NAND U4935 ( .A(n6261), .B(n4205), .Z(n4209) );
  NAND U4936 ( .A(n4207), .B(n4206), .Z(n4208) );
  NAND U4937 ( .A(n4209), .B(n4208), .Z(n4342) );
  XOR U4938 ( .A(n4343), .B(n4342), .Z(n4345) );
  AND U4939 ( .A(x[138]), .B(y[683]), .Z(n4211) );
  NAND U4940 ( .A(n4211), .B(n4210), .Z(n4215) );
  NAND U4941 ( .A(n4213), .B(n4212), .Z(n4214) );
  AND U4942 ( .A(n4215), .B(n4214), .Z(n4307) );
  AND U4943 ( .A(x[128]), .B(y[688]), .Z(n4325) );
  AND U4944 ( .A(x[144]), .B(y[672]), .Z(n4324) );
  XOR U4945 ( .A(n4325), .B(n4324), .Z(n4327) );
  AND U4946 ( .A(x[143]), .B(y[673]), .Z(n4316) );
  XOR U4947 ( .A(n4316), .B(o[48]), .Z(n4326) );
  XOR U4948 ( .A(n4327), .B(n4326), .Z(n4305) );
  NAND U4949 ( .A(y[681]), .B(x[135]), .Z(n4216) );
  XNOR U4950 ( .A(n4217), .B(n4216), .Z(n4321) );
  AND U4951 ( .A(x[138]), .B(y[678]), .Z(n4320) );
  XOR U4952 ( .A(n4321), .B(n4320), .Z(n4304) );
  XOR U4953 ( .A(n4305), .B(n4304), .Z(n4306) );
  XOR U4954 ( .A(n4345), .B(n4344), .Z(n4301) );
  NANDN U4955 ( .A(n4218), .B(n4319), .Z(n4222) );
  NANDN U4956 ( .A(n4220), .B(n4219), .Z(n4221) );
  AND U4957 ( .A(n4222), .B(n4221), .Z(n4299) );
  NAND U4958 ( .A(x[137]), .B(y[685]), .Z(n5042) );
  NANDN U4959 ( .A(n5042), .B(n4614), .Z(n4226) );
  NANDN U4960 ( .A(n4224), .B(n4223), .Z(n4225) );
  AND U4961 ( .A(n4226), .B(n4225), .Z(n4333) );
  AND U4962 ( .A(y[687]), .B(x[129]), .Z(n4228) );
  NAND U4963 ( .A(y[680]), .B(x[136]), .Z(n4227) );
  XNOR U4964 ( .A(n4228), .B(n4227), .Z(n4323) );
  ANDN U4965 ( .B(o[47]), .A(n4229), .Z(n4322) );
  XOR U4966 ( .A(n4323), .B(n4322), .Z(n4330) );
  AND U4967 ( .A(y[674]), .B(x[142]), .Z(n4231) );
  NAND U4968 ( .A(y[677]), .B(x[139]), .Z(n4230) );
  XNOR U4969 ( .A(n4231), .B(n4230), .Z(n4354) );
  NAND U4970 ( .A(x[132]), .B(y[684]), .Z(n4355) );
  XOR U4971 ( .A(n4354), .B(n4355), .Z(n4331) );
  XOR U4972 ( .A(n4333), .B(n4332), .Z(n4298) );
  XNOR U4973 ( .A(n4299), .B(n4298), .Z(n4300) );
  XNOR U4974 ( .A(n4301), .B(n4300), .Z(n4336) );
  NANDN U4975 ( .A(n4233), .B(n4232), .Z(n4237) );
  NAND U4976 ( .A(n4235), .B(n4234), .Z(n4236) );
  NAND U4977 ( .A(n4237), .B(n4236), .Z(n4337) );
  XNOR U4978 ( .A(n4336), .B(n4337), .Z(n4339) );
  NANDN U4979 ( .A(n4239), .B(n4238), .Z(n4243) );
  NAND U4980 ( .A(n4241), .B(n4240), .Z(n4242) );
  AND U4981 ( .A(n4243), .B(n4242), .Z(n4369) );
  AND U4982 ( .A(x[139]), .B(y[674]), .Z(n4851) );
  AND U4983 ( .A(x[141]), .B(y[676]), .Z(n4365) );
  NAND U4984 ( .A(n4851), .B(n4365), .Z(n4247) );
  NAND U4985 ( .A(n4245), .B(n4244), .Z(n4246) );
  AND U4986 ( .A(n4247), .B(n4246), .Z(n4351) );
  AND U4987 ( .A(y[679]), .B(x[137]), .Z(n4249) );
  NAND U4988 ( .A(y[686]), .B(x[130]), .Z(n4248) );
  XNOR U4989 ( .A(n4249), .B(n4248), .Z(n4358) );
  NAND U4990 ( .A(x[131]), .B(y[685]), .Z(n4359) );
  XNOR U4991 ( .A(n4358), .B(n4359), .Z(n4348) );
  AND U4992 ( .A(x[140]), .B(y[676]), .Z(n5030) );
  AND U4993 ( .A(y[683]), .B(x[133]), .Z(n4251) );
  NAND U4994 ( .A(y[675]), .B(x[141]), .Z(n4250) );
  XOR U4995 ( .A(n4251), .B(n4250), .Z(n4311) );
  XOR U4996 ( .A(n5030), .B(n4311), .Z(n4349) );
  NAND U4997 ( .A(n4253), .B(n4252), .Z(n4257) );
  NAND U4998 ( .A(n4255), .B(n4254), .Z(n4256) );
  AND U4999 ( .A(n4257), .B(n4256), .Z(n4367) );
  XOR U5000 ( .A(n4366), .B(n4367), .Z(n4368) );
  XOR U5001 ( .A(n4339), .B(n4338), .Z(n4376) );
  NAND U5002 ( .A(n4259), .B(n4258), .Z(n4263) );
  NANDN U5003 ( .A(n4261), .B(n4260), .Z(n4262) );
  AND U5004 ( .A(n4263), .B(n4262), .Z(n4375) );
  NANDN U5005 ( .A(n4265), .B(n4264), .Z(n4269) );
  NANDN U5006 ( .A(n4267), .B(n4266), .Z(n4268) );
  NAND U5007 ( .A(n4269), .B(n4268), .Z(n4294) );
  NAND U5008 ( .A(n4271), .B(n4270), .Z(n4275) );
  NANDN U5009 ( .A(n4273), .B(n4272), .Z(n4274) );
  NAND U5010 ( .A(n4275), .B(n4274), .Z(n4292) );
  NANDN U5011 ( .A(n4277), .B(n4276), .Z(n4281) );
  NAND U5012 ( .A(n4279), .B(n4278), .Z(n4280) );
  AND U5013 ( .A(n4281), .B(n4280), .Z(n4293) );
  XOR U5014 ( .A(n4292), .B(n4293), .Z(n4295) );
  XOR U5015 ( .A(n4294), .B(n4295), .Z(n4377) );
  XNOR U5016 ( .A(n4378), .B(n4377), .Z(n4374) );
  NAND U5017 ( .A(n4283), .B(n4282), .Z(n4287) );
  NANDN U5018 ( .A(n4285), .B(n4284), .Z(n4286) );
  NAND U5019 ( .A(n4287), .B(n4286), .Z(n4372) );
  XOR U5020 ( .A(n4372), .B(n4373), .Z(n4291) );
  XNOR U5021 ( .A(n4374), .B(n4291), .Z(N113) );
  NAND U5022 ( .A(n4293), .B(n4292), .Z(n4297) );
  NAND U5023 ( .A(n4295), .B(n4294), .Z(n4296) );
  NAND U5024 ( .A(n4297), .B(n4296), .Z(n4479) );
  NANDN U5025 ( .A(n4299), .B(n4298), .Z(n4303) );
  NANDN U5026 ( .A(n4301), .B(n4300), .Z(n4302) );
  AND U5027 ( .A(n4303), .B(n4302), .Z(n4391) );
  NAND U5028 ( .A(n4305), .B(n4304), .Z(n4309) );
  NANDN U5029 ( .A(n4307), .B(n4306), .Z(n4308) );
  NAND U5030 ( .A(n4309), .B(n4308), .Z(n4466) );
  AND U5031 ( .A(x[141]), .B(y[683]), .Z(n5282) );
  NAND U5032 ( .A(n5282), .B(n4310), .Z(n4313) );
  NANDN U5033 ( .A(n4311), .B(n5030), .Z(n4312) );
  NAND U5034 ( .A(n4313), .B(n4312), .Z(n4420) );
  AND U5035 ( .A(y[680]), .B(x[137]), .Z(n4315) );
  NAND U5036 ( .A(y[688]), .B(x[129]), .Z(n4314) );
  XNOR U5037 ( .A(n4315), .B(n4314), .Z(n4435) );
  NAND U5038 ( .A(n4316), .B(o[48]), .Z(n4436) );
  XNOR U5039 ( .A(n4435), .B(n4436), .Z(n4419) );
  AND U5040 ( .A(y[674]), .B(x[143]), .Z(n4318) );
  NAND U5041 ( .A(y[677]), .B(x[140]), .Z(n4317) );
  XNOR U5042 ( .A(n4318), .B(n4317), .Z(n4396) );
  AND U5043 ( .A(x[142]), .B(y[675]), .Z(n4395) );
  XOR U5044 ( .A(n4396), .B(n4395), .Z(n4418) );
  XOR U5045 ( .A(n4419), .B(n4418), .Z(n4421) );
  XOR U5046 ( .A(n4420), .B(n4421), .Z(n4465) );
  NAND U5047 ( .A(x[135]), .B(y[682]), .Z(n4447) );
  AND U5048 ( .A(x[136]), .B(y[687]), .Z(n5090) );
  XOR U5049 ( .A(n4426), .B(n4427), .Z(n4428) );
  AND U5050 ( .A(x[128]), .B(y[689]), .Z(n4410) );
  AND U5051 ( .A(x[145]), .B(y[672]), .Z(n4409) );
  XOR U5052 ( .A(n4410), .B(n4409), .Z(n4412) );
  AND U5053 ( .A(x[144]), .B(y[673]), .Z(n4406) );
  XOR U5054 ( .A(n4406), .B(o[49]), .Z(n4411) );
  XOR U5055 ( .A(n4412), .B(n4411), .Z(n4423) );
  AND U5056 ( .A(y[687]), .B(x[130]), .Z(n4329) );
  NAND U5057 ( .A(y[679]), .B(x[138]), .Z(n4328) );
  XNOR U5058 ( .A(n4329), .B(n4328), .Z(n4440) );
  NAND U5059 ( .A(x[131]), .B(y[686]), .Z(n4441) );
  XNOR U5060 ( .A(n4440), .B(n4441), .Z(n4422) );
  XOR U5061 ( .A(n4423), .B(n4422), .Z(n4424) );
  XNOR U5062 ( .A(n4425), .B(n4424), .Z(n4429) );
  XNOR U5063 ( .A(n4428), .B(n4429), .Z(n4464) );
  XOR U5064 ( .A(n4465), .B(n4464), .Z(n4467) );
  XNOR U5065 ( .A(n4466), .B(n4467), .Z(n4388) );
  NANDN U5066 ( .A(n4331), .B(n4330), .Z(n4335) );
  NANDN U5067 ( .A(n4333), .B(n4332), .Z(n4334) );
  AND U5068 ( .A(n4335), .B(n4334), .Z(n4389) );
  XOR U5069 ( .A(n4388), .B(n4389), .Z(n4390) );
  NANDN U5070 ( .A(n4337), .B(n4336), .Z(n4341) );
  NAND U5071 ( .A(n4339), .B(n4338), .Z(n4340) );
  NAND U5072 ( .A(n4341), .B(n4340), .Z(n4385) );
  NAND U5073 ( .A(n4343), .B(n4342), .Z(n4347) );
  NAND U5074 ( .A(n4345), .B(n4344), .Z(n4346) );
  AND U5075 ( .A(n4347), .B(n4346), .Z(n4461) );
  NANDN U5076 ( .A(n4349), .B(n4348), .Z(n4353) );
  NANDN U5077 ( .A(n4351), .B(n4350), .Z(n4352) );
  AND U5078 ( .A(n4353), .B(n4352), .Z(n4459) );
  NAND U5079 ( .A(x[142]), .B(y[677]), .Z(n4646) );
  NANDN U5080 ( .A(n4646), .B(n4851), .Z(n4357) );
  NANDN U5081 ( .A(n4355), .B(n4354), .Z(n4356) );
  AND U5082 ( .A(n4357), .B(n4356), .Z(n4453) );
  AND U5083 ( .A(y[686]), .B(x[137]), .Z(n5263) );
  NAND U5084 ( .A(n4439), .B(n5263), .Z(n4361) );
  NANDN U5085 ( .A(n4359), .B(n4358), .Z(n4360) );
  NAND U5086 ( .A(n4361), .B(n4360), .Z(n4452) );
  XNOR U5087 ( .A(n4453), .B(n4452), .Z(n4454) );
  AND U5088 ( .A(x[133]), .B(y[684]), .Z(n4502) );
  NAND U5089 ( .A(y[681]), .B(x[136]), .Z(n4362) );
  XNOR U5090 ( .A(n4502), .B(n4362), .Z(n4431) );
  XOR U5091 ( .A(n4431), .B(n4363), .Z(n4446) );
  XNOR U5092 ( .A(n4446), .B(n4447), .Z(n4448) );
  NAND U5093 ( .A(y[685]), .B(x[132]), .Z(n4364) );
  XNOR U5094 ( .A(n4365), .B(n4364), .Z(n4400) );
  NAND U5095 ( .A(x[139]), .B(y[678]), .Z(n4401) );
  XOR U5096 ( .A(n4400), .B(n4401), .Z(n4449) );
  XOR U5097 ( .A(n4448), .B(n4449), .Z(n4455) );
  XNOR U5098 ( .A(n4454), .B(n4455), .Z(n4458) );
  NAND U5099 ( .A(n4367), .B(n4366), .Z(n4371) );
  NANDN U5100 ( .A(n4369), .B(n4368), .Z(n4370) );
  NAND U5101 ( .A(n4371), .B(n4370), .Z(n4382) );
  XOR U5102 ( .A(n4383), .B(n4382), .Z(n4384) );
  XNOR U5103 ( .A(n4385), .B(n4384), .Z(n4477) );
  XOR U5104 ( .A(n4478), .B(n4477), .Z(n4480) );
  XOR U5105 ( .A(n4479), .B(n4480), .Z(n4473) );
  NANDN U5106 ( .A(n4376), .B(n4375), .Z(n4380) );
  NAND U5107 ( .A(n4378), .B(n4377), .Z(n4379) );
  NAND U5108 ( .A(n4380), .B(n4379), .Z(n4471) );
  IV U5109 ( .A(n4471), .Z(n4470) );
  XOR U5110 ( .A(n4472), .B(n4470), .Z(n4381) );
  XNOR U5111 ( .A(n4473), .B(n4381), .Z(N114) );
  NAND U5112 ( .A(n4383), .B(n4382), .Z(n4387) );
  NAND U5113 ( .A(n4385), .B(n4384), .Z(n4386) );
  AND U5114 ( .A(n4387), .B(n4386), .Z(n4584) );
  NAND U5115 ( .A(n4389), .B(n4388), .Z(n4393) );
  NANDN U5116 ( .A(n4391), .B(n4390), .Z(n4392) );
  AND U5117 ( .A(n4393), .B(n4392), .Z(n4582) );
  AND U5118 ( .A(x[143]), .B(y[677]), .Z(n4394) );
  NAND U5119 ( .A(n4394), .B(n4712), .Z(n4398) );
  NAND U5120 ( .A(n4396), .B(n4395), .Z(n4397) );
  NAND U5121 ( .A(n4398), .B(n4397), .Z(n4567) );
  NAND U5122 ( .A(n5605), .B(n4399), .Z(n4403) );
  NANDN U5123 ( .A(n4401), .B(n4400), .Z(n4402) );
  AND U5124 ( .A(n4403), .B(n4402), .Z(n4560) );
  AND U5125 ( .A(y[689]), .B(x[129]), .Z(n4405) );
  NAND U5126 ( .A(y[680]), .B(x[138]), .Z(n4404) );
  XNOR U5127 ( .A(n4405), .B(n4404), .Z(n4522) );
  NAND U5128 ( .A(n4406), .B(o[49]), .Z(n4523) );
  XNOR U5129 ( .A(n4522), .B(n4523), .Z(n4558) );
  NAND U5130 ( .A(y[675]), .B(x[143]), .Z(n4407) );
  XNOR U5131 ( .A(n4408), .B(n4407), .Z(n4513) );
  NAND U5132 ( .A(x[142]), .B(y[676]), .Z(n4514) );
  XNOR U5133 ( .A(n4513), .B(n4514), .Z(n4557) );
  XOR U5134 ( .A(n4558), .B(n4557), .Z(n4559) );
  XOR U5135 ( .A(n4567), .B(n4568), .Z(n4570) );
  AND U5136 ( .A(y[679]), .B(x[139]), .Z(n4414) );
  NAND U5137 ( .A(y[674]), .B(x[144]), .Z(n4413) );
  XNOR U5138 ( .A(n4414), .B(n4413), .Z(n4509) );
  NAND U5139 ( .A(x[130]), .B(y[688]), .Z(n4510) );
  XOR U5140 ( .A(n4576), .B(n4575), .Z(n4578) );
  AND U5141 ( .A(y[685]), .B(x[133]), .Z(n4630) );
  NAND U5142 ( .A(y[684]), .B(x[134]), .Z(n4415) );
  XNOR U5143 ( .A(n4630), .B(n4415), .Z(n4505) );
  AND U5144 ( .A(y[686]), .B(x[132]), .Z(n4417) );
  NAND U5145 ( .A(y[682]), .B(x[136]), .Z(n4416) );
  XNOR U5146 ( .A(n4417), .B(n4416), .Z(n4544) );
  NAND U5147 ( .A(x[135]), .B(y[683]), .Z(n4545) );
  XNOR U5148 ( .A(n4544), .B(n4545), .Z(n4504) );
  XOR U5149 ( .A(n4505), .B(n4504), .Z(n4577) );
  XOR U5150 ( .A(n4578), .B(n4577), .Z(n4569) );
  XOR U5151 ( .A(n4570), .B(n4569), .Z(n4491) );
  XOR U5152 ( .A(n4564), .B(n4563), .Z(n4566) );
  XOR U5153 ( .A(n4566), .B(n4565), .Z(n4490) );
  AND U5154 ( .A(x[136]), .B(y[684]), .Z(n4758) );
  NAND U5155 ( .A(n4758), .B(n4430), .Z(n4434) );
  NANDN U5156 ( .A(n4432), .B(n4431), .Z(n4433) );
  NAND U5157 ( .A(n4434), .B(n4433), .Z(n4571) );
  AND U5158 ( .A(x[137]), .B(y[688]), .Z(n5384) );
  NAND U5159 ( .A(n5384), .B(n4521), .Z(n4438) );
  NANDN U5160 ( .A(n4436), .B(n4435), .Z(n4437) );
  NAND U5161 ( .A(n4438), .B(n4437), .Z(n4572) );
  XOR U5162 ( .A(n4571), .B(n4572), .Z(n4574) );
  AND U5163 ( .A(x[138]), .B(y[687]), .Z(n5383) );
  NAND U5164 ( .A(n5383), .B(n4439), .Z(n4443) );
  NANDN U5165 ( .A(n4441), .B(n4440), .Z(n4442) );
  AND U5166 ( .A(n4443), .B(n4442), .Z(n4554) );
  AND U5167 ( .A(x[128]), .B(y[690]), .Z(n4526) );
  NAND U5168 ( .A(x[146]), .B(y[672]), .Z(n4527) );
  XNOR U5169 ( .A(n4526), .B(n4527), .Z(n4528) );
  NAND U5170 ( .A(x[145]), .B(y[673]), .Z(n4548) );
  XOR U5171 ( .A(o[50]), .B(n4548), .Z(n4529) );
  XNOR U5172 ( .A(n4528), .B(n4529), .Z(n4552) );
  AND U5173 ( .A(y[687]), .B(x[131]), .Z(n4445) );
  NAND U5174 ( .A(y[677]), .B(x[141]), .Z(n4444) );
  XNOR U5175 ( .A(n4445), .B(n4444), .Z(n4535) );
  NAND U5176 ( .A(x[140]), .B(y[678]), .Z(n4536) );
  XNOR U5177 ( .A(n4535), .B(n4536), .Z(n4551) );
  XOR U5178 ( .A(n4552), .B(n4551), .Z(n4553) );
  XOR U5179 ( .A(n4574), .B(n4573), .Z(n4497) );
  NANDN U5180 ( .A(n4447), .B(n4446), .Z(n4451) );
  NANDN U5181 ( .A(n4449), .B(n4448), .Z(n4450) );
  AND U5182 ( .A(n4451), .B(n4450), .Z(n4496) );
  XNOR U5183 ( .A(n4497), .B(n4496), .Z(n4499) );
  NANDN U5184 ( .A(n4453), .B(n4452), .Z(n4457) );
  NANDN U5185 ( .A(n4455), .B(n4454), .Z(n4456) );
  AND U5186 ( .A(n4457), .B(n4456), .Z(n4498) );
  XOR U5187 ( .A(n4499), .B(n4498), .Z(n4492) );
  XOR U5188 ( .A(n4493), .B(n4492), .Z(n4487) );
  NANDN U5189 ( .A(n4459), .B(n4458), .Z(n4463) );
  NANDN U5190 ( .A(n4461), .B(n4460), .Z(n4462) );
  NAND U5191 ( .A(n4463), .B(n4462), .Z(n4485) );
  NAND U5192 ( .A(n4465), .B(n4464), .Z(n4469) );
  NAND U5193 ( .A(n4467), .B(n4466), .Z(n4468) );
  NAND U5194 ( .A(n4469), .B(n4468), .Z(n4484) );
  XOR U5195 ( .A(n4485), .B(n4484), .Z(n4486) );
  XOR U5196 ( .A(n4582), .B(n4581), .Z(n4583) );
  XNOR U5197 ( .A(n4584), .B(n4583), .Z(n4589) );
  OR U5198 ( .A(n4472), .B(n4470), .Z(n4476) );
  ANDN U5199 ( .B(n4472), .A(n4471), .Z(n4474) );
  OR U5200 ( .A(n4474), .B(n4473), .Z(n4475) );
  AND U5201 ( .A(n4476), .B(n4475), .Z(n4588) );
  NANDN U5202 ( .A(n4478), .B(n4477), .Z(n4482) );
  NANDN U5203 ( .A(n4480), .B(n4479), .Z(n4481) );
  NAND U5204 ( .A(n4482), .B(n4481), .Z(n4587) );
  XNOR U5205 ( .A(n4588), .B(n4587), .Z(n4483) );
  XNOR U5206 ( .A(n4589), .B(n4483), .Z(N115) );
  NAND U5207 ( .A(n4485), .B(n4484), .Z(n4489) );
  NANDN U5208 ( .A(n4487), .B(n4486), .Z(n4488) );
  NAND U5209 ( .A(n4489), .B(n4488), .Z(n4698) );
  NANDN U5210 ( .A(n4491), .B(n4490), .Z(n4495) );
  NAND U5211 ( .A(n4493), .B(n4492), .Z(n4494) );
  AND U5212 ( .A(n4495), .B(n4494), .Z(n4697) );
  NANDN U5213 ( .A(n4497), .B(n4496), .Z(n4501) );
  NAND U5214 ( .A(n4499), .B(n4498), .Z(n4500) );
  AND U5215 ( .A(n4501), .B(n4500), .Z(n4594) );
  AND U5216 ( .A(x[134]), .B(y[685]), .Z(n4503) );
  NAND U5217 ( .A(n4503), .B(n4502), .Z(n4507) );
  NAND U5218 ( .A(n4505), .B(n4504), .Z(n4506) );
  AND U5219 ( .A(n4507), .B(n4506), .Z(n4669) );
  AND U5220 ( .A(x[144]), .B(y[679]), .Z(n4508) );
  NAND U5221 ( .A(n4508), .B(n4851), .Z(n4512) );
  NANDN U5222 ( .A(n4510), .B(n4509), .Z(n4511) );
  AND U5223 ( .A(n4512), .B(n4511), .Z(n4667) );
  AND U5224 ( .A(x[143]), .B(y[681]), .Z(n5299) );
  NAND U5225 ( .A(n5299), .B(n4609), .Z(n4516) );
  NANDN U5226 ( .A(n4514), .B(n4513), .Z(n4515) );
  AND U5227 ( .A(n4516), .B(n4515), .Z(n4600) );
  AND U5228 ( .A(y[690]), .B(x[129]), .Z(n4518) );
  NAND U5229 ( .A(y[683]), .B(x[136]), .Z(n4517) );
  XNOR U5230 ( .A(n4518), .B(n4517), .Z(n4645) );
  XNOR U5231 ( .A(n4645), .B(n4646), .Z(n4598) );
  AND U5232 ( .A(y[689]), .B(x[130]), .Z(n4520) );
  NAND U5233 ( .A(y[678]), .B(x[141]), .Z(n4519) );
  XNOR U5234 ( .A(n4520), .B(n4519), .Z(n4615) );
  XOR U5235 ( .A(n4598), .B(n4597), .Z(n4599) );
  XNOR U5236 ( .A(n4600), .B(n4599), .Z(n4666) );
  AND U5237 ( .A(x[138]), .B(y[689]), .Z(n5705) );
  IV U5238 ( .A(n5705), .Z(n5566) );
  NANDN U5239 ( .A(n5566), .B(n4521), .Z(n4525) );
  NANDN U5240 ( .A(n4523), .B(n4522), .Z(n4524) );
  AND U5241 ( .A(n4525), .B(n4524), .Z(n4657) );
  NANDN U5242 ( .A(n4527), .B(n4526), .Z(n4531) );
  NANDN U5243 ( .A(n4529), .B(n4528), .Z(n4530) );
  AND U5244 ( .A(n4531), .B(n4530), .Z(n4655) );
  AND U5245 ( .A(y[682]), .B(x[137]), .Z(n4533) );
  NAND U5246 ( .A(y[675]), .B(x[144]), .Z(n4532) );
  XNOR U5247 ( .A(n4533), .B(n4532), .Z(n4610) );
  NAND U5248 ( .A(x[143]), .B(y[676]), .Z(n4611) );
  XNOR U5249 ( .A(n4610), .B(n4611), .Z(n4654) );
  XNOR U5250 ( .A(n4655), .B(n4654), .Z(n4656) );
  XOR U5251 ( .A(n4657), .B(n4656), .Z(n4674) );
  AND U5252 ( .A(x[141]), .B(y[687]), .Z(n5887) );
  NANDN U5253 ( .A(n4534), .B(n5887), .Z(n4538) );
  NANDN U5254 ( .A(n4536), .B(n4535), .Z(n4537) );
  AND U5255 ( .A(n4538), .B(n4537), .Z(n4663) );
  AND U5256 ( .A(y[674]), .B(x[145]), .Z(n4540) );
  NAND U5257 ( .A(y[681]), .B(x[138]), .Z(n4539) );
  XNOR U5258 ( .A(n4540), .B(n4539), .Z(n4650) );
  NAND U5259 ( .A(x[146]), .B(y[673]), .Z(n4629) );
  XOR U5260 ( .A(o[51]), .B(n4629), .Z(n4651) );
  XNOR U5261 ( .A(n4650), .B(n4651), .Z(n4661) );
  AND U5262 ( .A(y[688]), .B(x[131]), .Z(n4542) );
  NAND U5263 ( .A(y[680]), .B(x[139]), .Z(n4541) );
  XNOR U5264 ( .A(n4542), .B(n4541), .Z(n4623) );
  XOR U5265 ( .A(n4661), .B(n4660), .Z(n4662) );
  XOR U5266 ( .A(n4663), .B(n4662), .Z(n4673) );
  NAND U5267 ( .A(n4895), .B(n4543), .Z(n4547) );
  NANDN U5268 ( .A(n4545), .B(n4544), .Z(n4546) );
  AND U5269 ( .A(n4547), .B(n4546), .Z(n4606) );
  AND U5270 ( .A(x[128]), .B(y[691]), .Z(n4634) );
  NAND U5271 ( .A(x[147]), .B(y[672]), .Z(n4635) );
  XNOR U5272 ( .A(n4634), .B(n4635), .Z(n4637) );
  ANDN U5273 ( .B(o[50]), .A(n4548), .Z(n4636) );
  XOR U5274 ( .A(n4637), .B(n4636), .Z(n4603) );
  AND U5275 ( .A(x[132]), .B(y[687]), .Z(n4772) );
  AND U5276 ( .A(y[686]), .B(x[133]), .Z(n4550) );
  NAND U5277 ( .A(y[685]), .B(x[134]), .Z(n4549) );
  XOR U5278 ( .A(n4550), .B(n4549), .Z(n4631) );
  XOR U5279 ( .A(n4772), .B(n4631), .Z(n4604) );
  XNOR U5280 ( .A(n4603), .B(n4604), .Z(n4605) );
  XOR U5281 ( .A(n4606), .B(n4605), .Z(n4672) );
  XOR U5282 ( .A(n4673), .B(n4672), .Z(n4675) );
  XNOR U5283 ( .A(n4674), .B(n4675), .Z(n4680) );
  NAND U5284 ( .A(n4552), .B(n4551), .Z(n4556) );
  NANDN U5285 ( .A(n4554), .B(n4553), .Z(n4555) );
  AND U5286 ( .A(n4556), .B(n4555), .Z(n4679) );
  NAND U5287 ( .A(n4558), .B(n4557), .Z(n4562) );
  NANDN U5288 ( .A(n4560), .B(n4559), .Z(n4561) );
  NAND U5289 ( .A(n4562), .B(n4561), .Z(n4678) );
  XNOR U5290 ( .A(n4680), .B(n4681), .Z(n4591) );
  XOR U5291 ( .A(n4592), .B(n4591), .Z(n4593) );
  NAND U5292 ( .A(n4576), .B(n4575), .Z(n4580) );
  NAND U5293 ( .A(n4578), .B(n4577), .Z(n4579) );
  NAND U5294 ( .A(n4580), .B(n4579), .Z(n4684) );
  XNOR U5295 ( .A(n4685), .B(n4684), .Z(n4687) );
  XOR U5296 ( .A(n4686), .B(n4687), .Z(n4691) );
  XNOR U5297 ( .A(n4690), .B(n4691), .Z(n4692) );
  XNOR U5298 ( .A(n4693), .B(n4692), .Z(n4696) );
  XOR U5299 ( .A(n4697), .B(n4696), .Z(n4699) );
  XNOR U5300 ( .A(n4698), .B(n4699), .Z(n4704) );
  NAND U5301 ( .A(n4582), .B(n4581), .Z(n4586) );
  NAND U5302 ( .A(n4584), .B(n4583), .Z(n4585) );
  NAND U5303 ( .A(n4586), .B(n4585), .Z(n4702) );
  XOR U5304 ( .A(n4702), .B(n4703), .Z(n4590) );
  XNOR U5305 ( .A(n4704), .B(n4590), .Z(N116) );
  NAND U5306 ( .A(n4592), .B(n4591), .Z(n4596) );
  NANDN U5307 ( .A(n4594), .B(n4593), .Z(n4595) );
  AND U5308 ( .A(n4596), .B(n4595), .Z(n4806) );
  NAND U5309 ( .A(n4598), .B(n4597), .Z(n4602) );
  NANDN U5310 ( .A(n4600), .B(n4599), .Z(n4601) );
  NAND U5311 ( .A(n4602), .B(n4601), .Z(n4707) );
  NANDN U5312 ( .A(n4604), .B(n4603), .Z(n4608) );
  NANDN U5313 ( .A(n4606), .B(n4605), .Z(n4607) );
  NAND U5314 ( .A(n4608), .B(n4607), .Z(n4706) );
  XOR U5315 ( .A(n4707), .B(n4706), .Z(n4709) );
  AND U5316 ( .A(x[144]), .B(y[682]), .Z(n5525) );
  NAND U5317 ( .A(n5525), .B(n4609), .Z(n4613) );
  NANDN U5318 ( .A(n4611), .B(n4610), .Z(n4612) );
  AND U5319 ( .A(n4613), .B(n4612), .Z(n4747) );
  AND U5320 ( .A(x[141]), .B(y[689]), .Z(n6086) );
  NAND U5321 ( .A(n6086), .B(n4614), .Z(n4618) );
  NANDN U5322 ( .A(n4616), .B(n4615), .Z(n4617) );
  AND U5323 ( .A(n4618), .B(n4617), .Z(n4790) );
  NAND U5324 ( .A(y[676]), .B(x[144]), .Z(n4619) );
  XNOR U5325 ( .A(n4620), .B(n4619), .Z(n4753) );
  NAND U5326 ( .A(x[130]), .B(y[690]), .Z(n4754) );
  XNOR U5327 ( .A(n4753), .B(n4754), .Z(n4787) );
  NAND U5328 ( .A(y[677]), .B(x[143]), .Z(n4621) );
  XNOR U5329 ( .A(n4622), .B(n4621), .Z(n4723) );
  NAND U5330 ( .A(x[142]), .B(y[678]), .Z(n4724) );
  XOR U5331 ( .A(n4723), .B(n4724), .Z(n4788) );
  XNOR U5332 ( .A(n4787), .B(n4788), .Z(n4789) );
  XNOR U5333 ( .A(n4790), .B(n4789), .Z(n4746) );
  XNOR U5334 ( .A(n4747), .B(n4746), .Z(n4749) );
  NAND U5335 ( .A(x[139]), .B(y[688]), .Z(n5706) );
  NANDN U5336 ( .A(n5706), .B(n4874), .Z(n4626) );
  NANDN U5337 ( .A(n4624), .B(n4623), .Z(n4625) );
  AND U5338 ( .A(n4626), .B(n4625), .Z(n4796) );
  AND U5339 ( .A(y[691]), .B(x[129]), .Z(n4628) );
  NAND U5340 ( .A(y[681]), .B(x[139]), .Z(n4627) );
  XNOR U5341 ( .A(n4628), .B(n4627), .Z(n4718) );
  NAND U5342 ( .A(x[147]), .B(y[673]), .Z(n4727) );
  XOR U5343 ( .A(o[52]), .B(n4727), .Z(n4719) );
  XNOR U5344 ( .A(n4718), .B(n4719), .Z(n4794) );
  AND U5345 ( .A(x[128]), .B(y[692]), .Z(n4777) );
  NAND U5346 ( .A(x[148]), .B(y[672]), .Z(n4778) );
  XNOR U5347 ( .A(n4777), .B(n4778), .Z(n4780) );
  ANDN U5348 ( .B(o[51]), .A(n4629), .Z(n4779) );
  XOR U5349 ( .A(n4780), .B(n4779), .Z(n4793) );
  XOR U5350 ( .A(n4794), .B(n4793), .Z(n4795) );
  XNOR U5351 ( .A(n4796), .B(n4795), .Z(n4748) );
  XOR U5352 ( .A(n4749), .B(n4748), .Z(n4708) );
  XOR U5353 ( .A(n4709), .B(n4708), .Z(n4800) );
  AND U5354 ( .A(x[134]), .B(y[686]), .Z(n4729) );
  NAND U5355 ( .A(n4729), .B(n4630), .Z(n4633) );
  NANDN U5356 ( .A(n4631), .B(n4772), .Z(n4632) );
  AND U5357 ( .A(n4633), .B(n4632), .Z(n4737) );
  AND U5358 ( .A(y[674]), .B(x[146]), .Z(n4639) );
  NAND U5359 ( .A(y[680]), .B(x[140]), .Z(n4638) );
  XNOR U5360 ( .A(n4639), .B(n4638), .Z(n4713) );
  NAND U5361 ( .A(x[145]), .B(y[675]), .Z(n4714) );
  XNOR U5362 ( .A(n4713), .B(n4714), .Z(n4734) );
  XNOR U5363 ( .A(n4735), .B(n4734), .Z(n4736) );
  XOR U5364 ( .A(n4737), .B(n4736), .Z(n4741) );
  AND U5365 ( .A(y[689]), .B(x[131]), .Z(n4641) );
  NAND U5366 ( .A(y[679]), .B(x[141]), .Z(n4640) );
  XNOR U5367 ( .A(n4641), .B(n4640), .Z(n4759) );
  XOR U5368 ( .A(n4759), .B(n4758), .Z(n4730) );
  AND U5369 ( .A(y[687]), .B(x[133]), .Z(n4643) );
  NAND U5370 ( .A(y[688]), .B(x[132]), .Z(n4642) );
  XNOR U5371 ( .A(n4643), .B(n4642), .Z(n4774) );
  AND U5372 ( .A(x[135]), .B(y[685]), .Z(n4773) );
  XNOR U5373 ( .A(n4774), .B(n4773), .Z(n4728) );
  XOR U5374 ( .A(n4729), .B(n4728), .Z(n4731) );
  XOR U5375 ( .A(n4730), .B(n4731), .Z(n4783) );
  AND U5376 ( .A(x[136]), .B(y[690]), .Z(n5851) );
  NAND U5377 ( .A(n5851), .B(n4644), .Z(n4648) );
  NANDN U5378 ( .A(n4646), .B(n4645), .Z(n4647) );
  AND U5379 ( .A(n4648), .B(n4647), .Z(n4782) );
  AND U5380 ( .A(x[145]), .B(y[681]), .Z(n5531) );
  AND U5381 ( .A(x[138]), .B(y[674]), .Z(n4649) );
  NAND U5382 ( .A(n5531), .B(n4649), .Z(n4653) );
  NANDN U5383 ( .A(n4651), .B(n4650), .Z(n4652) );
  NAND U5384 ( .A(n4653), .B(n4652), .Z(n4781) );
  XOR U5385 ( .A(n4782), .B(n4781), .Z(n4784) );
  XNOR U5386 ( .A(n4783), .B(n4784), .Z(n4740) );
  XOR U5387 ( .A(n4741), .B(n4740), .Z(n4743) );
  NANDN U5388 ( .A(n4655), .B(n4654), .Z(n4659) );
  NANDN U5389 ( .A(n4657), .B(n4656), .Z(n4658) );
  AND U5390 ( .A(n4659), .B(n4658), .Z(n4742) );
  XOR U5391 ( .A(n4743), .B(n4742), .Z(n4798) );
  NAND U5392 ( .A(n4661), .B(n4660), .Z(n4665) );
  NANDN U5393 ( .A(n4663), .B(n4662), .Z(n4664) );
  AND U5394 ( .A(n4665), .B(n4664), .Z(n4797) );
  XOR U5395 ( .A(n4798), .B(n4797), .Z(n4799) );
  XNOR U5396 ( .A(n4800), .B(n4799), .Z(n4804) );
  NANDN U5397 ( .A(n4667), .B(n4666), .Z(n4671) );
  NANDN U5398 ( .A(n4669), .B(n4668), .Z(n4670) );
  AND U5399 ( .A(n4671), .B(n4670), .Z(n4811) );
  NAND U5400 ( .A(n4673), .B(n4672), .Z(n4677) );
  NAND U5401 ( .A(n4675), .B(n4674), .Z(n4676) );
  NAND U5402 ( .A(n4677), .B(n4676), .Z(n4809) );
  NANDN U5403 ( .A(n4679), .B(n4678), .Z(n4683) );
  NAND U5404 ( .A(n4681), .B(n4680), .Z(n4682) );
  AND U5405 ( .A(n4683), .B(n4682), .Z(n4810) );
  XNOR U5406 ( .A(n4809), .B(n4810), .Z(n4812) );
  XOR U5407 ( .A(n4804), .B(n4803), .Z(n4805) );
  NAND U5408 ( .A(n4685), .B(n4684), .Z(n4689) );
  NANDN U5409 ( .A(n4687), .B(n4686), .Z(n4688) );
  AND U5410 ( .A(n4689), .B(n4688), .Z(n4819) );
  NANDN U5411 ( .A(n4691), .B(n4690), .Z(n4695) );
  NANDN U5412 ( .A(n4693), .B(n4692), .Z(n4694) );
  AND U5413 ( .A(n4695), .B(n4694), .Z(n4818) );
  XOR U5414 ( .A(n4819), .B(n4818), .Z(n4820) );
  XNOR U5415 ( .A(n4821), .B(n4820), .Z(n4817) );
  NAND U5416 ( .A(n4697), .B(n4696), .Z(n4701) );
  NAND U5417 ( .A(n4699), .B(n4698), .Z(n4700) );
  AND U5418 ( .A(n4701), .B(n4700), .Z(n4816) );
  XNOR U5419 ( .A(n4816), .B(n4815), .Z(n4705) );
  XNOR U5420 ( .A(n4817), .B(n4705), .Z(N117) );
  NAND U5421 ( .A(n4707), .B(n4706), .Z(n4711) );
  NAND U5422 ( .A(n4709), .B(n4708), .Z(n4710) );
  NAND U5423 ( .A(n4711), .B(n4710), .Z(n4831) );
  AND U5424 ( .A(x[146]), .B(y[680]), .Z(n5532) );
  NAND U5425 ( .A(n5532), .B(n4712), .Z(n4716) );
  NANDN U5426 ( .A(n4714), .B(n4713), .Z(n4715) );
  AND U5427 ( .A(n4716), .B(n4715), .Z(n4897) );
  AND U5428 ( .A(x[139]), .B(y[691]), .Z(n6233) );
  NAND U5429 ( .A(n6233), .B(n4717), .Z(n4721) );
  NANDN U5430 ( .A(n4719), .B(n4718), .Z(n4720) );
  NAND U5431 ( .A(n4721), .B(n4720), .Z(n4896) );
  XNOR U5432 ( .A(n4897), .B(n4896), .Z(n4899) );
  AND U5433 ( .A(x[143]), .B(y[683]), .Z(n5519) );
  NAND U5434 ( .A(n5519), .B(n4722), .Z(n4726) );
  NANDN U5435 ( .A(n4724), .B(n4723), .Z(n4725) );
  AND U5436 ( .A(n4726), .B(n4725), .Z(n4863) );
  AND U5437 ( .A(x[128]), .B(y[693]), .Z(n4880) );
  NAND U5438 ( .A(x[149]), .B(y[672]), .Z(n4881) );
  XNOR U5439 ( .A(n4880), .B(n4881), .Z(n4883) );
  ANDN U5440 ( .B(o[52]), .A(n4727), .Z(n4882) );
  XOR U5441 ( .A(n4883), .B(n4882), .Z(n4861) );
  AND U5442 ( .A(x[133]), .B(y[688]), .Z(n4865) );
  AND U5443 ( .A(x[144]), .B(y[677]), .Z(n4864) );
  XOR U5444 ( .A(n4865), .B(n4864), .Z(n4867) );
  NAND U5445 ( .A(x[143]), .B(y[678]), .Z(n4866) );
  XNOR U5446 ( .A(n4867), .B(n4866), .Z(n4860) );
  XOR U5447 ( .A(n4861), .B(n4860), .Z(n4862) );
  XNOR U5448 ( .A(n4863), .B(n4862), .Z(n4898) );
  XOR U5449 ( .A(n4899), .B(n4898), .Z(n4915) );
  NANDN U5450 ( .A(n4729), .B(n4728), .Z(n4733) );
  OR U5451 ( .A(n4731), .B(n4730), .Z(n4732) );
  NAND U5452 ( .A(n4733), .B(n4732), .Z(n4914) );
  XNOR U5453 ( .A(n4915), .B(n4914), .Z(n4916) );
  NANDN U5454 ( .A(n4735), .B(n4734), .Z(n4739) );
  NANDN U5455 ( .A(n4737), .B(n4736), .Z(n4738) );
  NAND U5456 ( .A(n4739), .B(n4738), .Z(n4917) );
  XOR U5457 ( .A(n4916), .B(n4917), .Z(n4829) );
  NAND U5458 ( .A(n4741), .B(n4740), .Z(n4745) );
  NAND U5459 ( .A(n4743), .B(n4742), .Z(n4744) );
  AND U5460 ( .A(n4745), .B(n4744), .Z(n4830) );
  XOR U5461 ( .A(n4829), .B(n4830), .Z(n4832) );
  XNOR U5462 ( .A(n4831), .B(n4832), .Z(n4825) );
  NANDN U5463 ( .A(n4747), .B(n4746), .Z(n4751) );
  NAND U5464 ( .A(n4749), .B(n4748), .Z(n4750) );
  AND U5465 ( .A(n4751), .B(n4750), .Z(n4923) );
  NAND U5466 ( .A(n5525), .B(n4752), .Z(n4756) );
  NANDN U5467 ( .A(n4754), .B(n4753), .Z(n4755) );
  AND U5468 ( .A(n4756), .B(n4755), .Z(n4836) );
  AND U5469 ( .A(x[131]), .B(y[679]), .Z(n4757) );
  NAND U5470 ( .A(n6086), .B(n4757), .Z(n4761) );
  NAND U5471 ( .A(n4759), .B(n4758), .Z(n4760) );
  AND U5472 ( .A(n4761), .B(n4760), .Z(n4911) );
  AND U5473 ( .A(y[674]), .B(x[147]), .Z(n4763) );
  NAND U5474 ( .A(y[682]), .B(x[139]), .Z(n4762) );
  XNOR U5475 ( .A(n4763), .B(n4762), .Z(n4852) );
  NAND U5476 ( .A(x[148]), .B(y[673]), .Z(n4879) );
  XOR U5477 ( .A(o[53]), .B(n4879), .Z(n4853) );
  XNOR U5478 ( .A(n4852), .B(n4853), .Z(n4908) );
  AND U5479 ( .A(y[675]), .B(x[146]), .Z(n4765) );
  NAND U5480 ( .A(y[683]), .B(x[138]), .Z(n4764) );
  XNOR U5481 ( .A(n4765), .B(n4764), .Z(n4887) );
  NAND U5482 ( .A(x[129]), .B(y[692]), .Z(n4888) );
  XOR U5483 ( .A(n4887), .B(n4888), .Z(n4909) );
  XNOR U5484 ( .A(n4908), .B(n4909), .Z(n4910) );
  XNOR U5485 ( .A(n4911), .B(n4910), .Z(n4835) );
  XNOR U5486 ( .A(n4836), .B(n4835), .Z(n4838) );
  AND U5487 ( .A(x[135]), .B(y[686]), .Z(n5089) );
  AND U5488 ( .A(y[679]), .B(x[142]), .Z(n4767) );
  NAND U5489 ( .A(y[687]), .B(x[134]), .Z(n4766) );
  XNOR U5490 ( .A(n4767), .B(n4766), .Z(n4891) );
  XOR U5491 ( .A(n5089), .B(n4891), .Z(n4842) );
  AND U5492 ( .A(x[137]), .B(y[684]), .Z(n4840) );
  NAND U5493 ( .A(x[136]), .B(y[685]), .Z(n4839) );
  XNOR U5494 ( .A(n4840), .B(n4839), .Z(n4841) );
  XOR U5495 ( .A(n4842), .B(n4841), .Z(n4859) );
  AND U5496 ( .A(y[676]), .B(x[145]), .Z(n4769) );
  NAND U5497 ( .A(y[681]), .B(x[140]), .Z(n4768) );
  XNOR U5498 ( .A(n4769), .B(n4768), .Z(n4845) );
  NAND U5499 ( .A(x[130]), .B(y[691]), .Z(n4846) );
  XNOR U5500 ( .A(n4845), .B(n4846), .Z(n4857) );
  AND U5501 ( .A(y[690]), .B(x[131]), .Z(n4771) );
  NAND U5502 ( .A(y[680]), .B(x[141]), .Z(n4770) );
  XNOR U5503 ( .A(n4771), .B(n4770), .Z(n4875) );
  NAND U5504 ( .A(x[132]), .B(y[689]), .Z(n4876) );
  XNOR U5505 ( .A(n4875), .B(n4876), .Z(n4856) );
  XOR U5506 ( .A(n4857), .B(n4856), .Z(n4858) );
  XOR U5507 ( .A(n4859), .B(n4858), .Z(n4905) );
  NAND U5508 ( .A(n4865), .B(n4772), .Z(n4776) );
  NAND U5509 ( .A(n4774), .B(n4773), .Z(n4775) );
  AND U5510 ( .A(n4776), .B(n4775), .Z(n4903) );
  XNOR U5511 ( .A(n4903), .B(n4902), .Z(n4904) );
  XOR U5512 ( .A(n4905), .B(n4904), .Z(n4837) );
  XOR U5513 ( .A(n4838), .B(n4837), .Z(n4921) );
  NANDN U5514 ( .A(n4782), .B(n4781), .Z(n4786) );
  OR U5515 ( .A(n4784), .B(n4783), .Z(n4785) );
  NAND U5516 ( .A(n4786), .B(n4785), .Z(n4926) );
  NANDN U5517 ( .A(n4788), .B(n4787), .Z(n4792) );
  NANDN U5518 ( .A(n4790), .B(n4789), .Z(n4791) );
  NAND U5519 ( .A(n4792), .B(n4791), .Z(n4925) );
  XOR U5520 ( .A(n4925), .B(n4924), .Z(n4927) );
  XOR U5521 ( .A(n4926), .B(n4927), .Z(n4920) );
  XOR U5522 ( .A(n4921), .B(n4920), .Z(n4922) );
  XOR U5523 ( .A(n4923), .B(n4922), .Z(n4824) );
  NAND U5524 ( .A(n4798), .B(n4797), .Z(n4802) );
  NANDN U5525 ( .A(n4800), .B(n4799), .Z(n4801) );
  NAND U5526 ( .A(n4802), .B(n4801), .Z(n4823) );
  XNOR U5527 ( .A(n4824), .B(n4823), .Z(n4826) );
  XOR U5528 ( .A(n4825), .B(n4826), .Z(n4935) );
  NAND U5529 ( .A(n4804), .B(n4803), .Z(n4808) );
  NANDN U5530 ( .A(n4806), .B(n4805), .Z(n4807) );
  AND U5531 ( .A(n4808), .B(n4807), .Z(n4933) );
  NAND U5532 ( .A(n4810), .B(n4809), .Z(n4814) );
  NANDN U5533 ( .A(n4812), .B(n4811), .Z(n4813) );
  NAND U5534 ( .A(n4814), .B(n4813), .Z(n4934) );
  XNOR U5535 ( .A(n4935), .B(n4936), .Z(n4932) );
  XOR U5536 ( .A(n4930), .B(n4931), .Z(n4822) );
  XNOR U5537 ( .A(n4932), .B(n4822), .Z(N118) );
  NAND U5538 ( .A(n4824), .B(n4823), .Z(n4828) );
  NANDN U5539 ( .A(n4826), .B(n4825), .Z(n4827) );
  AND U5540 ( .A(n4828), .B(n4827), .Z(n4943) );
  NAND U5541 ( .A(n4830), .B(n4829), .Z(n4834) );
  NAND U5542 ( .A(n4832), .B(n4831), .Z(n4833) );
  NAND U5543 ( .A(n4834), .B(n4833), .Z(n4940) );
  NANDN U5544 ( .A(n4840), .B(n4839), .Z(n4844) );
  NANDN U5545 ( .A(n4842), .B(n4841), .Z(n4843) );
  AND U5546 ( .A(n4844), .B(n4843), .Z(n4978) );
  NAND U5547 ( .A(n5531), .B(n5030), .Z(n4848) );
  NANDN U5548 ( .A(n4846), .B(n4845), .Z(n4847) );
  NAND U5549 ( .A(n4848), .B(n4847), .Z(n5007) );
  AND U5550 ( .A(x[133]), .B(y[689]), .Z(n5051) );
  NAND U5551 ( .A(x[145]), .B(y[677]), .Z(n5052) );
  XNOR U5552 ( .A(n5051), .B(n5052), .Z(n5053) );
  NAND U5553 ( .A(x[144]), .B(y[678]), .Z(n5054) );
  XNOR U5554 ( .A(n5053), .B(n5054), .Z(n5006) );
  AND U5555 ( .A(y[676]), .B(x[146]), .Z(n4850) );
  NAND U5556 ( .A(y[682]), .B(x[140]), .Z(n4849) );
  XNOR U5557 ( .A(n4850), .B(n4849), .Z(n5031) );
  NAND U5558 ( .A(x[132]), .B(y[690]), .Z(n5032) );
  XNOR U5559 ( .A(n5031), .B(n5032), .Z(n5005) );
  XOR U5560 ( .A(n5006), .B(n5005), .Z(n5008) );
  XNOR U5561 ( .A(n5007), .B(n5008), .Z(n4975) );
  NAND U5562 ( .A(x[147]), .B(y[682]), .Z(n6000) );
  NANDN U5563 ( .A(n6000), .B(n4851), .Z(n4855) );
  NANDN U5564 ( .A(n4853), .B(n4852), .Z(n4854) );
  AND U5565 ( .A(n4855), .B(n4854), .Z(n4976) );
  XOR U5566 ( .A(n4975), .B(n4976), .Z(n4977) );
  XOR U5567 ( .A(n4978), .B(n4977), .Z(n4958) );
  XNOR U5568 ( .A(n4964), .B(n4963), .Z(n4966) );
  NAND U5569 ( .A(n4865), .B(n4864), .Z(n4869) );
  ANDN U5570 ( .B(n4867), .A(n4866), .Z(n4868) );
  ANDN U5571 ( .B(n4869), .A(n4868), .Z(n5027) );
  AND U5572 ( .A(y[674]), .B(x[148]), .Z(n4871) );
  NAND U5573 ( .A(y[681]), .B(x[141]), .Z(n4870) );
  XNOR U5574 ( .A(n4871), .B(n4870), .Z(n5047) );
  NAND U5575 ( .A(x[130]), .B(y[692]), .Z(n5048) );
  XNOR U5576 ( .A(n5047), .B(n5048), .Z(n5025) );
  AND U5577 ( .A(y[688]), .B(x[134]), .Z(n4873) );
  NAND U5578 ( .A(y[679]), .B(x[143]), .Z(n4872) );
  XNOR U5579 ( .A(n4873), .B(n4872), .Z(n5059) );
  XOR U5580 ( .A(n5025), .B(n5024), .Z(n5026) );
  XNOR U5581 ( .A(n5027), .B(n5026), .Z(n4970) );
  AND U5582 ( .A(x[141]), .B(y[690]), .Z(n6230) );
  NAND U5583 ( .A(n4874), .B(n6230), .Z(n4878) );
  NANDN U5584 ( .A(n4876), .B(n4875), .Z(n4877) );
  AND U5585 ( .A(n4878), .B(n4877), .Z(n4996) );
  AND U5586 ( .A(x[129]), .B(y[693]), .Z(n5019) );
  XOR U5587 ( .A(n5020), .B(n5019), .Z(n5018) );
  ANDN U5588 ( .B(o[53]), .A(n4879), .Z(n5017) );
  XOR U5589 ( .A(n5018), .B(n5017), .Z(n4994) );
  AND U5590 ( .A(x[142]), .B(y[680]), .Z(n5011) );
  NAND U5591 ( .A(x[131]), .B(y[691]), .Z(n5012) );
  XNOR U5592 ( .A(n5011), .B(n5012), .Z(n5013) );
  NAND U5593 ( .A(x[147]), .B(y[675]), .Z(n5014) );
  XNOR U5594 ( .A(n5013), .B(n5014), .Z(n4993) );
  XOR U5595 ( .A(n4994), .B(n4993), .Z(n4995) );
  XNOR U5596 ( .A(n4996), .B(n4995), .Z(n4969) );
  XOR U5597 ( .A(n4970), .B(n4969), .Z(n4972) );
  NANDN U5598 ( .A(n4881), .B(n4880), .Z(n4885) );
  NAND U5599 ( .A(n4883), .B(n4882), .Z(n4884) );
  AND U5600 ( .A(n4885), .B(n4884), .Z(n4988) );
  NAND U5601 ( .A(x[146]), .B(y[683]), .Z(n6002) );
  NANDN U5602 ( .A(n6002), .B(n4886), .Z(n4890) );
  NANDN U5603 ( .A(n4888), .B(n4887), .Z(n4889) );
  NAND U5604 ( .A(n4890), .B(n4889), .Z(n4987) );
  XNOR U5605 ( .A(n4988), .B(n4987), .Z(n4990) );
  AND U5606 ( .A(x[142]), .B(y[687]), .Z(n6036) );
  NAND U5607 ( .A(n6036), .B(n5058), .Z(n4893) );
  NAND U5608 ( .A(n5089), .B(n4891), .Z(n4892) );
  AND U5609 ( .A(n4893), .B(n4892), .Z(n5002) );
  AND U5610 ( .A(x[128]), .B(y[694]), .Z(n5035) );
  NAND U5611 ( .A(x[150]), .B(y[672]), .Z(n5036) );
  XNOR U5612 ( .A(n5035), .B(n5036), .Z(n5038) );
  NAND U5613 ( .A(x[149]), .B(y[673]), .Z(n5057) );
  XNOR U5614 ( .A(o[54]), .B(n5057), .Z(n5037) );
  XOR U5615 ( .A(n5038), .B(n5037), .Z(n5000) );
  NAND U5616 ( .A(y[687]), .B(x[135]), .Z(n4894) );
  XNOR U5617 ( .A(n4895), .B(n4894), .Z(n5041) );
  XOR U5618 ( .A(n5000), .B(n4999), .Z(n5001) );
  XNOR U5619 ( .A(n5002), .B(n5001), .Z(n4989) );
  XOR U5620 ( .A(n4990), .B(n4989), .Z(n4971) );
  XOR U5621 ( .A(n4972), .B(n4971), .Z(n4965) );
  XOR U5622 ( .A(n4966), .B(n4965), .Z(n4957) );
  XOR U5623 ( .A(n4958), .B(n4957), .Z(n4959) );
  XOR U5624 ( .A(n4960), .B(n4959), .Z(n5065) );
  NANDN U5625 ( .A(n4897), .B(n4896), .Z(n4901) );
  NAND U5626 ( .A(n4899), .B(n4898), .Z(n4900) );
  AND U5627 ( .A(n4901), .B(n4900), .Z(n4983) );
  NANDN U5628 ( .A(n4903), .B(n4902), .Z(n4907) );
  NAND U5629 ( .A(n4905), .B(n4904), .Z(n4906) );
  AND U5630 ( .A(n4907), .B(n4906), .Z(n4982) );
  NANDN U5631 ( .A(n4909), .B(n4908), .Z(n4913) );
  NANDN U5632 ( .A(n4911), .B(n4910), .Z(n4912) );
  NAND U5633 ( .A(n4913), .B(n4912), .Z(n4981) );
  XOR U5634 ( .A(n4982), .B(n4981), .Z(n4984) );
  XOR U5635 ( .A(n4983), .B(n4984), .Z(n5064) );
  NANDN U5636 ( .A(n4915), .B(n4914), .Z(n4919) );
  NANDN U5637 ( .A(n4917), .B(n4916), .Z(n4918) );
  NAND U5638 ( .A(n4919), .B(n4918), .Z(n5063) );
  XOR U5639 ( .A(n5064), .B(n5063), .Z(n5066) );
  XOR U5640 ( .A(n5065), .B(n5066), .Z(n4955) );
  NAND U5641 ( .A(n4925), .B(n4924), .Z(n4929) );
  NAND U5642 ( .A(n4927), .B(n4926), .Z(n4928) );
  NAND U5643 ( .A(n4929), .B(n4928), .Z(n4953) );
  XNOR U5644 ( .A(n4954), .B(n4953), .Z(n4956) );
  XOR U5645 ( .A(n4955), .B(n4956), .Z(n4941) );
  XOR U5646 ( .A(n4940), .B(n4941), .Z(n4942) );
  XNOR U5647 ( .A(n4943), .B(n4942), .Z(n4949) );
  NANDN U5648 ( .A(n4934), .B(n4933), .Z(n4938) );
  NAND U5649 ( .A(n4936), .B(n4935), .Z(n4937) );
  NAND U5650 ( .A(n4938), .B(n4937), .Z(n4947) );
  IV U5651 ( .A(n4947), .Z(n4946) );
  XOR U5652 ( .A(n4948), .B(n4946), .Z(n4939) );
  XNOR U5653 ( .A(n4949), .B(n4939), .Z(N119) );
  NAND U5654 ( .A(n4941), .B(n4940), .Z(n4945) );
  NAND U5655 ( .A(n4943), .B(n4942), .Z(n4944) );
  NAND U5656 ( .A(n4945), .B(n4944), .Z(n5206) );
  OR U5657 ( .A(n4948), .B(n4946), .Z(n4952) );
  ANDN U5658 ( .B(n4948), .A(n4947), .Z(n4950) );
  OR U5659 ( .A(n4950), .B(n4949), .Z(n4951) );
  AND U5660 ( .A(n4952), .B(n4951), .Z(n5207) );
  NAND U5661 ( .A(n4958), .B(n4957), .Z(n4962) );
  NANDN U5662 ( .A(n4960), .B(n4959), .Z(n4961) );
  AND U5663 ( .A(n4962), .B(n4961), .Z(n5071) );
  NANDN U5664 ( .A(n4964), .B(n4963), .Z(n4968) );
  NAND U5665 ( .A(n4966), .B(n4965), .Z(n4967) );
  AND U5666 ( .A(n4968), .B(n4967), .Z(n5191) );
  NAND U5667 ( .A(n4970), .B(n4969), .Z(n4974) );
  NAND U5668 ( .A(n4972), .B(n4971), .Z(n4973) );
  AND U5669 ( .A(n4974), .B(n4973), .Z(n5189) );
  NAND U5670 ( .A(n4976), .B(n4975), .Z(n4980) );
  NANDN U5671 ( .A(n4978), .B(n4977), .Z(n4979) );
  AND U5672 ( .A(n4980), .B(n4979), .Z(n5188) );
  XNOR U5673 ( .A(n5189), .B(n5188), .Z(n5190) );
  XNOR U5674 ( .A(n5191), .B(n5190), .Z(n5070) );
  NANDN U5675 ( .A(n4982), .B(n4981), .Z(n4986) );
  OR U5676 ( .A(n4984), .B(n4983), .Z(n4985) );
  AND U5677 ( .A(n4986), .B(n4985), .Z(n5185) );
  NANDN U5678 ( .A(n4988), .B(n4987), .Z(n4992) );
  NAND U5679 ( .A(n4990), .B(n4989), .Z(n4991) );
  AND U5680 ( .A(n4992), .B(n4991), .Z(n5179) );
  NAND U5681 ( .A(n4994), .B(n4993), .Z(n4998) );
  NANDN U5682 ( .A(n4996), .B(n4995), .Z(n4997) );
  AND U5683 ( .A(n4998), .B(n4997), .Z(n5177) );
  NAND U5684 ( .A(n5000), .B(n4999), .Z(n5004) );
  NANDN U5685 ( .A(n5002), .B(n5001), .Z(n5003) );
  NAND U5686 ( .A(n5004), .B(n5003), .Z(n5176) );
  XNOR U5687 ( .A(n5177), .B(n5176), .Z(n5178) );
  XNOR U5688 ( .A(n5179), .B(n5178), .Z(n5197) );
  NAND U5689 ( .A(n5006), .B(n5005), .Z(n5010) );
  NAND U5690 ( .A(n5008), .B(n5007), .Z(n5009) );
  AND U5691 ( .A(n5010), .B(n5009), .Z(n5195) );
  NANDN U5692 ( .A(n5012), .B(n5011), .Z(n5016) );
  NANDN U5693 ( .A(n5014), .B(n5013), .Z(n5015) );
  AND U5694 ( .A(n5016), .B(n5015), .Z(n5123) );
  AND U5695 ( .A(n5018), .B(n5017), .Z(n5022) );
  NAND U5696 ( .A(n5020), .B(n5019), .Z(n5021) );
  NANDN U5697 ( .A(n5022), .B(n5021), .Z(n5122) );
  XNOR U5698 ( .A(n5123), .B(n5122), .Z(n5125) );
  NAND U5699 ( .A(y[688]), .B(x[135]), .Z(n5023) );
  XOR U5700 ( .A(n5263), .B(n5023), .Z(n5091) );
  XNOR U5701 ( .A(n5090), .B(n5091), .Z(n5128) );
  NAND U5702 ( .A(x[138]), .B(y[685]), .Z(n5129) );
  XNOR U5703 ( .A(n5128), .B(n5129), .Z(n5131) );
  AND U5704 ( .A(x[134]), .B(y[689]), .Z(n5081) );
  NAND U5705 ( .A(x[143]), .B(y[680]), .Z(n5082) );
  XNOR U5706 ( .A(n5081), .B(n5082), .Z(n5083) );
  NAND U5707 ( .A(x[139]), .B(y[684]), .Z(n5084) );
  XNOR U5708 ( .A(n5083), .B(n5084), .Z(n5130) );
  XOR U5709 ( .A(n5131), .B(n5130), .Z(n5124) );
  XOR U5710 ( .A(n5125), .B(n5124), .Z(n5194) );
  XNOR U5711 ( .A(n5195), .B(n5194), .Z(n5196) );
  XOR U5712 ( .A(n5197), .B(n5196), .Z(n5183) );
  NAND U5713 ( .A(n5025), .B(n5024), .Z(n5029) );
  NANDN U5714 ( .A(n5027), .B(n5026), .Z(n5028) );
  AND U5715 ( .A(n5029), .B(n5028), .Z(n5117) );
  AND U5716 ( .A(x[146]), .B(y[682]), .Z(n5873) );
  NAND U5717 ( .A(n5873), .B(n5030), .Z(n5034) );
  NANDN U5718 ( .A(n5032), .B(n5031), .Z(n5033) );
  AND U5719 ( .A(n5034), .B(n5033), .Z(n5165) );
  NANDN U5720 ( .A(n5036), .B(n5035), .Z(n5040) );
  NAND U5721 ( .A(n5038), .B(n5037), .Z(n5039) );
  NAND U5722 ( .A(n5040), .B(n5039), .Z(n5164) );
  XNOR U5723 ( .A(n5165), .B(n5164), .Z(n5167) );
  NAND U5724 ( .A(n5089), .B(n5090), .Z(n5044) );
  NANDN U5725 ( .A(n5042), .B(n5041), .Z(n5043) );
  AND U5726 ( .A(n5044), .B(n5043), .Z(n5161) );
  AND U5727 ( .A(x[128]), .B(y[695]), .Z(n5100) );
  NAND U5728 ( .A(x[151]), .B(y[672]), .Z(n5101) );
  XNOR U5729 ( .A(n5100), .B(n5101), .Z(n5103) );
  NAND U5730 ( .A(x[150]), .B(y[673]), .Z(n5080) );
  XNOR U5731 ( .A(o[55]), .B(n5080), .Z(n5102) );
  XOR U5732 ( .A(n5103), .B(n5102), .Z(n5159) );
  AND U5733 ( .A(y[675]), .B(x[148]), .Z(n5743) );
  NAND U5734 ( .A(y[679]), .B(x[144]), .Z(n5045) );
  XNOR U5735 ( .A(n5743), .B(n5045), .Z(n5076) );
  NAND U5736 ( .A(x[147]), .B(y[676]), .Z(n5077) );
  XNOR U5737 ( .A(n5076), .B(n5077), .Z(n5158) );
  XOR U5738 ( .A(n5159), .B(n5158), .Z(n5160) );
  XNOR U5739 ( .A(n5161), .B(n5160), .Z(n5166) );
  XOR U5740 ( .A(n5167), .B(n5166), .Z(n5116) );
  XNOR U5741 ( .A(n5117), .B(n5116), .Z(n5119) );
  NAND U5742 ( .A(x[148]), .B(y[681]), .Z(n6044) );
  NANDN U5743 ( .A(n6044), .B(n5046), .Z(n5050) );
  NANDN U5744 ( .A(n5048), .B(n5047), .Z(n5049) );
  AND U5745 ( .A(n5050), .B(n5049), .Z(n5111) );
  NANDN U5746 ( .A(n5052), .B(n5051), .Z(n5056) );
  NANDN U5747 ( .A(n5054), .B(n5053), .Z(n5055) );
  AND U5748 ( .A(n5056), .B(n5055), .Z(n5173) );
  AND U5749 ( .A(x[141]), .B(y[682]), .Z(n5146) );
  NAND U5750 ( .A(x[130]), .B(y[693]), .Z(n5147) );
  XNOR U5751 ( .A(n5146), .B(n5147), .Z(n5148) );
  NAND U5752 ( .A(x[149]), .B(y[674]), .Z(n5149) );
  XNOR U5753 ( .A(n5148), .B(n5149), .Z(n5171) );
  ANDN U5754 ( .B(o[54]), .A(n5057), .Z(n5097) );
  AND U5755 ( .A(x[140]), .B(y[683]), .Z(n5094) );
  NAND U5756 ( .A(x[129]), .B(y[694]), .Z(n5095) );
  XNOR U5757 ( .A(n5094), .B(n5095), .Z(n5096) );
  XOR U5758 ( .A(n5097), .B(n5096), .Z(n5170) );
  XOR U5759 ( .A(n5171), .B(n5170), .Z(n5172) );
  XNOR U5760 ( .A(n5173), .B(n5172), .Z(n5110) );
  XNOR U5761 ( .A(n5111), .B(n5110), .Z(n5113) );
  AND U5762 ( .A(x[143]), .B(y[688]), .Z(n6196) );
  NAND U5763 ( .A(n6196), .B(n5058), .Z(n5062) );
  NANDN U5764 ( .A(n5060), .B(n5059), .Z(n5061) );
  AND U5765 ( .A(n5062), .B(n5061), .Z(n5155) );
  AND U5766 ( .A(x[142]), .B(y[681]), .Z(n5140) );
  NAND U5767 ( .A(x[131]), .B(y[692]), .Z(n5141) );
  XNOR U5768 ( .A(n5140), .B(n5141), .Z(n5142) );
  NAND U5769 ( .A(x[132]), .B(y[691]), .Z(n5143) );
  XNOR U5770 ( .A(n5142), .B(n5143), .Z(n5153) );
  AND U5771 ( .A(x[133]), .B(y[690]), .Z(n5134) );
  NAND U5772 ( .A(x[146]), .B(y[677]), .Z(n5135) );
  XNOR U5773 ( .A(n5134), .B(n5135), .Z(n5136) );
  NAND U5774 ( .A(x[145]), .B(y[678]), .Z(n5137) );
  XNOR U5775 ( .A(n5136), .B(n5137), .Z(n5152) );
  XOR U5776 ( .A(n5153), .B(n5152), .Z(n5154) );
  XNOR U5777 ( .A(n5155), .B(n5154), .Z(n5112) );
  XOR U5778 ( .A(n5113), .B(n5112), .Z(n5118) );
  XOR U5779 ( .A(n5119), .B(n5118), .Z(n5182) );
  XOR U5780 ( .A(n5183), .B(n5182), .Z(n5184) );
  XNOR U5781 ( .A(n5185), .B(n5184), .Z(n5072) );
  XOR U5782 ( .A(n5073), .B(n5072), .Z(n5201) );
  NANDN U5783 ( .A(n5064), .B(n5063), .Z(n5068) );
  NANDN U5784 ( .A(n5066), .B(n5065), .Z(n5067) );
  NAND U5785 ( .A(n5068), .B(n5067), .Z(n5200) );
  XOR U5786 ( .A(n5201), .B(n5200), .Z(n5203) );
  XNOR U5787 ( .A(n5202), .B(n5203), .Z(n5208) );
  XNOR U5788 ( .A(n5207), .B(n5208), .Z(n5069) );
  XNOR U5789 ( .A(n5206), .B(n5069), .Z(N120) );
  NANDN U5790 ( .A(n5071), .B(n5070), .Z(n5075) );
  NAND U5791 ( .A(n5073), .B(n5072), .Z(n5074) );
  AND U5792 ( .A(n5075), .B(n5074), .Z(n5343) );
  AND U5793 ( .A(x[148]), .B(y[679]), .Z(n5629) );
  AND U5794 ( .A(x[144]), .B(y[675]), .Z(n5234) );
  NAND U5795 ( .A(n5629), .B(n5234), .Z(n5079) );
  NANDN U5796 ( .A(n5077), .B(n5076), .Z(n5078) );
  AND U5797 ( .A(n5079), .B(n5078), .Z(n5248) );
  AND U5798 ( .A(x[150]), .B(y[674]), .Z(n5273) );
  XOR U5799 ( .A(n5274), .B(n5273), .Z(n5276) );
  AND U5800 ( .A(x[130]), .B(y[694]), .Z(n5275) );
  XOR U5801 ( .A(n5276), .B(n5275), .Z(n5246) );
  AND U5802 ( .A(x[129]), .B(y[695]), .Z(n5281) );
  XOR U5803 ( .A(n5282), .B(n5281), .Z(n5280) );
  ANDN U5804 ( .B(o[55]), .A(n5080), .Z(n5279) );
  XOR U5805 ( .A(n5280), .B(n5279), .Z(n5245) );
  XOR U5806 ( .A(n5246), .B(n5245), .Z(n5247) );
  XNOR U5807 ( .A(n5248), .B(n5247), .Z(n5311) );
  NANDN U5808 ( .A(n5082), .B(n5081), .Z(n5086) );
  NANDN U5809 ( .A(n5084), .B(n5083), .Z(n5085) );
  AND U5810 ( .A(n5086), .B(n5085), .Z(n5254) );
  AND U5811 ( .A(y[675]), .B(x[149]), .Z(n5088) );
  NAND U5812 ( .A(y[680]), .B(x[144]), .Z(n5087) );
  XNOR U5813 ( .A(n5088), .B(n5087), .Z(n5236) );
  AND U5814 ( .A(x[133]), .B(y[691]), .Z(n5235) );
  XOR U5815 ( .A(n5236), .B(n5235), .Z(n5252) );
  AND U5816 ( .A(x[134]), .B(y[690]), .Z(n5616) );
  AND U5817 ( .A(x[148]), .B(y[676]), .Z(n5458) );
  XOR U5818 ( .A(n5616), .B(n5458), .Z(n5242) );
  AND U5819 ( .A(x[147]), .B(y[677]), .Z(n5241) );
  XOR U5820 ( .A(n5242), .B(n5241), .Z(n5251) );
  XOR U5821 ( .A(n5252), .B(n5251), .Z(n5253) );
  XNOR U5822 ( .A(n5254), .B(n5253), .Z(n5225) );
  NAND U5823 ( .A(n5384), .B(n5089), .Z(n5093) );
  NANDN U5824 ( .A(n5091), .B(n5090), .Z(n5092) );
  AND U5825 ( .A(n5093), .B(n5092), .Z(n5223) );
  NANDN U5826 ( .A(n5095), .B(n5094), .Z(n5099) );
  NAND U5827 ( .A(n5097), .B(n5096), .Z(n5098) );
  NAND U5828 ( .A(n5099), .B(n5098), .Z(n5222) );
  XNOR U5829 ( .A(n5223), .B(n5222), .Z(n5224) );
  XOR U5830 ( .A(n5225), .B(n5224), .Z(n5310) );
  XOR U5831 ( .A(n5311), .B(n5310), .Z(n5313) );
  NANDN U5832 ( .A(n5101), .B(n5100), .Z(n5105) );
  NAND U5833 ( .A(n5103), .B(n5102), .Z(n5104) );
  AND U5834 ( .A(n5105), .B(n5104), .Z(n5293) );
  AND U5835 ( .A(x[131]), .B(y[693]), .Z(n5298) );
  XOR U5836 ( .A(n5299), .B(n5298), .Z(n5301) );
  NAND U5837 ( .A(x[132]), .B(y[692]), .Z(n5300) );
  XNOR U5838 ( .A(n5301), .B(n5300), .Z(n5292) );
  AND U5839 ( .A(y[687]), .B(x[137]), .Z(n5107) );
  NAND U5840 ( .A(y[686]), .B(x[138]), .Z(n5106) );
  XNOR U5841 ( .A(n5107), .B(n5106), .Z(n5265) );
  AND U5842 ( .A(y[682]), .B(x[142]), .Z(n5109) );
  NAND U5843 ( .A(y[688]), .B(x[136]), .Z(n5108) );
  XNOR U5844 ( .A(n5109), .B(n5108), .Z(n5269) );
  NAND U5845 ( .A(x[139]), .B(y[685]), .Z(n5270) );
  XNOR U5846 ( .A(n5269), .B(n5270), .Z(n5264) );
  XOR U5847 ( .A(n5265), .B(n5264), .Z(n5294) );
  XOR U5848 ( .A(n5295), .B(n5294), .Z(n5312) );
  XOR U5849 ( .A(n5313), .B(n5312), .Z(n5323) );
  NANDN U5850 ( .A(n5111), .B(n5110), .Z(n5115) );
  NAND U5851 ( .A(n5113), .B(n5112), .Z(n5114) );
  AND U5852 ( .A(n5115), .B(n5114), .Z(n5322) );
  XNOR U5853 ( .A(n5323), .B(n5322), .Z(n5324) );
  NANDN U5854 ( .A(n5117), .B(n5116), .Z(n5121) );
  NAND U5855 ( .A(n5119), .B(n5118), .Z(n5120) );
  NAND U5856 ( .A(n5121), .B(n5120), .Z(n5325) );
  XNOR U5857 ( .A(n5324), .B(n5325), .Z(n5331) );
  NANDN U5858 ( .A(n5123), .B(n5122), .Z(n5127) );
  NAND U5859 ( .A(n5125), .B(n5124), .Z(n5126) );
  AND U5860 ( .A(n5127), .B(n5126), .Z(n5319) );
  NANDN U5861 ( .A(n5129), .B(n5128), .Z(n5133) );
  NAND U5862 ( .A(n5131), .B(n5130), .Z(n5132) );
  AND U5863 ( .A(n5133), .B(n5132), .Z(n5317) );
  NANDN U5864 ( .A(n5135), .B(n5134), .Z(n5139) );
  NANDN U5865 ( .A(n5137), .B(n5136), .Z(n5138) );
  AND U5866 ( .A(n5139), .B(n5138), .Z(n5231) );
  AND U5867 ( .A(x[128]), .B(y[696]), .Z(n5305) );
  AND U5868 ( .A(x[152]), .B(y[672]), .Z(n5304) );
  XOR U5869 ( .A(n5305), .B(n5304), .Z(n5307) );
  AND U5870 ( .A(x[151]), .B(y[673]), .Z(n5291) );
  XOR U5871 ( .A(n5291), .B(o[56]), .Z(n5306) );
  XOR U5872 ( .A(n5307), .B(n5306), .Z(n5229) );
  AND U5873 ( .A(x[135]), .B(y[689]), .Z(n5286) );
  AND U5874 ( .A(x[146]), .B(y[678]), .Z(n5285) );
  XOR U5875 ( .A(n5286), .B(n5285), .Z(n5288) );
  AND U5876 ( .A(x[145]), .B(y[679]), .Z(n5287) );
  XOR U5877 ( .A(n5288), .B(n5287), .Z(n5228) );
  XOR U5878 ( .A(n5229), .B(n5228), .Z(n5230) );
  XNOR U5879 ( .A(n5231), .B(n5230), .Z(n5219) );
  NANDN U5880 ( .A(n5141), .B(n5140), .Z(n5145) );
  NANDN U5881 ( .A(n5143), .B(n5142), .Z(n5144) );
  AND U5882 ( .A(n5145), .B(n5144), .Z(n5217) );
  NANDN U5883 ( .A(n5147), .B(n5146), .Z(n5151) );
  NANDN U5884 ( .A(n5149), .B(n5148), .Z(n5150) );
  NAND U5885 ( .A(n5151), .B(n5150), .Z(n5216) );
  XNOR U5886 ( .A(n5217), .B(n5216), .Z(n5218) );
  XOR U5887 ( .A(n5219), .B(n5218), .Z(n5316) );
  XNOR U5888 ( .A(n5317), .B(n5316), .Z(n5318) );
  XOR U5889 ( .A(n5319), .B(n5318), .Z(n5212) );
  NAND U5890 ( .A(n5153), .B(n5152), .Z(n5157) );
  NANDN U5891 ( .A(n5155), .B(n5154), .Z(n5156) );
  AND U5892 ( .A(n5157), .B(n5156), .Z(n5258) );
  NAND U5893 ( .A(n5159), .B(n5158), .Z(n5163) );
  NANDN U5894 ( .A(n5161), .B(n5160), .Z(n5162) );
  AND U5895 ( .A(n5163), .B(n5162), .Z(n5257) );
  XOR U5896 ( .A(n5258), .B(n5257), .Z(n5260) );
  NANDN U5897 ( .A(n5165), .B(n5164), .Z(n5169) );
  NAND U5898 ( .A(n5167), .B(n5166), .Z(n5168) );
  AND U5899 ( .A(n5169), .B(n5168), .Z(n5259) );
  XOR U5900 ( .A(n5260), .B(n5259), .Z(n5210) );
  NAND U5901 ( .A(n5171), .B(n5170), .Z(n5175) );
  NANDN U5902 ( .A(n5173), .B(n5172), .Z(n5174) );
  NAND U5903 ( .A(n5175), .B(n5174), .Z(n5211) );
  XNOR U5904 ( .A(n5210), .B(n5211), .Z(n5213) );
  XOR U5905 ( .A(n5212), .B(n5213), .Z(n5328) );
  NANDN U5906 ( .A(n5177), .B(n5176), .Z(n5181) );
  NANDN U5907 ( .A(n5179), .B(n5178), .Z(n5180) );
  NAND U5908 ( .A(n5181), .B(n5180), .Z(n5329) );
  XNOR U5909 ( .A(n5328), .B(n5329), .Z(n5330) );
  XOR U5910 ( .A(n5331), .B(n5330), .Z(n5341) );
  NAND U5911 ( .A(n5183), .B(n5182), .Z(n5187) );
  NANDN U5912 ( .A(n5185), .B(n5184), .Z(n5186) );
  AND U5913 ( .A(n5187), .B(n5186), .Z(n5337) );
  NANDN U5914 ( .A(n5189), .B(n5188), .Z(n5193) );
  NANDN U5915 ( .A(n5191), .B(n5190), .Z(n5192) );
  AND U5916 ( .A(n5193), .B(n5192), .Z(n5335) );
  NANDN U5917 ( .A(n5195), .B(n5194), .Z(n5199) );
  NAND U5918 ( .A(n5197), .B(n5196), .Z(n5198) );
  NAND U5919 ( .A(n5199), .B(n5198), .Z(n5334) );
  XNOR U5920 ( .A(n5335), .B(n5334), .Z(n5336) );
  XNOR U5921 ( .A(n5337), .B(n5336), .Z(n5340) );
  XOR U5922 ( .A(n5343), .B(n5342), .Z(n5348) );
  NANDN U5923 ( .A(n5201), .B(n5200), .Z(n5205) );
  NANDN U5924 ( .A(n5203), .B(n5202), .Z(n5204) );
  AND U5925 ( .A(n5205), .B(n5204), .Z(n5347) );
  XOR U5926 ( .A(n5347), .B(n5346), .Z(n5209) );
  XNOR U5927 ( .A(n5348), .B(n5209), .Z(N121) );
  NANDN U5928 ( .A(n5211), .B(n5210), .Z(n5215) );
  NAND U5929 ( .A(n5213), .B(n5212), .Z(n5214) );
  NAND U5930 ( .A(n5215), .B(n5214), .Z(n5367) );
  NANDN U5931 ( .A(n5217), .B(n5216), .Z(n5221) );
  NAND U5932 ( .A(n5219), .B(n5218), .Z(n5220) );
  AND U5933 ( .A(n5221), .B(n5220), .Z(n5372) );
  NANDN U5934 ( .A(n5223), .B(n5222), .Z(n5227) );
  NAND U5935 ( .A(n5225), .B(n5224), .Z(n5226) );
  NAND U5936 ( .A(n5227), .B(n5226), .Z(n5371) );
  XNOR U5937 ( .A(n5372), .B(n5371), .Z(n5374) );
  NAND U5938 ( .A(n5229), .B(n5228), .Z(n5233) );
  NANDN U5939 ( .A(n5231), .B(n5230), .Z(n5232) );
  AND U5940 ( .A(n5233), .B(n5232), .Z(n5404) );
  NAND U5941 ( .A(x[149]), .B(y[680]), .Z(n6283) );
  NANDN U5942 ( .A(n6283), .B(n5234), .Z(n5238) );
  NAND U5943 ( .A(n5236), .B(n5235), .Z(n5237) );
  NAND U5944 ( .A(n5238), .B(n5237), .Z(n5477) );
  NAND U5945 ( .A(x[150]), .B(y[675]), .Z(n5447) );
  NAND U5946 ( .A(x[133]), .B(y[692]), .Z(n5446) );
  NAND U5947 ( .A(x[145]), .B(y[680]), .Z(n5445) );
  XOR U5948 ( .A(n5446), .B(n5445), .Z(n5448) );
  XOR U5949 ( .A(n5447), .B(n5448), .Z(n5476) );
  AND U5950 ( .A(y[677]), .B(x[148]), .Z(n5240) );
  NAND U5951 ( .A(y[676]), .B(x[149]), .Z(n5239) );
  XNOR U5952 ( .A(n5240), .B(n5239), .Z(n5460) );
  AND U5953 ( .A(x[147]), .B(y[678]), .Z(n5459) );
  XOR U5954 ( .A(n5460), .B(n5459), .Z(n5475) );
  XNOR U5955 ( .A(n5476), .B(n5475), .Z(n5478) );
  XOR U5956 ( .A(n5477), .B(n5478), .Z(n5402) );
  NAND U5957 ( .A(n5616), .B(n5458), .Z(n5244) );
  NAND U5958 ( .A(n5242), .B(n5241), .Z(n5243) );
  NAND U5959 ( .A(n5244), .B(n5243), .Z(n5483) );
  NAND U5960 ( .A(x[143]), .B(y[682]), .Z(n5465) );
  NAND U5961 ( .A(x[146]), .B(y[679]), .Z(n5464) );
  NAND U5962 ( .A(x[134]), .B(y[691]), .Z(n5463) );
  XOR U5963 ( .A(n5464), .B(n5463), .Z(n5466) );
  XOR U5964 ( .A(n5465), .B(n5466), .Z(n5482) );
  NAND U5965 ( .A(x[151]), .B(y[674]), .Z(n5441) );
  NAND U5966 ( .A(x[132]), .B(y[693]), .Z(n5440) );
  NAND U5967 ( .A(x[144]), .B(y[681]), .Z(n5439) );
  XOR U5968 ( .A(n5440), .B(n5439), .Z(n5442) );
  XNOR U5969 ( .A(n5441), .B(n5442), .Z(n5481) );
  XOR U5970 ( .A(n5482), .B(n5481), .Z(n5484) );
  XOR U5971 ( .A(n5483), .B(n5484), .Z(n5401) );
  XOR U5972 ( .A(n5404), .B(n5403), .Z(n5416) );
  NAND U5973 ( .A(n5246), .B(n5245), .Z(n5250) );
  NANDN U5974 ( .A(n5248), .B(n5247), .Z(n5249) );
  AND U5975 ( .A(n5250), .B(n5249), .Z(n5414) );
  NAND U5976 ( .A(n5252), .B(n5251), .Z(n5256) );
  NANDN U5977 ( .A(n5254), .B(n5253), .Z(n5255) );
  NAND U5978 ( .A(n5256), .B(n5255), .Z(n5413) );
  XNOR U5979 ( .A(n5414), .B(n5413), .Z(n5415) );
  XNOR U5980 ( .A(n5416), .B(n5415), .Z(n5373) );
  XOR U5981 ( .A(n5374), .B(n5373), .Z(n5366) );
  NAND U5982 ( .A(n5258), .B(n5257), .Z(n5262) );
  NAND U5983 ( .A(n5260), .B(n5259), .Z(n5261) );
  NAND U5984 ( .A(n5262), .B(n5261), .Z(n5365) );
  XNOR U5985 ( .A(n5367), .B(n5368), .Z(n5361) );
  NAND U5986 ( .A(n5383), .B(n5263), .Z(n5267) );
  NAND U5987 ( .A(n5265), .B(n5264), .Z(n5266) );
  AND U5988 ( .A(n5267), .B(n5266), .Z(n5408) );
  AND U5989 ( .A(x[142]), .B(y[688]), .Z(n6269) );
  NAND U5990 ( .A(n6269), .B(n5268), .Z(n5272) );
  NANDN U5991 ( .A(n5270), .B(n5269), .Z(n5271) );
  AND U5992 ( .A(n5272), .B(n5271), .Z(n5436) );
  NAND U5993 ( .A(x[139]), .B(y[686]), .Z(n5454) );
  NAND U5994 ( .A(x[140]), .B(y[685]), .Z(n5453) );
  NAND U5995 ( .A(x[135]), .B(y[690]), .Z(n5452) );
  XNOR U5996 ( .A(n5453), .B(n5452), .Z(n5455) );
  XOR U5997 ( .A(n5454), .B(n5455), .Z(n5433) );
  AND U5998 ( .A(x[152]), .B(y[673]), .Z(n5451) );
  XOR U5999 ( .A(o[57]), .B(n5451), .Z(n5421) );
  NAND U6000 ( .A(x[129]), .B(y[696]), .Z(n5422) );
  XNOR U6001 ( .A(n5421), .B(n5422), .Z(n5423) );
  NAND U6002 ( .A(x[141]), .B(y[684]), .Z(n5424) );
  XNOR U6003 ( .A(n5423), .B(n5424), .Z(n5434) );
  XOR U6004 ( .A(n5433), .B(n5434), .Z(n5435) );
  XNOR U6005 ( .A(n5436), .B(n5435), .Z(n5407) );
  XNOR U6006 ( .A(n5408), .B(n5407), .Z(n5410) );
  NAND U6007 ( .A(n5274), .B(n5273), .Z(n5278) );
  AND U6008 ( .A(n5276), .B(n5275), .Z(n5277) );
  ANDN U6009 ( .B(n5278), .A(n5277), .Z(n5396) );
  AND U6010 ( .A(n5280), .B(n5279), .Z(n5284) );
  NAND U6011 ( .A(n5282), .B(n5281), .Z(n5283) );
  NANDN U6012 ( .A(n5284), .B(n5283), .Z(n5395) );
  XNOR U6013 ( .A(n5396), .B(n5395), .Z(n5398) );
  NAND U6014 ( .A(n5286), .B(n5285), .Z(n5290) );
  NAND U6015 ( .A(n5288), .B(n5287), .Z(n5289) );
  AND U6016 ( .A(n5290), .B(n5289), .Z(n5392) );
  AND U6017 ( .A(x[136]), .B(y[689]), .Z(n5386) );
  XOR U6018 ( .A(n5384), .B(n5383), .Z(n5385) );
  XOR U6019 ( .A(n5386), .B(n5385), .Z(n5390) );
  AND U6020 ( .A(n5291), .B(o[56]), .Z(n5380) );
  AND U6021 ( .A(x[153]), .B(y[672]), .Z(n5378) );
  NAND U6022 ( .A(x[128]), .B(y[697]), .Z(n5377) );
  XNOR U6023 ( .A(n5378), .B(n5377), .Z(n5379) );
  XOR U6024 ( .A(n5380), .B(n5379), .Z(n5389) );
  XOR U6025 ( .A(n5390), .B(n5389), .Z(n5391) );
  XNOR U6026 ( .A(n5392), .B(n5391), .Z(n5397) );
  XOR U6027 ( .A(n5398), .B(n5397), .Z(n5409) );
  XOR U6028 ( .A(n5410), .B(n5409), .Z(n5490) );
  NANDN U6029 ( .A(n5293), .B(n5292), .Z(n5297) );
  NAND U6030 ( .A(n5295), .B(n5294), .Z(n5296) );
  AND U6031 ( .A(n5297), .B(n5296), .Z(n5488) );
  NAND U6032 ( .A(n5299), .B(n5298), .Z(n5303) );
  ANDN U6033 ( .B(n5301), .A(n5300), .Z(n5302) );
  ANDN U6034 ( .B(n5303), .A(n5302), .Z(n5472) );
  NAND U6035 ( .A(n5305), .B(n5304), .Z(n5309) );
  NAND U6036 ( .A(n5307), .B(n5306), .Z(n5308) );
  AND U6037 ( .A(n5309), .B(n5308), .Z(n5470) );
  AND U6038 ( .A(x[142]), .B(y[683]), .Z(n5427) );
  NAND U6039 ( .A(x[130]), .B(y[695]), .Z(n5428) );
  XNOR U6040 ( .A(n5427), .B(n5428), .Z(n5429) );
  NAND U6041 ( .A(x[131]), .B(y[694]), .Z(n5430) );
  XNOR U6042 ( .A(n5429), .B(n5430), .Z(n5469) );
  XNOR U6043 ( .A(n5470), .B(n5469), .Z(n5471) );
  XOR U6044 ( .A(n5472), .B(n5471), .Z(n5487) );
  XOR U6045 ( .A(n5488), .B(n5487), .Z(n5489) );
  NAND U6046 ( .A(n5311), .B(n5310), .Z(n5315) );
  NAND U6047 ( .A(n5313), .B(n5312), .Z(n5314) );
  NAND U6048 ( .A(n5315), .B(n5314), .Z(n5494) );
  XNOR U6049 ( .A(n5493), .B(n5494), .Z(n5495) );
  NANDN U6050 ( .A(n5317), .B(n5316), .Z(n5321) );
  NANDN U6051 ( .A(n5319), .B(n5318), .Z(n5320) );
  NAND U6052 ( .A(n5321), .B(n5320), .Z(n5496) );
  XNOR U6053 ( .A(n5495), .B(n5496), .Z(n5360) );
  NANDN U6054 ( .A(n5323), .B(n5322), .Z(n5327) );
  NANDN U6055 ( .A(n5325), .B(n5324), .Z(n5326) );
  AND U6056 ( .A(n5327), .B(n5326), .Z(n5359) );
  XOR U6057 ( .A(n5361), .B(n5362), .Z(n5351) );
  NANDN U6058 ( .A(n5329), .B(n5328), .Z(n5333) );
  NAND U6059 ( .A(n5331), .B(n5330), .Z(n5332) );
  NAND U6060 ( .A(n5333), .B(n5332), .Z(n5350) );
  XOR U6061 ( .A(n5351), .B(n5350), .Z(n5352) );
  NANDN U6062 ( .A(n5335), .B(n5334), .Z(n5339) );
  NANDN U6063 ( .A(n5337), .B(n5336), .Z(n5338) );
  NAND U6064 ( .A(n5339), .B(n5338), .Z(n5353) );
  XNOR U6065 ( .A(n5352), .B(n5353), .Z(n5358) );
  NANDN U6066 ( .A(n5341), .B(n5340), .Z(n5345) );
  NANDN U6067 ( .A(n5343), .B(n5342), .Z(n5344) );
  NAND U6068 ( .A(n5345), .B(n5344), .Z(n5356) );
  XOR U6069 ( .A(n5356), .B(n5357), .Z(n5349) );
  XNOR U6070 ( .A(n5358), .B(n5349), .Z(N122) );
  NAND U6071 ( .A(n5351), .B(n5350), .Z(n5355) );
  NANDN U6072 ( .A(n5353), .B(n5352), .Z(n5354) );
  NAND U6073 ( .A(n5355), .B(n5354), .Z(n5650) );
  IV U6074 ( .A(n5650), .Z(n5648) );
  NANDN U6075 ( .A(n5360), .B(n5359), .Z(n5364) );
  NANDN U6076 ( .A(n5362), .B(n5361), .Z(n5363) );
  NAND U6077 ( .A(n5364), .B(n5363), .Z(n5655) );
  NANDN U6078 ( .A(n5366), .B(n5365), .Z(n5370) );
  NAND U6079 ( .A(n5368), .B(n5367), .Z(n5369) );
  AND U6080 ( .A(n5370), .B(n5369), .Z(n5656) );
  XOR U6081 ( .A(n5655), .B(n5656), .Z(n5658) );
  NANDN U6082 ( .A(n5372), .B(n5371), .Z(n5376) );
  NAND U6083 ( .A(n5374), .B(n5373), .Z(n5375) );
  AND U6084 ( .A(n5376), .B(n5375), .Z(n5645) );
  AND U6085 ( .A(x[130]), .B(y[696]), .Z(n5518) );
  XOR U6086 ( .A(n5519), .B(n5518), .Z(n5521) );
  AND U6087 ( .A(x[152]), .B(y[674]), .Z(n5520) );
  XOR U6088 ( .A(n5521), .B(n5520), .Z(n5555) );
  NANDN U6089 ( .A(n5378), .B(n5377), .Z(n5382) );
  NANDN U6090 ( .A(n5380), .B(n5379), .Z(n5381) );
  AND U6091 ( .A(n5382), .B(n5381), .Z(n5554) );
  XOR U6092 ( .A(n5555), .B(n5554), .Z(n5557) );
  OR U6093 ( .A(n5384), .B(n5383), .Z(n5388) );
  NANDN U6094 ( .A(n5386), .B(n5385), .Z(n5387) );
  AND U6095 ( .A(n5388), .B(n5387), .Z(n5556) );
  XOR U6096 ( .A(n5557), .B(n5556), .Z(n5593) );
  NAND U6097 ( .A(n5390), .B(n5389), .Z(n5394) );
  NANDN U6098 ( .A(n5392), .B(n5391), .Z(n5393) );
  AND U6099 ( .A(n5394), .B(n5393), .Z(n5592) );
  XNOR U6100 ( .A(n5593), .B(n5592), .Z(n5595) );
  NANDN U6101 ( .A(n5396), .B(n5395), .Z(n5400) );
  NAND U6102 ( .A(n5398), .B(n5397), .Z(n5399) );
  AND U6103 ( .A(n5400), .B(n5399), .Z(n5594) );
  XOR U6104 ( .A(n5595), .B(n5594), .Z(n5639) );
  NANDN U6105 ( .A(n5402), .B(n5401), .Z(n5406) );
  NAND U6106 ( .A(n5404), .B(n5403), .Z(n5405) );
  NAND U6107 ( .A(n5406), .B(n5405), .Z(n5636) );
  NANDN U6108 ( .A(n5408), .B(n5407), .Z(n5412) );
  NAND U6109 ( .A(n5410), .B(n5409), .Z(n5411) );
  AND U6110 ( .A(n5412), .B(n5411), .Z(n5637) );
  XOR U6111 ( .A(n5636), .B(n5637), .Z(n5638) );
  XOR U6112 ( .A(n5639), .B(n5638), .Z(n5643) );
  NANDN U6113 ( .A(n5414), .B(n5413), .Z(n5418) );
  NANDN U6114 ( .A(n5416), .B(n5415), .Z(n5417) );
  NAND U6115 ( .A(n5418), .B(n5417), .Z(n5588) );
  AND U6116 ( .A(y[692]), .B(x[134]), .Z(n5420) );
  NAND U6117 ( .A(y[690]), .B(x[136]), .Z(n5419) );
  XNOR U6118 ( .A(n5420), .B(n5419), .Z(n5618) );
  AND U6119 ( .A(x[137]), .B(y[689]), .Z(n5617) );
  XOR U6120 ( .A(n5618), .B(n5617), .Z(n5599) );
  AND U6121 ( .A(x[135]), .B(y[691]), .Z(n5598) );
  XOR U6122 ( .A(n5599), .B(n5598), .Z(n5601) );
  AND U6123 ( .A(x[140]), .B(y[686]), .Z(n5712) );
  AND U6124 ( .A(x[133]), .B(y[693]), .Z(n5569) );
  XOR U6125 ( .A(n5712), .B(n5569), .Z(n5571) );
  AND U6126 ( .A(x[138]), .B(y[688]), .Z(n5570) );
  XOR U6127 ( .A(n5571), .B(n5570), .Z(n5600) );
  XOR U6128 ( .A(n5601), .B(n5600), .Z(n5544) );
  NANDN U6129 ( .A(n5422), .B(n5421), .Z(n5426) );
  NANDN U6130 ( .A(n5424), .B(n5423), .Z(n5425) );
  NAND U6131 ( .A(n5426), .B(n5425), .Z(n5543) );
  NANDN U6132 ( .A(n5428), .B(n5427), .Z(n5432) );
  NANDN U6133 ( .A(n5430), .B(n5429), .Z(n5431) );
  NAND U6134 ( .A(n5432), .B(n5431), .Z(n5542) );
  XNOR U6135 ( .A(n5543), .B(n5542), .Z(n5545) );
  XNOR U6136 ( .A(n5544), .B(n5545), .Z(n5581) );
  NAND U6137 ( .A(n5434), .B(n5433), .Z(n5438) );
  NANDN U6138 ( .A(n5436), .B(n5435), .Z(n5437) );
  AND U6139 ( .A(n5438), .B(n5437), .Z(n5580) );
  XNOR U6140 ( .A(n5581), .B(n5580), .Z(n5582) );
  NAND U6141 ( .A(n5440), .B(n5439), .Z(n5444) );
  NAND U6142 ( .A(n5442), .B(n5441), .Z(n5443) );
  AND U6143 ( .A(n5444), .B(n5443), .Z(n5507) );
  NAND U6144 ( .A(n5446), .B(n5445), .Z(n5450) );
  NAND U6145 ( .A(n5448), .B(n5447), .Z(n5449) );
  AND U6146 ( .A(n5450), .B(n5449), .Z(n5506) );
  XOR U6147 ( .A(n5507), .B(n5506), .Z(n5509) );
  AND U6148 ( .A(n5451), .B(o[57]), .Z(n5611) );
  AND U6149 ( .A(x[142]), .B(y[684]), .Z(n5610) );
  XOR U6150 ( .A(n5611), .B(n5610), .Z(n5613) );
  AND U6151 ( .A(x[129]), .B(y[697]), .Z(n5612) );
  XOR U6152 ( .A(n5613), .B(n5612), .Z(n5561) );
  AND U6153 ( .A(x[153]), .B(y[673]), .Z(n5621) );
  XOR U6154 ( .A(o[58]), .B(n5621), .Z(n5575) );
  AND U6155 ( .A(x[154]), .B(y[672]), .Z(n5574) );
  XOR U6156 ( .A(n5575), .B(n5574), .Z(n5577) );
  AND U6157 ( .A(x[128]), .B(y[698]), .Z(n5576) );
  XOR U6158 ( .A(n5577), .B(n5576), .Z(n5560) );
  XOR U6159 ( .A(n5561), .B(n5560), .Z(n5563) );
  NAND U6160 ( .A(n5453), .B(n5452), .Z(n5457) );
  NANDN U6161 ( .A(n5455), .B(n5454), .Z(n5456) );
  AND U6162 ( .A(n5457), .B(n5456), .Z(n5562) );
  XOR U6163 ( .A(n5563), .B(n5562), .Z(n5508) );
  XNOR U6164 ( .A(n5509), .B(n5508), .Z(n5550) );
  NAND U6165 ( .A(x[149]), .B(y[677]), .Z(n5604) );
  NANDN U6166 ( .A(n5604), .B(n5458), .Z(n5462) );
  NAND U6167 ( .A(n5460), .B(n5459), .Z(n5461) );
  NAND U6168 ( .A(n5462), .B(n5461), .Z(n5538) );
  AND U6169 ( .A(x[148]), .B(y[678]), .Z(n5606) );
  XOR U6170 ( .A(n5607), .B(n5606), .Z(n5537) );
  AND U6171 ( .A(x[151]), .B(y[675]), .Z(n5524) );
  XOR U6172 ( .A(n5525), .B(n5524), .Z(n5527) );
  AND U6173 ( .A(x[150]), .B(y[676]), .Z(n5526) );
  XOR U6174 ( .A(n5527), .B(n5526), .Z(n5536) );
  XOR U6175 ( .A(n5537), .B(n5536), .Z(n5539) );
  XOR U6176 ( .A(n5538), .B(n5539), .Z(n5549) );
  AND U6177 ( .A(x[147]), .B(y[679]), .Z(n5623) );
  AND U6178 ( .A(x[131]), .B(y[695]), .Z(n5622) );
  XOR U6179 ( .A(n5623), .B(n5622), .Z(n5625) );
  AND U6180 ( .A(x[139]), .B(y[687]), .Z(n5624) );
  XOR U6181 ( .A(n5625), .B(n5624), .Z(n5513) );
  AND U6182 ( .A(x[132]), .B(y[694]), .Z(n5530) );
  XOR U6183 ( .A(n5531), .B(n5530), .Z(n5533) );
  XOR U6184 ( .A(n5533), .B(n5532), .Z(n5512) );
  XOR U6185 ( .A(n5513), .B(n5512), .Z(n5515) );
  NAND U6186 ( .A(n5464), .B(n5463), .Z(n5468) );
  NAND U6187 ( .A(n5466), .B(n5465), .Z(n5467) );
  AND U6188 ( .A(n5468), .B(n5467), .Z(n5514) );
  XNOR U6189 ( .A(n5515), .B(n5514), .Z(n5548) );
  XOR U6190 ( .A(n5549), .B(n5548), .Z(n5551) );
  XOR U6191 ( .A(n5550), .B(n5551), .Z(n5583) );
  XNOR U6192 ( .A(n5582), .B(n5583), .Z(n5587) );
  NANDN U6193 ( .A(n5470), .B(n5469), .Z(n5474) );
  NANDN U6194 ( .A(n5472), .B(n5471), .Z(n5473) );
  NAND U6195 ( .A(n5474), .B(n5473), .Z(n5632) );
  NANDN U6196 ( .A(n5476), .B(n5475), .Z(n5480) );
  NAND U6197 ( .A(n5478), .B(n5477), .Z(n5479) );
  NAND U6198 ( .A(n5480), .B(n5479), .Z(n5631) );
  NANDN U6199 ( .A(n5482), .B(n5481), .Z(n5486) );
  NANDN U6200 ( .A(n5484), .B(n5483), .Z(n5485) );
  NAND U6201 ( .A(n5486), .B(n5485), .Z(n5630) );
  XOR U6202 ( .A(n5631), .B(n5630), .Z(n5633) );
  XOR U6203 ( .A(n5632), .B(n5633), .Z(n5586) );
  XNOR U6204 ( .A(n5587), .B(n5586), .Z(n5589) );
  XOR U6205 ( .A(n5588), .B(n5589), .Z(n5642) );
  XNOR U6206 ( .A(n5643), .B(n5642), .Z(n5644) );
  XNOR U6207 ( .A(n5645), .B(n5644), .Z(n5503) );
  NAND U6208 ( .A(n5488), .B(n5487), .Z(n5492) );
  NANDN U6209 ( .A(n5490), .B(n5489), .Z(n5491) );
  AND U6210 ( .A(n5492), .B(n5491), .Z(n5500) );
  NANDN U6211 ( .A(n5494), .B(n5493), .Z(n5498) );
  NANDN U6212 ( .A(n5496), .B(n5495), .Z(n5497) );
  NAND U6213 ( .A(n5498), .B(n5497), .Z(n5501) );
  XNOR U6214 ( .A(n5500), .B(n5501), .Z(n5502) );
  XOR U6215 ( .A(n5503), .B(n5502), .Z(n5657) );
  XOR U6216 ( .A(n5658), .B(n5657), .Z(n5651) );
  XNOR U6217 ( .A(n5649), .B(n5651), .Z(n5499) );
  XOR U6218 ( .A(n5648), .B(n5499), .Z(N123) );
  NANDN U6219 ( .A(n5501), .B(n5500), .Z(n5505) );
  NAND U6220 ( .A(n5503), .B(n5502), .Z(n5504) );
  AND U6221 ( .A(n5505), .B(n5504), .Z(n5802) );
  NAND U6222 ( .A(n5507), .B(n5506), .Z(n5511) );
  NAND U6223 ( .A(n5509), .B(n5508), .Z(n5510) );
  NAND U6224 ( .A(n5511), .B(n5510), .Z(n5774) );
  NAND U6225 ( .A(n5513), .B(n5512), .Z(n5517) );
  NAND U6226 ( .A(n5515), .B(n5514), .Z(n5516) );
  NAND U6227 ( .A(n5517), .B(n5516), .Z(n5772) );
  AND U6228 ( .A(n5519), .B(n5518), .Z(n5523) );
  NAND U6229 ( .A(n5521), .B(n5520), .Z(n5522) );
  NANDN U6230 ( .A(n5523), .B(n5522), .Z(n5687) );
  NAND U6231 ( .A(n5525), .B(n5524), .Z(n5529) );
  NAND U6232 ( .A(n5527), .B(n5526), .Z(n5528) );
  NAND U6233 ( .A(n5529), .B(n5528), .Z(n5686) );
  XOR U6234 ( .A(n5687), .B(n5686), .Z(n5688) );
  NAND U6235 ( .A(n5531), .B(n5530), .Z(n5535) );
  NAND U6236 ( .A(n5533), .B(n5532), .Z(n5534) );
  NAND U6237 ( .A(n5535), .B(n5534), .Z(n5700) );
  AND U6238 ( .A(x[128]), .B(y[699]), .Z(n5755) );
  AND U6239 ( .A(x[155]), .B(y[672]), .Z(n5754) );
  XOR U6240 ( .A(n5755), .B(n5754), .Z(n5757) );
  AND U6241 ( .A(x[154]), .B(y[673]), .Z(n5762) );
  XOR U6242 ( .A(n5762), .B(o[59]), .Z(n5756) );
  XOR U6243 ( .A(n5757), .B(n5756), .Z(n5699) );
  AND U6244 ( .A(x[137]), .B(y[690]), .Z(n5759) );
  AND U6245 ( .A(x[149]), .B(y[678]), .Z(n5758) );
  XOR U6246 ( .A(n5759), .B(n5758), .Z(n5761) );
  AND U6247 ( .A(x[146]), .B(y[681]), .Z(n5760) );
  XOR U6248 ( .A(n5761), .B(n5760), .Z(n5698) );
  XOR U6249 ( .A(n5699), .B(n5698), .Z(n5701) );
  XNOR U6250 ( .A(n5700), .B(n5701), .Z(n5689) );
  XOR U6251 ( .A(n5772), .B(n5773), .Z(n5775) );
  XOR U6252 ( .A(n5774), .B(n5775), .Z(n5793) );
  NAND U6253 ( .A(n5537), .B(n5536), .Z(n5541) );
  NAND U6254 ( .A(n5539), .B(n5538), .Z(n5540) );
  AND U6255 ( .A(n5541), .B(n5540), .Z(n5791) );
  NAND U6256 ( .A(n5543), .B(n5542), .Z(n5547) );
  NANDN U6257 ( .A(n5545), .B(n5544), .Z(n5546) );
  AND U6258 ( .A(n5547), .B(n5546), .Z(n5790) );
  XOR U6259 ( .A(n5791), .B(n5790), .Z(n5792) );
  NANDN U6260 ( .A(n5549), .B(n5548), .Z(n5553) );
  NANDN U6261 ( .A(n5551), .B(n5550), .Z(n5552) );
  AND U6262 ( .A(n5553), .B(n5552), .Z(n5778) );
  NAND U6263 ( .A(n5555), .B(n5554), .Z(n5559) );
  NAND U6264 ( .A(n5557), .B(n5556), .Z(n5558) );
  NAND U6265 ( .A(n5559), .B(n5558), .Z(n5768) );
  NAND U6266 ( .A(n5561), .B(n5560), .Z(n5565) );
  NAND U6267 ( .A(n5563), .B(n5562), .Z(n5564) );
  NAND U6268 ( .A(n5565), .B(n5564), .Z(n5766) );
  AND U6269 ( .A(x[147]), .B(y[680]), .Z(n5747) );
  AND U6270 ( .A(x[153]), .B(y[674]), .Z(n5746) );
  XOR U6271 ( .A(n5747), .B(n5746), .Z(n5749) );
  AND U6272 ( .A(x[134]), .B(y[693]), .Z(n5748) );
  XOR U6273 ( .A(n5749), .B(n5748), .Z(n5738) );
  AND U6274 ( .A(x[143]), .B(y[684]), .Z(n5718) );
  AND U6275 ( .A(x[130]), .B(y[697]), .Z(n5717) );
  XOR U6276 ( .A(n5718), .B(n5717), .Z(n5720) );
  AND U6277 ( .A(x[131]), .B(y[696]), .Z(n5719) );
  XOR U6278 ( .A(n5720), .B(n5719), .Z(n5737) );
  XOR U6279 ( .A(n5738), .B(n5737), .Z(n5739) );
  NAND U6280 ( .A(x[144]), .B(y[683]), .Z(n5704) );
  XOR U6281 ( .A(n5704), .B(n5566), .Z(n5707) );
  XOR U6282 ( .A(n5706), .B(n5707), .Z(n5714) );
  AND U6283 ( .A(y[686]), .B(x[141]), .Z(n5568) );
  AND U6284 ( .A(y[687]), .B(x[140]), .Z(n5567) );
  XOR U6285 ( .A(n5568), .B(n5567), .Z(n5713) );
  XOR U6286 ( .A(n5714), .B(n5713), .Z(n5740) );
  AND U6287 ( .A(n5712), .B(n5569), .Z(n5573) );
  NAND U6288 ( .A(n5571), .B(n5570), .Z(n5572) );
  NANDN U6289 ( .A(n5573), .B(n5572), .Z(n5681) );
  NAND U6290 ( .A(n5575), .B(n5574), .Z(n5579) );
  NAND U6291 ( .A(n5577), .B(n5576), .Z(n5578) );
  NAND U6292 ( .A(n5579), .B(n5578), .Z(n5680) );
  XOR U6293 ( .A(n5681), .B(n5680), .Z(n5682) );
  XOR U6294 ( .A(n5683), .B(n5682), .Z(n5767) );
  XNOR U6295 ( .A(n5766), .B(n5767), .Z(n5769) );
  XNOR U6296 ( .A(n5778), .B(n5779), .Z(n5781) );
  NANDN U6297 ( .A(n5581), .B(n5580), .Z(n5585) );
  NANDN U6298 ( .A(n5583), .B(n5582), .Z(n5584) );
  AND U6299 ( .A(n5585), .B(n5584), .Z(n5780) );
  XOR U6300 ( .A(n5781), .B(n5780), .Z(n5668) );
  NANDN U6301 ( .A(n5587), .B(n5586), .Z(n5591) );
  NAND U6302 ( .A(n5589), .B(n5588), .Z(n5590) );
  NAND U6303 ( .A(n5591), .B(n5590), .Z(n5670) );
  XOR U6304 ( .A(n5671), .B(n5670), .Z(n5665) );
  NANDN U6305 ( .A(n5593), .B(n5592), .Z(n5597) );
  NAND U6306 ( .A(n5595), .B(n5594), .Z(n5596) );
  NAND U6307 ( .A(n5597), .B(n5596), .Z(n5675) );
  NAND U6308 ( .A(n5599), .B(n5598), .Z(n5603) );
  NAND U6309 ( .A(n5601), .B(n5600), .Z(n5602) );
  NAND U6310 ( .A(n5603), .B(n5602), .Z(n5786) );
  ANDN U6311 ( .B(n5605), .A(n5604), .Z(n5609) );
  NAND U6312 ( .A(n5607), .B(n5606), .Z(n5608) );
  NANDN U6313 ( .A(n5609), .B(n5608), .Z(n5726) );
  NAND U6314 ( .A(n5611), .B(n5610), .Z(n5615) );
  NAND U6315 ( .A(n5613), .B(n5612), .Z(n5614) );
  NAND U6316 ( .A(n5615), .B(n5614), .Z(n5725) );
  XOR U6317 ( .A(n5726), .B(n5725), .Z(n5727) );
  AND U6318 ( .A(x[136]), .B(y[692]), .Z(n5764) );
  NAND U6319 ( .A(n5764), .B(n5616), .Z(n5620) );
  NAND U6320 ( .A(n5618), .B(n5617), .Z(n5619) );
  NAND U6321 ( .A(n5620), .B(n5619), .Z(n5694) );
  AND U6322 ( .A(x[142]), .B(y[685]), .Z(n5722) );
  AND U6323 ( .A(x[129]), .B(y[698]), .Z(n5721) );
  XOR U6324 ( .A(n5722), .B(n5721), .Z(n5723) );
  XOR U6325 ( .A(n5723), .B(n5724), .Z(n5693) );
  AND U6326 ( .A(x[145]), .B(y[682]), .Z(n5751) );
  AND U6327 ( .A(x[132]), .B(y[695]), .Z(n5750) );
  XOR U6328 ( .A(n5751), .B(n5750), .Z(n5753) );
  AND U6329 ( .A(x[133]), .B(y[694]), .Z(n5752) );
  XOR U6330 ( .A(n5753), .B(n5752), .Z(n5692) );
  XOR U6331 ( .A(n5693), .B(n5692), .Z(n5695) );
  XNOR U6332 ( .A(n5694), .B(n5695), .Z(n5728) );
  NAND U6333 ( .A(n5623), .B(n5622), .Z(n5627) );
  NAND U6334 ( .A(n5625), .B(n5624), .Z(n5626) );
  NAND U6335 ( .A(n5627), .B(n5626), .Z(n5733) );
  NAND U6336 ( .A(y[675]), .B(x[152]), .Z(n5628) );
  XNOR U6337 ( .A(n5629), .B(n5628), .Z(n5745) );
  AND U6338 ( .A(x[135]), .B(y[692]), .Z(n5744) );
  XOR U6339 ( .A(n5745), .B(n5744), .Z(n5732) );
  AND U6340 ( .A(x[136]), .B(y[691]), .Z(n5709) );
  AND U6341 ( .A(x[151]), .B(y[676]), .Z(n5708) );
  XOR U6342 ( .A(n5709), .B(n5708), .Z(n5711) );
  AND U6343 ( .A(x[150]), .B(y[677]), .Z(n5710) );
  XOR U6344 ( .A(n5711), .B(n5710), .Z(n5731) );
  XOR U6345 ( .A(n5732), .B(n5731), .Z(n5734) );
  XOR U6346 ( .A(n5733), .B(n5734), .Z(n5784) );
  XOR U6347 ( .A(n5785), .B(n5784), .Z(n5787) );
  XNOR U6348 ( .A(n5786), .B(n5787), .Z(n5674) );
  XOR U6349 ( .A(n5675), .B(n5674), .Z(n5677) );
  NAND U6350 ( .A(n5631), .B(n5630), .Z(n5635) );
  NAND U6351 ( .A(n5633), .B(n5632), .Z(n5634) );
  AND U6352 ( .A(n5635), .B(n5634), .Z(n5676) );
  XOR U6353 ( .A(n5677), .B(n5676), .Z(n5663) );
  NAND U6354 ( .A(n5637), .B(n5636), .Z(n5641) );
  NAND U6355 ( .A(n5639), .B(n5638), .Z(n5640) );
  AND U6356 ( .A(n5641), .B(n5640), .Z(n5662) );
  XOR U6357 ( .A(n5665), .B(n5664), .Z(n5800) );
  NANDN U6358 ( .A(n5643), .B(n5642), .Z(n5647) );
  NANDN U6359 ( .A(n5645), .B(n5644), .Z(n5646) );
  AND U6360 ( .A(n5647), .B(n5646), .Z(n5799) );
  XNOR U6361 ( .A(n5800), .B(n5799), .Z(n5801) );
  XNOR U6362 ( .A(n5802), .B(n5801), .Z(n5798) );
  NANDN U6363 ( .A(n5648), .B(n5649), .Z(n5654) );
  NOR U6364 ( .A(n5650), .B(n5649), .Z(n5652) );
  OR U6365 ( .A(n5652), .B(n5651), .Z(n5653) );
  AND U6366 ( .A(n5654), .B(n5653), .Z(n5797) );
  NAND U6367 ( .A(n5656), .B(n5655), .Z(n5660) );
  NAND U6368 ( .A(n5658), .B(n5657), .Z(n5659) );
  AND U6369 ( .A(n5660), .B(n5659), .Z(n5796) );
  XOR U6370 ( .A(n5797), .B(n5796), .Z(n5661) );
  XNOR U6371 ( .A(n5798), .B(n5661), .Z(N124) );
  NANDN U6372 ( .A(n5663), .B(n5662), .Z(n5667) );
  NAND U6373 ( .A(n5665), .B(n5664), .Z(n5666) );
  NAND U6374 ( .A(n5667), .B(n5666), .Z(n5935) );
  NANDN U6375 ( .A(n5669), .B(n5668), .Z(n5673) );
  NAND U6376 ( .A(n5671), .B(n5670), .Z(n5672) );
  NAND U6377 ( .A(n5673), .B(n5672), .Z(n5934) );
  XOR U6378 ( .A(n5935), .B(n5934), .Z(n5937) );
  NAND U6379 ( .A(n5675), .B(n5674), .Z(n5679) );
  NAND U6380 ( .A(n5677), .B(n5676), .Z(n5678) );
  AND U6381 ( .A(n5679), .B(n5678), .Z(n5806) );
  NAND U6382 ( .A(n5681), .B(n5680), .Z(n5685) );
  NAND U6383 ( .A(n5683), .B(n5682), .Z(n5684) );
  NAND U6384 ( .A(n5685), .B(n5684), .Z(n5830) );
  NAND U6385 ( .A(n5687), .B(n5686), .Z(n5691) );
  NANDN U6386 ( .A(n5689), .B(n5688), .Z(n5690) );
  NAND U6387 ( .A(n5691), .B(n5690), .Z(n5912) );
  NAND U6388 ( .A(n5693), .B(n5692), .Z(n5697) );
  NAND U6389 ( .A(n5695), .B(n5694), .Z(n5696) );
  NAND U6390 ( .A(n5697), .B(n5696), .Z(n5911) );
  NAND U6391 ( .A(n5699), .B(n5698), .Z(n5703) );
  NAND U6392 ( .A(n5701), .B(n5700), .Z(n5702) );
  NAND U6393 ( .A(n5703), .B(n5702), .Z(n5910) );
  XOR U6394 ( .A(n5911), .B(n5910), .Z(n5913) );
  XOR U6395 ( .A(n5912), .B(n5913), .Z(n5831) );
  XOR U6396 ( .A(n5830), .B(n5831), .Z(n5833) );
  AND U6397 ( .A(x[135]), .B(y[693]), .Z(n5869) );
  AND U6398 ( .A(x[140]), .B(y[688]), .Z(n5868) );
  XOR U6399 ( .A(n5869), .B(n5868), .Z(n5871) );
  AND U6400 ( .A(x[139]), .B(y[689]), .Z(n5870) );
  XOR U6401 ( .A(n5871), .B(n5870), .Z(n5891) );
  AND U6402 ( .A(x[155]), .B(y[673]), .Z(n5879) );
  XOR U6403 ( .A(o[60]), .B(n5879), .Z(n5883) );
  AND U6404 ( .A(x[154]), .B(y[674]), .Z(n5882) );
  XOR U6405 ( .A(n5883), .B(n5882), .Z(n5885) );
  AND U6406 ( .A(x[143]), .B(y[685]), .Z(n5884) );
  XNOR U6407 ( .A(n5885), .B(n5884), .Z(n5890) );
  XNOR U6408 ( .A(n5891), .B(n5890), .Z(n5893) );
  XOR U6409 ( .A(n5892), .B(n5893), .Z(n5917) );
  AND U6410 ( .A(x[145]), .B(y[683]), .Z(n5841) );
  AND U6411 ( .A(x[150]), .B(y[678]), .Z(n5840) );
  XOR U6412 ( .A(n5841), .B(n5840), .Z(n5843) );
  AND U6413 ( .A(x[132]), .B(y[696]), .Z(n5842) );
  XOR U6414 ( .A(n5843), .B(n5842), .Z(n5895) );
  AND U6415 ( .A(x[134]), .B(y[694]), .Z(n6020) );
  AND U6416 ( .A(x[147]), .B(y[681]), .Z(n5872) );
  XOR U6417 ( .A(n6020), .B(n5872), .Z(n5874) );
  XOR U6418 ( .A(n5874), .B(n5873), .Z(n5894) );
  XOR U6419 ( .A(n5895), .B(n5894), .Z(n5897) );
  XOR U6420 ( .A(n5896), .B(n5897), .Z(n5916) );
  NAND U6421 ( .A(n5887), .B(n5712), .Z(n5716) );
  NANDN U6422 ( .A(n5714), .B(n5713), .Z(n5715) );
  NAND U6423 ( .A(n5716), .B(n5715), .Z(n5838) );
  XOR U6424 ( .A(n5836), .B(n5837), .Z(n5839) );
  XOR U6425 ( .A(n5838), .B(n5839), .Z(n5918) );
  XOR U6426 ( .A(n5919), .B(n5918), .Z(n5832) );
  XNOR U6427 ( .A(n5833), .B(n5832), .Z(n5827) );
  NAND U6428 ( .A(n5726), .B(n5725), .Z(n5730) );
  NANDN U6429 ( .A(n5728), .B(n5727), .Z(n5729) );
  NAND U6430 ( .A(n5730), .B(n5729), .Z(n5900) );
  NAND U6431 ( .A(n5732), .B(n5731), .Z(n5736) );
  NAND U6432 ( .A(n5734), .B(n5733), .Z(n5735) );
  NAND U6433 ( .A(n5736), .B(n5735), .Z(n5899) );
  NAND U6434 ( .A(n5738), .B(n5737), .Z(n5742) );
  NANDN U6435 ( .A(n5740), .B(n5739), .Z(n5741) );
  NAND U6436 ( .A(n5742), .B(n5741), .Z(n5898) );
  XOR U6437 ( .A(n5899), .B(n5898), .Z(n5901) );
  XOR U6438 ( .A(n5900), .B(n5901), .Z(n5825) );
  AND U6439 ( .A(x[152]), .B(y[679]), .Z(n6180) );
  AND U6440 ( .A(x[153]), .B(y[675]), .Z(n5866) );
  XOR U6441 ( .A(n5867), .B(n5866), .Z(n5865) );
  AND U6442 ( .A(x[129]), .B(y[699]), .Z(n5864) );
  XOR U6443 ( .A(n5865), .B(n5864), .Z(n5931) );
  AND U6444 ( .A(x[144]), .B(y[684]), .Z(n5861) );
  AND U6445 ( .A(x[152]), .B(y[676]), .Z(n5860) );
  XOR U6446 ( .A(n5861), .B(n5860), .Z(n5863) );
  AND U6447 ( .A(x[130]), .B(y[698]), .Z(n5862) );
  XOR U6448 ( .A(n5863), .B(n5862), .Z(n5930) );
  XOR U6449 ( .A(n5931), .B(n5930), .Z(n5933) );
  XOR U6450 ( .A(n5932), .B(n5933), .Z(n5907) );
  AND U6451 ( .A(x[131]), .B(y[697]), .Z(n5886) );
  XOR U6452 ( .A(n5887), .B(n5886), .Z(n5889) );
  AND U6453 ( .A(x[151]), .B(y[677]), .Z(n5888) );
  XOR U6454 ( .A(n5889), .B(n5888), .Z(n5927) );
  AND U6455 ( .A(x[133]), .B(y[695]), .Z(n5876) );
  AND U6456 ( .A(x[149]), .B(y[679]), .Z(n5875) );
  XOR U6457 ( .A(n5876), .B(n5875), .Z(n5878) );
  AND U6458 ( .A(x[148]), .B(y[680]), .Z(n5877) );
  XOR U6459 ( .A(n5878), .B(n5877), .Z(n5926) );
  XOR U6460 ( .A(n5927), .B(n5926), .Z(n5929) );
  XOR U6461 ( .A(n5928), .B(n5929), .Z(n5905) );
  IV U6462 ( .A(n5905), .Z(n5765) );
  XOR U6463 ( .A(n5922), .B(n5923), .Z(n5925) );
  AND U6464 ( .A(n5762), .B(o[59]), .Z(n5847) );
  AND U6465 ( .A(x[128]), .B(y[700]), .Z(n5845) );
  AND U6466 ( .A(x[156]), .B(y[672]), .Z(n5844) );
  XOR U6467 ( .A(n5845), .B(n5844), .Z(n5846) );
  XOR U6468 ( .A(n5847), .B(n5846), .Z(n5857) );
  NAND U6469 ( .A(y[690]), .B(x[138]), .Z(n5763) );
  XNOR U6470 ( .A(n5764), .B(n5763), .Z(n5853) );
  AND U6471 ( .A(x[137]), .B(y[691]), .Z(n5852) );
  XOR U6472 ( .A(n5853), .B(n5852), .Z(n5856) );
  XOR U6473 ( .A(n5857), .B(n5856), .Z(n5859) );
  XOR U6474 ( .A(n5858), .B(n5859), .Z(n5924) );
  XNOR U6475 ( .A(n5925), .B(n5924), .Z(n5904) );
  XOR U6476 ( .A(n5765), .B(n5904), .Z(n5906) );
  XNOR U6477 ( .A(n5827), .B(n5826), .Z(n5820) );
  NAND U6478 ( .A(n5767), .B(n5766), .Z(n5771) );
  NANDN U6479 ( .A(n5769), .B(n5768), .Z(n5770) );
  NAND U6480 ( .A(n5771), .B(n5770), .Z(n5819) );
  NAND U6481 ( .A(n5773), .B(n5772), .Z(n5777) );
  NAND U6482 ( .A(n5775), .B(n5774), .Z(n5776) );
  NAND U6483 ( .A(n5777), .B(n5776), .Z(n5818) );
  XNOR U6484 ( .A(n5819), .B(n5818), .Z(n5821) );
  XNOR U6485 ( .A(n5806), .B(n5807), .Z(n5808) );
  NANDN U6486 ( .A(n5779), .B(n5778), .Z(n5783) );
  NAND U6487 ( .A(n5781), .B(n5780), .Z(n5782) );
  NAND U6488 ( .A(n5783), .B(n5782), .Z(n5814) );
  NAND U6489 ( .A(n5785), .B(n5784), .Z(n5789) );
  NAND U6490 ( .A(n5787), .B(n5786), .Z(n5788) );
  NAND U6491 ( .A(n5789), .B(n5788), .Z(n5812) );
  NAND U6492 ( .A(n5791), .B(n5790), .Z(n5795) );
  NANDN U6493 ( .A(n5793), .B(n5792), .Z(n5794) );
  AND U6494 ( .A(n5795), .B(n5794), .Z(n5813) );
  XNOR U6495 ( .A(n5812), .B(n5813), .Z(n5815) );
  XNOR U6496 ( .A(n5808), .B(n5809), .Z(n5936) );
  XNOR U6497 ( .A(n5937), .B(n5936), .Z(n5942) );
  NANDN U6498 ( .A(n5800), .B(n5799), .Z(n5804) );
  NAND U6499 ( .A(n5802), .B(n5801), .Z(n5803) );
  AND U6500 ( .A(n5804), .B(n5803), .Z(n5941) );
  XOR U6501 ( .A(n5940), .B(n5941), .Z(n5805) );
  XNOR U6502 ( .A(n5942), .B(n5805), .Z(N125) );
  NANDN U6503 ( .A(n5807), .B(n5806), .Z(n5811) );
  NANDN U6504 ( .A(n5809), .B(n5808), .Z(n5810) );
  NAND U6505 ( .A(n5811), .B(n5810), .Z(n5949) );
  NAND U6506 ( .A(n5813), .B(n5812), .Z(n5817) );
  NANDN U6507 ( .A(n5815), .B(n5814), .Z(n5816) );
  NAND U6508 ( .A(n5817), .B(n5816), .Z(n5947) );
  NAND U6509 ( .A(n5819), .B(n5818), .Z(n5823) );
  NANDN U6510 ( .A(n5821), .B(n5820), .Z(n5822) );
  NAND U6511 ( .A(n5823), .B(n5822), .Z(n5953) );
  NANDN U6512 ( .A(n5825), .B(n5824), .Z(n5829) );
  NAND U6513 ( .A(n5827), .B(n5826), .Z(n5828) );
  AND U6514 ( .A(n5829), .B(n5828), .Z(n5954) );
  XOR U6515 ( .A(n5953), .B(n5954), .Z(n5956) );
  NAND U6516 ( .A(n5831), .B(n5830), .Z(n5835) );
  NAND U6517 ( .A(n5833), .B(n5832), .Z(n5834) );
  NAND U6518 ( .A(n5835), .B(n5834), .Z(n5971) );
  NAND U6519 ( .A(n5845), .B(n5844), .Z(n5850) );
  IV U6520 ( .A(n5846), .Z(n5848) );
  NANDN U6521 ( .A(n5848), .B(n5847), .Z(n5849) );
  NAND U6522 ( .A(n5850), .B(n5849), .Z(n6090) );
  XOR U6523 ( .A(n6089), .B(n6090), .Z(n6091) );
  AND U6524 ( .A(x[138]), .B(y[692]), .Z(n6087) );
  NAND U6525 ( .A(n5851), .B(n6087), .Z(n5855) );
  NAND U6526 ( .A(n5853), .B(n5852), .Z(n5854) );
  NAND U6527 ( .A(n5855), .B(n5854), .Z(n6064) );
  AND U6528 ( .A(x[150]), .B(y[679]), .Z(n6041) );
  AND U6529 ( .A(x[140]), .B(y[689]), .Z(n6231) );
  AND U6530 ( .A(x[129]), .B(y[700]), .Z(n6039) );
  XOR U6531 ( .A(n6231), .B(n6039), .Z(n6040) );
  XOR U6532 ( .A(n6041), .B(n6040), .Z(n6063) );
  AND U6533 ( .A(x[143]), .B(y[686]), .Z(n6042) );
  XOR U6534 ( .A(n6063), .B(n6062), .Z(n6065) );
  XNOR U6535 ( .A(n6064), .B(n6065), .Z(n6092) );
  XOR U6536 ( .A(n6091), .B(n6092), .Z(n6059) );
  XNOR U6537 ( .A(n6059), .B(n6058), .Z(n6061) );
  XOR U6538 ( .A(n6060), .B(n6061), .Z(n6056) );
  XOR U6539 ( .A(n6068), .B(n6069), .Z(n6070) );
  AND U6540 ( .A(x[139]), .B(y[690]), .Z(n6017) );
  AND U6541 ( .A(x[131]), .B(y[698]), .Z(n6015) );
  AND U6542 ( .A(x[145]), .B(y[684]), .Z(n6014) );
  XOR U6543 ( .A(n6015), .B(n6014), .Z(n6016) );
  XOR U6544 ( .A(n6017), .B(n6016), .Z(n5986) );
  AND U6545 ( .A(x[151]), .B(y[678]), .Z(n6011) );
  AND U6546 ( .A(x[141]), .B(y[688]), .Z(n6009) );
  AND U6547 ( .A(x[152]), .B(y[677]), .Z(n6211) );
  XOR U6548 ( .A(n6009), .B(n6211), .Z(n6010) );
  XOR U6549 ( .A(n6011), .B(n6010), .Z(n5985) );
  XOR U6550 ( .A(n5986), .B(n5985), .Z(n5987) );
  XNOR U6551 ( .A(n5988), .B(n5987), .Z(n6071) );
  XOR U6552 ( .A(n6070), .B(n6071), .Z(n5979) );
  AND U6553 ( .A(x[153]), .B(y[676]), .Z(n6038) );
  AND U6554 ( .A(x[154]), .B(y[675]), .Z(n6035) );
  XOR U6555 ( .A(n6036), .B(n6035), .Z(n6037) );
  XOR U6556 ( .A(n6038), .B(n6037), .Z(n6073) );
  AND U6557 ( .A(x[156]), .B(y[673]), .Z(n6049) );
  XOR U6558 ( .A(o[61]), .B(n6049), .Z(n6084) );
  AND U6559 ( .A(x[128]), .B(y[701]), .Z(n6082) );
  AND U6560 ( .A(x[157]), .B(y[672]), .Z(n6081) );
  XOR U6561 ( .A(n6082), .B(n6081), .Z(n6083) );
  XOR U6562 ( .A(n6084), .B(n6083), .Z(n6072) );
  XOR U6563 ( .A(n6073), .B(n6072), .Z(n6074) );
  XOR U6564 ( .A(n6075), .B(n6074), .Z(n5977) );
  AND U6565 ( .A(x[130]), .B(y[699]), .Z(n5999) );
  AND U6566 ( .A(o[60]), .B(n5879), .Z(n5992) );
  AND U6567 ( .A(x[144]), .B(y[685]), .Z(n5990) );
  AND U6568 ( .A(x[155]), .B(y[674]), .Z(n5989) );
  XOR U6569 ( .A(n5990), .B(n5989), .Z(n5991) );
  XOR U6570 ( .A(n5992), .B(n5991), .Z(n6027) );
  XOR U6571 ( .A(n6028), .B(n6027), .Z(n6031) );
  XOR U6572 ( .A(n6030), .B(n6031), .Z(n5978) );
  XNOR U6573 ( .A(n5977), .B(n5978), .Z(n5980) );
  XOR U6574 ( .A(n5979), .B(n5980), .Z(n5983) );
  AND U6575 ( .A(x[133]), .B(y[696]), .Z(n5995) );
  AND U6576 ( .A(x[132]), .B(y[697]), .Z(n5994) );
  AND U6577 ( .A(x[138]), .B(y[691]), .Z(n5993) );
  XOR U6578 ( .A(n5994), .B(n5993), .Z(n5996) );
  XOR U6579 ( .A(n5995), .B(n5996), .Z(n6078) );
  AND U6580 ( .A(x[136]), .B(y[693]), .Z(n6022) );
  AND U6581 ( .A(x[134]), .B(y[695]), .Z(n5881) );
  AND U6582 ( .A(y[694]), .B(x[135]), .Z(n5880) );
  XOR U6583 ( .A(n5881), .B(n5880), .Z(n6021) );
  XOR U6584 ( .A(n6022), .B(n6021), .Z(n6076) );
  AND U6585 ( .A(x[137]), .B(y[692]), .Z(n6132) );
  XOR U6586 ( .A(n6076), .B(n6132), .Z(n6077) );
  XOR U6587 ( .A(n6078), .B(n6077), .Z(n6007) );
  XNOR U6588 ( .A(n6005), .B(n6006), .Z(n6008) );
  XOR U6589 ( .A(n6007), .B(n6008), .Z(n5981) );
  XNOR U6590 ( .A(n5981), .B(n5982), .Z(n5984) );
  XOR U6591 ( .A(n5983), .B(n5984), .Z(n6054) );
  XOR U6592 ( .A(n6054), .B(n6055), .Z(n6057) );
  XOR U6593 ( .A(n6056), .B(n6057), .Z(n5972) );
  XOR U6594 ( .A(n5971), .B(n5972), .Z(n5974) );
  NAND U6595 ( .A(n5899), .B(n5898), .Z(n5903) );
  NAND U6596 ( .A(n5901), .B(n5900), .Z(n5902) );
  NAND U6597 ( .A(n5903), .B(n5902), .Z(n5965) );
  NANDN U6598 ( .A(n5905), .B(n5904), .Z(n5909) );
  NANDN U6599 ( .A(n5907), .B(n5906), .Z(n5908) );
  AND U6600 ( .A(n5909), .B(n5908), .Z(n5966) );
  XOR U6601 ( .A(n5965), .B(n5966), .Z(n5967) );
  NAND U6602 ( .A(n5911), .B(n5910), .Z(n5915) );
  NAND U6603 ( .A(n5913), .B(n5912), .Z(n5914) );
  NAND U6604 ( .A(n5915), .B(n5914), .Z(n5961) );
  NANDN U6605 ( .A(n5917), .B(n5916), .Z(n5921) );
  NAND U6606 ( .A(n5919), .B(n5918), .Z(n5920) );
  NAND U6607 ( .A(n5921), .B(n5920), .Z(n5959) );
  XNOR U6608 ( .A(n6050), .B(n6051), .Z(n6053) );
  XOR U6609 ( .A(n6052), .B(n6053), .Z(n5960) );
  XOR U6610 ( .A(n5961), .B(n5962), .Z(n5968) );
  XNOR U6611 ( .A(n5967), .B(n5968), .Z(n5973) );
  XOR U6612 ( .A(n5974), .B(n5973), .Z(n5955) );
  XOR U6613 ( .A(n5956), .B(n5955), .Z(n5948) );
  XOR U6614 ( .A(n5947), .B(n5948), .Z(n5950) );
  XOR U6615 ( .A(n5949), .B(n5950), .Z(n5946) );
  NAND U6616 ( .A(n5935), .B(n5934), .Z(n5939) );
  NAND U6617 ( .A(n5937), .B(n5936), .Z(n5938) );
  AND U6618 ( .A(n5939), .B(n5938), .Z(n5945) );
  XNOR U6619 ( .A(n5945), .B(n5944), .Z(n5943) );
  XNOR U6620 ( .A(n5946), .B(n5943), .Z(N126) );
  NAND U6621 ( .A(n5948), .B(n5947), .Z(n5952) );
  NAND U6622 ( .A(n5950), .B(n5949), .Z(n5951) );
  NAND U6623 ( .A(n5952), .B(n5951), .Z(n6357) );
  NAND U6624 ( .A(n5954), .B(n5953), .Z(n5958) );
  NAND U6625 ( .A(n5956), .B(n5955), .Z(n5957) );
  NAND U6626 ( .A(n5958), .B(n5957), .Z(n6362) );
  NANDN U6627 ( .A(n5960), .B(n5959), .Z(n5964) );
  NANDN U6628 ( .A(n5962), .B(n5961), .Z(n5963) );
  AND U6629 ( .A(n5964), .B(n5963), .Z(n6369) );
  NAND U6630 ( .A(n5966), .B(n5965), .Z(n5970) );
  NANDN U6631 ( .A(n5968), .B(n5967), .Z(n5969) );
  AND U6632 ( .A(n5970), .B(n5969), .Z(n6371) );
  NAND U6633 ( .A(n5972), .B(n5971), .Z(n5976) );
  NAND U6634 ( .A(n5974), .B(n5973), .Z(n5975) );
  AND U6635 ( .A(n5976), .B(n5975), .Z(n6370) );
  XOR U6636 ( .A(n6371), .B(n6370), .Z(n6368) );
  XOR U6637 ( .A(n6369), .B(n6368), .Z(n6365) );
  NAND U6638 ( .A(n5994), .B(n5993), .Z(n5998) );
  NAND U6639 ( .A(n5996), .B(n5995), .Z(n5997) );
  NAND U6640 ( .A(n5998), .B(n5997), .Z(n6109) );
  AND U6641 ( .A(x[134]), .B(y[696]), .Z(n6142) );
  AND U6642 ( .A(x[133]), .B(y[697]), .Z(n6144) );
  AND U6643 ( .A(x[147]), .B(y[683]), .Z(n6143) );
  XOR U6644 ( .A(n6144), .B(n6143), .Z(n6141) );
  XNOR U6645 ( .A(n6142), .B(n6141), .Z(n6112) );
  AND U6646 ( .A(x[132]), .B(y[698]), .Z(n6225) );
  AND U6647 ( .A(x[131]), .B(y[699]), .Z(n6227) );
  AND U6648 ( .A(x[146]), .B(y[684]), .Z(n6226) );
  XOR U6649 ( .A(n6227), .B(n6226), .Z(n6224) );
  XOR U6650 ( .A(n6225), .B(n6224), .Z(n6115) );
  NANDN U6651 ( .A(n6000), .B(n5999), .Z(n6004) );
  NANDN U6652 ( .A(n6002), .B(n6001), .Z(n6003) );
  AND U6653 ( .A(n6004), .B(n6003), .Z(n6114) );
  XOR U6654 ( .A(n6112), .B(n6113), .Z(n6108) );
  XOR U6655 ( .A(n6109), .B(n6108), .Z(n6107) );
  XOR U6656 ( .A(n6106), .B(n6107), .Z(n6097) );
  XOR U6657 ( .A(n6094), .B(n6093), .Z(n6336) );
  NAND U6658 ( .A(n6009), .B(n6211), .Z(n6013) );
  NAND U6659 ( .A(n6011), .B(n6010), .Z(n6012) );
  NAND U6660 ( .A(n6013), .B(n6012), .Z(n6103) );
  NAND U6661 ( .A(n6015), .B(n6014), .Z(n6019) );
  NAND U6662 ( .A(n6017), .B(n6016), .Z(n6018) );
  AND U6663 ( .A(n6019), .B(n6018), .Z(n6251) );
  AND U6664 ( .A(x[128]), .B(y[702]), .Z(n6150) );
  AND U6665 ( .A(x[157]), .B(y[673]), .Z(n6195) );
  XOR U6666 ( .A(o[62]), .B(n6195), .Z(n6152) );
  AND U6667 ( .A(x[158]), .B(y[672]), .Z(n6151) );
  XOR U6668 ( .A(n6152), .B(n6151), .Z(n6149) );
  XOR U6669 ( .A(n6150), .B(n6149), .Z(n6253) );
  AND U6670 ( .A(x[148]), .B(y[682]), .Z(n6268) );
  XOR U6671 ( .A(n6269), .B(n6268), .Z(n6267) );
  AND U6672 ( .A(x[136]), .B(y[694]), .Z(n6266) );
  XNOR U6673 ( .A(n6267), .B(n6266), .Z(n6252) );
  XNOR U6674 ( .A(n6251), .B(n6250), .Z(n6102) );
  XOR U6675 ( .A(n6103), .B(n6102), .Z(n6100) );
  AND U6676 ( .A(x[135]), .B(y[695]), .Z(n6281) );
  NAND U6677 ( .A(n6020), .B(n6281), .Z(n6024) );
  NAND U6678 ( .A(n6022), .B(n6021), .Z(n6023) );
  AND U6679 ( .A(n6024), .B(n6023), .Z(n6122) );
  AND U6680 ( .A(y[681]), .B(x[149]), .Z(n6026) );
  AND U6681 ( .A(y[680]), .B(x[150]), .Z(n6025) );
  XOR U6682 ( .A(n6026), .B(n6025), .Z(n6280) );
  XOR U6683 ( .A(n6281), .B(n6280), .Z(n6125) );
  AND U6684 ( .A(x[145]), .B(y[685]), .Z(n6275) );
  AND U6685 ( .A(x[130]), .B(y[700]), .Z(n6277) );
  AND U6686 ( .A(x[154]), .B(y[676]), .Z(n6276) );
  XOR U6687 ( .A(n6277), .B(n6276), .Z(n6274) );
  XNOR U6688 ( .A(n6275), .B(n6274), .Z(n6124) );
  XNOR U6689 ( .A(n6122), .B(n6123), .Z(n6101) );
  XNOR U6690 ( .A(n6100), .B(n6101), .Z(n6318) );
  IV U6691 ( .A(n6027), .Z(n6029) );
  NANDN U6692 ( .A(n6029), .B(n6028), .Z(n6034) );
  IV U6693 ( .A(n6030), .Z(n6032) );
  NANDN U6694 ( .A(n6032), .B(n6031), .Z(n6033) );
  NAND U6695 ( .A(n6034), .B(n6033), .Z(n6317) );
  XOR U6696 ( .A(n6318), .B(n6317), .Z(n6316) );
  NANDN U6697 ( .A(n6283), .B(n6042), .Z(n6046) );
  NANDN U6698 ( .A(n6044), .B(n6043), .Z(n6045) );
  AND U6699 ( .A(n6046), .B(n6045), .Z(n6245) );
  AND U6700 ( .A(x[151]), .B(y[679]), .Z(n6209) );
  AND U6701 ( .A(y[678]), .B(x[152]), .Z(n6048) );
  AND U6702 ( .A(y[677]), .B(x[153]), .Z(n6047) );
  XOR U6703 ( .A(n6048), .B(n6047), .Z(n6208) );
  XOR U6704 ( .A(n6209), .B(n6208), .Z(n6247) );
  AND U6705 ( .A(n6049), .B(o[61]), .Z(n6136) );
  AND U6706 ( .A(x[156]), .B(y[674]), .Z(n6138) );
  AND U6707 ( .A(x[144]), .B(y[686]), .Z(n6137) );
  XOR U6708 ( .A(n6138), .B(n6137), .Z(n6135) );
  XNOR U6709 ( .A(n6136), .B(n6135), .Z(n6246) );
  XNOR U6710 ( .A(n6245), .B(n6244), .Z(n6128) );
  XOR U6711 ( .A(n6129), .B(n6128), .Z(n6127) );
  XOR U6712 ( .A(n6126), .B(n6127), .Z(n6315) );
  XOR U6713 ( .A(n6316), .B(n6315), .Z(n6335) );
  XNOR U6714 ( .A(n6333), .B(n6334), .Z(n6348) );
  NAND U6715 ( .A(n6063), .B(n6062), .Z(n6067) );
  NAND U6716 ( .A(n6065), .B(n6064), .Z(n6066) );
  AND U6717 ( .A(n6067), .B(n6066), .Z(n6302) );
  XOR U6718 ( .A(n6302), .B(n6301), .Z(n6300) );
  XOR U6719 ( .A(n6300), .B(n6299), .Z(n6312) );
  NAND U6720 ( .A(n6076), .B(n6132), .Z(n6080) );
  NAND U6721 ( .A(n6078), .B(n6077), .Z(n6079) );
  AND U6722 ( .A(n6080), .B(n6079), .Z(n6295) );
  AND U6723 ( .A(y[690]), .B(x[140]), .Z(n6085) );
  XOR U6724 ( .A(n6086), .B(n6085), .Z(n6232) );
  XOR U6725 ( .A(n6233), .B(n6232), .Z(n6131) );
  AND U6726 ( .A(y[693]), .B(x[137]), .Z(n6088) );
  XOR U6727 ( .A(n6088), .B(n6087), .Z(n6130) );
  XOR U6728 ( .A(n6131), .B(n6130), .Z(n6121) );
  AND U6729 ( .A(x[155]), .B(y[675]), .Z(n6263) );
  AND U6730 ( .A(x[129]), .B(y[701]), .Z(n6262) );
  XOR U6731 ( .A(n6263), .B(n6262), .Z(n6260) );
  XOR U6732 ( .A(n6261), .B(n6260), .Z(n6120) );
  XOR U6733 ( .A(n6121), .B(n6120), .Z(n6119) );
  XOR U6734 ( .A(n6118), .B(n6119), .Z(n6296) );
  XNOR U6735 ( .A(n6293), .B(n6294), .Z(n6311) );
  XNOR U6736 ( .A(n6309), .B(n6310), .Z(n6330) );
  XOR U6737 ( .A(n6329), .B(n6330), .Z(n6327) );
  XOR U6738 ( .A(n6328), .B(n6327), .Z(n6364) );
  XOR U6739 ( .A(n6362), .B(n6363), .Z(n6354) );
  XNOR U6740 ( .A(n6355), .B(n6354), .Z(N127) );
  IV U6741 ( .A(n6093), .Z(n6095) );
  NANDN U6742 ( .A(n6095), .B(n6094), .Z(n6099) );
  NANDN U6743 ( .A(n6097), .B(n6096), .Z(n6098) );
  AND U6744 ( .A(n6099), .B(n6098), .Z(n6344) );
  NANDN U6745 ( .A(n6101), .B(n6100), .Z(n6105) );
  NAND U6746 ( .A(n6103), .B(n6102), .Z(n6104) );
  AND U6747 ( .A(n6105), .B(n6104), .Z(n6326) );
  NAND U6748 ( .A(n6107), .B(n6106), .Z(n6111) );
  NAND U6749 ( .A(n6109), .B(n6108), .Z(n6110) );
  AND U6750 ( .A(n6111), .B(n6110), .Z(n6308) );
  NANDN U6751 ( .A(n6113), .B(n6112), .Z(n6117) );
  NANDN U6752 ( .A(n6115), .B(n6114), .Z(n6116) );
  AND U6753 ( .A(n6117), .B(n6116), .Z(n6292) );
  NAND U6754 ( .A(n6131), .B(n6130), .Z(n6134) );
  AND U6755 ( .A(x[138]), .B(y[693]), .Z(n6169) );
  NAND U6756 ( .A(n6132), .B(n6169), .Z(n6133) );
  NAND U6757 ( .A(n6136), .B(n6135), .Z(n6140) );
  NAND U6758 ( .A(n6138), .B(n6137), .Z(n6139) );
  AND U6759 ( .A(n6140), .B(n6139), .Z(n6148) );
  NAND U6760 ( .A(n6142), .B(n6141), .Z(n6146) );
  NAND U6761 ( .A(n6144), .B(n6143), .Z(n6145) );
  NAND U6762 ( .A(n6146), .B(n6145), .Z(n6147) );
  XNOR U6763 ( .A(n6148), .B(n6147), .Z(n6205) );
  NAND U6764 ( .A(n6150), .B(n6149), .Z(n6154) );
  NAND U6765 ( .A(n6152), .B(n6151), .Z(n6153) );
  AND U6766 ( .A(n6154), .B(n6153), .Z(n6203) );
  AND U6767 ( .A(y[694]), .B(x[137]), .Z(n6156) );
  NAND U6768 ( .A(y[677]), .B(x[154]), .Z(n6155) );
  XNOR U6769 ( .A(n6156), .B(n6155), .Z(n6160) );
  AND U6770 ( .A(y[680]), .B(x[151]), .Z(n6158) );
  NAND U6771 ( .A(y[696]), .B(x[135]), .Z(n6157) );
  XNOR U6772 ( .A(n6158), .B(n6157), .Z(n6159) );
  XOR U6773 ( .A(n6160), .B(n6159), .Z(n6168) );
  AND U6774 ( .A(y[673]), .B(x[158]), .Z(n6162) );
  NAND U6775 ( .A(y[674]), .B(x[157]), .Z(n6161) );
  XNOR U6776 ( .A(n6162), .B(n6161), .Z(n6166) );
  AND U6777 ( .A(y[689]), .B(x[142]), .Z(n6164) );
  NAND U6778 ( .A(y[691]), .B(x[140]), .Z(n6163) );
  XNOR U6779 ( .A(n6164), .B(n6163), .Z(n6165) );
  XNOR U6780 ( .A(n6166), .B(n6165), .Z(n6167) );
  XNOR U6781 ( .A(n6168), .B(n6167), .Z(n6201) );
  XOR U6782 ( .A(n6169), .B(o[63]), .Z(n6171) );
  AND U6783 ( .A(x[150]), .B(y[681]), .Z(n6282) );
  XNOR U6784 ( .A(n6282), .B(n6230), .Z(n6170) );
  XNOR U6785 ( .A(n6171), .B(n6170), .Z(n6194) );
  AND U6786 ( .A(y[684]), .B(x[147]), .Z(n6173) );
  NAND U6787 ( .A(y[695]), .B(x[136]), .Z(n6172) );
  XNOR U6788 ( .A(n6173), .B(n6172), .Z(n6184) );
  AND U6789 ( .A(y[682]), .B(x[149]), .Z(n6175) );
  NAND U6790 ( .A(y[687]), .B(x[144]), .Z(n6174) );
  XNOR U6791 ( .A(n6175), .B(n6174), .Z(n6179) );
  AND U6792 ( .A(y[702]), .B(x[129]), .Z(n6177) );
  NAND U6793 ( .A(y[692]), .B(x[139]), .Z(n6176) );
  XNOR U6794 ( .A(n6177), .B(n6176), .Z(n6178) );
  XOR U6795 ( .A(n6179), .B(n6178), .Z(n6182) );
  AND U6796 ( .A(x[153]), .B(y[678]), .Z(n6210) );
  XNOR U6797 ( .A(n6180), .B(n6210), .Z(n6181) );
  XNOR U6798 ( .A(n6182), .B(n6181), .Z(n6183) );
  XOR U6799 ( .A(n6184), .B(n6183), .Z(n6192) );
  AND U6800 ( .A(y[675]), .B(x[156]), .Z(n6186) );
  NAND U6801 ( .A(y[703]), .B(x[128]), .Z(n6185) );
  XNOR U6802 ( .A(n6186), .B(n6185), .Z(n6190) );
  AND U6803 ( .A(y[672]), .B(x[159]), .Z(n6188) );
  NAND U6804 ( .A(y[683]), .B(x[148]), .Z(n6187) );
  XNOR U6805 ( .A(n6188), .B(n6187), .Z(n6189) );
  XNOR U6806 ( .A(n6190), .B(n6189), .Z(n6191) );
  XNOR U6807 ( .A(n6192), .B(n6191), .Z(n6193) );
  XOR U6808 ( .A(n6194), .B(n6193), .Z(n6199) );
  AND U6809 ( .A(n6195), .B(o[62]), .Z(n6197) );
  XNOR U6810 ( .A(n6197), .B(n6196), .Z(n6198) );
  XNOR U6811 ( .A(n6199), .B(n6198), .Z(n6200) );
  XNOR U6812 ( .A(n6201), .B(n6200), .Z(n6202) );
  XNOR U6813 ( .A(n6203), .B(n6202), .Z(n6204) );
  AND U6814 ( .A(y[701]), .B(x[130]), .Z(n6207) );
  NAND U6815 ( .A(y[686]), .B(x[145]), .Z(n6206) );
  XNOR U6816 ( .A(n6207), .B(n6206), .Z(n6223) );
  NAND U6817 ( .A(n6209), .B(n6208), .Z(n6213) );
  NAND U6818 ( .A(n6211), .B(n6210), .Z(n6212) );
  AND U6819 ( .A(n6213), .B(n6212), .Z(n6221) );
  AND U6820 ( .A(y[699]), .B(x[132]), .Z(n6215) );
  NAND U6821 ( .A(y[676]), .B(x[155]), .Z(n6214) );
  XNOR U6822 ( .A(n6215), .B(n6214), .Z(n6219) );
  AND U6823 ( .A(y[698]), .B(x[133]), .Z(n6217) );
  NAND U6824 ( .A(y[697]), .B(x[134]), .Z(n6216) );
  XNOR U6825 ( .A(n6217), .B(n6216), .Z(n6218) );
  XNOR U6826 ( .A(n6219), .B(n6218), .Z(n6220) );
  XNOR U6827 ( .A(n6221), .B(n6220), .Z(n6222) );
  XOR U6828 ( .A(n6223), .B(n6222), .Z(n6243) );
  NAND U6829 ( .A(n6225), .B(n6224), .Z(n6229) );
  NAND U6830 ( .A(n6227), .B(n6226), .Z(n6228) );
  AND U6831 ( .A(n6229), .B(n6228), .Z(n6237) );
  NAND U6832 ( .A(n6231), .B(n6230), .Z(n6235) );
  NAND U6833 ( .A(n6233), .B(n6232), .Z(n6234) );
  AND U6834 ( .A(n6235), .B(n6234), .Z(n6236) );
  XNOR U6835 ( .A(n6237), .B(n6236), .Z(n6241) );
  AND U6836 ( .A(y[700]), .B(x[131]), .Z(n6239) );
  NAND U6837 ( .A(y[685]), .B(x[146]), .Z(n6238) );
  XNOR U6838 ( .A(n6239), .B(n6238), .Z(n6240) );
  XOR U6839 ( .A(n6241), .B(n6240), .Z(n6242) );
  XNOR U6840 ( .A(n6243), .B(n6242), .Z(n6259) );
  NAND U6841 ( .A(n6245), .B(n6244), .Z(n6249) );
  NANDN U6842 ( .A(n6247), .B(n6246), .Z(n6248) );
  AND U6843 ( .A(n6249), .B(n6248), .Z(n6257) );
  NAND U6844 ( .A(n6251), .B(n6250), .Z(n6255) );
  NANDN U6845 ( .A(n6253), .B(n6252), .Z(n6254) );
  NAND U6846 ( .A(n6255), .B(n6254), .Z(n6256) );
  XNOR U6847 ( .A(n6257), .B(n6256), .Z(n6258) );
  NAND U6848 ( .A(n6261), .B(n6260), .Z(n6265) );
  NAND U6849 ( .A(n6263), .B(n6262), .Z(n6264) );
  AND U6850 ( .A(n6265), .B(n6264), .Z(n6273) );
  NAND U6851 ( .A(n6267), .B(n6266), .Z(n6271) );
  NAND U6852 ( .A(n6269), .B(n6268), .Z(n6270) );
  NAND U6853 ( .A(n6271), .B(n6270), .Z(n6272) );
  XNOR U6854 ( .A(n6273), .B(n6272), .Z(n6289) );
  NAND U6855 ( .A(n6275), .B(n6274), .Z(n6279) );
  NAND U6856 ( .A(n6277), .B(n6276), .Z(n6278) );
  AND U6857 ( .A(n6279), .B(n6278), .Z(n6287) );
  NAND U6858 ( .A(n6281), .B(n6280), .Z(n6285) );
  NANDN U6859 ( .A(n6283), .B(n6282), .Z(n6284) );
  NAND U6860 ( .A(n6285), .B(n6284), .Z(n6286) );
  XNOR U6861 ( .A(n6287), .B(n6286), .Z(n6288) );
  XNOR U6862 ( .A(n6289), .B(n6288), .Z(n6290) );
  XNOR U6863 ( .A(n6292), .B(n6291), .Z(n6306) );
  NAND U6864 ( .A(n6294), .B(n6293), .Z(n6298) );
  NANDN U6865 ( .A(n6296), .B(n6295), .Z(n6297) );
  AND U6866 ( .A(n6298), .B(n6297), .Z(n6304) );
  XNOR U6867 ( .A(n6304), .B(n6303), .Z(n6305) );
  XNOR U6868 ( .A(n6306), .B(n6305), .Z(n6307) );
  XNOR U6869 ( .A(n6308), .B(n6307), .Z(n6324) );
  NANDN U6870 ( .A(n6310), .B(n6309), .Z(n6314) );
  NANDN U6871 ( .A(n6312), .B(n6311), .Z(n6313) );
  AND U6872 ( .A(n6314), .B(n6313), .Z(n6322) );
  NAND U6873 ( .A(n6316), .B(n6315), .Z(n6320) );
  NAND U6874 ( .A(n6318), .B(n6317), .Z(n6319) );
  NAND U6875 ( .A(n6320), .B(n6319), .Z(n6321) );
  XNOR U6876 ( .A(n6322), .B(n6321), .Z(n6323) );
  XNOR U6877 ( .A(n6324), .B(n6323), .Z(n6325) );
  XNOR U6878 ( .A(n6326), .B(n6325), .Z(n6342) );
  NAND U6879 ( .A(n6328), .B(n6327), .Z(n6332) );
  NAND U6880 ( .A(n6330), .B(n6329), .Z(n6331) );
  AND U6881 ( .A(n6332), .B(n6331), .Z(n6340) );
  NANDN U6882 ( .A(n6334), .B(n6333), .Z(n6338) );
  NANDN U6883 ( .A(n6336), .B(n6335), .Z(n6337) );
  NAND U6884 ( .A(n6338), .B(n6337), .Z(n6339) );
  XNOR U6885 ( .A(n6340), .B(n6339), .Z(n6341) );
  XNOR U6886 ( .A(n6342), .B(n6341), .Z(n6343) );
  XNOR U6887 ( .A(n6344), .B(n6343), .Z(n6353) );
  IV U6888 ( .A(n6346), .Z(n6345) );
  OR U6889 ( .A(n6347), .B(n6345), .Z(n6351) );
  ANDN U6890 ( .B(n6347), .A(n6346), .Z(n6349) );
  NANDN U6891 ( .A(n6349), .B(n6348), .Z(n6350) );
  NAND U6892 ( .A(n6351), .B(n6350), .Z(n6352) );
  XNOR U6893 ( .A(n6353), .B(n6352), .Z(n6361) );
  NAND U6894 ( .A(n6355), .B(n6354), .Z(n6359) );
  NANDN U6895 ( .A(n6357), .B(n6356), .Z(n6358) );
  NAND U6896 ( .A(n6359), .B(n6358), .Z(n6360) );
  XNOR U6897 ( .A(n6361), .B(n6360), .Z(n6377) );
  NANDN U6898 ( .A(n6363), .B(n6362), .Z(n6367) );
  NANDN U6899 ( .A(n6365), .B(n6364), .Z(n6366) );
  AND U6900 ( .A(n6367), .B(n6366), .Z(n6375) );
  NAND U6901 ( .A(n6369), .B(n6368), .Z(n6373) );
  NAND U6902 ( .A(n6371), .B(n6370), .Z(n6372) );
  NAND U6903 ( .A(n6373), .B(n6372), .Z(n6374) );
  XNOR U6904 ( .A(n6375), .B(n6374), .Z(n6376) );
  XNOR U6905 ( .A(n6377), .B(n6376), .Z(N128) );
  AND U6906 ( .A(x[128]), .B(y[704]), .Z(n7019) );
  XOR U6907 ( .A(n7019), .B(o[64]), .Z(N161) );
  NAND U6908 ( .A(x[129]), .B(y[704]), .Z(n6387) );
  AND U6909 ( .A(x[128]), .B(y[705]), .Z(n6383) );
  XNOR U6910 ( .A(n6383), .B(o[65]), .Z(n6378) );
  XOR U6911 ( .A(n6387), .B(n6378), .Z(n6380) );
  NAND U6912 ( .A(n7019), .B(o[64]), .Z(n6379) );
  XNOR U6913 ( .A(n6380), .B(n6379), .Z(N162) );
  AND U6914 ( .A(x[128]), .B(y[706]), .Z(n6386) );
  XNOR U6915 ( .A(n6386), .B(o[66]), .Z(n6392) );
  XNOR U6916 ( .A(n6393), .B(n6392), .Z(n6395) );
  AND U6917 ( .A(y[705]), .B(x[129]), .Z(n6382) );
  NAND U6918 ( .A(y[704]), .B(x[130]), .Z(n6381) );
  XNOR U6919 ( .A(n6382), .B(n6381), .Z(n6389) );
  AND U6920 ( .A(n6383), .B(o[65]), .Z(n6388) );
  XNOR U6921 ( .A(n6389), .B(n6388), .Z(n6394) );
  XNOR U6922 ( .A(n6395), .B(n6394), .Z(N163) );
  AND U6923 ( .A(x[129]), .B(y[706]), .Z(n6506) );
  AND U6924 ( .A(x[130]), .B(y[705]), .Z(n6405) );
  XOR U6925 ( .A(n6405), .B(o[67]), .Z(n6410) );
  XOR U6926 ( .A(n6506), .B(n6410), .Z(n6412) );
  AND U6927 ( .A(y[707]), .B(x[128]), .Z(n6385) );
  NAND U6928 ( .A(y[704]), .B(x[131]), .Z(n6384) );
  XNOR U6929 ( .A(n6385), .B(n6384), .Z(n6399) );
  NAND U6930 ( .A(n6386), .B(o[66]), .Z(n6400) );
  XNOR U6931 ( .A(n6399), .B(n6400), .Z(n6411) );
  XNOR U6932 ( .A(n6412), .B(n6411), .Z(n6409) );
  NANDN U6933 ( .A(n6387), .B(n6405), .Z(n6391) );
  NAND U6934 ( .A(n6389), .B(n6388), .Z(n6390) );
  NAND U6935 ( .A(n6391), .B(n6390), .Z(n6407) );
  NANDN U6936 ( .A(n6393), .B(n6392), .Z(n6397) );
  NAND U6937 ( .A(n6395), .B(n6394), .Z(n6396) );
  AND U6938 ( .A(n6397), .B(n6396), .Z(n6408) );
  XOR U6939 ( .A(n6407), .B(n6408), .Z(n6398) );
  XNOR U6940 ( .A(n6409), .B(n6398), .Z(N164) );
  AND U6941 ( .A(x[131]), .B(y[707]), .Z(n6463) );
  NAND U6942 ( .A(n7019), .B(n6463), .Z(n6402) );
  NANDN U6943 ( .A(n6400), .B(n6399), .Z(n6401) );
  AND U6944 ( .A(n6402), .B(n6401), .Z(n6432) );
  AND U6945 ( .A(y[708]), .B(x[128]), .Z(n6404) );
  NAND U6946 ( .A(y[704]), .B(x[132]), .Z(n6403) );
  XNOR U6947 ( .A(n6404), .B(n6403), .Z(n6426) );
  AND U6948 ( .A(n6405), .B(o[67]), .Z(n6425) );
  XOR U6949 ( .A(n6426), .B(n6425), .Z(n6430) );
  AND U6950 ( .A(y[707]), .B(x[129]), .Z(n6611) );
  NAND U6951 ( .A(y[706]), .B(x[130]), .Z(n6406) );
  XNOR U6952 ( .A(n6611), .B(n6406), .Z(n6422) );
  AND U6953 ( .A(x[131]), .B(y[705]), .Z(n6417) );
  XOR U6954 ( .A(n6417), .B(o[68]), .Z(n6421) );
  XOR U6955 ( .A(n6422), .B(n6421), .Z(n6429) );
  XOR U6956 ( .A(n6430), .B(n6429), .Z(n6431) );
  XNOR U6957 ( .A(n6432), .B(n6431), .Z(n6436) );
  NAND U6958 ( .A(n6506), .B(n6410), .Z(n6414) );
  NAND U6959 ( .A(n6412), .B(n6411), .Z(n6413) );
  NAND U6960 ( .A(n6414), .B(n6413), .Z(n6433) );
  XNOR U6961 ( .A(n6434), .B(n6433), .Z(n6435) );
  XOR U6962 ( .A(n6436), .B(n6435), .Z(N165) );
  AND U6963 ( .A(y[709]), .B(x[128]), .Z(n6416) );
  NAND U6964 ( .A(y[704]), .B(x[133]), .Z(n6415) );
  XNOR U6965 ( .A(n6416), .B(n6415), .Z(n6455) );
  NAND U6966 ( .A(n6417), .B(o[68]), .Z(n6456) );
  XNOR U6967 ( .A(n6455), .B(n6456), .Z(n6454) );
  NAND U6968 ( .A(x[130]), .B(y[707]), .Z(n6514) );
  AND U6969 ( .A(y[708]), .B(x[129]), .Z(n6419) );
  NAND U6970 ( .A(y[706]), .B(x[131]), .Z(n6418) );
  XNOR U6971 ( .A(n6419), .B(n6418), .Z(n6450) );
  AND U6972 ( .A(x[132]), .B(y[705]), .Z(n6461) );
  XOR U6973 ( .A(n6461), .B(o[69]), .Z(n6449) );
  XOR U6974 ( .A(n6450), .B(n6449), .Z(n6453) );
  XOR U6975 ( .A(n6514), .B(n6453), .Z(n6420) );
  XNOR U6976 ( .A(n6454), .B(n6420), .Z(n6442) );
  NANDN U6977 ( .A(n6514), .B(n6506), .Z(n6424) );
  NAND U6978 ( .A(n6422), .B(n6421), .Z(n6423) );
  NAND U6979 ( .A(n6424), .B(n6423), .Z(n6441) );
  AND U6980 ( .A(x[132]), .B(y[708]), .Z(n7240) );
  NAND U6981 ( .A(n7240), .B(n7019), .Z(n6428) );
  NAND U6982 ( .A(n6426), .B(n6425), .Z(n6427) );
  NAND U6983 ( .A(n6428), .B(n6427), .Z(n6440) );
  XNOR U6984 ( .A(n6441), .B(n6440), .Z(n6443) );
  NANDN U6985 ( .A(n6434), .B(n6433), .Z(n6438) );
  NAND U6986 ( .A(n6436), .B(n6435), .Z(n6437) );
  AND U6987 ( .A(n6438), .B(n6437), .Z(n6446) );
  XOR U6988 ( .A(n6447), .B(n6446), .Z(n6439) );
  XNOR U6989 ( .A(n6448), .B(n6439), .Z(N166) );
  NAND U6990 ( .A(n6441), .B(n6440), .Z(n6445) );
  NANDN U6991 ( .A(n6443), .B(n6442), .Z(n6444) );
  AND U6992 ( .A(n6445), .B(n6444), .Z(n6496) );
  AND U6993 ( .A(x[131]), .B(y[708]), .Z(n6515) );
  NAND U6994 ( .A(n6515), .B(n6506), .Z(n6452) );
  NAND U6995 ( .A(n6450), .B(n6449), .Z(n6451) );
  AND U6996 ( .A(n6452), .B(n6451), .Z(n6491) );
  XNOR U6997 ( .A(n6491), .B(n6490), .Z(n6493) );
  AND U6998 ( .A(x[133]), .B(y[709]), .Z(n6687) );
  NAND U6999 ( .A(n7019), .B(n6687), .Z(n6458) );
  NANDN U7000 ( .A(n6456), .B(n6455), .Z(n6457) );
  AND U7001 ( .A(n6458), .B(n6457), .Z(n6467) );
  AND U7002 ( .A(y[710]), .B(x[128]), .Z(n6460) );
  NAND U7003 ( .A(y[704]), .B(x[134]), .Z(n6459) );
  XNOR U7004 ( .A(n6460), .B(n6459), .Z(n6473) );
  NAND U7005 ( .A(n6461), .B(o[69]), .Z(n6474) );
  XNOR U7006 ( .A(n6473), .B(n6474), .Z(n6466) );
  XNOR U7007 ( .A(n6467), .B(n6466), .Z(n6469) );
  NAND U7008 ( .A(y[708]), .B(x[130]), .Z(n6462) );
  XNOR U7009 ( .A(n6463), .B(n6462), .Z(n6478) );
  AND U7010 ( .A(y[709]), .B(x[129]), .Z(n6723) );
  NAND U7011 ( .A(y[706]), .B(x[132]), .Z(n6464) );
  XNOR U7012 ( .A(n6723), .B(n6464), .Z(n6482) );
  NAND U7013 ( .A(x[133]), .B(y[705]), .Z(n6489) );
  XNOR U7014 ( .A(o[70]), .B(n6489), .Z(n6481) );
  XOR U7015 ( .A(n6482), .B(n6481), .Z(n6477) );
  XOR U7016 ( .A(n6478), .B(n6477), .Z(n6468) );
  XOR U7017 ( .A(n6469), .B(n6468), .Z(n6492) );
  XOR U7018 ( .A(n6493), .B(n6492), .Z(n6498) );
  XNOR U7019 ( .A(n6497), .B(n6498), .Z(n6465) );
  XOR U7020 ( .A(n6496), .B(n6465), .Z(N167) );
  NANDN U7021 ( .A(n6467), .B(n6466), .Z(n6471) );
  NAND U7022 ( .A(n6469), .B(n6468), .Z(n6470) );
  AND U7023 ( .A(n6471), .B(n6470), .Z(n6538) );
  AND U7024 ( .A(y[706]), .B(x[133]), .Z(n6599) );
  NAND U7025 ( .A(y[710]), .B(x[129]), .Z(n6472) );
  XNOR U7026 ( .A(n6599), .B(n6472), .Z(n6508) );
  NAND U7027 ( .A(x[134]), .B(y[705]), .Z(n6511) );
  XNOR U7028 ( .A(o[71]), .B(n6511), .Z(n6507) );
  XOR U7029 ( .A(n6508), .B(n6507), .Z(n6527) );
  AND U7030 ( .A(x[134]), .B(y[710]), .Z(n6563) );
  NAND U7031 ( .A(n7019), .B(n6563), .Z(n6476) );
  NANDN U7032 ( .A(n6474), .B(n6473), .Z(n6475) );
  AND U7033 ( .A(n6476), .B(n6475), .Z(n6526) );
  NANDN U7034 ( .A(n6514), .B(n6515), .Z(n6480) );
  NAND U7035 ( .A(n6478), .B(n6477), .Z(n6479) );
  NAND U7036 ( .A(n6480), .B(n6479), .Z(n6529) );
  AND U7037 ( .A(x[132]), .B(y[709]), .Z(n7024) );
  NAND U7038 ( .A(n7024), .B(n6506), .Z(n6484) );
  NAND U7039 ( .A(n6482), .B(n6481), .Z(n6483) );
  AND U7040 ( .A(n6484), .B(n6483), .Z(n6503) );
  AND U7041 ( .A(y[709]), .B(x[130]), .Z(n6486) );
  NAND U7042 ( .A(y[707]), .B(x[132]), .Z(n6485) );
  XNOR U7043 ( .A(n6486), .B(n6485), .Z(n6516) );
  XOR U7044 ( .A(n6516), .B(n6515), .Z(n6501) );
  AND U7045 ( .A(y[711]), .B(x[128]), .Z(n6488) );
  NAND U7046 ( .A(y[704]), .B(x[135]), .Z(n6487) );
  XNOR U7047 ( .A(n6488), .B(n6487), .Z(n6521) );
  ANDN U7048 ( .B(o[70]), .A(n6489), .Z(n6520) );
  XNOR U7049 ( .A(n6521), .B(n6520), .Z(n6500) );
  XNOR U7050 ( .A(n6501), .B(n6500), .Z(n6502) );
  XOR U7051 ( .A(n6503), .B(n6502), .Z(n6535) );
  XOR U7052 ( .A(n6536), .B(n6535), .Z(n6537) );
  XOR U7053 ( .A(n6538), .B(n6537), .Z(n6534) );
  NANDN U7054 ( .A(n6491), .B(n6490), .Z(n6495) );
  NAND U7055 ( .A(n6493), .B(n6492), .Z(n6494) );
  NAND U7056 ( .A(n6495), .B(n6494), .Z(n6533) );
  XOR U7057 ( .A(n6533), .B(n6532), .Z(n6499) );
  XNOR U7058 ( .A(n6534), .B(n6499), .Z(N168) );
  NANDN U7059 ( .A(n6501), .B(n6500), .Z(n6505) );
  NAND U7060 ( .A(n6503), .B(n6502), .Z(n6504) );
  AND U7061 ( .A(n6505), .B(n6504), .Z(n6576) );
  AND U7062 ( .A(x[133]), .B(y[710]), .Z(n6679) );
  NAND U7063 ( .A(n6679), .B(n6506), .Z(n6510) );
  NAND U7064 ( .A(n6508), .B(n6507), .Z(n6509) );
  AND U7065 ( .A(n6510), .B(n6509), .Z(n6574) );
  ANDN U7066 ( .B(o[71]), .A(n6511), .Z(n6553) );
  AND U7067 ( .A(y[707]), .B(x[133]), .Z(n7164) );
  NAND U7068 ( .A(y[711]), .B(x[129]), .Z(n6512) );
  XNOR U7069 ( .A(n7164), .B(n6512), .Z(n6554) );
  XNOR U7070 ( .A(n6553), .B(n6554), .Z(n6558) );
  NAND U7071 ( .A(x[131]), .B(y[709]), .Z(n7370) );
  AND U7072 ( .A(y[710]), .B(x[130]), .Z(n7463) );
  AND U7073 ( .A(y[706]), .B(x[134]), .Z(n6513) );
  XOR U7074 ( .A(n7463), .B(n6513), .Z(n6564) );
  XNOR U7075 ( .A(n7240), .B(n6564), .Z(n6557) );
  XNOR U7076 ( .A(n7370), .B(n6557), .Z(n6559) );
  XOR U7077 ( .A(n6558), .B(n6559), .Z(n6573) );
  XNOR U7078 ( .A(n6574), .B(n6573), .Z(n6575) );
  XOR U7079 ( .A(n6576), .B(n6575), .Z(n6582) );
  NANDN U7080 ( .A(n6514), .B(n7024), .Z(n6518) );
  NAND U7081 ( .A(n6516), .B(n6515), .Z(n6517) );
  AND U7082 ( .A(n6518), .B(n6517), .Z(n6570) );
  AND U7083 ( .A(x[135]), .B(y[711]), .Z(n6519) );
  NAND U7084 ( .A(n7019), .B(n6519), .Z(n6523) );
  NAND U7085 ( .A(n6521), .B(n6520), .Z(n6522) );
  AND U7086 ( .A(n6523), .B(n6522), .Z(n6568) );
  AND U7087 ( .A(y[712]), .B(x[128]), .Z(n6525) );
  NAND U7088 ( .A(y[704]), .B(x[136]), .Z(n6524) );
  XNOR U7089 ( .A(n6525), .B(n6524), .Z(n6544) );
  NAND U7090 ( .A(x[135]), .B(y[705]), .Z(n6549) );
  XNOR U7091 ( .A(o[72]), .B(n6549), .Z(n6543) );
  XOR U7092 ( .A(n6544), .B(n6543), .Z(n6567) );
  XNOR U7093 ( .A(n6568), .B(n6567), .Z(n6569) );
  XOR U7094 ( .A(n6570), .B(n6569), .Z(n6580) );
  NANDN U7095 ( .A(n6527), .B(n6526), .Z(n6531) );
  NANDN U7096 ( .A(n6529), .B(n6528), .Z(n6530) );
  NAND U7097 ( .A(n6531), .B(n6530), .Z(n6579) );
  XOR U7098 ( .A(n6580), .B(n6579), .Z(n6581) );
  XOR U7099 ( .A(n6582), .B(n6581), .Z(n6588) );
  NAND U7100 ( .A(n6536), .B(n6535), .Z(n6540) );
  NAND U7101 ( .A(n6538), .B(n6537), .Z(n6539) );
  NAND U7102 ( .A(n6540), .B(n6539), .Z(n6587) );
  IV U7103 ( .A(n6587), .Z(n6585) );
  XOR U7104 ( .A(n6586), .B(n6585), .Z(n6541) );
  XNOR U7105 ( .A(n6588), .B(n6541), .Z(N169) );
  AND U7106 ( .A(x[136]), .B(y[712]), .Z(n6542) );
  NAND U7107 ( .A(n6542), .B(n7019), .Z(n6546) );
  NAND U7108 ( .A(n6544), .B(n6543), .Z(n6545) );
  AND U7109 ( .A(n6546), .B(n6545), .Z(n6628) );
  AND U7110 ( .A(y[708]), .B(x[133]), .Z(n6548) );
  NAND U7111 ( .A(y[706]), .B(x[135]), .Z(n6547) );
  XNOR U7112 ( .A(n6548), .B(n6547), .Z(n6602) );
  ANDN U7113 ( .B(o[72]), .A(n6549), .Z(n6601) );
  XOR U7114 ( .A(n6602), .B(n6601), .Z(n6626) );
  AND U7115 ( .A(y[704]), .B(x[137]), .Z(n6551) );
  NAND U7116 ( .A(y[713]), .B(x[128]), .Z(n6550) );
  XNOR U7117 ( .A(n6551), .B(n6550), .Z(n6608) );
  NAND U7118 ( .A(x[136]), .B(y[705]), .Z(n6617) );
  XNOR U7119 ( .A(o[73]), .B(n6617), .Z(n6607) );
  XNOR U7120 ( .A(n6608), .B(n6607), .Z(n6625) );
  XNOR U7121 ( .A(n6626), .B(n6625), .Z(n6627) );
  XNOR U7122 ( .A(n6628), .B(n6627), .Z(n6622) );
  AND U7123 ( .A(y[712]), .B(x[129]), .Z(n7357) );
  NAND U7124 ( .A(y[707]), .B(x[134]), .Z(n6552) );
  XNOR U7125 ( .A(n7357), .B(n6552), .Z(n6612) );
  XOR U7126 ( .A(n7024), .B(n6612), .Z(n6632) );
  NAND U7127 ( .A(x[130]), .B(y[711]), .Z(n7288) );
  NAND U7128 ( .A(x[131]), .B(y[710]), .Z(n6977) );
  XOR U7129 ( .A(n7288), .B(n6977), .Z(n6631) );
  XOR U7130 ( .A(n6632), .B(n6631), .Z(n6620) );
  NAND U7131 ( .A(x[133]), .B(y[711]), .Z(n6803) );
  NANDN U7132 ( .A(n6803), .B(n6611), .Z(n6556) );
  NAND U7133 ( .A(n6554), .B(n6553), .Z(n6555) );
  NAND U7134 ( .A(n6556), .B(n6555), .Z(n6619) );
  XOR U7135 ( .A(n6620), .B(n6619), .Z(n6621) );
  XNOR U7136 ( .A(n6622), .B(n6621), .Z(n6595) );
  NAND U7137 ( .A(n7370), .B(n6557), .Z(n6561) );
  NANDN U7138 ( .A(n6559), .B(n6558), .Z(n6560) );
  NAND U7139 ( .A(n6561), .B(n6560), .Z(n6593) );
  AND U7140 ( .A(x[130]), .B(y[706]), .Z(n6562) );
  NAND U7141 ( .A(n6563), .B(n6562), .Z(n6566) );
  NAND U7142 ( .A(n7240), .B(n6564), .Z(n6565) );
  AND U7143 ( .A(n6566), .B(n6565), .Z(n6594) );
  XNOR U7144 ( .A(n6593), .B(n6594), .Z(n6596) );
  NANDN U7145 ( .A(n6568), .B(n6567), .Z(n6572) );
  NANDN U7146 ( .A(n6570), .B(n6569), .Z(n6571) );
  AND U7147 ( .A(n6572), .B(n6571), .Z(n6636) );
  NANDN U7148 ( .A(n6574), .B(n6573), .Z(n6578) );
  NAND U7149 ( .A(n6576), .B(n6575), .Z(n6577) );
  NAND U7150 ( .A(n6578), .B(n6577), .Z(n6635) );
  XNOR U7151 ( .A(n6636), .B(n6635), .Z(n6638) );
  XOR U7152 ( .A(n6637), .B(n6638), .Z(n6643) );
  NAND U7153 ( .A(n6580), .B(n6579), .Z(n6584) );
  NANDN U7154 ( .A(n6582), .B(n6581), .Z(n6583) );
  NAND U7155 ( .A(n6584), .B(n6583), .Z(n6641) );
  NANDN U7156 ( .A(n6585), .B(n6586), .Z(n6591) );
  NOR U7157 ( .A(n6587), .B(n6586), .Z(n6589) );
  OR U7158 ( .A(n6589), .B(n6588), .Z(n6590) );
  AND U7159 ( .A(n6591), .B(n6590), .Z(n6642) );
  XOR U7160 ( .A(n6641), .B(n6642), .Z(n6592) );
  XNOR U7161 ( .A(n6643), .B(n6592), .Z(N170) );
  NAND U7162 ( .A(n6594), .B(n6593), .Z(n6598) );
  NANDN U7163 ( .A(n6596), .B(n6595), .Z(n6597) );
  NAND U7164 ( .A(n6598), .B(n6597), .Z(n6702) );
  AND U7165 ( .A(x[135]), .B(y[708]), .Z(n6600) );
  NAND U7166 ( .A(n6600), .B(n6599), .Z(n6604) );
  NAND U7167 ( .A(n6602), .B(n6601), .Z(n6603) );
  AND U7168 ( .A(n6604), .B(n6603), .Z(n6694) );
  AND U7169 ( .A(y[710]), .B(x[132]), .Z(n6606) );
  NAND U7170 ( .A(y[707]), .B(x[135]), .Z(n6605) );
  XNOR U7171 ( .A(n6606), .B(n6605), .Z(n6666) );
  AND U7172 ( .A(x[134]), .B(y[708]), .Z(n6665) );
  XOR U7173 ( .A(n6666), .B(n6665), .Z(n6692) );
  AND U7174 ( .A(x[136]), .B(y[706]), .Z(n6877) );
  NAND U7175 ( .A(x[137]), .B(y[705]), .Z(n6673) );
  XNOR U7176 ( .A(o[74]), .B(n6673), .Z(n6686) );
  XOR U7177 ( .A(n6877), .B(n6686), .Z(n6688) );
  XNOR U7178 ( .A(n6688), .B(n6687), .Z(n6691) );
  XOR U7179 ( .A(n6694), .B(n6693), .Z(n6654) );
  AND U7180 ( .A(x[137]), .B(y[713]), .Z(n7249) );
  NAND U7181 ( .A(n7249), .B(n7019), .Z(n6610) );
  NAND U7182 ( .A(n6608), .B(n6607), .Z(n6609) );
  AND U7183 ( .A(n6610), .B(n6609), .Z(n6652) );
  AND U7184 ( .A(x[134]), .B(y[712]), .Z(n6912) );
  NAND U7185 ( .A(n6912), .B(n6611), .Z(n6614) );
  NAND U7186 ( .A(n7024), .B(n6612), .Z(n6613) );
  AND U7187 ( .A(n6614), .B(n6613), .Z(n6660) );
  AND U7188 ( .A(y[714]), .B(x[128]), .Z(n6616) );
  NAND U7189 ( .A(y[704]), .B(x[138]), .Z(n6615) );
  XNOR U7190 ( .A(n6616), .B(n6615), .Z(n6670) );
  ANDN U7191 ( .B(o[73]), .A(n6617), .Z(n6669) );
  XOR U7192 ( .A(n6670), .B(n6669), .Z(n6658) );
  AND U7193 ( .A(y[713]), .B(x[129]), .Z(n7565) );
  NAND U7194 ( .A(y[711]), .B(x[131]), .Z(n6618) );
  XNOR U7195 ( .A(n7565), .B(n6618), .Z(n6682) );
  NAND U7196 ( .A(x[130]), .B(y[712]), .Z(n6683) );
  XNOR U7197 ( .A(n6682), .B(n6683), .Z(n6657) );
  XOR U7198 ( .A(n6658), .B(n6657), .Z(n6659) );
  XNOR U7199 ( .A(n6660), .B(n6659), .Z(n6651) );
  XNOR U7200 ( .A(n6652), .B(n6651), .Z(n6653) );
  XNOR U7201 ( .A(n6654), .B(n6653), .Z(n6701) );
  NAND U7202 ( .A(n6620), .B(n6619), .Z(n6624) );
  NAND U7203 ( .A(n6622), .B(n6621), .Z(n6623) );
  AND U7204 ( .A(n6624), .B(n6623), .Z(n6648) );
  NANDN U7205 ( .A(n6626), .B(n6625), .Z(n6630) );
  NAND U7206 ( .A(n6628), .B(n6627), .Z(n6629) );
  AND U7207 ( .A(n6630), .B(n6629), .Z(n6645) );
  AND U7208 ( .A(n7288), .B(n6977), .Z(n6634) );
  NANDN U7209 ( .A(n6632), .B(n6631), .Z(n6633) );
  NANDN U7210 ( .A(n6634), .B(n6633), .Z(n6646) );
  XNOR U7211 ( .A(n6645), .B(n6646), .Z(n6647) );
  XOR U7212 ( .A(n6648), .B(n6647), .Z(n6700) );
  XOR U7213 ( .A(n6702), .B(n6703), .Z(n6699) );
  NANDN U7214 ( .A(n6636), .B(n6635), .Z(n6640) );
  NAND U7215 ( .A(n6638), .B(n6637), .Z(n6639) );
  NAND U7216 ( .A(n6640), .B(n6639), .Z(n6698) );
  XOR U7217 ( .A(n6698), .B(n6697), .Z(n6644) );
  XNOR U7218 ( .A(n6699), .B(n6644), .Z(N171) );
  NANDN U7219 ( .A(n6646), .B(n6645), .Z(n6650) );
  NANDN U7220 ( .A(n6648), .B(n6647), .Z(n6649) );
  AND U7221 ( .A(n6650), .B(n6649), .Z(n6771) );
  NANDN U7222 ( .A(n6652), .B(n6651), .Z(n6656) );
  NANDN U7223 ( .A(n6654), .B(n6653), .Z(n6655) );
  AND U7224 ( .A(n6656), .B(n6655), .Z(n6769) );
  NAND U7225 ( .A(n6658), .B(n6657), .Z(n6662) );
  NANDN U7226 ( .A(n6660), .B(n6659), .Z(n6661) );
  AND U7227 ( .A(n6662), .B(n6661), .Z(n6758) );
  AND U7228 ( .A(x[135]), .B(y[710]), .Z(n6664) );
  AND U7229 ( .A(x[132]), .B(y[707]), .Z(n6663) );
  NAND U7230 ( .A(n6664), .B(n6663), .Z(n6668) );
  NAND U7231 ( .A(n6666), .B(n6665), .Z(n6667) );
  AND U7232 ( .A(n6668), .B(n6667), .Z(n6756) );
  AND U7233 ( .A(x[138]), .B(y[714]), .Z(n7469) );
  NAND U7234 ( .A(n7469), .B(n7019), .Z(n6672) );
  NAND U7235 ( .A(n6670), .B(n6669), .Z(n6671) );
  AND U7236 ( .A(n6672), .B(n6671), .Z(n6752) );
  ANDN U7237 ( .B(o[74]), .A(n6673), .Z(n6728) );
  AND U7238 ( .A(y[715]), .B(x[128]), .Z(n6675) );
  NAND U7239 ( .A(y[704]), .B(x[139]), .Z(n6674) );
  XOR U7240 ( .A(n6675), .B(n6674), .Z(n6729) );
  XNOR U7241 ( .A(n6728), .B(n6729), .Z(n6750) );
  AND U7242 ( .A(y[714]), .B(x[129]), .Z(n6677) );
  NAND U7243 ( .A(y[709]), .B(x[134]), .Z(n6676) );
  XNOR U7244 ( .A(n6677), .B(n6676), .Z(n6725) );
  NAND U7245 ( .A(x[138]), .B(y[705]), .Z(n6737) );
  XNOR U7246 ( .A(o[75]), .B(n6737), .Z(n6724) );
  XOR U7247 ( .A(n6725), .B(n6724), .Z(n6749) );
  XOR U7248 ( .A(n6750), .B(n6749), .Z(n6751) );
  XNOR U7249 ( .A(n6752), .B(n6751), .Z(n6755) );
  XNOR U7250 ( .A(n6756), .B(n6755), .Z(n6757) );
  XOR U7251 ( .A(n6758), .B(n6757), .Z(n6740) );
  NAND U7252 ( .A(x[131]), .B(y[712]), .Z(n7738) );
  NAND U7253 ( .A(y[713]), .B(x[130]), .Z(n6678) );
  XNOR U7254 ( .A(n6679), .B(n6678), .Z(n6720) );
  AND U7255 ( .A(x[132]), .B(y[711]), .Z(n6719) );
  XNOR U7256 ( .A(n6720), .B(n6719), .Z(n6744) );
  XOR U7257 ( .A(n7738), .B(n6744), .Z(n6746) );
  AND U7258 ( .A(y[706]), .B(x[137]), .Z(n6681) );
  NAND U7259 ( .A(y[708]), .B(x[135]), .Z(n6680) );
  XNOR U7260 ( .A(n6681), .B(n6680), .Z(n6733) );
  AND U7261 ( .A(x[136]), .B(y[707]), .Z(n6732) );
  XNOR U7262 ( .A(n6733), .B(n6732), .Z(n6745) );
  XOR U7263 ( .A(n6746), .B(n6745), .Z(n6710) );
  NAND U7264 ( .A(x[131]), .B(y[713]), .Z(n6794) );
  AND U7265 ( .A(x[129]), .B(y[711]), .Z(n7014) );
  NANDN U7266 ( .A(n6794), .B(n7014), .Z(n6685) );
  NANDN U7267 ( .A(n6683), .B(n6682), .Z(n6684) );
  AND U7268 ( .A(n6685), .B(n6684), .Z(n6708) );
  NAND U7269 ( .A(n6877), .B(n6686), .Z(n6690) );
  NAND U7270 ( .A(n6688), .B(n6687), .Z(n6689) );
  NAND U7271 ( .A(n6690), .B(n6689), .Z(n6707) );
  XNOR U7272 ( .A(n6708), .B(n6707), .Z(n6709) );
  XOR U7273 ( .A(n6710), .B(n6709), .Z(n6739) );
  NANDN U7274 ( .A(n6692), .B(n6691), .Z(n6696) );
  NAND U7275 ( .A(n6694), .B(n6693), .Z(n6695) );
  NAND U7276 ( .A(n6696), .B(n6695), .Z(n6738) );
  XOR U7277 ( .A(n6739), .B(n6738), .Z(n6741) );
  XNOR U7278 ( .A(n6740), .B(n6741), .Z(n6768) );
  XNOR U7279 ( .A(n6769), .B(n6768), .Z(n6770) );
  XOR U7280 ( .A(n6771), .B(n6770), .Z(n6764) );
  NANDN U7281 ( .A(n6701), .B(n6700), .Z(n6705) );
  NAND U7282 ( .A(n6703), .B(n6702), .Z(n6704) );
  AND U7283 ( .A(n6705), .B(n6704), .Z(n6762) );
  IV U7284 ( .A(n6762), .Z(n6761) );
  XOR U7285 ( .A(n6763), .B(n6761), .Z(n6706) );
  XNOR U7286 ( .A(n6764), .B(n6706), .Z(N172) );
  NANDN U7287 ( .A(n6708), .B(n6707), .Z(n6712) );
  NANDN U7288 ( .A(n6710), .B(n6709), .Z(n6711) );
  AND U7289 ( .A(n6712), .B(n6711), .Z(n6836) );
  AND U7290 ( .A(x[137]), .B(y[707]), .Z(n7458) );
  AND U7291 ( .A(y[712]), .B(x[132]), .Z(n6714) );
  NAND U7292 ( .A(y[706]), .B(x[138]), .Z(n6713) );
  XNOR U7293 ( .A(n6714), .B(n6713), .Z(n6826) );
  XOR U7294 ( .A(n7458), .B(n6826), .Z(n6805) );
  NAND U7295 ( .A(x[135]), .B(y[709]), .Z(n6802) );
  XOR U7296 ( .A(n6803), .B(n6802), .Z(n6804) );
  AND U7297 ( .A(y[716]), .B(x[128]), .Z(n6716) );
  NAND U7298 ( .A(y[704]), .B(x[140]), .Z(n6715) );
  XNOR U7299 ( .A(n6716), .B(n6715), .Z(n6819) );
  NAND U7300 ( .A(x[139]), .B(y[705]), .Z(n6799) );
  XNOR U7301 ( .A(o[76]), .B(n6799), .Z(n6818) );
  XOR U7302 ( .A(n6819), .B(n6818), .Z(n6788) );
  AND U7303 ( .A(y[714]), .B(x[130]), .Z(n6718) );
  NAND U7304 ( .A(y[708]), .B(x[136]), .Z(n6717) );
  XNOR U7305 ( .A(n6718), .B(n6717), .Z(n6793) );
  XOR U7306 ( .A(n6788), .B(n6787), .Z(n6790) );
  XOR U7307 ( .A(n6789), .B(n6790), .Z(n6784) );
  AND U7308 ( .A(x[133]), .B(y[713]), .Z(n7279) );
  NAND U7309 ( .A(n7463), .B(n7279), .Z(n6722) );
  NAND U7310 ( .A(n6720), .B(n6719), .Z(n6721) );
  AND U7311 ( .A(n6722), .B(n6721), .Z(n6782) );
  AND U7312 ( .A(x[134]), .B(y[714]), .Z(n7031) );
  NAND U7313 ( .A(n7031), .B(n6723), .Z(n6727) );
  NAND U7314 ( .A(n6725), .B(n6724), .Z(n6726) );
  NAND U7315 ( .A(n6727), .B(n6726), .Z(n6781) );
  XNOR U7316 ( .A(n6782), .B(n6781), .Z(n6783) );
  XOR U7317 ( .A(n6784), .B(n6783), .Z(n6834) );
  AND U7318 ( .A(x[139]), .B(y[715]), .Z(n7861) );
  NAND U7319 ( .A(n7861), .B(n7019), .Z(n6731) );
  NANDN U7320 ( .A(n6729), .B(n6728), .Z(n6730) );
  AND U7321 ( .A(n6731), .B(n6730), .Z(n6811) );
  AND U7322 ( .A(x[135]), .B(y[706]), .Z(n6953) );
  AND U7323 ( .A(x[137]), .B(y[708]), .Z(n6801) );
  NAND U7324 ( .A(n6953), .B(n6801), .Z(n6735) );
  NAND U7325 ( .A(n6733), .B(n6732), .Z(n6734) );
  AND U7326 ( .A(n6735), .B(n6734), .Z(n6809) );
  AND U7327 ( .A(y[715]), .B(x[129]), .Z(n7495) );
  NAND U7328 ( .A(y[710]), .B(x[134]), .Z(n6736) );
  XNOR U7329 ( .A(n7495), .B(n6736), .Z(n6815) );
  ANDN U7330 ( .B(o[75]), .A(n6737), .Z(n6814) );
  XOR U7331 ( .A(n6815), .B(n6814), .Z(n6808) );
  XNOR U7332 ( .A(n6809), .B(n6808), .Z(n6810) );
  XNOR U7333 ( .A(n6811), .B(n6810), .Z(n6833) );
  XOR U7334 ( .A(n6834), .B(n6833), .Z(n6835) );
  XOR U7335 ( .A(n6836), .B(n6835), .Z(n6840) );
  NAND U7336 ( .A(n6739), .B(n6738), .Z(n6743) );
  NAND U7337 ( .A(n6741), .B(n6740), .Z(n6742) );
  NAND U7338 ( .A(n6743), .B(n6742), .Z(n6839) );
  XOR U7339 ( .A(n6840), .B(n6839), .Z(n6842) );
  NAND U7340 ( .A(n7738), .B(n6744), .Z(n6748) );
  NAND U7341 ( .A(n6746), .B(n6745), .Z(n6747) );
  AND U7342 ( .A(n6748), .B(n6747), .Z(n6776) );
  NAND U7343 ( .A(n6750), .B(n6749), .Z(n6754) );
  NANDN U7344 ( .A(n6752), .B(n6751), .Z(n6753) );
  AND U7345 ( .A(n6754), .B(n6753), .Z(n6775) );
  XNOR U7346 ( .A(n6776), .B(n6775), .Z(n6777) );
  NANDN U7347 ( .A(n6756), .B(n6755), .Z(n6760) );
  NANDN U7348 ( .A(n6758), .B(n6757), .Z(n6759) );
  NAND U7349 ( .A(n6760), .B(n6759), .Z(n6778) );
  XNOR U7350 ( .A(n6777), .B(n6778), .Z(n6841) );
  XNOR U7351 ( .A(n6842), .B(n6841), .Z(n6848) );
  OR U7352 ( .A(n6763), .B(n6761), .Z(n6767) );
  ANDN U7353 ( .B(n6763), .A(n6762), .Z(n6765) );
  OR U7354 ( .A(n6765), .B(n6764), .Z(n6766) );
  AND U7355 ( .A(n6767), .B(n6766), .Z(n6846) );
  NANDN U7356 ( .A(n6769), .B(n6768), .Z(n6773) );
  NANDN U7357 ( .A(n6771), .B(n6770), .Z(n6772) );
  AND U7358 ( .A(n6773), .B(n6772), .Z(n6847) );
  IV U7359 ( .A(n6847), .Z(n6845) );
  XOR U7360 ( .A(n6846), .B(n6845), .Z(n6774) );
  XNOR U7361 ( .A(n6848), .B(n6774), .Z(N173) );
  NANDN U7362 ( .A(n6776), .B(n6775), .Z(n6780) );
  NANDN U7363 ( .A(n6778), .B(n6777), .Z(n6779) );
  AND U7364 ( .A(n6780), .B(n6779), .Z(n6925) );
  NANDN U7365 ( .A(n6782), .B(n6781), .Z(n6786) );
  NAND U7366 ( .A(n6784), .B(n6783), .Z(n6785) );
  AND U7367 ( .A(n6786), .B(n6785), .Z(n6860) );
  NAND U7368 ( .A(n6788), .B(n6787), .Z(n6792) );
  NAND U7369 ( .A(n6790), .B(n6789), .Z(n6791) );
  AND U7370 ( .A(n6792), .B(n6791), .Z(n6856) );
  AND U7371 ( .A(x[136]), .B(y[714]), .Z(n8147) );
  AND U7372 ( .A(x[130]), .B(y[708]), .Z(n6962) );
  NAND U7373 ( .A(n8147), .B(n6962), .Z(n6796) );
  NANDN U7374 ( .A(n6794), .B(n6793), .Z(n6795) );
  AND U7375 ( .A(n6796), .B(n6795), .Z(n6893) );
  AND U7376 ( .A(y[716]), .B(x[129]), .Z(n6798) );
  NAND U7377 ( .A(y[710]), .B(x[135]), .Z(n6797) );
  XNOR U7378 ( .A(n6798), .B(n6797), .Z(n6884) );
  ANDN U7379 ( .B(o[76]), .A(n6799), .Z(n6883) );
  XOR U7380 ( .A(n6884), .B(n6883), .Z(n6891) );
  AND U7381 ( .A(x[134]), .B(y[711]), .Z(n7899) );
  NAND U7382 ( .A(y[715]), .B(x[130]), .Z(n6800) );
  XOR U7383 ( .A(n6801), .B(n6800), .Z(n6896) );
  XNOR U7384 ( .A(n7899), .B(n6896), .Z(n6890) );
  XOR U7385 ( .A(n6891), .B(n6890), .Z(n6892) );
  XNOR U7386 ( .A(n6893), .B(n6892), .Z(n6853) );
  AND U7387 ( .A(n6803), .B(n6802), .Z(n6807) );
  NANDN U7388 ( .A(n6805), .B(n6804), .Z(n6806) );
  NANDN U7389 ( .A(n6807), .B(n6806), .Z(n6854) );
  NANDN U7390 ( .A(n6809), .B(n6808), .Z(n6813) );
  NANDN U7391 ( .A(n6811), .B(n6810), .Z(n6812) );
  AND U7392 ( .A(n6813), .B(n6812), .Z(n6868) );
  AND U7393 ( .A(x[134]), .B(y[715]), .Z(n7143) );
  IV U7394 ( .A(n7143), .Z(n7281) );
  AND U7395 ( .A(x[129]), .B(y[710]), .Z(n6882) );
  NANDN U7396 ( .A(n7281), .B(n6882), .Z(n6817) );
  NAND U7397 ( .A(n6815), .B(n6814), .Z(n6816) );
  AND U7398 ( .A(n6817), .B(n6816), .Z(n6874) );
  AND U7399 ( .A(x[140]), .B(y[716]), .Z(n8153) );
  NAND U7400 ( .A(n8153), .B(n7019), .Z(n6821) );
  NAND U7401 ( .A(n6819), .B(n6818), .Z(n6820) );
  AND U7402 ( .A(n6821), .B(n6820), .Z(n6872) );
  AND U7403 ( .A(x[138]), .B(y[707]), .Z(n7750) );
  AND U7404 ( .A(y[709]), .B(x[136]), .Z(n6823) );
  NAND U7405 ( .A(y[706]), .B(x[139]), .Z(n6822) );
  XOR U7406 ( .A(n6823), .B(n6822), .Z(n6879) );
  XNOR U7407 ( .A(n7750), .B(n6879), .Z(n6871) );
  XNOR U7408 ( .A(n6872), .B(n6871), .Z(n6873) );
  XNOR U7409 ( .A(n6874), .B(n6873), .Z(n6866) );
  AND U7410 ( .A(x[138]), .B(y[712]), .Z(n6825) );
  AND U7411 ( .A(x[132]), .B(y[706]), .Z(n6824) );
  NAND U7412 ( .A(n6825), .B(n6824), .Z(n6828) );
  NAND U7413 ( .A(n7458), .B(n6826), .Z(n6827) );
  AND U7414 ( .A(n6828), .B(n6827), .Z(n6916) );
  AND U7415 ( .A(y[717]), .B(x[128]), .Z(n6830) );
  NAND U7416 ( .A(y[704]), .B(x[141]), .Z(n6829) );
  XNOR U7417 ( .A(n6830), .B(n6829), .Z(n6908) );
  NAND U7418 ( .A(x[140]), .B(y[705]), .Z(n6901) );
  XNOR U7419 ( .A(o[77]), .B(n6901), .Z(n6907) );
  XOR U7420 ( .A(n6908), .B(n6907), .Z(n6914) );
  AND U7421 ( .A(y[712]), .B(x[133]), .Z(n6832) );
  NAND U7422 ( .A(y[714]), .B(x[131]), .Z(n6831) );
  XNOR U7423 ( .A(n6832), .B(n6831), .Z(n6903) );
  NAND U7424 ( .A(x[132]), .B(y[713]), .Z(n6904) );
  XNOR U7425 ( .A(n6903), .B(n6904), .Z(n6913) );
  XOR U7426 ( .A(n6914), .B(n6913), .Z(n6915) );
  XOR U7427 ( .A(n6866), .B(n6865), .Z(n6867) );
  XOR U7428 ( .A(n6862), .B(n6861), .Z(n6923) );
  NAND U7429 ( .A(n6834), .B(n6833), .Z(n6838) );
  NANDN U7430 ( .A(n6836), .B(n6835), .Z(n6837) );
  AND U7431 ( .A(n6838), .B(n6837), .Z(n6922) );
  XNOR U7432 ( .A(n6923), .B(n6922), .Z(n6924) );
  XOR U7433 ( .A(n6925), .B(n6924), .Z(n6921) );
  NAND U7434 ( .A(n6840), .B(n6839), .Z(n6844) );
  NAND U7435 ( .A(n6842), .B(n6841), .Z(n6843) );
  NAND U7436 ( .A(n6844), .B(n6843), .Z(n6919) );
  NANDN U7437 ( .A(n6845), .B(n6846), .Z(n6851) );
  NOR U7438 ( .A(n6847), .B(n6846), .Z(n6849) );
  OR U7439 ( .A(n6849), .B(n6848), .Z(n6850) );
  AND U7440 ( .A(n6851), .B(n6850), .Z(n6920) );
  XOR U7441 ( .A(n6919), .B(n6920), .Z(n6852) );
  XNOR U7442 ( .A(n6921), .B(n6852), .Z(N174) );
  NANDN U7443 ( .A(n6854), .B(n6853), .Z(n6858) );
  NANDN U7444 ( .A(n6856), .B(n6855), .Z(n6857) );
  AND U7445 ( .A(n6858), .B(n6857), .Z(n7008) );
  NANDN U7446 ( .A(n6860), .B(n6859), .Z(n6864) );
  NAND U7447 ( .A(n6862), .B(n6861), .Z(n6863) );
  NAND U7448 ( .A(n6864), .B(n6863), .Z(n7007) );
  NAND U7449 ( .A(n6866), .B(n6865), .Z(n6870) );
  NANDN U7450 ( .A(n6868), .B(n6867), .Z(n6869) );
  AND U7451 ( .A(n6870), .B(n6869), .Z(n6932) );
  NANDN U7452 ( .A(n6872), .B(n6871), .Z(n6876) );
  NANDN U7453 ( .A(n6874), .B(n6873), .Z(n6875) );
  AND U7454 ( .A(n6876), .B(n6875), .Z(n6938) );
  AND U7455 ( .A(x[139]), .B(y[709]), .Z(n6878) );
  NAND U7456 ( .A(n6878), .B(n6877), .Z(n6881) );
  NANDN U7457 ( .A(n6879), .B(n7750), .Z(n6880) );
  AND U7458 ( .A(n6881), .B(n6880), .Z(n6993) );
  NAND U7459 ( .A(x[135]), .B(y[716]), .Z(n7473) );
  NANDN U7460 ( .A(n7473), .B(n6882), .Z(n6886) );
  NAND U7461 ( .A(n6884), .B(n6883), .Z(n6885) );
  NAND U7462 ( .A(n6886), .B(n6885), .Z(n6992) );
  XNOR U7463 ( .A(n6993), .B(n6992), .Z(n6995) );
  AND U7464 ( .A(x[132]), .B(y[714]), .Z(n7379) );
  AND U7465 ( .A(y[715]), .B(x[131]), .Z(n6888) );
  NAND U7466 ( .A(y[710]), .B(x[136]), .Z(n6887) );
  XOR U7467 ( .A(n6888), .B(n6887), .Z(n6978) );
  XNOR U7468 ( .A(n7279), .B(n6978), .Z(n6987) );
  XOR U7469 ( .A(n7379), .B(n6987), .Z(n6989) );
  AND U7470 ( .A(x[137]), .B(y[709]), .Z(n7570) );
  AND U7471 ( .A(y[716]), .B(x[130]), .Z(n6889) );
  AND U7472 ( .A(y[708]), .B(x[138]), .Z(n7600) );
  XOR U7473 ( .A(n6889), .B(n7600), .Z(n6963) );
  XOR U7474 ( .A(n7570), .B(n6963), .Z(n6988) );
  XOR U7475 ( .A(n6989), .B(n6988), .Z(n6994) );
  XOR U7476 ( .A(n6995), .B(n6994), .Z(n6936) );
  NAND U7477 ( .A(n6891), .B(n6890), .Z(n6895) );
  NANDN U7478 ( .A(n6893), .B(n6892), .Z(n6894) );
  AND U7479 ( .A(n6895), .B(n6894), .Z(n6935) );
  XNOR U7480 ( .A(n6936), .B(n6935), .Z(n6937) );
  XOR U7481 ( .A(n6938), .B(n6937), .Z(n6930) );
  AND U7482 ( .A(x[137]), .B(y[715]), .Z(n7471) );
  NAND U7483 ( .A(n7471), .B(n6962), .Z(n6898) );
  NANDN U7484 ( .A(n6896), .B(n7899), .Z(n6897) );
  AND U7485 ( .A(n6898), .B(n6897), .Z(n6950) );
  AND U7486 ( .A(y[718]), .B(x[128]), .Z(n6900) );
  NAND U7487 ( .A(y[704]), .B(x[142]), .Z(n6899) );
  XNOR U7488 ( .A(n6900), .B(n6899), .Z(n6973) );
  ANDN U7489 ( .B(o[77]), .A(n6901), .Z(n6972) );
  XOR U7490 ( .A(n6973), .B(n6972), .Z(n6948) );
  AND U7491 ( .A(y[706]), .B(x[140]), .Z(n7560) );
  NAND U7492 ( .A(y[711]), .B(x[135]), .Z(n6902) );
  XNOR U7493 ( .A(n7560), .B(n6902), .Z(n6955) );
  NAND U7494 ( .A(x[141]), .B(y[705]), .Z(n6961) );
  XNOR U7495 ( .A(o[78]), .B(n6961), .Z(n6954) );
  XOR U7496 ( .A(n6955), .B(n6954), .Z(n6947) );
  XOR U7497 ( .A(n6948), .B(n6947), .Z(n6949) );
  XOR U7498 ( .A(n6950), .B(n6949), .Z(n6999) );
  AND U7499 ( .A(x[133]), .B(y[714]), .Z(n7032) );
  NANDN U7500 ( .A(n7738), .B(n7032), .Z(n6906) );
  NANDN U7501 ( .A(n6904), .B(n6903), .Z(n6905) );
  AND U7502 ( .A(n6906), .B(n6905), .Z(n6944) );
  AND U7503 ( .A(x[141]), .B(y[717]), .Z(n8488) );
  NAND U7504 ( .A(n8488), .B(n7019), .Z(n6910) );
  NAND U7505 ( .A(n6908), .B(n6907), .Z(n6909) );
  AND U7506 ( .A(n6910), .B(n6909), .Z(n6942) );
  NAND U7507 ( .A(y[707]), .B(x[139]), .Z(n6911) );
  XNOR U7508 ( .A(n6912), .B(n6911), .Z(n6968) );
  NAND U7509 ( .A(x[129]), .B(y[717]), .Z(n6969) );
  XNOR U7510 ( .A(n6942), .B(n6941), .Z(n6943) );
  XOR U7511 ( .A(n6944), .B(n6943), .Z(n6998) );
  XOR U7512 ( .A(n6999), .B(n6998), .Z(n7001) );
  NAND U7513 ( .A(n6914), .B(n6913), .Z(n6918) );
  NANDN U7514 ( .A(n6916), .B(n6915), .Z(n6917) );
  AND U7515 ( .A(n6918), .B(n6917), .Z(n7000) );
  XNOR U7516 ( .A(n7001), .B(n7000), .Z(n6929) );
  XNOR U7517 ( .A(n7010), .B(n7009), .Z(n7006) );
  NANDN U7518 ( .A(n6923), .B(n6922), .Z(n6927) );
  NANDN U7519 ( .A(n6925), .B(n6924), .Z(n6926) );
  AND U7520 ( .A(n6927), .B(n6926), .Z(n7005) );
  XOR U7521 ( .A(n7004), .B(n7005), .Z(n6928) );
  XNOR U7522 ( .A(n7006), .B(n6928), .Z(N175) );
  NANDN U7523 ( .A(n6930), .B(n6929), .Z(n6934) );
  NANDN U7524 ( .A(n6932), .B(n6931), .Z(n6933) );
  AND U7525 ( .A(n6934), .B(n6933), .Z(n7106) );
  NANDN U7526 ( .A(n6936), .B(n6935), .Z(n6940) );
  NAND U7527 ( .A(n6938), .B(n6937), .Z(n6939) );
  AND U7528 ( .A(n6940), .B(n6939), .Z(n7075) );
  NANDN U7529 ( .A(n6942), .B(n6941), .Z(n6946) );
  NANDN U7530 ( .A(n6944), .B(n6943), .Z(n6945) );
  AND U7531 ( .A(n6946), .B(n6945), .Z(n7081) );
  NAND U7532 ( .A(n6948), .B(n6947), .Z(n6952) );
  NANDN U7533 ( .A(n6950), .B(n6949), .Z(n6951) );
  AND U7534 ( .A(n6952), .B(n6951), .Z(n7079) );
  NAND U7535 ( .A(x[140]), .B(y[711]), .Z(n7465) );
  NANDN U7536 ( .A(n7465), .B(n6953), .Z(n6957) );
  NAND U7537 ( .A(n6955), .B(n6954), .Z(n6956) );
  AND U7538 ( .A(n6957), .B(n6956), .Z(n7055) );
  AND U7539 ( .A(y[706]), .B(x[141]), .Z(n7887) );
  NAND U7540 ( .A(y[708]), .B(x[139]), .Z(n6958) );
  XNOR U7541 ( .A(n7887), .B(n6958), .Z(n7059) );
  AND U7542 ( .A(x[140]), .B(y[707]), .Z(n7058) );
  XOR U7543 ( .A(n7059), .B(n7058), .Z(n7053) );
  AND U7544 ( .A(y[719]), .B(x[128]), .Z(n6960) );
  NAND U7545 ( .A(y[704]), .B(x[143]), .Z(n6959) );
  XNOR U7546 ( .A(n6960), .B(n6959), .Z(n7021) );
  ANDN U7547 ( .B(o[78]), .A(n6961), .Z(n7020) );
  XNOR U7548 ( .A(n7021), .B(n7020), .Z(n7052) );
  XNOR U7549 ( .A(n7053), .B(n7052), .Z(n7054) );
  XOR U7550 ( .A(n7055), .B(n7054), .Z(n7087) );
  AND U7551 ( .A(x[138]), .B(y[716]), .Z(n7900) );
  NAND U7552 ( .A(n7900), .B(n6962), .Z(n6965) );
  NAND U7553 ( .A(n7570), .B(n6963), .Z(n6964) );
  AND U7554 ( .A(n6965), .B(n6964), .Z(n7085) );
  AND U7555 ( .A(x[139]), .B(y[712]), .Z(n6967) );
  AND U7556 ( .A(x[134]), .B(y[707]), .Z(n6966) );
  NAND U7557 ( .A(n6967), .B(n6966), .Z(n6971) );
  NANDN U7558 ( .A(n6969), .B(n6968), .Z(n6970) );
  NAND U7559 ( .A(n6971), .B(n6970), .Z(n7084) );
  AND U7560 ( .A(x[142]), .B(y[718]), .Z(n8790) );
  NAND U7561 ( .A(n8790), .B(n7019), .Z(n6975) );
  NAND U7562 ( .A(n6973), .B(n6972), .Z(n6974) );
  AND U7563 ( .A(n6975), .B(n6974), .Z(n7047) );
  AND U7564 ( .A(x[136]), .B(y[715]), .Z(n6976) );
  NANDN U7565 ( .A(n6977), .B(n6976), .Z(n6980) );
  NANDN U7566 ( .A(n6978), .B(n7279), .Z(n6979) );
  NAND U7567 ( .A(n6980), .B(n6979), .Z(n7046) );
  XNOR U7568 ( .A(n7047), .B(n7046), .Z(n7049) );
  AND U7569 ( .A(y[715]), .B(x[132]), .Z(n6982) );
  NAND U7570 ( .A(y[709]), .B(x[138]), .Z(n6981) );
  XNOR U7571 ( .A(n6982), .B(n6981), .Z(n7027) );
  AND U7572 ( .A(x[135]), .B(y[712]), .Z(n7026) );
  XOR U7573 ( .A(n7027), .B(n7026), .Z(n7034) );
  NAND U7574 ( .A(x[134]), .B(y[713]), .Z(n7173) );
  XNOR U7575 ( .A(n7173), .B(n7032), .Z(n7033) );
  XOR U7576 ( .A(n7034), .B(n7033), .Z(n7068) );
  AND U7577 ( .A(y[710]), .B(x[137]), .Z(n6984) );
  NAND U7578 ( .A(y[717]), .B(x[130]), .Z(n6983) );
  XNOR U7579 ( .A(n6984), .B(n6983), .Z(n7037) );
  NAND U7580 ( .A(x[131]), .B(y[716]), .Z(n7038) );
  XNOR U7581 ( .A(n7037), .B(n7038), .Z(n7067) );
  AND U7582 ( .A(y[718]), .B(x[129]), .Z(n6986) );
  NAND U7583 ( .A(y[711]), .B(x[136]), .Z(n6985) );
  XNOR U7584 ( .A(n6986), .B(n6985), .Z(n7016) );
  NAND U7585 ( .A(x[142]), .B(y[705]), .Z(n7043) );
  XNOR U7586 ( .A(o[79]), .B(n7043), .Z(n7015) );
  XOR U7587 ( .A(n7016), .B(n7015), .Z(n7066) );
  XOR U7588 ( .A(n7067), .B(n7066), .Z(n7069) );
  XOR U7589 ( .A(n7068), .B(n7069), .Z(n7048) );
  XOR U7590 ( .A(n7049), .B(n7048), .Z(n7091) );
  NAND U7591 ( .A(n7379), .B(n6987), .Z(n6991) );
  NAND U7592 ( .A(n6989), .B(n6988), .Z(n6990) );
  AND U7593 ( .A(n6991), .B(n6990), .Z(n7090) );
  NANDN U7594 ( .A(n6993), .B(n6992), .Z(n6997) );
  NAND U7595 ( .A(n6995), .B(n6994), .Z(n6996) );
  NAND U7596 ( .A(n6997), .B(n6996), .Z(n7093) );
  XOR U7597 ( .A(n7072), .B(n7073), .Z(n7074) );
  XOR U7598 ( .A(n7075), .B(n7074), .Z(n7103) );
  NAND U7599 ( .A(n6999), .B(n6998), .Z(n7003) );
  NAND U7600 ( .A(n7001), .B(n7000), .Z(n7002) );
  AND U7601 ( .A(n7003), .B(n7002), .Z(n7104) );
  XOR U7602 ( .A(n7103), .B(n7104), .Z(n7105) );
  XOR U7603 ( .A(n7106), .B(n7105), .Z(n7099) );
  NANDN U7604 ( .A(n7008), .B(n7007), .Z(n7012) );
  NAND U7605 ( .A(n7010), .B(n7009), .Z(n7011) );
  NAND U7606 ( .A(n7012), .B(n7011), .Z(n7097) );
  IV U7607 ( .A(n7097), .Z(n7096) );
  XOR U7608 ( .A(n7098), .B(n7096), .Z(n7013) );
  XNOR U7609 ( .A(n7099), .B(n7013), .Z(N176) );
  AND U7610 ( .A(x[136]), .B(y[718]), .Z(n7759) );
  NAND U7611 ( .A(n7759), .B(n7014), .Z(n7018) );
  NAND U7612 ( .A(n7016), .B(n7015), .Z(n7017) );
  AND U7613 ( .A(n7018), .B(n7017), .Z(n7123) );
  AND U7614 ( .A(x[143]), .B(y[719]), .Z(n9201) );
  NAND U7615 ( .A(n9201), .B(n7019), .Z(n7023) );
  NAND U7616 ( .A(n7021), .B(n7020), .Z(n7022) );
  NAND U7617 ( .A(n7023), .B(n7022), .Z(n7122) );
  AND U7618 ( .A(x[138]), .B(y[715]), .Z(n7025) );
  NAND U7619 ( .A(n7025), .B(n7024), .Z(n7029) );
  NAND U7620 ( .A(n7027), .B(n7026), .Z(n7028) );
  NAND U7621 ( .A(n7029), .B(n7028), .Z(n7160) );
  AND U7622 ( .A(x[128]), .B(y[720]), .Z(n7182) );
  NAND U7623 ( .A(x[144]), .B(y[704]), .Z(n7183) );
  NAND U7624 ( .A(x[143]), .B(y[705]), .Z(n7170) );
  XNOR U7625 ( .A(o[80]), .B(n7170), .Z(n7184) );
  XOR U7626 ( .A(n7185), .B(n7184), .Z(n7159) );
  NAND U7627 ( .A(y[713]), .B(x[135]), .Z(n7030) );
  XNOR U7628 ( .A(n7031), .B(n7030), .Z(n7175) );
  AND U7629 ( .A(x[138]), .B(y[710]), .Z(n7174) );
  XOR U7630 ( .A(n7175), .B(n7174), .Z(n7158) );
  XOR U7631 ( .A(n7159), .B(n7158), .Z(n7161) );
  XOR U7632 ( .A(n7160), .B(n7161), .Z(n7124) );
  XOR U7633 ( .A(n7125), .B(n7124), .Z(n7155) );
  NANDN U7634 ( .A(n7032), .B(n7173), .Z(n7036) );
  NANDN U7635 ( .A(n7034), .B(n7033), .Z(n7035) );
  AND U7636 ( .A(n7036), .B(n7035), .Z(n7153) );
  AND U7637 ( .A(x[137]), .B(y[717]), .Z(n7871) );
  NAND U7638 ( .A(n7871), .B(n7463), .Z(n7040) );
  NANDN U7639 ( .A(n7038), .B(n7037), .Z(n7039) );
  AND U7640 ( .A(n7040), .B(n7039), .Z(n7193) );
  AND U7641 ( .A(y[719]), .B(x[129]), .Z(n7042) );
  NAND U7642 ( .A(y[712]), .B(x[136]), .Z(n7041) );
  XNOR U7643 ( .A(n7042), .B(n7041), .Z(n7179) );
  ANDN U7644 ( .B(o[79]), .A(n7043), .Z(n7178) );
  XOR U7645 ( .A(n7179), .B(n7178), .Z(n7191) );
  AND U7646 ( .A(y[706]), .B(x[142]), .Z(n7045) );
  NAND U7647 ( .A(y[709]), .B(x[139]), .Z(n7044) );
  XNOR U7648 ( .A(n7045), .B(n7044), .Z(n7134) );
  NAND U7649 ( .A(x[132]), .B(y[716]), .Z(n7135) );
  XNOR U7650 ( .A(n7134), .B(n7135), .Z(n7190) );
  XOR U7651 ( .A(n7191), .B(n7190), .Z(n7192) );
  XOR U7652 ( .A(n7193), .B(n7192), .Z(n7152) );
  XNOR U7653 ( .A(n7153), .B(n7152), .Z(n7154) );
  XNOR U7654 ( .A(n7155), .B(n7154), .Z(n7116) );
  NANDN U7655 ( .A(n7047), .B(n7046), .Z(n7051) );
  NAND U7656 ( .A(n7049), .B(n7048), .Z(n7050) );
  NAND U7657 ( .A(n7051), .B(n7050), .Z(n7117) );
  XNOR U7658 ( .A(n7116), .B(n7117), .Z(n7119) );
  NANDN U7659 ( .A(n7053), .B(n7052), .Z(n7057) );
  NAND U7660 ( .A(n7055), .B(n7054), .Z(n7056) );
  AND U7661 ( .A(n7057), .B(n7056), .Z(n7149) );
  AND U7662 ( .A(x[139]), .B(y[706]), .Z(n7711) );
  AND U7663 ( .A(x[141]), .B(y[708]), .Z(n7145) );
  NAND U7664 ( .A(n7711), .B(n7145), .Z(n7061) );
  NAND U7665 ( .A(n7059), .B(n7058), .Z(n7060) );
  AND U7666 ( .A(n7061), .B(n7060), .Z(n7131) );
  AND U7667 ( .A(y[711]), .B(x[137]), .Z(n7063) );
  NAND U7668 ( .A(y[718]), .B(x[130]), .Z(n7062) );
  XNOR U7669 ( .A(n7063), .B(n7062), .Z(n7138) );
  NAND U7670 ( .A(x[131]), .B(y[717]), .Z(n7139) );
  XNOR U7671 ( .A(n7138), .B(n7139), .Z(n7129) );
  AND U7672 ( .A(x[140]), .B(y[708]), .Z(n7876) );
  AND U7673 ( .A(y[715]), .B(x[133]), .Z(n7065) );
  NAND U7674 ( .A(y[707]), .B(x[141]), .Z(n7064) );
  XOR U7675 ( .A(n7065), .B(n7064), .Z(n7165) );
  XNOR U7676 ( .A(n7876), .B(n7165), .Z(n7128) );
  XOR U7677 ( .A(n7129), .B(n7128), .Z(n7130) );
  XOR U7678 ( .A(n7131), .B(n7130), .Z(n7146) );
  NAND U7679 ( .A(n7067), .B(n7066), .Z(n7071) );
  NAND U7680 ( .A(n7069), .B(n7068), .Z(n7070) );
  AND U7681 ( .A(n7071), .B(n7070), .Z(n7147) );
  XOR U7682 ( .A(n7146), .B(n7147), .Z(n7148) );
  XNOR U7683 ( .A(n7149), .B(n7148), .Z(n7118) );
  XOR U7684 ( .A(n7119), .B(n7118), .Z(n7204) );
  NAND U7685 ( .A(n7073), .B(n7072), .Z(n7077) );
  NANDN U7686 ( .A(n7075), .B(n7074), .Z(n7076) );
  AND U7687 ( .A(n7077), .B(n7076), .Z(n7203) );
  XNOR U7688 ( .A(n7204), .B(n7203), .Z(n7206) );
  NANDN U7689 ( .A(n7079), .B(n7078), .Z(n7083) );
  NANDN U7690 ( .A(n7081), .B(n7080), .Z(n7082) );
  AND U7691 ( .A(n7083), .B(n7082), .Z(n7113) );
  NANDN U7692 ( .A(n7085), .B(n7084), .Z(n7089) );
  NANDN U7693 ( .A(n7087), .B(n7086), .Z(n7088) );
  AND U7694 ( .A(n7089), .B(n7088), .Z(n7111) );
  NANDN U7695 ( .A(n7091), .B(n7090), .Z(n7095) );
  NANDN U7696 ( .A(n7093), .B(n7092), .Z(n7094) );
  AND U7697 ( .A(n7095), .B(n7094), .Z(n7110) );
  XNOR U7698 ( .A(n7206), .B(n7205), .Z(n7199) );
  OR U7699 ( .A(n7098), .B(n7096), .Z(n7102) );
  ANDN U7700 ( .B(n7098), .A(n7097), .Z(n7100) );
  OR U7701 ( .A(n7100), .B(n7099), .Z(n7101) );
  AND U7702 ( .A(n7102), .B(n7101), .Z(n7198) );
  NAND U7703 ( .A(n7104), .B(n7103), .Z(n7108) );
  NANDN U7704 ( .A(n7106), .B(n7105), .Z(n7107) );
  NAND U7705 ( .A(n7108), .B(n7107), .Z(n7197) );
  IV U7706 ( .A(n7197), .Z(n7196) );
  XOR U7707 ( .A(n7198), .B(n7196), .Z(n7109) );
  XNOR U7708 ( .A(n7199), .B(n7109), .Z(N177) );
  NANDN U7709 ( .A(n7111), .B(n7110), .Z(n7115) );
  NANDN U7710 ( .A(n7113), .B(n7112), .Z(n7114) );
  AND U7711 ( .A(n7115), .B(n7114), .Z(n7213) );
  NANDN U7712 ( .A(n7117), .B(n7116), .Z(n7121) );
  NAND U7713 ( .A(n7119), .B(n7118), .Z(n7120) );
  AND U7714 ( .A(n7121), .B(n7120), .Z(n7226) );
  NANDN U7715 ( .A(n7123), .B(n7122), .Z(n7127) );
  NAND U7716 ( .A(n7125), .B(n7124), .Z(n7126) );
  AND U7717 ( .A(n7127), .B(n7126), .Z(n7310) );
  NAND U7718 ( .A(n7129), .B(n7128), .Z(n7133) );
  NANDN U7719 ( .A(n7131), .B(n7130), .Z(n7132) );
  AND U7720 ( .A(n7133), .B(n7132), .Z(n7308) );
  NAND U7721 ( .A(x[142]), .B(y[709]), .Z(n7497) );
  NANDN U7722 ( .A(n7497), .B(n7711), .Z(n7137) );
  NANDN U7723 ( .A(n7135), .B(n7134), .Z(n7136) );
  AND U7724 ( .A(n7137), .B(n7136), .Z(n7302) );
  AND U7725 ( .A(y[718]), .B(x[137]), .Z(n8142) );
  NANDN U7726 ( .A(n7288), .B(n8142), .Z(n7141) );
  NANDN U7727 ( .A(n7139), .B(n7138), .Z(n7140) );
  NAND U7728 ( .A(n7141), .B(n7140), .Z(n7301) );
  XNOR U7729 ( .A(n7302), .B(n7301), .Z(n7304) );
  AND U7730 ( .A(x[135]), .B(y[714]), .Z(n7296) );
  AND U7731 ( .A(y[716]), .B(x[133]), .Z(n7338) );
  NAND U7732 ( .A(y[713]), .B(x[136]), .Z(n7142) );
  XNOR U7733 ( .A(n7338), .B(n7142), .Z(n7280) );
  XOR U7734 ( .A(n7280), .B(n7143), .Z(n7295) );
  XOR U7735 ( .A(n7296), .B(n7295), .Z(n7298) );
  NAND U7736 ( .A(y[717]), .B(x[132]), .Z(n7144) );
  XNOR U7737 ( .A(n7145), .B(n7144), .Z(n7241) );
  NAND U7738 ( .A(x[139]), .B(y[710]), .Z(n7242) );
  XNOR U7739 ( .A(n7241), .B(n7242), .Z(n7297) );
  XOR U7740 ( .A(n7298), .B(n7297), .Z(n7303) );
  XOR U7741 ( .A(n7304), .B(n7303), .Z(n7307) );
  XNOR U7742 ( .A(n7308), .B(n7307), .Z(n7309) );
  XOR U7743 ( .A(n7310), .B(n7309), .Z(n7224) );
  NAND U7744 ( .A(n7147), .B(n7146), .Z(n7151) );
  NANDN U7745 ( .A(n7149), .B(n7148), .Z(n7150) );
  NAND U7746 ( .A(n7151), .B(n7150), .Z(n7223) );
  XOR U7747 ( .A(n7224), .B(n7223), .Z(n7225) );
  XOR U7748 ( .A(n7226), .B(n7225), .Z(n7211) );
  NANDN U7749 ( .A(n7153), .B(n7152), .Z(n7157) );
  NANDN U7750 ( .A(n7155), .B(n7154), .Z(n7156) );
  AND U7751 ( .A(n7157), .B(n7156), .Z(n7232) );
  NAND U7752 ( .A(n7159), .B(n7158), .Z(n7163) );
  NAND U7753 ( .A(n7161), .B(n7160), .Z(n7162) );
  AND U7754 ( .A(n7163), .B(n7162), .Z(n7316) );
  AND U7755 ( .A(x[141]), .B(y[715]), .Z(n8161) );
  NAND U7756 ( .A(n8161), .B(n7164), .Z(n7167) );
  NANDN U7757 ( .A(n7165), .B(n7876), .Z(n7166) );
  AND U7758 ( .A(n7167), .B(n7166), .Z(n7264) );
  AND U7759 ( .A(y[712]), .B(x[137]), .Z(n7169) );
  NAND U7760 ( .A(y[720]), .B(x[129]), .Z(n7168) );
  XNOR U7761 ( .A(n7169), .B(n7168), .Z(n7285) );
  ANDN U7762 ( .B(o[80]), .A(n7170), .Z(n7284) );
  XOR U7763 ( .A(n7285), .B(n7284), .Z(n7262) );
  AND U7764 ( .A(y[706]), .B(x[143]), .Z(n7172) );
  NAND U7765 ( .A(y[709]), .B(x[140]), .Z(n7171) );
  XNOR U7766 ( .A(n7172), .B(n7171), .Z(n7237) );
  AND U7767 ( .A(x[142]), .B(y[707]), .Z(n7236) );
  XOR U7768 ( .A(n7237), .B(n7236), .Z(n7261) );
  XOR U7769 ( .A(n7262), .B(n7261), .Z(n7263) );
  NANDN U7770 ( .A(n7173), .B(n7296), .Z(n7177) );
  NAND U7771 ( .A(n7175), .B(n7174), .Z(n7176) );
  AND U7772 ( .A(n7177), .B(n7176), .Z(n7274) );
  AND U7773 ( .A(x[136]), .B(y[719]), .Z(n7971) );
  NAND U7774 ( .A(n7971), .B(n7357), .Z(n7181) );
  NAND U7775 ( .A(n7179), .B(n7178), .Z(n7180) );
  NAND U7776 ( .A(n7181), .B(n7180), .Z(n7273) );
  NANDN U7777 ( .A(n7183), .B(n7182), .Z(n7187) );
  NAND U7778 ( .A(n7185), .B(n7184), .Z(n7186) );
  AND U7779 ( .A(n7187), .B(n7186), .Z(n7270) );
  AND U7780 ( .A(x[128]), .B(y[721]), .Z(n7251) );
  AND U7781 ( .A(x[145]), .B(y[704]), .Z(n7250) );
  XOR U7782 ( .A(n7251), .B(n7250), .Z(n7253) );
  AND U7783 ( .A(x[144]), .B(y[705]), .Z(n7247) );
  XOR U7784 ( .A(n7247), .B(o[81]), .Z(n7252) );
  XOR U7785 ( .A(n7253), .B(n7252), .Z(n7268) );
  AND U7786 ( .A(y[719]), .B(x[130]), .Z(n7189) );
  NAND U7787 ( .A(y[711]), .B(x[138]), .Z(n7188) );
  XNOR U7788 ( .A(n7189), .B(n7188), .Z(n7289) );
  NAND U7789 ( .A(x[131]), .B(y[718]), .Z(n7290) );
  XNOR U7790 ( .A(n7289), .B(n7290), .Z(n7267) );
  XOR U7791 ( .A(n7268), .B(n7267), .Z(n7269) );
  XOR U7792 ( .A(n7276), .B(n7275), .Z(n7313) );
  XOR U7793 ( .A(n7314), .B(n7313), .Z(n7315) );
  NAND U7794 ( .A(n7191), .B(n7190), .Z(n7195) );
  NANDN U7795 ( .A(n7193), .B(n7192), .Z(n7194) );
  AND U7796 ( .A(n7195), .B(n7194), .Z(n7230) );
  XOR U7797 ( .A(n7229), .B(n7230), .Z(n7231) );
  XOR U7798 ( .A(n7232), .B(n7231), .Z(n7210) );
  XOR U7799 ( .A(n7211), .B(n7210), .Z(n7212) );
  OR U7800 ( .A(n7198), .B(n7196), .Z(n7202) );
  ANDN U7801 ( .B(n7198), .A(n7197), .Z(n7200) );
  OR U7802 ( .A(n7200), .B(n7199), .Z(n7201) );
  AND U7803 ( .A(n7202), .B(n7201), .Z(n7217) );
  NANDN U7804 ( .A(n7204), .B(n7203), .Z(n7208) );
  NAND U7805 ( .A(n7206), .B(n7205), .Z(n7207) );
  AND U7806 ( .A(n7208), .B(n7207), .Z(n7218) );
  IV U7807 ( .A(n7218), .Z(n7216) );
  XOR U7808 ( .A(n7217), .B(n7216), .Z(n7209) );
  XNOR U7809 ( .A(n7219), .B(n7209), .Z(N178) );
  NAND U7810 ( .A(n7211), .B(n7210), .Z(n7215) );
  NANDN U7811 ( .A(n7213), .B(n7212), .Z(n7214) );
  NAND U7812 ( .A(n7215), .B(n7214), .Z(n7433) );
  IV U7813 ( .A(n7433), .Z(n7429) );
  NANDN U7814 ( .A(n7216), .B(n7217), .Z(n7222) );
  NOR U7815 ( .A(n7218), .B(n7217), .Z(n7220) );
  OR U7816 ( .A(n7220), .B(n7219), .Z(n7221) );
  AND U7817 ( .A(n7222), .B(n7221), .Z(n7432) );
  NAND U7818 ( .A(n7224), .B(n7223), .Z(n7228) );
  NANDN U7819 ( .A(n7226), .B(n7225), .Z(n7227) );
  AND U7820 ( .A(n7228), .B(n7227), .Z(n7426) );
  NAND U7821 ( .A(n7230), .B(n7229), .Z(n7234) );
  NANDN U7822 ( .A(n7232), .B(n7231), .Z(n7233) );
  AND U7823 ( .A(n7234), .B(n7233), .Z(n7424) );
  AND U7824 ( .A(x[143]), .B(y[709]), .Z(n7235) );
  NAND U7825 ( .A(n7235), .B(n7560), .Z(n7239) );
  NAND U7826 ( .A(n7237), .B(n7236), .Z(n7238) );
  NAND U7827 ( .A(n7239), .B(n7238), .Z(n7405) );
  NAND U7828 ( .A(n8488), .B(n7240), .Z(n7244) );
  NANDN U7829 ( .A(n7242), .B(n7241), .Z(n7243) );
  AND U7830 ( .A(n7244), .B(n7243), .Z(n7396) );
  AND U7831 ( .A(y[721]), .B(x[129]), .Z(n7246) );
  NAND U7832 ( .A(y[712]), .B(x[138]), .Z(n7245) );
  XNOR U7833 ( .A(n7246), .B(n7245), .Z(n7358) );
  NAND U7834 ( .A(n7247), .B(o[81]), .Z(n7359) );
  XNOR U7835 ( .A(n7358), .B(n7359), .Z(n7394) );
  NAND U7836 ( .A(y[707]), .B(x[143]), .Z(n7248) );
  XNOR U7837 ( .A(n7249), .B(n7248), .Z(n7349) );
  NAND U7838 ( .A(x[142]), .B(y[708]), .Z(n7350) );
  XNOR U7839 ( .A(n7349), .B(n7350), .Z(n7393) );
  XOR U7840 ( .A(n7394), .B(n7393), .Z(n7395) );
  XNOR U7841 ( .A(n7396), .B(n7395), .Z(n7406) );
  XOR U7842 ( .A(n7405), .B(n7406), .Z(n7408) );
  NAND U7843 ( .A(n7251), .B(n7250), .Z(n7255) );
  NAND U7844 ( .A(n7253), .B(n7252), .Z(n7254) );
  NAND U7845 ( .A(n7255), .B(n7254), .Z(n7417) );
  AND U7846 ( .A(y[711]), .B(x[139]), .Z(n7257) );
  NAND U7847 ( .A(y[706]), .B(x[144]), .Z(n7256) );
  XNOR U7848 ( .A(n7257), .B(n7256), .Z(n7345) );
  NAND U7849 ( .A(x[130]), .B(y[720]), .Z(n7346) );
  XNOR U7850 ( .A(n7345), .B(n7346), .Z(n7418) );
  XOR U7851 ( .A(n7417), .B(n7418), .Z(n7420) );
  AND U7852 ( .A(y[717]), .B(x[133]), .Z(n7479) );
  NAND U7853 ( .A(y[716]), .B(x[134]), .Z(n7258) );
  XNOR U7854 ( .A(n7479), .B(n7258), .Z(n7341) );
  AND U7855 ( .A(y[718]), .B(x[132]), .Z(n7260) );
  NAND U7856 ( .A(y[714]), .B(x[136]), .Z(n7259) );
  XNOR U7857 ( .A(n7260), .B(n7259), .Z(n7380) );
  NAND U7858 ( .A(x[135]), .B(y[715]), .Z(n7381) );
  XNOR U7859 ( .A(n7380), .B(n7381), .Z(n7340) );
  XOR U7860 ( .A(n7341), .B(n7340), .Z(n7419) );
  XOR U7861 ( .A(n7420), .B(n7419), .Z(n7407) );
  XOR U7862 ( .A(n7408), .B(n7407), .Z(n7327) );
  NAND U7863 ( .A(n7262), .B(n7261), .Z(n7266) );
  NANDN U7864 ( .A(n7264), .B(n7263), .Z(n7265) );
  AND U7865 ( .A(n7266), .B(n7265), .Z(n7400) );
  NAND U7866 ( .A(n7268), .B(n7267), .Z(n7272) );
  NANDN U7867 ( .A(n7270), .B(n7269), .Z(n7271) );
  AND U7868 ( .A(n7272), .B(n7271), .Z(n7399) );
  XOR U7869 ( .A(n7400), .B(n7399), .Z(n7402) );
  NANDN U7870 ( .A(n7274), .B(n7273), .Z(n7278) );
  NAND U7871 ( .A(n7276), .B(n7275), .Z(n7277) );
  AND U7872 ( .A(n7278), .B(n7277), .Z(n7401) );
  XOR U7873 ( .A(n7402), .B(n7401), .Z(n7326) );
  AND U7874 ( .A(x[136]), .B(y[716]), .Z(n7606) );
  NAND U7875 ( .A(n7606), .B(n7279), .Z(n7283) );
  NANDN U7876 ( .A(n7281), .B(n7280), .Z(n7282) );
  NAND U7877 ( .A(n7283), .B(n7282), .Z(n7412) );
  AND U7878 ( .A(x[137]), .B(y[720]), .Z(n8261) );
  NAND U7879 ( .A(n8261), .B(n7357), .Z(n7287) );
  NAND U7880 ( .A(n7285), .B(n7284), .Z(n7286) );
  NAND U7881 ( .A(n7287), .B(n7286), .Z(n7411) );
  XOR U7882 ( .A(n7412), .B(n7411), .Z(n7414) );
  AND U7883 ( .A(x[138]), .B(y[719]), .Z(n8141) );
  NANDN U7884 ( .A(n7288), .B(n8141), .Z(n7292) );
  NANDN U7885 ( .A(n7290), .B(n7289), .Z(n7291) );
  AND U7886 ( .A(n7292), .B(n7291), .Z(n7390) );
  AND U7887 ( .A(x[128]), .B(y[722]), .Z(n7362) );
  NAND U7888 ( .A(x[146]), .B(y[704]), .Z(n7363) );
  XNOR U7889 ( .A(n7362), .B(n7363), .Z(n7365) );
  NAND U7890 ( .A(x[145]), .B(y[705]), .Z(n7384) );
  XNOR U7891 ( .A(o[82]), .B(n7384), .Z(n7364) );
  XOR U7892 ( .A(n7365), .B(n7364), .Z(n7388) );
  AND U7893 ( .A(y[719]), .B(x[131]), .Z(n7294) );
  NAND U7894 ( .A(y[709]), .B(x[141]), .Z(n7293) );
  XNOR U7895 ( .A(n7294), .B(n7293), .Z(n7371) );
  NAND U7896 ( .A(x[140]), .B(y[710]), .Z(n7372) );
  XNOR U7897 ( .A(n7371), .B(n7372), .Z(n7387) );
  XOR U7898 ( .A(n7388), .B(n7387), .Z(n7389) );
  XNOR U7899 ( .A(n7390), .B(n7389), .Z(n7413) );
  XOR U7900 ( .A(n7414), .B(n7413), .Z(n7333) );
  NAND U7901 ( .A(n7296), .B(n7295), .Z(n7300) );
  NAND U7902 ( .A(n7298), .B(n7297), .Z(n7299) );
  AND U7903 ( .A(n7300), .B(n7299), .Z(n7332) );
  XNOR U7904 ( .A(n7333), .B(n7332), .Z(n7334) );
  NANDN U7905 ( .A(n7302), .B(n7301), .Z(n7306) );
  NAND U7906 ( .A(n7304), .B(n7303), .Z(n7305) );
  NAND U7907 ( .A(n7306), .B(n7305), .Z(n7335) );
  XNOR U7908 ( .A(n7334), .B(n7335), .Z(n7328) );
  XOR U7909 ( .A(n7329), .B(n7328), .Z(n7323) );
  NANDN U7910 ( .A(n7308), .B(n7307), .Z(n7312) );
  NANDN U7911 ( .A(n7310), .B(n7309), .Z(n7311) );
  AND U7912 ( .A(n7312), .B(n7311), .Z(n7321) );
  NAND U7913 ( .A(n7314), .B(n7313), .Z(n7318) );
  NANDN U7914 ( .A(n7316), .B(n7315), .Z(n7317) );
  NAND U7915 ( .A(n7318), .B(n7317), .Z(n7320) );
  XOR U7916 ( .A(n7424), .B(n7423), .Z(n7425) );
  XOR U7917 ( .A(n7426), .B(n7425), .Z(n7430) );
  XNOR U7918 ( .A(n7432), .B(n7430), .Z(n7319) );
  XOR U7919 ( .A(n7429), .B(n7319), .Z(N179) );
  NANDN U7920 ( .A(n7321), .B(n7320), .Z(n7325) );
  NANDN U7921 ( .A(n7323), .B(n7322), .Z(n7324) );
  AND U7922 ( .A(n7325), .B(n7324), .Z(n7440) );
  NANDN U7923 ( .A(n7327), .B(n7326), .Z(n7331) );
  NAND U7924 ( .A(n7329), .B(n7328), .Z(n7330) );
  AND U7925 ( .A(n7331), .B(n7330), .Z(n7438) );
  NANDN U7926 ( .A(n7333), .B(n7332), .Z(n7337) );
  NANDN U7927 ( .A(n7335), .B(n7334), .Z(n7336) );
  AND U7928 ( .A(n7337), .B(n7336), .Z(n7538) );
  AND U7929 ( .A(x[134]), .B(y[717]), .Z(n7339) );
  NAND U7930 ( .A(n7339), .B(n7338), .Z(n7343) );
  NAND U7931 ( .A(n7341), .B(n7340), .Z(n7342) );
  AND U7932 ( .A(n7343), .B(n7342), .Z(n7532) );
  AND U7933 ( .A(x[144]), .B(y[711]), .Z(n7344) );
  NAND U7934 ( .A(n7344), .B(n7711), .Z(n7348) );
  NANDN U7935 ( .A(n7346), .B(n7345), .Z(n7347) );
  AND U7936 ( .A(n7348), .B(n7347), .Z(n7530) );
  AND U7937 ( .A(x[143]), .B(y[713]), .Z(n8172) );
  NAND U7938 ( .A(n8172), .B(n7458), .Z(n7352) );
  NANDN U7939 ( .A(n7350), .B(n7349), .Z(n7351) );
  AND U7940 ( .A(n7352), .B(n7351), .Z(n7449) );
  AND U7941 ( .A(y[722]), .B(x[129]), .Z(n7354) );
  NAND U7942 ( .A(y[715]), .B(x[136]), .Z(n7353) );
  XNOR U7943 ( .A(n7354), .B(n7353), .Z(n7496) );
  AND U7944 ( .A(y[721]), .B(x[130]), .Z(n7356) );
  NAND U7945 ( .A(y[710]), .B(x[141]), .Z(n7355) );
  XNOR U7946 ( .A(n7356), .B(n7355), .Z(n7464) );
  XOR U7947 ( .A(n7447), .B(n7446), .Z(n7448) );
  XNOR U7948 ( .A(n7449), .B(n7448), .Z(n7529) );
  XNOR U7949 ( .A(n7530), .B(n7529), .Z(n7531) );
  XOR U7950 ( .A(n7532), .B(n7531), .Z(n7536) );
  AND U7951 ( .A(x[138]), .B(y[721]), .Z(n8456) );
  IV U7952 ( .A(n8456), .Z(n8591) );
  NANDN U7953 ( .A(n8591), .B(n7357), .Z(n7361) );
  NANDN U7954 ( .A(n7359), .B(n7358), .Z(n7360) );
  AND U7955 ( .A(n7361), .B(n7360), .Z(n7508) );
  NANDN U7956 ( .A(n7363), .B(n7362), .Z(n7367) );
  NAND U7957 ( .A(n7365), .B(n7364), .Z(n7366) );
  AND U7958 ( .A(n7367), .B(n7366), .Z(n7506) );
  AND U7959 ( .A(y[714]), .B(x[137]), .Z(n7369) );
  NAND U7960 ( .A(y[707]), .B(x[144]), .Z(n7368) );
  XNOR U7961 ( .A(n7369), .B(n7368), .Z(n7459) );
  NAND U7962 ( .A(x[143]), .B(y[708]), .Z(n7460) );
  XNOR U7963 ( .A(n7459), .B(n7460), .Z(n7505) );
  XNOR U7964 ( .A(n7506), .B(n7505), .Z(n7507) );
  XOR U7965 ( .A(n7508), .B(n7507), .Z(n7525) );
  AND U7966 ( .A(x[141]), .B(y[719]), .Z(n8805) );
  NANDN U7967 ( .A(n7370), .B(n8805), .Z(n7374) );
  NANDN U7968 ( .A(n7372), .B(n7371), .Z(n7373) );
  AND U7969 ( .A(n7374), .B(n7373), .Z(n7514) );
  AND U7970 ( .A(y[706]), .B(x[145]), .Z(n7376) );
  NAND U7971 ( .A(y[713]), .B(x[138]), .Z(n7375) );
  XNOR U7972 ( .A(n7376), .B(n7375), .Z(n7502) );
  NAND U7973 ( .A(x[146]), .B(y[705]), .Z(n7478) );
  XNOR U7974 ( .A(o[83]), .B(n7478), .Z(n7501) );
  XOR U7975 ( .A(n7502), .B(n7501), .Z(n7512) );
  AND U7976 ( .A(y[720]), .B(x[131]), .Z(n7378) );
  NAND U7977 ( .A(y[712]), .B(x[139]), .Z(n7377) );
  XNOR U7978 ( .A(n7378), .B(n7377), .Z(n7472) );
  XOR U7979 ( .A(n7512), .B(n7511), .Z(n7513) );
  XOR U7980 ( .A(n7514), .B(n7513), .Z(n7524) );
  NAND U7981 ( .A(n7759), .B(n7379), .Z(n7383) );
  NANDN U7982 ( .A(n7381), .B(n7380), .Z(n7382) );
  AND U7983 ( .A(n7383), .B(n7382), .Z(n7455) );
  AND U7984 ( .A(x[128]), .B(y[723]), .Z(n7483) );
  NAND U7985 ( .A(x[147]), .B(y[704]), .Z(n7484) );
  XNOR U7986 ( .A(n7483), .B(n7484), .Z(n7486) );
  ANDN U7987 ( .B(o[82]), .A(n7384), .Z(n7485) );
  XOR U7988 ( .A(n7486), .B(n7485), .Z(n7453) );
  AND U7989 ( .A(x[132]), .B(y[719]), .Z(n7620) );
  AND U7990 ( .A(y[718]), .B(x[133]), .Z(n7386) );
  NAND U7991 ( .A(y[717]), .B(x[134]), .Z(n7385) );
  XOR U7992 ( .A(n7386), .B(n7385), .Z(n7480) );
  XNOR U7993 ( .A(n7620), .B(n7480), .Z(n7452) );
  XOR U7994 ( .A(n7453), .B(n7452), .Z(n7454) );
  XOR U7995 ( .A(n7455), .B(n7454), .Z(n7523) );
  XOR U7996 ( .A(n7524), .B(n7523), .Z(n7526) );
  XNOR U7997 ( .A(n7525), .B(n7526), .Z(n7519) );
  NAND U7998 ( .A(n7388), .B(n7387), .Z(n7392) );
  NANDN U7999 ( .A(n7390), .B(n7389), .Z(n7391) );
  AND U8000 ( .A(n7392), .B(n7391), .Z(n7518) );
  NAND U8001 ( .A(n7394), .B(n7393), .Z(n7398) );
  NANDN U8002 ( .A(n7396), .B(n7395), .Z(n7397) );
  NAND U8003 ( .A(n7398), .B(n7397), .Z(n7517) );
  XNOR U8004 ( .A(n7518), .B(n7517), .Z(n7520) );
  XNOR U8005 ( .A(n7519), .B(n7520), .Z(n7535) );
  XOR U8006 ( .A(n7536), .B(n7535), .Z(n7537) );
  XNOR U8007 ( .A(n7538), .B(n7537), .Z(n7550) );
  NAND U8008 ( .A(n7400), .B(n7399), .Z(n7404) );
  NAND U8009 ( .A(n7402), .B(n7401), .Z(n7403) );
  AND U8010 ( .A(n7404), .B(n7403), .Z(n7547) );
  NAND U8011 ( .A(n7406), .B(n7405), .Z(n7410) );
  NAND U8012 ( .A(n7408), .B(n7407), .Z(n7409) );
  NAND U8013 ( .A(n7410), .B(n7409), .Z(n7543) );
  NAND U8014 ( .A(n7412), .B(n7411), .Z(n7416) );
  NAND U8015 ( .A(n7414), .B(n7413), .Z(n7415) );
  NAND U8016 ( .A(n7416), .B(n7415), .Z(n7542) );
  NAND U8017 ( .A(n7418), .B(n7417), .Z(n7422) );
  NAND U8018 ( .A(n7420), .B(n7419), .Z(n7421) );
  NAND U8019 ( .A(n7422), .B(n7421), .Z(n7541) );
  XNOR U8020 ( .A(n7542), .B(n7541), .Z(n7544) );
  XNOR U8021 ( .A(n7547), .B(n7548), .Z(n7549) );
  XOR U8022 ( .A(n7438), .B(n7437), .Z(n7439) );
  XOR U8023 ( .A(n7440), .B(n7439), .Z(n7445) );
  NAND U8024 ( .A(n7424), .B(n7423), .Z(n7428) );
  NAND U8025 ( .A(n7426), .B(n7425), .Z(n7427) );
  NAND U8026 ( .A(n7428), .B(n7427), .Z(n7444) );
  ANDN U8027 ( .B(n7432), .A(n7429), .Z(n7431) );
  OR U8028 ( .A(n7431), .B(n7430), .Z(n7435) );
  NOR U8029 ( .A(n7433), .B(n7432), .Z(n7434) );
  ANDN U8030 ( .B(n7435), .A(n7434), .Z(n7443) );
  XOR U8031 ( .A(n7444), .B(n7443), .Z(n7436) );
  XNOR U8032 ( .A(n7445), .B(n7436), .Z(N180) );
  NAND U8033 ( .A(n7438), .B(n7437), .Z(n7442) );
  NANDN U8034 ( .A(n7440), .B(n7439), .Z(n7441) );
  NAND U8035 ( .A(n7442), .B(n7441), .Z(n7668) );
  IV U8036 ( .A(n7668), .Z(n7667) );
  NAND U8037 ( .A(n7447), .B(n7446), .Z(n7451) );
  NANDN U8038 ( .A(n7449), .B(n7448), .Z(n7450) );
  AND U8039 ( .A(n7451), .B(n7450), .Z(n7555) );
  NAND U8040 ( .A(n7453), .B(n7452), .Z(n7457) );
  NANDN U8041 ( .A(n7455), .B(n7454), .Z(n7456) );
  NAND U8042 ( .A(n7457), .B(n7456), .Z(n7554) );
  XNOR U8043 ( .A(n7555), .B(n7554), .Z(n7557) );
  AND U8044 ( .A(x[144]), .B(y[714]), .Z(n8414) );
  NAND U8045 ( .A(n8414), .B(n7458), .Z(n7462) );
  NANDN U8046 ( .A(n7460), .B(n7459), .Z(n7461) );
  AND U8047 ( .A(n7462), .B(n7461), .Z(n7595) );
  AND U8048 ( .A(x[141]), .B(y[721]), .Z(n9030) );
  NAND U8049 ( .A(n9030), .B(n7463), .Z(n7467) );
  NANDN U8050 ( .A(n7465), .B(n7464), .Z(n7466) );
  AND U8051 ( .A(n7467), .B(n7466), .Z(n7640) );
  NAND U8052 ( .A(y[708]), .B(x[144]), .Z(n7468) );
  XNOR U8053 ( .A(n7469), .B(n7468), .Z(n7601) );
  NAND U8054 ( .A(x[130]), .B(y[722]), .Z(n7602) );
  XNOR U8055 ( .A(n7601), .B(n7602), .Z(n7638) );
  NAND U8056 ( .A(y[709]), .B(x[143]), .Z(n7470) );
  XNOR U8057 ( .A(n7471), .B(n7470), .Z(n7571) );
  NAND U8058 ( .A(x[142]), .B(y[710]), .Z(n7572) );
  XNOR U8059 ( .A(n7571), .B(n7572), .Z(n7637) );
  XOR U8060 ( .A(n7638), .B(n7637), .Z(n7639) );
  XNOR U8061 ( .A(n7640), .B(n7639), .Z(n7594) );
  XNOR U8062 ( .A(n7595), .B(n7594), .Z(n7597) );
  AND U8063 ( .A(x[139]), .B(y[720]), .Z(n8594) );
  NANDN U8064 ( .A(n7738), .B(n8594), .Z(n7475) );
  NANDN U8065 ( .A(n7473), .B(n7472), .Z(n7474) );
  AND U8066 ( .A(n7475), .B(n7474), .Z(n7646) );
  AND U8067 ( .A(y[723]), .B(x[129]), .Z(n7477) );
  NAND U8068 ( .A(y[713]), .B(x[139]), .Z(n7476) );
  XNOR U8069 ( .A(n7477), .B(n7476), .Z(n7567) );
  NAND U8070 ( .A(x[147]), .B(y[705]), .Z(n7575) );
  XNOR U8071 ( .A(o[84]), .B(n7575), .Z(n7566) );
  XOR U8072 ( .A(n7567), .B(n7566), .Z(n7644) );
  AND U8073 ( .A(x[128]), .B(y[724]), .Z(n7625) );
  NAND U8074 ( .A(x[148]), .B(y[704]), .Z(n7626) );
  XNOR U8075 ( .A(n7625), .B(n7626), .Z(n7628) );
  ANDN U8076 ( .B(o[83]), .A(n7478), .Z(n7627) );
  XOR U8077 ( .A(n7628), .B(n7627), .Z(n7643) );
  XOR U8078 ( .A(n7644), .B(n7643), .Z(n7645) );
  XNOR U8079 ( .A(n7646), .B(n7645), .Z(n7596) );
  XOR U8080 ( .A(n7597), .B(n7596), .Z(n7556) );
  XOR U8081 ( .A(n7557), .B(n7556), .Z(n7652) );
  AND U8082 ( .A(x[134]), .B(y[718]), .Z(n7577) );
  NAND U8083 ( .A(n7577), .B(n7479), .Z(n7482) );
  NANDN U8084 ( .A(n7480), .B(n7620), .Z(n7481) );
  AND U8085 ( .A(n7482), .B(n7481), .Z(n7585) );
  NANDN U8086 ( .A(n7484), .B(n7483), .Z(n7488) );
  NAND U8087 ( .A(n7486), .B(n7485), .Z(n7487) );
  AND U8088 ( .A(n7488), .B(n7487), .Z(n7583) );
  AND U8089 ( .A(y[706]), .B(x[146]), .Z(n7490) );
  NAND U8090 ( .A(y[712]), .B(x[140]), .Z(n7489) );
  XNOR U8091 ( .A(n7490), .B(n7489), .Z(n7561) );
  NAND U8092 ( .A(x[145]), .B(y[707]), .Z(n7562) );
  XNOR U8093 ( .A(n7561), .B(n7562), .Z(n7582) );
  XNOR U8094 ( .A(n7583), .B(n7582), .Z(n7584) );
  XOR U8095 ( .A(n7585), .B(n7584), .Z(n7589) );
  AND U8096 ( .A(y[721]), .B(x[131]), .Z(n7492) );
  NAND U8097 ( .A(y[711]), .B(x[141]), .Z(n7491) );
  XNOR U8098 ( .A(n7492), .B(n7491), .Z(n7607) );
  XOR U8099 ( .A(n7607), .B(n7606), .Z(n7579) );
  AND U8100 ( .A(y[719]), .B(x[133]), .Z(n7494) );
  NAND U8101 ( .A(y[720]), .B(x[132]), .Z(n7493) );
  XNOR U8102 ( .A(n7494), .B(n7493), .Z(n7622) );
  AND U8103 ( .A(x[135]), .B(y[717]), .Z(n7621) );
  XNOR U8104 ( .A(n7622), .B(n7621), .Z(n7576) );
  XNOR U8105 ( .A(n7577), .B(n7576), .Z(n7578) );
  XOR U8106 ( .A(n7579), .B(n7578), .Z(n7633) );
  AND U8107 ( .A(x[136]), .B(y[722]), .Z(n8758) );
  NAND U8108 ( .A(n8758), .B(n7495), .Z(n7499) );
  NANDN U8109 ( .A(n7497), .B(n7496), .Z(n7498) );
  AND U8110 ( .A(n7499), .B(n7498), .Z(n7632) );
  AND U8111 ( .A(x[145]), .B(y[713]), .Z(n8420) );
  AND U8112 ( .A(x[138]), .B(y[706]), .Z(n7500) );
  NAND U8113 ( .A(n8420), .B(n7500), .Z(n7504) );
  NAND U8114 ( .A(n7502), .B(n7501), .Z(n7503) );
  NAND U8115 ( .A(n7504), .B(n7503), .Z(n7631) );
  XNOR U8116 ( .A(n7632), .B(n7631), .Z(n7634) );
  XNOR U8117 ( .A(n7633), .B(n7634), .Z(n7588) );
  XOR U8118 ( .A(n7589), .B(n7588), .Z(n7590) );
  NANDN U8119 ( .A(n7506), .B(n7505), .Z(n7510) );
  NANDN U8120 ( .A(n7508), .B(n7507), .Z(n7509) );
  NAND U8121 ( .A(n7510), .B(n7509), .Z(n7591) );
  XNOR U8122 ( .A(n7590), .B(n7591), .Z(n7649) );
  NAND U8123 ( .A(n7512), .B(n7511), .Z(n7516) );
  NANDN U8124 ( .A(n7514), .B(n7513), .Z(n7515) );
  NAND U8125 ( .A(n7516), .B(n7515), .Z(n7650) );
  XNOR U8126 ( .A(n7649), .B(n7650), .Z(n7651) );
  XOR U8127 ( .A(n7652), .B(n7651), .Z(n7656) );
  NANDN U8128 ( .A(n7518), .B(n7517), .Z(n7522) );
  NAND U8129 ( .A(n7520), .B(n7519), .Z(n7521) );
  AND U8130 ( .A(n7522), .B(n7521), .Z(n7664) );
  NAND U8131 ( .A(n7524), .B(n7523), .Z(n7528) );
  NAND U8132 ( .A(n7526), .B(n7525), .Z(n7527) );
  AND U8133 ( .A(n7528), .B(n7527), .Z(n7662) );
  NANDN U8134 ( .A(n7530), .B(n7529), .Z(n7534) );
  NANDN U8135 ( .A(n7532), .B(n7531), .Z(n7533) );
  AND U8136 ( .A(n7534), .B(n7533), .Z(n7661) );
  XNOR U8137 ( .A(n7664), .B(n7663), .Z(n7655) );
  XOR U8138 ( .A(n7656), .B(n7655), .Z(n7657) );
  NAND U8139 ( .A(n7536), .B(n7535), .Z(n7540) );
  NANDN U8140 ( .A(n7538), .B(n7537), .Z(n7539) );
  NAND U8141 ( .A(n7540), .B(n7539), .Z(n7658) );
  XNOR U8142 ( .A(n7657), .B(n7658), .Z(n7677) );
  NAND U8143 ( .A(n7542), .B(n7541), .Z(n7546) );
  NANDN U8144 ( .A(n7544), .B(n7543), .Z(n7545) );
  AND U8145 ( .A(n7546), .B(n7545), .Z(n7675) );
  NANDN U8146 ( .A(n7548), .B(n7547), .Z(n7552) );
  NANDN U8147 ( .A(n7550), .B(n7549), .Z(n7551) );
  AND U8148 ( .A(n7552), .B(n7551), .Z(n7674) );
  XOR U8149 ( .A(n7675), .B(n7674), .Z(n7676) );
  XNOR U8150 ( .A(n7669), .B(n7670), .Z(n7553) );
  XOR U8151 ( .A(n7667), .B(n7553), .Z(N181) );
  NANDN U8152 ( .A(n7555), .B(n7554), .Z(n7559) );
  NAND U8153 ( .A(n7557), .B(n7556), .Z(n7558) );
  AND U8154 ( .A(n7559), .B(n7558), .Z(n7690) );
  AND U8155 ( .A(x[146]), .B(y[712]), .Z(n8422) );
  NAND U8156 ( .A(n8422), .B(n7560), .Z(n7564) );
  NANDN U8157 ( .A(n7562), .B(n7561), .Z(n7563) );
  AND U8158 ( .A(n7564), .B(n7563), .Z(n7767) );
  AND U8159 ( .A(x[139]), .B(y[723]), .Z(n9083) );
  NAND U8160 ( .A(n9083), .B(n7565), .Z(n7569) );
  NAND U8161 ( .A(n7567), .B(n7566), .Z(n7568) );
  NAND U8162 ( .A(n7569), .B(n7568), .Z(n7766) );
  XNOR U8163 ( .A(n7767), .B(n7766), .Z(n7769) );
  AND U8164 ( .A(x[143]), .B(y[715]), .Z(n8409) );
  NAND U8165 ( .A(n8409), .B(n7570), .Z(n7574) );
  NANDN U8166 ( .A(n7572), .B(n7571), .Z(n7573) );
  AND U8167 ( .A(n7574), .B(n7573), .Z(n7725) );
  AND U8168 ( .A(x[128]), .B(y[725]), .Z(n7744) );
  NAND U8169 ( .A(x[149]), .B(y[704]), .Z(n7745) );
  XNOR U8170 ( .A(n7744), .B(n7745), .Z(n7747) );
  ANDN U8171 ( .B(o[84]), .A(n7575), .Z(n7746) );
  XOR U8172 ( .A(n7747), .B(n7746), .Z(n7723) );
  AND U8173 ( .A(x[133]), .B(y[720]), .Z(n7729) );
  AND U8174 ( .A(x[144]), .B(y[709]), .Z(n7728) );
  XOR U8175 ( .A(n7729), .B(n7728), .Z(n7731) );
  NAND U8176 ( .A(x[143]), .B(y[710]), .Z(n7730) );
  XNOR U8177 ( .A(n7731), .B(n7730), .Z(n7722) );
  XOR U8178 ( .A(n7723), .B(n7722), .Z(n7724) );
  XNOR U8179 ( .A(n7725), .B(n7724), .Z(n7768) );
  XOR U8180 ( .A(n7769), .B(n7768), .Z(n7761) );
  NANDN U8181 ( .A(n7577), .B(n7576), .Z(n7581) );
  NANDN U8182 ( .A(n7579), .B(n7578), .Z(n7580) );
  NAND U8183 ( .A(n7581), .B(n7580), .Z(n7760) );
  XNOR U8184 ( .A(n7761), .B(n7760), .Z(n7763) );
  NANDN U8185 ( .A(n7583), .B(n7582), .Z(n7587) );
  NANDN U8186 ( .A(n7585), .B(n7584), .Z(n7586) );
  AND U8187 ( .A(n7587), .B(n7586), .Z(n7762) );
  XOR U8188 ( .A(n7763), .B(n7762), .Z(n7688) );
  NAND U8189 ( .A(n7589), .B(n7588), .Z(n7593) );
  NANDN U8190 ( .A(n7591), .B(n7590), .Z(n7592) );
  AND U8191 ( .A(n7593), .B(n7592), .Z(n7687) );
  XNOR U8192 ( .A(n7688), .B(n7687), .Z(n7689) );
  XOR U8193 ( .A(n7690), .B(n7689), .Z(n7683) );
  NANDN U8194 ( .A(n7595), .B(n7594), .Z(n7599) );
  NAND U8195 ( .A(n7597), .B(n7596), .Z(n7598) );
  AND U8196 ( .A(n7599), .B(n7598), .Z(n7787) );
  NAND U8197 ( .A(n8414), .B(n7600), .Z(n7604) );
  NANDN U8198 ( .A(n7602), .B(n7601), .Z(n7603) );
  AND U8199 ( .A(n7604), .B(n7603), .Z(n7694) );
  AND U8200 ( .A(x[131]), .B(y[711]), .Z(n7605) );
  NAND U8201 ( .A(n9030), .B(n7605), .Z(n7609) );
  NAND U8202 ( .A(n7607), .B(n7606), .Z(n7608) );
  AND U8203 ( .A(n7609), .B(n7608), .Z(n7781) );
  AND U8204 ( .A(y[706]), .B(x[147]), .Z(n7611) );
  NAND U8205 ( .A(y[714]), .B(x[139]), .Z(n7610) );
  XNOR U8206 ( .A(n7611), .B(n7610), .Z(n7713) );
  NAND U8207 ( .A(x[148]), .B(y[705]), .Z(n7743) );
  XNOR U8208 ( .A(o[85]), .B(n7743), .Z(n7712) );
  XOR U8209 ( .A(n7713), .B(n7712), .Z(n7779) );
  AND U8210 ( .A(y[707]), .B(x[146]), .Z(n7613) );
  NAND U8211 ( .A(y[715]), .B(x[138]), .Z(n7612) );
  XNOR U8212 ( .A(n7613), .B(n7612), .Z(n7751) );
  NAND U8213 ( .A(x[129]), .B(y[724]), .Z(n7752) );
  XNOR U8214 ( .A(n7751), .B(n7752), .Z(n7778) );
  XOR U8215 ( .A(n7779), .B(n7778), .Z(n7780) );
  XNOR U8216 ( .A(n7781), .B(n7780), .Z(n7693) );
  XNOR U8217 ( .A(n7694), .B(n7693), .Z(n7696) );
  AND U8218 ( .A(x[135]), .B(y[718]), .Z(n7970) );
  AND U8219 ( .A(y[711]), .B(x[142]), .Z(n7615) );
  NAND U8220 ( .A(y[719]), .B(x[134]), .Z(n7614) );
  XNOR U8221 ( .A(n7615), .B(n7614), .Z(n7755) );
  XOR U8222 ( .A(n7970), .B(n7755), .Z(n7702) );
  AND U8223 ( .A(x[137]), .B(y[716]), .Z(n7700) );
  NAND U8224 ( .A(x[136]), .B(y[717]), .Z(n7699) );
  XNOR U8225 ( .A(n7700), .B(n7699), .Z(n7701) );
  XOR U8226 ( .A(n7702), .B(n7701), .Z(n7718) );
  AND U8227 ( .A(y[708]), .B(x[145]), .Z(n7617) );
  NAND U8228 ( .A(y[713]), .B(x[140]), .Z(n7616) );
  XNOR U8229 ( .A(n7617), .B(n7616), .Z(n7705) );
  NAND U8230 ( .A(x[130]), .B(y[723]), .Z(n7706) );
  XNOR U8231 ( .A(n7705), .B(n7706), .Z(n7717) );
  AND U8232 ( .A(y[722]), .B(x[131]), .Z(n7619) );
  NAND U8233 ( .A(y[712]), .B(x[141]), .Z(n7618) );
  XNOR U8234 ( .A(n7619), .B(n7618), .Z(n7739) );
  NAND U8235 ( .A(x[132]), .B(y[721]), .Z(n7740) );
  XNOR U8236 ( .A(n7739), .B(n7740), .Z(n7716) );
  XOR U8237 ( .A(n7717), .B(n7716), .Z(n7719) );
  XOR U8238 ( .A(n7718), .B(n7719), .Z(n7775) );
  NAND U8239 ( .A(n7729), .B(n7620), .Z(n7624) );
  NAND U8240 ( .A(n7622), .B(n7621), .Z(n7623) );
  AND U8241 ( .A(n7624), .B(n7623), .Z(n7773) );
  NANDN U8242 ( .A(n7626), .B(n7625), .Z(n7630) );
  NAND U8243 ( .A(n7628), .B(n7627), .Z(n7629) );
  NAND U8244 ( .A(n7630), .B(n7629), .Z(n7772) );
  XNOR U8245 ( .A(n7773), .B(n7772), .Z(n7774) );
  XOR U8246 ( .A(n7775), .B(n7774), .Z(n7695) );
  XOR U8247 ( .A(n7696), .B(n7695), .Z(n7785) );
  NANDN U8248 ( .A(n7632), .B(n7631), .Z(n7636) );
  NAND U8249 ( .A(n7634), .B(n7633), .Z(n7635) );
  NAND U8250 ( .A(n7636), .B(n7635), .Z(n7792) );
  NAND U8251 ( .A(n7638), .B(n7637), .Z(n7642) );
  NANDN U8252 ( .A(n7640), .B(n7639), .Z(n7641) );
  NAND U8253 ( .A(n7642), .B(n7641), .Z(n7791) );
  NAND U8254 ( .A(n7644), .B(n7643), .Z(n7648) );
  NANDN U8255 ( .A(n7646), .B(n7645), .Z(n7647) );
  NAND U8256 ( .A(n7648), .B(n7647), .Z(n7790) );
  XOR U8257 ( .A(n7791), .B(n7790), .Z(n7793) );
  XOR U8258 ( .A(n7792), .B(n7793), .Z(n7784) );
  XOR U8259 ( .A(n7785), .B(n7784), .Z(n7786) );
  XOR U8260 ( .A(n7787), .B(n7786), .Z(n7682) );
  NANDN U8261 ( .A(n7650), .B(n7649), .Z(n7654) );
  NANDN U8262 ( .A(n7652), .B(n7651), .Z(n7653) );
  NAND U8263 ( .A(n7654), .B(n7653), .Z(n7681) );
  XOR U8264 ( .A(n7682), .B(n7681), .Z(n7684) );
  XNOR U8265 ( .A(n7683), .B(n7684), .Z(n7805) );
  NAND U8266 ( .A(n7656), .B(n7655), .Z(n7660) );
  NANDN U8267 ( .A(n7658), .B(n7657), .Z(n7659) );
  AND U8268 ( .A(n7660), .B(n7659), .Z(n7804) );
  NANDN U8269 ( .A(n7662), .B(n7661), .Z(n7666) );
  NAND U8270 ( .A(n7664), .B(n7663), .Z(n7665) );
  AND U8271 ( .A(n7666), .B(n7665), .Z(n7803) );
  XNOR U8272 ( .A(n7804), .B(n7803), .Z(n7806) );
  XNOR U8273 ( .A(n7805), .B(n7806), .Z(n7799) );
  OR U8274 ( .A(n7669), .B(n7667), .Z(n7673) );
  ANDN U8275 ( .B(n7669), .A(n7668), .Z(n7671) );
  OR U8276 ( .A(n7671), .B(n7670), .Z(n7672) );
  AND U8277 ( .A(n7673), .B(n7672), .Z(n7798) );
  NAND U8278 ( .A(n7675), .B(n7674), .Z(n7679) );
  NANDN U8279 ( .A(n7677), .B(n7676), .Z(n7678) );
  AND U8280 ( .A(n7679), .B(n7678), .Z(n7797) );
  IV U8281 ( .A(n7797), .Z(n7796) );
  XOR U8282 ( .A(n7798), .B(n7796), .Z(n7680) );
  XNOR U8283 ( .A(n7799), .B(n7680), .Z(N182) );
  NAND U8284 ( .A(n7682), .B(n7681), .Z(n7686) );
  NAND U8285 ( .A(n7684), .B(n7683), .Z(n7685) );
  AND U8286 ( .A(n7686), .B(n7685), .Z(n7931) );
  NANDN U8287 ( .A(n7688), .B(n7687), .Z(n7692) );
  NANDN U8288 ( .A(n7690), .B(n7689), .Z(n7691) );
  AND U8289 ( .A(n7692), .B(n7691), .Z(n7929) );
  NANDN U8290 ( .A(n7694), .B(n7693), .Z(n7698) );
  NAND U8291 ( .A(n7696), .B(n7695), .Z(n7697) );
  AND U8292 ( .A(n7698), .B(n7697), .Z(n7925) );
  NANDN U8293 ( .A(n7700), .B(n7699), .Z(n7704) );
  NANDN U8294 ( .A(n7702), .B(n7701), .Z(n7703) );
  AND U8295 ( .A(n7704), .B(n7703), .Z(n7919) );
  NAND U8296 ( .A(n8420), .B(n7876), .Z(n7708) );
  NANDN U8297 ( .A(n7706), .B(n7705), .Z(n7707) );
  NAND U8298 ( .A(n7708), .B(n7707), .Z(n7848) );
  AND U8299 ( .A(x[133]), .B(y[721]), .Z(n7892) );
  NAND U8300 ( .A(x[145]), .B(y[709]), .Z(n7893) );
  XNOR U8301 ( .A(n7892), .B(n7893), .Z(n7894) );
  NAND U8302 ( .A(x[144]), .B(y[710]), .Z(n7895) );
  XNOR U8303 ( .A(n7894), .B(n7895), .Z(n7847) );
  AND U8304 ( .A(y[708]), .B(x[146]), .Z(n7710) );
  NAND U8305 ( .A(y[714]), .B(x[140]), .Z(n7709) );
  XNOR U8306 ( .A(n7710), .B(n7709), .Z(n7877) );
  NAND U8307 ( .A(x[132]), .B(y[722]), .Z(n7878) );
  XNOR U8308 ( .A(n7877), .B(n7878), .Z(n7846) );
  XOR U8309 ( .A(n7847), .B(n7846), .Z(n7849) );
  XNOR U8310 ( .A(n7848), .B(n7849), .Z(n7916) );
  AND U8311 ( .A(x[147]), .B(y[714]), .Z(n8917) );
  NAND U8312 ( .A(n8917), .B(n7711), .Z(n7715) );
  NAND U8313 ( .A(n7713), .B(n7712), .Z(n7714) );
  AND U8314 ( .A(n7715), .B(n7714), .Z(n7917) );
  XOR U8315 ( .A(n7916), .B(n7917), .Z(n7918) );
  XOR U8316 ( .A(n7919), .B(n7918), .Z(n7922) );
  NAND U8317 ( .A(n7717), .B(n7716), .Z(n7721) );
  NAND U8318 ( .A(n7719), .B(n7718), .Z(n7720) );
  AND U8319 ( .A(n7721), .B(n7720), .Z(n7905) );
  NAND U8320 ( .A(n7723), .B(n7722), .Z(n7727) );
  NANDN U8321 ( .A(n7725), .B(n7724), .Z(n7726) );
  NAND U8322 ( .A(n7727), .B(n7726), .Z(n7904) );
  XNOR U8323 ( .A(n7905), .B(n7904), .Z(n7907) );
  NAND U8324 ( .A(n7729), .B(n7728), .Z(n7733) );
  ANDN U8325 ( .B(n7731), .A(n7730), .Z(n7732) );
  ANDN U8326 ( .B(n7733), .A(n7732), .Z(n7868) );
  AND U8327 ( .A(y[706]), .B(x[148]), .Z(n7735) );
  NAND U8328 ( .A(y[713]), .B(x[141]), .Z(n7734) );
  XNOR U8329 ( .A(n7735), .B(n7734), .Z(n7888) );
  NAND U8330 ( .A(x[130]), .B(y[724]), .Z(n7889) );
  XNOR U8331 ( .A(n7888), .B(n7889), .Z(n7866) );
  AND U8332 ( .A(y[720]), .B(x[134]), .Z(n7737) );
  NAND U8333 ( .A(y[711]), .B(x[143]), .Z(n7736) );
  XOR U8334 ( .A(n7737), .B(n7736), .Z(n7901) );
  XNOR U8335 ( .A(n7900), .B(n7901), .Z(n7865) );
  XOR U8336 ( .A(n7866), .B(n7865), .Z(n7867) );
  XNOR U8337 ( .A(n7868), .B(n7867), .Z(n7911) );
  AND U8338 ( .A(x[141]), .B(y[722]), .Z(n9164) );
  NANDN U8339 ( .A(n7738), .B(n9164), .Z(n7742) );
  NANDN U8340 ( .A(n7740), .B(n7739), .Z(n7741) );
  AND U8341 ( .A(n7742), .B(n7741), .Z(n7837) );
  AND U8342 ( .A(x[129]), .B(y[725]), .Z(n7860) );
  XOR U8343 ( .A(n7861), .B(n7860), .Z(n7859) );
  ANDN U8344 ( .B(o[85]), .A(n7743), .Z(n7858) );
  XOR U8345 ( .A(n7859), .B(n7858), .Z(n7835) );
  AND U8346 ( .A(x[142]), .B(y[712]), .Z(n7852) );
  NAND U8347 ( .A(x[131]), .B(y[723]), .Z(n7853) );
  XNOR U8348 ( .A(n7852), .B(n7853), .Z(n7854) );
  NAND U8349 ( .A(x[147]), .B(y[707]), .Z(n7855) );
  XNOR U8350 ( .A(n7854), .B(n7855), .Z(n7834) );
  XOR U8351 ( .A(n7835), .B(n7834), .Z(n7836) );
  XNOR U8352 ( .A(n7837), .B(n7836), .Z(n7910) );
  XOR U8353 ( .A(n7911), .B(n7910), .Z(n7913) );
  NANDN U8354 ( .A(n7745), .B(n7744), .Z(n7749) );
  NAND U8355 ( .A(n7747), .B(n7746), .Z(n7748) );
  AND U8356 ( .A(n7749), .B(n7748), .Z(n7829) );
  AND U8357 ( .A(x[146]), .B(y[715]), .Z(n8920) );
  NAND U8358 ( .A(n8920), .B(n7750), .Z(n7754) );
  NANDN U8359 ( .A(n7752), .B(n7751), .Z(n7753) );
  NAND U8360 ( .A(n7754), .B(n7753), .Z(n7828) );
  XNOR U8361 ( .A(n7829), .B(n7828), .Z(n7831) );
  AND U8362 ( .A(x[142]), .B(y[719]), .Z(n8960) );
  NAND U8363 ( .A(n8960), .B(n7899), .Z(n7757) );
  NAND U8364 ( .A(n7970), .B(n7755), .Z(n7756) );
  AND U8365 ( .A(n7757), .B(n7756), .Z(n7843) );
  AND U8366 ( .A(x[128]), .B(y[726]), .Z(n7881) );
  NAND U8367 ( .A(x[150]), .B(y[704]), .Z(n7882) );
  XNOR U8368 ( .A(n7881), .B(n7882), .Z(n7884) );
  NAND U8369 ( .A(x[149]), .B(y[705]), .Z(n7898) );
  XNOR U8370 ( .A(o[86]), .B(n7898), .Z(n7883) );
  XOR U8371 ( .A(n7884), .B(n7883), .Z(n7841) );
  NAND U8372 ( .A(y[719]), .B(x[135]), .Z(n7758) );
  XOR U8373 ( .A(n7759), .B(n7758), .Z(n7872) );
  XNOR U8374 ( .A(n7871), .B(n7872), .Z(n7840) );
  XOR U8375 ( .A(n7841), .B(n7840), .Z(n7842) );
  XNOR U8376 ( .A(n7843), .B(n7842), .Z(n7830) );
  XOR U8377 ( .A(n7831), .B(n7830), .Z(n7912) );
  XOR U8378 ( .A(n7913), .B(n7912), .Z(n7906) );
  XOR U8379 ( .A(n7907), .B(n7906), .Z(n7923) );
  XOR U8380 ( .A(n7922), .B(n7923), .Z(n7924) );
  XOR U8381 ( .A(n7925), .B(n7924), .Z(n7818) );
  NANDN U8382 ( .A(n7761), .B(n7760), .Z(n7765) );
  NAND U8383 ( .A(n7763), .B(n7762), .Z(n7764) );
  AND U8384 ( .A(n7765), .B(n7764), .Z(n7817) );
  NANDN U8385 ( .A(n7767), .B(n7766), .Z(n7771) );
  NAND U8386 ( .A(n7769), .B(n7768), .Z(n7770) );
  AND U8387 ( .A(n7771), .B(n7770), .Z(n7825) );
  NANDN U8388 ( .A(n7773), .B(n7772), .Z(n7777) );
  NAND U8389 ( .A(n7775), .B(n7774), .Z(n7776) );
  AND U8390 ( .A(n7777), .B(n7776), .Z(n7823) );
  NAND U8391 ( .A(n7779), .B(n7778), .Z(n7783) );
  NANDN U8392 ( .A(n7781), .B(n7780), .Z(n7782) );
  NAND U8393 ( .A(n7783), .B(n7782), .Z(n7822) );
  XNOR U8394 ( .A(n7823), .B(n7822), .Z(n7824) );
  XOR U8395 ( .A(n7825), .B(n7824), .Z(n7816) );
  XNOR U8396 ( .A(n7817), .B(n7816), .Z(n7819) );
  XNOR U8397 ( .A(n7818), .B(n7819), .Z(n7812) );
  NAND U8398 ( .A(n7785), .B(n7784), .Z(n7789) );
  NANDN U8399 ( .A(n7787), .B(n7786), .Z(n7788) );
  AND U8400 ( .A(n7789), .B(n7788), .Z(n7811) );
  NAND U8401 ( .A(n7791), .B(n7790), .Z(n7795) );
  NAND U8402 ( .A(n7793), .B(n7792), .Z(n7794) );
  NAND U8403 ( .A(n7795), .B(n7794), .Z(n7810) );
  XNOR U8404 ( .A(n7811), .B(n7810), .Z(n7813) );
  XOR U8405 ( .A(n7812), .B(n7813), .Z(n7928) );
  XNOR U8406 ( .A(n7929), .B(n7928), .Z(n7930) );
  XOR U8407 ( .A(n7931), .B(n7930), .Z(n7937) );
  OR U8408 ( .A(n7798), .B(n7796), .Z(n7802) );
  ANDN U8409 ( .B(n7798), .A(n7797), .Z(n7800) );
  OR U8410 ( .A(n7800), .B(n7799), .Z(n7801) );
  AND U8411 ( .A(n7802), .B(n7801), .Z(n7935) );
  NANDN U8412 ( .A(n7804), .B(n7803), .Z(n7808) );
  NAND U8413 ( .A(n7806), .B(n7805), .Z(n7807) );
  AND U8414 ( .A(n7808), .B(n7807), .Z(n7936) );
  IV U8415 ( .A(n7936), .Z(n7934) );
  XOR U8416 ( .A(n7935), .B(n7934), .Z(n7809) );
  XNOR U8417 ( .A(n7937), .B(n7809), .Z(N183) );
  NANDN U8418 ( .A(n7811), .B(n7810), .Z(n7815) );
  NAND U8419 ( .A(n7813), .B(n7812), .Z(n7814) );
  AND U8420 ( .A(n7815), .B(n7814), .Z(n7945) );
  NANDN U8421 ( .A(n7817), .B(n7816), .Z(n7821) );
  NAND U8422 ( .A(n7819), .B(n7818), .Z(n7820) );
  AND U8423 ( .A(n7821), .B(n7820), .Z(n7943) );
  NANDN U8424 ( .A(n7823), .B(n7822), .Z(n7827) );
  NANDN U8425 ( .A(n7825), .B(n7824), .Z(n7826) );
  AND U8426 ( .A(n7827), .B(n7826), .Z(n8066) );
  NANDN U8427 ( .A(n7829), .B(n7828), .Z(n7833) );
  NAND U8428 ( .A(n7831), .B(n7830), .Z(n7832) );
  AND U8429 ( .A(n7833), .B(n7832), .Z(n8060) );
  NAND U8430 ( .A(n7835), .B(n7834), .Z(n7839) );
  NANDN U8431 ( .A(n7837), .B(n7836), .Z(n7838) );
  AND U8432 ( .A(n7839), .B(n7838), .Z(n8058) );
  NAND U8433 ( .A(n7841), .B(n7840), .Z(n7845) );
  NANDN U8434 ( .A(n7843), .B(n7842), .Z(n7844) );
  NAND U8435 ( .A(n7845), .B(n7844), .Z(n8057) );
  XNOR U8436 ( .A(n8058), .B(n8057), .Z(n8059) );
  XNOR U8437 ( .A(n8060), .B(n8059), .Z(n8078) );
  NAND U8438 ( .A(n7847), .B(n7846), .Z(n7851) );
  NAND U8439 ( .A(n7849), .B(n7848), .Z(n7850) );
  AND U8440 ( .A(n7851), .B(n7850), .Z(n8076) );
  NANDN U8441 ( .A(n7853), .B(n7852), .Z(n7857) );
  NANDN U8442 ( .A(n7855), .B(n7854), .Z(n7856) );
  AND U8443 ( .A(n7857), .B(n7856), .Z(n8004) );
  AND U8444 ( .A(n7859), .B(n7858), .Z(n7863) );
  NAND U8445 ( .A(n7861), .B(n7860), .Z(n7862) );
  NANDN U8446 ( .A(n7863), .B(n7862), .Z(n8003) );
  XNOR U8447 ( .A(n8004), .B(n8003), .Z(n8006) );
  NAND U8448 ( .A(y[720]), .B(x[135]), .Z(n7864) );
  XOR U8449 ( .A(n8142), .B(n7864), .Z(n7972) );
  XNOR U8450 ( .A(n7971), .B(n7972), .Z(n8009) );
  NAND U8451 ( .A(x[138]), .B(y[717]), .Z(n8010) );
  XNOR U8452 ( .A(n8009), .B(n8010), .Z(n8012) );
  AND U8453 ( .A(x[134]), .B(y[721]), .Z(n7962) );
  NAND U8454 ( .A(x[143]), .B(y[712]), .Z(n7963) );
  XNOR U8455 ( .A(n7962), .B(n7963), .Z(n7964) );
  NAND U8456 ( .A(x[139]), .B(y[716]), .Z(n7965) );
  XNOR U8457 ( .A(n7964), .B(n7965), .Z(n8011) );
  XOR U8458 ( .A(n8012), .B(n8011), .Z(n8005) );
  XOR U8459 ( .A(n8006), .B(n8005), .Z(n8075) );
  XNOR U8460 ( .A(n8076), .B(n8075), .Z(n8077) );
  XOR U8461 ( .A(n8078), .B(n8077), .Z(n8064) );
  NAND U8462 ( .A(n7866), .B(n7865), .Z(n7870) );
  NANDN U8463 ( .A(n7868), .B(n7867), .Z(n7869) );
  AND U8464 ( .A(n7870), .B(n7869), .Z(n7998) );
  NAND U8465 ( .A(n7970), .B(n7971), .Z(n7874) );
  NANDN U8466 ( .A(n7872), .B(n7871), .Z(n7873) );
  AND U8467 ( .A(n7874), .B(n7873), .Z(n8048) );
  AND U8468 ( .A(x[128]), .B(y[727]), .Z(n7981) );
  NAND U8469 ( .A(x[151]), .B(y[704]), .Z(n7982) );
  XNOR U8470 ( .A(n7981), .B(n7982), .Z(n7984) );
  NAND U8471 ( .A(x[150]), .B(y[705]), .Z(n7961) );
  XNOR U8472 ( .A(o[87]), .B(n7961), .Z(n7983) );
  XOR U8473 ( .A(n7984), .B(n7983), .Z(n8046) );
  AND U8474 ( .A(y[707]), .B(x[148]), .Z(n8634) );
  NAND U8475 ( .A(y[711]), .B(x[144]), .Z(n7875) );
  XNOR U8476 ( .A(n8634), .B(n7875), .Z(n7957) );
  NAND U8477 ( .A(x[147]), .B(y[708]), .Z(n7958) );
  XNOR U8478 ( .A(n7957), .B(n7958), .Z(n8045) );
  XOR U8479 ( .A(n8046), .B(n8045), .Z(n8047) );
  NAND U8480 ( .A(x[146]), .B(y[714]), .Z(n8771) );
  NANDN U8481 ( .A(n8771), .B(n7876), .Z(n7880) );
  NANDN U8482 ( .A(n7878), .B(n7877), .Z(n7879) );
  AND U8483 ( .A(n7880), .B(n7879), .Z(n8034) );
  NANDN U8484 ( .A(n7882), .B(n7881), .Z(n7886) );
  NAND U8485 ( .A(n7884), .B(n7883), .Z(n7885) );
  NAND U8486 ( .A(n7886), .B(n7885), .Z(n8033) );
  XOR U8487 ( .A(n8036), .B(n8035), .Z(n7997) );
  XNOR U8488 ( .A(n7998), .B(n7997), .Z(n8000) );
  NAND U8489 ( .A(x[148]), .B(y[713]), .Z(n8970) );
  NANDN U8490 ( .A(n8970), .B(n7887), .Z(n7891) );
  NANDN U8491 ( .A(n7889), .B(n7888), .Z(n7890) );
  AND U8492 ( .A(n7891), .B(n7890), .Z(n7992) );
  NANDN U8493 ( .A(n7893), .B(n7892), .Z(n7897) );
  NANDN U8494 ( .A(n7895), .B(n7894), .Z(n7896) );
  AND U8495 ( .A(n7897), .B(n7896), .Z(n8054) );
  AND U8496 ( .A(x[141]), .B(y[714]), .Z(n8027) );
  NAND U8497 ( .A(x[130]), .B(y[725]), .Z(n8028) );
  XNOR U8498 ( .A(n8027), .B(n8028), .Z(n8029) );
  NAND U8499 ( .A(x[149]), .B(y[706]), .Z(n8030) );
  XNOR U8500 ( .A(n8029), .B(n8030), .Z(n8052) );
  AND U8501 ( .A(x[140]), .B(y[715]), .Z(n7975) );
  NAND U8502 ( .A(x[129]), .B(y[726]), .Z(n7976) );
  XNOR U8503 ( .A(n7975), .B(n7976), .Z(n7978) );
  ANDN U8504 ( .B(o[86]), .A(n7898), .Z(n7977) );
  XOR U8505 ( .A(n7978), .B(n7977), .Z(n8051) );
  XOR U8506 ( .A(n8052), .B(n8051), .Z(n8053) );
  XNOR U8507 ( .A(n7992), .B(n7991), .Z(n7994) );
  AND U8508 ( .A(x[143]), .B(y[720]), .Z(n9158) );
  NAND U8509 ( .A(n9158), .B(n7899), .Z(n7903) );
  NANDN U8510 ( .A(n7901), .B(n7900), .Z(n7902) );
  AND U8511 ( .A(n7903), .B(n7902), .Z(n8042) );
  AND U8512 ( .A(x[142]), .B(y[713]), .Z(n8021) );
  NAND U8513 ( .A(x[131]), .B(y[724]), .Z(n8022) );
  XNOR U8514 ( .A(n8021), .B(n8022), .Z(n8023) );
  NAND U8515 ( .A(x[132]), .B(y[723]), .Z(n8024) );
  XNOR U8516 ( .A(n8023), .B(n8024), .Z(n8040) );
  AND U8517 ( .A(x[133]), .B(y[722]), .Z(n8015) );
  NAND U8518 ( .A(x[146]), .B(y[709]), .Z(n8016) );
  XNOR U8519 ( .A(n8015), .B(n8016), .Z(n8017) );
  NAND U8520 ( .A(x[145]), .B(y[710]), .Z(n8018) );
  XNOR U8521 ( .A(n8017), .B(n8018), .Z(n8039) );
  XOR U8522 ( .A(n8040), .B(n8039), .Z(n8041) );
  XOR U8523 ( .A(n7994), .B(n7993), .Z(n7999) );
  XOR U8524 ( .A(n8000), .B(n7999), .Z(n8063) );
  XOR U8525 ( .A(n8064), .B(n8063), .Z(n8065) );
  XOR U8526 ( .A(n8066), .B(n8065), .Z(n7953) );
  NANDN U8527 ( .A(n7905), .B(n7904), .Z(n7909) );
  NAND U8528 ( .A(n7907), .B(n7906), .Z(n7908) );
  AND U8529 ( .A(n7909), .B(n7908), .Z(n8072) );
  NAND U8530 ( .A(n7911), .B(n7910), .Z(n7915) );
  NAND U8531 ( .A(n7913), .B(n7912), .Z(n7914) );
  AND U8532 ( .A(n7915), .B(n7914), .Z(n8070) );
  NAND U8533 ( .A(n7917), .B(n7916), .Z(n7921) );
  NANDN U8534 ( .A(n7919), .B(n7918), .Z(n7920) );
  AND U8535 ( .A(n7921), .B(n7920), .Z(n8069) );
  XNOR U8536 ( .A(n8070), .B(n8069), .Z(n8071) );
  XOR U8537 ( .A(n8072), .B(n8071), .Z(n7951) );
  NAND U8538 ( .A(n7923), .B(n7922), .Z(n7927) );
  NANDN U8539 ( .A(n7925), .B(n7924), .Z(n7926) );
  AND U8540 ( .A(n7927), .B(n7926), .Z(n7952) );
  XOR U8541 ( .A(n7951), .B(n7952), .Z(n7954) );
  XOR U8542 ( .A(n7953), .B(n7954), .Z(n7942) );
  XNOR U8543 ( .A(n7943), .B(n7942), .Z(n7944) );
  XOR U8544 ( .A(n7945), .B(n7944), .Z(n7950) );
  NANDN U8545 ( .A(n7929), .B(n7928), .Z(n7933) );
  NAND U8546 ( .A(n7931), .B(n7930), .Z(n7932) );
  NAND U8547 ( .A(n7933), .B(n7932), .Z(n7949) );
  NANDN U8548 ( .A(n7934), .B(n7935), .Z(n7940) );
  NOR U8549 ( .A(n7936), .B(n7935), .Z(n7938) );
  OR U8550 ( .A(n7938), .B(n7937), .Z(n7939) );
  AND U8551 ( .A(n7940), .B(n7939), .Z(n7948) );
  XOR U8552 ( .A(n7949), .B(n7948), .Z(n7941) );
  XNOR U8553 ( .A(n7950), .B(n7941), .Z(N184) );
  NANDN U8554 ( .A(n7943), .B(n7942), .Z(n7947) );
  NAND U8555 ( .A(n7945), .B(n7944), .Z(n7946) );
  NAND U8556 ( .A(n7947), .B(n7946), .Z(n8221) );
  IV U8557 ( .A(n8221), .Z(n8219) );
  NAND U8558 ( .A(n7952), .B(n7951), .Z(n7956) );
  NAND U8559 ( .A(n7954), .B(n7953), .Z(n7955) );
  AND U8560 ( .A(n7956), .B(n7955), .Z(n8216) );
  AND U8561 ( .A(x[148]), .B(y[711]), .Z(n8513) );
  AND U8562 ( .A(x[144]), .B(y[707]), .Z(n8106) );
  NAND U8563 ( .A(n8513), .B(n8106), .Z(n7960) );
  NANDN U8564 ( .A(n7958), .B(n7957), .Z(n7959) );
  AND U8565 ( .A(n7960), .B(n7959), .Z(n8132) );
  AND U8566 ( .A(x[150]), .B(y[706]), .Z(n8152) );
  XOR U8567 ( .A(n8153), .B(n8152), .Z(n8155) );
  AND U8568 ( .A(x[130]), .B(y[726]), .Z(n8154) );
  XOR U8569 ( .A(n8155), .B(n8154), .Z(n8130) );
  AND U8570 ( .A(x[129]), .B(y[727]), .Z(n8160) );
  XOR U8571 ( .A(n8161), .B(n8160), .Z(n8159) );
  ANDN U8572 ( .B(o[87]), .A(n7961), .Z(n8158) );
  XOR U8573 ( .A(n8159), .B(n8158), .Z(n8129) );
  XOR U8574 ( .A(n8130), .B(n8129), .Z(n8131) );
  XNOR U8575 ( .A(n8132), .B(n8131), .Z(n8190) );
  NANDN U8576 ( .A(n7963), .B(n7962), .Z(n7967) );
  NANDN U8577 ( .A(n7965), .B(n7964), .Z(n7966) );
  AND U8578 ( .A(n7967), .B(n7966), .Z(n8126) );
  AND U8579 ( .A(y[707]), .B(x[149]), .Z(n7969) );
  NAND U8580 ( .A(y[712]), .B(x[144]), .Z(n7968) );
  XNOR U8581 ( .A(n7969), .B(n7968), .Z(n8108) );
  AND U8582 ( .A(x[133]), .B(y[723]), .Z(n8107) );
  XOR U8583 ( .A(n8108), .B(n8107), .Z(n8124) );
  AND U8584 ( .A(x[134]), .B(y[722]), .Z(n8500) );
  AND U8585 ( .A(x[148]), .B(y[708]), .Z(n8335) );
  XOR U8586 ( .A(n8500), .B(n8335), .Z(n8114) );
  AND U8587 ( .A(x[147]), .B(y[709]), .Z(n8113) );
  XOR U8588 ( .A(n8114), .B(n8113), .Z(n8123) );
  XOR U8589 ( .A(n8124), .B(n8123), .Z(n8125) );
  XNOR U8590 ( .A(n8126), .B(n8125), .Z(n8103) );
  NAND U8591 ( .A(n8261), .B(n7970), .Z(n7974) );
  NANDN U8592 ( .A(n7972), .B(n7971), .Z(n7973) );
  AND U8593 ( .A(n7974), .B(n7973), .Z(n8101) );
  NANDN U8594 ( .A(n7976), .B(n7975), .Z(n7980) );
  NAND U8595 ( .A(n7978), .B(n7977), .Z(n7979) );
  NAND U8596 ( .A(n7980), .B(n7979), .Z(n8100) );
  XNOR U8597 ( .A(n8101), .B(n8100), .Z(n8102) );
  XOR U8598 ( .A(n8103), .B(n8102), .Z(n8189) );
  XOR U8599 ( .A(n8190), .B(n8189), .Z(n8192) );
  NANDN U8600 ( .A(n7982), .B(n7981), .Z(n7986) );
  NAND U8601 ( .A(n7984), .B(n7983), .Z(n7985) );
  AND U8602 ( .A(n7986), .B(n7985), .Z(n8184) );
  AND U8603 ( .A(x[131]), .B(y[725]), .Z(n8171) );
  XOR U8604 ( .A(n8172), .B(n8171), .Z(n8174) );
  NAND U8605 ( .A(x[132]), .B(y[724]), .Z(n8173) );
  XNOR U8606 ( .A(n8174), .B(n8173), .Z(n8183) );
  AND U8607 ( .A(y[719]), .B(x[137]), .Z(n7988) );
  NAND U8608 ( .A(y[718]), .B(x[138]), .Z(n7987) );
  XNOR U8609 ( .A(n7988), .B(n7987), .Z(n8144) );
  AND U8610 ( .A(y[714]), .B(x[142]), .Z(n7990) );
  NAND U8611 ( .A(y[720]), .B(x[136]), .Z(n7989) );
  XNOR U8612 ( .A(n7990), .B(n7989), .Z(n8148) );
  NAND U8613 ( .A(x[139]), .B(y[717]), .Z(n8149) );
  XOR U8614 ( .A(n8144), .B(n8143), .Z(n8185) );
  XOR U8615 ( .A(n8186), .B(n8185), .Z(n8191) );
  XOR U8616 ( .A(n8192), .B(n8191), .Z(n8202) );
  NANDN U8617 ( .A(n7992), .B(n7991), .Z(n7996) );
  NAND U8618 ( .A(n7994), .B(n7993), .Z(n7995) );
  AND U8619 ( .A(n7996), .B(n7995), .Z(n8201) );
  XNOR U8620 ( .A(n8202), .B(n8201), .Z(n8203) );
  NANDN U8621 ( .A(n7998), .B(n7997), .Z(n8002) );
  NAND U8622 ( .A(n8000), .B(n7999), .Z(n8001) );
  NAND U8623 ( .A(n8002), .B(n8001), .Z(n8204) );
  XNOR U8624 ( .A(n8203), .B(n8204), .Z(n8210) );
  NANDN U8625 ( .A(n8004), .B(n8003), .Z(n8008) );
  NAND U8626 ( .A(n8006), .B(n8005), .Z(n8007) );
  AND U8627 ( .A(n8008), .B(n8007), .Z(n8198) );
  NANDN U8628 ( .A(n8010), .B(n8009), .Z(n8014) );
  NAND U8629 ( .A(n8012), .B(n8011), .Z(n8013) );
  AND U8630 ( .A(n8014), .B(n8013), .Z(n8196) );
  NANDN U8631 ( .A(n8016), .B(n8015), .Z(n8020) );
  NANDN U8632 ( .A(n8018), .B(n8017), .Z(n8019) );
  AND U8633 ( .A(n8020), .B(n8019), .Z(n8120) );
  AND U8634 ( .A(x[128]), .B(y[728]), .Z(n8178) );
  AND U8635 ( .A(x[152]), .B(y[704]), .Z(n8177) );
  XOR U8636 ( .A(n8178), .B(n8177), .Z(n8180) );
  AND U8637 ( .A(x[151]), .B(y[705]), .Z(n8170) );
  XOR U8638 ( .A(n8170), .B(o[88]), .Z(n8179) );
  XOR U8639 ( .A(n8180), .B(n8179), .Z(n8118) );
  AND U8640 ( .A(x[135]), .B(y[721]), .Z(n8165) );
  AND U8641 ( .A(x[146]), .B(y[710]), .Z(n8164) );
  XOR U8642 ( .A(n8165), .B(n8164), .Z(n8167) );
  AND U8643 ( .A(x[145]), .B(y[711]), .Z(n8166) );
  XOR U8644 ( .A(n8167), .B(n8166), .Z(n8117) );
  XOR U8645 ( .A(n8118), .B(n8117), .Z(n8119) );
  XNOR U8646 ( .A(n8120), .B(n8119), .Z(n8097) );
  NANDN U8647 ( .A(n8022), .B(n8021), .Z(n8026) );
  NANDN U8648 ( .A(n8024), .B(n8023), .Z(n8025) );
  AND U8649 ( .A(n8026), .B(n8025), .Z(n8095) );
  NANDN U8650 ( .A(n8028), .B(n8027), .Z(n8032) );
  NANDN U8651 ( .A(n8030), .B(n8029), .Z(n8031) );
  NAND U8652 ( .A(n8032), .B(n8031), .Z(n8094) );
  XNOR U8653 ( .A(n8095), .B(n8094), .Z(n8096) );
  XOR U8654 ( .A(n8097), .B(n8096), .Z(n8195) );
  XNOR U8655 ( .A(n8196), .B(n8195), .Z(n8197) );
  XOR U8656 ( .A(n8198), .B(n8197), .Z(n8137) );
  NANDN U8657 ( .A(n8034), .B(n8033), .Z(n8038) );
  NAND U8658 ( .A(n8036), .B(n8035), .Z(n8037) );
  AND U8659 ( .A(n8038), .B(n8037), .Z(n8091) );
  NAND U8660 ( .A(n8040), .B(n8039), .Z(n8044) );
  NANDN U8661 ( .A(n8042), .B(n8041), .Z(n8043) );
  AND U8662 ( .A(n8044), .B(n8043), .Z(n8088) );
  NAND U8663 ( .A(n8046), .B(n8045), .Z(n8050) );
  NANDN U8664 ( .A(n8048), .B(n8047), .Z(n8049) );
  NAND U8665 ( .A(n8050), .B(n8049), .Z(n8089) );
  XNOR U8666 ( .A(n8088), .B(n8089), .Z(n8090) );
  XOR U8667 ( .A(n8091), .B(n8090), .Z(n8135) );
  NAND U8668 ( .A(n8052), .B(n8051), .Z(n8056) );
  NANDN U8669 ( .A(n8054), .B(n8053), .Z(n8055) );
  NAND U8670 ( .A(n8056), .B(n8055), .Z(n8136) );
  XNOR U8671 ( .A(n8135), .B(n8136), .Z(n8138) );
  XOR U8672 ( .A(n8137), .B(n8138), .Z(n8207) );
  NANDN U8673 ( .A(n8058), .B(n8057), .Z(n8062) );
  NANDN U8674 ( .A(n8060), .B(n8059), .Z(n8061) );
  NAND U8675 ( .A(n8062), .B(n8061), .Z(n8208) );
  XNOR U8676 ( .A(n8207), .B(n8208), .Z(n8209) );
  XOR U8677 ( .A(n8210), .B(n8209), .Z(n8214) );
  NAND U8678 ( .A(n8064), .B(n8063), .Z(n8068) );
  NANDN U8679 ( .A(n8066), .B(n8065), .Z(n8067) );
  AND U8680 ( .A(n8068), .B(n8067), .Z(n8085) );
  NANDN U8681 ( .A(n8070), .B(n8069), .Z(n8074) );
  NANDN U8682 ( .A(n8072), .B(n8071), .Z(n8073) );
  AND U8683 ( .A(n8074), .B(n8073), .Z(n8083) );
  NANDN U8684 ( .A(n8076), .B(n8075), .Z(n8080) );
  NAND U8685 ( .A(n8078), .B(n8077), .Z(n8079) );
  NAND U8686 ( .A(n8080), .B(n8079), .Z(n8082) );
  XNOR U8687 ( .A(n8083), .B(n8082), .Z(n8084) );
  XNOR U8688 ( .A(n8085), .B(n8084), .Z(n8213) );
  XNOR U8689 ( .A(n8214), .B(n8213), .Z(n8215) );
  XOR U8690 ( .A(n8216), .B(n8215), .Z(n8222) );
  XNOR U8691 ( .A(n8220), .B(n8222), .Z(n8081) );
  XOR U8692 ( .A(n8219), .B(n8081), .Z(N185) );
  NANDN U8693 ( .A(n8083), .B(n8082), .Z(n8087) );
  NANDN U8694 ( .A(n8085), .B(n8084), .Z(n8086) );
  AND U8695 ( .A(n8087), .B(n8086), .Z(n8230) );
  NANDN U8696 ( .A(n8089), .B(n8088), .Z(n8093) );
  NAND U8697 ( .A(n8091), .B(n8090), .Z(n8092) );
  AND U8698 ( .A(n8093), .B(n8092), .Z(n8243) );
  NANDN U8699 ( .A(n8095), .B(n8094), .Z(n8099) );
  NAND U8700 ( .A(n8097), .B(n8096), .Z(n8098) );
  AND U8701 ( .A(n8099), .B(n8098), .Z(n8249) );
  NANDN U8702 ( .A(n8101), .B(n8100), .Z(n8105) );
  NAND U8703 ( .A(n8103), .B(n8102), .Z(n8104) );
  NAND U8704 ( .A(n8105), .B(n8104), .Z(n8248) );
  XNOR U8705 ( .A(n8249), .B(n8248), .Z(n8251) );
  NAND U8706 ( .A(x[149]), .B(y[712]), .Z(n9126) );
  NANDN U8707 ( .A(n9126), .B(n8106), .Z(n8110) );
  NAND U8708 ( .A(n8108), .B(n8107), .Z(n8109) );
  NAND U8709 ( .A(n8110), .B(n8109), .Z(n8355) );
  NAND U8710 ( .A(x[150]), .B(y[707]), .Z(n8324) );
  NAND U8711 ( .A(x[133]), .B(y[724]), .Z(n8323) );
  NAND U8712 ( .A(x[145]), .B(y[712]), .Z(n8322) );
  XOR U8713 ( .A(n8323), .B(n8322), .Z(n8325) );
  XOR U8714 ( .A(n8324), .B(n8325), .Z(n8354) );
  AND U8715 ( .A(y[709]), .B(x[148]), .Z(n8112) );
  NAND U8716 ( .A(y[708]), .B(x[149]), .Z(n8111) );
  XNOR U8717 ( .A(n8112), .B(n8111), .Z(n8337) );
  AND U8718 ( .A(x[147]), .B(y[710]), .Z(n8336) );
  XOR U8719 ( .A(n8337), .B(n8336), .Z(n8353) );
  XOR U8720 ( .A(n8355), .B(n8356), .Z(n8279) );
  NAND U8721 ( .A(n8500), .B(n8335), .Z(n8116) );
  NAND U8722 ( .A(n8114), .B(n8113), .Z(n8115) );
  NAND U8723 ( .A(n8116), .B(n8115), .Z(n8361) );
  NAND U8724 ( .A(x[143]), .B(y[714]), .Z(n8343) );
  NAND U8725 ( .A(x[146]), .B(y[711]), .Z(n8342) );
  NAND U8726 ( .A(x[134]), .B(y[723]), .Z(n8341) );
  XOR U8727 ( .A(n8342), .B(n8341), .Z(n8344) );
  XOR U8728 ( .A(n8343), .B(n8344), .Z(n8360) );
  NAND U8729 ( .A(x[151]), .B(y[706]), .Z(n8318) );
  NAND U8730 ( .A(x[132]), .B(y[725]), .Z(n8317) );
  NAND U8731 ( .A(x[144]), .B(y[713]), .Z(n8316) );
  XOR U8732 ( .A(n8317), .B(n8316), .Z(n8319) );
  XNOR U8733 ( .A(n8318), .B(n8319), .Z(n8359) );
  XOR U8734 ( .A(n8361), .B(n8362), .Z(n8278) );
  XNOR U8735 ( .A(n8279), .B(n8278), .Z(n8281) );
  NAND U8736 ( .A(n8118), .B(n8117), .Z(n8122) );
  NANDN U8737 ( .A(n8120), .B(n8119), .Z(n8121) );
  AND U8738 ( .A(n8122), .B(n8121), .Z(n8280) );
  XOR U8739 ( .A(n8281), .B(n8280), .Z(n8293) );
  NAND U8740 ( .A(n8124), .B(n8123), .Z(n8128) );
  NANDN U8741 ( .A(n8126), .B(n8125), .Z(n8127) );
  AND U8742 ( .A(n8128), .B(n8127), .Z(n8291) );
  NAND U8743 ( .A(n8130), .B(n8129), .Z(n8134) );
  NANDN U8744 ( .A(n8132), .B(n8131), .Z(n8133) );
  NAND U8745 ( .A(n8134), .B(n8133), .Z(n8290) );
  XNOR U8746 ( .A(n8291), .B(n8290), .Z(n8292) );
  XNOR U8747 ( .A(n8293), .B(n8292), .Z(n8250) );
  XNOR U8748 ( .A(n8251), .B(n8250), .Z(n8242) );
  NANDN U8749 ( .A(n8136), .B(n8135), .Z(n8140) );
  NAND U8750 ( .A(n8138), .B(n8137), .Z(n8139) );
  NAND U8751 ( .A(n8140), .B(n8139), .Z(n8244) );
  XOR U8752 ( .A(n8245), .B(n8244), .Z(n8239) );
  IV U8753 ( .A(n8141), .Z(n8260) );
  NANDN U8754 ( .A(n8260), .B(n8142), .Z(n8146) );
  NAND U8755 ( .A(n8144), .B(n8143), .Z(n8145) );
  AND U8756 ( .A(n8146), .B(n8145), .Z(n8285) );
  AND U8757 ( .A(x[142]), .B(y[720]), .Z(n9223) );
  NAND U8758 ( .A(n9223), .B(n8147), .Z(n8151) );
  NANDN U8759 ( .A(n8149), .B(n8148), .Z(n8150) );
  AND U8760 ( .A(n8151), .B(n8150), .Z(n8313) );
  NAND U8761 ( .A(x[139]), .B(y[718]), .Z(n8331) );
  NAND U8762 ( .A(x[140]), .B(y[717]), .Z(n8330) );
  NAND U8763 ( .A(x[135]), .B(y[722]), .Z(n8329) );
  XNOR U8764 ( .A(n8330), .B(n8329), .Z(n8332) );
  NAND U8765 ( .A(x[152]), .B(y[705]), .Z(n8328) );
  NAND U8766 ( .A(x[129]), .B(y[728]), .Z(n8299) );
  NAND U8767 ( .A(x[141]), .B(y[716]), .Z(n8301) );
  XOR U8768 ( .A(n8310), .B(n8311), .Z(n8312) );
  XNOR U8769 ( .A(n8285), .B(n8284), .Z(n8287) );
  NAND U8770 ( .A(n8153), .B(n8152), .Z(n8157) );
  AND U8771 ( .A(n8155), .B(n8154), .Z(n8156) );
  ANDN U8772 ( .B(n8157), .A(n8156), .Z(n8273) );
  AND U8773 ( .A(n8159), .B(n8158), .Z(n8163) );
  NAND U8774 ( .A(n8161), .B(n8160), .Z(n8162) );
  NANDN U8775 ( .A(n8163), .B(n8162), .Z(n8272) );
  XNOR U8776 ( .A(n8273), .B(n8272), .Z(n8275) );
  NAND U8777 ( .A(n8165), .B(n8164), .Z(n8169) );
  NAND U8778 ( .A(n8167), .B(n8166), .Z(n8168) );
  AND U8779 ( .A(n8169), .B(n8168), .Z(n8269) );
  AND U8780 ( .A(x[136]), .B(y[721]), .Z(n8263) );
  XNOR U8781 ( .A(n8261), .B(n8260), .Z(n8262) );
  XOR U8782 ( .A(n8263), .B(n8262), .Z(n8267) );
  AND U8783 ( .A(n8170), .B(o[88]), .Z(n8257) );
  AND U8784 ( .A(x[153]), .B(y[704]), .Z(n8255) );
  NAND U8785 ( .A(x[128]), .B(y[729]), .Z(n8254) );
  XNOR U8786 ( .A(n8255), .B(n8254), .Z(n8256) );
  XOR U8787 ( .A(n8257), .B(n8256), .Z(n8266) );
  XOR U8788 ( .A(n8267), .B(n8266), .Z(n8268) );
  XNOR U8789 ( .A(n8269), .B(n8268), .Z(n8274) );
  XOR U8790 ( .A(n8275), .B(n8274), .Z(n8286) );
  XOR U8791 ( .A(n8287), .B(n8286), .Z(n8368) );
  NAND U8792 ( .A(n8172), .B(n8171), .Z(n8176) );
  ANDN U8793 ( .B(n8174), .A(n8173), .Z(n8175) );
  ANDN U8794 ( .B(n8176), .A(n8175), .Z(n8350) );
  NAND U8795 ( .A(n8178), .B(n8177), .Z(n8182) );
  NAND U8796 ( .A(n8180), .B(n8179), .Z(n8181) );
  AND U8797 ( .A(n8182), .B(n8181), .Z(n8348) );
  AND U8798 ( .A(x[142]), .B(y[715]), .Z(n8304) );
  NAND U8799 ( .A(x[130]), .B(y[727]), .Z(n8305) );
  XNOR U8800 ( .A(n8304), .B(n8305), .Z(n8306) );
  NAND U8801 ( .A(x[131]), .B(y[726]), .Z(n8307) );
  XNOR U8802 ( .A(n8306), .B(n8307), .Z(n8347) );
  XNOR U8803 ( .A(n8348), .B(n8347), .Z(n8349) );
  XOR U8804 ( .A(n8350), .B(n8349), .Z(n8365) );
  NANDN U8805 ( .A(n8184), .B(n8183), .Z(n8188) );
  NAND U8806 ( .A(n8186), .B(n8185), .Z(n8187) );
  AND U8807 ( .A(n8188), .B(n8187), .Z(n8366) );
  XOR U8808 ( .A(n8365), .B(n8366), .Z(n8367) );
  NAND U8809 ( .A(n8190), .B(n8189), .Z(n8194) );
  NAND U8810 ( .A(n8192), .B(n8191), .Z(n8193) );
  NAND U8811 ( .A(n8194), .B(n8193), .Z(n8372) );
  XNOR U8812 ( .A(n8371), .B(n8372), .Z(n8374) );
  NANDN U8813 ( .A(n8196), .B(n8195), .Z(n8200) );
  NANDN U8814 ( .A(n8198), .B(n8197), .Z(n8199) );
  AND U8815 ( .A(n8200), .B(n8199), .Z(n8373) );
  XOR U8816 ( .A(n8374), .B(n8373), .Z(n8237) );
  NANDN U8817 ( .A(n8202), .B(n8201), .Z(n8206) );
  NANDN U8818 ( .A(n8204), .B(n8203), .Z(n8205) );
  AND U8819 ( .A(n8206), .B(n8205), .Z(n8236) );
  XNOR U8820 ( .A(n8237), .B(n8236), .Z(n8238) );
  XOR U8821 ( .A(n8239), .B(n8238), .Z(n8228) );
  NANDN U8822 ( .A(n8208), .B(n8207), .Z(n8212) );
  NAND U8823 ( .A(n8210), .B(n8209), .Z(n8211) );
  NAND U8824 ( .A(n8212), .B(n8211), .Z(n8227) );
  XOR U8825 ( .A(n8228), .B(n8227), .Z(n8229) );
  XOR U8826 ( .A(n8230), .B(n8229), .Z(n8235) );
  NANDN U8827 ( .A(n8214), .B(n8213), .Z(n8218) );
  NAND U8828 ( .A(n8216), .B(n8215), .Z(n8217) );
  NAND U8829 ( .A(n8218), .B(n8217), .Z(n8234) );
  NANDN U8830 ( .A(n8219), .B(n8220), .Z(n8225) );
  NOR U8831 ( .A(n8221), .B(n8220), .Z(n8223) );
  OR U8832 ( .A(n8223), .B(n8222), .Z(n8224) );
  AND U8833 ( .A(n8225), .B(n8224), .Z(n8233) );
  XOR U8834 ( .A(n8234), .B(n8233), .Z(n8226) );
  XNOR U8835 ( .A(n8235), .B(n8226), .Z(N186) );
  NAND U8836 ( .A(n8228), .B(n8227), .Z(n8232) );
  NAND U8837 ( .A(n8230), .B(n8229), .Z(n8231) );
  NAND U8838 ( .A(n8232), .B(n8231), .Z(n8534) );
  IV U8839 ( .A(n8534), .Z(n8532) );
  NANDN U8840 ( .A(n8237), .B(n8236), .Z(n8241) );
  NANDN U8841 ( .A(n8239), .B(n8238), .Z(n8240) );
  AND U8842 ( .A(n8241), .B(n8240), .Z(n8527) );
  NANDN U8843 ( .A(n8243), .B(n8242), .Z(n8247) );
  NAND U8844 ( .A(n8245), .B(n8244), .Z(n8246) );
  AND U8845 ( .A(n8247), .B(n8246), .Z(n8526) );
  XNOR U8846 ( .A(n8527), .B(n8526), .Z(n8529) );
  NANDN U8847 ( .A(n8249), .B(n8248), .Z(n8253) );
  NAND U8848 ( .A(n8251), .B(n8250), .Z(n8252) );
  AND U8849 ( .A(n8253), .B(n8252), .Z(n8387) );
  AND U8850 ( .A(x[130]), .B(y[728]), .Z(n8408) );
  XOR U8851 ( .A(n8409), .B(n8408), .Z(n8411) );
  NAND U8852 ( .A(x[152]), .B(y[706]), .Z(n8410) );
  NANDN U8853 ( .A(n8255), .B(n8254), .Z(n8259) );
  NANDN U8854 ( .A(n8257), .B(n8256), .Z(n8258) );
  AND U8855 ( .A(n8259), .B(n8258), .Z(n8444) );
  XOR U8856 ( .A(n8445), .B(n8444), .Z(n8447) );
  NANDN U8857 ( .A(n8261), .B(n8260), .Z(n8265) );
  NANDN U8858 ( .A(n8263), .B(n8262), .Z(n8264) );
  AND U8859 ( .A(n8265), .B(n8264), .Z(n8446) );
  XOR U8860 ( .A(n8447), .B(n8446), .Z(n8515) );
  NAND U8861 ( .A(n8267), .B(n8266), .Z(n8271) );
  NANDN U8862 ( .A(n8269), .B(n8268), .Z(n8270) );
  AND U8863 ( .A(n8271), .B(n8270), .Z(n8514) );
  NANDN U8864 ( .A(n8273), .B(n8272), .Z(n8277) );
  NAND U8865 ( .A(n8275), .B(n8274), .Z(n8276) );
  AND U8866 ( .A(n8277), .B(n8276), .Z(n8516) );
  XOR U8867 ( .A(n8517), .B(n8516), .Z(n8479) );
  NANDN U8868 ( .A(n8279), .B(n8278), .Z(n8283) );
  NAND U8869 ( .A(n8281), .B(n8280), .Z(n8282) );
  NAND U8870 ( .A(n8283), .B(n8282), .Z(n8476) );
  NANDN U8871 ( .A(n8285), .B(n8284), .Z(n8289) );
  NAND U8872 ( .A(n8287), .B(n8286), .Z(n8288) );
  AND U8873 ( .A(n8289), .B(n8288), .Z(n8477) );
  XOR U8874 ( .A(n8476), .B(n8477), .Z(n8478) );
  XOR U8875 ( .A(n8479), .B(n8478), .Z(n8385) );
  NANDN U8876 ( .A(n8291), .B(n8290), .Z(n8295) );
  NANDN U8877 ( .A(n8293), .B(n8292), .Z(n8294) );
  NAND U8878 ( .A(n8295), .B(n8294), .Z(n8392) );
  AND U8879 ( .A(x[140]), .B(y[718]), .Z(n8603) );
  AND U8880 ( .A(x[133]), .B(y[725]), .Z(n8459) );
  XOR U8881 ( .A(n8603), .B(n8459), .Z(n8461) );
  NAND U8882 ( .A(x[138]), .B(y[720]), .Z(n8460) );
  AND U8883 ( .A(x[135]), .B(y[723]), .Z(n8483) );
  AND U8884 ( .A(y[724]), .B(x[134]), .Z(n8297) );
  NAND U8885 ( .A(y[722]), .B(x[136]), .Z(n8296) );
  XNOR U8886 ( .A(n8297), .B(n8296), .Z(n8501) );
  NAND U8887 ( .A(x[137]), .B(y[721]), .Z(n8502) );
  XOR U8888 ( .A(n8483), .B(n8482), .Z(n8484) );
  XOR U8889 ( .A(n8485), .B(n8484), .Z(n8434) );
  NANDN U8890 ( .A(n8299), .B(n8298), .Z(n8303) );
  NANDN U8891 ( .A(n8301), .B(n8300), .Z(n8302) );
  NAND U8892 ( .A(n8303), .B(n8302), .Z(n8433) );
  NANDN U8893 ( .A(n8305), .B(n8304), .Z(n8309) );
  NANDN U8894 ( .A(n8307), .B(n8306), .Z(n8308) );
  NAND U8895 ( .A(n8309), .B(n8308), .Z(n8432) );
  XNOR U8896 ( .A(n8433), .B(n8432), .Z(n8435) );
  NAND U8897 ( .A(n8311), .B(n8310), .Z(n8315) );
  NANDN U8898 ( .A(n8313), .B(n8312), .Z(n8314) );
  AND U8899 ( .A(n8315), .B(n8314), .Z(n8470) );
  NAND U8900 ( .A(n8317), .B(n8316), .Z(n8321) );
  NAND U8901 ( .A(n8319), .B(n8318), .Z(n8320) );
  AND U8902 ( .A(n8321), .B(n8320), .Z(n8397) );
  NAND U8903 ( .A(n8323), .B(n8322), .Z(n8327) );
  NAND U8904 ( .A(n8325), .B(n8324), .Z(n8326) );
  AND U8905 ( .A(n8327), .B(n8326), .Z(n8396) );
  XOR U8906 ( .A(n8397), .B(n8396), .Z(n8399) );
  ANDN U8907 ( .B(o[89]), .A(n8328), .Z(n8494) );
  NAND U8908 ( .A(x[142]), .B(y[716]), .Z(n8495) );
  NAND U8909 ( .A(x[129]), .B(y[729]), .Z(n8497) );
  NAND U8910 ( .A(x[153]), .B(y[705]), .Z(n8505) );
  XNOR U8911 ( .A(o[90]), .B(n8505), .Z(n8464) );
  NAND U8912 ( .A(x[154]), .B(y[704]), .Z(n8465) );
  AND U8913 ( .A(x[128]), .B(y[730]), .Z(n8466) );
  XOR U8914 ( .A(n8467), .B(n8466), .Z(n8450) );
  XOR U8915 ( .A(n8451), .B(n8450), .Z(n8453) );
  NAND U8916 ( .A(n8330), .B(n8329), .Z(n8334) );
  NANDN U8917 ( .A(n8332), .B(n8331), .Z(n8333) );
  AND U8918 ( .A(n8334), .B(n8333), .Z(n8452) );
  XOR U8919 ( .A(n8453), .B(n8452), .Z(n8398) );
  XNOR U8920 ( .A(n8399), .B(n8398), .Z(n8440) );
  AND U8921 ( .A(x[149]), .B(y[709]), .Z(n8340) );
  IV U8922 ( .A(n8340), .Z(n8489) );
  NANDN U8923 ( .A(n8489), .B(n8335), .Z(n8339) );
  NAND U8924 ( .A(n8337), .B(n8336), .Z(n8338) );
  NAND U8925 ( .A(n8339), .B(n8338), .Z(n8428) );
  XOR U8926 ( .A(n8488), .B(n8340), .Z(n8491) );
  NAND U8927 ( .A(x[148]), .B(y[710]), .Z(n8490) );
  NAND U8928 ( .A(x[151]), .B(y[707]), .Z(n8415) );
  AND U8929 ( .A(x[150]), .B(y[708]), .Z(n8416) );
  XOR U8930 ( .A(n8417), .B(n8416), .Z(n8426) );
  XOR U8931 ( .A(n8427), .B(n8426), .Z(n8429) );
  XOR U8932 ( .A(n8428), .B(n8429), .Z(n8439) );
  AND U8933 ( .A(x[147]), .B(y[711]), .Z(n8506) );
  NAND U8934 ( .A(x[131]), .B(y[727]), .Z(n8507) );
  NAND U8935 ( .A(x[139]), .B(y[719]), .Z(n8509) );
  NAND U8936 ( .A(x[132]), .B(y[726]), .Z(n8421) );
  XOR U8937 ( .A(n8423), .B(n8422), .Z(n8402) );
  XOR U8938 ( .A(n8403), .B(n8402), .Z(n8405) );
  NAND U8939 ( .A(n8342), .B(n8341), .Z(n8346) );
  NAND U8940 ( .A(n8344), .B(n8343), .Z(n8345) );
  AND U8941 ( .A(n8346), .B(n8345), .Z(n8404) );
  XNOR U8942 ( .A(n8405), .B(n8404), .Z(n8438) );
  XOR U8943 ( .A(n8440), .B(n8441), .Z(n8473) );
  XNOR U8944 ( .A(n8472), .B(n8473), .Z(n8391) );
  NANDN U8945 ( .A(n8348), .B(n8347), .Z(n8352) );
  NANDN U8946 ( .A(n8350), .B(n8349), .Z(n8351) );
  NAND U8947 ( .A(n8352), .B(n8351), .Z(n8522) );
  NANDN U8948 ( .A(n8354), .B(n8353), .Z(n8358) );
  NAND U8949 ( .A(n8356), .B(n8355), .Z(n8357) );
  NAND U8950 ( .A(n8358), .B(n8357), .Z(n8521) );
  NANDN U8951 ( .A(n8360), .B(n8359), .Z(n8364) );
  NANDN U8952 ( .A(n8362), .B(n8361), .Z(n8363) );
  NAND U8953 ( .A(n8364), .B(n8363), .Z(n8520) );
  XOR U8954 ( .A(n8521), .B(n8520), .Z(n8523) );
  XOR U8955 ( .A(n8522), .B(n8523), .Z(n8390) );
  XOR U8956 ( .A(n8392), .B(n8393), .Z(n8384) );
  XNOR U8957 ( .A(n8385), .B(n8384), .Z(n8386) );
  XNOR U8958 ( .A(n8387), .B(n8386), .Z(n8381) );
  NAND U8959 ( .A(n8366), .B(n8365), .Z(n8370) );
  NANDN U8960 ( .A(n8368), .B(n8367), .Z(n8369) );
  AND U8961 ( .A(n8370), .B(n8369), .Z(n8378) );
  NANDN U8962 ( .A(n8372), .B(n8371), .Z(n8376) );
  NAND U8963 ( .A(n8374), .B(n8373), .Z(n8375) );
  NAND U8964 ( .A(n8376), .B(n8375), .Z(n8379) );
  XNOR U8965 ( .A(n8378), .B(n8379), .Z(n8380) );
  XOR U8966 ( .A(n8381), .B(n8380), .Z(n8528) );
  XOR U8967 ( .A(n8529), .B(n8528), .Z(n8535) );
  XNOR U8968 ( .A(n8533), .B(n8535), .Z(n8377) );
  XOR U8969 ( .A(n8532), .B(n8377), .Z(N187) );
  NANDN U8970 ( .A(n8379), .B(n8378), .Z(n8383) );
  NAND U8971 ( .A(n8381), .B(n8380), .Z(n8382) );
  AND U8972 ( .A(n8383), .B(n8382), .Z(n8543) );
  NANDN U8973 ( .A(n8385), .B(n8384), .Z(n8389) );
  NANDN U8974 ( .A(n8387), .B(n8386), .Z(n8388) );
  AND U8975 ( .A(n8389), .B(n8388), .Z(n8541) );
  NANDN U8976 ( .A(n8391), .B(n8390), .Z(n8395) );
  NAND U8977 ( .A(n8393), .B(n8392), .Z(n8394) );
  NAND U8978 ( .A(n8395), .B(n8394), .Z(n8551) );
  NAND U8979 ( .A(n8397), .B(n8396), .Z(n8401) );
  NAND U8980 ( .A(n8399), .B(n8398), .Z(n8400) );
  NAND U8981 ( .A(n8401), .B(n8400), .Z(n8674) );
  NAND U8982 ( .A(n8403), .B(n8402), .Z(n8407) );
  NAND U8983 ( .A(n8405), .B(n8404), .Z(n8406) );
  NAND U8984 ( .A(n8407), .B(n8406), .Z(n8672) );
  NAND U8985 ( .A(n8409), .B(n8408), .Z(n8413) );
  ANDN U8986 ( .B(n8411), .A(n8410), .Z(n8412) );
  ANDN U8987 ( .B(n8413), .A(n8412), .Z(n8574) );
  NANDN U8988 ( .A(n8415), .B(n8414), .Z(n8419) );
  NAND U8989 ( .A(n8417), .B(n8416), .Z(n8418) );
  NAND U8990 ( .A(n8419), .B(n8418), .Z(n8573) );
  NANDN U8991 ( .A(n8421), .B(n8420), .Z(n8425) );
  NAND U8992 ( .A(n8423), .B(n8422), .Z(n8424) );
  AND U8993 ( .A(n8425), .B(n8424), .Z(n8588) );
  AND U8994 ( .A(x[128]), .B(y[731]), .Z(n8651) );
  NAND U8995 ( .A(x[155]), .B(y[704]), .Z(n8652) );
  XNOR U8996 ( .A(n8651), .B(n8652), .Z(n8653) );
  NAND U8997 ( .A(x[154]), .B(y[705]), .Z(n8663) );
  XOR U8998 ( .A(o[91]), .B(n8663), .Z(n8654) );
  XNOR U8999 ( .A(n8653), .B(n8654), .Z(n8585) );
  AND U9000 ( .A(x[137]), .B(y[722]), .Z(n8657) );
  NAND U9001 ( .A(x[149]), .B(y[710]), .Z(n8658) );
  XNOR U9002 ( .A(n8657), .B(n8658), .Z(n8659) );
  NAND U9003 ( .A(x[146]), .B(y[713]), .Z(n8660) );
  XOR U9004 ( .A(n8659), .B(n8660), .Z(n8586) );
  XOR U9005 ( .A(n8576), .B(n8575), .Z(n8673) );
  XOR U9006 ( .A(n8672), .B(n8673), .Z(n8675) );
  XOR U9007 ( .A(n8674), .B(n8675), .Z(n8693) );
  NAND U9008 ( .A(n8427), .B(n8426), .Z(n8431) );
  NAND U9009 ( .A(n8429), .B(n8428), .Z(n8430) );
  AND U9010 ( .A(n8431), .B(n8430), .Z(n8691) );
  NAND U9011 ( .A(n8433), .B(n8432), .Z(n8437) );
  NANDN U9012 ( .A(n8435), .B(n8434), .Z(n8436) );
  AND U9013 ( .A(n8437), .B(n8436), .Z(n8690) );
  XOR U9014 ( .A(n8691), .B(n8690), .Z(n8692) );
  NANDN U9015 ( .A(n8439), .B(n8438), .Z(n8443) );
  NANDN U9016 ( .A(n8441), .B(n8440), .Z(n8442) );
  AND U9017 ( .A(n8443), .B(n8442), .Z(n8678) );
  NAND U9018 ( .A(n8445), .B(n8444), .Z(n8449) );
  NAND U9019 ( .A(n8447), .B(n8446), .Z(n8448) );
  NAND U9020 ( .A(n8449), .B(n8448), .Z(n8668) );
  NAND U9021 ( .A(n8451), .B(n8450), .Z(n8455) );
  NAND U9022 ( .A(n8453), .B(n8452), .Z(n8454) );
  NAND U9023 ( .A(n8455), .B(n8454), .Z(n8666) );
  AND U9024 ( .A(x[147]), .B(y[712]), .Z(n8639) );
  NAND U9025 ( .A(x[153]), .B(y[706]), .Z(n8640) );
  XNOR U9026 ( .A(n8639), .B(n8640), .Z(n8641) );
  NAND U9027 ( .A(x[134]), .B(y[725]), .Z(n8642) );
  XNOR U9028 ( .A(n8641), .B(n8642), .Z(n8628) );
  AND U9029 ( .A(x[143]), .B(y[716]), .Z(n8606) );
  NAND U9030 ( .A(x[130]), .B(y[729]), .Z(n8607) );
  XNOR U9031 ( .A(n8606), .B(n8607), .Z(n8608) );
  NAND U9032 ( .A(x[131]), .B(y[728]), .Z(n8609) );
  XOR U9033 ( .A(n8608), .B(n8609), .Z(n8629) );
  AND U9034 ( .A(x[144]), .B(y[715]), .Z(n8592) );
  XOR U9035 ( .A(n8592), .B(n8456), .Z(n8593) );
  XOR U9036 ( .A(n8594), .B(n8593), .Z(n8604) );
  AND U9037 ( .A(y[718]), .B(x[141]), .Z(n8458) );
  NAND U9038 ( .A(y[719]), .B(x[140]), .Z(n8457) );
  XNOR U9039 ( .A(n8458), .B(n8457), .Z(n8605) );
  XOR U9040 ( .A(n8604), .B(n8605), .Z(n8630) );
  XOR U9041 ( .A(n8631), .B(n8630), .Z(n8570) );
  NAND U9042 ( .A(n8603), .B(n8459), .Z(n8463) );
  ANDN U9043 ( .B(n8461), .A(n8460), .Z(n8462) );
  ANDN U9044 ( .B(n8463), .A(n8462), .Z(n8568) );
  NANDN U9045 ( .A(n8465), .B(n8464), .Z(n8469) );
  NAND U9046 ( .A(n8467), .B(n8466), .Z(n8468) );
  NAND U9047 ( .A(n8469), .B(n8468), .Z(n8567) );
  XOR U9048 ( .A(n8570), .B(n8569), .Z(n8667) );
  XNOR U9049 ( .A(n8666), .B(n8667), .Z(n8669) );
  XNOR U9050 ( .A(n8678), .B(n8679), .Z(n8681) );
  NANDN U9051 ( .A(n8471), .B(n8470), .Z(n8475) );
  NANDN U9052 ( .A(n8473), .B(n8472), .Z(n8474) );
  AND U9053 ( .A(n8475), .B(n8474), .Z(n8680) );
  XOR U9054 ( .A(n8681), .B(n8680), .Z(n8549) );
  XOR U9055 ( .A(n8551), .B(n8552), .Z(n8558) );
  NAND U9056 ( .A(n8477), .B(n8476), .Z(n8481) );
  NAND U9057 ( .A(n8479), .B(n8478), .Z(n8480) );
  NAND U9058 ( .A(n8481), .B(n8480), .Z(n8555) );
  NAND U9059 ( .A(n8483), .B(n8482), .Z(n8487) );
  NAND U9060 ( .A(n8485), .B(n8484), .Z(n8486) );
  NAND U9061 ( .A(n8487), .B(n8486), .Z(n8686) );
  NANDN U9062 ( .A(n8489), .B(n8488), .Z(n8493) );
  ANDN U9063 ( .B(n8491), .A(n8490), .Z(n8492) );
  ANDN U9064 ( .B(n8493), .A(n8492), .Z(n8617) );
  NANDN U9065 ( .A(n8495), .B(n8494), .Z(n8499) );
  NANDN U9066 ( .A(n8497), .B(n8496), .Z(n8498) );
  NAND U9067 ( .A(n8499), .B(n8498), .Z(n8616) );
  AND U9068 ( .A(x[136]), .B(y[724]), .Z(n8665) );
  NAND U9069 ( .A(n8500), .B(n8665), .Z(n8504) );
  NANDN U9070 ( .A(n8502), .B(n8501), .Z(n8503) );
  NAND U9071 ( .A(n8504), .B(n8503), .Z(n8581) );
  AND U9072 ( .A(x[142]), .B(y[717]), .Z(n8612) );
  NAND U9073 ( .A(x[129]), .B(y[730]), .Z(n8613) );
  XNOR U9074 ( .A(n8612), .B(n8613), .Z(n8615) );
  ANDN U9075 ( .B(o[90]), .A(n8505), .Z(n8614) );
  XOR U9076 ( .A(n8615), .B(n8614), .Z(n8580) );
  AND U9077 ( .A(x[145]), .B(y[714]), .Z(n8645) );
  NAND U9078 ( .A(x[132]), .B(y[727]), .Z(n8646) );
  XNOR U9079 ( .A(n8645), .B(n8646), .Z(n8648) );
  AND U9080 ( .A(x[133]), .B(y[726]), .Z(n8647) );
  XOR U9081 ( .A(n8648), .B(n8647), .Z(n8579) );
  XOR U9082 ( .A(n8580), .B(n8579), .Z(n8582) );
  XOR U9083 ( .A(n8581), .B(n8582), .Z(n8618) );
  XOR U9084 ( .A(n8619), .B(n8618), .Z(n8684) );
  NANDN U9085 ( .A(n8507), .B(n8506), .Z(n8511) );
  NANDN U9086 ( .A(n8509), .B(n8508), .Z(n8510) );
  AND U9087 ( .A(n8511), .B(n8510), .Z(n8625) );
  NAND U9088 ( .A(y[707]), .B(x[152]), .Z(n8512) );
  XNOR U9089 ( .A(n8513), .B(n8512), .Z(n8635) );
  NAND U9090 ( .A(x[135]), .B(y[724]), .Z(n8636) );
  XNOR U9091 ( .A(n8635), .B(n8636), .Z(n8622) );
  AND U9092 ( .A(x[136]), .B(y[723]), .Z(n8597) );
  NAND U9093 ( .A(x[151]), .B(y[708]), .Z(n8598) );
  XNOR U9094 ( .A(n8597), .B(n8598), .Z(n8599) );
  NAND U9095 ( .A(x[150]), .B(y[709]), .Z(n8600) );
  XOR U9096 ( .A(n8599), .B(n8600), .Z(n8623) );
  XNOR U9097 ( .A(n8684), .B(n8685), .Z(n8687) );
  XOR U9098 ( .A(n8686), .B(n8687), .Z(n8562) );
  NANDN U9099 ( .A(n8515), .B(n8514), .Z(n8519) );
  NAND U9100 ( .A(n8517), .B(n8516), .Z(n8518) );
  NAND U9101 ( .A(n8519), .B(n8518), .Z(n8561) );
  NAND U9102 ( .A(n8521), .B(n8520), .Z(n8525) );
  NAND U9103 ( .A(n8523), .B(n8522), .Z(n8524) );
  AND U9104 ( .A(n8525), .B(n8524), .Z(n8563) );
  XOR U9105 ( .A(n8564), .B(n8563), .Z(n8556) );
  XOR U9106 ( .A(n8555), .B(n8556), .Z(n8557) );
  XOR U9107 ( .A(n8541), .B(n8540), .Z(n8542) );
  XOR U9108 ( .A(n8543), .B(n8542), .Z(n8548) );
  NANDN U9109 ( .A(n8527), .B(n8526), .Z(n8531) );
  NAND U9110 ( .A(n8529), .B(n8528), .Z(n8530) );
  NAND U9111 ( .A(n8531), .B(n8530), .Z(n8547) );
  NANDN U9112 ( .A(n8532), .B(n8533), .Z(n8538) );
  NOR U9113 ( .A(n8534), .B(n8533), .Z(n8536) );
  OR U9114 ( .A(n8536), .B(n8535), .Z(n8537) );
  AND U9115 ( .A(n8538), .B(n8537), .Z(n8546) );
  XOR U9116 ( .A(n8547), .B(n8546), .Z(n8539) );
  XNOR U9117 ( .A(n8548), .B(n8539), .Z(N188) );
  NAND U9118 ( .A(n8541), .B(n8540), .Z(n8545) );
  NAND U9119 ( .A(n8543), .B(n8542), .Z(n8544) );
  NAND U9120 ( .A(n8545), .B(n8544), .Z(n8705) );
  IV U9121 ( .A(n8705), .Z(n8703) );
  NANDN U9122 ( .A(n8550), .B(n8549), .Z(n8554) );
  NAND U9123 ( .A(n8552), .B(n8551), .Z(n8553) );
  NAND U9124 ( .A(n8554), .B(n8553), .Z(n8697) );
  NAND U9125 ( .A(n8556), .B(n8555), .Z(n8560) );
  NANDN U9126 ( .A(n8558), .B(n8557), .Z(n8559) );
  AND U9127 ( .A(n8560), .B(n8559), .Z(n8698) );
  XOR U9128 ( .A(n8697), .B(n8698), .Z(n8700) );
  NANDN U9129 ( .A(n8562), .B(n8561), .Z(n8566) );
  NAND U9130 ( .A(n8564), .B(n8563), .Z(n8565) );
  AND U9131 ( .A(n8566), .B(n8565), .Z(n8710) );
  NANDN U9132 ( .A(n8568), .B(n8567), .Z(n8572) );
  NAND U9133 ( .A(n8570), .B(n8569), .Z(n8571) );
  AND U9134 ( .A(n8572), .B(n8571), .Z(n8735) );
  NANDN U9135 ( .A(n8574), .B(n8573), .Z(n8578) );
  NAND U9136 ( .A(n8576), .B(n8575), .Z(n8577) );
  AND U9137 ( .A(n8578), .B(n8577), .Z(n8838) );
  NAND U9138 ( .A(n8580), .B(n8579), .Z(n8584) );
  NAND U9139 ( .A(n8582), .B(n8581), .Z(n8583) );
  AND U9140 ( .A(n8584), .B(n8583), .Z(n8836) );
  NANDN U9141 ( .A(n8586), .B(n8585), .Z(n8590) );
  NANDN U9142 ( .A(n8588), .B(n8587), .Z(n8589) );
  NAND U9143 ( .A(n8590), .B(n8589), .Z(n8835) );
  NANDN U9144 ( .A(n8592), .B(n8591), .Z(n8596) );
  NANDN U9145 ( .A(n8594), .B(n8593), .Z(n8595) );
  AND U9146 ( .A(n8596), .B(n8595), .Z(n8801) );
  AND U9147 ( .A(x[135]), .B(y[725]), .Z(n8793) );
  NAND U9148 ( .A(x[140]), .B(y[720]), .Z(n8794) );
  XNOR U9149 ( .A(n8793), .B(n8794), .Z(n8796) );
  AND U9150 ( .A(x[139]), .B(y[721]), .Z(n8795) );
  XOR U9151 ( .A(n8796), .B(n8795), .Z(n8800) );
  NAND U9152 ( .A(x[155]), .B(y[705]), .Z(n8780) );
  XNOR U9153 ( .A(o[92]), .B(n8780), .Z(n8811) );
  NAND U9154 ( .A(x[154]), .B(y[706]), .Z(n8812) );
  XNOR U9155 ( .A(n8811), .B(n8812), .Z(n8814) );
  AND U9156 ( .A(x[143]), .B(y[717]), .Z(n8813) );
  XNOR U9157 ( .A(n8814), .B(n8813), .Z(n8799) );
  XOR U9158 ( .A(n8800), .B(n8799), .Z(n8802) );
  XOR U9159 ( .A(n8801), .B(n8802), .Z(n8842) );
  NANDN U9160 ( .A(n8598), .B(n8597), .Z(n8602) );
  NANDN U9161 ( .A(n8600), .B(n8599), .Z(n8601) );
  AND U9162 ( .A(n8602), .B(n8601), .Z(n8822) );
  AND U9163 ( .A(x[145]), .B(y[715]), .Z(n8746) );
  NAND U9164 ( .A(x[150]), .B(y[710]), .Z(n8747) );
  XNOR U9165 ( .A(n8746), .B(n8747), .Z(n8748) );
  NAND U9166 ( .A(x[132]), .B(y[728]), .Z(n8749) );
  XNOR U9167 ( .A(n8748), .B(n8749), .Z(n8820) );
  AND U9168 ( .A(x[134]), .B(y[726]), .Z(n8946) );
  NAND U9169 ( .A(x[147]), .B(y[713]), .Z(n8769) );
  XNOR U9170 ( .A(n8946), .B(n8769), .Z(n8770) );
  XOR U9171 ( .A(n8820), .B(n8819), .Z(n8821) );
  XNOR U9172 ( .A(n8822), .B(n8821), .Z(n8841) );
  NANDN U9173 ( .A(n8607), .B(n8606), .Z(n8611) );
  NANDN U9174 ( .A(n8609), .B(n8608), .Z(n8610) );
  AND U9175 ( .A(n8611), .B(n8610), .Z(n8741) );
  XNOR U9176 ( .A(n8741), .B(n8740), .Z(n8742) );
  XOR U9177 ( .A(n8743), .B(n8742), .Z(n8844) );
  XNOR U9178 ( .A(n8737), .B(n8736), .Z(n8731) );
  NANDN U9179 ( .A(n8617), .B(n8616), .Z(n8621) );
  NAND U9180 ( .A(n8619), .B(n8618), .Z(n8620) );
  AND U9181 ( .A(n8621), .B(n8620), .Z(n8826) );
  NANDN U9182 ( .A(n8623), .B(n8622), .Z(n8627) );
  NANDN U9183 ( .A(n8625), .B(n8624), .Z(n8626) );
  AND U9184 ( .A(n8627), .B(n8626), .Z(n8824) );
  NANDN U9185 ( .A(n8629), .B(n8628), .Z(n8633) );
  NAND U9186 ( .A(n8631), .B(n8630), .Z(n8632) );
  NAND U9187 ( .A(n8633), .B(n8632), .Z(n8823) );
  AND U9188 ( .A(x[152]), .B(y[711]), .Z(n9146) );
  NAND U9189 ( .A(n9146), .B(n8634), .Z(n8638) );
  NANDN U9190 ( .A(n8636), .B(n8635), .Z(n8637) );
  AND U9191 ( .A(n8638), .B(n8637), .Z(n8861) );
  AND U9192 ( .A(x[153]), .B(y[707]), .Z(n8789) );
  XOR U9193 ( .A(n8790), .B(n8789), .Z(n8788) );
  NAND U9194 ( .A(x[129]), .B(y[731]), .Z(n8787) );
  XNOR U9195 ( .A(n8788), .B(n8787), .Z(n8859) );
  AND U9196 ( .A(x[144]), .B(y[716]), .Z(n8781) );
  NAND U9197 ( .A(x[152]), .B(y[708]), .Z(n8782) );
  XNOR U9198 ( .A(n8781), .B(n8782), .Z(n8783) );
  NAND U9199 ( .A(x[130]), .B(y[730]), .Z(n8784) );
  XOR U9200 ( .A(n8783), .B(n8784), .Z(n8860) );
  XOR U9201 ( .A(n8859), .B(n8860), .Z(n8862) );
  XOR U9202 ( .A(n8861), .B(n8862), .Z(n8832) );
  NANDN U9203 ( .A(n8640), .B(n8639), .Z(n8644) );
  NANDN U9204 ( .A(n8642), .B(n8641), .Z(n8643) );
  AND U9205 ( .A(n8644), .B(n8643), .Z(n8855) );
  NAND U9206 ( .A(x[131]), .B(y[729]), .Z(n8806) );
  XNOR U9207 ( .A(n8805), .B(n8806), .Z(n8807) );
  NAND U9208 ( .A(x[151]), .B(y[709]), .Z(n8808) );
  XNOR U9209 ( .A(n8807), .B(n8808), .Z(n8853) );
  AND U9210 ( .A(x[133]), .B(y[727]), .Z(n8774) );
  NAND U9211 ( .A(x[149]), .B(y[711]), .Z(n8775) );
  XNOR U9212 ( .A(n8774), .B(n8775), .Z(n8776) );
  NAND U9213 ( .A(x[148]), .B(y[712]), .Z(n8777) );
  XOR U9214 ( .A(n8776), .B(n8777), .Z(n8854) );
  XOR U9215 ( .A(n8853), .B(n8854), .Z(n8856) );
  XOR U9216 ( .A(n8855), .B(n8856), .Z(n8830) );
  NANDN U9217 ( .A(n8646), .B(n8645), .Z(n8650) );
  NAND U9218 ( .A(n8648), .B(n8647), .Z(n8649) );
  AND U9219 ( .A(n8650), .B(n8649), .Z(n8848) );
  NANDN U9220 ( .A(n8652), .B(n8651), .Z(n8656) );
  NANDN U9221 ( .A(n8654), .B(n8653), .Z(n8655) );
  NAND U9222 ( .A(n8656), .B(n8655), .Z(n8847) );
  XNOR U9223 ( .A(n8848), .B(n8847), .Z(n8850) );
  NANDN U9224 ( .A(n8658), .B(n8657), .Z(n8662) );
  NANDN U9225 ( .A(n8660), .B(n8659), .Z(n8661) );
  AND U9226 ( .A(n8662), .B(n8661), .Z(n8766) );
  ANDN U9227 ( .B(o[91]), .A(n8663), .Z(n8754) );
  AND U9228 ( .A(x[128]), .B(y[732]), .Z(n8752) );
  NAND U9229 ( .A(x[156]), .B(y[704]), .Z(n8753) );
  XOR U9230 ( .A(n8752), .B(n8753), .Z(n8755) );
  XNOR U9231 ( .A(n8754), .B(n8755), .Z(n8763) );
  NAND U9232 ( .A(y[722]), .B(x[138]), .Z(n8664) );
  XNOR U9233 ( .A(n8665), .B(n8664), .Z(n8759) );
  NAND U9234 ( .A(x[137]), .B(y[723]), .Z(n8760) );
  XOR U9235 ( .A(n8759), .B(n8760), .Z(n8764) );
  XNOR U9236 ( .A(n8763), .B(n8764), .Z(n8765) );
  XNOR U9237 ( .A(n8766), .B(n8765), .Z(n8849) );
  XNOR U9238 ( .A(n8850), .B(n8849), .Z(n8829) );
  XNOR U9239 ( .A(n8731), .B(n8730), .Z(n8724) );
  NAND U9240 ( .A(n8667), .B(n8666), .Z(n8671) );
  NANDN U9241 ( .A(n8669), .B(n8668), .Z(n8670) );
  NAND U9242 ( .A(n8671), .B(n8670), .Z(n8723) );
  NAND U9243 ( .A(n8673), .B(n8672), .Z(n8677) );
  NAND U9244 ( .A(n8675), .B(n8674), .Z(n8676) );
  NAND U9245 ( .A(n8677), .B(n8676), .Z(n8722) );
  XNOR U9246 ( .A(n8723), .B(n8722), .Z(n8725) );
  XNOR U9247 ( .A(n8710), .B(n8711), .Z(n8713) );
  NANDN U9248 ( .A(n8679), .B(n8678), .Z(n8683) );
  NAND U9249 ( .A(n8681), .B(n8680), .Z(n8682) );
  NAND U9250 ( .A(n8683), .B(n8682), .Z(n8718) );
  NANDN U9251 ( .A(n8685), .B(n8684), .Z(n8689) );
  NAND U9252 ( .A(n8687), .B(n8686), .Z(n8688) );
  NAND U9253 ( .A(n8689), .B(n8688), .Z(n8716) );
  NAND U9254 ( .A(n8691), .B(n8690), .Z(n8695) );
  NANDN U9255 ( .A(n8693), .B(n8692), .Z(n8694) );
  AND U9256 ( .A(n8695), .B(n8694), .Z(n8717) );
  XOR U9257 ( .A(n8716), .B(n8717), .Z(n8719) );
  XOR U9258 ( .A(n8718), .B(n8719), .Z(n8712) );
  XOR U9259 ( .A(n8713), .B(n8712), .Z(n8699) );
  XOR U9260 ( .A(n8700), .B(n8699), .Z(n8706) );
  XNOR U9261 ( .A(n8704), .B(n8706), .Z(n8696) );
  XOR U9262 ( .A(n8703), .B(n8696), .Z(N189) );
  NAND U9263 ( .A(n8698), .B(n8697), .Z(n8702) );
  NAND U9264 ( .A(n8700), .B(n8699), .Z(n8701) );
  AND U9265 ( .A(n8702), .B(n8701), .Z(n8866) );
  NANDN U9266 ( .A(n8703), .B(n8704), .Z(n8709) );
  NOR U9267 ( .A(n8705), .B(n8704), .Z(n8707) );
  OR U9268 ( .A(n8707), .B(n8706), .Z(n8708) );
  AND U9269 ( .A(n8709), .B(n8708), .Z(n8867) );
  NANDN U9270 ( .A(n8711), .B(n8710), .Z(n8715) );
  NAND U9271 ( .A(n8713), .B(n8712), .Z(n8714) );
  NAND U9272 ( .A(n8715), .B(n8714), .Z(n8871) );
  NAND U9273 ( .A(n8717), .B(n8716), .Z(n8721) );
  NAND U9274 ( .A(n8719), .B(n8718), .Z(n8720) );
  NAND U9275 ( .A(n8721), .B(n8720), .Z(n8869) );
  NAND U9276 ( .A(n8723), .B(n8722), .Z(n8727) );
  NANDN U9277 ( .A(n8725), .B(n8724), .Z(n8726) );
  NAND U9278 ( .A(n8727), .B(n8726), .Z(n8875) );
  NANDN U9279 ( .A(n8729), .B(n8728), .Z(n8733) );
  NAND U9280 ( .A(n8731), .B(n8730), .Z(n8732) );
  AND U9281 ( .A(n8733), .B(n8732), .Z(n8876) );
  XOR U9282 ( .A(n8875), .B(n8876), .Z(n8878) );
  NANDN U9283 ( .A(n8735), .B(n8734), .Z(n8739) );
  NAND U9284 ( .A(n8737), .B(n8736), .Z(n8738) );
  AND U9285 ( .A(n8739), .B(n8738), .Z(n8888) );
  NANDN U9286 ( .A(n8741), .B(n8740), .Z(n8745) );
  NANDN U9287 ( .A(n8743), .B(n8742), .Z(n8744) );
  AND U9288 ( .A(n8745), .B(n8744), .Z(n8997) );
  NANDN U9289 ( .A(n8747), .B(n8746), .Z(n8751) );
  NANDN U9290 ( .A(n8749), .B(n8748), .Z(n8750) );
  AND U9291 ( .A(n8751), .B(n8750), .Z(n9034) );
  NANDN U9292 ( .A(n8753), .B(n8752), .Z(n8757) );
  NANDN U9293 ( .A(n8755), .B(n8754), .Z(n8756) );
  NAND U9294 ( .A(n8757), .B(n8756), .Z(n9033) );
  XNOR U9295 ( .A(n9034), .B(n9033), .Z(n9036) );
  AND U9296 ( .A(x[138]), .B(y[724]), .Z(n9031) );
  NAND U9297 ( .A(n8758), .B(n9031), .Z(n8762) );
  NANDN U9298 ( .A(n8760), .B(n8759), .Z(n8761) );
  AND U9299 ( .A(n8762), .B(n8761), .Z(n9003) );
  AND U9300 ( .A(x[150]), .B(y[711]), .Z(n8967) );
  AND U9301 ( .A(x[140]), .B(y[721]), .Z(n9085) );
  AND U9302 ( .A(x[129]), .B(y[732]), .Z(n8965) );
  XOR U9303 ( .A(n9085), .B(n8965), .Z(n8966) );
  XOR U9304 ( .A(n8967), .B(n8966), .Z(n9001) );
  AND U9305 ( .A(x[143]), .B(y[718]), .Z(n8968) );
  XOR U9306 ( .A(n9001), .B(n9000), .Z(n9002) );
  XOR U9307 ( .A(n9036), .B(n9035), .Z(n8995) );
  NANDN U9308 ( .A(n8764), .B(n8763), .Z(n8768) );
  NANDN U9309 ( .A(n8766), .B(n8765), .Z(n8767) );
  AND U9310 ( .A(n8768), .B(n8767), .Z(n8994) );
  XNOR U9311 ( .A(n8995), .B(n8994), .Z(n8996) );
  XOR U9312 ( .A(n8997), .B(n8996), .Z(n8991) );
  NANDN U9313 ( .A(n8769), .B(n8946), .Z(n8773) );
  NANDN U9314 ( .A(n8771), .B(n8770), .Z(n8772) );
  AND U9315 ( .A(n8773), .B(n8772), .Z(n9014) );
  AND U9316 ( .A(x[153]), .B(y[708]), .Z(n8962) );
  AND U9317 ( .A(x[154]), .B(y[707]), .Z(n8959) );
  XOR U9318 ( .A(n8960), .B(n8959), .Z(n8961) );
  XOR U9319 ( .A(n8962), .B(n8961), .Z(n9013) );
  NAND U9320 ( .A(x[156]), .B(y[705]), .Z(n8975) );
  XNOR U9321 ( .A(o[93]), .B(n8975), .Z(n9026) );
  AND U9322 ( .A(x[128]), .B(y[733]), .Z(n9024) );
  AND U9323 ( .A(x[157]), .B(y[704]), .Z(n9023) );
  XOR U9324 ( .A(n9024), .B(n9023), .Z(n9025) );
  XNOR U9325 ( .A(n9026), .B(n9025), .Z(n9012) );
  XNOR U9326 ( .A(n9014), .B(n9015), .Z(n8982) );
  NANDN U9327 ( .A(n8775), .B(n8774), .Z(n8779) );
  NANDN U9328 ( .A(n8777), .B(n8776), .Z(n8778) );
  AND U9329 ( .A(n8779), .B(n8778), .Z(n8956) );
  AND U9330 ( .A(x[130]), .B(y[731]), .Z(n8918) );
  XOR U9331 ( .A(n8918), .B(n8917), .Z(n8919) );
  XOR U9332 ( .A(n8920), .B(n8919), .Z(n8954) );
  ANDN U9333 ( .B(o[92]), .A(n8780), .Z(n8926) );
  AND U9334 ( .A(x[144]), .B(y[717]), .Z(n8924) );
  AND U9335 ( .A(x[155]), .B(y[706]), .Z(n8923) );
  XOR U9336 ( .A(n8924), .B(n8923), .Z(n8925) );
  XOR U9337 ( .A(n8926), .B(n8925), .Z(n8953) );
  XOR U9338 ( .A(n8954), .B(n8953), .Z(n8955) );
  XNOR U9339 ( .A(n8956), .B(n8955), .Z(n8983) );
  NANDN U9340 ( .A(n8782), .B(n8781), .Z(n8786) );
  NANDN U9341 ( .A(n8784), .B(n8783), .Z(n8785) );
  NAND U9342 ( .A(n8786), .B(n8785), .Z(n9007) );
  ANDN U9343 ( .B(n8788), .A(n8787), .Z(n8792) );
  NAND U9344 ( .A(n8790), .B(n8789), .Z(n8791) );
  NANDN U9345 ( .A(n8792), .B(n8791), .Z(n9006) );
  XOR U9346 ( .A(n9007), .B(n9006), .Z(n9008) );
  NANDN U9347 ( .A(n8794), .B(n8793), .Z(n8798) );
  NAND U9348 ( .A(n8796), .B(n8795), .Z(n8797) );
  AND U9349 ( .A(n8798), .B(n8797), .Z(n8908) );
  AND U9350 ( .A(x[139]), .B(y[722]), .Z(n8943) );
  AND U9351 ( .A(x[131]), .B(y[730]), .Z(n8940) );
  NAND U9352 ( .A(x[145]), .B(y[716]), .Z(n8941) );
  XOR U9353 ( .A(n8943), .B(n8942), .Z(n8906) );
  AND U9354 ( .A(x[151]), .B(y[710]), .Z(n8937) );
  AND U9355 ( .A(x[141]), .B(y[720]), .Z(n8935) );
  NAND U9356 ( .A(x[152]), .B(y[709]), .Z(n9090) );
  XOR U9357 ( .A(n8937), .B(n8936), .Z(n8905) );
  XOR U9358 ( .A(n8906), .B(n8905), .Z(n8907) );
  XOR U9359 ( .A(n8908), .B(n8907), .Z(n9009) );
  XNOR U9360 ( .A(n9008), .B(n9009), .Z(n8985) );
  NANDN U9361 ( .A(n8800), .B(n8799), .Z(n8804) );
  OR U9362 ( .A(n8802), .B(n8801), .Z(n8803) );
  AND U9363 ( .A(n8804), .B(n8803), .Z(n8900) );
  NANDN U9364 ( .A(n8806), .B(n8805), .Z(n8810) );
  NANDN U9365 ( .A(n8808), .B(n8807), .Z(n8809) );
  AND U9366 ( .A(n8810), .B(n8809), .Z(n8930) );
  NANDN U9367 ( .A(n8812), .B(n8811), .Z(n8816) );
  NAND U9368 ( .A(n8814), .B(n8813), .Z(n8815) );
  NAND U9369 ( .A(n8816), .B(n8815), .Z(n8929) );
  XNOR U9370 ( .A(n8930), .B(n8929), .Z(n8932) );
  AND U9371 ( .A(x[137]), .B(y[724]), .Z(n9121) );
  AND U9372 ( .A(x[136]), .B(y[725]), .Z(n8948) );
  AND U9373 ( .A(y[727]), .B(x[134]), .Z(n8818) );
  NAND U9374 ( .A(y[726]), .B(x[135]), .Z(n8817) );
  XNOR U9375 ( .A(n8818), .B(n8817), .Z(n8947) );
  XOR U9376 ( .A(n8948), .B(n8947), .Z(n9018) );
  XOR U9377 ( .A(n9121), .B(n9018), .Z(n9020) );
  AND U9378 ( .A(x[133]), .B(y[728]), .Z(n8914) );
  AND U9379 ( .A(x[132]), .B(y[729]), .Z(n8911) );
  NAND U9380 ( .A(x[138]), .B(y[723]), .Z(n8912) );
  XNOR U9381 ( .A(n8911), .B(n8912), .Z(n8913) );
  XOR U9382 ( .A(n8914), .B(n8913), .Z(n9019) );
  XOR U9383 ( .A(n9020), .B(n9019), .Z(n8931) );
  XNOR U9384 ( .A(n8932), .B(n8931), .Z(n8899) );
  XNOR U9385 ( .A(n8900), .B(n8899), .Z(n8901) );
  XOR U9386 ( .A(n8902), .B(n8901), .Z(n8989) );
  XNOR U9387 ( .A(n8989), .B(n8988), .Z(n8990) );
  XNOR U9388 ( .A(n8991), .B(n8990), .Z(n8887) );
  NANDN U9389 ( .A(n8824), .B(n8823), .Z(n8828) );
  NANDN U9390 ( .A(n8826), .B(n8825), .Z(n8827) );
  AND U9391 ( .A(n8828), .B(n8827), .Z(n8882) );
  NANDN U9392 ( .A(n8830), .B(n8829), .Z(n8834) );
  NANDN U9393 ( .A(n8832), .B(n8831), .Z(n8833) );
  AND U9394 ( .A(n8834), .B(n8833), .Z(n8881) );
  NANDN U9395 ( .A(n8836), .B(n8835), .Z(n8840) );
  NANDN U9396 ( .A(n8838), .B(n8837), .Z(n8839) );
  NAND U9397 ( .A(n8840), .B(n8839), .Z(n8895) );
  NANDN U9398 ( .A(n8842), .B(n8841), .Z(n8846) );
  NANDN U9399 ( .A(n8844), .B(n8843), .Z(n8845) );
  NAND U9400 ( .A(n8846), .B(n8845), .Z(n8893) );
  NANDN U9401 ( .A(n8848), .B(n8847), .Z(n8852) );
  NAND U9402 ( .A(n8850), .B(n8849), .Z(n8851) );
  AND U9403 ( .A(n8852), .B(n8851), .Z(n8979) );
  NANDN U9404 ( .A(n8854), .B(n8853), .Z(n8858) );
  OR U9405 ( .A(n8856), .B(n8855), .Z(n8857) );
  AND U9406 ( .A(n8858), .B(n8857), .Z(n8977) );
  NANDN U9407 ( .A(n8860), .B(n8859), .Z(n8864) );
  OR U9408 ( .A(n8862), .B(n8861), .Z(n8863) );
  NAND U9409 ( .A(n8864), .B(n8863), .Z(n8976) );
  XNOR U9410 ( .A(n8977), .B(n8976), .Z(n8978) );
  XNOR U9411 ( .A(n8979), .B(n8978), .Z(n8894) );
  XOR U9412 ( .A(n8893), .B(n8894), .Z(n8896) );
  XOR U9413 ( .A(n8895), .B(n8896), .Z(n8883) );
  XOR U9414 ( .A(n8884), .B(n8883), .Z(n8889) );
  XOR U9415 ( .A(n8890), .B(n8889), .Z(n8877) );
  XOR U9416 ( .A(n8878), .B(n8877), .Z(n8870) );
  XOR U9417 ( .A(n8869), .B(n8870), .Z(n8872) );
  XOR U9418 ( .A(n8871), .B(n8872), .Z(n8868) );
  XNOR U9419 ( .A(n8867), .B(n8868), .Z(n8865) );
  XOR U9420 ( .A(n8866), .B(n8865), .Z(N190) );
  NAND U9421 ( .A(n8870), .B(n8869), .Z(n8874) );
  NAND U9422 ( .A(n8872), .B(n8871), .Z(n8873) );
  AND U9423 ( .A(n8874), .B(n8873), .Z(n9291) );
  XNOR U9424 ( .A(n9292), .B(n9291), .Z(n9290) );
  NAND U9425 ( .A(n8876), .B(n8875), .Z(n8880) );
  NAND U9426 ( .A(n8878), .B(n8877), .Z(n8879) );
  NAND U9427 ( .A(n8880), .B(n8879), .Z(n9304) );
  NANDN U9428 ( .A(n8882), .B(n8881), .Z(n8886) );
  NAND U9429 ( .A(n8884), .B(n8883), .Z(n8885) );
  AND U9430 ( .A(n8886), .B(n8885), .Z(n9297) );
  NANDN U9431 ( .A(n8888), .B(n8887), .Z(n8892) );
  NAND U9432 ( .A(n8890), .B(n8889), .Z(n8891) );
  NAND U9433 ( .A(n8892), .B(n8891), .Z(n9298) );
  NAND U9434 ( .A(n8894), .B(n8893), .Z(n8898) );
  NAND U9435 ( .A(n8896), .B(n8895), .Z(n8897) );
  AND U9436 ( .A(n8898), .B(n8897), .Z(n9295) );
  XOR U9437 ( .A(n9296), .B(n9295), .Z(n9301) );
  NANDN U9438 ( .A(n8900), .B(n8899), .Z(n8904) );
  NAND U9439 ( .A(n8902), .B(n8901), .Z(n8903) );
  AND U9440 ( .A(n8904), .B(n8903), .Z(n9040) );
  NAND U9441 ( .A(n8906), .B(n8905), .Z(n8910) );
  NANDN U9442 ( .A(n8908), .B(n8907), .Z(n8909) );
  AND U9443 ( .A(n8910), .B(n8909), .Z(n9046) );
  NANDN U9444 ( .A(n8912), .B(n8911), .Z(n8916) );
  NAND U9445 ( .A(n8914), .B(n8913), .Z(n8915) );
  AND U9446 ( .A(n8916), .B(n8915), .Z(n9055) );
  AND U9447 ( .A(x[134]), .B(y[728]), .Z(n9094) );
  AND U9448 ( .A(x[133]), .B(y[729]), .Z(n9096) );
  AND U9449 ( .A(x[147]), .B(y[715]), .Z(n9095) );
  XOR U9450 ( .A(n9096), .B(n9095), .Z(n9093) );
  XNOR U9451 ( .A(n9094), .B(n9093), .Z(n9057) );
  AND U9452 ( .A(x[132]), .B(y[730]), .Z(n9130) );
  AND U9453 ( .A(x[131]), .B(y[731]), .Z(n9132) );
  AND U9454 ( .A(x[146]), .B(y[716]), .Z(n9131) );
  XOR U9455 ( .A(n9132), .B(n9131), .Z(n9129) );
  XOR U9456 ( .A(n9130), .B(n9129), .Z(n9060) );
  NAND U9457 ( .A(n8918), .B(n8917), .Z(n8922) );
  NAND U9458 ( .A(n8920), .B(n8919), .Z(n8921) );
  AND U9459 ( .A(n8922), .B(n8921), .Z(n9059) );
  XOR U9460 ( .A(n9057), .B(n9058), .Z(n9056) );
  XNOR U9461 ( .A(n9055), .B(n9056), .Z(n9054) );
  NAND U9462 ( .A(n8924), .B(n8923), .Z(n8928) );
  NAND U9463 ( .A(n8926), .B(n8925), .Z(n8927) );
  AND U9464 ( .A(n8928), .B(n8927), .Z(n9053) );
  XOR U9465 ( .A(n9054), .B(n9053), .Z(n9045) );
  XOR U9466 ( .A(n9046), .B(n9045), .Z(n9044) );
  NANDN U9467 ( .A(n8930), .B(n8929), .Z(n8934) );
  NAND U9468 ( .A(n8932), .B(n8931), .Z(n8933) );
  AND U9469 ( .A(n8934), .B(n8933), .Z(n9043) );
  XOR U9470 ( .A(n9044), .B(n9043), .Z(n9042) );
  NANDN U9471 ( .A(n9090), .B(n8935), .Z(n8939) );
  NAND U9472 ( .A(n8937), .B(n8936), .Z(n8938) );
  NAND U9473 ( .A(n8939), .B(n8938), .Z(n9050) );
  NANDN U9474 ( .A(n8941), .B(n8940), .Z(n8945) );
  NAND U9475 ( .A(n8943), .B(n8942), .Z(n8944) );
  AND U9476 ( .A(n8945), .B(n8944), .Z(n9240) );
  AND U9477 ( .A(x[128]), .B(y[734]), .Z(n9138) );
  AND U9478 ( .A(x[157]), .B(y[705]), .Z(n9143) );
  XOR U9479 ( .A(o[94]), .B(n9143), .Z(n9140) );
  AND U9480 ( .A(x[158]), .B(y[704]), .Z(n9139) );
  XOR U9481 ( .A(n9140), .B(n9139), .Z(n9137) );
  XOR U9482 ( .A(n9138), .B(n9137), .Z(n9242) );
  AND U9483 ( .A(x[148]), .B(y[714]), .Z(n9224) );
  XOR U9484 ( .A(n9224), .B(n9223), .Z(n9222) );
  AND U9485 ( .A(x[136]), .B(y[726]), .Z(n9221) );
  XNOR U9486 ( .A(n9222), .B(n9221), .Z(n9241) );
  XNOR U9487 ( .A(n9240), .B(n9239), .Z(n9049) );
  XOR U9488 ( .A(n9050), .B(n9049), .Z(n9047) );
  AND U9489 ( .A(x[135]), .B(y[727]), .Z(n9125) );
  NAND U9490 ( .A(n8946), .B(n9125), .Z(n8950) );
  NAND U9491 ( .A(n8948), .B(n8947), .Z(n8949) );
  AND U9492 ( .A(n8950), .B(n8949), .Z(n9233) );
  AND U9493 ( .A(y[713]), .B(x[149]), .Z(n8952) );
  AND U9494 ( .A(y[712]), .B(x[150]), .Z(n8951) );
  XOR U9495 ( .A(n8952), .B(n8951), .Z(n9124) );
  XOR U9496 ( .A(n9125), .B(n9124), .Z(n9236) );
  AND U9497 ( .A(x[145]), .B(y[717]), .Z(n9216) );
  AND U9498 ( .A(x[130]), .B(y[732]), .Z(n9218) );
  AND U9499 ( .A(x[154]), .B(y[708]), .Z(n9217) );
  XOR U9500 ( .A(n9218), .B(n9217), .Z(n9215) );
  XNOR U9501 ( .A(n9216), .B(n9215), .Z(n9235) );
  XNOR U9502 ( .A(n9233), .B(n9234), .Z(n9048) );
  NAND U9503 ( .A(n8954), .B(n8953), .Z(n8958) );
  NANDN U9504 ( .A(n8956), .B(n8955), .Z(n8957) );
  NAND U9505 ( .A(n8958), .B(n8957), .Z(n9271) );
  XOR U9506 ( .A(n9272), .B(n9271), .Z(n9269) );
  AND U9507 ( .A(n8960), .B(n8959), .Z(n8964) );
  NAND U9508 ( .A(n8962), .B(n8961), .Z(n8963) );
  NANDN U9509 ( .A(n8964), .B(n8963), .Z(n9077) );
  NANDN U9510 ( .A(n9126), .B(n8968), .Z(n8972) );
  NANDN U9511 ( .A(n8970), .B(n8969), .Z(n8971) );
  AND U9512 ( .A(n8972), .B(n8971), .Z(n9069) );
  AND U9513 ( .A(x[151]), .B(y[711]), .Z(n9089) );
  AND U9514 ( .A(y[710]), .B(x[152]), .Z(n8974) );
  AND U9515 ( .A(y[709]), .B(x[153]), .Z(n8973) );
  XOR U9516 ( .A(n8974), .B(n8973), .Z(n9088) );
  XOR U9517 ( .A(n9089), .B(n9088), .Z(n9072) );
  ANDN U9518 ( .B(o[93]), .A(n8975), .Z(n9208) );
  AND U9519 ( .A(x[156]), .B(y[706]), .Z(n9210) );
  AND U9520 ( .A(x[144]), .B(y[718]), .Z(n9209) );
  XOR U9521 ( .A(n9210), .B(n9209), .Z(n9207) );
  XNOR U9522 ( .A(n9208), .B(n9207), .Z(n9071) );
  XNOR U9523 ( .A(n9069), .B(n9070), .Z(n9080) );
  XOR U9524 ( .A(n9077), .B(n9078), .Z(n9270) );
  XNOR U9525 ( .A(n9269), .B(n9270), .Z(n9041) );
  XOR U9526 ( .A(n9040), .B(n9039), .Z(n9282) );
  NANDN U9527 ( .A(n8977), .B(n8976), .Z(n8981) );
  NANDN U9528 ( .A(n8979), .B(n8978), .Z(n8980) );
  AND U9529 ( .A(n8981), .B(n8980), .Z(n9284) );
  NANDN U9530 ( .A(n8983), .B(n8982), .Z(n8987) );
  NANDN U9531 ( .A(n8985), .B(n8984), .Z(n8986) );
  NAND U9532 ( .A(n8987), .B(n8986), .Z(n9283) );
  XOR U9533 ( .A(n9284), .B(n9283), .Z(n9281) );
  NANDN U9534 ( .A(n8989), .B(n8988), .Z(n8993) );
  NANDN U9535 ( .A(n8991), .B(n8990), .Z(n8992) );
  AND U9536 ( .A(n8993), .B(n8992), .Z(n9278) );
  NANDN U9537 ( .A(n8995), .B(n8994), .Z(n8999) );
  NAND U9538 ( .A(n8997), .B(n8996), .Z(n8998) );
  AND U9539 ( .A(n8999), .B(n8998), .Z(n9266) );
  NAND U9540 ( .A(n9001), .B(n9000), .Z(n9005) );
  NANDN U9541 ( .A(n9003), .B(n9002), .Z(n9004) );
  AND U9542 ( .A(n9005), .B(n9004), .Z(n9261) );
  NAND U9543 ( .A(n9007), .B(n9006), .Z(n9011) );
  NANDN U9544 ( .A(n9009), .B(n9008), .Z(n9010) );
  NAND U9545 ( .A(n9011), .B(n9010), .Z(n9262) );
  NANDN U9546 ( .A(n9013), .B(n9012), .Z(n9017) );
  NANDN U9547 ( .A(n9015), .B(n9014), .Z(n9016) );
  NAND U9548 ( .A(n9017), .B(n9016), .Z(n9259) );
  XOR U9549 ( .A(n9260), .B(n9259), .Z(n9268) );
  NAND U9550 ( .A(n9121), .B(n9018), .Z(n9022) );
  NAND U9551 ( .A(n9020), .B(n9019), .Z(n9021) );
  AND U9552 ( .A(n9022), .B(n9021), .Z(n9256) );
  NAND U9553 ( .A(n9024), .B(n9023), .Z(n9028) );
  NAND U9554 ( .A(n9026), .B(n9025), .Z(n9027) );
  AND U9555 ( .A(n9028), .B(n9027), .Z(n9064) );
  NAND U9556 ( .A(y[722]), .B(x[140]), .Z(n9029) );
  XNOR U9557 ( .A(n9030), .B(n9029), .Z(n9084) );
  XOR U9558 ( .A(n9084), .B(n9083), .Z(n9120) );
  AND U9559 ( .A(y[725]), .B(x[137]), .Z(n9032) );
  XOR U9560 ( .A(n9032), .B(n9031), .Z(n9119) );
  XOR U9561 ( .A(n9120), .B(n9119), .Z(n9066) );
  AND U9562 ( .A(x[155]), .B(y[707]), .Z(n9204) );
  AND U9563 ( .A(x[129]), .B(y[733]), .Z(n9203) );
  XOR U9564 ( .A(n9204), .B(n9203), .Z(n9202) );
  XOR U9565 ( .A(n9202), .B(n9201), .Z(n9065) );
  XOR U9566 ( .A(n9066), .B(n9065), .Z(n9063) );
  XOR U9567 ( .A(n9064), .B(n9063), .Z(n9255) );
  XOR U9568 ( .A(n9256), .B(n9255), .Z(n9254) );
  NANDN U9569 ( .A(n9034), .B(n9033), .Z(n9038) );
  NAND U9570 ( .A(n9036), .B(n9035), .Z(n9037) );
  AND U9571 ( .A(n9038), .B(n9037), .Z(n9253) );
  XNOR U9572 ( .A(n9254), .B(n9253), .Z(n9267) );
  XOR U9573 ( .A(n9266), .B(n9265), .Z(n9277) );
  XNOR U9574 ( .A(n9278), .B(n9277), .Z(n9276) );
  XOR U9575 ( .A(n9275), .B(n9276), .Z(n9302) );
  XOR U9576 ( .A(n9304), .B(n9303), .Z(n9289) );
  XNOR U9577 ( .A(n9290), .B(n9289), .Z(N191) );
  NANDN U9578 ( .A(n9048), .B(n9047), .Z(n9052) );
  NAND U9579 ( .A(n9050), .B(n9049), .Z(n9051) );
  AND U9580 ( .A(n9052), .B(n9051), .Z(n9274) );
  NANDN U9581 ( .A(n9058), .B(n9057), .Z(n9062) );
  NANDN U9582 ( .A(n9060), .B(n9059), .Z(n9061) );
  NANDN U9583 ( .A(n9064), .B(n9063), .Z(n9068) );
  NAND U9584 ( .A(n9066), .B(n9065), .Z(n9067) );
  AND U9585 ( .A(n9068), .B(n9067), .Z(n9076) );
  NANDN U9586 ( .A(n9070), .B(n9069), .Z(n9074) );
  NANDN U9587 ( .A(n9072), .B(n9071), .Z(n9073) );
  NAND U9588 ( .A(n9074), .B(n9073), .Z(n9075) );
  XNOR U9589 ( .A(n9076), .B(n9075), .Z(n9252) );
  NANDN U9590 ( .A(n9078), .B(n9077), .Z(n9082) );
  NANDN U9591 ( .A(n9080), .B(n9079), .Z(n9081) );
  AND U9592 ( .A(n9082), .B(n9081), .Z(n9250) );
  NAND U9593 ( .A(n9084), .B(n9083), .Z(n9087) );
  NAND U9594 ( .A(n9085), .B(n9164), .Z(n9086) );
  AND U9595 ( .A(n9087), .B(n9086), .Z(n9118) );
  NAND U9596 ( .A(n9089), .B(n9088), .Z(n9092) );
  AND U9597 ( .A(x[153]), .B(y[710]), .Z(n9144) );
  NANDN U9598 ( .A(n9090), .B(n9144), .Z(n9091) );
  AND U9599 ( .A(n9092), .B(n9091), .Z(n9100) );
  NAND U9600 ( .A(n9094), .B(n9093), .Z(n9098) );
  NAND U9601 ( .A(n9096), .B(n9095), .Z(n9097) );
  NAND U9602 ( .A(n9098), .B(n9097), .Z(n9099) );
  XNOR U9603 ( .A(n9100), .B(n9099), .Z(n9116) );
  AND U9604 ( .A(y[729]), .B(x[134]), .Z(n9102) );
  NAND U9605 ( .A(y[728]), .B(x[135]), .Z(n9101) );
  XNOR U9606 ( .A(n9102), .B(n9101), .Z(n9106) );
  AND U9607 ( .A(y[723]), .B(x[140]), .Z(n9104) );
  NAND U9608 ( .A(y[719]), .B(x[144]), .Z(n9103) );
  XNOR U9609 ( .A(n9104), .B(n9103), .Z(n9105) );
  XOR U9610 ( .A(n9106), .B(n9105), .Z(n9114) );
  AND U9611 ( .A(y[730]), .B(x[133]), .Z(n9108) );
  NAND U9612 ( .A(y[717]), .B(x[146]), .Z(n9107) );
  XNOR U9613 ( .A(n9108), .B(n9107), .Z(n9112) );
  AND U9614 ( .A(y[732]), .B(x[131]), .Z(n9110) );
  NAND U9615 ( .A(y[731]), .B(x[132]), .Z(n9109) );
  XNOR U9616 ( .A(n9110), .B(n9109), .Z(n9111) );
  XNOR U9617 ( .A(n9112), .B(n9111), .Z(n9113) );
  XNOR U9618 ( .A(n9114), .B(n9113), .Z(n9115) );
  XNOR U9619 ( .A(n9116), .B(n9115), .Z(n9117) );
  XNOR U9620 ( .A(n9118), .B(n9117), .Z(n9200) );
  NAND U9621 ( .A(n9120), .B(n9119), .Z(n9123) );
  AND U9622 ( .A(x[138]), .B(y[725]), .Z(n9163) );
  NAND U9623 ( .A(n9121), .B(n9163), .Z(n9122) );
  AND U9624 ( .A(n9123), .B(n9122), .Z(n9198) );
  NAND U9625 ( .A(n9125), .B(n9124), .Z(n9128) );
  AND U9626 ( .A(x[150]), .B(y[713]), .Z(n9145) );
  NANDN U9627 ( .A(n9126), .B(n9145), .Z(n9127) );
  AND U9628 ( .A(n9128), .B(n9127), .Z(n9136) );
  NAND U9629 ( .A(n9130), .B(n9129), .Z(n9134) );
  NAND U9630 ( .A(n9132), .B(n9131), .Z(n9133) );
  NAND U9631 ( .A(n9134), .B(n9133), .Z(n9135) );
  XNOR U9632 ( .A(n9136), .B(n9135), .Z(n9196) );
  NAND U9633 ( .A(n9138), .B(n9137), .Z(n9142) );
  NAND U9634 ( .A(n9140), .B(n9139), .Z(n9141) );
  AND U9635 ( .A(n9142), .B(n9141), .Z(n9194) );
  AND U9636 ( .A(y[708]), .B(x[155]), .Z(n9152) );
  AND U9637 ( .A(n9143), .B(o[94]), .Z(n9150) );
  XOR U9638 ( .A(n9144), .B(o[95]), .Z(n9148) );
  XNOR U9639 ( .A(n9146), .B(n9145), .Z(n9147) );
  XNOR U9640 ( .A(n9148), .B(n9147), .Z(n9149) );
  XNOR U9641 ( .A(n9150), .B(n9149), .Z(n9151) );
  XNOR U9642 ( .A(n9152), .B(n9151), .Z(n9192) );
  AND U9643 ( .A(y[716]), .B(x[147]), .Z(n9154) );
  NAND U9644 ( .A(y[727]), .B(x[136]), .Z(n9153) );
  XNOR U9645 ( .A(n9154), .B(n9153), .Z(n9162) );
  AND U9646 ( .A(y[714]), .B(x[149]), .Z(n9160) );
  AND U9647 ( .A(y[705]), .B(x[158]), .Z(n9156) );
  NAND U9648 ( .A(y[706]), .B(x[157]), .Z(n9155) );
  XNOR U9649 ( .A(n9156), .B(n9155), .Z(n9157) );
  XNOR U9650 ( .A(n9158), .B(n9157), .Z(n9159) );
  XNOR U9651 ( .A(n9160), .B(n9159), .Z(n9161) );
  XOR U9652 ( .A(n9162), .B(n9161), .Z(n9166) );
  XNOR U9653 ( .A(n9164), .B(n9163), .Z(n9165) );
  XNOR U9654 ( .A(n9166), .B(n9165), .Z(n9182) );
  AND U9655 ( .A(y[715]), .B(x[148]), .Z(n9168) );
  NAND U9656 ( .A(y[709]), .B(x[154]), .Z(n9167) );
  XNOR U9657 ( .A(n9168), .B(n9167), .Z(n9172) );
  AND U9658 ( .A(y[726]), .B(x[137]), .Z(n9170) );
  NAND U9659 ( .A(y[724]), .B(x[139]), .Z(n9169) );
  XNOR U9660 ( .A(n9170), .B(n9169), .Z(n9171) );
  XOR U9661 ( .A(n9172), .B(n9171), .Z(n9180) );
  AND U9662 ( .A(y[707]), .B(x[156]), .Z(n9174) );
  NAND U9663 ( .A(y[735]), .B(x[128]), .Z(n9173) );
  XNOR U9664 ( .A(n9174), .B(n9173), .Z(n9178) );
  AND U9665 ( .A(y[734]), .B(x[129]), .Z(n9176) );
  NAND U9666 ( .A(y[721]), .B(x[142]), .Z(n9175) );
  XNOR U9667 ( .A(n9176), .B(n9175), .Z(n9177) );
  XNOR U9668 ( .A(n9178), .B(n9177), .Z(n9179) );
  XNOR U9669 ( .A(n9180), .B(n9179), .Z(n9181) );
  XOR U9670 ( .A(n9182), .B(n9181), .Z(n9190) );
  AND U9671 ( .A(y[718]), .B(x[145]), .Z(n9184) );
  NAND U9672 ( .A(y[712]), .B(x[151]), .Z(n9183) );
  XNOR U9673 ( .A(n9184), .B(n9183), .Z(n9188) );
  AND U9674 ( .A(y[704]), .B(x[159]), .Z(n9186) );
  NAND U9675 ( .A(y[733]), .B(x[130]), .Z(n9185) );
  XNOR U9676 ( .A(n9186), .B(n9185), .Z(n9187) );
  XNOR U9677 ( .A(n9188), .B(n9187), .Z(n9189) );
  XNOR U9678 ( .A(n9190), .B(n9189), .Z(n9191) );
  XNOR U9679 ( .A(n9192), .B(n9191), .Z(n9193) );
  XNOR U9680 ( .A(n9194), .B(n9193), .Z(n9195) );
  XNOR U9681 ( .A(n9196), .B(n9195), .Z(n9197) );
  XNOR U9682 ( .A(n9198), .B(n9197), .Z(n9199) );
  XOR U9683 ( .A(n9200), .B(n9199), .Z(n9232) );
  NAND U9684 ( .A(n9202), .B(n9201), .Z(n9206) );
  NAND U9685 ( .A(n9204), .B(n9203), .Z(n9205) );
  AND U9686 ( .A(n9206), .B(n9205), .Z(n9214) );
  NAND U9687 ( .A(n9208), .B(n9207), .Z(n9212) );
  NAND U9688 ( .A(n9210), .B(n9209), .Z(n9211) );
  NAND U9689 ( .A(n9212), .B(n9211), .Z(n9213) );
  XNOR U9690 ( .A(n9214), .B(n9213), .Z(n9230) );
  NAND U9691 ( .A(n9216), .B(n9215), .Z(n9220) );
  NAND U9692 ( .A(n9218), .B(n9217), .Z(n9219) );
  AND U9693 ( .A(n9220), .B(n9219), .Z(n9228) );
  NAND U9694 ( .A(n9222), .B(n9221), .Z(n9226) );
  NAND U9695 ( .A(n9224), .B(n9223), .Z(n9225) );
  NAND U9696 ( .A(n9226), .B(n9225), .Z(n9227) );
  XNOR U9697 ( .A(n9228), .B(n9227), .Z(n9229) );
  XNOR U9698 ( .A(n9230), .B(n9229), .Z(n9231) );
  XNOR U9699 ( .A(n9232), .B(n9231), .Z(n9248) );
  NANDN U9700 ( .A(n9234), .B(n9233), .Z(n9238) );
  NANDN U9701 ( .A(n9236), .B(n9235), .Z(n9237) );
  AND U9702 ( .A(n9238), .B(n9237), .Z(n9246) );
  NAND U9703 ( .A(n9240), .B(n9239), .Z(n9244) );
  NANDN U9704 ( .A(n9242), .B(n9241), .Z(n9243) );
  NAND U9705 ( .A(n9244), .B(n9243), .Z(n9245) );
  XNOR U9706 ( .A(n9246), .B(n9245), .Z(n9247) );
  XNOR U9707 ( .A(n9248), .B(n9247), .Z(n9249) );
  XNOR U9708 ( .A(n9250), .B(n9249), .Z(n9251) );
  NAND U9709 ( .A(n9254), .B(n9253), .Z(n9258) );
  NAND U9710 ( .A(n9256), .B(n9255), .Z(n9257) );
  NAND U9711 ( .A(n9260), .B(n9259), .Z(n9264) );
  NANDN U9712 ( .A(n9262), .B(n9261), .Z(n9263) );
  NAND U9713 ( .A(n9276), .B(n9275), .Z(n9280) );
  NANDN U9714 ( .A(n9278), .B(n9277), .Z(n9279) );
  AND U9715 ( .A(n9280), .B(n9279), .Z(n9288) );
  NANDN U9716 ( .A(n9282), .B(n9281), .Z(n9286) );
  NAND U9717 ( .A(n9284), .B(n9283), .Z(n9285) );
  NAND U9718 ( .A(n9286), .B(n9285), .Z(n9287) );
  NAND U9719 ( .A(n9290), .B(n9289), .Z(n9294) );
  NANDN U9720 ( .A(n9292), .B(n9291), .Z(n9293) );
  NAND U9721 ( .A(n9296), .B(n9295), .Z(n9300) );
  NANDN U9722 ( .A(n9298), .B(n9297), .Z(n9299) );
  AND U9723 ( .A(x[128]), .B(y[736]), .Z(n9959) );
  XOR U9724 ( .A(n9959), .B(o[96]), .Z(N225) );
  AND U9725 ( .A(x[129]), .B(y[736]), .Z(n9313) );
  AND U9726 ( .A(x[128]), .B(y[737]), .Z(n9312) );
  XNOR U9727 ( .A(n9312), .B(o[97]), .Z(n9305) );
  XNOR U9728 ( .A(n9313), .B(n9305), .Z(n9307) );
  NAND U9729 ( .A(n9959), .B(o[96]), .Z(n9306) );
  XNOR U9730 ( .A(n9307), .B(n9306), .Z(N226) );
  NANDN U9731 ( .A(n9313), .B(n9305), .Z(n9309) );
  NAND U9732 ( .A(n9307), .B(n9306), .Z(n9308) );
  AND U9733 ( .A(n9309), .B(n9308), .Z(n9319) );
  AND U9734 ( .A(x[128]), .B(y[738]), .Z(n9326) );
  XNOR U9735 ( .A(n9326), .B(o[98]), .Z(n9318) );
  XNOR U9736 ( .A(n9319), .B(n9318), .Z(n9321) );
  AND U9737 ( .A(y[737]), .B(x[129]), .Z(n9311) );
  NAND U9738 ( .A(y[736]), .B(x[130]), .Z(n9310) );
  XNOR U9739 ( .A(n9311), .B(n9310), .Z(n9315) );
  AND U9740 ( .A(n9312), .B(o[97]), .Z(n9314) );
  XNOR U9741 ( .A(n9315), .B(n9314), .Z(n9320) );
  XNOR U9742 ( .A(n9321), .B(n9320), .Z(N227) );
  AND U9743 ( .A(x[130]), .B(y[737]), .Z(n9333) );
  NAND U9744 ( .A(n9333), .B(n9313), .Z(n9317) );
  NAND U9745 ( .A(n9315), .B(n9314), .Z(n9316) );
  AND U9746 ( .A(n9317), .B(n9316), .Z(n9336) );
  NANDN U9747 ( .A(n9319), .B(n9318), .Z(n9323) );
  NAND U9748 ( .A(n9321), .B(n9320), .Z(n9322) );
  AND U9749 ( .A(n9323), .B(n9322), .Z(n9335) );
  XNOR U9750 ( .A(n9336), .B(n9335), .Z(n9338) );
  AND U9751 ( .A(x[129]), .B(y[738]), .Z(n9455) );
  XOR U9752 ( .A(n9333), .B(o[99]), .Z(n9341) );
  XOR U9753 ( .A(n9455), .B(n9341), .Z(n9343) );
  AND U9754 ( .A(y[739]), .B(x[128]), .Z(n9325) );
  NAND U9755 ( .A(y[736]), .B(x[131]), .Z(n9324) );
  XNOR U9756 ( .A(n9325), .B(n9324), .Z(n9328) );
  AND U9757 ( .A(n9326), .B(o[98]), .Z(n9327) );
  XOR U9758 ( .A(n9328), .B(n9327), .Z(n9342) );
  XOR U9759 ( .A(n9343), .B(n9342), .Z(n9337) );
  XOR U9760 ( .A(n9338), .B(n9337), .Z(N228) );
  AND U9761 ( .A(x[131]), .B(y[739]), .Z(n9386) );
  NAND U9762 ( .A(n9959), .B(n9386), .Z(n9330) );
  NAND U9763 ( .A(n9328), .B(n9327), .Z(n9329) );
  AND U9764 ( .A(n9330), .B(n9329), .Z(n9364) );
  AND U9765 ( .A(y[740]), .B(x[128]), .Z(n9332) );
  NAND U9766 ( .A(y[736]), .B(x[132]), .Z(n9331) );
  XNOR U9767 ( .A(n9332), .B(n9331), .Z(n9357) );
  NAND U9768 ( .A(n9333), .B(o[99]), .Z(n9358) );
  AND U9769 ( .A(y[739]), .B(x[129]), .Z(n9547) );
  NAND U9770 ( .A(y[738]), .B(x[130]), .Z(n9334) );
  XNOR U9771 ( .A(n9547), .B(n9334), .Z(n9354) );
  NAND U9772 ( .A(x[131]), .B(y[737]), .Z(n9349) );
  XNOR U9773 ( .A(o[100]), .B(n9349), .Z(n9353) );
  XOR U9774 ( .A(n9354), .B(n9353), .Z(n9361) );
  XOR U9775 ( .A(n9362), .B(n9361), .Z(n9363) );
  XNOR U9776 ( .A(n9364), .B(n9363), .Z(n9368) );
  NANDN U9777 ( .A(n9336), .B(n9335), .Z(n9340) );
  NAND U9778 ( .A(n9338), .B(n9337), .Z(n9339) );
  NAND U9779 ( .A(n9340), .B(n9339), .Z(n9369) );
  NAND U9780 ( .A(n9455), .B(n9341), .Z(n9345) );
  NAND U9781 ( .A(n9343), .B(n9342), .Z(n9344) );
  NAND U9782 ( .A(n9345), .B(n9344), .Z(n9370) );
  IV U9783 ( .A(n9370), .Z(n9367) );
  XOR U9784 ( .A(n9369), .B(n9367), .Z(n9346) );
  XNOR U9785 ( .A(n9368), .B(n9346), .Z(N229) );
  AND U9786 ( .A(y[740]), .B(x[129]), .Z(n9348) );
  NAND U9787 ( .A(y[738]), .B(x[131]), .Z(n9347) );
  XNOR U9788 ( .A(n9348), .B(n9347), .Z(n9373) );
  AND U9789 ( .A(x[132]), .B(y[737]), .Z(n9382) );
  XOR U9790 ( .A(n9382), .B(o[101]), .Z(n9372) );
  XNOR U9791 ( .A(n9373), .B(n9372), .Z(n9376) );
  NAND U9792 ( .A(x[130]), .B(y[739]), .Z(n9463) );
  ANDN U9793 ( .B(o[100]), .A(n9349), .Z(n9378) );
  AND U9794 ( .A(y[741]), .B(x[128]), .Z(n9351) );
  NAND U9795 ( .A(y[736]), .B(x[133]), .Z(n9350) );
  XOR U9796 ( .A(n9351), .B(n9350), .Z(n9379) );
  XNOR U9797 ( .A(n9378), .B(n9379), .Z(n9377) );
  XOR U9798 ( .A(n9463), .B(n9377), .Z(n9352) );
  XOR U9799 ( .A(n9376), .B(n9352), .Z(n9394) );
  NANDN U9800 ( .A(n9463), .B(n9455), .Z(n9356) );
  NAND U9801 ( .A(n9354), .B(n9353), .Z(n9355) );
  AND U9802 ( .A(n9356), .B(n9355), .Z(n9392) );
  AND U9803 ( .A(x[132]), .B(y[740]), .Z(n10157) );
  NAND U9804 ( .A(n10157), .B(n9959), .Z(n9360) );
  NANDN U9805 ( .A(n9358), .B(n9357), .Z(n9359) );
  NAND U9806 ( .A(n9360), .B(n9359), .Z(n9391) );
  XNOR U9807 ( .A(n9394), .B(n9393), .Z(n9390) );
  NAND U9808 ( .A(n9362), .B(n9361), .Z(n9366) );
  NANDN U9809 ( .A(n9364), .B(n9363), .Z(n9365) );
  NAND U9810 ( .A(n9366), .B(n9365), .Z(n9389) );
  XOR U9811 ( .A(n9389), .B(n9388), .Z(n9371) );
  XNOR U9812 ( .A(n9390), .B(n9371), .Z(N230) );
  AND U9813 ( .A(x[131]), .B(y[740]), .Z(n9465) );
  NAND U9814 ( .A(n9455), .B(n9465), .Z(n9375) );
  NAND U9815 ( .A(n9373), .B(n9372), .Z(n9374) );
  AND U9816 ( .A(n9375), .B(n9374), .Z(n9430) );
  XNOR U9817 ( .A(n9430), .B(n9429), .Z(n9432) );
  AND U9818 ( .A(x[133]), .B(y[741]), .Z(n9627) );
  NAND U9819 ( .A(n9959), .B(n9627), .Z(n9381) );
  NANDN U9820 ( .A(n9379), .B(n9378), .Z(n9380) );
  AND U9821 ( .A(n9381), .B(n9380), .Z(n9399) );
  AND U9822 ( .A(n9382), .B(o[101]), .Z(n9405) );
  AND U9823 ( .A(y[742]), .B(x[128]), .Z(n9384) );
  NAND U9824 ( .A(y[736]), .B(x[134]), .Z(n9383) );
  XOR U9825 ( .A(n9384), .B(n9383), .Z(n9406) );
  XNOR U9826 ( .A(n9405), .B(n9406), .Z(n9398) );
  XNOR U9827 ( .A(n9399), .B(n9398), .Z(n9401) );
  NAND U9828 ( .A(y[740]), .B(x[130]), .Z(n9385) );
  XNOR U9829 ( .A(n9386), .B(n9385), .Z(n9410) );
  AND U9830 ( .A(y[741]), .B(x[129]), .Z(n9661) );
  NAND U9831 ( .A(y[738]), .B(x[132]), .Z(n9387) );
  XNOR U9832 ( .A(n9661), .B(n9387), .Z(n9414) );
  NAND U9833 ( .A(x[133]), .B(y[737]), .Z(n9419) );
  XNOR U9834 ( .A(o[102]), .B(n9419), .Z(n9413) );
  XOR U9835 ( .A(n9414), .B(n9413), .Z(n9409) );
  XOR U9836 ( .A(n9410), .B(n9409), .Z(n9400) );
  XOR U9837 ( .A(n9401), .B(n9400), .Z(n9431) );
  XNOR U9838 ( .A(n9432), .B(n9431), .Z(n9425) );
  NANDN U9839 ( .A(n9392), .B(n9391), .Z(n9396) );
  NAND U9840 ( .A(n9394), .B(n9393), .Z(n9395) );
  NAND U9841 ( .A(n9396), .B(n9395), .Z(n9423) );
  IV U9842 ( .A(n9423), .Z(n9422) );
  XOR U9843 ( .A(n9424), .B(n9422), .Z(n9397) );
  XNOR U9844 ( .A(n9425), .B(n9397), .Z(N231) );
  NANDN U9845 ( .A(n9399), .B(n9398), .Z(n9403) );
  NAND U9846 ( .A(n9401), .B(n9400), .Z(n9402) );
  AND U9847 ( .A(n9403), .B(n9402), .Z(n9439) );
  AND U9848 ( .A(y[738]), .B(x[133]), .Z(n9535) );
  NAND U9849 ( .A(y[742]), .B(x[129]), .Z(n9404) );
  XNOR U9850 ( .A(n9535), .B(n9404), .Z(n9457) );
  NAND U9851 ( .A(x[134]), .B(y[737]), .Z(n9460) );
  XNOR U9852 ( .A(o[103]), .B(n9460), .Z(n9456) );
  XOR U9853 ( .A(n9457), .B(n9456), .Z(n9476) );
  AND U9854 ( .A(x[134]), .B(y[742]), .Z(n9503) );
  NAND U9855 ( .A(n9959), .B(n9503), .Z(n9408) );
  NANDN U9856 ( .A(n9406), .B(n9405), .Z(n9407) );
  AND U9857 ( .A(n9408), .B(n9407), .Z(n9475) );
  NANDN U9858 ( .A(n9463), .B(n9465), .Z(n9412) );
  NAND U9859 ( .A(n9410), .B(n9409), .Z(n9411) );
  AND U9860 ( .A(n9412), .B(n9411), .Z(n9477) );
  XOR U9861 ( .A(n9478), .B(n9477), .Z(n9437) );
  AND U9862 ( .A(x[132]), .B(y[741]), .Z(n9964) );
  NAND U9863 ( .A(n9964), .B(n9455), .Z(n9416) );
  NAND U9864 ( .A(n9414), .B(n9413), .Z(n9415) );
  AND U9865 ( .A(n9416), .B(n9415), .Z(n9452) );
  AND U9866 ( .A(y[741]), .B(x[130]), .Z(n9418) );
  NAND U9867 ( .A(y[739]), .B(x[132]), .Z(n9417) );
  XNOR U9868 ( .A(n9418), .B(n9417), .Z(n9464) );
  XOR U9869 ( .A(n9465), .B(n9464), .Z(n9450) );
  ANDN U9870 ( .B(o[102]), .A(n9419), .Z(n9470) );
  AND U9871 ( .A(y[743]), .B(x[128]), .Z(n9421) );
  NAND U9872 ( .A(y[736]), .B(x[135]), .Z(n9420) );
  XNOR U9873 ( .A(n9421), .B(n9420), .Z(n9469) );
  XNOR U9874 ( .A(n9470), .B(n9469), .Z(n9449) );
  XNOR U9875 ( .A(n9450), .B(n9449), .Z(n9451) );
  XOR U9876 ( .A(n9452), .B(n9451), .Z(n9436) );
  XOR U9877 ( .A(n9437), .B(n9436), .Z(n9438) );
  XNOR U9878 ( .A(n9439), .B(n9438), .Z(n9445) );
  OR U9879 ( .A(n9424), .B(n9422), .Z(n9428) );
  ANDN U9880 ( .B(n9424), .A(n9423), .Z(n9426) );
  OR U9881 ( .A(n9426), .B(n9425), .Z(n9427) );
  AND U9882 ( .A(n9428), .B(n9427), .Z(n9443) );
  NANDN U9883 ( .A(n9430), .B(n9429), .Z(n9434) );
  NAND U9884 ( .A(n9432), .B(n9431), .Z(n9433) );
  AND U9885 ( .A(n9434), .B(n9433), .Z(n9444) );
  IV U9886 ( .A(n9444), .Z(n9442) );
  XOR U9887 ( .A(n9443), .B(n9442), .Z(n9435) );
  XNOR U9888 ( .A(n9445), .B(n9435), .Z(N232) );
  NAND U9889 ( .A(n9437), .B(n9436), .Z(n9441) );
  NAND U9890 ( .A(n9439), .B(n9438), .Z(n9440) );
  AND U9891 ( .A(n9441), .B(n9440), .Z(n9520) );
  NANDN U9892 ( .A(n9442), .B(n9443), .Z(n9448) );
  NOR U9893 ( .A(n9444), .B(n9443), .Z(n9446) );
  OR U9894 ( .A(n9446), .B(n9445), .Z(n9447) );
  AND U9895 ( .A(n9448), .B(n9447), .Z(n9519) );
  NANDN U9896 ( .A(n9450), .B(n9449), .Z(n9454) );
  NAND U9897 ( .A(n9452), .B(n9451), .Z(n9453) );
  AND U9898 ( .A(n9454), .B(n9453), .Z(n9516) );
  AND U9899 ( .A(x[133]), .B(y[742]), .Z(n9619) );
  NAND U9900 ( .A(n9619), .B(n9455), .Z(n9459) );
  NAND U9901 ( .A(n9457), .B(n9456), .Z(n9458) );
  AND U9902 ( .A(n9459), .B(n9458), .Z(n9514) );
  ANDN U9903 ( .B(o[103]), .A(n9460), .Z(n9494) );
  AND U9904 ( .A(y[739]), .B(x[133]), .Z(n10064) );
  NAND U9905 ( .A(y[743]), .B(x[129]), .Z(n9461) );
  XNOR U9906 ( .A(n10064), .B(n9461), .Z(n9493) );
  XOR U9907 ( .A(n9494), .B(n9493), .Z(n9499) );
  NAND U9908 ( .A(x[131]), .B(y[741]), .Z(n10278) );
  AND U9909 ( .A(y[742]), .B(x[130]), .Z(n10354) );
  NAND U9910 ( .A(y[738]), .B(x[134]), .Z(n9462) );
  XNOR U9911 ( .A(n10354), .B(n9462), .Z(n9504) );
  XNOR U9912 ( .A(n10157), .B(n9504), .Z(n9497) );
  XOR U9913 ( .A(n10278), .B(n9497), .Z(n9498) );
  XOR U9914 ( .A(n9499), .B(n9498), .Z(n9513) );
  XNOR U9915 ( .A(n9514), .B(n9513), .Z(n9515) );
  XOR U9916 ( .A(n9516), .B(n9515), .Z(n9525) );
  NANDN U9917 ( .A(n9463), .B(n9964), .Z(n9467) );
  NAND U9918 ( .A(n9465), .B(n9464), .Z(n9466) );
  AND U9919 ( .A(n9467), .B(n9466), .Z(n9510) );
  AND U9920 ( .A(x[135]), .B(y[743]), .Z(n9468) );
  NAND U9921 ( .A(n9959), .B(n9468), .Z(n9472) );
  NAND U9922 ( .A(n9470), .B(n9469), .Z(n9471) );
  AND U9923 ( .A(n9472), .B(n9471), .Z(n9508) );
  AND U9924 ( .A(y[744]), .B(x[128]), .Z(n9474) );
  NAND U9925 ( .A(y[736]), .B(x[136]), .Z(n9473) );
  XNOR U9926 ( .A(n9474), .B(n9473), .Z(n9484) );
  NAND U9927 ( .A(x[135]), .B(y[737]), .Z(n9489) );
  XNOR U9928 ( .A(o[104]), .B(n9489), .Z(n9483) );
  XOR U9929 ( .A(n9484), .B(n9483), .Z(n9507) );
  XNOR U9930 ( .A(n9508), .B(n9507), .Z(n9509) );
  XNOR U9931 ( .A(n9510), .B(n9509), .Z(n9523) );
  NANDN U9932 ( .A(n9476), .B(n9475), .Z(n9480) );
  NAND U9933 ( .A(n9478), .B(n9477), .Z(n9479) );
  NAND U9934 ( .A(n9480), .B(n9479), .Z(n9522) );
  XNOR U9935 ( .A(n9519), .B(n9521), .Z(n9481) );
  XOR U9936 ( .A(n9520), .B(n9481), .Z(N233) );
  AND U9937 ( .A(x[136]), .B(y[744]), .Z(n9482) );
  NAND U9938 ( .A(n9482), .B(n9959), .Z(n9486) );
  NAND U9939 ( .A(n9484), .B(n9483), .Z(n9485) );
  AND U9940 ( .A(n9486), .B(n9485), .Z(n9564) );
  AND U9941 ( .A(y[740]), .B(x[133]), .Z(n9488) );
  NAND U9942 ( .A(y[738]), .B(x[135]), .Z(n9487) );
  XNOR U9943 ( .A(n9488), .B(n9487), .Z(n9538) );
  ANDN U9944 ( .B(o[104]), .A(n9489), .Z(n9537) );
  XOR U9945 ( .A(n9538), .B(n9537), .Z(n9562) );
  AND U9946 ( .A(y[736]), .B(x[137]), .Z(n9491) );
  NAND U9947 ( .A(y[745]), .B(x[128]), .Z(n9490) );
  XNOR U9948 ( .A(n9491), .B(n9490), .Z(n9544) );
  NAND U9949 ( .A(x[136]), .B(y[737]), .Z(n9553) );
  XNOR U9950 ( .A(n9544), .B(n9543), .Z(n9561) );
  XNOR U9951 ( .A(n9562), .B(n9561), .Z(n9563) );
  XOR U9952 ( .A(n9564), .B(n9563), .Z(n9558) );
  AND U9953 ( .A(y[744]), .B(x[129]), .Z(n10267) );
  NAND U9954 ( .A(y[739]), .B(x[134]), .Z(n9492) );
  XNOR U9955 ( .A(n10267), .B(n9492), .Z(n9548) );
  XOR U9956 ( .A(n9964), .B(n9548), .Z(n9568) );
  NAND U9957 ( .A(x[130]), .B(y[743]), .Z(n10112) );
  IV U9958 ( .A(n10112), .Z(n10201) );
  NAND U9959 ( .A(x[131]), .B(y[742]), .Z(n9880) );
  XNOR U9960 ( .A(n10201), .B(n9880), .Z(n9567) );
  XOR U9961 ( .A(n9568), .B(n9567), .Z(n9556) );
  NAND U9962 ( .A(x[133]), .B(y[743]), .Z(n9743) );
  NANDN U9963 ( .A(n9743), .B(n9547), .Z(n9496) );
  NAND U9964 ( .A(n9494), .B(n9493), .Z(n9495) );
  NAND U9965 ( .A(n9496), .B(n9495), .Z(n9555) );
  XOR U9966 ( .A(n9556), .B(n9555), .Z(n9557) );
  XOR U9967 ( .A(n9558), .B(n9557), .Z(n9531) );
  NAND U9968 ( .A(n10278), .B(n9497), .Z(n9501) );
  NANDN U9969 ( .A(n9499), .B(n9498), .Z(n9500) );
  AND U9970 ( .A(n9501), .B(n9500), .Z(n9530) );
  AND U9971 ( .A(x[130]), .B(y[738]), .Z(n9502) );
  NAND U9972 ( .A(n9503), .B(n9502), .Z(n9506) );
  NAND U9973 ( .A(n10157), .B(n9504), .Z(n9505) );
  AND U9974 ( .A(n9506), .B(n9505), .Z(n9529) );
  XNOR U9975 ( .A(n9530), .B(n9529), .Z(n9532) );
  XNOR U9976 ( .A(n9531), .B(n9532), .Z(n9580) );
  NANDN U9977 ( .A(n9508), .B(n9507), .Z(n9512) );
  NANDN U9978 ( .A(n9510), .B(n9509), .Z(n9511) );
  AND U9979 ( .A(n9512), .B(n9511), .Z(n9579) );
  NANDN U9980 ( .A(n9514), .B(n9513), .Z(n9518) );
  NAND U9981 ( .A(n9516), .B(n9515), .Z(n9517) );
  NAND U9982 ( .A(n9518), .B(n9517), .Z(n9578) );
  XNOR U9983 ( .A(n9579), .B(n9578), .Z(n9581) );
  XNOR U9984 ( .A(n9580), .B(n9581), .Z(n9574) );
  NANDN U9985 ( .A(n9523), .B(n9522), .Z(n9527) );
  NANDN U9986 ( .A(n9525), .B(n9524), .Z(n9526) );
  AND U9987 ( .A(n9527), .B(n9526), .Z(n9572) );
  IV U9988 ( .A(n9572), .Z(n9571) );
  XOR U9989 ( .A(n9573), .B(n9571), .Z(n9528) );
  XNOR U9990 ( .A(n9574), .B(n9528), .Z(N234) );
  NANDN U9991 ( .A(n9530), .B(n9529), .Z(n9534) );
  NAND U9992 ( .A(n9532), .B(n9531), .Z(n9533) );
  AND U9993 ( .A(n9534), .B(n9533), .Z(n9647) );
  AND U9994 ( .A(x[135]), .B(y[740]), .Z(n9536) );
  NAND U9995 ( .A(n9536), .B(n9535), .Z(n9540) );
  NAND U9996 ( .A(n9538), .B(n9537), .Z(n9539) );
  AND U9997 ( .A(n9540), .B(n9539), .Z(n9634) );
  AND U9998 ( .A(y[742]), .B(x[132]), .Z(n9542) );
  NAND U9999 ( .A(y[739]), .B(x[135]), .Z(n9541) );
  XNOR U10000 ( .A(n9542), .B(n9541), .Z(n9606) );
  AND U10001 ( .A(x[134]), .B(y[740]), .Z(n9605) );
  XOR U10002 ( .A(n9606), .B(n9605), .Z(n9632) );
  AND U10003 ( .A(x[136]), .B(y[738]), .Z(n9817) );
  NAND U10004 ( .A(x[137]), .B(y[737]), .Z(n9615) );
  XNOR U10005 ( .A(o[106]), .B(n9615), .Z(n9626) );
  XOR U10006 ( .A(n9817), .B(n9626), .Z(n9628) );
  XNOR U10007 ( .A(n9628), .B(n9627), .Z(n9631) );
  XOR U10008 ( .A(n9634), .B(n9633), .Z(n9594) );
  AND U10009 ( .A(x[137]), .B(y[745]), .Z(n10166) );
  NAND U10010 ( .A(n10166), .B(n9959), .Z(n9546) );
  NAND U10011 ( .A(n9544), .B(n9543), .Z(n9545) );
  AND U10012 ( .A(n9546), .B(n9545), .Z(n9592) );
  AND U10013 ( .A(x[134]), .B(y[744]), .Z(n9852) );
  NAND U10014 ( .A(n9852), .B(n9547), .Z(n9550) );
  NAND U10015 ( .A(n9964), .B(n9548), .Z(n9549) );
  AND U10016 ( .A(n9550), .B(n9549), .Z(n9600) );
  AND U10017 ( .A(y[746]), .B(x[128]), .Z(n9552) );
  NAND U10018 ( .A(y[736]), .B(x[138]), .Z(n9551) );
  XNOR U10019 ( .A(n9552), .B(n9551), .Z(n9610) );
  ANDN U10020 ( .B(o[105]), .A(n9553), .Z(n9609) );
  XOR U10021 ( .A(n9610), .B(n9609), .Z(n9598) );
  AND U10022 ( .A(y[745]), .B(x[129]), .Z(n10460) );
  NAND U10023 ( .A(y[743]), .B(x[131]), .Z(n9554) );
  XNOR U10024 ( .A(n10460), .B(n9554), .Z(n9622) );
  NAND U10025 ( .A(x[130]), .B(y[744]), .Z(n9623) );
  XOR U10026 ( .A(n9598), .B(n9597), .Z(n9599) );
  XNOR U10027 ( .A(n9592), .B(n9591), .Z(n9593) );
  XOR U10028 ( .A(n9594), .B(n9593), .Z(n9645) );
  NAND U10029 ( .A(n9556), .B(n9555), .Z(n9560) );
  NANDN U10030 ( .A(n9558), .B(n9557), .Z(n9559) );
  AND U10031 ( .A(n9560), .B(n9559), .Z(n9588) );
  NANDN U10032 ( .A(n9562), .B(n9561), .Z(n9566) );
  NAND U10033 ( .A(n9564), .B(n9563), .Z(n9565) );
  AND U10034 ( .A(n9566), .B(n9565), .Z(n9585) );
  ANDN U10035 ( .B(n9880), .A(n10201), .Z(n9570) );
  NANDN U10036 ( .A(n9568), .B(n9567), .Z(n9569) );
  NANDN U10037 ( .A(n9570), .B(n9569), .Z(n9586) );
  XNOR U10038 ( .A(n9585), .B(n9586), .Z(n9587) );
  XOR U10039 ( .A(n9588), .B(n9587), .Z(n9644) );
  XOR U10040 ( .A(n9645), .B(n9644), .Z(n9646) );
  XOR U10041 ( .A(n9647), .B(n9646), .Z(n9640) );
  OR U10042 ( .A(n9573), .B(n9571), .Z(n9577) );
  ANDN U10043 ( .B(n9573), .A(n9572), .Z(n9575) );
  OR U10044 ( .A(n9575), .B(n9574), .Z(n9576) );
  AND U10045 ( .A(n9577), .B(n9576), .Z(n9638) );
  NANDN U10046 ( .A(n9579), .B(n9578), .Z(n9583) );
  NAND U10047 ( .A(n9581), .B(n9580), .Z(n9582) );
  AND U10048 ( .A(n9583), .B(n9582), .Z(n9639) );
  IV U10049 ( .A(n9639), .Z(n9637) );
  XOR U10050 ( .A(n9638), .B(n9637), .Z(n9584) );
  XNOR U10051 ( .A(n9640), .B(n9584), .Z(N235) );
  NANDN U10052 ( .A(n9586), .B(n9585), .Z(n9590) );
  NANDN U10053 ( .A(n9588), .B(n9587), .Z(n9589) );
  AND U10054 ( .A(n9590), .B(n9589), .Z(n9711) );
  NANDN U10055 ( .A(n9592), .B(n9591), .Z(n9596) );
  NANDN U10056 ( .A(n9594), .B(n9593), .Z(n9595) );
  AND U10057 ( .A(n9596), .B(n9595), .Z(n9709) );
  NAND U10058 ( .A(n9598), .B(n9597), .Z(n9602) );
  NANDN U10059 ( .A(n9600), .B(n9599), .Z(n9601) );
  AND U10060 ( .A(n9602), .B(n9601), .Z(n9702) );
  AND U10061 ( .A(x[135]), .B(y[742]), .Z(n9604) );
  AND U10062 ( .A(x[132]), .B(y[739]), .Z(n9603) );
  NAND U10063 ( .A(n9604), .B(n9603), .Z(n9608) );
  NAND U10064 ( .A(n9606), .B(n9605), .Z(n9607) );
  AND U10065 ( .A(n9608), .B(n9607), .Z(n9700) );
  AND U10066 ( .A(x[138]), .B(y[746]), .Z(n10360) );
  NAND U10067 ( .A(n10360), .B(n9959), .Z(n9612) );
  NAND U10068 ( .A(n9610), .B(n9609), .Z(n9611) );
  AND U10069 ( .A(n9612), .B(n9611), .Z(n9696) );
  AND U10070 ( .A(y[747]), .B(x[128]), .Z(n9614) );
  NAND U10071 ( .A(y[736]), .B(x[139]), .Z(n9613) );
  XNOR U10072 ( .A(n9614), .B(n9613), .Z(n9673) );
  ANDN U10073 ( .B(o[106]), .A(n9615), .Z(n9672) );
  XOR U10074 ( .A(n9673), .B(n9672), .Z(n9694) );
  AND U10075 ( .A(y[746]), .B(x[129]), .Z(n9617) );
  NAND U10076 ( .A(y[741]), .B(x[134]), .Z(n9616) );
  XNOR U10077 ( .A(n9617), .B(n9616), .Z(n9663) );
  NAND U10078 ( .A(x[138]), .B(y[737]), .Z(n9681) );
  XNOR U10079 ( .A(o[107]), .B(n9681), .Z(n9662) );
  XOR U10080 ( .A(n9663), .B(n9662), .Z(n9693) );
  XOR U10081 ( .A(n9694), .B(n9693), .Z(n9695) );
  NAND U10082 ( .A(x[131]), .B(y[744]), .Z(n10638) );
  NAND U10083 ( .A(y[745]), .B(x[130]), .Z(n9618) );
  XNOR U10084 ( .A(n9619), .B(n9618), .Z(n9658) );
  AND U10085 ( .A(x[132]), .B(y[743]), .Z(n9657) );
  XNOR U10086 ( .A(n9658), .B(n9657), .Z(n9688) );
  XOR U10087 ( .A(n10638), .B(n9688), .Z(n9690) );
  AND U10088 ( .A(y[738]), .B(x[137]), .Z(n9621) );
  NAND U10089 ( .A(y[740]), .B(x[135]), .Z(n9620) );
  XNOR U10090 ( .A(n9621), .B(n9620), .Z(n9677) );
  AND U10091 ( .A(x[136]), .B(y[739]), .Z(n9676) );
  XNOR U10092 ( .A(n9677), .B(n9676), .Z(n9689) );
  XOR U10093 ( .A(n9690), .B(n9689), .Z(n9654) );
  NAND U10094 ( .A(x[131]), .B(y[745]), .Z(n9734) );
  AND U10095 ( .A(x[129]), .B(y[743]), .Z(n9954) );
  NANDN U10096 ( .A(n9734), .B(n9954), .Z(n9625) );
  NANDN U10097 ( .A(n9623), .B(n9622), .Z(n9624) );
  AND U10098 ( .A(n9625), .B(n9624), .Z(n9652) );
  NAND U10099 ( .A(n9817), .B(n9626), .Z(n9630) );
  NAND U10100 ( .A(n9628), .B(n9627), .Z(n9629) );
  NAND U10101 ( .A(n9630), .B(n9629), .Z(n9651) );
  NANDN U10102 ( .A(n9632), .B(n9631), .Z(n9636) );
  NAND U10103 ( .A(n9634), .B(n9633), .Z(n9635) );
  NAND U10104 ( .A(n9636), .B(n9635), .Z(n9682) );
  XOR U10105 ( .A(n9683), .B(n9682), .Z(n9685) );
  XNOR U10106 ( .A(n9684), .B(n9685), .Z(n9708) );
  XNOR U10107 ( .A(n9709), .B(n9708), .Z(n9710) );
  XOR U10108 ( .A(n9711), .B(n9710), .Z(n9707) );
  NANDN U10109 ( .A(n9637), .B(n9638), .Z(n9643) );
  NOR U10110 ( .A(n9639), .B(n9638), .Z(n9641) );
  OR U10111 ( .A(n9641), .B(n9640), .Z(n9642) );
  AND U10112 ( .A(n9643), .B(n9642), .Z(n9705) );
  NAND U10113 ( .A(n9645), .B(n9644), .Z(n9649) );
  NANDN U10114 ( .A(n9647), .B(n9646), .Z(n9648) );
  AND U10115 ( .A(n9649), .B(n9648), .Z(n9706) );
  XOR U10116 ( .A(n9705), .B(n9706), .Z(n9650) );
  XNOR U10117 ( .A(n9707), .B(n9650), .Z(N236) );
  NANDN U10118 ( .A(n9652), .B(n9651), .Z(n9656) );
  NANDN U10119 ( .A(n9654), .B(n9653), .Z(n9655) );
  AND U10120 ( .A(n9656), .B(n9655), .Z(n9776) );
  AND U10121 ( .A(x[133]), .B(y[745]), .Z(n10194) );
  NAND U10122 ( .A(n10354), .B(n10194), .Z(n9660) );
  NAND U10123 ( .A(n9658), .B(n9657), .Z(n9659) );
  AND U10124 ( .A(n9660), .B(n9659), .Z(n9722) );
  AND U10125 ( .A(x[134]), .B(y[746]), .Z(n9971) );
  NAND U10126 ( .A(n9971), .B(n9661), .Z(n9665) );
  NAND U10127 ( .A(n9663), .B(n9662), .Z(n9664) );
  NAND U10128 ( .A(n9665), .B(n9664), .Z(n9721) );
  XNOR U10129 ( .A(n9722), .B(n9721), .Z(n9724) );
  AND U10130 ( .A(x[137]), .B(y[739]), .Z(n10349) );
  AND U10131 ( .A(y[744]), .B(x[132]), .Z(n9667) );
  NAND U10132 ( .A(y[738]), .B(x[138]), .Z(n9666) );
  XOR U10133 ( .A(n9667), .B(n9666), .Z(n9766) );
  NAND U10134 ( .A(x[135]), .B(y[741]), .Z(n9742) );
  XOR U10135 ( .A(n9743), .B(n9742), .Z(n9745) );
  AND U10136 ( .A(y[748]), .B(x[128]), .Z(n9669) );
  NAND U10137 ( .A(y[736]), .B(x[140]), .Z(n9668) );
  XNOR U10138 ( .A(n9669), .B(n9668), .Z(n9759) );
  NAND U10139 ( .A(x[139]), .B(y[737]), .Z(n9739) );
  XNOR U10140 ( .A(o[108]), .B(n9739), .Z(n9758) );
  XOR U10141 ( .A(n9759), .B(n9758), .Z(n9728) );
  AND U10142 ( .A(y[746]), .B(x[130]), .Z(n9671) );
  NAND U10143 ( .A(y[740]), .B(x[136]), .Z(n9670) );
  XNOR U10144 ( .A(n9671), .B(n9670), .Z(n9733) );
  XOR U10145 ( .A(n9728), .B(n9727), .Z(n9730) );
  XOR U10146 ( .A(n9729), .B(n9730), .Z(n9723) );
  XOR U10147 ( .A(n9724), .B(n9723), .Z(n9774) );
  AND U10148 ( .A(x[139]), .B(y[747]), .Z(n10748) );
  NAND U10149 ( .A(n10748), .B(n9959), .Z(n9675) );
  NAND U10150 ( .A(n9673), .B(n9672), .Z(n9674) );
  AND U10151 ( .A(n9675), .B(n9674), .Z(n9751) );
  AND U10152 ( .A(x[135]), .B(y[738]), .Z(n9913) );
  AND U10153 ( .A(x[137]), .B(y[740]), .Z(n9741) );
  NAND U10154 ( .A(n9913), .B(n9741), .Z(n9679) );
  NAND U10155 ( .A(n9677), .B(n9676), .Z(n9678) );
  AND U10156 ( .A(n9679), .B(n9678), .Z(n9749) );
  AND U10157 ( .A(y[747]), .B(x[129]), .Z(n10399) );
  NAND U10158 ( .A(y[742]), .B(x[134]), .Z(n9680) );
  XNOR U10159 ( .A(n10399), .B(n9680), .Z(n9755) );
  ANDN U10160 ( .B(o[107]), .A(n9681), .Z(n9754) );
  XOR U10161 ( .A(n9755), .B(n9754), .Z(n9748) );
  XNOR U10162 ( .A(n9749), .B(n9748), .Z(n9750) );
  XNOR U10163 ( .A(n9751), .B(n9750), .Z(n9773) );
  XOR U10164 ( .A(n9774), .B(n9773), .Z(n9775) );
  NAND U10165 ( .A(n9683), .B(n9682), .Z(n9687) );
  NAND U10166 ( .A(n9685), .B(n9684), .Z(n9686) );
  NAND U10167 ( .A(n9687), .B(n9686), .Z(n9779) );
  XOR U10168 ( .A(n9780), .B(n9779), .Z(n9782) );
  IV U10169 ( .A(n10638), .Z(n10363) );
  NANDN U10170 ( .A(n10363), .B(n9688), .Z(n9692) );
  NAND U10171 ( .A(n9690), .B(n9689), .Z(n9691) );
  AND U10172 ( .A(n9692), .B(n9691), .Z(n9716) );
  NAND U10173 ( .A(n9694), .B(n9693), .Z(n9698) );
  NANDN U10174 ( .A(n9696), .B(n9695), .Z(n9697) );
  AND U10175 ( .A(n9698), .B(n9697), .Z(n9715) );
  NANDN U10176 ( .A(n9700), .B(n9699), .Z(n9704) );
  NANDN U10177 ( .A(n9702), .B(n9701), .Z(n9703) );
  NAND U10178 ( .A(n9704), .B(n9703), .Z(n9718) );
  XNOR U10179 ( .A(n9782), .B(n9781), .Z(n9788) );
  NANDN U10180 ( .A(n9709), .B(n9708), .Z(n9713) );
  NANDN U10181 ( .A(n9711), .B(n9710), .Z(n9712) );
  AND U10182 ( .A(n9713), .B(n9712), .Z(n9787) );
  IV U10183 ( .A(n9787), .Z(n9785) );
  XOR U10184 ( .A(n9786), .B(n9785), .Z(n9714) );
  XNOR U10185 ( .A(n9788), .B(n9714), .Z(N237) );
  NANDN U10186 ( .A(n9716), .B(n9715), .Z(n9720) );
  NANDN U10187 ( .A(n9718), .B(n9717), .Z(n9719) );
  AND U10188 ( .A(n9720), .B(n9719), .Z(n9862) );
  NANDN U10189 ( .A(n9722), .B(n9721), .Z(n9726) );
  NAND U10190 ( .A(n9724), .B(n9723), .Z(n9725) );
  AND U10191 ( .A(n9726), .B(n9725), .Z(n9794) );
  NAND U10192 ( .A(n9728), .B(n9727), .Z(n9732) );
  NAND U10193 ( .A(n9730), .B(n9729), .Z(n9731) );
  NAND U10194 ( .A(n9732), .B(n9731), .Z(n9801) );
  AND U10195 ( .A(x[136]), .B(y[746]), .Z(n10991) );
  AND U10196 ( .A(x[130]), .B(y[740]), .Z(n9922) );
  NAND U10197 ( .A(n10991), .B(n9922), .Z(n9736) );
  NANDN U10198 ( .A(n9734), .B(n9733), .Z(n9735) );
  AND U10199 ( .A(n9736), .B(n9735), .Z(n9833) );
  AND U10200 ( .A(y[748]), .B(x[129]), .Z(n9738) );
  NAND U10201 ( .A(y[742]), .B(x[135]), .Z(n9737) );
  XNOR U10202 ( .A(n9738), .B(n9737), .Z(n9824) );
  ANDN U10203 ( .B(o[108]), .A(n9739), .Z(n9823) );
  XOR U10204 ( .A(n9824), .B(n9823), .Z(n9831) );
  AND U10205 ( .A(x[134]), .B(y[743]), .Z(n10787) );
  NAND U10206 ( .A(y[747]), .B(x[130]), .Z(n9740) );
  XOR U10207 ( .A(n9741), .B(n9740), .Z(n9836) );
  XNOR U10208 ( .A(n10787), .B(n9836), .Z(n9830) );
  XOR U10209 ( .A(n9831), .B(n9830), .Z(n9832) );
  XNOR U10210 ( .A(n9833), .B(n9832), .Z(n9800) );
  NAND U10211 ( .A(n9743), .B(n9742), .Z(n9747) );
  ANDN U10212 ( .B(n9745), .A(n9744), .Z(n9746) );
  ANDN U10213 ( .B(n9747), .A(n9746), .Z(n9799) );
  XOR U10214 ( .A(n9800), .B(n9799), .Z(n9802) );
  XOR U10215 ( .A(n9801), .B(n9802), .Z(n9793) );
  XNOR U10216 ( .A(n9794), .B(n9793), .Z(n9796) );
  NANDN U10217 ( .A(n9749), .B(n9748), .Z(n9753) );
  NANDN U10218 ( .A(n9751), .B(n9750), .Z(n9752) );
  AND U10219 ( .A(n9753), .B(n9752), .Z(n9808) );
  NAND U10220 ( .A(x[134]), .B(y[747]), .Z(n10196) );
  AND U10221 ( .A(x[129]), .B(y[742]), .Z(n9822) );
  NANDN U10222 ( .A(n10196), .B(n9822), .Z(n9757) );
  NAND U10223 ( .A(n9755), .B(n9754), .Z(n9756) );
  AND U10224 ( .A(n9757), .B(n9756), .Z(n9814) );
  AND U10225 ( .A(x[140]), .B(y[748]), .Z(n10997) );
  NAND U10226 ( .A(n10997), .B(n9959), .Z(n9761) );
  NAND U10227 ( .A(n9759), .B(n9758), .Z(n9760) );
  AND U10228 ( .A(n9761), .B(n9760), .Z(n9812) );
  AND U10229 ( .A(x[138]), .B(y[739]), .Z(n10650) );
  AND U10230 ( .A(y[741]), .B(x[136]), .Z(n9763) );
  NAND U10231 ( .A(y[738]), .B(x[139]), .Z(n9762) );
  XOR U10232 ( .A(n9763), .B(n9762), .Z(n9819) );
  XNOR U10233 ( .A(n10650), .B(n9819), .Z(n9811) );
  XNOR U10234 ( .A(n9812), .B(n9811), .Z(n9813) );
  XNOR U10235 ( .A(n9814), .B(n9813), .Z(n9806) );
  AND U10236 ( .A(x[138]), .B(y[744]), .Z(n9765) );
  AND U10237 ( .A(x[132]), .B(y[738]), .Z(n9764) );
  NAND U10238 ( .A(n9765), .B(n9764), .Z(n9768) );
  NANDN U10239 ( .A(n9766), .B(n10349), .Z(n9767) );
  AND U10240 ( .A(n9768), .B(n9767), .Z(n9856) );
  AND U10241 ( .A(y[749]), .B(x[128]), .Z(n9770) );
  NAND U10242 ( .A(y[736]), .B(x[141]), .Z(n9769) );
  XNOR U10243 ( .A(n9770), .B(n9769), .Z(n9848) );
  NAND U10244 ( .A(x[140]), .B(y[737]), .Z(n9841) );
  XNOR U10245 ( .A(o[109]), .B(n9841), .Z(n9847) );
  XOR U10246 ( .A(n9848), .B(n9847), .Z(n9854) );
  AND U10247 ( .A(y[744]), .B(x[133]), .Z(n9772) );
  NAND U10248 ( .A(y[746]), .B(x[131]), .Z(n9771) );
  XNOR U10249 ( .A(n9772), .B(n9771), .Z(n9843) );
  NAND U10250 ( .A(x[132]), .B(y[745]), .Z(n9844) );
  XNOR U10251 ( .A(n9843), .B(n9844), .Z(n9853) );
  XOR U10252 ( .A(n9854), .B(n9853), .Z(n9855) );
  XOR U10253 ( .A(n9806), .B(n9805), .Z(n9807) );
  XOR U10254 ( .A(n9796), .B(n9795), .Z(n9860) );
  NAND U10255 ( .A(n9774), .B(n9773), .Z(n9778) );
  NANDN U10256 ( .A(n9776), .B(n9775), .Z(n9777) );
  AND U10257 ( .A(n9778), .B(n9777), .Z(n9859) );
  XOR U10258 ( .A(n9862), .B(n9861), .Z(n9867) );
  NAND U10259 ( .A(n9780), .B(n9779), .Z(n9784) );
  NAND U10260 ( .A(n9782), .B(n9781), .Z(n9783) );
  NAND U10261 ( .A(n9784), .B(n9783), .Z(n9865) );
  NANDN U10262 ( .A(n9785), .B(n9786), .Z(n9791) );
  NOR U10263 ( .A(n9787), .B(n9786), .Z(n9789) );
  OR U10264 ( .A(n9789), .B(n9788), .Z(n9790) );
  AND U10265 ( .A(n9791), .B(n9790), .Z(n9866) );
  XOR U10266 ( .A(n9865), .B(n9866), .Z(n9792) );
  XNOR U10267 ( .A(n9867), .B(n9792), .Z(N238) );
  NANDN U10268 ( .A(n9794), .B(n9793), .Z(n9798) );
  NAND U10269 ( .A(n9796), .B(n9795), .Z(n9797) );
  AND U10270 ( .A(n9798), .B(n9797), .Z(n9945) );
  NAND U10271 ( .A(n9800), .B(n9799), .Z(n9804) );
  NAND U10272 ( .A(n9802), .B(n9801), .Z(n9803) );
  NAND U10273 ( .A(n9804), .B(n9803), .Z(n9944) );
  XNOR U10274 ( .A(n9945), .B(n9944), .Z(n9947) );
  NAND U10275 ( .A(n9806), .B(n9805), .Z(n9810) );
  NANDN U10276 ( .A(n9808), .B(n9807), .Z(n9809) );
  AND U10277 ( .A(n9810), .B(n9809), .Z(n9872) );
  NANDN U10278 ( .A(n9812), .B(n9811), .Z(n9816) );
  NANDN U10279 ( .A(n9814), .B(n9813), .Z(n9815) );
  AND U10280 ( .A(n9816), .B(n9815), .Z(n9935) );
  AND U10281 ( .A(x[139]), .B(y[741]), .Z(n9818) );
  NAND U10282 ( .A(n9818), .B(n9817), .Z(n9821) );
  NANDN U10283 ( .A(n9819), .B(n10650), .Z(n9820) );
  AND U10284 ( .A(n9821), .B(n9820), .Z(n9896) );
  NAND U10285 ( .A(x[135]), .B(y[748]), .Z(n10365) );
  NANDN U10286 ( .A(n10365), .B(n9822), .Z(n9826) );
  NAND U10287 ( .A(n9824), .B(n9823), .Z(n9825) );
  NAND U10288 ( .A(n9826), .B(n9825), .Z(n9895) );
  XNOR U10289 ( .A(n9896), .B(n9895), .Z(n9898) );
  AND U10290 ( .A(x[132]), .B(y[746]), .Z(n10287) );
  AND U10291 ( .A(y[747]), .B(x[131]), .Z(n9828) );
  NAND U10292 ( .A(y[742]), .B(x[136]), .Z(n9827) );
  XOR U10293 ( .A(n9828), .B(n9827), .Z(n9881) );
  XNOR U10294 ( .A(n10194), .B(n9881), .Z(n9890) );
  XOR U10295 ( .A(n10287), .B(n9890), .Z(n9892) );
  AND U10296 ( .A(x[137]), .B(y[741]), .Z(n10465) );
  AND U10297 ( .A(y[748]), .B(x[130]), .Z(n9829) );
  AND U10298 ( .A(y[740]), .B(x[138]), .Z(n10495) );
  XOR U10299 ( .A(n9829), .B(n10495), .Z(n9923) );
  XOR U10300 ( .A(n10465), .B(n9923), .Z(n9891) );
  XOR U10301 ( .A(n9892), .B(n9891), .Z(n9897) );
  XOR U10302 ( .A(n9898), .B(n9897), .Z(n9933) );
  NAND U10303 ( .A(n9831), .B(n9830), .Z(n9835) );
  NANDN U10304 ( .A(n9833), .B(n9832), .Z(n9834) );
  AND U10305 ( .A(n9835), .B(n9834), .Z(n9932) );
  XNOR U10306 ( .A(n9933), .B(n9932), .Z(n9934) );
  XOR U10307 ( .A(n9935), .B(n9934), .Z(n9870) );
  AND U10308 ( .A(x[137]), .B(y[747]), .Z(n10362) );
  NAND U10309 ( .A(n10362), .B(n9922), .Z(n9838) );
  NANDN U10310 ( .A(n9836), .B(n10787), .Z(n9837) );
  AND U10311 ( .A(n9838), .B(n9837), .Z(n9910) );
  AND U10312 ( .A(y[750]), .B(x[128]), .Z(n9840) );
  NAND U10313 ( .A(y[736]), .B(x[142]), .Z(n9839) );
  XNOR U10314 ( .A(n9840), .B(n9839), .Z(n9876) );
  ANDN U10315 ( .B(o[109]), .A(n9841), .Z(n9875) );
  XOR U10316 ( .A(n9876), .B(n9875), .Z(n9908) );
  AND U10317 ( .A(y[738]), .B(x[140]), .Z(n10455) );
  NAND U10318 ( .A(y[743]), .B(x[135]), .Z(n9842) );
  XNOR U10319 ( .A(n10455), .B(n9842), .Z(n9914) );
  NAND U10320 ( .A(x[141]), .B(y[737]), .Z(n9921) );
  XOR U10321 ( .A(o[110]), .B(n9921), .Z(n9915) );
  XNOR U10322 ( .A(n9914), .B(n9915), .Z(n9907) );
  XOR U10323 ( .A(n9908), .B(n9907), .Z(n9909) );
  XOR U10324 ( .A(n9910), .B(n9909), .Z(n9939) );
  AND U10325 ( .A(x[133]), .B(y[746]), .Z(n9972) );
  NANDN U10326 ( .A(n10638), .B(n9972), .Z(n9846) );
  NANDN U10327 ( .A(n9844), .B(n9843), .Z(n9845) );
  AND U10328 ( .A(n9846), .B(n9845), .Z(n9904) );
  AND U10329 ( .A(x[141]), .B(y[749]), .Z(n11388) );
  NAND U10330 ( .A(n11388), .B(n9959), .Z(n9850) );
  NAND U10331 ( .A(n9848), .B(n9847), .Z(n9849) );
  AND U10332 ( .A(n9850), .B(n9849), .Z(n9902) );
  NAND U10333 ( .A(y[739]), .B(x[139]), .Z(n9851) );
  XNOR U10334 ( .A(n9852), .B(n9851), .Z(n9928) );
  NAND U10335 ( .A(x[129]), .B(y[749]), .Z(n9929) );
  XNOR U10336 ( .A(n9928), .B(n9929), .Z(n9901) );
  XNOR U10337 ( .A(n9902), .B(n9901), .Z(n9903) );
  XOR U10338 ( .A(n9904), .B(n9903), .Z(n9938) );
  XOR U10339 ( .A(n9939), .B(n9938), .Z(n9941) );
  NAND U10340 ( .A(n9854), .B(n9853), .Z(n9858) );
  NANDN U10341 ( .A(n9856), .B(n9855), .Z(n9857) );
  AND U10342 ( .A(n9858), .B(n9857), .Z(n9940) );
  XNOR U10343 ( .A(n9941), .B(n9940), .Z(n9869) );
  XOR U10344 ( .A(n9947), .B(n9946), .Z(n9952) );
  NANDN U10345 ( .A(n9860), .B(n9859), .Z(n9864) );
  NANDN U10346 ( .A(n9862), .B(n9861), .Z(n9863) );
  NAND U10347 ( .A(n9864), .B(n9863), .Z(n9950) );
  XOR U10348 ( .A(n9950), .B(n9951), .Z(n9868) );
  XNOR U10349 ( .A(n9952), .B(n9868), .Z(N239) );
  NANDN U10350 ( .A(n9870), .B(n9869), .Z(n9874) );
  NANDN U10351 ( .A(n9872), .B(n9871), .Z(n9873) );
  AND U10352 ( .A(n9874), .B(n9873), .Z(n10042) );
  AND U10353 ( .A(x[142]), .B(y[750]), .Z(n11649) );
  NAND U10354 ( .A(n11649), .B(n9959), .Z(n9878) );
  NAND U10355 ( .A(n9876), .B(n9875), .Z(n9877) );
  AND U10356 ( .A(n9878), .B(n9877), .Z(n9987) );
  AND U10357 ( .A(x[136]), .B(y[747]), .Z(n9879) );
  NANDN U10358 ( .A(n9880), .B(n9879), .Z(n9883) );
  NANDN U10359 ( .A(n9881), .B(n10194), .Z(n9882) );
  NAND U10360 ( .A(n9883), .B(n9882), .Z(n9986) );
  XNOR U10361 ( .A(n9987), .B(n9986), .Z(n9989) );
  AND U10362 ( .A(y[747]), .B(x[132]), .Z(n9885) );
  NAND U10363 ( .A(y[741]), .B(x[138]), .Z(n9884) );
  XNOR U10364 ( .A(n9885), .B(n9884), .Z(n9967) );
  AND U10365 ( .A(x[135]), .B(y[744]), .Z(n9966) );
  XOR U10366 ( .A(n9967), .B(n9966), .Z(n9974) );
  NAND U10367 ( .A(x[134]), .B(y[745]), .Z(n10073) );
  XNOR U10368 ( .A(n10073), .B(n9972), .Z(n9973) );
  XNOR U10369 ( .A(n9974), .B(n9973), .Z(n10009) );
  AND U10370 ( .A(y[742]), .B(x[137]), .Z(n9887) );
  NAND U10371 ( .A(y[749]), .B(x[130]), .Z(n9886) );
  XNOR U10372 ( .A(n9887), .B(n9886), .Z(n9977) );
  NAND U10373 ( .A(x[131]), .B(y[748]), .Z(n9978) );
  XNOR U10374 ( .A(n9977), .B(n9978), .Z(n10007) );
  AND U10375 ( .A(y[750]), .B(x[129]), .Z(n9889) );
  NAND U10376 ( .A(y[743]), .B(x[136]), .Z(n9888) );
  XNOR U10377 ( .A(n9889), .B(n9888), .Z(n9956) );
  NAND U10378 ( .A(x[142]), .B(y[737]), .Z(n9983) );
  XNOR U10379 ( .A(o[111]), .B(n9983), .Z(n9955) );
  XOR U10380 ( .A(n9956), .B(n9955), .Z(n10006) );
  XOR U10381 ( .A(n10007), .B(n10006), .Z(n10008) );
  XNOR U10382 ( .A(n10009), .B(n10008), .Z(n9988) );
  XOR U10383 ( .A(n9989), .B(n9988), .Z(n10031) );
  NAND U10384 ( .A(n10287), .B(n9890), .Z(n9894) );
  NAND U10385 ( .A(n9892), .B(n9891), .Z(n9893) );
  AND U10386 ( .A(n9894), .B(n9893), .Z(n10030) );
  XNOR U10387 ( .A(n10031), .B(n10030), .Z(n10033) );
  NANDN U10388 ( .A(n9896), .B(n9895), .Z(n9900) );
  NAND U10389 ( .A(n9898), .B(n9897), .Z(n9899) );
  AND U10390 ( .A(n9900), .B(n9899), .Z(n10032) );
  XOR U10391 ( .A(n10033), .B(n10032), .Z(n10013) );
  NANDN U10392 ( .A(n9902), .B(n9901), .Z(n9906) );
  NANDN U10393 ( .A(n9904), .B(n9903), .Z(n9905) );
  AND U10394 ( .A(n9906), .B(n9905), .Z(n10021) );
  NAND U10395 ( .A(n9908), .B(n9907), .Z(n9912) );
  NANDN U10396 ( .A(n9910), .B(n9909), .Z(n9911) );
  AND U10397 ( .A(n9912), .B(n9911), .Z(n10019) );
  NAND U10398 ( .A(x[140]), .B(y[743]), .Z(n10356) );
  NANDN U10399 ( .A(n10356), .B(n9913), .Z(n9917) );
  NANDN U10400 ( .A(n9915), .B(n9914), .Z(n9916) );
  AND U10401 ( .A(n9917), .B(n9916), .Z(n9995) );
  AND U10402 ( .A(y[738]), .B(x[141]), .Z(n10775) );
  NAND U10403 ( .A(y[740]), .B(x[139]), .Z(n9918) );
  XNOR U10404 ( .A(n10775), .B(n9918), .Z(n9999) );
  AND U10405 ( .A(x[140]), .B(y[739]), .Z(n9998) );
  XOR U10406 ( .A(n9999), .B(n9998), .Z(n9993) );
  AND U10407 ( .A(y[751]), .B(x[128]), .Z(n9920) );
  NAND U10408 ( .A(y[736]), .B(x[143]), .Z(n9919) );
  XNOR U10409 ( .A(n9920), .B(n9919), .Z(n9961) );
  ANDN U10410 ( .B(o[110]), .A(n9921), .Z(n9960) );
  XNOR U10411 ( .A(n9961), .B(n9960), .Z(n9992) );
  XNOR U10412 ( .A(n9993), .B(n9992), .Z(n9994) );
  XOR U10413 ( .A(n9995), .B(n9994), .Z(n10027) );
  AND U10414 ( .A(x[138]), .B(y[748]), .Z(n10637) );
  IV U10415 ( .A(n10637), .Z(n10789) );
  NANDN U10416 ( .A(n10789), .B(n9922), .Z(n9925) );
  NAND U10417 ( .A(n10465), .B(n9923), .Z(n9924) );
  AND U10418 ( .A(n9925), .B(n9924), .Z(n10025) );
  AND U10419 ( .A(x[139]), .B(y[744]), .Z(n9927) );
  AND U10420 ( .A(x[134]), .B(y[739]), .Z(n9926) );
  NAND U10421 ( .A(n9927), .B(n9926), .Z(n9931) );
  NANDN U10422 ( .A(n9929), .B(n9928), .Z(n9930) );
  NAND U10423 ( .A(n9931), .B(n9930), .Z(n10024) );
  XNOR U10424 ( .A(n10025), .B(n10024), .Z(n10026) );
  XNOR U10425 ( .A(n10027), .B(n10026), .Z(n10018) );
  XNOR U10426 ( .A(n10019), .B(n10018), .Z(n10020) );
  XNOR U10427 ( .A(n10021), .B(n10020), .Z(n10012) );
  XNOR U10428 ( .A(n10013), .B(n10012), .Z(n10014) );
  NANDN U10429 ( .A(n9933), .B(n9932), .Z(n9937) );
  NAND U10430 ( .A(n9935), .B(n9934), .Z(n9936) );
  NAND U10431 ( .A(n9937), .B(n9936), .Z(n10015) );
  XNOR U10432 ( .A(n10014), .B(n10015), .Z(n10039) );
  NAND U10433 ( .A(n9939), .B(n9938), .Z(n9943) );
  NAND U10434 ( .A(n9941), .B(n9940), .Z(n9942) );
  NAND U10435 ( .A(n9943), .B(n9942), .Z(n10040) );
  XOR U10436 ( .A(n10042), .B(n10041), .Z(n10038) );
  NANDN U10437 ( .A(n9945), .B(n9944), .Z(n9949) );
  NAND U10438 ( .A(n9947), .B(n9946), .Z(n9948) );
  NAND U10439 ( .A(n9949), .B(n9948), .Z(n10037) );
  XOR U10440 ( .A(n10037), .B(n10036), .Z(n9953) );
  XNOR U10441 ( .A(n10038), .B(n9953), .Z(N240) );
  AND U10442 ( .A(x[136]), .B(y[750]), .Z(n10659) );
  NAND U10443 ( .A(n10659), .B(n9954), .Z(n9958) );
  NAND U10444 ( .A(n9956), .B(n9955), .Z(n9957) );
  NAND U10445 ( .A(n9958), .B(n9957), .Z(n10100) );
  AND U10446 ( .A(x[143]), .B(y[751]), .Z(n12002) );
  NAND U10447 ( .A(n12002), .B(n9959), .Z(n9963) );
  NAND U10448 ( .A(n9961), .B(n9960), .Z(n9962) );
  NAND U10449 ( .A(n9963), .B(n9962), .Z(n10101) );
  XOR U10450 ( .A(n10100), .B(n10101), .Z(n10103) );
  AND U10451 ( .A(x[138]), .B(y[747]), .Z(n9965) );
  NAND U10452 ( .A(n9965), .B(n9964), .Z(n9969) );
  NAND U10453 ( .A(n9967), .B(n9966), .Z(n9968) );
  NAND U10454 ( .A(n9969), .B(n9968), .Z(n10060) );
  AND U10455 ( .A(x[128]), .B(y[752]), .Z(n10080) );
  NAND U10456 ( .A(x[144]), .B(y[736]), .Z(n10081) );
  XNOR U10457 ( .A(n10080), .B(n10081), .Z(n10082) );
  NAND U10458 ( .A(x[143]), .B(y[737]), .Z(n10070) );
  XOR U10459 ( .A(o[112]), .B(n10070), .Z(n10083) );
  XNOR U10460 ( .A(n10082), .B(n10083), .Z(n10059) );
  NAND U10461 ( .A(y[745]), .B(x[135]), .Z(n9970) );
  XNOR U10462 ( .A(n9971), .B(n9970), .Z(n10075) );
  AND U10463 ( .A(x[138]), .B(y[742]), .Z(n10074) );
  XOR U10464 ( .A(n10075), .B(n10074), .Z(n10058) );
  XOR U10465 ( .A(n10059), .B(n10058), .Z(n10061) );
  XOR U10466 ( .A(n10060), .B(n10061), .Z(n10102) );
  XOR U10467 ( .A(n10103), .B(n10102), .Z(n10055) );
  NANDN U10468 ( .A(n9972), .B(n10073), .Z(n9976) );
  NANDN U10469 ( .A(n9974), .B(n9973), .Z(n9975) );
  AND U10470 ( .A(n9976), .B(n9975), .Z(n10053) );
  AND U10471 ( .A(x[137]), .B(y[749]), .Z(n10770) );
  NAND U10472 ( .A(n10770), .B(n10354), .Z(n9980) );
  NANDN U10473 ( .A(n9978), .B(n9977), .Z(n9979) );
  NAND U10474 ( .A(n9980), .B(n9979), .Z(n10090) );
  AND U10475 ( .A(y[751]), .B(x[129]), .Z(n9982) );
  NAND U10476 ( .A(y[744]), .B(x[136]), .Z(n9981) );
  XNOR U10477 ( .A(n9982), .B(n9981), .Z(n10079) );
  ANDN U10478 ( .B(o[111]), .A(n9983), .Z(n10078) );
  XOR U10479 ( .A(n10079), .B(n10078), .Z(n10089) );
  AND U10480 ( .A(y[738]), .B(x[142]), .Z(n9985) );
  NAND U10481 ( .A(y[741]), .B(x[139]), .Z(n9984) );
  XNOR U10482 ( .A(n9985), .B(n9984), .Z(n10108) );
  NAND U10483 ( .A(x[132]), .B(y[748]), .Z(n10109) );
  XNOR U10484 ( .A(n10108), .B(n10109), .Z(n10088) );
  XOR U10485 ( .A(n10089), .B(n10088), .Z(n10091) );
  XNOR U10486 ( .A(n10090), .B(n10091), .Z(n10052) );
  XNOR U10487 ( .A(n10053), .B(n10052), .Z(n10054) );
  XNOR U10488 ( .A(n10055), .B(n10054), .Z(n10094) );
  NANDN U10489 ( .A(n9987), .B(n9986), .Z(n9991) );
  NAND U10490 ( .A(n9989), .B(n9988), .Z(n9990) );
  NAND U10491 ( .A(n9991), .B(n9990), .Z(n10095) );
  XNOR U10492 ( .A(n10094), .B(n10095), .Z(n10097) );
  NANDN U10493 ( .A(n9993), .B(n9992), .Z(n9997) );
  NAND U10494 ( .A(n9995), .B(n9994), .Z(n9996) );
  NAND U10495 ( .A(n9997), .B(n9996), .Z(n10122) );
  AND U10496 ( .A(x[139]), .B(y[738]), .Z(n10660) );
  AND U10497 ( .A(x[141]), .B(y[740]), .Z(n10119) );
  NAND U10498 ( .A(n10660), .B(n10119), .Z(n10001) );
  NAND U10499 ( .A(n9999), .B(n9998), .Z(n10000) );
  NAND U10500 ( .A(n10001), .B(n10000), .Z(n10106) );
  AND U10501 ( .A(y[743]), .B(x[137]), .Z(n10003) );
  NAND U10502 ( .A(y[750]), .B(x[130]), .Z(n10002) );
  XNOR U10503 ( .A(n10003), .B(n10002), .Z(n10113) );
  NAND U10504 ( .A(x[131]), .B(y[749]), .Z(n10114) );
  XNOR U10505 ( .A(n10113), .B(n10114), .Z(n10105) );
  AND U10506 ( .A(x[140]), .B(y[740]), .Z(n10759) );
  AND U10507 ( .A(y[747]), .B(x[133]), .Z(n10005) );
  NAND U10508 ( .A(y[739]), .B(x[141]), .Z(n10004) );
  XNOR U10509 ( .A(n10005), .B(n10004), .Z(n10065) );
  XOR U10510 ( .A(n10759), .B(n10065), .Z(n10104) );
  XOR U10511 ( .A(n10105), .B(n10104), .Z(n10107) );
  XOR U10512 ( .A(n10106), .B(n10107), .Z(n10121) );
  NAND U10513 ( .A(n10007), .B(n10006), .Z(n10011) );
  NANDN U10514 ( .A(n10009), .B(n10008), .Z(n10010) );
  AND U10515 ( .A(n10011), .B(n10010), .Z(n10120) );
  XNOR U10516 ( .A(n10121), .B(n10120), .Z(n10123) );
  XOR U10517 ( .A(n10122), .B(n10123), .Z(n10096) );
  XOR U10518 ( .A(n10097), .B(n10096), .Z(n10134) );
  NANDN U10519 ( .A(n10013), .B(n10012), .Z(n10017) );
  NANDN U10520 ( .A(n10015), .B(n10014), .Z(n10016) );
  NAND U10521 ( .A(n10017), .B(n10016), .Z(n10133) );
  XNOR U10522 ( .A(n10134), .B(n10133), .Z(n10136) );
  NANDN U10523 ( .A(n10019), .B(n10018), .Z(n10023) );
  NANDN U10524 ( .A(n10021), .B(n10020), .Z(n10022) );
  AND U10525 ( .A(n10023), .B(n10022), .Z(n10049) );
  NANDN U10526 ( .A(n10025), .B(n10024), .Z(n10029) );
  NANDN U10527 ( .A(n10027), .B(n10026), .Z(n10028) );
  AND U10528 ( .A(n10029), .B(n10028), .Z(n10047) );
  NANDN U10529 ( .A(n10031), .B(n10030), .Z(n10035) );
  NAND U10530 ( .A(n10033), .B(n10032), .Z(n10034) );
  AND U10531 ( .A(n10035), .B(n10034), .Z(n10046) );
  XNOR U10532 ( .A(n10047), .B(n10046), .Z(n10048) );
  XNOR U10533 ( .A(n10049), .B(n10048), .Z(n10135) );
  XNOR U10534 ( .A(n10136), .B(n10135), .Z(n10129) );
  NANDN U10535 ( .A(n10040), .B(n10039), .Z(n10044) );
  NANDN U10536 ( .A(n10042), .B(n10041), .Z(n10043) );
  NAND U10537 ( .A(n10044), .B(n10043), .Z(n10127) );
  IV U10538 ( .A(n10127), .Z(n10126) );
  XOR U10539 ( .A(n10128), .B(n10126), .Z(n10045) );
  XNOR U10540 ( .A(n10129), .B(n10045), .Z(N241) );
  NANDN U10541 ( .A(n10047), .B(n10046), .Z(n10051) );
  NANDN U10542 ( .A(n10049), .B(n10048), .Z(n10050) );
  AND U10543 ( .A(n10051), .B(n10050), .Z(n10229) );
  NANDN U10544 ( .A(n10053), .B(n10052), .Z(n10057) );
  NANDN U10545 ( .A(n10055), .B(n10054), .Z(n10056) );
  NAND U10546 ( .A(n10057), .B(n10056), .Z(n10148) );
  NAND U10547 ( .A(n10059), .B(n10058), .Z(n10063) );
  NAND U10548 ( .A(n10061), .B(n10060), .Z(n10062) );
  NAND U10549 ( .A(n10063), .B(n10062), .Z(n10224) );
  AND U10550 ( .A(x[141]), .B(y[747]), .Z(n11005) );
  NAND U10551 ( .A(n11005), .B(n10064), .Z(n10067) );
  NAND U10552 ( .A(n10759), .B(n10065), .Z(n10066) );
  AND U10553 ( .A(n10067), .B(n10066), .Z(n10181) );
  AND U10554 ( .A(y[744]), .B(x[137]), .Z(n10069) );
  NAND U10555 ( .A(y[752]), .B(x[129]), .Z(n10068) );
  XNOR U10556 ( .A(n10069), .B(n10068), .Z(n10200) );
  ANDN U10557 ( .B(o[112]), .A(n10070), .Z(n10199) );
  XOR U10558 ( .A(n10200), .B(n10199), .Z(n10179) );
  AND U10559 ( .A(y[738]), .B(x[143]), .Z(n10072) );
  NAND U10560 ( .A(y[741]), .B(x[140]), .Z(n10071) );
  XNOR U10561 ( .A(n10072), .B(n10071), .Z(n10153) );
  NAND U10562 ( .A(x[142]), .B(y[739]), .Z(n10154) );
  XNOR U10563 ( .A(n10153), .B(n10154), .Z(n10178) );
  XOR U10564 ( .A(n10179), .B(n10178), .Z(n10180) );
  XNOR U10565 ( .A(n10181), .B(n10180), .Z(n10223) );
  AND U10566 ( .A(x[135]), .B(y[746]), .Z(n10209) );
  NANDN U10567 ( .A(n10073), .B(n10209), .Z(n10077) );
  NAND U10568 ( .A(n10075), .B(n10074), .Z(n10076) );
  AND U10569 ( .A(n10077), .B(n10076), .Z(n10189) );
  AND U10570 ( .A(x[136]), .B(y[751]), .Z(n10752) );
  IV U10571 ( .A(n10752), .Z(n10911) );
  XNOR U10572 ( .A(n10189), .B(n10188), .Z(n10191) );
  NANDN U10573 ( .A(n10081), .B(n10080), .Z(n10085) );
  NANDN U10574 ( .A(n10083), .B(n10082), .Z(n10084) );
  AND U10575 ( .A(n10085), .B(n10084), .Z(n10185) );
  AND U10576 ( .A(x[128]), .B(y[753]), .Z(n10167) );
  NAND U10577 ( .A(x[145]), .B(y[736]), .Z(n10168) );
  XNOR U10578 ( .A(n10167), .B(n10168), .Z(n10169) );
  NAND U10579 ( .A(x[144]), .B(y[737]), .Z(n10164) );
  XOR U10580 ( .A(o[113]), .B(n10164), .Z(n10170) );
  XNOR U10581 ( .A(n10169), .B(n10170), .Z(n10182) );
  AND U10582 ( .A(y[751]), .B(x[130]), .Z(n10087) );
  NAND U10583 ( .A(y[743]), .B(x[138]), .Z(n10086) );
  XNOR U10584 ( .A(n10087), .B(n10086), .Z(n10202) );
  NAND U10585 ( .A(x[131]), .B(y[750]), .Z(n10203) );
  XOR U10586 ( .A(n10202), .B(n10203), .Z(n10183) );
  XNOR U10587 ( .A(n10182), .B(n10183), .Z(n10184) );
  XNOR U10588 ( .A(n10185), .B(n10184), .Z(n10190) );
  XOR U10589 ( .A(n10191), .B(n10190), .Z(n10222) );
  XOR U10590 ( .A(n10223), .B(n10222), .Z(n10225) );
  XOR U10591 ( .A(n10224), .B(n10225), .Z(n10147) );
  NAND U10592 ( .A(n10089), .B(n10088), .Z(n10093) );
  NAND U10593 ( .A(n10091), .B(n10090), .Z(n10092) );
  AND U10594 ( .A(n10093), .B(n10092), .Z(n10146) );
  XOR U10595 ( .A(n10147), .B(n10146), .Z(n10149) );
  XOR U10596 ( .A(n10148), .B(n10149), .Z(n10227) );
  NANDN U10597 ( .A(n10095), .B(n10094), .Z(n10099) );
  NAND U10598 ( .A(n10097), .B(n10096), .Z(n10098) );
  NAND U10599 ( .A(n10099), .B(n10098), .Z(n10142) );
  NAND U10600 ( .A(x[142]), .B(y[741]), .Z(n10401) );
  NANDN U10601 ( .A(n10401), .B(n10660), .Z(n10111) );
  NANDN U10602 ( .A(n10109), .B(n10108), .Z(n10110) );
  AND U10603 ( .A(n10111), .B(n10110), .Z(n10213) );
  AND U10604 ( .A(y[750]), .B(x[137]), .Z(n10986) );
  NANDN U10605 ( .A(n10112), .B(n10986), .Z(n10116) );
  NANDN U10606 ( .A(n10114), .B(n10113), .Z(n10115) );
  NAND U10607 ( .A(n10116), .B(n10115), .Z(n10212) );
  XNOR U10608 ( .A(n10213), .B(n10212), .Z(n10214) );
  AND U10609 ( .A(y[748]), .B(x[133]), .Z(n10254) );
  NAND U10610 ( .A(y[745]), .B(x[136]), .Z(n10117) );
  XNOR U10611 ( .A(n10254), .B(n10117), .Z(n10195) );
  XOR U10612 ( .A(n10209), .B(n10208), .Z(n10210) );
  NAND U10613 ( .A(y[749]), .B(x[132]), .Z(n10118) );
  XNOR U10614 ( .A(n10119), .B(n10118), .Z(n10158) );
  NAND U10615 ( .A(x[139]), .B(y[742]), .Z(n10159) );
  XOR U10616 ( .A(n10158), .B(n10159), .Z(n10211) );
  XOR U10617 ( .A(n10210), .B(n10211), .Z(n10215) );
  XNOR U10618 ( .A(n10214), .B(n10215), .Z(n10219) );
  XOR U10619 ( .A(n10218), .B(n10219), .Z(n10221) );
  XOR U10620 ( .A(n10220), .B(n10221), .Z(n10141) );
  NANDN U10621 ( .A(n10121), .B(n10120), .Z(n10125) );
  NAND U10622 ( .A(n10123), .B(n10122), .Z(n10124) );
  NAND U10623 ( .A(n10125), .B(n10124), .Z(n10140) );
  XOR U10624 ( .A(n10141), .B(n10140), .Z(n10143) );
  XOR U10625 ( .A(n10142), .B(n10143), .Z(n10226) );
  XOR U10626 ( .A(n10227), .B(n10226), .Z(n10228) );
  XNOR U10627 ( .A(n10229), .B(n10228), .Z(n10235) );
  OR U10628 ( .A(n10128), .B(n10126), .Z(n10132) );
  ANDN U10629 ( .B(n10128), .A(n10127), .Z(n10130) );
  OR U10630 ( .A(n10130), .B(n10129), .Z(n10131) );
  AND U10631 ( .A(n10132), .B(n10131), .Z(n10233) );
  NANDN U10632 ( .A(n10134), .B(n10133), .Z(n10138) );
  NAND U10633 ( .A(n10136), .B(n10135), .Z(n10137) );
  AND U10634 ( .A(n10138), .B(n10137), .Z(n10234) );
  IV U10635 ( .A(n10234), .Z(n10232) );
  XOR U10636 ( .A(n10233), .B(n10232), .Z(n10139) );
  XNOR U10637 ( .A(n10235), .B(n10139), .Z(N242) );
  NANDN U10638 ( .A(n10141), .B(n10140), .Z(n10145) );
  NANDN U10639 ( .A(n10143), .B(n10142), .Z(n10144) );
  AND U10640 ( .A(n10145), .B(n10144), .Z(n10333) );
  NANDN U10641 ( .A(n10147), .B(n10146), .Z(n10151) );
  NANDN U10642 ( .A(n10149), .B(n10148), .Z(n10150) );
  AND U10643 ( .A(n10151), .B(n10150), .Z(n10331) );
  AND U10644 ( .A(x[143]), .B(y[741]), .Z(n10152) );
  NAND U10645 ( .A(n10455), .B(n10152), .Z(n10156) );
  NANDN U10646 ( .A(n10154), .B(n10153), .Z(n10155) );
  AND U10647 ( .A(n10156), .B(n10155), .Z(n10310) );
  NAND U10648 ( .A(n11388), .B(n10157), .Z(n10161) );
  NANDN U10649 ( .A(n10159), .B(n10158), .Z(n10160) );
  NAND U10650 ( .A(n10161), .B(n10160), .Z(n10301) );
  AND U10651 ( .A(y[753]), .B(x[129]), .Z(n10163) );
  NAND U10652 ( .A(y[744]), .B(x[138]), .Z(n10162) );
  XNOR U10653 ( .A(n10163), .B(n10162), .Z(n10269) );
  ANDN U10654 ( .B(o[113]), .A(n10164), .Z(n10268) );
  XOR U10655 ( .A(n10269), .B(n10268), .Z(n10300) );
  NAND U10656 ( .A(y[739]), .B(x[143]), .Z(n10165) );
  XNOR U10657 ( .A(n10166), .B(n10165), .Z(n10260) );
  AND U10658 ( .A(x[142]), .B(y[740]), .Z(n10259) );
  XOR U10659 ( .A(n10260), .B(n10259), .Z(n10299) );
  XOR U10660 ( .A(n10300), .B(n10299), .Z(n10302) );
  XOR U10661 ( .A(n10301), .B(n10302), .Z(n10309) );
  NANDN U10662 ( .A(n10168), .B(n10167), .Z(n10172) );
  NANDN U10663 ( .A(n10170), .B(n10169), .Z(n10171) );
  AND U10664 ( .A(n10172), .B(n10171), .Z(n10322) );
  AND U10665 ( .A(y[743]), .B(x[139]), .Z(n10174) );
  NAND U10666 ( .A(y[738]), .B(x[144]), .Z(n10173) );
  XNOR U10667 ( .A(n10174), .B(n10173), .Z(n10258) );
  AND U10668 ( .A(x[130]), .B(y[752]), .Z(n10257) );
  XOR U10669 ( .A(n10258), .B(n10257), .Z(n10321) );
  AND U10670 ( .A(y[749]), .B(x[133]), .Z(n10383) );
  NAND U10671 ( .A(y[748]), .B(x[134]), .Z(n10175) );
  XNOR U10672 ( .A(n10383), .B(n10175), .Z(n10256) );
  AND U10673 ( .A(y[750]), .B(x[132]), .Z(n10177) );
  NAND U10674 ( .A(y[746]), .B(x[136]), .Z(n10176) );
  XNOR U10675 ( .A(n10177), .B(n10176), .Z(n10289) );
  AND U10676 ( .A(x[135]), .B(y[747]), .Z(n10288) );
  XOR U10677 ( .A(n10289), .B(n10288), .Z(n10255) );
  XOR U10678 ( .A(n10256), .B(n10255), .Z(n10323) );
  XOR U10679 ( .A(n10324), .B(n10323), .Z(n10311) );
  XOR U10680 ( .A(n10312), .B(n10311), .Z(n10245) );
  NANDN U10681 ( .A(n10183), .B(n10182), .Z(n10187) );
  NANDN U10682 ( .A(n10185), .B(n10184), .Z(n10186) );
  NAND U10683 ( .A(n10187), .B(n10186), .Z(n10304) );
  NANDN U10684 ( .A(n10189), .B(n10188), .Z(n10193) );
  NAND U10685 ( .A(n10191), .B(n10190), .Z(n10192) );
  NAND U10686 ( .A(n10193), .B(n10192), .Z(n10306) );
  XNOR U10687 ( .A(n10245), .B(n10244), .Z(n10247) );
  AND U10688 ( .A(x[136]), .B(y[748]), .Z(n10501) );
  NAND U10689 ( .A(n10501), .B(n10194), .Z(n10198) );
  NANDN U10690 ( .A(n10196), .B(n10195), .Z(n10197) );
  AND U10691 ( .A(n10198), .B(n10197), .Z(n10316) );
  NAND U10692 ( .A(x[137]), .B(y[752]), .Z(n11139) );
  NAND U10693 ( .A(x[138]), .B(y[751]), .Z(n11138) );
  NANDN U10694 ( .A(n11138), .B(n10201), .Z(n10205) );
  NANDN U10695 ( .A(n10203), .B(n10202), .Z(n10204) );
  NAND U10696 ( .A(n10205), .B(n10204), .Z(n10297) );
  AND U10697 ( .A(x[128]), .B(y[754]), .Z(n10270) );
  NAND U10698 ( .A(x[146]), .B(y[736]), .Z(n10271) );
  XNOR U10699 ( .A(n10270), .B(n10271), .Z(n10272) );
  NAND U10700 ( .A(x[145]), .B(y[737]), .Z(n10292) );
  XOR U10701 ( .A(o[114]), .B(n10292), .Z(n10273) );
  XNOR U10702 ( .A(n10272), .B(n10273), .Z(n10296) );
  AND U10703 ( .A(y[751]), .B(x[131]), .Z(n10207) );
  NAND U10704 ( .A(y[741]), .B(x[141]), .Z(n10206) );
  XNOR U10705 ( .A(n10207), .B(n10206), .Z(n10280) );
  AND U10706 ( .A(x[140]), .B(y[742]), .Z(n10279) );
  XOR U10707 ( .A(n10280), .B(n10279), .Z(n10295) );
  XOR U10708 ( .A(n10296), .B(n10295), .Z(n10298) );
  XOR U10709 ( .A(n10297), .B(n10298), .Z(n10317) );
  XOR U10710 ( .A(n10318), .B(n10317), .Z(n10249) );
  XNOR U10711 ( .A(n10249), .B(n10248), .Z(n10251) );
  NANDN U10712 ( .A(n10213), .B(n10212), .Z(n10217) );
  NANDN U10713 ( .A(n10215), .B(n10214), .Z(n10216) );
  AND U10714 ( .A(n10217), .B(n10216), .Z(n10250) );
  XOR U10715 ( .A(n10251), .B(n10250), .Z(n10246) );
  XOR U10716 ( .A(n10247), .B(n10246), .Z(n10242) );
  XNOR U10717 ( .A(n10240), .B(n10241), .Z(n10243) );
  XOR U10718 ( .A(n10242), .B(n10243), .Z(n10330) );
  XOR U10719 ( .A(n10331), .B(n10330), .Z(n10332) );
  XNOR U10720 ( .A(n10333), .B(n10332), .Z(n10329) );
  NAND U10721 ( .A(n10227), .B(n10226), .Z(n10231) );
  NANDN U10722 ( .A(n10229), .B(n10228), .Z(n10230) );
  NAND U10723 ( .A(n10231), .B(n10230), .Z(n10328) );
  NANDN U10724 ( .A(n10232), .B(n10233), .Z(n10238) );
  NOR U10725 ( .A(n10234), .B(n10233), .Z(n10236) );
  OR U10726 ( .A(n10236), .B(n10235), .Z(n10237) );
  AND U10727 ( .A(n10238), .B(n10237), .Z(n10327) );
  XOR U10728 ( .A(n10328), .B(n10327), .Z(n10239) );
  XNOR U10729 ( .A(n10329), .B(n10239), .Z(N243) );
  NANDN U10730 ( .A(n10249), .B(n10248), .Z(n10253) );
  NAND U10731 ( .A(n10251), .B(n10250), .Z(n10252) );
  NAND U10732 ( .A(n10253), .B(n10252), .Z(n10426) );
  AND U10733 ( .A(x[143]), .B(y[745]), .Z(n11022) );
  NAND U10734 ( .A(n11022), .B(n10349), .Z(n10262) );
  NAND U10735 ( .A(n10260), .B(n10259), .Z(n10261) );
  AND U10736 ( .A(n10262), .B(n10261), .Z(n10340) );
  AND U10737 ( .A(y[754]), .B(x[129]), .Z(n10264) );
  NAND U10738 ( .A(y[747]), .B(x[136]), .Z(n10263) );
  XNOR U10739 ( .A(n10264), .B(n10263), .Z(n10400) );
  AND U10740 ( .A(y[753]), .B(x[130]), .Z(n10266) );
  NAND U10741 ( .A(y[742]), .B(x[141]), .Z(n10265) );
  XNOR U10742 ( .A(n10266), .B(n10265), .Z(n10355) );
  XOR U10743 ( .A(n10338), .B(n10337), .Z(n10339) );
  XNOR U10744 ( .A(n10340), .B(n10339), .Z(n10420) );
  XOR U10745 ( .A(n10419), .B(n10420), .Z(n10422) );
  XOR U10746 ( .A(n10421), .B(n10422), .Z(n10424) );
  AND U10747 ( .A(x[138]), .B(y[753]), .Z(n11445) );
  IV U10748 ( .A(n11445), .Z(n11349) );
  NANDN U10749 ( .A(n10271), .B(n10270), .Z(n10275) );
  NANDN U10750 ( .A(n10273), .B(n10272), .Z(n10274) );
  AND U10751 ( .A(n10275), .B(n10274), .Z(n10378) );
  AND U10752 ( .A(y[746]), .B(x[137]), .Z(n10277) );
  NAND U10753 ( .A(y[739]), .B(x[144]), .Z(n10276) );
  XNOR U10754 ( .A(n10277), .B(n10276), .Z(n10350) );
  NAND U10755 ( .A(x[143]), .B(y[740]), .Z(n10351) );
  XNOR U10756 ( .A(n10378), .B(n10377), .Z(n10379) );
  XNOR U10757 ( .A(n10380), .B(n10379), .Z(n10416) );
  AND U10758 ( .A(x[141]), .B(y[751]), .Z(n11671) );
  NANDN U10759 ( .A(n10278), .B(n11671), .Z(n10282) );
  NAND U10760 ( .A(n10280), .B(n10279), .Z(n10281) );
  AND U10761 ( .A(n10282), .B(n10281), .Z(n10374) );
  AND U10762 ( .A(y[738]), .B(x[145]), .Z(n10284) );
  NAND U10763 ( .A(y[745]), .B(x[138]), .Z(n10283) );
  XNOR U10764 ( .A(n10284), .B(n10283), .Z(n10406) );
  NAND U10765 ( .A(x[146]), .B(y[737]), .Z(n10370) );
  XNOR U10766 ( .A(o[115]), .B(n10370), .Z(n10405) );
  XOR U10767 ( .A(n10406), .B(n10405), .Z(n10372) );
  AND U10768 ( .A(y[752]), .B(x[131]), .Z(n10286) );
  NAND U10769 ( .A(y[744]), .B(x[139]), .Z(n10285) );
  XNOR U10770 ( .A(n10286), .B(n10285), .Z(n10364) );
  XOR U10771 ( .A(n10372), .B(n10371), .Z(n10373) );
  XNOR U10772 ( .A(n10374), .B(n10373), .Z(n10414) );
  NAND U10773 ( .A(n10659), .B(n10287), .Z(n10291) );
  NAND U10774 ( .A(n10289), .B(n10288), .Z(n10290) );
  AND U10775 ( .A(n10291), .B(n10290), .Z(n10346) );
  AND U10776 ( .A(x[128]), .B(y[755]), .Z(n10387) );
  NAND U10777 ( .A(x[147]), .B(y[736]), .Z(n10388) );
  XNOR U10778 ( .A(n10387), .B(n10388), .Z(n10390) );
  ANDN U10779 ( .B(o[114]), .A(n10292), .Z(n10389) );
  XOR U10780 ( .A(n10390), .B(n10389), .Z(n10344) );
  AND U10781 ( .A(x[132]), .B(y[751]), .Z(n10515) );
  AND U10782 ( .A(y[750]), .B(x[133]), .Z(n10294) );
  NAND U10783 ( .A(y[749]), .B(x[134]), .Z(n10293) );
  XOR U10784 ( .A(n10294), .B(n10293), .Z(n10384) );
  XNOR U10785 ( .A(n10515), .B(n10384), .Z(n10343) );
  XOR U10786 ( .A(n10344), .B(n10343), .Z(n10345) );
  XOR U10787 ( .A(n10346), .B(n10345), .Z(n10413) );
  XNOR U10788 ( .A(n10414), .B(n10413), .Z(n10415) );
  XOR U10789 ( .A(n10416), .B(n10415), .Z(n10411) );
  XOR U10790 ( .A(n10409), .B(n10410), .Z(n10412) );
  XOR U10791 ( .A(n10411), .B(n10412), .Z(n10423) );
  XOR U10792 ( .A(n10424), .B(n10423), .Z(n10425) );
  XNOR U10793 ( .A(n10426), .B(n10425), .Z(n10435) );
  NANDN U10794 ( .A(n10304), .B(n10303), .Z(n10308) );
  NANDN U10795 ( .A(n10306), .B(n10305), .Z(n10307) );
  AND U10796 ( .A(n10308), .B(n10307), .Z(n10434) );
  NANDN U10797 ( .A(n10310), .B(n10309), .Z(n10314) );
  NAND U10798 ( .A(n10312), .B(n10311), .Z(n10313) );
  AND U10799 ( .A(n10314), .B(n10313), .Z(n10430) );
  NANDN U10800 ( .A(n10316), .B(n10315), .Z(n10320) );
  NAND U10801 ( .A(n10318), .B(n10317), .Z(n10319) );
  AND U10802 ( .A(n10320), .B(n10319), .Z(n10428) );
  NANDN U10803 ( .A(n10322), .B(n10321), .Z(n10326) );
  NAND U10804 ( .A(n10324), .B(n10323), .Z(n10325) );
  NAND U10805 ( .A(n10326), .B(n10325), .Z(n10427) );
  XOR U10806 ( .A(n10434), .B(n10433), .Z(n10436) );
  XOR U10807 ( .A(n10435), .B(n10436), .Z(n10442) );
  XNOR U10808 ( .A(n10443), .B(n10442), .Z(n10445) );
  XOR U10809 ( .A(n10444), .B(n10445), .Z(n10441) );
  NAND U10810 ( .A(n10331), .B(n10330), .Z(n10335) );
  NAND U10811 ( .A(n10333), .B(n10332), .Z(n10334) );
  NAND U10812 ( .A(n10335), .B(n10334), .Z(n10439) );
  XNOR U10813 ( .A(n10440), .B(n10439), .Z(n10336) );
  XNOR U10814 ( .A(n10441), .B(n10336), .Z(N244) );
  NAND U10815 ( .A(n10338), .B(n10337), .Z(n10342) );
  NANDN U10816 ( .A(n10340), .B(n10339), .Z(n10341) );
  AND U10817 ( .A(n10342), .B(n10341), .Z(n10450) );
  NAND U10818 ( .A(n10344), .B(n10343), .Z(n10348) );
  NANDN U10819 ( .A(n10346), .B(n10345), .Z(n10347) );
  NAND U10820 ( .A(n10348), .B(n10347), .Z(n10449) );
  XNOR U10821 ( .A(n10450), .B(n10449), .Z(n10452) );
  AND U10822 ( .A(x[144]), .B(y[746]), .Z(n11307) );
  NAND U10823 ( .A(n11307), .B(n10349), .Z(n10353) );
  NANDN U10824 ( .A(n10351), .B(n10350), .Z(n10352) );
  AND U10825 ( .A(n10353), .B(n10352), .Z(n10490) );
  AND U10826 ( .A(x[141]), .B(y[753]), .Z(n11924) );
  NAND U10827 ( .A(n11924), .B(n10354), .Z(n10358) );
  NANDN U10828 ( .A(n10356), .B(n10355), .Z(n10357) );
  AND U10829 ( .A(n10358), .B(n10357), .Z(n10535) );
  NAND U10830 ( .A(y[740]), .B(x[144]), .Z(n10359) );
  XNOR U10831 ( .A(n10360), .B(n10359), .Z(n10496) );
  NAND U10832 ( .A(x[130]), .B(y[754]), .Z(n10497) );
  XNOR U10833 ( .A(n10496), .B(n10497), .Z(n10533) );
  NAND U10834 ( .A(y[741]), .B(x[143]), .Z(n10361) );
  XNOR U10835 ( .A(n10362), .B(n10361), .Z(n10466) );
  NAND U10836 ( .A(x[142]), .B(y[742]), .Z(n10467) );
  XNOR U10837 ( .A(n10466), .B(n10467), .Z(n10532) );
  XOR U10838 ( .A(n10533), .B(n10532), .Z(n10534) );
  NAND U10839 ( .A(x[139]), .B(y[752]), .Z(n11446) );
  NANDN U10840 ( .A(n11446), .B(n10363), .Z(n10367) );
  NANDN U10841 ( .A(n10365), .B(n10364), .Z(n10366) );
  AND U10842 ( .A(n10367), .B(n10366), .Z(n10541) );
  AND U10843 ( .A(y[755]), .B(x[129]), .Z(n10369) );
  NAND U10844 ( .A(y[745]), .B(x[139]), .Z(n10368) );
  XNOR U10845 ( .A(n10369), .B(n10368), .Z(n10462) );
  NAND U10846 ( .A(x[147]), .B(y[737]), .Z(n10470) );
  XNOR U10847 ( .A(o[116]), .B(n10470), .Z(n10461) );
  XOR U10848 ( .A(n10462), .B(n10461), .Z(n10539) );
  AND U10849 ( .A(x[128]), .B(y[756]), .Z(n10520) );
  NAND U10850 ( .A(x[148]), .B(y[736]), .Z(n10521) );
  XNOR U10851 ( .A(n10520), .B(n10521), .Z(n10523) );
  ANDN U10852 ( .B(o[115]), .A(n10370), .Z(n10522) );
  XOR U10853 ( .A(n10523), .B(n10522), .Z(n10538) );
  XOR U10854 ( .A(n10539), .B(n10538), .Z(n10540) );
  XOR U10855 ( .A(n10492), .B(n10491), .Z(n10451) );
  XOR U10856 ( .A(n10452), .B(n10451), .Z(n10547) );
  NAND U10857 ( .A(n10372), .B(n10371), .Z(n10376) );
  NANDN U10858 ( .A(n10374), .B(n10373), .Z(n10375) );
  AND U10859 ( .A(n10376), .B(n10375), .Z(n10545) );
  NANDN U10860 ( .A(n10378), .B(n10377), .Z(n10382) );
  NANDN U10861 ( .A(n10380), .B(n10379), .Z(n10381) );
  AND U10862 ( .A(n10382), .B(n10381), .Z(n10486) );
  AND U10863 ( .A(x[134]), .B(y[750]), .Z(n10472) );
  NAND U10864 ( .A(n10472), .B(n10383), .Z(n10386) );
  NANDN U10865 ( .A(n10384), .B(n10515), .Z(n10385) );
  AND U10866 ( .A(n10386), .B(n10385), .Z(n10480) );
  NANDN U10867 ( .A(n10388), .B(n10387), .Z(n10392) );
  NAND U10868 ( .A(n10390), .B(n10389), .Z(n10391) );
  AND U10869 ( .A(n10392), .B(n10391), .Z(n10478) );
  AND U10870 ( .A(y[738]), .B(x[146]), .Z(n10394) );
  NAND U10871 ( .A(y[744]), .B(x[140]), .Z(n10393) );
  XNOR U10872 ( .A(n10394), .B(n10393), .Z(n10456) );
  NAND U10873 ( .A(x[145]), .B(y[739]), .Z(n10457) );
  XNOR U10874 ( .A(n10456), .B(n10457), .Z(n10477) );
  XNOR U10875 ( .A(n10478), .B(n10477), .Z(n10479) );
  XOR U10876 ( .A(n10480), .B(n10479), .Z(n10484) );
  AND U10877 ( .A(y[753]), .B(x[131]), .Z(n10396) );
  NAND U10878 ( .A(y[743]), .B(x[141]), .Z(n10395) );
  XNOR U10879 ( .A(n10396), .B(n10395), .Z(n10502) );
  XOR U10880 ( .A(n10502), .B(n10501), .Z(n10474) );
  AND U10881 ( .A(y[751]), .B(x[133]), .Z(n10398) );
  NAND U10882 ( .A(y[752]), .B(x[132]), .Z(n10397) );
  XNOR U10883 ( .A(n10398), .B(n10397), .Z(n10517) );
  AND U10884 ( .A(x[135]), .B(y[749]), .Z(n10516) );
  XNOR U10885 ( .A(n10517), .B(n10516), .Z(n10471) );
  XNOR U10886 ( .A(n10472), .B(n10471), .Z(n10473) );
  XOR U10887 ( .A(n10474), .B(n10473), .Z(n10528) );
  AND U10888 ( .A(x[136]), .B(y[754]), .Z(n11623) );
  NAND U10889 ( .A(n11623), .B(n10399), .Z(n10403) );
  NANDN U10890 ( .A(n10401), .B(n10400), .Z(n10402) );
  AND U10891 ( .A(n10403), .B(n10402), .Z(n10527) );
  AND U10892 ( .A(x[145]), .B(y[745]), .Z(n11314) );
  AND U10893 ( .A(x[138]), .B(y[738]), .Z(n10404) );
  NAND U10894 ( .A(n11314), .B(n10404), .Z(n10408) );
  NAND U10895 ( .A(n10406), .B(n10405), .Z(n10407) );
  NAND U10896 ( .A(n10408), .B(n10407), .Z(n10526) );
  XNOR U10897 ( .A(n10528), .B(n10529), .Z(n10483) );
  XOR U10898 ( .A(n10484), .B(n10483), .Z(n10485) );
  XOR U10899 ( .A(n10486), .B(n10485), .Z(n10544) );
  XOR U10900 ( .A(n10545), .B(n10544), .Z(n10546) );
  XNOR U10901 ( .A(n10547), .B(n10546), .Z(n10551) );
  NANDN U10902 ( .A(n10414), .B(n10413), .Z(n10418) );
  NANDN U10903 ( .A(n10416), .B(n10415), .Z(n10417) );
  NAND U10904 ( .A(n10418), .B(n10417), .Z(n10557) );
  XOR U10905 ( .A(n10557), .B(n10556), .Z(n10558) );
  XNOR U10906 ( .A(n10559), .B(n10558), .Z(n10550) );
  XNOR U10907 ( .A(n10551), .B(n10550), .Z(n10553) );
  XOR U10908 ( .A(n10553), .B(n10552), .Z(n10565) );
  NANDN U10909 ( .A(n10428), .B(n10427), .Z(n10432) );
  NANDN U10910 ( .A(n10430), .B(n10429), .Z(n10431) );
  AND U10911 ( .A(n10432), .B(n10431), .Z(n10562) );
  NAND U10912 ( .A(n10434), .B(n10433), .Z(n10438) );
  NAND U10913 ( .A(n10436), .B(n10435), .Z(n10437) );
  NAND U10914 ( .A(n10438), .B(n10437), .Z(n10563) );
  XOR U10915 ( .A(n10565), .B(n10564), .Z(n10571) );
  NAND U10916 ( .A(n10443), .B(n10442), .Z(n10447) );
  NANDN U10917 ( .A(n10445), .B(n10444), .Z(n10446) );
  AND U10918 ( .A(n10447), .B(n10446), .Z(n10570) );
  IV U10919 ( .A(n10570), .Z(n10568) );
  XOR U10920 ( .A(n10569), .B(n10568), .Z(n10448) );
  XNOR U10921 ( .A(n10571), .B(n10448), .Z(N245) );
  NANDN U10922 ( .A(n10450), .B(n10449), .Z(n10454) );
  NAND U10923 ( .A(n10452), .B(n10451), .Z(n10453) );
  AND U10924 ( .A(n10454), .B(n10453), .Z(n10582) );
  AND U10925 ( .A(x[146]), .B(y[744]), .Z(n11316) );
  NAND U10926 ( .A(n11316), .B(n10455), .Z(n10459) );
  NANDN U10927 ( .A(n10457), .B(n10456), .Z(n10458) );
  AND U10928 ( .A(n10459), .B(n10458), .Z(n10592) );
  AND U10929 ( .A(x[139]), .B(y[755]), .Z(n11997) );
  NAND U10930 ( .A(n11997), .B(n10460), .Z(n10464) );
  NAND U10931 ( .A(n10462), .B(n10461), .Z(n10463) );
  NAND U10932 ( .A(n10464), .B(n10463), .Z(n10591) );
  XNOR U10933 ( .A(n10592), .B(n10591), .Z(n10594) );
  AND U10934 ( .A(x[143]), .B(y[747]), .Z(n11302) );
  NAND U10935 ( .A(n11302), .B(n10465), .Z(n10469) );
  NANDN U10936 ( .A(n10467), .B(n10466), .Z(n10468) );
  NAND U10937 ( .A(n10469), .B(n10468), .Z(n10623) );
  AND U10938 ( .A(x[128]), .B(y[757]), .Z(n10644) );
  NAND U10939 ( .A(x[149]), .B(y[736]), .Z(n10645) );
  XNOR U10940 ( .A(n10644), .B(n10645), .Z(n10647) );
  ANDN U10941 ( .B(o[116]), .A(n10470), .Z(n10646) );
  XOR U10942 ( .A(n10647), .B(n10646), .Z(n10622) );
  AND U10943 ( .A(x[133]), .B(y[752]), .Z(n10628) );
  AND U10944 ( .A(x[144]), .B(y[741]), .Z(n10627) );
  XOR U10945 ( .A(n10628), .B(n10627), .Z(n10630) );
  AND U10946 ( .A(x[143]), .B(y[742]), .Z(n10629) );
  XOR U10947 ( .A(n10630), .B(n10629), .Z(n10621) );
  XOR U10948 ( .A(n10622), .B(n10621), .Z(n10624) );
  XOR U10949 ( .A(n10623), .B(n10624), .Z(n10593) );
  XOR U10950 ( .A(n10594), .B(n10593), .Z(n10586) );
  NANDN U10951 ( .A(n10472), .B(n10471), .Z(n10476) );
  NANDN U10952 ( .A(n10474), .B(n10473), .Z(n10475) );
  NAND U10953 ( .A(n10476), .B(n10475), .Z(n10585) );
  NANDN U10954 ( .A(n10478), .B(n10477), .Z(n10482) );
  NANDN U10955 ( .A(n10480), .B(n10479), .Z(n10481) );
  AND U10956 ( .A(n10482), .B(n10481), .Z(n10587) );
  XOR U10957 ( .A(n10588), .B(n10587), .Z(n10580) );
  NAND U10958 ( .A(n10484), .B(n10483), .Z(n10488) );
  NAND U10959 ( .A(n10486), .B(n10485), .Z(n10487) );
  AND U10960 ( .A(n10488), .B(n10487), .Z(n10579) );
  XNOR U10961 ( .A(n10580), .B(n10579), .Z(n10581) );
  XOR U10962 ( .A(n10582), .B(n10581), .Z(n10575) );
  NANDN U10963 ( .A(n10490), .B(n10489), .Z(n10494) );
  NAND U10964 ( .A(n10492), .B(n10491), .Z(n10493) );
  AND U10965 ( .A(n10494), .B(n10493), .Z(n10680) );
  NAND U10966 ( .A(n11307), .B(n10495), .Z(n10499) );
  NANDN U10967 ( .A(n10497), .B(n10496), .Z(n10498) );
  AND U10968 ( .A(n10499), .B(n10498), .Z(n10610) );
  AND U10969 ( .A(x[131]), .B(y[743]), .Z(n10500) );
  NAND U10970 ( .A(n11924), .B(n10500), .Z(n10504) );
  NAND U10971 ( .A(n10502), .B(n10501), .Z(n10503) );
  AND U10972 ( .A(n10504), .B(n10503), .Z(n10606) );
  AND U10973 ( .A(y[738]), .B(x[147]), .Z(n10506) );
  NAND U10974 ( .A(y[746]), .B(x[139]), .Z(n10505) );
  XNOR U10975 ( .A(n10506), .B(n10505), .Z(n10662) );
  AND U10976 ( .A(x[148]), .B(y[737]), .Z(n10643) );
  XOR U10977 ( .A(n10643), .B(o[117]), .Z(n10661) );
  XOR U10978 ( .A(n10662), .B(n10661), .Z(n10604) );
  AND U10979 ( .A(y[739]), .B(x[146]), .Z(n10508) );
  NAND U10980 ( .A(y[747]), .B(x[138]), .Z(n10507) );
  XNOR U10981 ( .A(n10508), .B(n10507), .Z(n10651) );
  NAND U10982 ( .A(x[129]), .B(y[756]), .Z(n10652) );
  XNOR U10983 ( .A(n10651), .B(n10652), .Z(n10603) );
  XOR U10984 ( .A(n10604), .B(n10603), .Z(n10605) );
  XNOR U10985 ( .A(n10606), .B(n10605), .Z(n10609) );
  XNOR U10986 ( .A(n10610), .B(n10609), .Z(n10612) );
  AND U10987 ( .A(x[135]), .B(y[750]), .Z(n10909) );
  AND U10988 ( .A(y[743]), .B(x[142]), .Z(n10510) );
  NAND U10989 ( .A(y[751]), .B(x[134]), .Z(n10509) );
  XOR U10990 ( .A(n10510), .B(n10509), .Z(n10655) );
  XNOR U10991 ( .A(n10909), .B(n10655), .Z(n10674) );
  NAND U10992 ( .A(x[137]), .B(y[748]), .Z(n10672) );
  NAND U10993 ( .A(x[136]), .B(y[749]), .Z(n10671) );
  XOR U10994 ( .A(n10672), .B(n10671), .Z(n10673) );
  AND U10995 ( .A(y[740]), .B(x[145]), .Z(n10512) );
  NAND U10996 ( .A(y[745]), .B(x[140]), .Z(n10511) );
  XNOR U10997 ( .A(n10512), .B(n10511), .Z(n10665) );
  NAND U10998 ( .A(x[130]), .B(y[755]), .Z(n10666) );
  XNOR U10999 ( .A(n10665), .B(n10666), .Z(n10616) );
  AND U11000 ( .A(y[754]), .B(x[131]), .Z(n10514) );
  NAND U11001 ( .A(y[744]), .B(x[141]), .Z(n10513) );
  XNOR U11002 ( .A(n10514), .B(n10513), .Z(n10640) );
  AND U11003 ( .A(x[132]), .B(y[753]), .Z(n10639) );
  XOR U11004 ( .A(n10640), .B(n10639), .Z(n10615) );
  XOR U11005 ( .A(n10616), .B(n10615), .Z(n10617) );
  NAND U11006 ( .A(n10628), .B(n10515), .Z(n10519) );
  NAND U11007 ( .A(n10517), .B(n10516), .Z(n10518) );
  AND U11008 ( .A(n10519), .B(n10518), .Z(n10598) );
  NANDN U11009 ( .A(n10521), .B(n10520), .Z(n10525) );
  NAND U11010 ( .A(n10523), .B(n10522), .Z(n10524) );
  NAND U11011 ( .A(n10525), .B(n10524), .Z(n10597) );
  XNOR U11012 ( .A(n10598), .B(n10597), .Z(n10599) );
  XOR U11013 ( .A(n10600), .B(n10599), .Z(n10611) );
  XOR U11014 ( .A(n10612), .B(n10611), .Z(n10678) );
  NANDN U11015 ( .A(n10527), .B(n10526), .Z(n10531) );
  NAND U11016 ( .A(n10529), .B(n10528), .Z(n10530) );
  NAND U11017 ( .A(n10531), .B(n10530), .Z(n10685) );
  NAND U11018 ( .A(n10533), .B(n10532), .Z(n10537) );
  NANDN U11019 ( .A(n10535), .B(n10534), .Z(n10536) );
  NAND U11020 ( .A(n10537), .B(n10536), .Z(n10684) );
  NAND U11021 ( .A(n10539), .B(n10538), .Z(n10543) );
  NANDN U11022 ( .A(n10541), .B(n10540), .Z(n10542) );
  NAND U11023 ( .A(n10543), .B(n10542), .Z(n10683) );
  XOR U11024 ( .A(n10684), .B(n10683), .Z(n10686) );
  XOR U11025 ( .A(n10685), .B(n10686), .Z(n10677) );
  XOR U11026 ( .A(n10678), .B(n10677), .Z(n10679) );
  XOR U11027 ( .A(n10680), .B(n10679), .Z(n10574) );
  NAND U11028 ( .A(n10545), .B(n10544), .Z(n10549) );
  NANDN U11029 ( .A(n10547), .B(n10546), .Z(n10548) );
  NAND U11030 ( .A(n10549), .B(n10548), .Z(n10573) );
  XOR U11031 ( .A(n10574), .B(n10573), .Z(n10576) );
  XOR U11032 ( .A(n10575), .B(n10576), .Z(n10692) );
  NANDN U11033 ( .A(n10551), .B(n10550), .Z(n10555) );
  NAND U11034 ( .A(n10553), .B(n10552), .Z(n10554) );
  NAND U11035 ( .A(n10555), .B(n10554), .Z(n10689) );
  NAND U11036 ( .A(n10557), .B(n10556), .Z(n10561) );
  NAND U11037 ( .A(n10559), .B(n10558), .Z(n10560) );
  AND U11038 ( .A(n10561), .B(n10560), .Z(n10690) );
  XOR U11039 ( .A(n10689), .B(n10690), .Z(n10691) );
  XNOR U11040 ( .A(n10692), .B(n10691), .Z(n10695) );
  NANDN U11041 ( .A(n10563), .B(n10562), .Z(n10567) );
  NANDN U11042 ( .A(n10565), .B(n10564), .Z(n10566) );
  NAND U11043 ( .A(n10567), .B(n10566), .Z(n10693) );
  XOR U11044 ( .A(n10693), .B(n10694), .Z(n10572) );
  XNOR U11045 ( .A(n10695), .B(n10572), .Z(N246) );
  NAND U11046 ( .A(n10574), .B(n10573), .Z(n10578) );
  NAND U11047 ( .A(n10576), .B(n10575), .Z(n10577) );
  AND U11048 ( .A(n10578), .B(n10577), .Z(n10826) );
  NANDN U11049 ( .A(n10580), .B(n10579), .Z(n10584) );
  NANDN U11050 ( .A(n10582), .B(n10581), .Z(n10583) );
  AND U11051 ( .A(n10584), .B(n10583), .Z(n10824) );
  NANDN U11052 ( .A(n10586), .B(n10585), .Z(n10590) );
  NAND U11053 ( .A(n10588), .B(n10587), .Z(n10589) );
  AND U11054 ( .A(n10590), .B(n10589), .Z(n10704) );
  NANDN U11055 ( .A(n10592), .B(n10591), .Z(n10596) );
  NAND U11056 ( .A(n10594), .B(n10593), .Z(n10595) );
  AND U11057 ( .A(n10596), .B(n10595), .Z(n10712) );
  NANDN U11058 ( .A(n10598), .B(n10597), .Z(n10602) );
  NAND U11059 ( .A(n10600), .B(n10599), .Z(n10601) );
  AND U11060 ( .A(n10602), .B(n10601), .Z(n10710) );
  NAND U11061 ( .A(n10604), .B(n10603), .Z(n10608) );
  NANDN U11062 ( .A(n10606), .B(n10605), .Z(n10607) );
  NAND U11063 ( .A(n10608), .B(n10607), .Z(n10709) );
  XNOR U11064 ( .A(n10710), .B(n10709), .Z(n10711) );
  XOR U11065 ( .A(n10712), .B(n10711), .Z(n10703) );
  NANDN U11066 ( .A(n10610), .B(n10609), .Z(n10614) );
  NAND U11067 ( .A(n10612), .B(n10611), .Z(n10613) );
  AND U11068 ( .A(n10614), .B(n10613), .Z(n10813) );
  NAND U11069 ( .A(n10616), .B(n10615), .Z(n10620) );
  NANDN U11070 ( .A(n10618), .B(n10617), .Z(n10619) );
  AND U11071 ( .A(n10620), .B(n10619), .Z(n10793) );
  NAND U11072 ( .A(n10622), .B(n10621), .Z(n10626) );
  NAND U11073 ( .A(n10624), .B(n10623), .Z(n10625) );
  NAND U11074 ( .A(n10626), .B(n10625), .Z(n10792) );
  XNOR U11075 ( .A(n10793), .B(n10792), .Z(n10795) );
  NAND U11076 ( .A(n10628), .B(n10627), .Z(n10632) );
  AND U11077 ( .A(n10630), .B(n10629), .Z(n10631) );
  ANDN U11078 ( .B(n10632), .A(n10631), .Z(n10756) );
  AND U11079 ( .A(y[738]), .B(x[148]), .Z(n10634) );
  NAND U11080 ( .A(y[745]), .B(x[141]), .Z(n10633) );
  XNOR U11081 ( .A(n10634), .B(n10633), .Z(n10777) );
  AND U11082 ( .A(x[130]), .B(y[756]), .Z(n10776) );
  XOR U11083 ( .A(n10777), .B(n10776), .Z(n10754) );
  AND U11084 ( .A(y[752]), .B(x[134]), .Z(n10636) );
  NAND U11085 ( .A(y[743]), .B(x[143]), .Z(n10635) );
  XNOR U11086 ( .A(n10636), .B(n10635), .Z(n10788) );
  XOR U11087 ( .A(n10788), .B(n10637), .Z(n10753) );
  XOR U11088 ( .A(n10754), .B(n10753), .Z(n10755) );
  XNOR U11089 ( .A(n10756), .B(n10755), .Z(n10799) );
  AND U11090 ( .A(x[141]), .B(y[754]), .Z(n12100) );
  NANDN U11091 ( .A(n10638), .B(n12100), .Z(n10642) );
  NAND U11092 ( .A(n10640), .B(n10639), .Z(n10641) );
  AND U11093 ( .A(n10642), .B(n10641), .Z(n10724) );
  AND U11094 ( .A(x[129]), .B(y[757]), .Z(n10747) );
  XOR U11095 ( .A(n10748), .B(n10747), .Z(n10746) );
  AND U11096 ( .A(n10643), .B(o[117]), .Z(n10745) );
  XOR U11097 ( .A(n10746), .B(n10745), .Z(n10722) );
  AND U11098 ( .A(x[142]), .B(y[744]), .Z(n10740) );
  AND U11099 ( .A(x[131]), .B(y[755]), .Z(n10739) );
  XOR U11100 ( .A(n10740), .B(n10739), .Z(n10742) );
  AND U11101 ( .A(x[147]), .B(y[739]), .Z(n10741) );
  XOR U11102 ( .A(n10742), .B(n10741), .Z(n10721) );
  XOR U11103 ( .A(n10722), .B(n10721), .Z(n10723) );
  XNOR U11104 ( .A(n10724), .B(n10723), .Z(n10798) );
  XOR U11105 ( .A(n10799), .B(n10798), .Z(n10801) );
  NANDN U11106 ( .A(n10645), .B(n10644), .Z(n10649) );
  NAND U11107 ( .A(n10647), .B(n10646), .Z(n10648) );
  AND U11108 ( .A(n10649), .B(n10648), .Z(n10716) );
  AND U11109 ( .A(x[146]), .B(y[747]), .Z(n11824) );
  NAND U11110 ( .A(n11824), .B(n10650), .Z(n10654) );
  NANDN U11111 ( .A(n10652), .B(n10651), .Z(n10653) );
  NAND U11112 ( .A(n10654), .B(n10653), .Z(n10715) );
  XNOR U11113 ( .A(n10716), .B(n10715), .Z(n10718) );
  AND U11114 ( .A(x[142]), .B(y[751]), .Z(n11858) );
  NAND U11115 ( .A(n11858), .B(n10787), .Z(n10657) );
  NANDN U11116 ( .A(n10655), .B(n10909), .Z(n10656) );
  NAND U11117 ( .A(n10657), .B(n10656), .Z(n10729) );
  AND U11118 ( .A(x[128]), .B(y[758]), .Z(n10765) );
  AND U11119 ( .A(x[150]), .B(y[736]), .Z(n10764) );
  XOR U11120 ( .A(n10765), .B(n10764), .Z(n10767) );
  AND U11121 ( .A(x[149]), .B(y[737]), .Z(n10786) );
  XOR U11122 ( .A(n10786), .B(o[118]), .Z(n10766) );
  XOR U11123 ( .A(n10767), .B(n10766), .Z(n10728) );
  NAND U11124 ( .A(y[751]), .B(x[135]), .Z(n10658) );
  XNOR U11125 ( .A(n10659), .B(n10658), .Z(n10771) );
  XOR U11126 ( .A(n10771), .B(n10770), .Z(n10727) );
  XOR U11127 ( .A(n10728), .B(n10727), .Z(n10730) );
  XOR U11128 ( .A(n10729), .B(n10730), .Z(n10717) );
  XOR U11129 ( .A(n10718), .B(n10717), .Z(n10800) );
  XOR U11130 ( .A(n10801), .B(n10800), .Z(n10794) );
  XOR U11131 ( .A(n10795), .B(n10794), .Z(n10811) );
  AND U11132 ( .A(x[147]), .B(y[746]), .Z(n11821) );
  NAND U11133 ( .A(n11821), .B(n10660), .Z(n10664) );
  NAND U11134 ( .A(n10662), .B(n10661), .Z(n10663) );
  AND U11135 ( .A(n10664), .B(n10663), .Z(n10805) );
  NAND U11136 ( .A(n11314), .B(n10759), .Z(n10668) );
  NANDN U11137 ( .A(n10666), .B(n10665), .Z(n10667) );
  AND U11138 ( .A(n10668), .B(n10667), .Z(n10736) );
  AND U11139 ( .A(x[133]), .B(y[753]), .Z(n10781) );
  AND U11140 ( .A(x[145]), .B(y[741]), .Z(n10780) );
  XOR U11141 ( .A(n10781), .B(n10780), .Z(n10783) );
  AND U11142 ( .A(x[144]), .B(y[742]), .Z(n10782) );
  XOR U11143 ( .A(n10783), .B(n10782), .Z(n10734) );
  AND U11144 ( .A(y[740]), .B(x[146]), .Z(n10670) );
  NAND U11145 ( .A(y[746]), .B(x[140]), .Z(n10669) );
  XNOR U11146 ( .A(n10670), .B(n10669), .Z(n10761) );
  AND U11147 ( .A(x[132]), .B(y[754]), .Z(n10760) );
  XOR U11148 ( .A(n10761), .B(n10760), .Z(n10733) );
  XOR U11149 ( .A(n10734), .B(n10733), .Z(n10735) );
  XNOR U11150 ( .A(n10736), .B(n10735), .Z(n10804) );
  XNOR U11151 ( .A(n10805), .B(n10804), .Z(n10807) );
  NAND U11152 ( .A(n10672), .B(n10671), .Z(n10676) );
  NANDN U11153 ( .A(n10674), .B(n10673), .Z(n10675) );
  AND U11154 ( .A(n10676), .B(n10675), .Z(n10806) );
  XNOR U11155 ( .A(n10807), .B(n10806), .Z(n10810) );
  XNOR U11156 ( .A(n10811), .B(n10810), .Z(n10812) );
  XOR U11157 ( .A(n10813), .B(n10812), .Z(n10705) );
  XOR U11158 ( .A(n10706), .B(n10705), .Z(n10700) );
  NAND U11159 ( .A(n10678), .B(n10677), .Z(n10682) );
  NANDN U11160 ( .A(n10680), .B(n10679), .Z(n10681) );
  AND U11161 ( .A(n10682), .B(n10681), .Z(n10698) );
  NAND U11162 ( .A(n10684), .B(n10683), .Z(n10688) );
  NAND U11163 ( .A(n10686), .B(n10685), .Z(n10687) );
  NAND U11164 ( .A(n10688), .B(n10687), .Z(n10697) );
  XNOR U11165 ( .A(n10824), .B(n10823), .Z(n10825) );
  XNOR U11166 ( .A(n10826), .B(n10825), .Z(n10817) );
  IV U11167 ( .A(n10819), .Z(n10816) );
  XOR U11168 ( .A(n10816), .B(n10820), .Z(n10696) );
  XNOR U11169 ( .A(n10817), .B(n10696), .Z(N247) );
  NANDN U11170 ( .A(n10698), .B(n10697), .Z(n10702) );
  NANDN U11171 ( .A(n10700), .B(n10699), .Z(n10701) );
  AND U11172 ( .A(n10702), .B(n10701), .Z(n10963) );
  NANDN U11173 ( .A(n10704), .B(n10703), .Z(n10708) );
  NAND U11174 ( .A(n10706), .B(n10705), .Z(n10707) );
  AND U11175 ( .A(n10708), .B(n10707), .Z(n10961) );
  NANDN U11176 ( .A(n10710), .B(n10709), .Z(n10714) );
  NANDN U11177 ( .A(n10712), .B(n10711), .Z(n10713) );
  AND U11178 ( .A(n10714), .B(n10713), .Z(n10945) );
  NANDN U11179 ( .A(n10716), .B(n10715), .Z(n10720) );
  NAND U11180 ( .A(n10718), .B(n10717), .Z(n10719) );
  NAND U11181 ( .A(n10720), .B(n10719), .Z(n10892) );
  NAND U11182 ( .A(n10722), .B(n10721), .Z(n10726) );
  NANDN U11183 ( .A(n10724), .B(n10723), .Z(n10725) );
  NAND U11184 ( .A(n10726), .B(n10725), .Z(n10891) );
  NAND U11185 ( .A(n10728), .B(n10727), .Z(n10732) );
  NAND U11186 ( .A(n10730), .B(n10729), .Z(n10731) );
  NAND U11187 ( .A(n10732), .B(n10731), .Z(n10890) );
  XOR U11188 ( .A(n10891), .B(n10890), .Z(n10893) );
  XOR U11189 ( .A(n10892), .B(n10893), .Z(n10956) );
  NAND U11190 ( .A(n10734), .B(n10733), .Z(n10738) );
  NANDN U11191 ( .A(n10736), .B(n10735), .Z(n10737) );
  NAND U11192 ( .A(n10738), .B(n10737), .Z(n10954) );
  NAND U11193 ( .A(n10740), .B(n10739), .Z(n10744) );
  NAND U11194 ( .A(n10742), .B(n10741), .Z(n10743) );
  NAND U11195 ( .A(n10744), .B(n10743), .Z(n10837) );
  AND U11196 ( .A(n10746), .B(n10745), .Z(n10750) );
  NAND U11197 ( .A(n10748), .B(n10747), .Z(n10749) );
  NANDN U11198 ( .A(n10750), .B(n10749), .Z(n10836) );
  XOR U11199 ( .A(n10837), .B(n10836), .Z(n10839) );
  NAND U11200 ( .A(y[752]), .B(x[135]), .Z(n10751) );
  XNOR U11201 ( .A(n10986), .B(n10751), .Z(n10910) );
  XOR U11202 ( .A(n10910), .B(n10752), .Z(n10843) );
  AND U11203 ( .A(x[138]), .B(y[749]), .Z(n10842) );
  XOR U11204 ( .A(n10843), .B(n10842), .Z(n10845) );
  AND U11205 ( .A(x[134]), .B(y[753]), .Z(n10901) );
  NAND U11206 ( .A(x[143]), .B(y[744]), .Z(n10902) );
  XNOR U11207 ( .A(n10901), .B(n10902), .Z(n10904) );
  AND U11208 ( .A(x[139]), .B(y[748]), .Z(n10903) );
  XOR U11209 ( .A(n10904), .B(n10903), .Z(n10844) );
  XOR U11210 ( .A(n10845), .B(n10844), .Z(n10838) );
  XOR U11211 ( .A(n10839), .B(n10838), .Z(n10955) );
  XNOR U11212 ( .A(n10954), .B(n10955), .Z(n10957) );
  NAND U11213 ( .A(n10754), .B(n10753), .Z(n10758) );
  NANDN U11214 ( .A(n10756), .B(n10755), .Z(n10757) );
  NAND U11215 ( .A(n10758), .B(n10757), .Z(n10936) );
  AND U11216 ( .A(x[146]), .B(y[746]), .Z(n11659) );
  NAND U11217 ( .A(n11659), .B(n10759), .Z(n10763) );
  NAND U11218 ( .A(n10761), .B(n10760), .Z(n10762) );
  NAND U11219 ( .A(n10763), .B(n10762), .Z(n10867) );
  NAND U11220 ( .A(n10765), .B(n10764), .Z(n10769) );
  NAND U11221 ( .A(n10767), .B(n10766), .Z(n10768) );
  NAND U11222 ( .A(n10769), .B(n10768), .Z(n10866) );
  XOR U11223 ( .A(n10867), .B(n10866), .Z(n10868) );
  NANDN U11224 ( .A(n10911), .B(n10909), .Z(n10773) );
  NAND U11225 ( .A(n10771), .B(n10770), .Z(n10772) );
  NAND U11226 ( .A(n10773), .B(n10772), .Z(n10880) );
  AND U11227 ( .A(x[128]), .B(y[759]), .Z(n10921) );
  AND U11228 ( .A(x[151]), .B(y[736]), .Z(n10920) );
  XOR U11229 ( .A(n10921), .B(n10920), .Z(n10923) );
  AND U11230 ( .A(x[150]), .B(y[737]), .Z(n10900) );
  XOR U11231 ( .A(n10900), .B(o[119]), .Z(n10922) );
  XOR U11232 ( .A(n10923), .B(n10922), .Z(n10879) );
  AND U11233 ( .A(x[148]), .B(y[739]), .Z(n11515) );
  NAND U11234 ( .A(y[743]), .B(x[144]), .Z(n10774) );
  XNOR U11235 ( .A(n11515), .B(n10774), .Z(n10896) );
  NAND U11236 ( .A(x[147]), .B(y[740]), .Z(n10897) );
  XNOR U11237 ( .A(n10896), .B(n10897), .Z(n10878) );
  XOR U11238 ( .A(n10879), .B(n10878), .Z(n10881) );
  XNOR U11239 ( .A(n10880), .B(n10881), .Z(n10869) );
  XOR U11240 ( .A(n10936), .B(n10937), .Z(n10939) );
  NAND U11241 ( .A(x[148]), .B(y[745]), .Z(n11870) );
  NANDN U11242 ( .A(n11870), .B(n10775), .Z(n10779) );
  NAND U11243 ( .A(n10777), .B(n10776), .Z(n10778) );
  NAND U11244 ( .A(n10779), .B(n10778), .Z(n10930) );
  NAND U11245 ( .A(n10781), .B(n10780), .Z(n10785) );
  NAND U11246 ( .A(n10783), .B(n10782), .Z(n10784) );
  NAND U11247 ( .A(n10785), .B(n10784), .Z(n10886) );
  AND U11248 ( .A(x[141]), .B(y[746]), .Z(n10861) );
  AND U11249 ( .A(x[130]), .B(y[757]), .Z(n10860) );
  XOR U11250 ( .A(n10861), .B(n10860), .Z(n10863) );
  AND U11251 ( .A(x[149]), .B(y[738]), .Z(n10862) );
  XOR U11252 ( .A(n10863), .B(n10862), .Z(n10885) );
  AND U11253 ( .A(n10786), .B(o[118]), .Z(n10917) );
  AND U11254 ( .A(x[140]), .B(y[747]), .Z(n10915) );
  AND U11255 ( .A(x[129]), .B(y[758]), .Z(n10914) );
  XOR U11256 ( .A(n10915), .B(n10914), .Z(n10916) );
  XOR U11257 ( .A(n10917), .B(n10916), .Z(n10884) );
  XOR U11258 ( .A(n10885), .B(n10884), .Z(n10887) );
  XOR U11259 ( .A(n10886), .B(n10887), .Z(n10931) );
  XOR U11260 ( .A(n10930), .B(n10931), .Z(n10933) );
  AND U11261 ( .A(x[143]), .B(y[752]), .Z(n12088) );
  NAND U11262 ( .A(n12088), .B(n10787), .Z(n10791) );
  NANDN U11263 ( .A(n10789), .B(n10788), .Z(n10790) );
  NAND U11264 ( .A(n10791), .B(n10790), .Z(n10874) );
  AND U11265 ( .A(x[142]), .B(y[745]), .Z(n10855) );
  AND U11266 ( .A(x[131]), .B(y[756]), .Z(n10854) );
  XOR U11267 ( .A(n10855), .B(n10854), .Z(n10857) );
  AND U11268 ( .A(x[132]), .B(y[755]), .Z(n10856) );
  XOR U11269 ( .A(n10857), .B(n10856), .Z(n10873) );
  AND U11270 ( .A(x[133]), .B(y[754]), .Z(n10848) );
  NAND U11271 ( .A(x[146]), .B(y[741]), .Z(n10849) );
  XNOR U11272 ( .A(n10848), .B(n10849), .Z(n10851) );
  AND U11273 ( .A(x[145]), .B(y[742]), .Z(n10850) );
  XOR U11274 ( .A(n10851), .B(n10850), .Z(n10872) );
  XOR U11275 ( .A(n10873), .B(n10872), .Z(n10875) );
  XOR U11276 ( .A(n10874), .B(n10875), .Z(n10932) );
  XOR U11277 ( .A(n10933), .B(n10932), .Z(n10938) );
  XOR U11278 ( .A(n10939), .B(n10938), .Z(n10942) );
  XOR U11279 ( .A(n10943), .B(n10942), .Z(n10944) );
  XOR U11280 ( .A(n10945), .B(n10944), .Z(n10832) );
  NANDN U11281 ( .A(n10793), .B(n10792), .Z(n10797) );
  NAND U11282 ( .A(n10795), .B(n10794), .Z(n10796) );
  AND U11283 ( .A(n10797), .B(n10796), .Z(n10951) );
  NAND U11284 ( .A(n10799), .B(n10798), .Z(n10803) );
  NAND U11285 ( .A(n10801), .B(n10800), .Z(n10802) );
  AND U11286 ( .A(n10803), .B(n10802), .Z(n10949) );
  NANDN U11287 ( .A(n10805), .B(n10804), .Z(n10809) );
  NAND U11288 ( .A(n10807), .B(n10806), .Z(n10808) );
  NAND U11289 ( .A(n10809), .B(n10808), .Z(n10948) );
  XNOR U11290 ( .A(n10949), .B(n10948), .Z(n10950) );
  XOR U11291 ( .A(n10951), .B(n10950), .Z(n10831) );
  NANDN U11292 ( .A(n10811), .B(n10810), .Z(n10815) );
  NAND U11293 ( .A(n10813), .B(n10812), .Z(n10814) );
  NAND U11294 ( .A(n10815), .B(n10814), .Z(n10830) );
  XOR U11295 ( .A(n10831), .B(n10830), .Z(n10833) );
  XOR U11296 ( .A(n10832), .B(n10833), .Z(n10960) );
  XNOR U11297 ( .A(n10963), .B(n10962), .Z(n10969) );
  NOR U11298 ( .A(n10816), .B(n10820), .Z(n10818) );
  OR U11299 ( .A(n10818), .B(n10817), .Z(n10822) );
  ANDN U11300 ( .B(n10820), .A(n10819), .Z(n10821) );
  ANDN U11301 ( .B(n10822), .A(n10821), .Z(n10967) );
  NANDN U11302 ( .A(n10824), .B(n10823), .Z(n10828) );
  NAND U11303 ( .A(n10826), .B(n10825), .Z(n10827) );
  AND U11304 ( .A(n10828), .B(n10827), .Z(n10968) );
  IV U11305 ( .A(n10968), .Z(n10966) );
  XOR U11306 ( .A(n10967), .B(n10966), .Z(n10829) );
  XNOR U11307 ( .A(n10969), .B(n10829), .Z(N248) );
  NAND U11308 ( .A(n10831), .B(n10830), .Z(n10835) );
  NAND U11309 ( .A(n10833), .B(n10832), .Z(n10834) );
  AND U11310 ( .A(n10835), .B(n10834), .Z(n11107) );
  NAND U11311 ( .A(n10837), .B(n10836), .Z(n10841) );
  NAND U11312 ( .A(n10839), .B(n10838), .Z(n10840) );
  NAND U11313 ( .A(n10841), .B(n10840), .Z(n11041) );
  NAND U11314 ( .A(n10843), .B(n10842), .Z(n10847) );
  NAND U11315 ( .A(n10845), .B(n10844), .Z(n10846) );
  NAND U11316 ( .A(n10847), .B(n10846), .Z(n11039) );
  NANDN U11317 ( .A(n10849), .B(n10848), .Z(n10853) );
  NAND U11318 ( .A(n10851), .B(n10850), .Z(n10852) );
  AND U11319 ( .A(n10853), .B(n10852), .Z(n11077) );
  AND U11320 ( .A(x[128]), .B(y[760]), .Z(n11027) );
  NAND U11321 ( .A(x[152]), .B(y[736]), .Z(n11028) );
  XNOR U11322 ( .A(n11027), .B(n11028), .Z(n11030) );
  NAND U11323 ( .A(x[151]), .B(y[737]), .Z(n11014) );
  XNOR U11324 ( .A(o[120]), .B(n11014), .Z(n11029) );
  XOR U11325 ( .A(n11030), .B(n11029), .Z(n11075) );
  AND U11326 ( .A(x[135]), .B(y[753]), .Z(n11008) );
  NAND U11327 ( .A(x[146]), .B(y[742]), .Z(n11009) );
  NAND U11328 ( .A(x[145]), .B(y[743]), .Z(n11011) );
  XOR U11329 ( .A(n11075), .B(n11074), .Z(n11076) );
  XNOR U11330 ( .A(n11077), .B(n11076), .Z(n11053) );
  NAND U11331 ( .A(n10855), .B(n10854), .Z(n10859) );
  NAND U11332 ( .A(n10857), .B(n10856), .Z(n10858) );
  NAND U11333 ( .A(n10859), .B(n10858), .Z(n11052) );
  NAND U11334 ( .A(n10861), .B(n10860), .Z(n10865) );
  NAND U11335 ( .A(n10863), .B(n10862), .Z(n10864) );
  NAND U11336 ( .A(n10865), .B(n10864), .Z(n11051) );
  XNOR U11337 ( .A(n11052), .B(n11051), .Z(n11054) );
  XOR U11338 ( .A(n11039), .B(n11040), .Z(n11042) );
  XOR U11339 ( .A(n11041), .B(n11042), .Z(n11048) );
  NAND U11340 ( .A(n10867), .B(n10866), .Z(n10871) );
  NANDN U11341 ( .A(n10869), .B(n10868), .Z(n10870) );
  AND U11342 ( .A(n10871), .B(n10870), .Z(n11095) );
  NAND U11343 ( .A(n10873), .B(n10872), .Z(n10877) );
  NAND U11344 ( .A(n10875), .B(n10874), .Z(n10876) );
  AND U11345 ( .A(n10877), .B(n10876), .Z(n11093) );
  NAND U11346 ( .A(n10879), .B(n10878), .Z(n10883) );
  NAND U11347 ( .A(n10881), .B(n10880), .Z(n10882) );
  AND U11348 ( .A(n10883), .B(n10882), .Z(n11092) );
  XOR U11349 ( .A(n11093), .B(n11092), .Z(n11094) );
  XOR U11350 ( .A(n11095), .B(n11094), .Z(n11046) );
  NAND U11351 ( .A(n10885), .B(n10884), .Z(n10889) );
  NAND U11352 ( .A(n10887), .B(n10886), .Z(n10888) );
  AND U11353 ( .A(n10889), .B(n10888), .Z(n11045) );
  XOR U11354 ( .A(n11046), .B(n11045), .Z(n11047) );
  XNOR U11355 ( .A(n11048), .B(n11047), .Z(n10975) );
  NAND U11356 ( .A(n10891), .B(n10890), .Z(n10895) );
  NAND U11357 ( .A(n10893), .B(n10892), .Z(n10894) );
  AND U11358 ( .A(n10895), .B(n10894), .Z(n10974) );
  XOR U11359 ( .A(n10975), .B(n10974), .Z(n10977) );
  AND U11360 ( .A(x[148]), .B(y[743]), .Z(n11412) );
  AND U11361 ( .A(x[144]), .B(y[739]), .Z(n11063) );
  NAND U11362 ( .A(n11412), .B(n11063), .Z(n10899) );
  NANDN U11363 ( .A(n10897), .B(n10896), .Z(n10898) );
  AND U11364 ( .A(n10899), .B(n10898), .Z(n11083) );
  AND U11365 ( .A(x[150]), .B(y[738]), .Z(n10996) );
  XOR U11366 ( .A(n10997), .B(n10996), .Z(n10999) );
  NAND U11367 ( .A(x[130]), .B(y[758]), .Z(n10998) );
  AND U11368 ( .A(n10900), .B(o[119]), .Z(n11003) );
  AND U11369 ( .A(x[129]), .B(y[759]), .Z(n11004) );
  XOR U11370 ( .A(n11005), .B(n11004), .Z(n11002) );
  XOR U11371 ( .A(n11003), .B(n11002), .Z(n11080) );
  XOR U11372 ( .A(n11081), .B(n11080), .Z(n11082) );
  XNOR U11373 ( .A(n11083), .B(n11082), .Z(n11034) );
  NANDN U11374 ( .A(n10902), .B(n10901), .Z(n10906) );
  NAND U11375 ( .A(n10904), .B(n10903), .Z(n10905) );
  AND U11376 ( .A(n10906), .B(n10905), .Z(n11089) );
  AND U11377 ( .A(y[739]), .B(x[149]), .Z(n10908) );
  NAND U11378 ( .A(y[744]), .B(x[144]), .Z(n10907) );
  XNOR U11379 ( .A(n10908), .B(n10907), .Z(n11064) );
  NAND U11380 ( .A(x[133]), .B(y[755]), .Z(n11065) );
  XNOR U11381 ( .A(n11064), .B(n11065), .Z(n11087) );
  AND U11382 ( .A(x[134]), .B(y[754]), .Z(n11399) );
  NAND U11383 ( .A(x[148]), .B(y[740]), .Z(n11213) );
  XNOR U11384 ( .A(n11399), .B(n11213), .Z(n11070) );
  NAND U11385 ( .A(x[147]), .B(y[741]), .Z(n11071) );
  XNOR U11386 ( .A(n11070), .B(n11071), .Z(n11086) );
  XOR U11387 ( .A(n11087), .B(n11086), .Z(n11088) );
  XNOR U11388 ( .A(n11089), .B(n11088), .Z(n11060) );
  NANDN U11389 ( .A(n11139), .B(n10909), .Z(n10913) );
  NANDN U11390 ( .A(n10911), .B(n10910), .Z(n10912) );
  NAND U11391 ( .A(n10913), .B(n10912), .Z(n11058) );
  NAND U11392 ( .A(n10915), .B(n10914), .Z(n10919) );
  NAND U11393 ( .A(n10917), .B(n10916), .Z(n10918) );
  NAND U11394 ( .A(n10919), .B(n10918), .Z(n11057) );
  XOR U11395 ( .A(n11058), .B(n11057), .Z(n11059) );
  XOR U11396 ( .A(n11060), .B(n11059), .Z(n11033) );
  XOR U11397 ( .A(n11034), .B(n11033), .Z(n11036) );
  NAND U11398 ( .A(n10921), .B(n10920), .Z(n10925) );
  NAND U11399 ( .A(n10923), .B(n10922), .Z(n10924) );
  NAND U11400 ( .A(n10925), .B(n10924), .Z(n11015) );
  AND U11401 ( .A(x[131]), .B(y[757]), .Z(n11021) );
  XOR U11402 ( .A(n11022), .B(n11021), .Z(n11024) );
  NAND U11403 ( .A(x[132]), .B(y[756]), .Z(n11023) );
  XNOR U11404 ( .A(n11024), .B(n11023), .Z(n11016) );
  XOR U11405 ( .A(n11015), .B(n11016), .Z(n11018) );
  AND U11406 ( .A(y[751]), .B(x[137]), .Z(n10927) );
  NAND U11407 ( .A(y[750]), .B(x[138]), .Z(n10926) );
  XNOR U11408 ( .A(n10927), .B(n10926), .Z(n10988) );
  AND U11409 ( .A(y[746]), .B(x[142]), .Z(n10929) );
  NAND U11410 ( .A(y[752]), .B(x[136]), .Z(n10928) );
  XNOR U11411 ( .A(n10929), .B(n10928), .Z(n10992) );
  NAND U11412 ( .A(x[139]), .B(y[749]), .Z(n10993) );
  XNOR U11413 ( .A(n10992), .B(n10993), .Z(n10987) );
  XOR U11414 ( .A(n10988), .B(n10987), .Z(n11017) );
  XOR U11415 ( .A(n11018), .B(n11017), .Z(n11035) );
  XOR U11416 ( .A(n11036), .B(n11035), .Z(n10981) );
  NAND U11417 ( .A(n10931), .B(n10930), .Z(n10935) );
  NAND U11418 ( .A(n10933), .B(n10932), .Z(n10934) );
  AND U11419 ( .A(n10935), .B(n10934), .Z(n10980) );
  XNOR U11420 ( .A(n10981), .B(n10980), .Z(n10983) );
  NAND U11421 ( .A(n10937), .B(n10936), .Z(n10941) );
  NAND U11422 ( .A(n10939), .B(n10938), .Z(n10940) );
  AND U11423 ( .A(n10941), .B(n10940), .Z(n10982) );
  XOR U11424 ( .A(n10983), .B(n10982), .Z(n10976) );
  XOR U11425 ( .A(n10977), .B(n10976), .Z(n11105) );
  NAND U11426 ( .A(n10943), .B(n10942), .Z(n10947) );
  NANDN U11427 ( .A(n10945), .B(n10944), .Z(n10946) );
  NAND U11428 ( .A(n10947), .B(n10946), .Z(n11100) );
  NANDN U11429 ( .A(n10949), .B(n10948), .Z(n10953) );
  NANDN U11430 ( .A(n10951), .B(n10950), .Z(n10952) );
  NAND U11431 ( .A(n10953), .B(n10952), .Z(n11099) );
  NAND U11432 ( .A(n10955), .B(n10954), .Z(n10959) );
  NANDN U11433 ( .A(n10957), .B(n10956), .Z(n10958) );
  NAND U11434 ( .A(n10959), .B(n10958), .Z(n11098) );
  XOR U11435 ( .A(n11099), .B(n11098), .Z(n11101) );
  XOR U11436 ( .A(n11100), .B(n11101), .Z(n11104) );
  XNOR U11437 ( .A(n11105), .B(n11104), .Z(n11106) );
  XOR U11438 ( .A(n11107), .B(n11106), .Z(n11112) );
  NANDN U11439 ( .A(n10961), .B(n10960), .Z(n10965) );
  NAND U11440 ( .A(n10963), .B(n10962), .Z(n10964) );
  NAND U11441 ( .A(n10965), .B(n10964), .Z(n11110) );
  NANDN U11442 ( .A(n10966), .B(n10967), .Z(n10972) );
  NOR U11443 ( .A(n10968), .B(n10967), .Z(n10970) );
  OR U11444 ( .A(n10970), .B(n10969), .Z(n10971) );
  AND U11445 ( .A(n10972), .B(n10971), .Z(n11111) );
  XOR U11446 ( .A(n11110), .B(n11111), .Z(n10973) );
  XNOR U11447 ( .A(n11112), .B(n10973), .Z(N249) );
  NAND U11448 ( .A(n10975), .B(n10974), .Z(n10979) );
  NAND U11449 ( .A(n10977), .B(n10976), .Z(n10978) );
  NAND U11450 ( .A(n10979), .B(n10978), .Z(n11257) );
  NANDN U11451 ( .A(n10981), .B(n10980), .Z(n10985) );
  NAND U11452 ( .A(n10983), .B(n10982), .Z(n10984) );
  NAND U11453 ( .A(n10985), .B(n10984), .Z(n11114) );
  NANDN U11454 ( .A(n11138), .B(n10986), .Z(n10990) );
  NAND U11455 ( .A(n10988), .B(n10987), .Z(n10989) );
  AND U11456 ( .A(n10990), .B(n10989), .Z(n11163) );
  AND U11457 ( .A(x[142]), .B(y[752]), .Z(n12064) );
  NAND U11458 ( .A(n12064), .B(n10991), .Z(n10995) );
  NANDN U11459 ( .A(n10993), .B(n10992), .Z(n10994) );
  NAND U11460 ( .A(n10995), .B(n10994), .Z(n11190) );
  NAND U11461 ( .A(x[139]), .B(y[750]), .Z(n11209) );
  NAND U11462 ( .A(x[140]), .B(y[749]), .Z(n11208) );
  NAND U11463 ( .A(x[135]), .B(y[754]), .Z(n11207) );
  XOR U11464 ( .A(n11208), .B(n11207), .Z(n11210) );
  XOR U11465 ( .A(n11209), .B(n11210), .Z(n11189) );
  NAND U11466 ( .A(x[152]), .B(y[737]), .Z(n11206) );
  XNOR U11467 ( .A(o[121]), .B(n11206), .Z(n11177) );
  AND U11468 ( .A(x[129]), .B(y[760]), .Z(n11176) );
  XOR U11469 ( .A(n11177), .B(n11176), .Z(n11179) );
  AND U11470 ( .A(x[141]), .B(y[748]), .Z(n11178) );
  XOR U11471 ( .A(n11179), .B(n11178), .Z(n11188) );
  XNOR U11472 ( .A(n11189), .B(n11188), .Z(n11191) );
  XOR U11473 ( .A(n11190), .B(n11191), .Z(n11162) );
  XNOR U11474 ( .A(n11163), .B(n11162), .Z(n11165) );
  NAND U11475 ( .A(n10997), .B(n10996), .Z(n11001) );
  ANDN U11476 ( .B(n10999), .A(n10998), .Z(n11000) );
  ANDN U11477 ( .B(n11001), .A(n11000), .Z(n11151) );
  AND U11478 ( .A(n11003), .B(n11002), .Z(n11007) );
  NAND U11479 ( .A(n11005), .B(n11004), .Z(n11006) );
  NANDN U11480 ( .A(n11007), .B(n11006), .Z(n11150) );
  NANDN U11481 ( .A(n11009), .B(n11008), .Z(n11013) );
  NANDN U11482 ( .A(n11011), .B(n11010), .Z(n11012) );
  AND U11483 ( .A(n11013), .B(n11012), .Z(n11147) );
  NAND U11484 ( .A(x[136]), .B(y[753]), .Z(n11140) );
  XNOR U11485 ( .A(n11139), .B(n11138), .Z(n11141) );
  XOR U11486 ( .A(n11140), .B(n11141), .Z(n11145) );
  NANDN U11487 ( .A(n11014), .B(o[120]), .Z(n11134) );
  NAND U11488 ( .A(x[153]), .B(y[736]), .Z(n11133) );
  NAND U11489 ( .A(x[128]), .B(y[761]), .Z(n11132) );
  XNOR U11490 ( .A(n11133), .B(n11132), .Z(n11135) );
  XOR U11491 ( .A(n11134), .B(n11135), .Z(n11144) );
  XOR U11492 ( .A(n11145), .B(n11144), .Z(n11146) );
  XOR U11493 ( .A(n11153), .B(n11152), .Z(n11164) );
  XOR U11494 ( .A(n11165), .B(n11164), .Z(n11245) );
  NAND U11495 ( .A(n11016), .B(n11015), .Z(n11020) );
  NAND U11496 ( .A(n11018), .B(n11017), .Z(n11019) );
  AND U11497 ( .A(n11020), .B(n11019), .Z(n11242) );
  NAND U11498 ( .A(n11022), .B(n11021), .Z(n11026) );
  ANDN U11499 ( .B(n11024), .A(n11023), .Z(n11025) );
  ANDN U11500 ( .B(n11026), .A(n11025), .Z(n11227) );
  NANDN U11501 ( .A(n11028), .B(n11027), .Z(n11032) );
  NAND U11502 ( .A(n11030), .B(n11029), .Z(n11031) );
  AND U11503 ( .A(n11032), .B(n11031), .Z(n11225) );
  AND U11504 ( .A(x[142]), .B(y[747]), .Z(n11183) );
  AND U11505 ( .A(x[130]), .B(y[759]), .Z(n11182) );
  XOR U11506 ( .A(n11183), .B(n11182), .Z(n11185) );
  AND U11507 ( .A(x[131]), .B(y[758]), .Z(n11184) );
  XOR U11508 ( .A(n11185), .B(n11184), .Z(n11224) );
  XNOR U11509 ( .A(n11225), .B(n11224), .Z(n11226) );
  XNOR U11510 ( .A(n11227), .B(n11226), .Z(n11243) );
  NAND U11511 ( .A(n11034), .B(n11033), .Z(n11038) );
  NAND U11512 ( .A(n11036), .B(n11035), .Z(n11037) );
  AND U11513 ( .A(n11038), .B(n11037), .Z(n11248) );
  XOR U11514 ( .A(n11249), .B(n11248), .Z(n11251) );
  NAND U11515 ( .A(n11040), .B(n11039), .Z(n11044) );
  NAND U11516 ( .A(n11042), .B(n11041), .Z(n11043) );
  AND U11517 ( .A(n11044), .B(n11043), .Z(n11250) );
  XOR U11518 ( .A(n11251), .B(n11250), .Z(n11115) );
  XOR U11519 ( .A(n11114), .B(n11115), .Z(n11116) );
  NAND U11520 ( .A(n11046), .B(n11045), .Z(n11050) );
  NANDN U11521 ( .A(n11048), .B(n11047), .Z(n11049) );
  NAND U11522 ( .A(n11050), .B(n11049), .Z(n11122) );
  NAND U11523 ( .A(n11052), .B(n11051), .Z(n11056) );
  NANDN U11524 ( .A(n11054), .B(n11053), .Z(n11055) );
  NAND U11525 ( .A(n11056), .B(n11055), .Z(n11127) );
  NAND U11526 ( .A(n11058), .B(n11057), .Z(n11062) );
  NAND U11527 ( .A(n11060), .B(n11059), .Z(n11061) );
  NAND U11528 ( .A(n11062), .B(n11061), .Z(n11126) );
  XOR U11529 ( .A(n11127), .B(n11126), .Z(n11128) );
  AND U11530 ( .A(x[149]), .B(y[744]), .Z(n12033) );
  NAND U11531 ( .A(n12033), .B(n11063), .Z(n11067) );
  NANDN U11532 ( .A(n11065), .B(n11064), .Z(n11066) );
  AND U11533 ( .A(n11067), .B(n11066), .Z(n11233) );
  NAND U11534 ( .A(x[150]), .B(y[739]), .Z(n11202) );
  NAND U11535 ( .A(x[133]), .B(y[756]), .Z(n11201) );
  NAND U11536 ( .A(x[145]), .B(y[744]), .Z(n11200) );
  XNOR U11537 ( .A(n11201), .B(n11200), .Z(n11203) );
  XOR U11538 ( .A(n11202), .B(n11203), .Z(n11230) );
  AND U11539 ( .A(y[741]), .B(x[148]), .Z(n11069) );
  NAND U11540 ( .A(y[740]), .B(x[149]), .Z(n11068) );
  XNOR U11541 ( .A(n11069), .B(n11068), .Z(n11215) );
  AND U11542 ( .A(x[147]), .B(y[742]), .Z(n11214) );
  XOR U11543 ( .A(n11215), .B(n11214), .Z(n11231) );
  XOR U11544 ( .A(n11230), .B(n11231), .Z(n11232) );
  XOR U11545 ( .A(n11233), .B(n11232), .Z(n11157) );
  NANDN U11546 ( .A(n11213), .B(n11399), .Z(n11073) );
  NANDN U11547 ( .A(n11071), .B(n11070), .Z(n11072) );
  AND U11548 ( .A(n11073), .B(n11072), .Z(n11239) );
  NAND U11549 ( .A(x[143]), .B(y[746]), .Z(n11220) );
  NAND U11550 ( .A(x[146]), .B(y[743]), .Z(n11219) );
  NAND U11551 ( .A(x[134]), .B(y[755]), .Z(n11218) );
  XNOR U11552 ( .A(n11219), .B(n11218), .Z(n11221) );
  XOR U11553 ( .A(n11220), .B(n11221), .Z(n11237) );
  NAND U11554 ( .A(x[151]), .B(y[738]), .Z(n11196) );
  NAND U11555 ( .A(x[132]), .B(y[757]), .Z(n11195) );
  NAND U11556 ( .A(x[144]), .B(y[745]), .Z(n11194) );
  XNOR U11557 ( .A(n11195), .B(n11194), .Z(n11197) );
  XOR U11558 ( .A(n11196), .B(n11197), .Z(n11236) );
  XOR U11559 ( .A(n11237), .B(n11236), .Z(n11238) );
  XOR U11560 ( .A(n11239), .B(n11238), .Z(n11156) );
  XOR U11561 ( .A(n11157), .B(n11156), .Z(n11159) );
  NAND U11562 ( .A(n11075), .B(n11074), .Z(n11079) );
  NANDN U11563 ( .A(n11077), .B(n11076), .Z(n11078) );
  AND U11564 ( .A(n11079), .B(n11078), .Z(n11158) );
  XOR U11565 ( .A(n11159), .B(n11158), .Z(n11171) );
  NAND U11566 ( .A(n11081), .B(n11080), .Z(n11085) );
  NANDN U11567 ( .A(n11083), .B(n11082), .Z(n11084) );
  AND U11568 ( .A(n11085), .B(n11084), .Z(n11169) );
  NAND U11569 ( .A(n11087), .B(n11086), .Z(n11091) );
  NANDN U11570 ( .A(n11089), .B(n11088), .Z(n11090) );
  NAND U11571 ( .A(n11091), .B(n11090), .Z(n11168) );
  XNOR U11572 ( .A(n11169), .B(n11168), .Z(n11170) );
  XOR U11573 ( .A(n11171), .B(n11170), .Z(n11129) );
  XNOR U11574 ( .A(n11128), .B(n11129), .Z(n11121) );
  NAND U11575 ( .A(n11093), .B(n11092), .Z(n11097) );
  NAND U11576 ( .A(n11095), .B(n11094), .Z(n11096) );
  NAND U11577 ( .A(n11097), .B(n11096), .Z(n11120) );
  XOR U11578 ( .A(n11122), .B(n11123), .Z(n11117) );
  XNOR U11579 ( .A(n11116), .B(n11117), .Z(n11258) );
  XOR U11580 ( .A(n11257), .B(n11258), .Z(n11260) );
  NAND U11581 ( .A(n11099), .B(n11098), .Z(n11103) );
  NAND U11582 ( .A(n11101), .B(n11100), .Z(n11102) );
  AND U11583 ( .A(n11103), .B(n11102), .Z(n11259) );
  XOR U11584 ( .A(n11260), .B(n11259), .Z(n11256) );
  NANDN U11585 ( .A(n11105), .B(n11104), .Z(n11109) );
  NAND U11586 ( .A(n11107), .B(n11106), .Z(n11108) );
  NAND U11587 ( .A(n11109), .B(n11108), .Z(n11255) );
  XOR U11588 ( .A(n11255), .B(n11254), .Z(n11113) );
  XNOR U11589 ( .A(n11256), .B(n11113), .Z(N250) );
  NAND U11590 ( .A(n11115), .B(n11114), .Z(n11119) );
  NANDN U11591 ( .A(n11117), .B(n11116), .Z(n11118) );
  AND U11592 ( .A(n11119), .B(n11118), .Z(n11265) );
  NANDN U11593 ( .A(n11121), .B(n11120), .Z(n11125) );
  NANDN U11594 ( .A(n11123), .B(n11122), .Z(n11124) );
  AND U11595 ( .A(n11125), .B(n11124), .Z(n11264) );
  XOR U11596 ( .A(n11265), .B(n11264), .Z(n11267) );
  NAND U11597 ( .A(n11127), .B(n11126), .Z(n11131) );
  NANDN U11598 ( .A(n11129), .B(n11128), .Z(n11130) );
  NAND U11599 ( .A(n11131), .B(n11130), .Z(n11285) );
  AND U11600 ( .A(x[130]), .B(y[760]), .Z(n11301) );
  XOR U11601 ( .A(n11302), .B(n11301), .Z(n11304) );
  AND U11602 ( .A(x[152]), .B(y[738]), .Z(n11303) );
  XOR U11603 ( .A(n11304), .B(n11303), .Z(n11338) );
  NAND U11604 ( .A(n11133), .B(n11132), .Z(n11137) );
  NANDN U11605 ( .A(n11135), .B(n11134), .Z(n11136) );
  AND U11606 ( .A(n11137), .B(n11136), .Z(n11337) );
  XOR U11607 ( .A(n11338), .B(n11337), .Z(n11340) );
  NAND U11608 ( .A(n11139), .B(n11138), .Z(n11143) );
  NANDN U11609 ( .A(n11141), .B(n11140), .Z(n11142) );
  AND U11610 ( .A(n11143), .B(n11142), .Z(n11339) );
  XOR U11611 ( .A(n11340), .B(n11339), .Z(n11414) );
  NAND U11612 ( .A(n11145), .B(n11144), .Z(n11149) );
  NANDN U11613 ( .A(n11147), .B(n11146), .Z(n11148) );
  AND U11614 ( .A(n11149), .B(n11148), .Z(n11413) );
  NANDN U11615 ( .A(n11151), .B(n11150), .Z(n11155) );
  NAND U11616 ( .A(n11153), .B(n11152), .Z(n11154) );
  NAND U11617 ( .A(n11155), .B(n11154), .Z(n11416) );
  NAND U11618 ( .A(n11157), .B(n11156), .Z(n11161) );
  NAND U11619 ( .A(n11159), .B(n11158), .Z(n11160) );
  AND U11620 ( .A(n11161), .B(n11160), .Z(n11376) );
  NANDN U11621 ( .A(n11163), .B(n11162), .Z(n11167) );
  NAND U11622 ( .A(n11165), .B(n11164), .Z(n11166) );
  AND U11623 ( .A(n11167), .B(n11166), .Z(n11375) );
  XNOR U11624 ( .A(n11376), .B(n11375), .Z(n11377) );
  XOR U11625 ( .A(n11378), .B(n11377), .Z(n11284) );
  NANDN U11626 ( .A(n11169), .B(n11168), .Z(n11173) );
  NANDN U11627 ( .A(n11171), .B(n11170), .Z(n11172) );
  AND U11628 ( .A(n11173), .B(n11172), .Z(n11372) );
  AND U11629 ( .A(x[140]), .B(y[750]), .Z(n11456) );
  AND U11630 ( .A(x[133]), .B(y[757]), .Z(n11352) );
  XOR U11631 ( .A(n11456), .B(n11352), .Z(n11354) );
  AND U11632 ( .A(x[138]), .B(y[752]), .Z(n11353) );
  XOR U11633 ( .A(n11354), .B(n11353), .Z(n11384) );
  AND U11634 ( .A(x[135]), .B(y[755]), .Z(n11382) );
  AND U11635 ( .A(y[756]), .B(x[134]), .Z(n11175) );
  NAND U11636 ( .A(y[754]), .B(x[136]), .Z(n11174) );
  XNOR U11637 ( .A(n11175), .B(n11174), .Z(n11401) );
  AND U11638 ( .A(x[137]), .B(y[753]), .Z(n11400) );
  XOR U11639 ( .A(n11401), .B(n11400), .Z(n11381) );
  XOR U11640 ( .A(n11382), .B(n11381), .Z(n11383) );
  XOR U11641 ( .A(n11384), .B(n11383), .Z(n11328) );
  NAND U11642 ( .A(n11177), .B(n11176), .Z(n11181) );
  NAND U11643 ( .A(n11179), .B(n11178), .Z(n11180) );
  AND U11644 ( .A(n11181), .B(n11180), .Z(n11326) );
  NAND U11645 ( .A(n11183), .B(n11182), .Z(n11187) );
  NAND U11646 ( .A(n11185), .B(n11184), .Z(n11186) );
  NAND U11647 ( .A(n11187), .B(n11186), .Z(n11325) );
  XNOR U11648 ( .A(n11326), .B(n11325), .Z(n11327) );
  XOR U11649 ( .A(n11328), .B(n11327), .Z(n11364) );
  NANDN U11650 ( .A(n11189), .B(n11188), .Z(n11193) );
  NAND U11651 ( .A(n11191), .B(n11190), .Z(n11192) );
  AND U11652 ( .A(n11193), .B(n11192), .Z(n11363) );
  XNOR U11653 ( .A(n11364), .B(n11363), .Z(n11366) );
  NAND U11654 ( .A(n11195), .B(n11194), .Z(n11199) );
  NANDN U11655 ( .A(n11197), .B(n11196), .Z(n11198) );
  AND U11656 ( .A(n11199), .B(n11198), .Z(n11289) );
  NAND U11657 ( .A(n11201), .B(n11200), .Z(n11205) );
  NANDN U11658 ( .A(n11203), .B(n11202), .Z(n11204) );
  NAND U11659 ( .A(n11205), .B(n11204), .Z(n11290) );
  XNOR U11660 ( .A(n11289), .B(n11290), .Z(n11292) );
  ANDN U11661 ( .B(o[121]), .A(n11206), .Z(n11393) );
  NAND U11662 ( .A(x[142]), .B(y[748]), .Z(n11394) );
  NAND U11663 ( .A(x[129]), .B(y[761]), .Z(n11396) );
  NAND U11664 ( .A(x[153]), .B(y[737]), .Z(n11404) );
  AND U11665 ( .A(x[154]), .B(y[736]), .Z(n11357) );
  XOR U11666 ( .A(n11358), .B(n11357), .Z(n11360) );
  AND U11667 ( .A(x[128]), .B(y[762]), .Z(n11359) );
  XOR U11668 ( .A(n11360), .B(n11359), .Z(n11343) );
  XOR U11669 ( .A(n11344), .B(n11343), .Z(n11346) );
  NAND U11670 ( .A(n11208), .B(n11207), .Z(n11212) );
  NAND U11671 ( .A(n11210), .B(n11209), .Z(n11211) );
  AND U11672 ( .A(n11212), .B(n11211), .Z(n11345) );
  XOR U11673 ( .A(n11346), .B(n11345), .Z(n11291) );
  XOR U11674 ( .A(n11292), .B(n11291), .Z(n11334) );
  AND U11675 ( .A(x[149]), .B(y[741]), .Z(n11387) );
  NANDN U11676 ( .A(n11213), .B(n11387), .Z(n11217) );
  NAND U11677 ( .A(n11215), .B(n11214), .Z(n11216) );
  AND U11678 ( .A(n11217), .B(n11216), .Z(n11322) );
  XOR U11679 ( .A(n11388), .B(n11387), .Z(n11389) );
  NAND U11680 ( .A(x[148]), .B(y[742]), .Z(n11390) );
  NAND U11681 ( .A(x[151]), .B(y[739]), .Z(n11308) );
  XNOR U11682 ( .A(n11307), .B(n11308), .Z(n11309) );
  NAND U11683 ( .A(x[150]), .B(y[740]), .Z(n11310) );
  XNOR U11684 ( .A(n11309), .B(n11310), .Z(n11319) );
  XOR U11685 ( .A(n11320), .B(n11319), .Z(n11321) );
  XOR U11686 ( .A(n11322), .B(n11321), .Z(n11332) );
  AND U11687 ( .A(x[131]), .B(y[759]), .Z(n11405) );
  NAND U11688 ( .A(x[147]), .B(y[743]), .Z(n11406) );
  NAND U11689 ( .A(x[139]), .B(y[751]), .Z(n11408) );
  AND U11690 ( .A(x[132]), .B(y[758]), .Z(n11313) );
  XOR U11691 ( .A(n11314), .B(n11313), .Z(n11315) );
  XOR U11692 ( .A(n11315), .B(n11316), .Z(n11295) );
  XOR U11693 ( .A(n11296), .B(n11295), .Z(n11298) );
  NAND U11694 ( .A(n11219), .B(n11218), .Z(n11223) );
  NANDN U11695 ( .A(n11221), .B(n11220), .Z(n11222) );
  AND U11696 ( .A(n11223), .B(n11222), .Z(n11297) );
  XNOR U11697 ( .A(n11298), .B(n11297), .Z(n11331) );
  XOR U11698 ( .A(n11332), .B(n11331), .Z(n11333) );
  XNOR U11699 ( .A(n11334), .B(n11333), .Z(n11365) );
  XOR U11700 ( .A(n11366), .B(n11365), .Z(n11370) );
  NANDN U11701 ( .A(n11225), .B(n11224), .Z(n11229) );
  NANDN U11702 ( .A(n11227), .B(n11226), .Z(n11228) );
  AND U11703 ( .A(n11229), .B(n11228), .Z(n11422) );
  NAND U11704 ( .A(n11231), .B(n11230), .Z(n11235) );
  NANDN U11705 ( .A(n11233), .B(n11232), .Z(n11234) );
  AND U11706 ( .A(n11235), .B(n11234), .Z(n11420) );
  NAND U11707 ( .A(n11237), .B(n11236), .Z(n11241) );
  NANDN U11708 ( .A(n11239), .B(n11238), .Z(n11240) );
  NAND U11709 ( .A(n11241), .B(n11240), .Z(n11419) );
  XNOR U11710 ( .A(n11370), .B(n11369), .Z(n11371) );
  XNOR U11711 ( .A(n11372), .B(n11371), .Z(n11283) );
  XOR U11712 ( .A(n11285), .B(n11286), .Z(n11280) );
  NANDN U11713 ( .A(n11243), .B(n11242), .Z(n11247) );
  NANDN U11714 ( .A(n11245), .B(n11244), .Z(n11246) );
  AND U11715 ( .A(n11247), .B(n11246), .Z(n11278) );
  NAND U11716 ( .A(n11249), .B(n11248), .Z(n11253) );
  NAND U11717 ( .A(n11251), .B(n11250), .Z(n11252) );
  AND U11718 ( .A(n11253), .B(n11252), .Z(n11277) );
  XOR U11719 ( .A(n11278), .B(n11277), .Z(n11279) );
  XOR U11720 ( .A(n11280), .B(n11279), .Z(n11266) );
  XNOR U11721 ( .A(n11267), .B(n11266), .Z(n11273) );
  NAND U11722 ( .A(n11258), .B(n11257), .Z(n11262) );
  NAND U11723 ( .A(n11260), .B(n11259), .Z(n11261) );
  AND U11724 ( .A(n11262), .B(n11261), .Z(n11271) );
  IV U11725 ( .A(n11271), .Z(n11270) );
  XOR U11726 ( .A(n11272), .B(n11270), .Z(n11263) );
  XNOR U11727 ( .A(n11273), .B(n11263), .Z(N251) );
  NAND U11728 ( .A(n11265), .B(n11264), .Z(n11269) );
  NAND U11729 ( .A(n11267), .B(n11266), .Z(n11268) );
  NAND U11730 ( .A(n11269), .B(n11268), .Z(n11577) );
  OR U11731 ( .A(n11272), .B(n11270), .Z(n11276) );
  ANDN U11732 ( .B(n11272), .A(n11271), .Z(n11274) );
  OR U11733 ( .A(n11274), .B(n11273), .Z(n11275) );
  AND U11734 ( .A(n11276), .B(n11275), .Z(n11578) );
  NAND U11735 ( .A(n11278), .B(n11277), .Z(n11282) );
  NAND U11736 ( .A(n11280), .B(n11279), .Z(n11281) );
  AND U11737 ( .A(n11282), .B(n11281), .Z(n11583) );
  NANDN U11738 ( .A(n11284), .B(n11283), .Z(n11288) );
  NAND U11739 ( .A(n11286), .B(n11285), .Z(n11287) );
  AND U11740 ( .A(n11288), .B(n11287), .Z(n11581) );
  NANDN U11741 ( .A(n11290), .B(n11289), .Z(n11294) );
  NAND U11742 ( .A(n11292), .B(n11291), .Z(n11293) );
  NAND U11743 ( .A(n11294), .B(n11293), .Z(n11555) );
  NAND U11744 ( .A(n11296), .B(n11295), .Z(n11300) );
  NAND U11745 ( .A(n11298), .B(n11297), .Z(n11299) );
  NAND U11746 ( .A(n11300), .B(n11299), .Z(n11553) );
  AND U11747 ( .A(n11302), .B(n11301), .Z(n11306) );
  NAND U11748 ( .A(n11304), .B(n11303), .Z(n11305) );
  NANDN U11749 ( .A(n11306), .B(n11305), .Z(n11480) );
  NANDN U11750 ( .A(n11308), .B(n11307), .Z(n11312) );
  NANDN U11751 ( .A(n11310), .B(n11309), .Z(n11311) );
  NAND U11752 ( .A(n11312), .B(n11311), .Z(n11479) );
  XOR U11753 ( .A(n11480), .B(n11479), .Z(n11481) );
  NAND U11754 ( .A(n11314), .B(n11313), .Z(n11318) );
  NAND U11755 ( .A(n11316), .B(n11315), .Z(n11317) );
  NAND U11756 ( .A(n11318), .B(n11317), .Z(n11493) );
  AND U11757 ( .A(x[128]), .B(y[763]), .Z(n11533) );
  AND U11758 ( .A(x[155]), .B(y[736]), .Z(n11532) );
  XOR U11759 ( .A(n11533), .B(n11532), .Z(n11535) );
  AND U11760 ( .A(x[154]), .B(y[737]), .Z(n11544) );
  XOR U11761 ( .A(n11544), .B(o[123]), .Z(n11534) );
  XOR U11762 ( .A(n11535), .B(n11534), .Z(n11492) );
  AND U11763 ( .A(x[137]), .B(y[754]), .Z(n11539) );
  AND U11764 ( .A(x[149]), .B(y[742]), .Z(n11538) );
  XOR U11765 ( .A(n11539), .B(n11538), .Z(n11541) );
  AND U11766 ( .A(x[146]), .B(y[745]), .Z(n11540) );
  XOR U11767 ( .A(n11541), .B(n11540), .Z(n11491) );
  XOR U11768 ( .A(n11492), .B(n11491), .Z(n11494) );
  XNOR U11769 ( .A(n11493), .B(n11494), .Z(n11482) );
  XOR U11770 ( .A(n11553), .B(n11554), .Z(n11556) );
  XOR U11771 ( .A(n11555), .B(n11556), .Z(n11574) );
  NAND U11772 ( .A(n11320), .B(n11319), .Z(n11324) );
  NANDN U11773 ( .A(n11322), .B(n11321), .Z(n11323) );
  AND U11774 ( .A(n11324), .B(n11323), .Z(n11572) );
  NANDN U11775 ( .A(n11326), .B(n11325), .Z(n11330) );
  NAND U11776 ( .A(n11328), .B(n11327), .Z(n11329) );
  AND U11777 ( .A(n11330), .B(n11329), .Z(n11571) );
  XOR U11778 ( .A(n11572), .B(n11571), .Z(n11573) );
  NAND U11779 ( .A(n11332), .B(n11331), .Z(n11336) );
  NANDN U11780 ( .A(n11334), .B(n11333), .Z(n11335) );
  AND U11781 ( .A(n11336), .B(n11335), .Z(n11559) );
  NAND U11782 ( .A(n11338), .B(n11337), .Z(n11342) );
  NAND U11783 ( .A(n11340), .B(n11339), .Z(n11341) );
  NAND U11784 ( .A(n11342), .B(n11341), .Z(n11549) );
  NAND U11785 ( .A(n11344), .B(n11343), .Z(n11348) );
  NAND U11786 ( .A(n11346), .B(n11345), .Z(n11347) );
  NAND U11787 ( .A(n11348), .B(n11347), .Z(n11547) );
  AND U11788 ( .A(x[134]), .B(y[757]), .Z(n11523) );
  AND U11789 ( .A(x[147]), .B(y[744]), .Z(n11521) );
  AND U11790 ( .A(x[153]), .B(y[738]), .Z(n11520) );
  XOR U11791 ( .A(n11521), .B(n11520), .Z(n11522) );
  XOR U11792 ( .A(n11523), .B(n11522), .Z(n11510) );
  AND U11793 ( .A(x[143]), .B(y[748]), .Z(n11468) );
  AND U11794 ( .A(x[130]), .B(y[761]), .Z(n11467) );
  XOR U11795 ( .A(n11468), .B(n11467), .Z(n11470) );
  AND U11796 ( .A(x[131]), .B(y[760]), .Z(n11469) );
  XOR U11797 ( .A(n11470), .B(n11469), .Z(n11509) );
  XOR U11798 ( .A(n11510), .B(n11509), .Z(n11511) );
  NAND U11799 ( .A(x[144]), .B(y[747]), .Z(n11444) );
  XOR U11800 ( .A(n11444), .B(n11349), .Z(n11447) );
  XOR U11801 ( .A(n11446), .B(n11447), .Z(n11458) );
  AND U11802 ( .A(y[750]), .B(x[141]), .Z(n11351) );
  AND U11803 ( .A(y[751]), .B(x[140]), .Z(n11350) );
  XOR U11804 ( .A(n11351), .B(n11350), .Z(n11457) );
  XNOR U11805 ( .A(n11511), .B(n11512), .Z(n11476) );
  AND U11806 ( .A(n11456), .B(n11352), .Z(n11356) );
  NAND U11807 ( .A(n11354), .B(n11353), .Z(n11355) );
  NANDN U11808 ( .A(n11356), .B(n11355), .Z(n11474) );
  NAND U11809 ( .A(n11358), .B(n11357), .Z(n11362) );
  NAND U11810 ( .A(n11360), .B(n11359), .Z(n11361) );
  NAND U11811 ( .A(n11362), .B(n11361), .Z(n11473) );
  XOR U11812 ( .A(n11474), .B(n11473), .Z(n11475) );
  XOR U11813 ( .A(n11476), .B(n11475), .Z(n11548) );
  XNOR U11814 ( .A(n11547), .B(n11548), .Z(n11550) );
  XNOR U11815 ( .A(n11559), .B(n11560), .Z(n11562) );
  NANDN U11816 ( .A(n11364), .B(n11363), .Z(n11368) );
  NAND U11817 ( .A(n11366), .B(n11365), .Z(n11367) );
  AND U11818 ( .A(n11368), .B(n11367), .Z(n11561) );
  XOR U11819 ( .A(n11562), .B(n11561), .Z(n11426) );
  XNOR U11820 ( .A(n11427), .B(n11426), .Z(n11429) );
  NANDN U11821 ( .A(n11370), .B(n11369), .Z(n11374) );
  NANDN U11822 ( .A(n11372), .B(n11371), .Z(n11373) );
  NAND U11823 ( .A(n11374), .B(n11373), .Z(n11428) );
  XOR U11824 ( .A(n11429), .B(n11428), .Z(n11435) );
  NANDN U11825 ( .A(n11376), .B(n11375), .Z(n11380) );
  NAND U11826 ( .A(n11378), .B(n11377), .Z(n11379) );
  AND U11827 ( .A(n11380), .B(n11379), .Z(n11433) );
  NAND U11828 ( .A(n11382), .B(n11381), .Z(n11386) );
  NAND U11829 ( .A(n11384), .B(n11383), .Z(n11385) );
  NAND U11830 ( .A(n11386), .B(n11385), .Z(n11567) );
  AND U11831 ( .A(n11388), .B(n11387), .Z(n11392) );
  NANDN U11832 ( .A(n11390), .B(n11389), .Z(n11391) );
  NANDN U11833 ( .A(n11392), .B(n11391), .Z(n11498) );
  NANDN U11834 ( .A(n11394), .B(n11393), .Z(n11398) );
  NANDN U11835 ( .A(n11396), .B(n11395), .Z(n11397) );
  NAND U11836 ( .A(n11398), .B(n11397), .Z(n11497) );
  XOR U11837 ( .A(n11498), .B(n11497), .Z(n11499) );
  AND U11838 ( .A(y[756]), .B(x[136]), .Z(n11546) );
  NAND U11839 ( .A(n11399), .B(n11546), .Z(n11403) );
  NAND U11840 ( .A(n11401), .B(n11400), .Z(n11402) );
  NAND U11841 ( .A(n11403), .B(n11402), .Z(n11487) );
  ANDN U11842 ( .B(o[122]), .A(n11404), .Z(n11464) );
  AND U11843 ( .A(x[129]), .B(y[762]), .Z(n11462) );
  AND U11844 ( .A(x[142]), .B(y[749]), .Z(n11461) );
  XOR U11845 ( .A(n11462), .B(n11461), .Z(n11463) );
  XOR U11846 ( .A(n11464), .B(n11463), .Z(n11486) );
  AND U11847 ( .A(x[145]), .B(y[746]), .Z(n11527) );
  AND U11848 ( .A(x[132]), .B(y[759]), .Z(n11526) );
  XOR U11849 ( .A(n11527), .B(n11526), .Z(n11529) );
  AND U11850 ( .A(x[133]), .B(y[758]), .Z(n11528) );
  XOR U11851 ( .A(n11529), .B(n11528), .Z(n11485) );
  XOR U11852 ( .A(n11486), .B(n11485), .Z(n11488) );
  XNOR U11853 ( .A(n11487), .B(n11488), .Z(n11500) );
  NANDN U11854 ( .A(n11406), .B(n11405), .Z(n11410) );
  NANDN U11855 ( .A(n11408), .B(n11407), .Z(n11409) );
  NAND U11856 ( .A(n11410), .B(n11409), .Z(n11505) );
  AND U11857 ( .A(x[135]), .B(y[756]), .Z(n11517) );
  AND U11858 ( .A(y[739]), .B(x[152]), .Z(n11411) );
  XOR U11859 ( .A(n11412), .B(n11411), .Z(n11516) );
  XOR U11860 ( .A(n11517), .B(n11516), .Z(n11504) );
  AND U11861 ( .A(x[150]), .B(y[741]), .Z(n11453) );
  AND U11862 ( .A(x[136]), .B(y[755]), .Z(n11451) );
  AND U11863 ( .A(x[151]), .B(y[740]), .Z(n11450) );
  XOR U11864 ( .A(n11451), .B(n11450), .Z(n11452) );
  XOR U11865 ( .A(n11453), .B(n11452), .Z(n11503) );
  XOR U11866 ( .A(n11504), .B(n11503), .Z(n11506) );
  XNOR U11867 ( .A(n11505), .B(n11506), .Z(n11566) );
  XOR U11868 ( .A(n11567), .B(n11568), .Z(n11439) );
  NANDN U11869 ( .A(n11414), .B(n11413), .Z(n11418) );
  NANDN U11870 ( .A(n11416), .B(n11415), .Z(n11417) );
  NAND U11871 ( .A(n11418), .B(n11417), .Z(n11438) );
  NANDN U11872 ( .A(n11420), .B(n11419), .Z(n11424) );
  NANDN U11873 ( .A(n11422), .B(n11421), .Z(n11423) );
  AND U11874 ( .A(n11424), .B(n11423), .Z(n11440) );
  XOR U11875 ( .A(n11441), .B(n11440), .Z(n11432) );
  XNOR U11876 ( .A(n11433), .B(n11432), .Z(n11434) );
  XNOR U11877 ( .A(n11435), .B(n11434), .Z(n11580) );
  XOR U11878 ( .A(n11581), .B(n11580), .Z(n11582) );
  XOR U11879 ( .A(n11583), .B(n11582), .Z(n11579) );
  XNOR U11880 ( .A(n11578), .B(n11579), .Z(n11425) );
  XNOR U11881 ( .A(n11577), .B(n11425), .Z(N252) );
  NANDN U11882 ( .A(n11427), .B(n11426), .Z(n11431) );
  NAND U11883 ( .A(n11429), .B(n11428), .Z(n11430) );
  AND U11884 ( .A(n11431), .B(n11430), .Z(n11748) );
  NANDN U11885 ( .A(n11433), .B(n11432), .Z(n11437) );
  NANDN U11886 ( .A(n11435), .B(n11434), .Z(n11436) );
  AND U11887 ( .A(n11437), .B(n11436), .Z(n11747) );
  XNOR U11888 ( .A(n11748), .B(n11747), .Z(n11750) );
  NANDN U11889 ( .A(n11439), .B(n11438), .Z(n11443) );
  NAND U11890 ( .A(n11441), .B(n11440), .Z(n11442) );
  AND U11891 ( .A(n11443), .B(n11442), .Z(n11587) );
  NANDN U11892 ( .A(n11445), .B(n11444), .Z(n11449) );
  NAND U11893 ( .A(n11447), .B(n11446), .Z(n11448) );
  NAND U11894 ( .A(n11449), .B(n11448), .Z(n11686) );
  AND U11895 ( .A(x[135]), .B(y[757]), .Z(n11653) );
  AND U11896 ( .A(x[140]), .B(y[752]), .Z(n11652) );
  XOR U11897 ( .A(n11653), .B(n11652), .Z(n11655) );
  AND U11898 ( .A(x[139]), .B(y[753]), .Z(n11654) );
  XOR U11899 ( .A(n11655), .B(n11654), .Z(n11685) );
  AND U11900 ( .A(x[143]), .B(y[749]), .Z(n11679) );
  AND U11901 ( .A(x[155]), .B(y[737]), .Z(n11669) );
  XOR U11902 ( .A(o[124]), .B(n11669), .Z(n11677) );
  AND U11903 ( .A(x[154]), .B(y[738]), .Z(n11676) );
  XOR U11904 ( .A(n11677), .B(n11676), .Z(n11678) );
  XNOR U11905 ( .A(n11679), .B(n11678), .Z(n11684) );
  XOR U11906 ( .A(n11686), .B(n11687), .Z(n11727) );
  NAND U11907 ( .A(n11451), .B(n11450), .Z(n11455) );
  NAND U11908 ( .A(n11453), .B(n11452), .Z(n11454) );
  NAND U11909 ( .A(n11455), .B(n11454), .Z(n11636) );
  AND U11910 ( .A(x[145]), .B(y[747]), .Z(n11612) );
  AND U11911 ( .A(x[150]), .B(y[742]), .Z(n11611) );
  XOR U11912 ( .A(n11612), .B(n11611), .Z(n11614) );
  AND U11913 ( .A(x[132]), .B(y[760]), .Z(n11613) );
  XOR U11914 ( .A(n11614), .B(n11613), .Z(n11635) );
  AND U11915 ( .A(x[134]), .B(y[758]), .Z(n11844) );
  AND U11916 ( .A(x[147]), .B(y[745]), .Z(n11658) );
  XOR U11917 ( .A(n11844), .B(n11658), .Z(n11660) );
  XOR U11918 ( .A(n11660), .B(n11659), .Z(n11634) );
  XOR U11919 ( .A(n11635), .B(n11634), .Z(n11637) );
  XOR U11920 ( .A(n11636), .B(n11637), .Z(n11726) );
  NAND U11921 ( .A(n11456), .B(n11671), .Z(n11460) );
  NANDN U11922 ( .A(n11458), .B(n11457), .Z(n11459) );
  NAND U11923 ( .A(n11460), .B(n11459), .Z(n11630) );
  NAND U11924 ( .A(n11462), .B(n11461), .Z(n11466) );
  NAND U11925 ( .A(n11464), .B(n11463), .Z(n11465) );
  NAND U11926 ( .A(n11466), .B(n11465), .Z(n11629) );
  NAND U11927 ( .A(n11468), .B(n11467), .Z(n11472) );
  NAND U11928 ( .A(n11470), .B(n11469), .Z(n11471) );
  NAND U11929 ( .A(n11472), .B(n11471), .Z(n11628) );
  XNOR U11930 ( .A(n11629), .B(n11628), .Z(n11631) );
  XNOR U11931 ( .A(n11728), .B(n11729), .Z(n11601) );
  NAND U11932 ( .A(n11474), .B(n11473), .Z(n11478) );
  NAND U11933 ( .A(n11476), .B(n11475), .Z(n11477) );
  NAND U11934 ( .A(n11478), .B(n11477), .Z(n11599) );
  NAND U11935 ( .A(n11480), .B(n11479), .Z(n11484) );
  NANDN U11936 ( .A(n11482), .B(n11481), .Z(n11483) );
  NAND U11937 ( .A(n11484), .B(n11483), .Z(n11704) );
  NAND U11938 ( .A(n11486), .B(n11485), .Z(n11490) );
  NAND U11939 ( .A(n11488), .B(n11487), .Z(n11489) );
  NAND U11940 ( .A(n11490), .B(n11489), .Z(n11703) );
  NAND U11941 ( .A(n11492), .B(n11491), .Z(n11496) );
  NAND U11942 ( .A(n11494), .B(n11493), .Z(n11495) );
  NAND U11943 ( .A(n11496), .B(n11495), .Z(n11702) );
  XNOR U11944 ( .A(n11703), .B(n11702), .Z(n11705) );
  XOR U11945 ( .A(n11599), .B(n11600), .Z(n11602) );
  XOR U11946 ( .A(n11601), .B(n11602), .Z(n11735) );
  NAND U11947 ( .A(n11498), .B(n11497), .Z(n11502) );
  NANDN U11948 ( .A(n11500), .B(n11499), .Z(n11501) );
  NAND U11949 ( .A(n11502), .B(n11501), .Z(n11692) );
  NAND U11950 ( .A(n11504), .B(n11503), .Z(n11508) );
  NAND U11951 ( .A(n11506), .B(n11505), .Z(n11507) );
  NAND U11952 ( .A(n11508), .B(n11507), .Z(n11691) );
  NAND U11953 ( .A(n11510), .B(n11509), .Z(n11514) );
  NANDN U11954 ( .A(n11512), .B(n11511), .Z(n11513) );
  NAND U11955 ( .A(n11514), .B(n11513), .Z(n11690) );
  XOR U11956 ( .A(n11691), .B(n11690), .Z(n11693) );
  XOR U11957 ( .A(n11692), .B(n11693), .Z(n11733) );
  AND U11958 ( .A(x[152]), .B(y[743]), .Z(n12078) );
  NAND U11959 ( .A(n12078), .B(n11515), .Z(n11519) );
  NAND U11960 ( .A(n11517), .B(n11516), .Z(n11518) );
  NAND U11961 ( .A(n11519), .B(n11518), .Z(n11716) );
  AND U11962 ( .A(x[153]), .B(y[739]), .Z(n11648) );
  XOR U11963 ( .A(n11649), .B(n11648), .Z(n11647) );
  AND U11964 ( .A(x[129]), .B(y[763]), .Z(n11646) );
  XOR U11965 ( .A(n11647), .B(n11646), .Z(n11715) );
  AND U11966 ( .A(x[144]), .B(y[748]), .Z(n11641) );
  AND U11967 ( .A(x[152]), .B(y[740]), .Z(n11640) );
  XOR U11968 ( .A(n11641), .B(n11640), .Z(n11643) );
  AND U11969 ( .A(x[130]), .B(y[762]), .Z(n11642) );
  XOR U11970 ( .A(n11643), .B(n11642), .Z(n11714) );
  XOR U11971 ( .A(n11715), .B(n11714), .Z(n11717) );
  XOR U11972 ( .A(n11716), .B(n11717), .Z(n11699) );
  NAND U11973 ( .A(n11521), .B(n11520), .Z(n11525) );
  NAND U11974 ( .A(n11523), .B(n11522), .Z(n11524) );
  NAND U11975 ( .A(n11525), .B(n11524), .Z(n11722) );
  AND U11976 ( .A(x[131]), .B(y[761]), .Z(n11670) );
  XOR U11977 ( .A(n11671), .B(n11670), .Z(n11673) );
  AND U11978 ( .A(x[151]), .B(y[741]), .Z(n11672) );
  XOR U11979 ( .A(n11673), .B(n11672), .Z(n11721) );
  AND U11980 ( .A(x[133]), .B(y[759]), .Z(n11664) );
  AND U11981 ( .A(x[149]), .B(y[743]), .Z(n11663) );
  XOR U11982 ( .A(n11664), .B(n11663), .Z(n11666) );
  AND U11983 ( .A(x[148]), .B(y[744]), .Z(n11665) );
  XOR U11984 ( .A(n11666), .B(n11665), .Z(n11720) );
  XOR U11985 ( .A(n11721), .B(n11720), .Z(n11723) );
  XOR U11986 ( .A(n11722), .B(n11723), .Z(n11697) );
  NAND U11987 ( .A(n11527), .B(n11526), .Z(n11531) );
  NAND U11988 ( .A(n11529), .B(n11528), .Z(n11530) );
  NAND U11989 ( .A(n11531), .B(n11530), .Z(n11709) );
  NAND U11990 ( .A(n11533), .B(n11532), .Z(n11537) );
  NAND U11991 ( .A(n11535), .B(n11534), .Z(n11536) );
  NAND U11992 ( .A(n11537), .B(n11536), .Z(n11708) );
  XOR U11993 ( .A(n11709), .B(n11708), .Z(n11711) );
  NAND U11994 ( .A(n11539), .B(n11538), .Z(n11543) );
  NAND U11995 ( .A(n11541), .B(n11540), .Z(n11542) );
  NAND U11996 ( .A(n11543), .B(n11542), .Z(n11607) );
  AND U11997 ( .A(n11544), .B(o[123]), .Z(n11620) );
  AND U11998 ( .A(x[128]), .B(y[764]), .Z(n11618) );
  AND U11999 ( .A(x[156]), .B(y[736]), .Z(n11617) );
  XOR U12000 ( .A(n11618), .B(n11617), .Z(n11619) );
  XOR U12001 ( .A(n11620), .B(n11619), .Z(n11606) );
  NAND U12002 ( .A(y[754]), .B(x[138]), .Z(n11545) );
  XNOR U12003 ( .A(n11546), .B(n11545), .Z(n11625) );
  AND U12004 ( .A(x[137]), .B(y[755]), .Z(n11624) );
  XOR U12005 ( .A(n11625), .B(n11624), .Z(n11605) );
  XOR U12006 ( .A(n11606), .B(n11605), .Z(n11608) );
  XOR U12007 ( .A(n11607), .B(n11608), .Z(n11710) );
  XNOR U12008 ( .A(n11711), .B(n11710), .Z(n11696) );
  XNOR U12009 ( .A(n11735), .B(n11734), .Z(n11740) );
  NAND U12010 ( .A(n11548), .B(n11547), .Z(n11552) );
  NANDN U12011 ( .A(n11550), .B(n11549), .Z(n11551) );
  NAND U12012 ( .A(n11552), .B(n11551), .Z(n11739) );
  NAND U12013 ( .A(n11554), .B(n11553), .Z(n11558) );
  NAND U12014 ( .A(n11556), .B(n11555), .Z(n11557) );
  NAND U12015 ( .A(n11558), .B(n11557), .Z(n11738) );
  XNOR U12016 ( .A(n11739), .B(n11738), .Z(n11741) );
  XNOR U12017 ( .A(n11587), .B(n11588), .Z(n11589) );
  NANDN U12018 ( .A(n11560), .B(n11559), .Z(n11564) );
  NAND U12019 ( .A(n11562), .B(n11561), .Z(n11563) );
  NAND U12020 ( .A(n11564), .B(n11563), .Z(n11595) );
  NANDN U12021 ( .A(n11566), .B(n11565), .Z(n11570) );
  NAND U12022 ( .A(n11568), .B(n11567), .Z(n11569) );
  NAND U12023 ( .A(n11570), .B(n11569), .Z(n11593) );
  NAND U12024 ( .A(n11572), .B(n11571), .Z(n11576) );
  NANDN U12025 ( .A(n11574), .B(n11573), .Z(n11575) );
  AND U12026 ( .A(n11576), .B(n11575), .Z(n11594) );
  XNOR U12027 ( .A(n11593), .B(n11594), .Z(n11596) );
  XNOR U12028 ( .A(n11589), .B(n11590), .Z(n11749) );
  XNOR U12029 ( .A(n11750), .B(n11749), .Z(n11746) );
  NAND U12030 ( .A(n11581), .B(n11580), .Z(n11585) );
  NAND U12031 ( .A(n11583), .B(n11582), .Z(n11584) );
  AND U12032 ( .A(n11585), .B(n11584), .Z(n11745) );
  XOR U12033 ( .A(n11744), .B(n11745), .Z(n11586) );
  XNOR U12034 ( .A(n11746), .B(n11586), .Z(N253) );
  NANDN U12035 ( .A(n11588), .B(n11587), .Z(n11592) );
  NANDN U12036 ( .A(n11590), .B(n11589), .Z(n11591) );
  NAND U12037 ( .A(n11592), .B(n11591), .Z(n11763) );
  NAND U12038 ( .A(n11594), .B(n11593), .Z(n11598) );
  NANDN U12039 ( .A(n11596), .B(n11595), .Z(n11597) );
  NAND U12040 ( .A(n11598), .B(n11597), .Z(n11762) );
  NANDN U12041 ( .A(n11600), .B(n11599), .Z(n11604) );
  NANDN U12042 ( .A(n11602), .B(n11601), .Z(n11603) );
  NAND U12043 ( .A(n11604), .B(n11603), .Z(n11779) );
  NAND U12044 ( .A(n11606), .B(n11605), .Z(n11610) );
  NAND U12045 ( .A(n11608), .B(n11607), .Z(n11609) );
  AND U12046 ( .A(n11610), .B(n11609), .Z(n11888) );
  NAND U12047 ( .A(n11612), .B(n11611), .Z(n11616) );
  NAND U12048 ( .A(n11614), .B(n11613), .Z(n11615) );
  NAND U12049 ( .A(n11616), .B(n11615), .Z(n11928) );
  NAND U12050 ( .A(n11618), .B(n11617), .Z(n11622) );
  NAND U12051 ( .A(n11620), .B(n11619), .Z(n11621) );
  NAND U12052 ( .A(n11622), .B(n11621), .Z(n11927) );
  XOR U12053 ( .A(n11928), .B(n11927), .Z(n11929) );
  AND U12054 ( .A(y[756]), .B(x[138]), .Z(n11925) );
  NAND U12055 ( .A(n11623), .B(n11925), .Z(n11627) );
  NAND U12056 ( .A(n11625), .B(n11624), .Z(n11626) );
  NAND U12057 ( .A(n11627), .B(n11626), .Z(n11896) );
  AND U12058 ( .A(x[150]), .B(y[743]), .Z(n11865) );
  AND U12059 ( .A(x[129]), .B(y[764]), .Z(n11863) );
  AND U12060 ( .A(x[140]), .B(y[753]), .Z(n11998) );
  XOR U12061 ( .A(n11863), .B(n11998), .Z(n11864) );
  XOR U12062 ( .A(n11865), .B(n11864), .Z(n11895) );
  AND U12063 ( .A(x[143]), .B(y[750]), .Z(n11868) );
  XOR U12064 ( .A(n12033), .B(n11868), .Z(n11869) );
  XOR U12065 ( .A(n11895), .B(n11894), .Z(n11897) );
  XNOR U12066 ( .A(n11896), .B(n11897), .Z(n11930) );
  NAND U12067 ( .A(n11629), .B(n11628), .Z(n11633) );
  NANDN U12068 ( .A(n11631), .B(n11630), .Z(n11632) );
  AND U12069 ( .A(n11633), .B(n11632), .Z(n11890) );
  XOR U12070 ( .A(n11891), .B(n11890), .Z(n11885) );
  NAND U12071 ( .A(n11635), .B(n11634), .Z(n11639) );
  NAND U12072 ( .A(n11637), .B(n11636), .Z(n11638) );
  NAND U12073 ( .A(n11639), .B(n11638), .Z(n11883) );
  NAND U12074 ( .A(n11641), .B(n11640), .Z(n11645) );
  NAND U12075 ( .A(n11643), .B(n11642), .Z(n11644) );
  NAND U12076 ( .A(n11645), .B(n11644), .Z(n11901) );
  AND U12077 ( .A(n11647), .B(n11646), .Z(n11651) );
  NAND U12078 ( .A(n11649), .B(n11648), .Z(n11650) );
  NANDN U12079 ( .A(n11651), .B(n11650), .Z(n11900) );
  XOR U12080 ( .A(n11901), .B(n11900), .Z(n11902) );
  NAND U12081 ( .A(n11653), .B(n11652), .Z(n11657) );
  NAND U12082 ( .A(n11655), .B(n11654), .Z(n11656) );
  NAND U12083 ( .A(n11657), .B(n11656), .Z(n11805) );
  AND U12084 ( .A(x[139]), .B(y[754]), .Z(n11841) );
  AND U12085 ( .A(x[131]), .B(y[762]), .Z(n11839) );
  AND U12086 ( .A(x[145]), .B(y[748]), .Z(n11838) );
  XOR U12087 ( .A(n11839), .B(n11838), .Z(n11840) );
  XOR U12088 ( .A(n11841), .B(n11840), .Z(n11804) );
  AND U12089 ( .A(x[151]), .B(y[742]), .Z(n11835) );
  AND U12090 ( .A(x[141]), .B(y[752]), .Z(n11833) );
  AND U12091 ( .A(x[152]), .B(y[741]), .Z(n11983) );
  XOR U12092 ( .A(n11833), .B(n11983), .Z(n11834) );
  XOR U12093 ( .A(n11835), .B(n11834), .Z(n11803) );
  XOR U12094 ( .A(n11804), .B(n11803), .Z(n11806) );
  XNOR U12095 ( .A(n11805), .B(n11806), .Z(n11903) );
  NAND U12096 ( .A(n11844), .B(n11658), .Z(n11662) );
  NAND U12097 ( .A(n11660), .B(n11659), .Z(n11661) );
  NAND U12098 ( .A(n11662), .B(n11661), .Z(n11909) );
  AND U12099 ( .A(x[156]), .B(y[737]), .Z(n11875) );
  XOR U12100 ( .A(o[125]), .B(n11875), .Z(n11920) );
  AND U12101 ( .A(x[128]), .B(y[765]), .Z(n11918) );
  AND U12102 ( .A(x[157]), .B(y[736]), .Z(n11917) );
  XOR U12103 ( .A(n11918), .B(n11917), .Z(n11919) );
  XOR U12104 ( .A(n11920), .B(n11919), .Z(n11907) );
  AND U12105 ( .A(x[153]), .B(y[740]), .Z(n11860) );
  AND U12106 ( .A(x[154]), .B(y[739]), .Z(n11857) );
  XOR U12107 ( .A(n11858), .B(n11857), .Z(n11859) );
  XOR U12108 ( .A(n11860), .B(n11859), .Z(n11906) );
  XOR U12109 ( .A(n11907), .B(n11906), .Z(n11908) );
  XNOR U12110 ( .A(n11909), .B(n11908), .Z(n11792) );
  NAND U12111 ( .A(n11664), .B(n11663), .Z(n11668) );
  NAND U12112 ( .A(n11666), .B(n11665), .Z(n11667) );
  NAND U12113 ( .A(n11668), .B(n11667), .Z(n11853) );
  AND U12114 ( .A(n11669), .B(o[124]), .Z(n11812) );
  AND U12115 ( .A(x[144]), .B(y[749]), .Z(n11810) );
  AND U12116 ( .A(x[155]), .B(y[738]), .Z(n11809) );
  XOR U12117 ( .A(n11810), .B(n11809), .Z(n11811) );
  XOR U12118 ( .A(n11812), .B(n11811), .Z(n11852) );
  AND U12119 ( .A(x[130]), .B(y[763]), .Z(n11822) );
  XOR U12120 ( .A(n11822), .B(n11821), .Z(n11823) );
  XOR U12121 ( .A(n11824), .B(n11823), .Z(n11851) );
  XOR U12122 ( .A(n11852), .B(n11851), .Z(n11854) );
  XNOR U12123 ( .A(n11853), .B(n11854), .Z(n11791) );
  XOR U12124 ( .A(n11792), .B(n11791), .Z(n11793) );
  NAND U12125 ( .A(n11671), .B(n11670), .Z(n11675) );
  NAND U12126 ( .A(n11673), .B(n11672), .Z(n11674) );
  NAND U12127 ( .A(n11675), .B(n11674), .Z(n11828) );
  NAND U12128 ( .A(n11677), .B(n11676), .Z(n11681) );
  NAND U12129 ( .A(n11679), .B(n11678), .Z(n11680) );
  NAND U12130 ( .A(n11681), .B(n11680), .Z(n11827) );
  XOR U12131 ( .A(n11828), .B(n11827), .Z(n11830) );
  AND U12132 ( .A(x[136]), .B(y[757]), .Z(n11846) );
  AND U12133 ( .A(x[134]), .B(y[759]), .Z(n11683) );
  AND U12134 ( .A(y[758]), .B(x[135]), .Z(n11682) );
  XOR U12135 ( .A(n11683), .B(n11682), .Z(n11845) );
  XOR U12136 ( .A(n11846), .B(n11845), .Z(n11912) );
  AND U12137 ( .A(x[137]), .B(y[756]), .Z(n12052) );
  XOR U12138 ( .A(n11912), .B(n12052), .Z(n11914) );
  AND U12139 ( .A(x[133]), .B(y[760]), .Z(n11818) );
  AND U12140 ( .A(x[132]), .B(y[761]), .Z(n11816) );
  AND U12141 ( .A(x[138]), .B(y[755]), .Z(n11815) );
  XOR U12142 ( .A(n11816), .B(n11815), .Z(n11817) );
  XOR U12143 ( .A(n11818), .B(n11817), .Z(n11913) );
  XOR U12144 ( .A(n11914), .B(n11913), .Z(n11829) );
  XOR U12145 ( .A(n11830), .B(n11829), .Z(n11798) );
  NANDN U12146 ( .A(n11685), .B(n11684), .Z(n11689) );
  NAND U12147 ( .A(n11687), .B(n11686), .Z(n11688) );
  NAND U12148 ( .A(n11689), .B(n11688), .Z(n11797) );
  XNOR U12149 ( .A(n11800), .B(n11799), .Z(n11882) );
  XOR U12150 ( .A(n11883), .B(n11882), .Z(n11884) );
  XOR U12151 ( .A(n11779), .B(n11780), .Z(n11782) );
  NAND U12152 ( .A(n11691), .B(n11690), .Z(n11695) );
  NAND U12153 ( .A(n11693), .B(n11692), .Z(n11694) );
  NAND U12154 ( .A(n11695), .B(n11694), .Z(n11773) );
  NANDN U12155 ( .A(n11697), .B(n11696), .Z(n11701) );
  NANDN U12156 ( .A(n11699), .B(n11698), .Z(n11700) );
  AND U12157 ( .A(n11701), .B(n11700), .Z(n11774) );
  XOR U12158 ( .A(n11773), .B(n11774), .Z(n11776) );
  NAND U12159 ( .A(n11703), .B(n11702), .Z(n11707) );
  NANDN U12160 ( .A(n11705), .B(n11704), .Z(n11706) );
  NAND U12161 ( .A(n11707), .B(n11706), .Z(n11787) );
  NAND U12162 ( .A(n11709), .B(n11708), .Z(n11713) );
  NAND U12163 ( .A(n11711), .B(n11710), .Z(n11712) );
  NAND U12164 ( .A(n11713), .B(n11712), .Z(n11878) );
  NAND U12165 ( .A(n11715), .B(n11714), .Z(n11719) );
  NAND U12166 ( .A(n11717), .B(n11716), .Z(n11718) );
  NAND U12167 ( .A(n11719), .B(n11718), .Z(n11877) );
  NAND U12168 ( .A(n11721), .B(n11720), .Z(n11725) );
  NAND U12169 ( .A(n11723), .B(n11722), .Z(n11724) );
  NAND U12170 ( .A(n11725), .B(n11724), .Z(n11876) );
  XOR U12171 ( .A(n11877), .B(n11876), .Z(n11879) );
  XOR U12172 ( .A(n11878), .B(n11879), .Z(n11786) );
  NANDN U12173 ( .A(n11727), .B(n11726), .Z(n11731) );
  NANDN U12174 ( .A(n11729), .B(n11728), .Z(n11730) );
  NAND U12175 ( .A(n11731), .B(n11730), .Z(n11785) );
  XOR U12176 ( .A(n11786), .B(n11785), .Z(n11788) );
  XOR U12177 ( .A(n11787), .B(n11788), .Z(n11775) );
  XOR U12178 ( .A(n11776), .B(n11775), .Z(n11781) );
  XNOR U12179 ( .A(n11782), .B(n11781), .Z(n11769) );
  NANDN U12180 ( .A(n11733), .B(n11732), .Z(n11737) );
  NAND U12181 ( .A(n11735), .B(n11734), .Z(n11736) );
  NAND U12182 ( .A(n11737), .B(n11736), .Z(n11767) );
  NAND U12183 ( .A(n11739), .B(n11738), .Z(n11743) );
  NANDN U12184 ( .A(n11741), .B(n11740), .Z(n11742) );
  AND U12185 ( .A(n11743), .B(n11742), .Z(n11768) );
  XNOR U12186 ( .A(n11767), .B(n11768), .Z(n11770) );
  XOR U12187 ( .A(n11769), .B(n11770), .Z(n11761) );
  XOR U12188 ( .A(n11762), .B(n11761), .Z(n11764) );
  XOR U12189 ( .A(n11763), .B(n11764), .Z(n11757) );
  NANDN U12190 ( .A(n11748), .B(n11747), .Z(n11752) );
  NAND U12191 ( .A(n11750), .B(n11749), .Z(n11751) );
  AND U12192 ( .A(n11752), .B(n11751), .Z(n11756) );
  IV U12193 ( .A(n11756), .Z(n11754) );
  XOR U12194 ( .A(n11755), .B(n11754), .Z(n11753) );
  XNOR U12195 ( .A(n11757), .B(n11753), .Z(N254) );
  NANDN U12196 ( .A(n11754), .B(n11755), .Z(n11760) );
  NOR U12197 ( .A(n11756), .B(n11755), .Z(n11758) );
  OR U12198 ( .A(n11758), .B(n11757), .Z(n11759) );
  AND U12199 ( .A(n11760), .B(n11759), .Z(n11936) );
  NAND U12200 ( .A(n11762), .B(n11761), .Z(n11766) );
  NAND U12201 ( .A(n11764), .B(n11763), .Z(n11765) );
  AND U12202 ( .A(n11766), .B(n11765), .Z(n11935) );
  XNOR U12203 ( .A(n11936), .B(n11935), .Z(n11934) );
  NAND U12204 ( .A(n11768), .B(n11767), .Z(n11772) );
  NANDN U12205 ( .A(n11770), .B(n11769), .Z(n11771) );
  AND U12206 ( .A(n11772), .B(n11771), .Z(n12220) );
  NAND U12207 ( .A(n11774), .B(n11773), .Z(n11778) );
  NAND U12208 ( .A(n11776), .B(n11775), .Z(n11777) );
  AND U12209 ( .A(n11778), .B(n11777), .Z(n12228) );
  NAND U12210 ( .A(n11780), .B(n11779), .Z(n11784) );
  NAND U12211 ( .A(n11782), .B(n11781), .Z(n11783) );
  AND U12212 ( .A(n11784), .B(n11783), .Z(n12227) );
  XOR U12213 ( .A(n12228), .B(n12227), .Z(n12226) );
  NAND U12214 ( .A(n11786), .B(n11785), .Z(n11790) );
  NAND U12215 ( .A(n11788), .B(n11787), .Z(n11789) );
  AND U12216 ( .A(n11790), .B(n11789), .Z(n12225) );
  XOR U12217 ( .A(n12226), .B(n12225), .Z(n12222) );
  NAND U12218 ( .A(n11792), .B(n11791), .Z(n11796) );
  NANDN U12219 ( .A(n11794), .B(n11793), .Z(n11795) );
  AND U12220 ( .A(n11796), .B(n11795), .Z(n12207) );
  NANDN U12221 ( .A(n11798), .B(n11797), .Z(n11802) );
  NAND U12222 ( .A(n11800), .B(n11799), .Z(n11801) );
  AND U12223 ( .A(n11802), .B(n11801), .Z(n12199) );
  NAND U12224 ( .A(n11804), .B(n11803), .Z(n11808) );
  NAND U12225 ( .A(n11806), .B(n11805), .Z(n11807) );
  AND U12226 ( .A(n11808), .B(n11807), .Z(n12183) );
  NAND U12227 ( .A(n11810), .B(n11809), .Z(n11814) );
  NAND U12228 ( .A(n11812), .B(n11811), .Z(n11813) );
  NAND U12229 ( .A(n11814), .B(n11813), .Z(n12141) );
  NAND U12230 ( .A(n11816), .B(n11815), .Z(n11820) );
  NAND U12231 ( .A(n11818), .B(n11817), .Z(n11819) );
  NAND U12232 ( .A(n11820), .B(n11819), .Z(n12144) );
  AND U12233 ( .A(x[134]), .B(y[760]), .Z(n11991) );
  AND U12234 ( .A(x[133]), .B(y[761]), .Z(n11989) );
  AND U12235 ( .A(x[147]), .B(y[747]), .Z(n11988) );
  XOR U12236 ( .A(n11989), .B(n11988), .Z(n11990) );
  XNOR U12237 ( .A(n11991), .B(n11990), .Z(n11971) );
  AND U12238 ( .A(x[132]), .B(y[762]), .Z(n12041) );
  AND U12239 ( .A(x[131]), .B(y[763]), .Z(n12039) );
  AND U12240 ( .A(x[146]), .B(y[748]), .Z(n12038) );
  XOR U12241 ( .A(n12039), .B(n12038), .Z(n12040) );
  XOR U12242 ( .A(n12041), .B(n12040), .Z(n11974) );
  NAND U12243 ( .A(n11822), .B(n11821), .Z(n11826) );
  NAND U12244 ( .A(n11824), .B(n11823), .Z(n11825) );
  AND U12245 ( .A(n11826), .B(n11825), .Z(n11973) );
  XOR U12246 ( .A(n11971), .B(n11972), .Z(n12143) );
  XOR U12247 ( .A(n12144), .B(n12143), .Z(n12142) );
  XOR U12248 ( .A(n12141), .B(n12142), .Z(n12184) );
  NAND U12249 ( .A(n11828), .B(n11827), .Z(n11832) );
  NAND U12250 ( .A(n11830), .B(n11829), .Z(n11831) );
  AND U12251 ( .A(n11832), .B(n11831), .Z(n12181) );
  XOR U12252 ( .A(n12182), .B(n12181), .Z(n12202) );
  NAND U12253 ( .A(n11833), .B(n11983), .Z(n11837) );
  NAND U12254 ( .A(n11835), .B(n11834), .Z(n11836) );
  NAND U12255 ( .A(n11837), .B(n11836), .Z(n11948) );
  NAND U12256 ( .A(n11839), .B(n11838), .Z(n11843) );
  NAND U12257 ( .A(n11841), .B(n11840), .Z(n11842) );
  AND U12258 ( .A(n11843), .B(n11842), .Z(n11952) );
  AND U12259 ( .A(x[128]), .B(y[766]), .Z(n12070) );
  AND U12260 ( .A(x[157]), .B(y[737]), .Z(n12075) );
  XOR U12261 ( .A(o[126]), .B(n12075), .Z(n12072) );
  AND U12262 ( .A(x[158]), .B(y[736]), .Z(n12071) );
  XOR U12263 ( .A(n12072), .B(n12071), .Z(n12069) );
  XOR U12264 ( .A(n12070), .B(n12069), .Z(n11954) );
  AND U12265 ( .A(x[148]), .B(y[746]), .Z(n12063) );
  XOR U12266 ( .A(n12064), .B(n12063), .Z(n12062) );
  AND U12267 ( .A(x[136]), .B(y[758]), .Z(n12061) );
  XNOR U12268 ( .A(n12062), .B(n12061), .Z(n11953) );
  XNOR U12269 ( .A(n11952), .B(n11951), .Z(n11947) );
  XOR U12270 ( .A(n11948), .B(n11947), .Z(n11945) );
  AND U12271 ( .A(x[135]), .B(y[759]), .Z(n12035) );
  NAND U12272 ( .A(n11844), .B(n12035), .Z(n11848) );
  NAND U12273 ( .A(n11846), .B(n11845), .Z(n11847) );
  AND U12274 ( .A(n11848), .B(n11847), .Z(n11963) );
  AND U12275 ( .A(y[745]), .B(x[149]), .Z(n11850) );
  AND U12276 ( .A(y[744]), .B(x[150]), .Z(n11849) );
  XOR U12277 ( .A(n11850), .B(n11849), .Z(n12034) );
  XOR U12278 ( .A(n12035), .B(n12034), .Z(n11966) );
  AND U12279 ( .A(x[145]), .B(y[749]), .Z(n12056) );
  AND U12280 ( .A(x[130]), .B(y[764]), .Z(n12058) );
  AND U12281 ( .A(x[154]), .B(y[740]), .Z(n12057) );
  XOR U12282 ( .A(n12058), .B(n12057), .Z(n12055) );
  XNOR U12283 ( .A(n12056), .B(n12055), .Z(n11965) );
  XNOR U12284 ( .A(n11963), .B(n11964), .Z(n11946) );
  NAND U12285 ( .A(n11852), .B(n11851), .Z(n11856) );
  NAND U12286 ( .A(n11854), .B(n11853), .Z(n11855) );
  NAND U12287 ( .A(n11856), .B(n11855), .Z(n12177) );
  XOR U12288 ( .A(n12178), .B(n12177), .Z(n12176) );
  AND U12289 ( .A(n11858), .B(n11857), .Z(n11862) );
  NAND U12290 ( .A(n11860), .B(n11859), .Z(n11861) );
  NANDN U12291 ( .A(n11862), .B(n11861), .Z(n12135) );
  NAND U12292 ( .A(n11863), .B(n11998), .Z(n11867) );
  NAND U12293 ( .A(n11865), .B(n11864), .Z(n11866) );
  NAND U12294 ( .A(n11867), .B(n11866), .Z(n12138) );
  NAND U12295 ( .A(n12033), .B(n11868), .Z(n11872) );
  NANDN U12296 ( .A(n11870), .B(n11869), .Z(n11871) );
  AND U12297 ( .A(n11872), .B(n11871), .Z(n11958) );
  AND U12298 ( .A(x[151]), .B(y[743]), .Z(n11985) );
  AND U12299 ( .A(y[742]), .B(x[152]), .Z(n11874) );
  AND U12300 ( .A(y[741]), .B(x[153]), .Z(n11873) );
  XOR U12301 ( .A(n11874), .B(n11873), .Z(n11984) );
  XOR U12302 ( .A(n11985), .B(n11984), .Z(n11960) );
  AND U12303 ( .A(n11875), .B(o[125]), .Z(n12008) );
  AND U12304 ( .A(x[156]), .B(y[738]), .Z(n12010) );
  AND U12305 ( .A(x[144]), .B(y[750]), .Z(n12009) );
  XOR U12306 ( .A(n12010), .B(n12009), .Z(n12007) );
  XNOR U12307 ( .A(n12008), .B(n12007), .Z(n11959) );
  XNOR U12308 ( .A(n11958), .B(n11957), .Z(n12137) );
  XOR U12309 ( .A(n12138), .B(n12137), .Z(n12136) );
  XOR U12310 ( .A(n12135), .B(n12136), .Z(n12175) );
  XOR U12311 ( .A(n12176), .B(n12175), .Z(n12201) );
  XNOR U12312 ( .A(n12199), .B(n12200), .Z(n12209) );
  NAND U12313 ( .A(n11877), .B(n11876), .Z(n11881) );
  NAND U12314 ( .A(n11879), .B(n11878), .Z(n11880) );
  AND U12315 ( .A(n11881), .B(n11880), .Z(n12208) );
  NAND U12316 ( .A(n11883), .B(n11882), .Z(n11887) );
  NANDN U12317 ( .A(n11885), .B(n11884), .Z(n11886) );
  NAND U12318 ( .A(n11887), .B(n11886), .Z(n12195) );
  NANDN U12319 ( .A(n11889), .B(n11888), .Z(n11893) );
  NAND U12320 ( .A(n11891), .B(n11890), .Z(n11892) );
  AND U12321 ( .A(n11893), .B(n11892), .Z(n11940) );
  NAND U12322 ( .A(n11895), .B(n11894), .Z(n11899) );
  NAND U12323 ( .A(n11897), .B(n11896), .Z(n11898) );
  AND U12324 ( .A(n11899), .B(n11898), .Z(n12166) );
  NAND U12325 ( .A(n11901), .B(n11900), .Z(n11905) );
  NANDN U12326 ( .A(n11903), .B(n11902), .Z(n11904) );
  AND U12327 ( .A(n11905), .B(n11904), .Z(n12165) );
  XOR U12328 ( .A(n12166), .B(n12165), .Z(n12164) );
  NAND U12329 ( .A(n11907), .B(n11906), .Z(n11911) );
  NAND U12330 ( .A(n11909), .B(n11908), .Z(n11910) );
  AND U12331 ( .A(n11911), .B(n11910), .Z(n12163) );
  XOR U12332 ( .A(n12164), .B(n12163), .Z(n11942) );
  NAND U12333 ( .A(n11912), .B(n12052), .Z(n11916) );
  NAND U12334 ( .A(n11914), .B(n11913), .Z(n11915) );
  AND U12335 ( .A(n11916), .B(n11915), .Z(n12159) );
  NAND U12336 ( .A(n11918), .B(n11917), .Z(n11922) );
  NAND U12337 ( .A(n11920), .B(n11919), .Z(n11921) );
  NAND U12338 ( .A(n11922), .B(n11921), .Z(n11977) );
  AND U12339 ( .A(y[754]), .B(x[140]), .Z(n11923) );
  XOR U12340 ( .A(n11924), .B(n11923), .Z(n11996) );
  XOR U12341 ( .A(n11997), .B(n11996), .Z(n12051) );
  AND U12342 ( .A(y[757]), .B(x[137]), .Z(n11926) );
  XOR U12343 ( .A(n11926), .B(n11925), .Z(n12050) );
  XOR U12344 ( .A(n12051), .B(n12050), .Z(n11980) );
  AND U12345 ( .A(x[155]), .B(y[739]), .Z(n12004) );
  AND U12346 ( .A(x[129]), .B(y[765]), .Z(n12003) );
  XOR U12347 ( .A(n12004), .B(n12003), .Z(n12001) );
  XOR U12348 ( .A(n12002), .B(n12001), .Z(n11979) );
  XOR U12349 ( .A(n11980), .B(n11979), .Z(n11978) );
  XOR U12350 ( .A(n11977), .B(n11978), .Z(n12160) );
  NAND U12351 ( .A(n11928), .B(n11927), .Z(n11932) );
  NANDN U12352 ( .A(n11930), .B(n11929), .Z(n11931) );
  AND U12353 ( .A(n11932), .B(n11931), .Z(n12157) );
  XNOR U12354 ( .A(n12158), .B(n12157), .Z(n11941) );
  XOR U12355 ( .A(n11940), .B(n11939), .Z(n12196) );
  XNOR U12356 ( .A(n12195), .B(n12196), .Z(n12194) );
  XNOR U12357 ( .A(n12220), .B(n12219), .Z(n11933) );
  XNOR U12358 ( .A(n11934), .B(n11933), .Z(N255) );
  NAND U12359 ( .A(n11934), .B(n11933), .Z(n11938) );
  NANDN U12360 ( .A(n11936), .B(n11935), .Z(n11937) );
  AND U12361 ( .A(n11938), .B(n11937), .Z(n12218) );
  NAND U12362 ( .A(n11940), .B(n11939), .Z(n11944) );
  NANDN U12363 ( .A(n11942), .B(n11941), .Z(n11943) );
  AND U12364 ( .A(n11944), .B(n11943), .Z(n12192) );
  NANDN U12365 ( .A(n11946), .B(n11945), .Z(n11950) );
  NAND U12366 ( .A(n11948), .B(n11947), .Z(n11949) );
  AND U12367 ( .A(n11950), .B(n11949), .Z(n12174) );
  NAND U12368 ( .A(n11952), .B(n11951), .Z(n11956) );
  NANDN U12369 ( .A(n11954), .B(n11953), .Z(n11955) );
  AND U12370 ( .A(n11956), .B(n11955), .Z(n12156) );
  NAND U12371 ( .A(n11958), .B(n11957), .Z(n11962) );
  NANDN U12372 ( .A(n11960), .B(n11959), .Z(n11961) );
  AND U12373 ( .A(n11962), .B(n11961), .Z(n11970) );
  NANDN U12374 ( .A(n11964), .B(n11963), .Z(n11968) );
  NANDN U12375 ( .A(n11966), .B(n11965), .Z(n11967) );
  NAND U12376 ( .A(n11968), .B(n11967), .Z(n11969) );
  XNOR U12377 ( .A(n11970), .B(n11969), .Z(n12154) );
  NANDN U12378 ( .A(n11972), .B(n11971), .Z(n11976) );
  NANDN U12379 ( .A(n11974), .B(n11973), .Z(n11975) );
  AND U12380 ( .A(n11976), .B(n11975), .Z(n12152) );
  NAND U12381 ( .A(n11978), .B(n11977), .Z(n11982) );
  NAND U12382 ( .A(n11980), .B(n11979), .Z(n11981) );
  AND U12383 ( .A(n11982), .B(n11981), .Z(n12134) );
  AND U12384 ( .A(x[153]), .B(y[742]), .Z(n12076) );
  AND U12385 ( .A(n11983), .B(n12076), .Z(n11987) );
  AND U12386 ( .A(n11985), .B(n11984), .Z(n11986) );
  NOR U12387 ( .A(n11987), .B(n11986), .Z(n11995) );
  NAND U12388 ( .A(n11989), .B(n11988), .Z(n11993) );
  NAND U12389 ( .A(n11991), .B(n11990), .Z(n11992) );
  AND U12390 ( .A(n11993), .B(n11992), .Z(n11994) );
  XNOR U12391 ( .A(n11995), .B(n11994), .Z(n12049) );
  NAND U12392 ( .A(n11997), .B(n11996), .Z(n12000) );
  NAND U12393 ( .A(n11998), .B(n12100), .Z(n11999) );
  AND U12394 ( .A(n12000), .B(n11999), .Z(n12032) );
  NAND U12395 ( .A(n12002), .B(n12001), .Z(n12006) );
  NAND U12396 ( .A(n12004), .B(n12003), .Z(n12005) );
  AND U12397 ( .A(n12006), .B(n12005), .Z(n12014) );
  NAND U12398 ( .A(n12008), .B(n12007), .Z(n12012) );
  NAND U12399 ( .A(n12010), .B(n12009), .Z(n12011) );
  NAND U12400 ( .A(n12012), .B(n12011), .Z(n12013) );
  XNOR U12401 ( .A(n12014), .B(n12013), .Z(n12030) );
  AND U12402 ( .A(y[767]), .B(x[128]), .Z(n12016) );
  NAND U12403 ( .A(y[763]), .B(x[132]), .Z(n12015) );
  XNOR U12404 ( .A(n12016), .B(n12015), .Z(n12020) );
  AND U12405 ( .A(y[739]), .B(x[156]), .Z(n12018) );
  NAND U12406 ( .A(y[766]), .B(x[129]), .Z(n12017) );
  XNOR U12407 ( .A(n12018), .B(n12017), .Z(n12019) );
  XOR U12408 ( .A(n12020), .B(n12019), .Z(n12028) );
  AND U12409 ( .A(y[736]), .B(x[159]), .Z(n12022) );
  NAND U12410 ( .A(y[749]), .B(x[146]), .Z(n12021) );
  XNOR U12411 ( .A(n12022), .B(n12021), .Z(n12026) );
  AND U12412 ( .A(y[764]), .B(x[131]), .Z(n12024) );
  NAND U12413 ( .A(y[761]), .B(x[134]), .Z(n12023) );
  XNOR U12414 ( .A(n12024), .B(n12023), .Z(n12025) );
  XNOR U12415 ( .A(n12026), .B(n12025), .Z(n12027) );
  XNOR U12416 ( .A(n12028), .B(n12027), .Z(n12029) );
  XNOR U12417 ( .A(n12030), .B(n12029), .Z(n12031) );
  XNOR U12418 ( .A(n12032), .B(n12031), .Z(n12047) );
  AND U12419 ( .A(x[150]), .B(y[745]), .Z(n12077) );
  AND U12420 ( .A(n12033), .B(n12077), .Z(n12037) );
  AND U12421 ( .A(n12035), .B(n12034), .Z(n12036) );
  NOR U12422 ( .A(n12037), .B(n12036), .Z(n12045) );
  NAND U12423 ( .A(n12039), .B(n12038), .Z(n12043) );
  NAND U12424 ( .A(n12041), .B(n12040), .Z(n12042) );
  AND U12425 ( .A(n12043), .B(n12042), .Z(n12044) );
  XNOR U12426 ( .A(n12045), .B(n12044), .Z(n12046) );
  XNOR U12427 ( .A(n12047), .B(n12046), .Z(n12048) );
  XNOR U12428 ( .A(n12049), .B(n12048), .Z(n12132) );
  NAND U12429 ( .A(n12051), .B(n12050), .Z(n12054) );
  AND U12430 ( .A(x[138]), .B(y[757]), .Z(n12099) );
  NAND U12431 ( .A(n12052), .B(n12099), .Z(n12053) );
  AND U12432 ( .A(n12054), .B(n12053), .Z(n12130) );
  NAND U12433 ( .A(n12056), .B(n12055), .Z(n12060) );
  NAND U12434 ( .A(n12058), .B(n12057), .Z(n12059) );
  AND U12435 ( .A(n12060), .B(n12059), .Z(n12068) );
  NAND U12436 ( .A(n12062), .B(n12061), .Z(n12066) );
  NAND U12437 ( .A(n12064), .B(n12063), .Z(n12065) );
  NAND U12438 ( .A(n12066), .B(n12065), .Z(n12067) );
  XNOR U12439 ( .A(n12068), .B(n12067), .Z(n12128) );
  NAND U12440 ( .A(n12070), .B(n12069), .Z(n12074) );
  NAND U12441 ( .A(n12072), .B(n12071), .Z(n12073) );
  AND U12442 ( .A(n12074), .B(n12073), .Z(n12126) );
  AND U12443 ( .A(y[748]), .B(x[147]), .Z(n12084) );
  AND U12444 ( .A(n12075), .B(o[126]), .Z(n12082) );
  XOR U12445 ( .A(n12076), .B(o[127]), .Z(n12080) );
  XNOR U12446 ( .A(n12078), .B(n12077), .Z(n12079) );
  XNOR U12447 ( .A(n12080), .B(n12079), .Z(n12081) );
  XNOR U12448 ( .A(n12082), .B(n12081), .Z(n12083) );
  XNOR U12449 ( .A(n12084), .B(n12083), .Z(n12124) );
  AND U12450 ( .A(y[765]), .B(x[130]), .Z(n12090) );
  AND U12451 ( .A(y[758]), .B(x[137]), .Z(n12086) );
  NAND U12452 ( .A(y[753]), .B(x[142]), .Z(n12085) );
  XNOR U12453 ( .A(n12086), .B(n12085), .Z(n12087) );
  XNOR U12454 ( .A(n12088), .B(n12087), .Z(n12089) );
  XNOR U12455 ( .A(n12090), .B(n12089), .Z(n12114) );
  AND U12456 ( .A(y[755]), .B(x[140]), .Z(n12092) );
  NAND U12457 ( .A(y[756]), .B(x[139]), .Z(n12091) );
  XNOR U12458 ( .A(n12092), .B(n12091), .Z(n12104) );
  AND U12459 ( .A(y[741]), .B(x[154]), .Z(n12094) );
  NAND U12460 ( .A(y[751]), .B(x[144]), .Z(n12093) );
  XNOR U12461 ( .A(n12094), .B(n12093), .Z(n12098) );
  AND U12462 ( .A(y[738]), .B(x[157]), .Z(n12096) );
  NAND U12463 ( .A(y[747]), .B(x[148]), .Z(n12095) );
  XNOR U12464 ( .A(n12096), .B(n12095), .Z(n12097) );
  XOR U12465 ( .A(n12098), .B(n12097), .Z(n12102) );
  XNOR U12466 ( .A(n12100), .B(n12099), .Z(n12101) );
  XNOR U12467 ( .A(n12102), .B(n12101), .Z(n12103) );
  XOR U12468 ( .A(n12104), .B(n12103), .Z(n12112) );
  AND U12469 ( .A(y[746]), .B(x[149]), .Z(n12106) );
  NAND U12470 ( .A(y[759]), .B(x[136]), .Z(n12105) );
  XNOR U12471 ( .A(n12106), .B(n12105), .Z(n12110) );
  AND U12472 ( .A(y[762]), .B(x[133]), .Z(n12108) );
  NAND U12473 ( .A(y[760]), .B(x[135]), .Z(n12107) );
  XNOR U12474 ( .A(n12108), .B(n12107), .Z(n12109) );
  XNOR U12475 ( .A(n12110), .B(n12109), .Z(n12111) );
  XNOR U12476 ( .A(n12112), .B(n12111), .Z(n12113) );
  XOR U12477 ( .A(n12114), .B(n12113), .Z(n12122) );
  AND U12478 ( .A(y[737]), .B(x[158]), .Z(n12116) );
  NAND U12479 ( .A(y[740]), .B(x[155]), .Z(n12115) );
  XNOR U12480 ( .A(n12116), .B(n12115), .Z(n12120) );
  AND U12481 ( .A(y[750]), .B(x[145]), .Z(n12118) );
  NAND U12482 ( .A(y[744]), .B(x[151]), .Z(n12117) );
  XNOR U12483 ( .A(n12118), .B(n12117), .Z(n12119) );
  XNOR U12484 ( .A(n12120), .B(n12119), .Z(n12121) );
  XNOR U12485 ( .A(n12122), .B(n12121), .Z(n12123) );
  XNOR U12486 ( .A(n12124), .B(n12123), .Z(n12125) );
  XNOR U12487 ( .A(n12126), .B(n12125), .Z(n12127) );
  XNOR U12488 ( .A(n12128), .B(n12127), .Z(n12129) );
  XNOR U12489 ( .A(n12130), .B(n12129), .Z(n12131) );
  XNOR U12490 ( .A(n12132), .B(n12131), .Z(n12133) );
  XNOR U12491 ( .A(n12134), .B(n12133), .Z(n12150) );
  NAND U12492 ( .A(n12136), .B(n12135), .Z(n12140) );
  NAND U12493 ( .A(n12138), .B(n12137), .Z(n12139) );
  AND U12494 ( .A(n12140), .B(n12139), .Z(n12148) );
  NAND U12495 ( .A(n12142), .B(n12141), .Z(n12146) );
  NAND U12496 ( .A(n12144), .B(n12143), .Z(n12145) );
  NAND U12497 ( .A(n12146), .B(n12145), .Z(n12147) );
  XNOR U12498 ( .A(n12148), .B(n12147), .Z(n12149) );
  XNOR U12499 ( .A(n12150), .B(n12149), .Z(n12151) );
  XNOR U12500 ( .A(n12152), .B(n12151), .Z(n12153) );
  XNOR U12501 ( .A(n12154), .B(n12153), .Z(n12155) );
  XNOR U12502 ( .A(n12156), .B(n12155), .Z(n12172) );
  NAND U12503 ( .A(n12158), .B(n12157), .Z(n12162) );
  NANDN U12504 ( .A(n12160), .B(n12159), .Z(n12161) );
  AND U12505 ( .A(n12162), .B(n12161), .Z(n12170) );
  NAND U12506 ( .A(n12164), .B(n12163), .Z(n12168) );
  NAND U12507 ( .A(n12166), .B(n12165), .Z(n12167) );
  NAND U12508 ( .A(n12168), .B(n12167), .Z(n12169) );
  XNOR U12509 ( .A(n12170), .B(n12169), .Z(n12171) );
  XNOR U12510 ( .A(n12172), .B(n12171), .Z(n12173) );
  XNOR U12511 ( .A(n12174), .B(n12173), .Z(n12190) );
  NAND U12512 ( .A(n12176), .B(n12175), .Z(n12180) );
  NAND U12513 ( .A(n12178), .B(n12177), .Z(n12179) );
  AND U12514 ( .A(n12180), .B(n12179), .Z(n12188) );
  NAND U12515 ( .A(n12182), .B(n12181), .Z(n12186) );
  NANDN U12516 ( .A(n12184), .B(n12183), .Z(n12185) );
  NAND U12517 ( .A(n12186), .B(n12185), .Z(n12187) );
  XNOR U12518 ( .A(n12188), .B(n12187), .Z(n12189) );
  XNOR U12519 ( .A(n12190), .B(n12189), .Z(n12191) );
  XNOR U12520 ( .A(n12192), .B(n12191), .Z(n12216) );
  NANDN U12521 ( .A(n12194), .B(n12193), .Z(n12198) );
  NAND U12522 ( .A(n12196), .B(n12195), .Z(n12197) );
  AND U12523 ( .A(n12198), .B(n12197), .Z(n12206) );
  NANDN U12524 ( .A(n12200), .B(n12199), .Z(n12204) );
  NANDN U12525 ( .A(n12202), .B(n12201), .Z(n12203) );
  NAND U12526 ( .A(n12204), .B(n12203), .Z(n12205) );
  XNOR U12527 ( .A(n12206), .B(n12205), .Z(n12214) );
  ANDN U12528 ( .B(n12208), .A(n12207), .Z(n12210) );
  NANDN U12529 ( .A(n12210), .B(n12209), .Z(n12211) );
  NAND U12530 ( .A(n12212), .B(n12211), .Z(n12213) );
  XNOR U12531 ( .A(n12214), .B(n12213), .Z(n12215) );
  XNOR U12532 ( .A(n12216), .B(n12215), .Z(n12217) );
  XNOR U12533 ( .A(n12218), .B(n12217), .Z(n12234) );
  NAND U12534 ( .A(n12220), .B(n12219), .Z(n12224) );
  NANDN U12535 ( .A(n12222), .B(n12221), .Z(n12223) );
  AND U12536 ( .A(n12224), .B(n12223), .Z(n12232) );
  NAND U12537 ( .A(n12226), .B(n12225), .Z(n12230) );
  NAND U12538 ( .A(n12228), .B(n12227), .Z(n12229) );
  NAND U12539 ( .A(n12230), .B(n12229), .Z(n12231) );
  XNOR U12540 ( .A(n12232), .B(n12231), .Z(n12233) );
  XNOR U12541 ( .A(n12234), .B(n12233), .Z(N256) );
  AND U12542 ( .A(x[128]), .B(y[768]), .Z(n12891) );
  XOR U12543 ( .A(n12891), .B(o[128]), .Z(N289) );
  AND U12544 ( .A(x[129]), .B(y[768]), .Z(n12243) );
  AND U12545 ( .A(x[128]), .B(y[769]), .Z(n12242) );
  XNOR U12546 ( .A(n12242), .B(o[129]), .Z(n12235) );
  XNOR U12547 ( .A(n12243), .B(n12235), .Z(n12237) );
  NAND U12548 ( .A(n12891), .B(o[128]), .Z(n12236) );
  XNOR U12549 ( .A(n12237), .B(n12236), .Z(N290) );
  NANDN U12550 ( .A(n12243), .B(n12235), .Z(n12239) );
  NAND U12551 ( .A(n12237), .B(n12236), .Z(n12238) );
  AND U12552 ( .A(n12239), .B(n12238), .Z(n12249) );
  AND U12553 ( .A(x[128]), .B(y[770]), .Z(n12256) );
  XNOR U12554 ( .A(n12256), .B(o[130]), .Z(n12248) );
  XNOR U12555 ( .A(n12249), .B(n12248), .Z(n12251) );
  AND U12556 ( .A(y[769]), .B(x[129]), .Z(n12241) );
  NAND U12557 ( .A(y[768]), .B(x[130]), .Z(n12240) );
  XNOR U12558 ( .A(n12241), .B(n12240), .Z(n12245) );
  AND U12559 ( .A(n12242), .B(o[129]), .Z(n12244) );
  XNOR U12560 ( .A(n12245), .B(n12244), .Z(n12250) );
  XNOR U12561 ( .A(n12251), .B(n12250), .Z(N291) );
  AND U12562 ( .A(x[130]), .B(y[769]), .Z(n12263) );
  NAND U12563 ( .A(n12263), .B(n12243), .Z(n12247) );
  NAND U12564 ( .A(n12245), .B(n12244), .Z(n12246) );
  AND U12565 ( .A(n12247), .B(n12246), .Z(n12266) );
  NANDN U12566 ( .A(n12249), .B(n12248), .Z(n12253) );
  NAND U12567 ( .A(n12251), .B(n12250), .Z(n12252) );
  AND U12568 ( .A(n12253), .B(n12252), .Z(n12265) );
  XNOR U12569 ( .A(n12266), .B(n12265), .Z(n12268) );
  AND U12570 ( .A(x[129]), .B(y[770]), .Z(n12372) );
  XOR U12571 ( .A(n12263), .B(o[131]), .Z(n12271) );
  XOR U12572 ( .A(n12372), .B(n12271), .Z(n12273) );
  AND U12573 ( .A(y[771]), .B(x[128]), .Z(n12255) );
  NAND U12574 ( .A(y[768]), .B(x[131]), .Z(n12254) );
  XNOR U12575 ( .A(n12255), .B(n12254), .Z(n12258) );
  AND U12576 ( .A(n12256), .B(o[130]), .Z(n12257) );
  XOR U12577 ( .A(n12258), .B(n12257), .Z(n12272) );
  XOR U12578 ( .A(n12273), .B(n12272), .Z(n12267) );
  XOR U12579 ( .A(n12268), .B(n12267), .Z(N292) );
  AND U12580 ( .A(x[131]), .B(y[771]), .Z(n12316) );
  NAND U12581 ( .A(n12891), .B(n12316), .Z(n12260) );
  NAND U12582 ( .A(n12258), .B(n12257), .Z(n12259) );
  AND U12583 ( .A(n12260), .B(n12259), .Z(n12294) );
  AND U12584 ( .A(y[772]), .B(x[128]), .Z(n12262) );
  NAND U12585 ( .A(y[768]), .B(x[132]), .Z(n12261) );
  XNOR U12586 ( .A(n12262), .B(n12261), .Z(n12287) );
  NAND U12587 ( .A(n12263), .B(o[131]), .Z(n12288) );
  AND U12588 ( .A(y[771]), .B(x[129]), .Z(n12479) );
  NAND U12589 ( .A(y[770]), .B(x[130]), .Z(n12264) );
  XNOR U12590 ( .A(n12479), .B(n12264), .Z(n12284) );
  NAND U12591 ( .A(x[131]), .B(y[769]), .Z(n12279) );
  XOR U12592 ( .A(n12284), .B(n12283), .Z(n12291) );
  XOR U12593 ( .A(n12292), .B(n12291), .Z(n12293) );
  XNOR U12594 ( .A(n12294), .B(n12293), .Z(n12298) );
  NANDN U12595 ( .A(n12266), .B(n12265), .Z(n12270) );
  NAND U12596 ( .A(n12268), .B(n12267), .Z(n12269) );
  NAND U12597 ( .A(n12270), .B(n12269), .Z(n12299) );
  NAND U12598 ( .A(n12372), .B(n12271), .Z(n12275) );
  NAND U12599 ( .A(n12273), .B(n12272), .Z(n12274) );
  NAND U12600 ( .A(n12275), .B(n12274), .Z(n12300) );
  IV U12601 ( .A(n12300), .Z(n12297) );
  XOR U12602 ( .A(n12299), .B(n12297), .Z(n12276) );
  XNOR U12603 ( .A(n12298), .B(n12276), .Z(N293) );
  AND U12604 ( .A(y[773]), .B(x[128]), .Z(n12278) );
  NAND U12605 ( .A(y[768]), .B(x[133]), .Z(n12277) );
  XNOR U12606 ( .A(n12278), .B(n12277), .Z(n12309) );
  ANDN U12607 ( .B(o[132]), .A(n12279), .Z(n12308) );
  XOR U12608 ( .A(n12309), .B(n12308), .Z(n12307) );
  NAND U12609 ( .A(x[130]), .B(y[771]), .Z(n12380) );
  AND U12610 ( .A(y[772]), .B(x[129]), .Z(n12281) );
  NAND U12611 ( .A(y[770]), .B(x[131]), .Z(n12280) );
  XNOR U12612 ( .A(n12281), .B(n12280), .Z(n12303) );
  AND U12613 ( .A(x[132]), .B(y[769]), .Z(n12314) );
  XOR U12614 ( .A(n12314), .B(o[133]), .Z(n12302) );
  XOR U12615 ( .A(n12303), .B(n12302), .Z(n12306) );
  XOR U12616 ( .A(n12380), .B(n12306), .Z(n12282) );
  XNOR U12617 ( .A(n12307), .B(n12282), .Z(n12324) );
  NANDN U12618 ( .A(n12380), .B(n12372), .Z(n12286) );
  NAND U12619 ( .A(n12284), .B(n12283), .Z(n12285) );
  AND U12620 ( .A(n12286), .B(n12285), .Z(n12322) );
  AND U12621 ( .A(x[132]), .B(y[772]), .Z(n13118) );
  NAND U12622 ( .A(n13118), .B(n12891), .Z(n12290) );
  NANDN U12623 ( .A(n12288), .B(n12287), .Z(n12289) );
  NAND U12624 ( .A(n12290), .B(n12289), .Z(n12321) );
  XNOR U12625 ( .A(n12324), .B(n12323), .Z(n12320) );
  NAND U12626 ( .A(n12292), .B(n12291), .Z(n12296) );
  NANDN U12627 ( .A(n12294), .B(n12293), .Z(n12295) );
  NAND U12628 ( .A(n12296), .B(n12295), .Z(n12319) );
  XOR U12629 ( .A(n12319), .B(n12318), .Z(n12301) );
  XNOR U12630 ( .A(n12320), .B(n12301), .Z(N294) );
  AND U12631 ( .A(x[131]), .B(y[772]), .Z(n12381) );
  NAND U12632 ( .A(n12381), .B(n12372), .Z(n12305) );
  NAND U12633 ( .A(n12303), .B(n12302), .Z(n12304) );
  AND U12634 ( .A(n12305), .B(n12304), .Z(n12329) );
  AND U12635 ( .A(x[133]), .B(y[773]), .Z(n12559) );
  NAND U12636 ( .A(n12891), .B(n12559), .Z(n12311) );
  NAND U12637 ( .A(n12309), .B(n12308), .Z(n12310) );
  NAND U12638 ( .A(n12311), .B(n12310), .Z(n12341) );
  AND U12639 ( .A(y[774]), .B(x[128]), .Z(n12313) );
  NAND U12640 ( .A(y[768]), .B(x[134]), .Z(n12312) );
  XNOR U12641 ( .A(n12313), .B(n12312), .Z(n12348) );
  NAND U12642 ( .A(n12314), .B(o[133]), .Z(n12349) );
  XNOR U12643 ( .A(n12348), .B(n12349), .Z(n12342) );
  XOR U12644 ( .A(n12341), .B(n12342), .Z(n12344) );
  NAND U12645 ( .A(y[772]), .B(x[130]), .Z(n12315) );
  XNOR U12646 ( .A(n12316), .B(n12315), .Z(n12353) );
  AND U12647 ( .A(y[773]), .B(x[129]), .Z(n12589) );
  NAND U12648 ( .A(y[770]), .B(x[132]), .Z(n12317) );
  XNOR U12649 ( .A(n12589), .B(n12317), .Z(n12357) );
  AND U12650 ( .A(x[133]), .B(y[769]), .Z(n12364) );
  XOR U12651 ( .A(n12364), .B(o[134]), .Z(n12356) );
  XOR U12652 ( .A(n12357), .B(n12356), .Z(n12352) );
  XOR U12653 ( .A(n12353), .B(n12352), .Z(n12343) );
  XOR U12654 ( .A(n12344), .B(n12343), .Z(n12330) );
  XNOR U12655 ( .A(n12331), .B(n12330), .Z(n12337) );
  NANDN U12656 ( .A(n12322), .B(n12321), .Z(n12326) );
  NAND U12657 ( .A(n12324), .B(n12323), .Z(n12325) );
  NAND U12658 ( .A(n12326), .B(n12325), .Z(n12335) );
  IV U12659 ( .A(n12335), .Z(n12334) );
  XOR U12660 ( .A(n12336), .B(n12334), .Z(n12327) );
  XNOR U12661 ( .A(n12337), .B(n12327), .Z(N295) );
  NANDN U12662 ( .A(n12329), .B(n12328), .Z(n12333) );
  NAND U12663 ( .A(n12331), .B(n12330), .Z(n12332) );
  NAND U12664 ( .A(n12333), .B(n12332), .Z(n12399) );
  IV U12665 ( .A(n12399), .Z(n12398) );
  OR U12666 ( .A(n12336), .B(n12334), .Z(n12340) );
  ANDN U12667 ( .B(n12336), .A(n12335), .Z(n12338) );
  OR U12668 ( .A(n12338), .B(n12337), .Z(n12339) );
  AND U12669 ( .A(n12340), .B(n12339), .Z(n12400) );
  NAND U12670 ( .A(n12342), .B(n12341), .Z(n12346) );
  NAND U12671 ( .A(n12344), .B(n12343), .Z(n12345) );
  AND U12672 ( .A(n12346), .B(n12345), .Z(n12408) );
  AND U12673 ( .A(y[770]), .B(x[133]), .Z(n12467) );
  NAND U12674 ( .A(y[774]), .B(x[129]), .Z(n12347) );
  XNOR U12675 ( .A(n12467), .B(n12347), .Z(n12374) );
  NAND U12676 ( .A(x[134]), .B(y[769]), .Z(n12377) );
  XNOR U12677 ( .A(o[135]), .B(n12377), .Z(n12373) );
  XOR U12678 ( .A(n12374), .B(n12373), .Z(n12393) );
  AND U12679 ( .A(x[134]), .B(y[774]), .Z(n12426) );
  NAND U12680 ( .A(n12891), .B(n12426), .Z(n12351) );
  NANDN U12681 ( .A(n12349), .B(n12348), .Z(n12350) );
  AND U12682 ( .A(n12351), .B(n12350), .Z(n12392) );
  XNOR U12683 ( .A(n12393), .B(n12392), .Z(n12394) );
  NANDN U12684 ( .A(n12380), .B(n12381), .Z(n12355) );
  NAND U12685 ( .A(n12353), .B(n12352), .Z(n12354) );
  NAND U12686 ( .A(n12355), .B(n12354), .Z(n12395) );
  XNOR U12687 ( .A(n12394), .B(n12395), .Z(n12406) );
  AND U12688 ( .A(x[132]), .B(y[773]), .Z(n12896) );
  NAND U12689 ( .A(n12896), .B(n12372), .Z(n12359) );
  NAND U12690 ( .A(n12357), .B(n12356), .Z(n12358) );
  AND U12691 ( .A(n12359), .B(n12358), .Z(n12369) );
  AND U12692 ( .A(y[773]), .B(x[130]), .Z(n12361) );
  NAND U12693 ( .A(y[771]), .B(x[132]), .Z(n12360) );
  XNOR U12694 ( .A(n12361), .B(n12360), .Z(n12382) );
  XOR U12695 ( .A(n12382), .B(n12381), .Z(n12367) );
  AND U12696 ( .A(y[775]), .B(x[128]), .Z(n12363) );
  NAND U12697 ( .A(y[768]), .B(x[135]), .Z(n12362) );
  XNOR U12698 ( .A(n12363), .B(n12362), .Z(n12387) );
  AND U12699 ( .A(n12364), .B(o[134]), .Z(n12386) );
  XNOR U12700 ( .A(n12387), .B(n12386), .Z(n12366) );
  XNOR U12701 ( .A(n12367), .B(n12366), .Z(n12368) );
  XOR U12702 ( .A(n12369), .B(n12368), .Z(n12405) );
  XOR U12703 ( .A(n12406), .B(n12405), .Z(n12407) );
  XOR U12704 ( .A(n12408), .B(n12407), .Z(n12401) );
  XNOR U12705 ( .A(n12400), .B(n12401), .Z(n12365) );
  XOR U12706 ( .A(n12398), .B(n12365), .Z(N296) );
  NANDN U12707 ( .A(n12367), .B(n12366), .Z(n12371) );
  NAND U12708 ( .A(n12369), .B(n12368), .Z(n12370) );
  AND U12709 ( .A(n12371), .B(n12370), .Z(n12457) );
  AND U12710 ( .A(x[133]), .B(y[774]), .Z(n12551) );
  NAND U12711 ( .A(n12551), .B(n12372), .Z(n12376) );
  NAND U12712 ( .A(n12374), .B(n12373), .Z(n12375) );
  NAND U12713 ( .A(n12376), .B(n12375), .Z(n12455) );
  ANDN U12714 ( .B(o[135]), .A(n12377), .Z(n12445) );
  AND U12715 ( .A(y[771]), .B(x[133]), .Z(n12996) );
  NAND U12716 ( .A(y[775]), .B(x[129]), .Z(n12378) );
  XNOR U12717 ( .A(n12996), .B(n12378), .Z(n12444) );
  XOR U12718 ( .A(n12445), .B(n12444), .Z(n12432) );
  NAND U12719 ( .A(x[131]), .B(y[773]), .Z(n13232) );
  AND U12720 ( .A(y[774]), .B(x[130]), .Z(n13314) );
  NAND U12721 ( .A(y[770]), .B(x[134]), .Z(n12379) );
  XNOR U12722 ( .A(n13314), .B(n12379), .Z(n12427) );
  XNOR U12723 ( .A(n13118), .B(n12427), .Z(n12430) );
  XOR U12724 ( .A(n13232), .B(n12430), .Z(n12431) );
  XOR U12725 ( .A(n12432), .B(n12431), .Z(n12454) );
  XOR U12726 ( .A(n12455), .B(n12454), .Z(n12456) );
  XOR U12727 ( .A(n12457), .B(n12456), .Z(n12415) );
  NANDN U12728 ( .A(n12380), .B(n12896), .Z(n12384) );
  NAND U12729 ( .A(n12382), .B(n12381), .Z(n12383) );
  NAND U12730 ( .A(n12384), .B(n12383), .Z(n12450) );
  AND U12731 ( .A(x[135]), .B(y[775]), .Z(n12385) );
  NAND U12732 ( .A(n12891), .B(n12385), .Z(n12389) );
  NAND U12733 ( .A(n12387), .B(n12386), .Z(n12388) );
  NAND U12734 ( .A(n12389), .B(n12388), .Z(n12448) );
  AND U12735 ( .A(y[776]), .B(x[128]), .Z(n12391) );
  NAND U12736 ( .A(y[768]), .B(x[136]), .Z(n12390) );
  XNOR U12737 ( .A(n12391), .B(n12390), .Z(n12435) );
  NAND U12738 ( .A(x[135]), .B(y[769]), .Z(n12438) );
  XNOR U12739 ( .A(o[136]), .B(n12438), .Z(n12434) );
  XOR U12740 ( .A(n12435), .B(n12434), .Z(n12449) );
  XNOR U12741 ( .A(n12448), .B(n12449), .Z(n12451) );
  NANDN U12742 ( .A(n12393), .B(n12392), .Z(n12397) );
  NANDN U12743 ( .A(n12395), .B(n12394), .Z(n12396) );
  NAND U12744 ( .A(n12397), .B(n12396), .Z(n12412) );
  XOR U12745 ( .A(n12413), .B(n12412), .Z(n12414) );
  XNOR U12746 ( .A(n12415), .B(n12414), .Z(n12421) );
  OR U12747 ( .A(n12400), .B(n12398), .Z(n12404) );
  ANDN U12748 ( .B(n12400), .A(n12399), .Z(n12402) );
  OR U12749 ( .A(n12402), .B(n12401), .Z(n12403) );
  AND U12750 ( .A(n12404), .B(n12403), .Z(n12420) );
  NAND U12751 ( .A(n12406), .B(n12405), .Z(n12410) );
  NAND U12752 ( .A(n12408), .B(n12407), .Z(n12409) );
  AND U12753 ( .A(n12410), .B(n12409), .Z(n12419) );
  IV U12754 ( .A(n12419), .Z(n12418) );
  XOR U12755 ( .A(n12420), .B(n12418), .Z(n12411) );
  XNOR U12756 ( .A(n12421), .B(n12411), .Z(N297) );
  NAND U12757 ( .A(n12413), .B(n12412), .Z(n12417) );
  NANDN U12758 ( .A(n12415), .B(n12414), .Z(n12416) );
  NAND U12759 ( .A(n12417), .B(n12416), .Z(n12505) );
  IV U12760 ( .A(n12505), .Z(n12503) );
  OR U12761 ( .A(n12420), .B(n12418), .Z(n12424) );
  ANDN U12762 ( .B(n12420), .A(n12419), .Z(n12422) );
  OR U12763 ( .A(n12422), .B(n12421), .Z(n12423) );
  AND U12764 ( .A(n12424), .B(n12423), .Z(n12504) );
  AND U12765 ( .A(x[130]), .B(y[770]), .Z(n12425) );
  NAND U12766 ( .A(n12426), .B(n12425), .Z(n12429) );
  NAND U12767 ( .A(n13118), .B(n12427), .Z(n12428) );
  AND U12768 ( .A(n12429), .B(n12428), .Z(n12462) );
  XNOR U12769 ( .A(n12462), .B(n12461), .Z(n12464) );
  AND U12770 ( .A(x[136]), .B(y[776]), .Z(n12433) );
  NAND U12771 ( .A(n12433), .B(n12891), .Z(n12437) );
  NAND U12772 ( .A(n12435), .B(n12434), .Z(n12436) );
  AND U12773 ( .A(n12437), .B(n12436), .Z(n12496) );
  ANDN U12774 ( .B(o[136]), .A(n12438), .Z(n12470) );
  AND U12775 ( .A(y[772]), .B(x[133]), .Z(n12440) );
  NAND U12776 ( .A(y[770]), .B(x[135]), .Z(n12439) );
  XNOR U12777 ( .A(n12440), .B(n12439), .Z(n12469) );
  XOR U12778 ( .A(n12470), .B(n12469), .Z(n12494) );
  AND U12779 ( .A(y[768]), .B(x[137]), .Z(n12442) );
  NAND U12780 ( .A(y[777]), .B(x[128]), .Z(n12441) );
  XNOR U12781 ( .A(n12442), .B(n12441), .Z(n12476) );
  NAND U12782 ( .A(x[136]), .B(y[769]), .Z(n12485) );
  XNOR U12783 ( .A(o[137]), .B(n12485), .Z(n12475) );
  XNOR U12784 ( .A(n12476), .B(n12475), .Z(n12493) );
  XNOR U12785 ( .A(n12494), .B(n12493), .Z(n12495) );
  XOR U12786 ( .A(n12496), .B(n12495), .Z(n12490) );
  AND U12787 ( .A(y[776]), .B(x[129]), .Z(n13219) );
  NAND U12788 ( .A(y[771]), .B(x[134]), .Z(n12443) );
  XNOR U12789 ( .A(n13219), .B(n12443), .Z(n12480) );
  XOR U12790 ( .A(n12896), .B(n12480), .Z(n12500) );
  NAND U12791 ( .A(x[130]), .B(y[775]), .Z(n13094) );
  NAND U12792 ( .A(x[131]), .B(y[774]), .Z(n12858) );
  XOR U12793 ( .A(n13094), .B(n12858), .Z(n12499) );
  XOR U12794 ( .A(n12500), .B(n12499), .Z(n12488) );
  NAND U12795 ( .A(x[133]), .B(y[775]), .Z(n12684) );
  NANDN U12796 ( .A(n12684), .B(n12479), .Z(n12447) );
  NAND U12797 ( .A(n12445), .B(n12444), .Z(n12446) );
  NAND U12798 ( .A(n12447), .B(n12446), .Z(n12487) );
  XOR U12799 ( .A(n12488), .B(n12487), .Z(n12489) );
  XNOR U12800 ( .A(n12490), .B(n12489), .Z(n12463) );
  XOR U12801 ( .A(n12464), .B(n12463), .Z(n12512) );
  NAND U12802 ( .A(n12449), .B(n12448), .Z(n12453) );
  NANDN U12803 ( .A(n12451), .B(n12450), .Z(n12452) );
  NAND U12804 ( .A(n12453), .B(n12452), .Z(n12511) );
  NAND U12805 ( .A(n12455), .B(n12454), .Z(n12459) );
  NAND U12806 ( .A(n12457), .B(n12456), .Z(n12458) );
  NAND U12807 ( .A(n12459), .B(n12458), .Z(n12510) );
  XNOR U12808 ( .A(n12511), .B(n12510), .Z(n12513) );
  XNOR U12809 ( .A(n12504), .B(n12506), .Z(n12460) );
  XOR U12810 ( .A(n12503), .B(n12460), .Z(N298) );
  NANDN U12811 ( .A(n12462), .B(n12461), .Z(n12466) );
  NAND U12812 ( .A(n12464), .B(n12463), .Z(n12465) );
  AND U12813 ( .A(n12466), .B(n12465), .Z(n12575) );
  AND U12814 ( .A(x[135]), .B(y[772]), .Z(n12468) );
  NAND U12815 ( .A(n12468), .B(n12467), .Z(n12472) );
  NAND U12816 ( .A(n12470), .B(n12469), .Z(n12471) );
  AND U12817 ( .A(n12472), .B(n12471), .Z(n12566) );
  AND U12818 ( .A(y[774]), .B(x[132]), .Z(n12474) );
  NAND U12819 ( .A(y[771]), .B(x[135]), .Z(n12473) );
  XNOR U12820 ( .A(n12474), .B(n12473), .Z(n12538) );
  AND U12821 ( .A(x[134]), .B(y[772]), .Z(n12537) );
  XOR U12822 ( .A(n12538), .B(n12537), .Z(n12564) );
  AND U12823 ( .A(x[136]), .B(y[770]), .Z(n12742) );
  NAND U12824 ( .A(x[137]), .B(y[769]), .Z(n12547) );
  XNOR U12825 ( .A(o[138]), .B(n12547), .Z(n12558) );
  XOR U12826 ( .A(n12742), .B(n12558), .Z(n12560) );
  XNOR U12827 ( .A(n12560), .B(n12559), .Z(n12563) );
  XNOR U12828 ( .A(n12564), .B(n12563), .Z(n12565) );
  XOR U12829 ( .A(n12566), .B(n12565), .Z(n12526) );
  AND U12830 ( .A(x[137]), .B(y[777]), .Z(n13127) );
  NAND U12831 ( .A(n13127), .B(n12891), .Z(n12478) );
  NAND U12832 ( .A(n12476), .B(n12475), .Z(n12477) );
  AND U12833 ( .A(n12478), .B(n12477), .Z(n12524) );
  AND U12834 ( .A(x[134]), .B(y[776]), .Z(n12777) );
  NAND U12835 ( .A(n12777), .B(n12479), .Z(n12482) );
  NAND U12836 ( .A(n12896), .B(n12480), .Z(n12481) );
  AND U12837 ( .A(n12482), .B(n12481), .Z(n12532) );
  AND U12838 ( .A(y[778]), .B(x[128]), .Z(n12484) );
  NAND U12839 ( .A(y[768]), .B(x[138]), .Z(n12483) );
  XNOR U12840 ( .A(n12484), .B(n12483), .Z(n12542) );
  ANDN U12841 ( .B(o[137]), .A(n12485), .Z(n12541) );
  XOR U12842 ( .A(n12542), .B(n12541), .Z(n12530) );
  AND U12843 ( .A(y[777]), .B(x[129]), .Z(n13422) );
  NAND U12844 ( .A(y[775]), .B(x[131]), .Z(n12486) );
  XNOR U12845 ( .A(n13422), .B(n12486), .Z(n12554) );
  NAND U12846 ( .A(x[130]), .B(y[776]), .Z(n12555) );
  XNOR U12847 ( .A(n12554), .B(n12555), .Z(n12529) );
  XOR U12848 ( .A(n12530), .B(n12529), .Z(n12531) );
  XNOR U12849 ( .A(n12532), .B(n12531), .Z(n12523) );
  XNOR U12850 ( .A(n12524), .B(n12523), .Z(n12525) );
  XOR U12851 ( .A(n12526), .B(n12525), .Z(n12573) );
  NAND U12852 ( .A(n12488), .B(n12487), .Z(n12492) );
  NANDN U12853 ( .A(n12490), .B(n12489), .Z(n12491) );
  AND U12854 ( .A(n12492), .B(n12491), .Z(n12520) );
  NANDN U12855 ( .A(n12494), .B(n12493), .Z(n12498) );
  NAND U12856 ( .A(n12496), .B(n12495), .Z(n12497) );
  AND U12857 ( .A(n12498), .B(n12497), .Z(n12517) );
  AND U12858 ( .A(n13094), .B(n12858), .Z(n12502) );
  NANDN U12859 ( .A(n12500), .B(n12499), .Z(n12501) );
  NANDN U12860 ( .A(n12502), .B(n12501), .Z(n12518) );
  XNOR U12861 ( .A(n12517), .B(n12518), .Z(n12519) );
  XOR U12862 ( .A(n12520), .B(n12519), .Z(n12572) );
  XOR U12863 ( .A(n12573), .B(n12572), .Z(n12574) );
  XNOR U12864 ( .A(n12575), .B(n12574), .Z(n12571) );
  NANDN U12865 ( .A(n12503), .B(n12504), .Z(n12509) );
  NOR U12866 ( .A(n12505), .B(n12504), .Z(n12507) );
  OR U12867 ( .A(n12507), .B(n12506), .Z(n12508) );
  AND U12868 ( .A(n12509), .B(n12508), .Z(n12570) );
  NAND U12869 ( .A(n12511), .B(n12510), .Z(n12515) );
  NANDN U12870 ( .A(n12513), .B(n12512), .Z(n12514) );
  AND U12871 ( .A(n12515), .B(n12514), .Z(n12569) );
  XOR U12872 ( .A(n12570), .B(n12569), .Z(n12516) );
  XNOR U12873 ( .A(n12571), .B(n12516), .Z(N299) );
  NANDN U12874 ( .A(n12518), .B(n12517), .Z(n12522) );
  NANDN U12875 ( .A(n12520), .B(n12519), .Z(n12521) );
  AND U12876 ( .A(n12522), .B(n12521), .Z(n12639) );
  NANDN U12877 ( .A(n12524), .B(n12523), .Z(n12528) );
  NANDN U12878 ( .A(n12526), .B(n12525), .Z(n12527) );
  AND U12879 ( .A(n12528), .B(n12527), .Z(n12637) );
  NAND U12880 ( .A(n12530), .B(n12529), .Z(n12534) );
  NANDN U12881 ( .A(n12532), .B(n12531), .Z(n12533) );
  AND U12882 ( .A(n12534), .B(n12533), .Z(n12630) );
  AND U12883 ( .A(x[135]), .B(y[774]), .Z(n12536) );
  AND U12884 ( .A(x[132]), .B(y[771]), .Z(n12535) );
  NAND U12885 ( .A(n12536), .B(n12535), .Z(n12540) );
  NAND U12886 ( .A(n12538), .B(n12537), .Z(n12539) );
  AND U12887 ( .A(n12540), .B(n12539), .Z(n12628) );
  AND U12888 ( .A(x[138]), .B(y[778]), .Z(n13320) );
  NAND U12889 ( .A(n13320), .B(n12891), .Z(n12544) );
  NAND U12890 ( .A(n12542), .B(n12541), .Z(n12543) );
  AND U12891 ( .A(n12544), .B(n12543), .Z(n12624) );
  AND U12892 ( .A(y[779]), .B(x[128]), .Z(n12546) );
  NAND U12893 ( .A(y[768]), .B(x[139]), .Z(n12545) );
  XNOR U12894 ( .A(n12546), .B(n12545), .Z(n12601) );
  ANDN U12895 ( .B(o[138]), .A(n12547), .Z(n12600) );
  XOR U12896 ( .A(n12601), .B(n12600), .Z(n12622) );
  AND U12897 ( .A(y[778]), .B(x[129]), .Z(n12549) );
  NAND U12898 ( .A(y[773]), .B(x[134]), .Z(n12548) );
  XNOR U12899 ( .A(n12549), .B(n12548), .Z(n12591) );
  NAND U12900 ( .A(x[138]), .B(y[769]), .Z(n12609) );
  XNOR U12901 ( .A(o[139]), .B(n12609), .Z(n12590) );
  XOR U12902 ( .A(n12591), .B(n12590), .Z(n12621) );
  XOR U12903 ( .A(n12622), .B(n12621), .Z(n12623) );
  XNOR U12904 ( .A(n12624), .B(n12623), .Z(n12627) );
  XNOR U12905 ( .A(n12628), .B(n12627), .Z(n12629) );
  XOR U12906 ( .A(n12630), .B(n12629), .Z(n12612) );
  NAND U12907 ( .A(x[131]), .B(y[776]), .Z(n13590) );
  NAND U12908 ( .A(y[777]), .B(x[130]), .Z(n12550) );
  XNOR U12909 ( .A(n12551), .B(n12550), .Z(n12586) );
  AND U12910 ( .A(x[132]), .B(y[775]), .Z(n12585) );
  XNOR U12911 ( .A(n12586), .B(n12585), .Z(n12616) );
  XOR U12912 ( .A(n13590), .B(n12616), .Z(n12618) );
  AND U12913 ( .A(y[770]), .B(x[137]), .Z(n12553) );
  NAND U12914 ( .A(y[772]), .B(x[135]), .Z(n12552) );
  XNOR U12915 ( .A(n12553), .B(n12552), .Z(n12605) );
  AND U12916 ( .A(x[136]), .B(y[771]), .Z(n12604) );
  XNOR U12917 ( .A(n12605), .B(n12604), .Z(n12617) );
  XOR U12918 ( .A(n12618), .B(n12617), .Z(n12582) );
  NAND U12919 ( .A(x[131]), .B(y[777]), .Z(n12675) );
  AND U12920 ( .A(x[129]), .B(y[775]), .Z(n12886) );
  NANDN U12921 ( .A(n12675), .B(n12886), .Z(n12557) );
  NANDN U12922 ( .A(n12555), .B(n12554), .Z(n12556) );
  AND U12923 ( .A(n12557), .B(n12556), .Z(n12580) );
  NAND U12924 ( .A(n12742), .B(n12558), .Z(n12562) );
  NAND U12925 ( .A(n12560), .B(n12559), .Z(n12561) );
  NAND U12926 ( .A(n12562), .B(n12561), .Z(n12579) );
  XNOR U12927 ( .A(n12580), .B(n12579), .Z(n12581) );
  XOR U12928 ( .A(n12582), .B(n12581), .Z(n12611) );
  NANDN U12929 ( .A(n12564), .B(n12563), .Z(n12568) );
  NAND U12930 ( .A(n12566), .B(n12565), .Z(n12567) );
  NAND U12931 ( .A(n12568), .B(n12567), .Z(n12610) );
  XOR U12932 ( .A(n12611), .B(n12610), .Z(n12613) );
  XNOR U12933 ( .A(n12612), .B(n12613), .Z(n12636) );
  XNOR U12934 ( .A(n12637), .B(n12636), .Z(n12638) );
  XOR U12935 ( .A(n12639), .B(n12638), .Z(n12635) );
  NAND U12936 ( .A(n12573), .B(n12572), .Z(n12577) );
  NAND U12937 ( .A(n12575), .B(n12574), .Z(n12576) );
  AND U12938 ( .A(n12577), .B(n12576), .Z(n12634) );
  XOR U12939 ( .A(n12633), .B(n12634), .Z(n12578) );
  XNOR U12940 ( .A(n12635), .B(n12578), .Z(N300) );
  NANDN U12941 ( .A(n12580), .B(n12579), .Z(n12584) );
  NANDN U12942 ( .A(n12582), .B(n12581), .Z(n12583) );
  AND U12943 ( .A(n12584), .B(n12583), .Z(n12717) );
  AND U12944 ( .A(x[133]), .B(y[777]), .Z(n13085) );
  NAND U12945 ( .A(n13314), .B(n13085), .Z(n12588) );
  NAND U12946 ( .A(n12586), .B(n12585), .Z(n12587) );
  NAND U12947 ( .A(n12588), .B(n12587), .Z(n12663) );
  AND U12948 ( .A(x[134]), .B(y[778]), .Z(n12903) );
  NAND U12949 ( .A(n12903), .B(n12589), .Z(n12593) );
  NAND U12950 ( .A(n12591), .B(n12590), .Z(n12592) );
  NAND U12951 ( .A(n12593), .B(n12592), .Z(n12662) );
  XOR U12952 ( .A(n12663), .B(n12662), .Z(n12664) );
  AND U12953 ( .A(x[137]), .B(y[771]), .Z(n13311) );
  AND U12954 ( .A(y[776]), .B(x[132]), .Z(n12595) );
  NAND U12955 ( .A(y[770]), .B(x[138]), .Z(n12594) );
  XOR U12956 ( .A(n12595), .B(n12594), .Z(n12707) );
  XNOR U12957 ( .A(n13311), .B(n12707), .Z(n12685) );
  NAND U12958 ( .A(x[135]), .B(y[773]), .Z(n12683) );
  XOR U12959 ( .A(n12684), .B(n12683), .Z(n12686) );
  AND U12960 ( .A(y[780]), .B(x[128]), .Z(n12597) );
  NAND U12961 ( .A(y[768]), .B(x[140]), .Z(n12596) );
  XNOR U12962 ( .A(n12597), .B(n12596), .Z(n12700) );
  NAND U12963 ( .A(x[139]), .B(y[769]), .Z(n12680) );
  XNOR U12964 ( .A(o[140]), .B(n12680), .Z(n12699) );
  XOR U12965 ( .A(n12700), .B(n12699), .Z(n12669) );
  AND U12966 ( .A(y[778]), .B(x[130]), .Z(n12599) );
  NAND U12967 ( .A(y[772]), .B(x[136]), .Z(n12598) );
  XNOR U12968 ( .A(n12599), .B(n12598), .Z(n12674) );
  XOR U12969 ( .A(n12669), .B(n12668), .Z(n12670) );
  XNOR U12970 ( .A(n12664), .B(n12665), .Z(n12715) );
  AND U12971 ( .A(x[139]), .B(y[779]), .Z(n13686) );
  NAND U12972 ( .A(n13686), .B(n12891), .Z(n12603) );
  NAND U12973 ( .A(n12601), .B(n12600), .Z(n12602) );
  AND U12974 ( .A(n12603), .B(n12602), .Z(n12692) );
  AND U12975 ( .A(x[135]), .B(y[770]), .Z(n12834) );
  AND U12976 ( .A(x[137]), .B(y[772]), .Z(n12682) );
  NAND U12977 ( .A(n12834), .B(n12682), .Z(n12607) );
  NAND U12978 ( .A(n12605), .B(n12604), .Z(n12606) );
  AND U12979 ( .A(n12607), .B(n12606), .Z(n12690) );
  AND U12980 ( .A(y[779]), .B(x[129]), .Z(n13342) );
  NAND U12981 ( .A(y[774]), .B(x[134]), .Z(n12608) );
  XNOR U12982 ( .A(n13342), .B(n12608), .Z(n12696) );
  ANDN U12983 ( .B(o[139]), .A(n12609), .Z(n12695) );
  XOR U12984 ( .A(n12696), .B(n12695), .Z(n12689) );
  XNOR U12985 ( .A(n12690), .B(n12689), .Z(n12691) );
  XNOR U12986 ( .A(n12692), .B(n12691), .Z(n12714) );
  XOR U12987 ( .A(n12715), .B(n12714), .Z(n12716) );
  XOR U12988 ( .A(n12717), .B(n12716), .Z(n12644) );
  NAND U12989 ( .A(n12611), .B(n12610), .Z(n12615) );
  NAND U12990 ( .A(n12613), .B(n12612), .Z(n12614) );
  NAND U12991 ( .A(n12615), .B(n12614), .Z(n12643) );
  XOR U12992 ( .A(n12644), .B(n12643), .Z(n12646) );
  NAND U12993 ( .A(n13590), .B(n12616), .Z(n12620) );
  NAND U12994 ( .A(n12618), .B(n12617), .Z(n12619) );
  AND U12995 ( .A(n12620), .B(n12619), .Z(n12657) );
  NAND U12996 ( .A(n12622), .B(n12621), .Z(n12626) );
  NANDN U12997 ( .A(n12624), .B(n12623), .Z(n12625) );
  AND U12998 ( .A(n12626), .B(n12625), .Z(n12656) );
  XNOR U12999 ( .A(n12657), .B(n12656), .Z(n12658) );
  NANDN U13000 ( .A(n12628), .B(n12627), .Z(n12632) );
  NANDN U13001 ( .A(n12630), .B(n12629), .Z(n12631) );
  NAND U13002 ( .A(n12632), .B(n12631), .Z(n12659) );
  XNOR U13003 ( .A(n12658), .B(n12659), .Z(n12645) );
  XNOR U13004 ( .A(n12646), .B(n12645), .Z(n12652) );
  NANDN U13005 ( .A(n12637), .B(n12636), .Z(n12641) );
  NANDN U13006 ( .A(n12639), .B(n12638), .Z(n12640) );
  AND U13007 ( .A(n12641), .B(n12640), .Z(n12651) );
  IV U13008 ( .A(n12651), .Z(n12649) );
  XOR U13009 ( .A(n12650), .B(n12649), .Z(n12642) );
  XNOR U13010 ( .A(n12652), .B(n12642), .Z(N301) );
  NAND U13011 ( .A(n12644), .B(n12643), .Z(n12648) );
  NAND U13012 ( .A(n12646), .B(n12645), .Z(n12647) );
  AND U13013 ( .A(n12648), .B(n12647), .Z(n12728) );
  NANDN U13014 ( .A(n12649), .B(n12650), .Z(n12655) );
  NOR U13015 ( .A(n12651), .B(n12650), .Z(n12653) );
  OR U13016 ( .A(n12653), .B(n12652), .Z(n12654) );
  AND U13017 ( .A(n12655), .B(n12654), .Z(n12727) );
  NANDN U13018 ( .A(n12657), .B(n12656), .Z(n12661) );
  NANDN U13019 ( .A(n12659), .B(n12658), .Z(n12660) );
  AND U13020 ( .A(n12661), .B(n12660), .Z(n12724) );
  NAND U13021 ( .A(n12663), .B(n12662), .Z(n12667) );
  NANDN U13022 ( .A(n12665), .B(n12664), .Z(n12666) );
  NAND U13023 ( .A(n12667), .B(n12666), .Z(n12784) );
  NAND U13024 ( .A(n12669), .B(n12668), .Z(n12673) );
  NANDN U13025 ( .A(n12671), .B(n12670), .Z(n12672) );
  NAND U13026 ( .A(n12673), .B(n12672), .Z(n12792) );
  AND U13027 ( .A(x[136]), .B(y[778]), .Z(n13929) );
  AND U13028 ( .A(x[130]), .B(y[772]), .Z(n12843) );
  NAND U13029 ( .A(n13929), .B(n12843), .Z(n12677) );
  NANDN U13030 ( .A(n12675), .B(n12674), .Z(n12676) );
  AND U13031 ( .A(n12677), .B(n12676), .Z(n12758) );
  AND U13032 ( .A(y[780]), .B(x[129]), .Z(n12679) );
  NAND U13033 ( .A(y[774]), .B(x[135]), .Z(n12678) );
  XNOR U13034 ( .A(n12679), .B(n12678), .Z(n12749) );
  ANDN U13035 ( .B(o[140]), .A(n12680), .Z(n12748) );
  XOR U13036 ( .A(n12749), .B(n12748), .Z(n12756) );
  AND U13037 ( .A(x[134]), .B(y[775]), .Z(n13720) );
  NAND U13038 ( .A(y[779]), .B(x[130]), .Z(n12681) );
  XOR U13039 ( .A(n12682), .B(n12681), .Z(n12761) );
  XNOR U13040 ( .A(n13720), .B(n12761), .Z(n12755) );
  XOR U13041 ( .A(n12756), .B(n12755), .Z(n12757) );
  XNOR U13042 ( .A(n12758), .B(n12757), .Z(n12791) );
  NAND U13043 ( .A(n12684), .B(n12683), .Z(n12688) );
  ANDN U13044 ( .B(n12686), .A(n12685), .Z(n12687) );
  ANDN U13045 ( .B(n12688), .A(n12687), .Z(n12790) );
  XOR U13046 ( .A(n12791), .B(n12790), .Z(n12793) );
  XOR U13047 ( .A(n12792), .B(n12793), .Z(n12785) );
  XOR U13048 ( .A(n12784), .B(n12785), .Z(n12787) );
  NANDN U13049 ( .A(n12690), .B(n12689), .Z(n12694) );
  NANDN U13050 ( .A(n12692), .B(n12691), .Z(n12693) );
  AND U13051 ( .A(n12694), .B(n12693), .Z(n12733) );
  NAND U13052 ( .A(x[134]), .B(y[779]), .Z(n13087) );
  AND U13053 ( .A(x[129]), .B(y[774]), .Z(n12747) );
  NANDN U13054 ( .A(n13087), .B(n12747), .Z(n12698) );
  NAND U13055 ( .A(n12696), .B(n12695), .Z(n12697) );
  AND U13056 ( .A(n12698), .B(n12697), .Z(n12739) );
  AND U13057 ( .A(x[140]), .B(y[780]), .Z(n13935) );
  NAND U13058 ( .A(n12891), .B(n13935), .Z(n12702) );
  NAND U13059 ( .A(n12700), .B(n12699), .Z(n12701) );
  AND U13060 ( .A(n12702), .B(n12701), .Z(n12737) );
  AND U13061 ( .A(x[138]), .B(y[771]), .Z(n13602) );
  AND U13062 ( .A(y[773]), .B(x[136]), .Z(n12704) );
  NAND U13063 ( .A(y[770]), .B(x[139]), .Z(n12703) );
  XOR U13064 ( .A(n12704), .B(n12703), .Z(n12744) );
  XNOR U13065 ( .A(n13602), .B(n12744), .Z(n12736) );
  XNOR U13066 ( .A(n12737), .B(n12736), .Z(n12738) );
  XNOR U13067 ( .A(n12739), .B(n12738), .Z(n12731) );
  AND U13068 ( .A(x[138]), .B(y[776]), .Z(n12706) );
  AND U13069 ( .A(x[132]), .B(y[770]), .Z(n12705) );
  NAND U13070 ( .A(n12706), .B(n12705), .Z(n12709) );
  NANDN U13071 ( .A(n12707), .B(n13311), .Z(n12708) );
  AND U13072 ( .A(n12709), .B(n12708), .Z(n12781) );
  AND U13073 ( .A(y[781]), .B(x[128]), .Z(n12711) );
  NAND U13074 ( .A(y[768]), .B(x[141]), .Z(n12710) );
  XNOR U13075 ( .A(n12711), .B(n12710), .Z(n12773) );
  NAND U13076 ( .A(x[140]), .B(y[769]), .Z(n12766) );
  XNOR U13077 ( .A(o[141]), .B(n12766), .Z(n12772) );
  XOR U13078 ( .A(n12773), .B(n12772), .Z(n12779) );
  AND U13079 ( .A(y[776]), .B(x[133]), .Z(n12713) );
  NAND U13080 ( .A(y[778]), .B(x[131]), .Z(n12712) );
  XNOR U13081 ( .A(n12713), .B(n12712), .Z(n12768) );
  NAND U13082 ( .A(x[132]), .B(y[777]), .Z(n12769) );
  XNOR U13083 ( .A(n12768), .B(n12769), .Z(n12778) );
  XOR U13084 ( .A(n12779), .B(n12778), .Z(n12780) );
  XNOR U13085 ( .A(n12781), .B(n12780), .Z(n12730) );
  XOR U13086 ( .A(n12731), .B(n12730), .Z(n12732) );
  XNOR U13087 ( .A(n12733), .B(n12732), .Z(n12786) );
  XOR U13088 ( .A(n12787), .B(n12786), .Z(n12722) );
  NAND U13089 ( .A(n12715), .B(n12714), .Z(n12719) );
  NANDN U13090 ( .A(n12717), .B(n12716), .Z(n12718) );
  AND U13091 ( .A(n12719), .B(n12718), .Z(n12721) );
  XNOR U13092 ( .A(n12722), .B(n12721), .Z(n12723) );
  XNOR U13093 ( .A(n12724), .B(n12723), .Z(n12729) );
  XNOR U13094 ( .A(n12727), .B(n12729), .Z(n12720) );
  XOR U13095 ( .A(n12728), .B(n12720), .Z(N302) );
  NANDN U13096 ( .A(n12722), .B(n12721), .Z(n12726) );
  NANDN U13097 ( .A(n12724), .B(n12723), .Z(n12725) );
  NAND U13098 ( .A(n12726), .B(n12725), .Z(n12805) );
  IV U13099 ( .A(n12805), .Z(n12803) );
  NAND U13100 ( .A(n12731), .B(n12730), .Z(n12735) );
  NANDN U13101 ( .A(n12733), .B(n12732), .Z(n12734) );
  AND U13102 ( .A(n12735), .B(n12734), .Z(n12813) );
  NANDN U13103 ( .A(n12737), .B(n12736), .Z(n12741) );
  NANDN U13104 ( .A(n12739), .B(n12738), .Z(n12740) );
  AND U13105 ( .A(n12741), .B(n12740), .Z(n12819) );
  AND U13106 ( .A(x[139]), .B(y[773]), .Z(n12743) );
  NAND U13107 ( .A(n12743), .B(n12742), .Z(n12746) );
  NANDN U13108 ( .A(n12744), .B(n13602), .Z(n12745) );
  AND U13109 ( .A(n12746), .B(n12745), .Z(n12874) );
  AND U13110 ( .A(x[135]), .B(y[780]), .Z(n13323) );
  NAND U13111 ( .A(n13323), .B(n12747), .Z(n12751) );
  NAND U13112 ( .A(n12749), .B(n12748), .Z(n12750) );
  NAND U13113 ( .A(n12751), .B(n12750), .Z(n12873) );
  AND U13114 ( .A(x[132]), .B(y[778]), .Z(n13241) );
  AND U13115 ( .A(y[779]), .B(x[131]), .Z(n12753) );
  NAND U13116 ( .A(y[774]), .B(x[136]), .Z(n12752) );
  XOR U13117 ( .A(n12753), .B(n12752), .Z(n12859) );
  XOR U13118 ( .A(n13241), .B(n12868), .Z(n12870) );
  AND U13119 ( .A(x[137]), .B(y[773]), .Z(n13425) );
  AND U13120 ( .A(y[780]), .B(x[130]), .Z(n12754) );
  AND U13121 ( .A(y[772]), .B(x[138]), .Z(n13449) );
  XOR U13122 ( .A(n12754), .B(n13449), .Z(n12844) );
  XOR U13123 ( .A(n13425), .B(n12844), .Z(n12869) );
  XOR U13124 ( .A(n12870), .B(n12869), .Z(n12875) );
  XOR U13125 ( .A(n12876), .B(n12875), .Z(n12817) );
  NAND U13126 ( .A(n12756), .B(n12755), .Z(n12760) );
  NANDN U13127 ( .A(n12758), .B(n12757), .Z(n12759) );
  AND U13128 ( .A(n12760), .B(n12759), .Z(n12816) );
  XNOR U13129 ( .A(n12817), .B(n12816), .Z(n12818) );
  XOR U13130 ( .A(n12819), .B(n12818), .Z(n12811) );
  AND U13131 ( .A(x[137]), .B(y[779]), .Z(n13322) );
  NAND U13132 ( .A(n13322), .B(n12843), .Z(n12763) );
  NANDN U13133 ( .A(n12761), .B(n13720), .Z(n12762) );
  AND U13134 ( .A(n12763), .B(n12762), .Z(n12831) );
  AND U13135 ( .A(y[782]), .B(x[128]), .Z(n12765) );
  NAND U13136 ( .A(y[768]), .B(x[142]), .Z(n12764) );
  XNOR U13137 ( .A(n12765), .B(n12764), .Z(n12854) );
  ANDN U13138 ( .B(o[141]), .A(n12766), .Z(n12853) );
  XOR U13139 ( .A(n12854), .B(n12853), .Z(n12829) );
  AND U13140 ( .A(y[770]), .B(x[140]), .Z(n13417) );
  NAND U13141 ( .A(y[775]), .B(x[135]), .Z(n12767) );
  XNOR U13142 ( .A(n13417), .B(n12767), .Z(n12836) );
  NAND U13143 ( .A(x[141]), .B(y[769]), .Z(n12842) );
  XNOR U13144 ( .A(o[142]), .B(n12842), .Z(n12835) );
  XOR U13145 ( .A(n12836), .B(n12835), .Z(n12828) );
  XOR U13146 ( .A(n12829), .B(n12828), .Z(n12830) );
  AND U13147 ( .A(x[133]), .B(y[778]), .Z(n12904) );
  NANDN U13148 ( .A(n13590), .B(n12904), .Z(n12771) );
  NANDN U13149 ( .A(n12769), .B(n12768), .Z(n12770) );
  AND U13150 ( .A(n12771), .B(n12770), .Z(n12825) );
  AND U13151 ( .A(x[141]), .B(y[781]), .Z(n14167) );
  NAND U13152 ( .A(n14167), .B(n12891), .Z(n12775) );
  NAND U13153 ( .A(n12773), .B(n12772), .Z(n12774) );
  AND U13154 ( .A(n12775), .B(n12774), .Z(n12823) );
  NAND U13155 ( .A(y[771]), .B(x[139]), .Z(n12776) );
  XNOR U13156 ( .A(n12777), .B(n12776), .Z(n12849) );
  NAND U13157 ( .A(x[129]), .B(y[781]), .Z(n12850) );
  XOR U13158 ( .A(n12825), .B(n12824), .Z(n12879) );
  XOR U13159 ( .A(n12880), .B(n12879), .Z(n12882) );
  NAND U13160 ( .A(n12779), .B(n12778), .Z(n12783) );
  NANDN U13161 ( .A(n12781), .B(n12780), .Z(n12782) );
  AND U13162 ( .A(n12783), .B(n12782), .Z(n12881) );
  XNOR U13163 ( .A(n12882), .B(n12881), .Z(n12810) );
  XNOR U13164 ( .A(n12811), .B(n12810), .Z(n12812) );
  XNOR U13165 ( .A(n12813), .B(n12812), .Z(n12799) );
  NAND U13166 ( .A(n12785), .B(n12784), .Z(n12789) );
  NAND U13167 ( .A(n12787), .B(n12786), .Z(n12788) );
  NAND U13168 ( .A(n12789), .B(n12788), .Z(n12798) );
  NAND U13169 ( .A(n12791), .B(n12790), .Z(n12795) );
  NAND U13170 ( .A(n12793), .B(n12792), .Z(n12794) );
  NAND U13171 ( .A(n12795), .B(n12794), .Z(n12797) );
  XNOR U13172 ( .A(n12798), .B(n12797), .Z(n12800) );
  XNOR U13173 ( .A(n12804), .B(n12806), .Z(n12796) );
  XOR U13174 ( .A(n12803), .B(n12796), .Z(N303) );
  NAND U13175 ( .A(n12798), .B(n12797), .Z(n12802) );
  NANDN U13176 ( .A(n12800), .B(n12799), .Z(n12801) );
  AND U13177 ( .A(n12802), .B(n12801), .Z(n12974) );
  NANDN U13178 ( .A(n12803), .B(n12804), .Z(n12809) );
  NOR U13179 ( .A(n12805), .B(n12804), .Z(n12807) );
  OR U13180 ( .A(n12807), .B(n12806), .Z(n12808) );
  AND U13181 ( .A(n12809), .B(n12808), .Z(n12975) );
  NANDN U13182 ( .A(n12811), .B(n12810), .Z(n12815) );
  NANDN U13183 ( .A(n12813), .B(n12812), .Z(n12814) );
  AND U13184 ( .A(n12815), .B(n12814), .Z(n12971) );
  NANDN U13185 ( .A(n12817), .B(n12816), .Z(n12821) );
  NAND U13186 ( .A(n12819), .B(n12818), .Z(n12820) );
  AND U13187 ( .A(n12821), .B(n12820), .Z(n12947) );
  NANDN U13188 ( .A(n12823), .B(n12822), .Z(n12827) );
  NANDN U13189 ( .A(n12825), .B(n12824), .Z(n12826) );
  AND U13190 ( .A(n12827), .B(n12826), .Z(n12953) );
  NAND U13191 ( .A(n12829), .B(n12828), .Z(n12833) );
  NANDN U13192 ( .A(n12831), .B(n12830), .Z(n12832) );
  AND U13193 ( .A(n12833), .B(n12832), .Z(n12951) );
  AND U13194 ( .A(x[140]), .B(y[775]), .Z(n13315) );
  NAND U13195 ( .A(n13315), .B(n12834), .Z(n12838) );
  NAND U13196 ( .A(n12836), .B(n12835), .Z(n12837) );
  AND U13197 ( .A(n12838), .B(n12837), .Z(n12927) );
  AND U13198 ( .A(y[770]), .B(x[141]), .Z(n13708) );
  NAND U13199 ( .A(y[772]), .B(x[139]), .Z(n12839) );
  XNOR U13200 ( .A(n13708), .B(n12839), .Z(n12931) );
  AND U13201 ( .A(x[140]), .B(y[771]), .Z(n12930) );
  XOR U13202 ( .A(n12931), .B(n12930), .Z(n12925) );
  AND U13203 ( .A(y[783]), .B(x[128]), .Z(n12841) );
  NAND U13204 ( .A(y[768]), .B(x[143]), .Z(n12840) );
  XNOR U13205 ( .A(n12841), .B(n12840), .Z(n12893) );
  ANDN U13206 ( .B(o[142]), .A(n12842), .Z(n12892) );
  XNOR U13207 ( .A(n12893), .B(n12892), .Z(n12924) );
  XOR U13208 ( .A(n12927), .B(n12926), .Z(n12959) );
  NAND U13209 ( .A(x[138]), .B(y[780]), .Z(n13722) );
  NANDN U13210 ( .A(n13722), .B(n12843), .Z(n12846) );
  NAND U13211 ( .A(n13425), .B(n12844), .Z(n12845) );
  AND U13212 ( .A(n12846), .B(n12845), .Z(n12957) );
  AND U13213 ( .A(x[139]), .B(y[776]), .Z(n12848) );
  AND U13214 ( .A(x[134]), .B(y[771]), .Z(n12847) );
  NAND U13215 ( .A(n12848), .B(n12847), .Z(n12852) );
  NANDN U13216 ( .A(n12850), .B(n12849), .Z(n12851) );
  NAND U13217 ( .A(n12852), .B(n12851), .Z(n12956) );
  AND U13218 ( .A(x[142]), .B(y[782]), .Z(n14521) );
  NAND U13219 ( .A(n14521), .B(n12891), .Z(n12856) );
  NAND U13220 ( .A(n12854), .B(n12853), .Z(n12855) );
  AND U13221 ( .A(n12856), .B(n12855), .Z(n12919) );
  AND U13222 ( .A(x[136]), .B(y[779]), .Z(n12857) );
  NANDN U13223 ( .A(n12858), .B(n12857), .Z(n12861) );
  NANDN U13224 ( .A(n12859), .B(n13085), .Z(n12860) );
  NAND U13225 ( .A(n12861), .B(n12860), .Z(n12918) );
  AND U13226 ( .A(y[779]), .B(x[132]), .Z(n12863) );
  NAND U13227 ( .A(y[773]), .B(x[138]), .Z(n12862) );
  XNOR U13228 ( .A(n12863), .B(n12862), .Z(n12899) );
  AND U13229 ( .A(x[135]), .B(y[776]), .Z(n12898) );
  XOR U13230 ( .A(n12899), .B(n12898), .Z(n12906) );
  NAND U13231 ( .A(x[134]), .B(y[777]), .Z(n13005) );
  XNOR U13232 ( .A(n13005), .B(n12904), .Z(n12905) );
  AND U13233 ( .A(y[774]), .B(x[137]), .Z(n12865) );
  NAND U13234 ( .A(y[781]), .B(x[130]), .Z(n12864) );
  XNOR U13235 ( .A(n12865), .B(n12864), .Z(n12909) );
  NAND U13236 ( .A(x[131]), .B(y[780]), .Z(n12910) );
  AND U13237 ( .A(y[782]), .B(x[129]), .Z(n12867) );
  NAND U13238 ( .A(y[775]), .B(x[136]), .Z(n12866) );
  XNOR U13239 ( .A(n12867), .B(n12866), .Z(n12888) );
  NAND U13240 ( .A(x[142]), .B(y[769]), .Z(n12915) );
  XNOR U13241 ( .A(o[143]), .B(n12915), .Z(n12887) );
  XOR U13242 ( .A(n12888), .B(n12887), .Z(n12938) );
  XOR U13243 ( .A(n12939), .B(n12938), .Z(n12941) );
  XOR U13244 ( .A(n12940), .B(n12941), .Z(n12920) );
  XOR U13245 ( .A(n12921), .B(n12920), .Z(n12963) );
  NAND U13246 ( .A(n13241), .B(n12868), .Z(n12872) );
  NAND U13247 ( .A(n12870), .B(n12869), .Z(n12871) );
  AND U13248 ( .A(n12872), .B(n12871), .Z(n12962) );
  NANDN U13249 ( .A(n12874), .B(n12873), .Z(n12878) );
  NAND U13250 ( .A(n12876), .B(n12875), .Z(n12877) );
  NAND U13251 ( .A(n12878), .B(n12877), .Z(n12965) );
  XOR U13252 ( .A(n12944), .B(n12945), .Z(n12946) );
  NAND U13253 ( .A(n12880), .B(n12879), .Z(n12884) );
  NAND U13254 ( .A(n12882), .B(n12881), .Z(n12883) );
  AND U13255 ( .A(n12884), .B(n12883), .Z(n12969) );
  XOR U13256 ( .A(n12968), .B(n12969), .Z(n12970) );
  XNOR U13257 ( .A(n12971), .B(n12970), .Z(n12976) );
  XNOR U13258 ( .A(n12975), .B(n12976), .Z(n12885) );
  XOR U13259 ( .A(n12974), .B(n12885), .Z(N304) );
  AND U13260 ( .A(x[136]), .B(y[782]), .Z(n13611) );
  NAND U13261 ( .A(n13611), .B(n12886), .Z(n12890) );
  NAND U13262 ( .A(n12888), .B(n12887), .Z(n12889) );
  AND U13263 ( .A(n12890), .B(n12889), .Z(n13035) );
  AND U13264 ( .A(x[143]), .B(y[783]), .Z(n14840) );
  NAND U13265 ( .A(n14840), .B(n12891), .Z(n12895) );
  NAND U13266 ( .A(n12893), .B(n12892), .Z(n12894) );
  NAND U13267 ( .A(n12895), .B(n12894), .Z(n13034) );
  XNOR U13268 ( .A(n13035), .B(n13034), .Z(n13037) );
  AND U13269 ( .A(x[138]), .B(y[779]), .Z(n12897) );
  NAND U13270 ( .A(n12897), .B(n12896), .Z(n12901) );
  NAND U13271 ( .A(n12899), .B(n12898), .Z(n12900) );
  NAND U13272 ( .A(n12901), .B(n12900), .Z(n12992) );
  AND U13273 ( .A(x[128]), .B(y[784]), .Z(n13014) );
  NAND U13274 ( .A(x[144]), .B(y[768]), .Z(n13015) );
  XNOR U13275 ( .A(n13014), .B(n13015), .Z(n13017) );
  NAND U13276 ( .A(x[143]), .B(y[769]), .Z(n13002) );
  XNOR U13277 ( .A(o[144]), .B(n13002), .Z(n13016) );
  XOR U13278 ( .A(n13017), .B(n13016), .Z(n12991) );
  NAND U13279 ( .A(y[777]), .B(x[135]), .Z(n12902) );
  XNOR U13280 ( .A(n12903), .B(n12902), .Z(n13007) );
  AND U13281 ( .A(x[138]), .B(y[774]), .Z(n13006) );
  XOR U13282 ( .A(n13007), .B(n13006), .Z(n12990) );
  XOR U13283 ( .A(n12991), .B(n12990), .Z(n12993) );
  XOR U13284 ( .A(n12992), .B(n12993), .Z(n13036) );
  XOR U13285 ( .A(n13037), .B(n13036), .Z(n12987) );
  NANDN U13286 ( .A(n12904), .B(n13005), .Z(n12908) );
  NANDN U13287 ( .A(n12906), .B(n12905), .Z(n12907) );
  AND U13288 ( .A(n12908), .B(n12907), .Z(n12985) );
  NAND U13289 ( .A(x[137]), .B(y[781]), .Z(n13704) );
  NANDN U13290 ( .A(n13704), .B(n13314), .Z(n12912) );
  NANDN U13291 ( .A(n12910), .B(n12909), .Z(n12911) );
  AND U13292 ( .A(n12912), .B(n12911), .Z(n13025) );
  AND U13293 ( .A(y[783]), .B(x[129]), .Z(n12914) );
  NAND U13294 ( .A(y[776]), .B(x[136]), .Z(n12913) );
  XNOR U13295 ( .A(n12914), .B(n12913), .Z(n13011) );
  ANDN U13296 ( .B(o[143]), .A(n12915), .Z(n13010) );
  XOR U13297 ( .A(n13011), .B(n13010), .Z(n13023) );
  AND U13298 ( .A(y[770]), .B(x[142]), .Z(n12917) );
  NAND U13299 ( .A(y[773]), .B(x[139]), .Z(n12916) );
  XNOR U13300 ( .A(n12917), .B(n12916), .Z(n13046) );
  NAND U13301 ( .A(x[132]), .B(y[780]), .Z(n13047) );
  XNOR U13302 ( .A(n13046), .B(n13047), .Z(n13022) );
  XOR U13303 ( .A(n13023), .B(n13022), .Z(n13024) );
  XOR U13304 ( .A(n13025), .B(n13024), .Z(n12984) );
  NANDN U13305 ( .A(n12919), .B(n12918), .Z(n12923) );
  NAND U13306 ( .A(n12921), .B(n12920), .Z(n12922) );
  NAND U13307 ( .A(n12923), .B(n12922), .Z(n13029) );
  NANDN U13308 ( .A(n12925), .B(n12924), .Z(n12929) );
  NAND U13309 ( .A(n12927), .B(n12926), .Z(n12928) );
  AND U13310 ( .A(n12929), .B(n12928), .Z(n13060) );
  AND U13311 ( .A(x[139]), .B(y[770]), .Z(n13563) );
  AND U13312 ( .A(x[141]), .B(y[772]), .Z(n13056) );
  NAND U13313 ( .A(n13563), .B(n13056), .Z(n12933) );
  NAND U13314 ( .A(n12931), .B(n12930), .Z(n12932) );
  AND U13315 ( .A(n12933), .B(n12932), .Z(n13043) );
  AND U13316 ( .A(y[775]), .B(x[137]), .Z(n12935) );
  NAND U13317 ( .A(y[782]), .B(x[130]), .Z(n12934) );
  XNOR U13318 ( .A(n12935), .B(n12934), .Z(n13050) );
  NAND U13319 ( .A(x[131]), .B(y[781]), .Z(n13051) );
  XNOR U13320 ( .A(n13050), .B(n13051), .Z(n13041) );
  AND U13321 ( .A(x[140]), .B(y[772]), .Z(n13692) );
  AND U13322 ( .A(y[779]), .B(x[133]), .Z(n12937) );
  NAND U13323 ( .A(y[771]), .B(x[141]), .Z(n12936) );
  XOR U13324 ( .A(n12937), .B(n12936), .Z(n12997) );
  XNOR U13325 ( .A(n13692), .B(n12997), .Z(n13040) );
  XOR U13326 ( .A(n13041), .B(n13040), .Z(n13042) );
  XOR U13327 ( .A(n13043), .B(n13042), .Z(n13057) );
  NAND U13328 ( .A(n12939), .B(n12938), .Z(n12943) );
  NAND U13329 ( .A(n12941), .B(n12940), .Z(n12942) );
  AND U13330 ( .A(n12943), .B(n12942), .Z(n13058) );
  XOR U13331 ( .A(n13057), .B(n13058), .Z(n13059) );
  XOR U13332 ( .A(n13031), .B(n13030), .Z(n13067) );
  NAND U13333 ( .A(n12945), .B(n12944), .Z(n12949) );
  NANDN U13334 ( .A(n12947), .B(n12946), .Z(n12948) );
  AND U13335 ( .A(n12949), .B(n12948), .Z(n13066) );
  NANDN U13336 ( .A(n12951), .B(n12950), .Z(n12955) );
  NANDN U13337 ( .A(n12953), .B(n12952), .Z(n12954) );
  AND U13338 ( .A(n12955), .B(n12954), .Z(n12981) );
  NANDN U13339 ( .A(n12957), .B(n12956), .Z(n12961) );
  NANDN U13340 ( .A(n12959), .B(n12958), .Z(n12960) );
  AND U13341 ( .A(n12961), .B(n12960), .Z(n12979) );
  NANDN U13342 ( .A(n12963), .B(n12962), .Z(n12967) );
  NANDN U13343 ( .A(n12965), .B(n12964), .Z(n12966) );
  AND U13344 ( .A(n12967), .B(n12966), .Z(n12978) );
  XNOR U13345 ( .A(n13069), .B(n13068), .Z(n13065) );
  NAND U13346 ( .A(n12969), .B(n12968), .Z(n12973) );
  NANDN U13347 ( .A(n12971), .B(n12970), .Z(n12972) );
  NAND U13348 ( .A(n12973), .B(n12972), .Z(n13064) );
  XOR U13349 ( .A(n13064), .B(n13063), .Z(n12977) );
  XNOR U13350 ( .A(n13065), .B(n12977), .Z(N305) );
  NANDN U13351 ( .A(n12979), .B(n12978), .Z(n12983) );
  NANDN U13352 ( .A(n12981), .B(n12980), .Z(n12982) );
  AND U13353 ( .A(n12983), .B(n12982), .Z(n13179) );
  NANDN U13354 ( .A(n12985), .B(n12984), .Z(n12989) );
  NANDN U13355 ( .A(n12987), .B(n12986), .Z(n12988) );
  AND U13356 ( .A(n12989), .B(n12988), .Z(n13082) );
  NAND U13357 ( .A(n12991), .B(n12990), .Z(n12995) );
  NAND U13358 ( .A(n12993), .B(n12992), .Z(n12994) );
  AND U13359 ( .A(n12995), .B(n12994), .Z(n13166) );
  AND U13360 ( .A(x[141]), .B(y[779]), .Z(n13941) );
  NAND U13361 ( .A(n13941), .B(n12996), .Z(n12999) );
  NANDN U13362 ( .A(n12997), .B(n13692), .Z(n12998) );
  AND U13363 ( .A(n12999), .B(n12998), .Z(n13142) );
  AND U13364 ( .A(y[776]), .B(x[137]), .Z(n13001) );
  NAND U13365 ( .A(y[784]), .B(x[129]), .Z(n13000) );
  XNOR U13366 ( .A(n13001), .B(n13000), .Z(n13091) );
  ANDN U13367 ( .B(o[144]), .A(n13002), .Z(n13090) );
  XOR U13368 ( .A(n13091), .B(n13090), .Z(n13140) );
  AND U13369 ( .A(y[770]), .B(x[143]), .Z(n13004) );
  NAND U13370 ( .A(y[773]), .B(x[140]), .Z(n13003) );
  XNOR U13371 ( .A(n13004), .B(n13003), .Z(n13114) );
  NAND U13372 ( .A(x[142]), .B(y[771]), .Z(n13115) );
  XNOR U13373 ( .A(n13114), .B(n13115), .Z(n13139) );
  XOR U13374 ( .A(n13140), .B(n13139), .Z(n13141) );
  XNOR U13375 ( .A(n13142), .B(n13141), .Z(n13164) );
  AND U13376 ( .A(x[135]), .B(y[778]), .Z(n13102) );
  NANDN U13377 ( .A(n13005), .B(n13102), .Z(n13009) );
  NAND U13378 ( .A(n13007), .B(n13006), .Z(n13008) );
  AND U13379 ( .A(n13009), .B(n13008), .Z(n13152) );
  AND U13380 ( .A(x[136]), .B(y[783]), .Z(n13772) );
  NAND U13381 ( .A(n13219), .B(n13772), .Z(n13013) );
  NAND U13382 ( .A(n13011), .B(n13010), .Z(n13012) );
  NAND U13383 ( .A(n13013), .B(n13012), .Z(n13151) );
  XNOR U13384 ( .A(n13152), .B(n13151), .Z(n13154) );
  NANDN U13385 ( .A(n13015), .B(n13014), .Z(n13019) );
  NAND U13386 ( .A(n13017), .B(n13016), .Z(n13018) );
  AND U13387 ( .A(n13019), .B(n13018), .Z(n13148) );
  AND U13388 ( .A(x[128]), .B(y[785]), .Z(n13128) );
  NAND U13389 ( .A(x[145]), .B(y[768]), .Z(n13129) );
  XNOR U13390 ( .A(n13128), .B(n13129), .Z(n13131) );
  AND U13391 ( .A(x[144]), .B(y[769]), .Z(n13125) );
  XOR U13392 ( .A(o[145]), .B(n13125), .Z(n13130) );
  XOR U13393 ( .A(n13131), .B(n13130), .Z(n13146) );
  AND U13394 ( .A(y[783]), .B(x[130]), .Z(n13021) );
  NAND U13395 ( .A(y[775]), .B(x[138]), .Z(n13020) );
  XNOR U13396 ( .A(n13021), .B(n13020), .Z(n13095) );
  NAND U13397 ( .A(x[131]), .B(y[782]), .Z(n13096) );
  XOR U13398 ( .A(n13146), .B(n13145), .Z(n13147) );
  XNOR U13399 ( .A(n13148), .B(n13147), .Z(n13153) );
  XOR U13400 ( .A(n13154), .B(n13153), .Z(n13163) );
  XOR U13401 ( .A(n13164), .B(n13163), .Z(n13165) );
  XOR U13402 ( .A(n13166), .B(n13165), .Z(n13079) );
  NAND U13403 ( .A(n13023), .B(n13022), .Z(n13027) );
  NANDN U13404 ( .A(n13025), .B(n13024), .Z(n13026) );
  AND U13405 ( .A(n13027), .B(n13026), .Z(n13080) );
  XOR U13406 ( .A(n13079), .B(n13080), .Z(n13081) );
  NANDN U13407 ( .A(n13029), .B(n13028), .Z(n13033) );
  NAND U13408 ( .A(n13031), .B(n13030), .Z(n13032) );
  AND U13409 ( .A(n13033), .B(n13032), .Z(n13076) );
  NANDN U13410 ( .A(n13035), .B(n13034), .Z(n13039) );
  NAND U13411 ( .A(n13037), .B(n13036), .Z(n13038) );
  AND U13412 ( .A(n13039), .B(n13038), .Z(n13160) );
  NAND U13413 ( .A(n13041), .B(n13040), .Z(n13045) );
  NANDN U13414 ( .A(n13043), .B(n13042), .Z(n13044) );
  AND U13415 ( .A(n13045), .B(n13044), .Z(n13158) );
  NAND U13416 ( .A(x[142]), .B(y[773]), .Z(n13344) );
  NANDN U13417 ( .A(n13344), .B(n13563), .Z(n13049) );
  NANDN U13418 ( .A(n13047), .B(n13046), .Z(n13048) );
  AND U13419 ( .A(n13049), .B(n13048), .Z(n13108) );
  AND U13420 ( .A(y[782]), .B(x[137]), .Z(n13926) );
  NANDN U13421 ( .A(n13094), .B(n13926), .Z(n13053) );
  NANDN U13422 ( .A(n13051), .B(n13050), .Z(n13052) );
  NAND U13423 ( .A(n13053), .B(n13052), .Z(n13107) );
  XNOR U13424 ( .A(n13108), .B(n13107), .Z(n13110) );
  AND U13425 ( .A(x[133]), .B(y[780]), .Z(n13201) );
  NAND U13426 ( .A(y[777]), .B(x[136]), .Z(n13054) );
  XNOR U13427 ( .A(n13201), .B(n13054), .Z(n13086) );
  XOR U13428 ( .A(n13102), .B(n13101), .Z(n13104) );
  NAND U13429 ( .A(y[781]), .B(x[132]), .Z(n13055) );
  XNOR U13430 ( .A(n13056), .B(n13055), .Z(n13119) );
  NAND U13431 ( .A(x[139]), .B(y[774]), .Z(n13120) );
  XNOR U13432 ( .A(n13119), .B(n13120), .Z(n13103) );
  XOR U13433 ( .A(n13104), .B(n13103), .Z(n13109) );
  XOR U13434 ( .A(n13110), .B(n13109), .Z(n13157) );
  XNOR U13435 ( .A(n13158), .B(n13157), .Z(n13159) );
  XOR U13436 ( .A(n13160), .B(n13159), .Z(n13074) );
  NAND U13437 ( .A(n13058), .B(n13057), .Z(n13062) );
  NANDN U13438 ( .A(n13060), .B(n13059), .Z(n13061) );
  NAND U13439 ( .A(n13062), .B(n13061), .Z(n13073) );
  XOR U13440 ( .A(n13074), .B(n13073), .Z(n13075) );
  XOR U13441 ( .A(n13076), .B(n13075), .Z(n13176) );
  XOR U13442 ( .A(n13177), .B(n13176), .Z(n13178) );
  XOR U13443 ( .A(n13179), .B(n13178), .Z(n13172) );
  NANDN U13444 ( .A(n13067), .B(n13066), .Z(n13071) );
  NAND U13445 ( .A(n13069), .B(n13068), .Z(n13070) );
  NAND U13446 ( .A(n13071), .B(n13070), .Z(n13170) );
  IV U13447 ( .A(n13170), .Z(n13169) );
  XOR U13448 ( .A(n13171), .B(n13169), .Z(n13072) );
  XNOR U13449 ( .A(n13172), .B(n13072), .Z(N306) );
  NAND U13450 ( .A(n13074), .B(n13073), .Z(n13078) );
  NANDN U13451 ( .A(n13076), .B(n13075), .Z(n13077) );
  AND U13452 ( .A(n13078), .B(n13077), .Z(n13295) );
  NAND U13453 ( .A(n13080), .B(n13079), .Z(n13084) );
  NANDN U13454 ( .A(n13082), .B(n13081), .Z(n13083) );
  AND U13455 ( .A(n13084), .B(n13083), .Z(n13293) );
  NAND U13456 ( .A(x[136]), .B(y[780]), .Z(n13456) );
  NANDN U13457 ( .A(n13456), .B(n13085), .Z(n13089) );
  NANDN U13458 ( .A(n13087), .B(n13086), .Z(n13088) );
  AND U13459 ( .A(n13089), .B(n13088), .Z(n13274) );
  AND U13460 ( .A(x[137]), .B(y[784]), .Z(n14021) );
  NAND U13461 ( .A(n14021), .B(n13219), .Z(n13093) );
  NAND U13462 ( .A(n13091), .B(n13090), .Z(n13092) );
  NAND U13463 ( .A(n13093), .B(n13092), .Z(n13273) );
  AND U13464 ( .A(x[138]), .B(y[783]), .Z(n13946) );
  NANDN U13465 ( .A(n13094), .B(n13946), .Z(n13098) );
  NANDN U13466 ( .A(n13096), .B(n13095), .Z(n13097) );
  NAND U13467 ( .A(n13098), .B(n13097), .Z(n13251) );
  AND U13468 ( .A(y[783]), .B(x[131]), .Z(n13100) );
  NAND U13469 ( .A(y[773]), .B(x[141]), .Z(n13099) );
  XNOR U13470 ( .A(n13100), .B(n13099), .Z(n13234) );
  AND U13471 ( .A(x[140]), .B(y[774]), .Z(n13233) );
  XOR U13472 ( .A(n13234), .B(n13233), .Z(n13250) );
  AND U13473 ( .A(x[128]), .B(y[786]), .Z(n13225) );
  AND U13474 ( .A(x[146]), .B(y[768]), .Z(n13224) );
  XOR U13475 ( .A(n13225), .B(n13224), .Z(n13227) );
  AND U13476 ( .A(x[145]), .B(y[769]), .Z(n13246) );
  XOR U13477 ( .A(o[146]), .B(n13246), .Z(n13226) );
  XOR U13478 ( .A(n13227), .B(n13226), .Z(n13249) );
  XOR U13479 ( .A(n13250), .B(n13249), .Z(n13252) );
  XOR U13480 ( .A(n13251), .B(n13252), .Z(n13275) );
  XOR U13481 ( .A(n13276), .B(n13275), .Z(n13196) );
  NAND U13482 ( .A(n13102), .B(n13101), .Z(n13106) );
  NAND U13483 ( .A(n13104), .B(n13103), .Z(n13105) );
  AND U13484 ( .A(n13106), .B(n13105), .Z(n13195) );
  NANDN U13485 ( .A(n13108), .B(n13107), .Z(n13112) );
  NAND U13486 ( .A(n13110), .B(n13109), .Z(n13111) );
  NAND U13487 ( .A(n13112), .B(n13111), .Z(n13198) );
  AND U13488 ( .A(x[143]), .B(y[773]), .Z(n13113) );
  NAND U13489 ( .A(n13417), .B(n13113), .Z(n13117) );
  NANDN U13490 ( .A(n13115), .B(n13114), .Z(n13116) );
  AND U13491 ( .A(n13117), .B(n13116), .Z(n13268) );
  NAND U13492 ( .A(n14167), .B(n13118), .Z(n13122) );
  NANDN U13493 ( .A(n13120), .B(n13119), .Z(n13121) );
  NAND U13494 ( .A(n13122), .B(n13121), .Z(n13257) );
  AND U13495 ( .A(y[785]), .B(x[129]), .Z(n13124) );
  NAND U13496 ( .A(y[776]), .B(x[138]), .Z(n13123) );
  XNOR U13497 ( .A(n13124), .B(n13123), .Z(n13221) );
  AND U13498 ( .A(n13125), .B(o[145]), .Z(n13220) );
  XOR U13499 ( .A(n13221), .B(n13220), .Z(n13256) );
  NAND U13500 ( .A(y[771]), .B(x[143]), .Z(n13126) );
  XNOR U13501 ( .A(n13127), .B(n13126), .Z(n13212) );
  AND U13502 ( .A(x[142]), .B(y[772]), .Z(n13211) );
  XOR U13503 ( .A(n13212), .B(n13211), .Z(n13255) );
  XOR U13504 ( .A(n13256), .B(n13255), .Z(n13258) );
  XOR U13505 ( .A(n13257), .B(n13258), .Z(n13267) );
  NANDN U13506 ( .A(n13129), .B(n13128), .Z(n13133) );
  NAND U13507 ( .A(n13131), .B(n13130), .Z(n13132) );
  AND U13508 ( .A(n13133), .B(n13132), .Z(n13280) );
  AND U13509 ( .A(y[775]), .B(x[139]), .Z(n13135) );
  NAND U13510 ( .A(y[770]), .B(x[144]), .Z(n13134) );
  XNOR U13511 ( .A(n13135), .B(n13134), .Z(n13208) );
  AND U13512 ( .A(x[130]), .B(y[784]), .Z(n13207) );
  XOR U13513 ( .A(n13208), .B(n13207), .Z(n13279) );
  AND U13514 ( .A(y[781]), .B(x[133]), .Z(n13330) );
  NAND U13515 ( .A(y[780]), .B(x[134]), .Z(n13136) );
  XNOR U13516 ( .A(n13330), .B(n13136), .Z(n13203) );
  AND U13517 ( .A(y[782]), .B(x[132]), .Z(n13138) );
  NAND U13518 ( .A(y[778]), .B(x[136]), .Z(n13137) );
  XNOR U13519 ( .A(n13138), .B(n13137), .Z(n13243) );
  AND U13520 ( .A(x[135]), .B(y[779]), .Z(n13242) );
  XOR U13521 ( .A(n13243), .B(n13242), .Z(n13202) );
  XOR U13522 ( .A(n13203), .B(n13202), .Z(n13281) );
  XOR U13523 ( .A(n13282), .B(n13281), .Z(n13269) );
  XOR U13524 ( .A(n13270), .B(n13269), .Z(n13190) );
  NAND U13525 ( .A(n13140), .B(n13139), .Z(n13144) );
  NANDN U13526 ( .A(n13142), .B(n13141), .Z(n13143) );
  AND U13527 ( .A(n13144), .B(n13143), .Z(n13261) );
  NAND U13528 ( .A(n13146), .B(n13145), .Z(n13150) );
  NANDN U13529 ( .A(n13148), .B(n13147), .Z(n13149) );
  NAND U13530 ( .A(n13150), .B(n13149), .Z(n13262) );
  NANDN U13531 ( .A(n13152), .B(n13151), .Z(n13156) );
  NAND U13532 ( .A(n13154), .B(n13153), .Z(n13155) );
  NAND U13533 ( .A(n13156), .B(n13155), .Z(n13264) );
  XNOR U13534 ( .A(n13190), .B(n13189), .Z(n13191) );
  XOR U13535 ( .A(n13192), .B(n13191), .Z(n13186) );
  NANDN U13536 ( .A(n13158), .B(n13157), .Z(n13162) );
  NANDN U13537 ( .A(n13160), .B(n13159), .Z(n13161) );
  AND U13538 ( .A(n13162), .B(n13161), .Z(n13184) );
  NAND U13539 ( .A(n13164), .B(n13163), .Z(n13168) );
  NANDN U13540 ( .A(n13166), .B(n13165), .Z(n13167) );
  NAND U13541 ( .A(n13168), .B(n13167), .Z(n13183) );
  XNOR U13542 ( .A(n13184), .B(n13183), .Z(n13185) );
  XNOR U13543 ( .A(n13186), .B(n13185), .Z(n13292) );
  XOR U13544 ( .A(n13293), .B(n13292), .Z(n13294) );
  XNOR U13545 ( .A(n13295), .B(n13294), .Z(n13288) );
  OR U13546 ( .A(n13171), .B(n13169), .Z(n13175) );
  ANDN U13547 ( .B(n13171), .A(n13170), .Z(n13173) );
  OR U13548 ( .A(n13173), .B(n13172), .Z(n13174) );
  AND U13549 ( .A(n13175), .B(n13174), .Z(n13287) );
  NAND U13550 ( .A(n13177), .B(n13176), .Z(n13181) );
  NANDN U13551 ( .A(n13179), .B(n13178), .Z(n13180) );
  NAND U13552 ( .A(n13181), .B(n13180), .Z(n13286) );
  IV U13553 ( .A(n13286), .Z(n13285) );
  XOR U13554 ( .A(n13287), .B(n13285), .Z(n13182) );
  XNOR U13555 ( .A(n13288), .B(n13182), .Z(N307) );
  NANDN U13556 ( .A(n13184), .B(n13183), .Z(n13188) );
  NANDN U13557 ( .A(n13186), .B(n13185), .Z(n13187) );
  AND U13558 ( .A(n13188), .B(n13187), .Z(n13407) );
  NANDN U13559 ( .A(n13190), .B(n13189), .Z(n13194) );
  NAND U13560 ( .A(n13192), .B(n13191), .Z(n13193) );
  AND U13561 ( .A(n13194), .B(n13193), .Z(n13405) );
  NANDN U13562 ( .A(n13196), .B(n13195), .Z(n13200) );
  NANDN U13563 ( .A(n13198), .B(n13197), .Z(n13199) );
  NAND U13564 ( .A(n13200), .B(n13199), .Z(n13381) );
  AND U13565 ( .A(x[134]), .B(y[781]), .Z(n13247) );
  NAND U13566 ( .A(n13247), .B(n13201), .Z(n13205) );
  NAND U13567 ( .A(n13203), .B(n13202), .Z(n13204) );
  NAND U13568 ( .A(n13205), .B(n13204), .Z(n13375) );
  AND U13569 ( .A(x[144]), .B(y[775]), .Z(n13206) );
  NAND U13570 ( .A(n13563), .B(n13206), .Z(n13210) );
  NAND U13571 ( .A(n13208), .B(n13207), .Z(n13209) );
  NAND U13572 ( .A(n13210), .B(n13209), .Z(n13373) );
  AND U13573 ( .A(x[143]), .B(y[777]), .Z(n13949) );
  NAND U13574 ( .A(n13311), .B(n13949), .Z(n13214) );
  NAND U13575 ( .A(n13212), .B(n13211), .Z(n13213) );
  NAND U13576 ( .A(n13214), .B(n13213), .Z(n13301) );
  AND U13577 ( .A(y[786]), .B(x[129]), .Z(n13216) );
  NAND U13578 ( .A(y[779]), .B(x[136]), .Z(n13215) );
  XNOR U13579 ( .A(n13216), .B(n13215), .Z(n13343) );
  XNOR U13580 ( .A(n13343), .B(n13344), .Z(n13300) );
  AND U13581 ( .A(y[785]), .B(x[130]), .Z(n13218) );
  NAND U13582 ( .A(y[774]), .B(x[141]), .Z(n13217) );
  XNOR U13583 ( .A(n13218), .B(n13217), .Z(n13316) );
  XOR U13584 ( .A(n13316), .B(n13315), .Z(n13299) );
  XOR U13585 ( .A(n13300), .B(n13299), .Z(n13302) );
  XOR U13586 ( .A(n13301), .B(n13302), .Z(n13374) );
  XOR U13587 ( .A(n13373), .B(n13374), .Z(n13376) );
  XOR U13588 ( .A(n13375), .B(n13376), .Z(n13380) );
  AND U13589 ( .A(x[138]), .B(y[785]), .Z(n14334) );
  NAND U13590 ( .A(n14334), .B(n13219), .Z(n13223) );
  NAND U13591 ( .A(n13221), .B(n13220), .Z(n13222) );
  NAND U13592 ( .A(n13223), .B(n13222), .Z(n13351) );
  NAND U13593 ( .A(n13225), .B(n13224), .Z(n13229) );
  NAND U13594 ( .A(n13227), .B(n13226), .Z(n13228) );
  NAND U13595 ( .A(n13229), .B(n13228), .Z(n13349) );
  AND U13596 ( .A(y[778]), .B(x[137]), .Z(n13231) );
  NAND U13597 ( .A(y[771]), .B(x[144]), .Z(n13230) );
  XNOR U13598 ( .A(n13231), .B(n13230), .Z(n13313) );
  AND U13599 ( .A(x[143]), .B(y[772]), .Z(n13312) );
  XOR U13600 ( .A(n13313), .B(n13312), .Z(n13350) );
  XOR U13601 ( .A(n13349), .B(n13350), .Z(n13352) );
  XOR U13602 ( .A(n13351), .B(n13352), .Z(n13370) );
  AND U13603 ( .A(x[141]), .B(y[783]), .Z(n14548) );
  NANDN U13604 ( .A(n13232), .B(n14548), .Z(n13236) );
  NAND U13605 ( .A(n13234), .B(n13233), .Z(n13235) );
  NAND U13606 ( .A(n13236), .B(n13235), .Z(n13357) );
  AND U13607 ( .A(y[770]), .B(x[145]), .Z(n13238) );
  NAND U13608 ( .A(y[777]), .B(x[138]), .Z(n13237) );
  XNOR U13609 ( .A(n13238), .B(n13237), .Z(n13348) );
  AND U13610 ( .A(x[146]), .B(y[769]), .Z(n13329) );
  XOR U13611 ( .A(n13329), .B(o[147]), .Z(n13347) );
  XOR U13612 ( .A(n13348), .B(n13347), .Z(n13356) );
  AND U13613 ( .A(y[784]), .B(x[131]), .Z(n13240) );
  NAND U13614 ( .A(y[776]), .B(x[139]), .Z(n13239) );
  XNOR U13615 ( .A(n13240), .B(n13239), .Z(n13324) );
  XOR U13616 ( .A(n13324), .B(n13323), .Z(n13355) );
  XOR U13617 ( .A(n13356), .B(n13355), .Z(n13358) );
  XOR U13618 ( .A(n13357), .B(n13358), .Z(n13368) );
  NAND U13619 ( .A(n13241), .B(n13611), .Z(n13245) );
  NAND U13620 ( .A(n13243), .B(n13242), .Z(n13244) );
  NAND U13621 ( .A(n13245), .B(n13244), .Z(n13307) );
  AND U13622 ( .A(x[128]), .B(y[787]), .Z(n13333) );
  AND U13623 ( .A(x[147]), .B(y[768]), .Z(n13332) );
  XOR U13624 ( .A(n13333), .B(n13332), .Z(n13334) );
  XOR U13625 ( .A(n13334), .B(n13335), .Z(n13306) );
  AND U13626 ( .A(x[132]), .B(y[783]), .Z(n13469) );
  AND U13627 ( .A(y[782]), .B(x[133]), .Z(n13248) );
  XOR U13628 ( .A(n13248), .B(n13247), .Z(n13331) );
  XOR U13629 ( .A(n13469), .B(n13331), .Z(n13305) );
  XOR U13630 ( .A(n13306), .B(n13305), .Z(n13308) );
  XNOR U13631 ( .A(n13307), .B(n13308), .Z(n13367) );
  NAND U13632 ( .A(n13250), .B(n13249), .Z(n13254) );
  NAND U13633 ( .A(n13252), .B(n13251), .Z(n13253) );
  NAND U13634 ( .A(n13254), .B(n13253), .Z(n13362) );
  NAND U13635 ( .A(n13256), .B(n13255), .Z(n13260) );
  NAND U13636 ( .A(n13258), .B(n13257), .Z(n13259) );
  NAND U13637 ( .A(n13260), .B(n13259), .Z(n13361) );
  XOR U13638 ( .A(n13362), .B(n13361), .Z(n13363) );
  XNOR U13639 ( .A(n13364), .B(n13363), .Z(n13379) );
  XOR U13640 ( .A(n13381), .B(n13382), .Z(n13393) );
  NANDN U13641 ( .A(n13262), .B(n13261), .Z(n13266) );
  NANDN U13642 ( .A(n13264), .B(n13263), .Z(n13265) );
  AND U13643 ( .A(n13266), .B(n13265), .Z(n13392) );
  NANDN U13644 ( .A(n13268), .B(n13267), .Z(n13272) );
  NAND U13645 ( .A(n13270), .B(n13269), .Z(n13271) );
  AND U13646 ( .A(n13272), .B(n13271), .Z(n13388) );
  NANDN U13647 ( .A(n13274), .B(n13273), .Z(n13278) );
  NAND U13648 ( .A(n13276), .B(n13275), .Z(n13277) );
  AND U13649 ( .A(n13278), .B(n13277), .Z(n13386) );
  NANDN U13650 ( .A(n13280), .B(n13279), .Z(n13284) );
  NAND U13651 ( .A(n13282), .B(n13281), .Z(n13283) );
  NAND U13652 ( .A(n13284), .B(n13283), .Z(n13385) );
  XOR U13653 ( .A(n13392), .B(n13391), .Z(n13394) );
  XOR U13654 ( .A(n13393), .B(n13394), .Z(n13404) );
  XOR U13655 ( .A(n13405), .B(n13404), .Z(n13406) );
  XOR U13656 ( .A(n13407), .B(n13406), .Z(n13400) );
  OR U13657 ( .A(n13287), .B(n13285), .Z(n13291) );
  ANDN U13658 ( .B(n13287), .A(n13286), .Z(n13289) );
  OR U13659 ( .A(n13289), .B(n13288), .Z(n13290) );
  AND U13660 ( .A(n13291), .B(n13290), .Z(n13399) );
  NAND U13661 ( .A(n13293), .B(n13292), .Z(n13297) );
  NAND U13662 ( .A(n13295), .B(n13294), .Z(n13296) );
  NAND U13663 ( .A(n13297), .B(n13296), .Z(n13398) );
  IV U13664 ( .A(n13398), .Z(n13397) );
  XOR U13665 ( .A(n13399), .B(n13397), .Z(n13298) );
  XNOR U13666 ( .A(n13400), .B(n13298), .Z(N308) );
  NAND U13667 ( .A(n13300), .B(n13299), .Z(n13304) );
  NAND U13668 ( .A(n13302), .B(n13301), .Z(n13303) );
  NAND U13669 ( .A(n13304), .B(n13303), .Z(n13412) );
  NAND U13670 ( .A(n13306), .B(n13305), .Z(n13310) );
  NAND U13671 ( .A(n13308), .B(n13307), .Z(n13309) );
  NAND U13672 ( .A(n13310), .B(n13309), .Z(n13411) );
  XOR U13673 ( .A(n13412), .B(n13411), .Z(n13414) );
  AND U13674 ( .A(x[144]), .B(y[778]), .Z(n14208) );
  AND U13675 ( .A(x[141]), .B(y[785]), .Z(n14775) );
  NAND U13676 ( .A(n14775), .B(n13314), .Z(n13318) );
  NAND U13677 ( .A(n13316), .B(n13315), .Z(n13317) );
  NAND U13678 ( .A(n13318), .B(n13317), .Z(n13486) );
  NAND U13679 ( .A(y[772]), .B(x[144]), .Z(n13319) );
  XNOR U13680 ( .A(n13320), .B(n13319), .Z(n13450) );
  NAND U13681 ( .A(x[130]), .B(y[786]), .Z(n13451) );
  XNOR U13682 ( .A(n13450), .B(n13451), .Z(n13485) );
  NAND U13683 ( .A(y[773]), .B(x[143]), .Z(n13321) );
  XNOR U13684 ( .A(n13322), .B(n13321), .Z(n13427) );
  AND U13685 ( .A(x[142]), .B(y[774]), .Z(n13426) );
  XOR U13686 ( .A(n13427), .B(n13426), .Z(n13484) );
  XOR U13687 ( .A(n13485), .B(n13484), .Z(n13487) );
  XOR U13688 ( .A(n13486), .B(n13487), .Z(n13446) );
  XOR U13689 ( .A(n13445), .B(n13446), .Z(n13448) );
  AND U13690 ( .A(x[139]), .B(y[784]), .Z(n14337) );
  NANDN U13691 ( .A(n13590), .B(n14337), .Z(n13326) );
  NAND U13692 ( .A(n13324), .B(n13323), .Z(n13325) );
  NAND U13693 ( .A(n13326), .B(n13325), .Z(n13490) );
  AND U13694 ( .A(y[787]), .B(x[129]), .Z(n13328) );
  NAND U13695 ( .A(y[777]), .B(x[139]), .Z(n13327) );
  XNOR U13696 ( .A(n13328), .B(n13327), .Z(n13424) );
  NAND U13697 ( .A(x[147]), .B(y[769]), .Z(n13430) );
  XNOR U13698 ( .A(o[148]), .B(n13430), .Z(n13423) );
  XOR U13699 ( .A(n13424), .B(n13423), .Z(n13489) );
  AND U13700 ( .A(n13329), .B(o[147]), .Z(n13477) );
  AND U13701 ( .A(x[128]), .B(y[788]), .Z(n13474) );
  NAND U13702 ( .A(x[148]), .B(y[768]), .Z(n13475) );
  XNOR U13703 ( .A(n13474), .B(n13475), .Z(n13476) );
  XOR U13704 ( .A(n13477), .B(n13476), .Z(n13488) );
  XOR U13705 ( .A(n13489), .B(n13488), .Z(n13491) );
  XOR U13706 ( .A(n13490), .B(n13491), .Z(n13447) );
  XOR U13707 ( .A(n13448), .B(n13447), .Z(n13413) );
  XOR U13708 ( .A(n13414), .B(n13413), .Z(n13495) );
  NAND U13709 ( .A(x[134]), .B(y[782]), .Z(n13431) );
  AND U13710 ( .A(y[770]), .B(x[146]), .Z(n13337) );
  NAND U13711 ( .A(y[776]), .B(x[140]), .Z(n13336) );
  XNOR U13712 ( .A(n13337), .B(n13336), .Z(n13418) );
  NAND U13713 ( .A(x[145]), .B(y[771]), .Z(n13419) );
  XNOR U13714 ( .A(n13418), .B(n13419), .Z(n13436) );
  XOR U13715 ( .A(n13435), .B(n13436), .Z(n13438) );
  XOR U13716 ( .A(n13437), .B(n13438), .Z(n13440) );
  AND U13717 ( .A(y[785]), .B(x[131]), .Z(n13339) );
  NAND U13718 ( .A(y[775]), .B(x[141]), .Z(n13338) );
  XNOR U13719 ( .A(n13339), .B(n13338), .Z(n13455) );
  AND U13720 ( .A(y[783]), .B(x[133]), .Z(n13341) );
  NAND U13721 ( .A(y[784]), .B(x[132]), .Z(n13340) );
  XNOR U13722 ( .A(n13341), .B(n13340), .Z(n13471) );
  AND U13723 ( .A(x[135]), .B(y[781]), .Z(n13470) );
  XNOR U13724 ( .A(n13471), .B(n13470), .Z(n13432) );
  XOR U13725 ( .A(n13431), .B(n13432), .Z(n13433) );
  XOR U13726 ( .A(n13434), .B(n13433), .Z(n13482) );
  AND U13727 ( .A(x[136]), .B(y[786]), .Z(n14501) );
  NAND U13728 ( .A(n14501), .B(n13342), .Z(n13346) );
  NANDN U13729 ( .A(n13344), .B(n13343), .Z(n13345) );
  NAND U13730 ( .A(n13346), .B(n13345), .Z(n13480) );
  AND U13731 ( .A(x[145]), .B(y[777]), .Z(n14214) );
  XNOR U13732 ( .A(n13480), .B(n13481), .Z(n13483) );
  XOR U13733 ( .A(n13482), .B(n13483), .Z(n13439) );
  XNOR U13734 ( .A(n13440), .B(n13439), .Z(n13442) );
  NAND U13735 ( .A(n13350), .B(n13349), .Z(n13354) );
  NAND U13736 ( .A(n13352), .B(n13351), .Z(n13353) );
  AND U13737 ( .A(n13354), .B(n13353), .Z(n13441) );
  XOR U13738 ( .A(n13442), .B(n13441), .Z(n13493) );
  NAND U13739 ( .A(n13356), .B(n13355), .Z(n13360) );
  NAND U13740 ( .A(n13358), .B(n13357), .Z(n13359) );
  AND U13741 ( .A(n13360), .B(n13359), .Z(n13492) );
  XOR U13742 ( .A(n13493), .B(n13492), .Z(n13494) );
  XNOR U13743 ( .A(n13495), .B(n13494), .Z(n13499) );
  NAND U13744 ( .A(n13362), .B(n13361), .Z(n13366) );
  NAND U13745 ( .A(n13364), .B(n13363), .Z(n13365) );
  AND U13746 ( .A(n13366), .B(n13365), .Z(n13507) );
  NANDN U13747 ( .A(n13368), .B(n13367), .Z(n13372) );
  NANDN U13748 ( .A(n13370), .B(n13369), .Z(n13371) );
  NAND U13749 ( .A(n13372), .B(n13371), .Z(n13504) );
  NAND U13750 ( .A(n13374), .B(n13373), .Z(n13378) );
  NAND U13751 ( .A(n13376), .B(n13375), .Z(n13377) );
  AND U13752 ( .A(n13378), .B(n13377), .Z(n13505) );
  XOR U13753 ( .A(n13504), .B(n13505), .Z(n13506) );
  XNOR U13754 ( .A(n13507), .B(n13506), .Z(n13498) );
  NANDN U13755 ( .A(n13380), .B(n13379), .Z(n13384) );
  NANDN U13756 ( .A(n13382), .B(n13381), .Z(n13383) );
  AND U13757 ( .A(n13384), .B(n13383), .Z(n13500) );
  XOR U13758 ( .A(n13501), .B(n13500), .Z(n13513) );
  NANDN U13759 ( .A(n13386), .B(n13385), .Z(n13390) );
  NANDN U13760 ( .A(n13388), .B(n13387), .Z(n13389) );
  AND U13761 ( .A(n13390), .B(n13389), .Z(n13510) );
  NAND U13762 ( .A(n13392), .B(n13391), .Z(n13396) );
  NAND U13763 ( .A(n13394), .B(n13393), .Z(n13395) );
  NAND U13764 ( .A(n13396), .B(n13395), .Z(n13511) );
  XOR U13765 ( .A(n13513), .B(n13512), .Z(n13519) );
  OR U13766 ( .A(n13399), .B(n13397), .Z(n13403) );
  ANDN U13767 ( .B(n13399), .A(n13398), .Z(n13401) );
  OR U13768 ( .A(n13401), .B(n13400), .Z(n13402) );
  AND U13769 ( .A(n13403), .B(n13402), .Z(n13517) );
  NAND U13770 ( .A(n13405), .B(n13404), .Z(n13409) );
  NANDN U13771 ( .A(n13407), .B(n13406), .Z(n13408) );
  AND U13772 ( .A(n13409), .B(n13408), .Z(n13518) );
  IV U13773 ( .A(n13518), .Z(n13516) );
  XOR U13774 ( .A(n13517), .B(n13516), .Z(n13410) );
  XNOR U13775 ( .A(n13519), .B(n13410), .Z(N309) );
  NAND U13776 ( .A(n13412), .B(n13411), .Z(n13416) );
  NAND U13777 ( .A(n13414), .B(n13413), .Z(n13415) );
  NAND U13778 ( .A(n13416), .B(n13415), .Z(n13541) );
  NAND U13779 ( .A(x[146]), .B(y[776]), .Z(n14217) );
  NANDN U13780 ( .A(n14217), .B(n13417), .Z(n13421) );
  NANDN U13781 ( .A(n13419), .B(n13418), .Z(n13420) );
  AND U13782 ( .A(n13421), .B(n13420), .Z(n13617) );
  AND U13783 ( .A(x[139]), .B(y[787]), .Z(n14835) );
  XNOR U13784 ( .A(n13617), .B(n13616), .Z(n13619) );
  AND U13785 ( .A(x[143]), .B(y[779]), .Z(n14203) );
  NAND U13786 ( .A(n14203), .B(n13425), .Z(n13429) );
  NAND U13787 ( .A(n13427), .B(n13426), .Z(n13428) );
  AND U13788 ( .A(n13429), .B(n13428), .Z(n13577) );
  ANDN U13789 ( .B(o[148]), .A(n13430), .Z(n13599) );
  AND U13790 ( .A(x[128]), .B(y[789]), .Z(n13596) );
  NAND U13791 ( .A(x[149]), .B(y[768]), .Z(n13597) );
  XNOR U13792 ( .A(n13596), .B(n13597), .Z(n13598) );
  XOR U13793 ( .A(n13599), .B(n13598), .Z(n13575) );
  AND U13794 ( .A(x[133]), .B(y[784]), .Z(n13581) );
  AND U13795 ( .A(x[144]), .B(y[773]), .Z(n13580) );
  XOR U13796 ( .A(n13581), .B(n13580), .Z(n13583) );
  NAND U13797 ( .A(x[143]), .B(y[774]), .Z(n13582) );
  XNOR U13798 ( .A(n13583), .B(n13582), .Z(n13574) );
  XOR U13799 ( .A(n13575), .B(n13574), .Z(n13576) );
  XNOR U13800 ( .A(n13577), .B(n13576), .Z(n13618) );
  XOR U13801 ( .A(n13619), .B(n13618), .Z(n13613) );
  XNOR U13802 ( .A(n13613), .B(n13612), .Z(n13615) );
  XOR U13803 ( .A(n13615), .B(n13614), .Z(n13540) );
  NANDN U13804 ( .A(n13440), .B(n13439), .Z(n13444) );
  NAND U13805 ( .A(n13442), .B(n13441), .Z(n13443) );
  AND U13806 ( .A(n13444), .B(n13443), .Z(n13539) );
  XNOR U13807 ( .A(n13540), .B(n13539), .Z(n13542) );
  XOR U13808 ( .A(n13541), .B(n13542), .Z(n13536) );
  NAND U13809 ( .A(n14208), .B(n13449), .Z(n13453) );
  NANDN U13810 ( .A(n13451), .B(n13450), .Z(n13452) );
  AND U13811 ( .A(n13453), .B(n13452), .Z(n13546) );
  AND U13812 ( .A(x[131]), .B(y[775]), .Z(n13454) );
  NAND U13813 ( .A(n14775), .B(n13454), .Z(n13458) );
  NANDN U13814 ( .A(n13456), .B(n13455), .Z(n13457) );
  AND U13815 ( .A(n13458), .B(n13457), .Z(n13629) );
  AND U13816 ( .A(y[770]), .B(x[147]), .Z(n13460) );
  NAND U13817 ( .A(y[778]), .B(x[139]), .Z(n13459) );
  XNOR U13818 ( .A(n13460), .B(n13459), .Z(n13564) );
  NAND U13819 ( .A(x[148]), .B(y[769]), .Z(n13595) );
  XOR U13820 ( .A(o[149]), .B(n13595), .Z(n13565) );
  XNOR U13821 ( .A(n13564), .B(n13565), .Z(n13627) );
  AND U13822 ( .A(y[771]), .B(x[146]), .Z(n13462) );
  NAND U13823 ( .A(y[779]), .B(x[138]), .Z(n13461) );
  XNOR U13824 ( .A(n13462), .B(n13461), .Z(n13603) );
  NAND U13825 ( .A(x[129]), .B(y[788]), .Z(n13604) );
  XNOR U13826 ( .A(n13603), .B(n13604), .Z(n13626) );
  XOR U13827 ( .A(n13627), .B(n13626), .Z(n13628) );
  XNOR U13828 ( .A(n13629), .B(n13628), .Z(n13545) );
  XNOR U13829 ( .A(n13546), .B(n13545), .Z(n13547) );
  AND U13830 ( .A(x[135]), .B(y[782]), .Z(n13770) );
  AND U13831 ( .A(y[775]), .B(x[142]), .Z(n13464) );
  NAND U13832 ( .A(y[783]), .B(x[134]), .Z(n13463) );
  XNOR U13833 ( .A(n13464), .B(n13463), .Z(n13607) );
  XOR U13834 ( .A(n13770), .B(n13607), .Z(n13554) );
  AND U13835 ( .A(x[137]), .B(y[780]), .Z(n13552) );
  NAND U13836 ( .A(x[136]), .B(y[781]), .Z(n13551) );
  XNOR U13837 ( .A(n13552), .B(n13551), .Z(n13553) );
  XOR U13838 ( .A(n13554), .B(n13553), .Z(n13570) );
  AND U13839 ( .A(y[772]), .B(x[145]), .Z(n13466) );
  NAND U13840 ( .A(y[777]), .B(x[140]), .Z(n13465) );
  XNOR U13841 ( .A(n13466), .B(n13465), .Z(n13557) );
  NAND U13842 ( .A(x[130]), .B(y[787]), .Z(n13558) );
  XNOR U13843 ( .A(n13557), .B(n13558), .Z(n13569) );
  AND U13844 ( .A(y[786]), .B(x[131]), .Z(n13468) );
  NAND U13845 ( .A(y[776]), .B(x[141]), .Z(n13467) );
  XNOR U13846 ( .A(n13468), .B(n13467), .Z(n13591) );
  NAND U13847 ( .A(x[132]), .B(y[785]), .Z(n13592) );
  XNOR U13848 ( .A(n13591), .B(n13592), .Z(n13568) );
  XOR U13849 ( .A(n13569), .B(n13568), .Z(n13571) );
  XOR U13850 ( .A(n13570), .B(n13571), .Z(n13622) );
  NAND U13851 ( .A(n13581), .B(n13469), .Z(n13473) );
  NAND U13852 ( .A(n13471), .B(n13470), .Z(n13472) );
  AND U13853 ( .A(n13473), .B(n13472), .Z(n13621) );
  NANDN U13854 ( .A(n13475), .B(n13474), .Z(n13479) );
  NAND U13855 ( .A(n13477), .B(n13476), .Z(n13478) );
  NAND U13856 ( .A(n13479), .B(n13478), .Z(n13620) );
  XOR U13857 ( .A(n13621), .B(n13620), .Z(n13623) );
  XOR U13858 ( .A(n13622), .B(n13623), .Z(n13548) );
  XNOR U13859 ( .A(n13547), .B(n13548), .Z(n13630) );
  XNOR U13860 ( .A(n13635), .B(n13634), .Z(n13637) );
  XNOR U13861 ( .A(n13630), .B(n13631), .Z(n13633) );
  XOR U13862 ( .A(n13632), .B(n13633), .Z(n13534) );
  NAND U13863 ( .A(n13493), .B(n13492), .Z(n13497) );
  NANDN U13864 ( .A(n13495), .B(n13494), .Z(n13496) );
  NAND U13865 ( .A(n13497), .B(n13496), .Z(n13533) );
  XNOR U13866 ( .A(n13534), .B(n13533), .Z(n13535) );
  XNOR U13867 ( .A(n13536), .B(n13535), .Z(n13527) );
  NANDN U13868 ( .A(n13499), .B(n13498), .Z(n13503) );
  NAND U13869 ( .A(n13501), .B(n13500), .Z(n13502) );
  NAND U13870 ( .A(n13503), .B(n13502), .Z(n13524) );
  NAND U13871 ( .A(n13505), .B(n13504), .Z(n13509) );
  NAND U13872 ( .A(n13507), .B(n13506), .Z(n13508) );
  AND U13873 ( .A(n13509), .B(n13508), .Z(n13525) );
  XOR U13874 ( .A(n13524), .B(n13525), .Z(n13526) );
  NANDN U13875 ( .A(n13511), .B(n13510), .Z(n13515) );
  NANDN U13876 ( .A(n13513), .B(n13512), .Z(n13514) );
  NAND U13877 ( .A(n13515), .B(n13514), .Z(n13530) );
  NANDN U13878 ( .A(n13516), .B(n13517), .Z(n13522) );
  NOR U13879 ( .A(n13518), .B(n13517), .Z(n13520) );
  OR U13880 ( .A(n13520), .B(n13519), .Z(n13521) );
  AND U13881 ( .A(n13522), .B(n13521), .Z(n13531) );
  XOR U13882 ( .A(n13530), .B(n13531), .Z(n13523) );
  XNOR U13883 ( .A(n13532), .B(n13523), .Z(N310) );
  NAND U13884 ( .A(n13525), .B(n13524), .Z(n13529) );
  NANDN U13885 ( .A(n13527), .B(n13526), .Z(n13528) );
  AND U13886 ( .A(n13529), .B(n13528), .Z(n13745) );
  NANDN U13887 ( .A(n13534), .B(n13533), .Z(n13538) );
  NANDN U13888 ( .A(n13536), .B(n13535), .Z(n13537) );
  AND U13889 ( .A(n13538), .B(n13537), .Z(n13750) );
  NANDN U13890 ( .A(n13540), .B(n13539), .Z(n13544) );
  NAND U13891 ( .A(n13542), .B(n13541), .Z(n13543) );
  NAND U13892 ( .A(n13544), .B(n13543), .Z(n13748) );
  NANDN U13893 ( .A(n13546), .B(n13545), .Z(n13550) );
  NANDN U13894 ( .A(n13548), .B(n13547), .Z(n13549) );
  AND U13895 ( .A(n13550), .B(n13549), .Z(n13744) );
  NANDN U13896 ( .A(n13552), .B(n13551), .Z(n13556) );
  NANDN U13897 ( .A(n13554), .B(n13553), .Z(n13555) );
  AND U13898 ( .A(n13556), .B(n13555), .Z(n13738) );
  NAND U13899 ( .A(n14214), .B(n13692), .Z(n13560) );
  NANDN U13900 ( .A(n13558), .B(n13557), .Z(n13559) );
  NAND U13901 ( .A(n13560), .B(n13559), .Z(n13673) );
  AND U13902 ( .A(x[133]), .B(y[785]), .Z(n13713) );
  NAND U13903 ( .A(x[145]), .B(y[773]), .Z(n13714) );
  XNOR U13904 ( .A(n13713), .B(n13714), .Z(n13715) );
  NAND U13905 ( .A(x[144]), .B(y[774]), .Z(n13716) );
  XNOR U13906 ( .A(n13715), .B(n13716), .Z(n13672) );
  AND U13907 ( .A(y[772]), .B(x[146]), .Z(n13562) );
  NAND U13908 ( .A(y[778]), .B(x[140]), .Z(n13561) );
  XNOR U13909 ( .A(n13562), .B(n13561), .Z(n13693) );
  NAND U13910 ( .A(x[132]), .B(y[786]), .Z(n13694) );
  XNOR U13911 ( .A(n13693), .B(n13694), .Z(n13671) );
  XOR U13912 ( .A(n13672), .B(n13671), .Z(n13674) );
  XNOR U13913 ( .A(n13673), .B(n13674), .Z(n13736) );
  AND U13914 ( .A(x[147]), .B(y[778]), .Z(n14668) );
  NAND U13915 ( .A(n14668), .B(n13563), .Z(n13567) );
  NANDN U13916 ( .A(n13565), .B(n13564), .Z(n13566) );
  AND U13917 ( .A(n13567), .B(n13566), .Z(n13735) );
  XOR U13918 ( .A(n13736), .B(n13735), .Z(n13737) );
  XOR U13919 ( .A(n13738), .B(n13737), .Z(n13741) );
  NAND U13920 ( .A(n13569), .B(n13568), .Z(n13573) );
  NAND U13921 ( .A(n13571), .B(n13570), .Z(n13572) );
  AND U13922 ( .A(n13573), .B(n13572), .Z(n13726) );
  NAND U13923 ( .A(n13575), .B(n13574), .Z(n13579) );
  NANDN U13924 ( .A(n13577), .B(n13576), .Z(n13578) );
  NAND U13925 ( .A(n13579), .B(n13578), .Z(n13725) );
  XNOR U13926 ( .A(n13726), .B(n13725), .Z(n13728) );
  NAND U13927 ( .A(n13581), .B(n13580), .Z(n13585) );
  ANDN U13928 ( .B(n13583), .A(n13582), .Z(n13584) );
  ANDN U13929 ( .B(n13585), .A(n13584), .Z(n13691) );
  AND U13930 ( .A(y[770]), .B(x[148]), .Z(n13587) );
  NAND U13931 ( .A(y[777]), .B(x[141]), .Z(n13586) );
  XNOR U13932 ( .A(n13587), .B(n13586), .Z(n13709) );
  NAND U13933 ( .A(x[130]), .B(y[788]), .Z(n13710) );
  XNOR U13934 ( .A(n13709), .B(n13710), .Z(n13689) );
  AND U13935 ( .A(y[784]), .B(x[134]), .Z(n13589) );
  NAND U13936 ( .A(y[775]), .B(x[143]), .Z(n13588) );
  XNOR U13937 ( .A(n13589), .B(n13588), .Z(n13721) );
  XOR U13938 ( .A(n13689), .B(n13688), .Z(n13690) );
  XNOR U13939 ( .A(n13691), .B(n13690), .Z(n13729) );
  AND U13940 ( .A(x[141]), .B(y[786]), .Z(n14919) );
  NANDN U13941 ( .A(n13590), .B(n14919), .Z(n13594) );
  NANDN U13942 ( .A(n13592), .B(n13591), .Z(n13593) );
  AND U13943 ( .A(n13594), .B(n13593), .Z(n13662) );
  ANDN U13944 ( .B(o[149]), .A(n13595), .Z(n13684) );
  AND U13945 ( .A(x[129]), .B(y[789]), .Z(n13685) );
  XOR U13946 ( .A(n13686), .B(n13685), .Z(n13683) );
  XOR U13947 ( .A(n13684), .B(n13683), .Z(n13659) );
  AND U13948 ( .A(x[142]), .B(y[776]), .Z(n13677) );
  NAND U13949 ( .A(x[131]), .B(y[787]), .Z(n13678) );
  XNOR U13950 ( .A(n13677), .B(n13678), .Z(n13679) );
  NAND U13951 ( .A(x[147]), .B(y[771]), .Z(n13680) );
  XOR U13952 ( .A(n13679), .B(n13680), .Z(n13660) );
  XNOR U13953 ( .A(n13659), .B(n13660), .Z(n13661) );
  XOR U13954 ( .A(n13662), .B(n13661), .Z(n13730) );
  XNOR U13955 ( .A(n13729), .B(n13730), .Z(n13732) );
  NANDN U13956 ( .A(n13597), .B(n13596), .Z(n13601) );
  NAND U13957 ( .A(n13599), .B(n13598), .Z(n13600) );
  AND U13958 ( .A(n13601), .B(n13600), .Z(n13656) );
  AND U13959 ( .A(x[146]), .B(y[779]), .Z(n14671) );
  NAND U13960 ( .A(n14671), .B(n13602), .Z(n13606) );
  NANDN U13961 ( .A(n13604), .B(n13603), .Z(n13605) );
  NAND U13962 ( .A(n13606), .B(n13605), .Z(n13655) );
  XNOR U13963 ( .A(n13656), .B(n13655), .Z(n13658) );
  AND U13964 ( .A(x[142]), .B(y[783]), .Z(n14687) );
  NAND U13965 ( .A(n14687), .B(n13720), .Z(n13609) );
  NAND U13966 ( .A(n13770), .B(n13607), .Z(n13608) );
  AND U13967 ( .A(n13609), .B(n13608), .Z(n13668) );
  AND U13968 ( .A(x[128]), .B(y[790]), .Z(n13697) );
  NAND U13969 ( .A(x[150]), .B(y[768]), .Z(n13698) );
  XNOR U13970 ( .A(n13697), .B(n13698), .Z(n13700) );
  AND U13971 ( .A(x[149]), .B(y[769]), .Z(n13719) );
  XOR U13972 ( .A(o[150]), .B(n13719), .Z(n13699) );
  XOR U13973 ( .A(n13700), .B(n13699), .Z(n13666) );
  NAND U13974 ( .A(y[783]), .B(x[135]), .Z(n13610) );
  XNOR U13975 ( .A(n13611), .B(n13610), .Z(n13703) );
  XOR U13976 ( .A(n13666), .B(n13665), .Z(n13667) );
  XNOR U13977 ( .A(n13668), .B(n13667), .Z(n13657) );
  XOR U13978 ( .A(n13658), .B(n13657), .Z(n13731) );
  XOR U13979 ( .A(n13732), .B(n13731), .Z(n13727) );
  XOR U13980 ( .A(n13728), .B(n13727), .Z(n13742) );
  XOR U13981 ( .A(n13741), .B(n13742), .Z(n13743) );
  XOR U13982 ( .A(n13744), .B(n13743), .Z(n13647) );
  NANDN U13983 ( .A(n13621), .B(n13620), .Z(n13625) );
  NANDN U13984 ( .A(n13623), .B(n13622), .Z(n13624) );
  AND U13985 ( .A(n13625), .B(n13624), .Z(n13650) );
  XOR U13986 ( .A(n13650), .B(n13649), .Z(n13652) );
  XNOR U13987 ( .A(n13651), .B(n13652), .Z(n13646) );
  XOR U13988 ( .A(n13645), .B(n13646), .Z(n13648) );
  XOR U13989 ( .A(n13647), .B(n13648), .Z(n13643) );
  NAND U13990 ( .A(n13635), .B(n13634), .Z(n13639) );
  NANDN U13991 ( .A(n13637), .B(n13636), .Z(n13638) );
  NAND U13992 ( .A(n13639), .B(n13638), .Z(n13642) );
  XNOR U13993 ( .A(n13641), .B(n13642), .Z(n13644) );
  XOR U13994 ( .A(n13643), .B(n13644), .Z(n13749) );
  XNOR U13995 ( .A(n13748), .B(n13749), .Z(n13751) );
  XNOR U13996 ( .A(n13750), .B(n13751), .Z(n13747) );
  XNOR U13997 ( .A(n13746), .B(n13747), .Z(n13640) );
  XOR U13998 ( .A(n13745), .B(n13640), .Z(N311) );
  NANDN U13999 ( .A(n13650), .B(n13649), .Z(n13654) );
  OR U14000 ( .A(n13652), .B(n13651), .Z(n13653) );
  AND U14001 ( .A(n13654), .B(n13653), .Z(n13850) );
  NANDN U14002 ( .A(n13660), .B(n13659), .Z(n13664) );
  NANDN U14003 ( .A(n13662), .B(n13661), .Z(n13663) );
  AND U14004 ( .A(n13664), .B(n13663), .Z(n13842) );
  NAND U14005 ( .A(n13666), .B(n13665), .Z(n13670) );
  NANDN U14006 ( .A(n13668), .B(n13667), .Z(n13669) );
  NAND U14007 ( .A(n13670), .B(n13669), .Z(n13841) );
  XNOR U14008 ( .A(n13842), .B(n13841), .Z(n13843) );
  XNOR U14009 ( .A(n13844), .B(n13843), .Z(n13862) );
  NAND U14010 ( .A(n13672), .B(n13671), .Z(n13676) );
  NAND U14011 ( .A(n13674), .B(n13673), .Z(n13675) );
  AND U14012 ( .A(n13676), .B(n13675), .Z(n13860) );
  NANDN U14013 ( .A(n13678), .B(n13677), .Z(n13682) );
  NANDN U14014 ( .A(n13680), .B(n13679), .Z(n13681) );
  AND U14015 ( .A(n13682), .B(n13681), .Z(n13798) );
  XNOR U14016 ( .A(n13798), .B(n13797), .Z(n13800) );
  AND U14017 ( .A(y[784]), .B(x[135]), .Z(n13687) );
  XOR U14018 ( .A(n13926), .B(n13687), .Z(n13771) );
  XOR U14019 ( .A(n13772), .B(n13771), .Z(n13802) );
  AND U14020 ( .A(x[138]), .B(y[781]), .Z(n13801) );
  XOR U14021 ( .A(n13802), .B(n13801), .Z(n13804) );
  AND U14022 ( .A(x[134]), .B(y[785]), .Z(n13765) );
  AND U14023 ( .A(x[143]), .B(y[776]), .Z(n13764) );
  XOR U14024 ( .A(n13765), .B(n13764), .Z(n13767) );
  AND U14025 ( .A(x[139]), .B(y[780]), .Z(n13766) );
  XOR U14026 ( .A(n13767), .B(n13766), .Z(n13803) );
  XOR U14027 ( .A(n13804), .B(n13803), .Z(n13799) );
  XOR U14028 ( .A(n13800), .B(n13799), .Z(n13859) );
  XNOR U14029 ( .A(n13860), .B(n13859), .Z(n13861) );
  XOR U14030 ( .A(n13862), .B(n13861), .Z(n13848) );
  NAND U14031 ( .A(x[146]), .B(y[778]), .Z(n14532) );
  NANDN U14032 ( .A(n14532), .B(n13692), .Z(n13696) );
  NANDN U14033 ( .A(n13694), .B(n13693), .Z(n13695) );
  AND U14034 ( .A(n13696), .B(n13695), .Z(n13830) );
  NANDN U14035 ( .A(n13698), .B(n13697), .Z(n13702) );
  NAND U14036 ( .A(n13700), .B(n13699), .Z(n13701) );
  NAND U14037 ( .A(n13702), .B(n13701), .Z(n13829) );
  XNOR U14038 ( .A(n13830), .B(n13829), .Z(n13832) );
  NAND U14039 ( .A(n13770), .B(n13772), .Z(n13706) );
  NANDN U14040 ( .A(n13704), .B(n13703), .Z(n13705) );
  AND U14041 ( .A(n13706), .B(n13705), .Z(n13826) );
  AND U14042 ( .A(x[128]), .B(y[791]), .Z(n13778) );
  AND U14043 ( .A(x[151]), .B(y[768]), .Z(n13777) );
  XOR U14044 ( .A(n13778), .B(n13777), .Z(n13780) );
  AND U14045 ( .A(x[150]), .B(y[769]), .Z(n13763) );
  XOR U14046 ( .A(n13763), .B(o[151]), .Z(n13779) );
  XOR U14047 ( .A(n13780), .B(n13779), .Z(n13824) );
  AND U14048 ( .A(y[771]), .B(x[148]), .Z(n14381) );
  NAND U14049 ( .A(y[775]), .B(x[144]), .Z(n13707) );
  XNOR U14050 ( .A(n14381), .B(n13707), .Z(n13762) );
  AND U14051 ( .A(x[147]), .B(y[772]), .Z(n13761) );
  XOR U14052 ( .A(n13762), .B(n13761), .Z(n13823) );
  XOR U14053 ( .A(n13824), .B(n13823), .Z(n13825) );
  XNOR U14054 ( .A(n13826), .B(n13825), .Z(n13831) );
  XOR U14055 ( .A(n13832), .B(n13831), .Z(n13791) );
  XNOR U14056 ( .A(n13792), .B(n13791), .Z(n13794) );
  NAND U14057 ( .A(x[148]), .B(y[777]), .Z(n14699) );
  NANDN U14058 ( .A(n14699), .B(n13708), .Z(n13712) );
  NANDN U14059 ( .A(n13710), .B(n13709), .Z(n13711) );
  AND U14060 ( .A(n13712), .B(n13711), .Z(n13786) );
  NANDN U14061 ( .A(n13714), .B(n13713), .Z(n13718) );
  NANDN U14062 ( .A(n13716), .B(n13715), .Z(n13717) );
  AND U14063 ( .A(n13718), .B(n13717), .Z(n13838) );
  AND U14064 ( .A(x[141]), .B(y[778]), .Z(n13814) );
  AND U14065 ( .A(x[130]), .B(y[789]), .Z(n13813) );
  XOR U14066 ( .A(n13814), .B(n13813), .Z(n13816) );
  AND U14067 ( .A(x[149]), .B(y[770]), .Z(n13815) );
  XOR U14068 ( .A(n13816), .B(n13815), .Z(n13836) );
  AND U14069 ( .A(x[140]), .B(y[779]), .Z(n13774) );
  AND U14070 ( .A(x[129]), .B(y[790]), .Z(n13773) );
  XOR U14071 ( .A(n13774), .B(n13773), .Z(n13775) );
  XOR U14072 ( .A(n13776), .B(n13775), .Z(n13835) );
  XOR U14073 ( .A(n13836), .B(n13835), .Z(n13837) );
  XNOR U14074 ( .A(n13838), .B(n13837), .Z(n13785) );
  XNOR U14075 ( .A(n13786), .B(n13785), .Z(n13788) );
  AND U14076 ( .A(x[143]), .B(y[784]), .Z(n14907) );
  NAND U14077 ( .A(n13720), .B(n14907), .Z(n13724) );
  NANDN U14078 ( .A(n13722), .B(n13721), .Z(n13723) );
  AND U14079 ( .A(n13724), .B(n13723), .Z(n13820) );
  AND U14080 ( .A(x[142]), .B(y[777]), .Z(n13810) );
  AND U14081 ( .A(x[131]), .B(y[788]), .Z(n13809) );
  XOR U14082 ( .A(n13810), .B(n13809), .Z(n13812) );
  AND U14083 ( .A(x[132]), .B(y[787]), .Z(n13811) );
  XOR U14084 ( .A(n13812), .B(n13811), .Z(n13818) );
  AND U14085 ( .A(x[133]), .B(y[786]), .Z(n13806) );
  AND U14086 ( .A(x[146]), .B(y[773]), .Z(n13805) );
  XOR U14087 ( .A(n13806), .B(n13805), .Z(n13808) );
  AND U14088 ( .A(x[145]), .B(y[774]), .Z(n13807) );
  XOR U14089 ( .A(n13808), .B(n13807), .Z(n13817) );
  XOR U14090 ( .A(n13818), .B(n13817), .Z(n13819) );
  XNOR U14091 ( .A(n13820), .B(n13819), .Z(n13787) );
  XOR U14092 ( .A(n13788), .B(n13787), .Z(n13793) );
  XOR U14093 ( .A(n13794), .B(n13793), .Z(n13847) );
  XOR U14094 ( .A(n13848), .B(n13847), .Z(n13849) );
  XOR U14095 ( .A(n13850), .B(n13849), .Z(n13757) );
  NANDN U14096 ( .A(n13730), .B(n13729), .Z(n13734) );
  NAND U14097 ( .A(n13732), .B(n13731), .Z(n13733) );
  AND U14098 ( .A(n13734), .B(n13733), .Z(n13854) );
  NAND U14099 ( .A(n13736), .B(n13735), .Z(n13740) );
  NANDN U14100 ( .A(n13738), .B(n13737), .Z(n13739) );
  AND U14101 ( .A(n13740), .B(n13739), .Z(n13853) );
  XNOR U14102 ( .A(n13854), .B(n13853), .Z(n13855) );
  XOR U14103 ( .A(n13856), .B(n13855), .Z(n13755) );
  XOR U14104 ( .A(n13755), .B(n13756), .Z(n13758) );
  XOR U14105 ( .A(n13757), .B(n13758), .Z(n13869) );
  XOR U14106 ( .A(n13868), .B(n13869), .Z(n13870) );
  XNOR U14107 ( .A(n13871), .B(n13870), .Z(n13867) );
  NAND U14108 ( .A(n13749), .B(n13748), .Z(n13753) );
  NANDN U14109 ( .A(n13751), .B(n13750), .Z(n13752) );
  AND U14110 ( .A(n13753), .B(n13752), .Z(n13865) );
  XOR U14111 ( .A(n13866), .B(n13865), .Z(n13754) );
  XNOR U14112 ( .A(n13867), .B(n13754), .Z(N312) );
  NAND U14113 ( .A(n13756), .B(n13755), .Z(n13760) );
  NAND U14114 ( .A(n13758), .B(n13757), .Z(n13759) );
  AND U14115 ( .A(n13760), .B(n13759), .Z(n13994) );
  AND U14116 ( .A(x[148]), .B(y[775]), .Z(n14165) );
  AND U14117 ( .A(x[144]), .B(y[771]), .Z(n13899) );
  AND U14118 ( .A(x[150]), .B(y[770]), .Z(n13934) );
  XOR U14119 ( .A(n13935), .B(n13934), .Z(n13937) );
  AND U14120 ( .A(x[130]), .B(y[790]), .Z(n13936) );
  XOR U14121 ( .A(n13937), .B(n13936), .Z(n13914) );
  AND U14122 ( .A(n13763), .B(o[151]), .Z(n13939) );
  AND U14123 ( .A(x[129]), .B(y[791]), .Z(n13940) );
  XOR U14124 ( .A(n13941), .B(n13940), .Z(n13938) );
  XOR U14125 ( .A(n13939), .B(n13938), .Z(n13913) );
  XOR U14126 ( .A(n13914), .B(n13913), .Z(n13916) );
  XNOR U14127 ( .A(n13917), .B(n13916), .Z(n13966) );
  AND U14128 ( .A(y[771]), .B(x[149]), .Z(n13769) );
  NAND U14129 ( .A(y[776]), .B(x[144]), .Z(n13768) );
  XNOR U14130 ( .A(n13769), .B(n13768), .Z(n13901) );
  AND U14131 ( .A(x[133]), .B(y[787]), .Z(n13900) );
  XOR U14132 ( .A(n13901), .B(n13900), .Z(n13910) );
  AND U14133 ( .A(x[134]), .B(y[786]), .Z(n14178) );
  AND U14134 ( .A(x[148]), .B(y[772]), .Z(n13904) );
  XOR U14135 ( .A(n14178), .B(n13904), .Z(n13906) );
  AND U14136 ( .A(x[147]), .B(y[773]), .Z(n13905) );
  XOR U14137 ( .A(n13906), .B(n13905), .Z(n13909) );
  XOR U14138 ( .A(n13910), .B(n13909), .Z(n13912) );
  XOR U14139 ( .A(n13911), .B(n13912), .Z(n13891) );
  XOR U14140 ( .A(n13890), .B(n13889), .Z(n13892) );
  XOR U14141 ( .A(n13891), .B(n13892), .Z(n13967) );
  XNOR U14142 ( .A(n13966), .B(n13967), .Z(n13969) );
  AND U14143 ( .A(x[131]), .B(y[789]), .Z(n13948) );
  XOR U14144 ( .A(n13949), .B(n13948), .Z(n13950) );
  NAND U14145 ( .A(x[132]), .B(y[788]), .Z(n13951) );
  XNOR U14146 ( .A(n13950), .B(n13951), .Z(n13960) );
  XNOR U14147 ( .A(n13961), .B(n13960), .Z(n13962) );
  AND U14148 ( .A(y[783]), .B(x[137]), .Z(n13782) );
  NAND U14149 ( .A(y[782]), .B(x[138]), .Z(n13781) );
  XNOR U14150 ( .A(n13782), .B(n13781), .Z(n13928) );
  AND U14151 ( .A(y[778]), .B(x[142]), .Z(n13784) );
  NAND U14152 ( .A(y[784]), .B(x[136]), .Z(n13783) );
  XNOR U14153 ( .A(n13784), .B(n13783), .Z(n13930) );
  AND U14154 ( .A(x[139]), .B(y[781]), .Z(n13931) );
  XOR U14155 ( .A(n13930), .B(n13931), .Z(n13927) );
  XOR U14156 ( .A(n13928), .B(n13927), .Z(n13963) );
  XOR U14157 ( .A(n13962), .B(n13963), .Z(n13968) );
  XOR U14158 ( .A(n13969), .B(n13968), .Z(n13977) );
  NANDN U14159 ( .A(n13786), .B(n13785), .Z(n13790) );
  NAND U14160 ( .A(n13788), .B(n13787), .Z(n13789) );
  AND U14161 ( .A(n13790), .B(n13789), .Z(n13976) );
  XNOR U14162 ( .A(n13977), .B(n13976), .Z(n13978) );
  NANDN U14163 ( .A(n13792), .B(n13791), .Z(n13796) );
  NAND U14164 ( .A(n13794), .B(n13793), .Z(n13795) );
  NAND U14165 ( .A(n13796), .B(n13795), .Z(n13979) );
  XNOR U14166 ( .A(n13978), .B(n13979), .Z(n13985) );
  AND U14167 ( .A(x[128]), .B(y[792]), .Z(n13955) );
  AND U14168 ( .A(x[152]), .B(y[768]), .Z(n13954) );
  XOR U14169 ( .A(n13955), .B(n13954), .Z(n13957) );
  AND U14170 ( .A(x[151]), .B(y[769]), .Z(n13947) );
  XOR U14171 ( .A(n13947), .B(o[152]), .Z(n13956) );
  XOR U14172 ( .A(n13957), .B(n13956), .Z(n13896) );
  AND U14173 ( .A(x[135]), .B(y[785]), .Z(n13943) );
  AND U14174 ( .A(x[146]), .B(y[774]), .Z(n13942) );
  XOR U14175 ( .A(n13943), .B(n13942), .Z(n13945) );
  AND U14176 ( .A(x[145]), .B(y[775]), .Z(n13944) );
  XOR U14177 ( .A(n13945), .B(n13944), .Z(n13895) );
  XOR U14178 ( .A(n13896), .B(n13895), .Z(n13898) );
  XOR U14179 ( .A(n13897), .B(n13898), .Z(n13888) );
  XOR U14180 ( .A(n13885), .B(n13886), .Z(n13887) );
  XOR U14181 ( .A(n13888), .B(n13887), .Z(n13972) );
  XNOR U14182 ( .A(n13973), .B(n13972), .Z(n13975) );
  XOR U14183 ( .A(n13974), .B(n13975), .Z(n13881) );
  NAND U14184 ( .A(n13818), .B(n13817), .Z(n13822) );
  NANDN U14185 ( .A(n13820), .B(n13819), .Z(n13821) );
  AND U14186 ( .A(n13822), .B(n13821), .Z(n13921) );
  NAND U14187 ( .A(n13824), .B(n13823), .Z(n13828) );
  NANDN U14188 ( .A(n13826), .B(n13825), .Z(n13827) );
  AND U14189 ( .A(n13828), .B(n13827), .Z(n13920) );
  XOR U14190 ( .A(n13921), .B(n13920), .Z(n13923) );
  NANDN U14191 ( .A(n13830), .B(n13829), .Z(n13834) );
  NAND U14192 ( .A(n13832), .B(n13831), .Z(n13833) );
  AND U14193 ( .A(n13834), .B(n13833), .Z(n13922) );
  XOR U14194 ( .A(n13923), .B(n13922), .Z(n13879) );
  NAND U14195 ( .A(n13836), .B(n13835), .Z(n13840) );
  NANDN U14196 ( .A(n13838), .B(n13837), .Z(n13839) );
  NAND U14197 ( .A(n13840), .B(n13839), .Z(n13880) );
  XNOR U14198 ( .A(n13879), .B(n13880), .Z(n13882) );
  XOR U14199 ( .A(n13881), .B(n13882), .Z(n13982) );
  NANDN U14200 ( .A(n13842), .B(n13841), .Z(n13846) );
  NANDN U14201 ( .A(n13844), .B(n13843), .Z(n13845) );
  NAND U14202 ( .A(n13846), .B(n13845), .Z(n13983) );
  XNOR U14203 ( .A(n13982), .B(n13983), .Z(n13984) );
  XOR U14204 ( .A(n13985), .B(n13984), .Z(n13992) );
  NAND U14205 ( .A(n13848), .B(n13847), .Z(n13852) );
  NANDN U14206 ( .A(n13850), .B(n13849), .Z(n13851) );
  AND U14207 ( .A(n13852), .B(n13851), .Z(n13876) );
  NANDN U14208 ( .A(n13854), .B(n13853), .Z(n13858) );
  NANDN U14209 ( .A(n13856), .B(n13855), .Z(n13857) );
  AND U14210 ( .A(n13858), .B(n13857), .Z(n13874) );
  NANDN U14211 ( .A(n13860), .B(n13859), .Z(n13864) );
  NAND U14212 ( .A(n13862), .B(n13861), .Z(n13863) );
  NAND U14213 ( .A(n13864), .B(n13863), .Z(n13873) );
  XNOR U14214 ( .A(n13874), .B(n13873), .Z(n13875) );
  XNOR U14215 ( .A(n13876), .B(n13875), .Z(n13991) );
  XNOR U14216 ( .A(n13992), .B(n13991), .Z(n13993) );
  XNOR U14217 ( .A(n13994), .B(n13993), .Z(n13990) );
  XOR U14218 ( .A(n13988), .B(n13989), .Z(n13872) );
  XNOR U14219 ( .A(n13990), .B(n13872), .Z(N313) );
  NANDN U14220 ( .A(n13874), .B(n13873), .Z(n13878) );
  NANDN U14221 ( .A(n13876), .B(n13875), .Z(n13877) );
  AND U14222 ( .A(n13878), .B(n13877), .Z(n14136) );
  NANDN U14223 ( .A(n13880), .B(n13879), .Z(n13884) );
  NAND U14224 ( .A(n13882), .B(n13881), .Z(n13883) );
  NAND U14225 ( .A(n13884), .B(n13883), .Z(n14006) );
  NANDN U14226 ( .A(n13890), .B(n13889), .Z(n13894) );
  NANDN U14227 ( .A(n13892), .B(n13891), .Z(n13893) );
  NAND U14228 ( .A(n13894), .B(n13893), .Z(n14011) );
  XOR U14229 ( .A(n14010), .B(n14011), .Z(n14013) );
  NAND U14230 ( .A(x[149]), .B(y[776]), .Z(n14878) );
  AND U14231 ( .A(x[150]), .B(y[771]), .Z(n14079) );
  AND U14232 ( .A(x[133]), .B(y[788]), .Z(n14077) );
  NAND U14233 ( .A(x[145]), .B(y[776]), .Z(n14076) );
  XNOR U14234 ( .A(n14077), .B(n14076), .Z(n14078) );
  XOR U14235 ( .A(n14079), .B(n14078), .Z(n14104) );
  AND U14236 ( .A(y[773]), .B(x[148]), .Z(n13903) );
  NAND U14237 ( .A(y[772]), .B(x[149]), .Z(n13902) );
  XNOR U14238 ( .A(n13903), .B(n13902), .Z(n14091) );
  AND U14239 ( .A(x[147]), .B(y[774]), .Z(n14090) );
  XOR U14240 ( .A(n14091), .B(n14090), .Z(n14105) );
  XOR U14241 ( .A(n14104), .B(n14105), .Z(n14107) );
  XOR U14242 ( .A(n14106), .B(n14107), .Z(n14039) );
  IV U14243 ( .A(n13904), .Z(n14089) );
  NANDN U14244 ( .A(n14089), .B(n14178), .Z(n13908) );
  NAND U14245 ( .A(n13906), .B(n13905), .Z(n13907) );
  NAND U14246 ( .A(n13908), .B(n13907), .Z(n14112) );
  AND U14247 ( .A(x[143]), .B(y[778]), .Z(n14097) );
  AND U14248 ( .A(x[146]), .B(y[775]), .Z(n14095) );
  NAND U14249 ( .A(x[134]), .B(y[787]), .Z(n14094) );
  XNOR U14250 ( .A(n14095), .B(n14094), .Z(n14096) );
  XOR U14251 ( .A(n14097), .B(n14096), .Z(n14111) );
  AND U14252 ( .A(x[151]), .B(y[770]), .Z(n14072) );
  AND U14253 ( .A(x[132]), .B(y[789]), .Z(n14071) );
  NAND U14254 ( .A(x[144]), .B(y[777]), .Z(n14070) );
  XOR U14255 ( .A(n14071), .B(n14070), .Z(n14073) );
  XNOR U14256 ( .A(n14072), .B(n14073), .Z(n14110) );
  XOR U14257 ( .A(n14111), .B(n14110), .Z(n14113) );
  XOR U14258 ( .A(n14112), .B(n14113), .Z(n14038) );
  XOR U14259 ( .A(n14039), .B(n14038), .Z(n14040) );
  XOR U14260 ( .A(n14041), .B(n14040), .Z(n14048) );
  IV U14261 ( .A(n13913), .Z(n13915) );
  NANDN U14262 ( .A(n13915), .B(n13914), .Z(n13919) );
  NANDN U14263 ( .A(n13917), .B(n13916), .Z(n13918) );
  NAND U14264 ( .A(n13919), .B(n13918), .Z(n14047) );
  XNOR U14265 ( .A(n14046), .B(n14047), .Z(n14049) );
  XOR U14266 ( .A(n14048), .B(n14049), .Z(n14012) );
  XOR U14267 ( .A(n14013), .B(n14012), .Z(n14005) );
  NAND U14268 ( .A(n13921), .B(n13920), .Z(n13925) );
  NAND U14269 ( .A(n13923), .B(n13922), .Z(n13924) );
  NAND U14270 ( .A(n13925), .B(n13924), .Z(n14004) );
  XNOR U14271 ( .A(n14005), .B(n14004), .Z(n14007) );
  XNOR U14272 ( .A(n14006), .B(n14007), .Z(n14000) );
  IV U14273 ( .A(n13946), .Z(n14020) );
  AND U14274 ( .A(x[142]), .B(y[784]), .Z(n14969) );
  NAND U14275 ( .A(n14969), .B(n13929), .Z(n13933) );
  NAND U14276 ( .A(n13931), .B(n13930), .Z(n13932) );
  NAND U14277 ( .A(n13933), .B(n13932), .Z(n14066) );
  AND U14278 ( .A(x[139]), .B(y[782]), .Z(n14086) );
  AND U14279 ( .A(x[140]), .B(y[781]), .Z(n14084) );
  NAND U14280 ( .A(x[135]), .B(y[786]), .Z(n14083) );
  XNOR U14281 ( .A(n14084), .B(n14083), .Z(n14085) );
  XOR U14282 ( .A(n14086), .B(n14085), .Z(n14064) );
  NAND U14283 ( .A(x[152]), .B(y[769]), .Z(n14082) );
  XNOR U14284 ( .A(o[153]), .B(n14082), .Z(n14053) );
  AND U14285 ( .A(x[129]), .B(y[792]), .Z(n14052) );
  XOR U14286 ( .A(n14053), .B(n14052), .Z(n14055) );
  AND U14287 ( .A(x[141]), .B(y[780]), .Z(n14054) );
  XOR U14288 ( .A(n14055), .B(n14054), .Z(n14065) );
  XOR U14289 ( .A(n14064), .B(n14065), .Z(n14067) );
  XOR U14290 ( .A(n14066), .B(n14067), .Z(n14043) );
  XOR U14291 ( .A(n14042), .B(n14043), .Z(n14045) );
  XOR U14292 ( .A(n14033), .B(n14032), .Z(n14035) );
  AND U14293 ( .A(x[136]), .B(y[785]), .Z(n14023) );
  XOR U14294 ( .A(n14021), .B(n13946), .Z(n14022) );
  XOR U14295 ( .A(n14023), .B(n14022), .Z(n14027) );
  AND U14296 ( .A(n13947), .B(o[152]), .Z(n14016) );
  AND U14297 ( .A(x[153]), .B(y[768]), .Z(n14015) );
  NAND U14298 ( .A(x[128]), .B(y[793]), .Z(n14014) );
  XOR U14299 ( .A(n14015), .B(n14014), .Z(n14017) );
  XNOR U14300 ( .A(n14016), .B(n14017), .Z(n14026) );
  XOR U14301 ( .A(n14027), .B(n14026), .Z(n14029) );
  XOR U14302 ( .A(n14028), .B(n14029), .Z(n14034) );
  XOR U14303 ( .A(n14035), .B(n14034), .Z(n14044) );
  XOR U14304 ( .A(n14045), .B(n14044), .Z(n14123) );
  AND U14305 ( .A(n13949), .B(n13948), .Z(n13953) );
  NANDN U14306 ( .A(n13951), .B(n13950), .Z(n13952) );
  NANDN U14307 ( .A(n13953), .B(n13952), .Z(n14102) );
  NAND U14308 ( .A(n13955), .B(n13954), .Z(n13959) );
  NAND U14309 ( .A(n13957), .B(n13956), .Z(n13958) );
  NAND U14310 ( .A(n13959), .B(n13958), .Z(n14100) );
  AND U14311 ( .A(x[142]), .B(y[779]), .Z(n14059) );
  AND U14312 ( .A(x[130]), .B(y[791]), .Z(n14058) );
  XOR U14313 ( .A(n14059), .B(n14058), .Z(n14061) );
  AND U14314 ( .A(x[131]), .B(y[790]), .Z(n14060) );
  XOR U14315 ( .A(n14061), .B(n14060), .Z(n14101) );
  XOR U14316 ( .A(n14100), .B(n14101), .Z(n14103) );
  XOR U14317 ( .A(n14102), .B(n14103), .Z(n14121) );
  NANDN U14318 ( .A(n13961), .B(n13960), .Z(n13965) );
  NAND U14319 ( .A(n13963), .B(n13962), .Z(n13964) );
  AND U14320 ( .A(n13965), .B(n13964), .Z(n14120) );
  NANDN U14321 ( .A(n13967), .B(n13966), .Z(n13971) );
  NAND U14322 ( .A(n13969), .B(n13968), .Z(n13970) );
  AND U14323 ( .A(n13971), .B(n13970), .Z(n14116) );
  XOR U14324 ( .A(n14117), .B(n14116), .Z(n14119) );
  XOR U14325 ( .A(n14119), .B(n14118), .Z(n13999) );
  NANDN U14326 ( .A(n13977), .B(n13976), .Z(n13981) );
  NANDN U14327 ( .A(n13979), .B(n13978), .Z(n13980) );
  AND U14328 ( .A(n13981), .B(n13980), .Z(n13998) );
  XOR U14329 ( .A(n13999), .B(n13998), .Z(n14001) );
  XOR U14330 ( .A(n14000), .B(n14001), .Z(n14134) );
  NANDN U14331 ( .A(n13983), .B(n13982), .Z(n13987) );
  NAND U14332 ( .A(n13985), .B(n13984), .Z(n13986) );
  NAND U14333 ( .A(n13987), .B(n13986), .Z(n14133) );
  XOR U14334 ( .A(n14134), .B(n14133), .Z(n14135) );
  XNOR U14335 ( .A(n14136), .B(n14135), .Z(n14129) );
  NANDN U14336 ( .A(n13992), .B(n13991), .Z(n13996) );
  NAND U14337 ( .A(n13994), .B(n13993), .Z(n13995) );
  AND U14338 ( .A(n13996), .B(n13995), .Z(n14128) );
  IV U14339 ( .A(n14128), .Z(n14126) );
  XOR U14340 ( .A(n14127), .B(n14126), .Z(n13997) );
  XNOR U14341 ( .A(n14129), .B(n13997), .Z(N314) );
  NANDN U14342 ( .A(n13999), .B(n13998), .Z(n14003) );
  NANDN U14343 ( .A(n14001), .B(n14000), .Z(n14002) );
  NAND U14344 ( .A(n14003), .B(n14002), .Z(n14276) );
  NANDN U14345 ( .A(n14005), .B(n14004), .Z(n14009) );
  NAND U14346 ( .A(n14007), .B(n14006), .Z(n14008) );
  AND U14347 ( .A(n14009), .B(n14008), .Z(n14277) );
  XOR U14348 ( .A(n14276), .B(n14277), .Z(n14279) );
  AND U14349 ( .A(x[130]), .B(y[792]), .Z(n14202) );
  XOR U14350 ( .A(n14203), .B(n14202), .Z(n14205) );
  NAND U14351 ( .A(x[152]), .B(y[770]), .Z(n14204) );
  XNOR U14352 ( .A(n14205), .B(n14204), .Z(n14238) );
  NANDN U14353 ( .A(n14015), .B(n14014), .Z(n14019) );
  OR U14354 ( .A(n14017), .B(n14016), .Z(n14018) );
  NAND U14355 ( .A(n14019), .B(n14018), .Z(n14239) );
  XNOR U14356 ( .A(n14238), .B(n14239), .Z(n14240) );
  NANDN U14357 ( .A(n14021), .B(n14020), .Z(n14025) );
  NANDN U14358 ( .A(n14023), .B(n14022), .Z(n14024) );
  NAND U14359 ( .A(n14025), .B(n14024), .Z(n14241) );
  XOR U14360 ( .A(n14240), .B(n14241), .Z(n14148) );
  NAND U14361 ( .A(n14027), .B(n14026), .Z(n14031) );
  NAND U14362 ( .A(n14029), .B(n14028), .Z(n14030) );
  AND U14363 ( .A(n14031), .B(n14030), .Z(n14149) );
  XOR U14364 ( .A(n14148), .B(n14149), .Z(n14151) );
  NAND U14365 ( .A(n14033), .B(n14032), .Z(n14037) );
  NAND U14366 ( .A(n14035), .B(n14034), .Z(n14036) );
  AND U14367 ( .A(n14037), .B(n14036), .Z(n14150) );
  XOR U14368 ( .A(n14151), .B(n14150), .Z(n14146) );
  XNOR U14369 ( .A(n14145), .B(n14144), .Z(n14147) );
  XOR U14370 ( .A(n14146), .B(n14147), .Z(n14269) );
  AND U14371 ( .A(x[140]), .B(y[782]), .Z(n14346) );
  AND U14372 ( .A(x[133]), .B(y[789]), .Z(n14252) );
  XOR U14373 ( .A(n14346), .B(n14252), .Z(n14254) );
  NAND U14374 ( .A(x[138]), .B(y[784]), .Z(n14253) );
  XNOR U14375 ( .A(n14254), .B(n14253), .Z(n14157) );
  AND U14376 ( .A(x[135]), .B(y[787]), .Z(n14155) );
  AND U14377 ( .A(y[788]), .B(x[134]), .Z(n14051) );
  NAND U14378 ( .A(y[786]), .B(x[136]), .Z(n14050) );
  XNOR U14379 ( .A(n14051), .B(n14050), .Z(n14179) );
  NAND U14380 ( .A(x[137]), .B(y[785]), .Z(n14180) );
  XNOR U14381 ( .A(n14179), .B(n14180), .Z(n14154) );
  XOR U14382 ( .A(n14155), .B(n14154), .Z(n14156) );
  XOR U14383 ( .A(n14157), .B(n14156), .Z(n14228) );
  NAND U14384 ( .A(n14053), .B(n14052), .Z(n14057) );
  NAND U14385 ( .A(n14055), .B(n14054), .Z(n14056) );
  NAND U14386 ( .A(n14057), .B(n14056), .Z(n14227) );
  NAND U14387 ( .A(n14059), .B(n14058), .Z(n14063) );
  NAND U14388 ( .A(n14061), .B(n14060), .Z(n14062) );
  NAND U14389 ( .A(n14063), .B(n14062), .Z(n14226) );
  XNOR U14390 ( .A(n14227), .B(n14226), .Z(n14229) );
  NAND U14391 ( .A(n14065), .B(n14064), .Z(n14069) );
  NAND U14392 ( .A(n14067), .B(n14066), .Z(n14068) );
  AND U14393 ( .A(n14069), .B(n14068), .Z(n14263) );
  NANDN U14394 ( .A(n14071), .B(n14070), .Z(n14075) );
  OR U14395 ( .A(n14073), .B(n14072), .Z(n14074) );
  AND U14396 ( .A(n14075), .B(n14074), .Z(n14192) );
  NANDN U14397 ( .A(n14077), .B(n14076), .Z(n14081) );
  NANDN U14398 ( .A(n14079), .B(n14078), .Z(n14080) );
  NAND U14399 ( .A(n14081), .B(n14080), .Z(n14193) );
  XNOR U14400 ( .A(n14192), .B(n14193), .Z(n14194) );
  ANDN U14401 ( .B(o[153]), .A(n14082), .Z(n14172) );
  NAND U14402 ( .A(x[142]), .B(y[780]), .Z(n14173) );
  XNOR U14403 ( .A(n14172), .B(n14173), .Z(n14174) );
  NAND U14404 ( .A(x[129]), .B(y[793]), .Z(n14175) );
  XNOR U14405 ( .A(n14174), .B(n14175), .Z(n14244) );
  NAND U14406 ( .A(x[153]), .B(y[769]), .Z(n14183) );
  XNOR U14407 ( .A(o[154]), .B(n14183), .Z(n14257) );
  NAND U14408 ( .A(x[154]), .B(y[768]), .Z(n14258) );
  XNOR U14409 ( .A(n14257), .B(n14258), .Z(n14259) );
  NAND U14410 ( .A(x[128]), .B(y[794]), .Z(n14260) );
  XOR U14411 ( .A(n14259), .B(n14260), .Z(n14245) );
  XNOR U14412 ( .A(n14244), .B(n14245), .Z(n14246) );
  NANDN U14413 ( .A(n14084), .B(n14083), .Z(n14088) );
  NANDN U14414 ( .A(n14086), .B(n14085), .Z(n14087) );
  NAND U14415 ( .A(n14088), .B(n14087), .Z(n14247) );
  XOR U14416 ( .A(n14246), .B(n14247), .Z(n14195) );
  XOR U14417 ( .A(n14194), .B(n14195), .Z(n14234) );
  AND U14418 ( .A(x[149]), .B(y[773]), .Z(n14166) );
  NANDN U14419 ( .A(n14089), .B(n14166), .Z(n14093) );
  NAND U14420 ( .A(n14091), .B(n14090), .Z(n14092) );
  NAND U14421 ( .A(n14093), .B(n14092), .Z(n14222) );
  XOR U14422 ( .A(n14167), .B(n14166), .Z(n14169) );
  NAND U14423 ( .A(x[148]), .B(y[774]), .Z(n14168) );
  XNOR U14424 ( .A(n14169), .B(n14168), .Z(n14221) );
  NAND U14425 ( .A(x[151]), .B(y[771]), .Z(n14209) );
  XNOR U14426 ( .A(n14208), .B(n14209), .Z(n14211) );
  AND U14427 ( .A(x[150]), .B(y[772]), .Z(n14210) );
  XOR U14428 ( .A(n14211), .B(n14210), .Z(n14220) );
  XOR U14429 ( .A(n14221), .B(n14220), .Z(n14223) );
  XOR U14430 ( .A(n14222), .B(n14223), .Z(n14233) );
  AND U14431 ( .A(x[131]), .B(y[791]), .Z(n14158) );
  NAND U14432 ( .A(x[139]), .B(y[783]), .Z(n14159) );
  XNOR U14433 ( .A(n14158), .B(n14159), .Z(n14160) );
  NAND U14434 ( .A(x[147]), .B(y[775]), .Z(n14161) );
  XNOR U14435 ( .A(n14160), .B(n14161), .Z(n14199) );
  NAND U14436 ( .A(x[132]), .B(y[790]), .Z(n14215) );
  XNOR U14437 ( .A(n14214), .B(n14215), .Z(n14216) );
  XOR U14438 ( .A(n14199), .B(n14198), .Z(n14200) );
  NANDN U14439 ( .A(n14095), .B(n14094), .Z(n14099) );
  NANDN U14440 ( .A(n14097), .B(n14096), .Z(n14098) );
  NAND U14441 ( .A(n14099), .B(n14098), .Z(n14201) );
  XOR U14442 ( .A(n14200), .B(n14201), .Z(n14232) );
  XOR U14443 ( .A(n14234), .B(n14235), .Z(n14266) );
  XNOR U14444 ( .A(n14265), .B(n14266), .Z(n14189) );
  NAND U14445 ( .A(n14105), .B(n14104), .Z(n14109) );
  NAND U14446 ( .A(n14107), .B(n14106), .Z(n14108) );
  NAND U14447 ( .A(n14109), .B(n14108), .Z(n14184) );
  NAND U14448 ( .A(n14111), .B(n14110), .Z(n14115) );
  NAND U14449 ( .A(n14113), .B(n14112), .Z(n14114) );
  NAND U14450 ( .A(n14115), .B(n14114), .Z(n14185) );
  XOR U14451 ( .A(n14184), .B(n14185), .Z(n14187) );
  XOR U14452 ( .A(n14186), .B(n14187), .Z(n14188) );
  XNOR U14453 ( .A(n14189), .B(n14188), .Z(n14191) );
  XOR U14454 ( .A(n14190), .B(n14191), .Z(n14270) );
  XOR U14455 ( .A(n14269), .B(n14270), .Z(n14272) );
  XOR U14456 ( .A(n14271), .B(n14272), .Z(n14143) );
  NANDN U14457 ( .A(n14121), .B(n14120), .Z(n14125) );
  NANDN U14458 ( .A(n14123), .B(n14122), .Z(n14124) );
  AND U14459 ( .A(n14125), .B(n14124), .Z(n14140) );
  XOR U14460 ( .A(n14141), .B(n14140), .Z(n14142) );
  XOR U14461 ( .A(n14143), .B(n14142), .Z(n14278) );
  XNOR U14462 ( .A(n14279), .B(n14278), .Z(n14275) );
  NANDN U14463 ( .A(n14126), .B(n14127), .Z(n14132) );
  NOR U14464 ( .A(n14128), .B(n14127), .Z(n14130) );
  OR U14465 ( .A(n14130), .B(n14129), .Z(n14131) );
  AND U14466 ( .A(n14132), .B(n14131), .Z(n14273) );
  NAND U14467 ( .A(n14134), .B(n14133), .Z(n14138) );
  NAND U14468 ( .A(n14136), .B(n14135), .Z(n14137) );
  AND U14469 ( .A(n14138), .B(n14137), .Z(n14274) );
  XOR U14470 ( .A(n14273), .B(n14274), .Z(n14139) );
  XNOR U14471 ( .A(n14275), .B(n14139), .Z(N315) );
  NAND U14472 ( .A(n14149), .B(n14148), .Z(n14153) );
  NAND U14473 ( .A(n14151), .B(n14150), .Z(n14152) );
  NAND U14474 ( .A(n14153), .B(n14152), .Z(n14304) );
  NANDN U14475 ( .A(n14159), .B(n14158), .Z(n14163) );
  NANDN U14476 ( .A(n14161), .B(n14160), .Z(n14162) );
  AND U14477 ( .A(n14163), .B(n14162), .Z(n14372) );
  NAND U14478 ( .A(y[771]), .B(x[152]), .Z(n14164) );
  XNOR U14479 ( .A(n14165), .B(n14164), .Z(n14382) );
  NAND U14480 ( .A(x[135]), .B(y[788]), .Z(n14383) );
  XNOR U14481 ( .A(n14382), .B(n14383), .Z(n14369) );
  AND U14482 ( .A(x[136]), .B(y[787]), .Z(n14340) );
  NAND U14483 ( .A(x[151]), .B(y[772]), .Z(n14341) );
  XNOR U14484 ( .A(n14340), .B(n14341), .Z(n14342) );
  NAND U14485 ( .A(x[150]), .B(y[773]), .Z(n14343) );
  XOR U14486 ( .A(n14342), .B(n14343), .Z(n14370) );
  XNOR U14487 ( .A(n14369), .B(n14370), .Z(n14371) );
  XOR U14488 ( .A(n14372), .B(n14371), .Z(n14432) );
  NAND U14489 ( .A(n14167), .B(n14166), .Z(n14171) );
  ANDN U14490 ( .B(n14169), .A(n14168), .Z(n14170) );
  ANDN U14491 ( .B(n14171), .A(n14170), .Z(n14364) );
  NANDN U14492 ( .A(n14173), .B(n14172), .Z(n14177) );
  NANDN U14493 ( .A(n14175), .B(n14174), .Z(n14176) );
  NAND U14494 ( .A(n14177), .B(n14176), .Z(n14363) );
  XNOR U14495 ( .A(n14364), .B(n14363), .Z(n14365) );
  AND U14496 ( .A(y[788]), .B(x[136]), .Z(n14412) );
  NAND U14497 ( .A(n14412), .B(n14178), .Z(n14182) );
  NANDN U14498 ( .A(n14180), .B(n14179), .Z(n14181) );
  AND U14499 ( .A(n14182), .B(n14181), .Z(n14325) );
  AND U14500 ( .A(x[142]), .B(y[781]), .Z(n14357) );
  NAND U14501 ( .A(x[129]), .B(y[794]), .Z(n14358) );
  XNOR U14502 ( .A(n14357), .B(n14358), .Z(n14359) );
  ANDN U14503 ( .B(o[154]), .A(n14183), .Z(n14360) );
  XOR U14504 ( .A(n14359), .B(n14360), .Z(n14322) );
  AND U14505 ( .A(x[145]), .B(y[778]), .Z(n14392) );
  NAND U14506 ( .A(x[132]), .B(y[791]), .Z(n14393) );
  XNOR U14507 ( .A(n14392), .B(n14393), .Z(n14394) );
  NAND U14508 ( .A(x[133]), .B(y[790]), .Z(n14395) );
  XOR U14509 ( .A(n14394), .B(n14395), .Z(n14323) );
  XNOR U14510 ( .A(n14322), .B(n14323), .Z(n14324) );
  XOR U14511 ( .A(n14325), .B(n14324), .Z(n14366) );
  XOR U14512 ( .A(n14365), .B(n14366), .Z(n14431) );
  XNOR U14513 ( .A(n14432), .B(n14431), .Z(n14434) );
  XOR U14514 ( .A(n14304), .B(n14305), .Z(n14307) );
  XOR U14515 ( .A(n14307), .B(n14306), .Z(n14299) );
  XOR U14516 ( .A(n14298), .B(n14299), .Z(n14301) );
  NANDN U14517 ( .A(n14193), .B(n14192), .Z(n14197) );
  NANDN U14518 ( .A(n14195), .B(n14194), .Z(n14196) );
  AND U14519 ( .A(n14197), .B(n14196), .Z(n14422) );
  NAND U14520 ( .A(n14203), .B(n14202), .Z(n14207) );
  ANDN U14521 ( .B(n14205), .A(n14204), .Z(n14206) );
  ANDN U14522 ( .B(n14207), .A(n14206), .Z(n14317) );
  NANDN U14523 ( .A(n14209), .B(n14208), .Z(n14213) );
  NAND U14524 ( .A(n14211), .B(n14210), .Z(n14212) );
  NAND U14525 ( .A(n14213), .B(n14212), .Z(n14316) );
  XNOR U14526 ( .A(n14317), .B(n14316), .Z(n14318) );
  NANDN U14527 ( .A(n14215), .B(n14214), .Z(n14219) );
  NANDN U14528 ( .A(n14217), .B(n14216), .Z(n14218) );
  AND U14529 ( .A(n14219), .B(n14218), .Z(n14331) );
  AND U14530 ( .A(x[128]), .B(y[795]), .Z(n14398) );
  NAND U14531 ( .A(x[155]), .B(y[768]), .Z(n14399) );
  XNOR U14532 ( .A(n14398), .B(n14399), .Z(n14400) );
  AND U14533 ( .A(x[154]), .B(y[769]), .Z(n14410) );
  XOR U14534 ( .A(o[155]), .B(n14410), .Z(n14401) );
  XOR U14535 ( .A(n14400), .B(n14401), .Z(n14328) );
  AND U14536 ( .A(x[137]), .B(y[786]), .Z(n14404) );
  NAND U14537 ( .A(x[149]), .B(y[774]), .Z(n14405) );
  XNOR U14538 ( .A(n14404), .B(n14405), .Z(n14406) );
  NAND U14539 ( .A(x[146]), .B(y[777]), .Z(n14407) );
  XOR U14540 ( .A(n14406), .B(n14407), .Z(n14329) );
  XNOR U14541 ( .A(n14328), .B(n14329), .Z(n14330) );
  XOR U14542 ( .A(n14331), .B(n14330), .Z(n14319) );
  XNOR U14543 ( .A(n14318), .B(n14319), .Z(n14419) );
  XNOR U14544 ( .A(n14420), .B(n14419), .Z(n14421) );
  XOR U14545 ( .A(n14422), .B(n14421), .Z(n14439) );
  NAND U14546 ( .A(n14221), .B(n14220), .Z(n14225) );
  NAND U14547 ( .A(n14223), .B(n14222), .Z(n14224) );
  AND U14548 ( .A(n14225), .B(n14224), .Z(n14438) );
  NAND U14549 ( .A(n14227), .B(n14226), .Z(n14231) );
  NANDN U14550 ( .A(n14229), .B(n14228), .Z(n14230) );
  AND U14551 ( .A(n14231), .B(n14230), .Z(n14437) );
  XOR U14552 ( .A(n14438), .B(n14437), .Z(n14440) );
  XOR U14553 ( .A(n14439), .B(n14440), .Z(n14292) );
  NANDN U14554 ( .A(n14233), .B(n14232), .Z(n14237) );
  NANDN U14555 ( .A(n14235), .B(n14234), .Z(n14236) );
  AND U14556 ( .A(n14237), .B(n14236), .Z(n14426) );
  NANDN U14557 ( .A(n14239), .B(n14238), .Z(n14243) );
  NANDN U14558 ( .A(n14241), .B(n14240), .Z(n14242) );
  AND U14559 ( .A(n14243), .B(n14242), .Z(n14415) );
  NANDN U14560 ( .A(n14245), .B(n14244), .Z(n14249) );
  NANDN U14561 ( .A(n14247), .B(n14246), .Z(n14248) );
  AND U14562 ( .A(n14249), .B(n14248), .Z(n14414) );
  AND U14563 ( .A(x[147]), .B(y[776]), .Z(n14386) );
  NAND U14564 ( .A(x[153]), .B(y[770]), .Z(n14387) );
  XNOR U14565 ( .A(n14386), .B(n14387), .Z(n14388) );
  NAND U14566 ( .A(x[134]), .B(y[789]), .Z(n14389) );
  XNOR U14567 ( .A(n14388), .B(n14389), .Z(n14375) );
  AND U14568 ( .A(x[143]), .B(y[780]), .Z(n14351) );
  NAND U14569 ( .A(x[130]), .B(y[793]), .Z(n14352) );
  XNOR U14570 ( .A(n14351), .B(n14352), .Z(n14353) );
  NAND U14571 ( .A(x[131]), .B(y[792]), .Z(n14354) );
  XOR U14572 ( .A(n14353), .B(n14354), .Z(n14376) );
  XNOR U14573 ( .A(n14375), .B(n14376), .Z(n14377) );
  AND U14574 ( .A(x[144]), .B(y[779]), .Z(n14335) );
  XOR U14575 ( .A(n14335), .B(n14334), .Z(n14336) );
  XOR U14576 ( .A(n14337), .B(n14336), .Z(n14348) );
  AND U14577 ( .A(y[782]), .B(x[141]), .Z(n14251) );
  NAND U14578 ( .A(y[783]), .B(x[140]), .Z(n14250) );
  XNOR U14579 ( .A(n14251), .B(n14250), .Z(n14347) );
  XOR U14580 ( .A(n14348), .B(n14347), .Z(n14378) );
  XOR U14581 ( .A(n14377), .B(n14378), .Z(n14312) );
  NAND U14582 ( .A(n14346), .B(n14252), .Z(n14256) );
  ANDN U14583 ( .B(n14254), .A(n14253), .Z(n14255) );
  ANDN U14584 ( .B(n14256), .A(n14255), .Z(n14311) );
  NANDN U14585 ( .A(n14258), .B(n14257), .Z(n14262) );
  NANDN U14586 ( .A(n14260), .B(n14259), .Z(n14261) );
  NAND U14587 ( .A(n14262), .B(n14261), .Z(n14310) );
  XOR U14588 ( .A(n14311), .B(n14310), .Z(n14313) );
  XNOR U14589 ( .A(n14312), .B(n14313), .Z(n14413) );
  XOR U14590 ( .A(n14414), .B(n14413), .Z(n14416) );
  XOR U14591 ( .A(n14415), .B(n14416), .Z(n14425) );
  XOR U14592 ( .A(n14426), .B(n14425), .Z(n14428) );
  NANDN U14593 ( .A(n14264), .B(n14263), .Z(n14268) );
  NANDN U14594 ( .A(n14266), .B(n14265), .Z(n14267) );
  AND U14595 ( .A(n14268), .B(n14267), .Z(n14427) );
  XOR U14596 ( .A(n14428), .B(n14427), .Z(n14293) );
  XOR U14597 ( .A(n14295), .B(n14294), .Z(n14300) );
  XOR U14598 ( .A(n14301), .B(n14300), .Z(n14284) );
  XOR U14599 ( .A(n14284), .B(n14283), .Z(n14286) );
  XOR U14600 ( .A(n14285), .B(n14286), .Z(n14291) );
  NAND U14601 ( .A(n14277), .B(n14276), .Z(n14281) );
  NAND U14602 ( .A(n14279), .B(n14278), .Z(n14280) );
  NAND U14603 ( .A(n14281), .B(n14280), .Z(n14289) );
  XNOR U14604 ( .A(n14290), .B(n14289), .Z(n14282) );
  XNOR U14605 ( .A(n14291), .B(n14282), .Z(N316) );
  NANDN U14606 ( .A(n14284), .B(n14283), .Z(n14288) );
  NANDN U14607 ( .A(n14286), .B(n14285), .Z(n14287) );
  AND U14608 ( .A(n14288), .B(n14287), .Z(n14451) );
  NANDN U14609 ( .A(n14293), .B(n14292), .Z(n14297) );
  NAND U14610 ( .A(n14295), .B(n14294), .Z(n14296) );
  AND U14611 ( .A(n14297), .B(n14296), .Z(n14445) );
  NAND U14612 ( .A(n14299), .B(n14298), .Z(n14303) );
  NAND U14613 ( .A(n14301), .B(n14300), .Z(n14302) );
  AND U14614 ( .A(n14303), .B(n14302), .Z(n14444) );
  XOR U14615 ( .A(n14445), .B(n14444), .Z(n14447) );
  NAND U14616 ( .A(n14305), .B(n14304), .Z(n14309) );
  NAND U14617 ( .A(n14307), .B(n14306), .Z(n14308) );
  AND U14618 ( .A(n14309), .B(n14308), .Z(n14454) );
  NANDN U14619 ( .A(n14311), .B(n14310), .Z(n14315) );
  NANDN U14620 ( .A(n14313), .B(n14312), .Z(n14314) );
  AND U14621 ( .A(n14315), .B(n14314), .Z(n14478) );
  NANDN U14622 ( .A(n14317), .B(n14316), .Z(n14321) );
  NANDN U14623 ( .A(n14319), .B(n14318), .Z(n14320) );
  AND U14624 ( .A(n14321), .B(n14320), .Z(n14583) );
  NANDN U14625 ( .A(n14323), .B(n14322), .Z(n14327) );
  NANDN U14626 ( .A(n14325), .B(n14324), .Z(n14326) );
  AND U14627 ( .A(n14327), .B(n14326), .Z(n14581) );
  NANDN U14628 ( .A(n14329), .B(n14328), .Z(n14333) );
  NANDN U14629 ( .A(n14331), .B(n14330), .Z(n14332) );
  NAND U14630 ( .A(n14333), .B(n14332), .Z(n14580) );
  XNOR U14631 ( .A(n14581), .B(n14580), .Z(n14582) );
  XNOR U14632 ( .A(n14583), .B(n14582), .Z(n14477) );
  XNOR U14633 ( .A(n14478), .B(n14477), .Z(n14480) );
  OR U14634 ( .A(n14335), .B(n14334), .Z(n14339) );
  NANDN U14635 ( .A(n14337), .B(n14336), .Z(n14338) );
  AND U14636 ( .A(n14339), .B(n14338), .Z(n14545) );
  AND U14637 ( .A(x[135]), .B(y[789]), .Z(n14525) );
  AND U14638 ( .A(x[140]), .B(y[784]), .Z(n14524) );
  XOR U14639 ( .A(n14525), .B(n14524), .Z(n14527) );
  AND U14640 ( .A(x[139]), .B(y[785]), .Z(n14526) );
  XOR U14641 ( .A(n14527), .B(n14526), .Z(n14543) );
  AND U14642 ( .A(x[155]), .B(y[769]), .Z(n14541) );
  XOR U14643 ( .A(o[156]), .B(n14541), .Z(n14555) );
  AND U14644 ( .A(x[154]), .B(y[770]), .Z(n14554) );
  XOR U14645 ( .A(n14555), .B(n14554), .Z(n14557) );
  AND U14646 ( .A(x[143]), .B(y[781]), .Z(n14556) );
  XNOR U14647 ( .A(n14557), .B(n14556), .Z(n14542) );
  NANDN U14648 ( .A(n14341), .B(n14340), .Z(n14345) );
  NANDN U14649 ( .A(n14343), .B(n14342), .Z(n14344) );
  AND U14650 ( .A(n14345), .B(n14344), .Z(n14565) );
  AND U14651 ( .A(x[145]), .B(y[779]), .Z(n14490) );
  AND U14652 ( .A(x[150]), .B(y[774]), .Z(n14489) );
  XOR U14653 ( .A(n14490), .B(n14489), .Z(n14492) );
  AND U14654 ( .A(x[132]), .B(y[792]), .Z(n14491) );
  XOR U14655 ( .A(n14492), .B(n14491), .Z(n14563) );
  AND U14656 ( .A(x[134]), .B(y[790]), .Z(n14722) );
  NAND U14657 ( .A(x[147]), .B(y[777]), .Z(n14530) );
  XOR U14658 ( .A(n14563), .B(n14562), .Z(n14564) );
  XOR U14659 ( .A(n14587), .B(n14586), .Z(n14588) );
  NAND U14660 ( .A(n14548), .B(n14346), .Z(n14350) );
  NAND U14661 ( .A(n14348), .B(n14347), .Z(n14349) );
  AND U14662 ( .A(n14350), .B(n14349), .Z(n14509) );
  NANDN U14663 ( .A(n14352), .B(n14351), .Z(n14356) );
  NANDN U14664 ( .A(n14354), .B(n14353), .Z(n14355) );
  AND U14665 ( .A(n14356), .B(n14355), .Z(n14507) );
  NANDN U14666 ( .A(n14358), .B(n14357), .Z(n14362) );
  NAND U14667 ( .A(n14360), .B(n14359), .Z(n14361) );
  NAND U14668 ( .A(n14362), .B(n14361), .Z(n14506) );
  XOR U14669 ( .A(n14588), .B(n14589), .Z(n14479) );
  XOR U14670 ( .A(n14480), .B(n14479), .Z(n14473) );
  NANDN U14671 ( .A(n14364), .B(n14363), .Z(n14368) );
  NANDN U14672 ( .A(n14366), .B(n14365), .Z(n14367) );
  AND U14673 ( .A(n14368), .B(n14367), .Z(n14570) );
  NANDN U14674 ( .A(n14370), .B(n14369), .Z(n14374) );
  NANDN U14675 ( .A(n14372), .B(n14371), .Z(n14373) );
  AND U14676 ( .A(n14374), .B(n14373), .Z(n14569) );
  NANDN U14677 ( .A(n14376), .B(n14375), .Z(n14380) );
  NAND U14678 ( .A(n14378), .B(n14377), .Z(n14379) );
  NAND U14679 ( .A(n14380), .B(n14379), .Z(n14568) );
  XOR U14680 ( .A(n14569), .B(n14568), .Z(n14571) );
  XOR U14681 ( .A(n14570), .B(n14571), .Z(n14472) );
  AND U14682 ( .A(x[152]), .B(y[775]), .Z(n14897) );
  NAND U14683 ( .A(n14897), .B(n14381), .Z(n14385) );
  NANDN U14684 ( .A(n14383), .B(n14382), .Z(n14384) );
  AND U14685 ( .A(n14385), .B(n14384), .Z(n14607) );
  AND U14686 ( .A(x[153]), .B(y[771]), .Z(n14520) );
  XOR U14687 ( .A(n14521), .B(n14520), .Z(n14519) );
  NAND U14688 ( .A(x[129]), .B(y[795]), .Z(n14518) );
  AND U14689 ( .A(x[144]), .B(y[780]), .Z(n14512) );
  NAND U14690 ( .A(x[152]), .B(y[772]), .Z(n14513) );
  NAND U14691 ( .A(x[130]), .B(y[794]), .Z(n14515) );
  XOR U14692 ( .A(n14604), .B(n14605), .Z(n14606) );
  XOR U14693 ( .A(n14607), .B(n14606), .Z(n14577) );
  NANDN U14694 ( .A(n14387), .B(n14386), .Z(n14391) );
  NANDN U14695 ( .A(n14389), .B(n14388), .Z(n14390) );
  AND U14696 ( .A(n14391), .B(n14390), .Z(n14601) );
  NAND U14697 ( .A(x[131]), .B(y[793]), .Z(n14549) );
  NAND U14698 ( .A(x[151]), .B(y[773]), .Z(n14551) );
  AND U14699 ( .A(x[133]), .B(y[791]), .Z(n14535) );
  NAND U14700 ( .A(x[149]), .B(y[775]), .Z(n14536) );
  NAND U14701 ( .A(x[148]), .B(y[776]), .Z(n14538) );
  XOR U14702 ( .A(n14598), .B(n14599), .Z(n14600) );
  XOR U14703 ( .A(n14601), .B(n14600), .Z(n14575) );
  NANDN U14704 ( .A(n14393), .B(n14392), .Z(n14397) );
  NANDN U14705 ( .A(n14395), .B(n14394), .Z(n14396) );
  AND U14706 ( .A(n14397), .B(n14396), .Z(n14593) );
  NANDN U14707 ( .A(n14399), .B(n14398), .Z(n14403) );
  NAND U14708 ( .A(n14401), .B(n14400), .Z(n14402) );
  NAND U14709 ( .A(n14403), .B(n14402), .Z(n14592) );
  XNOR U14710 ( .A(n14593), .B(n14592), .Z(n14595) );
  NANDN U14711 ( .A(n14405), .B(n14404), .Z(n14409) );
  NANDN U14712 ( .A(n14407), .B(n14406), .Z(n14408) );
  NAND U14713 ( .A(n14409), .B(n14408), .Z(n14485) );
  AND U14714 ( .A(n14410), .B(o[155]), .Z(n14498) );
  AND U14715 ( .A(x[128]), .B(y[796]), .Z(n14496) );
  AND U14716 ( .A(x[156]), .B(y[768]), .Z(n14495) );
  XOR U14717 ( .A(n14496), .B(n14495), .Z(n14497) );
  XOR U14718 ( .A(n14498), .B(n14497), .Z(n14484) );
  NAND U14719 ( .A(y[786]), .B(x[138]), .Z(n14411) );
  XNOR U14720 ( .A(n14412), .B(n14411), .Z(n14503) );
  AND U14721 ( .A(x[137]), .B(y[787]), .Z(n14502) );
  XOR U14722 ( .A(n14503), .B(n14502), .Z(n14483) );
  XOR U14723 ( .A(n14484), .B(n14483), .Z(n14486) );
  XOR U14724 ( .A(n14485), .B(n14486), .Z(n14594) );
  XNOR U14725 ( .A(n14595), .B(n14594), .Z(n14574) );
  XOR U14726 ( .A(n14575), .B(n14574), .Z(n14576) );
  XOR U14727 ( .A(n14577), .B(n14576), .Z(n14471) );
  XOR U14728 ( .A(n14472), .B(n14471), .Z(n14474) );
  XOR U14729 ( .A(n14473), .B(n14474), .Z(n14467) );
  NANDN U14730 ( .A(n14414), .B(n14413), .Z(n14418) );
  OR U14731 ( .A(n14416), .B(n14415), .Z(n14417) );
  AND U14732 ( .A(n14418), .B(n14417), .Z(n14466) );
  NANDN U14733 ( .A(n14420), .B(n14419), .Z(n14424) );
  NANDN U14734 ( .A(n14422), .B(n14421), .Z(n14423) );
  NAND U14735 ( .A(n14424), .B(n14423), .Z(n14465) );
  XOR U14736 ( .A(n14466), .B(n14465), .Z(n14468) );
  XOR U14737 ( .A(n14467), .B(n14468), .Z(n14453) );
  XOR U14738 ( .A(n14454), .B(n14453), .Z(n14456) );
  NAND U14739 ( .A(n14426), .B(n14425), .Z(n14430) );
  NAND U14740 ( .A(n14428), .B(n14427), .Z(n14429) );
  NAND U14741 ( .A(n14430), .B(n14429), .Z(n14461) );
  NAND U14742 ( .A(n14432), .B(n14431), .Z(n14436) );
  NANDN U14743 ( .A(n14434), .B(n14433), .Z(n14435) );
  AND U14744 ( .A(n14436), .B(n14435), .Z(n14460) );
  NAND U14745 ( .A(n14438), .B(n14437), .Z(n14442) );
  NAND U14746 ( .A(n14440), .B(n14439), .Z(n14441) );
  AND U14747 ( .A(n14442), .B(n14441), .Z(n14459) );
  XOR U14748 ( .A(n14460), .B(n14459), .Z(n14462) );
  XOR U14749 ( .A(n14461), .B(n14462), .Z(n14455) );
  XOR U14750 ( .A(n14456), .B(n14455), .Z(n14446) );
  XOR U14751 ( .A(n14447), .B(n14446), .Z(n14452) );
  XOR U14752 ( .A(n14450), .B(n14452), .Z(n14443) );
  XOR U14753 ( .A(n14451), .B(n14443), .Z(N317) );
  NAND U14754 ( .A(n14445), .B(n14444), .Z(n14449) );
  NAND U14755 ( .A(n14447), .B(n14446), .Z(n14448) );
  AND U14756 ( .A(n14449), .B(n14448), .Z(n14611) );
  NAND U14757 ( .A(n14454), .B(n14453), .Z(n14458) );
  NAND U14758 ( .A(n14456), .B(n14455), .Z(n14457) );
  NAND U14759 ( .A(n14458), .B(n14457), .Z(n14616) );
  NAND U14760 ( .A(n14460), .B(n14459), .Z(n14464) );
  NAND U14761 ( .A(n14462), .B(n14461), .Z(n14463) );
  NAND U14762 ( .A(n14464), .B(n14463), .Z(n14614) );
  NANDN U14763 ( .A(n14466), .B(n14465), .Z(n14470) );
  OR U14764 ( .A(n14468), .B(n14467), .Z(n14469) );
  AND U14765 ( .A(n14470), .B(n14469), .Z(n14621) );
  NANDN U14766 ( .A(n14472), .B(n14471), .Z(n14476) );
  OR U14767 ( .A(n14474), .B(n14473), .Z(n14475) );
  AND U14768 ( .A(n14476), .B(n14475), .Z(n14620) );
  XNOR U14769 ( .A(n14621), .B(n14620), .Z(n14622) );
  NANDN U14770 ( .A(n14478), .B(n14477), .Z(n14482) );
  NAND U14771 ( .A(n14480), .B(n14479), .Z(n14481) );
  AND U14772 ( .A(n14482), .B(n14481), .Z(n14639) );
  NAND U14773 ( .A(n14484), .B(n14483), .Z(n14488) );
  NAND U14774 ( .A(n14486), .B(n14485), .Z(n14487) );
  AND U14775 ( .A(n14488), .B(n14487), .Z(n14742) );
  NAND U14776 ( .A(n14490), .B(n14489), .Z(n14494) );
  NAND U14777 ( .A(n14492), .B(n14491), .Z(n14493) );
  NAND U14778 ( .A(n14494), .B(n14493), .Z(n14779) );
  NAND U14779 ( .A(n14496), .B(n14495), .Z(n14500) );
  NAND U14780 ( .A(n14498), .B(n14497), .Z(n14499) );
  NAND U14781 ( .A(n14500), .B(n14499), .Z(n14778) );
  XOR U14782 ( .A(n14779), .B(n14778), .Z(n14780) );
  AND U14783 ( .A(y[788]), .B(x[138]), .Z(n14776) );
  NAND U14784 ( .A(n14776), .B(n14501), .Z(n14505) );
  NAND U14785 ( .A(n14503), .B(n14502), .Z(n14504) );
  NAND U14786 ( .A(n14505), .B(n14504), .Z(n14750) );
  AND U14787 ( .A(x[150]), .B(y[775]), .Z(n14694) );
  AND U14788 ( .A(x[140]), .B(y[785]), .Z(n14836) );
  AND U14789 ( .A(x[129]), .B(y[796]), .Z(n14692) );
  XOR U14790 ( .A(n14836), .B(n14692), .Z(n14693) );
  XOR U14791 ( .A(n14694), .B(n14693), .Z(n14749) );
  AND U14792 ( .A(x[143]), .B(y[782]), .Z(n14697) );
  XOR U14793 ( .A(n14749), .B(n14748), .Z(n14751) );
  XNOR U14794 ( .A(n14750), .B(n14751), .Z(n14781) );
  NANDN U14795 ( .A(n14507), .B(n14506), .Z(n14511) );
  NANDN U14796 ( .A(n14509), .B(n14508), .Z(n14510) );
  AND U14797 ( .A(n14511), .B(n14510), .Z(n14744) );
  XOR U14798 ( .A(n14745), .B(n14744), .Z(n14739) );
  NANDN U14799 ( .A(n14513), .B(n14512), .Z(n14517) );
  NANDN U14800 ( .A(n14515), .B(n14514), .Z(n14516) );
  NAND U14801 ( .A(n14517), .B(n14516), .Z(n14755) );
  ANDN U14802 ( .B(n14519), .A(n14518), .Z(n14523) );
  NAND U14803 ( .A(n14521), .B(n14520), .Z(n14522) );
  NANDN U14804 ( .A(n14523), .B(n14522), .Z(n14754) );
  XOR U14805 ( .A(n14755), .B(n14754), .Z(n14756) );
  NAND U14806 ( .A(n14525), .B(n14524), .Z(n14529) );
  NAND U14807 ( .A(n14527), .B(n14526), .Z(n14528) );
  NAND U14808 ( .A(n14529), .B(n14528), .Z(n14658) );
  AND U14809 ( .A(x[139]), .B(y[786]), .Z(n14719) );
  AND U14810 ( .A(x[131]), .B(y[794]), .Z(n14717) );
  AND U14811 ( .A(x[145]), .B(y[780]), .Z(n14716) );
  XOR U14812 ( .A(n14717), .B(n14716), .Z(n14718) );
  XOR U14813 ( .A(n14719), .B(n14718), .Z(n14657) );
  AND U14814 ( .A(x[151]), .B(y[774]), .Z(n14713) );
  AND U14815 ( .A(x[141]), .B(y[784]), .Z(n14711) );
  AND U14816 ( .A(x[152]), .B(y[773]), .Z(n14975) );
  XOR U14817 ( .A(n14711), .B(n14975), .Z(n14712) );
  XOR U14818 ( .A(n14713), .B(n14712), .Z(n14656) );
  XOR U14819 ( .A(n14657), .B(n14656), .Z(n14659) );
  XNOR U14820 ( .A(n14658), .B(n14659), .Z(n14757) );
  NANDN U14821 ( .A(n14530), .B(n14722), .Z(n14534) );
  NANDN U14822 ( .A(n14532), .B(n14531), .Z(n14533) );
  NAND U14823 ( .A(n14534), .B(n14533), .Z(n14763) );
  AND U14824 ( .A(x[153]), .B(y[772]), .Z(n14689) );
  AND U14825 ( .A(x[154]), .B(y[771]), .Z(n14686) );
  XOR U14826 ( .A(n14687), .B(n14686), .Z(n14688) );
  XOR U14827 ( .A(n14689), .B(n14688), .Z(n14761) );
  AND U14828 ( .A(x[156]), .B(y[769]), .Z(n14704) );
  XOR U14829 ( .A(o[157]), .B(n14704), .Z(n14771) );
  AND U14830 ( .A(x[128]), .B(y[797]), .Z(n14769) );
  AND U14831 ( .A(x[157]), .B(y[768]), .Z(n14768) );
  XOR U14832 ( .A(n14769), .B(n14768), .Z(n14770) );
  XNOR U14833 ( .A(n14771), .B(n14770), .Z(n14760) );
  XOR U14834 ( .A(n14763), .B(n14762), .Z(n14644) );
  NANDN U14835 ( .A(n14536), .B(n14535), .Z(n14540) );
  NANDN U14836 ( .A(n14538), .B(n14537), .Z(n14539) );
  NAND U14837 ( .A(n14540), .B(n14539), .Z(n14707) );
  AND U14838 ( .A(x[130]), .B(y[795]), .Z(n14669) );
  XOR U14839 ( .A(n14669), .B(n14668), .Z(n14670) );
  XOR U14840 ( .A(n14671), .B(n14670), .Z(n14706) );
  AND U14841 ( .A(n14541), .B(o[156]), .Z(n14677) );
  AND U14842 ( .A(x[144]), .B(y[781]), .Z(n14675) );
  AND U14843 ( .A(x[155]), .B(y[770]), .Z(n14674) );
  XOR U14844 ( .A(n14675), .B(n14674), .Z(n14676) );
  XOR U14845 ( .A(n14677), .B(n14676), .Z(n14705) );
  XOR U14846 ( .A(n14706), .B(n14705), .Z(n14708) );
  XOR U14847 ( .A(n14707), .B(n14708), .Z(n14645) );
  NANDN U14848 ( .A(n14543), .B(n14542), .Z(n14547) );
  NANDN U14849 ( .A(n14545), .B(n14544), .Z(n14546) );
  AND U14850 ( .A(n14547), .B(n14546), .Z(n14651) );
  NANDN U14851 ( .A(n14549), .B(n14548), .Z(n14553) );
  NANDN U14852 ( .A(n14551), .B(n14550), .Z(n14552) );
  NAND U14853 ( .A(n14553), .B(n14552), .Z(n14681) );
  NAND U14854 ( .A(n14555), .B(n14554), .Z(n14559) );
  NAND U14855 ( .A(n14557), .B(n14556), .Z(n14558) );
  NAND U14856 ( .A(n14559), .B(n14558), .Z(n14680) );
  XOR U14857 ( .A(n14681), .B(n14680), .Z(n14683) );
  AND U14858 ( .A(x[136]), .B(y[789]), .Z(n14724) );
  AND U14859 ( .A(y[791]), .B(x[134]), .Z(n14561) );
  AND U14860 ( .A(y[790]), .B(x[135]), .Z(n14560) );
  XOR U14861 ( .A(n14561), .B(n14560), .Z(n14723) );
  XOR U14862 ( .A(n14724), .B(n14723), .Z(n14766) );
  AND U14863 ( .A(x[133]), .B(y[792]), .Z(n14665) );
  AND U14864 ( .A(x[132]), .B(y[793]), .Z(n14663) );
  AND U14865 ( .A(x[138]), .B(y[787]), .Z(n14662) );
  XOR U14866 ( .A(n14663), .B(n14662), .Z(n14664) );
  XOR U14867 ( .A(n14665), .B(n14664), .Z(n14767) );
  NAND U14868 ( .A(x[137]), .B(y[788]), .Z(n14873) );
  XNOR U14869 ( .A(n14683), .B(n14682), .Z(n14650) );
  XOR U14870 ( .A(n14653), .B(n14652), .Z(n14737) );
  NAND U14871 ( .A(n14563), .B(n14562), .Z(n14567) );
  NANDN U14872 ( .A(n14565), .B(n14564), .Z(n14566) );
  NAND U14873 ( .A(n14567), .B(n14566), .Z(n14736) );
  XNOR U14874 ( .A(n14639), .B(n14638), .Z(n14640) );
  NANDN U14875 ( .A(n14569), .B(n14568), .Z(n14573) );
  OR U14876 ( .A(n14571), .B(n14570), .Z(n14572) );
  AND U14877 ( .A(n14573), .B(n14572), .Z(n14633) );
  NAND U14878 ( .A(n14575), .B(n14574), .Z(n14579) );
  NAND U14879 ( .A(n14577), .B(n14576), .Z(n14578) );
  AND U14880 ( .A(n14579), .B(n14578), .Z(n14632) );
  XNOR U14881 ( .A(n14633), .B(n14632), .Z(n14634) );
  NANDN U14882 ( .A(n14581), .B(n14580), .Z(n14585) );
  NANDN U14883 ( .A(n14583), .B(n14582), .Z(n14584) );
  AND U14884 ( .A(n14585), .B(n14584), .Z(n14629) );
  NAND U14885 ( .A(n14587), .B(n14586), .Z(n14591) );
  NAND U14886 ( .A(n14589), .B(n14588), .Z(n14590) );
  AND U14887 ( .A(n14591), .B(n14590), .Z(n14627) );
  NANDN U14888 ( .A(n14593), .B(n14592), .Z(n14597) );
  NAND U14889 ( .A(n14595), .B(n14594), .Z(n14596) );
  AND U14890 ( .A(n14597), .B(n14596), .Z(n14732) );
  NAND U14891 ( .A(n14599), .B(n14598), .Z(n14603) );
  NANDN U14892 ( .A(n14601), .B(n14600), .Z(n14602) );
  AND U14893 ( .A(n14603), .B(n14602), .Z(n14730) );
  NAND U14894 ( .A(n14605), .B(n14604), .Z(n14609) );
  NANDN U14895 ( .A(n14607), .B(n14606), .Z(n14608) );
  NAND U14896 ( .A(n14609), .B(n14608), .Z(n14729) );
  XNOR U14897 ( .A(n14627), .B(n14626), .Z(n14628) );
  XOR U14898 ( .A(n14629), .B(n14628), .Z(n14635) );
  XOR U14899 ( .A(n14634), .B(n14635), .Z(n14641) );
  XOR U14900 ( .A(n14640), .B(n14641), .Z(n14623) );
  XNOR U14901 ( .A(n14622), .B(n14623), .Z(n14615) );
  XOR U14902 ( .A(n14614), .B(n14615), .Z(n14617) );
  XOR U14903 ( .A(n14616), .B(n14617), .Z(n14613) );
  XNOR U14904 ( .A(n14612), .B(n14613), .Z(n14610) );
  XOR U14905 ( .A(n14611), .B(n14610), .Z(N318) );
  NAND U14906 ( .A(n14615), .B(n14614), .Z(n14619) );
  NAND U14907 ( .A(n14617), .B(n14616), .Z(n14618) );
  AND U14908 ( .A(n14619), .B(n14618), .Z(n15070) );
  XNOR U14909 ( .A(n15071), .B(n15070), .Z(n15069) );
  NANDN U14910 ( .A(n14621), .B(n14620), .Z(n14625) );
  NANDN U14911 ( .A(n14623), .B(n14622), .Z(n14624) );
  AND U14912 ( .A(n14625), .B(n14624), .Z(n14785) );
  NANDN U14913 ( .A(n14627), .B(n14626), .Z(n14631) );
  NANDN U14914 ( .A(n14629), .B(n14628), .Z(n14630) );
  AND U14915 ( .A(n14631), .B(n14630), .Z(n15075) );
  NANDN U14916 ( .A(n14633), .B(n14632), .Z(n14637) );
  NANDN U14917 ( .A(n14635), .B(n14634), .Z(n14636) );
  AND U14918 ( .A(n14637), .B(n14636), .Z(n15077) );
  NANDN U14919 ( .A(n14639), .B(n14638), .Z(n14643) );
  NANDN U14920 ( .A(n14641), .B(n14640), .Z(n14642) );
  AND U14921 ( .A(n14643), .B(n14642), .Z(n15076) );
  XOR U14922 ( .A(n15077), .B(n15076), .Z(n15074) );
  XOR U14923 ( .A(n15075), .B(n15074), .Z(n14787) );
  NANDN U14924 ( .A(n14645), .B(n14644), .Z(n14649) );
  NANDN U14925 ( .A(n14647), .B(n14646), .Z(n14648) );
  AND U14926 ( .A(n14649), .B(n14648), .Z(n15061) );
  NANDN U14927 ( .A(n14651), .B(n14650), .Z(n14655) );
  NAND U14928 ( .A(n14653), .B(n14652), .Z(n14654) );
  AND U14929 ( .A(n14655), .B(n14654), .Z(n15048) );
  NAND U14930 ( .A(n14657), .B(n14656), .Z(n14661) );
  NAND U14931 ( .A(n14659), .B(n14658), .Z(n14660) );
  AND U14932 ( .A(n14661), .B(n14660), .Z(n14792) );
  NAND U14933 ( .A(n14663), .B(n14662), .Z(n14667) );
  NAND U14934 ( .A(n14665), .B(n14664), .Z(n14666) );
  NAND U14935 ( .A(n14667), .B(n14666), .Z(n14805) );
  AND U14936 ( .A(x[134]), .B(y[792]), .Z(n14846) );
  AND U14937 ( .A(x[133]), .B(y[793]), .Z(n14848) );
  AND U14938 ( .A(x[147]), .B(y[779]), .Z(n14847) );
  XOR U14939 ( .A(n14848), .B(n14847), .Z(n14845) );
  XNOR U14940 ( .A(n14846), .B(n14845), .Z(n14808) );
  AND U14941 ( .A(x[132]), .B(y[794]), .Z(n14882) );
  AND U14942 ( .A(x[131]), .B(y[795]), .Z(n14884) );
  AND U14943 ( .A(x[146]), .B(y[780]), .Z(n14883) );
  XOR U14944 ( .A(n14884), .B(n14883), .Z(n14881) );
  XOR U14945 ( .A(n14882), .B(n14881), .Z(n14811) );
  NAND U14946 ( .A(n14669), .B(n14668), .Z(n14673) );
  NAND U14947 ( .A(n14671), .B(n14670), .Z(n14672) );
  AND U14948 ( .A(n14673), .B(n14672), .Z(n14810) );
  XOR U14949 ( .A(n14808), .B(n14809), .Z(n14804) );
  XOR U14950 ( .A(n14805), .B(n14804), .Z(n14803) );
  NAND U14951 ( .A(n14675), .B(n14674), .Z(n14679) );
  NAND U14952 ( .A(n14677), .B(n14676), .Z(n14678) );
  NAND U14953 ( .A(n14679), .B(n14678), .Z(n14802) );
  XOR U14954 ( .A(n14803), .B(n14802), .Z(n14793) );
  NAND U14955 ( .A(n14681), .B(n14680), .Z(n14685) );
  NAND U14956 ( .A(n14683), .B(n14682), .Z(n14684) );
  AND U14957 ( .A(n14685), .B(n14684), .Z(n14790) );
  XOR U14958 ( .A(n14791), .B(n14790), .Z(n15051) );
  AND U14959 ( .A(n14687), .B(n14686), .Z(n14691) );
  NAND U14960 ( .A(n14689), .B(n14688), .Z(n14690) );
  NANDN U14961 ( .A(n14691), .B(n14690), .Z(n14828) );
  AND U14962 ( .A(n14836), .B(n14692), .Z(n14696) );
  NAND U14963 ( .A(n14694), .B(n14693), .Z(n14695) );
  NANDN U14964 ( .A(n14696), .B(n14695), .Z(n14831) );
  NANDN U14965 ( .A(n14878), .B(n14697), .Z(n14701) );
  NANDN U14966 ( .A(n14699), .B(n14698), .Z(n14700) );
  AND U14967 ( .A(n14701), .B(n14700), .Z(n14991) );
  AND U14968 ( .A(x[151]), .B(y[775]), .Z(n14973) );
  AND U14969 ( .A(y[774]), .B(x[152]), .Z(n14703) );
  AND U14970 ( .A(y[773]), .B(x[153]), .Z(n14702) );
  XOR U14971 ( .A(n14703), .B(n14702), .Z(n14972) );
  XOR U14972 ( .A(n14973), .B(n14972), .Z(n14993) );
  AND U14973 ( .A(n14704), .B(o[157]), .Z(n14959) );
  AND U14974 ( .A(x[156]), .B(y[770]), .Z(n14961) );
  AND U14975 ( .A(x[144]), .B(y[782]), .Z(n14960) );
  XOR U14976 ( .A(n14961), .B(n14960), .Z(n14958) );
  XNOR U14977 ( .A(n14959), .B(n14958), .Z(n14992) );
  XNOR U14978 ( .A(n14991), .B(n14990), .Z(n14830) );
  XOR U14979 ( .A(n14831), .B(n14830), .Z(n14829) );
  XOR U14980 ( .A(n14828), .B(n14829), .Z(n15031) );
  NAND U14981 ( .A(n14706), .B(n14705), .Z(n14710) );
  NAND U14982 ( .A(n14708), .B(n14707), .Z(n14709) );
  NAND U14983 ( .A(n14710), .B(n14709), .Z(n15032) );
  NAND U14984 ( .A(n14711), .B(n14975), .Z(n14715) );
  NAND U14985 ( .A(n14713), .B(n14712), .Z(n14714) );
  NAND U14986 ( .A(n14715), .B(n14714), .Z(n14799) );
  NAND U14987 ( .A(n14717), .B(n14716), .Z(n14721) );
  NAND U14988 ( .A(n14719), .B(n14718), .Z(n14720) );
  AND U14989 ( .A(n14721), .B(n14720), .Z(n14985) );
  AND U14990 ( .A(x[128]), .B(y[798]), .Z(n14890) );
  AND U14991 ( .A(x[157]), .B(y[769]), .Z(n14895) );
  XOR U14992 ( .A(o[158]), .B(n14895), .Z(n14892) );
  AND U14993 ( .A(x[158]), .B(y[768]), .Z(n14891) );
  XOR U14994 ( .A(n14892), .B(n14891), .Z(n14889) );
  XOR U14995 ( .A(n14890), .B(n14889), .Z(n14987) );
  AND U14996 ( .A(x[148]), .B(y[778]), .Z(n14968) );
  XOR U14997 ( .A(n14969), .B(n14968), .Z(n14967) );
  AND U14998 ( .A(x[136]), .B(y[790]), .Z(n14966) );
  XNOR U14999 ( .A(n14967), .B(n14966), .Z(n14986) );
  XNOR U15000 ( .A(n14985), .B(n14984), .Z(n14798) );
  XOR U15001 ( .A(n14799), .B(n14798), .Z(n14796) );
  AND U15002 ( .A(x[135]), .B(y[791]), .Z(n14877) );
  NAND U15003 ( .A(n14722), .B(n14877), .Z(n14726) );
  NAND U15004 ( .A(n14724), .B(n14723), .Z(n14725) );
  AND U15005 ( .A(n14726), .B(n14725), .Z(n14820) );
  AND U15006 ( .A(x[149]), .B(y[777]), .Z(n14728) );
  AND U15007 ( .A(y[776]), .B(x[150]), .Z(n14727) );
  XOR U15008 ( .A(n14728), .B(n14727), .Z(n14876) );
  XOR U15009 ( .A(n14877), .B(n14876), .Z(n14823) );
  AND U15010 ( .A(x[145]), .B(y[781]), .Z(n14953) );
  AND U15011 ( .A(x[130]), .B(y[796]), .Z(n14955) );
  AND U15012 ( .A(x[154]), .B(y[772]), .Z(n14954) );
  XOR U15013 ( .A(n14955), .B(n14954), .Z(n14952) );
  XNOR U15014 ( .A(n14953), .B(n14952), .Z(n14822) );
  XNOR U15015 ( .A(n14820), .B(n14821), .Z(n14797) );
  XOR U15016 ( .A(n15032), .B(n15033), .Z(n15030) );
  XOR U15017 ( .A(n15031), .B(n15030), .Z(n15050) );
  XNOR U15018 ( .A(n15048), .B(n15049), .Z(n15063) );
  NANDN U15019 ( .A(n14730), .B(n14729), .Z(n14734) );
  NANDN U15020 ( .A(n14732), .B(n14731), .Z(n14733) );
  NAND U15021 ( .A(n14734), .B(n14733), .Z(n15060) );
  XOR U15022 ( .A(n15063), .B(n15060), .Z(n14735) );
  XOR U15023 ( .A(n15061), .B(n14735), .Z(n15042) );
  NANDN U15024 ( .A(n14737), .B(n14736), .Z(n14741) );
  NANDN U15025 ( .A(n14739), .B(n14738), .Z(n14740) );
  NAND U15026 ( .A(n14741), .B(n14740), .Z(n15044) );
  NANDN U15027 ( .A(n14743), .B(n14742), .Z(n14747) );
  NAND U15028 ( .A(n14745), .B(n14744), .Z(n14746) );
  AND U15029 ( .A(n14747), .B(n14746), .Z(n15025) );
  NAND U15030 ( .A(n14749), .B(n14748), .Z(n14753) );
  NAND U15031 ( .A(n14751), .B(n14750), .Z(n14752) );
  AND U15032 ( .A(n14753), .B(n14752), .Z(n15015) );
  NAND U15033 ( .A(n14755), .B(n14754), .Z(n14759) );
  NANDN U15034 ( .A(n14757), .B(n14756), .Z(n14758) );
  AND U15035 ( .A(n14759), .B(n14758), .Z(n15014) );
  XOR U15036 ( .A(n15015), .B(n15014), .Z(n15013) );
  NANDN U15037 ( .A(n14761), .B(n14760), .Z(n14765) );
  OR U15038 ( .A(n14763), .B(n14762), .Z(n14764) );
  NAND U15039 ( .A(n14765), .B(n14764), .Z(n15012) );
  XOR U15040 ( .A(n15013), .B(n15012), .Z(n15027) );
  NAND U15041 ( .A(n14769), .B(n14768), .Z(n14773) );
  NAND U15042 ( .A(n14771), .B(n14770), .Z(n14772) );
  NAND U15043 ( .A(n14773), .B(n14772), .Z(n14814) );
  AND U15044 ( .A(y[786]), .B(x[140]), .Z(n14774) );
  XOR U15045 ( .A(n14775), .B(n14774), .Z(n14834) );
  XOR U15046 ( .A(n14835), .B(n14834), .Z(n14872) );
  AND U15047 ( .A(x[137]), .B(y[789]), .Z(n14777) );
  XOR U15048 ( .A(n14777), .B(n14776), .Z(n14871) );
  XOR U15049 ( .A(n14872), .B(n14871), .Z(n14817) );
  AND U15050 ( .A(x[155]), .B(y[771]), .Z(n14842) );
  AND U15051 ( .A(x[129]), .B(y[797]), .Z(n14841) );
  XOR U15052 ( .A(n14842), .B(n14841), .Z(n14839) );
  XOR U15053 ( .A(n14840), .B(n14839), .Z(n14816) );
  XOR U15054 ( .A(n14817), .B(n14816), .Z(n14815) );
  XOR U15055 ( .A(n14814), .B(n14815), .Z(n15009) );
  NAND U15056 ( .A(n14779), .B(n14778), .Z(n14783) );
  NANDN U15057 ( .A(n14781), .B(n14780), .Z(n14782) );
  AND U15058 ( .A(n14783), .B(n14782), .Z(n15006) );
  XNOR U15059 ( .A(n15007), .B(n15006), .Z(n15026) );
  XOR U15060 ( .A(n15025), .B(n15024), .Z(n15045) );
  XNOR U15061 ( .A(n15044), .B(n15045), .Z(n15043) );
  XOR U15062 ( .A(n14785), .B(n14784), .Z(n15068) );
  XNOR U15063 ( .A(n15069), .B(n15068), .Z(N319) );
  NANDN U15064 ( .A(n14785), .B(n14784), .Z(n14789) );
  NANDN U15065 ( .A(n14787), .B(n14786), .Z(n14788) );
  AND U15066 ( .A(n14789), .B(n14788), .Z(n15085) );
  NAND U15067 ( .A(n14791), .B(n14790), .Z(n14795) );
  NANDN U15068 ( .A(n14793), .B(n14792), .Z(n14794) );
  AND U15069 ( .A(n14795), .B(n14794), .Z(n15059) );
  NANDN U15070 ( .A(n14797), .B(n14796), .Z(n14801) );
  NAND U15071 ( .A(n14799), .B(n14798), .Z(n14800) );
  AND U15072 ( .A(n14801), .B(n14800), .Z(n15041) );
  NAND U15073 ( .A(n14803), .B(n14802), .Z(n14807) );
  NAND U15074 ( .A(n14805), .B(n14804), .Z(n14806) );
  AND U15075 ( .A(n14807), .B(n14806), .Z(n15023) );
  NANDN U15076 ( .A(n14809), .B(n14808), .Z(n14813) );
  NANDN U15077 ( .A(n14811), .B(n14810), .Z(n14812) );
  AND U15078 ( .A(n14813), .B(n14812), .Z(n15005) );
  NAND U15079 ( .A(n14815), .B(n14814), .Z(n14819) );
  NAND U15080 ( .A(n14817), .B(n14816), .Z(n14818) );
  AND U15081 ( .A(n14819), .B(n14818), .Z(n14827) );
  NANDN U15082 ( .A(n14821), .B(n14820), .Z(n14825) );
  NANDN U15083 ( .A(n14823), .B(n14822), .Z(n14824) );
  NAND U15084 ( .A(n14825), .B(n14824), .Z(n14826) );
  XNOR U15085 ( .A(n14827), .B(n14826), .Z(n15003) );
  NAND U15086 ( .A(n14829), .B(n14828), .Z(n14833) );
  NAND U15087 ( .A(n14831), .B(n14830), .Z(n14832) );
  AND U15088 ( .A(n14833), .B(n14832), .Z(n15001) );
  NAND U15089 ( .A(n14835), .B(n14834), .Z(n14838) );
  NAND U15090 ( .A(n14836), .B(n14919), .Z(n14837) );
  AND U15091 ( .A(n14838), .B(n14837), .Z(n14870) );
  NAND U15092 ( .A(n14840), .B(n14839), .Z(n14844) );
  NAND U15093 ( .A(n14842), .B(n14841), .Z(n14843) );
  AND U15094 ( .A(n14844), .B(n14843), .Z(n14852) );
  NAND U15095 ( .A(n14846), .B(n14845), .Z(n14850) );
  NAND U15096 ( .A(n14848), .B(n14847), .Z(n14849) );
  NAND U15097 ( .A(n14850), .B(n14849), .Z(n14851) );
  XNOR U15098 ( .A(n14852), .B(n14851), .Z(n14868) );
  AND U15099 ( .A(y[771]), .B(x[156]), .Z(n14854) );
  NAND U15100 ( .A(y[773]), .B(x[154]), .Z(n14853) );
  XNOR U15101 ( .A(n14854), .B(n14853), .Z(n14858) );
  AND U15102 ( .A(y[787]), .B(x[140]), .Z(n14856) );
  NAND U15103 ( .A(y[788]), .B(x[139]), .Z(n14855) );
  XNOR U15104 ( .A(n14856), .B(n14855), .Z(n14857) );
  XOR U15105 ( .A(n14858), .B(n14857), .Z(n14866) );
  AND U15106 ( .A(y[799]), .B(x[128]), .Z(n14860) );
  NAND U15107 ( .A(y[798]), .B(x[129]), .Z(n14859) );
  XNOR U15108 ( .A(n14860), .B(n14859), .Z(n14864) );
  AND U15109 ( .A(y[778]), .B(x[149]), .Z(n14862) );
  NAND U15110 ( .A(y[783]), .B(x[144]), .Z(n14861) );
  XNOR U15111 ( .A(n14862), .B(n14861), .Z(n14863) );
  XNOR U15112 ( .A(n14864), .B(n14863), .Z(n14865) );
  XNOR U15113 ( .A(n14866), .B(n14865), .Z(n14867) );
  XNOR U15114 ( .A(n14868), .B(n14867), .Z(n14869) );
  XNOR U15115 ( .A(n14870), .B(n14869), .Z(n14951) );
  NAND U15116 ( .A(n14872), .B(n14871), .Z(n14875) );
  AND U15117 ( .A(x[138]), .B(y[789]), .Z(n14918) );
  NANDN U15118 ( .A(n14873), .B(n14918), .Z(n14874) );
  AND U15119 ( .A(n14875), .B(n14874), .Z(n14949) );
  NAND U15120 ( .A(n14877), .B(n14876), .Z(n14880) );
  AND U15121 ( .A(x[150]), .B(y[777]), .Z(n14896) );
  NANDN U15122 ( .A(n14878), .B(n14896), .Z(n14879) );
  AND U15123 ( .A(n14880), .B(n14879), .Z(n14888) );
  NAND U15124 ( .A(n14882), .B(n14881), .Z(n14886) );
  NAND U15125 ( .A(n14884), .B(n14883), .Z(n14885) );
  NAND U15126 ( .A(n14886), .B(n14885), .Z(n14887) );
  XNOR U15127 ( .A(n14888), .B(n14887), .Z(n14947) );
  NAND U15128 ( .A(n14890), .B(n14889), .Z(n14894) );
  NAND U15129 ( .A(n14892), .B(n14891), .Z(n14893) );
  AND U15130 ( .A(n14894), .B(n14893), .Z(n14945) );
  AND U15131 ( .A(y[785]), .B(x[142]), .Z(n14903) );
  AND U15132 ( .A(n14895), .B(o[158]), .Z(n14901) );
  XOR U15133 ( .A(n14896), .B(o[159]), .Z(n14899) );
  AND U15134 ( .A(x[153]), .B(y[774]), .Z(n14974) );
  XNOR U15135 ( .A(n14897), .B(n14974), .Z(n14898) );
  XNOR U15136 ( .A(n14899), .B(n14898), .Z(n14900) );
  XNOR U15137 ( .A(n14901), .B(n14900), .Z(n14902) );
  XNOR U15138 ( .A(n14903), .B(n14902), .Z(n14943) );
  AND U15139 ( .A(y[780]), .B(x[147]), .Z(n14909) );
  AND U15140 ( .A(y[782]), .B(x[145]), .Z(n14905) );
  NAND U15141 ( .A(y[791]), .B(x[136]), .Z(n14904) );
  XNOR U15142 ( .A(n14905), .B(n14904), .Z(n14906) );
  XNOR U15143 ( .A(n14907), .B(n14906), .Z(n14908) );
  XNOR U15144 ( .A(n14909), .B(n14908), .Z(n14933) );
  AND U15145 ( .A(y[793]), .B(x[134]), .Z(n14911) );
  NAND U15146 ( .A(y[792]), .B(x[135]), .Z(n14910) );
  XNOR U15147 ( .A(n14911), .B(n14910), .Z(n14923) );
  AND U15148 ( .A(y[794]), .B(x[133]), .Z(n14913) );
  NAND U15149 ( .A(y[781]), .B(x[146]), .Z(n14912) );
  XNOR U15150 ( .A(n14913), .B(n14912), .Z(n14917) );
  AND U15151 ( .A(y[796]), .B(x[131]), .Z(n14915) );
  NAND U15152 ( .A(y[795]), .B(x[132]), .Z(n14914) );
  XNOR U15153 ( .A(n14915), .B(n14914), .Z(n14916) );
  XOR U15154 ( .A(n14917), .B(n14916), .Z(n14921) );
  XNOR U15155 ( .A(n14919), .B(n14918), .Z(n14920) );
  XNOR U15156 ( .A(n14921), .B(n14920), .Z(n14922) );
  XOR U15157 ( .A(n14923), .B(n14922), .Z(n14931) );
  AND U15158 ( .A(y[769]), .B(x[158]), .Z(n14925) );
  NAND U15159 ( .A(y[790]), .B(x[137]), .Z(n14924) );
  XNOR U15160 ( .A(n14925), .B(n14924), .Z(n14929) );
  AND U15161 ( .A(y[770]), .B(x[157]), .Z(n14927) );
  NAND U15162 ( .A(y[779]), .B(x[148]), .Z(n14926) );
  XNOR U15163 ( .A(n14927), .B(n14926), .Z(n14928) );
  XNOR U15164 ( .A(n14929), .B(n14928), .Z(n14930) );
  XNOR U15165 ( .A(n14931), .B(n14930), .Z(n14932) );
  XOR U15166 ( .A(n14933), .B(n14932), .Z(n14941) );
  AND U15167 ( .A(y[768]), .B(x[159]), .Z(n14935) );
  NAND U15168 ( .A(y[772]), .B(x[155]), .Z(n14934) );
  XNOR U15169 ( .A(n14935), .B(n14934), .Z(n14939) );
  AND U15170 ( .A(y[797]), .B(x[130]), .Z(n14937) );
  NAND U15171 ( .A(y[776]), .B(x[151]), .Z(n14936) );
  XNOR U15172 ( .A(n14937), .B(n14936), .Z(n14938) );
  XNOR U15173 ( .A(n14939), .B(n14938), .Z(n14940) );
  XNOR U15174 ( .A(n14941), .B(n14940), .Z(n14942) );
  XNOR U15175 ( .A(n14943), .B(n14942), .Z(n14944) );
  XNOR U15176 ( .A(n14945), .B(n14944), .Z(n14946) );
  XNOR U15177 ( .A(n14947), .B(n14946), .Z(n14948) );
  XNOR U15178 ( .A(n14949), .B(n14948), .Z(n14950) );
  XOR U15179 ( .A(n14951), .B(n14950), .Z(n14983) );
  NAND U15180 ( .A(n14953), .B(n14952), .Z(n14957) );
  NAND U15181 ( .A(n14955), .B(n14954), .Z(n14956) );
  AND U15182 ( .A(n14957), .B(n14956), .Z(n14965) );
  NAND U15183 ( .A(n14959), .B(n14958), .Z(n14963) );
  NAND U15184 ( .A(n14961), .B(n14960), .Z(n14962) );
  NAND U15185 ( .A(n14963), .B(n14962), .Z(n14964) );
  XNOR U15186 ( .A(n14965), .B(n14964), .Z(n14981) );
  NAND U15187 ( .A(n14967), .B(n14966), .Z(n14971) );
  NAND U15188 ( .A(n14969), .B(n14968), .Z(n14970) );
  AND U15189 ( .A(n14971), .B(n14970), .Z(n14979) );
  NAND U15190 ( .A(n14973), .B(n14972), .Z(n14977) );
  NAND U15191 ( .A(n14975), .B(n14974), .Z(n14976) );
  NAND U15192 ( .A(n14977), .B(n14976), .Z(n14978) );
  XNOR U15193 ( .A(n14979), .B(n14978), .Z(n14980) );
  XNOR U15194 ( .A(n14981), .B(n14980), .Z(n14982) );
  XNOR U15195 ( .A(n14983), .B(n14982), .Z(n14999) );
  NAND U15196 ( .A(n14985), .B(n14984), .Z(n14989) );
  NANDN U15197 ( .A(n14987), .B(n14986), .Z(n14988) );
  AND U15198 ( .A(n14989), .B(n14988), .Z(n14997) );
  NAND U15199 ( .A(n14991), .B(n14990), .Z(n14995) );
  NANDN U15200 ( .A(n14993), .B(n14992), .Z(n14994) );
  NAND U15201 ( .A(n14995), .B(n14994), .Z(n14996) );
  XNOR U15202 ( .A(n14997), .B(n14996), .Z(n14998) );
  XNOR U15203 ( .A(n14999), .B(n14998), .Z(n15000) );
  XNOR U15204 ( .A(n15001), .B(n15000), .Z(n15002) );
  XNOR U15205 ( .A(n15003), .B(n15002), .Z(n15004) );
  XNOR U15206 ( .A(n15005), .B(n15004), .Z(n15021) );
  NAND U15207 ( .A(n15007), .B(n15006), .Z(n15011) );
  NANDN U15208 ( .A(n15009), .B(n15008), .Z(n15010) );
  AND U15209 ( .A(n15011), .B(n15010), .Z(n15019) );
  NAND U15210 ( .A(n15013), .B(n15012), .Z(n15017) );
  NAND U15211 ( .A(n15015), .B(n15014), .Z(n15016) );
  NAND U15212 ( .A(n15017), .B(n15016), .Z(n15018) );
  XNOR U15213 ( .A(n15019), .B(n15018), .Z(n15020) );
  XNOR U15214 ( .A(n15021), .B(n15020), .Z(n15022) );
  XNOR U15215 ( .A(n15023), .B(n15022), .Z(n15039) );
  NAND U15216 ( .A(n15025), .B(n15024), .Z(n15029) );
  NANDN U15217 ( .A(n15027), .B(n15026), .Z(n15028) );
  AND U15218 ( .A(n15029), .B(n15028), .Z(n15037) );
  NAND U15219 ( .A(n15031), .B(n15030), .Z(n15035) );
  NAND U15220 ( .A(n15033), .B(n15032), .Z(n15034) );
  NAND U15221 ( .A(n15035), .B(n15034), .Z(n15036) );
  XNOR U15222 ( .A(n15037), .B(n15036), .Z(n15038) );
  XNOR U15223 ( .A(n15039), .B(n15038), .Z(n15040) );
  XNOR U15224 ( .A(n15041), .B(n15040), .Z(n15057) );
  NANDN U15225 ( .A(n15043), .B(n15042), .Z(n15047) );
  NAND U15226 ( .A(n15045), .B(n15044), .Z(n15046) );
  AND U15227 ( .A(n15047), .B(n15046), .Z(n15055) );
  NANDN U15228 ( .A(n15049), .B(n15048), .Z(n15053) );
  NANDN U15229 ( .A(n15051), .B(n15050), .Z(n15052) );
  NAND U15230 ( .A(n15053), .B(n15052), .Z(n15054) );
  XNOR U15231 ( .A(n15055), .B(n15054), .Z(n15056) );
  XNOR U15232 ( .A(n15057), .B(n15056), .Z(n15058) );
  XNOR U15233 ( .A(n15059), .B(n15058), .Z(n15067) );
  OR U15234 ( .A(n15060), .B(n15061), .Z(n15065) );
  AND U15235 ( .A(n15061), .B(n15060), .Z(n15062) );
  OR U15236 ( .A(n15063), .B(n15062), .Z(n15064) );
  NAND U15237 ( .A(n15065), .B(n15064), .Z(n15066) );
  XNOR U15238 ( .A(n15067), .B(n15066), .Z(n15083) );
  NAND U15239 ( .A(n15069), .B(n15068), .Z(n15073) );
  NANDN U15240 ( .A(n15071), .B(n15070), .Z(n15072) );
  AND U15241 ( .A(n15073), .B(n15072), .Z(n15081) );
  NAND U15242 ( .A(n15075), .B(n15074), .Z(n15079) );
  NAND U15243 ( .A(n15077), .B(n15076), .Z(n15078) );
  NAND U15244 ( .A(n15079), .B(n15078), .Z(n15080) );
  XNOR U15245 ( .A(n15081), .B(n15080), .Z(n15082) );
  XNOR U15246 ( .A(n15083), .B(n15082), .Z(n15084) );
  XNOR U15247 ( .A(n15085), .B(n15084), .Z(N320) );
endmodule

