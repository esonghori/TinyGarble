
module hamming_N16000_CC64_DW01_add_0 ( A, B, CI, SUM, CO );
  input [13:0] A;
  input [13:0] B;
  output [13:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41;

  XOR U1 ( .A(A[9]), .B(n1), .Z(SUM[9]) );
  XOR U2 ( .A(A[8]), .B(n2), .Z(SUM[8]) );
  XOR U3 ( .A(n3), .B(n4), .Z(SUM[7]) );
  XNOR U4 ( .A(B[7]), .B(A[7]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[5]) );
  XNOR U8 ( .A(B[5]), .B(A[5]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U14 ( .A(B[2]), .B(A[2]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[1]) );
  XOR U16 ( .A(B[1]), .B(A[1]), .Z(n16) );
  XOR U17 ( .A(A[13]), .B(n17), .Z(SUM[13]) );
  ANDN U18 ( .B(A[12]), .A(n18), .Z(n17) );
  XNOR U19 ( .A(A[12]), .B(n18), .Z(SUM[12]) );
  NAND U20 ( .A(n19), .B(A[11]), .Z(n18) );
  XOR U21 ( .A(A[11]), .B(n19), .Z(SUM[11]) );
  ANDN U22 ( .B(A[10]), .A(n20), .Z(n19) );
  XNOR U23 ( .A(A[10]), .B(n20), .Z(SUM[10]) );
  NAND U24 ( .A(n1), .B(A[9]), .Z(n20) );
  AND U25 ( .A(A[8]), .B(n2), .Z(n1) );
  NAND U26 ( .A(n21), .B(n22), .Z(n2) );
  NAND U27 ( .A(n23), .B(B[7]), .Z(n22) );
  NANDN U28 ( .A(A[7]), .B(n3), .Z(n23) );
  NANDN U29 ( .A(n3), .B(A[7]), .Z(n21) );
  AND U30 ( .A(n24), .B(n25), .Z(n3) );
  NAND U31 ( .A(n26), .B(B[6]), .Z(n25) );
  NANDN U32 ( .A(A[6]), .B(n5), .Z(n26) );
  NANDN U33 ( .A(n5), .B(A[6]), .Z(n24) );
  AND U34 ( .A(n27), .B(n28), .Z(n5) );
  NAND U35 ( .A(n29), .B(B[5]), .Z(n28) );
  NANDN U36 ( .A(A[5]), .B(n7), .Z(n29) );
  NANDN U37 ( .A(n7), .B(A[5]), .Z(n27) );
  AND U38 ( .A(n30), .B(n31), .Z(n7) );
  NAND U39 ( .A(n32), .B(B[4]), .Z(n31) );
  NANDN U40 ( .A(A[4]), .B(n9), .Z(n32) );
  NANDN U41 ( .A(n9), .B(A[4]), .Z(n30) );
  AND U42 ( .A(n33), .B(n34), .Z(n9) );
  NAND U43 ( .A(n35), .B(B[3]), .Z(n34) );
  NANDN U44 ( .A(A[3]), .B(n11), .Z(n35) );
  NANDN U45 ( .A(n11), .B(A[3]), .Z(n33) );
  AND U46 ( .A(n36), .B(n37), .Z(n11) );
  NAND U47 ( .A(n38), .B(B[2]), .Z(n37) );
  NANDN U48 ( .A(A[2]), .B(n13), .Z(n38) );
  NANDN U49 ( .A(n13), .B(A[2]), .Z(n36) );
  AND U50 ( .A(n39), .B(n40), .Z(n13) );
  NAND U51 ( .A(n41), .B(B[1]), .Z(n40) );
  OR U52 ( .A(n15), .B(A[1]), .Z(n41) );
  NAND U53 ( .A(n15), .B(A[1]), .Z(n39) );
  AND U54 ( .A(B[0]), .B(A[0]), .Z(n15) );
  XOR U55 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC64_DW01_add_1 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32;

  IV U1 ( .A(B[7]), .Z(n1) );
  XOR U2 ( .A(n2), .B(n1), .Z(SUM[7]) );
  AND U3 ( .A(n3), .B(n4), .Z(n2) );
  NAND U4 ( .A(n5), .B(B[6]), .Z(n4) );
  NANDN U5 ( .A(A[6]), .B(n6), .Z(n5) );
  NANDN U6 ( .A(n6), .B(A[6]), .Z(n3) );
  XOR U7 ( .A(n6), .B(n7), .Z(SUM[6]) );
  XNOR U8 ( .A(B[6]), .B(A[6]), .Z(n7) );
  AND U9 ( .A(n8), .B(n9), .Z(n6) );
  NAND U10 ( .A(n10), .B(B[5]), .Z(n9) );
  NANDN U11 ( .A(A[5]), .B(n11), .Z(n10) );
  NANDN U12 ( .A(n11), .B(A[5]), .Z(n8) );
  XOR U13 ( .A(n11), .B(n12), .Z(SUM[5]) );
  XNOR U14 ( .A(B[5]), .B(A[5]), .Z(n12) );
  AND U15 ( .A(n13), .B(n14), .Z(n11) );
  NAND U16 ( .A(n15), .B(B[4]), .Z(n14) );
  NANDN U17 ( .A(A[4]), .B(n16), .Z(n15) );
  NANDN U18 ( .A(n16), .B(A[4]), .Z(n13) );
  XOR U19 ( .A(n16), .B(n17), .Z(SUM[4]) );
  XNOR U20 ( .A(B[4]), .B(A[4]), .Z(n17) );
  AND U21 ( .A(n18), .B(n19), .Z(n16) );
  NAND U22 ( .A(n20), .B(B[3]), .Z(n19) );
  NANDN U23 ( .A(A[3]), .B(n21), .Z(n20) );
  NANDN U24 ( .A(n21), .B(A[3]), .Z(n18) );
  XOR U25 ( .A(n21), .B(n22), .Z(SUM[3]) );
  XNOR U26 ( .A(B[3]), .B(A[3]), .Z(n22) );
  AND U27 ( .A(n23), .B(n24), .Z(n21) );
  NAND U28 ( .A(n25), .B(B[2]), .Z(n24) );
  NANDN U29 ( .A(A[2]), .B(n26), .Z(n25) );
  NANDN U30 ( .A(n26), .B(A[2]), .Z(n23) );
  XOR U31 ( .A(n26), .B(n27), .Z(SUM[2]) );
  XNOR U32 ( .A(B[2]), .B(A[2]), .Z(n27) );
  AND U33 ( .A(n28), .B(n29), .Z(n26) );
  NAND U34 ( .A(n30), .B(B[1]), .Z(n29) );
  OR U35 ( .A(n31), .B(A[1]), .Z(n30) );
  NAND U36 ( .A(n31), .B(A[1]), .Z(n28) );
  XOR U37 ( .A(n31), .B(n32), .Z(SUM[1]) );
  XOR U38 ( .A(B[1]), .B(A[1]), .Z(n32) );
  AND U39 ( .A(B[0]), .B(A[0]), .Z(n31) );
  XOR U40 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC64_DW01_add_2 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[7]) );
  NAND U2 ( .A(n4), .B(B[6]), .Z(n3) );
  NANDN U3 ( .A(A[6]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[6]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[6]) );
  XNOR U6 ( .A(B[6]), .B(A[6]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[5]), .Z(n8) );
  NANDN U9 ( .A(A[5]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[5]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[5]) );
  XNOR U12 ( .A(B[5]), .B(A[5]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[4]), .Z(n13) );
  NANDN U15 ( .A(A[4]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[4]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[4]) );
  XNOR U18 ( .A(B[4]), .B(A[4]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[3]), .Z(n18) );
  NANDN U21 ( .A(A[3]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[3]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[3]) );
  XNOR U24 ( .A(B[3]), .B(A[3]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[2]), .Z(n23) );
  NANDN U27 ( .A(A[2]), .B(n25), .Z(n24) );
  NANDN U28 ( .A(n25), .B(A[2]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[2]) );
  XNOR U30 ( .A(B[2]), .B(A[2]), .Z(n26) );
  AND U31 ( .A(n27), .B(n28), .Z(n25) );
  NAND U32 ( .A(n29), .B(B[1]), .Z(n28) );
  OR U33 ( .A(n30), .B(A[1]), .Z(n29) );
  NAND U34 ( .A(n30), .B(A[1]), .Z(n27) );
  XOR U35 ( .A(n30), .B(n31), .Z(SUM[1]) );
  XOR U36 ( .A(B[1]), .B(A[1]), .Z(n31) );
  AND U37 ( .A(B[0]), .B(A[0]), .Z(n30) );
  XOR U38 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC64_DW01_add_3 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC64_DW01_add_4 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[6]) );
  NAND U2 ( .A(n4), .B(B[5]), .Z(n3) );
  NANDN U3 ( .A(A[5]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[5]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[5]) );
  XNOR U6 ( .A(B[5]), .B(A[5]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[4]), .Z(n8) );
  NANDN U9 ( .A(A[4]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[4]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[4]) );
  XNOR U12 ( .A(B[4]), .B(A[4]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[3]), .Z(n13) );
  NANDN U15 ( .A(A[3]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[3]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[3]) );
  XNOR U18 ( .A(B[3]), .B(A[3]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[2]), .Z(n18) );
  NANDN U21 ( .A(A[2]), .B(n20), .Z(n19) );
  NANDN U22 ( .A(n20), .B(A[2]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[2]) );
  XNOR U24 ( .A(B[2]), .B(A[2]), .Z(n21) );
  AND U25 ( .A(n22), .B(n23), .Z(n20) );
  NAND U26 ( .A(n24), .B(B[1]), .Z(n23) );
  OR U27 ( .A(n25), .B(A[1]), .Z(n24) );
  NAND U28 ( .A(n25), .B(A[1]), .Z(n22) );
  XOR U29 ( .A(n25), .B(n26), .Z(SUM[1]) );
  XOR U30 ( .A(B[1]), .B(A[1]), .Z(n26) );
  AND U31 ( .A(B[0]), .B(A[0]), .Z(n25) );
  XOR U32 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC64_DW01_add_5 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;

  AND U1 ( .A(n2), .B(B[5]), .Z(SUM[6]) );
  IV U2 ( .A(n4), .Z(n2) );
  IV U3 ( .A(B[5]), .Z(n3) );
  XOR U4 ( .A(n4), .B(n3), .Z(SUM[5]) );
  AND U5 ( .A(n5), .B(n6), .Z(n4) );
  NAND U6 ( .A(n7), .B(B[4]), .Z(n6) );
  NANDN U7 ( .A(A[4]), .B(n8), .Z(n7) );
  NANDN U8 ( .A(n8), .B(A[4]), .Z(n5) );
  XOR U9 ( .A(n8), .B(n9), .Z(SUM[4]) );
  XNOR U10 ( .A(B[4]), .B(A[4]), .Z(n9) );
  AND U11 ( .A(n10), .B(n11), .Z(n8) );
  NAND U12 ( .A(n12), .B(B[3]), .Z(n11) );
  NANDN U13 ( .A(A[3]), .B(n13), .Z(n12) );
  NANDN U14 ( .A(n13), .B(A[3]), .Z(n10) );
  XOR U15 ( .A(n13), .B(n14), .Z(SUM[3]) );
  XNOR U16 ( .A(B[3]), .B(A[3]), .Z(n14) );
  AND U17 ( .A(n15), .B(n16), .Z(n13) );
  NAND U18 ( .A(n17), .B(B[2]), .Z(n16) );
  NANDN U19 ( .A(A[2]), .B(n18), .Z(n17) );
  NANDN U20 ( .A(n18), .B(A[2]), .Z(n15) );
  XOR U21 ( .A(n18), .B(n19), .Z(SUM[2]) );
  XNOR U22 ( .A(B[2]), .B(A[2]), .Z(n19) );
  AND U23 ( .A(n20), .B(n21), .Z(n18) );
  NAND U24 ( .A(n22), .B(B[1]), .Z(n21) );
  OR U25 ( .A(n23), .B(A[1]), .Z(n22) );
  NAND U26 ( .A(n23), .B(A[1]), .Z(n20) );
  XOR U27 ( .A(n23), .B(n24), .Z(SUM[1]) );
  XOR U28 ( .A(B[1]), .B(A[1]), .Z(n24) );
  AND U29 ( .A(B[0]), .B(A[0]), .Z(n23) );
  XOR U30 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC64_DW01_add_6 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC64_DW01_add_7 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC64_DW01_add_8 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC64_DW01_add_9 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  NAND U1 ( .A(n2), .B(n3), .Z(SUM[5]) );
  NAND U2 ( .A(n4), .B(B[4]), .Z(n3) );
  NANDN U3 ( .A(A[4]), .B(n5), .Z(n4) );
  NANDN U4 ( .A(n5), .B(A[4]), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[4]) );
  XNOR U6 ( .A(B[4]), .B(A[4]), .Z(n6) );
  AND U7 ( .A(n7), .B(n8), .Z(n5) );
  NAND U8 ( .A(n9), .B(B[3]), .Z(n8) );
  NANDN U9 ( .A(A[3]), .B(n10), .Z(n9) );
  NANDN U10 ( .A(n10), .B(A[3]), .Z(n7) );
  XOR U11 ( .A(n10), .B(n11), .Z(SUM[3]) );
  XNOR U12 ( .A(B[3]), .B(A[3]), .Z(n11) );
  AND U13 ( .A(n12), .B(n13), .Z(n10) );
  NAND U14 ( .A(n14), .B(B[2]), .Z(n13) );
  NANDN U15 ( .A(A[2]), .B(n15), .Z(n14) );
  NANDN U16 ( .A(n15), .B(A[2]), .Z(n12) );
  XOR U17 ( .A(n15), .B(n16), .Z(SUM[2]) );
  XNOR U18 ( .A(B[2]), .B(A[2]), .Z(n16) );
  AND U19 ( .A(n17), .B(n18), .Z(n15) );
  NAND U20 ( .A(n19), .B(B[1]), .Z(n18) );
  OR U21 ( .A(n20), .B(A[1]), .Z(n19) );
  NAND U22 ( .A(n20), .B(A[1]), .Z(n17) );
  XOR U23 ( .A(n20), .B(n21), .Z(SUM[1]) );
  XOR U24 ( .A(B[1]), .B(A[1]), .Z(n21) );
  AND U25 ( .A(B[0]), .B(A[0]), .Z(n20) );
  XOR U26 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC64_DW01_add_10 ( A, B, CI, SUM, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19;

  AND U1 ( .A(n3), .B(B[4]), .Z(SUM[5]) );
  IV U2 ( .A(B[4]), .Z(n2) );
  IV U3 ( .A(n4), .Z(n3) );
  XOR U4 ( .A(n4), .B(n2), .Z(SUM[4]) );
  AND U5 ( .A(n5), .B(n6), .Z(n4) );
  NAND U6 ( .A(n7), .B(B[3]), .Z(n6) );
  NANDN U7 ( .A(A[3]), .B(n8), .Z(n7) );
  NANDN U8 ( .A(n8), .B(A[3]), .Z(n5) );
  XOR U9 ( .A(n8), .B(n9), .Z(SUM[3]) );
  XNOR U10 ( .A(B[3]), .B(A[3]), .Z(n9) );
  AND U11 ( .A(n10), .B(n11), .Z(n8) );
  NAND U12 ( .A(n12), .B(B[2]), .Z(n11) );
  NANDN U13 ( .A(A[2]), .B(n13), .Z(n12) );
  NANDN U14 ( .A(n13), .B(A[2]), .Z(n10) );
  XOR U15 ( .A(n13), .B(n14), .Z(SUM[2]) );
  XNOR U16 ( .A(B[2]), .B(A[2]), .Z(n14) );
  AND U17 ( .A(n15), .B(n16), .Z(n13) );
  NAND U18 ( .A(n17), .B(B[1]), .Z(n16) );
  OR U19 ( .A(n18), .B(A[1]), .Z(n17) );
  NAND U20 ( .A(n18), .B(A[1]), .Z(n15) );
  XOR U21 ( .A(n18), .B(n19), .Z(SUM[1]) );
  XOR U22 ( .A(B[1]), .B(A[1]), .Z(n19) );
  AND U23 ( .A(B[0]), .B(A[0]), .Z(n18) );
  XOR U24 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
endmodule


module hamming_N16000_CC64 ( clk, rst, x, y, o );
  input [249:0] x;
  input [249:0] y;
  output [13:0] o;
  input clk, rst;
  wire   N1131, N1132, N1133, N1134, N1139, N1140, N1141, N1142, N1143, N1147,
         N1148, N1149, N1150, N1151, N1155, N1156, N1157, N1158, N1159, N1163,
         N1164, N1165, N1166, N1167, N1171, N1172, N1173, N1174, N1175, N1179,
         N1180, N1181, N1182, N1183, N1187, N1188, N1189, N1190, N1191, N1195,
         N1196, N1197, N1198, N1199, N1203, N1204, N1205, N1206, N1207, N1211,
         N1212, N1213, N1214, N1215, N1219, N1220, N1221, N1222, N1223, N1224,
         N1227, N1228, N1229, N1230, N1231, N1232, N1235, N1236, N1237, N1238,
         N1239, N1240, N1243, N1244, N1245, N1246, N1247, N1248, N1251, N1252,
         N1253, N1254, N1255, N1256, N1259, N1260, N1261, N1262, N1263, N1264,
         N1265, N1267, N1268, N1269, N1270, N1271, N1272, N1273, N1275, N1276,
         N1277, N1278, N1279, N1280, N1281, N1283, N1284, N1285, N1286, N1287,
         N1288, N1289, N1290, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704;
  wire   [7:0] olocal;
  wire   [13:0] oglobal;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12;

  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  hamming_N16000_CC64_DW01_add_0 add_97 ( .A(oglobal), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, olocal}), .CI(1'b0), .SUM(o) );
  hamming_N16000_CC64_DW01_add_1 add_84_root_add_47_I250 ( .A({1'b0, N1281, 
        N1280, N1279, N1278, N1277, N1276, N1275}), .B({N1290, N1289, N1288, 
        N1287, N1286, N1285, N1284, N1283}), .CI(1'b0), .SUM(olocal) );
  hamming_N16000_CC64_DW01_add_2 add_85_root_add_47_I250 ( .A({1'b0, N1265, 
        N1264, N1263, N1262, N1261, N1260, N1259}), .B({1'b0, N1273, N1272, 
        N1271, N1270, N1269, N1268, N1267}), .CI(1'b0), .SUM({N1290, N1289, 
        N1288, N1287, N1286, N1285, N1284, N1283}) );
  hamming_N16000_CC64_DW01_add_3 add_86_root_add_47_I250 ( .A({1'b0, 1'b0, 
        N1248, N1247, N1246, N1245, N1244, N1243}), .B({1'b0, 1'b0, N1256, 
        N1255, N1254, N1253, N1252, N1251}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__0, N1281, N1280, N1279, N1278, N1277, N1276, 
        N1275}) );
  hamming_N16000_CC64_DW01_add_4 add_87_root_add_47_I250 ( .A({1'b0, 1'b0, 
        N1232, N1231, N1230, N1229, N1228, N1227}), .B({1'b0, 1'b0, N1240, 
        N1239, N1238, N1237, N1236, N1235}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__1, N1273, N1272, N1271, N1270, N1269, N1268, 
        N1267}) );
  hamming_N16000_CC64_DW01_add_5 add_88_root_add_47_I250 ( .A({1'b0, 1'b0, 
        1'b0, N1215, N1214, N1213, N1212, N1211}), .B({1'b0, 1'b0, N1224, 
        N1223, N1222, N1221, N1220, N1219}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__2, N1265, N1264, N1263, N1262, N1261, N1260, 
        N1259}) );
  hamming_N16000_CC64_DW01_add_6 add_89_root_add_47_I250 ( .A({1'b0, 1'b0, 
        1'b0, N1199, N1198, N1197, N1196, N1195}), .B({1'b0, 1'b0, 1'b0, N1207, 
        N1206, N1205, N1204, N1203}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, N1256, N1255, N1254, N1253, N1252, N1251}) );
  hamming_N16000_CC64_DW01_add_7 add_90_root_add_47_I250 ( .A({1'b0, 1'b0, 
        1'b0, N1183, N1182, N1181, N1180, N1179}), .B({1'b0, 1'b0, 1'b0, N1191, 
        N1190, N1189, N1188, N1187}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, N1248, N1247, N1246, N1245, N1244, N1243}) );
  hamming_N16000_CC64_DW01_add_8 add_91_root_add_47_I250 ( .A({1'b0, 1'b0, 
        1'b0, N1167, N1166, N1165, N1164, N1163}), .B({1'b0, 1'b0, 1'b0, N1175, 
        N1174, N1173, N1172, N1171}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, N1240, N1239, N1238, N1237, N1236, N1235}) );
  hamming_N16000_CC64_DW01_add_9 add_92_root_add_47_I250 ( .A({1'b0, 1'b0, 
        1'b0, N1151, N1150, N1149, N1148, N1147}), .B({1'b0, 1'b0, 1'b0, N1159, 
        N1158, N1157, N1156, N1155}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, N1232, N1231, N1230, N1229, N1228, N1227})
         );
  hamming_N16000_CC64_DW01_add_10 add_93_root_add_47_I250 ( .A({1'b0, 1'b0, 
        1'b0, 1'b0, N1134, N1133, N1132, N1131}), .B({1'b0, 1'b0, 1'b0, N1143, 
        N1142, N1141, N1140, N1139}), .CI(1'b0), .SUM({
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, N1224, N1223, 
        N1222, N1221, N1220, N1219}) );
  NAND U436 ( .A(n187), .B(n188), .Z(N1215) );
  NANDN U437 ( .A(n189), .B(n190), .Z(n188) );
  OR U438 ( .A(n191), .B(n192), .Z(n190) );
  NAND U439 ( .A(n191), .B(n192), .Z(n187) );
  XOR U440 ( .A(n191), .B(n193), .Z(N1214) );
  XNOR U441 ( .A(n189), .B(n192), .Z(n193) );
  AND U442 ( .A(n194), .B(n195), .Z(n192) );
  NANDN U443 ( .A(n196), .B(n197), .Z(n195) );
  NANDN U444 ( .A(n198), .B(n199), .Z(n197) );
  NANDN U445 ( .A(n199), .B(n198), .Z(n194) );
  NAND U446 ( .A(n200), .B(n201), .Z(n189) );
  NANDN U447 ( .A(n202), .B(n203), .Z(n201) );
  OR U448 ( .A(n204), .B(n205), .Z(n203) );
  NAND U449 ( .A(n205), .B(n204), .Z(n200) );
  AND U450 ( .A(n206), .B(n207), .Z(n191) );
  NANDN U451 ( .A(n208), .B(n209), .Z(n207) );
  NANDN U452 ( .A(n210), .B(n211), .Z(n209) );
  NANDN U453 ( .A(n211), .B(n210), .Z(n206) );
  XOR U454 ( .A(n205), .B(n212), .Z(N1213) );
  XOR U455 ( .A(n202), .B(n204), .Z(n212) );
  XNOR U456 ( .A(n198), .B(n213), .Z(n204) );
  XNOR U457 ( .A(n196), .B(n199), .Z(n213) );
  NAND U458 ( .A(n214), .B(n215), .Z(n199) );
  NAND U459 ( .A(n216), .B(n217), .Z(n215) );
  OR U460 ( .A(n218), .B(n219), .Z(n216) );
  NANDN U461 ( .A(n220), .B(n218), .Z(n214) );
  IV U462 ( .A(n219), .Z(n220) );
  NAND U463 ( .A(n221), .B(n222), .Z(n196) );
  NAND U464 ( .A(n223), .B(n224), .Z(n222) );
  NANDN U465 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U466 ( .A(n226), .B(n225), .Z(n221) );
  AND U467 ( .A(n227), .B(n228), .Z(n198) );
  NAND U468 ( .A(n229), .B(n230), .Z(n228) );
  OR U469 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U470 ( .A(n233), .B(n231), .Z(n227) );
  NAND U471 ( .A(n234), .B(n235), .Z(n202) );
  NANDN U472 ( .A(n236), .B(n237), .Z(n235) );
  OR U473 ( .A(n238), .B(n239), .Z(n237) );
  NANDN U474 ( .A(n240), .B(n238), .Z(n234) );
  IV U475 ( .A(n239), .Z(n240) );
  XNOR U476 ( .A(n210), .B(n241), .Z(n205) );
  XNOR U477 ( .A(n208), .B(n211), .Z(n241) );
  NAND U478 ( .A(n242), .B(n243), .Z(n211) );
  NAND U479 ( .A(n244), .B(n245), .Z(n243) );
  OR U480 ( .A(n246), .B(n247), .Z(n244) );
  NANDN U481 ( .A(n248), .B(n246), .Z(n242) );
  IV U482 ( .A(n247), .Z(n248) );
  NAND U483 ( .A(n249), .B(n250), .Z(n208) );
  NAND U484 ( .A(n251), .B(n252), .Z(n250) );
  NANDN U485 ( .A(n253), .B(n254), .Z(n251) );
  NANDN U486 ( .A(n254), .B(n253), .Z(n249) );
  AND U487 ( .A(n255), .B(n256), .Z(n210) );
  NAND U488 ( .A(n257), .B(n258), .Z(n256) );
  OR U489 ( .A(n259), .B(n260), .Z(n257) );
  NANDN U490 ( .A(n261), .B(n259), .Z(n255) );
  XNOR U491 ( .A(n236), .B(n262), .Z(N1212) );
  XOR U492 ( .A(n238), .B(n239), .Z(n262) );
  XNOR U493 ( .A(n252), .B(n263), .Z(n239) );
  XOR U494 ( .A(n253), .B(n254), .Z(n263) );
  XOR U495 ( .A(n259), .B(n264), .Z(n254) );
  XOR U496 ( .A(n258), .B(n261), .Z(n264) );
  IV U497 ( .A(n260), .Z(n261) );
  NAND U498 ( .A(n265), .B(n266), .Z(n260) );
  OR U499 ( .A(n267), .B(n268), .Z(n266) );
  OR U500 ( .A(n269), .B(n270), .Z(n265) );
  NAND U501 ( .A(n271), .B(n272), .Z(n258) );
  OR U502 ( .A(n273), .B(n274), .Z(n272) );
  OR U503 ( .A(n275), .B(n276), .Z(n271) );
  NOR U504 ( .A(n277), .B(n278), .Z(n259) );
  ANDN U505 ( .B(n279), .A(n280), .Z(n253) );
  XNOR U506 ( .A(n246), .B(n281), .Z(n252) );
  XNOR U507 ( .A(n245), .B(n247), .Z(n281) );
  NAND U508 ( .A(n282), .B(n283), .Z(n247) );
  OR U509 ( .A(n284), .B(n285), .Z(n283) );
  OR U510 ( .A(n286), .B(n287), .Z(n282) );
  NAND U511 ( .A(n288), .B(n289), .Z(n245) );
  OR U512 ( .A(n290), .B(n291), .Z(n289) );
  OR U513 ( .A(n292), .B(n293), .Z(n288) );
  ANDN U514 ( .B(n294), .A(n295), .Z(n246) );
  IV U515 ( .A(n296), .Z(n294) );
  ANDN U516 ( .B(n297), .A(n298), .Z(n238) );
  XOR U517 ( .A(n224), .B(n299), .Z(n236) );
  XOR U518 ( .A(n225), .B(n226), .Z(n299) );
  XOR U519 ( .A(n231), .B(n300), .Z(n226) );
  XOR U520 ( .A(n230), .B(n233), .Z(n300) );
  IV U521 ( .A(n232), .Z(n233) );
  NAND U522 ( .A(n301), .B(n302), .Z(n232) );
  OR U523 ( .A(n303), .B(n304), .Z(n302) );
  OR U524 ( .A(n305), .B(n306), .Z(n301) );
  NAND U525 ( .A(n307), .B(n308), .Z(n230) );
  OR U526 ( .A(n309), .B(n310), .Z(n308) );
  OR U527 ( .A(n311), .B(n312), .Z(n307) );
  NOR U528 ( .A(n313), .B(n314), .Z(n231) );
  ANDN U529 ( .B(n315), .A(n316), .Z(n225) );
  IV U530 ( .A(n317), .Z(n315) );
  XNOR U531 ( .A(n218), .B(n318), .Z(n224) );
  XNOR U532 ( .A(n217), .B(n219), .Z(n318) );
  NAND U533 ( .A(n319), .B(n320), .Z(n219) );
  OR U534 ( .A(n321), .B(n322), .Z(n320) );
  OR U535 ( .A(n323), .B(n324), .Z(n319) );
  NAND U536 ( .A(n325), .B(n326), .Z(n217) );
  OR U537 ( .A(n327), .B(n328), .Z(n326) );
  OR U538 ( .A(n329), .B(n330), .Z(n325) );
  ANDN U539 ( .B(n331), .A(n332), .Z(n218) );
  IV U540 ( .A(n333), .Z(n331) );
  XNOR U541 ( .A(n298), .B(n297), .Z(N1211) );
  XOR U542 ( .A(n317), .B(n316), .Z(n297) );
  XNOR U543 ( .A(n332), .B(n333), .Z(n316) );
  XNOR U544 ( .A(n327), .B(n328), .Z(n333) );
  XNOR U545 ( .A(n329), .B(n330), .Z(n328) );
  XNOR U546 ( .A(y[232]), .B(x[232]), .Z(n330) );
  XNOR U547 ( .A(y[233]), .B(x[233]), .Z(n329) );
  XNOR U548 ( .A(y[231]), .B(x[231]), .Z(n327) );
  XNOR U549 ( .A(n321), .B(n322), .Z(n332) );
  XNOR U550 ( .A(y[228]), .B(x[228]), .Z(n322) );
  XNOR U551 ( .A(n323), .B(n324), .Z(n321) );
  XNOR U552 ( .A(y[229]), .B(x[229]), .Z(n324) );
  XNOR U553 ( .A(y[230]), .B(x[230]), .Z(n323) );
  XNOR U554 ( .A(n314), .B(n313), .Z(n317) );
  XNOR U555 ( .A(n309), .B(n310), .Z(n313) );
  XNOR U556 ( .A(y[225]), .B(x[225]), .Z(n310) );
  XNOR U557 ( .A(n311), .B(n312), .Z(n309) );
  XNOR U558 ( .A(y[226]), .B(x[226]), .Z(n312) );
  XNOR U559 ( .A(y[227]), .B(x[227]), .Z(n311) );
  XNOR U560 ( .A(n303), .B(n304), .Z(n314) );
  XNOR U561 ( .A(y[222]), .B(x[222]), .Z(n304) );
  XNOR U562 ( .A(n305), .B(n306), .Z(n303) );
  XNOR U563 ( .A(y[223]), .B(x[223]), .Z(n306) );
  XNOR U564 ( .A(y[224]), .B(x[224]), .Z(n305) );
  XOR U565 ( .A(n279), .B(n280), .Z(n298) );
  XNOR U566 ( .A(n295), .B(n296), .Z(n280) );
  XNOR U567 ( .A(n290), .B(n291), .Z(n296) );
  XNOR U568 ( .A(n292), .B(n293), .Z(n291) );
  XNOR U569 ( .A(y[220]), .B(x[220]), .Z(n293) );
  XNOR U570 ( .A(y[221]), .B(x[221]), .Z(n292) );
  XNOR U571 ( .A(y[219]), .B(x[219]), .Z(n290) );
  XNOR U572 ( .A(n284), .B(n285), .Z(n295) );
  XNOR U573 ( .A(y[216]), .B(x[216]), .Z(n285) );
  XNOR U574 ( .A(n286), .B(n287), .Z(n284) );
  XNOR U575 ( .A(y[217]), .B(x[217]), .Z(n287) );
  XNOR U576 ( .A(y[218]), .B(x[218]), .Z(n286) );
  XOR U577 ( .A(n278), .B(n277), .Z(n279) );
  XNOR U578 ( .A(n273), .B(n274), .Z(n277) );
  XNOR U579 ( .A(y[213]), .B(x[213]), .Z(n274) );
  XNOR U580 ( .A(n275), .B(n276), .Z(n273) );
  XNOR U581 ( .A(y[214]), .B(x[214]), .Z(n276) );
  XNOR U582 ( .A(y[215]), .B(x[215]), .Z(n275) );
  XNOR U583 ( .A(n267), .B(n268), .Z(n278) );
  XNOR U584 ( .A(y[210]), .B(x[210]), .Z(n268) );
  XNOR U585 ( .A(n269), .B(n270), .Z(n267) );
  XNOR U586 ( .A(y[211]), .B(x[211]), .Z(n270) );
  XNOR U587 ( .A(y[212]), .B(x[212]), .Z(n269) );
  NAND U588 ( .A(n334), .B(n335), .Z(N1207) );
  NANDN U589 ( .A(n336), .B(n337), .Z(n335) );
  OR U590 ( .A(n338), .B(n339), .Z(n337) );
  NAND U591 ( .A(n338), .B(n339), .Z(n334) );
  XOR U592 ( .A(n338), .B(n340), .Z(N1206) );
  XNOR U593 ( .A(n336), .B(n339), .Z(n340) );
  AND U594 ( .A(n341), .B(n342), .Z(n339) );
  NANDN U595 ( .A(n343), .B(n344), .Z(n342) );
  NANDN U596 ( .A(n345), .B(n346), .Z(n344) );
  NANDN U597 ( .A(n346), .B(n345), .Z(n341) );
  NAND U598 ( .A(n347), .B(n348), .Z(n336) );
  NANDN U599 ( .A(n349), .B(n350), .Z(n348) );
  OR U600 ( .A(n351), .B(n352), .Z(n350) );
  NAND U601 ( .A(n352), .B(n351), .Z(n347) );
  AND U602 ( .A(n353), .B(n354), .Z(n338) );
  NANDN U603 ( .A(n355), .B(n356), .Z(n354) );
  NANDN U604 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U605 ( .A(n358), .B(n357), .Z(n353) );
  XOR U606 ( .A(n352), .B(n359), .Z(N1205) );
  XOR U607 ( .A(n349), .B(n351), .Z(n359) );
  XNOR U608 ( .A(n345), .B(n360), .Z(n351) );
  XNOR U609 ( .A(n343), .B(n346), .Z(n360) );
  NAND U610 ( .A(n361), .B(n362), .Z(n346) );
  NAND U611 ( .A(n363), .B(n364), .Z(n362) );
  OR U612 ( .A(n365), .B(n366), .Z(n363) );
  NANDN U613 ( .A(n367), .B(n365), .Z(n361) );
  IV U614 ( .A(n366), .Z(n367) );
  NAND U615 ( .A(n368), .B(n369), .Z(n343) );
  NAND U616 ( .A(n370), .B(n371), .Z(n369) );
  NANDN U617 ( .A(n372), .B(n373), .Z(n370) );
  NANDN U618 ( .A(n373), .B(n372), .Z(n368) );
  AND U619 ( .A(n374), .B(n375), .Z(n345) );
  NAND U620 ( .A(n376), .B(n377), .Z(n375) );
  OR U621 ( .A(n378), .B(n379), .Z(n376) );
  NANDN U622 ( .A(n380), .B(n378), .Z(n374) );
  NAND U623 ( .A(n381), .B(n382), .Z(n349) );
  NANDN U624 ( .A(n383), .B(n384), .Z(n382) );
  OR U625 ( .A(n385), .B(n386), .Z(n384) );
  NANDN U626 ( .A(n387), .B(n385), .Z(n381) );
  IV U627 ( .A(n386), .Z(n387) );
  XNOR U628 ( .A(n357), .B(n388), .Z(n352) );
  XNOR U629 ( .A(n355), .B(n358), .Z(n388) );
  NAND U630 ( .A(n389), .B(n390), .Z(n358) );
  NAND U631 ( .A(n391), .B(n392), .Z(n390) );
  OR U632 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U633 ( .A(n395), .B(n393), .Z(n389) );
  IV U634 ( .A(n394), .Z(n395) );
  NAND U635 ( .A(n396), .B(n397), .Z(n355) );
  NAND U636 ( .A(n398), .B(n399), .Z(n397) );
  NANDN U637 ( .A(n400), .B(n401), .Z(n398) );
  NANDN U638 ( .A(n401), .B(n400), .Z(n396) );
  AND U639 ( .A(n402), .B(n403), .Z(n357) );
  NAND U640 ( .A(n404), .B(n405), .Z(n403) );
  OR U641 ( .A(n406), .B(n407), .Z(n404) );
  NANDN U642 ( .A(n408), .B(n406), .Z(n402) );
  XNOR U643 ( .A(n383), .B(n409), .Z(N1204) );
  XOR U644 ( .A(n385), .B(n386), .Z(n409) );
  XNOR U645 ( .A(n399), .B(n410), .Z(n386) );
  XOR U646 ( .A(n400), .B(n401), .Z(n410) );
  XOR U647 ( .A(n406), .B(n411), .Z(n401) );
  XOR U648 ( .A(n405), .B(n408), .Z(n411) );
  IV U649 ( .A(n407), .Z(n408) );
  NAND U650 ( .A(n412), .B(n413), .Z(n407) );
  OR U651 ( .A(n414), .B(n415), .Z(n413) );
  OR U652 ( .A(n416), .B(n417), .Z(n412) );
  NAND U653 ( .A(n418), .B(n419), .Z(n405) );
  OR U654 ( .A(n420), .B(n421), .Z(n419) );
  OR U655 ( .A(n422), .B(n423), .Z(n418) );
  NOR U656 ( .A(n424), .B(n425), .Z(n406) );
  ANDN U657 ( .B(n426), .A(n427), .Z(n400) );
  XNOR U658 ( .A(n393), .B(n428), .Z(n399) );
  XNOR U659 ( .A(n392), .B(n394), .Z(n428) );
  NAND U660 ( .A(n429), .B(n430), .Z(n394) );
  OR U661 ( .A(n431), .B(n432), .Z(n430) );
  OR U662 ( .A(n433), .B(n434), .Z(n429) );
  NAND U663 ( .A(n435), .B(n436), .Z(n392) );
  OR U664 ( .A(n437), .B(n438), .Z(n436) );
  OR U665 ( .A(n439), .B(n440), .Z(n435) );
  ANDN U666 ( .B(n441), .A(n442), .Z(n393) );
  IV U667 ( .A(n443), .Z(n441) );
  ANDN U668 ( .B(n444), .A(n445), .Z(n385) );
  XOR U669 ( .A(n371), .B(n446), .Z(n383) );
  XOR U670 ( .A(n372), .B(n373), .Z(n446) );
  XOR U671 ( .A(n378), .B(n447), .Z(n373) );
  XOR U672 ( .A(n377), .B(n380), .Z(n447) );
  IV U673 ( .A(n379), .Z(n380) );
  NAND U674 ( .A(n448), .B(n449), .Z(n379) );
  OR U675 ( .A(n450), .B(n451), .Z(n449) );
  OR U676 ( .A(n452), .B(n453), .Z(n448) );
  NAND U677 ( .A(n454), .B(n455), .Z(n377) );
  OR U678 ( .A(n456), .B(n457), .Z(n455) );
  OR U679 ( .A(n458), .B(n459), .Z(n454) );
  NOR U680 ( .A(n460), .B(n461), .Z(n378) );
  ANDN U681 ( .B(n462), .A(n463), .Z(n372) );
  IV U682 ( .A(n464), .Z(n462) );
  XNOR U683 ( .A(n365), .B(n465), .Z(n371) );
  XNOR U684 ( .A(n364), .B(n366), .Z(n465) );
  NAND U685 ( .A(n466), .B(n467), .Z(n366) );
  OR U686 ( .A(n468), .B(n469), .Z(n467) );
  OR U687 ( .A(n470), .B(n471), .Z(n466) );
  NAND U688 ( .A(n472), .B(n473), .Z(n364) );
  OR U689 ( .A(n474), .B(n475), .Z(n473) );
  OR U690 ( .A(n476), .B(n477), .Z(n472) );
  ANDN U691 ( .B(n478), .A(n479), .Z(n365) );
  IV U692 ( .A(n480), .Z(n478) );
  XNOR U693 ( .A(n445), .B(n444), .Z(N1203) );
  XOR U694 ( .A(n464), .B(n463), .Z(n444) );
  XNOR U695 ( .A(n479), .B(n480), .Z(n463) );
  XNOR U696 ( .A(n474), .B(n475), .Z(n480) );
  XNOR U697 ( .A(n476), .B(n477), .Z(n475) );
  XNOR U698 ( .A(y[208]), .B(x[208]), .Z(n477) );
  XNOR U699 ( .A(y[209]), .B(x[209]), .Z(n476) );
  XNOR U700 ( .A(y[207]), .B(x[207]), .Z(n474) );
  XNOR U701 ( .A(n468), .B(n469), .Z(n479) );
  XNOR U702 ( .A(y[204]), .B(x[204]), .Z(n469) );
  XNOR U703 ( .A(n470), .B(n471), .Z(n468) );
  XNOR U704 ( .A(y[205]), .B(x[205]), .Z(n471) );
  XNOR U705 ( .A(y[206]), .B(x[206]), .Z(n470) );
  XNOR U706 ( .A(n461), .B(n460), .Z(n464) );
  XNOR U707 ( .A(n456), .B(n457), .Z(n460) );
  XNOR U708 ( .A(y[201]), .B(x[201]), .Z(n457) );
  XNOR U709 ( .A(n458), .B(n459), .Z(n456) );
  XNOR U710 ( .A(y[202]), .B(x[202]), .Z(n459) );
  XNOR U711 ( .A(y[203]), .B(x[203]), .Z(n458) );
  XNOR U712 ( .A(n450), .B(n451), .Z(n461) );
  XNOR U713 ( .A(y[198]), .B(x[198]), .Z(n451) );
  XNOR U714 ( .A(n452), .B(n453), .Z(n450) );
  XNOR U715 ( .A(y[199]), .B(x[199]), .Z(n453) );
  XNOR U716 ( .A(y[200]), .B(x[200]), .Z(n452) );
  XOR U717 ( .A(n426), .B(n427), .Z(n445) );
  XNOR U718 ( .A(n442), .B(n443), .Z(n427) );
  XNOR U719 ( .A(n437), .B(n438), .Z(n443) );
  XNOR U720 ( .A(n439), .B(n440), .Z(n438) );
  XNOR U721 ( .A(y[196]), .B(x[196]), .Z(n440) );
  XNOR U722 ( .A(y[197]), .B(x[197]), .Z(n439) );
  XNOR U723 ( .A(y[195]), .B(x[195]), .Z(n437) );
  XNOR U724 ( .A(n431), .B(n432), .Z(n442) );
  XNOR U725 ( .A(y[192]), .B(x[192]), .Z(n432) );
  XNOR U726 ( .A(n433), .B(n434), .Z(n431) );
  XNOR U727 ( .A(y[193]), .B(x[193]), .Z(n434) );
  XNOR U728 ( .A(y[194]), .B(x[194]), .Z(n433) );
  XOR U729 ( .A(n425), .B(n424), .Z(n426) );
  XNOR U730 ( .A(n420), .B(n421), .Z(n424) );
  XNOR U731 ( .A(y[189]), .B(x[189]), .Z(n421) );
  XNOR U732 ( .A(n422), .B(n423), .Z(n420) );
  XNOR U733 ( .A(y[190]), .B(x[190]), .Z(n423) );
  XNOR U734 ( .A(y[191]), .B(x[191]), .Z(n422) );
  XNOR U735 ( .A(n414), .B(n415), .Z(n425) );
  XNOR U736 ( .A(y[186]), .B(x[186]), .Z(n415) );
  XNOR U737 ( .A(n416), .B(n417), .Z(n414) );
  XNOR U738 ( .A(y[187]), .B(x[187]), .Z(n417) );
  XNOR U739 ( .A(y[188]), .B(x[188]), .Z(n416) );
  NAND U740 ( .A(n481), .B(n482), .Z(N1199) );
  NANDN U741 ( .A(n483), .B(n484), .Z(n482) );
  OR U742 ( .A(n485), .B(n486), .Z(n484) );
  NAND U743 ( .A(n485), .B(n486), .Z(n481) );
  XOR U744 ( .A(n485), .B(n487), .Z(N1198) );
  XNOR U745 ( .A(n483), .B(n486), .Z(n487) );
  AND U746 ( .A(n488), .B(n489), .Z(n486) );
  NANDN U747 ( .A(n490), .B(n491), .Z(n489) );
  NANDN U748 ( .A(n492), .B(n493), .Z(n491) );
  NANDN U749 ( .A(n493), .B(n492), .Z(n488) );
  NAND U750 ( .A(n494), .B(n495), .Z(n483) );
  NANDN U751 ( .A(n496), .B(n497), .Z(n495) );
  OR U752 ( .A(n498), .B(n499), .Z(n497) );
  NAND U753 ( .A(n499), .B(n498), .Z(n494) );
  AND U754 ( .A(n500), .B(n501), .Z(n485) );
  NANDN U755 ( .A(n502), .B(n503), .Z(n501) );
  NANDN U756 ( .A(n504), .B(n505), .Z(n503) );
  NANDN U757 ( .A(n505), .B(n504), .Z(n500) );
  XOR U758 ( .A(n499), .B(n506), .Z(N1197) );
  XOR U759 ( .A(n496), .B(n498), .Z(n506) );
  XNOR U760 ( .A(n492), .B(n507), .Z(n498) );
  XNOR U761 ( .A(n490), .B(n493), .Z(n507) );
  NAND U762 ( .A(n508), .B(n509), .Z(n493) );
  NAND U763 ( .A(n510), .B(n511), .Z(n509) );
  OR U764 ( .A(n512), .B(n513), .Z(n510) );
  NANDN U765 ( .A(n514), .B(n512), .Z(n508) );
  IV U766 ( .A(n513), .Z(n514) );
  NAND U767 ( .A(n515), .B(n516), .Z(n490) );
  NAND U768 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U769 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U770 ( .A(n520), .B(n519), .Z(n515) );
  AND U771 ( .A(n521), .B(n522), .Z(n492) );
  NAND U772 ( .A(n523), .B(n524), .Z(n522) );
  OR U773 ( .A(n525), .B(n526), .Z(n523) );
  NANDN U774 ( .A(n527), .B(n525), .Z(n521) );
  NAND U775 ( .A(n528), .B(n529), .Z(n496) );
  NANDN U776 ( .A(n530), .B(n531), .Z(n529) );
  OR U777 ( .A(n532), .B(n533), .Z(n531) );
  NANDN U778 ( .A(n534), .B(n532), .Z(n528) );
  IV U779 ( .A(n533), .Z(n534) );
  XNOR U780 ( .A(n504), .B(n535), .Z(n499) );
  XNOR U781 ( .A(n502), .B(n505), .Z(n535) );
  NAND U782 ( .A(n536), .B(n537), .Z(n505) );
  NAND U783 ( .A(n538), .B(n539), .Z(n537) );
  OR U784 ( .A(n540), .B(n541), .Z(n538) );
  NANDN U785 ( .A(n542), .B(n540), .Z(n536) );
  IV U786 ( .A(n541), .Z(n542) );
  NAND U787 ( .A(n543), .B(n544), .Z(n502) );
  NAND U788 ( .A(n545), .B(n546), .Z(n544) );
  NANDN U789 ( .A(n547), .B(n548), .Z(n545) );
  NANDN U790 ( .A(n548), .B(n547), .Z(n543) );
  AND U791 ( .A(n549), .B(n550), .Z(n504) );
  NAND U792 ( .A(n551), .B(n552), .Z(n550) );
  OR U793 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U794 ( .A(n555), .B(n553), .Z(n549) );
  XNOR U795 ( .A(n530), .B(n556), .Z(N1196) );
  XOR U796 ( .A(n532), .B(n533), .Z(n556) );
  XNOR U797 ( .A(n546), .B(n557), .Z(n533) );
  XOR U798 ( .A(n547), .B(n548), .Z(n557) );
  XOR U799 ( .A(n553), .B(n558), .Z(n548) );
  XOR U800 ( .A(n552), .B(n555), .Z(n558) );
  IV U801 ( .A(n554), .Z(n555) );
  NAND U802 ( .A(n559), .B(n560), .Z(n554) );
  OR U803 ( .A(n561), .B(n562), .Z(n560) );
  OR U804 ( .A(n563), .B(n564), .Z(n559) );
  NAND U805 ( .A(n565), .B(n566), .Z(n552) );
  OR U806 ( .A(n567), .B(n568), .Z(n566) );
  OR U807 ( .A(n569), .B(n570), .Z(n565) );
  NOR U808 ( .A(n571), .B(n572), .Z(n553) );
  ANDN U809 ( .B(n573), .A(n574), .Z(n547) );
  XNOR U810 ( .A(n540), .B(n575), .Z(n546) );
  XNOR U811 ( .A(n539), .B(n541), .Z(n575) );
  NAND U812 ( .A(n576), .B(n577), .Z(n541) );
  OR U813 ( .A(n578), .B(n579), .Z(n577) );
  OR U814 ( .A(n580), .B(n581), .Z(n576) );
  NAND U815 ( .A(n582), .B(n583), .Z(n539) );
  OR U816 ( .A(n584), .B(n585), .Z(n583) );
  OR U817 ( .A(n586), .B(n587), .Z(n582) );
  ANDN U818 ( .B(n588), .A(n589), .Z(n540) );
  IV U819 ( .A(n590), .Z(n588) );
  ANDN U820 ( .B(n591), .A(n592), .Z(n532) );
  XOR U821 ( .A(n518), .B(n593), .Z(n530) );
  XOR U822 ( .A(n519), .B(n520), .Z(n593) );
  XOR U823 ( .A(n525), .B(n594), .Z(n520) );
  XOR U824 ( .A(n524), .B(n527), .Z(n594) );
  IV U825 ( .A(n526), .Z(n527) );
  NAND U826 ( .A(n595), .B(n596), .Z(n526) );
  OR U827 ( .A(n597), .B(n598), .Z(n596) );
  OR U828 ( .A(n599), .B(n600), .Z(n595) );
  NAND U829 ( .A(n601), .B(n602), .Z(n524) );
  OR U830 ( .A(n603), .B(n604), .Z(n602) );
  OR U831 ( .A(n605), .B(n606), .Z(n601) );
  NOR U832 ( .A(n607), .B(n608), .Z(n525) );
  ANDN U833 ( .B(n609), .A(n610), .Z(n519) );
  IV U834 ( .A(n611), .Z(n609) );
  XNOR U835 ( .A(n512), .B(n612), .Z(n518) );
  XNOR U836 ( .A(n511), .B(n513), .Z(n612) );
  NAND U837 ( .A(n613), .B(n614), .Z(n513) );
  OR U838 ( .A(n615), .B(n616), .Z(n614) );
  OR U839 ( .A(n617), .B(n618), .Z(n613) );
  NAND U840 ( .A(n619), .B(n620), .Z(n511) );
  OR U841 ( .A(n621), .B(n622), .Z(n620) );
  OR U842 ( .A(n623), .B(n624), .Z(n619) );
  ANDN U843 ( .B(n625), .A(n626), .Z(n512) );
  IV U844 ( .A(n627), .Z(n625) );
  XNOR U845 ( .A(n592), .B(n591), .Z(N1195) );
  XOR U846 ( .A(n611), .B(n610), .Z(n591) );
  XNOR U847 ( .A(n626), .B(n627), .Z(n610) );
  XNOR U848 ( .A(n621), .B(n622), .Z(n627) );
  XNOR U849 ( .A(n623), .B(n624), .Z(n622) );
  XNOR U850 ( .A(y[184]), .B(x[184]), .Z(n624) );
  XNOR U851 ( .A(y[185]), .B(x[185]), .Z(n623) );
  XNOR U852 ( .A(y[183]), .B(x[183]), .Z(n621) );
  XNOR U853 ( .A(n615), .B(n616), .Z(n626) );
  XNOR U854 ( .A(y[180]), .B(x[180]), .Z(n616) );
  XNOR U855 ( .A(n617), .B(n618), .Z(n615) );
  XNOR U856 ( .A(y[181]), .B(x[181]), .Z(n618) );
  XNOR U857 ( .A(y[182]), .B(x[182]), .Z(n617) );
  XNOR U858 ( .A(n608), .B(n607), .Z(n611) );
  XNOR U859 ( .A(n603), .B(n604), .Z(n607) );
  XNOR U860 ( .A(y[177]), .B(x[177]), .Z(n604) );
  XNOR U861 ( .A(n605), .B(n606), .Z(n603) );
  XNOR U862 ( .A(y[178]), .B(x[178]), .Z(n606) );
  XNOR U863 ( .A(y[179]), .B(x[179]), .Z(n605) );
  XNOR U864 ( .A(n597), .B(n598), .Z(n608) );
  XNOR U865 ( .A(y[174]), .B(x[174]), .Z(n598) );
  XNOR U866 ( .A(n599), .B(n600), .Z(n597) );
  XNOR U867 ( .A(y[175]), .B(x[175]), .Z(n600) );
  XNOR U868 ( .A(y[176]), .B(x[176]), .Z(n599) );
  XOR U869 ( .A(n573), .B(n574), .Z(n592) );
  XNOR U870 ( .A(n589), .B(n590), .Z(n574) );
  XNOR U871 ( .A(n584), .B(n585), .Z(n590) );
  XNOR U872 ( .A(n586), .B(n587), .Z(n585) );
  XNOR U873 ( .A(y[172]), .B(x[172]), .Z(n587) );
  XNOR U874 ( .A(y[173]), .B(x[173]), .Z(n586) );
  XNOR U875 ( .A(y[171]), .B(x[171]), .Z(n584) );
  XNOR U876 ( .A(n578), .B(n579), .Z(n589) );
  XNOR U877 ( .A(y[168]), .B(x[168]), .Z(n579) );
  XNOR U878 ( .A(n580), .B(n581), .Z(n578) );
  XNOR U879 ( .A(y[169]), .B(x[169]), .Z(n581) );
  XNOR U880 ( .A(y[170]), .B(x[170]), .Z(n580) );
  XOR U881 ( .A(n572), .B(n571), .Z(n573) );
  XNOR U882 ( .A(n567), .B(n568), .Z(n571) );
  XNOR U883 ( .A(y[165]), .B(x[165]), .Z(n568) );
  XNOR U884 ( .A(n569), .B(n570), .Z(n567) );
  XNOR U885 ( .A(y[166]), .B(x[166]), .Z(n570) );
  XNOR U886 ( .A(y[167]), .B(x[167]), .Z(n569) );
  XNOR U887 ( .A(n561), .B(n562), .Z(n572) );
  XNOR U888 ( .A(y[162]), .B(x[162]), .Z(n562) );
  XNOR U889 ( .A(n563), .B(n564), .Z(n561) );
  XNOR U890 ( .A(y[163]), .B(x[163]), .Z(n564) );
  XNOR U891 ( .A(y[164]), .B(x[164]), .Z(n563) );
  NAND U892 ( .A(n628), .B(n629), .Z(N1191) );
  NANDN U893 ( .A(n630), .B(n631), .Z(n629) );
  OR U894 ( .A(n632), .B(n633), .Z(n631) );
  NAND U895 ( .A(n632), .B(n633), .Z(n628) );
  XOR U896 ( .A(n632), .B(n634), .Z(N1190) );
  XNOR U897 ( .A(n630), .B(n633), .Z(n634) );
  AND U898 ( .A(n635), .B(n636), .Z(n633) );
  NANDN U899 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U900 ( .A(n639), .B(n640), .Z(n638) );
  NANDN U901 ( .A(n640), .B(n639), .Z(n635) );
  NAND U902 ( .A(n641), .B(n642), .Z(n630) );
  NANDN U903 ( .A(n643), .B(n644), .Z(n642) );
  OR U904 ( .A(n645), .B(n646), .Z(n644) );
  NAND U905 ( .A(n646), .B(n645), .Z(n641) );
  AND U906 ( .A(n647), .B(n648), .Z(n632) );
  NANDN U907 ( .A(n649), .B(n650), .Z(n648) );
  NANDN U908 ( .A(n651), .B(n652), .Z(n650) );
  NANDN U909 ( .A(n652), .B(n651), .Z(n647) );
  XOR U910 ( .A(n646), .B(n653), .Z(N1189) );
  XOR U911 ( .A(n643), .B(n645), .Z(n653) );
  XNOR U912 ( .A(n639), .B(n654), .Z(n645) );
  XNOR U913 ( .A(n637), .B(n640), .Z(n654) );
  NAND U914 ( .A(n655), .B(n656), .Z(n640) );
  NAND U915 ( .A(n657), .B(n658), .Z(n656) );
  OR U916 ( .A(n659), .B(n660), .Z(n657) );
  NANDN U917 ( .A(n661), .B(n659), .Z(n655) );
  IV U918 ( .A(n660), .Z(n661) );
  NAND U919 ( .A(n662), .B(n663), .Z(n637) );
  NAND U920 ( .A(n664), .B(n665), .Z(n663) );
  NANDN U921 ( .A(n666), .B(n667), .Z(n664) );
  NANDN U922 ( .A(n667), .B(n666), .Z(n662) );
  AND U923 ( .A(n668), .B(n669), .Z(n639) );
  NAND U924 ( .A(n670), .B(n671), .Z(n669) );
  OR U925 ( .A(n672), .B(n673), .Z(n670) );
  NANDN U926 ( .A(n674), .B(n672), .Z(n668) );
  NAND U927 ( .A(n675), .B(n676), .Z(n643) );
  NANDN U928 ( .A(n677), .B(n678), .Z(n676) );
  OR U929 ( .A(n679), .B(n680), .Z(n678) );
  NANDN U930 ( .A(n681), .B(n679), .Z(n675) );
  IV U931 ( .A(n680), .Z(n681) );
  XNOR U932 ( .A(n651), .B(n682), .Z(n646) );
  XNOR U933 ( .A(n649), .B(n652), .Z(n682) );
  NAND U934 ( .A(n683), .B(n684), .Z(n652) );
  NAND U935 ( .A(n685), .B(n686), .Z(n684) );
  OR U936 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U937 ( .A(n689), .B(n687), .Z(n683) );
  IV U938 ( .A(n688), .Z(n689) );
  NAND U939 ( .A(n690), .B(n691), .Z(n649) );
  NAND U940 ( .A(n692), .B(n693), .Z(n691) );
  NANDN U941 ( .A(n694), .B(n695), .Z(n692) );
  NANDN U942 ( .A(n695), .B(n694), .Z(n690) );
  AND U943 ( .A(n696), .B(n697), .Z(n651) );
  NAND U944 ( .A(n698), .B(n699), .Z(n697) );
  OR U945 ( .A(n700), .B(n701), .Z(n698) );
  NANDN U946 ( .A(n702), .B(n700), .Z(n696) );
  XNOR U947 ( .A(n677), .B(n703), .Z(N1188) );
  XOR U948 ( .A(n679), .B(n680), .Z(n703) );
  XNOR U949 ( .A(n693), .B(n704), .Z(n680) );
  XOR U950 ( .A(n694), .B(n695), .Z(n704) );
  XOR U951 ( .A(n700), .B(n705), .Z(n695) );
  XOR U952 ( .A(n699), .B(n702), .Z(n705) );
  IV U953 ( .A(n701), .Z(n702) );
  NAND U954 ( .A(n706), .B(n707), .Z(n701) );
  OR U955 ( .A(n708), .B(n709), .Z(n707) );
  OR U956 ( .A(n710), .B(n711), .Z(n706) );
  NAND U957 ( .A(n712), .B(n713), .Z(n699) );
  OR U958 ( .A(n714), .B(n715), .Z(n713) );
  OR U959 ( .A(n716), .B(n717), .Z(n712) );
  NOR U960 ( .A(n718), .B(n719), .Z(n700) );
  ANDN U961 ( .B(n720), .A(n721), .Z(n694) );
  XNOR U962 ( .A(n687), .B(n722), .Z(n693) );
  XNOR U963 ( .A(n686), .B(n688), .Z(n722) );
  NAND U964 ( .A(n723), .B(n724), .Z(n688) );
  OR U965 ( .A(n725), .B(n726), .Z(n724) );
  OR U966 ( .A(n727), .B(n728), .Z(n723) );
  NAND U967 ( .A(n729), .B(n730), .Z(n686) );
  OR U968 ( .A(n731), .B(n732), .Z(n730) );
  OR U969 ( .A(n733), .B(n734), .Z(n729) );
  ANDN U970 ( .B(n735), .A(n736), .Z(n687) );
  IV U971 ( .A(n737), .Z(n735) );
  ANDN U972 ( .B(n738), .A(n739), .Z(n679) );
  XOR U973 ( .A(n665), .B(n740), .Z(n677) );
  XOR U974 ( .A(n666), .B(n667), .Z(n740) );
  XOR U975 ( .A(n672), .B(n741), .Z(n667) );
  XOR U976 ( .A(n671), .B(n674), .Z(n741) );
  IV U977 ( .A(n673), .Z(n674) );
  NAND U978 ( .A(n742), .B(n743), .Z(n673) );
  OR U979 ( .A(n744), .B(n745), .Z(n743) );
  OR U980 ( .A(n746), .B(n747), .Z(n742) );
  NAND U981 ( .A(n748), .B(n749), .Z(n671) );
  OR U982 ( .A(n750), .B(n751), .Z(n749) );
  OR U983 ( .A(n752), .B(n753), .Z(n748) );
  NOR U984 ( .A(n754), .B(n755), .Z(n672) );
  ANDN U985 ( .B(n756), .A(n757), .Z(n666) );
  IV U986 ( .A(n758), .Z(n756) );
  XNOR U987 ( .A(n659), .B(n759), .Z(n665) );
  XNOR U988 ( .A(n658), .B(n660), .Z(n759) );
  NAND U989 ( .A(n760), .B(n761), .Z(n660) );
  OR U990 ( .A(n762), .B(n763), .Z(n761) );
  OR U991 ( .A(n764), .B(n765), .Z(n760) );
  NAND U992 ( .A(n766), .B(n767), .Z(n658) );
  OR U993 ( .A(n768), .B(n769), .Z(n767) );
  OR U994 ( .A(n770), .B(n771), .Z(n766) );
  ANDN U995 ( .B(n772), .A(n773), .Z(n659) );
  IV U996 ( .A(n774), .Z(n772) );
  XNOR U997 ( .A(n739), .B(n738), .Z(N1187) );
  XOR U998 ( .A(n758), .B(n757), .Z(n738) );
  XNOR U999 ( .A(n773), .B(n774), .Z(n757) );
  XNOR U1000 ( .A(n768), .B(n769), .Z(n774) );
  XNOR U1001 ( .A(n770), .B(n771), .Z(n769) );
  XNOR U1002 ( .A(y[160]), .B(x[160]), .Z(n771) );
  XNOR U1003 ( .A(y[161]), .B(x[161]), .Z(n770) );
  XNOR U1004 ( .A(y[159]), .B(x[159]), .Z(n768) );
  XNOR U1005 ( .A(n762), .B(n763), .Z(n773) );
  XNOR U1006 ( .A(y[156]), .B(x[156]), .Z(n763) );
  XNOR U1007 ( .A(n764), .B(n765), .Z(n762) );
  XNOR U1008 ( .A(y[157]), .B(x[157]), .Z(n765) );
  XNOR U1009 ( .A(y[158]), .B(x[158]), .Z(n764) );
  XNOR U1010 ( .A(n755), .B(n754), .Z(n758) );
  XNOR U1011 ( .A(n750), .B(n751), .Z(n754) );
  XNOR U1012 ( .A(y[153]), .B(x[153]), .Z(n751) );
  XNOR U1013 ( .A(n752), .B(n753), .Z(n750) );
  XNOR U1014 ( .A(y[154]), .B(x[154]), .Z(n753) );
  XNOR U1015 ( .A(y[155]), .B(x[155]), .Z(n752) );
  XNOR U1016 ( .A(n744), .B(n745), .Z(n755) );
  XNOR U1017 ( .A(y[150]), .B(x[150]), .Z(n745) );
  XNOR U1018 ( .A(n746), .B(n747), .Z(n744) );
  XNOR U1019 ( .A(y[151]), .B(x[151]), .Z(n747) );
  XNOR U1020 ( .A(y[152]), .B(x[152]), .Z(n746) );
  XOR U1021 ( .A(n720), .B(n721), .Z(n739) );
  XNOR U1022 ( .A(n736), .B(n737), .Z(n721) );
  XNOR U1023 ( .A(n731), .B(n732), .Z(n737) );
  XNOR U1024 ( .A(n733), .B(n734), .Z(n732) );
  XNOR U1025 ( .A(y[148]), .B(x[148]), .Z(n734) );
  XNOR U1026 ( .A(y[149]), .B(x[149]), .Z(n733) );
  XNOR U1027 ( .A(y[147]), .B(x[147]), .Z(n731) );
  XNOR U1028 ( .A(n725), .B(n726), .Z(n736) );
  XNOR U1029 ( .A(y[144]), .B(x[144]), .Z(n726) );
  XNOR U1030 ( .A(n727), .B(n728), .Z(n725) );
  XNOR U1031 ( .A(y[145]), .B(x[145]), .Z(n728) );
  XNOR U1032 ( .A(y[146]), .B(x[146]), .Z(n727) );
  XOR U1033 ( .A(n719), .B(n718), .Z(n720) );
  XNOR U1034 ( .A(n714), .B(n715), .Z(n718) );
  XNOR U1035 ( .A(y[141]), .B(x[141]), .Z(n715) );
  XNOR U1036 ( .A(n716), .B(n717), .Z(n714) );
  XNOR U1037 ( .A(y[142]), .B(x[142]), .Z(n717) );
  XNOR U1038 ( .A(y[143]), .B(x[143]), .Z(n716) );
  XNOR U1039 ( .A(n708), .B(n709), .Z(n719) );
  XNOR U1040 ( .A(y[138]), .B(x[138]), .Z(n709) );
  XNOR U1041 ( .A(n710), .B(n711), .Z(n708) );
  XNOR U1042 ( .A(y[139]), .B(x[139]), .Z(n711) );
  XNOR U1043 ( .A(y[140]), .B(x[140]), .Z(n710) );
  NAND U1044 ( .A(n775), .B(n776), .Z(N1183) );
  NANDN U1045 ( .A(n777), .B(n778), .Z(n776) );
  OR U1046 ( .A(n779), .B(n780), .Z(n778) );
  NAND U1047 ( .A(n779), .B(n780), .Z(n775) );
  XOR U1048 ( .A(n779), .B(n781), .Z(N1182) );
  XNOR U1049 ( .A(n777), .B(n780), .Z(n781) );
  AND U1050 ( .A(n782), .B(n783), .Z(n780) );
  NANDN U1051 ( .A(n784), .B(n785), .Z(n783) );
  NANDN U1052 ( .A(n786), .B(n787), .Z(n785) );
  NANDN U1053 ( .A(n787), .B(n786), .Z(n782) );
  NAND U1054 ( .A(n788), .B(n789), .Z(n777) );
  NANDN U1055 ( .A(n790), .B(n791), .Z(n789) );
  OR U1056 ( .A(n792), .B(n793), .Z(n791) );
  NAND U1057 ( .A(n793), .B(n792), .Z(n788) );
  AND U1058 ( .A(n794), .B(n795), .Z(n779) );
  NANDN U1059 ( .A(n796), .B(n797), .Z(n795) );
  NANDN U1060 ( .A(n798), .B(n799), .Z(n797) );
  NANDN U1061 ( .A(n799), .B(n798), .Z(n794) );
  XOR U1062 ( .A(n793), .B(n800), .Z(N1181) );
  XOR U1063 ( .A(n790), .B(n792), .Z(n800) );
  XNOR U1064 ( .A(n786), .B(n801), .Z(n792) );
  XNOR U1065 ( .A(n784), .B(n787), .Z(n801) );
  NAND U1066 ( .A(n802), .B(n803), .Z(n787) );
  NAND U1067 ( .A(n804), .B(n805), .Z(n803) );
  OR U1068 ( .A(n806), .B(n807), .Z(n804) );
  NANDN U1069 ( .A(n808), .B(n806), .Z(n802) );
  IV U1070 ( .A(n807), .Z(n808) );
  NAND U1071 ( .A(n809), .B(n810), .Z(n784) );
  NAND U1072 ( .A(n811), .B(n812), .Z(n810) );
  NANDN U1073 ( .A(n813), .B(n814), .Z(n811) );
  NANDN U1074 ( .A(n814), .B(n813), .Z(n809) );
  AND U1075 ( .A(n815), .B(n816), .Z(n786) );
  NAND U1076 ( .A(n817), .B(n818), .Z(n816) );
  OR U1077 ( .A(n819), .B(n820), .Z(n817) );
  NANDN U1078 ( .A(n821), .B(n819), .Z(n815) );
  NAND U1079 ( .A(n822), .B(n823), .Z(n790) );
  NANDN U1080 ( .A(n824), .B(n825), .Z(n823) );
  OR U1081 ( .A(n826), .B(n827), .Z(n825) );
  NANDN U1082 ( .A(n828), .B(n826), .Z(n822) );
  IV U1083 ( .A(n827), .Z(n828) );
  XNOR U1084 ( .A(n798), .B(n829), .Z(n793) );
  XNOR U1085 ( .A(n796), .B(n799), .Z(n829) );
  NAND U1086 ( .A(n830), .B(n831), .Z(n799) );
  NAND U1087 ( .A(n832), .B(n833), .Z(n831) );
  OR U1088 ( .A(n834), .B(n835), .Z(n832) );
  NANDN U1089 ( .A(n836), .B(n834), .Z(n830) );
  IV U1090 ( .A(n835), .Z(n836) );
  NAND U1091 ( .A(n837), .B(n838), .Z(n796) );
  NAND U1092 ( .A(n839), .B(n840), .Z(n838) );
  NANDN U1093 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U1094 ( .A(n842), .B(n841), .Z(n837) );
  AND U1095 ( .A(n843), .B(n844), .Z(n798) );
  NAND U1096 ( .A(n845), .B(n846), .Z(n844) );
  OR U1097 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U1098 ( .A(n849), .B(n847), .Z(n843) );
  XNOR U1099 ( .A(n824), .B(n850), .Z(N1180) );
  XOR U1100 ( .A(n826), .B(n827), .Z(n850) );
  XNOR U1101 ( .A(n840), .B(n851), .Z(n827) );
  XOR U1102 ( .A(n841), .B(n842), .Z(n851) );
  XOR U1103 ( .A(n847), .B(n852), .Z(n842) );
  XOR U1104 ( .A(n846), .B(n849), .Z(n852) );
  IV U1105 ( .A(n848), .Z(n849) );
  NAND U1106 ( .A(n853), .B(n854), .Z(n848) );
  OR U1107 ( .A(n855), .B(n856), .Z(n854) );
  OR U1108 ( .A(n857), .B(n858), .Z(n853) );
  NAND U1109 ( .A(n859), .B(n860), .Z(n846) );
  OR U1110 ( .A(n861), .B(n862), .Z(n860) );
  OR U1111 ( .A(n863), .B(n864), .Z(n859) );
  NOR U1112 ( .A(n865), .B(n866), .Z(n847) );
  ANDN U1113 ( .B(n867), .A(n868), .Z(n841) );
  XNOR U1114 ( .A(n834), .B(n869), .Z(n840) );
  XNOR U1115 ( .A(n833), .B(n835), .Z(n869) );
  NAND U1116 ( .A(n870), .B(n871), .Z(n835) );
  OR U1117 ( .A(n872), .B(n873), .Z(n871) );
  OR U1118 ( .A(n874), .B(n875), .Z(n870) );
  NAND U1119 ( .A(n876), .B(n877), .Z(n833) );
  OR U1120 ( .A(n878), .B(n879), .Z(n877) );
  OR U1121 ( .A(n880), .B(n881), .Z(n876) );
  ANDN U1122 ( .B(n882), .A(n883), .Z(n834) );
  IV U1123 ( .A(n884), .Z(n882) );
  ANDN U1124 ( .B(n885), .A(n886), .Z(n826) );
  XOR U1125 ( .A(n812), .B(n887), .Z(n824) );
  XOR U1126 ( .A(n813), .B(n814), .Z(n887) );
  XOR U1127 ( .A(n819), .B(n888), .Z(n814) );
  XOR U1128 ( .A(n818), .B(n821), .Z(n888) );
  IV U1129 ( .A(n820), .Z(n821) );
  NAND U1130 ( .A(n889), .B(n890), .Z(n820) );
  OR U1131 ( .A(n891), .B(n892), .Z(n890) );
  OR U1132 ( .A(n893), .B(n894), .Z(n889) );
  NAND U1133 ( .A(n895), .B(n896), .Z(n818) );
  OR U1134 ( .A(n897), .B(n898), .Z(n896) );
  OR U1135 ( .A(n899), .B(n900), .Z(n895) );
  NOR U1136 ( .A(n901), .B(n902), .Z(n819) );
  ANDN U1137 ( .B(n903), .A(n904), .Z(n813) );
  IV U1138 ( .A(n905), .Z(n903) );
  XNOR U1139 ( .A(n806), .B(n906), .Z(n812) );
  XNOR U1140 ( .A(n805), .B(n807), .Z(n906) );
  NAND U1141 ( .A(n907), .B(n908), .Z(n807) );
  OR U1142 ( .A(n909), .B(n910), .Z(n908) );
  OR U1143 ( .A(n911), .B(n912), .Z(n907) );
  NAND U1144 ( .A(n913), .B(n914), .Z(n805) );
  OR U1145 ( .A(n915), .B(n916), .Z(n914) );
  OR U1146 ( .A(n917), .B(n918), .Z(n913) );
  ANDN U1147 ( .B(n919), .A(n920), .Z(n806) );
  IV U1148 ( .A(n921), .Z(n919) );
  XNOR U1149 ( .A(n886), .B(n885), .Z(N1179) );
  XOR U1150 ( .A(n905), .B(n904), .Z(n885) );
  XNOR U1151 ( .A(n920), .B(n921), .Z(n904) );
  XNOR U1152 ( .A(n915), .B(n916), .Z(n921) );
  XNOR U1153 ( .A(n917), .B(n918), .Z(n916) );
  XNOR U1154 ( .A(y[136]), .B(x[136]), .Z(n918) );
  XNOR U1155 ( .A(y[137]), .B(x[137]), .Z(n917) );
  XNOR U1156 ( .A(y[135]), .B(x[135]), .Z(n915) );
  XNOR U1157 ( .A(n909), .B(n910), .Z(n920) );
  XNOR U1158 ( .A(y[132]), .B(x[132]), .Z(n910) );
  XNOR U1159 ( .A(n911), .B(n912), .Z(n909) );
  XNOR U1160 ( .A(y[133]), .B(x[133]), .Z(n912) );
  XNOR U1161 ( .A(y[134]), .B(x[134]), .Z(n911) );
  XNOR U1162 ( .A(n902), .B(n901), .Z(n905) );
  XNOR U1163 ( .A(n897), .B(n898), .Z(n901) );
  XNOR U1164 ( .A(y[129]), .B(x[129]), .Z(n898) );
  XNOR U1165 ( .A(n899), .B(n900), .Z(n897) );
  XNOR U1166 ( .A(y[130]), .B(x[130]), .Z(n900) );
  XNOR U1167 ( .A(y[131]), .B(x[131]), .Z(n899) );
  XNOR U1168 ( .A(n891), .B(n892), .Z(n902) );
  XNOR U1169 ( .A(y[126]), .B(x[126]), .Z(n892) );
  XNOR U1170 ( .A(n893), .B(n894), .Z(n891) );
  XNOR U1171 ( .A(y[127]), .B(x[127]), .Z(n894) );
  XNOR U1172 ( .A(y[128]), .B(x[128]), .Z(n893) );
  XOR U1173 ( .A(n867), .B(n868), .Z(n886) );
  XNOR U1174 ( .A(n883), .B(n884), .Z(n868) );
  XNOR U1175 ( .A(n878), .B(n879), .Z(n884) );
  XNOR U1176 ( .A(n880), .B(n881), .Z(n879) );
  XNOR U1177 ( .A(y[124]), .B(x[124]), .Z(n881) );
  XNOR U1178 ( .A(y[125]), .B(x[125]), .Z(n880) );
  XNOR U1179 ( .A(y[123]), .B(x[123]), .Z(n878) );
  XNOR U1180 ( .A(n872), .B(n873), .Z(n883) );
  XNOR U1181 ( .A(y[120]), .B(x[120]), .Z(n873) );
  XNOR U1182 ( .A(n874), .B(n875), .Z(n872) );
  XNOR U1183 ( .A(y[121]), .B(x[121]), .Z(n875) );
  XNOR U1184 ( .A(y[122]), .B(x[122]), .Z(n874) );
  XOR U1185 ( .A(n866), .B(n865), .Z(n867) );
  XNOR U1186 ( .A(n861), .B(n862), .Z(n865) );
  XNOR U1187 ( .A(y[117]), .B(x[117]), .Z(n862) );
  XNOR U1188 ( .A(n863), .B(n864), .Z(n861) );
  XNOR U1189 ( .A(y[118]), .B(x[118]), .Z(n864) );
  XNOR U1190 ( .A(y[119]), .B(x[119]), .Z(n863) );
  XNOR U1191 ( .A(n855), .B(n856), .Z(n866) );
  XNOR U1192 ( .A(y[114]), .B(x[114]), .Z(n856) );
  XNOR U1193 ( .A(n857), .B(n858), .Z(n855) );
  XNOR U1194 ( .A(y[115]), .B(x[115]), .Z(n858) );
  XNOR U1195 ( .A(y[116]), .B(x[116]), .Z(n857) );
  NAND U1196 ( .A(n922), .B(n923), .Z(N1175) );
  NANDN U1197 ( .A(n924), .B(n925), .Z(n923) );
  OR U1198 ( .A(n926), .B(n927), .Z(n925) );
  NAND U1199 ( .A(n926), .B(n927), .Z(n922) );
  XOR U1200 ( .A(n926), .B(n928), .Z(N1174) );
  XNOR U1201 ( .A(n924), .B(n927), .Z(n928) );
  AND U1202 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U1203 ( .A(n931), .B(n932), .Z(n930) );
  NANDN U1204 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U1205 ( .A(n934), .B(n933), .Z(n929) );
  NAND U1206 ( .A(n935), .B(n936), .Z(n924) );
  NANDN U1207 ( .A(n937), .B(n938), .Z(n936) );
  OR U1208 ( .A(n939), .B(n940), .Z(n938) );
  NAND U1209 ( .A(n940), .B(n939), .Z(n935) );
  AND U1210 ( .A(n941), .B(n942), .Z(n926) );
  NANDN U1211 ( .A(n943), .B(n944), .Z(n942) );
  NANDN U1212 ( .A(n945), .B(n946), .Z(n944) );
  NANDN U1213 ( .A(n946), .B(n945), .Z(n941) );
  XOR U1214 ( .A(n940), .B(n947), .Z(N1173) );
  XOR U1215 ( .A(n937), .B(n939), .Z(n947) );
  XNOR U1216 ( .A(n933), .B(n948), .Z(n939) );
  XNOR U1217 ( .A(n931), .B(n934), .Z(n948) );
  NAND U1218 ( .A(n949), .B(n950), .Z(n934) );
  NAND U1219 ( .A(n951), .B(n952), .Z(n950) );
  OR U1220 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U1221 ( .A(n955), .B(n953), .Z(n949) );
  IV U1222 ( .A(n954), .Z(n955) );
  NAND U1223 ( .A(n956), .B(n957), .Z(n931) );
  NAND U1224 ( .A(n958), .B(n959), .Z(n957) );
  NANDN U1225 ( .A(n960), .B(n961), .Z(n958) );
  NANDN U1226 ( .A(n961), .B(n960), .Z(n956) );
  AND U1227 ( .A(n962), .B(n963), .Z(n933) );
  NAND U1228 ( .A(n964), .B(n965), .Z(n963) );
  OR U1229 ( .A(n966), .B(n967), .Z(n964) );
  NANDN U1230 ( .A(n968), .B(n966), .Z(n962) );
  NAND U1231 ( .A(n969), .B(n970), .Z(n937) );
  NANDN U1232 ( .A(n971), .B(n972), .Z(n970) );
  OR U1233 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U1234 ( .A(n975), .B(n973), .Z(n969) );
  IV U1235 ( .A(n974), .Z(n975) );
  XNOR U1236 ( .A(n945), .B(n976), .Z(n940) );
  XNOR U1237 ( .A(n943), .B(n946), .Z(n976) );
  NAND U1238 ( .A(n977), .B(n978), .Z(n946) );
  NAND U1239 ( .A(n979), .B(n980), .Z(n978) );
  OR U1240 ( .A(n981), .B(n982), .Z(n979) );
  NANDN U1241 ( .A(n983), .B(n981), .Z(n977) );
  IV U1242 ( .A(n982), .Z(n983) );
  NAND U1243 ( .A(n984), .B(n985), .Z(n943) );
  NAND U1244 ( .A(n986), .B(n987), .Z(n985) );
  NANDN U1245 ( .A(n988), .B(n989), .Z(n986) );
  NANDN U1246 ( .A(n989), .B(n988), .Z(n984) );
  AND U1247 ( .A(n990), .B(n991), .Z(n945) );
  NAND U1248 ( .A(n992), .B(n993), .Z(n991) );
  OR U1249 ( .A(n994), .B(n995), .Z(n992) );
  NANDN U1250 ( .A(n996), .B(n994), .Z(n990) );
  XNOR U1251 ( .A(n971), .B(n997), .Z(N1172) );
  XOR U1252 ( .A(n973), .B(n974), .Z(n997) );
  XNOR U1253 ( .A(n987), .B(n998), .Z(n974) );
  XOR U1254 ( .A(n988), .B(n989), .Z(n998) );
  XOR U1255 ( .A(n994), .B(n999), .Z(n989) );
  XOR U1256 ( .A(n993), .B(n996), .Z(n999) );
  IV U1257 ( .A(n995), .Z(n996) );
  NAND U1258 ( .A(n1000), .B(n1001), .Z(n995) );
  OR U1259 ( .A(n1002), .B(n1003), .Z(n1001) );
  OR U1260 ( .A(n1004), .B(n1005), .Z(n1000) );
  NAND U1261 ( .A(n1006), .B(n1007), .Z(n993) );
  OR U1262 ( .A(n1008), .B(n1009), .Z(n1007) );
  OR U1263 ( .A(n1010), .B(n1011), .Z(n1006) );
  NOR U1264 ( .A(n1012), .B(n1013), .Z(n994) );
  ANDN U1265 ( .B(n1014), .A(n1015), .Z(n988) );
  XNOR U1266 ( .A(n981), .B(n1016), .Z(n987) );
  XNOR U1267 ( .A(n980), .B(n982), .Z(n1016) );
  NAND U1268 ( .A(n1017), .B(n1018), .Z(n982) );
  OR U1269 ( .A(n1019), .B(n1020), .Z(n1018) );
  OR U1270 ( .A(n1021), .B(n1022), .Z(n1017) );
  NAND U1271 ( .A(n1023), .B(n1024), .Z(n980) );
  OR U1272 ( .A(n1025), .B(n1026), .Z(n1024) );
  OR U1273 ( .A(n1027), .B(n1028), .Z(n1023) );
  ANDN U1274 ( .B(n1029), .A(n1030), .Z(n981) );
  IV U1275 ( .A(n1031), .Z(n1029) );
  ANDN U1276 ( .B(n1032), .A(n1033), .Z(n973) );
  XOR U1277 ( .A(n959), .B(n1034), .Z(n971) );
  XOR U1278 ( .A(n960), .B(n961), .Z(n1034) );
  XOR U1279 ( .A(n966), .B(n1035), .Z(n961) );
  XOR U1280 ( .A(n965), .B(n968), .Z(n1035) );
  IV U1281 ( .A(n967), .Z(n968) );
  NAND U1282 ( .A(n1036), .B(n1037), .Z(n967) );
  OR U1283 ( .A(n1038), .B(n1039), .Z(n1037) );
  OR U1284 ( .A(n1040), .B(n1041), .Z(n1036) );
  NAND U1285 ( .A(n1042), .B(n1043), .Z(n965) );
  OR U1286 ( .A(n1044), .B(n1045), .Z(n1043) );
  OR U1287 ( .A(n1046), .B(n1047), .Z(n1042) );
  NOR U1288 ( .A(n1048), .B(n1049), .Z(n966) );
  ANDN U1289 ( .B(n1050), .A(n1051), .Z(n960) );
  IV U1290 ( .A(n1052), .Z(n1050) );
  XNOR U1291 ( .A(n953), .B(n1053), .Z(n959) );
  XNOR U1292 ( .A(n952), .B(n954), .Z(n1053) );
  NAND U1293 ( .A(n1054), .B(n1055), .Z(n954) );
  OR U1294 ( .A(n1056), .B(n1057), .Z(n1055) );
  OR U1295 ( .A(n1058), .B(n1059), .Z(n1054) );
  NAND U1296 ( .A(n1060), .B(n1061), .Z(n952) );
  OR U1297 ( .A(n1062), .B(n1063), .Z(n1061) );
  OR U1298 ( .A(n1064), .B(n1065), .Z(n1060) );
  ANDN U1299 ( .B(n1066), .A(n1067), .Z(n953) );
  IV U1300 ( .A(n1068), .Z(n1066) );
  XNOR U1301 ( .A(n1033), .B(n1032), .Z(N1171) );
  XOR U1302 ( .A(n1052), .B(n1051), .Z(n1032) );
  XNOR U1303 ( .A(n1067), .B(n1068), .Z(n1051) );
  XNOR U1304 ( .A(n1062), .B(n1063), .Z(n1068) );
  XNOR U1305 ( .A(n1064), .B(n1065), .Z(n1063) );
  XNOR U1306 ( .A(y[112]), .B(x[112]), .Z(n1065) );
  XNOR U1307 ( .A(y[113]), .B(x[113]), .Z(n1064) );
  XNOR U1308 ( .A(y[111]), .B(x[111]), .Z(n1062) );
  XNOR U1309 ( .A(n1056), .B(n1057), .Z(n1067) );
  XNOR U1310 ( .A(y[108]), .B(x[108]), .Z(n1057) );
  XNOR U1311 ( .A(n1058), .B(n1059), .Z(n1056) );
  XNOR U1312 ( .A(y[109]), .B(x[109]), .Z(n1059) );
  XNOR U1313 ( .A(y[110]), .B(x[110]), .Z(n1058) );
  XNOR U1314 ( .A(n1049), .B(n1048), .Z(n1052) );
  XNOR U1315 ( .A(n1044), .B(n1045), .Z(n1048) );
  XNOR U1316 ( .A(y[105]), .B(x[105]), .Z(n1045) );
  XNOR U1317 ( .A(n1046), .B(n1047), .Z(n1044) );
  XNOR U1318 ( .A(y[106]), .B(x[106]), .Z(n1047) );
  XNOR U1319 ( .A(y[107]), .B(x[107]), .Z(n1046) );
  XNOR U1320 ( .A(n1038), .B(n1039), .Z(n1049) );
  XNOR U1321 ( .A(y[102]), .B(x[102]), .Z(n1039) );
  XNOR U1322 ( .A(n1040), .B(n1041), .Z(n1038) );
  XNOR U1323 ( .A(y[103]), .B(x[103]), .Z(n1041) );
  XNOR U1324 ( .A(y[104]), .B(x[104]), .Z(n1040) );
  XOR U1325 ( .A(n1014), .B(n1015), .Z(n1033) );
  XNOR U1326 ( .A(n1030), .B(n1031), .Z(n1015) );
  XNOR U1327 ( .A(n1025), .B(n1026), .Z(n1031) );
  XNOR U1328 ( .A(n1027), .B(n1028), .Z(n1026) );
  XNOR U1329 ( .A(y[100]), .B(x[100]), .Z(n1028) );
  XNOR U1330 ( .A(y[101]), .B(x[101]), .Z(n1027) );
  XNOR U1331 ( .A(y[99]), .B(x[99]), .Z(n1025) );
  XNOR U1332 ( .A(n1019), .B(n1020), .Z(n1030) );
  XNOR U1333 ( .A(y[96]), .B(x[96]), .Z(n1020) );
  XNOR U1334 ( .A(n1021), .B(n1022), .Z(n1019) );
  XNOR U1335 ( .A(y[97]), .B(x[97]), .Z(n1022) );
  XNOR U1336 ( .A(y[98]), .B(x[98]), .Z(n1021) );
  XOR U1337 ( .A(n1013), .B(n1012), .Z(n1014) );
  XNOR U1338 ( .A(n1008), .B(n1009), .Z(n1012) );
  XNOR U1339 ( .A(y[93]), .B(x[93]), .Z(n1009) );
  XNOR U1340 ( .A(n1010), .B(n1011), .Z(n1008) );
  XNOR U1341 ( .A(y[94]), .B(x[94]), .Z(n1011) );
  XNOR U1342 ( .A(y[95]), .B(x[95]), .Z(n1010) );
  XNOR U1343 ( .A(n1002), .B(n1003), .Z(n1013) );
  XNOR U1344 ( .A(y[90]), .B(x[90]), .Z(n1003) );
  XNOR U1345 ( .A(n1004), .B(n1005), .Z(n1002) );
  XNOR U1346 ( .A(y[91]), .B(x[91]), .Z(n1005) );
  XNOR U1347 ( .A(y[92]), .B(x[92]), .Z(n1004) );
  NAND U1348 ( .A(n1069), .B(n1070), .Z(N1167) );
  NANDN U1349 ( .A(n1071), .B(n1072), .Z(n1070) );
  OR U1350 ( .A(n1073), .B(n1074), .Z(n1072) );
  NAND U1351 ( .A(n1073), .B(n1074), .Z(n1069) );
  XOR U1352 ( .A(n1073), .B(n1075), .Z(N1166) );
  XNOR U1353 ( .A(n1071), .B(n1074), .Z(n1075) );
  AND U1354 ( .A(n1076), .B(n1077), .Z(n1074) );
  NANDN U1355 ( .A(n1078), .B(n1079), .Z(n1077) );
  NANDN U1356 ( .A(n1080), .B(n1081), .Z(n1079) );
  NANDN U1357 ( .A(n1081), .B(n1080), .Z(n1076) );
  NAND U1358 ( .A(n1082), .B(n1083), .Z(n1071) );
  NANDN U1359 ( .A(n1084), .B(n1085), .Z(n1083) );
  OR U1360 ( .A(n1086), .B(n1087), .Z(n1085) );
  NAND U1361 ( .A(n1087), .B(n1086), .Z(n1082) );
  AND U1362 ( .A(n1088), .B(n1089), .Z(n1073) );
  NANDN U1363 ( .A(n1090), .B(n1091), .Z(n1089) );
  NANDN U1364 ( .A(n1092), .B(n1093), .Z(n1091) );
  NANDN U1365 ( .A(n1093), .B(n1092), .Z(n1088) );
  XOR U1366 ( .A(n1087), .B(n1094), .Z(N1165) );
  XOR U1367 ( .A(n1084), .B(n1086), .Z(n1094) );
  XNOR U1368 ( .A(n1080), .B(n1095), .Z(n1086) );
  XNOR U1369 ( .A(n1078), .B(n1081), .Z(n1095) );
  NAND U1370 ( .A(n1096), .B(n1097), .Z(n1081) );
  NAND U1371 ( .A(n1098), .B(n1099), .Z(n1097) );
  OR U1372 ( .A(n1100), .B(n1101), .Z(n1098) );
  NANDN U1373 ( .A(n1102), .B(n1100), .Z(n1096) );
  IV U1374 ( .A(n1101), .Z(n1102) );
  NAND U1375 ( .A(n1103), .B(n1104), .Z(n1078) );
  NAND U1376 ( .A(n1105), .B(n1106), .Z(n1104) );
  NANDN U1377 ( .A(n1107), .B(n1108), .Z(n1105) );
  NANDN U1378 ( .A(n1108), .B(n1107), .Z(n1103) );
  AND U1379 ( .A(n1109), .B(n1110), .Z(n1080) );
  NAND U1380 ( .A(n1111), .B(n1112), .Z(n1110) );
  OR U1381 ( .A(n1113), .B(n1114), .Z(n1111) );
  NANDN U1382 ( .A(n1115), .B(n1113), .Z(n1109) );
  NAND U1383 ( .A(n1116), .B(n1117), .Z(n1084) );
  NANDN U1384 ( .A(n1118), .B(n1119), .Z(n1117) );
  OR U1385 ( .A(n1120), .B(n1121), .Z(n1119) );
  NANDN U1386 ( .A(n1122), .B(n1120), .Z(n1116) );
  IV U1387 ( .A(n1121), .Z(n1122) );
  XNOR U1388 ( .A(n1092), .B(n1123), .Z(n1087) );
  XNOR U1389 ( .A(n1090), .B(n1093), .Z(n1123) );
  NAND U1390 ( .A(n1124), .B(n1125), .Z(n1093) );
  NAND U1391 ( .A(n1126), .B(n1127), .Z(n1125) );
  OR U1392 ( .A(n1128), .B(n1129), .Z(n1126) );
  NANDN U1393 ( .A(n1130), .B(n1128), .Z(n1124) );
  IV U1394 ( .A(n1129), .Z(n1130) );
  NAND U1395 ( .A(n1131), .B(n1132), .Z(n1090) );
  NAND U1396 ( .A(n1133), .B(n1134), .Z(n1132) );
  NANDN U1397 ( .A(n1135), .B(n1136), .Z(n1133) );
  NANDN U1398 ( .A(n1136), .B(n1135), .Z(n1131) );
  AND U1399 ( .A(n1137), .B(n1138), .Z(n1092) );
  NAND U1400 ( .A(n1139), .B(n1140), .Z(n1138) );
  OR U1401 ( .A(n1141), .B(n1142), .Z(n1139) );
  NANDN U1402 ( .A(n1143), .B(n1141), .Z(n1137) );
  XNOR U1403 ( .A(n1118), .B(n1144), .Z(N1164) );
  XOR U1404 ( .A(n1120), .B(n1121), .Z(n1144) );
  XNOR U1405 ( .A(n1134), .B(n1145), .Z(n1121) );
  XOR U1406 ( .A(n1135), .B(n1136), .Z(n1145) );
  XOR U1407 ( .A(n1141), .B(n1146), .Z(n1136) );
  XOR U1408 ( .A(n1140), .B(n1143), .Z(n1146) );
  IV U1409 ( .A(n1142), .Z(n1143) );
  NAND U1410 ( .A(n1147), .B(n1148), .Z(n1142) );
  OR U1411 ( .A(n1149), .B(n1150), .Z(n1148) );
  OR U1412 ( .A(n1151), .B(n1152), .Z(n1147) );
  NAND U1413 ( .A(n1153), .B(n1154), .Z(n1140) );
  OR U1414 ( .A(n1155), .B(n1156), .Z(n1154) );
  OR U1415 ( .A(n1157), .B(n1158), .Z(n1153) );
  NOR U1416 ( .A(n1159), .B(n1160), .Z(n1141) );
  ANDN U1417 ( .B(n1161), .A(n1162), .Z(n1135) );
  XNOR U1418 ( .A(n1128), .B(n1163), .Z(n1134) );
  XNOR U1419 ( .A(n1127), .B(n1129), .Z(n1163) );
  NAND U1420 ( .A(n1164), .B(n1165), .Z(n1129) );
  OR U1421 ( .A(n1166), .B(n1167), .Z(n1165) );
  OR U1422 ( .A(n1168), .B(n1169), .Z(n1164) );
  NAND U1423 ( .A(n1170), .B(n1171), .Z(n1127) );
  OR U1424 ( .A(n1172), .B(n1173), .Z(n1171) );
  OR U1425 ( .A(n1174), .B(n1175), .Z(n1170) );
  ANDN U1426 ( .B(n1176), .A(n1177), .Z(n1128) );
  IV U1427 ( .A(n1178), .Z(n1176) );
  ANDN U1428 ( .B(n1179), .A(n1180), .Z(n1120) );
  XOR U1429 ( .A(n1106), .B(n1181), .Z(n1118) );
  XOR U1430 ( .A(n1107), .B(n1108), .Z(n1181) );
  XOR U1431 ( .A(n1113), .B(n1182), .Z(n1108) );
  XOR U1432 ( .A(n1112), .B(n1115), .Z(n1182) );
  IV U1433 ( .A(n1114), .Z(n1115) );
  NAND U1434 ( .A(n1183), .B(n1184), .Z(n1114) );
  OR U1435 ( .A(n1185), .B(n1186), .Z(n1184) );
  OR U1436 ( .A(n1187), .B(n1188), .Z(n1183) );
  NAND U1437 ( .A(n1189), .B(n1190), .Z(n1112) );
  OR U1438 ( .A(n1191), .B(n1192), .Z(n1190) );
  OR U1439 ( .A(n1193), .B(n1194), .Z(n1189) );
  NOR U1440 ( .A(n1195), .B(n1196), .Z(n1113) );
  ANDN U1441 ( .B(n1197), .A(n1198), .Z(n1107) );
  IV U1442 ( .A(n1199), .Z(n1197) );
  XNOR U1443 ( .A(n1100), .B(n1200), .Z(n1106) );
  XNOR U1444 ( .A(n1099), .B(n1101), .Z(n1200) );
  NAND U1445 ( .A(n1201), .B(n1202), .Z(n1101) );
  OR U1446 ( .A(n1203), .B(n1204), .Z(n1202) );
  OR U1447 ( .A(n1205), .B(n1206), .Z(n1201) );
  NAND U1448 ( .A(n1207), .B(n1208), .Z(n1099) );
  OR U1449 ( .A(n1209), .B(n1210), .Z(n1208) );
  OR U1450 ( .A(n1211), .B(n1212), .Z(n1207) );
  ANDN U1451 ( .B(n1213), .A(n1214), .Z(n1100) );
  IV U1452 ( .A(n1215), .Z(n1213) );
  XNOR U1453 ( .A(n1180), .B(n1179), .Z(N1163) );
  XOR U1454 ( .A(n1199), .B(n1198), .Z(n1179) );
  XNOR U1455 ( .A(n1214), .B(n1215), .Z(n1198) );
  XNOR U1456 ( .A(n1209), .B(n1210), .Z(n1215) );
  XNOR U1457 ( .A(n1211), .B(n1212), .Z(n1210) );
  XNOR U1458 ( .A(y[88]), .B(x[88]), .Z(n1212) );
  XNOR U1459 ( .A(y[89]), .B(x[89]), .Z(n1211) );
  XNOR U1460 ( .A(y[87]), .B(x[87]), .Z(n1209) );
  XNOR U1461 ( .A(n1203), .B(n1204), .Z(n1214) );
  XNOR U1462 ( .A(y[84]), .B(x[84]), .Z(n1204) );
  XNOR U1463 ( .A(n1205), .B(n1206), .Z(n1203) );
  XNOR U1464 ( .A(y[85]), .B(x[85]), .Z(n1206) );
  XNOR U1465 ( .A(y[86]), .B(x[86]), .Z(n1205) );
  XNOR U1466 ( .A(n1196), .B(n1195), .Z(n1199) );
  XNOR U1467 ( .A(n1191), .B(n1192), .Z(n1195) );
  XNOR U1468 ( .A(y[81]), .B(x[81]), .Z(n1192) );
  XNOR U1469 ( .A(n1193), .B(n1194), .Z(n1191) );
  XNOR U1470 ( .A(y[82]), .B(x[82]), .Z(n1194) );
  XNOR U1471 ( .A(y[83]), .B(x[83]), .Z(n1193) );
  XNOR U1472 ( .A(n1185), .B(n1186), .Z(n1196) );
  XNOR U1473 ( .A(y[78]), .B(x[78]), .Z(n1186) );
  XNOR U1474 ( .A(n1187), .B(n1188), .Z(n1185) );
  XNOR U1475 ( .A(y[79]), .B(x[79]), .Z(n1188) );
  XNOR U1476 ( .A(y[80]), .B(x[80]), .Z(n1187) );
  XOR U1477 ( .A(n1161), .B(n1162), .Z(n1180) );
  XNOR U1478 ( .A(n1177), .B(n1178), .Z(n1162) );
  XNOR U1479 ( .A(n1172), .B(n1173), .Z(n1178) );
  XNOR U1480 ( .A(n1174), .B(n1175), .Z(n1173) );
  XNOR U1481 ( .A(y[76]), .B(x[76]), .Z(n1175) );
  XNOR U1482 ( .A(y[77]), .B(x[77]), .Z(n1174) );
  XNOR U1483 ( .A(y[75]), .B(x[75]), .Z(n1172) );
  XNOR U1484 ( .A(n1166), .B(n1167), .Z(n1177) );
  XNOR U1485 ( .A(y[72]), .B(x[72]), .Z(n1167) );
  XNOR U1486 ( .A(n1168), .B(n1169), .Z(n1166) );
  XNOR U1487 ( .A(y[73]), .B(x[73]), .Z(n1169) );
  XNOR U1488 ( .A(y[74]), .B(x[74]), .Z(n1168) );
  XOR U1489 ( .A(n1160), .B(n1159), .Z(n1161) );
  XNOR U1490 ( .A(n1155), .B(n1156), .Z(n1159) );
  XNOR U1491 ( .A(y[69]), .B(x[69]), .Z(n1156) );
  XNOR U1492 ( .A(n1157), .B(n1158), .Z(n1155) );
  XNOR U1493 ( .A(y[70]), .B(x[70]), .Z(n1158) );
  XNOR U1494 ( .A(y[71]), .B(x[71]), .Z(n1157) );
  XNOR U1495 ( .A(n1149), .B(n1150), .Z(n1160) );
  XNOR U1496 ( .A(y[66]), .B(x[66]), .Z(n1150) );
  XNOR U1497 ( .A(n1151), .B(n1152), .Z(n1149) );
  XNOR U1498 ( .A(y[67]), .B(x[67]), .Z(n1152) );
  XNOR U1499 ( .A(y[68]), .B(x[68]), .Z(n1151) );
  NAND U1500 ( .A(n1216), .B(n1217), .Z(N1159) );
  NANDN U1501 ( .A(n1218), .B(n1219), .Z(n1217) );
  OR U1502 ( .A(n1220), .B(n1221), .Z(n1219) );
  NAND U1503 ( .A(n1220), .B(n1221), .Z(n1216) );
  XOR U1504 ( .A(n1220), .B(n1222), .Z(N1158) );
  XNOR U1505 ( .A(n1218), .B(n1221), .Z(n1222) );
  AND U1506 ( .A(n1223), .B(n1224), .Z(n1221) );
  NANDN U1507 ( .A(n1225), .B(n1226), .Z(n1224) );
  NANDN U1508 ( .A(n1227), .B(n1228), .Z(n1226) );
  NANDN U1509 ( .A(n1228), .B(n1227), .Z(n1223) );
  NAND U1510 ( .A(n1229), .B(n1230), .Z(n1218) );
  NANDN U1511 ( .A(n1231), .B(n1232), .Z(n1230) );
  OR U1512 ( .A(n1233), .B(n1234), .Z(n1232) );
  NAND U1513 ( .A(n1234), .B(n1233), .Z(n1229) );
  AND U1514 ( .A(n1235), .B(n1236), .Z(n1220) );
  NANDN U1515 ( .A(n1237), .B(n1238), .Z(n1236) );
  NANDN U1516 ( .A(n1239), .B(n1240), .Z(n1238) );
  NANDN U1517 ( .A(n1240), .B(n1239), .Z(n1235) );
  XOR U1518 ( .A(n1234), .B(n1241), .Z(N1157) );
  XOR U1519 ( .A(n1231), .B(n1233), .Z(n1241) );
  XNOR U1520 ( .A(n1227), .B(n1242), .Z(n1233) );
  XNOR U1521 ( .A(n1225), .B(n1228), .Z(n1242) );
  NAND U1522 ( .A(n1243), .B(n1244), .Z(n1228) );
  NAND U1523 ( .A(n1245), .B(n1246), .Z(n1244) );
  OR U1524 ( .A(n1247), .B(n1248), .Z(n1245) );
  NANDN U1525 ( .A(n1249), .B(n1247), .Z(n1243) );
  IV U1526 ( .A(n1248), .Z(n1249) );
  NAND U1527 ( .A(n1250), .B(n1251), .Z(n1225) );
  NAND U1528 ( .A(n1252), .B(n1253), .Z(n1251) );
  NANDN U1529 ( .A(n1254), .B(n1255), .Z(n1252) );
  NANDN U1530 ( .A(n1255), .B(n1254), .Z(n1250) );
  AND U1531 ( .A(n1256), .B(n1257), .Z(n1227) );
  NAND U1532 ( .A(n1258), .B(n1259), .Z(n1257) );
  OR U1533 ( .A(n1260), .B(n1261), .Z(n1258) );
  NANDN U1534 ( .A(n1262), .B(n1260), .Z(n1256) );
  NAND U1535 ( .A(n1263), .B(n1264), .Z(n1231) );
  NANDN U1536 ( .A(n1265), .B(n1266), .Z(n1264) );
  OR U1537 ( .A(n1267), .B(n1268), .Z(n1266) );
  NANDN U1538 ( .A(n1269), .B(n1267), .Z(n1263) );
  IV U1539 ( .A(n1268), .Z(n1269) );
  XNOR U1540 ( .A(n1239), .B(n1270), .Z(n1234) );
  XNOR U1541 ( .A(n1237), .B(n1240), .Z(n1270) );
  NAND U1542 ( .A(n1271), .B(n1272), .Z(n1240) );
  NAND U1543 ( .A(n1273), .B(n1274), .Z(n1272) );
  OR U1544 ( .A(n1275), .B(n1276), .Z(n1273) );
  NANDN U1545 ( .A(n1277), .B(n1275), .Z(n1271) );
  IV U1546 ( .A(n1276), .Z(n1277) );
  NAND U1547 ( .A(n1278), .B(n1279), .Z(n1237) );
  NAND U1548 ( .A(n1280), .B(n1281), .Z(n1279) );
  NANDN U1549 ( .A(n1282), .B(n1283), .Z(n1280) );
  NANDN U1550 ( .A(n1283), .B(n1282), .Z(n1278) );
  AND U1551 ( .A(n1284), .B(n1285), .Z(n1239) );
  NAND U1552 ( .A(n1286), .B(n1287), .Z(n1285) );
  OR U1553 ( .A(n1288), .B(n1289), .Z(n1286) );
  NANDN U1554 ( .A(n1290), .B(n1288), .Z(n1284) );
  XNOR U1555 ( .A(n1265), .B(n1291), .Z(N1156) );
  XOR U1556 ( .A(n1267), .B(n1268), .Z(n1291) );
  XNOR U1557 ( .A(n1281), .B(n1292), .Z(n1268) );
  XOR U1558 ( .A(n1282), .B(n1283), .Z(n1292) );
  XOR U1559 ( .A(n1288), .B(n1293), .Z(n1283) );
  XOR U1560 ( .A(n1287), .B(n1290), .Z(n1293) );
  IV U1561 ( .A(n1289), .Z(n1290) );
  NAND U1562 ( .A(n1294), .B(n1295), .Z(n1289) );
  OR U1563 ( .A(n1296), .B(n1297), .Z(n1295) );
  OR U1564 ( .A(n1298), .B(n1299), .Z(n1294) );
  NAND U1565 ( .A(n1300), .B(n1301), .Z(n1287) );
  OR U1566 ( .A(n1302), .B(n1303), .Z(n1301) );
  OR U1567 ( .A(n1304), .B(n1305), .Z(n1300) );
  NOR U1568 ( .A(n1306), .B(n1307), .Z(n1288) );
  ANDN U1569 ( .B(n1308), .A(n1309), .Z(n1282) );
  XNOR U1570 ( .A(n1275), .B(n1310), .Z(n1281) );
  XNOR U1571 ( .A(n1274), .B(n1276), .Z(n1310) );
  NAND U1572 ( .A(n1311), .B(n1312), .Z(n1276) );
  OR U1573 ( .A(n1313), .B(n1314), .Z(n1312) );
  OR U1574 ( .A(n1315), .B(n1316), .Z(n1311) );
  NAND U1575 ( .A(n1317), .B(n1318), .Z(n1274) );
  OR U1576 ( .A(n1319), .B(n1320), .Z(n1318) );
  OR U1577 ( .A(n1321), .B(n1322), .Z(n1317) );
  ANDN U1578 ( .B(n1323), .A(n1324), .Z(n1275) );
  IV U1579 ( .A(n1325), .Z(n1323) );
  ANDN U1580 ( .B(n1326), .A(n1327), .Z(n1267) );
  XOR U1581 ( .A(n1253), .B(n1328), .Z(n1265) );
  XOR U1582 ( .A(n1254), .B(n1255), .Z(n1328) );
  XOR U1583 ( .A(n1260), .B(n1329), .Z(n1255) );
  XOR U1584 ( .A(n1259), .B(n1262), .Z(n1329) );
  IV U1585 ( .A(n1261), .Z(n1262) );
  NAND U1586 ( .A(n1330), .B(n1331), .Z(n1261) );
  OR U1587 ( .A(n1332), .B(n1333), .Z(n1331) );
  OR U1588 ( .A(n1334), .B(n1335), .Z(n1330) );
  NAND U1589 ( .A(n1336), .B(n1337), .Z(n1259) );
  OR U1590 ( .A(n1338), .B(n1339), .Z(n1337) );
  OR U1591 ( .A(n1340), .B(n1341), .Z(n1336) );
  NOR U1592 ( .A(n1342), .B(n1343), .Z(n1260) );
  ANDN U1593 ( .B(n1344), .A(n1345), .Z(n1254) );
  IV U1594 ( .A(n1346), .Z(n1344) );
  XNOR U1595 ( .A(n1247), .B(n1347), .Z(n1253) );
  XNOR U1596 ( .A(n1246), .B(n1248), .Z(n1347) );
  NAND U1597 ( .A(n1348), .B(n1349), .Z(n1248) );
  OR U1598 ( .A(n1350), .B(n1351), .Z(n1349) );
  OR U1599 ( .A(n1352), .B(n1353), .Z(n1348) );
  NAND U1600 ( .A(n1354), .B(n1355), .Z(n1246) );
  OR U1601 ( .A(n1356), .B(n1357), .Z(n1355) );
  OR U1602 ( .A(n1358), .B(n1359), .Z(n1354) );
  ANDN U1603 ( .B(n1360), .A(n1361), .Z(n1247) );
  IV U1604 ( .A(n1362), .Z(n1360) );
  XNOR U1605 ( .A(n1327), .B(n1326), .Z(N1155) );
  XOR U1606 ( .A(n1346), .B(n1345), .Z(n1326) );
  XNOR U1607 ( .A(n1361), .B(n1362), .Z(n1345) );
  XNOR U1608 ( .A(n1356), .B(n1357), .Z(n1362) );
  XNOR U1609 ( .A(n1358), .B(n1359), .Z(n1357) );
  XNOR U1610 ( .A(y[64]), .B(x[64]), .Z(n1359) );
  XNOR U1611 ( .A(y[65]), .B(x[65]), .Z(n1358) );
  XNOR U1612 ( .A(y[63]), .B(x[63]), .Z(n1356) );
  XNOR U1613 ( .A(n1350), .B(n1351), .Z(n1361) );
  XNOR U1614 ( .A(y[60]), .B(x[60]), .Z(n1351) );
  XNOR U1615 ( .A(n1352), .B(n1353), .Z(n1350) );
  XNOR U1616 ( .A(y[61]), .B(x[61]), .Z(n1353) );
  XNOR U1617 ( .A(y[62]), .B(x[62]), .Z(n1352) );
  XNOR U1618 ( .A(n1343), .B(n1342), .Z(n1346) );
  XNOR U1619 ( .A(n1338), .B(n1339), .Z(n1342) );
  XNOR U1620 ( .A(y[57]), .B(x[57]), .Z(n1339) );
  XNOR U1621 ( .A(n1340), .B(n1341), .Z(n1338) );
  XNOR U1622 ( .A(y[58]), .B(x[58]), .Z(n1341) );
  XNOR U1623 ( .A(y[59]), .B(x[59]), .Z(n1340) );
  XNOR U1624 ( .A(n1332), .B(n1333), .Z(n1343) );
  XNOR U1625 ( .A(y[54]), .B(x[54]), .Z(n1333) );
  XNOR U1626 ( .A(n1334), .B(n1335), .Z(n1332) );
  XNOR U1627 ( .A(y[55]), .B(x[55]), .Z(n1335) );
  XNOR U1628 ( .A(y[56]), .B(x[56]), .Z(n1334) );
  XOR U1629 ( .A(n1308), .B(n1309), .Z(n1327) );
  XNOR U1630 ( .A(n1324), .B(n1325), .Z(n1309) );
  XNOR U1631 ( .A(n1319), .B(n1320), .Z(n1325) );
  XNOR U1632 ( .A(n1321), .B(n1322), .Z(n1320) );
  XNOR U1633 ( .A(y[52]), .B(x[52]), .Z(n1322) );
  XNOR U1634 ( .A(y[53]), .B(x[53]), .Z(n1321) );
  XNOR U1635 ( .A(y[51]), .B(x[51]), .Z(n1319) );
  XNOR U1636 ( .A(n1313), .B(n1314), .Z(n1324) );
  XNOR U1637 ( .A(y[48]), .B(x[48]), .Z(n1314) );
  XNOR U1638 ( .A(n1315), .B(n1316), .Z(n1313) );
  XNOR U1639 ( .A(y[49]), .B(x[49]), .Z(n1316) );
  XNOR U1640 ( .A(y[50]), .B(x[50]), .Z(n1315) );
  XOR U1641 ( .A(n1307), .B(n1306), .Z(n1308) );
  XNOR U1642 ( .A(n1302), .B(n1303), .Z(n1306) );
  XNOR U1643 ( .A(y[45]), .B(x[45]), .Z(n1303) );
  XNOR U1644 ( .A(n1304), .B(n1305), .Z(n1302) );
  XNOR U1645 ( .A(y[46]), .B(x[46]), .Z(n1305) );
  XNOR U1646 ( .A(y[47]), .B(x[47]), .Z(n1304) );
  XNOR U1647 ( .A(n1296), .B(n1297), .Z(n1307) );
  XNOR U1648 ( .A(y[42]), .B(x[42]), .Z(n1297) );
  XNOR U1649 ( .A(n1298), .B(n1299), .Z(n1296) );
  XNOR U1650 ( .A(y[43]), .B(x[43]), .Z(n1299) );
  XNOR U1651 ( .A(y[44]), .B(x[44]), .Z(n1298) );
  NAND U1652 ( .A(n1363), .B(n1364), .Z(N1151) );
  NANDN U1653 ( .A(n1365), .B(n1366), .Z(n1364) );
  OR U1654 ( .A(n1367), .B(n1368), .Z(n1366) );
  NAND U1655 ( .A(n1367), .B(n1368), .Z(n1363) );
  XOR U1656 ( .A(n1367), .B(n1369), .Z(N1150) );
  XNOR U1657 ( .A(n1365), .B(n1368), .Z(n1369) );
  AND U1658 ( .A(n1370), .B(n1371), .Z(n1368) );
  NANDN U1659 ( .A(n1372), .B(n1373), .Z(n1371) );
  NANDN U1660 ( .A(n1374), .B(n1375), .Z(n1373) );
  NANDN U1661 ( .A(n1375), .B(n1374), .Z(n1370) );
  NAND U1662 ( .A(n1376), .B(n1377), .Z(n1365) );
  NANDN U1663 ( .A(n1378), .B(n1379), .Z(n1377) );
  OR U1664 ( .A(n1380), .B(n1381), .Z(n1379) );
  NAND U1665 ( .A(n1381), .B(n1380), .Z(n1376) );
  AND U1666 ( .A(n1382), .B(n1383), .Z(n1367) );
  NANDN U1667 ( .A(n1384), .B(n1385), .Z(n1383) );
  NANDN U1668 ( .A(n1386), .B(n1387), .Z(n1385) );
  NANDN U1669 ( .A(n1387), .B(n1386), .Z(n1382) );
  XOR U1670 ( .A(n1381), .B(n1388), .Z(N1149) );
  XOR U1671 ( .A(n1378), .B(n1380), .Z(n1388) );
  XNOR U1672 ( .A(n1374), .B(n1389), .Z(n1380) );
  XNOR U1673 ( .A(n1372), .B(n1375), .Z(n1389) );
  NAND U1674 ( .A(n1390), .B(n1391), .Z(n1375) );
  NAND U1675 ( .A(n1392), .B(n1393), .Z(n1391) );
  OR U1676 ( .A(n1394), .B(n1395), .Z(n1392) );
  NANDN U1677 ( .A(n1396), .B(n1394), .Z(n1390) );
  IV U1678 ( .A(n1395), .Z(n1396) );
  NAND U1679 ( .A(n1397), .B(n1398), .Z(n1372) );
  NAND U1680 ( .A(n1399), .B(n1400), .Z(n1398) );
  NANDN U1681 ( .A(n1401), .B(n1402), .Z(n1399) );
  NANDN U1682 ( .A(n1402), .B(n1401), .Z(n1397) );
  AND U1683 ( .A(n1403), .B(n1404), .Z(n1374) );
  NAND U1684 ( .A(n1405), .B(n1406), .Z(n1404) );
  OR U1685 ( .A(n1407), .B(n1408), .Z(n1405) );
  NANDN U1686 ( .A(n1409), .B(n1407), .Z(n1403) );
  NAND U1687 ( .A(n1410), .B(n1411), .Z(n1378) );
  NANDN U1688 ( .A(n1412), .B(n1413), .Z(n1411) );
  OR U1689 ( .A(n1414), .B(n1415), .Z(n1413) );
  NANDN U1690 ( .A(n1416), .B(n1414), .Z(n1410) );
  IV U1691 ( .A(n1415), .Z(n1416) );
  XNOR U1692 ( .A(n1386), .B(n1417), .Z(n1381) );
  XNOR U1693 ( .A(n1384), .B(n1387), .Z(n1417) );
  NAND U1694 ( .A(n1418), .B(n1419), .Z(n1387) );
  NAND U1695 ( .A(n1420), .B(n1421), .Z(n1419) );
  OR U1696 ( .A(n1422), .B(n1423), .Z(n1420) );
  NANDN U1697 ( .A(n1424), .B(n1422), .Z(n1418) );
  IV U1698 ( .A(n1423), .Z(n1424) );
  NAND U1699 ( .A(n1425), .B(n1426), .Z(n1384) );
  NAND U1700 ( .A(n1427), .B(n1428), .Z(n1426) );
  NANDN U1701 ( .A(n1429), .B(n1430), .Z(n1427) );
  NANDN U1702 ( .A(n1430), .B(n1429), .Z(n1425) );
  AND U1703 ( .A(n1431), .B(n1432), .Z(n1386) );
  NAND U1704 ( .A(n1433), .B(n1434), .Z(n1432) );
  OR U1705 ( .A(n1435), .B(n1436), .Z(n1433) );
  NANDN U1706 ( .A(n1437), .B(n1435), .Z(n1431) );
  XNOR U1707 ( .A(n1412), .B(n1438), .Z(N1148) );
  XOR U1708 ( .A(n1414), .B(n1415), .Z(n1438) );
  XNOR U1709 ( .A(n1428), .B(n1439), .Z(n1415) );
  XOR U1710 ( .A(n1429), .B(n1430), .Z(n1439) );
  XOR U1711 ( .A(n1435), .B(n1440), .Z(n1430) );
  XOR U1712 ( .A(n1434), .B(n1437), .Z(n1440) );
  IV U1713 ( .A(n1436), .Z(n1437) );
  NAND U1714 ( .A(n1441), .B(n1442), .Z(n1436) );
  OR U1715 ( .A(n1443), .B(n1444), .Z(n1442) );
  OR U1716 ( .A(n1445), .B(n1446), .Z(n1441) );
  NAND U1717 ( .A(n1447), .B(n1448), .Z(n1434) );
  OR U1718 ( .A(n1449), .B(n1450), .Z(n1448) );
  OR U1719 ( .A(n1451), .B(n1452), .Z(n1447) );
  NOR U1720 ( .A(n1453), .B(n1454), .Z(n1435) );
  ANDN U1721 ( .B(n1455), .A(n1456), .Z(n1429) );
  XNOR U1722 ( .A(n1422), .B(n1457), .Z(n1428) );
  XNOR U1723 ( .A(n1421), .B(n1423), .Z(n1457) );
  NAND U1724 ( .A(n1458), .B(n1459), .Z(n1423) );
  OR U1725 ( .A(n1460), .B(n1461), .Z(n1459) );
  OR U1726 ( .A(n1462), .B(n1463), .Z(n1458) );
  NAND U1727 ( .A(n1464), .B(n1465), .Z(n1421) );
  OR U1728 ( .A(n1466), .B(n1467), .Z(n1465) );
  OR U1729 ( .A(n1468), .B(n1469), .Z(n1464) );
  ANDN U1730 ( .B(n1470), .A(n1471), .Z(n1422) );
  IV U1731 ( .A(n1472), .Z(n1470) );
  ANDN U1732 ( .B(n1473), .A(n1474), .Z(n1414) );
  XOR U1733 ( .A(n1400), .B(n1475), .Z(n1412) );
  XOR U1734 ( .A(n1401), .B(n1402), .Z(n1475) );
  XOR U1735 ( .A(n1407), .B(n1476), .Z(n1402) );
  XOR U1736 ( .A(n1406), .B(n1409), .Z(n1476) );
  IV U1737 ( .A(n1408), .Z(n1409) );
  NAND U1738 ( .A(n1477), .B(n1478), .Z(n1408) );
  OR U1739 ( .A(n1479), .B(n1480), .Z(n1478) );
  OR U1740 ( .A(n1481), .B(n1482), .Z(n1477) );
  NAND U1741 ( .A(n1483), .B(n1484), .Z(n1406) );
  OR U1742 ( .A(n1485), .B(n1486), .Z(n1484) );
  OR U1743 ( .A(n1487), .B(n1488), .Z(n1483) );
  NOR U1744 ( .A(n1489), .B(n1490), .Z(n1407) );
  ANDN U1745 ( .B(n1491), .A(n1492), .Z(n1401) );
  IV U1746 ( .A(n1493), .Z(n1491) );
  XNOR U1747 ( .A(n1394), .B(n1494), .Z(n1400) );
  XNOR U1748 ( .A(n1393), .B(n1395), .Z(n1494) );
  NAND U1749 ( .A(n1495), .B(n1496), .Z(n1395) );
  OR U1750 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1751 ( .A(n1499), .B(n1500), .Z(n1495) );
  NAND U1752 ( .A(n1501), .B(n1502), .Z(n1393) );
  OR U1753 ( .A(n1503), .B(n1504), .Z(n1502) );
  OR U1754 ( .A(n1505), .B(n1506), .Z(n1501) );
  ANDN U1755 ( .B(n1507), .A(n1508), .Z(n1394) );
  IV U1756 ( .A(n1509), .Z(n1507) );
  XNOR U1757 ( .A(n1474), .B(n1473), .Z(N1147) );
  XOR U1758 ( .A(n1493), .B(n1492), .Z(n1473) );
  XNOR U1759 ( .A(n1508), .B(n1509), .Z(n1492) );
  XNOR U1760 ( .A(n1503), .B(n1504), .Z(n1509) );
  XNOR U1761 ( .A(n1505), .B(n1506), .Z(n1504) );
  XNOR U1762 ( .A(y[40]), .B(x[40]), .Z(n1506) );
  XNOR U1763 ( .A(y[41]), .B(x[41]), .Z(n1505) );
  XNOR U1764 ( .A(y[39]), .B(x[39]), .Z(n1503) );
  XNOR U1765 ( .A(n1497), .B(n1498), .Z(n1508) );
  XNOR U1766 ( .A(y[36]), .B(x[36]), .Z(n1498) );
  XNOR U1767 ( .A(n1499), .B(n1500), .Z(n1497) );
  XNOR U1768 ( .A(y[37]), .B(x[37]), .Z(n1500) );
  XNOR U1769 ( .A(y[38]), .B(x[38]), .Z(n1499) );
  XNOR U1770 ( .A(n1490), .B(n1489), .Z(n1493) );
  XNOR U1771 ( .A(n1485), .B(n1486), .Z(n1489) );
  XNOR U1772 ( .A(y[33]), .B(x[33]), .Z(n1486) );
  XNOR U1773 ( .A(n1487), .B(n1488), .Z(n1485) );
  XNOR U1774 ( .A(y[34]), .B(x[34]), .Z(n1488) );
  XNOR U1775 ( .A(y[35]), .B(x[35]), .Z(n1487) );
  XNOR U1776 ( .A(n1479), .B(n1480), .Z(n1490) );
  XNOR U1777 ( .A(y[30]), .B(x[30]), .Z(n1480) );
  XNOR U1778 ( .A(n1481), .B(n1482), .Z(n1479) );
  XNOR U1779 ( .A(y[31]), .B(x[31]), .Z(n1482) );
  XNOR U1780 ( .A(y[32]), .B(x[32]), .Z(n1481) );
  XOR U1781 ( .A(n1455), .B(n1456), .Z(n1474) );
  XNOR U1782 ( .A(n1471), .B(n1472), .Z(n1456) );
  XNOR U1783 ( .A(n1466), .B(n1467), .Z(n1472) );
  XNOR U1784 ( .A(n1468), .B(n1469), .Z(n1467) );
  XNOR U1785 ( .A(y[28]), .B(x[28]), .Z(n1469) );
  XNOR U1786 ( .A(y[29]), .B(x[29]), .Z(n1468) );
  XNOR U1787 ( .A(y[27]), .B(x[27]), .Z(n1466) );
  XNOR U1788 ( .A(n1460), .B(n1461), .Z(n1471) );
  XNOR U1789 ( .A(y[24]), .B(x[24]), .Z(n1461) );
  XNOR U1790 ( .A(n1462), .B(n1463), .Z(n1460) );
  XNOR U1791 ( .A(y[25]), .B(x[25]), .Z(n1463) );
  XNOR U1792 ( .A(y[26]), .B(x[26]), .Z(n1462) );
  XOR U1793 ( .A(n1454), .B(n1453), .Z(n1455) );
  XNOR U1794 ( .A(n1449), .B(n1450), .Z(n1453) );
  XNOR U1795 ( .A(y[21]), .B(x[21]), .Z(n1450) );
  XNOR U1796 ( .A(n1451), .B(n1452), .Z(n1449) );
  XNOR U1797 ( .A(y[22]), .B(x[22]), .Z(n1452) );
  XNOR U1798 ( .A(y[23]), .B(x[23]), .Z(n1451) );
  XNOR U1799 ( .A(n1443), .B(n1444), .Z(n1454) );
  XNOR U1800 ( .A(y[18]), .B(x[18]), .Z(n1444) );
  XNOR U1801 ( .A(n1445), .B(n1446), .Z(n1443) );
  XNOR U1802 ( .A(y[19]), .B(x[19]), .Z(n1446) );
  XNOR U1803 ( .A(y[20]), .B(x[20]), .Z(n1445) );
  NANDN U1804 ( .A(n1510), .B(n1511), .Z(N1143) );
  NANDN U1805 ( .A(n1512), .B(n1513), .Z(n1511) );
  XNOR U1806 ( .A(n1512), .B(n1514), .Z(N1142) );
  ANDN U1807 ( .B(n1513), .A(n1510), .Z(n1514) );
  ANDN U1808 ( .B(n1515), .A(n1516), .Z(n1510) );
  NOR U1809 ( .A(n1517), .B(n1518), .Z(n1515) );
  NAND U1810 ( .A(n1519), .B(n1516), .Z(n1513) );
  NAND U1811 ( .A(n1520), .B(n1521), .Z(n1516) );
  NANDN U1812 ( .A(n1522), .B(n1523), .Z(n1521) );
  NANDN U1813 ( .A(n1524), .B(n1525), .Z(n1523) );
  NANDN U1814 ( .A(n1525), .B(n1524), .Z(n1520) );
  OR U1815 ( .A(n1518), .B(n1517), .Z(n1519) );
  IV U1816 ( .A(n1526), .Z(n1517) );
  NAND U1817 ( .A(n1527), .B(n1528), .Z(n1512) );
  NANDN U1818 ( .A(n1529), .B(n1530), .Z(n1528) );
  OR U1819 ( .A(n1531), .B(n1532), .Z(n1530) );
  NANDN U1820 ( .A(n1533), .B(n1531), .Z(n1527) );
  XOR U1821 ( .A(n1531), .B(n1534), .Z(N1141) );
  XNOR U1822 ( .A(n1529), .B(n1533), .Z(n1534) );
  IV U1823 ( .A(n1532), .Z(n1533) );
  XOR U1824 ( .A(n1518), .B(n1526), .Z(n1532) );
  NAND U1825 ( .A(n1535), .B(n1536), .Z(n1526) );
  OR U1826 ( .A(n1537), .B(n1538), .Z(n1536) );
  OR U1827 ( .A(n1539), .B(n1540), .Z(n1535) );
  AND U1828 ( .A(n1541), .B(n1542), .Z(n1518) );
  NAND U1829 ( .A(n1543), .B(n1544), .Z(n1542) );
  NAND U1830 ( .A(n1545), .B(n1546), .Z(n1543) );
  OR U1831 ( .A(n1545), .B(n1546), .Z(n1541) );
  NAND U1832 ( .A(n1547), .B(n1548), .Z(n1529) );
  NANDN U1833 ( .A(n1549), .B(n1550), .Z(n1548) );
  OR U1834 ( .A(n1551), .B(n1552), .Z(n1550) );
  NAND U1835 ( .A(n1552), .B(n1551), .Z(n1547) );
  XNOR U1836 ( .A(n1524), .B(n1553), .Z(n1531) );
  XNOR U1837 ( .A(n1522), .B(n1525), .Z(n1553) );
  NAND U1838 ( .A(n1554), .B(n1555), .Z(n1525) );
  NAND U1839 ( .A(n1556), .B(n1557), .Z(n1555) );
  OR U1840 ( .A(n1558), .B(n1559), .Z(n1556) );
  NANDN U1841 ( .A(n1560), .B(n1558), .Z(n1554) );
  IV U1842 ( .A(n1559), .Z(n1560) );
  NAND U1843 ( .A(n1561), .B(n1562), .Z(n1522) );
  NAND U1844 ( .A(n1563), .B(n1564), .Z(n1562) );
  NANDN U1845 ( .A(n1565), .B(n1566), .Z(n1563) );
  NANDN U1846 ( .A(n1566), .B(n1565), .Z(n1561) );
  AND U1847 ( .A(n1567), .B(n1568), .Z(n1524) );
  NAND U1848 ( .A(n1569), .B(n1570), .Z(n1568) );
  OR U1849 ( .A(n1571), .B(n1572), .Z(n1569) );
  NANDN U1850 ( .A(n1573), .B(n1571), .Z(n1567) );
  IV U1851 ( .A(n1572), .Z(n1573) );
  XNOR U1852 ( .A(n1549), .B(n1574), .Z(N1140) );
  XOR U1853 ( .A(n1551), .B(n1552), .Z(n1574) );
  XOR U1854 ( .A(n1544), .B(n1575), .Z(n1552) );
  XOR U1855 ( .A(n1546), .B(n1545), .Z(n1575) );
  OR U1856 ( .A(n1576), .B(n1577), .Z(n1545) );
  AND U1857 ( .A(n1578), .B(n1579), .Z(n1546) );
  OR U1858 ( .A(n1580), .B(n1581), .Z(n1579) );
  OR U1859 ( .A(n1582), .B(n1583), .Z(n1578) );
  XOR U1860 ( .A(n1537), .B(n1538), .Z(n1544) );
  XOR U1861 ( .A(n1584), .B(n1539), .Z(n1538) );
  AND U1862 ( .A(n1585), .B(n1586), .Z(n1539) );
  NANDN U1863 ( .A(n1587), .B(n1588), .Z(n1586) );
  OR U1864 ( .A(n1589), .B(n1590), .Z(n1585) );
  IV U1865 ( .A(n1540), .Z(n1584) );
  AND U1866 ( .A(n1591), .B(n1592), .Z(n1540) );
  NANDN U1867 ( .A(n1593), .B(n1594), .Z(n1592) );
  OR U1868 ( .A(n1595), .B(n1596), .Z(n1591) );
  AND U1869 ( .A(n1597), .B(n1598), .Z(n1537) );
  OR U1870 ( .A(n1599), .B(n1600), .Z(n1598) );
  NANDN U1871 ( .A(n1601), .B(n1602), .Z(n1597) );
  ANDN U1872 ( .B(n1603), .A(n1604), .Z(n1551) );
  XOR U1873 ( .A(n1564), .B(n1605), .Z(n1549) );
  XOR U1874 ( .A(n1565), .B(n1566), .Z(n1605) );
  XOR U1875 ( .A(n1571), .B(n1606), .Z(n1566) );
  XNOR U1876 ( .A(n1570), .B(n1572), .Z(n1606) );
  NAND U1877 ( .A(n1607), .B(n1608), .Z(n1572) );
  OR U1878 ( .A(n1609), .B(n1610), .Z(n1608) );
  IV U1879 ( .A(n1611), .Z(n1610) );
  OR U1880 ( .A(n1612), .B(n1613), .Z(n1607) );
  NAND U1881 ( .A(n1614), .B(n1615), .Z(n1570) );
  OR U1882 ( .A(n1616), .B(n1617), .Z(n1615) );
  OR U1883 ( .A(n1618), .B(n1619), .Z(n1614) );
  ANDN U1884 ( .B(n1620), .A(n1621), .Z(n1571) );
  IV U1885 ( .A(n1622), .Z(n1620) );
  NOR U1886 ( .A(n1623), .B(n1624), .Z(n1565) );
  XNOR U1887 ( .A(n1558), .B(n1625), .Z(n1564) );
  XNOR U1888 ( .A(n1557), .B(n1559), .Z(n1625) );
  NAND U1889 ( .A(n1626), .B(n1627), .Z(n1559) );
  OR U1890 ( .A(n1628), .B(n1629), .Z(n1627) );
  OR U1891 ( .A(n1630), .B(n1631), .Z(n1626) );
  NAND U1892 ( .A(n1632), .B(n1633), .Z(n1557) );
  OR U1893 ( .A(n1634), .B(n1635), .Z(n1633) );
  OR U1894 ( .A(n1636), .B(n1637), .Z(n1632) );
  ANDN U1895 ( .B(n1638), .A(n1639), .Z(n1558) );
  IV U1896 ( .A(n1640), .Z(n1638) );
  XNOR U1897 ( .A(n1604), .B(n1603), .Z(N1139) );
  XOR U1898 ( .A(n1623), .B(n1624), .Z(n1603) );
  XNOR U1899 ( .A(n1639), .B(n1640), .Z(n1624) );
  XNOR U1900 ( .A(n1634), .B(n1635), .Z(n1640) );
  XNOR U1901 ( .A(n1636), .B(n1637), .Z(n1635) );
  XNOR U1902 ( .A(y[16]), .B(x[16]), .Z(n1637) );
  XNOR U1903 ( .A(y[17]), .B(x[17]), .Z(n1636) );
  XNOR U1904 ( .A(y[15]), .B(x[15]), .Z(n1634) );
  XNOR U1905 ( .A(n1628), .B(n1629), .Z(n1639) );
  XNOR U1906 ( .A(y[12]), .B(x[12]), .Z(n1629) );
  XNOR U1907 ( .A(n1630), .B(n1631), .Z(n1628) );
  XNOR U1908 ( .A(y[13]), .B(x[13]), .Z(n1631) );
  XNOR U1909 ( .A(y[14]), .B(x[14]), .Z(n1630) );
  XNOR U1910 ( .A(n1622), .B(n1621), .Z(n1623) );
  XNOR U1911 ( .A(n1616), .B(n1617), .Z(n1621) );
  XNOR U1912 ( .A(y[9]), .B(x[9]), .Z(n1617) );
  XNOR U1913 ( .A(n1618), .B(n1619), .Z(n1616) );
  XNOR U1914 ( .A(y[10]), .B(x[10]), .Z(n1619) );
  XNOR U1915 ( .A(y[11]), .B(x[11]), .Z(n1618) );
  XOR U1916 ( .A(n1609), .B(n1611), .Z(n1622) );
  XOR U1917 ( .A(n1612), .B(n1613), .Z(n1611) );
  XNOR U1918 ( .A(y[7]), .B(x[7]), .Z(n1613) );
  XNOR U1919 ( .A(y[8]), .B(x[8]), .Z(n1612) );
  XNOR U1920 ( .A(y[6]), .B(x[6]), .Z(n1609) );
  XNOR U1921 ( .A(n1577), .B(n1576), .Z(n1604) );
  XOR U1922 ( .A(n1641), .B(n1599), .Z(n1576) );
  XNOR U1923 ( .A(y[249]), .B(x[249]), .Z(n1599) );
  IV U1924 ( .A(n1600), .Z(n1641) );
  XOR U1925 ( .A(n1602), .B(n1601), .Z(n1600) );
  XOR U1926 ( .A(n1587), .B(n1588), .Z(n1601) );
  XOR U1927 ( .A(n1590), .B(n1589), .Z(n1588) );
  XNOR U1928 ( .A(y[1]), .B(x[1]), .Z(n1589) );
  XNOR U1929 ( .A(y[2]), .B(x[2]), .Z(n1590) );
  XNOR U1930 ( .A(y[0]), .B(x[0]), .Z(n1587) );
  XNOR U1931 ( .A(n1593), .B(n1594), .Z(n1602) );
  XOR U1932 ( .A(n1596), .B(n1595), .Z(n1594) );
  XNOR U1933 ( .A(y[4]), .B(x[4]), .Z(n1595) );
  XNOR U1934 ( .A(y[5]), .B(x[5]), .Z(n1596) );
  XNOR U1935 ( .A(y[3]), .B(x[3]), .Z(n1593) );
  XNOR U1936 ( .A(n1580), .B(n1581), .Z(n1577) );
  XNOR U1937 ( .A(y[246]), .B(x[246]), .Z(n1581) );
  XNOR U1938 ( .A(n1582), .B(n1583), .Z(n1580) );
  XNOR U1939 ( .A(y[247]), .B(x[247]), .Z(n1583) );
  XNOR U1940 ( .A(y[248]), .B(x[248]), .Z(n1582) );
  NAND U1941 ( .A(n1642), .B(n1643), .Z(N1134) );
  NAND U1942 ( .A(n1644), .B(n1645), .Z(n1643) );
  OR U1943 ( .A(n1646), .B(n1647), .Z(n1644) );
  NANDN U1944 ( .A(n1648), .B(n1646), .Z(n1642) );
  XNOR U1945 ( .A(n1646), .B(n1649), .Z(N1133) );
  XOR U1946 ( .A(n1645), .B(n1648), .Z(n1649) );
  IV U1947 ( .A(n1647), .Z(n1648) );
  NAND U1948 ( .A(n1650), .B(n1651), .Z(n1647) );
  NAND U1949 ( .A(n1652), .B(n1653), .Z(n1651) );
  OR U1950 ( .A(n1654), .B(n1655), .Z(n1652) );
  NANDN U1951 ( .A(n1656), .B(n1654), .Z(n1650) );
  IV U1952 ( .A(n1655), .Z(n1656) );
  NAND U1953 ( .A(n1657), .B(n1658), .Z(n1645) );
  NAND U1954 ( .A(n1659), .B(n1660), .Z(n1658) );
  OR U1955 ( .A(n1661), .B(n1662), .Z(n1659) );
  NAND U1956 ( .A(n1662), .B(n1661), .Z(n1657) );
  NAND U1957 ( .A(n1663), .B(n1664), .Z(n1646) );
  NAND U1958 ( .A(n1665), .B(n1666), .Z(n1664) );
  OR U1959 ( .A(n1667), .B(n1668), .Z(n1665) );
  NANDN U1960 ( .A(n1669), .B(n1667), .Z(n1663) );
  XOR U1961 ( .A(n1660), .B(n1670), .Z(N1132) );
  XOR U1962 ( .A(n1661), .B(n1662), .Z(n1670) );
  XNOR U1963 ( .A(n1667), .B(n1671), .Z(n1662) );
  XOR U1964 ( .A(n1666), .B(n1669), .Z(n1671) );
  IV U1965 ( .A(n1668), .Z(n1669) );
  NAND U1966 ( .A(n1672), .B(n1673), .Z(n1668) );
  OR U1967 ( .A(n1674), .B(n1675), .Z(n1673) );
  OR U1968 ( .A(n1676), .B(n1677), .Z(n1672) );
  NAND U1969 ( .A(n1678), .B(n1679), .Z(n1666) );
  OR U1970 ( .A(n1680), .B(n1681), .Z(n1679) );
  OR U1971 ( .A(n1682), .B(n1683), .Z(n1678) );
  NOR U1972 ( .A(n1684), .B(n1685), .Z(n1667) );
  ANDN U1973 ( .B(n1686), .A(n1687), .Z(n1661) );
  XNOR U1974 ( .A(n1654), .B(n1688), .Z(n1660) );
  XNOR U1975 ( .A(n1653), .B(n1655), .Z(n1688) );
  NAND U1976 ( .A(n1689), .B(n1690), .Z(n1655) );
  OR U1977 ( .A(n1691), .B(n1692), .Z(n1690) );
  IV U1978 ( .A(n1693), .Z(n1692) );
  OR U1979 ( .A(n1694), .B(n1695), .Z(n1689) );
  NAND U1980 ( .A(n1696), .B(n1697), .Z(n1653) );
  OR U1981 ( .A(n1698), .B(n1699), .Z(n1697) );
  OR U1982 ( .A(n1700), .B(n1701), .Z(n1696) );
  AND U1983 ( .A(n1702), .B(n1703), .Z(n1654) );
  IV U1984 ( .A(n1704), .Z(n1703) );
  XNOR U1985 ( .A(n1687), .B(n1686), .Z(N1131) );
  XNOR U1986 ( .A(n1704), .B(n1702), .Z(n1686) );
  XOR U1987 ( .A(n1698), .B(n1699), .Z(n1702) );
  XNOR U1988 ( .A(n1700), .B(n1701), .Z(n1699) );
  XNOR U1989 ( .A(y[244]), .B(x[244]), .Z(n1701) );
  XNOR U1990 ( .A(y[245]), .B(x[245]), .Z(n1700) );
  XNOR U1991 ( .A(y[243]), .B(x[243]), .Z(n1698) );
  XOR U1992 ( .A(n1691), .B(n1693), .Z(n1704) );
  XOR U1993 ( .A(n1694), .B(n1695), .Z(n1693) );
  XNOR U1994 ( .A(y[241]), .B(x[241]), .Z(n1695) );
  XNOR U1995 ( .A(y[242]), .B(x[242]), .Z(n1694) );
  XNOR U1996 ( .A(y[240]), .B(x[240]), .Z(n1691) );
  XNOR U1997 ( .A(n1685), .B(n1684), .Z(n1687) );
  XNOR U1998 ( .A(n1680), .B(n1681), .Z(n1684) );
  XNOR U1999 ( .A(y[237]), .B(x[237]), .Z(n1681) );
  XNOR U2000 ( .A(n1682), .B(n1683), .Z(n1680) );
  XNOR U2001 ( .A(y[238]), .B(x[238]), .Z(n1683) );
  XNOR U2002 ( .A(y[239]), .B(x[239]), .Z(n1682) );
  XNOR U2003 ( .A(n1674), .B(n1675), .Z(n1685) );
  XNOR U2004 ( .A(y[234]), .B(x[234]), .Z(n1675) );
  XNOR U2005 ( .A(n1676), .B(n1677), .Z(n1674) );
  XNOR U2006 ( .A(y[235]), .B(x[235]), .Z(n1677) );
  XNOR U2007 ( .A(y[236]), .B(x[236]), .Z(n1676) );
endmodule

